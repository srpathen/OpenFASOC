* NGSPICE file created from opamp458.ext - technology: sky130A

.subckt opamp458 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 CSoutput.t167 a_n7636_8799.t36 vdd.t265 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 a_n2140_13878.t23 a_n2318_13878.t52 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2140_13878.t15 a_n2318_13878.t20 a_n2318_13878.t21 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t264 a_n7636_8799.t37 CSoutput.t166 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 outputibias.t1 outputibias.t0 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X5 a_n3827_n3924.t17 diffpairibias.t20 gnd.t351 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X6 gnd.t167 commonsourceibias.t80 CSoutput.t51 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t349 gnd.t347 gnd.t348 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 CSoutput.t165 a_n7636_8799.t38 vdd.t263 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 commonsourceibias.t79 commonsourceibias.t78 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X10 commonsourceibias.t77 commonsourceibias.t76 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t346 gnd.t344 gnd.t345 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X12 vdd.t125 vdd.t123 vdd.t124 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X13 vdd.t39 CSoutput.t176 output.t19 gnd.t224 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X14 a_n2318_8322.t23 a_n2318_13878.t53 a_n7636_8799.t32 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 gnd.t343 gnd.t341 gnd.t342 gnd.t259 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X16 CSoutput.t52 commonsourceibias.t81 gnd.t168 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t164 a_n7636_8799.t39 vdd.t262 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t75 commonsourceibias.t74 commonsourceibias.t75 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t340 gnd.t338 plus.t4 gnd.t339 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X20 CSoutput.t54 commonsourceibias.t82 gnd.t171 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 a_n7636_8799.t33 plus.t5 a_n3827_n3924.t43 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X22 vdd.t261 a_n7636_8799.t40 CSoutput.t163 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 gnd.t337 gnd.t335 gnd.t336 gnd.t259 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X24 minus.t4 gnd.t332 gnd.t334 gnd.t333 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 commonsourceibias.t73 commonsourceibias.t72 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 vdd.t40 CSoutput.t177 output.t18 gnd.t223 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X27 a_n7636_8799.t8 a_n2318_13878.t54 a_n2318_8322.t22 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X28 CSoutput.t55 commonsourceibias.t83 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 vdd.t260 a_n7636_8799.t41 CSoutput.t162 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 CSoutput.t161 a_n7636_8799.t42 vdd.t259 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 vdd.t258 a_n7636_8799.t43 CSoutput.t160 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 a_n7636_8799.t7 a_n2318_13878.t55 a_n2318_8322.t21 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 a_n7636_8799.t34 plus.t6 a_n3827_n3924.t44 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X34 gnd.t331 gnd.t328 gnd.t330 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X35 commonsourceibias.t71 commonsourceibias.t70 gnd.t76 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 vdd.t122 vdd.t120 vdd.t121 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X37 CSoutput.t159 a_n7636_8799.t44 vdd.t257 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n3827_n3924.t16 diffpairibias.t21 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X39 CSoutput.t45 commonsourceibias.t84 gnd.t159 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n3827_n3924.t42 minus.t5 a_n2318_13878.t47 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X41 CSoutput.t158 a_n7636_8799.t45 vdd.t256 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X42 gnd.t161 commonsourceibias.t85 CSoutput.t46 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n3827_n3924.t49 plus.t7 a_n7636_8799.t35 gnd.t126 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X44 gnd.t327 gnd.t325 gnd.t326 gnd.t247 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X45 gnd.t88 commonsourceibias.t68 commonsourceibias.t69 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 a_n2318_13878.t46 minus.t6 a_n3827_n3924.t41 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X47 a_n3827_n3924.t33 plus.t8 a_n7636_8799.t20 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X48 a_n3827_n3924.t29 minus.t7 a_n2318_13878.t41 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X49 CSoutput.t157 a_n7636_8799.t46 vdd.t255 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 commonsourceibias.t67 commonsourceibias.t66 gnd.t226 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 gnd.t201 commonsourceibias.t86 CSoutput.t68 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2140_13878.t14 a_n2318_13878.t12 a_n2318_13878.t13 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 vdd.t119 vdd.t117 vdd.t118 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X54 gnd.t202 commonsourceibias.t87 CSoutput.t69 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 a_n2318_13878.t7 a_n2318_13878.t6 a_n2140_13878.t13 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X56 gnd.t199 commonsourceibias.t88 CSoutput.t66 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 CSoutput.t156 a_n7636_8799.t47 vdd.t254 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 output.t17 CSoutput.t178 vdd.t41 gnd.t222 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X59 a_n3827_n3924.t1 minus.t8 a_n2318_13878.t0 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X60 vdd.t116 vdd.t114 vdd.t115 vdd.t97 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X61 vdd.t253 a_n7636_8799.t48 CSoutput.t155 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 gnd.t165 commonsourceibias.t64 commonsourceibias.t65 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 diffpairibias.t19 diffpairibias.t18 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X64 commonsourceibias.t63 commonsourceibias.t62 gnd.t227 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t324 gnd.t322 gnd.t323 gnd.t267 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X66 a_n7636_8799.t21 a_n2318_13878.t56 a_n2318_8322.t20 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t154 a_n7636_8799.t49 vdd.t252 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 commonsourceibias.t61 commonsourceibias.t60 gnd.t228 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 gnd.t321 gnd.t320 plus.t3 gnd.t267 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X70 vdd.t251 a_n7636_8799.t50 CSoutput.t153 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t250 a_n7636_8799.t51 CSoutput.t152 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 minus.t3 gnd.t317 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X73 gnd.t316 gnd.t313 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X74 diffpairibias.t17 diffpairibias.t16 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 gnd.t225 commonsourceibias.t58 commonsourceibias.t59 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 CSoutput.t151 a_n7636_8799.t52 vdd.t249 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 CSoutput.t67 commonsourceibias.t89 gnd.t200 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 vdd.t248 a_n7636_8799.t53 CSoutput.t150 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 CSoutput.t149 a_n7636_8799.t54 vdd.t247 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t64 commonsourceibias.t90 gnd.t197 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 CSoutput.t148 a_n7636_8799.t55 vdd.t246 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X82 CSoutput.t147 a_n7636_8799.t56 vdd.t245 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X83 CSoutput.t146 a_n7636_8799.t57 vdd.t244 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 gnd.t229 commonsourceibias.t56 commonsourceibias.t57 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 vdd.t42 CSoutput.t179 output.t16 gnd.t221 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X86 CSoutput.t65 commonsourceibias.t91 gnd.t198 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t171 commonsourceibias.t92 gnd.t239 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 a_n7636_8799.t2 plus.t9 a_n3827_n3924.t3 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X89 CSoutput.t172 commonsourceibias.t93 gnd.t240 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t174 commonsourceibias.t94 gnd.t357 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n3827_n3924.t15 diffpairibias.t22 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X92 vdd.t243 a_n7636_8799.t58 CSoutput.t145 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n3827_n3924.t28 minus.t9 a_n2318_13878.t40 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X94 a_n2318_13878.t15 a_n2318_13878.t14 a_n2140_13878.t12 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 vdd.t242 a_n7636_8799.t59 CSoutput.t144 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 output.t15 CSoutput.t180 vdd.t135 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X97 a_n7636_8799.t1 a_n2318_13878.t57 a_n2318_8322.t19 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t241 a_n7636_8799.t60 CSoutput.t143 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n2318_13878.t9 a_n2318_13878.t8 a_n2140_13878.t11 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 a_n2318_13878.t45 minus.t10 a_n3827_n3924.t38 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X101 gnd.t230 commonsourceibias.t54 commonsourceibias.t55 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 gnd.t231 commonsourceibias.t52 commonsourceibias.t53 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 a_n3827_n3924.t7 plus.t10 a_n7636_8799.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X104 gnd.t146 commonsourceibias.t50 commonsourceibias.t51 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 output.t3 outputibias.t8 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X106 CSoutput.t181 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X107 vdd.t240 a_n7636_8799.t61 CSoutput.t142 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 CSoutput.t141 a_n7636_8799.t62 vdd.t239 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 gnd.t312 gnd.t309 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X110 diffpairibias.t15 diffpairibias.t14 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X111 a_n3827_n3924.t37 minus.t11 a_n2318_13878.t44 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X112 output.t2 outputibias.t9 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X113 vdd.t113 vdd.t111 vdd.t112 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 vdd.t110 vdd.t108 vdd.t109 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X115 CSoutput.t140 a_n7636_8799.t63 vdd.t238 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t358 commonsourceibias.t95 CSoutput.t175 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t107 vdd.t104 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t176 commonsourceibias.t96 CSoutput.t57 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t177 commonsourceibias.t97 CSoutput.t58 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t163 commonsourceibias.t98 CSoutput.t48 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 gnd.t164 commonsourceibias.t99 CSoutput.t49 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 output.t14 CSoutput.t182 vdd.t136 gnd.t219 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X123 vdd.t43 CSoutput.t183 output.t13 gnd.t218 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X124 vdd.t6 a_n2318_13878.t58 a_n2318_8322.t7 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n2318_13878.t29 a_n2318_13878.t28 a_n2140_13878.t10 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd.t144 commonsourceibias.t100 CSoutput.t42 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t308 gnd.t306 gnd.t307 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X128 a_n2318_8322.t6 a_n2318_13878.t59 vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n3827_n3924.t14 diffpairibias.t23 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 CSoutput.t139 a_n7636_8799.t64 vdd.t237 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 CSoutput.t138 a_n7636_8799.t65 vdd.t235 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X132 a_n2318_13878.t51 minus.t12 a_n3827_n3924.t48 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X133 CSoutput.t43 commonsourceibias.t101 gnd.t145 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X134 gnd.t147 commonsourceibias.t48 commonsourceibias.t49 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 a_n3827_n3924.t20 plus.t11 a_n7636_8799.t11 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X136 vdd.t35 a_n2318_13878.t60 a_n2140_13878.t22 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 gnd.t54 commonsourceibias.t102 CSoutput.t16 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t103 vdd.t100 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X139 vdd.t234 a_n7636_8799.t66 CSoutput.t137 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 gnd.t149 commonsourceibias.t46 commonsourceibias.t47 gnd.t148 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 a_n7636_8799.t22 plus.t12 a_n3827_n3924.t34 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X142 vdd.t99 vdd.t96 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X143 a_n2318_8322.t5 a_n2318_13878.t61 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X144 a_n2318_13878.t43 minus.t13 a_n3827_n3924.t31 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X145 a_n7636_8799.t6 a_n2318_13878.t62 a_n2318_8322.t18 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 CSoutput.t136 a_n7636_8799.t67 vdd.t232 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 diffpairibias.t13 diffpairibias.t12 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X148 CSoutput.t184 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X149 vdd.t231 a_n7636_8799.t68 CSoutput.t135 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 CSoutput.t17 commonsourceibias.t103 gnd.t55 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 a_n2318_13878.t25 a_n2318_13878.t24 a_n2140_13878.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 vdd.t229 a_n7636_8799.t69 CSoutput.t134 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X153 a_n7636_8799.t29 a_n2318_13878.t63 a_n2318_8322.t17 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 CSoutput.t133 a_n7636_8799.t70 vdd.t228 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 CSoutput.t40 commonsourceibias.t104 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 a_n2140_13878.t8 a_n2318_13878.t10 a_n2318_13878.t11 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 commonsourceibias.t45 commonsourceibias.t44 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 CSoutput.t41 commonsourceibias.t105 gnd.t143 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 vdd.t95 vdd.t93 vdd.t94 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X160 gnd.t113 commonsourceibias.t106 CSoutput.t33 gnd.t3 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t34 commonsourceibias.t107 gnd.t114 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t44 CSoutput.t185 output.t12 gnd.t217 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X163 plus.t2 gnd.t303 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X164 CSoutput.t3 commonsourceibias.t108 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 gnd.t302 gnd.t300 minus.t2 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X166 gnd.t16 commonsourceibias.t109 CSoutput.t4 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput.t132 a_n7636_8799.t71 vdd.t227 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X168 gnd.t185 commonsourceibias.t42 commonsourceibias.t43 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2318_13878.t1 minus.t14 a_n3827_n3924.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X170 vdd.t38 a_n2318_13878.t64 a_n2318_8322.t4 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X171 a_n2140_13878.t7 a_n2318_13878.t18 a_n2318_13878.t19 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X172 gnd.t51 commonsourceibias.t110 CSoutput.t14 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd.t226 a_n7636_8799.t72 CSoutput.t131 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 a_n2318_13878.t35 a_n2318_13878.t34 a_n2140_13878.t6 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 commonsourceibias.t41 commonsourceibias.t40 gnd.t186 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 gnd.t152 commonsourceibias.t38 commonsourceibias.t39 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 vdd.t225 a_n7636_8799.t73 CSoutput.t130 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 gnd.t120 commonsourceibias.t36 commonsourceibias.t37 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 a_n3827_n3924.t13 diffpairibias.t24 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X180 commonsourceibias.t35 commonsourceibias.t34 gnd.t178 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 a_n3827_n3924.t12 diffpairibias.t25 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X182 gnd.t53 commonsourceibias.t111 CSoutput.t15 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n2318_13878.t3 minus.t15 a_n3827_n3924.t5 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X184 vdd.t224 a_n7636_8799.t74 CSoutput.t129 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 vdd.t223 a_n7636_8799.t75 CSoutput.t128 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X186 gnd.t110 commonsourceibias.t112 CSoutput.t31 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 gnd.t112 commonsourceibias.t113 CSoutput.t32 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 gnd.t28 commonsourceibias.t114 CSoutput.t6 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 gnd.t299 gnd.t297 minus.t1 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X190 gnd.t30 commonsourceibias.t115 CSoutput.t7 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X191 CSoutput.t186 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X192 CSoutput.t19 commonsourceibias.t116 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 gnd.t296 gnd.t294 gnd.t295 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X194 CSoutput.t127 a_n7636_8799.t76 vdd.t222 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 commonsourceibias.t33 commonsourceibias.t32 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t20 commonsourceibias.t117 gnd.t83 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X197 CSoutput.t126 a_n7636_8799.t77 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 a_n2318_13878.t39 minus.t16 a_n3827_n3924.t26 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X199 CSoutput.t125 a_n7636_8799.t78 vdd.t219 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 CSoutput.t187 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X201 gnd.t47 commonsourceibias.t118 CSoutput.t12 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 CSoutput.t13 commonsourceibias.t119 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 gnd.t293 gnd.t291 gnd.t292 gnd.t247 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 diffpairibias.t11 diffpairibias.t10 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 a_n2140_13878.t21 a_n2318_13878.t65 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 gnd.t10 commonsourceibias.t120 CSoutput.t1 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 vdd.t18 a_n2318_13878.t66 a_n2140_13878.t20 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X208 output.t1 outputibias.t10 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X209 vdd.t92 vdd.t90 vdd.t91 vdd.t80 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X210 gnd.t241 commonsourceibias.t30 commonsourceibias.t31 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 CSoutput.t124 a_n7636_8799.t79 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 gnd.t153 commonsourceibias.t28 commonsourceibias.t29 gnd.t3 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X213 a_n3827_n3924.t35 plus.t13 a_n7636_8799.t24 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X214 vdd.t216 a_n7636_8799.t80 CSoutput.t123 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 commonsourceibias.t27 commonsourceibias.t26 gnd.t205 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 vdd.t89 vdd.t87 vdd.t88 vdd.t80 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X217 CSoutput.t2 commonsourceibias.t121 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 a_n3827_n3924.t24 minus.t17 a_n2318_13878.t37 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X219 a_n2140_13878.t5 a_n2318_13878.t22 a_n2318_13878.t23 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X220 diffpairibias.t9 diffpairibias.t8 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X221 a_n3827_n3924.t40 plus.t14 a_n7636_8799.t27 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X222 a_n3827_n3924.t47 minus.t18 a_n2318_13878.t50 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X223 a_n7636_8799.t4 plus.t15 a_n3827_n3924.t6 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X224 vdd.t214 a_n7636_8799.t81 CSoutput.t122 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 gnd.t6 commonsourceibias.t24 commonsourceibias.t25 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 CSoutput.t22 commonsourceibias.t122 gnd.t92 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X227 a_n2318_8322.t16 a_n2318_13878.t67 a_n7636_8799.t19 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 CSoutput.t121 a_n7636_8799.t82 vdd.t213 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 diffpairibias.t7 diffpairibias.t6 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X230 vdd.t212 a_n7636_8799.t83 CSoutput.t120 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 gnd.t4 commonsourceibias.t123 CSoutput.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X232 vdd.t27 a_n2318_13878.t68 a_n2318_8322.t3 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X233 vdd.t210 a_n7636_8799.t84 CSoutput.t119 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X234 vdd.t207 a_n7636_8799.t85 CSoutput.t118 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 vdd.t137 CSoutput.t188 output.t11 gnd.t216 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X236 CSoutput.t170 commonsourceibias.t124 gnd.t238 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 CSoutput.t173 commonsourceibias.t125 gnd.t356 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t290 gnd.t287 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X239 gnd.t175 commonsourceibias.t126 CSoutput.t56 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 gnd.t286 gnd.t283 gnd.t285 gnd.t284 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X241 gnd.t140 commonsourceibias.t127 CSoutput.t39 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 a_n2140_13878.t19 a_n2318_13878.t69 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X243 CSoutput.t38 commonsourceibias.t128 gnd.t139 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 commonsourceibias.t23 commonsourceibias.t22 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 plus.t1 gnd.t280 gnd.t282 gnd.t281 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X246 CSoutput.t30 commonsourceibias.t129 gnd.t109 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 vdd.t209 a_n7636_8799.t86 CSoutput.t117 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t116 a_n7636_8799.t87 vdd.t208 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 CSoutput.t115 a_n7636_8799.t88 vdd.t205 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 gnd.t279 gnd.t277 minus.t0 gnd.t278 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X251 gnd.t276 gnd.t274 gnd.t275 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X252 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X253 a_n3827_n3924.t11 diffpairibias.t26 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X254 vdd.t82 vdd.t79 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X255 vdd.t127 a_n2318_13878.t70 a_n2318_8322.t2 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X256 a_n2318_8322.t15 a_n2318_13878.t71 a_n7636_8799.t23 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X257 CSoutput.t114 a_n7636_8799.t89 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 gnd.t128 commonsourceibias.t130 CSoutput.t35 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 vdd.t202 a_n7636_8799.t90 CSoutput.t113 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 CSoutput.t112 a_n7636_8799.t91 vdd.t201 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 vdd.t200 a_n7636_8799.t92 CSoutput.t111 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 vdd.t199 a_n7636_8799.t93 CSoutput.t110 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 gnd.t108 commonsourceibias.t131 CSoutput.t29 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 CSoutput.t37 commonsourceibias.t132 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 vdd.t78 vdd.t76 vdd.t77 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X266 a_n3827_n3924.t0 plus.t16 a_n7636_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X267 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X268 CSoutput.t28 commonsourceibias.t133 gnd.t106 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 vdd.t198 a_n7636_8799.t94 CSoutput.t109 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X270 a_n7636_8799.t26 plus.t17 a_n3827_n3924.t39 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X271 CSoutput.t108 a_n7636_8799.t95 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X272 gnd.t136 commonsourceibias.t134 CSoutput.t36 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 a_n3827_n3924.t30 minus.t19 a_n2318_13878.t42 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X274 gnd.t105 commonsourceibias.t135 CSoutput.t27 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2140_13878.t4 a_n2318_13878.t4 a_n2318_13878.t5 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 CSoutput.t107 a_n7636_8799.t96 vdd.t192 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 vdd.t128 CSoutput.t189 output.t10 gnd.t215 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X278 CSoutput.t18 commonsourceibias.t136 gnd.t72 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 a_n2318_8322.t14 a_n2318_13878.t72 a_n7636_8799.t30 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 diffpairibias.t5 diffpairibias.t4 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 a_n3827_n3924.t25 minus.t20 a_n2318_13878.t38 gnd.t126 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X282 a_n7636_8799.t13 plus.t18 a_n3827_n3924.t21 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X283 commonsourceibias.t21 commonsourceibias.t20 gnd.t187 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 gnd.t273 gnd.t270 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X285 gnd.t45 commonsourceibias.t137 CSoutput.t11 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t26 commonsourceibias.t138 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t20 commonsourceibias.t18 commonsourceibias.t19 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 CSoutput.t106 a_n7636_8799.t97 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t105 a_n7636_8799.t98 vdd.t191 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 a_n3827_n3924.t10 diffpairibias.t27 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X291 vdd.t193 a_n7636_8799.t99 CSoutput.t104 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t21 commonsourceibias.t139 gnd.t91 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 CSoutput.t190 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X294 vdd.t190 a_n7636_8799.t100 CSoutput.t103 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 a_n2318_8322.t1 a_n2318_13878.t73 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X296 CSoutput.t102 a_n7636_8799.t101 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 CSoutput.t10 commonsourceibias.t140 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X298 a_n3827_n3924.t27 plus.t19 a_n7636_8799.t15 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X299 vdd.t71 vdd.t69 vdd.t70 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X300 vdd.t49 a_n2318_13878.t74 a_n2140_13878.t18 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X301 gnd.t188 commonsourceibias.t16 commonsourceibias.t17 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 output.t0 outputibias.t11 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X303 CSoutput.t101 a_n7636_8799.t102 vdd.t183 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t25 commonsourceibias.t141 gnd.t100 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 CSoutput.t100 a_n7636_8799.t103 vdd.t186 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 gnd.t184 commonsourceibias.t142 CSoutput.t62 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t269 gnd.t266 gnd.t268 gnd.t267 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X308 vdd.t185 a_n7636_8799.t104 CSoutput.t99 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 vdd.t181 a_n7636_8799.t105 CSoutput.t98 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 CSoutput.t24 commonsourceibias.t143 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 a_n3827_n3924.t23 minus.t21 a_n2318_13878.t36 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X312 vdd.t68 vdd.t66 vdd.t67 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X313 commonsourceibias.t15 commonsourceibias.t14 gnd.t208 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X314 commonsourceibias.t13 commonsourceibias.t12 gnd.t121 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n2318_8322.t13 a_n2318_13878.t75 a_n7636_8799.t31 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 CSoutput.t97 a_n7636_8799.t106 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X317 CSoutput.t61 commonsourceibias.t144 gnd.t182 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 a_n7636_8799.t28 a_n2318_13878.t76 a_n2318_8322.t12 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X319 gnd.t179 commonsourceibias.t10 commonsourceibias.t11 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 output.t9 CSoutput.t191 vdd.t129 gnd.t214 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X321 vdd.t178 a_n7636_8799.t107 CSoutput.t96 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X322 a_n2140_13878.t17 a_n2318_13878.t77 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X323 gnd.t170 commonsourceibias.t145 CSoutput.t53 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 CSoutput.t50 commonsourceibias.t146 gnd.t166 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t176 a_n7636_8799.t108 CSoutput.t95 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 CSoutput.t94 a_n7636_8799.t109 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 gnd.t265 gnd.t262 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X328 a_n7636_8799.t25 plus.t20 a_n3827_n3924.t36 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X329 commonsourceibias.t9 commonsourceibias.t8 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n2318_8322.t11 a_n2318_13878.t78 a_n7636_8799.t18 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X331 a_n2318_13878.t49 minus.t22 a_n3827_n3924.t46 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X332 vdd.t173 a_n7636_8799.t110 CSoutput.t93 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t92 a_n7636_8799.t111 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 CSoutput.t91 a_n7636_8799.t112 vdd.t169 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t242 commonsourceibias.t6 commonsourceibias.t7 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 CSoutput.t90 a_n7636_8799.t113 vdd.t168 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 a_n2140_13878.t3 a_n2318_13878.t32 a_n2318_13878.t33 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X338 commonsourceibias.t5 commonsourceibias.t4 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 vdd.t167 a_n7636_8799.t114 CSoutput.t89 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 gnd.t162 commonsourceibias.t147 CSoutput.t47 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 CSoutput.t44 commonsourceibias.t148 gnd.t158 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 vdd.t65 vdd.t62 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X343 CSoutput.t192 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X344 vdd.t61 vdd.t58 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 output.t8 CSoutput.t193 vdd.t130 gnd.t213 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X346 gnd.t18 commonsourceibias.t149 CSoutput.t5 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n7636_8799.t9 plus.t21 a_n3827_n3924.t18 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X348 a_n3827_n3924.t9 diffpairibias.t28 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X349 vdd.t166 a_n7636_8799.t115 CSoutput.t88 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X350 vdd.t165 a_n7636_8799.t116 CSoutput.t87 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 gnd.t41 commonsourceibias.t150 CSoutput.t9 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 CSoutput.t86 a_n7636_8799.t117 vdd.t164 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 a_n2318_13878.t27 a_n2318_13878.t26 a_n2140_13878.t2 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X354 gnd.t261 gnd.t258 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X355 a_n7636_8799.t16 a_n2318_13878.t79 a_n2318_8322.t10 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X356 vdd.t163 a_n7636_8799.t118 CSoutput.t85 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 output.t7 CSoutput.t194 vdd.t131 gnd.t212 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X358 gnd.t232 commonsourceibias.t151 CSoutput.t168 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 CSoutput.t84 a_n7636_8799.t119 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 a_n3827_n3924.t22 plus.t22 a_n7636_8799.t14 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X361 vdd.t132 CSoutput.t195 output.t6 gnd.t211 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X362 vdd.t160 a_n7636_8799.t120 CSoutput.t83 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 gnd.t257 gnd.t254 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X364 CSoutput.t169 commonsourceibias.t152 gnd.t233 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 CSoutput.t71 commonsourceibias.t153 gnd.t207 gnd.t101 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 commonsourceibias.t3 commonsourceibias.t2 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 outputibias.t7 outputibias.t6 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X368 diffpairibias.t3 diffpairibias.t2 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X369 vdd.t159 a_n7636_8799.t121 CSoutput.t82 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 CSoutput.t81 a_n7636_8799.t122 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n2318_8322.t9 a_n2318_13878.t80 a_n7636_8799.t3 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X372 vdd.t155 a_n7636_8799.t123 CSoutput.t80 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 outputibias.t5 outputibias.t4 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X374 diffpairibias.t1 diffpairibias.t0 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X375 a_n7636_8799.t17 plus.t23 a_n3827_n3924.t32 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X376 CSoutput.t8 commonsourceibias.t154 gnd.t39 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 outputibias.t3 outputibias.t2 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X378 gnd.t253 gnd.t250 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X379 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X380 vdd.t30 a_n2318_13878.t81 a_n2140_13878.t16 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X381 gnd.t206 commonsourceibias.t155 CSoutput.t70 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 CSoutput.t79 a_n7636_8799.t124 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X384 vdd.t151 a_n7636_8799.t125 CSoutput.t78 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 vdd.t149 a_n7636_8799.t126 CSoutput.t77 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 CSoutput.t23 commonsourceibias.t156 gnd.t97 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 CSoutput.t76 a_n7636_8799.t127 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 output.t5 CSoutput.t196 vdd.t133 gnd.t210 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X389 gnd.t181 commonsourceibias.t157 CSoutput.t60 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 gnd.t249 gnd.t246 gnd.t248 gnd.t247 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X391 a_n2318_13878.t48 minus.t23 a_n3827_n3924.t45 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X392 gnd.t180 commonsourceibias.t158 CSoutput.t59 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 a_n2318_8322.t8 a_n2318_13878.t82 a_n7636_8799.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X394 vdd.t145 a_n7636_8799.t128 CSoutput.t75 vdd.t144 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X395 vdd.t143 a_n7636_8799.t129 CSoutput.t74 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 CSoutput.t73 a_n7636_8799.t130 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 output.t4 CSoutput.t197 vdd.t134 gnd.t209 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X398 gnd.t196 commonsourceibias.t159 CSoutput.t63 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 gnd.t245 gnd.t243 plus.t0 gnd.t244 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X400 a_n3827_n3924.t19 plus.t24 a_n7636_8799.t10 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X401 a_n2318_8322.t0 a_n2318_13878.t83 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X402 a_n2318_13878.t2 minus.t24 a_n3827_n3924.t4 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X403 a_n2140_13878.t1 a_n2318_13878.t16 a_n2318_13878.t17 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X404 vdd.t139 a_n7636_8799.t131 CSoutput.t72 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 commonsourceibias.t1 commonsourceibias.t0 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 a_n3827_n3924.t8 diffpairibias.t29 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X407 a_n2318_13878.t31 a_n2318_13878.t30 a_n2140_13878.t0 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n7636_8799.n179 a_n7636_8799.t56 485.149
R1 a_n7636_8799.n195 a_n7636_8799.t65 485.149
R2 a_n7636_8799.n212 a_n7636_8799.t95 485.149
R3 a_n7636_8799.n128 a_n7636_8799.t115 485.149
R4 a_n7636_8799.n144 a_n7636_8799.t128 485.149
R5 a_n7636_8799.n161 a_n7636_8799.t94 485.149
R6 a_n7636_8799.n189 a_n7636_8799.t75 464.166
R7 a_n7636_8799.n188 a_n7636_8799.t57 464.166
R8 a_n7636_8799.n174 a_n7636_8799.t120 464.166
R9 a_n7636_8799.n187 a_n7636_8799.t88 464.166
R10 a_n7636_8799.n186 a_n7636_8799.t86 464.166
R11 a_n7636_8799.n175 a_n7636_8799.t38 464.166
R12 a_n7636_8799.n185 a_n7636_8799.t92 464.166
R13 a_n7636_8799.n184 a_n7636_8799.t91 464.166
R14 a_n7636_8799.n176 a_n7636_8799.t40 464.166
R15 a_n7636_8799.n183 a_n7636_8799.t39 464.166
R16 a_n7636_8799.n182 a_n7636_8799.t108 464.166
R17 a_n7636_8799.n177 a_n7636_8799.t52 464.166
R18 a_n7636_8799.n181 a_n7636_8799.t43 464.166
R19 a_n7636_8799.n180 a_n7636_8799.t112 464.166
R20 a_n7636_8799.n178 a_n7636_8799.t74 464.166
R21 a_n7636_8799.n205 a_n7636_8799.t84 464.166
R22 a_n7636_8799.n204 a_n7636_8799.t64 464.166
R23 a_n7636_8799.n190 a_n7636_8799.t131 464.166
R24 a_n7636_8799.n203 a_n7636_8799.t101 464.166
R25 a_n7636_8799.n202 a_n7636_8799.t100 464.166
R26 a_n7636_8799.n191 a_n7636_8799.t46 464.166
R27 a_n7636_8799.n201 a_n7636_8799.t104 464.166
R28 a_n7636_8799.n200 a_n7636_8799.t103 464.166
R29 a_n7636_8799.n192 a_n7636_8799.t48 464.166
R30 a_n7636_8799.n199 a_n7636_8799.t47 464.166
R31 a_n7636_8799.n198 a_n7636_8799.t123 464.166
R32 a_n7636_8799.n193 a_n7636_8799.t63 464.166
R33 a_n7636_8799.n197 a_n7636_8799.t51 464.166
R34 a_n7636_8799.n196 a_n7636_8799.t124 464.166
R35 a_n7636_8799.n194 a_n7636_8799.t85 464.166
R36 a_n7636_8799.n222 a_n7636_8799.t107 464.166
R37 a_n7636_8799.n221 a_n7636_8799.t54 464.166
R38 a_n7636_8799.n207 a_n7636_8799.t90 464.166
R39 a_n7636_8799.n220 a_n7636_8799.t42 464.166
R40 a_n7636_8799.n219 a_n7636_8799.t59 464.166
R41 a_n7636_8799.n208 a_n7636_8799.t127 464.166
R42 a_n7636_8799.n218 a_n7636_8799.t99 464.166
R43 a_n7636_8799.n217 a_n7636_8799.t122 464.166
R44 a_n7636_8799.n209 a_n7636_8799.t83 464.166
R45 a_n7636_8799.n216 a_n7636_8799.t102 464.166
R46 a_n7636_8799.n215 a_n7636_8799.t50 464.166
R47 a_n7636_8799.n210 a_n7636_8799.t119 464.166
R48 a_n7636_8799.n214 a_n7636_8799.t68 464.166
R49 a_n7636_8799.n213 a_n7636_8799.t113 464.166
R50 a_n7636_8799.n211 a_n7636_8799.t58 464.166
R51 a_n7636_8799.n127 a_n7636_8799.t117 464.166
R52 a_n7636_8799.n130 a_n7636_8799.t73 464.166
R53 a_n7636_8799.n126 a_n7636_8799.t98 464.166
R54 a_n7636_8799.n131 a_n7636_8799.t114 464.166
R55 a_n7636_8799.n132 a_n7636_8799.t71 464.166
R56 a_n7636_8799.n133 a_n7636_8799.t72 464.166
R57 a_n7636_8799.n134 a_n7636_8799.t96 464.166
R58 a_n7636_8799.n125 a_n7636_8799.t61 464.166
R59 a_n7636_8799.n135 a_n7636_8799.t62 464.166
R60 a_n7636_8799.n136 a_n7636_8799.t93 464.166
R61 a_n7636_8799.n137 a_n7636_8799.t36 464.166
R62 a_n7636_8799.n138 a_n7636_8799.t60 464.166
R63 a_n7636_8799.n124 a_n7636_8799.t78 464.166
R64 a_n7636_8799.n139 a_n7636_8799.t116 464.166
R65 a_n7636_8799.n143 a_n7636_8799.t130 464.166
R66 a_n7636_8799.n146 a_n7636_8799.t81 464.166
R67 a_n7636_8799.n142 a_n7636_8799.t111 464.166
R68 a_n7636_8799.n147 a_n7636_8799.t126 464.166
R69 a_n7636_8799.n148 a_n7636_8799.t79 464.166
R70 a_n7636_8799.n149 a_n7636_8799.t80 464.166
R71 a_n7636_8799.n150 a_n7636_8799.t109 464.166
R72 a_n7636_8799.n141 a_n7636_8799.t69 464.166
R73 a_n7636_8799.n151 a_n7636_8799.t70 464.166
R74 a_n7636_8799.n152 a_n7636_8799.t105 464.166
R75 a_n7636_8799.n153 a_n7636_8799.t44 464.166
R76 a_n7636_8799.n154 a_n7636_8799.t66 464.166
R77 a_n7636_8799.n140 a_n7636_8799.t87 464.166
R78 a_n7636_8799.n155 a_n7636_8799.t129 464.166
R79 a_n7636_8799.n160 a_n7636_8799.t76 464.166
R80 a_n7636_8799.n163 a_n7636_8799.t110 464.166
R81 a_n7636_8799.n159 a_n7636_8799.t67 464.166
R82 a_n7636_8799.n164 a_n7636_8799.t118 464.166
R83 a_n7636_8799.n165 a_n7636_8799.t49 464.166
R84 a_n7636_8799.n166 a_n7636_8799.t37 464.166
R85 a_n7636_8799.n167 a_n7636_8799.t82 464.166
R86 a_n7636_8799.n158 a_n7636_8799.t121 464.166
R87 a_n7636_8799.n168 a_n7636_8799.t97 464.166
R88 a_n7636_8799.n169 a_n7636_8799.t125 464.166
R89 a_n7636_8799.n170 a_n7636_8799.t77 464.166
R90 a_n7636_8799.n171 a_n7636_8799.t41 464.166
R91 a_n7636_8799.n157 a_n7636_8799.t89 464.166
R92 a_n7636_8799.n172 a_n7636_8799.t53 464.166
R93 a_n7636_8799.n52 a_n7636_8799.n30 74.4178
R94 a_n7636_8799.n180 a_n7636_8799.n52 12.4674
R95 a_n7636_8799.n51 a_n7636_8799.n30 80.107
R96 a_n7636_8799.n51 a_n7636_8799.n181 1.08907
R97 a_n7636_8799.n31 a_n7636_8799.n50 75.3623
R98 a_n7636_8799.n49 a_n7636_8799.n31 70.3058
R99 a_n7636_8799.n33 a_n7636_8799.n48 70.1674
R100 a_n7636_8799.n48 a_n7636_8799.n176 20.9683
R101 a_n7636_8799.n47 a_n7636_8799.n33 75.0448
R102 a_n7636_8799.n184 a_n7636_8799.n47 11.2134
R103 a_n7636_8799.n46 a_n7636_8799.n32 80.4688
R104 a_n7636_8799.n32 a_n7636_8799.n45 74.73
R105 a_n7636_8799.n44 a_n7636_8799.n34 70.1674
R106 a_n7636_8799.n187 a_n7636_8799.n44 20.9683
R107 a_n7636_8799.n34 a_n7636_8799.n43 70.5844
R108 a_n7636_8799.n43 a_n7636_8799.n174 20.1342
R109 a_n7636_8799.n42 a_n7636_8799.n35 75.6825
R110 a_n7636_8799.n188 a_n7636_8799.n42 9.93802
R111 a_n7636_8799.n35 a_n7636_8799.n189 161.3
R112 a_n7636_8799.n63 a_n7636_8799.n24 74.4178
R113 a_n7636_8799.n196 a_n7636_8799.n63 12.4674
R114 a_n7636_8799.n62 a_n7636_8799.n24 80.107
R115 a_n7636_8799.n62 a_n7636_8799.n197 1.08907
R116 a_n7636_8799.n25 a_n7636_8799.n61 75.3623
R117 a_n7636_8799.n60 a_n7636_8799.n25 70.3058
R118 a_n7636_8799.n27 a_n7636_8799.n59 70.1674
R119 a_n7636_8799.n59 a_n7636_8799.n192 20.9683
R120 a_n7636_8799.n58 a_n7636_8799.n27 75.0448
R121 a_n7636_8799.n200 a_n7636_8799.n58 11.2134
R122 a_n7636_8799.n57 a_n7636_8799.n26 80.4688
R123 a_n7636_8799.n26 a_n7636_8799.n56 74.73
R124 a_n7636_8799.n55 a_n7636_8799.n28 70.1674
R125 a_n7636_8799.n203 a_n7636_8799.n55 20.9683
R126 a_n7636_8799.n28 a_n7636_8799.n54 70.5844
R127 a_n7636_8799.n54 a_n7636_8799.n190 20.1342
R128 a_n7636_8799.n53 a_n7636_8799.n29 75.6825
R129 a_n7636_8799.n204 a_n7636_8799.n53 9.93802
R130 a_n7636_8799.n29 a_n7636_8799.n205 161.3
R131 a_n7636_8799.n74 a_n7636_8799.n18 74.4178
R132 a_n7636_8799.n213 a_n7636_8799.n74 12.4674
R133 a_n7636_8799.n73 a_n7636_8799.n18 80.107
R134 a_n7636_8799.n73 a_n7636_8799.n214 1.08907
R135 a_n7636_8799.n19 a_n7636_8799.n72 75.3623
R136 a_n7636_8799.n71 a_n7636_8799.n19 70.3058
R137 a_n7636_8799.n21 a_n7636_8799.n70 70.1674
R138 a_n7636_8799.n70 a_n7636_8799.n209 20.9683
R139 a_n7636_8799.n69 a_n7636_8799.n21 75.0448
R140 a_n7636_8799.n217 a_n7636_8799.n69 11.2134
R141 a_n7636_8799.n68 a_n7636_8799.n20 80.4688
R142 a_n7636_8799.n20 a_n7636_8799.n67 74.73
R143 a_n7636_8799.n66 a_n7636_8799.n22 70.1674
R144 a_n7636_8799.n220 a_n7636_8799.n66 20.9683
R145 a_n7636_8799.n22 a_n7636_8799.n65 70.5844
R146 a_n7636_8799.n65 a_n7636_8799.n207 20.1342
R147 a_n7636_8799.n64 a_n7636_8799.n23 75.6825
R148 a_n7636_8799.n221 a_n7636_8799.n64 9.93802
R149 a_n7636_8799.n23 a_n7636_8799.n222 161.3
R150 a_n7636_8799.n13 a_n7636_8799.n85 70.1674
R151 a_n7636_8799.n139 a_n7636_8799.n85 20.9683
R152 a_n7636_8799.n84 a_n7636_8799.n13 74.4178
R153 a_n7636_8799.n84 a_n7636_8799.n124 12.4674
R154 a_n7636_8799.n12 a_n7636_8799.n83 80.107
R155 a_n7636_8799.n138 a_n7636_8799.n83 1.08907
R156 a_n7636_8799.n82 a_n7636_8799.n12 75.3623
R157 a_n7636_8799.n14 a_n7636_8799.n81 70.3058
R158 a_n7636_8799.n80 a_n7636_8799.n14 70.1674
R159 a_n7636_8799.n80 a_n7636_8799.n125 20.9683
R160 a_n7636_8799.n15 a_n7636_8799.n79 75.0448
R161 a_n7636_8799.n134 a_n7636_8799.n79 11.2134
R162 a_n7636_8799.n78 a_n7636_8799.n15 80.4688
R163 a_n7636_8799.n16 a_n7636_8799.n77 74.73
R164 a_n7636_8799.n76 a_n7636_8799.n16 70.1674
R165 a_n7636_8799.n76 a_n7636_8799.n126 20.9683
R166 a_n7636_8799.n17 a_n7636_8799.n75 70.5844
R167 a_n7636_8799.n130 a_n7636_8799.n75 20.1342
R168 a_n7636_8799.n129 a_n7636_8799.n17 161.3
R169 a_n7636_8799.n7 a_n7636_8799.n96 70.1674
R170 a_n7636_8799.n155 a_n7636_8799.n96 20.9683
R171 a_n7636_8799.n95 a_n7636_8799.n7 74.4178
R172 a_n7636_8799.n95 a_n7636_8799.n140 12.4674
R173 a_n7636_8799.n6 a_n7636_8799.n94 80.107
R174 a_n7636_8799.n154 a_n7636_8799.n94 1.08907
R175 a_n7636_8799.n93 a_n7636_8799.n6 75.3623
R176 a_n7636_8799.n8 a_n7636_8799.n92 70.3058
R177 a_n7636_8799.n91 a_n7636_8799.n8 70.1674
R178 a_n7636_8799.n91 a_n7636_8799.n141 20.9683
R179 a_n7636_8799.n9 a_n7636_8799.n90 75.0448
R180 a_n7636_8799.n150 a_n7636_8799.n90 11.2134
R181 a_n7636_8799.n89 a_n7636_8799.n9 80.4688
R182 a_n7636_8799.n10 a_n7636_8799.n88 74.73
R183 a_n7636_8799.n87 a_n7636_8799.n10 70.1674
R184 a_n7636_8799.n87 a_n7636_8799.n142 20.9683
R185 a_n7636_8799.n11 a_n7636_8799.n86 70.5844
R186 a_n7636_8799.n146 a_n7636_8799.n86 20.1342
R187 a_n7636_8799.n145 a_n7636_8799.n11 161.3
R188 a_n7636_8799.n1 a_n7636_8799.n107 70.1674
R189 a_n7636_8799.n172 a_n7636_8799.n107 20.9683
R190 a_n7636_8799.n106 a_n7636_8799.n1 74.4178
R191 a_n7636_8799.n106 a_n7636_8799.n157 12.4674
R192 a_n7636_8799.n0 a_n7636_8799.n105 80.107
R193 a_n7636_8799.n171 a_n7636_8799.n105 1.08907
R194 a_n7636_8799.n104 a_n7636_8799.n0 75.3623
R195 a_n7636_8799.n2 a_n7636_8799.n103 70.3058
R196 a_n7636_8799.n102 a_n7636_8799.n2 70.1674
R197 a_n7636_8799.n102 a_n7636_8799.n158 20.9683
R198 a_n7636_8799.n3 a_n7636_8799.n101 75.0448
R199 a_n7636_8799.n167 a_n7636_8799.n101 11.2134
R200 a_n7636_8799.n100 a_n7636_8799.n3 80.4688
R201 a_n7636_8799.n4 a_n7636_8799.n99 74.73
R202 a_n7636_8799.n98 a_n7636_8799.n4 70.1674
R203 a_n7636_8799.n98 a_n7636_8799.n159 20.9683
R204 a_n7636_8799.n5 a_n7636_8799.n97 70.5844
R205 a_n7636_8799.n163 a_n7636_8799.n97 20.1342
R206 a_n7636_8799.n162 a_n7636_8799.n5 161.3
R207 a_n7636_8799.n229 a_n7636_8799.n108 98.9633
R208 a_n7636_8799.n40 a_n7636_8799.n109 98.9631
R209 a_n7636_8799.n41 a_n7636_8799.n227 98.6055
R210 a_n7636_8799.n41 a_n7636_8799.n228 98.6055
R211 a_n7636_8799.n40 a_n7636_8799.n110 98.6055
R212 a_n7636_8799.n40 a_n7636_8799.n111 98.6055
R213 a_n7636_8799.n113 a_n7636_8799.n112 98.6055
R214 a_n7636_8799.n230 a_n7636_8799.n229 98.6054
R215 a_n7636_8799.n39 a_n7636_8799.n114 81.2902
R216 a_n7636_8799.n37 a_n7636_8799.n120 81.2902
R217 a_n7636_8799.n36 a_n7636_8799.n117 81.2902
R218 a_n7636_8799.n38 a_n7636_8799.n122 80.9324
R219 a_n7636_8799.n38 a_n7636_8799.n123 80.9324
R220 a_n7636_8799.n39 a_n7636_8799.n116 80.9324
R221 a_n7636_8799.n39 a_n7636_8799.n115 80.9324
R222 a_n7636_8799.n37 a_n7636_8799.n121 80.9324
R223 a_n7636_8799.n37 a_n7636_8799.n119 80.9324
R224 a_n7636_8799.n36 a_n7636_8799.n118 80.9324
R225 a_n7636_8799.n30 a_n7636_8799.n179 70.4033
R226 a_n7636_8799.n24 a_n7636_8799.n195 70.4033
R227 a_n7636_8799.n18 a_n7636_8799.n212 70.4033
R228 a_n7636_8799.n17 a_n7636_8799.n128 70.4033
R229 a_n7636_8799.n11 a_n7636_8799.n144 70.4033
R230 a_n7636_8799.n5 a_n7636_8799.n161 70.4033
R231 a_n7636_8799.n189 a_n7636_8799.n188 48.2005
R232 a_n7636_8799.n44 a_n7636_8799.n186 20.9683
R233 a_n7636_8799.n185 a_n7636_8799.n184 48.2005
R234 a_n7636_8799.n183 a_n7636_8799.n48 20.9683
R235 a_n7636_8799.n181 a_n7636_8799.n177 48.2005
R236 a_n7636_8799.n205 a_n7636_8799.n204 48.2005
R237 a_n7636_8799.n55 a_n7636_8799.n202 20.9683
R238 a_n7636_8799.n201 a_n7636_8799.n200 48.2005
R239 a_n7636_8799.n199 a_n7636_8799.n59 20.9683
R240 a_n7636_8799.n197 a_n7636_8799.n193 48.2005
R241 a_n7636_8799.n222 a_n7636_8799.n221 48.2005
R242 a_n7636_8799.n66 a_n7636_8799.n219 20.9683
R243 a_n7636_8799.n218 a_n7636_8799.n217 48.2005
R244 a_n7636_8799.n216 a_n7636_8799.n70 20.9683
R245 a_n7636_8799.n214 a_n7636_8799.n210 48.2005
R246 a_n7636_8799.n131 a_n7636_8799.n76 20.9683
R247 a_n7636_8799.n134 a_n7636_8799.n133 48.2005
R248 a_n7636_8799.n135 a_n7636_8799.n80 20.9683
R249 a_n7636_8799.n138 a_n7636_8799.n137 48.2005
R250 a_n7636_8799.t45 a_n7636_8799.n85 485.135
R251 a_n7636_8799.n147 a_n7636_8799.n87 20.9683
R252 a_n7636_8799.n150 a_n7636_8799.n149 48.2005
R253 a_n7636_8799.n151 a_n7636_8799.n91 20.9683
R254 a_n7636_8799.n154 a_n7636_8799.n153 48.2005
R255 a_n7636_8799.t55 a_n7636_8799.n96 485.135
R256 a_n7636_8799.n164 a_n7636_8799.n98 20.9683
R257 a_n7636_8799.n167 a_n7636_8799.n166 48.2005
R258 a_n7636_8799.n168 a_n7636_8799.n102 20.9683
R259 a_n7636_8799.n171 a_n7636_8799.n170 48.2005
R260 a_n7636_8799.t106 a_n7636_8799.n107 485.135
R261 a_n7636_8799.n46 a_n7636_8799.n175 47.835
R262 a_n7636_8799.n49 a_n7636_8799.n182 20.6913
R263 a_n7636_8799.n57 a_n7636_8799.n191 47.835
R264 a_n7636_8799.n60 a_n7636_8799.n198 20.6913
R265 a_n7636_8799.n68 a_n7636_8799.n208 47.835
R266 a_n7636_8799.n71 a_n7636_8799.n215 20.6913
R267 a_n7636_8799.n132 a_n7636_8799.n78 47.835
R268 a_n7636_8799.n136 a_n7636_8799.n81 20.6913
R269 a_n7636_8799.n148 a_n7636_8799.n89 47.835
R270 a_n7636_8799.n152 a_n7636_8799.n92 20.6913
R271 a_n7636_8799.n165 a_n7636_8799.n100 47.835
R272 a_n7636_8799.n169 a_n7636_8799.n103 20.6913
R273 a_n7636_8799.n187 a_n7636_8799.n43 22.3251
R274 a_n7636_8799.n203 a_n7636_8799.n54 22.3251
R275 a_n7636_8799.n220 a_n7636_8799.n65 22.3251
R276 a_n7636_8799.n126 a_n7636_8799.n75 22.3251
R277 a_n7636_8799.n142 a_n7636_8799.n86 22.3251
R278 a_n7636_8799.n159 a_n7636_8799.n97 22.3251
R279 a_n7636_8799.n38 a_n7636_8799.n37 31.9767
R280 a_n7636_8799.n226 a_n7636_8799.n113 31.5713
R281 a_n7636_8799.n52 a_n7636_8799.n178 33.6462
R282 a_n7636_8799.n63 a_n7636_8799.n194 33.6462
R283 a_n7636_8799.n74 a_n7636_8799.n211 33.6462
R284 a_n7636_8799.n130 a_n7636_8799.n129 27.0217
R285 a_n7636_8799.n139 a_n7636_8799.n84 33.6462
R286 a_n7636_8799.n146 a_n7636_8799.n145 27.0217
R287 a_n7636_8799.n155 a_n7636_8799.n95 33.6462
R288 a_n7636_8799.n163 a_n7636_8799.n162 27.0217
R289 a_n7636_8799.n172 a_n7636_8799.n106 33.6462
R290 a_n7636_8799.n45 a_n7636_8799.n175 11.843
R291 a_n7636_8799.n182 a_n7636_8799.n50 36.139
R292 a_n7636_8799.n56 a_n7636_8799.n191 11.843
R293 a_n7636_8799.n198 a_n7636_8799.n61 36.139
R294 a_n7636_8799.n67 a_n7636_8799.n208 11.843
R295 a_n7636_8799.n215 a_n7636_8799.n72 36.139
R296 a_n7636_8799.n132 a_n7636_8799.n77 11.843
R297 a_n7636_8799.n136 a_n7636_8799.n82 36.139
R298 a_n7636_8799.n148 a_n7636_8799.n88 11.843
R299 a_n7636_8799.n152 a_n7636_8799.n93 36.139
R300 a_n7636_8799.n165 a_n7636_8799.n99 11.843
R301 a_n7636_8799.n169 a_n7636_8799.n104 36.139
R302 a_n7636_8799.n47 a_n7636_8799.n176 35.3134
R303 a_n7636_8799.n58 a_n7636_8799.n192 35.3134
R304 a_n7636_8799.n69 a_n7636_8799.n209 35.3134
R305 a_n7636_8799.n125 a_n7636_8799.n79 35.3134
R306 a_n7636_8799.n141 a_n7636_8799.n90 35.3134
R307 a_n7636_8799.n158 a_n7636_8799.n101 35.3134
R308 a_n7636_8799.n186 a_n7636_8799.n45 34.4824
R309 a_n7636_8799.n50 a_n7636_8799.n177 10.5784
R310 a_n7636_8799.n202 a_n7636_8799.n56 34.4824
R311 a_n7636_8799.n61 a_n7636_8799.n193 10.5784
R312 a_n7636_8799.n219 a_n7636_8799.n67 34.4824
R313 a_n7636_8799.n72 a_n7636_8799.n210 10.5784
R314 a_n7636_8799.n77 a_n7636_8799.n131 34.4824
R315 a_n7636_8799.n137 a_n7636_8799.n82 10.5784
R316 a_n7636_8799.n88 a_n7636_8799.n147 34.4824
R317 a_n7636_8799.n153 a_n7636_8799.n93 10.5784
R318 a_n7636_8799.n99 a_n7636_8799.n164 34.4824
R319 a_n7636_8799.n170 a_n7636_8799.n104 10.5784
R320 a_n7636_8799.n42 a_n7636_8799.n174 36.9592
R321 a_n7636_8799.n53 a_n7636_8799.n190 36.9592
R322 a_n7636_8799.n64 a_n7636_8799.n207 36.9592
R323 a_n7636_8799.n129 a_n7636_8799.n127 21.1793
R324 a_n7636_8799.n145 a_n7636_8799.n143 21.1793
R325 a_n7636_8799.n162 a_n7636_8799.n160 21.1793
R326 a_n7636_8799.n179 a_n7636_8799.n178 20.9576
R327 a_n7636_8799.n195 a_n7636_8799.n194 20.9576
R328 a_n7636_8799.n212 a_n7636_8799.n211 20.9576
R329 a_n7636_8799.n128 a_n7636_8799.n127 20.9576
R330 a_n7636_8799.n144 a_n7636_8799.n143 20.9576
R331 a_n7636_8799.n161 a_n7636_8799.n160 20.9576
R332 a_n7636_8799.n41 a_n7636_8799.n226 19.0249
R333 a_n7636_8799.n225 a_n7636_8799.n39 12.3339
R334 a_n7636_8799.n226 a_n7636_8799.n225 11.4887
R335 a_n7636_8799.n206 a_n7636_8799.n35 9.07815
R336 a_n7636_8799.n156 a_n7636_8799.n13 9.07815
R337 a_n7636_8799.n224 a_n7636_8799.n173 6.94254
R338 a_n7636_8799.n224 a_n7636_8799.n223 6.64832
R339 a_n7636_8799.n206 a_n7636_8799.n29 4.9702
R340 a_n7636_8799.n223 a_n7636_8799.n23 4.9702
R341 a_n7636_8799.n156 a_n7636_8799.n7 4.9702
R342 a_n7636_8799.n173 a_n7636_8799.n1 4.9702
R343 a_n7636_8799.n223 a_n7636_8799.n206 4.10845
R344 a_n7636_8799.n173 a_n7636_8799.n156 4.10845
R345 a_n7636_8799.n227 a_n7636_8799.t3 3.61217
R346 a_n7636_8799.n227 a_n7636_8799.t8 3.61217
R347 a_n7636_8799.n228 a_n7636_8799.t30 3.61217
R348 a_n7636_8799.n228 a_n7636_8799.t16 3.61217
R349 a_n7636_8799.n108 a_n7636_8799.t12 3.61217
R350 a_n7636_8799.n108 a_n7636_8799.t29 3.61217
R351 a_n7636_8799.n109 a_n7636_8799.t23 3.61217
R352 a_n7636_8799.n109 a_n7636_8799.t7 3.61217
R353 a_n7636_8799.n110 a_n7636_8799.t32 3.61217
R354 a_n7636_8799.n110 a_n7636_8799.t6 3.61217
R355 a_n7636_8799.n111 a_n7636_8799.t31 3.61217
R356 a_n7636_8799.n111 a_n7636_8799.t28 3.61217
R357 a_n7636_8799.n112 a_n7636_8799.t18 3.61217
R358 a_n7636_8799.n112 a_n7636_8799.t21 3.61217
R359 a_n7636_8799.n230 a_n7636_8799.t19 3.61217
R360 a_n7636_8799.t1 a_n7636_8799.n230 3.61217
R361 a_n7636_8799.n225 a_n7636_8799.n224 3.4105
R362 a_n7636_8799.n122 a_n7636_8799.t20 2.82907
R363 a_n7636_8799.n122 a_n7636_8799.t4 2.82907
R364 a_n7636_8799.n123 a_n7636_8799.t5 2.82907
R365 a_n7636_8799.n123 a_n7636_8799.t13 2.82907
R366 a_n7636_8799.n116 a_n7636_8799.t11 2.82907
R367 a_n7636_8799.n116 a_n7636_8799.t34 2.82907
R368 a_n7636_8799.n115 a_n7636_8799.t15 2.82907
R369 a_n7636_8799.n115 a_n7636_8799.t17 2.82907
R370 a_n7636_8799.n114 a_n7636_8799.t14 2.82907
R371 a_n7636_8799.n114 a_n7636_8799.t33 2.82907
R372 a_n7636_8799.n120 a_n7636_8799.t27 2.82907
R373 a_n7636_8799.n120 a_n7636_8799.t22 2.82907
R374 a_n7636_8799.n121 a_n7636_8799.t0 2.82907
R375 a_n7636_8799.n121 a_n7636_8799.t2 2.82907
R376 a_n7636_8799.n119 a_n7636_8799.t24 2.82907
R377 a_n7636_8799.n119 a_n7636_8799.t9 2.82907
R378 a_n7636_8799.n118 a_n7636_8799.t35 2.82907
R379 a_n7636_8799.n118 a_n7636_8799.t26 2.82907
R380 a_n7636_8799.n117 a_n7636_8799.t10 2.82907
R381 a_n7636_8799.n117 a_n7636_8799.t25 2.82907
R382 a_n7636_8799.n51 a_n7636_8799.n180 47.0982
R383 a_n7636_8799.n62 a_n7636_8799.n196 47.0982
R384 a_n7636_8799.n73 a_n7636_8799.n213 47.0982
R385 a_n7636_8799.n124 a_n7636_8799.n83 47.0982
R386 a_n7636_8799.n140 a_n7636_8799.n94 47.0982
R387 a_n7636_8799.n157 a_n7636_8799.n105 47.0982
R388 a_n7636_8799.n46 a_n7636_8799.n185 0.365327
R389 a_n7636_8799.n183 a_n7636_8799.n49 21.4216
R390 a_n7636_8799.n57 a_n7636_8799.n201 0.365327
R391 a_n7636_8799.n199 a_n7636_8799.n60 21.4216
R392 a_n7636_8799.n68 a_n7636_8799.n218 0.365327
R393 a_n7636_8799.n216 a_n7636_8799.n71 21.4216
R394 a_n7636_8799.n133 a_n7636_8799.n78 0.365327
R395 a_n7636_8799.n81 a_n7636_8799.n135 21.4216
R396 a_n7636_8799.n149 a_n7636_8799.n89 0.365327
R397 a_n7636_8799.n92 a_n7636_8799.n151 21.4216
R398 a_n7636_8799.n166 a_n7636_8799.n100 0.365327
R399 a_n7636_8799.n103 a_n7636_8799.n168 21.4216
R400 a_n7636_8799.n31 a_n7636_8799.n30 1.13686
R401 a_n7636_8799.n25 a_n7636_8799.n24 1.13686
R402 a_n7636_8799.n19 a_n7636_8799.n18 1.13686
R403 a_n7636_8799.n13 a_n7636_8799.n12 1.13686
R404 a_n7636_8799.n7 a_n7636_8799.n6 1.13686
R405 a_n7636_8799.n1 a_n7636_8799.n0 1.13686
R406 a_n7636_8799.n39 a_n7636_8799.n38 1.07378
R407 a_n7636_8799.n35 a_n7636_8799.n34 0.758076
R408 a_n7636_8799.n32 a_n7636_8799.n34 0.758076
R409 a_n7636_8799.n33 a_n7636_8799.n32 0.758076
R410 a_n7636_8799.n33 a_n7636_8799.n31 0.758076
R411 a_n7636_8799.n29 a_n7636_8799.n28 0.758076
R412 a_n7636_8799.n26 a_n7636_8799.n28 0.758076
R413 a_n7636_8799.n27 a_n7636_8799.n26 0.758076
R414 a_n7636_8799.n27 a_n7636_8799.n25 0.758076
R415 a_n7636_8799.n23 a_n7636_8799.n22 0.758076
R416 a_n7636_8799.n20 a_n7636_8799.n22 0.758076
R417 a_n7636_8799.n21 a_n7636_8799.n20 0.758076
R418 a_n7636_8799.n21 a_n7636_8799.n19 0.758076
R419 a_n7636_8799.n16 a_n7636_8799.n17 0.758076
R420 a_n7636_8799.n15 a_n7636_8799.n16 0.758076
R421 a_n7636_8799.n14 a_n7636_8799.n15 0.758076
R422 a_n7636_8799.n12 a_n7636_8799.n14 0.758076
R423 a_n7636_8799.n10 a_n7636_8799.n11 0.758076
R424 a_n7636_8799.n9 a_n7636_8799.n10 0.758076
R425 a_n7636_8799.n8 a_n7636_8799.n9 0.758076
R426 a_n7636_8799.n6 a_n7636_8799.n8 0.758076
R427 a_n7636_8799.n4 a_n7636_8799.n5 0.758076
R428 a_n7636_8799.n3 a_n7636_8799.n4 0.758076
R429 a_n7636_8799.n2 a_n7636_8799.n3 0.758076
R430 a_n7636_8799.n0 a_n7636_8799.n2 0.758076
R431 a_n7636_8799.n229 a_n7636_8799.n41 0.716017
R432 a_n7636_8799.n113 a_n7636_8799.n40 0.716017
R433 a_n7636_8799.n37 a_n7636_8799.n36 0.716017
R434 vdd.n315 vdd.n279 756.745
R435 vdd.n260 vdd.n224 756.745
R436 vdd.n217 vdd.n181 756.745
R437 vdd.n162 vdd.n126 756.745
R438 vdd.n120 vdd.n84 756.745
R439 vdd.n65 vdd.n29 756.745
R440 vdd.n2046 vdd.n2010 756.745
R441 vdd.n2101 vdd.n2065 756.745
R442 vdd.n1948 vdd.n1912 756.745
R443 vdd.n2003 vdd.n1967 756.745
R444 vdd.n1851 vdd.n1815 756.745
R445 vdd.n1906 vdd.n1870 756.745
R446 vdd.n1224 vdd.t54 640.208
R447 vdd.n952 vdd.t96 640.208
R448 vdd.n1244 vdd.t69 640.208
R449 vdd.n943 vdd.t114 640.208
R450 vdd.n843 vdd.t72 640.208
R451 vdd.n2621 vdd.t111 640.208
R452 vdd.n804 vdd.t120 640.208
R453 vdd.n2618 vdd.t100 640.208
R454 vdd.n768 vdd.t50 640.208
R455 vdd.n1014 vdd.t104 640.208
R456 vdd.n1510 vdd.t87 592.009
R457 vdd.n1666 vdd.t79 592.009
R458 vdd.n1702 vdd.t90 592.009
R459 vdd.n2186 vdd.t62 592.009
R460 vdd.n1161 vdd.t93 592.009
R461 vdd.n1121 vdd.t108 592.009
R462 vdd.n405 vdd.t83 592.009
R463 vdd.n419 vdd.t117 592.009
R464 vdd.n431 vdd.t123 592.009
R465 vdd.n723 vdd.t66 592.009
R466 vdd.n686 vdd.t76 592.009
R467 vdd.n3105 vdd.t58 592.009
R468 vdd.n316 vdd.n315 585
R469 vdd.n314 vdd.n281 585
R470 vdd.n313 vdd.n312 585
R471 vdd.n284 vdd.n282 585
R472 vdd.n307 vdd.n306 585
R473 vdd.n305 vdd.n304 585
R474 vdd.n288 vdd.n287 585
R475 vdd.n299 vdd.n298 585
R476 vdd.n297 vdd.n296 585
R477 vdd.n292 vdd.n291 585
R478 vdd.n261 vdd.n260 585
R479 vdd.n259 vdd.n226 585
R480 vdd.n258 vdd.n257 585
R481 vdd.n229 vdd.n227 585
R482 vdd.n252 vdd.n251 585
R483 vdd.n250 vdd.n249 585
R484 vdd.n233 vdd.n232 585
R485 vdd.n244 vdd.n243 585
R486 vdd.n242 vdd.n241 585
R487 vdd.n237 vdd.n236 585
R488 vdd.n218 vdd.n217 585
R489 vdd.n216 vdd.n183 585
R490 vdd.n215 vdd.n214 585
R491 vdd.n186 vdd.n184 585
R492 vdd.n209 vdd.n208 585
R493 vdd.n207 vdd.n206 585
R494 vdd.n190 vdd.n189 585
R495 vdd.n201 vdd.n200 585
R496 vdd.n199 vdd.n198 585
R497 vdd.n194 vdd.n193 585
R498 vdd.n163 vdd.n162 585
R499 vdd.n161 vdd.n128 585
R500 vdd.n160 vdd.n159 585
R501 vdd.n131 vdd.n129 585
R502 vdd.n154 vdd.n153 585
R503 vdd.n152 vdd.n151 585
R504 vdd.n135 vdd.n134 585
R505 vdd.n146 vdd.n145 585
R506 vdd.n144 vdd.n143 585
R507 vdd.n139 vdd.n138 585
R508 vdd.n121 vdd.n120 585
R509 vdd.n119 vdd.n86 585
R510 vdd.n118 vdd.n117 585
R511 vdd.n89 vdd.n87 585
R512 vdd.n112 vdd.n111 585
R513 vdd.n110 vdd.n109 585
R514 vdd.n93 vdd.n92 585
R515 vdd.n104 vdd.n103 585
R516 vdd.n102 vdd.n101 585
R517 vdd.n97 vdd.n96 585
R518 vdd.n66 vdd.n65 585
R519 vdd.n64 vdd.n31 585
R520 vdd.n63 vdd.n62 585
R521 vdd.n34 vdd.n32 585
R522 vdd.n57 vdd.n56 585
R523 vdd.n55 vdd.n54 585
R524 vdd.n38 vdd.n37 585
R525 vdd.n49 vdd.n48 585
R526 vdd.n47 vdd.n46 585
R527 vdd.n42 vdd.n41 585
R528 vdd.n2047 vdd.n2046 585
R529 vdd.n2045 vdd.n2012 585
R530 vdd.n2044 vdd.n2043 585
R531 vdd.n2015 vdd.n2013 585
R532 vdd.n2038 vdd.n2037 585
R533 vdd.n2036 vdd.n2035 585
R534 vdd.n2019 vdd.n2018 585
R535 vdd.n2030 vdd.n2029 585
R536 vdd.n2028 vdd.n2027 585
R537 vdd.n2023 vdd.n2022 585
R538 vdd.n2102 vdd.n2101 585
R539 vdd.n2100 vdd.n2067 585
R540 vdd.n2099 vdd.n2098 585
R541 vdd.n2070 vdd.n2068 585
R542 vdd.n2093 vdd.n2092 585
R543 vdd.n2091 vdd.n2090 585
R544 vdd.n2074 vdd.n2073 585
R545 vdd.n2085 vdd.n2084 585
R546 vdd.n2083 vdd.n2082 585
R547 vdd.n2078 vdd.n2077 585
R548 vdd.n1949 vdd.n1948 585
R549 vdd.n1947 vdd.n1914 585
R550 vdd.n1946 vdd.n1945 585
R551 vdd.n1917 vdd.n1915 585
R552 vdd.n1940 vdd.n1939 585
R553 vdd.n1938 vdd.n1937 585
R554 vdd.n1921 vdd.n1920 585
R555 vdd.n1932 vdd.n1931 585
R556 vdd.n1930 vdd.n1929 585
R557 vdd.n1925 vdd.n1924 585
R558 vdd.n2004 vdd.n2003 585
R559 vdd.n2002 vdd.n1969 585
R560 vdd.n2001 vdd.n2000 585
R561 vdd.n1972 vdd.n1970 585
R562 vdd.n1995 vdd.n1994 585
R563 vdd.n1993 vdd.n1992 585
R564 vdd.n1976 vdd.n1975 585
R565 vdd.n1987 vdd.n1986 585
R566 vdd.n1985 vdd.n1984 585
R567 vdd.n1980 vdd.n1979 585
R568 vdd.n1852 vdd.n1851 585
R569 vdd.n1850 vdd.n1817 585
R570 vdd.n1849 vdd.n1848 585
R571 vdd.n1820 vdd.n1818 585
R572 vdd.n1843 vdd.n1842 585
R573 vdd.n1841 vdd.n1840 585
R574 vdd.n1824 vdd.n1823 585
R575 vdd.n1835 vdd.n1834 585
R576 vdd.n1833 vdd.n1832 585
R577 vdd.n1828 vdd.n1827 585
R578 vdd.n1907 vdd.n1906 585
R579 vdd.n1905 vdd.n1872 585
R580 vdd.n1904 vdd.n1903 585
R581 vdd.n1875 vdd.n1873 585
R582 vdd.n1898 vdd.n1897 585
R583 vdd.n1896 vdd.n1895 585
R584 vdd.n1879 vdd.n1878 585
R585 vdd.n1890 vdd.n1889 585
R586 vdd.n1888 vdd.n1887 585
R587 vdd.n1883 vdd.n1882 585
R588 vdd.n445 vdd.n370 462.44
R589 vdd.n3343 vdd.n372 462.44
R590 vdd.n3238 vdd.n657 462.44
R591 vdd.n3236 vdd.n660 462.44
R592 vdd.n2181 vdd.n1409 462.44
R593 vdd.n2184 vdd.n2183 462.44
R594 vdd.n1737 vdd.n1507 462.44
R595 vdd.n1734 vdd.n1505 462.44
R596 vdd.n293 vdd.t245 329.043
R597 vdd.n238 vdd.t223 329.043
R598 vdd.n195 vdd.t235 329.043
R599 vdd.n140 vdd.t210 329.043
R600 vdd.n98 vdd.t197 329.043
R601 vdd.n43 vdd.t178 329.043
R602 vdd.n2024 vdd.t256 329.043
R603 vdd.n2079 vdd.t166 329.043
R604 vdd.n1926 vdd.t246 329.043
R605 vdd.n1981 vdd.t145 329.043
R606 vdd.n1829 vdd.t180 329.043
R607 vdd.n1884 vdd.t198 329.043
R608 vdd.n1510 vdd.t89 319.788
R609 vdd.n1666 vdd.t82 319.788
R610 vdd.n1702 vdd.t92 319.788
R611 vdd.n2186 vdd.t64 319.788
R612 vdd.n1161 vdd.t94 319.788
R613 vdd.n1121 vdd.t109 319.788
R614 vdd.n405 vdd.t85 319.788
R615 vdd.n419 vdd.t118 319.788
R616 vdd.n431 vdd.t124 319.788
R617 vdd.n723 vdd.t68 319.788
R618 vdd.n686 vdd.t78 319.788
R619 vdd.n3105 vdd.t61 319.788
R620 vdd.n1511 vdd.t88 303.69
R621 vdd.n1667 vdd.t81 303.69
R622 vdd.n1703 vdd.t91 303.69
R623 vdd.n2187 vdd.t65 303.69
R624 vdd.n1162 vdd.t95 303.69
R625 vdd.n1122 vdd.t110 303.69
R626 vdd.n406 vdd.t86 303.69
R627 vdd.n420 vdd.t119 303.69
R628 vdd.n432 vdd.t125 303.69
R629 vdd.n724 vdd.t67 303.69
R630 vdd.n687 vdd.t77 303.69
R631 vdd.n3106 vdd.t60 303.69
R632 vdd.n2853 vdd.n898 291.221
R633 vdd.n3067 vdd.n778 291.221
R634 vdd.n3004 vdd.n775 291.221
R635 vdd.n2785 vdd.n2784 291.221
R636 vdd.n2581 vdd.n940 291.221
R637 vdd.n2512 vdd.n2511 291.221
R638 vdd.n1280 vdd.n1279 291.221
R639 vdd.n2332 vdd.n1046 291.221
R640 vdd.n2983 vdd.n776 291.221
R641 vdd.n3070 vdd.n3069 291.221
R642 vdd.n2689 vdd.n2615 291.221
R643 vdd.n2857 vdd.n902 291.221
R644 vdd.n2509 vdd.n950 291.221
R645 vdd.n948 vdd.n922 291.221
R646 vdd.n1358 vdd.n1087 291.221
R647 vdd.n2336 vdd.n1051 291.221
R648 vdd.n2985 vdd.n776 185
R649 vdd.n3068 vdd.n776 185
R650 vdd.n2987 vdd.n2986 185
R651 vdd.n2986 vdd.n774 185
R652 vdd.n2988 vdd.n810 185
R653 vdd.n2998 vdd.n810 185
R654 vdd.n2989 vdd.n819 185
R655 vdd.n819 vdd.n817 185
R656 vdd.n2991 vdd.n2990 185
R657 vdd.n2992 vdd.n2991 185
R658 vdd.n2944 vdd.n818 185
R659 vdd.n818 vdd.n814 185
R660 vdd.n2943 vdd.n2942 185
R661 vdd.n2942 vdd.n2941 185
R662 vdd.n821 vdd.n820 185
R663 vdd.n822 vdd.n821 185
R664 vdd.n2934 vdd.n2933 185
R665 vdd.n2935 vdd.n2934 185
R666 vdd.n2932 vdd.n831 185
R667 vdd.n831 vdd.n828 185
R668 vdd.n2931 vdd.n2930 185
R669 vdd.n2930 vdd.n2929 185
R670 vdd.n833 vdd.n832 185
R671 vdd.n841 vdd.n833 185
R672 vdd.n2922 vdd.n2921 185
R673 vdd.n2923 vdd.n2922 185
R674 vdd.n2919 vdd.n842 185
R675 vdd.n849 vdd.n842 185
R676 vdd.n2918 vdd.n2917 185
R677 vdd.n2917 vdd.n2916 185
R678 vdd.n845 vdd.n844 185
R679 vdd.n846 vdd.n845 185
R680 vdd.n2909 vdd.n2908 185
R681 vdd.n2910 vdd.n2909 185
R682 vdd.n2907 vdd.n856 185
R683 vdd.n856 vdd.n853 185
R684 vdd.n2906 vdd.n2905 185
R685 vdd.n2905 vdd.n2904 185
R686 vdd.n858 vdd.n857 185
R687 vdd.n866 vdd.n858 185
R688 vdd.n2897 vdd.n2896 185
R689 vdd.n2898 vdd.n2897 185
R690 vdd.n2895 vdd.n867 185
R691 vdd.n872 vdd.n867 185
R692 vdd.n2894 vdd.n2893 185
R693 vdd.n2893 vdd.n2892 185
R694 vdd.n869 vdd.n868 185
R695 vdd.n2764 vdd.n869 185
R696 vdd.n2885 vdd.n2884 185
R697 vdd.n2886 vdd.n2885 185
R698 vdd.n2883 vdd.n879 185
R699 vdd.n879 vdd.n876 185
R700 vdd.n2882 vdd.n2881 185
R701 vdd.n2881 vdd.n2880 185
R702 vdd.n881 vdd.n880 185
R703 vdd.n882 vdd.n881 185
R704 vdd.n2873 vdd.n2872 185
R705 vdd.n2874 vdd.n2873 185
R706 vdd.n2871 vdd.n891 185
R707 vdd.n891 vdd.n888 185
R708 vdd.n2870 vdd.n2869 185
R709 vdd.n2869 vdd.n2868 185
R710 vdd.n893 vdd.n892 185
R711 vdd.n2779 vdd.n893 185
R712 vdd.n2861 vdd.n2860 185
R713 vdd.n2862 vdd.n2861 185
R714 vdd.n2859 vdd.n902 185
R715 vdd.n902 vdd.n899 185
R716 vdd.n2858 vdd.n2857 185
R717 vdd.n904 vdd.n903 185
R718 vdd.n2625 vdd.n2624 185
R719 vdd.n2627 vdd.n2626 185
R720 vdd.n2629 vdd.n2628 185
R721 vdd.n2631 vdd.n2630 185
R722 vdd.n2633 vdd.n2632 185
R723 vdd.n2635 vdd.n2634 185
R724 vdd.n2637 vdd.n2636 185
R725 vdd.n2639 vdd.n2638 185
R726 vdd.n2641 vdd.n2640 185
R727 vdd.n2643 vdd.n2642 185
R728 vdd.n2645 vdd.n2644 185
R729 vdd.n2647 vdd.n2646 185
R730 vdd.n2649 vdd.n2648 185
R731 vdd.n2651 vdd.n2650 185
R732 vdd.n2653 vdd.n2652 185
R733 vdd.n2655 vdd.n2654 185
R734 vdd.n2657 vdd.n2656 185
R735 vdd.n2659 vdd.n2658 185
R736 vdd.n2661 vdd.n2660 185
R737 vdd.n2663 vdd.n2662 185
R738 vdd.n2665 vdd.n2664 185
R739 vdd.n2667 vdd.n2666 185
R740 vdd.n2669 vdd.n2668 185
R741 vdd.n2671 vdd.n2670 185
R742 vdd.n2673 vdd.n2672 185
R743 vdd.n2675 vdd.n2674 185
R744 vdd.n2677 vdd.n2676 185
R745 vdd.n2679 vdd.n2678 185
R746 vdd.n2681 vdd.n2680 185
R747 vdd.n2683 vdd.n2682 185
R748 vdd.n2685 vdd.n2684 185
R749 vdd.n2687 vdd.n2686 185
R750 vdd.n2688 vdd.n2615 185
R751 vdd.n2855 vdd.n2615 185
R752 vdd.n3071 vdd.n3070 185
R753 vdd.n3072 vdd.n767 185
R754 vdd.n3074 vdd.n3073 185
R755 vdd.n3076 vdd.n765 185
R756 vdd.n3078 vdd.n3077 185
R757 vdd.n3079 vdd.n764 185
R758 vdd.n3081 vdd.n3080 185
R759 vdd.n3083 vdd.n762 185
R760 vdd.n3085 vdd.n3084 185
R761 vdd.n3086 vdd.n761 185
R762 vdd.n3088 vdd.n3087 185
R763 vdd.n3090 vdd.n759 185
R764 vdd.n3092 vdd.n3091 185
R765 vdd.n3093 vdd.n758 185
R766 vdd.n3095 vdd.n3094 185
R767 vdd.n3097 vdd.n757 185
R768 vdd.n3098 vdd.n754 185
R769 vdd.n3101 vdd.n3100 185
R770 vdd.n755 vdd.n753 185
R771 vdd.n2957 vdd.n2956 185
R772 vdd.n2959 vdd.n2958 185
R773 vdd.n2961 vdd.n2953 185
R774 vdd.n2963 vdd.n2962 185
R775 vdd.n2964 vdd.n2952 185
R776 vdd.n2966 vdd.n2965 185
R777 vdd.n2968 vdd.n2950 185
R778 vdd.n2970 vdd.n2969 185
R779 vdd.n2971 vdd.n2949 185
R780 vdd.n2973 vdd.n2972 185
R781 vdd.n2975 vdd.n2947 185
R782 vdd.n2977 vdd.n2976 185
R783 vdd.n2978 vdd.n2946 185
R784 vdd.n2980 vdd.n2979 185
R785 vdd.n2982 vdd.n2945 185
R786 vdd.n2984 vdd.n2983 185
R787 vdd.n2983 vdd.n756 185
R788 vdd.n3069 vdd.n771 185
R789 vdd.n3069 vdd.n3068 185
R790 vdd.n2692 vdd.n773 185
R791 vdd.n774 vdd.n773 185
R792 vdd.n2693 vdd.n809 185
R793 vdd.n2998 vdd.n809 185
R794 vdd.n2695 vdd.n2694 185
R795 vdd.n2694 vdd.n817 185
R796 vdd.n2696 vdd.n816 185
R797 vdd.n2992 vdd.n816 185
R798 vdd.n2698 vdd.n2697 185
R799 vdd.n2697 vdd.n814 185
R800 vdd.n2699 vdd.n824 185
R801 vdd.n2941 vdd.n824 185
R802 vdd.n2701 vdd.n2700 185
R803 vdd.n2700 vdd.n822 185
R804 vdd.n2702 vdd.n830 185
R805 vdd.n2935 vdd.n830 185
R806 vdd.n2704 vdd.n2703 185
R807 vdd.n2703 vdd.n828 185
R808 vdd.n2705 vdd.n835 185
R809 vdd.n2929 vdd.n835 185
R810 vdd.n2707 vdd.n2706 185
R811 vdd.n2706 vdd.n841 185
R812 vdd.n2708 vdd.n840 185
R813 vdd.n2923 vdd.n840 185
R814 vdd.n2710 vdd.n2709 185
R815 vdd.n2709 vdd.n849 185
R816 vdd.n2711 vdd.n848 185
R817 vdd.n2916 vdd.n848 185
R818 vdd.n2713 vdd.n2712 185
R819 vdd.n2712 vdd.n846 185
R820 vdd.n2714 vdd.n855 185
R821 vdd.n2910 vdd.n855 185
R822 vdd.n2716 vdd.n2715 185
R823 vdd.n2715 vdd.n853 185
R824 vdd.n2717 vdd.n860 185
R825 vdd.n2904 vdd.n860 185
R826 vdd.n2719 vdd.n2718 185
R827 vdd.n2718 vdd.n866 185
R828 vdd.n2720 vdd.n865 185
R829 vdd.n2898 vdd.n865 185
R830 vdd.n2722 vdd.n2721 185
R831 vdd.n2721 vdd.n872 185
R832 vdd.n2723 vdd.n871 185
R833 vdd.n2892 vdd.n871 185
R834 vdd.n2766 vdd.n2765 185
R835 vdd.n2765 vdd.n2764 185
R836 vdd.n2767 vdd.n878 185
R837 vdd.n2886 vdd.n878 185
R838 vdd.n2769 vdd.n2768 185
R839 vdd.n2768 vdd.n876 185
R840 vdd.n2770 vdd.n884 185
R841 vdd.n2880 vdd.n884 185
R842 vdd.n2772 vdd.n2771 185
R843 vdd.n2771 vdd.n882 185
R844 vdd.n2773 vdd.n890 185
R845 vdd.n2874 vdd.n890 185
R846 vdd.n2775 vdd.n2774 185
R847 vdd.n2774 vdd.n888 185
R848 vdd.n2776 vdd.n895 185
R849 vdd.n2868 vdd.n895 185
R850 vdd.n2778 vdd.n2777 185
R851 vdd.n2779 vdd.n2778 185
R852 vdd.n2691 vdd.n901 185
R853 vdd.n2862 vdd.n901 185
R854 vdd.n2690 vdd.n2689 185
R855 vdd.n2689 vdd.n899 185
R856 vdd.n2181 vdd.n2180 185
R857 vdd.n2182 vdd.n2181 185
R858 vdd.n1410 vdd.n1408 185
R859 vdd.n1408 vdd.n1407 185
R860 vdd.n2176 vdd.n2175 185
R861 vdd.n2175 vdd.n2174 185
R862 vdd.n1413 vdd.n1412 185
R863 vdd.n1414 vdd.n1413 185
R864 vdd.n2163 vdd.n2162 185
R865 vdd.n2164 vdd.n2163 185
R866 vdd.n1422 vdd.n1421 185
R867 vdd.n2155 vdd.n1421 185
R868 vdd.n2158 vdd.n2157 185
R869 vdd.n2157 vdd.n2156 185
R870 vdd.n1425 vdd.n1424 185
R871 vdd.n1431 vdd.n1425 185
R872 vdd.n2146 vdd.n2145 185
R873 vdd.n2147 vdd.n2146 185
R874 vdd.n1433 vdd.n1432 185
R875 vdd.n2138 vdd.n1432 185
R876 vdd.n2141 vdd.n2140 185
R877 vdd.n2140 vdd.n2139 185
R878 vdd.n1436 vdd.n1435 185
R879 vdd.n1437 vdd.n1436 185
R880 vdd.n2129 vdd.n2128 185
R881 vdd.n2130 vdd.n2129 185
R882 vdd.n1445 vdd.n1444 185
R883 vdd.n1444 vdd.n1443 185
R884 vdd.n2124 vdd.n2123 185
R885 vdd.n2123 vdd.n2122 185
R886 vdd.n1448 vdd.n1447 185
R887 vdd.n1454 vdd.n1448 185
R888 vdd.n2113 vdd.n2112 185
R889 vdd.n2114 vdd.n2113 185
R890 vdd.n1456 vdd.n1455 185
R891 vdd.n1810 vdd.n1455 185
R892 vdd.n1813 vdd.n1812 185
R893 vdd.n1812 vdd.n1811 185
R894 vdd.n1459 vdd.n1458 185
R895 vdd.n1466 vdd.n1459 185
R896 vdd.n1801 vdd.n1800 185
R897 vdd.n1802 vdd.n1801 185
R898 vdd.n1468 vdd.n1467 185
R899 vdd.n1467 vdd.n1465 185
R900 vdd.n1796 vdd.n1795 185
R901 vdd.n1795 vdd.n1794 185
R902 vdd.n1471 vdd.n1470 185
R903 vdd.n1472 vdd.n1471 185
R904 vdd.n1785 vdd.n1784 185
R905 vdd.n1786 vdd.n1785 185
R906 vdd.n1479 vdd.n1478 185
R907 vdd.n1777 vdd.n1478 185
R908 vdd.n1780 vdd.n1779 185
R909 vdd.n1779 vdd.n1778 185
R910 vdd.n1482 vdd.n1481 185
R911 vdd.n1488 vdd.n1482 185
R912 vdd.n1768 vdd.n1767 185
R913 vdd.n1769 vdd.n1768 185
R914 vdd.n1490 vdd.n1489 185
R915 vdd.n1760 vdd.n1489 185
R916 vdd.n1763 vdd.n1762 185
R917 vdd.n1762 vdd.n1761 185
R918 vdd.n1493 vdd.n1492 185
R919 vdd.n1494 vdd.n1493 185
R920 vdd.n1751 vdd.n1750 185
R921 vdd.n1752 vdd.n1751 185
R922 vdd.n1502 vdd.n1501 185
R923 vdd.n1501 vdd.n1500 185
R924 vdd.n1746 vdd.n1745 185
R925 vdd.n1745 vdd.n1744 185
R926 vdd.n1505 vdd.n1504 185
R927 vdd.n1506 vdd.n1505 185
R928 vdd.n1734 vdd.n1733 185
R929 vdd.n1732 vdd.n1545 185
R930 vdd.n1547 vdd.n1544 185
R931 vdd.n1736 vdd.n1544 185
R932 vdd.n1728 vdd.n1549 185
R933 vdd.n1727 vdd.n1550 185
R934 vdd.n1726 vdd.n1551 185
R935 vdd.n1554 vdd.n1552 185
R936 vdd.n1722 vdd.n1555 185
R937 vdd.n1721 vdd.n1556 185
R938 vdd.n1720 vdd.n1557 185
R939 vdd.n1560 vdd.n1558 185
R940 vdd.n1716 vdd.n1561 185
R941 vdd.n1715 vdd.n1562 185
R942 vdd.n1714 vdd.n1563 185
R943 vdd.n1566 vdd.n1564 185
R944 vdd.n1710 vdd.n1567 185
R945 vdd.n1709 vdd.n1568 185
R946 vdd.n1708 vdd.n1569 185
R947 vdd.n1700 vdd.n1570 185
R948 vdd.n1704 vdd.n1701 185
R949 vdd.n1699 vdd.n1572 185
R950 vdd.n1698 vdd.n1573 185
R951 vdd.n1576 vdd.n1574 185
R952 vdd.n1694 vdd.n1577 185
R953 vdd.n1693 vdd.n1578 185
R954 vdd.n1692 vdd.n1579 185
R955 vdd.n1582 vdd.n1580 185
R956 vdd.n1688 vdd.n1583 185
R957 vdd.n1687 vdd.n1584 185
R958 vdd.n1686 vdd.n1585 185
R959 vdd.n1588 vdd.n1586 185
R960 vdd.n1682 vdd.n1589 185
R961 vdd.n1681 vdd.n1590 185
R962 vdd.n1680 vdd.n1591 185
R963 vdd.n1594 vdd.n1592 185
R964 vdd.n1676 vdd.n1595 185
R965 vdd.n1675 vdd.n1596 185
R966 vdd.n1674 vdd.n1597 185
R967 vdd.n1600 vdd.n1598 185
R968 vdd.n1670 vdd.n1601 185
R969 vdd.n1669 vdd.n1602 185
R970 vdd.n1668 vdd.n1665 185
R971 vdd.n1605 vdd.n1603 185
R972 vdd.n1661 vdd.n1606 185
R973 vdd.n1660 vdd.n1607 185
R974 vdd.n1659 vdd.n1608 185
R975 vdd.n1611 vdd.n1609 185
R976 vdd.n1655 vdd.n1612 185
R977 vdd.n1654 vdd.n1613 185
R978 vdd.n1653 vdd.n1614 185
R979 vdd.n1617 vdd.n1615 185
R980 vdd.n1649 vdd.n1618 185
R981 vdd.n1648 vdd.n1619 185
R982 vdd.n1647 vdd.n1620 185
R983 vdd.n1623 vdd.n1621 185
R984 vdd.n1643 vdd.n1624 185
R985 vdd.n1642 vdd.n1625 185
R986 vdd.n1641 vdd.n1626 185
R987 vdd.n1629 vdd.n1627 185
R988 vdd.n1637 vdd.n1630 185
R989 vdd.n1636 vdd.n1631 185
R990 vdd.n1635 vdd.n1632 185
R991 vdd.n1633 vdd.n1513 185
R992 vdd.n1738 vdd.n1737 185
R993 vdd.n1737 vdd.n1736 185
R994 vdd.n2185 vdd.n2184 185
R995 vdd.n2189 vdd.n1403 185
R996 vdd.n1402 vdd.n1396 185
R997 vdd.n1400 vdd.n1399 185
R998 vdd.n1398 vdd.n1192 185
R999 vdd.n2193 vdd.n1189 185
R1000 vdd.n2195 vdd.n2194 185
R1001 vdd.n2197 vdd.n1187 185
R1002 vdd.n2199 vdd.n2198 185
R1003 vdd.n2200 vdd.n1182 185
R1004 vdd.n2202 vdd.n2201 185
R1005 vdd.n2204 vdd.n1180 185
R1006 vdd.n2206 vdd.n2205 185
R1007 vdd.n2207 vdd.n1175 185
R1008 vdd.n2209 vdd.n2208 185
R1009 vdd.n2211 vdd.n1173 185
R1010 vdd.n2213 vdd.n2212 185
R1011 vdd.n2214 vdd.n1169 185
R1012 vdd.n2216 vdd.n2215 185
R1013 vdd.n2218 vdd.n1166 185
R1014 vdd.n2220 vdd.n2219 185
R1015 vdd.n1167 vdd.n1160 185
R1016 vdd.n2224 vdd.n1164 185
R1017 vdd.n2225 vdd.n1156 185
R1018 vdd.n2227 vdd.n2226 185
R1019 vdd.n2229 vdd.n1154 185
R1020 vdd.n2231 vdd.n2230 185
R1021 vdd.n2232 vdd.n1149 185
R1022 vdd.n2234 vdd.n2233 185
R1023 vdd.n2236 vdd.n1147 185
R1024 vdd.n2238 vdd.n2237 185
R1025 vdd.n2239 vdd.n1142 185
R1026 vdd.n2241 vdd.n2240 185
R1027 vdd.n2243 vdd.n1140 185
R1028 vdd.n2245 vdd.n2244 185
R1029 vdd.n2246 vdd.n1135 185
R1030 vdd.n2248 vdd.n2247 185
R1031 vdd.n2250 vdd.n1133 185
R1032 vdd.n2252 vdd.n2251 185
R1033 vdd.n2253 vdd.n1129 185
R1034 vdd.n2255 vdd.n2254 185
R1035 vdd.n2257 vdd.n1126 185
R1036 vdd.n2259 vdd.n2258 185
R1037 vdd.n1127 vdd.n1120 185
R1038 vdd.n2263 vdd.n1124 185
R1039 vdd.n2264 vdd.n1116 185
R1040 vdd.n2266 vdd.n2265 185
R1041 vdd.n2268 vdd.n1114 185
R1042 vdd.n2270 vdd.n2269 185
R1043 vdd.n2271 vdd.n1109 185
R1044 vdd.n2273 vdd.n2272 185
R1045 vdd.n2275 vdd.n1107 185
R1046 vdd.n2277 vdd.n2276 185
R1047 vdd.n2278 vdd.n1102 185
R1048 vdd.n2280 vdd.n2279 185
R1049 vdd.n2282 vdd.n1100 185
R1050 vdd.n2284 vdd.n2283 185
R1051 vdd.n2285 vdd.n1098 185
R1052 vdd.n2287 vdd.n2286 185
R1053 vdd.n2290 vdd.n2289 185
R1054 vdd.n2292 vdd.n2291 185
R1055 vdd.n2294 vdd.n1096 185
R1056 vdd.n2296 vdd.n2295 185
R1057 vdd.n1409 vdd.n1095 185
R1058 vdd.n2183 vdd.n1406 185
R1059 vdd.n2183 vdd.n2182 185
R1060 vdd.n1417 vdd.n1405 185
R1061 vdd.n1407 vdd.n1405 185
R1062 vdd.n2173 vdd.n2172 185
R1063 vdd.n2174 vdd.n2173 185
R1064 vdd.n1416 vdd.n1415 185
R1065 vdd.n1415 vdd.n1414 185
R1066 vdd.n2166 vdd.n2165 185
R1067 vdd.n2165 vdd.n2164 185
R1068 vdd.n1420 vdd.n1419 185
R1069 vdd.n2155 vdd.n1420 185
R1070 vdd.n2154 vdd.n2153 185
R1071 vdd.n2156 vdd.n2154 185
R1072 vdd.n1427 vdd.n1426 185
R1073 vdd.n1431 vdd.n1426 185
R1074 vdd.n2149 vdd.n2148 185
R1075 vdd.n2148 vdd.n2147 185
R1076 vdd.n1430 vdd.n1429 185
R1077 vdd.n2138 vdd.n1430 185
R1078 vdd.n2137 vdd.n2136 185
R1079 vdd.n2139 vdd.n2137 185
R1080 vdd.n1439 vdd.n1438 185
R1081 vdd.n1438 vdd.n1437 185
R1082 vdd.n2132 vdd.n2131 185
R1083 vdd.n2131 vdd.n2130 185
R1084 vdd.n1442 vdd.n1441 185
R1085 vdd.n1443 vdd.n1442 185
R1086 vdd.n2121 vdd.n2120 185
R1087 vdd.n2122 vdd.n2121 185
R1088 vdd.n1450 vdd.n1449 185
R1089 vdd.n1454 vdd.n1449 185
R1090 vdd.n2116 vdd.n2115 185
R1091 vdd.n2115 vdd.n2114 185
R1092 vdd.n1453 vdd.n1452 185
R1093 vdd.n1810 vdd.n1453 185
R1094 vdd.n1809 vdd.n1808 185
R1095 vdd.n1811 vdd.n1809 185
R1096 vdd.n1461 vdd.n1460 185
R1097 vdd.n1466 vdd.n1460 185
R1098 vdd.n1804 vdd.n1803 185
R1099 vdd.n1803 vdd.n1802 185
R1100 vdd.n1464 vdd.n1463 185
R1101 vdd.n1465 vdd.n1464 185
R1102 vdd.n1793 vdd.n1792 185
R1103 vdd.n1794 vdd.n1793 185
R1104 vdd.n1474 vdd.n1473 185
R1105 vdd.n1473 vdd.n1472 185
R1106 vdd.n1788 vdd.n1787 185
R1107 vdd.n1787 vdd.n1786 185
R1108 vdd.n1477 vdd.n1476 185
R1109 vdd.n1777 vdd.n1477 185
R1110 vdd.n1776 vdd.n1775 185
R1111 vdd.n1778 vdd.n1776 185
R1112 vdd.n1484 vdd.n1483 185
R1113 vdd.n1488 vdd.n1483 185
R1114 vdd.n1771 vdd.n1770 185
R1115 vdd.n1770 vdd.n1769 185
R1116 vdd.n1487 vdd.n1486 185
R1117 vdd.n1760 vdd.n1487 185
R1118 vdd.n1759 vdd.n1758 185
R1119 vdd.n1761 vdd.n1759 185
R1120 vdd.n1496 vdd.n1495 185
R1121 vdd.n1495 vdd.n1494 185
R1122 vdd.n1754 vdd.n1753 185
R1123 vdd.n1753 vdd.n1752 185
R1124 vdd.n1499 vdd.n1498 185
R1125 vdd.n1500 vdd.n1499 185
R1126 vdd.n1743 vdd.n1742 185
R1127 vdd.n1744 vdd.n1743 185
R1128 vdd.n1508 vdd.n1507 185
R1129 vdd.n1507 vdd.n1506 185
R1130 vdd.n942 vdd.n940 185
R1131 vdd.n2510 vdd.n940 185
R1132 vdd.n2432 vdd.n960 185
R1133 vdd.n960 vdd.n947 185
R1134 vdd.n2434 vdd.n2433 185
R1135 vdd.n2435 vdd.n2434 185
R1136 vdd.n2431 vdd.n959 185
R1137 vdd.n1309 vdd.n959 185
R1138 vdd.n2430 vdd.n2429 185
R1139 vdd.n2429 vdd.n2428 185
R1140 vdd.n962 vdd.n961 185
R1141 vdd.n963 vdd.n962 185
R1142 vdd.n2419 vdd.n2418 185
R1143 vdd.n2420 vdd.n2419 185
R1144 vdd.n2417 vdd.n973 185
R1145 vdd.n973 vdd.n970 185
R1146 vdd.n2416 vdd.n2415 185
R1147 vdd.n2415 vdd.n2414 185
R1148 vdd.n975 vdd.n974 185
R1149 vdd.n976 vdd.n975 185
R1150 vdd.n2407 vdd.n2406 185
R1151 vdd.n2408 vdd.n2407 185
R1152 vdd.n2405 vdd.n984 185
R1153 vdd.n989 vdd.n984 185
R1154 vdd.n2404 vdd.n2403 185
R1155 vdd.n2403 vdd.n2402 185
R1156 vdd.n986 vdd.n985 185
R1157 vdd.n995 vdd.n986 185
R1158 vdd.n2395 vdd.n2394 185
R1159 vdd.n2396 vdd.n2395 185
R1160 vdd.n2393 vdd.n996 185
R1161 vdd.n1330 vdd.n996 185
R1162 vdd.n2392 vdd.n2391 185
R1163 vdd.n2391 vdd.n2390 185
R1164 vdd.n998 vdd.n997 185
R1165 vdd.n999 vdd.n998 185
R1166 vdd.n2383 vdd.n2382 185
R1167 vdd.n2384 vdd.n2383 185
R1168 vdd.n2381 vdd.n1008 185
R1169 vdd.n1008 vdd.n1005 185
R1170 vdd.n2380 vdd.n2379 185
R1171 vdd.n2379 vdd.n2378 185
R1172 vdd.n1010 vdd.n1009 185
R1173 vdd.n1019 vdd.n1010 185
R1174 vdd.n2370 vdd.n2369 185
R1175 vdd.n2371 vdd.n2370 185
R1176 vdd.n2368 vdd.n1020 185
R1177 vdd.n1026 vdd.n1020 185
R1178 vdd.n2367 vdd.n2366 185
R1179 vdd.n2366 vdd.n2365 185
R1180 vdd.n1022 vdd.n1021 185
R1181 vdd.n1023 vdd.n1022 185
R1182 vdd.n2358 vdd.n2357 185
R1183 vdd.n2359 vdd.n2358 185
R1184 vdd.n2356 vdd.n1033 185
R1185 vdd.n1033 vdd.n1030 185
R1186 vdd.n2355 vdd.n2354 185
R1187 vdd.n2354 vdd.n2353 185
R1188 vdd.n1035 vdd.n1034 185
R1189 vdd.n1036 vdd.n1035 185
R1190 vdd.n2346 vdd.n2345 185
R1191 vdd.n2347 vdd.n2346 185
R1192 vdd.n2344 vdd.n1044 185
R1193 vdd.n1050 vdd.n1044 185
R1194 vdd.n2343 vdd.n2342 185
R1195 vdd.n2342 vdd.n2341 185
R1196 vdd.n1046 vdd.n1045 185
R1197 vdd.n1047 vdd.n1046 185
R1198 vdd.n2332 vdd.n2331 185
R1199 vdd.n2330 vdd.n1089 185
R1200 vdd.n2329 vdd.n1088 185
R1201 vdd.n2334 vdd.n1088 185
R1202 vdd.n2328 vdd.n2327 185
R1203 vdd.n2326 vdd.n2325 185
R1204 vdd.n2324 vdd.n2323 185
R1205 vdd.n2322 vdd.n2321 185
R1206 vdd.n2320 vdd.n2319 185
R1207 vdd.n2318 vdd.n2317 185
R1208 vdd.n2316 vdd.n2315 185
R1209 vdd.n2314 vdd.n2313 185
R1210 vdd.n2312 vdd.n2311 185
R1211 vdd.n2310 vdd.n2309 185
R1212 vdd.n2308 vdd.n2307 185
R1213 vdd.n2306 vdd.n2305 185
R1214 vdd.n2304 vdd.n2303 185
R1215 vdd.n2302 vdd.n2301 185
R1216 vdd.n2300 vdd.n2299 185
R1217 vdd.n1246 vdd.n1090 185
R1218 vdd.n1248 vdd.n1247 185
R1219 vdd.n1250 vdd.n1249 185
R1220 vdd.n1252 vdd.n1251 185
R1221 vdd.n1254 vdd.n1253 185
R1222 vdd.n1256 vdd.n1255 185
R1223 vdd.n1258 vdd.n1257 185
R1224 vdd.n1260 vdd.n1259 185
R1225 vdd.n1262 vdd.n1261 185
R1226 vdd.n1264 vdd.n1263 185
R1227 vdd.n1266 vdd.n1265 185
R1228 vdd.n1268 vdd.n1267 185
R1229 vdd.n1270 vdd.n1269 185
R1230 vdd.n1272 vdd.n1271 185
R1231 vdd.n1275 vdd.n1274 185
R1232 vdd.n1277 vdd.n1276 185
R1233 vdd.n1279 vdd.n1278 185
R1234 vdd.n2513 vdd.n2512 185
R1235 vdd.n2515 vdd.n2514 185
R1236 vdd.n2517 vdd.n2516 185
R1237 vdd.n2520 vdd.n2519 185
R1238 vdd.n2522 vdd.n2521 185
R1239 vdd.n2524 vdd.n2523 185
R1240 vdd.n2526 vdd.n2525 185
R1241 vdd.n2528 vdd.n2527 185
R1242 vdd.n2530 vdd.n2529 185
R1243 vdd.n2532 vdd.n2531 185
R1244 vdd.n2534 vdd.n2533 185
R1245 vdd.n2536 vdd.n2535 185
R1246 vdd.n2538 vdd.n2537 185
R1247 vdd.n2540 vdd.n2539 185
R1248 vdd.n2542 vdd.n2541 185
R1249 vdd.n2544 vdd.n2543 185
R1250 vdd.n2546 vdd.n2545 185
R1251 vdd.n2548 vdd.n2547 185
R1252 vdd.n2550 vdd.n2549 185
R1253 vdd.n2552 vdd.n2551 185
R1254 vdd.n2554 vdd.n2553 185
R1255 vdd.n2556 vdd.n2555 185
R1256 vdd.n2558 vdd.n2557 185
R1257 vdd.n2560 vdd.n2559 185
R1258 vdd.n2562 vdd.n2561 185
R1259 vdd.n2564 vdd.n2563 185
R1260 vdd.n2566 vdd.n2565 185
R1261 vdd.n2568 vdd.n2567 185
R1262 vdd.n2570 vdd.n2569 185
R1263 vdd.n2572 vdd.n2571 185
R1264 vdd.n2574 vdd.n2573 185
R1265 vdd.n2576 vdd.n2575 185
R1266 vdd.n2578 vdd.n2577 185
R1267 vdd.n2579 vdd.n941 185
R1268 vdd.n2581 vdd.n2580 185
R1269 vdd.n2582 vdd.n2581 185
R1270 vdd.n2511 vdd.n945 185
R1271 vdd.n2511 vdd.n2510 185
R1272 vdd.n1307 vdd.n946 185
R1273 vdd.n947 vdd.n946 185
R1274 vdd.n1308 vdd.n957 185
R1275 vdd.n2435 vdd.n957 185
R1276 vdd.n1311 vdd.n1310 185
R1277 vdd.n1310 vdd.n1309 185
R1278 vdd.n1312 vdd.n964 185
R1279 vdd.n2428 vdd.n964 185
R1280 vdd.n1314 vdd.n1313 185
R1281 vdd.n1313 vdd.n963 185
R1282 vdd.n1315 vdd.n971 185
R1283 vdd.n2420 vdd.n971 185
R1284 vdd.n1317 vdd.n1316 185
R1285 vdd.n1316 vdd.n970 185
R1286 vdd.n1318 vdd.n977 185
R1287 vdd.n2414 vdd.n977 185
R1288 vdd.n1320 vdd.n1319 185
R1289 vdd.n1319 vdd.n976 185
R1290 vdd.n1321 vdd.n982 185
R1291 vdd.n2408 vdd.n982 185
R1292 vdd.n1323 vdd.n1322 185
R1293 vdd.n1322 vdd.n989 185
R1294 vdd.n1324 vdd.n987 185
R1295 vdd.n2402 vdd.n987 185
R1296 vdd.n1326 vdd.n1325 185
R1297 vdd.n1325 vdd.n995 185
R1298 vdd.n1327 vdd.n993 185
R1299 vdd.n2396 vdd.n993 185
R1300 vdd.n1329 vdd.n1328 185
R1301 vdd.n1330 vdd.n1329 185
R1302 vdd.n1306 vdd.n1000 185
R1303 vdd.n2390 vdd.n1000 185
R1304 vdd.n1305 vdd.n1304 185
R1305 vdd.n1304 vdd.n999 185
R1306 vdd.n1303 vdd.n1006 185
R1307 vdd.n2384 vdd.n1006 185
R1308 vdd.n1302 vdd.n1301 185
R1309 vdd.n1301 vdd.n1005 185
R1310 vdd.n1300 vdd.n1011 185
R1311 vdd.n2378 vdd.n1011 185
R1312 vdd.n1299 vdd.n1298 185
R1313 vdd.n1298 vdd.n1019 185
R1314 vdd.n1297 vdd.n1017 185
R1315 vdd.n2371 vdd.n1017 185
R1316 vdd.n1296 vdd.n1295 185
R1317 vdd.n1295 vdd.n1026 185
R1318 vdd.n1294 vdd.n1024 185
R1319 vdd.n2365 vdd.n1024 185
R1320 vdd.n1293 vdd.n1292 185
R1321 vdd.n1292 vdd.n1023 185
R1322 vdd.n1291 vdd.n1031 185
R1323 vdd.n2359 vdd.n1031 185
R1324 vdd.n1290 vdd.n1289 185
R1325 vdd.n1289 vdd.n1030 185
R1326 vdd.n1288 vdd.n1037 185
R1327 vdd.n2353 vdd.n1037 185
R1328 vdd.n1287 vdd.n1286 185
R1329 vdd.n1286 vdd.n1036 185
R1330 vdd.n1285 vdd.n1042 185
R1331 vdd.n2347 vdd.n1042 185
R1332 vdd.n1284 vdd.n1283 185
R1333 vdd.n1283 vdd.n1050 185
R1334 vdd.n1282 vdd.n1048 185
R1335 vdd.n2341 vdd.n1048 185
R1336 vdd.n1281 vdd.n1280 185
R1337 vdd.n1280 vdd.n1047 185
R1338 vdd.n370 vdd.n369 185
R1339 vdd.n3346 vdd.n370 185
R1340 vdd.n3349 vdd.n3348 185
R1341 vdd.n3348 vdd.n3347 185
R1342 vdd.n3350 vdd.n364 185
R1343 vdd.n364 vdd.n363 185
R1344 vdd.n3352 vdd.n3351 185
R1345 vdd.n3353 vdd.n3352 185
R1346 vdd.n359 vdd.n358 185
R1347 vdd.n3354 vdd.n359 185
R1348 vdd.n3357 vdd.n3356 185
R1349 vdd.n3356 vdd.n3355 185
R1350 vdd.n3358 vdd.n353 185
R1351 vdd.n3328 vdd.n353 185
R1352 vdd.n3360 vdd.n3359 185
R1353 vdd.n3361 vdd.n3360 185
R1354 vdd.n348 vdd.n347 185
R1355 vdd.n3362 vdd.n348 185
R1356 vdd.n3365 vdd.n3364 185
R1357 vdd.n3364 vdd.n3363 185
R1358 vdd.n3366 vdd.n342 185
R1359 vdd.n349 vdd.n342 185
R1360 vdd.n3368 vdd.n3367 185
R1361 vdd.n3369 vdd.n3368 185
R1362 vdd.n338 vdd.n337 185
R1363 vdd.n3370 vdd.n338 185
R1364 vdd.n3373 vdd.n3372 185
R1365 vdd.n3372 vdd.n3371 185
R1366 vdd.n3374 vdd.n333 185
R1367 vdd.n333 vdd.n332 185
R1368 vdd.n3376 vdd.n3375 185
R1369 vdd.n3377 vdd.n3376 185
R1370 vdd.n327 vdd.n325 185
R1371 vdd.n3378 vdd.n327 185
R1372 vdd.n3381 vdd.n3380 185
R1373 vdd.n3380 vdd.n3379 185
R1374 vdd.n326 vdd.n324 185
R1375 vdd.n328 vdd.n326 185
R1376 vdd.n3304 vdd.n3303 185
R1377 vdd.n3305 vdd.n3304 185
R1378 vdd.n615 vdd.n614 185
R1379 vdd.n614 vdd.n613 185
R1380 vdd.n3299 vdd.n3298 185
R1381 vdd.n3298 vdd.n3297 185
R1382 vdd.n618 vdd.n617 185
R1383 vdd.n624 vdd.n618 185
R1384 vdd.n3285 vdd.n3284 185
R1385 vdd.n3286 vdd.n3285 185
R1386 vdd.n626 vdd.n625 185
R1387 vdd.n3277 vdd.n625 185
R1388 vdd.n3280 vdd.n3279 185
R1389 vdd.n3279 vdd.n3278 185
R1390 vdd.n629 vdd.n628 185
R1391 vdd.n636 vdd.n629 185
R1392 vdd.n3268 vdd.n3267 185
R1393 vdd.n3269 vdd.n3268 185
R1394 vdd.n638 vdd.n637 185
R1395 vdd.n637 vdd.n635 185
R1396 vdd.n3263 vdd.n3262 185
R1397 vdd.n3262 vdd.n3261 185
R1398 vdd.n641 vdd.n640 185
R1399 vdd.n642 vdd.n641 185
R1400 vdd.n3252 vdd.n3251 185
R1401 vdd.n3253 vdd.n3252 185
R1402 vdd.n650 vdd.n649 185
R1403 vdd.n649 vdd.n648 185
R1404 vdd.n3247 vdd.n3246 185
R1405 vdd.n3246 vdd.n3245 185
R1406 vdd.n653 vdd.n652 185
R1407 vdd.n659 vdd.n653 185
R1408 vdd.n3236 vdd.n3235 185
R1409 vdd.n3237 vdd.n3236 185
R1410 vdd.n3232 vdd.n660 185
R1411 vdd.n3231 vdd.n3230 185
R1412 vdd.n3228 vdd.n662 185
R1413 vdd.n3228 vdd.n658 185
R1414 vdd.n3227 vdd.n3226 185
R1415 vdd.n3225 vdd.n3224 185
R1416 vdd.n3223 vdd.n3222 185
R1417 vdd.n3221 vdd.n3220 185
R1418 vdd.n3219 vdd.n668 185
R1419 vdd.n3217 vdd.n3216 185
R1420 vdd.n3215 vdd.n669 185
R1421 vdd.n3214 vdd.n3213 185
R1422 vdd.n3211 vdd.n674 185
R1423 vdd.n3209 vdd.n3208 185
R1424 vdd.n3207 vdd.n675 185
R1425 vdd.n3206 vdd.n3205 185
R1426 vdd.n3203 vdd.n680 185
R1427 vdd.n3201 vdd.n3200 185
R1428 vdd.n3199 vdd.n681 185
R1429 vdd.n3198 vdd.n3197 185
R1430 vdd.n3195 vdd.n688 185
R1431 vdd.n3193 vdd.n3192 185
R1432 vdd.n3191 vdd.n689 185
R1433 vdd.n3190 vdd.n3189 185
R1434 vdd.n3187 vdd.n694 185
R1435 vdd.n3185 vdd.n3184 185
R1436 vdd.n3183 vdd.n695 185
R1437 vdd.n3182 vdd.n3181 185
R1438 vdd.n3179 vdd.n700 185
R1439 vdd.n3177 vdd.n3176 185
R1440 vdd.n3175 vdd.n701 185
R1441 vdd.n3174 vdd.n3173 185
R1442 vdd.n3171 vdd.n706 185
R1443 vdd.n3169 vdd.n3168 185
R1444 vdd.n3167 vdd.n707 185
R1445 vdd.n3166 vdd.n3165 185
R1446 vdd.n3163 vdd.n712 185
R1447 vdd.n3161 vdd.n3160 185
R1448 vdd.n3159 vdd.n713 185
R1449 vdd.n3158 vdd.n3157 185
R1450 vdd.n3155 vdd.n718 185
R1451 vdd.n3153 vdd.n3152 185
R1452 vdd.n3151 vdd.n719 185
R1453 vdd.n728 vdd.n722 185
R1454 vdd.n3147 vdd.n3146 185
R1455 vdd.n3144 vdd.n726 185
R1456 vdd.n3143 vdd.n3142 185
R1457 vdd.n3141 vdd.n3140 185
R1458 vdd.n3139 vdd.n732 185
R1459 vdd.n3137 vdd.n3136 185
R1460 vdd.n3135 vdd.n733 185
R1461 vdd.n3134 vdd.n3133 185
R1462 vdd.n3131 vdd.n738 185
R1463 vdd.n3129 vdd.n3128 185
R1464 vdd.n3127 vdd.n739 185
R1465 vdd.n3126 vdd.n3125 185
R1466 vdd.n3123 vdd.n744 185
R1467 vdd.n3121 vdd.n3120 185
R1468 vdd.n3119 vdd.n745 185
R1469 vdd.n3118 vdd.n3117 185
R1470 vdd.n3115 vdd.n3114 185
R1471 vdd.n3113 vdd.n3112 185
R1472 vdd.n3111 vdd.n3110 185
R1473 vdd.n3109 vdd.n3108 185
R1474 vdd.n3104 vdd.n657 185
R1475 vdd.n658 vdd.n657 185
R1476 vdd.n3343 vdd.n3342 185
R1477 vdd.n599 vdd.n404 185
R1478 vdd.n598 vdd.n597 185
R1479 vdd.n596 vdd.n595 185
R1480 vdd.n594 vdd.n409 185
R1481 vdd.n590 vdd.n589 185
R1482 vdd.n588 vdd.n587 185
R1483 vdd.n586 vdd.n585 185
R1484 vdd.n584 vdd.n411 185
R1485 vdd.n580 vdd.n579 185
R1486 vdd.n578 vdd.n577 185
R1487 vdd.n576 vdd.n575 185
R1488 vdd.n574 vdd.n413 185
R1489 vdd.n570 vdd.n569 185
R1490 vdd.n568 vdd.n567 185
R1491 vdd.n566 vdd.n565 185
R1492 vdd.n564 vdd.n415 185
R1493 vdd.n560 vdd.n559 185
R1494 vdd.n558 vdd.n557 185
R1495 vdd.n556 vdd.n555 185
R1496 vdd.n554 vdd.n417 185
R1497 vdd.n550 vdd.n549 185
R1498 vdd.n548 vdd.n547 185
R1499 vdd.n546 vdd.n545 185
R1500 vdd.n544 vdd.n421 185
R1501 vdd.n540 vdd.n539 185
R1502 vdd.n538 vdd.n537 185
R1503 vdd.n536 vdd.n535 185
R1504 vdd.n534 vdd.n423 185
R1505 vdd.n530 vdd.n529 185
R1506 vdd.n528 vdd.n527 185
R1507 vdd.n526 vdd.n525 185
R1508 vdd.n524 vdd.n425 185
R1509 vdd.n520 vdd.n519 185
R1510 vdd.n518 vdd.n517 185
R1511 vdd.n516 vdd.n515 185
R1512 vdd.n514 vdd.n427 185
R1513 vdd.n510 vdd.n509 185
R1514 vdd.n508 vdd.n507 185
R1515 vdd.n506 vdd.n505 185
R1516 vdd.n504 vdd.n429 185
R1517 vdd.n500 vdd.n499 185
R1518 vdd.n498 vdd.n497 185
R1519 vdd.n496 vdd.n495 185
R1520 vdd.n494 vdd.n433 185
R1521 vdd.n490 vdd.n489 185
R1522 vdd.n488 vdd.n487 185
R1523 vdd.n486 vdd.n485 185
R1524 vdd.n484 vdd.n435 185
R1525 vdd.n480 vdd.n479 185
R1526 vdd.n478 vdd.n477 185
R1527 vdd.n476 vdd.n475 185
R1528 vdd.n474 vdd.n437 185
R1529 vdd.n470 vdd.n469 185
R1530 vdd.n468 vdd.n467 185
R1531 vdd.n466 vdd.n465 185
R1532 vdd.n464 vdd.n439 185
R1533 vdd.n460 vdd.n459 185
R1534 vdd.n458 vdd.n457 185
R1535 vdd.n456 vdd.n455 185
R1536 vdd.n454 vdd.n441 185
R1537 vdd.n450 vdd.n449 185
R1538 vdd.n448 vdd.n447 185
R1539 vdd.n446 vdd.n445 185
R1540 vdd.n3339 vdd.n372 185
R1541 vdd.n3346 vdd.n372 185
R1542 vdd.n3338 vdd.n371 185
R1543 vdd.n3347 vdd.n371 185
R1544 vdd.n3337 vdd.n3336 185
R1545 vdd.n3336 vdd.n363 185
R1546 vdd.n602 vdd.n362 185
R1547 vdd.n3353 vdd.n362 185
R1548 vdd.n3332 vdd.n361 185
R1549 vdd.n3354 vdd.n361 185
R1550 vdd.n3331 vdd.n360 185
R1551 vdd.n3355 vdd.n360 185
R1552 vdd.n3330 vdd.n3329 185
R1553 vdd.n3329 vdd.n3328 185
R1554 vdd.n604 vdd.n352 185
R1555 vdd.n3361 vdd.n352 185
R1556 vdd.n3324 vdd.n351 185
R1557 vdd.n3362 vdd.n351 185
R1558 vdd.n3323 vdd.n350 185
R1559 vdd.n3363 vdd.n350 185
R1560 vdd.n3322 vdd.n3321 185
R1561 vdd.n3321 vdd.n349 185
R1562 vdd.n606 vdd.n341 185
R1563 vdd.n3369 vdd.n341 185
R1564 vdd.n3317 vdd.n340 185
R1565 vdd.n3370 vdd.n340 185
R1566 vdd.n3316 vdd.n339 185
R1567 vdd.n3371 vdd.n339 185
R1568 vdd.n3315 vdd.n3314 185
R1569 vdd.n3314 vdd.n332 185
R1570 vdd.n608 vdd.n331 185
R1571 vdd.n3377 vdd.n331 185
R1572 vdd.n3310 vdd.n330 185
R1573 vdd.n3378 vdd.n330 185
R1574 vdd.n3309 vdd.n329 185
R1575 vdd.n3379 vdd.n329 185
R1576 vdd.n3308 vdd.n3307 185
R1577 vdd.n3307 vdd.n328 185
R1578 vdd.n3306 vdd.n610 185
R1579 vdd.n3306 vdd.n3305 185
R1580 vdd.n3294 vdd.n612 185
R1581 vdd.n613 vdd.n612 185
R1582 vdd.n3296 vdd.n3295 185
R1583 vdd.n3297 vdd.n3296 185
R1584 vdd.n620 vdd.n619 185
R1585 vdd.n624 vdd.n619 185
R1586 vdd.n3288 vdd.n3287 185
R1587 vdd.n3287 vdd.n3286 185
R1588 vdd.n623 vdd.n622 185
R1589 vdd.n3277 vdd.n623 185
R1590 vdd.n3276 vdd.n3275 185
R1591 vdd.n3278 vdd.n3276 185
R1592 vdd.n631 vdd.n630 185
R1593 vdd.n636 vdd.n630 185
R1594 vdd.n3271 vdd.n3270 185
R1595 vdd.n3270 vdd.n3269 185
R1596 vdd.n634 vdd.n633 185
R1597 vdd.n635 vdd.n634 185
R1598 vdd.n3260 vdd.n3259 185
R1599 vdd.n3261 vdd.n3260 185
R1600 vdd.n644 vdd.n643 185
R1601 vdd.n643 vdd.n642 185
R1602 vdd.n3255 vdd.n3254 185
R1603 vdd.n3254 vdd.n3253 185
R1604 vdd.n647 vdd.n646 185
R1605 vdd.n648 vdd.n647 185
R1606 vdd.n3244 vdd.n3243 185
R1607 vdd.n3245 vdd.n3244 185
R1608 vdd.n655 vdd.n654 185
R1609 vdd.n659 vdd.n654 185
R1610 vdd.n3239 vdd.n3238 185
R1611 vdd.n3238 vdd.n3237 185
R1612 vdd.n2853 vdd.n2852 185
R1613 vdd.n2851 vdd.n2617 185
R1614 vdd.n2850 vdd.n2616 185
R1615 vdd.n2855 vdd.n2616 185
R1616 vdd.n2849 vdd.n2848 185
R1617 vdd.n2847 vdd.n2846 185
R1618 vdd.n2845 vdd.n2844 185
R1619 vdd.n2843 vdd.n2842 185
R1620 vdd.n2841 vdd.n2840 185
R1621 vdd.n2839 vdd.n2838 185
R1622 vdd.n2837 vdd.n2836 185
R1623 vdd.n2835 vdd.n2834 185
R1624 vdd.n2833 vdd.n2832 185
R1625 vdd.n2831 vdd.n2830 185
R1626 vdd.n2829 vdd.n2828 185
R1627 vdd.n2827 vdd.n2826 185
R1628 vdd.n2825 vdd.n2824 185
R1629 vdd.n2823 vdd.n2822 185
R1630 vdd.n2821 vdd.n2820 185
R1631 vdd.n2819 vdd.n2818 185
R1632 vdd.n2817 vdd.n2816 185
R1633 vdd.n2815 vdd.n2814 185
R1634 vdd.n2813 vdd.n2812 185
R1635 vdd.n2811 vdd.n2810 185
R1636 vdd.n2809 vdd.n2808 185
R1637 vdd.n2807 vdd.n2806 185
R1638 vdd.n2805 vdd.n2804 185
R1639 vdd.n2803 vdd.n2802 185
R1640 vdd.n2801 vdd.n2800 185
R1641 vdd.n2799 vdd.n2798 185
R1642 vdd.n2797 vdd.n2796 185
R1643 vdd.n2795 vdd.n2794 185
R1644 vdd.n2793 vdd.n2792 185
R1645 vdd.n2790 vdd.n2789 185
R1646 vdd.n2788 vdd.n2787 185
R1647 vdd.n2786 vdd.n2785 185
R1648 vdd.n3005 vdd.n3004 185
R1649 vdd.n3006 vdd.n803 185
R1650 vdd.n3008 vdd.n3007 185
R1651 vdd.n3010 vdd.n801 185
R1652 vdd.n3012 vdd.n3011 185
R1653 vdd.n3013 vdd.n800 185
R1654 vdd.n3015 vdd.n3014 185
R1655 vdd.n3017 vdd.n798 185
R1656 vdd.n3019 vdd.n3018 185
R1657 vdd.n3020 vdd.n797 185
R1658 vdd.n3022 vdd.n3021 185
R1659 vdd.n3024 vdd.n795 185
R1660 vdd.n3026 vdd.n3025 185
R1661 vdd.n3027 vdd.n794 185
R1662 vdd.n3029 vdd.n3028 185
R1663 vdd.n3031 vdd.n792 185
R1664 vdd.n3033 vdd.n3032 185
R1665 vdd.n3035 vdd.n791 185
R1666 vdd.n3037 vdd.n3036 185
R1667 vdd.n3039 vdd.n789 185
R1668 vdd.n3041 vdd.n3040 185
R1669 vdd.n3042 vdd.n788 185
R1670 vdd.n3044 vdd.n3043 185
R1671 vdd.n3046 vdd.n786 185
R1672 vdd.n3048 vdd.n3047 185
R1673 vdd.n3049 vdd.n785 185
R1674 vdd.n3051 vdd.n3050 185
R1675 vdd.n3053 vdd.n783 185
R1676 vdd.n3055 vdd.n3054 185
R1677 vdd.n3056 vdd.n782 185
R1678 vdd.n3058 vdd.n3057 185
R1679 vdd.n3060 vdd.n781 185
R1680 vdd.n3061 vdd.n780 185
R1681 vdd.n3064 vdd.n3063 185
R1682 vdd.n3065 vdd.n778 185
R1683 vdd.n778 vdd.n756 185
R1684 vdd.n3002 vdd.n775 185
R1685 vdd.n3068 vdd.n775 185
R1686 vdd.n3001 vdd.n3000 185
R1687 vdd.n3000 vdd.n774 185
R1688 vdd.n2999 vdd.n807 185
R1689 vdd.n2999 vdd.n2998 185
R1690 vdd.n2733 vdd.n808 185
R1691 vdd.n817 vdd.n808 185
R1692 vdd.n2734 vdd.n815 185
R1693 vdd.n2992 vdd.n815 185
R1694 vdd.n2736 vdd.n2735 185
R1695 vdd.n2735 vdd.n814 185
R1696 vdd.n2737 vdd.n823 185
R1697 vdd.n2941 vdd.n823 185
R1698 vdd.n2739 vdd.n2738 185
R1699 vdd.n2738 vdd.n822 185
R1700 vdd.n2740 vdd.n829 185
R1701 vdd.n2935 vdd.n829 185
R1702 vdd.n2742 vdd.n2741 185
R1703 vdd.n2741 vdd.n828 185
R1704 vdd.n2743 vdd.n834 185
R1705 vdd.n2929 vdd.n834 185
R1706 vdd.n2745 vdd.n2744 185
R1707 vdd.n2744 vdd.n841 185
R1708 vdd.n2746 vdd.n839 185
R1709 vdd.n2923 vdd.n839 185
R1710 vdd.n2748 vdd.n2747 185
R1711 vdd.n2747 vdd.n849 185
R1712 vdd.n2749 vdd.n847 185
R1713 vdd.n2916 vdd.n847 185
R1714 vdd.n2751 vdd.n2750 185
R1715 vdd.n2750 vdd.n846 185
R1716 vdd.n2752 vdd.n854 185
R1717 vdd.n2910 vdd.n854 185
R1718 vdd.n2754 vdd.n2753 185
R1719 vdd.n2753 vdd.n853 185
R1720 vdd.n2755 vdd.n859 185
R1721 vdd.n2904 vdd.n859 185
R1722 vdd.n2757 vdd.n2756 185
R1723 vdd.n2756 vdd.n866 185
R1724 vdd.n2758 vdd.n864 185
R1725 vdd.n2898 vdd.n864 185
R1726 vdd.n2760 vdd.n2759 185
R1727 vdd.n2759 vdd.n872 185
R1728 vdd.n2761 vdd.n870 185
R1729 vdd.n2892 vdd.n870 185
R1730 vdd.n2763 vdd.n2762 185
R1731 vdd.n2764 vdd.n2763 185
R1732 vdd.n2732 vdd.n877 185
R1733 vdd.n2886 vdd.n877 185
R1734 vdd.n2731 vdd.n2730 185
R1735 vdd.n2730 vdd.n876 185
R1736 vdd.n2729 vdd.n883 185
R1737 vdd.n2880 vdd.n883 185
R1738 vdd.n2728 vdd.n2727 185
R1739 vdd.n2727 vdd.n882 185
R1740 vdd.n2726 vdd.n889 185
R1741 vdd.n2874 vdd.n889 185
R1742 vdd.n2725 vdd.n2724 185
R1743 vdd.n2724 vdd.n888 185
R1744 vdd.n2620 vdd.n894 185
R1745 vdd.n2868 vdd.n894 185
R1746 vdd.n2781 vdd.n2780 185
R1747 vdd.n2780 vdd.n2779 185
R1748 vdd.n2782 vdd.n900 185
R1749 vdd.n2862 vdd.n900 185
R1750 vdd.n2784 vdd.n2783 185
R1751 vdd.n2784 vdd.n899 185
R1752 vdd.n898 vdd.n897 185
R1753 vdd.n899 vdd.n898 185
R1754 vdd.n2864 vdd.n2863 185
R1755 vdd.n2863 vdd.n2862 185
R1756 vdd.n2865 vdd.n896 185
R1757 vdd.n2779 vdd.n896 185
R1758 vdd.n2867 vdd.n2866 185
R1759 vdd.n2868 vdd.n2867 185
R1760 vdd.n887 vdd.n886 185
R1761 vdd.n888 vdd.n887 185
R1762 vdd.n2876 vdd.n2875 185
R1763 vdd.n2875 vdd.n2874 185
R1764 vdd.n2877 vdd.n885 185
R1765 vdd.n885 vdd.n882 185
R1766 vdd.n2879 vdd.n2878 185
R1767 vdd.n2880 vdd.n2879 185
R1768 vdd.n875 vdd.n874 185
R1769 vdd.n876 vdd.n875 185
R1770 vdd.n2888 vdd.n2887 185
R1771 vdd.n2887 vdd.n2886 185
R1772 vdd.n2889 vdd.n873 185
R1773 vdd.n2764 vdd.n873 185
R1774 vdd.n2891 vdd.n2890 185
R1775 vdd.n2892 vdd.n2891 185
R1776 vdd.n863 vdd.n862 185
R1777 vdd.n872 vdd.n863 185
R1778 vdd.n2900 vdd.n2899 185
R1779 vdd.n2899 vdd.n2898 185
R1780 vdd.n2901 vdd.n861 185
R1781 vdd.n866 vdd.n861 185
R1782 vdd.n2903 vdd.n2902 185
R1783 vdd.n2904 vdd.n2903 185
R1784 vdd.n852 vdd.n851 185
R1785 vdd.n853 vdd.n852 185
R1786 vdd.n2912 vdd.n2911 185
R1787 vdd.n2911 vdd.n2910 185
R1788 vdd.n2913 vdd.n850 185
R1789 vdd.n850 vdd.n846 185
R1790 vdd.n2915 vdd.n2914 185
R1791 vdd.n2916 vdd.n2915 185
R1792 vdd.n838 vdd.n837 185
R1793 vdd.n849 vdd.n838 185
R1794 vdd.n2925 vdd.n2924 185
R1795 vdd.n2924 vdd.n2923 185
R1796 vdd.n2926 vdd.n836 185
R1797 vdd.n841 vdd.n836 185
R1798 vdd.n2928 vdd.n2927 185
R1799 vdd.n2929 vdd.n2928 185
R1800 vdd.n827 vdd.n826 185
R1801 vdd.n828 vdd.n827 185
R1802 vdd.n2937 vdd.n2936 185
R1803 vdd.n2936 vdd.n2935 185
R1804 vdd.n2938 vdd.n825 185
R1805 vdd.n825 vdd.n822 185
R1806 vdd.n2940 vdd.n2939 185
R1807 vdd.n2941 vdd.n2940 185
R1808 vdd.n813 vdd.n812 185
R1809 vdd.n814 vdd.n813 185
R1810 vdd.n2994 vdd.n2993 185
R1811 vdd.n2993 vdd.n2992 185
R1812 vdd.n2995 vdd.n811 185
R1813 vdd.n817 vdd.n811 185
R1814 vdd.n2997 vdd.n2996 185
R1815 vdd.n2998 vdd.n2997 185
R1816 vdd.n779 vdd.n777 185
R1817 vdd.n777 vdd.n774 185
R1818 vdd.n3067 vdd.n3066 185
R1819 vdd.n3068 vdd.n3067 185
R1820 vdd.n2509 vdd.n2508 185
R1821 vdd.n2510 vdd.n2509 185
R1822 vdd.n951 vdd.n949 185
R1823 vdd.n949 vdd.n947 185
R1824 vdd.n2424 vdd.n958 185
R1825 vdd.n2435 vdd.n958 185
R1826 vdd.n2425 vdd.n967 185
R1827 vdd.n1309 vdd.n967 185
R1828 vdd.n2427 vdd.n2426 185
R1829 vdd.n2428 vdd.n2427 185
R1830 vdd.n2423 vdd.n966 185
R1831 vdd.n966 vdd.n963 185
R1832 vdd.n2422 vdd.n2421 185
R1833 vdd.n2421 vdd.n2420 185
R1834 vdd.n969 vdd.n968 185
R1835 vdd.n970 vdd.n969 185
R1836 vdd.n2413 vdd.n2412 185
R1837 vdd.n2414 vdd.n2413 185
R1838 vdd.n2411 vdd.n979 185
R1839 vdd.n979 vdd.n976 185
R1840 vdd.n2410 vdd.n2409 185
R1841 vdd.n2409 vdd.n2408 185
R1842 vdd.n981 vdd.n980 185
R1843 vdd.n989 vdd.n981 185
R1844 vdd.n2401 vdd.n2400 185
R1845 vdd.n2402 vdd.n2401 185
R1846 vdd.n2399 vdd.n990 185
R1847 vdd.n995 vdd.n990 185
R1848 vdd.n2398 vdd.n2397 185
R1849 vdd.n2397 vdd.n2396 185
R1850 vdd.n992 vdd.n991 185
R1851 vdd.n1330 vdd.n992 185
R1852 vdd.n2389 vdd.n2388 185
R1853 vdd.n2390 vdd.n2389 185
R1854 vdd.n2387 vdd.n1002 185
R1855 vdd.n1002 vdd.n999 185
R1856 vdd.n2386 vdd.n2385 185
R1857 vdd.n2385 vdd.n2384 185
R1858 vdd.n1004 vdd.n1003 185
R1859 vdd.n1005 vdd.n1004 185
R1860 vdd.n2377 vdd.n2376 185
R1861 vdd.n2378 vdd.n2377 185
R1862 vdd.n2374 vdd.n1013 185
R1863 vdd.n1019 vdd.n1013 185
R1864 vdd.n2373 vdd.n2372 185
R1865 vdd.n2372 vdd.n2371 185
R1866 vdd.n1016 vdd.n1015 185
R1867 vdd.n1026 vdd.n1016 185
R1868 vdd.n2364 vdd.n2363 185
R1869 vdd.n2365 vdd.n2364 185
R1870 vdd.n2362 vdd.n1027 185
R1871 vdd.n1027 vdd.n1023 185
R1872 vdd.n2361 vdd.n2360 185
R1873 vdd.n2360 vdd.n2359 185
R1874 vdd.n1029 vdd.n1028 185
R1875 vdd.n1030 vdd.n1029 185
R1876 vdd.n2352 vdd.n2351 185
R1877 vdd.n2353 vdd.n2352 185
R1878 vdd.n2350 vdd.n1039 185
R1879 vdd.n1039 vdd.n1036 185
R1880 vdd.n2349 vdd.n2348 185
R1881 vdd.n2348 vdd.n2347 185
R1882 vdd.n1041 vdd.n1040 185
R1883 vdd.n1050 vdd.n1041 185
R1884 vdd.n2340 vdd.n2339 185
R1885 vdd.n2341 vdd.n2340 185
R1886 vdd.n2338 vdd.n1051 185
R1887 vdd.n1051 vdd.n1047 185
R1888 vdd.n2440 vdd.n922 185
R1889 vdd.n2582 vdd.n922 185
R1890 vdd.n2442 vdd.n2441 185
R1891 vdd.n2444 vdd.n2443 185
R1892 vdd.n2446 vdd.n2445 185
R1893 vdd.n2448 vdd.n2447 185
R1894 vdd.n2450 vdd.n2449 185
R1895 vdd.n2452 vdd.n2451 185
R1896 vdd.n2454 vdd.n2453 185
R1897 vdd.n2456 vdd.n2455 185
R1898 vdd.n2458 vdd.n2457 185
R1899 vdd.n2460 vdd.n2459 185
R1900 vdd.n2462 vdd.n2461 185
R1901 vdd.n2464 vdd.n2463 185
R1902 vdd.n2466 vdd.n2465 185
R1903 vdd.n2468 vdd.n2467 185
R1904 vdd.n2470 vdd.n2469 185
R1905 vdd.n2472 vdd.n2471 185
R1906 vdd.n2474 vdd.n2473 185
R1907 vdd.n2476 vdd.n2475 185
R1908 vdd.n2478 vdd.n2477 185
R1909 vdd.n2480 vdd.n2479 185
R1910 vdd.n2482 vdd.n2481 185
R1911 vdd.n2484 vdd.n2483 185
R1912 vdd.n2486 vdd.n2485 185
R1913 vdd.n2488 vdd.n2487 185
R1914 vdd.n2490 vdd.n2489 185
R1915 vdd.n2492 vdd.n2491 185
R1916 vdd.n2494 vdd.n2493 185
R1917 vdd.n2496 vdd.n2495 185
R1918 vdd.n2498 vdd.n2497 185
R1919 vdd.n2500 vdd.n2499 185
R1920 vdd.n2502 vdd.n2501 185
R1921 vdd.n2504 vdd.n2503 185
R1922 vdd.n2506 vdd.n2505 185
R1923 vdd.n2507 vdd.n950 185
R1924 vdd.n2439 vdd.n948 185
R1925 vdd.n2510 vdd.n948 185
R1926 vdd.n2438 vdd.n2437 185
R1927 vdd.n2437 vdd.n947 185
R1928 vdd.n2436 vdd.n955 185
R1929 vdd.n2436 vdd.n2435 185
R1930 vdd.n1227 vdd.n956 185
R1931 vdd.n1309 vdd.n956 185
R1932 vdd.n1228 vdd.n965 185
R1933 vdd.n2428 vdd.n965 185
R1934 vdd.n1230 vdd.n1229 185
R1935 vdd.n1229 vdd.n963 185
R1936 vdd.n1231 vdd.n972 185
R1937 vdd.n2420 vdd.n972 185
R1938 vdd.n1233 vdd.n1232 185
R1939 vdd.n1232 vdd.n970 185
R1940 vdd.n1234 vdd.n978 185
R1941 vdd.n2414 vdd.n978 185
R1942 vdd.n1236 vdd.n1235 185
R1943 vdd.n1235 vdd.n976 185
R1944 vdd.n1237 vdd.n983 185
R1945 vdd.n2408 vdd.n983 185
R1946 vdd.n1239 vdd.n1238 185
R1947 vdd.n1238 vdd.n989 185
R1948 vdd.n1240 vdd.n988 185
R1949 vdd.n2402 vdd.n988 185
R1950 vdd.n1242 vdd.n1241 185
R1951 vdd.n1241 vdd.n995 185
R1952 vdd.n1243 vdd.n994 185
R1953 vdd.n2396 vdd.n994 185
R1954 vdd.n1332 vdd.n1331 185
R1955 vdd.n1331 vdd.n1330 185
R1956 vdd.n1333 vdd.n1001 185
R1957 vdd.n2390 vdd.n1001 185
R1958 vdd.n1335 vdd.n1334 185
R1959 vdd.n1334 vdd.n999 185
R1960 vdd.n1336 vdd.n1007 185
R1961 vdd.n2384 vdd.n1007 185
R1962 vdd.n1338 vdd.n1337 185
R1963 vdd.n1337 vdd.n1005 185
R1964 vdd.n1339 vdd.n1012 185
R1965 vdd.n2378 vdd.n1012 185
R1966 vdd.n1341 vdd.n1340 185
R1967 vdd.n1340 vdd.n1019 185
R1968 vdd.n1342 vdd.n1018 185
R1969 vdd.n2371 vdd.n1018 185
R1970 vdd.n1344 vdd.n1343 185
R1971 vdd.n1343 vdd.n1026 185
R1972 vdd.n1345 vdd.n1025 185
R1973 vdd.n2365 vdd.n1025 185
R1974 vdd.n1347 vdd.n1346 185
R1975 vdd.n1346 vdd.n1023 185
R1976 vdd.n1348 vdd.n1032 185
R1977 vdd.n2359 vdd.n1032 185
R1978 vdd.n1350 vdd.n1349 185
R1979 vdd.n1349 vdd.n1030 185
R1980 vdd.n1351 vdd.n1038 185
R1981 vdd.n2353 vdd.n1038 185
R1982 vdd.n1353 vdd.n1352 185
R1983 vdd.n1352 vdd.n1036 185
R1984 vdd.n1354 vdd.n1043 185
R1985 vdd.n2347 vdd.n1043 185
R1986 vdd.n1356 vdd.n1355 185
R1987 vdd.n1355 vdd.n1050 185
R1988 vdd.n1357 vdd.n1049 185
R1989 vdd.n2341 vdd.n1049 185
R1990 vdd.n1359 vdd.n1358 185
R1991 vdd.n1358 vdd.n1047 185
R1992 vdd.n2337 vdd.n2336 185
R1993 vdd.n1053 vdd.n1052 185
R1994 vdd.n1194 vdd.n1193 185
R1995 vdd.n1196 vdd.n1195 185
R1996 vdd.n1198 vdd.n1197 185
R1997 vdd.n1200 vdd.n1199 185
R1998 vdd.n1202 vdd.n1201 185
R1999 vdd.n1204 vdd.n1203 185
R2000 vdd.n1206 vdd.n1205 185
R2001 vdd.n1208 vdd.n1207 185
R2002 vdd.n1210 vdd.n1209 185
R2003 vdd.n1212 vdd.n1211 185
R2004 vdd.n1214 vdd.n1213 185
R2005 vdd.n1216 vdd.n1215 185
R2006 vdd.n1218 vdd.n1217 185
R2007 vdd.n1220 vdd.n1219 185
R2008 vdd.n1222 vdd.n1221 185
R2009 vdd.n1393 vdd.n1223 185
R2010 vdd.n1392 vdd.n1391 185
R2011 vdd.n1390 vdd.n1389 185
R2012 vdd.n1388 vdd.n1387 185
R2013 vdd.n1386 vdd.n1385 185
R2014 vdd.n1384 vdd.n1383 185
R2015 vdd.n1382 vdd.n1381 185
R2016 vdd.n1380 vdd.n1379 185
R2017 vdd.n1378 vdd.n1377 185
R2018 vdd.n1376 vdd.n1375 185
R2019 vdd.n1374 vdd.n1373 185
R2020 vdd.n1372 vdd.n1371 185
R2021 vdd.n1370 vdd.n1369 185
R2022 vdd.n1368 vdd.n1367 185
R2023 vdd.n1366 vdd.n1365 185
R2024 vdd.n1364 vdd.n1363 185
R2025 vdd.n1362 vdd.n1361 185
R2026 vdd.n1360 vdd.n1087 185
R2027 vdd.n2334 vdd.n1087 185
R2028 vdd.n2334 vdd.n1054 179.345
R2029 vdd.n756 vdd.n658 179.345
R2030 vdd.n315 vdd.n314 171.744
R2031 vdd.n314 vdd.n313 171.744
R2032 vdd.n313 vdd.n282 171.744
R2033 vdd.n306 vdd.n282 171.744
R2034 vdd.n306 vdd.n305 171.744
R2035 vdd.n305 vdd.n287 171.744
R2036 vdd.n298 vdd.n287 171.744
R2037 vdd.n298 vdd.n297 171.744
R2038 vdd.n297 vdd.n291 171.744
R2039 vdd.n260 vdd.n259 171.744
R2040 vdd.n259 vdd.n258 171.744
R2041 vdd.n258 vdd.n227 171.744
R2042 vdd.n251 vdd.n227 171.744
R2043 vdd.n251 vdd.n250 171.744
R2044 vdd.n250 vdd.n232 171.744
R2045 vdd.n243 vdd.n232 171.744
R2046 vdd.n243 vdd.n242 171.744
R2047 vdd.n242 vdd.n236 171.744
R2048 vdd.n217 vdd.n216 171.744
R2049 vdd.n216 vdd.n215 171.744
R2050 vdd.n215 vdd.n184 171.744
R2051 vdd.n208 vdd.n184 171.744
R2052 vdd.n208 vdd.n207 171.744
R2053 vdd.n207 vdd.n189 171.744
R2054 vdd.n200 vdd.n189 171.744
R2055 vdd.n200 vdd.n199 171.744
R2056 vdd.n199 vdd.n193 171.744
R2057 vdd.n162 vdd.n161 171.744
R2058 vdd.n161 vdd.n160 171.744
R2059 vdd.n160 vdd.n129 171.744
R2060 vdd.n153 vdd.n129 171.744
R2061 vdd.n153 vdd.n152 171.744
R2062 vdd.n152 vdd.n134 171.744
R2063 vdd.n145 vdd.n134 171.744
R2064 vdd.n145 vdd.n144 171.744
R2065 vdd.n144 vdd.n138 171.744
R2066 vdd.n120 vdd.n119 171.744
R2067 vdd.n119 vdd.n118 171.744
R2068 vdd.n118 vdd.n87 171.744
R2069 vdd.n111 vdd.n87 171.744
R2070 vdd.n111 vdd.n110 171.744
R2071 vdd.n110 vdd.n92 171.744
R2072 vdd.n103 vdd.n92 171.744
R2073 vdd.n103 vdd.n102 171.744
R2074 vdd.n102 vdd.n96 171.744
R2075 vdd.n65 vdd.n64 171.744
R2076 vdd.n64 vdd.n63 171.744
R2077 vdd.n63 vdd.n32 171.744
R2078 vdd.n56 vdd.n32 171.744
R2079 vdd.n56 vdd.n55 171.744
R2080 vdd.n55 vdd.n37 171.744
R2081 vdd.n48 vdd.n37 171.744
R2082 vdd.n48 vdd.n47 171.744
R2083 vdd.n47 vdd.n41 171.744
R2084 vdd.n2046 vdd.n2045 171.744
R2085 vdd.n2045 vdd.n2044 171.744
R2086 vdd.n2044 vdd.n2013 171.744
R2087 vdd.n2037 vdd.n2013 171.744
R2088 vdd.n2037 vdd.n2036 171.744
R2089 vdd.n2036 vdd.n2018 171.744
R2090 vdd.n2029 vdd.n2018 171.744
R2091 vdd.n2029 vdd.n2028 171.744
R2092 vdd.n2028 vdd.n2022 171.744
R2093 vdd.n2101 vdd.n2100 171.744
R2094 vdd.n2100 vdd.n2099 171.744
R2095 vdd.n2099 vdd.n2068 171.744
R2096 vdd.n2092 vdd.n2068 171.744
R2097 vdd.n2092 vdd.n2091 171.744
R2098 vdd.n2091 vdd.n2073 171.744
R2099 vdd.n2084 vdd.n2073 171.744
R2100 vdd.n2084 vdd.n2083 171.744
R2101 vdd.n2083 vdd.n2077 171.744
R2102 vdd.n1948 vdd.n1947 171.744
R2103 vdd.n1947 vdd.n1946 171.744
R2104 vdd.n1946 vdd.n1915 171.744
R2105 vdd.n1939 vdd.n1915 171.744
R2106 vdd.n1939 vdd.n1938 171.744
R2107 vdd.n1938 vdd.n1920 171.744
R2108 vdd.n1931 vdd.n1920 171.744
R2109 vdd.n1931 vdd.n1930 171.744
R2110 vdd.n1930 vdd.n1924 171.744
R2111 vdd.n2003 vdd.n2002 171.744
R2112 vdd.n2002 vdd.n2001 171.744
R2113 vdd.n2001 vdd.n1970 171.744
R2114 vdd.n1994 vdd.n1970 171.744
R2115 vdd.n1994 vdd.n1993 171.744
R2116 vdd.n1993 vdd.n1975 171.744
R2117 vdd.n1986 vdd.n1975 171.744
R2118 vdd.n1986 vdd.n1985 171.744
R2119 vdd.n1985 vdd.n1979 171.744
R2120 vdd.n1851 vdd.n1850 171.744
R2121 vdd.n1850 vdd.n1849 171.744
R2122 vdd.n1849 vdd.n1818 171.744
R2123 vdd.n1842 vdd.n1818 171.744
R2124 vdd.n1842 vdd.n1841 171.744
R2125 vdd.n1841 vdd.n1823 171.744
R2126 vdd.n1834 vdd.n1823 171.744
R2127 vdd.n1834 vdd.n1833 171.744
R2128 vdd.n1833 vdd.n1827 171.744
R2129 vdd.n1906 vdd.n1905 171.744
R2130 vdd.n1905 vdd.n1904 171.744
R2131 vdd.n1904 vdd.n1873 171.744
R2132 vdd.n1897 vdd.n1873 171.744
R2133 vdd.n1897 vdd.n1896 171.744
R2134 vdd.n1896 vdd.n1878 171.744
R2135 vdd.n1889 vdd.n1878 171.744
R2136 vdd.n1889 vdd.n1888 171.744
R2137 vdd.n1888 vdd.n1882 171.744
R2138 vdd.n449 vdd.n448 146.341
R2139 vdd.n455 vdd.n454 146.341
R2140 vdd.n459 vdd.n458 146.341
R2141 vdd.n465 vdd.n464 146.341
R2142 vdd.n469 vdd.n468 146.341
R2143 vdd.n475 vdd.n474 146.341
R2144 vdd.n479 vdd.n478 146.341
R2145 vdd.n485 vdd.n484 146.341
R2146 vdd.n489 vdd.n488 146.341
R2147 vdd.n495 vdd.n494 146.341
R2148 vdd.n499 vdd.n498 146.341
R2149 vdd.n505 vdd.n504 146.341
R2150 vdd.n509 vdd.n508 146.341
R2151 vdd.n515 vdd.n514 146.341
R2152 vdd.n519 vdd.n518 146.341
R2153 vdd.n525 vdd.n524 146.341
R2154 vdd.n529 vdd.n528 146.341
R2155 vdd.n535 vdd.n534 146.341
R2156 vdd.n539 vdd.n538 146.341
R2157 vdd.n545 vdd.n544 146.341
R2158 vdd.n549 vdd.n548 146.341
R2159 vdd.n555 vdd.n554 146.341
R2160 vdd.n559 vdd.n558 146.341
R2161 vdd.n565 vdd.n564 146.341
R2162 vdd.n569 vdd.n568 146.341
R2163 vdd.n575 vdd.n574 146.341
R2164 vdd.n579 vdd.n578 146.341
R2165 vdd.n585 vdd.n584 146.341
R2166 vdd.n589 vdd.n588 146.341
R2167 vdd.n595 vdd.n594 146.341
R2168 vdd.n597 vdd.n404 146.341
R2169 vdd.n3238 vdd.n654 146.341
R2170 vdd.n3244 vdd.n654 146.341
R2171 vdd.n3244 vdd.n647 146.341
R2172 vdd.n3254 vdd.n647 146.341
R2173 vdd.n3254 vdd.n643 146.341
R2174 vdd.n3260 vdd.n643 146.341
R2175 vdd.n3260 vdd.n634 146.341
R2176 vdd.n3270 vdd.n634 146.341
R2177 vdd.n3270 vdd.n630 146.341
R2178 vdd.n3276 vdd.n630 146.341
R2179 vdd.n3276 vdd.n623 146.341
R2180 vdd.n3287 vdd.n623 146.341
R2181 vdd.n3287 vdd.n619 146.341
R2182 vdd.n3296 vdd.n619 146.341
R2183 vdd.n3296 vdd.n612 146.341
R2184 vdd.n3306 vdd.n612 146.341
R2185 vdd.n3307 vdd.n3306 146.341
R2186 vdd.n3307 vdd.n329 146.341
R2187 vdd.n330 vdd.n329 146.341
R2188 vdd.n331 vdd.n330 146.341
R2189 vdd.n3314 vdd.n331 146.341
R2190 vdd.n3314 vdd.n339 146.341
R2191 vdd.n340 vdd.n339 146.341
R2192 vdd.n341 vdd.n340 146.341
R2193 vdd.n3321 vdd.n341 146.341
R2194 vdd.n3321 vdd.n350 146.341
R2195 vdd.n351 vdd.n350 146.341
R2196 vdd.n352 vdd.n351 146.341
R2197 vdd.n3329 vdd.n352 146.341
R2198 vdd.n3329 vdd.n360 146.341
R2199 vdd.n361 vdd.n360 146.341
R2200 vdd.n362 vdd.n361 146.341
R2201 vdd.n3336 vdd.n362 146.341
R2202 vdd.n3336 vdd.n371 146.341
R2203 vdd.n372 vdd.n371 146.341
R2204 vdd.n3230 vdd.n3228 146.341
R2205 vdd.n3228 vdd.n3227 146.341
R2206 vdd.n3224 vdd.n3223 146.341
R2207 vdd.n3220 vdd.n3219 146.341
R2208 vdd.n3217 vdd.n669 146.341
R2209 vdd.n3213 vdd.n3211 146.341
R2210 vdd.n3209 vdd.n675 146.341
R2211 vdd.n3205 vdd.n3203 146.341
R2212 vdd.n3201 vdd.n681 146.341
R2213 vdd.n3197 vdd.n3195 146.341
R2214 vdd.n3193 vdd.n689 146.341
R2215 vdd.n3189 vdd.n3187 146.341
R2216 vdd.n3185 vdd.n695 146.341
R2217 vdd.n3181 vdd.n3179 146.341
R2218 vdd.n3177 vdd.n701 146.341
R2219 vdd.n3173 vdd.n3171 146.341
R2220 vdd.n3169 vdd.n707 146.341
R2221 vdd.n3165 vdd.n3163 146.341
R2222 vdd.n3161 vdd.n713 146.341
R2223 vdd.n3157 vdd.n3155 146.341
R2224 vdd.n3153 vdd.n719 146.341
R2225 vdd.n3146 vdd.n728 146.341
R2226 vdd.n3144 vdd.n3143 146.341
R2227 vdd.n3140 vdd.n3139 146.341
R2228 vdd.n3137 vdd.n733 146.341
R2229 vdd.n3133 vdd.n3131 146.341
R2230 vdd.n3129 vdd.n739 146.341
R2231 vdd.n3125 vdd.n3123 146.341
R2232 vdd.n3121 vdd.n745 146.341
R2233 vdd.n3117 vdd.n3115 146.341
R2234 vdd.n3112 vdd.n3111 146.341
R2235 vdd.n3108 vdd.n657 146.341
R2236 vdd.n3236 vdd.n653 146.341
R2237 vdd.n3246 vdd.n653 146.341
R2238 vdd.n3246 vdd.n649 146.341
R2239 vdd.n3252 vdd.n649 146.341
R2240 vdd.n3252 vdd.n641 146.341
R2241 vdd.n3262 vdd.n641 146.341
R2242 vdd.n3262 vdd.n637 146.341
R2243 vdd.n3268 vdd.n637 146.341
R2244 vdd.n3268 vdd.n629 146.341
R2245 vdd.n3279 vdd.n629 146.341
R2246 vdd.n3279 vdd.n625 146.341
R2247 vdd.n3285 vdd.n625 146.341
R2248 vdd.n3285 vdd.n618 146.341
R2249 vdd.n3298 vdd.n618 146.341
R2250 vdd.n3298 vdd.n614 146.341
R2251 vdd.n3304 vdd.n614 146.341
R2252 vdd.n3304 vdd.n326 146.341
R2253 vdd.n3380 vdd.n326 146.341
R2254 vdd.n3380 vdd.n327 146.341
R2255 vdd.n3376 vdd.n327 146.341
R2256 vdd.n3376 vdd.n333 146.341
R2257 vdd.n3372 vdd.n333 146.341
R2258 vdd.n3372 vdd.n338 146.341
R2259 vdd.n3368 vdd.n338 146.341
R2260 vdd.n3368 vdd.n342 146.341
R2261 vdd.n3364 vdd.n342 146.341
R2262 vdd.n3364 vdd.n348 146.341
R2263 vdd.n3360 vdd.n348 146.341
R2264 vdd.n3360 vdd.n353 146.341
R2265 vdd.n3356 vdd.n353 146.341
R2266 vdd.n3356 vdd.n359 146.341
R2267 vdd.n3352 vdd.n359 146.341
R2268 vdd.n3352 vdd.n364 146.341
R2269 vdd.n3348 vdd.n364 146.341
R2270 vdd.n3348 vdd.n370 146.341
R2271 vdd.n2295 vdd.n2294 146.341
R2272 vdd.n2292 vdd.n2289 146.341
R2273 vdd.n2287 vdd.n1098 146.341
R2274 vdd.n2283 vdd.n2282 146.341
R2275 vdd.n2280 vdd.n1102 146.341
R2276 vdd.n2276 vdd.n2275 146.341
R2277 vdd.n2273 vdd.n1109 146.341
R2278 vdd.n2269 vdd.n2268 146.341
R2279 vdd.n2266 vdd.n1116 146.341
R2280 vdd.n1127 vdd.n1124 146.341
R2281 vdd.n2258 vdd.n2257 146.341
R2282 vdd.n2255 vdd.n1129 146.341
R2283 vdd.n2251 vdd.n2250 146.341
R2284 vdd.n2248 vdd.n1135 146.341
R2285 vdd.n2244 vdd.n2243 146.341
R2286 vdd.n2241 vdd.n1142 146.341
R2287 vdd.n2237 vdd.n2236 146.341
R2288 vdd.n2234 vdd.n1149 146.341
R2289 vdd.n2230 vdd.n2229 146.341
R2290 vdd.n2227 vdd.n1156 146.341
R2291 vdd.n1167 vdd.n1164 146.341
R2292 vdd.n2219 vdd.n2218 146.341
R2293 vdd.n2216 vdd.n1169 146.341
R2294 vdd.n2212 vdd.n2211 146.341
R2295 vdd.n2209 vdd.n1175 146.341
R2296 vdd.n2205 vdd.n2204 146.341
R2297 vdd.n2202 vdd.n1182 146.341
R2298 vdd.n2198 vdd.n2197 146.341
R2299 vdd.n2195 vdd.n1189 146.341
R2300 vdd.n1400 vdd.n1398 146.341
R2301 vdd.n1403 vdd.n1402 146.341
R2302 vdd.n1743 vdd.n1507 146.341
R2303 vdd.n1743 vdd.n1499 146.341
R2304 vdd.n1753 vdd.n1499 146.341
R2305 vdd.n1753 vdd.n1495 146.341
R2306 vdd.n1759 vdd.n1495 146.341
R2307 vdd.n1759 vdd.n1487 146.341
R2308 vdd.n1770 vdd.n1487 146.341
R2309 vdd.n1770 vdd.n1483 146.341
R2310 vdd.n1776 vdd.n1483 146.341
R2311 vdd.n1776 vdd.n1477 146.341
R2312 vdd.n1787 vdd.n1477 146.341
R2313 vdd.n1787 vdd.n1473 146.341
R2314 vdd.n1793 vdd.n1473 146.341
R2315 vdd.n1793 vdd.n1464 146.341
R2316 vdd.n1803 vdd.n1464 146.341
R2317 vdd.n1803 vdd.n1460 146.341
R2318 vdd.n1809 vdd.n1460 146.341
R2319 vdd.n1809 vdd.n1453 146.341
R2320 vdd.n2115 vdd.n1453 146.341
R2321 vdd.n2115 vdd.n1449 146.341
R2322 vdd.n2121 vdd.n1449 146.341
R2323 vdd.n2121 vdd.n1442 146.341
R2324 vdd.n2131 vdd.n1442 146.341
R2325 vdd.n2131 vdd.n1438 146.341
R2326 vdd.n2137 vdd.n1438 146.341
R2327 vdd.n2137 vdd.n1430 146.341
R2328 vdd.n2148 vdd.n1430 146.341
R2329 vdd.n2148 vdd.n1426 146.341
R2330 vdd.n2154 vdd.n1426 146.341
R2331 vdd.n2154 vdd.n1420 146.341
R2332 vdd.n2165 vdd.n1420 146.341
R2333 vdd.n2165 vdd.n1415 146.341
R2334 vdd.n2173 vdd.n1415 146.341
R2335 vdd.n2173 vdd.n1405 146.341
R2336 vdd.n2183 vdd.n1405 146.341
R2337 vdd.n1545 vdd.n1544 146.341
R2338 vdd.n1549 vdd.n1544 146.341
R2339 vdd.n1551 vdd.n1550 146.341
R2340 vdd.n1555 vdd.n1554 146.341
R2341 vdd.n1557 vdd.n1556 146.341
R2342 vdd.n1561 vdd.n1560 146.341
R2343 vdd.n1563 vdd.n1562 146.341
R2344 vdd.n1567 vdd.n1566 146.341
R2345 vdd.n1569 vdd.n1568 146.341
R2346 vdd.n1701 vdd.n1700 146.341
R2347 vdd.n1573 vdd.n1572 146.341
R2348 vdd.n1577 vdd.n1576 146.341
R2349 vdd.n1579 vdd.n1578 146.341
R2350 vdd.n1583 vdd.n1582 146.341
R2351 vdd.n1585 vdd.n1584 146.341
R2352 vdd.n1589 vdd.n1588 146.341
R2353 vdd.n1591 vdd.n1590 146.341
R2354 vdd.n1595 vdd.n1594 146.341
R2355 vdd.n1597 vdd.n1596 146.341
R2356 vdd.n1601 vdd.n1600 146.341
R2357 vdd.n1665 vdd.n1602 146.341
R2358 vdd.n1606 vdd.n1605 146.341
R2359 vdd.n1608 vdd.n1607 146.341
R2360 vdd.n1612 vdd.n1611 146.341
R2361 vdd.n1614 vdd.n1613 146.341
R2362 vdd.n1618 vdd.n1617 146.341
R2363 vdd.n1620 vdd.n1619 146.341
R2364 vdd.n1624 vdd.n1623 146.341
R2365 vdd.n1626 vdd.n1625 146.341
R2366 vdd.n1630 vdd.n1629 146.341
R2367 vdd.n1632 vdd.n1631 146.341
R2368 vdd.n1737 vdd.n1513 146.341
R2369 vdd.n1745 vdd.n1505 146.341
R2370 vdd.n1745 vdd.n1501 146.341
R2371 vdd.n1751 vdd.n1501 146.341
R2372 vdd.n1751 vdd.n1493 146.341
R2373 vdd.n1762 vdd.n1493 146.341
R2374 vdd.n1762 vdd.n1489 146.341
R2375 vdd.n1768 vdd.n1489 146.341
R2376 vdd.n1768 vdd.n1482 146.341
R2377 vdd.n1779 vdd.n1482 146.341
R2378 vdd.n1779 vdd.n1478 146.341
R2379 vdd.n1785 vdd.n1478 146.341
R2380 vdd.n1785 vdd.n1471 146.341
R2381 vdd.n1795 vdd.n1471 146.341
R2382 vdd.n1795 vdd.n1467 146.341
R2383 vdd.n1801 vdd.n1467 146.341
R2384 vdd.n1801 vdd.n1459 146.341
R2385 vdd.n1812 vdd.n1459 146.341
R2386 vdd.n1812 vdd.n1455 146.341
R2387 vdd.n2113 vdd.n1455 146.341
R2388 vdd.n2113 vdd.n1448 146.341
R2389 vdd.n2123 vdd.n1448 146.341
R2390 vdd.n2123 vdd.n1444 146.341
R2391 vdd.n2129 vdd.n1444 146.341
R2392 vdd.n2129 vdd.n1436 146.341
R2393 vdd.n2140 vdd.n1436 146.341
R2394 vdd.n2140 vdd.n1432 146.341
R2395 vdd.n2146 vdd.n1432 146.341
R2396 vdd.n2146 vdd.n1425 146.341
R2397 vdd.n2157 vdd.n1425 146.341
R2398 vdd.n2157 vdd.n1421 146.341
R2399 vdd.n2163 vdd.n1421 146.341
R2400 vdd.n2163 vdd.n1413 146.341
R2401 vdd.n2175 vdd.n1413 146.341
R2402 vdd.n2175 vdd.n1408 146.341
R2403 vdd.n2181 vdd.n1408 146.341
R2404 vdd.n1224 vdd.t57 127.284
R2405 vdd.n952 vdd.t98 127.284
R2406 vdd.n1244 vdd.t71 127.284
R2407 vdd.n943 vdd.t115 127.284
R2408 vdd.n843 vdd.t74 127.284
R2409 vdd.n843 vdd.t75 127.284
R2410 vdd.n2621 vdd.t113 127.284
R2411 vdd.n804 vdd.t121 127.284
R2412 vdd.n2618 vdd.t103 127.284
R2413 vdd.n768 vdd.t52 127.284
R2414 vdd.n1014 vdd.t106 127.284
R2415 vdd.n1014 vdd.t107 127.284
R2416 vdd.n22 vdd.n20 117.314
R2417 vdd.n17 vdd.n15 117.314
R2418 vdd.n27 vdd.n26 116.927
R2419 vdd.n24 vdd.n23 116.927
R2420 vdd.n22 vdd.n21 116.927
R2421 vdd.n17 vdd.n16 116.927
R2422 vdd.n19 vdd.n18 116.927
R2423 vdd.n27 vdd.n25 116.927
R2424 vdd.n1225 vdd.t56 111.188
R2425 vdd.n953 vdd.t99 111.188
R2426 vdd.n1245 vdd.t70 111.188
R2427 vdd.n944 vdd.t116 111.188
R2428 vdd.n2622 vdd.t112 111.188
R2429 vdd.n805 vdd.t122 111.188
R2430 vdd.n2619 vdd.t102 111.188
R2431 vdd.n769 vdd.t53 111.188
R2432 vdd.n2863 vdd.n898 99.5127
R2433 vdd.n2863 vdd.n896 99.5127
R2434 vdd.n2867 vdd.n896 99.5127
R2435 vdd.n2867 vdd.n887 99.5127
R2436 vdd.n2875 vdd.n887 99.5127
R2437 vdd.n2875 vdd.n885 99.5127
R2438 vdd.n2879 vdd.n885 99.5127
R2439 vdd.n2879 vdd.n875 99.5127
R2440 vdd.n2887 vdd.n875 99.5127
R2441 vdd.n2887 vdd.n873 99.5127
R2442 vdd.n2891 vdd.n873 99.5127
R2443 vdd.n2891 vdd.n863 99.5127
R2444 vdd.n2899 vdd.n863 99.5127
R2445 vdd.n2899 vdd.n861 99.5127
R2446 vdd.n2903 vdd.n861 99.5127
R2447 vdd.n2903 vdd.n852 99.5127
R2448 vdd.n2911 vdd.n852 99.5127
R2449 vdd.n2911 vdd.n850 99.5127
R2450 vdd.n2915 vdd.n850 99.5127
R2451 vdd.n2915 vdd.n838 99.5127
R2452 vdd.n2924 vdd.n838 99.5127
R2453 vdd.n2924 vdd.n836 99.5127
R2454 vdd.n2928 vdd.n836 99.5127
R2455 vdd.n2928 vdd.n827 99.5127
R2456 vdd.n2936 vdd.n827 99.5127
R2457 vdd.n2936 vdd.n825 99.5127
R2458 vdd.n2940 vdd.n825 99.5127
R2459 vdd.n2940 vdd.n813 99.5127
R2460 vdd.n2993 vdd.n813 99.5127
R2461 vdd.n2993 vdd.n811 99.5127
R2462 vdd.n2997 vdd.n811 99.5127
R2463 vdd.n2997 vdd.n777 99.5127
R2464 vdd.n3067 vdd.n777 99.5127
R2465 vdd.n3063 vdd.n778 99.5127
R2466 vdd.n3061 vdd.n3060 99.5127
R2467 vdd.n3058 vdd.n782 99.5127
R2468 vdd.n3054 vdd.n3053 99.5127
R2469 vdd.n3051 vdd.n785 99.5127
R2470 vdd.n3047 vdd.n3046 99.5127
R2471 vdd.n3044 vdd.n788 99.5127
R2472 vdd.n3040 vdd.n3039 99.5127
R2473 vdd.n3037 vdd.n791 99.5127
R2474 vdd.n3032 vdd.n3031 99.5127
R2475 vdd.n3029 vdd.n794 99.5127
R2476 vdd.n3025 vdd.n3024 99.5127
R2477 vdd.n3022 vdd.n797 99.5127
R2478 vdd.n3018 vdd.n3017 99.5127
R2479 vdd.n3015 vdd.n800 99.5127
R2480 vdd.n3011 vdd.n3010 99.5127
R2481 vdd.n3008 vdd.n803 99.5127
R2482 vdd.n2784 vdd.n900 99.5127
R2483 vdd.n2780 vdd.n900 99.5127
R2484 vdd.n2780 vdd.n894 99.5127
R2485 vdd.n2724 vdd.n894 99.5127
R2486 vdd.n2724 vdd.n889 99.5127
R2487 vdd.n2727 vdd.n889 99.5127
R2488 vdd.n2727 vdd.n883 99.5127
R2489 vdd.n2730 vdd.n883 99.5127
R2490 vdd.n2730 vdd.n877 99.5127
R2491 vdd.n2763 vdd.n877 99.5127
R2492 vdd.n2763 vdd.n870 99.5127
R2493 vdd.n2759 vdd.n870 99.5127
R2494 vdd.n2759 vdd.n864 99.5127
R2495 vdd.n2756 vdd.n864 99.5127
R2496 vdd.n2756 vdd.n859 99.5127
R2497 vdd.n2753 vdd.n859 99.5127
R2498 vdd.n2753 vdd.n854 99.5127
R2499 vdd.n2750 vdd.n854 99.5127
R2500 vdd.n2750 vdd.n847 99.5127
R2501 vdd.n2747 vdd.n847 99.5127
R2502 vdd.n2747 vdd.n839 99.5127
R2503 vdd.n2744 vdd.n839 99.5127
R2504 vdd.n2744 vdd.n834 99.5127
R2505 vdd.n2741 vdd.n834 99.5127
R2506 vdd.n2741 vdd.n829 99.5127
R2507 vdd.n2738 vdd.n829 99.5127
R2508 vdd.n2738 vdd.n823 99.5127
R2509 vdd.n2735 vdd.n823 99.5127
R2510 vdd.n2735 vdd.n815 99.5127
R2511 vdd.n815 vdd.n808 99.5127
R2512 vdd.n2999 vdd.n808 99.5127
R2513 vdd.n3000 vdd.n2999 99.5127
R2514 vdd.n3000 vdd.n775 99.5127
R2515 vdd.n2617 vdd.n2616 99.5127
R2516 vdd.n2848 vdd.n2616 99.5127
R2517 vdd.n2846 vdd.n2845 99.5127
R2518 vdd.n2842 vdd.n2841 99.5127
R2519 vdd.n2838 vdd.n2837 99.5127
R2520 vdd.n2834 vdd.n2833 99.5127
R2521 vdd.n2830 vdd.n2829 99.5127
R2522 vdd.n2826 vdd.n2825 99.5127
R2523 vdd.n2822 vdd.n2821 99.5127
R2524 vdd.n2818 vdd.n2817 99.5127
R2525 vdd.n2814 vdd.n2813 99.5127
R2526 vdd.n2810 vdd.n2809 99.5127
R2527 vdd.n2806 vdd.n2805 99.5127
R2528 vdd.n2802 vdd.n2801 99.5127
R2529 vdd.n2798 vdd.n2797 99.5127
R2530 vdd.n2794 vdd.n2793 99.5127
R2531 vdd.n2789 vdd.n2788 99.5127
R2532 vdd.n2581 vdd.n941 99.5127
R2533 vdd.n2577 vdd.n2576 99.5127
R2534 vdd.n2573 vdd.n2572 99.5127
R2535 vdd.n2569 vdd.n2568 99.5127
R2536 vdd.n2565 vdd.n2564 99.5127
R2537 vdd.n2561 vdd.n2560 99.5127
R2538 vdd.n2557 vdd.n2556 99.5127
R2539 vdd.n2553 vdd.n2552 99.5127
R2540 vdd.n2549 vdd.n2548 99.5127
R2541 vdd.n2545 vdd.n2544 99.5127
R2542 vdd.n2541 vdd.n2540 99.5127
R2543 vdd.n2537 vdd.n2536 99.5127
R2544 vdd.n2533 vdd.n2532 99.5127
R2545 vdd.n2529 vdd.n2528 99.5127
R2546 vdd.n2525 vdd.n2524 99.5127
R2547 vdd.n2521 vdd.n2520 99.5127
R2548 vdd.n2516 vdd.n2515 99.5127
R2549 vdd.n1280 vdd.n1048 99.5127
R2550 vdd.n1283 vdd.n1048 99.5127
R2551 vdd.n1283 vdd.n1042 99.5127
R2552 vdd.n1286 vdd.n1042 99.5127
R2553 vdd.n1286 vdd.n1037 99.5127
R2554 vdd.n1289 vdd.n1037 99.5127
R2555 vdd.n1289 vdd.n1031 99.5127
R2556 vdd.n1292 vdd.n1031 99.5127
R2557 vdd.n1292 vdd.n1024 99.5127
R2558 vdd.n1295 vdd.n1024 99.5127
R2559 vdd.n1295 vdd.n1017 99.5127
R2560 vdd.n1298 vdd.n1017 99.5127
R2561 vdd.n1298 vdd.n1011 99.5127
R2562 vdd.n1301 vdd.n1011 99.5127
R2563 vdd.n1301 vdd.n1006 99.5127
R2564 vdd.n1304 vdd.n1006 99.5127
R2565 vdd.n1304 vdd.n1000 99.5127
R2566 vdd.n1329 vdd.n1000 99.5127
R2567 vdd.n1329 vdd.n993 99.5127
R2568 vdd.n1325 vdd.n993 99.5127
R2569 vdd.n1325 vdd.n987 99.5127
R2570 vdd.n1322 vdd.n987 99.5127
R2571 vdd.n1322 vdd.n982 99.5127
R2572 vdd.n1319 vdd.n982 99.5127
R2573 vdd.n1319 vdd.n977 99.5127
R2574 vdd.n1316 vdd.n977 99.5127
R2575 vdd.n1316 vdd.n971 99.5127
R2576 vdd.n1313 vdd.n971 99.5127
R2577 vdd.n1313 vdd.n964 99.5127
R2578 vdd.n1310 vdd.n964 99.5127
R2579 vdd.n1310 vdd.n957 99.5127
R2580 vdd.n957 vdd.n946 99.5127
R2581 vdd.n2511 vdd.n946 99.5127
R2582 vdd.n1089 vdd.n1088 99.5127
R2583 vdd.n2327 vdd.n1088 99.5127
R2584 vdd.n2325 vdd.n2324 99.5127
R2585 vdd.n2321 vdd.n2320 99.5127
R2586 vdd.n2317 vdd.n2316 99.5127
R2587 vdd.n2313 vdd.n2312 99.5127
R2588 vdd.n2309 vdd.n2308 99.5127
R2589 vdd.n2305 vdd.n2304 99.5127
R2590 vdd.n2301 vdd.n2300 99.5127
R2591 vdd.n1247 vdd.n1246 99.5127
R2592 vdd.n1251 vdd.n1250 99.5127
R2593 vdd.n1255 vdd.n1254 99.5127
R2594 vdd.n1259 vdd.n1258 99.5127
R2595 vdd.n1263 vdd.n1262 99.5127
R2596 vdd.n1267 vdd.n1266 99.5127
R2597 vdd.n1271 vdd.n1270 99.5127
R2598 vdd.n1276 vdd.n1275 99.5127
R2599 vdd.n2342 vdd.n1046 99.5127
R2600 vdd.n2342 vdd.n1044 99.5127
R2601 vdd.n2346 vdd.n1044 99.5127
R2602 vdd.n2346 vdd.n1035 99.5127
R2603 vdd.n2354 vdd.n1035 99.5127
R2604 vdd.n2354 vdd.n1033 99.5127
R2605 vdd.n2358 vdd.n1033 99.5127
R2606 vdd.n2358 vdd.n1022 99.5127
R2607 vdd.n2366 vdd.n1022 99.5127
R2608 vdd.n2366 vdd.n1020 99.5127
R2609 vdd.n2370 vdd.n1020 99.5127
R2610 vdd.n2370 vdd.n1010 99.5127
R2611 vdd.n2379 vdd.n1010 99.5127
R2612 vdd.n2379 vdd.n1008 99.5127
R2613 vdd.n2383 vdd.n1008 99.5127
R2614 vdd.n2383 vdd.n998 99.5127
R2615 vdd.n2391 vdd.n998 99.5127
R2616 vdd.n2391 vdd.n996 99.5127
R2617 vdd.n2395 vdd.n996 99.5127
R2618 vdd.n2395 vdd.n986 99.5127
R2619 vdd.n2403 vdd.n986 99.5127
R2620 vdd.n2403 vdd.n984 99.5127
R2621 vdd.n2407 vdd.n984 99.5127
R2622 vdd.n2407 vdd.n975 99.5127
R2623 vdd.n2415 vdd.n975 99.5127
R2624 vdd.n2415 vdd.n973 99.5127
R2625 vdd.n2419 vdd.n973 99.5127
R2626 vdd.n2419 vdd.n962 99.5127
R2627 vdd.n2429 vdd.n962 99.5127
R2628 vdd.n2429 vdd.n959 99.5127
R2629 vdd.n2434 vdd.n959 99.5127
R2630 vdd.n2434 vdd.n960 99.5127
R2631 vdd.n960 vdd.n940 99.5127
R2632 vdd.n2983 vdd.n2982 99.5127
R2633 vdd.n2980 vdd.n2946 99.5127
R2634 vdd.n2976 vdd.n2975 99.5127
R2635 vdd.n2973 vdd.n2949 99.5127
R2636 vdd.n2969 vdd.n2968 99.5127
R2637 vdd.n2966 vdd.n2952 99.5127
R2638 vdd.n2962 vdd.n2961 99.5127
R2639 vdd.n2959 vdd.n2956 99.5127
R2640 vdd.n3100 vdd.n755 99.5127
R2641 vdd.n3098 vdd.n3097 99.5127
R2642 vdd.n3095 vdd.n758 99.5127
R2643 vdd.n3091 vdd.n3090 99.5127
R2644 vdd.n3088 vdd.n761 99.5127
R2645 vdd.n3084 vdd.n3083 99.5127
R2646 vdd.n3081 vdd.n764 99.5127
R2647 vdd.n3077 vdd.n3076 99.5127
R2648 vdd.n3074 vdd.n767 99.5127
R2649 vdd.n2689 vdd.n901 99.5127
R2650 vdd.n2778 vdd.n901 99.5127
R2651 vdd.n2778 vdd.n895 99.5127
R2652 vdd.n2774 vdd.n895 99.5127
R2653 vdd.n2774 vdd.n890 99.5127
R2654 vdd.n2771 vdd.n890 99.5127
R2655 vdd.n2771 vdd.n884 99.5127
R2656 vdd.n2768 vdd.n884 99.5127
R2657 vdd.n2768 vdd.n878 99.5127
R2658 vdd.n2765 vdd.n878 99.5127
R2659 vdd.n2765 vdd.n871 99.5127
R2660 vdd.n2721 vdd.n871 99.5127
R2661 vdd.n2721 vdd.n865 99.5127
R2662 vdd.n2718 vdd.n865 99.5127
R2663 vdd.n2718 vdd.n860 99.5127
R2664 vdd.n2715 vdd.n860 99.5127
R2665 vdd.n2715 vdd.n855 99.5127
R2666 vdd.n2712 vdd.n855 99.5127
R2667 vdd.n2712 vdd.n848 99.5127
R2668 vdd.n2709 vdd.n848 99.5127
R2669 vdd.n2709 vdd.n840 99.5127
R2670 vdd.n2706 vdd.n840 99.5127
R2671 vdd.n2706 vdd.n835 99.5127
R2672 vdd.n2703 vdd.n835 99.5127
R2673 vdd.n2703 vdd.n830 99.5127
R2674 vdd.n2700 vdd.n830 99.5127
R2675 vdd.n2700 vdd.n824 99.5127
R2676 vdd.n2697 vdd.n824 99.5127
R2677 vdd.n2697 vdd.n816 99.5127
R2678 vdd.n2694 vdd.n816 99.5127
R2679 vdd.n2694 vdd.n809 99.5127
R2680 vdd.n809 vdd.n773 99.5127
R2681 vdd.n3069 vdd.n773 99.5127
R2682 vdd.n2624 vdd.n904 99.5127
R2683 vdd.n2628 vdd.n2627 99.5127
R2684 vdd.n2632 vdd.n2631 99.5127
R2685 vdd.n2636 vdd.n2635 99.5127
R2686 vdd.n2640 vdd.n2639 99.5127
R2687 vdd.n2644 vdd.n2643 99.5127
R2688 vdd.n2648 vdd.n2647 99.5127
R2689 vdd.n2652 vdd.n2651 99.5127
R2690 vdd.n2656 vdd.n2655 99.5127
R2691 vdd.n2660 vdd.n2659 99.5127
R2692 vdd.n2664 vdd.n2663 99.5127
R2693 vdd.n2668 vdd.n2667 99.5127
R2694 vdd.n2672 vdd.n2671 99.5127
R2695 vdd.n2676 vdd.n2675 99.5127
R2696 vdd.n2680 vdd.n2679 99.5127
R2697 vdd.n2684 vdd.n2683 99.5127
R2698 vdd.n2686 vdd.n2615 99.5127
R2699 vdd.n2861 vdd.n902 99.5127
R2700 vdd.n2861 vdd.n893 99.5127
R2701 vdd.n2869 vdd.n893 99.5127
R2702 vdd.n2869 vdd.n891 99.5127
R2703 vdd.n2873 vdd.n891 99.5127
R2704 vdd.n2873 vdd.n881 99.5127
R2705 vdd.n2881 vdd.n881 99.5127
R2706 vdd.n2881 vdd.n879 99.5127
R2707 vdd.n2885 vdd.n879 99.5127
R2708 vdd.n2885 vdd.n869 99.5127
R2709 vdd.n2893 vdd.n869 99.5127
R2710 vdd.n2893 vdd.n867 99.5127
R2711 vdd.n2897 vdd.n867 99.5127
R2712 vdd.n2897 vdd.n858 99.5127
R2713 vdd.n2905 vdd.n858 99.5127
R2714 vdd.n2905 vdd.n856 99.5127
R2715 vdd.n2909 vdd.n856 99.5127
R2716 vdd.n2909 vdd.n845 99.5127
R2717 vdd.n2917 vdd.n845 99.5127
R2718 vdd.n2917 vdd.n842 99.5127
R2719 vdd.n2922 vdd.n842 99.5127
R2720 vdd.n2922 vdd.n833 99.5127
R2721 vdd.n2930 vdd.n833 99.5127
R2722 vdd.n2930 vdd.n831 99.5127
R2723 vdd.n2934 vdd.n831 99.5127
R2724 vdd.n2934 vdd.n821 99.5127
R2725 vdd.n2942 vdd.n821 99.5127
R2726 vdd.n2942 vdd.n818 99.5127
R2727 vdd.n2991 vdd.n818 99.5127
R2728 vdd.n2991 vdd.n819 99.5127
R2729 vdd.n819 vdd.n810 99.5127
R2730 vdd.n2986 vdd.n810 99.5127
R2731 vdd.n2986 vdd.n776 99.5127
R2732 vdd.n2505 vdd.n2504 99.5127
R2733 vdd.n2501 vdd.n2500 99.5127
R2734 vdd.n2497 vdd.n2496 99.5127
R2735 vdd.n2493 vdd.n2492 99.5127
R2736 vdd.n2489 vdd.n2488 99.5127
R2737 vdd.n2485 vdd.n2484 99.5127
R2738 vdd.n2481 vdd.n2480 99.5127
R2739 vdd.n2477 vdd.n2476 99.5127
R2740 vdd.n2473 vdd.n2472 99.5127
R2741 vdd.n2469 vdd.n2468 99.5127
R2742 vdd.n2465 vdd.n2464 99.5127
R2743 vdd.n2461 vdd.n2460 99.5127
R2744 vdd.n2457 vdd.n2456 99.5127
R2745 vdd.n2453 vdd.n2452 99.5127
R2746 vdd.n2449 vdd.n2448 99.5127
R2747 vdd.n2445 vdd.n2444 99.5127
R2748 vdd.n2441 vdd.n922 99.5127
R2749 vdd.n1358 vdd.n1049 99.5127
R2750 vdd.n1355 vdd.n1049 99.5127
R2751 vdd.n1355 vdd.n1043 99.5127
R2752 vdd.n1352 vdd.n1043 99.5127
R2753 vdd.n1352 vdd.n1038 99.5127
R2754 vdd.n1349 vdd.n1038 99.5127
R2755 vdd.n1349 vdd.n1032 99.5127
R2756 vdd.n1346 vdd.n1032 99.5127
R2757 vdd.n1346 vdd.n1025 99.5127
R2758 vdd.n1343 vdd.n1025 99.5127
R2759 vdd.n1343 vdd.n1018 99.5127
R2760 vdd.n1340 vdd.n1018 99.5127
R2761 vdd.n1340 vdd.n1012 99.5127
R2762 vdd.n1337 vdd.n1012 99.5127
R2763 vdd.n1337 vdd.n1007 99.5127
R2764 vdd.n1334 vdd.n1007 99.5127
R2765 vdd.n1334 vdd.n1001 99.5127
R2766 vdd.n1331 vdd.n1001 99.5127
R2767 vdd.n1331 vdd.n994 99.5127
R2768 vdd.n1241 vdd.n994 99.5127
R2769 vdd.n1241 vdd.n988 99.5127
R2770 vdd.n1238 vdd.n988 99.5127
R2771 vdd.n1238 vdd.n983 99.5127
R2772 vdd.n1235 vdd.n983 99.5127
R2773 vdd.n1235 vdd.n978 99.5127
R2774 vdd.n1232 vdd.n978 99.5127
R2775 vdd.n1232 vdd.n972 99.5127
R2776 vdd.n1229 vdd.n972 99.5127
R2777 vdd.n1229 vdd.n965 99.5127
R2778 vdd.n965 vdd.n956 99.5127
R2779 vdd.n2436 vdd.n956 99.5127
R2780 vdd.n2437 vdd.n2436 99.5127
R2781 vdd.n2437 vdd.n948 99.5127
R2782 vdd.n1193 vdd.n1053 99.5127
R2783 vdd.n1197 vdd.n1196 99.5127
R2784 vdd.n1201 vdd.n1200 99.5127
R2785 vdd.n1205 vdd.n1204 99.5127
R2786 vdd.n1209 vdd.n1208 99.5127
R2787 vdd.n1213 vdd.n1212 99.5127
R2788 vdd.n1217 vdd.n1216 99.5127
R2789 vdd.n1221 vdd.n1220 99.5127
R2790 vdd.n1391 vdd.n1223 99.5127
R2791 vdd.n1389 vdd.n1388 99.5127
R2792 vdd.n1385 vdd.n1384 99.5127
R2793 vdd.n1381 vdd.n1380 99.5127
R2794 vdd.n1377 vdd.n1376 99.5127
R2795 vdd.n1373 vdd.n1372 99.5127
R2796 vdd.n1369 vdd.n1368 99.5127
R2797 vdd.n1365 vdd.n1364 99.5127
R2798 vdd.n1361 vdd.n1087 99.5127
R2799 vdd.n2340 vdd.n1051 99.5127
R2800 vdd.n2340 vdd.n1041 99.5127
R2801 vdd.n2348 vdd.n1041 99.5127
R2802 vdd.n2348 vdd.n1039 99.5127
R2803 vdd.n2352 vdd.n1039 99.5127
R2804 vdd.n2352 vdd.n1029 99.5127
R2805 vdd.n2360 vdd.n1029 99.5127
R2806 vdd.n2360 vdd.n1027 99.5127
R2807 vdd.n2364 vdd.n1027 99.5127
R2808 vdd.n2364 vdd.n1016 99.5127
R2809 vdd.n2372 vdd.n1016 99.5127
R2810 vdd.n2372 vdd.n1013 99.5127
R2811 vdd.n2377 vdd.n1013 99.5127
R2812 vdd.n2377 vdd.n1004 99.5127
R2813 vdd.n2385 vdd.n1004 99.5127
R2814 vdd.n2385 vdd.n1002 99.5127
R2815 vdd.n2389 vdd.n1002 99.5127
R2816 vdd.n2389 vdd.n992 99.5127
R2817 vdd.n2397 vdd.n992 99.5127
R2818 vdd.n2397 vdd.n990 99.5127
R2819 vdd.n2401 vdd.n990 99.5127
R2820 vdd.n2401 vdd.n981 99.5127
R2821 vdd.n2409 vdd.n981 99.5127
R2822 vdd.n2409 vdd.n979 99.5127
R2823 vdd.n2413 vdd.n979 99.5127
R2824 vdd.n2413 vdd.n969 99.5127
R2825 vdd.n2421 vdd.n969 99.5127
R2826 vdd.n2421 vdd.n966 99.5127
R2827 vdd.n2427 vdd.n966 99.5127
R2828 vdd.n2427 vdd.n967 99.5127
R2829 vdd.n967 vdd.n958 99.5127
R2830 vdd.n958 vdd.n949 99.5127
R2831 vdd.n2509 vdd.n949 99.5127
R2832 vdd.n9 vdd.n7 98.9633
R2833 vdd.n2 vdd.n0 98.9633
R2834 vdd.n9 vdd.n8 98.6055
R2835 vdd.n11 vdd.n10 98.6055
R2836 vdd.n13 vdd.n12 98.6055
R2837 vdd.n6 vdd.n5 98.6055
R2838 vdd.n4 vdd.n3 98.6055
R2839 vdd.n2 vdd.n1 98.6055
R2840 vdd.t245 vdd.n291 85.8723
R2841 vdd.t223 vdd.n236 85.8723
R2842 vdd.t235 vdd.n193 85.8723
R2843 vdd.t210 vdd.n138 85.8723
R2844 vdd.t197 vdd.n96 85.8723
R2845 vdd.t178 vdd.n41 85.8723
R2846 vdd.t256 vdd.n2022 85.8723
R2847 vdd.t166 vdd.n2077 85.8723
R2848 vdd.t246 vdd.n1924 85.8723
R2849 vdd.t145 vdd.n1979 85.8723
R2850 vdd.t180 vdd.n1827 85.8723
R2851 vdd.t198 vdd.n1882 85.8723
R2852 vdd.n2920 vdd.n843 78.546
R2853 vdd.n2375 vdd.n1014 78.546
R2854 vdd.n278 vdd.n277 75.1835
R2855 vdd.n276 vdd.n275 75.1835
R2856 vdd.n274 vdd.n273 75.1835
R2857 vdd.n272 vdd.n271 75.1835
R2858 vdd.n270 vdd.n269 75.1835
R2859 vdd.n268 vdd.n267 75.1835
R2860 vdd.n266 vdd.n265 75.1835
R2861 vdd.n180 vdd.n179 75.1835
R2862 vdd.n178 vdd.n177 75.1835
R2863 vdd.n176 vdd.n175 75.1835
R2864 vdd.n174 vdd.n173 75.1835
R2865 vdd.n172 vdd.n171 75.1835
R2866 vdd.n170 vdd.n169 75.1835
R2867 vdd.n168 vdd.n167 75.1835
R2868 vdd.n83 vdd.n82 75.1835
R2869 vdd.n81 vdd.n80 75.1835
R2870 vdd.n79 vdd.n78 75.1835
R2871 vdd.n77 vdd.n76 75.1835
R2872 vdd.n75 vdd.n74 75.1835
R2873 vdd.n73 vdd.n72 75.1835
R2874 vdd.n71 vdd.n70 75.1835
R2875 vdd.n2052 vdd.n2051 75.1835
R2876 vdd.n2054 vdd.n2053 75.1835
R2877 vdd.n2056 vdd.n2055 75.1835
R2878 vdd.n2058 vdd.n2057 75.1835
R2879 vdd.n2060 vdd.n2059 75.1835
R2880 vdd.n2062 vdd.n2061 75.1835
R2881 vdd.n2064 vdd.n2063 75.1835
R2882 vdd.n1954 vdd.n1953 75.1835
R2883 vdd.n1956 vdd.n1955 75.1835
R2884 vdd.n1958 vdd.n1957 75.1835
R2885 vdd.n1960 vdd.n1959 75.1835
R2886 vdd.n1962 vdd.n1961 75.1835
R2887 vdd.n1964 vdd.n1963 75.1835
R2888 vdd.n1966 vdd.n1965 75.1835
R2889 vdd.n1857 vdd.n1856 75.1835
R2890 vdd.n1859 vdd.n1858 75.1835
R2891 vdd.n1861 vdd.n1860 75.1835
R2892 vdd.n1863 vdd.n1862 75.1835
R2893 vdd.n1865 vdd.n1864 75.1835
R2894 vdd.n1867 vdd.n1866 75.1835
R2895 vdd.n1869 vdd.n1868 75.1835
R2896 vdd.n2856 vdd.n2855 72.8958
R2897 vdd.n2855 vdd.n2599 72.8958
R2898 vdd.n2855 vdd.n2600 72.8958
R2899 vdd.n2855 vdd.n2601 72.8958
R2900 vdd.n2855 vdd.n2602 72.8958
R2901 vdd.n2855 vdd.n2603 72.8958
R2902 vdd.n2855 vdd.n2604 72.8958
R2903 vdd.n2855 vdd.n2605 72.8958
R2904 vdd.n2855 vdd.n2606 72.8958
R2905 vdd.n2855 vdd.n2607 72.8958
R2906 vdd.n2855 vdd.n2608 72.8958
R2907 vdd.n2855 vdd.n2609 72.8958
R2908 vdd.n2855 vdd.n2610 72.8958
R2909 vdd.n2855 vdd.n2611 72.8958
R2910 vdd.n2855 vdd.n2612 72.8958
R2911 vdd.n2855 vdd.n2613 72.8958
R2912 vdd.n2855 vdd.n2614 72.8958
R2913 vdd.n772 vdd.n756 72.8958
R2914 vdd.n3075 vdd.n756 72.8958
R2915 vdd.n766 vdd.n756 72.8958
R2916 vdd.n3082 vdd.n756 72.8958
R2917 vdd.n763 vdd.n756 72.8958
R2918 vdd.n3089 vdd.n756 72.8958
R2919 vdd.n760 vdd.n756 72.8958
R2920 vdd.n3096 vdd.n756 72.8958
R2921 vdd.n3099 vdd.n756 72.8958
R2922 vdd.n2955 vdd.n756 72.8958
R2923 vdd.n2960 vdd.n756 72.8958
R2924 vdd.n2954 vdd.n756 72.8958
R2925 vdd.n2967 vdd.n756 72.8958
R2926 vdd.n2951 vdd.n756 72.8958
R2927 vdd.n2974 vdd.n756 72.8958
R2928 vdd.n2948 vdd.n756 72.8958
R2929 vdd.n2981 vdd.n756 72.8958
R2930 vdd.n2334 vdd.n2333 72.8958
R2931 vdd.n2334 vdd.n1055 72.8958
R2932 vdd.n2334 vdd.n1056 72.8958
R2933 vdd.n2334 vdd.n1057 72.8958
R2934 vdd.n2334 vdd.n1058 72.8958
R2935 vdd.n2334 vdd.n1059 72.8958
R2936 vdd.n2334 vdd.n1060 72.8958
R2937 vdd.n2334 vdd.n1061 72.8958
R2938 vdd.n2334 vdd.n1062 72.8958
R2939 vdd.n2334 vdd.n1063 72.8958
R2940 vdd.n2334 vdd.n1064 72.8958
R2941 vdd.n2334 vdd.n1065 72.8958
R2942 vdd.n2334 vdd.n1066 72.8958
R2943 vdd.n2334 vdd.n1067 72.8958
R2944 vdd.n2334 vdd.n1068 72.8958
R2945 vdd.n2334 vdd.n1069 72.8958
R2946 vdd.n2334 vdd.n1070 72.8958
R2947 vdd.n2582 vdd.n923 72.8958
R2948 vdd.n2582 vdd.n924 72.8958
R2949 vdd.n2582 vdd.n925 72.8958
R2950 vdd.n2582 vdd.n926 72.8958
R2951 vdd.n2582 vdd.n927 72.8958
R2952 vdd.n2582 vdd.n928 72.8958
R2953 vdd.n2582 vdd.n929 72.8958
R2954 vdd.n2582 vdd.n930 72.8958
R2955 vdd.n2582 vdd.n931 72.8958
R2956 vdd.n2582 vdd.n932 72.8958
R2957 vdd.n2582 vdd.n933 72.8958
R2958 vdd.n2582 vdd.n934 72.8958
R2959 vdd.n2582 vdd.n935 72.8958
R2960 vdd.n2582 vdd.n936 72.8958
R2961 vdd.n2582 vdd.n937 72.8958
R2962 vdd.n2582 vdd.n938 72.8958
R2963 vdd.n2582 vdd.n939 72.8958
R2964 vdd.n2855 vdd.n2854 72.8958
R2965 vdd.n2855 vdd.n2583 72.8958
R2966 vdd.n2855 vdd.n2584 72.8958
R2967 vdd.n2855 vdd.n2585 72.8958
R2968 vdd.n2855 vdd.n2586 72.8958
R2969 vdd.n2855 vdd.n2587 72.8958
R2970 vdd.n2855 vdd.n2588 72.8958
R2971 vdd.n2855 vdd.n2589 72.8958
R2972 vdd.n2855 vdd.n2590 72.8958
R2973 vdd.n2855 vdd.n2591 72.8958
R2974 vdd.n2855 vdd.n2592 72.8958
R2975 vdd.n2855 vdd.n2593 72.8958
R2976 vdd.n2855 vdd.n2594 72.8958
R2977 vdd.n2855 vdd.n2595 72.8958
R2978 vdd.n2855 vdd.n2596 72.8958
R2979 vdd.n2855 vdd.n2597 72.8958
R2980 vdd.n2855 vdd.n2598 72.8958
R2981 vdd.n3003 vdd.n756 72.8958
R2982 vdd.n3009 vdd.n756 72.8958
R2983 vdd.n802 vdd.n756 72.8958
R2984 vdd.n3016 vdd.n756 72.8958
R2985 vdd.n799 vdd.n756 72.8958
R2986 vdd.n3023 vdd.n756 72.8958
R2987 vdd.n796 vdd.n756 72.8958
R2988 vdd.n3030 vdd.n756 72.8958
R2989 vdd.n793 vdd.n756 72.8958
R2990 vdd.n3038 vdd.n756 72.8958
R2991 vdd.n790 vdd.n756 72.8958
R2992 vdd.n3045 vdd.n756 72.8958
R2993 vdd.n787 vdd.n756 72.8958
R2994 vdd.n3052 vdd.n756 72.8958
R2995 vdd.n784 vdd.n756 72.8958
R2996 vdd.n3059 vdd.n756 72.8958
R2997 vdd.n3062 vdd.n756 72.8958
R2998 vdd.n2582 vdd.n921 72.8958
R2999 vdd.n2582 vdd.n920 72.8958
R3000 vdd.n2582 vdd.n919 72.8958
R3001 vdd.n2582 vdd.n918 72.8958
R3002 vdd.n2582 vdd.n917 72.8958
R3003 vdd.n2582 vdd.n916 72.8958
R3004 vdd.n2582 vdd.n915 72.8958
R3005 vdd.n2582 vdd.n914 72.8958
R3006 vdd.n2582 vdd.n913 72.8958
R3007 vdd.n2582 vdd.n912 72.8958
R3008 vdd.n2582 vdd.n911 72.8958
R3009 vdd.n2582 vdd.n910 72.8958
R3010 vdd.n2582 vdd.n909 72.8958
R3011 vdd.n2582 vdd.n908 72.8958
R3012 vdd.n2582 vdd.n907 72.8958
R3013 vdd.n2582 vdd.n906 72.8958
R3014 vdd.n2582 vdd.n905 72.8958
R3015 vdd.n2335 vdd.n2334 72.8958
R3016 vdd.n2334 vdd.n1071 72.8958
R3017 vdd.n2334 vdd.n1072 72.8958
R3018 vdd.n2334 vdd.n1073 72.8958
R3019 vdd.n2334 vdd.n1074 72.8958
R3020 vdd.n2334 vdd.n1075 72.8958
R3021 vdd.n2334 vdd.n1076 72.8958
R3022 vdd.n2334 vdd.n1077 72.8958
R3023 vdd.n2334 vdd.n1078 72.8958
R3024 vdd.n2334 vdd.n1079 72.8958
R3025 vdd.n2334 vdd.n1080 72.8958
R3026 vdd.n2334 vdd.n1081 72.8958
R3027 vdd.n2334 vdd.n1082 72.8958
R3028 vdd.n2334 vdd.n1083 72.8958
R3029 vdd.n2334 vdd.n1084 72.8958
R3030 vdd.n2334 vdd.n1085 72.8958
R3031 vdd.n2334 vdd.n1086 72.8958
R3032 vdd.n1736 vdd.n1735 66.2847
R3033 vdd.n1736 vdd.n1514 66.2847
R3034 vdd.n1736 vdd.n1515 66.2847
R3035 vdd.n1736 vdd.n1516 66.2847
R3036 vdd.n1736 vdd.n1517 66.2847
R3037 vdd.n1736 vdd.n1518 66.2847
R3038 vdd.n1736 vdd.n1519 66.2847
R3039 vdd.n1736 vdd.n1520 66.2847
R3040 vdd.n1736 vdd.n1521 66.2847
R3041 vdd.n1736 vdd.n1522 66.2847
R3042 vdd.n1736 vdd.n1523 66.2847
R3043 vdd.n1736 vdd.n1524 66.2847
R3044 vdd.n1736 vdd.n1525 66.2847
R3045 vdd.n1736 vdd.n1526 66.2847
R3046 vdd.n1736 vdd.n1527 66.2847
R3047 vdd.n1736 vdd.n1528 66.2847
R3048 vdd.n1736 vdd.n1529 66.2847
R3049 vdd.n1736 vdd.n1530 66.2847
R3050 vdd.n1736 vdd.n1531 66.2847
R3051 vdd.n1736 vdd.n1532 66.2847
R3052 vdd.n1736 vdd.n1533 66.2847
R3053 vdd.n1736 vdd.n1534 66.2847
R3054 vdd.n1736 vdd.n1535 66.2847
R3055 vdd.n1736 vdd.n1536 66.2847
R3056 vdd.n1736 vdd.n1537 66.2847
R3057 vdd.n1736 vdd.n1538 66.2847
R3058 vdd.n1736 vdd.n1539 66.2847
R3059 vdd.n1736 vdd.n1540 66.2847
R3060 vdd.n1736 vdd.n1541 66.2847
R3061 vdd.n1736 vdd.n1542 66.2847
R3062 vdd.n1736 vdd.n1543 66.2847
R3063 vdd.n1404 vdd.n1054 66.2847
R3064 vdd.n1401 vdd.n1054 66.2847
R3065 vdd.n1397 vdd.n1054 66.2847
R3066 vdd.n2196 vdd.n1054 66.2847
R3067 vdd.n1188 vdd.n1054 66.2847
R3068 vdd.n2203 vdd.n1054 66.2847
R3069 vdd.n1181 vdd.n1054 66.2847
R3070 vdd.n2210 vdd.n1054 66.2847
R3071 vdd.n1174 vdd.n1054 66.2847
R3072 vdd.n2217 vdd.n1054 66.2847
R3073 vdd.n1168 vdd.n1054 66.2847
R3074 vdd.n1163 vdd.n1054 66.2847
R3075 vdd.n2228 vdd.n1054 66.2847
R3076 vdd.n1155 vdd.n1054 66.2847
R3077 vdd.n2235 vdd.n1054 66.2847
R3078 vdd.n1148 vdd.n1054 66.2847
R3079 vdd.n2242 vdd.n1054 66.2847
R3080 vdd.n1141 vdd.n1054 66.2847
R3081 vdd.n2249 vdd.n1054 66.2847
R3082 vdd.n1134 vdd.n1054 66.2847
R3083 vdd.n2256 vdd.n1054 66.2847
R3084 vdd.n1128 vdd.n1054 66.2847
R3085 vdd.n1123 vdd.n1054 66.2847
R3086 vdd.n2267 vdd.n1054 66.2847
R3087 vdd.n1115 vdd.n1054 66.2847
R3088 vdd.n2274 vdd.n1054 66.2847
R3089 vdd.n1108 vdd.n1054 66.2847
R3090 vdd.n2281 vdd.n1054 66.2847
R3091 vdd.n1101 vdd.n1054 66.2847
R3092 vdd.n2288 vdd.n1054 66.2847
R3093 vdd.n2293 vdd.n1054 66.2847
R3094 vdd.n1097 vdd.n1054 66.2847
R3095 vdd.n3229 vdd.n658 66.2847
R3096 vdd.n663 vdd.n658 66.2847
R3097 vdd.n666 vdd.n658 66.2847
R3098 vdd.n3218 vdd.n658 66.2847
R3099 vdd.n3212 vdd.n658 66.2847
R3100 vdd.n3210 vdd.n658 66.2847
R3101 vdd.n3204 vdd.n658 66.2847
R3102 vdd.n3202 vdd.n658 66.2847
R3103 vdd.n3196 vdd.n658 66.2847
R3104 vdd.n3194 vdd.n658 66.2847
R3105 vdd.n3188 vdd.n658 66.2847
R3106 vdd.n3186 vdd.n658 66.2847
R3107 vdd.n3180 vdd.n658 66.2847
R3108 vdd.n3178 vdd.n658 66.2847
R3109 vdd.n3172 vdd.n658 66.2847
R3110 vdd.n3170 vdd.n658 66.2847
R3111 vdd.n3164 vdd.n658 66.2847
R3112 vdd.n3162 vdd.n658 66.2847
R3113 vdd.n3156 vdd.n658 66.2847
R3114 vdd.n3154 vdd.n658 66.2847
R3115 vdd.n727 vdd.n658 66.2847
R3116 vdd.n3145 vdd.n658 66.2847
R3117 vdd.n729 vdd.n658 66.2847
R3118 vdd.n3138 vdd.n658 66.2847
R3119 vdd.n3132 vdd.n658 66.2847
R3120 vdd.n3130 vdd.n658 66.2847
R3121 vdd.n3124 vdd.n658 66.2847
R3122 vdd.n3122 vdd.n658 66.2847
R3123 vdd.n3116 vdd.n658 66.2847
R3124 vdd.n750 vdd.n658 66.2847
R3125 vdd.n752 vdd.n658 66.2847
R3126 vdd.n3345 vdd.n3344 66.2847
R3127 vdd.n3345 vdd.n403 66.2847
R3128 vdd.n3345 vdd.n402 66.2847
R3129 vdd.n3345 vdd.n401 66.2847
R3130 vdd.n3345 vdd.n400 66.2847
R3131 vdd.n3345 vdd.n399 66.2847
R3132 vdd.n3345 vdd.n398 66.2847
R3133 vdd.n3345 vdd.n397 66.2847
R3134 vdd.n3345 vdd.n396 66.2847
R3135 vdd.n3345 vdd.n395 66.2847
R3136 vdd.n3345 vdd.n394 66.2847
R3137 vdd.n3345 vdd.n393 66.2847
R3138 vdd.n3345 vdd.n392 66.2847
R3139 vdd.n3345 vdd.n391 66.2847
R3140 vdd.n3345 vdd.n390 66.2847
R3141 vdd.n3345 vdd.n389 66.2847
R3142 vdd.n3345 vdd.n388 66.2847
R3143 vdd.n3345 vdd.n387 66.2847
R3144 vdd.n3345 vdd.n386 66.2847
R3145 vdd.n3345 vdd.n385 66.2847
R3146 vdd.n3345 vdd.n384 66.2847
R3147 vdd.n3345 vdd.n383 66.2847
R3148 vdd.n3345 vdd.n382 66.2847
R3149 vdd.n3345 vdd.n381 66.2847
R3150 vdd.n3345 vdd.n380 66.2847
R3151 vdd.n3345 vdd.n379 66.2847
R3152 vdd.n3345 vdd.n378 66.2847
R3153 vdd.n3345 vdd.n377 66.2847
R3154 vdd.n3345 vdd.n376 66.2847
R3155 vdd.n3345 vdd.n375 66.2847
R3156 vdd.n3345 vdd.n374 66.2847
R3157 vdd.n3345 vdd.n373 66.2847
R3158 vdd.n448 vdd.n373 52.4337
R3159 vdd.n454 vdd.n374 52.4337
R3160 vdd.n458 vdd.n375 52.4337
R3161 vdd.n464 vdd.n376 52.4337
R3162 vdd.n468 vdd.n377 52.4337
R3163 vdd.n474 vdd.n378 52.4337
R3164 vdd.n478 vdd.n379 52.4337
R3165 vdd.n484 vdd.n380 52.4337
R3166 vdd.n488 vdd.n381 52.4337
R3167 vdd.n494 vdd.n382 52.4337
R3168 vdd.n498 vdd.n383 52.4337
R3169 vdd.n504 vdd.n384 52.4337
R3170 vdd.n508 vdd.n385 52.4337
R3171 vdd.n514 vdd.n386 52.4337
R3172 vdd.n518 vdd.n387 52.4337
R3173 vdd.n524 vdd.n388 52.4337
R3174 vdd.n528 vdd.n389 52.4337
R3175 vdd.n534 vdd.n390 52.4337
R3176 vdd.n538 vdd.n391 52.4337
R3177 vdd.n544 vdd.n392 52.4337
R3178 vdd.n548 vdd.n393 52.4337
R3179 vdd.n554 vdd.n394 52.4337
R3180 vdd.n558 vdd.n395 52.4337
R3181 vdd.n564 vdd.n396 52.4337
R3182 vdd.n568 vdd.n397 52.4337
R3183 vdd.n574 vdd.n398 52.4337
R3184 vdd.n578 vdd.n399 52.4337
R3185 vdd.n584 vdd.n400 52.4337
R3186 vdd.n588 vdd.n401 52.4337
R3187 vdd.n594 vdd.n402 52.4337
R3188 vdd.n597 vdd.n403 52.4337
R3189 vdd.n3344 vdd.n3343 52.4337
R3190 vdd.n3229 vdd.n660 52.4337
R3191 vdd.n3227 vdd.n663 52.4337
R3192 vdd.n3223 vdd.n666 52.4337
R3193 vdd.n3219 vdd.n3218 52.4337
R3194 vdd.n3212 vdd.n669 52.4337
R3195 vdd.n3211 vdd.n3210 52.4337
R3196 vdd.n3204 vdd.n675 52.4337
R3197 vdd.n3203 vdd.n3202 52.4337
R3198 vdd.n3196 vdd.n681 52.4337
R3199 vdd.n3195 vdd.n3194 52.4337
R3200 vdd.n3188 vdd.n689 52.4337
R3201 vdd.n3187 vdd.n3186 52.4337
R3202 vdd.n3180 vdd.n695 52.4337
R3203 vdd.n3179 vdd.n3178 52.4337
R3204 vdd.n3172 vdd.n701 52.4337
R3205 vdd.n3171 vdd.n3170 52.4337
R3206 vdd.n3164 vdd.n707 52.4337
R3207 vdd.n3163 vdd.n3162 52.4337
R3208 vdd.n3156 vdd.n713 52.4337
R3209 vdd.n3155 vdd.n3154 52.4337
R3210 vdd.n727 vdd.n719 52.4337
R3211 vdd.n3146 vdd.n3145 52.4337
R3212 vdd.n3143 vdd.n729 52.4337
R3213 vdd.n3139 vdd.n3138 52.4337
R3214 vdd.n3132 vdd.n733 52.4337
R3215 vdd.n3131 vdd.n3130 52.4337
R3216 vdd.n3124 vdd.n739 52.4337
R3217 vdd.n3123 vdd.n3122 52.4337
R3218 vdd.n3116 vdd.n745 52.4337
R3219 vdd.n3115 vdd.n750 52.4337
R3220 vdd.n3111 vdd.n752 52.4337
R3221 vdd.n2295 vdd.n1097 52.4337
R3222 vdd.n2293 vdd.n2292 52.4337
R3223 vdd.n2288 vdd.n2287 52.4337
R3224 vdd.n2283 vdd.n1101 52.4337
R3225 vdd.n2281 vdd.n2280 52.4337
R3226 vdd.n2276 vdd.n1108 52.4337
R3227 vdd.n2274 vdd.n2273 52.4337
R3228 vdd.n2269 vdd.n1115 52.4337
R3229 vdd.n2267 vdd.n2266 52.4337
R3230 vdd.n1124 vdd.n1123 52.4337
R3231 vdd.n2258 vdd.n1128 52.4337
R3232 vdd.n2256 vdd.n2255 52.4337
R3233 vdd.n2251 vdd.n1134 52.4337
R3234 vdd.n2249 vdd.n2248 52.4337
R3235 vdd.n2244 vdd.n1141 52.4337
R3236 vdd.n2242 vdd.n2241 52.4337
R3237 vdd.n2237 vdd.n1148 52.4337
R3238 vdd.n2235 vdd.n2234 52.4337
R3239 vdd.n2230 vdd.n1155 52.4337
R3240 vdd.n2228 vdd.n2227 52.4337
R3241 vdd.n1164 vdd.n1163 52.4337
R3242 vdd.n2219 vdd.n1168 52.4337
R3243 vdd.n2217 vdd.n2216 52.4337
R3244 vdd.n2212 vdd.n1174 52.4337
R3245 vdd.n2210 vdd.n2209 52.4337
R3246 vdd.n2205 vdd.n1181 52.4337
R3247 vdd.n2203 vdd.n2202 52.4337
R3248 vdd.n2198 vdd.n1188 52.4337
R3249 vdd.n2196 vdd.n2195 52.4337
R3250 vdd.n1398 vdd.n1397 52.4337
R3251 vdd.n1402 vdd.n1401 52.4337
R3252 vdd.n2184 vdd.n1404 52.4337
R3253 vdd.n1735 vdd.n1734 52.4337
R3254 vdd.n1549 vdd.n1514 52.4337
R3255 vdd.n1551 vdd.n1515 52.4337
R3256 vdd.n1555 vdd.n1516 52.4337
R3257 vdd.n1557 vdd.n1517 52.4337
R3258 vdd.n1561 vdd.n1518 52.4337
R3259 vdd.n1563 vdd.n1519 52.4337
R3260 vdd.n1567 vdd.n1520 52.4337
R3261 vdd.n1569 vdd.n1521 52.4337
R3262 vdd.n1701 vdd.n1522 52.4337
R3263 vdd.n1573 vdd.n1523 52.4337
R3264 vdd.n1577 vdd.n1524 52.4337
R3265 vdd.n1579 vdd.n1525 52.4337
R3266 vdd.n1583 vdd.n1526 52.4337
R3267 vdd.n1585 vdd.n1527 52.4337
R3268 vdd.n1589 vdd.n1528 52.4337
R3269 vdd.n1591 vdd.n1529 52.4337
R3270 vdd.n1595 vdd.n1530 52.4337
R3271 vdd.n1597 vdd.n1531 52.4337
R3272 vdd.n1601 vdd.n1532 52.4337
R3273 vdd.n1665 vdd.n1533 52.4337
R3274 vdd.n1606 vdd.n1534 52.4337
R3275 vdd.n1608 vdd.n1535 52.4337
R3276 vdd.n1612 vdd.n1536 52.4337
R3277 vdd.n1614 vdd.n1537 52.4337
R3278 vdd.n1618 vdd.n1538 52.4337
R3279 vdd.n1620 vdd.n1539 52.4337
R3280 vdd.n1624 vdd.n1540 52.4337
R3281 vdd.n1626 vdd.n1541 52.4337
R3282 vdd.n1630 vdd.n1542 52.4337
R3283 vdd.n1632 vdd.n1543 52.4337
R3284 vdd.n1735 vdd.n1545 52.4337
R3285 vdd.n1550 vdd.n1514 52.4337
R3286 vdd.n1554 vdd.n1515 52.4337
R3287 vdd.n1556 vdd.n1516 52.4337
R3288 vdd.n1560 vdd.n1517 52.4337
R3289 vdd.n1562 vdd.n1518 52.4337
R3290 vdd.n1566 vdd.n1519 52.4337
R3291 vdd.n1568 vdd.n1520 52.4337
R3292 vdd.n1700 vdd.n1521 52.4337
R3293 vdd.n1572 vdd.n1522 52.4337
R3294 vdd.n1576 vdd.n1523 52.4337
R3295 vdd.n1578 vdd.n1524 52.4337
R3296 vdd.n1582 vdd.n1525 52.4337
R3297 vdd.n1584 vdd.n1526 52.4337
R3298 vdd.n1588 vdd.n1527 52.4337
R3299 vdd.n1590 vdd.n1528 52.4337
R3300 vdd.n1594 vdd.n1529 52.4337
R3301 vdd.n1596 vdd.n1530 52.4337
R3302 vdd.n1600 vdd.n1531 52.4337
R3303 vdd.n1602 vdd.n1532 52.4337
R3304 vdd.n1605 vdd.n1533 52.4337
R3305 vdd.n1607 vdd.n1534 52.4337
R3306 vdd.n1611 vdd.n1535 52.4337
R3307 vdd.n1613 vdd.n1536 52.4337
R3308 vdd.n1617 vdd.n1537 52.4337
R3309 vdd.n1619 vdd.n1538 52.4337
R3310 vdd.n1623 vdd.n1539 52.4337
R3311 vdd.n1625 vdd.n1540 52.4337
R3312 vdd.n1629 vdd.n1541 52.4337
R3313 vdd.n1631 vdd.n1542 52.4337
R3314 vdd.n1543 vdd.n1513 52.4337
R3315 vdd.n1404 vdd.n1403 52.4337
R3316 vdd.n1401 vdd.n1400 52.4337
R3317 vdd.n1397 vdd.n1189 52.4337
R3318 vdd.n2197 vdd.n2196 52.4337
R3319 vdd.n1188 vdd.n1182 52.4337
R3320 vdd.n2204 vdd.n2203 52.4337
R3321 vdd.n1181 vdd.n1175 52.4337
R3322 vdd.n2211 vdd.n2210 52.4337
R3323 vdd.n1174 vdd.n1169 52.4337
R3324 vdd.n2218 vdd.n2217 52.4337
R3325 vdd.n1168 vdd.n1167 52.4337
R3326 vdd.n1163 vdd.n1156 52.4337
R3327 vdd.n2229 vdd.n2228 52.4337
R3328 vdd.n1155 vdd.n1149 52.4337
R3329 vdd.n2236 vdd.n2235 52.4337
R3330 vdd.n1148 vdd.n1142 52.4337
R3331 vdd.n2243 vdd.n2242 52.4337
R3332 vdd.n1141 vdd.n1135 52.4337
R3333 vdd.n2250 vdd.n2249 52.4337
R3334 vdd.n1134 vdd.n1129 52.4337
R3335 vdd.n2257 vdd.n2256 52.4337
R3336 vdd.n1128 vdd.n1127 52.4337
R3337 vdd.n1123 vdd.n1116 52.4337
R3338 vdd.n2268 vdd.n2267 52.4337
R3339 vdd.n1115 vdd.n1109 52.4337
R3340 vdd.n2275 vdd.n2274 52.4337
R3341 vdd.n1108 vdd.n1102 52.4337
R3342 vdd.n2282 vdd.n2281 52.4337
R3343 vdd.n1101 vdd.n1098 52.4337
R3344 vdd.n2289 vdd.n2288 52.4337
R3345 vdd.n2294 vdd.n2293 52.4337
R3346 vdd.n1409 vdd.n1097 52.4337
R3347 vdd.n3230 vdd.n3229 52.4337
R3348 vdd.n3224 vdd.n663 52.4337
R3349 vdd.n3220 vdd.n666 52.4337
R3350 vdd.n3218 vdd.n3217 52.4337
R3351 vdd.n3213 vdd.n3212 52.4337
R3352 vdd.n3210 vdd.n3209 52.4337
R3353 vdd.n3205 vdd.n3204 52.4337
R3354 vdd.n3202 vdd.n3201 52.4337
R3355 vdd.n3197 vdd.n3196 52.4337
R3356 vdd.n3194 vdd.n3193 52.4337
R3357 vdd.n3189 vdd.n3188 52.4337
R3358 vdd.n3186 vdd.n3185 52.4337
R3359 vdd.n3181 vdd.n3180 52.4337
R3360 vdd.n3178 vdd.n3177 52.4337
R3361 vdd.n3173 vdd.n3172 52.4337
R3362 vdd.n3170 vdd.n3169 52.4337
R3363 vdd.n3165 vdd.n3164 52.4337
R3364 vdd.n3162 vdd.n3161 52.4337
R3365 vdd.n3157 vdd.n3156 52.4337
R3366 vdd.n3154 vdd.n3153 52.4337
R3367 vdd.n728 vdd.n727 52.4337
R3368 vdd.n3145 vdd.n3144 52.4337
R3369 vdd.n3140 vdd.n729 52.4337
R3370 vdd.n3138 vdd.n3137 52.4337
R3371 vdd.n3133 vdd.n3132 52.4337
R3372 vdd.n3130 vdd.n3129 52.4337
R3373 vdd.n3125 vdd.n3124 52.4337
R3374 vdd.n3122 vdd.n3121 52.4337
R3375 vdd.n3117 vdd.n3116 52.4337
R3376 vdd.n3112 vdd.n750 52.4337
R3377 vdd.n3108 vdd.n752 52.4337
R3378 vdd.n3344 vdd.n404 52.4337
R3379 vdd.n595 vdd.n403 52.4337
R3380 vdd.n589 vdd.n402 52.4337
R3381 vdd.n585 vdd.n401 52.4337
R3382 vdd.n579 vdd.n400 52.4337
R3383 vdd.n575 vdd.n399 52.4337
R3384 vdd.n569 vdd.n398 52.4337
R3385 vdd.n565 vdd.n397 52.4337
R3386 vdd.n559 vdd.n396 52.4337
R3387 vdd.n555 vdd.n395 52.4337
R3388 vdd.n549 vdd.n394 52.4337
R3389 vdd.n545 vdd.n393 52.4337
R3390 vdd.n539 vdd.n392 52.4337
R3391 vdd.n535 vdd.n391 52.4337
R3392 vdd.n529 vdd.n390 52.4337
R3393 vdd.n525 vdd.n389 52.4337
R3394 vdd.n519 vdd.n388 52.4337
R3395 vdd.n515 vdd.n387 52.4337
R3396 vdd.n509 vdd.n386 52.4337
R3397 vdd.n505 vdd.n385 52.4337
R3398 vdd.n499 vdd.n384 52.4337
R3399 vdd.n495 vdd.n383 52.4337
R3400 vdd.n489 vdd.n382 52.4337
R3401 vdd.n485 vdd.n381 52.4337
R3402 vdd.n479 vdd.n380 52.4337
R3403 vdd.n475 vdd.n379 52.4337
R3404 vdd.n469 vdd.n378 52.4337
R3405 vdd.n465 vdd.n377 52.4337
R3406 vdd.n459 vdd.n376 52.4337
R3407 vdd.n455 vdd.n375 52.4337
R3408 vdd.n449 vdd.n374 52.4337
R3409 vdd.n445 vdd.n373 52.4337
R3410 vdd.t14 vdd.t26 51.4683
R3411 vdd.n266 vdd.n264 42.0461
R3412 vdd.n168 vdd.n166 42.0461
R3413 vdd.n71 vdd.n69 42.0461
R3414 vdd.n2052 vdd.n2050 42.0461
R3415 vdd.n1954 vdd.n1952 42.0461
R3416 vdd.n1857 vdd.n1855 42.0461
R3417 vdd.n320 vdd.n319 41.6884
R3418 vdd.n222 vdd.n221 41.6884
R3419 vdd.n125 vdd.n124 41.6884
R3420 vdd.n2106 vdd.n2105 41.6884
R3421 vdd.n2008 vdd.n2007 41.6884
R3422 vdd.n1911 vdd.n1910 41.6884
R3423 vdd.n1512 vdd.n1511 41.1157
R3424 vdd.n1668 vdd.n1667 41.1157
R3425 vdd.n1704 vdd.n1703 41.1157
R3426 vdd.n407 vdd.n406 41.1157
R3427 vdd.n547 vdd.n420 41.1157
R3428 vdd.n433 vdd.n432 41.1157
R3429 vdd.n3062 vdd.n3061 39.2114
R3430 vdd.n3059 vdd.n3058 39.2114
R3431 vdd.n3054 vdd.n784 39.2114
R3432 vdd.n3052 vdd.n3051 39.2114
R3433 vdd.n3047 vdd.n787 39.2114
R3434 vdd.n3045 vdd.n3044 39.2114
R3435 vdd.n3040 vdd.n790 39.2114
R3436 vdd.n3038 vdd.n3037 39.2114
R3437 vdd.n3032 vdd.n793 39.2114
R3438 vdd.n3030 vdd.n3029 39.2114
R3439 vdd.n3025 vdd.n796 39.2114
R3440 vdd.n3023 vdd.n3022 39.2114
R3441 vdd.n3018 vdd.n799 39.2114
R3442 vdd.n3016 vdd.n3015 39.2114
R3443 vdd.n3011 vdd.n802 39.2114
R3444 vdd.n3009 vdd.n3008 39.2114
R3445 vdd.n3004 vdd.n3003 39.2114
R3446 vdd.n2854 vdd.n2853 39.2114
R3447 vdd.n2848 vdd.n2583 39.2114
R3448 vdd.n2845 vdd.n2584 39.2114
R3449 vdd.n2841 vdd.n2585 39.2114
R3450 vdd.n2837 vdd.n2586 39.2114
R3451 vdd.n2833 vdd.n2587 39.2114
R3452 vdd.n2829 vdd.n2588 39.2114
R3453 vdd.n2825 vdd.n2589 39.2114
R3454 vdd.n2821 vdd.n2590 39.2114
R3455 vdd.n2817 vdd.n2591 39.2114
R3456 vdd.n2813 vdd.n2592 39.2114
R3457 vdd.n2809 vdd.n2593 39.2114
R3458 vdd.n2805 vdd.n2594 39.2114
R3459 vdd.n2801 vdd.n2595 39.2114
R3460 vdd.n2797 vdd.n2596 39.2114
R3461 vdd.n2793 vdd.n2597 39.2114
R3462 vdd.n2788 vdd.n2598 39.2114
R3463 vdd.n2577 vdd.n939 39.2114
R3464 vdd.n2573 vdd.n938 39.2114
R3465 vdd.n2569 vdd.n937 39.2114
R3466 vdd.n2565 vdd.n936 39.2114
R3467 vdd.n2561 vdd.n935 39.2114
R3468 vdd.n2557 vdd.n934 39.2114
R3469 vdd.n2553 vdd.n933 39.2114
R3470 vdd.n2549 vdd.n932 39.2114
R3471 vdd.n2545 vdd.n931 39.2114
R3472 vdd.n2541 vdd.n930 39.2114
R3473 vdd.n2537 vdd.n929 39.2114
R3474 vdd.n2533 vdd.n928 39.2114
R3475 vdd.n2529 vdd.n927 39.2114
R3476 vdd.n2525 vdd.n926 39.2114
R3477 vdd.n2521 vdd.n925 39.2114
R3478 vdd.n2516 vdd.n924 39.2114
R3479 vdd.n2512 vdd.n923 39.2114
R3480 vdd.n2333 vdd.n2332 39.2114
R3481 vdd.n2327 vdd.n1055 39.2114
R3482 vdd.n2324 vdd.n1056 39.2114
R3483 vdd.n2320 vdd.n1057 39.2114
R3484 vdd.n2316 vdd.n1058 39.2114
R3485 vdd.n2312 vdd.n1059 39.2114
R3486 vdd.n2308 vdd.n1060 39.2114
R3487 vdd.n2304 vdd.n1061 39.2114
R3488 vdd.n2300 vdd.n1062 39.2114
R3489 vdd.n1247 vdd.n1063 39.2114
R3490 vdd.n1251 vdd.n1064 39.2114
R3491 vdd.n1255 vdd.n1065 39.2114
R3492 vdd.n1259 vdd.n1066 39.2114
R3493 vdd.n1263 vdd.n1067 39.2114
R3494 vdd.n1267 vdd.n1068 39.2114
R3495 vdd.n1271 vdd.n1069 39.2114
R3496 vdd.n1276 vdd.n1070 39.2114
R3497 vdd.n2981 vdd.n2980 39.2114
R3498 vdd.n2976 vdd.n2948 39.2114
R3499 vdd.n2974 vdd.n2973 39.2114
R3500 vdd.n2969 vdd.n2951 39.2114
R3501 vdd.n2967 vdd.n2966 39.2114
R3502 vdd.n2962 vdd.n2954 39.2114
R3503 vdd.n2960 vdd.n2959 39.2114
R3504 vdd.n2955 vdd.n755 39.2114
R3505 vdd.n3099 vdd.n3098 39.2114
R3506 vdd.n3096 vdd.n3095 39.2114
R3507 vdd.n3091 vdd.n760 39.2114
R3508 vdd.n3089 vdd.n3088 39.2114
R3509 vdd.n3084 vdd.n763 39.2114
R3510 vdd.n3082 vdd.n3081 39.2114
R3511 vdd.n3077 vdd.n766 39.2114
R3512 vdd.n3075 vdd.n3074 39.2114
R3513 vdd.n3070 vdd.n772 39.2114
R3514 vdd.n2857 vdd.n2856 39.2114
R3515 vdd.n2624 vdd.n2599 39.2114
R3516 vdd.n2628 vdd.n2600 39.2114
R3517 vdd.n2632 vdd.n2601 39.2114
R3518 vdd.n2636 vdd.n2602 39.2114
R3519 vdd.n2640 vdd.n2603 39.2114
R3520 vdd.n2644 vdd.n2604 39.2114
R3521 vdd.n2648 vdd.n2605 39.2114
R3522 vdd.n2652 vdd.n2606 39.2114
R3523 vdd.n2656 vdd.n2607 39.2114
R3524 vdd.n2660 vdd.n2608 39.2114
R3525 vdd.n2664 vdd.n2609 39.2114
R3526 vdd.n2668 vdd.n2610 39.2114
R3527 vdd.n2672 vdd.n2611 39.2114
R3528 vdd.n2676 vdd.n2612 39.2114
R3529 vdd.n2680 vdd.n2613 39.2114
R3530 vdd.n2684 vdd.n2614 39.2114
R3531 vdd.n2856 vdd.n904 39.2114
R3532 vdd.n2627 vdd.n2599 39.2114
R3533 vdd.n2631 vdd.n2600 39.2114
R3534 vdd.n2635 vdd.n2601 39.2114
R3535 vdd.n2639 vdd.n2602 39.2114
R3536 vdd.n2643 vdd.n2603 39.2114
R3537 vdd.n2647 vdd.n2604 39.2114
R3538 vdd.n2651 vdd.n2605 39.2114
R3539 vdd.n2655 vdd.n2606 39.2114
R3540 vdd.n2659 vdd.n2607 39.2114
R3541 vdd.n2663 vdd.n2608 39.2114
R3542 vdd.n2667 vdd.n2609 39.2114
R3543 vdd.n2671 vdd.n2610 39.2114
R3544 vdd.n2675 vdd.n2611 39.2114
R3545 vdd.n2679 vdd.n2612 39.2114
R3546 vdd.n2683 vdd.n2613 39.2114
R3547 vdd.n2686 vdd.n2614 39.2114
R3548 vdd.n772 vdd.n767 39.2114
R3549 vdd.n3076 vdd.n3075 39.2114
R3550 vdd.n766 vdd.n764 39.2114
R3551 vdd.n3083 vdd.n3082 39.2114
R3552 vdd.n763 vdd.n761 39.2114
R3553 vdd.n3090 vdd.n3089 39.2114
R3554 vdd.n760 vdd.n758 39.2114
R3555 vdd.n3097 vdd.n3096 39.2114
R3556 vdd.n3100 vdd.n3099 39.2114
R3557 vdd.n2956 vdd.n2955 39.2114
R3558 vdd.n2961 vdd.n2960 39.2114
R3559 vdd.n2954 vdd.n2952 39.2114
R3560 vdd.n2968 vdd.n2967 39.2114
R3561 vdd.n2951 vdd.n2949 39.2114
R3562 vdd.n2975 vdd.n2974 39.2114
R3563 vdd.n2948 vdd.n2946 39.2114
R3564 vdd.n2982 vdd.n2981 39.2114
R3565 vdd.n2333 vdd.n1089 39.2114
R3566 vdd.n2325 vdd.n1055 39.2114
R3567 vdd.n2321 vdd.n1056 39.2114
R3568 vdd.n2317 vdd.n1057 39.2114
R3569 vdd.n2313 vdd.n1058 39.2114
R3570 vdd.n2309 vdd.n1059 39.2114
R3571 vdd.n2305 vdd.n1060 39.2114
R3572 vdd.n2301 vdd.n1061 39.2114
R3573 vdd.n1246 vdd.n1062 39.2114
R3574 vdd.n1250 vdd.n1063 39.2114
R3575 vdd.n1254 vdd.n1064 39.2114
R3576 vdd.n1258 vdd.n1065 39.2114
R3577 vdd.n1262 vdd.n1066 39.2114
R3578 vdd.n1266 vdd.n1067 39.2114
R3579 vdd.n1270 vdd.n1068 39.2114
R3580 vdd.n1275 vdd.n1069 39.2114
R3581 vdd.n1279 vdd.n1070 39.2114
R3582 vdd.n2515 vdd.n923 39.2114
R3583 vdd.n2520 vdd.n924 39.2114
R3584 vdd.n2524 vdd.n925 39.2114
R3585 vdd.n2528 vdd.n926 39.2114
R3586 vdd.n2532 vdd.n927 39.2114
R3587 vdd.n2536 vdd.n928 39.2114
R3588 vdd.n2540 vdd.n929 39.2114
R3589 vdd.n2544 vdd.n930 39.2114
R3590 vdd.n2548 vdd.n931 39.2114
R3591 vdd.n2552 vdd.n932 39.2114
R3592 vdd.n2556 vdd.n933 39.2114
R3593 vdd.n2560 vdd.n934 39.2114
R3594 vdd.n2564 vdd.n935 39.2114
R3595 vdd.n2568 vdd.n936 39.2114
R3596 vdd.n2572 vdd.n937 39.2114
R3597 vdd.n2576 vdd.n938 39.2114
R3598 vdd.n941 vdd.n939 39.2114
R3599 vdd.n2854 vdd.n2617 39.2114
R3600 vdd.n2846 vdd.n2583 39.2114
R3601 vdd.n2842 vdd.n2584 39.2114
R3602 vdd.n2838 vdd.n2585 39.2114
R3603 vdd.n2834 vdd.n2586 39.2114
R3604 vdd.n2830 vdd.n2587 39.2114
R3605 vdd.n2826 vdd.n2588 39.2114
R3606 vdd.n2822 vdd.n2589 39.2114
R3607 vdd.n2818 vdd.n2590 39.2114
R3608 vdd.n2814 vdd.n2591 39.2114
R3609 vdd.n2810 vdd.n2592 39.2114
R3610 vdd.n2806 vdd.n2593 39.2114
R3611 vdd.n2802 vdd.n2594 39.2114
R3612 vdd.n2798 vdd.n2595 39.2114
R3613 vdd.n2794 vdd.n2596 39.2114
R3614 vdd.n2789 vdd.n2597 39.2114
R3615 vdd.n2785 vdd.n2598 39.2114
R3616 vdd.n3003 vdd.n803 39.2114
R3617 vdd.n3010 vdd.n3009 39.2114
R3618 vdd.n802 vdd.n800 39.2114
R3619 vdd.n3017 vdd.n3016 39.2114
R3620 vdd.n799 vdd.n797 39.2114
R3621 vdd.n3024 vdd.n3023 39.2114
R3622 vdd.n796 vdd.n794 39.2114
R3623 vdd.n3031 vdd.n3030 39.2114
R3624 vdd.n793 vdd.n791 39.2114
R3625 vdd.n3039 vdd.n3038 39.2114
R3626 vdd.n790 vdd.n788 39.2114
R3627 vdd.n3046 vdd.n3045 39.2114
R3628 vdd.n787 vdd.n785 39.2114
R3629 vdd.n3053 vdd.n3052 39.2114
R3630 vdd.n784 vdd.n782 39.2114
R3631 vdd.n3060 vdd.n3059 39.2114
R3632 vdd.n3063 vdd.n3062 39.2114
R3633 vdd.n950 vdd.n905 39.2114
R3634 vdd.n2504 vdd.n906 39.2114
R3635 vdd.n2500 vdd.n907 39.2114
R3636 vdd.n2496 vdd.n908 39.2114
R3637 vdd.n2492 vdd.n909 39.2114
R3638 vdd.n2488 vdd.n910 39.2114
R3639 vdd.n2484 vdd.n911 39.2114
R3640 vdd.n2480 vdd.n912 39.2114
R3641 vdd.n2476 vdd.n913 39.2114
R3642 vdd.n2472 vdd.n914 39.2114
R3643 vdd.n2468 vdd.n915 39.2114
R3644 vdd.n2464 vdd.n916 39.2114
R3645 vdd.n2460 vdd.n917 39.2114
R3646 vdd.n2456 vdd.n918 39.2114
R3647 vdd.n2452 vdd.n919 39.2114
R3648 vdd.n2448 vdd.n920 39.2114
R3649 vdd.n2444 vdd.n921 39.2114
R3650 vdd.n2336 vdd.n2335 39.2114
R3651 vdd.n1193 vdd.n1071 39.2114
R3652 vdd.n1197 vdd.n1072 39.2114
R3653 vdd.n1201 vdd.n1073 39.2114
R3654 vdd.n1205 vdd.n1074 39.2114
R3655 vdd.n1209 vdd.n1075 39.2114
R3656 vdd.n1213 vdd.n1076 39.2114
R3657 vdd.n1217 vdd.n1077 39.2114
R3658 vdd.n1221 vdd.n1078 39.2114
R3659 vdd.n1391 vdd.n1079 39.2114
R3660 vdd.n1388 vdd.n1080 39.2114
R3661 vdd.n1384 vdd.n1081 39.2114
R3662 vdd.n1380 vdd.n1082 39.2114
R3663 vdd.n1376 vdd.n1083 39.2114
R3664 vdd.n1372 vdd.n1084 39.2114
R3665 vdd.n1368 vdd.n1085 39.2114
R3666 vdd.n1364 vdd.n1086 39.2114
R3667 vdd.n2441 vdd.n921 39.2114
R3668 vdd.n2445 vdd.n920 39.2114
R3669 vdd.n2449 vdd.n919 39.2114
R3670 vdd.n2453 vdd.n918 39.2114
R3671 vdd.n2457 vdd.n917 39.2114
R3672 vdd.n2461 vdd.n916 39.2114
R3673 vdd.n2465 vdd.n915 39.2114
R3674 vdd.n2469 vdd.n914 39.2114
R3675 vdd.n2473 vdd.n913 39.2114
R3676 vdd.n2477 vdd.n912 39.2114
R3677 vdd.n2481 vdd.n911 39.2114
R3678 vdd.n2485 vdd.n910 39.2114
R3679 vdd.n2489 vdd.n909 39.2114
R3680 vdd.n2493 vdd.n908 39.2114
R3681 vdd.n2497 vdd.n907 39.2114
R3682 vdd.n2501 vdd.n906 39.2114
R3683 vdd.n2505 vdd.n905 39.2114
R3684 vdd.n2335 vdd.n1053 39.2114
R3685 vdd.n1196 vdd.n1071 39.2114
R3686 vdd.n1200 vdd.n1072 39.2114
R3687 vdd.n1204 vdd.n1073 39.2114
R3688 vdd.n1208 vdd.n1074 39.2114
R3689 vdd.n1212 vdd.n1075 39.2114
R3690 vdd.n1216 vdd.n1076 39.2114
R3691 vdd.n1220 vdd.n1077 39.2114
R3692 vdd.n1223 vdd.n1078 39.2114
R3693 vdd.n1389 vdd.n1079 39.2114
R3694 vdd.n1385 vdd.n1080 39.2114
R3695 vdd.n1381 vdd.n1081 39.2114
R3696 vdd.n1377 vdd.n1082 39.2114
R3697 vdd.n1373 vdd.n1083 39.2114
R3698 vdd.n1369 vdd.n1084 39.2114
R3699 vdd.n1365 vdd.n1085 39.2114
R3700 vdd.n1361 vdd.n1086 39.2114
R3701 vdd.n2188 vdd.n2187 37.2369
R3702 vdd.n2224 vdd.n1162 37.2369
R3703 vdd.n2263 vdd.n1122 37.2369
R3704 vdd.n3151 vdd.n724 37.2369
R3705 vdd.n688 vdd.n687 37.2369
R3706 vdd.n3107 vdd.n3106 37.2369
R3707 vdd.n2331 vdd.n1045 31.0639
R3708 vdd.n2580 vdd.n942 31.0639
R3709 vdd.n2513 vdd.n945 31.0639
R3710 vdd.n1281 vdd.n1278 31.0639
R3711 vdd.n2786 vdd.n2783 31.0639
R3712 vdd.n3005 vdd.n3002 31.0639
R3713 vdd.n2852 vdd.n897 31.0639
R3714 vdd.n3066 vdd.n3065 31.0639
R3715 vdd.n2985 vdd.n2984 31.0639
R3716 vdd.n3071 vdd.n771 31.0639
R3717 vdd.n2690 vdd.n2688 31.0639
R3718 vdd.n2859 vdd.n2858 31.0639
R3719 vdd.n2338 vdd.n2337 31.0639
R3720 vdd.n2508 vdd.n2507 31.0639
R3721 vdd.n2440 vdd.n2439 31.0639
R3722 vdd.n1360 vdd.n1359 31.0639
R3723 vdd.n1226 vdd.n1225 30.449
R3724 vdd.n954 vdd.n953 30.449
R3725 vdd.n1273 vdd.n1245 30.449
R3726 vdd.n2518 vdd.n944 30.449
R3727 vdd.n2623 vdd.n2622 30.449
R3728 vdd.n806 vdd.n805 30.449
R3729 vdd.n2791 vdd.n2619 30.449
R3730 vdd.n770 vdd.n769 30.449
R3731 vdd.n1742 vdd.n1508 19.3944
R3732 vdd.n1742 vdd.n1498 19.3944
R3733 vdd.n1754 vdd.n1498 19.3944
R3734 vdd.n1754 vdd.n1496 19.3944
R3735 vdd.n1758 vdd.n1496 19.3944
R3736 vdd.n1758 vdd.n1486 19.3944
R3737 vdd.n1771 vdd.n1486 19.3944
R3738 vdd.n1771 vdd.n1484 19.3944
R3739 vdd.n1775 vdd.n1484 19.3944
R3740 vdd.n1775 vdd.n1476 19.3944
R3741 vdd.n1788 vdd.n1476 19.3944
R3742 vdd.n1788 vdd.n1474 19.3944
R3743 vdd.n1792 vdd.n1474 19.3944
R3744 vdd.n1792 vdd.n1463 19.3944
R3745 vdd.n1804 vdd.n1463 19.3944
R3746 vdd.n1804 vdd.n1461 19.3944
R3747 vdd.n1808 vdd.n1461 19.3944
R3748 vdd.n1808 vdd.n1452 19.3944
R3749 vdd.n2116 vdd.n1452 19.3944
R3750 vdd.n2116 vdd.n1450 19.3944
R3751 vdd.n2120 vdd.n1450 19.3944
R3752 vdd.n2120 vdd.n1441 19.3944
R3753 vdd.n2132 vdd.n1441 19.3944
R3754 vdd.n2132 vdd.n1439 19.3944
R3755 vdd.n2136 vdd.n1439 19.3944
R3756 vdd.n2136 vdd.n1429 19.3944
R3757 vdd.n2149 vdd.n1429 19.3944
R3758 vdd.n2149 vdd.n1427 19.3944
R3759 vdd.n2153 vdd.n1427 19.3944
R3760 vdd.n2153 vdd.n1419 19.3944
R3761 vdd.n2166 vdd.n1419 19.3944
R3762 vdd.n2166 vdd.n1416 19.3944
R3763 vdd.n2172 vdd.n1416 19.3944
R3764 vdd.n2172 vdd.n1417 19.3944
R3765 vdd.n1417 vdd.n1406 19.3944
R3766 vdd.n1661 vdd.n1603 19.3944
R3767 vdd.n1661 vdd.n1660 19.3944
R3768 vdd.n1660 vdd.n1659 19.3944
R3769 vdd.n1659 vdd.n1609 19.3944
R3770 vdd.n1655 vdd.n1609 19.3944
R3771 vdd.n1655 vdd.n1654 19.3944
R3772 vdd.n1654 vdd.n1653 19.3944
R3773 vdd.n1653 vdd.n1615 19.3944
R3774 vdd.n1649 vdd.n1615 19.3944
R3775 vdd.n1649 vdd.n1648 19.3944
R3776 vdd.n1648 vdd.n1647 19.3944
R3777 vdd.n1647 vdd.n1621 19.3944
R3778 vdd.n1643 vdd.n1621 19.3944
R3779 vdd.n1643 vdd.n1642 19.3944
R3780 vdd.n1642 vdd.n1641 19.3944
R3781 vdd.n1641 vdd.n1627 19.3944
R3782 vdd.n1637 vdd.n1627 19.3944
R3783 vdd.n1637 vdd.n1636 19.3944
R3784 vdd.n1636 vdd.n1635 19.3944
R3785 vdd.n1635 vdd.n1633 19.3944
R3786 vdd.n1699 vdd.n1698 19.3944
R3787 vdd.n1698 vdd.n1574 19.3944
R3788 vdd.n1694 vdd.n1574 19.3944
R3789 vdd.n1694 vdd.n1693 19.3944
R3790 vdd.n1693 vdd.n1692 19.3944
R3791 vdd.n1692 vdd.n1580 19.3944
R3792 vdd.n1688 vdd.n1580 19.3944
R3793 vdd.n1688 vdd.n1687 19.3944
R3794 vdd.n1687 vdd.n1686 19.3944
R3795 vdd.n1686 vdd.n1586 19.3944
R3796 vdd.n1682 vdd.n1586 19.3944
R3797 vdd.n1682 vdd.n1681 19.3944
R3798 vdd.n1681 vdd.n1680 19.3944
R3799 vdd.n1680 vdd.n1592 19.3944
R3800 vdd.n1676 vdd.n1592 19.3944
R3801 vdd.n1676 vdd.n1675 19.3944
R3802 vdd.n1675 vdd.n1674 19.3944
R3803 vdd.n1674 vdd.n1598 19.3944
R3804 vdd.n1670 vdd.n1598 19.3944
R3805 vdd.n1670 vdd.n1669 19.3944
R3806 vdd.n1733 vdd.n1732 19.3944
R3807 vdd.n1732 vdd.n1547 19.3944
R3808 vdd.n1728 vdd.n1547 19.3944
R3809 vdd.n1728 vdd.n1727 19.3944
R3810 vdd.n1727 vdd.n1726 19.3944
R3811 vdd.n1726 vdd.n1552 19.3944
R3812 vdd.n1722 vdd.n1552 19.3944
R3813 vdd.n1722 vdd.n1721 19.3944
R3814 vdd.n1721 vdd.n1720 19.3944
R3815 vdd.n1720 vdd.n1558 19.3944
R3816 vdd.n1716 vdd.n1558 19.3944
R3817 vdd.n1716 vdd.n1715 19.3944
R3818 vdd.n1715 vdd.n1714 19.3944
R3819 vdd.n1714 vdd.n1564 19.3944
R3820 vdd.n1710 vdd.n1564 19.3944
R3821 vdd.n1710 vdd.n1709 19.3944
R3822 vdd.n1709 vdd.n1708 19.3944
R3823 vdd.n1708 vdd.n1570 19.3944
R3824 vdd.n2220 vdd.n1160 19.3944
R3825 vdd.n2220 vdd.n1166 19.3944
R3826 vdd.n2215 vdd.n1166 19.3944
R3827 vdd.n2215 vdd.n2214 19.3944
R3828 vdd.n2214 vdd.n2213 19.3944
R3829 vdd.n2213 vdd.n1173 19.3944
R3830 vdd.n2208 vdd.n1173 19.3944
R3831 vdd.n2208 vdd.n2207 19.3944
R3832 vdd.n2207 vdd.n2206 19.3944
R3833 vdd.n2206 vdd.n1180 19.3944
R3834 vdd.n2201 vdd.n1180 19.3944
R3835 vdd.n2201 vdd.n2200 19.3944
R3836 vdd.n2200 vdd.n2199 19.3944
R3837 vdd.n2199 vdd.n1187 19.3944
R3838 vdd.n2194 vdd.n1187 19.3944
R3839 vdd.n2194 vdd.n2193 19.3944
R3840 vdd.n1399 vdd.n1192 19.3944
R3841 vdd.n2189 vdd.n1396 19.3944
R3842 vdd.n2259 vdd.n1120 19.3944
R3843 vdd.n2259 vdd.n1126 19.3944
R3844 vdd.n2254 vdd.n1126 19.3944
R3845 vdd.n2254 vdd.n2253 19.3944
R3846 vdd.n2253 vdd.n2252 19.3944
R3847 vdd.n2252 vdd.n1133 19.3944
R3848 vdd.n2247 vdd.n1133 19.3944
R3849 vdd.n2247 vdd.n2246 19.3944
R3850 vdd.n2246 vdd.n2245 19.3944
R3851 vdd.n2245 vdd.n1140 19.3944
R3852 vdd.n2240 vdd.n1140 19.3944
R3853 vdd.n2240 vdd.n2239 19.3944
R3854 vdd.n2239 vdd.n2238 19.3944
R3855 vdd.n2238 vdd.n1147 19.3944
R3856 vdd.n2233 vdd.n1147 19.3944
R3857 vdd.n2233 vdd.n2232 19.3944
R3858 vdd.n2232 vdd.n2231 19.3944
R3859 vdd.n2231 vdd.n1154 19.3944
R3860 vdd.n2226 vdd.n1154 19.3944
R3861 vdd.n2226 vdd.n2225 19.3944
R3862 vdd.n2296 vdd.n1095 19.3944
R3863 vdd.n2296 vdd.n1096 19.3944
R3864 vdd.n2291 vdd.n2290 19.3944
R3865 vdd.n2286 vdd.n2285 19.3944
R3866 vdd.n2285 vdd.n2284 19.3944
R3867 vdd.n2284 vdd.n1100 19.3944
R3868 vdd.n2279 vdd.n1100 19.3944
R3869 vdd.n2279 vdd.n2278 19.3944
R3870 vdd.n2278 vdd.n2277 19.3944
R3871 vdd.n2277 vdd.n1107 19.3944
R3872 vdd.n2272 vdd.n1107 19.3944
R3873 vdd.n2272 vdd.n2271 19.3944
R3874 vdd.n2271 vdd.n2270 19.3944
R3875 vdd.n2270 vdd.n1114 19.3944
R3876 vdd.n2265 vdd.n1114 19.3944
R3877 vdd.n2265 vdd.n2264 19.3944
R3878 vdd.n1746 vdd.n1504 19.3944
R3879 vdd.n1746 vdd.n1502 19.3944
R3880 vdd.n1750 vdd.n1502 19.3944
R3881 vdd.n1750 vdd.n1492 19.3944
R3882 vdd.n1763 vdd.n1492 19.3944
R3883 vdd.n1763 vdd.n1490 19.3944
R3884 vdd.n1767 vdd.n1490 19.3944
R3885 vdd.n1767 vdd.n1481 19.3944
R3886 vdd.n1780 vdd.n1481 19.3944
R3887 vdd.n1780 vdd.n1479 19.3944
R3888 vdd.n1784 vdd.n1479 19.3944
R3889 vdd.n1784 vdd.n1470 19.3944
R3890 vdd.n1796 vdd.n1470 19.3944
R3891 vdd.n1796 vdd.n1468 19.3944
R3892 vdd.n1800 vdd.n1468 19.3944
R3893 vdd.n1800 vdd.n1458 19.3944
R3894 vdd.n1813 vdd.n1458 19.3944
R3895 vdd.n1813 vdd.n1456 19.3944
R3896 vdd.n2112 vdd.n1456 19.3944
R3897 vdd.n2112 vdd.n1447 19.3944
R3898 vdd.n2124 vdd.n1447 19.3944
R3899 vdd.n2124 vdd.n1445 19.3944
R3900 vdd.n2128 vdd.n1445 19.3944
R3901 vdd.n2128 vdd.n1435 19.3944
R3902 vdd.n2141 vdd.n1435 19.3944
R3903 vdd.n2141 vdd.n1433 19.3944
R3904 vdd.n2145 vdd.n1433 19.3944
R3905 vdd.n2145 vdd.n1424 19.3944
R3906 vdd.n2158 vdd.n1424 19.3944
R3907 vdd.n2158 vdd.n1422 19.3944
R3908 vdd.n2162 vdd.n1422 19.3944
R3909 vdd.n2162 vdd.n1412 19.3944
R3910 vdd.n2176 vdd.n1412 19.3944
R3911 vdd.n2176 vdd.n1410 19.3944
R3912 vdd.n2180 vdd.n1410 19.3944
R3913 vdd.n3239 vdd.n655 19.3944
R3914 vdd.n3243 vdd.n655 19.3944
R3915 vdd.n3243 vdd.n646 19.3944
R3916 vdd.n3255 vdd.n646 19.3944
R3917 vdd.n3255 vdd.n644 19.3944
R3918 vdd.n3259 vdd.n644 19.3944
R3919 vdd.n3259 vdd.n633 19.3944
R3920 vdd.n3271 vdd.n633 19.3944
R3921 vdd.n3271 vdd.n631 19.3944
R3922 vdd.n3275 vdd.n631 19.3944
R3923 vdd.n3275 vdd.n622 19.3944
R3924 vdd.n3288 vdd.n622 19.3944
R3925 vdd.n3288 vdd.n620 19.3944
R3926 vdd.n3295 vdd.n620 19.3944
R3927 vdd.n3295 vdd.n3294 19.3944
R3928 vdd.n3294 vdd.n610 19.3944
R3929 vdd.n3308 vdd.n610 19.3944
R3930 vdd.n3309 vdd.n3308 19.3944
R3931 vdd.n3310 vdd.n3309 19.3944
R3932 vdd.n3310 vdd.n608 19.3944
R3933 vdd.n3315 vdd.n608 19.3944
R3934 vdd.n3316 vdd.n3315 19.3944
R3935 vdd.n3317 vdd.n3316 19.3944
R3936 vdd.n3317 vdd.n606 19.3944
R3937 vdd.n3322 vdd.n606 19.3944
R3938 vdd.n3323 vdd.n3322 19.3944
R3939 vdd.n3324 vdd.n3323 19.3944
R3940 vdd.n3324 vdd.n604 19.3944
R3941 vdd.n3330 vdd.n604 19.3944
R3942 vdd.n3331 vdd.n3330 19.3944
R3943 vdd.n3332 vdd.n3331 19.3944
R3944 vdd.n3332 vdd.n602 19.3944
R3945 vdd.n3337 vdd.n602 19.3944
R3946 vdd.n3338 vdd.n3337 19.3944
R3947 vdd.n3339 vdd.n3338 19.3944
R3948 vdd.n550 vdd.n417 19.3944
R3949 vdd.n556 vdd.n417 19.3944
R3950 vdd.n557 vdd.n556 19.3944
R3951 vdd.n560 vdd.n557 19.3944
R3952 vdd.n560 vdd.n415 19.3944
R3953 vdd.n566 vdd.n415 19.3944
R3954 vdd.n567 vdd.n566 19.3944
R3955 vdd.n570 vdd.n567 19.3944
R3956 vdd.n570 vdd.n413 19.3944
R3957 vdd.n576 vdd.n413 19.3944
R3958 vdd.n577 vdd.n576 19.3944
R3959 vdd.n580 vdd.n577 19.3944
R3960 vdd.n580 vdd.n411 19.3944
R3961 vdd.n586 vdd.n411 19.3944
R3962 vdd.n587 vdd.n586 19.3944
R3963 vdd.n590 vdd.n587 19.3944
R3964 vdd.n590 vdd.n409 19.3944
R3965 vdd.n596 vdd.n409 19.3944
R3966 vdd.n598 vdd.n596 19.3944
R3967 vdd.n599 vdd.n598 19.3944
R3968 vdd.n497 vdd.n496 19.3944
R3969 vdd.n500 vdd.n497 19.3944
R3970 vdd.n500 vdd.n429 19.3944
R3971 vdd.n506 vdd.n429 19.3944
R3972 vdd.n507 vdd.n506 19.3944
R3973 vdd.n510 vdd.n507 19.3944
R3974 vdd.n510 vdd.n427 19.3944
R3975 vdd.n516 vdd.n427 19.3944
R3976 vdd.n517 vdd.n516 19.3944
R3977 vdd.n520 vdd.n517 19.3944
R3978 vdd.n520 vdd.n425 19.3944
R3979 vdd.n526 vdd.n425 19.3944
R3980 vdd.n527 vdd.n526 19.3944
R3981 vdd.n530 vdd.n527 19.3944
R3982 vdd.n530 vdd.n423 19.3944
R3983 vdd.n536 vdd.n423 19.3944
R3984 vdd.n537 vdd.n536 19.3944
R3985 vdd.n540 vdd.n537 19.3944
R3986 vdd.n540 vdd.n421 19.3944
R3987 vdd.n546 vdd.n421 19.3944
R3988 vdd.n447 vdd.n446 19.3944
R3989 vdd.n450 vdd.n447 19.3944
R3990 vdd.n450 vdd.n441 19.3944
R3991 vdd.n456 vdd.n441 19.3944
R3992 vdd.n457 vdd.n456 19.3944
R3993 vdd.n460 vdd.n457 19.3944
R3994 vdd.n460 vdd.n439 19.3944
R3995 vdd.n466 vdd.n439 19.3944
R3996 vdd.n467 vdd.n466 19.3944
R3997 vdd.n470 vdd.n467 19.3944
R3998 vdd.n470 vdd.n437 19.3944
R3999 vdd.n476 vdd.n437 19.3944
R4000 vdd.n477 vdd.n476 19.3944
R4001 vdd.n480 vdd.n477 19.3944
R4002 vdd.n480 vdd.n435 19.3944
R4003 vdd.n486 vdd.n435 19.3944
R4004 vdd.n487 vdd.n486 19.3944
R4005 vdd.n490 vdd.n487 19.3944
R4006 vdd.n3235 vdd.n652 19.3944
R4007 vdd.n3247 vdd.n652 19.3944
R4008 vdd.n3247 vdd.n650 19.3944
R4009 vdd.n3251 vdd.n650 19.3944
R4010 vdd.n3251 vdd.n640 19.3944
R4011 vdd.n3263 vdd.n640 19.3944
R4012 vdd.n3263 vdd.n638 19.3944
R4013 vdd.n3267 vdd.n638 19.3944
R4014 vdd.n3267 vdd.n628 19.3944
R4015 vdd.n3280 vdd.n628 19.3944
R4016 vdd.n3280 vdd.n626 19.3944
R4017 vdd.n3284 vdd.n626 19.3944
R4018 vdd.n3284 vdd.n617 19.3944
R4019 vdd.n3299 vdd.n617 19.3944
R4020 vdd.n3299 vdd.n615 19.3944
R4021 vdd.n3303 vdd.n615 19.3944
R4022 vdd.n3303 vdd.n324 19.3944
R4023 vdd.n3381 vdd.n324 19.3944
R4024 vdd.n3381 vdd.n325 19.3944
R4025 vdd.n3375 vdd.n325 19.3944
R4026 vdd.n3375 vdd.n3374 19.3944
R4027 vdd.n3374 vdd.n3373 19.3944
R4028 vdd.n3373 vdd.n337 19.3944
R4029 vdd.n3367 vdd.n337 19.3944
R4030 vdd.n3367 vdd.n3366 19.3944
R4031 vdd.n3366 vdd.n3365 19.3944
R4032 vdd.n3365 vdd.n347 19.3944
R4033 vdd.n3359 vdd.n347 19.3944
R4034 vdd.n3359 vdd.n3358 19.3944
R4035 vdd.n3358 vdd.n3357 19.3944
R4036 vdd.n3357 vdd.n358 19.3944
R4037 vdd.n3351 vdd.n358 19.3944
R4038 vdd.n3351 vdd.n3350 19.3944
R4039 vdd.n3350 vdd.n3349 19.3944
R4040 vdd.n3349 vdd.n369 19.3944
R4041 vdd.n3192 vdd.n3191 19.3944
R4042 vdd.n3191 vdd.n3190 19.3944
R4043 vdd.n3190 vdd.n694 19.3944
R4044 vdd.n3184 vdd.n694 19.3944
R4045 vdd.n3184 vdd.n3183 19.3944
R4046 vdd.n3183 vdd.n3182 19.3944
R4047 vdd.n3182 vdd.n700 19.3944
R4048 vdd.n3176 vdd.n700 19.3944
R4049 vdd.n3176 vdd.n3175 19.3944
R4050 vdd.n3175 vdd.n3174 19.3944
R4051 vdd.n3174 vdd.n706 19.3944
R4052 vdd.n3168 vdd.n706 19.3944
R4053 vdd.n3168 vdd.n3167 19.3944
R4054 vdd.n3167 vdd.n3166 19.3944
R4055 vdd.n3166 vdd.n712 19.3944
R4056 vdd.n3160 vdd.n712 19.3944
R4057 vdd.n3160 vdd.n3159 19.3944
R4058 vdd.n3159 vdd.n3158 19.3944
R4059 vdd.n3158 vdd.n718 19.3944
R4060 vdd.n3152 vdd.n718 19.3944
R4061 vdd.n3232 vdd.n3231 19.3944
R4062 vdd.n3231 vdd.n662 19.3944
R4063 vdd.n3226 vdd.n3225 19.3944
R4064 vdd.n3222 vdd.n3221 19.3944
R4065 vdd.n3221 vdd.n668 19.3944
R4066 vdd.n3216 vdd.n668 19.3944
R4067 vdd.n3216 vdd.n3215 19.3944
R4068 vdd.n3215 vdd.n3214 19.3944
R4069 vdd.n3214 vdd.n674 19.3944
R4070 vdd.n3208 vdd.n674 19.3944
R4071 vdd.n3208 vdd.n3207 19.3944
R4072 vdd.n3207 vdd.n3206 19.3944
R4073 vdd.n3206 vdd.n680 19.3944
R4074 vdd.n3200 vdd.n680 19.3944
R4075 vdd.n3200 vdd.n3199 19.3944
R4076 vdd.n3199 vdd.n3198 19.3944
R4077 vdd.n3147 vdd.n722 19.3944
R4078 vdd.n3147 vdd.n726 19.3944
R4079 vdd.n3142 vdd.n726 19.3944
R4080 vdd.n3142 vdd.n3141 19.3944
R4081 vdd.n3141 vdd.n732 19.3944
R4082 vdd.n3136 vdd.n732 19.3944
R4083 vdd.n3136 vdd.n3135 19.3944
R4084 vdd.n3135 vdd.n3134 19.3944
R4085 vdd.n3134 vdd.n738 19.3944
R4086 vdd.n3128 vdd.n738 19.3944
R4087 vdd.n3128 vdd.n3127 19.3944
R4088 vdd.n3127 vdd.n3126 19.3944
R4089 vdd.n3126 vdd.n744 19.3944
R4090 vdd.n3120 vdd.n744 19.3944
R4091 vdd.n3120 vdd.n3119 19.3944
R4092 vdd.n3119 vdd.n3118 19.3944
R4093 vdd.n3114 vdd.n3113 19.3944
R4094 vdd.n3110 vdd.n3109 19.3944
R4095 vdd.n1668 vdd.n1603 19.0066
R4096 vdd.n2224 vdd.n1160 19.0066
R4097 vdd.n550 vdd.n547 19.0066
R4098 vdd.n3151 vdd.n722 19.0066
R4099 vdd.n1736 vdd.n1506 18.5924
R4100 vdd.n2182 vdd.n1054 18.5924
R4101 vdd.n3237 vdd.n658 18.5924
R4102 vdd.n3346 vdd.n3345 18.5924
R4103 vdd.n1225 vdd.n1224 16.0975
R4104 vdd.n953 vdd.n952 16.0975
R4105 vdd.n1511 vdd.n1510 16.0975
R4106 vdd.n1667 vdd.n1666 16.0975
R4107 vdd.n1703 vdd.n1702 16.0975
R4108 vdd.n2187 vdd.n2186 16.0975
R4109 vdd.n1162 vdd.n1161 16.0975
R4110 vdd.n1122 vdd.n1121 16.0975
R4111 vdd.n1245 vdd.n1244 16.0975
R4112 vdd.n944 vdd.n943 16.0975
R4113 vdd.n2622 vdd.n2621 16.0975
R4114 vdd.n406 vdd.n405 16.0975
R4115 vdd.n420 vdd.n419 16.0975
R4116 vdd.n432 vdd.n431 16.0975
R4117 vdd.n724 vdd.n723 16.0975
R4118 vdd.n687 vdd.n686 16.0975
R4119 vdd.n805 vdd.n804 16.0975
R4120 vdd.n2619 vdd.n2618 16.0975
R4121 vdd.n3106 vdd.n3105 16.0975
R4122 vdd.n769 vdd.n768 16.0975
R4123 vdd.t26 vdd.n2582 15.4182
R4124 vdd.n2855 vdd.t14 15.4182
R4125 vdd.n28 vdd.n27 15.0023
R4126 vdd.n2334 vdd.n1047 14.0578
R4127 vdd.n3068 vdd.n756 14.0578
R4128 vdd.n316 vdd.n281 13.1884
R4129 vdd.n261 vdd.n226 13.1884
R4130 vdd.n218 vdd.n183 13.1884
R4131 vdd.n163 vdd.n128 13.1884
R4132 vdd.n121 vdd.n86 13.1884
R4133 vdd.n66 vdd.n31 13.1884
R4134 vdd.n2047 vdd.n2012 13.1884
R4135 vdd.n2102 vdd.n2067 13.1884
R4136 vdd.n1949 vdd.n1914 13.1884
R4137 vdd.n2004 vdd.n1969 13.1884
R4138 vdd.n1852 vdd.n1817 13.1884
R4139 vdd.n1907 vdd.n1872 13.1884
R4140 vdd.n1704 vdd.n1699 12.9944
R4141 vdd.n1704 vdd.n1570 12.9944
R4142 vdd.n2263 vdd.n1120 12.9944
R4143 vdd.n2264 vdd.n2263 12.9944
R4144 vdd.n496 vdd.n433 12.9944
R4145 vdd.n490 vdd.n433 12.9944
R4146 vdd.n3192 vdd.n688 12.9944
R4147 vdd.n3198 vdd.n688 12.9944
R4148 vdd.n317 vdd.n279 12.8005
R4149 vdd.n312 vdd.n283 12.8005
R4150 vdd.n262 vdd.n224 12.8005
R4151 vdd.n257 vdd.n228 12.8005
R4152 vdd.n219 vdd.n181 12.8005
R4153 vdd.n214 vdd.n185 12.8005
R4154 vdd.n164 vdd.n126 12.8005
R4155 vdd.n159 vdd.n130 12.8005
R4156 vdd.n122 vdd.n84 12.8005
R4157 vdd.n117 vdd.n88 12.8005
R4158 vdd.n67 vdd.n29 12.8005
R4159 vdd.n62 vdd.n33 12.8005
R4160 vdd.n2048 vdd.n2010 12.8005
R4161 vdd.n2043 vdd.n2014 12.8005
R4162 vdd.n2103 vdd.n2065 12.8005
R4163 vdd.n2098 vdd.n2069 12.8005
R4164 vdd.n1950 vdd.n1912 12.8005
R4165 vdd.n1945 vdd.n1916 12.8005
R4166 vdd.n2005 vdd.n1967 12.8005
R4167 vdd.n2000 vdd.n1971 12.8005
R4168 vdd.n1853 vdd.n1815 12.8005
R4169 vdd.n1848 vdd.n1819 12.8005
R4170 vdd.n1908 vdd.n1870 12.8005
R4171 vdd.n1903 vdd.n1874 12.8005
R4172 vdd.n311 vdd.n284 12.0247
R4173 vdd.n256 vdd.n229 12.0247
R4174 vdd.n213 vdd.n186 12.0247
R4175 vdd.n158 vdd.n131 12.0247
R4176 vdd.n116 vdd.n89 12.0247
R4177 vdd.n61 vdd.n34 12.0247
R4178 vdd.n2042 vdd.n2015 12.0247
R4179 vdd.n2097 vdd.n2070 12.0247
R4180 vdd.n1944 vdd.n1917 12.0247
R4181 vdd.n1999 vdd.n1972 12.0247
R4182 vdd.n1847 vdd.n1820 12.0247
R4183 vdd.n1902 vdd.n1875 12.0247
R4184 vdd.n1744 vdd.n1506 11.337
R4185 vdd.n1752 vdd.n1500 11.337
R4186 vdd.n1752 vdd.n1494 11.337
R4187 vdd.n1761 vdd.n1494 11.337
R4188 vdd.n1769 vdd.n1488 11.337
R4189 vdd.n1778 vdd.n1777 11.337
R4190 vdd.n1794 vdd.n1472 11.337
R4191 vdd.n1802 vdd.n1465 11.337
R4192 vdd.n1811 vdd.n1810 11.337
R4193 vdd.n2114 vdd.n1454 11.337
R4194 vdd.n2130 vdd.n1443 11.337
R4195 vdd.n2139 vdd.n1437 11.337
R4196 vdd.n2147 vdd.n1431 11.337
R4197 vdd.n2156 vdd.n2155 11.337
R4198 vdd.n2164 vdd.n1414 11.337
R4199 vdd.n2174 vdd.n1414 11.337
R4200 vdd.n2182 vdd.n1407 11.337
R4201 vdd.n3237 vdd.n659 11.337
R4202 vdd.n3245 vdd.n648 11.337
R4203 vdd.n3253 vdd.n648 11.337
R4204 vdd.n3261 vdd.n642 11.337
R4205 vdd.n3269 vdd.n635 11.337
R4206 vdd.n3278 vdd.n3277 11.337
R4207 vdd.n3286 vdd.n624 11.337
R4208 vdd.n3305 vdd.n613 11.337
R4209 vdd.n3379 vdd.n328 11.337
R4210 vdd.n3377 vdd.n332 11.337
R4211 vdd.n3371 vdd.n3370 11.337
R4212 vdd.n3363 vdd.n349 11.337
R4213 vdd.n3362 vdd.n3361 11.337
R4214 vdd.n3355 vdd.n3354 11.337
R4215 vdd.n3354 vdd.n3353 11.337
R4216 vdd.n3353 vdd.n363 11.337
R4217 vdd.n3347 vdd.n3346 11.337
R4218 vdd.n308 vdd.n307 11.249
R4219 vdd.n253 vdd.n252 11.249
R4220 vdd.n210 vdd.n209 11.249
R4221 vdd.n155 vdd.n154 11.249
R4222 vdd.n113 vdd.n112 11.249
R4223 vdd.n58 vdd.n57 11.249
R4224 vdd.n2039 vdd.n2038 11.249
R4225 vdd.n2094 vdd.n2093 11.249
R4226 vdd.n1941 vdd.n1940 11.249
R4227 vdd.n1996 vdd.n1995 11.249
R4228 vdd.n1844 vdd.n1843 11.249
R4229 vdd.n1899 vdd.n1898 11.249
R4230 vdd.n2164 vdd.t179 10.7702
R4231 vdd.n3253 vdd.t177 10.7702
R4232 vdd.n293 vdd.n292 10.7238
R4233 vdd.n238 vdd.n237 10.7238
R4234 vdd.n195 vdd.n194 10.7238
R4235 vdd.n140 vdd.n139 10.7238
R4236 vdd.n98 vdd.n97 10.7238
R4237 vdd.n43 vdd.n42 10.7238
R4238 vdd.n2024 vdd.n2023 10.7238
R4239 vdd.n2079 vdd.n2078 10.7238
R4240 vdd.n1926 vdd.n1925 10.7238
R4241 vdd.n1981 vdd.n1980 10.7238
R4242 vdd.n1829 vdd.n1828 10.7238
R4243 vdd.n1884 vdd.n1883 10.7238
R4244 vdd.n2510 vdd.t266 10.6568
R4245 vdd.t17 vdd.n899 10.6568
R4246 vdd.n2343 vdd.n1045 10.6151
R4247 vdd.n2344 vdd.n2343 10.6151
R4248 vdd.n2345 vdd.n2344 10.6151
R4249 vdd.n2345 vdd.n1034 10.6151
R4250 vdd.n2355 vdd.n1034 10.6151
R4251 vdd.n2356 vdd.n2355 10.6151
R4252 vdd.n2357 vdd.n2356 10.6151
R4253 vdd.n2357 vdd.n1021 10.6151
R4254 vdd.n2367 vdd.n1021 10.6151
R4255 vdd.n2368 vdd.n2367 10.6151
R4256 vdd.n2369 vdd.n2368 10.6151
R4257 vdd.n2369 vdd.n1009 10.6151
R4258 vdd.n2380 vdd.n1009 10.6151
R4259 vdd.n2381 vdd.n2380 10.6151
R4260 vdd.n2382 vdd.n2381 10.6151
R4261 vdd.n2382 vdd.n997 10.6151
R4262 vdd.n2392 vdd.n997 10.6151
R4263 vdd.n2393 vdd.n2392 10.6151
R4264 vdd.n2394 vdd.n2393 10.6151
R4265 vdd.n2394 vdd.n985 10.6151
R4266 vdd.n2404 vdd.n985 10.6151
R4267 vdd.n2405 vdd.n2404 10.6151
R4268 vdd.n2406 vdd.n2405 10.6151
R4269 vdd.n2406 vdd.n974 10.6151
R4270 vdd.n2416 vdd.n974 10.6151
R4271 vdd.n2417 vdd.n2416 10.6151
R4272 vdd.n2418 vdd.n2417 10.6151
R4273 vdd.n2418 vdd.n961 10.6151
R4274 vdd.n2430 vdd.n961 10.6151
R4275 vdd.n2431 vdd.n2430 10.6151
R4276 vdd.n2433 vdd.n2431 10.6151
R4277 vdd.n2433 vdd.n2432 10.6151
R4278 vdd.n2432 vdd.n942 10.6151
R4279 vdd.n2580 vdd.n2579 10.6151
R4280 vdd.n2579 vdd.n2578 10.6151
R4281 vdd.n2578 vdd.n2575 10.6151
R4282 vdd.n2575 vdd.n2574 10.6151
R4283 vdd.n2574 vdd.n2571 10.6151
R4284 vdd.n2571 vdd.n2570 10.6151
R4285 vdd.n2570 vdd.n2567 10.6151
R4286 vdd.n2567 vdd.n2566 10.6151
R4287 vdd.n2566 vdd.n2563 10.6151
R4288 vdd.n2563 vdd.n2562 10.6151
R4289 vdd.n2562 vdd.n2559 10.6151
R4290 vdd.n2559 vdd.n2558 10.6151
R4291 vdd.n2558 vdd.n2555 10.6151
R4292 vdd.n2555 vdd.n2554 10.6151
R4293 vdd.n2554 vdd.n2551 10.6151
R4294 vdd.n2551 vdd.n2550 10.6151
R4295 vdd.n2550 vdd.n2547 10.6151
R4296 vdd.n2547 vdd.n2546 10.6151
R4297 vdd.n2546 vdd.n2543 10.6151
R4298 vdd.n2543 vdd.n2542 10.6151
R4299 vdd.n2542 vdd.n2539 10.6151
R4300 vdd.n2539 vdd.n2538 10.6151
R4301 vdd.n2538 vdd.n2535 10.6151
R4302 vdd.n2535 vdd.n2534 10.6151
R4303 vdd.n2534 vdd.n2531 10.6151
R4304 vdd.n2531 vdd.n2530 10.6151
R4305 vdd.n2530 vdd.n2527 10.6151
R4306 vdd.n2527 vdd.n2526 10.6151
R4307 vdd.n2526 vdd.n2523 10.6151
R4308 vdd.n2523 vdd.n2522 10.6151
R4309 vdd.n2522 vdd.n2519 10.6151
R4310 vdd.n2517 vdd.n2514 10.6151
R4311 vdd.n2514 vdd.n2513 10.6151
R4312 vdd.n1282 vdd.n1281 10.6151
R4313 vdd.n1284 vdd.n1282 10.6151
R4314 vdd.n1285 vdd.n1284 10.6151
R4315 vdd.n1287 vdd.n1285 10.6151
R4316 vdd.n1288 vdd.n1287 10.6151
R4317 vdd.n1290 vdd.n1288 10.6151
R4318 vdd.n1291 vdd.n1290 10.6151
R4319 vdd.n1293 vdd.n1291 10.6151
R4320 vdd.n1294 vdd.n1293 10.6151
R4321 vdd.n1296 vdd.n1294 10.6151
R4322 vdd.n1297 vdd.n1296 10.6151
R4323 vdd.n1299 vdd.n1297 10.6151
R4324 vdd.n1300 vdd.n1299 10.6151
R4325 vdd.n1302 vdd.n1300 10.6151
R4326 vdd.n1303 vdd.n1302 10.6151
R4327 vdd.n1305 vdd.n1303 10.6151
R4328 vdd.n1306 vdd.n1305 10.6151
R4329 vdd.n1328 vdd.n1306 10.6151
R4330 vdd.n1328 vdd.n1327 10.6151
R4331 vdd.n1327 vdd.n1326 10.6151
R4332 vdd.n1326 vdd.n1324 10.6151
R4333 vdd.n1324 vdd.n1323 10.6151
R4334 vdd.n1323 vdd.n1321 10.6151
R4335 vdd.n1321 vdd.n1320 10.6151
R4336 vdd.n1320 vdd.n1318 10.6151
R4337 vdd.n1318 vdd.n1317 10.6151
R4338 vdd.n1317 vdd.n1315 10.6151
R4339 vdd.n1315 vdd.n1314 10.6151
R4340 vdd.n1314 vdd.n1312 10.6151
R4341 vdd.n1312 vdd.n1311 10.6151
R4342 vdd.n1311 vdd.n1308 10.6151
R4343 vdd.n1308 vdd.n1307 10.6151
R4344 vdd.n1307 vdd.n945 10.6151
R4345 vdd.n2331 vdd.n2330 10.6151
R4346 vdd.n2330 vdd.n2329 10.6151
R4347 vdd.n2329 vdd.n2328 10.6151
R4348 vdd.n2328 vdd.n2326 10.6151
R4349 vdd.n2326 vdd.n2323 10.6151
R4350 vdd.n2323 vdd.n2322 10.6151
R4351 vdd.n2322 vdd.n2319 10.6151
R4352 vdd.n2319 vdd.n2318 10.6151
R4353 vdd.n2318 vdd.n2315 10.6151
R4354 vdd.n2315 vdd.n2314 10.6151
R4355 vdd.n2314 vdd.n2311 10.6151
R4356 vdd.n2311 vdd.n2310 10.6151
R4357 vdd.n2310 vdd.n2307 10.6151
R4358 vdd.n2307 vdd.n2306 10.6151
R4359 vdd.n2306 vdd.n2303 10.6151
R4360 vdd.n2303 vdd.n2302 10.6151
R4361 vdd.n2302 vdd.n2299 10.6151
R4362 vdd.n2299 vdd.n1090 10.6151
R4363 vdd.n1248 vdd.n1090 10.6151
R4364 vdd.n1249 vdd.n1248 10.6151
R4365 vdd.n1252 vdd.n1249 10.6151
R4366 vdd.n1253 vdd.n1252 10.6151
R4367 vdd.n1256 vdd.n1253 10.6151
R4368 vdd.n1257 vdd.n1256 10.6151
R4369 vdd.n1260 vdd.n1257 10.6151
R4370 vdd.n1261 vdd.n1260 10.6151
R4371 vdd.n1264 vdd.n1261 10.6151
R4372 vdd.n1265 vdd.n1264 10.6151
R4373 vdd.n1268 vdd.n1265 10.6151
R4374 vdd.n1269 vdd.n1268 10.6151
R4375 vdd.n1272 vdd.n1269 10.6151
R4376 vdd.n1277 vdd.n1274 10.6151
R4377 vdd.n1278 vdd.n1277 10.6151
R4378 vdd.n2783 vdd.n2782 10.6151
R4379 vdd.n2782 vdd.n2781 10.6151
R4380 vdd.n2781 vdd.n2620 10.6151
R4381 vdd.n2725 vdd.n2620 10.6151
R4382 vdd.n2726 vdd.n2725 10.6151
R4383 vdd.n2728 vdd.n2726 10.6151
R4384 vdd.n2729 vdd.n2728 10.6151
R4385 vdd.n2731 vdd.n2729 10.6151
R4386 vdd.n2732 vdd.n2731 10.6151
R4387 vdd.n2762 vdd.n2732 10.6151
R4388 vdd.n2762 vdd.n2761 10.6151
R4389 vdd.n2761 vdd.n2760 10.6151
R4390 vdd.n2760 vdd.n2758 10.6151
R4391 vdd.n2758 vdd.n2757 10.6151
R4392 vdd.n2757 vdd.n2755 10.6151
R4393 vdd.n2755 vdd.n2754 10.6151
R4394 vdd.n2754 vdd.n2752 10.6151
R4395 vdd.n2752 vdd.n2751 10.6151
R4396 vdd.n2751 vdd.n2749 10.6151
R4397 vdd.n2749 vdd.n2748 10.6151
R4398 vdd.n2748 vdd.n2746 10.6151
R4399 vdd.n2746 vdd.n2745 10.6151
R4400 vdd.n2745 vdd.n2743 10.6151
R4401 vdd.n2743 vdd.n2742 10.6151
R4402 vdd.n2742 vdd.n2740 10.6151
R4403 vdd.n2740 vdd.n2739 10.6151
R4404 vdd.n2739 vdd.n2737 10.6151
R4405 vdd.n2737 vdd.n2736 10.6151
R4406 vdd.n2736 vdd.n2734 10.6151
R4407 vdd.n2734 vdd.n2733 10.6151
R4408 vdd.n2733 vdd.n807 10.6151
R4409 vdd.n3001 vdd.n807 10.6151
R4410 vdd.n3002 vdd.n3001 10.6151
R4411 vdd.n2852 vdd.n2851 10.6151
R4412 vdd.n2851 vdd.n2850 10.6151
R4413 vdd.n2850 vdd.n2849 10.6151
R4414 vdd.n2849 vdd.n2847 10.6151
R4415 vdd.n2847 vdd.n2844 10.6151
R4416 vdd.n2844 vdd.n2843 10.6151
R4417 vdd.n2843 vdd.n2840 10.6151
R4418 vdd.n2840 vdd.n2839 10.6151
R4419 vdd.n2839 vdd.n2836 10.6151
R4420 vdd.n2836 vdd.n2835 10.6151
R4421 vdd.n2835 vdd.n2832 10.6151
R4422 vdd.n2832 vdd.n2831 10.6151
R4423 vdd.n2831 vdd.n2828 10.6151
R4424 vdd.n2828 vdd.n2827 10.6151
R4425 vdd.n2827 vdd.n2824 10.6151
R4426 vdd.n2824 vdd.n2823 10.6151
R4427 vdd.n2823 vdd.n2820 10.6151
R4428 vdd.n2820 vdd.n2819 10.6151
R4429 vdd.n2819 vdd.n2816 10.6151
R4430 vdd.n2816 vdd.n2815 10.6151
R4431 vdd.n2815 vdd.n2812 10.6151
R4432 vdd.n2812 vdd.n2811 10.6151
R4433 vdd.n2811 vdd.n2808 10.6151
R4434 vdd.n2808 vdd.n2807 10.6151
R4435 vdd.n2807 vdd.n2804 10.6151
R4436 vdd.n2804 vdd.n2803 10.6151
R4437 vdd.n2803 vdd.n2800 10.6151
R4438 vdd.n2800 vdd.n2799 10.6151
R4439 vdd.n2799 vdd.n2796 10.6151
R4440 vdd.n2796 vdd.n2795 10.6151
R4441 vdd.n2795 vdd.n2792 10.6151
R4442 vdd.n2790 vdd.n2787 10.6151
R4443 vdd.n2787 vdd.n2786 10.6151
R4444 vdd.n2864 vdd.n897 10.6151
R4445 vdd.n2865 vdd.n2864 10.6151
R4446 vdd.n2866 vdd.n2865 10.6151
R4447 vdd.n2866 vdd.n886 10.6151
R4448 vdd.n2876 vdd.n886 10.6151
R4449 vdd.n2877 vdd.n2876 10.6151
R4450 vdd.n2878 vdd.n2877 10.6151
R4451 vdd.n2878 vdd.n874 10.6151
R4452 vdd.n2888 vdd.n874 10.6151
R4453 vdd.n2889 vdd.n2888 10.6151
R4454 vdd.n2890 vdd.n2889 10.6151
R4455 vdd.n2890 vdd.n862 10.6151
R4456 vdd.n2900 vdd.n862 10.6151
R4457 vdd.n2901 vdd.n2900 10.6151
R4458 vdd.n2902 vdd.n2901 10.6151
R4459 vdd.n2902 vdd.n851 10.6151
R4460 vdd.n2912 vdd.n851 10.6151
R4461 vdd.n2913 vdd.n2912 10.6151
R4462 vdd.n2914 vdd.n2913 10.6151
R4463 vdd.n2914 vdd.n837 10.6151
R4464 vdd.n2925 vdd.n837 10.6151
R4465 vdd.n2926 vdd.n2925 10.6151
R4466 vdd.n2927 vdd.n2926 10.6151
R4467 vdd.n2927 vdd.n826 10.6151
R4468 vdd.n2937 vdd.n826 10.6151
R4469 vdd.n2938 vdd.n2937 10.6151
R4470 vdd.n2939 vdd.n2938 10.6151
R4471 vdd.n2939 vdd.n812 10.6151
R4472 vdd.n2994 vdd.n812 10.6151
R4473 vdd.n2995 vdd.n2994 10.6151
R4474 vdd.n2996 vdd.n2995 10.6151
R4475 vdd.n2996 vdd.n779 10.6151
R4476 vdd.n3066 vdd.n779 10.6151
R4477 vdd.n3065 vdd.n3064 10.6151
R4478 vdd.n3064 vdd.n780 10.6151
R4479 vdd.n781 vdd.n780 10.6151
R4480 vdd.n3057 vdd.n781 10.6151
R4481 vdd.n3057 vdd.n3056 10.6151
R4482 vdd.n3056 vdd.n3055 10.6151
R4483 vdd.n3055 vdd.n783 10.6151
R4484 vdd.n3050 vdd.n783 10.6151
R4485 vdd.n3050 vdd.n3049 10.6151
R4486 vdd.n3049 vdd.n3048 10.6151
R4487 vdd.n3048 vdd.n786 10.6151
R4488 vdd.n3043 vdd.n786 10.6151
R4489 vdd.n3043 vdd.n3042 10.6151
R4490 vdd.n3042 vdd.n3041 10.6151
R4491 vdd.n3041 vdd.n789 10.6151
R4492 vdd.n3036 vdd.n789 10.6151
R4493 vdd.n3036 vdd.n3035 10.6151
R4494 vdd.n3035 vdd.n3033 10.6151
R4495 vdd.n3033 vdd.n792 10.6151
R4496 vdd.n3028 vdd.n792 10.6151
R4497 vdd.n3028 vdd.n3027 10.6151
R4498 vdd.n3027 vdd.n3026 10.6151
R4499 vdd.n3026 vdd.n795 10.6151
R4500 vdd.n3021 vdd.n795 10.6151
R4501 vdd.n3021 vdd.n3020 10.6151
R4502 vdd.n3020 vdd.n3019 10.6151
R4503 vdd.n3019 vdd.n798 10.6151
R4504 vdd.n3014 vdd.n798 10.6151
R4505 vdd.n3014 vdd.n3013 10.6151
R4506 vdd.n3013 vdd.n3012 10.6151
R4507 vdd.n3012 vdd.n801 10.6151
R4508 vdd.n3007 vdd.n3006 10.6151
R4509 vdd.n3006 vdd.n3005 10.6151
R4510 vdd.n2984 vdd.n2945 10.6151
R4511 vdd.n2979 vdd.n2945 10.6151
R4512 vdd.n2979 vdd.n2978 10.6151
R4513 vdd.n2978 vdd.n2977 10.6151
R4514 vdd.n2977 vdd.n2947 10.6151
R4515 vdd.n2972 vdd.n2947 10.6151
R4516 vdd.n2972 vdd.n2971 10.6151
R4517 vdd.n2971 vdd.n2970 10.6151
R4518 vdd.n2970 vdd.n2950 10.6151
R4519 vdd.n2965 vdd.n2950 10.6151
R4520 vdd.n2965 vdd.n2964 10.6151
R4521 vdd.n2964 vdd.n2963 10.6151
R4522 vdd.n2963 vdd.n2953 10.6151
R4523 vdd.n2958 vdd.n2953 10.6151
R4524 vdd.n2958 vdd.n2957 10.6151
R4525 vdd.n2957 vdd.n753 10.6151
R4526 vdd.n3101 vdd.n753 10.6151
R4527 vdd.n3101 vdd.n754 10.6151
R4528 vdd.n757 vdd.n754 10.6151
R4529 vdd.n3094 vdd.n757 10.6151
R4530 vdd.n3094 vdd.n3093 10.6151
R4531 vdd.n3093 vdd.n3092 10.6151
R4532 vdd.n3092 vdd.n759 10.6151
R4533 vdd.n3087 vdd.n759 10.6151
R4534 vdd.n3087 vdd.n3086 10.6151
R4535 vdd.n3086 vdd.n3085 10.6151
R4536 vdd.n3085 vdd.n762 10.6151
R4537 vdd.n3080 vdd.n762 10.6151
R4538 vdd.n3080 vdd.n3079 10.6151
R4539 vdd.n3079 vdd.n3078 10.6151
R4540 vdd.n3078 vdd.n765 10.6151
R4541 vdd.n3073 vdd.n3072 10.6151
R4542 vdd.n3072 vdd.n3071 10.6151
R4543 vdd.n2691 vdd.n2690 10.6151
R4544 vdd.n2777 vdd.n2691 10.6151
R4545 vdd.n2777 vdd.n2776 10.6151
R4546 vdd.n2776 vdd.n2775 10.6151
R4547 vdd.n2775 vdd.n2773 10.6151
R4548 vdd.n2773 vdd.n2772 10.6151
R4549 vdd.n2772 vdd.n2770 10.6151
R4550 vdd.n2770 vdd.n2769 10.6151
R4551 vdd.n2769 vdd.n2767 10.6151
R4552 vdd.n2767 vdd.n2766 10.6151
R4553 vdd.n2766 vdd.n2723 10.6151
R4554 vdd.n2723 vdd.n2722 10.6151
R4555 vdd.n2722 vdd.n2720 10.6151
R4556 vdd.n2720 vdd.n2719 10.6151
R4557 vdd.n2719 vdd.n2717 10.6151
R4558 vdd.n2717 vdd.n2716 10.6151
R4559 vdd.n2716 vdd.n2714 10.6151
R4560 vdd.n2714 vdd.n2713 10.6151
R4561 vdd.n2713 vdd.n2711 10.6151
R4562 vdd.n2711 vdd.n2710 10.6151
R4563 vdd.n2710 vdd.n2708 10.6151
R4564 vdd.n2708 vdd.n2707 10.6151
R4565 vdd.n2707 vdd.n2705 10.6151
R4566 vdd.n2705 vdd.n2704 10.6151
R4567 vdd.n2704 vdd.n2702 10.6151
R4568 vdd.n2702 vdd.n2701 10.6151
R4569 vdd.n2701 vdd.n2699 10.6151
R4570 vdd.n2699 vdd.n2698 10.6151
R4571 vdd.n2698 vdd.n2696 10.6151
R4572 vdd.n2696 vdd.n2695 10.6151
R4573 vdd.n2695 vdd.n2693 10.6151
R4574 vdd.n2693 vdd.n2692 10.6151
R4575 vdd.n2692 vdd.n771 10.6151
R4576 vdd.n2858 vdd.n903 10.6151
R4577 vdd.n2625 vdd.n903 10.6151
R4578 vdd.n2626 vdd.n2625 10.6151
R4579 vdd.n2629 vdd.n2626 10.6151
R4580 vdd.n2630 vdd.n2629 10.6151
R4581 vdd.n2633 vdd.n2630 10.6151
R4582 vdd.n2634 vdd.n2633 10.6151
R4583 vdd.n2637 vdd.n2634 10.6151
R4584 vdd.n2638 vdd.n2637 10.6151
R4585 vdd.n2641 vdd.n2638 10.6151
R4586 vdd.n2642 vdd.n2641 10.6151
R4587 vdd.n2645 vdd.n2642 10.6151
R4588 vdd.n2646 vdd.n2645 10.6151
R4589 vdd.n2649 vdd.n2646 10.6151
R4590 vdd.n2650 vdd.n2649 10.6151
R4591 vdd.n2653 vdd.n2650 10.6151
R4592 vdd.n2654 vdd.n2653 10.6151
R4593 vdd.n2657 vdd.n2654 10.6151
R4594 vdd.n2658 vdd.n2657 10.6151
R4595 vdd.n2661 vdd.n2658 10.6151
R4596 vdd.n2662 vdd.n2661 10.6151
R4597 vdd.n2665 vdd.n2662 10.6151
R4598 vdd.n2666 vdd.n2665 10.6151
R4599 vdd.n2669 vdd.n2666 10.6151
R4600 vdd.n2670 vdd.n2669 10.6151
R4601 vdd.n2673 vdd.n2670 10.6151
R4602 vdd.n2674 vdd.n2673 10.6151
R4603 vdd.n2677 vdd.n2674 10.6151
R4604 vdd.n2678 vdd.n2677 10.6151
R4605 vdd.n2681 vdd.n2678 10.6151
R4606 vdd.n2682 vdd.n2681 10.6151
R4607 vdd.n2687 vdd.n2685 10.6151
R4608 vdd.n2688 vdd.n2687 10.6151
R4609 vdd.n2860 vdd.n2859 10.6151
R4610 vdd.n2860 vdd.n892 10.6151
R4611 vdd.n2870 vdd.n892 10.6151
R4612 vdd.n2871 vdd.n2870 10.6151
R4613 vdd.n2872 vdd.n2871 10.6151
R4614 vdd.n2872 vdd.n880 10.6151
R4615 vdd.n2882 vdd.n880 10.6151
R4616 vdd.n2883 vdd.n2882 10.6151
R4617 vdd.n2884 vdd.n2883 10.6151
R4618 vdd.n2884 vdd.n868 10.6151
R4619 vdd.n2894 vdd.n868 10.6151
R4620 vdd.n2895 vdd.n2894 10.6151
R4621 vdd.n2896 vdd.n2895 10.6151
R4622 vdd.n2896 vdd.n857 10.6151
R4623 vdd.n2906 vdd.n857 10.6151
R4624 vdd.n2907 vdd.n2906 10.6151
R4625 vdd.n2908 vdd.n2907 10.6151
R4626 vdd.n2908 vdd.n844 10.6151
R4627 vdd.n2918 vdd.n844 10.6151
R4628 vdd.n2919 vdd.n2918 10.6151
R4629 vdd.n2921 vdd.n832 10.6151
R4630 vdd.n2931 vdd.n832 10.6151
R4631 vdd.n2932 vdd.n2931 10.6151
R4632 vdd.n2933 vdd.n2932 10.6151
R4633 vdd.n2933 vdd.n820 10.6151
R4634 vdd.n2943 vdd.n820 10.6151
R4635 vdd.n2944 vdd.n2943 10.6151
R4636 vdd.n2990 vdd.n2944 10.6151
R4637 vdd.n2990 vdd.n2989 10.6151
R4638 vdd.n2989 vdd.n2988 10.6151
R4639 vdd.n2988 vdd.n2987 10.6151
R4640 vdd.n2987 vdd.n2985 10.6151
R4641 vdd.n2339 vdd.n2338 10.6151
R4642 vdd.n2339 vdd.n1040 10.6151
R4643 vdd.n2349 vdd.n1040 10.6151
R4644 vdd.n2350 vdd.n2349 10.6151
R4645 vdd.n2351 vdd.n2350 10.6151
R4646 vdd.n2351 vdd.n1028 10.6151
R4647 vdd.n2361 vdd.n1028 10.6151
R4648 vdd.n2362 vdd.n2361 10.6151
R4649 vdd.n2363 vdd.n2362 10.6151
R4650 vdd.n2363 vdd.n1015 10.6151
R4651 vdd.n2373 vdd.n1015 10.6151
R4652 vdd.n2374 vdd.n2373 10.6151
R4653 vdd.n2376 vdd.n1003 10.6151
R4654 vdd.n2386 vdd.n1003 10.6151
R4655 vdd.n2387 vdd.n2386 10.6151
R4656 vdd.n2388 vdd.n2387 10.6151
R4657 vdd.n2388 vdd.n991 10.6151
R4658 vdd.n2398 vdd.n991 10.6151
R4659 vdd.n2399 vdd.n2398 10.6151
R4660 vdd.n2400 vdd.n2399 10.6151
R4661 vdd.n2400 vdd.n980 10.6151
R4662 vdd.n2410 vdd.n980 10.6151
R4663 vdd.n2411 vdd.n2410 10.6151
R4664 vdd.n2412 vdd.n2411 10.6151
R4665 vdd.n2412 vdd.n968 10.6151
R4666 vdd.n2422 vdd.n968 10.6151
R4667 vdd.n2423 vdd.n2422 10.6151
R4668 vdd.n2426 vdd.n2423 10.6151
R4669 vdd.n2426 vdd.n2425 10.6151
R4670 vdd.n2425 vdd.n2424 10.6151
R4671 vdd.n2424 vdd.n951 10.6151
R4672 vdd.n2508 vdd.n951 10.6151
R4673 vdd.n2507 vdd.n2506 10.6151
R4674 vdd.n2506 vdd.n2503 10.6151
R4675 vdd.n2503 vdd.n2502 10.6151
R4676 vdd.n2502 vdd.n2499 10.6151
R4677 vdd.n2499 vdd.n2498 10.6151
R4678 vdd.n2498 vdd.n2495 10.6151
R4679 vdd.n2495 vdd.n2494 10.6151
R4680 vdd.n2494 vdd.n2491 10.6151
R4681 vdd.n2491 vdd.n2490 10.6151
R4682 vdd.n2490 vdd.n2487 10.6151
R4683 vdd.n2487 vdd.n2486 10.6151
R4684 vdd.n2486 vdd.n2483 10.6151
R4685 vdd.n2483 vdd.n2482 10.6151
R4686 vdd.n2482 vdd.n2479 10.6151
R4687 vdd.n2479 vdd.n2478 10.6151
R4688 vdd.n2478 vdd.n2475 10.6151
R4689 vdd.n2475 vdd.n2474 10.6151
R4690 vdd.n2474 vdd.n2471 10.6151
R4691 vdd.n2471 vdd.n2470 10.6151
R4692 vdd.n2470 vdd.n2467 10.6151
R4693 vdd.n2467 vdd.n2466 10.6151
R4694 vdd.n2466 vdd.n2463 10.6151
R4695 vdd.n2463 vdd.n2462 10.6151
R4696 vdd.n2462 vdd.n2459 10.6151
R4697 vdd.n2459 vdd.n2458 10.6151
R4698 vdd.n2458 vdd.n2455 10.6151
R4699 vdd.n2455 vdd.n2454 10.6151
R4700 vdd.n2454 vdd.n2451 10.6151
R4701 vdd.n2451 vdd.n2450 10.6151
R4702 vdd.n2450 vdd.n2447 10.6151
R4703 vdd.n2447 vdd.n2446 10.6151
R4704 vdd.n2443 vdd.n2442 10.6151
R4705 vdd.n2442 vdd.n2440 10.6151
R4706 vdd.n1359 vdd.n1357 10.6151
R4707 vdd.n1357 vdd.n1356 10.6151
R4708 vdd.n1356 vdd.n1354 10.6151
R4709 vdd.n1354 vdd.n1353 10.6151
R4710 vdd.n1353 vdd.n1351 10.6151
R4711 vdd.n1351 vdd.n1350 10.6151
R4712 vdd.n1350 vdd.n1348 10.6151
R4713 vdd.n1348 vdd.n1347 10.6151
R4714 vdd.n1347 vdd.n1345 10.6151
R4715 vdd.n1345 vdd.n1344 10.6151
R4716 vdd.n1344 vdd.n1342 10.6151
R4717 vdd.n1342 vdd.n1341 10.6151
R4718 vdd.n1341 vdd.n1339 10.6151
R4719 vdd.n1339 vdd.n1338 10.6151
R4720 vdd.n1338 vdd.n1336 10.6151
R4721 vdd.n1336 vdd.n1335 10.6151
R4722 vdd.n1335 vdd.n1333 10.6151
R4723 vdd.n1333 vdd.n1332 10.6151
R4724 vdd.n1332 vdd.n1243 10.6151
R4725 vdd.n1243 vdd.n1242 10.6151
R4726 vdd.n1242 vdd.n1240 10.6151
R4727 vdd.n1240 vdd.n1239 10.6151
R4728 vdd.n1239 vdd.n1237 10.6151
R4729 vdd.n1237 vdd.n1236 10.6151
R4730 vdd.n1236 vdd.n1234 10.6151
R4731 vdd.n1234 vdd.n1233 10.6151
R4732 vdd.n1233 vdd.n1231 10.6151
R4733 vdd.n1231 vdd.n1230 10.6151
R4734 vdd.n1230 vdd.n1228 10.6151
R4735 vdd.n1228 vdd.n1227 10.6151
R4736 vdd.n1227 vdd.n955 10.6151
R4737 vdd.n2438 vdd.n955 10.6151
R4738 vdd.n2439 vdd.n2438 10.6151
R4739 vdd.n2337 vdd.n1052 10.6151
R4740 vdd.n1194 vdd.n1052 10.6151
R4741 vdd.n1195 vdd.n1194 10.6151
R4742 vdd.n1198 vdd.n1195 10.6151
R4743 vdd.n1199 vdd.n1198 10.6151
R4744 vdd.n1202 vdd.n1199 10.6151
R4745 vdd.n1203 vdd.n1202 10.6151
R4746 vdd.n1206 vdd.n1203 10.6151
R4747 vdd.n1207 vdd.n1206 10.6151
R4748 vdd.n1210 vdd.n1207 10.6151
R4749 vdd.n1211 vdd.n1210 10.6151
R4750 vdd.n1214 vdd.n1211 10.6151
R4751 vdd.n1215 vdd.n1214 10.6151
R4752 vdd.n1218 vdd.n1215 10.6151
R4753 vdd.n1219 vdd.n1218 10.6151
R4754 vdd.n1222 vdd.n1219 10.6151
R4755 vdd.n1393 vdd.n1222 10.6151
R4756 vdd.n1393 vdd.n1392 10.6151
R4757 vdd.n1392 vdd.n1390 10.6151
R4758 vdd.n1390 vdd.n1387 10.6151
R4759 vdd.n1387 vdd.n1386 10.6151
R4760 vdd.n1386 vdd.n1383 10.6151
R4761 vdd.n1383 vdd.n1382 10.6151
R4762 vdd.n1382 vdd.n1379 10.6151
R4763 vdd.n1379 vdd.n1378 10.6151
R4764 vdd.n1378 vdd.n1375 10.6151
R4765 vdd.n1375 vdd.n1374 10.6151
R4766 vdd.n1374 vdd.n1371 10.6151
R4767 vdd.n1371 vdd.n1370 10.6151
R4768 vdd.n1370 vdd.n1367 10.6151
R4769 vdd.n1367 vdd.n1366 10.6151
R4770 vdd.n1363 vdd.n1362 10.6151
R4771 vdd.n1362 vdd.n1360 10.6151
R4772 vdd.t233 vdd.n2138 10.5435
R4773 vdd.n636 vdd.t187 10.5435
R4774 vdd.n304 vdd.n286 10.4732
R4775 vdd.n249 vdd.n231 10.4732
R4776 vdd.n206 vdd.n188 10.4732
R4777 vdd.n151 vdd.n133 10.4732
R4778 vdd.n109 vdd.n91 10.4732
R4779 vdd.n54 vdd.n36 10.4732
R4780 vdd.n2035 vdd.n2017 10.4732
R4781 vdd.n2090 vdd.n2072 10.4732
R4782 vdd.n1937 vdd.n1919 10.4732
R4783 vdd.n1992 vdd.n1974 10.4732
R4784 vdd.n1840 vdd.n1822 10.4732
R4785 vdd.n1895 vdd.n1877 10.4732
R4786 vdd.n2122 vdd.t194 10.3167
R4787 vdd.n3297 vdd.t184 10.3167
R4788 vdd.t215 vdd.n1466 10.09
R4789 vdd.n2174 vdd.t63 10.09
R4790 vdd.n3245 vdd.t59 10.09
R4791 vdd.n3378 vdd.t182 10.09
R4792 vdd.n1786 vdd.t170 9.86327
R4793 vdd.n3369 vdd.t230 9.86327
R4794 vdd.n2299 vdd.n2298 9.78206
R4795 vdd.n3035 vdd.n3034 9.78206
R4796 vdd.n3102 vdd.n3101 9.78206
R4797 vdd.n2191 vdd.n1393 9.78206
R4798 vdd.n303 vdd.n288 9.69747
R4799 vdd.n248 vdd.n233 9.69747
R4800 vdd.n205 vdd.n190 9.69747
R4801 vdd.n150 vdd.n135 9.69747
R4802 vdd.n108 vdd.n93 9.69747
R4803 vdd.n53 vdd.n38 9.69747
R4804 vdd.n2034 vdd.n2019 9.69747
R4805 vdd.n2089 vdd.n2074 9.69747
R4806 vdd.n1936 vdd.n1921 9.69747
R4807 vdd.n1991 vdd.n1976 9.69747
R4808 vdd.n1839 vdd.n1824 9.69747
R4809 vdd.n1894 vdd.n1879 9.69747
R4810 vdd.t144 vdd.n1760 9.63654
R4811 vdd.n3328 vdd.t196 9.63654
R4812 vdd.n319 vdd.n318 9.45567
R4813 vdd.n264 vdd.n263 9.45567
R4814 vdd.n221 vdd.n220 9.45567
R4815 vdd.n166 vdd.n165 9.45567
R4816 vdd.n124 vdd.n123 9.45567
R4817 vdd.n69 vdd.n68 9.45567
R4818 vdd.n2050 vdd.n2049 9.45567
R4819 vdd.n2105 vdd.n2104 9.45567
R4820 vdd.n1952 vdd.n1951 9.45567
R4821 vdd.n2007 vdd.n2006 9.45567
R4822 vdd.n1855 vdd.n1854 9.45567
R4823 vdd.n1910 vdd.n1909 9.45567
R4824 vdd.n2261 vdd.n1120 9.3005
R4825 vdd.n2260 vdd.n2259 9.3005
R4826 vdd.n1126 vdd.n1125 9.3005
R4827 vdd.n2254 vdd.n1130 9.3005
R4828 vdd.n2253 vdd.n1131 9.3005
R4829 vdd.n2252 vdd.n1132 9.3005
R4830 vdd.n1136 vdd.n1133 9.3005
R4831 vdd.n2247 vdd.n1137 9.3005
R4832 vdd.n2246 vdd.n1138 9.3005
R4833 vdd.n2245 vdd.n1139 9.3005
R4834 vdd.n1143 vdd.n1140 9.3005
R4835 vdd.n2240 vdd.n1144 9.3005
R4836 vdd.n2239 vdd.n1145 9.3005
R4837 vdd.n2238 vdd.n1146 9.3005
R4838 vdd.n1150 vdd.n1147 9.3005
R4839 vdd.n2233 vdd.n1151 9.3005
R4840 vdd.n2232 vdd.n1152 9.3005
R4841 vdd.n2231 vdd.n1153 9.3005
R4842 vdd.n1157 vdd.n1154 9.3005
R4843 vdd.n2226 vdd.n1158 9.3005
R4844 vdd.n2225 vdd.n1159 9.3005
R4845 vdd.n2224 vdd.n2223 9.3005
R4846 vdd.n2222 vdd.n1160 9.3005
R4847 vdd.n2221 vdd.n2220 9.3005
R4848 vdd.n1166 vdd.n1165 9.3005
R4849 vdd.n2215 vdd.n1170 9.3005
R4850 vdd.n2214 vdd.n1171 9.3005
R4851 vdd.n2213 vdd.n1172 9.3005
R4852 vdd.n1176 vdd.n1173 9.3005
R4853 vdd.n2208 vdd.n1177 9.3005
R4854 vdd.n2207 vdd.n1178 9.3005
R4855 vdd.n2206 vdd.n1179 9.3005
R4856 vdd.n1183 vdd.n1180 9.3005
R4857 vdd.n2201 vdd.n1184 9.3005
R4858 vdd.n2200 vdd.n1185 9.3005
R4859 vdd.n2199 vdd.n1186 9.3005
R4860 vdd.n1190 vdd.n1187 9.3005
R4861 vdd.n2194 vdd.n1191 9.3005
R4862 vdd.n2263 vdd.n2262 9.3005
R4863 vdd.n2285 vdd.n1091 9.3005
R4864 vdd.n2284 vdd.n1099 9.3005
R4865 vdd.n1103 vdd.n1100 9.3005
R4866 vdd.n2279 vdd.n1104 9.3005
R4867 vdd.n2278 vdd.n1105 9.3005
R4868 vdd.n2277 vdd.n1106 9.3005
R4869 vdd.n1110 vdd.n1107 9.3005
R4870 vdd.n2272 vdd.n1111 9.3005
R4871 vdd.n2271 vdd.n1112 9.3005
R4872 vdd.n2270 vdd.n1113 9.3005
R4873 vdd.n1117 vdd.n1114 9.3005
R4874 vdd.n2265 vdd.n1118 9.3005
R4875 vdd.n2264 vdd.n1119 9.3005
R4876 vdd.n2297 vdd.n2296 9.3005
R4877 vdd.n1095 vdd.n1094 9.3005
R4878 vdd.n2110 vdd.n1456 9.3005
R4879 vdd.n2112 vdd.n2111 9.3005
R4880 vdd.n1447 vdd.n1446 9.3005
R4881 vdd.n2125 vdd.n2124 9.3005
R4882 vdd.n2126 vdd.n1445 9.3005
R4883 vdd.n2128 vdd.n2127 9.3005
R4884 vdd.n1435 vdd.n1434 9.3005
R4885 vdd.n2142 vdd.n2141 9.3005
R4886 vdd.n2143 vdd.n1433 9.3005
R4887 vdd.n2145 vdd.n2144 9.3005
R4888 vdd.n1424 vdd.n1423 9.3005
R4889 vdd.n2159 vdd.n2158 9.3005
R4890 vdd.n2160 vdd.n1422 9.3005
R4891 vdd.n2162 vdd.n2161 9.3005
R4892 vdd.n1412 vdd.n1411 9.3005
R4893 vdd.n2177 vdd.n2176 9.3005
R4894 vdd.n2178 vdd.n1410 9.3005
R4895 vdd.n2180 vdd.n2179 9.3005
R4896 vdd.n295 vdd.n294 9.3005
R4897 vdd.n290 vdd.n289 9.3005
R4898 vdd.n301 vdd.n300 9.3005
R4899 vdd.n303 vdd.n302 9.3005
R4900 vdd.n286 vdd.n285 9.3005
R4901 vdd.n309 vdd.n308 9.3005
R4902 vdd.n311 vdd.n310 9.3005
R4903 vdd.n283 vdd.n280 9.3005
R4904 vdd.n318 vdd.n317 9.3005
R4905 vdd.n240 vdd.n239 9.3005
R4906 vdd.n235 vdd.n234 9.3005
R4907 vdd.n246 vdd.n245 9.3005
R4908 vdd.n248 vdd.n247 9.3005
R4909 vdd.n231 vdd.n230 9.3005
R4910 vdd.n254 vdd.n253 9.3005
R4911 vdd.n256 vdd.n255 9.3005
R4912 vdd.n228 vdd.n225 9.3005
R4913 vdd.n263 vdd.n262 9.3005
R4914 vdd.n197 vdd.n196 9.3005
R4915 vdd.n192 vdd.n191 9.3005
R4916 vdd.n203 vdd.n202 9.3005
R4917 vdd.n205 vdd.n204 9.3005
R4918 vdd.n188 vdd.n187 9.3005
R4919 vdd.n211 vdd.n210 9.3005
R4920 vdd.n213 vdd.n212 9.3005
R4921 vdd.n185 vdd.n182 9.3005
R4922 vdd.n220 vdd.n219 9.3005
R4923 vdd.n142 vdd.n141 9.3005
R4924 vdd.n137 vdd.n136 9.3005
R4925 vdd.n148 vdd.n147 9.3005
R4926 vdd.n150 vdd.n149 9.3005
R4927 vdd.n133 vdd.n132 9.3005
R4928 vdd.n156 vdd.n155 9.3005
R4929 vdd.n158 vdd.n157 9.3005
R4930 vdd.n130 vdd.n127 9.3005
R4931 vdd.n165 vdd.n164 9.3005
R4932 vdd.n100 vdd.n99 9.3005
R4933 vdd.n95 vdd.n94 9.3005
R4934 vdd.n106 vdd.n105 9.3005
R4935 vdd.n108 vdd.n107 9.3005
R4936 vdd.n91 vdd.n90 9.3005
R4937 vdd.n114 vdd.n113 9.3005
R4938 vdd.n116 vdd.n115 9.3005
R4939 vdd.n88 vdd.n85 9.3005
R4940 vdd.n123 vdd.n122 9.3005
R4941 vdd.n45 vdd.n44 9.3005
R4942 vdd.n40 vdd.n39 9.3005
R4943 vdd.n51 vdd.n50 9.3005
R4944 vdd.n53 vdd.n52 9.3005
R4945 vdd.n36 vdd.n35 9.3005
R4946 vdd.n59 vdd.n58 9.3005
R4947 vdd.n61 vdd.n60 9.3005
R4948 vdd.n33 vdd.n30 9.3005
R4949 vdd.n68 vdd.n67 9.3005
R4950 vdd.n3151 vdd.n3150 9.3005
R4951 vdd.n3152 vdd.n721 9.3005
R4952 vdd.n720 vdd.n718 9.3005
R4953 vdd.n3158 vdd.n717 9.3005
R4954 vdd.n3159 vdd.n716 9.3005
R4955 vdd.n3160 vdd.n715 9.3005
R4956 vdd.n714 vdd.n712 9.3005
R4957 vdd.n3166 vdd.n711 9.3005
R4958 vdd.n3167 vdd.n710 9.3005
R4959 vdd.n3168 vdd.n709 9.3005
R4960 vdd.n708 vdd.n706 9.3005
R4961 vdd.n3174 vdd.n705 9.3005
R4962 vdd.n3175 vdd.n704 9.3005
R4963 vdd.n3176 vdd.n703 9.3005
R4964 vdd.n702 vdd.n700 9.3005
R4965 vdd.n3182 vdd.n699 9.3005
R4966 vdd.n3183 vdd.n698 9.3005
R4967 vdd.n3184 vdd.n697 9.3005
R4968 vdd.n696 vdd.n694 9.3005
R4969 vdd.n3190 vdd.n693 9.3005
R4970 vdd.n3191 vdd.n692 9.3005
R4971 vdd.n3192 vdd.n691 9.3005
R4972 vdd.n690 vdd.n688 9.3005
R4973 vdd.n3198 vdd.n685 9.3005
R4974 vdd.n3199 vdd.n684 9.3005
R4975 vdd.n3200 vdd.n683 9.3005
R4976 vdd.n682 vdd.n680 9.3005
R4977 vdd.n3206 vdd.n679 9.3005
R4978 vdd.n3207 vdd.n678 9.3005
R4979 vdd.n3208 vdd.n677 9.3005
R4980 vdd.n676 vdd.n674 9.3005
R4981 vdd.n3214 vdd.n673 9.3005
R4982 vdd.n3215 vdd.n672 9.3005
R4983 vdd.n3216 vdd.n671 9.3005
R4984 vdd.n670 vdd.n668 9.3005
R4985 vdd.n3221 vdd.n667 9.3005
R4986 vdd.n3231 vdd.n661 9.3005
R4987 vdd.n3233 vdd.n3232 9.3005
R4988 vdd.n652 vdd.n651 9.3005
R4989 vdd.n3248 vdd.n3247 9.3005
R4990 vdd.n3249 vdd.n650 9.3005
R4991 vdd.n3251 vdd.n3250 9.3005
R4992 vdd.n640 vdd.n639 9.3005
R4993 vdd.n3264 vdd.n3263 9.3005
R4994 vdd.n3265 vdd.n638 9.3005
R4995 vdd.n3267 vdd.n3266 9.3005
R4996 vdd.n628 vdd.n627 9.3005
R4997 vdd.n3281 vdd.n3280 9.3005
R4998 vdd.n3282 vdd.n626 9.3005
R4999 vdd.n3284 vdd.n3283 9.3005
R5000 vdd.n617 vdd.n616 9.3005
R5001 vdd.n3300 vdd.n3299 9.3005
R5002 vdd.n3301 vdd.n615 9.3005
R5003 vdd.n3303 vdd.n3302 9.3005
R5004 vdd.n324 vdd.n322 9.3005
R5005 vdd.n3235 vdd.n3234 9.3005
R5006 vdd.n3382 vdd.n3381 9.3005
R5007 vdd.n325 vdd.n323 9.3005
R5008 vdd.n3375 vdd.n334 9.3005
R5009 vdd.n3374 vdd.n335 9.3005
R5010 vdd.n3373 vdd.n336 9.3005
R5011 vdd.n343 vdd.n337 9.3005
R5012 vdd.n3367 vdd.n344 9.3005
R5013 vdd.n3366 vdd.n345 9.3005
R5014 vdd.n3365 vdd.n346 9.3005
R5015 vdd.n354 vdd.n347 9.3005
R5016 vdd.n3359 vdd.n355 9.3005
R5017 vdd.n3358 vdd.n356 9.3005
R5018 vdd.n3357 vdd.n357 9.3005
R5019 vdd.n365 vdd.n358 9.3005
R5020 vdd.n3351 vdd.n366 9.3005
R5021 vdd.n3350 vdd.n367 9.3005
R5022 vdd.n3349 vdd.n368 9.3005
R5023 vdd.n443 vdd.n369 9.3005
R5024 vdd.n447 vdd.n442 9.3005
R5025 vdd.n451 vdd.n450 9.3005
R5026 vdd.n452 vdd.n441 9.3005
R5027 vdd.n456 vdd.n453 9.3005
R5028 vdd.n457 vdd.n440 9.3005
R5029 vdd.n461 vdd.n460 9.3005
R5030 vdd.n462 vdd.n439 9.3005
R5031 vdd.n466 vdd.n463 9.3005
R5032 vdd.n467 vdd.n438 9.3005
R5033 vdd.n471 vdd.n470 9.3005
R5034 vdd.n472 vdd.n437 9.3005
R5035 vdd.n476 vdd.n473 9.3005
R5036 vdd.n477 vdd.n436 9.3005
R5037 vdd.n481 vdd.n480 9.3005
R5038 vdd.n482 vdd.n435 9.3005
R5039 vdd.n486 vdd.n483 9.3005
R5040 vdd.n487 vdd.n434 9.3005
R5041 vdd.n491 vdd.n490 9.3005
R5042 vdd.n492 vdd.n433 9.3005
R5043 vdd.n496 vdd.n493 9.3005
R5044 vdd.n497 vdd.n430 9.3005
R5045 vdd.n501 vdd.n500 9.3005
R5046 vdd.n502 vdd.n429 9.3005
R5047 vdd.n506 vdd.n503 9.3005
R5048 vdd.n507 vdd.n428 9.3005
R5049 vdd.n511 vdd.n510 9.3005
R5050 vdd.n512 vdd.n427 9.3005
R5051 vdd.n516 vdd.n513 9.3005
R5052 vdd.n517 vdd.n426 9.3005
R5053 vdd.n521 vdd.n520 9.3005
R5054 vdd.n522 vdd.n425 9.3005
R5055 vdd.n526 vdd.n523 9.3005
R5056 vdd.n527 vdd.n424 9.3005
R5057 vdd.n531 vdd.n530 9.3005
R5058 vdd.n532 vdd.n423 9.3005
R5059 vdd.n536 vdd.n533 9.3005
R5060 vdd.n537 vdd.n422 9.3005
R5061 vdd.n541 vdd.n540 9.3005
R5062 vdd.n542 vdd.n421 9.3005
R5063 vdd.n546 vdd.n543 9.3005
R5064 vdd.n547 vdd.n418 9.3005
R5065 vdd.n551 vdd.n550 9.3005
R5066 vdd.n552 vdd.n417 9.3005
R5067 vdd.n556 vdd.n553 9.3005
R5068 vdd.n557 vdd.n416 9.3005
R5069 vdd.n561 vdd.n560 9.3005
R5070 vdd.n562 vdd.n415 9.3005
R5071 vdd.n566 vdd.n563 9.3005
R5072 vdd.n567 vdd.n414 9.3005
R5073 vdd.n571 vdd.n570 9.3005
R5074 vdd.n572 vdd.n413 9.3005
R5075 vdd.n576 vdd.n573 9.3005
R5076 vdd.n577 vdd.n412 9.3005
R5077 vdd.n581 vdd.n580 9.3005
R5078 vdd.n582 vdd.n411 9.3005
R5079 vdd.n586 vdd.n583 9.3005
R5080 vdd.n587 vdd.n410 9.3005
R5081 vdd.n591 vdd.n590 9.3005
R5082 vdd.n592 vdd.n409 9.3005
R5083 vdd.n596 vdd.n593 9.3005
R5084 vdd.n598 vdd.n408 9.3005
R5085 vdd.n600 vdd.n599 9.3005
R5086 vdd.n3342 vdd.n3341 9.3005
R5087 vdd.n446 vdd.n444 9.3005
R5088 vdd.n3241 vdd.n655 9.3005
R5089 vdd.n3243 vdd.n3242 9.3005
R5090 vdd.n646 vdd.n645 9.3005
R5091 vdd.n3256 vdd.n3255 9.3005
R5092 vdd.n3257 vdd.n644 9.3005
R5093 vdd.n3259 vdd.n3258 9.3005
R5094 vdd.n633 vdd.n632 9.3005
R5095 vdd.n3272 vdd.n3271 9.3005
R5096 vdd.n3273 vdd.n631 9.3005
R5097 vdd.n3275 vdd.n3274 9.3005
R5098 vdd.n622 vdd.n621 9.3005
R5099 vdd.n3289 vdd.n3288 9.3005
R5100 vdd.n3290 vdd.n620 9.3005
R5101 vdd.n3295 vdd.n3291 9.3005
R5102 vdd.n3294 vdd.n3293 9.3005
R5103 vdd.n3292 vdd.n610 9.3005
R5104 vdd.n3308 vdd.n611 9.3005
R5105 vdd.n3309 vdd.n609 9.3005
R5106 vdd.n3311 vdd.n3310 9.3005
R5107 vdd.n3312 vdd.n608 9.3005
R5108 vdd.n3315 vdd.n3313 9.3005
R5109 vdd.n3316 vdd.n607 9.3005
R5110 vdd.n3318 vdd.n3317 9.3005
R5111 vdd.n3319 vdd.n606 9.3005
R5112 vdd.n3322 vdd.n3320 9.3005
R5113 vdd.n3323 vdd.n605 9.3005
R5114 vdd.n3325 vdd.n3324 9.3005
R5115 vdd.n3326 vdd.n604 9.3005
R5116 vdd.n3330 vdd.n3327 9.3005
R5117 vdd.n3331 vdd.n603 9.3005
R5118 vdd.n3333 vdd.n3332 9.3005
R5119 vdd.n3334 vdd.n602 9.3005
R5120 vdd.n3337 vdd.n3335 9.3005
R5121 vdd.n3338 vdd.n601 9.3005
R5122 vdd.n3340 vdd.n3339 9.3005
R5123 vdd.n3240 vdd.n3239 9.3005
R5124 vdd.n3104 vdd.n656 9.3005
R5125 vdd.n3109 vdd.n3103 9.3005
R5126 vdd.n3119 vdd.n748 9.3005
R5127 vdd.n3120 vdd.n747 9.3005
R5128 vdd.n746 vdd.n744 9.3005
R5129 vdd.n3126 vdd.n743 9.3005
R5130 vdd.n3127 vdd.n742 9.3005
R5131 vdd.n3128 vdd.n741 9.3005
R5132 vdd.n740 vdd.n738 9.3005
R5133 vdd.n3134 vdd.n737 9.3005
R5134 vdd.n3135 vdd.n736 9.3005
R5135 vdd.n3136 vdd.n735 9.3005
R5136 vdd.n734 vdd.n732 9.3005
R5137 vdd.n3141 vdd.n731 9.3005
R5138 vdd.n3142 vdd.n730 9.3005
R5139 vdd.n726 vdd.n725 9.3005
R5140 vdd.n3148 vdd.n3147 9.3005
R5141 vdd.n3149 vdd.n722 9.3005
R5142 vdd.n2190 vdd.n2189 9.3005
R5143 vdd.n2185 vdd.n1395 9.3005
R5144 vdd.n1742 vdd.n1741 9.3005
R5145 vdd.n1498 vdd.n1497 9.3005
R5146 vdd.n1755 vdd.n1754 9.3005
R5147 vdd.n1756 vdd.n1496 9.3005
R5148 vdd.n1758 vdd.n1757 9.3005
R5149 vdd.n1486 vdd.n1485 9.3005
R5150 vdd.n1772 vdd.n1771 9.3005
R5151 vdd.n1773 vdd.n1484 9.3005
R5152 vdd.n1775 vdd.n1774 9.3005
R5153 vdd.n1476 vdd.n1475 9.3005
R5154 vdd.n1789 vdd.n1788 9.3005
R5155 vdd.n1790 vdd.n1474 9.3005
R5156 vdd.n1792 vdd.n1791 9.3005
R5157 vdd.n1463 vdd.n1462 9.3005
R5158 vdd.n1805 vdd.n1804 9.3005
R5159 vdd.n1806 vdd.n1461 9.3005
R5160 vdd.n1808 vdd.n1807 9.3005
R5161 vdd.n1452 vdd.n1451 9.3005
R5162 vdd.n2117 vdd.n2116 9.3005
R5163 vdd.n2118 vdd.n1450 9.3005
R5164 vdd.n2120 vdd.n2119 9.3005
R5165 vdd.n1441 vdd.n1440 9.3005
R5166 vdd.n2133 vdd.n2132 9.3005
R5167 vdd.n2134 vdd.n1439 9.3005
R5168 vdd.n2136 vdd.n2135 9.3005
R5169 vdd.n1429 vdd.n1428 9.3005
R5170 vdd.n2150 vdd.n2149 9.3005
R5171 vdd.n2151 vdd.n1427 9.3005
R5172 vdd.n2153 vdd.n2152 9.3005
R5173 vdd.n1419 vdd.n1418 9.3005
R5174 vdd.n2167 vdd.n2166 9.3005
R5175 vdd.n2168 vdd.n1416 9.3005
R5176 vdd.n2172 vdd.n2171 9.3005
R5177 vdd.n2170 vdd.n1417 9.3005
R5178 vdd.n2169 vdd.n1406 9.3005
R5179 vdd.n1740 vdd.n1508 9.3005
R5180 vdd.n1633 vdd.n1509 9.3005
R5181 vdd.n1635 vdd.n1634 9.3005
R5182 vdd.n1636 vdd.n1628 9.3005
R5183 vdd.n1638 vdd.n1637 9.3005
R5184 vdd.n1639 vdd.n1627 9.3005
R5185 vdd.n1641 vdd.n1640 9.3005
R5186 vdd.n1642 vdd.n1622 9.3005
R5187 vdd.n1644 vdd.n1643 9.3005
R5188 vdd.n1645 vdd.n1621 9.3005
R5189 vdd.n1647 vdd.n1646 9.3005
R5190 vdd.n1648 vdd.n1616 9.3005
R5191 vdd.n1650 vdd.n1649 9.3005
R5192 vdd.n1651 vdd.n1615 9.3005
R5193 vdd.n1653 vdd.n1652 9.3005
R5194 vdd.n1654 vdd.n1610 9.3005
R5195 vdd.n1656 vdd.n1655 9.3005
R5196 vdd.n1657 vdd.n1609 9.3005
R5197 vdd.n1659 vdd.n1658 9.3005
R5198 vdd.n1660 vdd.n1604 9.3005
R5199 vdd.n1662 vdd.n1661 9.3005
R5200 vdd.n1663 vdd.n1603 9.3005
R5201 vdd.n1668 vdd.n1664 9.3005
R5202 vdd.n1669 vdd.n1599 9.3005
R5203 vdd.n1671 vdd.n1670 9.3005
R5204 vdd.n1672 vdd.n1598 9.3005
R5205 vdd.n1674 vdd.n1673 9.3005
R5206 vdd.n1675 vdd.n1593 9.3005
R5207 vdd.n1677 vdd.n1676 9.3005
R5208 vdd.n1678 vdd.n1592 9.3005
R5209 vdd.n1680 vdd.n1679 9.3005
R5210 vdd.n1681 vdd.n1587 9.3005
R5211 vdd.n1683 vdd.n1682 9.3005
R5212 vdd.n1684 vdd.n1586 9.3005
R5213 vdd.n1686 vdd.n1685 9.3005
R5214 vdd.n1687 vdd.n1581 9.3005
R5215 vdd.n1689 vdd.n1688 9.3005
R5216 vdd.n1690 vdd.n1580 9.3005
R5217 vdd.n1692 vdd.n1691 9.3005
R5218 vdd.n1693 vdd.n1575 9.3005
R5219 vdd.n1695 vdd.n1694 9.3005
R5220 vdd.n1696 vdd.n1574 9.3005
R5221 vdd.n1698 vdd.n1697 9.3005
R5222 vdd.n1699 vdd.n1571 9.3005
R5223 vdd.n1705 vdd.n1704 9.3005
R5224 vdd.n1706 vdd.n1570 9.3005
R5225 vdd.n1708 vdd.n1707 9.3005
R5226 vdd.n1709 vdd.n1565 9.3005
R5227 vdd.n1711 vdd.n1710 9.3005
R5228 vdd.n1712 vdd.n1564 9.3005
R5229 vdd.n1714 vdd.n1713 9.3005
R5230 vdd.n1715 vdd.n1559 9.3005
R5231 vdd.n1717 vdd.n1716 9.3005
R5232 vdd.n1718 vdd.n1558 9.3005
R5233 vdd.n1720 vdd.n1719 9.3005
R5234 vdd.n1721 vdd.n1553 9.3005
R5235 vdd.n1723 vdd.n1722 9.3005
R5236 vdd.n1724 vdd.n1552 9.3005
R5237 vdd.n1726 vdd.n1725 9.3005
R5238 vdd.n1727 vdd.n1548 9.3005
R5239 vdd.n1729 vdd.n1728 9.3005
R5240 vdd.n1730 vdd.n1547 9.3005
R5241 vdd.n1732 vdd.n1731 9.3005
R5242 vdd.n1733 vdd.n1546 9.3005
R5243 vdd.n1739 vdd.n1738 9.3005
R5244 vdd.n1747 vdd.n1746 9.3005
R5245 vdd.n1748 vdd.n1502 9.3005
R5246 vdd.n1750 vdd.n1749 9.3005
R5247 vdd.n1492 vdd.n1491 9.3005
R5248 vdd.n1764 vdd.n1763 9.3005
R5249 vdd.n1765 vdd.n1490 9.3005
R5250 vdd.n1767 vdd.n1766 9.3005
R5251 vdd.n1481 vdd.n1480 9.3005
R5252 vdd.n1781 vdd.n1780 9.3005
R5253 vdd.n1782 vdd.n1479 9.3005
R5254 vdd.n1784 vdd.n1783 9.3005
R5255 vdd.n1470 vdd.n1469 9.3005
R5256 vdd.n1797 vdd.n1796 9.3005
R5257 vdd.n1798 vdd.n1468 9.3005
R5258 vdd.n1800 vdd.n1799 9.3005
R5259 vdd.n1458 vdd.n1457 9.3005
R5260 vdd.n1814 vdd.n1813 9.3005
R5261 vdd.n1504 vdd.n1503 9.3005
R5262 vdd.n2026 vdd.n2025 9.3005
R5263 vdd.n2021 vdd.n2020 9.3005
R5264 vdd.n2032 vdd.n2031 9.3005
R5265 vdd.n2034 vdd.n2033 9.3005
R5266 vdd.n2017 vdd.n2016 9.3005
R5267 vdd.n2040 vdd.n2039 9.3005
R5268 vdd.n2042 vdd.n2041 9.3005
R5269 vdd.n2014 vdd.n2011 9.3005
R5270 vdd.n2049 vdd.n2048 9.3005
R5271 vdd.n2081 vdd.n2080 9.3005
R5272 vdd.n2076 vdd.n2075 9.3005
R5273 vdd.n2087 vdd.n2086 9.3005
R5274 vdd.n2089 vdd.n2088 9.3005
R5275 vdd.n2072 vdd.n2071 9.3005
R5276 vdd.n2095 vdd.n2094 9.3005
R5277 vdd.n2097 vdd.n2096 9.3005
R5278 vdd.n2069 vdd.n2066 9.3005
R5279 vdd.n2104 vdd.n2103 9.3005
R5280 vdd.n1928 vdd.n1927 9.3005
R5281 vdd.n1923 vdd.n1922 9.3005
R5282 vdd.n1934 vdd.n1933 9.3005
R5283 vdd.n1936 vdd.n1935 9.3005
R5284 vdd.n1919 vdd.n1918 9.3005
R5285 vdd.n1942 vdd.n1941 9.3005
R5286 vdd.n1944 vdd.n1943 9.3005
R5287 vdd.n1916 vdd.n1913 9.3005
R5288 vdd.n1951 vdd.n1950 9.3005
R5289 vdd.n1983 vdd.n1982 9.3005
R5290 vdd.n1978 vdd.n1977 9.3005
R5291 vdd.n1989 vdd.n1988 9.3005
R5292 vdd.n1991 vdd.n1990 9.3005
R5293 vdd.n1974 vdd.n1973 9.3005
R5294 vdd.n1997 vdd.n1996 9.3005
R5295 vdd.n1999 vdd.n1998 9.3005
R5296 vdd.n1971 vdd.n1968 9.3005
R5297 vdd.n2006 vdd.n2005 9.3005
R5298 vdd.n1831 vdd.n1830 9.3005
R5299 vdd.n1826 vdd.n1825 9.3005
R5300 vdd.n1837 vdd.n1836 9.3005
R5301 vdd.n1839 vdd.n1838 9.3005
R5302 vdd.n1822 vdd.n1821 9.3005
R5303 vdd.n1845 vdd.n1844 9.3005
R5304 vdd.n1847 vdd.n1846 9.3005
R5305 vdd.n1819 vdd.n1816 9.3005
R5306 vdd.n1854 vdd.n1853 9.3005
R5307 vdd.n1886 vdd.n1885 9.3005
R5308 vdd.n1881 vdd.n1880 9.3005
R5309 vdd.n1892 vdd.n1891 9.3005
R5310 vdd.n1894 vdd.n1893 9.3005
R5311 vdd.n1877 vdd.n1876 9.3005
R5312 vdd.n1900 vdd.n1899 9.3005
R5313 vdd.n1902 vdd.n1901 9.3005
R5314 vdd.n1874 vdd.n1871 9.3005
R5315 vdd.n1909 vdd.n1908 9.3005
R5316 vdd.n1760 vdd.t140 9.18308
R5317 vdd.n3328 vdd.t206 9.18308
R5318 vdd.n1786 vdd.t148 8.95635
R5319 vdd.t161 vdd.n3369 8.95635
R5320 vdd.n300 vdd.n299 8.92171
R5321 vdd.n245 vdd.n244 8.92171
R5322 vdd.n202 vdd.n201 8.92171
R5323 vdd.n147 vdd.n146 8.92171
R5324 vdd.n105 vdd.n104 8.92171
R5325 vdd.n50 vdd.n49 8.92171
R5326 vdd.n2031 vdd.n2030 8.92171
R5327 vdd.n2086 vdd.n2085 8.92171
R5328 vdd.n1933 vdd.n1932 8.92171
R5329 vdd.n1988 vdd.n1987 8.92171
R5330 vdd.n1836 vdd.n1835 8.92171
R5331 vdd.n1891 vdd.n1890 8.92171
R5332 vdd.n223 vdd.n125 8.81535
R5333 vdd.n2009 vdd.n1911 8.81535
R5334 vdd.n1466 vdd.t174 8.72962
R5335 vdd.t211 vdd.n3378 8.72962
R5336 vdd.n2122 vdd.t150 8.50289
R5337 vdd.n3297 vdd.t146 8.50289
R5338 vdd.n28 vdd.n14 8.42249
R5339 vdd.n2138 vdd.t203 8.27616
R5340 vdd.t138 vdd.n636 8.27616
R5341 vdd.n3384 vdd.n3383 8.16225
R5342 vdd.n2109 vdd.n2108 8.16225
R5343 vdd.n296 vdd.n290 8.14595
R5344 vdd.n241 vdd.n235 8.14595
R5345 vdd.n198 vdd.n192 8.14595
R5346 vdd.n143 vdd.n137 8.14595
R5347 vdd.n101 vdd.n95 8.14595
R5348 vdd.n46 vdd.n40 8.14595
R5349 vdd.n2027 vdd.n2021 8.14595
R5350 vdd.n2082 vdd.n2076 8.14595
R5351 vdd.n1929 vdd.n1923 8.14595
R5352 vdd.n1984 vdd.n1978 8.14595
R5353 vdd.n1832 vdd.n1826 8.14595
R5354 vdd.n1887 vdd.n1881 8.14595
R5355 vdd.t80 vdd.n1500 7.8227
R5356 vdd.t84 vdd.n363 7.8227
R5357 vdd.n2341 vdd.n1047 7.70933
R5358 vdd.n2341 vdd.n1050 7.70933
R5359 vdd.n2347 vdd.n1036 7.70933
R5360 vdd.n2353 vdd.n1036 7.70933
R5361 vdd.n2353 vdd.n1030 7.70933
R5362 vdd.n2359 vdd.n1030 7.70933
R5363 vdd.n2365 vdd.n1023 7.70933
R5364 vdd.n2365 vdd.n1026 7.70933
R5365 vdd.n2371 vdd.n1019 7.70933
R5366 vdd.n2378 vdd.n1005 7.70933
R5367 vdd.n2384 vdd.n1005 7.70933
R5368 vdd.n2390 vdd.n999 7.70933
R5369 vdd.n2396 vdd.n995 7.70933
R5370 vdd.n2402 vdd.n989 7.70933
R5371 vdd.n2414 vdd.n976 7.70933
R5372 vdd.n2420 vdd.n970 7.70933
R5373 vdd.n2420 vdd.n963 7.70933
R5374 vdd.n2428 vdd.n963 7.70933
R5375 vdd.n2510 vdd.n947 7.70933
R5376 vdd.n2862 vdd.n899 7.70933
R5377 vdd.n2874 vdd.n888 7.70933
R5378 vdd.n2874 vdd.n882 7.70933
R5379 vdd.n2880 vdd.n882 7.70933
R5380 vdd.n2886 vdd.n876 7.70933
R5381 vdd.n2892 vdd.n872 7.70933
R5382 vdd.n2898 vdd.n866 7.70933
R5383 vdd.n2910 vdd.n853 7.70933
R5384 vdd.n2916 vdd.n846 7.70933
R5385 vdd.n2916 vdd.n849 7.70933
R5386 vdd.n2923 vdd.n841 7.70933
R5387 vdd.n2929 vdd.n828 7.70933
R5388 vdd.n2935 vdd.n828 7.70933
R5389 vdd.n2941 vdd.n822 7.70933
R5390 vdd.n2941 vdd.n814 7.70933
R5391 vdd.n2992 vdd.n814 7.70933
R5392 vdd.n2992 vdd.n817 7.70933
R5393 vdd.n2998 vdd.n774 7.70933
R5394 vdd.n3068 vdd.n774 7.70933
R5395 vdd.n2921 vdd.n2920 7.49318
R5396 vdd.n2375 vdd.n2374 7.49318
R5397 vdd.n295 vdd.n292 7.3702
R5398 vdd.n240 vdd.n237 7.3702
R5399 vdd.n197 vdd.n194 7.3702
R5400 vdd.n142 vdd.n139 7.3702
R5401 vdd.n100 vdd.n97 7.3702
R5402 vdd.n45 vdd.n42 7.3702
R5403 vdd.n2026 vdd.n2023 7.3702
R5404 vdd.n2081 vdd.n2078 7.3702
R5405 vdd.n1928 vdd.n1925 7.3702
R5406 vdd.n1983 vdd.n1980 7.3702
R5407 vdd.n1831 vdd.n1828 7.3702
R5408 vdd.n1886 vdd.n1883 7.3702
R5409 vdd.n2359 vdd.t28 7.36923
R5410 vdd.t10 vdd.n822 7.36923
R5411 vdd.n2435 vdd.t5 7.25587
R5412 vdd.n2779 vdd.t31 7.25587
R5413 vdd.n1669 vdd.n1668 6.98232
R5414 vdd.n2225 vdd.n2224 6.98232
R5415 vdd.n547 vdd.n546 6.98232
R5416 vdd.n3152 vdd.n3151 6.98232
R5417 vdd.n2156 vdd.t142 6.91577
R5418 vdd.n3261 vdd.t236 6.91577
R5419 vdd.t220 vdd.n1437 6.68904
R5420 vdd.n3277 vdd.t189 6.68904
R5421 vdd.n2114 vdd.t158 6.46231
R5422 vdd.n3305 vdd.t156 6.46231
R5423 vdd.n3384 vdd.n321 6.32949
R5424 vdd.n2108 vdd.n2107 6.32949
R5425 vdd.t217 vdd.n1465 6.23558
R5426 vdd.t154 vdd.n332 6.23558
R5427 vdd.n1778 vdd.t172 6.00885
R5428 vdd.n3363 vdd.t152 6.00885
R5429 vdd.t2 vdd.n976 5.89549
R5430 vdd.n2886 vdd.t34 5.89549
R5431 vdd.n296 vdd.n295 5.81868
R5432 vdd.n241 vdd.n240 5.81868
R5433 vdd.n198 vdd.n197 5.81868
R5434 vdd.n143 vdd.n142 5.81868
R5435 vdd.n101 vdd.n100 5.81868
R5436 vdd.n46 vdd.n45 5.81868
R5437 vdd.n2027 vdd.n2026 5.81868
R5438 vdd.n2082 vdd.n2081 5.81868
R5439 vdd.n1929 vdd.n1928 5.81868
R5440 vdd.n1984 vdd.n1983 5.81868
R5441 vdd.n1832 vdd.n1831 5.81868
R5442 vdd.n1887 vdd.n1886 5.81868
R5443 vdd.n2518 vdd.n2517 5.77611
R5444 vdd.n1274 vdd.n1273 5.77611
R5445 vdd.n2791 vdd.n2790 5.77611
R5446 vdd.n3007 vdd.n806 5.77611
R5447 vdd.n3073 vdd.n770 5.77611
R5448 vdd.n2685 vdd.n2623 5.77611
R5449 vdd.n2443 vdd.n954 5.77611
R5450 vdd.n1363 vdd.n1226 5.77611
R5451 vdd.n1738 vdd.n1512 5.62474
R5452 vdd.n2188 vdd.n2185 5.62474
R5453 vdd.n3342 vdd.n407 5.62474
R5454 vdd.n3107 vdd.n3104 5.62474
R5455 vdd.t23 vdd.n999 5.55539
R5456 vdd.n2390 vdd.t0 5.55539
R5457 vdd.t1 vdd.n853 5.55539
R5458 vdd.n2910 vdd.t36 5.55539
R5459 vdd.n1019 vdd.t105 5.44203
R5460 vdd.n2923 vdd.t73 5.44203
R5461 vdd.n1488 vdd.t172 5.32866
R5462 vdd.n2347 vdd.t55 5.32866
R5463 vdd.n1309 vdd.t97 5.32866
R5464 vdd.n2868 vdd.t101 5.32866
R5465 vdd.n817 vdd.t51 5.32866
R5466 vdd.t152 vdd.n3362 5.32866
R5467 vdd.n1794 vdd.t217 5.10193
R5468 vdd.n3371 vdd.t154 5.10193
R5469 vdd.n299 vdd.n290 5.04292
R5470 vdd.n244 vdd.n235 5.04292
R5471 vdd.n201 vdd.n192 5.04292
R5472 vdd.n146 vdd.n137 5.04292
R5473 vdd.n104 vdd.n95 5.04292
R5474 vdd.n49 vdd.n40 5.04292
R5475 vdd.n2030 vdd.n2021 5.04292
R5476 vdd.n2085 vdd.n2076 5.04292
R5477 vdd.n1932 vdd.n1923 5.04292
R5478 vdd.n1987 vdd.n1978 5.04292
R5479 vdd.n1835 vdd.n1826 5.04292
R5480 vdd.n1890 vdd.n1881 5.04292
R5481 vdd.n2396 vdd.t24 4.98857
R5482 vdd.n866 vdd.t48 4.98857
R5483 vdd.n1810 vdd.t158 4.8752
R5484 vdd.t4 vdd.t126 4.8752
R5485 vdd.t9 vdd.t37 4.8752
R5486 vdd.t12 vdd.t11 4.8752
R5487 vdd.t20 vdd.t33 4.8752
R5488 vdd.t156 vdd.n328 4.8752
R5489 vdd.n2519 vdd.n2518 4.83952
R5490 vdd.n1273 vdd.n1272 4.83952
R5491 vdd.n2792 vdd.n2791 4.83952
R5492 vdd.n806 vdd.n801 4.83952
R5493 vdd.n770 vdd.n765 4.83952
R5494 vdd.n2682 vdd.n2623 4.83952
R5495 vdd.n2446 vdd.n954 4.83952
R5496 vdd.n1366 vdd.n1226 4.83952
R5497 vdd.n2193 vdd.n2192 4.74817
R5498 vdd.n1399 vdd.n1394 4.74817
R5499 vdd.n1096 vdd.n1093 4.74817
R5500 vdd.n2286 vdd.n1092 4.74817
R5501 vdd.n2291 vdd.n1093 4.74817
R5502 vdd.n2290 vdd.n1092 4.74817
R5503 vdd.n664 vdd.n662 4.74817
R5504 vdd.n3222 vdd.n665 4.74817
R5505 vdd.n3225 vdd.n665 4.74817
R5506 vdd.n3226 vdd.n664 4.74817
R5507 vdd.n3114 vdd.n749 4.74817
R5508 vdd.n3110 vdd.n751 4.74817
R5509 vdd.n3113 vdd.n751 4.74817
R5510 vdd.n3118 vdd.n749 4.74817
R5511 vdd.n2192 vdd.n1192 4.74817
R5512 vdd.n1396 vdd.n1394 4.74817
R5513 vdd.n321 vdd.n320 4.7074
R5514 vdd.n223 vdd.n222 4.7074
R5515 vdd.n2107 vdd.n2106 4.7074
R5516 vdd.n2009 vdd.n2008 4.7074
R5517 vdd.n2130 vdd.t220 4.64847
R5518 vdd.n2371 vdd.t16 4.64847
R5519 vdd.n989 vdd.t8 4.64847
R5520 vdd.n2892 vdd.t45 4.64847
R5521 vdd.n841 vdd.t7 4.64847
R5522 vdd.n3286 vdd.t189 4.64847
R5523 vdd.n1431 vdd.t142 4.42174
R5524 vdd.t236 vdd.n635 4.42174
R5525 vdd.n300 vdd.n288 4.26717
R5526 vdd.n245 vdd.n233 4.26717
R5527 vdd.n202 vdd.n190 4.26717
R5528 vdd.n147 vdd.n135 4.26717
R5529 vdd.n105 vdd.n93 4.26717
R5530 vdd.n50 vdd.n38 4.26717
R5531 vdd.n2031 vdd.n2019 4.26717
R5532 vdd.n2086 vdd.n2074 4.26717
R5533 vdd.n1933 vdd.n1921 4.26717
R5534 vdd.n1988 vdd.n1976 4.26717
R5535 vdd.n1836 vdd.n1824 4.26717
R5536 vdd.n1891 vdd.n1879 4.26717
R5537 vdd.n321 vdd.n223 4.10845
R5538 vdd.n2107 vdd.n2009 4.10845
R5539 vdd.n277 vdd.t169 4.06363
R5540 vdd.n277 vdd.t224 4.06363
R5541 vdd.n275 vdd.t249 4.06363
R5542 vdd.n275 vdd.t258 4.06363
R5543 vdd.n273 vdd.t262 4.06363
R5544 vdd.n273 vdd.t176 4.06363
R5545 vdd.n271 vdd.t201 4.06363
R5546 vdd.n271 vdd.t261 4.06363
R5547 vdd.n269 vdd.t263 4.06363
R5548 vdd.n269 vdd.t200 4.06363
R5549 vdd.n267 vdd.t205 4.06363
R5550 vdd.n267 vdd.t209 4.06363
R5551 vdd.n265 vdd.t244 4.06363
R5552 vdd.n265 vdd.t160 4.06363
R5553 vdd.n179 vdd.t153 4.06363
R5554 vdd.n179 vdd.t207 4.06363
R5555 vdd.n177 vdd.t238 4.06363
R5556 vdd.n177 vdd.t250 4.06363
R5557 vdd.n175 vdd.t254 4.06363
R5558 vdd.n175 vdd.t155 4.06363
R5559 vdd.n173 vdd.t186 4.06363
R5560 vdd.n173 vdd.t253 4.06363
R5561 vdd.n171 vdd.t255 4.06363
R5562 vdd.n171 vdd.t185 4.06363
R5563 vdd.n169 vdd.t188 4.06363
R5564 vdd.n169 vdd.t190 4.06363
R5565 vdd.n167 vdd.t237 4.06363
R5566 vdd.n167 vdd.t139 4.06363
R5567 vdd.n82 vdd.t168 4.06363
R5568 vdd.n82 vdd.t243 4.06363
R5569 vdd.n80 vdd.t162 4.06363
R5570 vdd.n80 vdd.t231 4.06363
R5571 vdd.n78 vdd.t183 4.06363
R5572 vdd.n78 vdd.t251 4.06363
R5573 vdd.n76 vdd.t157 4.06363
R5574 vdd.n76 vdd.t212 4.06363
R5575 vdd.n74 vdd.t147 4.06363
R5576 vdd.n74 vdd.t193 4.06363
R5577 vdd.n72 vdd.t259 4.06363
R5578 vdd.n72 vdd.t242 4.06363
R5579 vdd.n70 vdd.t247 4.06363
R5580 vdd.n70 vdd.t202 4.06363
R5581 vdd.n2051 vdd.t219 4.06363
R5582 vdd.n2051 vdd.t165 4.06363
R5583 vdd.n2053 vdd.t265 4.06363
R5584 vdd.n2053 vdd.t241 4.06363
R5585 vdd.n2055 vdd.t239 4.06363
R5586 vdd.n2055 vdd.t199 4.06363
R5587 vdd.n2057 vdd.t192 4.06363
R5588 vdd.n2057 vdd.t240 4.06363
R5589 vdd.n2059 vdd.t227 4.06363
R5590 vdd.n2059 vdd.t226 4.06363
R5591 vdd.n2061 vdd.t191 4.06363
R5592 vdd.n2061 vdd.t167 4.06363
R5593 vdd.n2063 vdd.t164 4.06363
R5594 vdd.n2063 vdd.t225 4.06363
R5595 vdd.n1953 vdd.t208 4.06363
R5596 vdd.n1953 vdd.t143 4.06363
R5597 vdd.n1955 vdd.t257 4.06363
R5598 vdd.n1955 vdd.t234 4.06363
R5599 vdd.n1957 vdd.t228 4.06363
R5600 vdd.n1957 vdd.t181 4.06363
R5601 vdd.n1959 vdd.t175 4.06363
R5602 vdd.n1959 vdd.t229 4.06363
R5603 vdd.n1961 vdd.t218 4.06363
R5604 vdd.n1961 vdd.t216 4.06363
R5605 vdd.n1963 vdd.t171 4.06363
R5606 vdd.n1963 vdd.t149 4.06363
R5607 vdd.n1965 vdd.t141 4.06363
R5608 vdd.n1965 vdd.t214 4.06363
R5609 vdd.n1856 vdd.t204 4.06363
R5610 vdd.n1856 vdd.t248 4.06363
R5611 vdd.n1858 vdd.t221 4.06363
R5612 vdd.n1858 vdd.t260 4.06363
R5613 vdd.n1860 vdd.t195 4.06363
R5614 vdd.n1860 vdd.t151 4.06363
R5615 vdd.n1862 vdd.t213 4.06363
R5616 vdd.n1862 vdd.t159 4.06363
R5617 vdd.n1864 vdd.t252 4.06363
R5618 vdd.n1864 vdd.t264 4.06363
R5619 vdd.n1866 vdd.t232 4.06363
R5620 vdd.n1866 vdd.t163 4.06363
R5621 vdd.n1868 vdd.t222 4.06363
R5622 vdd.n1868 vdd.t173 4.06363
R5623 vdd.n26 vdd.t136 3.9605
R5624 vdd.n26 vdd.t132 3.9605
R5625 vdd.n23 vdd.t41 3.9605
R5626 vdd.n23 vdd.t42 3.9605
R5627 vdd.n21 vdd.t131 3.9605
R5628 vdd.n21 vdd.t128 3.9605
R5629 vdd.n20 vdd.t135 3.9605
R5630 vdd.n20 vdd.t40 3.9605
R5631 vdd.n15 vdd.t130 3.9605
R5632 vdd.n15 vdd.t43 3.9605
R5633 vdd.n16 vdd.t134 3.9605
R5634 vdd.n16 vdd.t39 3.9605
R5635 vdd.n18 vdd.t133 3.9605
R5636 vdd.n18 vdd.t44 3.9605
R5637 vdd.n25 vdd.t129 3.9605
R5638 vdd.n25 vdd.t137 3.9605
R5639 vdd.n2428 vdd.t46 3.85492
R5640 vdd.n1309 vdd.t46 3.85492
R5641 vdd.n2868 vdd.t29 3.85492
R5642 vdd.t29 vdd.n888 3.85492
R5643 vdd.n7 vdd.t21 3.61217
R5644 vdd.n7 vdd.t49 3.61217
R5645 vdd.n8 vdd.t13 3.61217
R5646 vdd.n8 vdd.t35 3.61217
R5647 vdd.n10 vdd.t32 3.61217
R5648 vdd.n10 vdd.t30 3.61217
R5649 vdd.n12 vdd.t15 3.61217
R5650 vdd.n12 vdd.t18 3.61217
R5651 vdd.n5 vdd.t267 3.61217
R5652 vdd.n5 vdd.t27 3.61217
R5653 vdd.n3 vdd.t47 3.61217
R5654 vdd.n3 vdd.t6 3.61217
R5655 vdd.n1 vdd.t3 3.61217
R5656 vdd.n1 vdd.t38 3.61217
R5657 vdd.n0 vdd.t25 3.61217
R5658 vdd.n0 vdd.t127 3.61217
R5659 vdd.n1744 vdd.t80 3.51482
R5660 vdd.n3347 vdd.t84 3.51482
R5661 vdd.n304 vdd.n303 3.49141
R5662 vdd.n249 vdd.n248 3.49141
R5663 vdd.n206 vdd.n205 3.49141
R5664 vdd.n151 vdd.n150 3.49141
R5665 vdd.n109 vdd.n108 3.49141
R5666 vdd.n54 vdd.n53 3.49141
R5667 vdd.n2035 vdd.n2034 3.49141
R5668 vdd.n2090 vdd.n2089 3.49141
R5669 vdd.n1937 vdd.n1936 3.49141
R5670 vdd.n1992 vdd.n1991 3.49141
R5671 vdd.n1840 vdd.n1839 3.49141
R5672 vdd.n1895 vdd.n1894 3.49141
R5673 vdd.n2582 vdd.t266 3.40145
R5674 vdd.n2855 vdd.t17 3.40145
R5675 vdd.n2920 vdd.n2919 3.12245
R5676 vdd.n2376 vdd.n2375 3.12245
R5677 vdd.n2147 vdd.t203 3.06136
R5678 vdd.n1026 vdd.t16 3.06136
R5679 vdd.n2408 vdd.t8 3.06136
R5680 vdd.n2764 vdd.t45 3.06136
R5681 vdd.n2929 vdd.t7 3.06136
R5682 vdd.n3269 vdd.t138 3.06136
R5683 vdd.t150 vdd.n1443 2.83463
R5684 vdd.n624 vdd.t146 2.83463
R5685 vdd.n1330 vdd.t24 2.72126
R5686 vdd.n2904 vdd.t48 2.72126
R5687 vdd.n307 vdd.n286 2.71565
R5688 vdd.n252 vdd.n231 2.71565
R5689 vdd.n209 vdd.n188 2.71565
R5690 vdd.n154 vdd.n133 2.71565
R5691 vdd.n112 vdd.n91 2.71565
R5692 vdd.n57 vdd.n36 2.71565
R5693 vdd.n2038 vdd.n2017 2.71565
R5694 vdd.n2093 vdd.n2072 2.71565
R5695 vdd.n1940 vdd.n1919 2.71565
R5696 vdd.n1995 vdd.n1974 2.71565
R5697 vdd.n1843 vdd.n1822 2.71565
R5698 vdd.n1898 vdd.n1877 2.71565
R5699 vdd.n1811 vdd.t174 2.6079
R5700 vdd.n3379 vdd.t211 2.6079
R5701 vdd.t37 vdd.n970 2.49453
R5702 vdd.n2880 vdd.t12 2.49453
R5703 vdd.n294 vdd.n293 2.4129
R5704 vdd.n239 vdd.n238 2.4129
R5705 vdd.n196 vdd.n195 2.4129
R5706 vdd.n141 vdd.n140 2.4129
R5707 vdd.n99 vdd.n98 2.4129
R5708 vdd.n44 vdd.n43 2.4129
R5709 vdd.n2025 vdd.n2024 2.4129
R5710 vdd.n2080 vdd.n2079 2.4129
R5711 vdd.n1927 vdd.n1926 2.4129
R5712 vdd.n1982 vdd.n1981 2.4129
R5713 vdd.n1830 vdd.n1829 2.4129
R5714 vdd.n1885 vdd.n1884 2.4129
R5715 vdd.t148 vdd.n1472 2.38117
R5716 vdd.n1050 vdd.t55 2.38117
R5717 vdd.n2435 vdd.t97 2.38117
R5718 vdd.n2779 vdd.t101 2.38117
R5719 vdd.n2998 vdd.t51 2.38117
R5720 vdd.n3370 vdd.t161 2.38117
R5721 vdd.n2298 vdd.n1093 2.27742
R5722 vdd.n2298 vdd.n1092 2.27742
R5723 vdd.n3034 vdd.n665 2.27742
R5724 vdd.n3034 vdd.n664 2.27742
R5725 vdd.n3102 vdd.n751 2.27742
R5726 vdd.n3102 vdd.n749 2.27742
R5727 vdd.n2192 vdd.n2191 2.27742
R5728 vdd.n2191 vdd.n1394 2.27742
R5729 vdd.n1769 vdd.t140 2.15444
R5730 vdd.n2384 vdd.t23 2.15444
R5731 vdd.n1330 vdd.t0 2.15444
R5732 vdd.n2904 vdd.t1 2.15444
R5733 vdd.t36 vdd.n846 2.15444
R5734 vdd.n3361 vdd.t206 2.15444
R5735 vdd.n308 vdd.n284 1.93989
R5736 vdd.n253 vdd.n229 1.93989
R5737 vdd.n210 vdd.n186 1.93989
R5738 vdd.n155 vdd.n131 1.93989
R5739 vdd.n113 vdd.n89 1.93989
R5740 vdd.n58 vdd.n34 1.93989
R5741 vdd.n2039 vdd.n2015 1.93989
R5742 vdd.n2094 vdd.n2070 1.93989
R5743 vdd.n1941 vdd.n1917 1.93989
R5744 vdd.n1996 vdd.n1972 1.93989
R5745 vdd.n1844 vdd.n1820 1.93989
R5746 vdd.n1899 vdd.n1875 1.93989
R5747 vdd.n2408 vdd.t2 1.81434
R5748 vdd.n2764 vdd.t34 1.81434
R5749 vdd.n1761 vdd.t144 1.70098
R5750 vdd.n3355 vdd.t196 1.70098
R5751 vdd.n2402 vdd.t126 1.58761
R5752 vdd.n872 vdd.t20 1.58761
R5753 vdd.n1777 vdd.t170 1.47425
R5754 vdd.n349 vdd.t230 1.47425
R5755 vdd.n1802 vdd.t215 1.24752
R5756 vdd.t63 vdd.n1407 1.24752
R5757 vdd.n2378 vdd.t22 1.24752
R5758 vdd.n995 vdd.t4 1.24752
R5759 vdd.n2898 vdd.t33 1.24752
R5760 vdd.n849 vdd.t19 1.24752
R5761 vdd.n659 vdd.t59 1.24752
R5762 vdd.t182 vdd.n3377 1.24752
R5763 vdd.n319 vdd.n279 1.16414
R5764 vdd.n312 vdd.n311 1.16414
R5765 vdd.n264 vdd.n224 1.16414
R5766 vdd.n257 vdd.n256 1.16414
R5767 vdd.n221 vdd.n181 1.16414
R5768 vdd.n214 vdd.n213 1.16414
R5769 vdd.n166 vdd.n126 1.16414
R5770 vdd.n159 vdd.n158 1.16414
R5771 vdd.n124 vdd.n84 1.16414
R5772 vdd.n117 vdd.n116 1.16414
R5773 vdd.n69 vdd.n29 1.16414
R5774 vdd.n62 vdd.n61 1.16414
R5775 vdd.n2050 vdd.n2010 1.16414
R5776 vdd.n2043 vdd.n2042 1.16414
R5777 vdd.n2105 vdd.n2065 1.16414
R5778 vdd.n2098 vdd.n2097 1.16414
R5779 vdd.n1952 vdd.n1912 1.16414
R5780 vdd.n1945 vdd.n1944 1.16414
R5781 vdd.n2007 vdd.n1967 1.16414
R5782 vdd.n2000 vdd.n1999 1.16414
R5783 vdd.n1855 vdd.n1815 1.16414
R5784 vdd.n1848 vdd.n1847 1.16414
R5785 vdd.n1910 vdd.n1870 1.16414
R5786 vdd.n1903 vdd.n1902 1.16414
R5787 vdd.n1454 vdd.t194 1.02079
R5788 vdd.t105 vdd.t22 1.02079
R5789 vdd.t19 vdd.t73 1.02079
R5790 vdd.t184 vdd.n613 1.02079
R5791 vdd.n1633 vdd.n1512 0.970197
R5792 vdd.n2189 vdd.n2188 0.970197
R5793 vdd.n599 vdd.n407 0.970197
R5794 vdd.n3109 vdd.n3107 0.970197
R5795 vdd.n2108 vdd.n28 0.956323
R5796 vdd vdd.n3384 0.94849
R5797 vdd.n2139 vdd.t233 0.794056
R5798 vdd.n3278 vdd.t187 0.794056
R5799 vdd.n2155 vdd.t179 0.567326
R5800 vdd.t177 vdd.n642 0.567326
R5801 vdd.n2179 vdd.n1094 0.482207
R5802 vdd.n3234 vdd.n3233 0.482207
R5803 vdd.n444 vdd.n443 0.482207
R5804 vdd.n3341 vdd.n3340 0.482207
R5805 vdd.n3240 vdd.n656 0.482207
R5806 vdd.n2169 vdd.n1395 0.482207
R5807 vdd.n1740 vdd.n1739 0.482207
R5808 vdd.n1546 vdd.n1503 0.482207
R5809 vdd.n4 vdd.n2 0.459552
R5810 vdd.n11 vdd.n9 0.459552
R5811 vdd.t5 vdd.n947 0.453961
R5812 vdd.n2862 vdd.t31 0.453961
R5813 vdd.n317 vdd.n316 0.388379
R5814 vdd.n283 vdd.n281 0.388379
R5815 vdd.n262 vdd.n261 0.388379
R5816 vdd.n228 vdd.n226 0.388379
R5817 vdd.n219 vdd.n218 0.388379
R5818 vdd.n185 vdd.n183 0.388379
R5819 vdd.n164 vdd.n163 0.388379
R5820 vdd.n130 vdd.n128 0.388379
R5821 vdd.n122 vdd.n121 0.388379
R5822 vdd.n88 vdd.n86 0.388379
R5823 vdd.n67 vdd.n66 0.388379
R5824 vdd.n33 vdd.n31 0.388379
R5825 vdd.n2048 vdd.n2047 0.388379
R5826 vdd.n2014 vdd.n2012 0.388379
R5827 vdd.n2103 vdd.n2102 0.388379
R5828 vdd.n2069 vdd.n2067 0.388379
R5829 vdd.n1950 vdd.n1949 0.388379
R5830 vdd.n1916 vdd.n1914 0.388379
R5831 vdd.n2005 vdd.n2004 0.388379
R5832 vdd.n1971 vdd.n1969 0.388379
R5833 vdd.n1853 vdd.n1852 0.388379
R5834 vdd.n1819 vdd.n1817 0.388379
R5835 vdd.n1908 vdd.n1907 0.388379
R5836 vdd.n1874 vdd.n1872 0.388379
R5837 vdd.n19 vdd.n17 0.387128
R5838 vdd.n24 vdd.n22 0.387128
R5839 vdd.n6 vdd.n4 0.358259
R5840 vdd.n13 vdd.n11 0.358259
R5841 vdd.n268 vdd.n266 0.358259
R5842 vdd.n270 vdd.n268 0.358259
R5843 vdd.n272 vdd.n270 0.358259
R5844 vdd.n274 vdd.n272 0.358259
R5845 vdd.n276 vdd.n274 0.358259
R5846 vdd.n278 vdd.n276 0.358259
R5847 vdd.n320 vdd.n278 0.358259
R5848 vdd.n170 vdd.n168 0.358259
R5849 vdd.n172 vdd.n170 0.358259
R5850 vdd.n174 vdd.n172 0.358259
R5851 vdd.n176 vdd.n174 0.358259
R5852 vdd.n178 vdd.n176 0.358259
R5853 vdd.n180 vdd.n178 0.358259
R5854 vdd.n222 vdd.n180 0.358259
R5855 vdd.n73 vdd.n71 0.358259
R5856 vdd.n75 vdd.n73 0.358259
R5857 vdd.n77 vdd.n75 0.358259
R5858 vdd.n79 vdd.n77 0.358259
R5859 vdd.n81 vdd.n79 0.358259
R5860 vdd.n83 vdd.n81 0.358259
R5861 vdd.n125 vdd.n83 0.358259
R5862 vdd.n2106 vdd.n2064 0.358259
R5863 vdd.n2064 vdd.n2062 0.358259
R5864 vdd.n2062 vdd.n2060 0.358259
R5865 vdd.n2060 vdd.n2058 0.358259
R5866 vdd.n2058 vdd.n2056 0.358259
R5867 vdd.n2056 vdd.n2054 0.358259
R5868 vdd.n2054 vdd.n2052 0.358259
R5869 vdd.n2008 vdd.n1966 0.358259
R5870 vdd.n1966 vdd.n1964 0.358259
R5871 vdd.n1964 vdd.n1962 0.358259
R5872 vdd.n1962 vdd.n1960 0.358259
R5873 vdd.n1960 vdd.n1958 0.358259
R5874 vdd.n1958 vdd.n1956 0.358259
R5875 vdd.n1956 vdd.n1954 0.358259
R5876 vdd.n1911 vdd.n1869 0.358259
R5877 vdd.n1869 vdd.n1867 0.358259
R5878 vdd.n1867 vdd.n1865 0.358259
R5879 vdd.n1865 vdd.n1863 0.358259
R5880 vdd.n1863 vdd.n1861 0.358259
R5881 vdd.n1861 vdd.n1859 0.358259
R5882 vdd.n1859 vdd.n1857 0.358259
R5883 vdd.t28 vdd.n1023 0.340595
R5884 vdd.n2414 vdd.t9 0.340595
R5885 vdd.t11 vdd.n876 0.340595
R5886 vdd.n2935 vdd.t10 0.340595
R5887 vdd.n14 vdd.n6 0.334552
R5888 vdd.n14 vdd.n13 0.334552
R5889 vdd.n27 vdd.n19 0.21707
R5890 vdd.n27 vdd.n24 0.21707
R5891 vdd.n318 vdd.n280 0.155672
R5892 vdd.n310 vdd.n280 0.155672
R5893 vdd.n310 vdd.n309 0.155672
R5894 vdd.n309 vdd.n285 0.155672
R5895 vdd.n302 vdd.n285 0.155672
R5896 vdd.n302 vdd.n301 0.155672
R5897 vdd.n301 vdd.n289 0.155672
R5898 vdd.n294 vdd.n289 0.155672
R5899 vdd.n263 vdd.n225 0.155672
R5900 vdd.n255 vdd.n225 0.155672
R5901 vdd.n255 vdd.n254 0.155672
R5902 vdd.n254 vdd.n230 0.155672
R5903 vdd.n247 vdd.n230 0.155672
R5904 vdd.n247 vdd.n246 0.155672
R5905 vdd.n246 vdd.n234 0.155672
R5906 vdd.n239 vdd.n234 0.155672
R5907 vdd.n220 vdd.n182 0.155672
R5908 vdd.n212 vdd.n182 0.155672
R5909 vdd.n212 vdd.n211 0.155672
R5910 vdd.n211 vdd.n187 0.155672
R5911 vdd.n204 vdd.n187 0.155672
R5912 vdd.n204 vdd.n203 0.155672
R5913 vdd.n203 vdd.n191 0.155672
R5914 vdd.n196 vdd.n191 0.155672
R5915 vdd.n165 vdd.n127 0.155672
R5916 vdd.n157 vdd.n127 0.155672
R5917 vdd.n157 vdd.n156 0.155672
R5918 vdd.n156 vdd.n132 0.155672
R5919 vdd.n149 vdd.n132 0.155672
R5920 vdd.n149 vdd.n148 0.155672
R5921 vdd.n148 vdd.n136 0.155672
R5922 vdd.n141 vdd.n136 0.155672
R5923 vdd.n123 vdd.n85 0.155672
R5924 vdd.n115 vdd.n85 0.155672
R5925 vdd.n115 vdd.n114 0.155672
R5926 vdd.n114 vdd.n90 0.155672
R5927 vdd.n107 vdd.n90 0.155672
R5928 vdd.n107 vdd.n106 0.155672
R5929 vdd.n106 vdd.n94 0.155672
R5930 vdd.n99 vdd.n94 0.155672
R5931 vdd.n68 vdd.n30 0.155672
R5932 vdd.n60 vdd.n30 0.155672
R5933 vdd.n60 vdd.n59 0.155672
R5934 vdd.n59 vdd.n35 0.155672
R5935 vdd.n52 vdd.n35 0.155672
R5936 vdd.n52 vdd.n51 0.155672
R5937 vdd.n51 vdd.n39 0.155672
R5938 vdd.n44 vdd.n39 0.155672
R5939 vdd.n2049 vdd.n2011 0.155672
R5940 vdd.n2041 vdd.n2011 0.155672
R5941 vdd.n2041 vdd.n2040 0.155672
R5942 vdd.n2040 vdd.n2016 0.155672
R5943 vdd.n2033 vdd.n2016 0.155672
R5944 vdd.n2033 vdd.n2032 0.155672
R5945 vdd.n2032 vdd.n2020 0.155672
R5946 vdd.n2025 vdd.n2020 0.155672
R5947 vdd.n2104 vdd.n2066 0.155672
R5948 vdd.n2096 vdd.n2066 0.155672
R5949 vdd.n2096 vdd.n2095 0.155672
R5950 vdd.n2095 vdd.n2071 0.155672
R5951 vdd.n2088 vdd.n2071 0.155672
R5952 vdd.n2088 vdd.n2087 0.155672
R5953 vdd.n2087 vdd.n2075 0.155672
R5954 vdd.n2080 vdd.n2075 0.155672
R5955 vdd.n1951 vdd.n1913 0.155672
R5956 vdd.n1943 vdd.n1913 0.155672
R5957 vdd.n1943 vdd.n1942 0.155672
R5958 vdd.n1942 vdd.n1918 0.155672
R5959 vdd.n1935 vdd.n1918 0.155672
R5960 vdd.n1935 vdd.n1934 0.155672
R5961 vdd.n1934 vdd.n1922 0.155672
R5962 vdd.n1927 vdd.n1922 0.155672
R5963 vdd.n2006 vdd.n1968 0.155672
R5964 vdd.n1998 vdd.n1968 0.155672
R5965 vdd.n1998 vdd.n1997 0.155672
R5966 vdd.n1997 vdd.n1973 0.155672
R5967 vdd.n1990 vdd.n1973 0.155672
R5968 vdd.n1990 vdd.n1989 0.155672
R5969 vdd.n1989 vdd.n1977 0.155672
R5970 vdd.n1982 vdd.n1977 0.155672
R5971 vdd.n1854 vdd.n1816 0.155672
R5972 vdd.n1846 vdd.n1816 0.155672
R5973 vdd.n1846 vdd.n1845 0.155672
R5974 vdd.n1845 vdd.n1821 0.155672
R5975 vdd.n1838 vdd.n1821 0.155672
R5976 vdd.n1838 vdd.n1837 0.155672
R5977 vdd.n1837 vdd.n1825 0.155672
R5978 vdd.n1830 vdd.n1825 0.155672
R5979 vdd.n1909 vdd.n1871 0.155672
R5980 vdd.n1901 vdd.n1871 0.155672
R5981 vdd.n1901 vdd.n1900 0.155672
R5982 vdd.n1900 vdd.n1876 0.155672
R5983 vdd.n1893 vdd.n1876 0.155672
R5984 vdd.n1893 vdd.n1892 0.155672
R5985 vdd.n1892 vdd.n1880 0.155672
R5986 vdd.n1885 vdd.n1880 0.155672
R5987 vdd.n1099 vdd.n1091 0.152939
R5988 vdd.n1103 vdd.n1099 0.152939
R5989 vdd.n1104 vdd.n1103 0.152939
R5990 vdd.n1105 vdd.n1104 0.152939
R5991 vdd.n1106 vdd.n1105 0.152939
R5992 vdd.n1110 vdd.n1106 0.152939
R5993 vdd.n1111 vdd.n1110 0.152939
R5994 vdd.n1112 vdd.n1111 0.152939
R5995 vdd.n1113 vdd.n1112 0.152939
R5996 vdd.n1117 vdd.n1113 0.152939
R5997 vdd.n1118 vdd.n1117 0.152939
R5998 vdd.n1119 vdd.n1118 0.152939
R5999 vdd.n2262 vdd.n1119 0.152939
R6000 vdd.n2262 vdd.n2261 0.152939
R6001 vdd.n2261 vdd.n2260 0.152939
R6002 vdd.n2260 vdd.n1125 0.152939
R6003 vdd.n1130 vdd.n1125 0.152939
R6004 vdd.n1131 vdd.n1130 0.152939
R6005 vdd.n1132 vdd.n1131 0.152939
R6006 vdd.n1136 vdd.n1132 0.152939
R6007 vdd.n1137 vdd.n1136 0.152939
R6008 vdd.n1138 vdd.n1137 0.152939
R6009 vdd.n1139 vdd.n1138 0.152939
R6010 vdd.n1143 vdd.n1139 0.152939
R6011 vdd.n1144 vdd.n1143 0.152939
R6012 vdd.n1145 vdd.n1144 0.152939
R6013 vdd.n1146 vdd.n1145 0.152939
R6014 vdd.n1150 vdd.n1146 0.152939
R6015 vdd.n1151 vdd.n1150 0.152939
R6016 vdd.n1152 vdd.n1151 0.152939
R6017 vdd.n1153 vdd.n1152 0.152939
R6018 vdd.n1157 vdd.n1153 0.152939
R6019 vdd.n1158 vdd.n1157 0.152939
R6020 vdd.n1159 vdd.n1158 0.152939
R6021 vdd.n2223 vdd.n1159 0.152939
R6022 vdd.n2223 vdd.n2222 0.152939
R6023 vdd.n2222 vdd.n2221 0.152939
R6024 vdd.n2221 vdd.n1165 0.152939
R6025 vdd.n1170 vdd.n1165 0.152939
R6026 vdd.n1171 vdd.n1170 0.152939
R6027 vdd.n1172 vdd.n1171 0.152939
R6028 vdd.n1176 vdd.n1172 0.152939
R6029 vdd.n1177 vdd.n1176 0.152939
R6030 vdd.n1178 vdd.n1177 0.152939
R6031 vdd.n1179 vdd.n1178 0.152939
R6032 vdd.n1183 vdd.n1179 0.152939
R6033 vdd.n1184 vdd.n1183 0.152939
R6034 vdd.n1185 vdd.n1184 0.152939
R6035 vdd.n1186 vdd.n1185 0.152939
R6036 vdd.n1190 vdd.n1186 0.152939
R6037 vdd.n1191 vdd.n1190 0.152939
R6038 vdd.n2297 vdd.n1094 0.152939
R6039 vdd.n2111 vdd.n2110 0.152939
R6040 vdd.n2111 vdd.n1446 0.152939
R6041 vdd.n2125 vdd.n1446 0.152939
R6042 vdd.n2126 vdd.n2125 0.152939
R6043 vdd.n2127 vdd.n2126 0.152939
R6044 vdd.n2127 vdd.n1434 0.152939
R6045 vdd.n2142 vdd.n1434 0.152939
R6046 vdd.n2143 vdd.n2142 0.152939
R6047 vdd.n2144 vdd.n2143 0.152939
R6048 vdd.n2144 vdd.n1423 0.152939
R6049 vdd.n2159 vdd.n1423 0.152939
R6050 vdd.n2160 vdd.n2159 0.152939
R6051 vdd.n2161 vdd.n2160 0.152939
R6052 vdd.n2161 vdd.n1411 0.152939
R6053 vdd.n2177 vdd.n1411 0.152939
R6054 vdd.n2178 vdd.n2177 0.152939
R6055 vdd.n2179 vdd.n2178 0.152939
R6056 vdd.n670 vdd.n667 0.152939
R6057 vdd.n671 vdd.n670 0.152939
R6058 vdd.n672 vdd.n671 0.152939
R6059 vdd.n673 vdd.n672 0.152939
R6060 vdd.n676 vdd.n673 0.152939
R6061 vdd.n677 vdd.n676 0.152939
R6062 vdd.n678 vdd.n677 0.152939
R6063 vdd.n679 vdd.n678 0.152939
R6064 vdd.n682 vdd.n679 0.152939
R6065 vdd.n683 vdd.n682 0.152939
R6066 vdd.n684 vdd.n683 0.152939
R6067 vdd.n685 vdd.n684 0.152939
R6068 vdd.n690 vdd.n685 0.152939
R6069 vdd.n691 vdd.n690 0.152939
R6070 vdd.n692 vdd.n691 0.152939
R6071 vdd.n693 vdd.n692 0.152939
R6072 vdd.n696 vdd.n693 0.152939
R6073 vdd.n697 vdd.n696 0.152939
R6074 vdd.n698 vdd.n697 0.152939
R6075 vdd.n699 vdd.n698 0.152939
R6076 vdd.n702 vdd.n699 0.152939
R6077 vdd.n703 vdd.n702 0.152939
R6078 vdd.n704 vdd.n703 0.152939
R6079 vdd.n705 vdd.n704 0.152939
R6080 vdd.n708 vdd.n705 0.152939
R6081 vdd.n709 vdd.n708 0.152939
R6082 vdd.n710 vdd.n709 0.152939
R6083 vdd.n711 vdd.n710 0.152939
R6084 vdd.n714 vdd.n711 0.152939
R6085 vdd.n715 vdd.n714 0.152939
R6086 vdd.n716 vdd.n715 0.152939
R6087 vdd.n717 vdd.n716 0.152939
R6088 vdd.n720 vdd.n717 0.152939
R6089 vdd.n721 vdd.n720 0.152939
R6090 vdd.n3150 vdd.n721 0.152939
R6091 vdd.n3150 vdd.n3149 0.152939
R6092 vdd.n3149 vdd.n3148 0.152939
R6093 vdd.n3148 vdd.n725 0.152939
R6094 vdd.n730 vdd.n725 0.152939
R6095 vdd.n731 vdd.n730 0.152939
R6096 vdd.n734 vdd.n731 0.152939
R6097 vdd.n735 vdd.n734 0.152939
R6098 vdd.n736 vdd.n735 0.152939
R6099 vdd.n737 vdd.n736 0.152939
R6100 vdd.n740 vdd.n737 0.152939
R6101 vdd.n741 vdd.n740 0.152939
R6102 vdd.n742 vdd.n741 0.152939
R6103 vdd.n743 vdd.n742 0.152939
R6104 vdd.n746 vdd.n743 0.152939
R6105 vdd.n747 vdd.n746 0.152939
R6106 vdd.n748 vdd.n747 0.152939
R6107 vdd.n3233 vdd.n661 0.152939
R6108 vdd.n3234 vdd.n651 0.152939
R6109 vdd.n3248 vdd.n651 0.152939
R6110 vdd.n3249 vdd.n3248 0.152939
R6111 vdd.n3250 vdd.n3249 0.152939
R6112 vdd.n3250 vdd.n639 0.152939
R6113 vdd.n3264 vdd.n639 0.152939
R6114 vdd.n3265 vdd.n3264 0.152939
R6115 vdd.n3266 vdd.n3265 0.152939
R6116 vdd.n3266 vdd.n627 0.152939
R6117 vdd.n3281 vdd.n627 0.152939
R6118 vdd.n3282 vdd.n3281 0.152939
R6119 vdd.n3283 vdd.n3282 0.152939
R6120 vdd.n3283 vdd.n616 0.152939
R6121 vdd.n3300 vdd.n616 0.152939
R6122 vdd.n3301 vdd.n3300 0.152939
R6123 vdd.n3302 vdd.n3301 0.152939
R6124 vdd.n3302 vdd.n322 0.152939
R6125 vdd.n3382 vdd.n323 0.152939
R6126 vdd.n334 vdd.n323 0.152939
R6127 vdd.n335 vdd.n334 0.152939
R6128 vdd.n336 vdd.n335 0.152939
R6129 vdd.n343 vdd.n336 0.152939
R6130 vdd.n344 vdd.n343 0.152939
R6131 vdd.n345 vdd.n344 0.152939
R6132 vdd.n346 vdd.n345 0.152939
R6133 vdd.n354 vdd.n346 0.152939
R6134 vdd.n355 vdd.n354 0.152939
R6135 vdd.n356 vdd.n355 0.152939
R6136 vdd.n357 vdd.n356 0.152939
R6137 vdd.n365 vdd.n357 0.152939
R6138 vdd.n366 vdd.n365 0.152939
R6139 vdd.n367 vdd.n366 0.152939
R6140 vdd.n368 vdd.n367 0.152939
R6141 vdd.n443 vdd.n368 0.152939
R6142 vdd.n444 vdd.n442 0.152939
R6143 vdd.n451 vdd.n442 0.152939
R6144 vdd.n452 vdd.n451 0.152939
R6145 vdd.n453 vdd.n452 0.152939
R6146 vdd.n453 vdd.n440 0.152939
R6147 vdd.n461 vdd.n440 0.152939
R6148 vdd.n462 vdd.n461 0.152939
R6149 vdd.n463 vdd.n462 0.152939
R6150 vdd.n463 vdd.n438 0.152939
R6151 vdd.n471 vdd.n438 0.152939
R6152 vdd.n472 vdd.n471 0.152939
R6153 vdd.n473 vdd.n472 0.152939
R6154 vdd.n473 vdd.n436 0.152939
R6155 vdd.n481 vdd.n436 0.152939
R6156 vdd.n482 vdd.n481 0.152939
R6157 vdd.n483 vdd.n482 0.152939
R6158 vdd.n483 vdd.n434 0.152939
R6159 vdd.n491 vdd.n434 0.152939
R6160 vdd.n492 vdd.n491 0.152939
R6161 vdd.n493 vdd.n492 0.152939
R6162 vdd.n493 vdd.n430 0.152939
R6163 vdd.n501 vdd.n430 0.152939
R6164 vdd.n502 vdd.n501 0.152939
R6165 vdd.n503 vdd.n502 0.152939
R6166 vdd.n503 vdd.n428 0.152939
R6167 vdd.n511 vdd.n428 0.152939
R6168 vdd.n512 vdd.n511 0.152939
R6169 vdd.n513 vdd.n512 0.152939
R6170 vdd.n513 vdd.n426 0.152939
R6171 vdd.n521 vdd.n426 0.152939
R6172 vdd.n522 vdd.n521 0.152939
R6173 vdd.n523 vdd.n522 0.152939
R6174 vdd.n523 vdd.n424 0.152939
R6175 vdd.n531 vdd.n424 0.152939
R6176 vdd.n532 vdd.n531 0.152939
R6177 vdd.n533 vdd.n532 0.152939
R6178 vdd.n533 vdd.n422 0.152939
R6179 vdd.n541 vdd.n422 0.152939
R6180 vdd.n542 vdd.n541 0.152939
R6181 vdd.n543 vdd.n542 0.152939
R6182 vdd.n543 vdd.n418 0.152939
R6183 vdd.n551 vdd.n418 0.152939
R6184 vdd.n552 vdd.n551 0.152939
R6185 vdd.n553 vdd.n552 0.152939
R6186 vdd.n553 vdd.n416 0.152939
R6187 vdd.n561 vdd.n416 0.152939
R6188 vdd.n562 vdd.n561 0.152939
R6189 vdd.n563 vdd.n562 0.152939
R6190 vdd.n563 vdd.n414 0.152939
R6191 vdd.n571 vdd.n414 0.152939
R6192 vdd.n572 vdd.n571 0.152939
R6193 vdd.n573 vdd.n572 0.152939
R6194 vdd.n573 vdd.n412 0.152939
R6195 vdd.n581 vdd.n412 0.152939
R6196 vdd.n582 vdd.n581 0.152939
R6197 vdd.n583 vdd.n582 0.152939
R6198 vdd.n583 vdd.n410 0.152939
R6199 vdd.n591 vdd.n410 0.152939
R6200 vdd.n592 vdd.n591 0.152939
R6201 vdd.n593 vdd.n592 0.152939
R6202 vdd.n593 vdd.n408 0.152939
R6203 vdd.n600 vdd.n408 0.152939
R6204 vdd.n3341 vdd.n600 0.152939
R6205 vdd.n3241 vdd.n3240 0.152939
R6206 vdd.n3242 vdd.n3241 0.152939
R6207 vdd.n3242 vdd.n645 0.152939
R6208 vdd.n3256 vdd.n645 0.152939
R6209 vdd.n3257 vdd.n3256 0.152939
R6210 vdd.n3258 vdd.n3257 0.152939
R6211 vdd.n3258 vdd.n632 0.152939
R6212 vdd.n3272 vdd.n632 0.152939
R6213 vdd.n3273 vdd.n3272 0.152939
R6214 vdd.n3274 vdd.n3273 0.152939
R6215 vdd.n3274 vdd.n621 0.152939
R6216 vdd.n3289 vdd.n621 0.152939
R6217 vdd.n3290 vdd.n3289 0.152939
R6218 vdd.n3291 vdd.n3290 0.152939
R6219 vdd.n3293 vdd.n3291 0.152939
R6220 vdd.n3293 vdd.n3292 0.152939
R6221 vdd.n3292 vdd.n611 0.152939
R6222 vdd.n611 vdd.n609 0.152939
R6223 vdd.n3311 vdd.n609 0.152939
R6224 vdd.n3312 vdd.n3311 0.152939
R6225 vdd.n3313 vdd.n3312 0.152939
R6226 vdd.n3313 vdd.n607 0.152939
R6227 vdd.n3318 vdd.n607 0.152939
R6228 vdd.n3319 vdd.n3318 0.152939
R6229 vdd.n3320 vdd.n3319 0.152939
R6230 vdd.n3320 vdd.n605 0.152939
R6231 vdd.n3325 vdd.n605 0.152939
R6232 vdd.n3326 vdd.n3325 0.152939
R6233 vdd.n3327 vdd.n3326 0.152939
R6234 vdd.n3327 vdd.n603 0.152939
R6235 vdd.n3333 vdd.n603 0.152939
R6236 vdd.n3334 vdd.n3333 0.152939
R6237 vdd.n3335 vdd.n3334 0.152939
R6238 vdd.n3335 vdd.n601 0.152939
R6239 vdd.n3340 vdd.n601 0.152939
R6240 vdd.n3103 vdd.n656 0.152939
R6241 vdd.n2190 vdd.n1395 0.152939
R6242 vdd.n1741 vdd.n1740 0.152939
R6243 vdd.n1741 vdd.n1497 0.152939
R6244 vdd.n1755 vdd.n1497 0.152939
R6245 vdd.n1756 vdd.n1755 0.152939
R6246 vdd.n1757 vdd.n1756 0.152939
R6247 vdd.n1757 vdd.n1485 0.152939
R6248 vdd.n1772 vdd.n1485 0.152939
R6249 vdd.n1773 vdd.n1772 0.152939
R6250 vdd.n1774 vdd.n1773 0.152939
R6251 vdd.n1774 vdd.n1475 0.152939
R6252 vdd.n1789 vdd.n1475 0.152939
R6253 vdd.n1790 vdd.n1789 0.152939
R6254 vdd.n1791 vdd.n1790 0.152939
R6255 vdd.n1791 vdd.n1462 0.152939
R6256 vdd.n1805 vdd.n1462 0.152939
R6257 vdd.n1806 vdd.n1805 0.152939
R6258 vdd.n1807 vdd.n1806 0.152939
R6259 vdd.n1807 vdd.n1451 0.152939
R6260 vdd.n2117 vdd.n1451 0.152939
R6261 vdd.n2118 vdd.n2117 0.152939
R6262 vdd.n2119 vdd.n2118 0.152939
R6263 vdd.n2119 vdd.n1440 0.152939
R6264 vdd.n2133 vdd.n1440 0.152939
R6265 vdd.n2134 vdd.n2133 0.152939
R6266 vdd.n2135 vdd.n2134 0.152939
R6267 vdd.n2135 vdd.n1428 0.152939
R6268 vdd.n2150 vdd.n1428 0.152939
R6269 vdd.n2151 vdd.n2150 0.152939
R6270 vdd.n2152 vdd.n2151 0.152939
R6271 vdd.n2152 vdd.n1418 0.152939
R6272 vdd.n2167 vdd.n1418 0.152939
R6273 vdd.n2168 vdd.n2167 0.152939
R6274 vdd.n2171 vdd.n2168 0.152939
R6275 vdd.n2171 vdd.n2170 0.152939
R6276 vdd.n2170 vdd.n2169 0.152939
R6277 vdd.n1731 vdd.n1546 0.152939
R6278 vdd.n1731 vdd.n1730 0.152939
R6279 vdd.n1730 vdd.n1729 0.152939
R6280 vdd.n1729 vdd.n1548 0.152939
R6281 vdd.n1725 vdd.n1548 0.152939
R6282 vdd.n1725 vdd.n1724 0.152939
R6283 vdd.n1724 vdd.n1723 0.152939
R6284 vdd.n1723 vdd.n1553 0.152939
R6285 vdd.n1719 vdd.n1553 0.152939
R6286 vdd.n1719 vdd.n1718 0.152939
R6287 vdd.n1718 vdd.n1717 0.152939
R6288 vdd.n1717 vdd.n1559 0.152939
R6289 vdd.n1713 vdd.n1559 0.152939
R6290 vdd.n1713 vdd.n1712 0.152939
R6291 vdd.n1712 vdd.n1711 0.152939
R6292 vdd.n1711 vdd.n1565 0.152939
R6293 vdd.n1707 vdd.n1565 0.152939
R6294 vdd.n1707 vdd.n1706 0.152939
R6295 vdd.n1706 vdd.n1705 0.152939
R6296 vdd.n1705 vdd.n1571 0.152939
R6297 vdd.n1697 vdd.n1571 0.152939
R6298 vdd.n1697 vdd.n1696 0.152939
R6299 vdd.n1696 vdd.n1695 0.152939
R6300 vdd.n1695 vdd.n1575 0.152939
R6301 vdd.n1691 vdd.n1575 0.152939
R6302 vdd.n1691 vdd.n1690 0.152939
R6303 vdd.n1690 vdd.n1689 0.152939
R6304 vdd.n1689 vdd.n1581 0.152939
R6305 vdd.n1685 vdd.n1581 0.152939
R6306 vdd.n1685 vdd.n1684 0.152939
R6307 vdd.n1684 vdd.n1683 0.152939
R6308 vdd.n1683 vdd.n1587 0.152939
R6309 vdd.n1679 vdd.n1587 0.152939
R6310 vdd.n1679 vdd.n1678 0.152939
R6311 vdd.n1678 vdd.n1677 0.152939
R6312 vdd.n1677 vdd.n1593 0.152939
R6313 vdd.n1673 vdd.n1593 0.152939
R6314 vdd.n1673 vdd.n1672 0.152939
R6315 vdd.n1672 vdd.n1671 0.152939
R6316 vdd.n1671 vdd.n1599 0.152939
R6317 vdd.n1664 vdd.n1599 0.152939
R6318 vdd.n1664 vdd.n1663 0.152939
R6319 vdd.n1663 vdd.n1662 0.152939
R6320 vdd.n1662 vdd.n1604 0.152939
R6321 vdd.n1658 vdd.n1604 0.152939
R6322 vdd.n1658 vdd.n1657 0.152939
R6323 vdd.n1657 vdd.n1656 0.152939
R6324 vdd.n1656 vdd.n1610 0.152939
R6325 vdd.n1652 vdd.n1610 0.152939
R6326 vdd.n1652 vdd.n1651 0.152939
R6327 vdd.n1651 vdd.n1650 0.152939
R6328 vdd.n1650 vdd.n1616 0.152939
R6329 vdd.n1646 vdd.n1616 0.152939
R6330 vdd.n1646 vdd.n1645 0.152939
R6331 vdd.n1645 vdd.n1644 0.152939
R6332 vdd.n1644 vdd.n1622 0.152939
R6333 vdd.n1640 vdd.n1622 0.152939
R6334 vdd.n1640 vdd.n1639 0.152939
R6335 vdd.n1639 vdd.n1638 0.152939
R6336 vdd.n1638 vdd.n1628 0.152939
R6337 vdd.n1634 vdd.n1628 0.152939
R6338 vdd.n1634 vdd.n1509 0.152939
R6339 vdd.n1739 vdd.n1509 0.152939
R6340 vdd.n1747 vdd.n1503 0.152939
R6341 vdd.n1748 vdd.n1747 0.152939
R6342 vdd.n1749 vdd.n1748 0.152939
R6343 vdd.n1749 vdd.n1491 0.152939
R6344 vdd.n1764 vdd.n1491 0.152939
R6345 vdd.n1765 vdd.n1764 0.152939
R6346 vdd.n1766 vdd.n1765 0.152939
R6347 vdd.n1766 vdd.n1480 0.152939
R6348 vdd.n1781 vdd.n1480 0.152939
R6349 vdd.n1782 vdd.n1781 0.152939
R6350 vdd.n1783 vdd.n1782 0.152939
R6351 vdd.n1783 vdd.n1469 0.152939
R6352 vdd.n1797 vdd.n1469 0.152939
R6353 vdd.n1798 vdd.n1797 0.152939
R6354 vdd.n1799 vdd.n1798 0.152939
R6355 vdd.n1799 vdd.n1457 0.152939
R6356 vdd.n1814 vdd.n1457 0.152939
R6357 vdd.n2298 vdd.n2297 0.110256
R6358 vdd.n3034 vdd.n661 0.110256
R6359 vdd.n3103 vdd.n3102 0.110256
R6360 vdd.n2191 vdd.n2190 0.110256
R6361 vdd.n2110 vdd.n2109 0.0695946
R6362 vdd.n3383 vdd.n322 0.0695946
R6363 vdd.n3383 vdd.n3382 0.0695946
R6364 vdd.n2109 vdd.n1814 0.0695946
R6365 vdd.n2298 vdd.n1091 0.0431829
R6366 vdd.n2191 vdd.n1191 0.0431829
R6367 vdd.n3034 vdd.n667 0.0431829
R6368 vdd.n3102 vdd.n748 0.0431829
R6369 vdd vdd.n28 0.00833333
R6370 CSoutput.n19 CSoutput.t180 184.661
R6371 CSoutput.n78 CSoutput.n77 165.8
R6372 CSoutput.n76 CSoutput.n0 165.8
R6373 CSoutput.n75 CSoutput.n74 165.8
R6374 CSoutput.n73 CSoutput.n72 165.8
R6375 CSoutput.n71 CSoutput.n2 165.8
R6376 CSoutput.n69 CSoutput.n68 165.8
R6377 CSoutput.n67 CSoutput.n3 165.8
R6378 CSoutput.n66 CSoutput.n65 165.8
R6379 CSoutput.n63 CSoutput.n4 165.8
R6380 CSoutput.n61 CSoutput.n60 165.8
R6381 CSoutput.n59 CSoutput.n5 165.8
R6382 CSoutput.n58 CSoutput.n57 165.8
R6383 CSoutput.n55 CSoutput.n6 165.8
R6384 CSoutput.n54 CSoutput.n53 165.8
R6385 CSoutput.n52 CSoutput.n51 165.8
R6386 CSoutput.n50 CSoutput.n8 165.8
R6387 CSoutput.n48 CSoutput.n47 165.8
R6388 CSoutput.n46 CSoutput.n9 165.8
R6389 CSoutput.n45 CSoutput.n44 165.8
R6390 CSoutput.n42 CSoutput.n10 165.8
R6391 CSoutput.n41 CSoutput.n40 165.8
R6392 CSoutput.n39 CSoutput.n38 165.8
R6393 CSoutput.n37 CSoutput.n12 165.8
R6394 CSoutput.n35 CSoutput.n34 165.8
R6395 CSoutput.n33 CSoutput.n13 165.8
R6396 CSoutput.n32 CSoutput.n31 165.8
R6397 CSoutput.n29 CSoutput.n14 165.8
R6398 CSoutput.n28 CSoutput.n27 165.8
R6399 CSoutput.n26 CSoutput.n25 165.8
R6400 CSoutput.n24 CSoutput.n16 165.8
R6401 CSoutput.n22 CSoutput.n21 165.8
R6402 CSoutput.n20 CSoutput.n17 165.8
R6403 CSoutput.n77 CSoutput.t183 162.194
R6404 CSoutput.n18 CSoutput.t177 120.501
R6405 CSoutput.n23 CSoutput.t194 120.501
R6406 CSoutput.n15 CSoutput.t189 120.501
R6407 CSoutput.n30 CSoutput.t178 120.501
R6408 CSoutput.n36 CSoutput.t179 120.501
R6409 CSoutput.n11 CSoutput.t191 120.501
R6410 CSoutput.n43 CSoutput.t188 120.501
R6411 CSoutput.n49 CSoutput.t182 120.501
R6412 CSoutput.n7 CSoutput.t195 120.501
R6413 CSoutput.n56 CSoutput.t196 120.501
R6414 CSoutput.n62 CSoutput.t185 120.501
R6415 CSoutput.n64 CSoutput.t197 120.501
R6416 CSoutput.n70 CSoutput.t176 120.501
R6417 CSoutput.n1 CSoutput.t193 120.501
R6418 CSoutput.n310 CSoutput.n308 103.469
R6419 CSoutput.n294 CSoutput.n292 103.469
R6420 CSoutput.n279 CSoutput.n277 103.469
R6421 CSoutput.n112 CSoutput.n110 103.469
R6422 CSoutput.n96 CSoutput.n94 103.469
R6423 CSoutput.n81 CSoutput.n79 103.469
R6424 CSoutput.n320 CSoutput.n319 103.111
R6425 CSoutput.n318 CSoutput.n317 103.111
R6426 CSoutput.n316 CSoutput.n315 103.111
R6427 CSoutput.n314 CSoutput.n313 103.111
R6428 CSoutput.n312 CSoutput.n311 103.111
R6429 CSoutput.n310 CSoutput.n309 103.111
R6430 CSoutput.n306 CSoutput.n305 103.111
R6431 CSoutput.n304 CSoutput.n303 103.111
R6432 CSoutput.n302 CSoutput.n301 103.111
R6433 CSoutput.n300 CSoutput.n299 103.111
R6434 CSoutput.n298 CSoutput.n297 103.111
R6435 CSoutput.n296 CSoutput.n295 103.111
R6436 CSoutput.n294 CSoutput.n293 103.111
R6437 CSoutput.n291 CSoutput.n290 103.111
R6438 CSoutput.n289 CSoutput.n288 103.111
R6439 CSoutput.n287 CSoutput.n286 103.111
R6440 CSoutput.n285 CSoutput.n284 103.111
R6441 CSoutput.n283 CSoutput.n282 103.111
R6442 CSoutput.n281 CSoutput.n280 103.111
R6443 CSoutput.n279 CSoutput.n278 103.111
R6444 CSoutput.n112 CSoutput.n111 103.111
R6445 CSoutput.n114 CSoutput.n113 103.111
R6446 CSoutput.n116 CSoutput.n115 103.111
R6447 CSoutput.n118 CSoutput.n117 103.111
R6448 CSoutput.n120 CSoutput.n119 103.111
R6449 CSoutput.n122 CSoutput.n121 103.111
R6450 CSoutput.n124 CSoutput.n123 103.111
R6451 CSoutput.n96 CSoutput.n95 103.111
R6452 CSoutput.n98 CSoutput.n97 103.111
R6453 CSoutput.n100 CSoutput.n99 103.111
R6454 CSoutput.n102 CSoutput.n101 103.111
R6455 CSoutput.n104 CSoutput.n103 103.111
R6456 CSoutput.n106 CSoutput.n105 103.111
R6457 CSoutput.n108 CSoutput.n107 103.111
R6458 CSoutput.n81 CSoutput.n80 103.111
R6459 CSoutput.n83 CSoutput.n82 103.111
R6460 CSoutput.n85 CSoutput.n84 103.111
R6461 CSoutput.n87 CSoutput.n86 103.111
R6462 CSoutput.n89 CSoutput.n88 103.111
R6463 CSoutput.n91 CSoutput.n90 103.111
R6464 CSoutput.n93 CSoutput.n92 103.111
R6465 CSoutput.n322 CSoutput.n321 103.111
R6466 CSoutput.n346 CSoutput.n344 81.5057
R6467 CSoutput.n327 CSoutput.n325 81.5057
R6468 CSoutput.n386 CSoutput.n384 81.5057
R6469 CSoutput.n367 CSoutput.n365 81.5057
R6470 CSoutput.n362 CSoutput.n361 80.9324
R6471 CSoutput.n360 CSoutput.n359 80.9324
R6472 CSoutput.n358 CSoutput.n357 80.9324
R6473 CSoutput.n356 CSoutput.n355 80.9324
R6474 CSoutput.n354 CSoutput.n353 80.9324
R6475 CSoutput.n352 CSoutput.n351 80.9324
R6476 CSoutput.n350 CSoutput.n349 80.9324
R6477 CSoutput.n348 CSoutput.n347 80.9324
R6478 CSoutput.n346 CSoutput.n345 80.9324
R6479 CSoutput.n343 CSoutput.n342 80.9324
R6480 CSoutput.n341 CSoutput.n340 80.9324
R6481 CSoutput.n339 CSoutput.n338 80.9324
R6482 CSoutput.n337 CSoutput.n336 80.9324
R6483 CSoutput.n335 CSoutput.n334 80.9324
R6484 CSoutput.n333 CSoutput.n332 80.9324
R6485 CSoutput.n331 CSoutput.n330 80.9324
R6486 CSoutput.n329 CSoutput.n328 80.9324
R6487 CSoutput.n327 CSoutput.n326 80.9324
R6488 CSoutput.n386 CSoutput.n385 80.9324
R6489 CSoutput.n388 CSoutput.n387 80.9324
R6490 CSoutput.n390 CSoutput.n389 80.9324
R6491 CSoutput.n392 CSoutput.n391 80.9324
R6492 CSoutput.n394 CSoutput.n393 80.9324
R6493 CSoutput.n396 CSoutput.n395 80.9324
R6494 CSoutput.n398 CSoutput.n397 80.9324
R6495 CSoutput.n400 CSoutput.n399 80.9324
R6496 CSoutput.n402 CSoutput.n401 80.9324
R6497 CSoutput.n367 CSoutput.n366 80.9324
R6498 CSoutput.n369 CSoutput.n368 80.9324
R6499 CSoutput.n371 CSoutput.n370 80.9324
R6500 CSoutput.n373 CSoutput.n372 80.9324
R6501 CSoutput.n375 CSoutput.n374 80.9324
R6502 CSoutput.n377 CSoutput.n376 80.9324
R6503 CSoutput.n379 CSoutput.n378 80.9324
R6504 CSoutput.n381 CSoutput.n380 80.9324
R6505 CSoutput.n383 CSoutput.n382 80.9324
R6506 CSoutput.n25 CSoutput.n24 48.1486
R6507 CSoutput.n69 CSoutput.n3 48.1486
R6508 CSoutput.n38 CSoutput.n37 48.1486
R6509 CSoutput.n42 CSoutput.n41 48.1486
R6510 CSoutput.n51 CSoutput.n50 48.1486
R6511 CSoutput.n55 CSoutput.n54 48.1486
R6512 CSoutput.n22 CSoutput.n17 46.462
R6513 CSoutput.n72 CSoutput.n71 46.462
R6514 CSoutput.n20 CSoutput.n19 44.9055
R6515 CSoutput.n29 CSoutput.n28 43.7635
R6516 CSoutput.n65 CSoutput.n63 43.7635
R6517 CSoutput.n35 CSoutput.n13 41.7396
R6518 CSoutput.n57 CSoutput.n5 41.7396
R6519 CSoutput.n44 CSoutput.n9 37.0171
R6520 CSoutput.n48 CSoutput.n9 37.0171
R6521 CSoutput.n76 CSoutput.n75 34.9932
R6522 CSoutput.n31 CSoutput.n13 32.2947
R6523 CSoutput.n61 CSoutput.n5 32.2947
R6524 CSoutput.n30 CSoutput.n29 29.6014
R6525 CSoutput.n63 CSoutput.n62 29.6014
R6526 CSoutput.n19 CSoutput.n18 28.4085
R6527 CSoutput.n18 CSoutput.n17 25.1176
R6528 CSoutput.n72 CSoutput.n1 25.1176
R6529 CSoutput.n43 CSoutput.n42 22.0922
R6530 CSoutput.n50 CSoutput.n49 22.0922
R6531 CSoutput.n77 CSoutput.n76 21.8586
R6532 CSoutput.n37 CSoutput.n36 18.9681
R6533 CSoutput.n56 CSoutput.n55 18.9681
R6534 CSoutput.n25 CSoutput.n15 17.6292
R6535 CSoutput.n64 CSoutput.n3 17.6292
R6536 CSoutput.n24 CSoutput.n23 15.844
R6537 CSoutput.n70 CSoutput.n69 15.844
R6538 CSoutput.n38 CSoutput.n11 14.5051
R6539 CSoutput.n54 CSoutput.n7 14.5051
R6540 CSoutput.n405 CSoutput.n78 11.6139
R6541 CSoutput.n41 CSoutput.n11 11.3811
R6542 CSoutput.n51 CSoutput.n7 11.3811
R6543 CSoutput.n23 CSoutput.n22 10.0422
R6544 CSoutput.n71 CSoutput.n70 10.0422
R6545 CSoutput.n307 CSoutput.n291 9.25285
R6546 CSoutput.n109 CSoutput.n93 9.25285
R6547 CSoutput.n364 CSoutput.n324 9.09467
R6548 CSoutput.n363 CSoutput.n343 8.97993
R6549 CSoutput.n403 CSoutput.n383 8.97993
R6550 CSoutput.n28 CSoutput.n15 8.25698
R6551 CSoutput.n65 CSoutput.n64 8.25698
R6552 CSoutput.n364 CSoutput.n363 7.89345
R6553 CSoutput.n404 CSoutput.n403 7.89345
R6554 CSoutput.n324 CSoutput.n323 7.12641
R6555 CSoutput.n126 CSoutput.n125 7.12641
R6556 CSoutput.n36 CSoutput.n35 6.91809
R6557 CSoutput.n57 CSoutput.n56 6.91809
R6558 CSoutput.n405 CSoutput.n126 5.50223
R6559 CSoutput.n363 CSoutput.n362 5.25266
R6560 CSoutput.n403 CSoutput.n402 5.25266
R6561 CSoutput.n323 CSoutput.n322 5.1449
R6562 CSoutput.n307 CSoutput.n306 5.1449
R6563 CSoutput.n125 CSoutput.n124 5.1449
R6564 CSoutput.n109 CSoutput.n108 5.1449
R6565 CSoutput.n217 CSoutput.n170 4.5005
R6566 CSoutput.n186 CSoutput.n170 4.5005
R6567 CSoutput.n181 CSoutput.n165 4.5005
R6568 CSoutput.n181 CSoutput.n167 4.5005
R6569 CSoutput.n181 CSoutput.n164 4.5005
R6570 CSoutput.n181 CSoutput.n168 4.5005
R6571 CSoutput.n181 CSoutput.n163 4.5005
R6572 CSoutput.n181 CSoutput.t184 4.5005
R6573 CSoutput.n181 CSoutput.n162 4.5005
R6574 CSoutput.n181 CSoutput.n169 4.5005
R6575 CSoutput.n181 CSoutput.n170 4.5005
R6576 CSoutput.n179 CSoutput.n165 4.5005
R6577 CSoutput.n179 CSoutput.n167 4.5005
R6578 CSoutput.n179 CSoutput.n164 4.5005
R6579 CSoutput.n179 CSoutput.n168 4.5005
R6580 CSoutput.n179 CSoutput.n163 4.5005
R6581 CSoutput.n179 CSoutput.t184 4.5005
R6582 CSoutput.n179 CSoutput.n162 4.5005
R6583 CSoutput.n179 CSoutput.n169 4.5005
R6584 CSoutput.n179 CSoutput.n170 4.5005
R6585 CSoutput.n178 CSoutput.n165 4.5005
R6586 CSoutput.n178 CSoutput.n167 4.5005
R6587 CSoutput.n178 CSoutput.n164 4.5005
R6588 CSoutput.n178 CSoutput.n168 4.5005
R6589 CSoutput.n178 CSoutput.n163 4.5005
R6590 CSoutput.n178 CSoutput.t184 4.5005
R6591 CSoutput.n178 CSoutput.n162 4.5005
R6592 CSoutput.n178 CSoutput.n169 4.5005
R6593 CSoutput.n178 CSoutput.n170 4.5005
R6594 CSoutput.n263 CSoutput.n165 4.5005
R6595 CSoutput.n263 CSoutput.n167 4.5005
R6596 CSoutput.n263 CSoutput.n164 4.5005
R6597 CSoutput.n263 CSoutput.n168 4.5005
R6598 CSoutput.n263 CSoutput.n163 4.5005
R6599 CSoutput.n263 CSoutput.t184 4.5005
R6600 CSoutput.n263 CSoutput.n162 4.5005
R6601 CSoutput.n263 CSoutput.n169 4.5005
R6602 CSoutput.n263 CSoutput.n170 4.5005
R6603 CSoutput.n261 CSoutput.n165 4.5005
R6604 CSoutput.n261 CSoutput.n167 4.5005
R6605 CSoutput.n261 CSoutput.n164 4.5005
R6606 CSoutput.n261 CSoutput.n168 4.5005
R6607 CSoutput.n261 CSoutput.n163 4.5005
R6608 CSoutput.n261 CSoutput.t184 4.5005
R6609 CSoutput.n261 CSoutput.n162 4.5005
R6610 CSoutput.n261 CSoutput.n169 4.5005
R6611 CSoutput.n259 CSoutput.n165 4.5005
R6612 CSoutput.n259 CSoutput.n167 4.5005
R6613 CSoutput.n259 CSoutput.n164 4.5005
R6614 CSoutput.n259 CSoutput.n168 4.5005
R6615 CSoutput.n259 CSoutput.n163 4.5005
R6616 CSoutput.n259 CSoutput.t184 4.5005
R6617 CSoutput.n259 CSoutput.n162 4.5005
R6618 CSoutput.n259 CSoutput.n169 4.5005
R6619 CSoutput.n189 CSoutput.n165 4.5005
R6620 CSoutput.n189 CSoutput.n167 4.5005
R6621 CSoutput.n189 CSoutput.n164 4.5005
R6622 CSoutput.n189 CSoutput.n168 4.5005
R6623 CSoutput.n189 CSoutput.n163 4.5005
R6624 CSoutput.n189 CSoutput.t184 4.5005
R6625 CSoutput.n189 CSoutput.n162 4.5005
R6626 CSoutput.n189 CSoutput.n169 4.5005
R6627 CSoutput.n189 CSoutput.n170 4.5005
R6628 CSoutput.n188 CSoutput.n165 4.5005
R6629 CSoutput.n188 CSoutput.n167 4.5005
R6630 CSoutput.n188 CSoutput.n164 4.5005
R6631 CSoutput.n188 CSoutput.n168 4.5005
R6632 CSoutput.n188 CSoutput.n163 4.5005
R6633 CSoutput.n188 CSoutput.t184 4.5005
R6634 CSoutput.n188 CSoutput.n162 4.5005
R6635 CSoutput.n188 CSoutput.n169 4.5005
R6636 CSoutput.n188 CSoutput.n170 4.5005
R6637 CSoutput.n192 CSoutput.n165 4.5005
R6638 CSoutput.n192 CSoutput.n167 4.5005
R6639 CSoutput.n192 CSoutput.n164 4.5005
R6640 CSoutput.n192 CSoutput.n168 4.5005
R6641 CSoutput.n192 CSoutput.n163 4.5005
R6642 CSoutput.n192 CSoutput.t184 4.5005
R6643 CSoutput.n192 CSoutput.n162 4.5005
R6644 CSoutput.n192 CSoutput.n169 4.5005
R6645 CSoutput.n192 CSoutput.n170 4.5005
R6646 CSoutput.n191 CSoutput.n165 4.5005
R6647 CSoutput.n191 CSoutput.n167 4.5005
R6648 CSoutput.n191 CSoutput.n164 4.5005
R6649 CSoutput.n191 CSoutput.n168 4.5005
R6650 CSoutput.n191 CSoutput.n163 4.5005
R6651 CSoutput.n191 CSoutput.t184 4.5005
R6652 CSoutput.n191 CSoutput.n162 4.5005
R6653 CSoutput.n191 CSoutput.n169 4.5005
R6654 CSoutput.n191 CSoutput.n170 4.5005
R6655 CSoutput.n174 CSoutput.n165 4.5005
R6656 CSoutput.n174 CSoutput.n167 4.5005
R6657 CSoutput.n174 CSoutput.n164 4.5005
R6658 CSoutput.n174 CSoutput.n168 4.5005
R6659 CSoutput.n174 CSoutput.n163 4.5005
R6660 CSoutput.n174 CSoutput.t184 4.5005
R6661 CSoutput.n174 CSoutput.n162 4.5005
R6662 CSoutput.n174 CSoutput.n169 4.5005
R6663 CSoutput.n174 CSoutput.n170 4.5005
R6664 CSoutput.n266 CSoutput.n165 4.5005
R6665 CSoutput.n266 CSoutput.n167 4.5005
R6666 CSoutput.n266 CSoutput.n164 4.5005
R6667 CSoutput.n266 CSoutput.n168 4.5005
R6668 CSoutput.n266 CSoutput.n163 4.5005
R6669 CSoutput.n266 CSoutput.t184 4.5005
R6670 CSoutput.n266 CSoutput.n162 4.5005
R6671 CSoutput.n266 CSoutput.n169 4.5005
R6672 CSoutput.n266 CSoutput.n170 4.5005
R6673 CSoutput.n253 CSoutput.n224 4.5005
R6674 CSoutput.n253 CSoutput.n230 4.5005
R6675 CSoutput.n211 CSoutput.n200 4.5005
R6676 CSoutput.n211 CSoutput.n202 4.5005
R6677 CSoutput.n211 CSoutput.n199 4.5005
R6678 CSoutput.n211 CSoutput.n203 4.5005
R6679 CSoutput.n211 CSoutput.n198 4.5005
R6680 CSoutput.n211 CSoutput.t186 4.5005
R6681 CSoutput.n211 CSoutput.n197 4.5005
R6682 CSoutput.n211 CSoutput.n204 4.5005
R6683 CSoutput.n253 CSoutput.n211 4.5005
R6684 CSoutput.n232 CSoutput.n200 4.5005
R6685 CSoutput.n232 CSoutput.n202 4.5005
R6686 CSoutput.n232 CSoutput.n199 4.5005
R6687 CSoutput.n232 CSoutput.n203 4.5005
R6688 CSoutput.n232 CSoutput.n198 4.5005
R6689 CSoutput.n232 CSoutput.t186 4.5005
R6690 CSoutput.n232 CSoutput.n197 4.5005
R6691 CSoutput.n232 CSoutput.n204 4.5005
R6692 CSoutput.n253 CSoutput.n232 4.5005
R6693 CSoutput.n210 CSoutput.n200 4.5005
R6694 CSoutput.n210 CSoutput.n202 4.5005
R6695 CSoutput.n210 CSoutput.n199 4.5005
R6696 CSoutput.n210 CSoutput.n203 4.5005
R6697 CSoutput.n210 CSoutput.n198 4.5005
R6698 CSoutput.n210 CSoutput.t186 4.5005
R6699 CSoutput.n210 CSoutput.n197 4.5005
R6700 CSoutput.n210 CSoutput.n204 4.5005
R6701 CSoutput.n253 CSoutput.n210 4.5005
R6702 CSoutput.n234 CSoutput.n200 4.5005
R6703 CSoutput.n234 CSoutput.n202 4.5005
R6704 CSoutput.n234 CSoutput.n199 4.5005
R6705 CSoutput.n234 CSoutput.n203 4.5005
R6706 CSoutput.n234 CSoutput.n198 4.5005
R6707 CSoutput.n234 CSoutput.t186 4.5005
R6708 CSoutput.n234 CSoutput.n197 4.5005
R6709 CSoutput.n234 CSoutput.n204 4.5005
R6710 CSoutput.n253 CSoutput.n234 4.5005
R6711 CSoutput.n200 CSoutput.n195 4.5005
R6712 CSoutput.n202 CSoutput.n195 4.5005
R6713 CSoutput.n199 CSoutput.n195 4.5005
R6714 CSoutput.n203 CSoutput.n195 4.5005
R6715 CSoutput.n198 CSoutput.n195 4.5005
R6716 CSoutput.t186 CSoutput.n195 4.5005
R6717 CSoutput.n197 CSoutput.n195 4.5005
R6718 CSoutput.n204 CSoutput.n195 4.5005
R6719 CSoutput.n256 CSoutput.n200 4.5005
R6720 CSoutput.n256 CSoutput.n202 4.5005
R6721 CSoutput.n256 CSoutput.n199 4.5005
R6722 CSoutput.n256 CSoutput.n203 4.5005
R6723 CSoutput.n256 CSoutput.n198 4.5005
R6724 CSoutput.n256 CSoutput.t186 4.5005
R6725 CSoutput.n256 CSoutput.n197 4.5005
R6726 CSoutput.n256 CSoutput.n204 4.5005
R6727 CSoutput.n254 CSoutput.n200 4.5005
R6728 CSoutput.n254 CSoutput.n202 4.5005
R6729 CSoutput.n254 CSoutput.n199 4.5005
R6730 CSoutput.n254 CSoutput.n203 4.5005
R6731 CSoutput.n254 CSoutput.n198 4.5005
R6732 CSoutput.n254 CSoutput.t186 4.5005
R6733 CSoutput.n254 CSoutput.n197 4.5005
R6734 CSoutput.n254 CSoutput.n204 4.5005
R6735 CSoutput.n254 CSoutput.n253 4.5005
R6736 CSoutput.n236 CSoutput.n200 4.5005
R6737 CSoutput.n236 CSoutput.n202 4.5005
R6738 CSoutput.n236 CSoutput.n199 4.5005
R6739 CSoutput.n236 CSoutput.n203 4.5005
R6740 CSoutput.n236 CSoutput.n198 4.5005
R6741 CSoutput.n236 CSoutput.t186 4.5005
R6742 CSoutput.n236 CSoutput.n197 4.5005
R6743 CSoutput.n236 CSoutput.n204 4.5005
R6744 CSoutput.n253 CSoutput.n236 4.5005
R6745 CSoutput.n208 CSoutput.n200 4.5005
R6746 CSoutput.n208 CSoutput.n202 4.5005
R6747 CSoutput.n208 CSoutput.n199 4.5005
R6748 CSoutput.n208 CSoutput.n203 4.5005
R6749 CSoutput.n208 CSoutput.n198 4.5005
R6750 CSoutput.n208 CSoutput.t186 4.5005
R6751 CSoutput.n208 CSoutput.n197 4.5005
R6752 CSoutput.n208 CSoutput.n204 4.5005
R6753 CSoutput.n253 CSoutput.n208 4.5005
R6754 CSoutput.n238 CSoutput.n200 4.5005
R6755 CSoutput.n238 CSoutput.n202 4.5005
R6756 CSoutput.n238 CSoutput.n199 4.5005
R6757 CSoutput.n238 CSoutput.n203 4.5005
R6758 CSoutput.n238 CSoutput.n198 4.5005
R6759 CSoutput.n238 CSoutput.t186 4.5005
R6760 CSoutput.n238 CSoutput.n197 4.5005
R6761 CSoutput.n238 CSoutput.n204 4.5005
R6762 CSoutput.n253 CSoutput.n238 4.5005
R6763 CSoutput.n207 CSoutput.n200 4.5005
R6764 CSoutput.n207 CSoutput.n202 4.5005
R6765 CSoutput.n207 CSoutput.n199 4.5005
R6766 CSoutput.n207 CSoutput.n203 4.5005
R6767 CSoutput.n207 CSoutput.n198 4.5005
R6768 CSoutput.n207 CSoutput.t186 4.5005
R6769 CSoutput.n207 CSoutput.n197 4.5005
R6770 CSoutput.n207 CSoutput.n204 4.5005
R6771 CSoutput.n253 CSoutput.n207 4.5005
R6772 CSoutput.n252 CSoutput.n200 4.5005
R6773 CSoutput.n252 CSoutput.n202 4.5005
R6774 CSoutput.n252 CSoutput.n199 4.5005
R6775 CSoutput.n252 CSoutput.n203 4.5005
R6776 CSoutput.n252 CSoutput.n198 4.5005
R6777 CSoutput.n252 CSoutput.t186 4.5005
R6778 CSoutput.n252 CSoutput.n197 4.5005
R6779 CSoutput.n252 CSoutput.n204 4.5005
R6780 CSoutput.n253 CSoutput.n252 4.5005
R6781 CSoutput.n251 CSoutput.n136 4.5005
R6782 CSoutput.n152 CSoutput.n136 4.5005
R6783 CSoutput.n147 CSoutput.n131 4.5005
R6784 CSoutput.n147 CSoutput.n133 4.5005
R6785 CSoutput.n147 CSoutput.n130 4.5005
R6786 CSoutput.n147 CSoutput.n134 4.5005
R6787 CSoutput.n147 CSoutput.n129 4.5005
R6788 CSoutput.n147 CSoutput.t187 4.5005
R6789 CSoutput.n147 CSoutput.n128 4.5005
R6790 CSoutput.n147 CSoutput.n135 4.5005
R6791 CSoutput.n147 CSoutput.n136 4.5005
R6792 CSoutput.n145 CSoutput.n131 4.5005
R6793 CSoutput.n145 CSoutput.n133 4.5005
R6794 CSoutput.n145 CSoutput.n130 4.5005
R6795 CSoutput.n145 CSoutput.n134 4.5005
R6796 CSoutput.n145 CSoutput.n129 4.5005
R6797 CSoutput.n145 CSoutput.t187 4.5005
R6798 CSoutput.n145 CSoutput.n128 4.5005
R6799 CSoutput.n145 CSoutput.n135 4.5005
R6800 CSoutput.n145 CSoutput.n136 4.5005
R6801 CSoutput.n144 CSoutput.n131 4.5005
R6802 CSoutput.n144 CSoutput.n133 4.5005
R6803 CSoutput.n144 CSoutput.n130 4.5005
R6804 CSoutput.n144 CSoutput.n134 4.5005
R6805 CSoutput.n144 CSoutput.n129 4.5005
R6806 CSoutput.n144 CSoutput.t187 4.5005
R6807 CSoutput.n144 CSoutput.n128 4.5005
R6808 CSoutput.n144 CSoutput.n135 4.5005
R6809 CSoutput.n144 CSoutput.n136 4.5005
R6810 CSoutput.n273 CSoutput.n131 4.5005
R6811 CSoutput.n273 CSoutput.n133 4.5005
R6812 CSoutput.n273 CSoutput.n130 4.5005
R6813 CSoutput.n273 CSoutput.n134 4.5005
R6814 CSoutput.n273 CSoutput.n129 4.5005
R6815 CSoutput.n273 CSoutput.t187 4.5005
R6816 CSoutput.n273 CSoutput.n128 4.5005
R6817 CSoutput.n273 CSoutput.n135 4.5005
R6818 CSoutput.n273 CSoutput.n136 4.5005
R6819 CSoutput.n271 CSoutput.n131 4.5005
R6820 CSoutput.n271 CSoutput.n133 4.5005
R6821 CSoutput.n271 CSoutput.n130 4.5005
R6822 CSoutput.n271 CSoutput.n134 4.5005
R6823 CSoutput.n271 CSoutput.n129 4.5005
R6824 CSoutput.n271 CSoutput.t187 4.5005
R6825 CSoutput.n271 CSoutput.n128 4.5005
R6826 CSoutput.n271 CSoutput.n135 4.5005
R6827 CSoutput.n269 CSoutput.n131 4.5005
R6828 CSoutput.n269 CSoutput.n133 4.5005
R6829 CSoutput.n269 CSoutput.n130 4.5005
R6830 CSoutput.n269 CSoutput.n134 4.5005
R6831 CSoutput.n269 CSoutput.n129 4.5005
R6832 CSoutput.n269 CSoutput.t187 4.5005
R6833 CSoutput.n269 CSoutput.n128 4.5005
R6834 CSoutput.n269 CSoutput.n135 4.5005
R6835 CSoutput.n155 CSoutput.n131 4.5005
R6836 CSoutput.n155 CSoutput.n133 4.5005
R6837 CSoutput.n155 CSoutput.n130 4.5005
R6838 CSoutput.n155 CSoutput.n134 4.5005
R6839 CSoutput.n155 CSoutput.n129 4.5005
R6840 CSoutput.n155 CSoutput.t187 4.5005
R6841 CSoutput.n155 CSoutput.n128 4.5005
R6842 CSoutput.n155 CSoutput.n135 4.5005
R6843 CSoutput.n155 CSoutput.n136 4.5005
R6844 CSoutput.n154 CSoutput.n131 4.5005
R6845 CSoutput.n154 CSoutput.n133 4.5005
R6846 CSoutput.n154 CSoutput.n130 4.5005
R6847 CSoutput.n154 CSoutput.n134 4.5005
R6848 CSoutput.n154 CSoutput.n129 4.5005
R6849 CSoutput.n154 CSoutput.t187 4.5005
R6850 CSoutput.n154 CSoutput.n128 4.5005
R6851 CSoutput.n154 CSoutput.n135 4.5005
R6852 CSoutput.n154 CSoutput.n136 4.5005
R6853 CSoutput.n158 CSoutput.n131 4.5005
R6854 CSoutput.n158 CSoutput.n133 4.5005
R6855 CSoutput.n158 CSoutput.n130 4.5005
R6856 CSoutput.n158 CSoutput.n134 4.5005
R6857 CSoutput.n158 CSoutput.n129 4.5005
R6858 CSoutput.n158 CSoutput.t187 4.5005
R6859 CSoutput.n158 CSoutput.n128 4.5005
R6860 CSoutput.n158 CSoutput.n135 4.5005
R6861 CSoutput.n158 CSoutput.n136 4.5005
R6862 CSoutput.n157 CSoutput.n131 4.5005
R6863 CSoutput.n157 CSoutput.n133 4.5005
R6864 CSoutput.n157 CSoutput.n130 4.5005
R6865 CSoutput.n157 CSoutput.n134 4.5005
R6866 CSoutput.n157 CSoutput.n129 4.5005
R6867 CSoutput.n157 CSoutput.t187 4.5005
R6868 CSoutput.n157 CSoutput.n128 4.5005
R6869 CSoutput.n157 CSoutput.n135 4.5005
R6870 CSoutput.n157 CSoutput.n136 4.5005
R6871 CSoutput.n140 CSoutput.n131 4.5005
R6872 CSoutput.n140 CSoutput.n133 4.5005
R6873 CSoutput.n140 CSoutput.n130 4.5005
R6874 CSoutput.n140 CSoutput.n134 4.5005
R6875 CSoutput.n140 CSoutput.n129 4.5005
R6876 CSoutput.n140 CSoutput.t187 4.5005
R6877 CSoutput.n140 CSoutput.n128 4.5005
R6878 CSoutput.n140 CSoutput.n135 4.5005
R6879 CSoutput.n140 CSoutput.n136 4.5005
R6880 CSoutput.n276 CSoutput.n131 4.5005
R6881 CSoutput.n276 CSoutput.n133 4.5005
R6882 CSoutput.n276 CSoutput.n130 4.5005
R6883 CSoutput.n276 CSoutput.n134 4.5005
R6884 CSoutput.n276 CSoutput.n129 4.5005
R6885 CSoutput.n276 CSoutput.t187 4.5005
R6886 CSoutput.n276 CSoutput.n128 4.5005
R6887 CSoutput.n276 CSoutput.n135 4.5005
R6888 CSoutput.n276 CSoutput.n136 4.5005
R6889 CSoutput.n323 CSoutput.n307 4.10845
R6890 CSoutput.n125 CSoutput.n109 4.10845
R6891 CSoutput.n321 CSoutput.t129 4.06363
R6892 CSoutput.n321 CSoutput.t147 4.06363
R6893 CSoutput.n319 CSoutput.t160 4.06363
R6894 CSoutput.n319 CSoutput.t91 4.06363
R6895 CSoutput.n317 CSoutput.t95 4.06363
R6896 CSoutput.n317 CSoutput.t151 4.06363
R6897 CSoutput.n315 CSoutput.t163 4.06363
R6898 CSoutput.n315 CSoutput.t164 4.06363
R6899 CSoutput.n313 CSoutput.t111 4.06363
R6900 CSoutput.n313 CSoutput.t112 4.06363
R6901 CSoutput.n311 CSoutput.t117 4.06363
R6902 CSoutput.n311 CSoutput.t165 4.06363
R6903 CSoutput.n309 CSoutput.t83 4.06363
R6904 CSoutput.n309 CSoutput.t115 4.06363
R6905 CSoutput.n308 CSoutput.t128 4.06363
R6906 CSoutput.n308 CSoutput.t146 4.06363
R6907 CSoutput.n305 CSoutput.t118 4.06363
R6908 CSoutput.n305 CSoutput.t138 4.06363
R6909 CSoutput.n303 CSoutput.t152 4.06363
R6910 CSoutput.n303 CSoutput.t79 4.06363
R6911 CSoutput.n301 CSoutput.t80 4.06363
R6912 CSoutput.n301 CSoutput.t140 4.06363
R6913 CSoutput.n299 CSoutput.t155 4.06363
R6914 CSoutput.n299 CSoutput.t156 4.06363
R6915 CSoutput.n297 CSoutput.t99 4.06363
R6916 CSoutput.n297 CSoutput.t100 4.06363
R6917 CSoutput.n295 CSoutput.t103 4.06363
R6918 CSoutput.n295 CSoutput.t157 4.06363
R6919 CSoutput.n293 CSoutput.t72 4.06363
R6920 CSoutput.n293 CSoutput.t102 4.06363
R6921 CSoutput.n292 CSoutput.t119 4.06363
R6922 CSoutput.n292 CSoutput.t139 4.06363
R6923 CSoutput.n290 CSoutput.t145 4.06363
R6924 CSoutput.n290 CSoutput.t108 4.06363
R6925 CSoutput.n288 CSoutput.t135 4.06363
R6926 CSoutput.n288 CSoutput.t90 4.06363
R6927 CSoutput.n286 CSoutput.t153 4.06363
R6928 CSoutput.n286 CSoutput.t84 4.06363
R6929 CSoutput.n284 CSoutput.t120 4.06363
R6930 CSoutput.n284 CSoutput.t101 4.06363
R6931 CSoutput.n282 CSoutput.t104 4.06363
R6932 CSoutput.n282 CSoutput.t81 4.06363
R6933 CSoutput.n280 CSoutput.t144 4.06363
R6934 CSoutput.n280 CSoutput.t76 4.06363
R6935 CSoutput.n278 CSoutput.t113 4.06363
R6936 CSoutput.n278 CSoutput.t161 4.06363
R6937 CSoutput.n277 CSoutput.t96 4.06363
R6938 CSoutput.n277 CSoutput.t149 4.06363
R6939 CSoutput.n110 CSoutput.t87 4.06363
R6940 CSoutput.n110 CSoutput.t158 4.06363
R6941 CSoutput.n111 CSoutput.t143 4.06363
R6942 CSoutput.n111 CSoutput.t125 4.06363
R6943 CSoutput.n113 CSoutput.t110 4.06363
R6944 CSoutput.n113 CSoutput.t167 4.06363
R6945 CSoutput.n115 CSoutput.t142 4.06363
R6946 CSoutput.n115 CSoutput.t141 4.06363
R6947 CSoutput.n117 CSoutput.t131 4.06363
R6948 CSoutput.n117 CSoutput.t107 4.06363
R6949 CSoutput.n119 CSoutput.t89 4.06363
R6950 CSoutput.n119 CSoutput.t132 4.06363
R6951 CSoutput.n121 CSoutput.t130 4.06363
R6952 CSoutput.n121 CSoutput.t105 4.06363
R6953 CSoutput.n123 CSoutput.t88 4.06363
R6954 CSoutput.n123 CSoutput.t86 4.06363
R6955 CSoutput.n94 CSoutput.t74 4.06363
R6956 CSoutput.n94 CSoutput.t148 4.06363
R6957 CSoutput.n95 CSoutput.t137 4.06363
R6958 CSoutput.n95 CSoutput.t116 4.06363
R6959 CSoutput.n97 CSoutput.t98 4.06363
R6960 CSoutput.n97 CSoutput.t159 4.06363
R6961 CSoutput.n99 CSoutput.t134 4.06363
R6962 CSoutput.n99 CSoutput.t133 4.06363
R6963 CSoutput.n101 CSoutput.t123 4.06363
R6964 CSoutput.n101 CSoutput.t94 4.06363
R6965 CSoutput.n103 CSoutput.t77 4.06363
R6966 CSoutput.n103 CSoutput.t124 4.06363
R6967 CSoutput.n105 CSoutput.t122 4.06363
R6968 CSoutput.n105 CSoutput.t92 4.06363
R6969 CSoutput.n107 CSoutput.t75 4.06363
R6970 CSoutput.n107 CSoutput.t73 4.06363
R6971 CSoutput.n79 CSoutput.t150 4.06363
R6972 CSoutput.n79 CSoutput.t97 4.06363
R6973 CSoutput.n80 CSoutput.t162 4.06363
R6974 CSoutput.n80 CSoutput.t114 4.06363
R6975 CSoutput.n82 CSoutput.t78 4.06363
R6976 CSoutput.n82 CSoutput.t126 4.06363
R6977 CSoutput.n84 CSoutput.t82 4.06363
R6978 CSoutput.n84 CSoutput.t106 4.06363
R6979 CSoutput.n86 CSoutput.t166 4.06363
R6980 CSoutput.n86 CSoutput.t121 4.06363
R6981 CSoutput.n88 CSoutput.t85 4.06363
R6982 CSoutput.n88 CSoutput.t154 4.06363
R6983 CSoutput.n90 CSoutput.t93 4.06363
R6984 CSoutput.n90 CSoutput.t136 4.06363
R6985 CSoutput.n92 CSoutput.t109 4.06363
R6986 CSoutput.n92 CSoutput.t127 4.06363
R6987 CSoutput.n44 CSoutput.n43 3.79402
R6988 CSoutput.n49 CSoutput.n48 3.79402
R6989 CSoutput.n404 CSoutput.n364 3.71319
R6990 CSoutput.n405 CSoutput.n404 3.57343
R6991 CSoutput.n361 CSoutput.t69 2.82907
R6992 CSoutput.n361 CSoutput.t43 2.82907
R6993 CSoutput.n359 CSoutput.t14 2.82907
R6994 CSoutput.n359 CSoutput.t30 2.82907
R6995 CSoutput.n357 CSoutput.t175 2.82907
R6996 CSoutput.n357 CSoutput.t172 2.82907
R6997 CSoutput.n355 CSoutput.t16 2.82907
R6998 CSoutput.n355 CSoutput.t2 2.82907
R6999 CSoutput.n353 CSoutput.t63 2.82907
R7000 CSoutput.n353 CSoutput.t3 2.82907
R7001 CSoutput.n351 CSoutput.t12 2.82907
R7002 CSoutput.n351 CSoutput.t26 2.82907
R7003 CSoutput.n349 CSoutput.t68 2.82907
R7004 CSoutput.n349 CSoutput.t55 2.82907
R7005 CSoutput.n347 CSoutput.t4 2.82907
R7006 CSoutput.n347 CSoutput.t38 2.82907
R7007 CSoutput.n345 CSoutput.t11 2.82907
R7008 CSoutput.n345 CSoutput.t171 2.82907
R7009 CSoutput.n344 CSoutput.t42 2.82907
R7010 CSoutput.n344 CSoutput.t13 2.82907
R7011 CSoutput.n342 CSoutput.t49 2.82907
R7012 CSoutput.n342 CSoutput.t20 2.82907
R7013 CSoutput.n340 CSoutput.t39 2.82907
R7014 CSoutput.n340 CSoutput.t50 2.82907
R7015 CSoutput.n338 CSoutput.t31 2.82907
R7016 CSoutput.n338 CSoutput.t34 2.82907
R7017 CSoutput.n336 CSoutput.t1 2.82907
R7018 CSoutput.n336 CSoutput.t21 2.82907
R7019 CSoutput.n334 CSoutput.t66 2.82907
R7020 CSoutput.n334 CSoutput.t173 2.82907
R7021 CSoutput.n332 CSoutput.t27 2.82907
R7022 CSoutput.n332 CSoutput.t71 2.82907
R7023 CSoutput.n330 CSoutput.t48 2.82907
R7024 CSoutput.n330 CSoutput.t174 2.82907
R7025 CSoutput.n328 CSoutput.t56 2.82907
R7026 CSoutput.n328 CSoutput.t61 2.82907
R7027 CSoutput.n326 CSoutput.t168 2.82907
R7028 CSoutput.n326 CSoutput.t41 2.82907
R7029 CSoutput.n325 CSoutput.t7 2.82907
R7030 CSoutput.n325 CSoutput.t18 2.82907
R7031 CSoutput.n384 CSoutput.t62 2.82907
R7032 CSoutput.n384 CSoutput.t22 2.82907
R7033 CSoutput.n385 CSoutput.t15 2.82907
R7034 CSoutput.n385 CSoutput.t23 2.82907
R7035 CSoutput.n387 CSoutput.t5 2.82907
R7036 CSoutput.n387 CSoutput.t37 2.82907
R7037 CSoutput.n389 CSoutput.t58 2.82907
R7038 CSoutput.n389 CSoutput.t52 2.82907
R7039 CSoutput.n391 CSoutput.t60 2.82907
R7040 CSoutput.n391 CSoutput.t25 2.82907
R7041 CSoutput.n393 CSoutput.t29 2.82907
R7042 CSoutput.n393 CSoutput.t169 2.82907
R7043 CSoutput.n395 CSoutput.t53 2.82907
R7044 CSoutput.n395 CSoutput.t170 2.82907
R7045 CSoutput.n397 CSoutput.t57 2.82907
R7046 CSoutput.n397 CSoutput.t65 2.82907
R7047 CSoutput.n399 CSoutput.t36 2.82907
R7048 CSoutput.n399 CSoutput.t19 2.82907
R7049 CSoutput.n401 CSoutput.t33 2.82907
R7050 CSoutput.n401 CSoutput.t64 2.82907
R7051 CSoutput.n365 CSoutput.t70 2.82907
R7052 CSoutput.n365 CSoutput.t10 2.82907
R7053 CSoutput.n366 CSoutput.t35 2.82907
R7054 CSoutput.n366 CSoutput.t45 2.82907
R7055 CSoutput.n368 CSoutput.t51 2.82907
R7056 CSoutput.n368 CSoutput.t44 2.82907
R7057 CSoutput.n370 CSoutput.t32 2.82907
R7058 CSoutput.n370 CSoutput.t67 2.82907
R7059 CSoutput.n372 CSoutput.t46 2.82907
R7060 CSoutput.n372 CSoutput.t8 2.82907
R7061 CSoutput.n374 CSoutput.t47 2.82907
R7062 CSoutput.n374 CSoutput.t54 2.82907
R7063 CSoutput.n376 CSoutput.t59 2.82907
R7064 CSoutput.n376 CSoutput.t24 2.82907
R7065 CSoutput.n378 CSoutput.t6 2.82907
R7066 CSoutput.n378 CSoutput.t40 2.82907
R7067 CSoutput.n380 CSoutput.t9 2.82907
R7068 CSoutput.n380 CSoutput.t28 2.82907
R7069 CSoutput.n382 CSoutput.t0 2.82907
R7070 CSoutput.n382 CSoutput.t17 2.82907
R7071 CSoutput.n324 CSoutput.n126 2.57547
R7072 CSoutput.n75 CSoutput.n1 2.45513
R7073 CSoutput.n217 CSoutput.n215 2.251
R7074 CSoutput.n217 CSoutput.n214 2.251
R7075 CSoutput.n217 CSoutput.n213 2.251
R7076 CSoutput.n217 CSoutput.n212 2.251
R7077 CSoutput.n186 CSoutput.n185 2.251
R7078 CSoutput.n186 CSoutput.n184 2.251
R7079 CSoutput.n186 CSoutput.n183 2.251
R7080 CSoutput.n186 CSoutput.n182 2.251
R7081 CSoutput.n259 CSoutput.n258 2.251
R7082 CSoutput.n224 CSoutput.n222 2.251
R7083 CSoutput.n224 CSoutput.n221 2.251
R7084 CSoutput.n224 CSoutput.n220 2.251
R7085 CSoutput.n242 CSoutput.n224 2.251
R7086 CSoutput.n230 CSoutput.n229 2.251
R7087 CSoutput.n230 CSoutput.n228 2.251
R7088 CSoutput.n230 CSoutput.n227 2.251
R7089 CSoutput.n230 CSoutput.n226 2.251
R7090 CSoutput.n256 CSoutput.n196 2.251
R7091 CSoutput.n251 CSoutput.n249 2.251
R7092 CSoutput.n251 CSoutput.n248 2.251
R7093 CSoutput.n251 CSoutput.n247 2.251
R7094 CSoutput.n251 CSoutput.n246 2.251
R7095 CSoutput.n152 CSoutput.n151 2.251
R7096 CSoutput.n152 CSoutput.n150 2.251
R7097 CSoutput.n152 CSoutput.n149 2.251
R7098 CSoutput.n152 CSoutput.n148 2.251
R7099 CSoutput.n269 CSoutput.n268 2.251
R7100 CSoutput.n186 CSoutput.n166 2.2505
R7101 CSoutput.n181 CSoutput.n166 2.2505
R7102 CSoutput.n179 CSoutput.n166 2.2505
R7103 CSoutput.n178 CSoutput.n166 2.2505
R7104 CSoutput.n263 CSoutput.n166 2.2505
R7105 CSoutput.n261 CSoutput.n166 2.2505
R7106 CSoutput.n259 CSoutput.n166 2.2505
R7107 CSoutput.n189 CSoutput.n166 2.2505
R7108 CSoutput.n188 CSoutput.n166 2.2505
R7109 CSoutput.n192 CSoutput.n166 2.2505
R7110 CSoutput.n191 CSoutput.n166 2.2505
R7111 CSoutput.n174 CSoutput.n166 2.2505
R7112 CSoutput.n266 CSoutput.n166 2.2505
R7113 CSoutput.n266 CSoutput.n265 2.2505
R7114 CSoutput.n230 CSoutput.n201 2.2505
R7115 CSoutput.n211 CSoutput.n201 2.2505
R7116 CSoutput.n232 CSoutput.n201 2.2505
R7117 CSoutput.n210 CSoutput.n201 2.2505
R7118 CSoutput.n234 CSoutput.n201 2.2505
R7119 CSoutput.n201 CSoutput.n195 2.2505
R7120 CSoutput.n256 CSoutput.n201 2.2505
R7121 CSoutput.n254 CSoutput.n201 2.2505
R7122 CSoutput.n236 CSoutput.n201 2.2505
R7123 CSoutput.n208 CSoutput.n201 2.2505
R7124 CSoutput.n238 CSoutput.n201 2.2505
R7125 CSoutput.n207 CSoutput.n201 2.2505
R7126 CSoutput.n252 CSoutput.n201 2.2505
R7127 CSoutput.n252 CSoutput.n205 2.2505
R7128 CSoutput.n152 CSoutput.n132 2.2505
R7129 CSoutput.n147 CSoutput.n132 2.2505
R7130 CSoutput.n145 CSoutput.n132 2.2505
R7131 CSoutput.n144 CSoutput.n132 2.2505
R7132 CSoutput.n273 CSoutput.n132 2.2505
R7133 CSoutput.n271 CSoutput.n132 2.2505
R7134 CSoutput.n269 CSoutput.n132 2.2505
R7135 CSoutput.n155 CSoutput.n132 2.2505
R7136 CSoutput.n154 CSoutput.n132 2.2505
R7137 CSoutput.n158 CSoutput.n132 2.2505
R7138 CSoutput.n157 CSoutput.n132 2.2505
R7139 CSoutput.n140 CSoutput.n132 2.2505
R7140 CSoutput.n276 CSoutput.n132 2.2505
R7141 CSoutput.n276 CSoutput.n275 2.2505
R7142 CSoutput.n194 CSoutput.n187 2.25024
R7143 CSoutput.n194 CSoutput.n180 2.25024
R7144 CSoutput.n262 CSoutput.n194 2.25024
R7145 CSoutput.n194 CSoutput.n190 2.25024
R7146 CSoutput.n194 CSoutput.n193 2.25024
R7147 CSoutput.n194 CSoutput.n161 2.25024
R7148 CSoutput.n244 CSoutput.n241 2.25024
R7149 CSoutput.n244 CSoutput.n240 2.25024
R7150 CSoutput.n244 CSoutput.n239 2.25024
R7151 CSoutput.n244 CSoutput.n206 2.25024
R7152 CSoutput.n244 CSoutput.n243 2.25024
R7153 CSoutput.n245 CSoutput.n244 2.25024
R7154 CSoutput.n160 CSoutput.n153 2.25024
R7155 CSoutput.n160 CSoutput.n146 2.25024
R7156 CSoutput.n272 CSoutput.n160 2.25024
R7157 CSoutput.n160 CSoutput.n156 2.25024
R7158 CSoutput.n160 CSoutput.n159 2.25024
R7159 CSoutput.n160 CSoutput.n127 2.25024
R7160 CSoutput.n261 CSoutput.n171 1.50111
R7161 CSoutput.n209 CSoutput.n195 1.50111
R7162 CSoutput.n271 CSoutput.n137 1.50111
R7163 CSoutput.n217 CSoutput.n216 1.501
R7164 CSoutput.n224 CSoutput.n223 1.501
R7165 CSoutput.n251 CSoutput.n250 1.501
R7166 CSoutput.n265 CSoutput.n176 1.12536
R7167 CSoutput.n265 CSoutput.n177 1.12536
R7168 CSoutput.n265 CSoutput.n264 1.12536
R7169 CSoutput.n225 CSoutput.n205 1.12536
R7170 CSoutput.n231 CSoutput.n205 1.12536
R7171 CSoutput.n233 CSoutput.n205 1.12536
R7172 CSoutput.n275 CSoutput.n142 1.12536
R7173 CSoutput.n275 CSoutput.n143 1.12536
R7174 CSoutput.n275 CSoutput.n274 1.12536
R7175 CSoutput.n265 CSoutput.n172 1.12536
R7176 CSoutput.n265 CSoutput.n173 1.12536
R7177 CSoutput.n265 CSoutput.n175 1.12536
R7178 CSoutput.n255 CSoutput.n205 1.12536
R7179 CSoutput.n235 CSoutput.n205 1.12536
R7180 CSoutput.n237 CSoutput.n205 1.12536
R7181 CSoutput.n275 CSoutput.n138 1.12536
R7182 CSoutput.n275 CSoutput.n139 1.12536
R7183 CSoutput.n275 CSoutput.n141 1.12536
R7184 CSoutput.n31 CSoutput.n30 0.669944
R7185 CSoutput.n62 CSoutput.n61 0.669944
R7186 CSoutput.n348 CSoutput.n346 0.573776
R7187 CSoutput.n350 CSoutput.n348 0.573776
R7188 CSoutput.n352 CSoutput.n350 0.573776
R7189 CSoutput.n354 CSoutput.n352 0.573776
R7190 CSoutput.n356 CSoutput.n354 0.573776
R7191 CSoutput.n358 CSoutput.n356 0.573776
R7192 CSoutput.n360 CSoutput.n358 0.573776
R7193 CSoutput.n362 CSoutput.n360 0.573776
R7194 CSoutput.n329 CSoutput.n327 0.573776
R7195 CSoutput.n331 CSoutput.n329 0.573776
R7196 CSoutput.n333 CSoutput.n331 0.573776
R7197 CSoutput.n335 CSoutput.n333 0.573776
R7198 CSoutput.n337 CSoutput.n335 0.573776
R7199 CSoutput.n339 CSoutput.n337 0.573776
R7200 CSoutput.n341 CSoutput.n339 0.573776
R7201 CSoutput.n343 CSoutput.n341 0.573776
R7202 CSoutput.n402 CSoutput.n400 0.573776
R7203 CSoutput.n400 CSoutput.n398 0.573776
R7204 CSoutput.n398 CSoutput.n396 0.573776
R7205 CSoutput.n396 CSoutput.n394 0.573776
R7206 CSoutput.n394 CSoutput.n392 0.573776
R7207 CSoutput.n392 CSoutput.n390 0.573776
R7208 CSoutput.n390 CSoutput.n388 0.573776
R7209 CSoutput.n388 CSoutput.n386 0.573776
R7210 CSoutput.n383 CSoutput.n381 0.573776
R7211 CSoutput.n381 CSoutput.n379 0.573776
R7212 CSoutput.n379 CSoutput.n377 0.573776
R7213 CSoutput.n377 CSoutput.n375 0.573776
R7214 CSoutput.n375 CSoutput.n373 0.573776
R7215 CSoutput.n373 CSoutput.n371 0.573776
R7216 CSoutput.n371 CSoutput.n369 0.573776
R7217 CSoutput.n369 CSoutput.n367 0.573776
R7218 CSoutput.n405 CSoutput.n276 0.53442
R7219 CSoutput.n312 CSoutput.n310 0.358259
R7220 CSoutput.n314 CSoutput.n312 0.358259
R7221 CSoutput.n316 CSoutput.n314 0.358259
R7222 CSoutput.n318 CSoutput.n316 0.358259
R7223 CSoutput.n320 CSoutput.n318 0.358259
R7224 CSoutput.n322 CSoutput.n320 0.358259
R7225 CSoutput.n296 CSoutput.n294 0.358259
R7226 CSoutput.n298 CSoutput.n296 0.358259
R7227 CSoutput.n300 CSoutput.n298 0.358259
R7228 CSoutput.n302 CSoutput.n300 0.358259
R7229 CSoutput.n304 CSoutput.n302 0.358259
R7230 CSoutput.n306 CSoutput.n304 0.358259
R7231 CSoutput.n281 CSoutput.n279 0.358259
R7232 CSoutput.n283 CSoutput.n281 0.358259
R7233 CSoutput.n285 CSoutput.n283 0.358259
R7234 CSoutput.n287 CSoutput.n285 0.358259
R7235 CSoutput.n289 CSoutput.n287 0.358259
R7236 CSoutput.n291 CSoutput.n289 0.358259
R7237 CSoutput.n124 CSoutput.n122 0.358259
R7238 CSoutput.n122 CSoutput.n120 0.358259
R7239 CSoutput.n120 CSoutput.n118 0.358259
R7240 CSoutput.n118 CSoutput.n116 0.358259
R7241 CSoutput.n116 CSoutput.n114 0.358259
R7242 CSoutput.n114 CSoutput.n112 0.358259
R7243 CSoutput.n108 CSoutput.n106 0.358259
R7244 CSoutput.n106 CSoutput.n104 0.358259
R7245 CSoutput.n104 CSoutput.n102 0.358259
R7246 CSoutput.n102 CSoutput.n100 0.358259
R7247 CSoutput.n100 CSoutput.n98 0.358259
R7248 CSoutput.n98 CSoutput.n96 0.358259
R7249 CSoutput.n93 CSoutput.n91 0.358259
R7250 CSoutput.n91 CSoutput.n89 0.358259
R7251 CSoutput.n89 CSoutput.n87 0.358259
R7252 CSoutput.n87 CSoutput.n85 0.358259
R7253 CSoutput.n85 CSoutput.n83 0.358259
R7254 CSoutput.n83 CSoutput.n81 0.358259
R7255 CSoutput.n21 CSoutput.n20 0.169105
R7256 CSoutput.n21 CSoutput.n16 0.169105
R7257 CSoutput.n26 CSoutput.n16 0.169105
R7258 CSoutput.n27 CSoutput.n26 0.169105
R7259 CSoutput.n27 CSoutput.n14 0.169105
R7260 CSoutput.n32 CSoutput.n14 0.169105
R7261 CSoutput.n33 CSoutput.n32 0.169105
R7262 CSoutput.n34 CSoutput.n33 0.169105
R7263 CSoutput.n34 CSoutput.n12 0.169105
R7264 CSoutput.n39 CSoutput.n12 0.169105
R7265 CSoutput.n40 CSoutput.n39 0.169105
R7266 CSoutput.n40 CSoutput.n10 0.169105
R7267 CSoutput.n45 CSoutput.n10 0.169105
R7268 CSoutput.n46 CSoutput.n45 0.169105
R7269 CSoutput.n47 CSoutput.n46 0.169105
R7270 CSoutput.n47 CSoutput.n8 0.169105
R7271 CSoutput.n52 CSoutput.n8 0.169105
R7272 CSoutput.n53 CSoutput.n52 0.169105
R7273 CSoutput.n53 CSoutput.n6 0.169105
R7274 CSoutput.n58 CSoutput.n6 0.169105
R7275 CSoutput.n59 CSoutput.n58 0.169105
R7276 CSoutput.n60 CSoutput.n59 0.169105
R7277 CSoutput.n60 CSoutput.n4 0.169105
R7278 CSoutput.n66 CSoutput.n4 0.169105
R7279 CSoutput.n67 CSoutput.n66 0.169105
R7280 CSoutput.n68 CSoutput.n67 0.169105
R7281 CSoutput.n68 CSoutput.n2 0.169105
R7282 CSoutput.n73 CSoutput.n2 0.169105
R7283 CSoutput.n74 CSoutput.n73 0.169105
R7284 CSoutput.n74 CSoutput.n0 0.169105
R7285 CSoutput.n78 CSoutput.n0 0.169105
R7286 CSoutput.n219 CSoutput.n218 0.0910737
R7287 CSoutput.n270 CSoutput.n267 0.0723685
R7288 CSoutput.n224 CSoutput.n219 0.0522944
R7289 CSoutput.n267 CSoutput.n266 0.0499135
R7290 CSoutput.n218 CSoutput.n217 0.0499135
R7291 CSoutput.n252 CSoutput.n251 0.0464294
R7292 CSoutput.n260 CSoutput.n257 0.0391444
R7293 CSoutput.n219 CSoutput.t192 0.023435
R7294 CSoutput.n267 CSoutput.t181 0.02262
R7295 CSoutput.n218 CSoutput.t190 0.02262
R7296 CSoutput CSoutput.n405 0.0052
R7297 CSoutput.n189 CSoutput.n172 0.00365111
R7298 CSoutput.n192 CSoutput.n173 0.00365111
R7299 CSoutput.n175 CSoutput.n174 0.00365111
R7300 CSoutput.n217 CSoutput.n176 0.00365111
R7301 CSoutput.n181 CSoutput.n177 0.00365111
R7302 CSoutput.n264 CSoutput.n178 0.00365111
R7303 CSoutput.n255 CSoutput.n254 0.00365111
R7304 CSoutput.n235 CSoutput.n208 0.00365111
R7305 CSoutput.n237 CSoutput.n207 0.00365111
R7306 CSoutput.n225 CSoutput.n224 0.00365111
R7307 CSoutput.n231 CSoutput.n211 0.00365111
R7308 CSoutput.n233 CSoutput.n210 0.00365111
R7309 CSoutput.n155 CSoutput.n138 0.00365111
R7310 CSoutput.n158 CSoutput.n139 0.00365111
R7311 CSoutput.n141 CSoutput.n140 0.00365111
R7312 CSoutput.n251 CSoutput.n142 0.00365111
R7313 CSoutput.n147 CSoutput.n143 0.00365111
R7314 CSoutput.n274 CSoutput.n144 0.00365111
R7315 CSoutput.n186 CSoutput.n176 0.00340054
R7316 CSoutput.n179 CSoutput.n177 0.00340054
R7317 CSoutput.n264 CSoutput.n263 0.00340054
R7318 CSoutput.n259 CSoutput.n172 0.00340054
R7319 CSoutput.n188 CSoutput.n173 0.00340054
R7320 CSoutput.n191 CSoutput.n175 0.00340054
R7321 CSoutput.n230 CSoutput.n225 0.00340054
R7322 CSoutput.n232 CSoutput.n231 0.00340054
R7323 CSoutput.n234 CSoutput.n233 0.00340054
R7324 CSoutput.n256 CSoutput.n255 0.00340054
R7325 CSoutput.n236 CSoutput.n235 0.00340054
R7326 CSoutput.n238 CSoutput.n237 0.00340054
R7327 CSoutput.n152 CSoutput.n142 0.00340054
R7328 CSoutput.n145 CSoutput.n143 0.00340054
R7329 CSoutput.n274 CSoutput.n273 0.00340054
R7330 CSoutput.n269 CSoutput.n138 0.00340054
R7331 CSoutput.n154 CSoutput.n139 0.00340054
R7332 CSoutput.n157 CSoutput.n141 0.00340054
R7333 CSoutput.n187 CSoutput.n181 0.00252698
R7334 CSoutput.n180 CSoutput.n178 0.00252698
R7335 CSoutput.n262 CSoutput.n261 0.00252698
R7336 CSoutput.n190 CSoutput.n188 0.00252698
R7337 CSoutput.n193 CSoutput.n191 0.00252698
R7338 CSoutput.n266 CSoutput.n161 0.00252698
R7339 CSoutput.n187 CSoutput.n186 0.00252698
R7340 CSoutput.n180 CSoutput.n179 0.00252698
R7341 CSoutput.n263 CSoutput.n262 0.00252698
R7342 CSoutput.n190 CSoutput.n189 0.00252698
R7343 CSoutput.n193 CSoutput.n192 0.00252698
R7344 CSoutput.n174 CSoutput.n161 0.00252698
R7345 CSoutput.n241 CSoutput.n211 0.00252698
R7346 CSoutput.n240 CSoutput.n210 0.00252698
R7347 CSoutput.n239 CSoutput.n195 0.00252698
R7348 CSoutput.n236 CSoutput.n206 0.00252698
R7349 CSoutput.n243 CSoutput.n238 0.00252698
R7350 CSoutput.n252 CSoutput.n245 0.00252698
R7351 CSoutput.n241 CSoutput.n230 0.00252698
R7352 CSoutput.n240 CSoutput.n232 0.00252698
R7353 CSoutput.n239 CSoutput.n234 0.00252698
R7354 CSoutput.n254 CSoutput.n206 0.00252698
R7355 CSoutput.n243 CSoutput.n208 0.00252698
R7356 CSoutput.n245 CSoutput.n207 0.00252698
R7357 CSoutput.n153 CSoutput.n147 0.00252698
R7358 CSoutput.n146 CSoutput.n144 0.00252698
R7359 CSoutput.n272 CSoutput.n271 0.00252698
R7360 CSoutput.n156 CSoutput.n154 0.00252698
R7361 CSoutput.n159 CSoutput.n157 0.00252698
R7362 CSoutput.n276 CSoutput.n127 0.00252698
R7363 CSoutput.n153 CSoutput.n152 0.00252698
R7364 CSoutput.n146 CSoutput.n145 0.00252698
R7365 CSoutput.n273 CSoutput.n272 0.00252698
R7366 CSoutput.n156 CSoutput.n155 0.00252698
R7367 CSoutput.n159 CSoutput.n158 0.00252698
R7368 CSoutput.n140 CSoutput.n127 0.00252698
R7369 CSoutput.n261 CSoutput.n260 0.0020275
R7370 CSoutput.n260 CSoutput.n259 0.0020275
R7371 CSoutput.n257 CSoutput.n195 0.0020275
R7372 CSoutput.n257 CSoutput.n256 0.0020275
R7373 CSoutput.n271 CSoutput.n270 0.0020275
R7374 CSoutput.n270 CSoutput.n269 0.0020275
R7375 CSoutput.n171 CSoutput.n170 0.00166668
R7376 CSoutput.n253 CSoutput.n209 0.00166668
R7377 CSoutput.n137 CSoutput.n136 0.00166668
R7378 CSoutput.n275 CSoutput.n137 0.00133328
R7379 CSoutput.n209 CSoutput.n205 0.00133328
R7380 CSoutput.n265 CSoutput.n171 0.00133328
R7381 CSoutput.n268 CSoutput.n160 0.001
R7382 CSoutput.n246 CSoutput.n160 0.001
R7383 CSoutput.n148 CSoutput.n128 0.001
R7384 CSoutput.n247 CSoutput.n128 0.001
R7385 CSoutput.n149 CSoutput.n129 0.001
R7386 CSoutput.n248 CSoutput.n129 0.001
R7387 CSoutput.n150 CSoutput.n130 0.001
R7388 CSoutput.n249 CSoutput.n130 0.001
R7389 CSoutput.n151 CSoutput.n131 0.001
R7390 CSoutput.n250 CSoutput.n131 0.001
R7391 CSoutput.n244 CSoutput.n196 0.001
R7392 CSoutput.n244 CSoutput.n242 0.001
R7393 CSoutput.n226 CSoutput.n197 0.001
R7394 CSoutput.n220 CSoutput.n197 0.001
R7395 CSoutput.n227 CSoutput.n198 0.001
R7396 CSoutput.n221 CSoutput.n198 0.001
R7397 CSoutput.n228 CSoutput.n199 0.001
R7398 CSoutput.n222 CSoutput.n199 0.001
R7399 CSoutput.n229 CSoutput.n200 0.001
R7400 CSoutput.n223 CSoutput.n200 0.001
R7401 CSoutput.n258 CSoutput.n194 0.001
R7402 CSoutput.n212 CSoutput.n194 0.001
R7403 CSoutput.n182 CSoutput.n162 0.001
R7404 CSoutput.n213 CSoutput.n162 0.001
R7405 CSoutput.n183 CSoutput.n163 0.001
R7406 CSoutput.n214 CSoutput.n163 0.001
R7407 CSoutput.n184 CSoutput.n164 0.001
R7408 CSoutput.n215 CSoutput.n164 0.001
R7409 CSoutput.n185 CSoutput.n165 0.001
R7410 CSoutput.n216 CSoutput.n165 0.001
R7411 CSoutput.n216 CSoutput.n166 0.001
R7412 CSoutput.n215 CSoutput.n167 0.001
R7413 CSoutput.n214 CSoutput.n168 0.001
R7414 CSoutput.n213 CSoutput.t184 0.001
R7415 CSoutput.n212 CSoutput.n169 0.001
R7416 CSoutput.n185 CSoutput.n167 0.001
R7417 CSoutput.n184 CSoutput.n168 0.001
R7418 CSoutput.n183 CSoutput.t184 0.001
R7419 CSoutput.n182 CSoutput.n169 0.001
R7420 CSoutput.n258 CSoutput.n170 0.001
R7421 CSoutput.n223 CSoutput.n201 0.001
R7422 CSoutput.n222 CSoutput.n202 0.001
R7423 CSoutput.n221 CSoutput.n203 0.001
R7424 CSoutput.n220 CSoutput.t186 0.001
R7425 CSoutput.n242 CSoutput.n204 0.001
R7426 CSoutput.n229 CSoutput.n202 0.001
R7427 CSoutput.n228 CSoutput.n203 0.001
R7428 CSoutput.n227 CSoutput.t186 0.001
R7429 CSoutput.n226 CSoutput.n204 0.001
R7430 CSoutput.n253 CSoutput.n196 0.001
R7431 CSoutput.n250 CSoutput.n132 0.001
R7432 CSoutput.n249 CSoutput.n133 0.001
R7433 CSoutput.n248 CSoutput.n134 0.001
R7434 CSoutput.n247 CSoutput.t187 0.001
R7435 CSoutput.n246 CSoutput.n135 0.001
R7436 CSoutput.n151 CSoutput.n133 0.001
R7437 CSoutput.n150 CSoutput.n134 0.001
R7438 CSoutput.n149 CSoutput.t187 0.001
R7439 CSoutput.n148 CSoutput.n135 0.001
R7440 CSoutput.n268 CSoutput.n136 0.001
R7441 a_n2318_13878.n59 a_n2318_13878.t28 533.335
R7442 a_n2318_13878.n115 a_n2318_13878.t22 512.366
R7443 a_n2318_13878.n65 a_n2318_13878.t26 512.366
R7444 a_n2318_13878.n114 a_n2318_13878.t4 512.366
R7445 a_n2318_13878.n113 a_n2318_13878.t14 512.366
R7446 a_n2318_13878.n66 a_n2318_13878.t32 512.366
R7447 a_n2318_13878.n112 a_n2318_13878.t24 512.366
R7448 a_n2318_13878.n53 a_n2318_13878.t82 533.335
R7449 a_n2318_13878.n101 a_n2318_13878.t63 512.366
R7450 a_n2318_13878.n67 a_n2318_13878.t67 512.366
R7451 a_n2318_13878.n100 a_n2318_13878.t57 512.366
R7452 a_n2318_13878.n99 a_n2318_13878.t72 512.366
R7453 a_n2318_13878.n68 a_n2318_13878.t79 512.366
R7454 a_n2318_13878.n98 a_n2318_13878.t80 512.366
R7455 a_n2318_13878.n38 a_n2318_13878.t8 533.335
R7456 a_n2318_13878.n79 a_n2318_13878.t20 512.366
R7457 a_n2318_13878.n80 a_n2318_13878.t30 512.366
R7458 a_n2318_13878.n81 a_n2318_13878.t10 512.366
R7459 a_n2318_13878.n82 a_n2318_13878.t6 512.366
R7460 a_n2318_13878.n72 a_n2318_13878.t12 512.366
R7461 a_n2318_13878.n83 a_n2318_13878.t34 512.366
R7462 a_n2318_13878.n31 a_n2318_13878.t78 533.335
R7463 a_n2318_13878.n74 a_n2318_13878.t56 512.366
R7464 a_n2318_13878.n75 a_n2318_13878.t75 512.366
R7465 a_n2318_13878.n76 a_n2318_13878.t76 512.366
R7466 a_n2318_13878.n77 a_n2318_13878.t53 512.366
R7467 a_n2318_13878.n73 a_n2318_13878.t62 512.366
R7468 a_n2318_13878.n78 a_n2318_13878.t71 512.366
R7469 a_n2318_13878.n95 a_n2318_13878.t69 512.366
R7470 a_n2318_13878.n85 a_n2318_13878.t60 512.366
R7471 a_n2318_13878.n96 a_n2318_13878.t52 512.366
R7472 a_n2318_13878.n93 a_n2318_13878.t77 512.366
R7473 a_n2318_13878.n86 a_n2318_13878.t66 512.366
R7474 a_n2318_13878.n94 a_n2318_13878.t65 512.366
R7475 a_n2318_13878.n91 a_n2318_13878.t73 512.366
R7476 a_n2318_13878.n87 a_n2318_13878.t58 512.366
R7477 a_n2318_13878.n92 a_n2318_13878.t59 512.366
R7478 a_n2318_13878.n89 a_n2318_13878.t61 512.366
R7479 a_n2318_13878.n88 a_n2318_13878.t70 512.366
R7480 a_n2318_13878.n90 a_n2318_13878.t83 512.366
R7481 a_n2318_13878.n64 a_n2318_13878.n1 70.1674
R7482 a_n2318_13878.n58 a_n2318_13878.n5 70.1674
R7483 a_n2318_13878.n17 a_n2318_13878.n44 70.1674
R7484 a_n2318_13878.n20 a_n2318_13878.n37 70.1674
R7485 a_n2318_13878.n78 a_n2318_13878.n37 20.9683
R7486 a_n2318_13878.n36 a_n2318_13878.n21 72.3034
R7487 a_n2318_13878.n36 a_n2318_13878.n73 16.6962
R7488 a_n2318_13878.n21 a_n2318_13878.n35 77.6622
R7489 a_n2318_13878.n77 a_n2318_13878.n35 5.97853
R7490 a_n2318_13878.n34 a_n2318_13878.n22 77.6622
R7491 a_n2318_13878.n22 a_n2318_13878.n33 72.3034
R7492 a_n2318_13878.n74 a_n2318_13878.n31 20.9683
R7493 a_n2318_13878.n32 a_n2318_13878.n31 70.1674
R7494 a_n2318_13878.n83 a_n2318_13878.n44 20.9683
R7495 a_n2318_13878.n43 a_n2318_13878.n18 72.3034
R7496 a_n2318_13878.n43 a_n2318_13878.n72 16.6962
R7497 a_n2318_13878.n18 a_n2318_13878.n42 77.6622
R7498 a_n2318_13878.n82 a_n2318_13878.n42 5.97853
R7499 a_n2318_13878.n41 a_n2318_13878.n19 77.6622
R7500 a_n2318_13878.n19 a_n2318_13878.n40 72.3034
R7501 a_n2318_13878.n79 a_n2318_13878.n38 20.9683
R7502 a_n2318_13878.n39 a_n2318_13878.n38 70.1674
R7503 a_n2318_13878.n8 a_n2318_13878.n52 70.1674
R7504 a_n2318_13878.n10 a_n2318_13878.n50 70.1674
R7505 a_n2318_13878.n12 a_n2318_13878.n48 70.1674
R7506 a_n2318_13878.n15 a_n2318_13878.n46 70.1674
R7507 a_n2318_13878.n90 a_n2318_13878.n46 20.9683
R7508 a_n2318_13878.n45 a_n2318_13878.n16 75.0448
R7509 a_n2318_13878.n45 a_n2318_13878.n88 11.2134
R7510 a_n2318_13878.n16 a_n2318_13878.n89 161.3
R7511 a_n2318_13878.n92 a_n2318_13878.n48 20.9683
R7512 a_n2318_13878.n47 a_n2318_13878.n13 75.0448
R7513 a_n2318_13878.n47 a_n2318_13878.n87 11.2134
R7514 a_n2318_13878.n13 a_n2318_13878.n91 161.3
R7515 a_n2318_13878.n94 a_n2318_13878.n50 20.9683
R7516 a_n2318_13878.n49 a_n2318_13878.n11 75.0448
R7517 a_n2318_13878.n49 a_n2318_13878.n86 11.2134
R7518 a_n2318_13878.n11 a_n2318_13878.n93 161.3
R7519 a_n2318_13878.n96 a_n2318_13878.n52 20.9683
R7520 a_n2318_13878.n51 a_n2318_13878.n9 75.0448
R7521 a_n2318_13878.n51 a_n2318_13878.n85 11.2134
R7522 a_n2318_13878.n9 a_n2318_13878.n95 161.3
R7523 a_n2318_13878.n98 a_n2318_13878.n58 20.9683
R7524 a_n2318_13878.n6 a_n2318_13878.n57 72.3034
R7525 a_n2318_13878.n57 a_n2318_13878.n68 16.6962
R7526 a_n2318_13878.n56 a_n2318_13878.n6 77.6622
R7527 a_n2318_13878.n99 a_n2318_13878.n56 5.97853
R7528 a_n2318_13878.n55 a_n2318_13878.n4 77.6622
R7529 a_n2318_13878.n4 a_n2318_13878.n54 72.3034
R7530 a_n2318_13878.n101 a_n2318_13878.n53 20.9683
R7531 a_n2318_13878.n7 a_n2318_13878.n53 70.1674
R7532 a_n2318_13878.n112 a_n2318_13878.n64 20.9683
R7533 a_n2318_13878.n2 a_n2318_13878.n63 72.3034
R7534 a_n2318_13878.n63 a_n2318_13878.n66 16.6962
R7535 a_n2318_13878.n62 a_n2318_13878.n2 77.6622
R7536 a_n2318_13878.n113 a_n2318_13878.n62 5.97853
R7537 a_n2318_13878.n61 a_n2318_13878.n0 77.6622
R7538 a_n2318_13878.n0 a_n2318_13878.n60 72.3034
R7539 a_n2318_13878.n115 a_n2318_13878.n59 20.9683
R7540 a_n2318_13878.n3 a_n2318_13878.n59 70.1674
R7541 a_n2318_13878.n26 a_n2318_13878.n110 81.2902
R7542 a_n2318_13878.n24 a_n2318_13878.n105 81.2902
R7543 a_n2318_13878.n23 a_n2318_13878.n102 81.2902
R7544 a_n2318_13878.n26 a_n2318_13878.n111 80.9324
R7545 a_n2318_13878.n26 a_n2318_13878.n109 80.9324
R7546 a_n2318_13878.n25 a_n2318_13878.n108 80.9324
R7547 a_n2318_13878.n25 a_n2318_13878.n107 80.9324
R7548 a_n2318_13878.n24 a_n2318_13878.n106 80.9324
R7549 a_n2318_13878.n24 a_n2318_13878.n104 80.9324
R7550 a_n2318_13878.n23 a_n2318_13878.n103 80.9324
R7551 a_n2318_13878.n30 a_n2318_13878.t17 74.6477
R7552 a_n2318_13878.n27 a_n2318_13878.t9 74.6477
R7553 a_n2318_13878.n29 a_n2318_13878.t29 74.2899
R7554 a_n2318_13878.n28 a_n2318_13878.t19 74.2897
R7555 a_n2318_13878.n30 a_n2318_13878.n118 70.6783
R7556 a_n2318_13878.n29 a_n2318_13878.n117 70.6783
R7557 a_n2318_13878.n28 a_n2318_13878.n71 70.6783
R7558 a_n2318_13878.n27 a_n2318_13878.n70 70.6783
R7559 a_n2318_13878.n27 a_n2318_13878.n69 70.6783
R7560 a_n2318_13878.n119 a_n2318_13878.n30 70.6782
R7561 a_n2318_13878.n114 a_n2318_13878.n113 48.2005
R7562 a_n2318_13878.n64 a_n2318_13878.t16 533.335
R7563 a_n2318_13878.n100 a_n2318_13878.n99 48.2005
R7564 a_n2318_13878.n58 a_n2318_13878.t54 533.335
R7565 a_n2318_13878.n82 a_n2318_13878.n81 48.2005
R7566 a_n2318_13878.t18 a_n2318_13878.n44 533.335
R7567 a_n2318_13878.n77 a_n2318_13878.n76 48.2005
R7568 a_n2318_13878.t55 a_n2318_13878.n37 533.335
R7569 a_n2318_13878.n95 a_n2318_13878.n85 48.2005
R7570 a_n2318_13878.t74 a_n2318_13878.n52 533.335
R7571 a_n2318_13878.n93 a_n2318_13878.n86 48.2005
R7572 a_n2318_13878.t81 a_n2318_13878.n50 533.335
R7573 a_n2318_13878.n91 a_n2318_13878.n87 48.2005
R7574 a_n2318_13878.t68 a_n2318_13878.n48 533.335
R7575 a_n2318_13878.n89 a_n2318_13878.n88 48.2005
R7576 a_n2318_13878.t64 a_n2318_13878.n46 533.335
R7577 a_n2318_13878.n60 a_n2318_13878.n65 16.6962
R7578 a_n2318_13878.n112 a_n2318_13878.n63 27.6507
R7579 a_n2318_13878.n54 a_n2318_13878.n67 16.6962
R7580 a_n2318_13878.n98 a_n2318_13878.n57 27.6507
R7581 a_n2318_13878.n80 a_n2318_13878.n40 16.6962
R7582 a_n2318_13878.n83 a_n2318_13878.n43 27.6507
R7583 a_n2318_13878.n75 a_n2318_13878.n33 16.6962
R7584 a_n2318_13878.n78 a_n2318_13878.n36 27.6507
R7585 a_n2318_13878.n61 a_n2318_13878.n65 41.7634
R7586 a_n2318_13878.n55 a_n2318_13878.n67 41.7634
R7587 a_n2318_13878.n80 a_n2318_13878.n41 41.7634
R7588 a_n2318_13878.n75 a_n2318_13878.n34 41.7634
R7589 a_n2318_13878.n25 a_n2318_13878.n24 31.238
R7590 a_n2318_13878.n96 a_n2318_13878.n51 35.3134
R7591 a_n2318_13878.n94 a_n2318_13878.n49 35.3134
R7592 a_n2318_13878.n92 a_n2318_13878.n47 35.3134
R7593 a_n2318_13878.n90 a_n2318_13878.n45 35.3134
R7594 a_n2318_13878.n1 a_n2318_13878.n26 23.891
R7595 a_n2318_13878.n32 a_n2318_13878.n14 12.705
R7596 a_n2318_13878.n5 a_n2318_13878.n97 12.5005
R7597 a_n2318_13878.n61 a_n2318_13878.n114 5.97853
R7598 a_n2318_13878.n62 a_n2318_13878.n66 41.7634
R7599 a_n2318_13878.n55 a_n2318_13878.n100 5.97853
R7600 a_n2318_13878.n56 a_n2318_13878.n68 41.7634
R7601 a_n2318_13878.n81 a_n2318_13878.n41 5.97853
R7602 a_n2318_13878.n72 a_n2318_13878.n42 41.7634
R7603 a_n2318_13878.n76 a_n2318_13878.n34 5.97853
R7604 a_n2318_13878.n73 a_n2318_13878.n35 41.7634
R7605 a_n2318_13878.n116 a_n2318_13878.n3 11.1956
R7606 a_n2318_13878.n115 a_n2318_13878.n60 27.6507
R7607 a_n2318_13878.n101 a_n2318_13878.n54 27.6507
R7608 a_n2318_13878.n40 a_n2318_13878.n79 27.6507
R7609 a_n2318_13878.n33 a_n2318_13878.n74 27.6507
R7610 a_n2318_13878.n84 a_n2318_13878.n28 9.85898
R7611 a_n2318_13878.n16 a_n2318_13878.n14 8.73345
R7612 a_n2318_13878.n97 a_n2318_13878.n8 8.73345
R7613 a_n2318_13878.n84 a_n2318_13878.n17 7.36035
R7614 a_n2318_13878.n29 a_n2318_13878.n116 6.01559
R7615 a_n2318_13878.n97 a_n2318_13878.n84 5.3452
R7616 a_n2318_13878.n39 a_n2318_13878.n20 4.01186
R7617 a_n2318_13878.n1 a_n2318_13878.n7 3.76565
R7618 a_n2318_13878.n118 a_n2318_13878.t33 3.61217
R7619 a_n2318_13878.n118 a_n2318_13878.t25 3.61217
R7620 a_n2318_13878.n117 a_n2318_13878.t23 3.61217
R7621 a_n2318_13878.n117 a_n2318_13878.t27 3.61217
R7622 a_n2318_13878.n71 a_n2318_13878.t13 3.61217
R7623 a_n2318_13878.n71 a_n2318_13878.t35 3.61217
R7624 a_n2318_13878.n70 a_n2318_13878.t11 3.61217
R7625 a_n2318_13878.n70 a_n2318_13878.t7 3.61217
R7626 a_n2318_13878.n69 a_n2318_13878.t21 3.61217
R7627 a_n2318_13878.n69 a_n2318_13878.t31 3.61217
R7628 a_n2318_13878.t5 a_n2318_13878.n119 3.61217
R7629 a_n2318_13878.n119 a_n2318_13878.t15 3.61217
R7630 a_n2318_13878.n110 a_n2318_13878.t41 2.82907
R7631 a_n2318_13878.n110 a_n2318_13878.t48 2.82907
R7632 a_n2318_13878.n111 a_n2318_13878.t40 2.82907
R7633 a_n2318_13878.n111 a_n2318_13878.t49 2.82907
R7634 a_n2318_13878.n109 a_n2318_13878.t47 2.82907
R7635 a_n2318_13878.n109 a_n2318_13878.t1 2.82907
R7636 a_n2318_13878.n108 a_n2318_13878.t38 2.82907
R7637 a_n2318_13878.n108 a_n2318_13878.t45 2.82907
R7638 a_n2318_13878.n107 a_n2318_13878.t50 2.82907
R7639 a_n2318_13878.n107 a_n2318_13878.t43 2.82907
R7640 a_n2318_13878.n105 a_n2318_13878.t37 2.82907
R7641 a_n2318_13878.n105 a_n2318_13878.t2 2.82907
R7642 a_n2318_13878.n106 a_n2318_13878.t42 2.82907
R7643 a_n2318_13878.n106 a_n2318_13878.t46 2.82907
R7644 a_n2318_13878.n104 a_n2318_13878.t36 2.82907
R7645 a_n2318_13878.n104 a_n2318_13878.t39 2.82907
R7646 a_n2318_13878.n103 a_n2318_13878.t0 2.82907
R7647 a_n2318_13878.n103 a_n2318_13878.t51 2.82907
R7648 a_n2318_13878.n102 a_n2318_13878.t44 2.82907
R7649 a_n2318_13878.n102 a_n2318_13878.t3 2.82907
R7650 a_n2318_13878.n116 a_n2318_13878.n14 1.30542
R7651 a_n2318_13878.n30 a_n2318_13878.n29 1.07378
R7652 a_n2318_13878.n28 a_n2318_13878.n27 1.07378
R7653 a_n2318_13878.n26 a_n2318_13878.n25 1.07378
R7654 a_n2318_13878.n11 a_n2318_13878.n12 1.04595
R7655 a_n2318_13878.n2 a_n2318_13878.n1 0.966409
R7656 a_n2318_13878.n22 a_n2318_13878.n21 0.758076
R7657 a_n2318_13878.n21 a_n2318_13878.n20 0.758076
R7658 a_n2318_13878.n19 a_n2318_13878.n18 0.758076
R7659 a_n2318_13878.n18 a_n2318_13878.n17 0.758076
R7660 a_n2318_13878.n16 a_n2318_13878.n15 0.758076
R7661 a_n2318_13878.n13 a_n2318_13878.n12 0.758076
R7662 a_n2318_13878.n11 a_n2318_13878.n10 0.758076
R7663 a_n2318_13878.n9 a_n2318_13878.n8 0.758076
R7664 a_n2318_13878.n6 a_n2318_13878.n4 0.758076
R7665 a_n2318_13878.n6 a_n2318_13878.n5 0.758076
R7666 a_n2318_13878.n2 a_n2318_13878.n0 0.758076
R7667 a_n2318_13878.n24 a_n2318_13878.n23 0.716017
R7668 a_n2318_13878.n13 a_n2318_13878.n15 0.67853
R7669 a_n2318_13878.n9 a_n2318_13878.n10 0.67853
R7670 a_n2318_13878.n0 a_n2318_13878.n3 0.568682
R7671 a_n2318_13878.n4 a_n2318_13878.n7 0.568682
R7672 a_n2318_13878.n39 a_n2318_13878.n19 0.568682
R7673 a_n2318_13878.n32 a_n2318_13878.n22 0.568682
R7674 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R7675 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R7676 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R7677 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R7678 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R7679 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R7680 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R7681 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R7682 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R7683 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R7684 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R7685 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R7686 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R7687 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R7688 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R7689 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R7690 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R7691 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R7692 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R7693 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R7694 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R7695 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R7696 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R7697 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R7698 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R7699 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R7700 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R7701 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R7702 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R7703 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R7704 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R7705 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R7706 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R7707 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R7708 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R7709 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R7710 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R7711 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R7712 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R7713 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R7714 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R7715 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R7716 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R7717 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R7718 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R7719 outputibias.n27 outputibias.n1 289.615
R7720 outputibias.n58 outputibias.n32 289.615
R7721 outputibias.n90 outputibias.n64 289.615
R7722 outputibias.n122 outputibias.n96 289.615
R7723 outputibias.n28 outputibias.n27 185
R7724 outputibias.n26 outputibias.n25 185
R7725 outputibias.n5 outputibias.n4 185
R7726 outputibias.n20 outputibias.n19 185
R7727 outputibias.n18 outputibias.n17 185
R7728 outputibias.n9 outputibias.n8 185
R7729 outputibias.n12 outputibias.n11 185
R7730 outputibias.n59 outputibias.n58 185
R7731 outputibias.n57 outputibias.n56 185
R7732 outputibias.n36 outputibias.n35 185
R7733 outputibias.n51 outputibias.n50 185
R7734 outputibias.n49 outputibias.n48 185
R7735 outputibias.n40 outputibias.n39 185
R7736 outputibias.n43 outputibias.n42 185
R7737 outputibias.n91 outputibias.n90 185
R7738 outputibias.n89 outputibias.n88 185
R7739 outputibias.n68 outputibias.n67 185
R7740 outputibias.n83 outputibias.n82 185
R7741 outputibias.n81 outputibias.n80 185
R7742 outputibias.n72 outputibias.n71 185
R7743 outputibias.n75 outputibias.n74 185
R7744 outputibias.n123 outputibias.n122 185
R7745 outputibias.n121 outputibias.n120 185
R7746 outputibias.n100 outputibias.n99 185
R7747 outputibias.n115 outputibias.n114 185
R7748 outputibias.n113 outputibias.n112 185
R7749 outputibias.n104 outputibias.n103 185
R7750 outputibias.n107 outputibias.n106 185
R7751 outputibias.n0 outputibias.t8 178.945
R7752 outputibias.n133 outputibias.t9 177.018
R7753 outputibias.n132 outputibias.t11 177.018
R7754 outputibias.n0 outputibias.t10 177.018
R7755 outputibias.t7 outputibias.n10 147.661
R7756 outputibias.t5 outputibias.n41 147.661
R7757 outputibias.t3 outputibias.n73 147.661
R7758 outputibias.t1 outputibias.n105 147.661
R7759 outputibias.n128 outputibias.t6 132.363
R7760 outputibias.n128 outputibias.t4 130.436
R7761 outputibias.n129 outputibias.t2 130.436
R7762 outputibias.n130 outputibias.t0 130.436
R7763 outputibias.n27 outputibias.n26 104.615
R7764 outputibias.n26 outputibias.n4 104.615
R7765 outputibias.n19 outputibias.n4 104.615
R7766 outputibias.n19 outputibias.n18 104.615
R7767 outputibias.n18 outputibias.n8 104.615
R7768 outputibias.n11 outputibias.n8 104.615
R7769 outputibias.n58 outputibias.n57 104.615
R7770 outputibias.n57 outputibias.n35 104.615
R7771 outputibias.n50 outputibias.n35 104.615
R7772 outputibias.n50 outputibias.n49 104.615
R7773 outputibias.n49 outputibias.n39 104.615
R7774 outputibias.n42 outputibias.n39 104.615
R7775 outputibias.n90 outputibias.n89 104.615
R7776 outputibias.n89 outputibias.n67 104.615
R7777 outputibias.n82 outputibias.n67 104.615
R7778 outputibias.n82 outputibias.n81 104.615
R7779 outputibias.n81 outputibias.n71 104.615
R7780 outputibias.n74 outputibias.n71 104.615
R7781 outputibias.n122 outputibias.n121 104.615
R7782 outputibias.n121 outputibias.n99 104.615
R7783 outputibias.n114 outputibias.n99 104.615
R7784 outputibias.n114 outputibias.n113 104.615
R7785 outputibias.n113 outputibias.n103 104.615
R7786 outputibias.n106 outputibias.n103 104.615
R7787 outputibias.n63 outputibias.n31 95.6354
R7788 outputibias.n63 outputibias.n62 94.6732
R7789 outputibias.n95 outputibias.n94 94.6732
R7790 outputibias.n127 outputibias.n126 94.6732
R7791 outputibias.n11 outputibias.t7 52.3082
R7792 outputibias.n42 outputibias.t5 52.3082
R7793 outputibias.n74 outputibias.t3 52.3082
R7794 outputibias.n106 outputibias.t1 52.3082
R7795 outputibias.n12 outputibias.n10 15.6674
R7796 outputibias.n43 outputibias.n41 15.6674
R7797 outputibias.n75 outputibias.n73 15.6674
R7798 outputibias.n107 outputibias.n105 15.6674
R7799 outputibias.n13 outputibias.n9 12.8005
R7800 outputibias.n44 outputibias.n40 12.8005
R7801 outputibias.n76 outputibias.n72 12.8005
R7802 outputibias.n108 outputibias.n104 12.8005
R7803 outputibias.n17 outputibias.n16 12.0247
R7804 outputibias.n48 outputibias.n47 12.0247
R7805 outputibias.n80 outputibias.n79 12.0247
R7806 outputibias.n112 outputibias.n111 12.0247
R7807 outputibias.n20 outputibias.n7 11.249
R7808 outputibias.n51 outputibias.n38 11.249
R7809 outputibias.n83 outputibias.n70 11.249
R7810 outputibias.n115 outputibias.n102 11.249
R7811 outputibias.n21 outputibias.n5 10.4732
R7812 outputibias.n52 outputibias.n36 10.4732
R7813 outputibias.n84 outputibias.n68 10.4732
R7814 outputibias.n116 outputibias.n100 10.4732
R7815 outputibias.n25 outputibias.n24 9.69747
R7816 outputibias.n56 outputibias.n55 9.69747
R7817 outputibias.n88 outputibias.n87 9.69747
R7818 outputibias.n120 outputibias.n119 9.69747
R7819 outputibias.n31 outputibias.n30 9.45567
R7820 outputibias.n62 outputibias.n61 9.45567
R7821 outputibias.n94 outputibias.n93 9.45567
R7822 outputibias.n126 outputibias.n125 9.45567
R7823 outputibias.n30 outputibias.n29 9.3005
R7824 outputibias.n3 outputibias.n2 9.3005
R7825 outputibias.n24 outputibias.n23 9.3005
R7826 outputibias.n22 outputibias.n21 9.3005
R7827 outputibias.n7 outputibias.n6 9.3005
R7828 outputibias.n16 outputibias.n15 9.3005
R7829 outputibias.n14 outputibias.n13 9.3005
R7830 outputibias.n61 outputibias.n60 9.3005
R7831 outputibias.n34 outputibias.n33 9.3005
R7832 outputibias.n55 outputibias.n54 9.3005
R7833 outputibias.n53 outputibias.n52 9.3005
R7834 outputibias.n38 outputibias.n37 9.3005
R7835 outputibias.n47 outputibias.n46 9.3005
R7836 outputibias.n45 outputibias.n44 9.3005
R7837 outputibias.n93 outputibias.n92 9.3005
R7838 outputibias.n66 outputibias.n65 9.3005
R7839 outputibias.n87 outputibias.n86 9.3005
R7840 outputibias.n85 outputibias.n84 9.3005
R7841 outputibias.n70 outputibias.n69 9.3005
R7842 outputibias.n79 outputibias.n78 9.3005
R7843 outputibias.n77 outputibias.n76 9.3005
R7844 outputibias.n125 outputibias.n124 9.3005
R7845 outputibias.n98 outputibias.n97 9.3005
R7846 outputibias.n119 outputibias.n118 9.3005
R7847 outputibias.n117 outputibias.n116 9.3005
R7848 outputibias.n102 outputibias.n101 9.3005
R7849 outputibias.n111 outputibias.n110 9.3005
R7850 outputibias.n109 outputibias.n108 9.3005
R7851 outputibias.n28 outputibias.n3 8.92171
R7852 outputibias.n59 outputibias.n34 8.92171
R7853 outputibias.n91 outputibias.n66 8.92171
R7854 outputibias.n123 outputibias.n98 8.92171
R7855 outputibias.n29 outputibias.n1 8.14595
R7856 outputibias.n60 outputibias.n32 8.14595
R7857 outputibias.n92 outputibias.n64 8.14595
R7858 outputibias.n124 outputibias.n96 8.14595
R7859 outputibias.n31 outputibias.n1 5.81868
R7860 outputibias.n62 outputibias.n32 5.81868
R7861 outputibias.n94 outputibias.n64 5.81868
R7862 outputibias.n126 outputibias.n96 5.81868
R7863 outputibias.n131 outputibias.n130 5.20947
R7864 outputibias.n29 outputibias.n28 5.04292
R7865 outputibias.n60 outputibias.n59 5.04292
R7866 outputibias.n92 outputibias.n91 5.04292
R7867 outputibias.n124 outputibias.n123 5.04292
R7868 outputibias.n131 outputibias.n127 4.42209
R7869 outputibias.n14 outputibias.n10 4.38594
R7870 outputibias.n45 outputibias.n41 4.38594
R7871 outputibias.n77 outputibias.n73 4.38594
R7872 outputibias.n109 outputibias.n105 4.38594
R7873 outputibias.n132 outputibias.n131 4.28454
R7874 outputibias.n25 outputibias.n3 4.26717
R7875 outputibias.n56 outputibias.n34 4.26717
R7876 outputibias.n88 outputibias.n66 4.26717
R7877 outputibias.n120 outputibias.n98 4.26717
R7878 outputibias.n24 outputibias.n5 3.49141
R7879 outputibias.n55 outputibias.n36 3.49141
R7880 outputibias.n87 outputibias.n68 3.49141
R7881 outputibias.n119 outputibias.n100 3.49141
R7882 outputibias.n21 outputibias.n20 2.71565
R7883 outputibias.n52 outputibias.n51 2.71565
R7884 outputibias.n84 outputibias.n83 2.71565
R7885 outputibias.n116 outputibias.n115 2.71565
R7886 outputibias.n17 outputibias.n7 1.93989
R7887 outputibias.n48 outputibias.n38 1.93989
R7888 outputibias.n80 outputibias.n70 1.93989
R7889 outputibias.n112 outputibias.n102 1.93989
R7890 outputibias.n130 outputibias.n129 1.9266
R7891 outputibias.n129 outputibias.n128 1.9266
R7892 outputibias.n133 outputibias.n132 1.92658
R7893 outputibias.n134 outputibias.n133 1.29913
R7894 outputibias.n16 outputibias.n9 1.16414
R7895 outputibias.n47 outputibias.n40 1.16414
R7896 outputibias.n79 outputibias.n72 1.16414
R7897 outputibias.n111 outputibias.n104 1.16414
R7898 outputibias.n127 outputibias.n95 0.962709
R7899 outputibias.n95 outputibias.n63 0.962709
R7900 outputibias.n13 outputibias.n12 0.388379
R7901 outputibias.n44 outputibias.n43 0.388379
R7902 outputibias.n76 outputibias.n75 0.388379
R7903 outputibias.n108 outputibias.n107 0.388379
R7904 outputibias.n134 outputibias.n0 0.337251
R7905 outputibias outputibias.n134 0.302375
R7906 outputibias.n30 outputibias.n2 0.155672
R7907 outputibias.n23 outputibias.n2 0.155672
R7908 outputibias.n23 outputibias.n22 0.155672
R7909 outputibias.n22 outputibias.n6 0.155672
R7910 outputibias.n15 outputibias.n6 0.155672
R7911 outputibias.n15 outputibias.n14 0.155672
R7912 outputibias.n61 outputibias.n33 0.155672
R7913 outputibias.n54 outputibias.n33 0.155672
R7914 outputibias.n54 outputibias.n53 0.155672
R7915 outputibias.n53 outputibias.n37 0.155672
R7916 outputibias.n46 outputibias.n37 0.155672
R7917 outputibias.n46 outputibias.n45 0.155672
R7918 outputibias.n93 outputibias.n65 0.155672
R7919 outputibias.n86 outputibias.n65 0.155672
R7920 outputibias.n86 outputibias.n85 0.155672
R7921 outputibias.n85 outputibias.n69 0.155672
R7922 outputibias.n78 outputibias.n69 0.155672
R7923 outputibias.n78 outputibias.n77 0.155672
R7924 outputibias.n125 outputibias.n97 0.155672
R7925 outputibias.n118 outputibias.n97 0.155672
R7926 outputibias.n118 outputibias.n117 0.155672
R7927 outputibias.n117 outputibias.n101 0.155672
R7928 outputibias.n110 outputibias.n101 0.155672
R7929 outputibias.n110 outputibias.n109 0.155672
R7930 gnd.n6940 gnd.n546 965.481
R7931 gnd.n3793 gnd.n3792 939.716
R7932 gnd.n3700 gnd.n2319 766.379
R7933 gnd.n3703 gnd.n3702 766.379
R7934 gnd.n2942 gnd.n2845 766.379
R7935 gnd.n2938 gnd.n2843 766.379
R7936 gnd.n3791 gnd.n2341 756.769
R7937 gnd.n3694 gnd.n3693 756.769
R7938 gnd.n3035 gnd.n2752 756.769
R7939 gnd.n3033 gnd.n2755 756.769
R7940 gnd.n6518 gnd.n798 756.769
R7941 gnd.n6939 gnd.n547 756.769
R7942 gnd.n7151 gnd.n7150 756.769
R7943 gnd.n6341 gnd.n963 756.769
R7944 gnd.n7446 gnd.n129 751.963
R7945 gnd.n7604 gnd.n7603 751.963
R7946 gnd.n1337 gnd.n1284 751.963
R7947 gnd.n6015 gnd.n1339 751.963
R7948 gnd.n6260 gnd.n1113 751.963
R7949 gnd.n5356 gnd.n1111 751.963
R7950 gnd.n3860 gnd.n3795 751.963
R7951 gnd.n4180 gnd.n2318 751.963
R7952 gnd.n7601 gnd.n131 732.745
R7953 gnd.n199 gnd.n127 732.745
R7954 gnd.n6018 gnd.n6017 732.745
R7955 gnd.n6090 gnd.n1288 732.745
R7956 gnd.n6262 gnd.n1108 732.745
R7957 gnd.n2103 gnd.n1110 732.745
R7958 gnd.n4099 gnd.n3794 732.745
R7959 gnd.n4178 gnd.n3958 732.745
R7960 gnd.n5402 gnd.n1118 711.122
R7961 gnd.n6102 gnd.n1244 711.122
R7962 gnd.n5406 gnd.n1953 711.122
R7963 gnd.n5820 gnd.n1247 711.122
R7964 gnd.n6514 gnd.n798 585
R7965 gnd.n798 gnd.n797 585
R7966 gnd.n6513 gnd.n6512 585
R7967 gnd.n6512 gnd.n6511 585
R7968 gnd.n801 gnd.n800 585
R7969 gnd.n6510 gnd.n801 585
R7970 gnd.n6508 gnd.n6507 585
R7971 gnd.n6509 gnd.n6508 585
R7972 gnd.n6506 gnd.n803 585
R7973 gnd.n803 gnd.n802 585
R7974 gnd.n6505 gnd.n6504 585
R7975 gnd.n6504 gnd.n6503 585
R7976 gnd.n809 gnd.n808 585
R7977 gnd.n6502 gnd.n809 585
R7978 gnd.n6500 gnd.n6499 585
R7979 gnd.n6501 gnd.n6500 585
R7980 gnd.n6498 gnd.n811 585
R7981 gnd.n811 gnd.n810 585
R7982 gnd.n6497 gnd.n6496 585
R7983 gnd.n6496 gnd.n6495 585
R7984 gnd.n817 gnd.n816 585
R7985 gnd.n6494 gnd.n817 585
R7986 gnd.n6492 gnd.n6491 585
R7987 gnd.n6493 gnd.n6492 585
R7988 gnd.n6490 gnd.n819 585
R7989 gnd.n819 gnd.n818 585
R7990 gnd.n6489 gnd.n6488 585
R7991 gnd.n6488 gnd.n6487 585
R7992 gnd.n825 gnd.n824 585
R7993 gnd.n6486 gnd.n825 585
R7994 gnd.n6484 gnd.n6483 585
R7995 gnd.n6485 gnd.n6484 585
R7996 gnd.n6482 gnd.n827 585
R7997 gnd.n827 gnd.n826 585
R7998 gnd.n6481 gnd.n6480 585
R7999 gnd.n6480 gnd.n6479 585
R8000 gnd.n833 gnd.n832 585
R8001 gnd.n6478 gnd.n833 585
R8002 gnd.n6476 gnd.n6475 585
R8003 gnd.n6477 gnd.n6476 585
R8004 gnd.n6474 gnd.n835 585
R8005 gnd.n835 gnd.n834 585
R8006 gnd.n6473 gnd.n6472 585
R8007 gnd.n6472 gnd.n6471 585
R8008 gnd.n841 gnd.n840 585
R8009 gnd.n6470 gnd.n841 585
R8010 gnd.n6468 gnd.n6467 585
R8011 gnd.n6469 gnd.n6468 585
R8012 gnd.n6466 gnd.n843 585
R8013 gnd.n843 gnd.n842 585
R8014 gnd.n6465 gnd.n6464 585
R8015 gnd.n6464 gnd.n6463 585
R8016 gnd.n849 gnd.n848 585
R8017 gnd.n6462 gnd.n849 585
R8018 gnd.n6460 gnd.n6459 585
R8019 gnd.n6461 gnd.n6460 585
R8020 gnd.n6458 gnd.n851 585
R8021 gnd.n851 gnd.n850 585
R8022 gnd.n6457 gnd.n6456 585
R8023 gnd.n6456 gnd.n6455 585
R8024 gnd.n857 gnd.n856 585
R8025 gnd.n6454 gnd.n857 585
R8026 gnd.n6452 gnd.n6451 585
R8027 gnd.n6453 gnd.n6452 585
R8028 gnd.n6450 gnd.n859 585
R8029 gnd.n859 gnd.n858 585
R8030 gnd.n6449 gnd.n6448 585
R8031 gnd.n6448 gnd.n6447 585
R8032 gnd.n865 gnd.n864 585
R8033 gnd.n6446 gnd.n865 585
R8034 gnd.n6444 gnd.n6443 585
R8035 gnd.n6445 gnd.n6444 585
R8036 gnd.n6442 gnd.n867 585
R8037 gnd.n867 gnd.n866 585
R8038 gnd.n6441 gnd.n6440 585
R8039 gnd.n6440 gnd.n6439 585
R8040 gnd.n873 gnd.n872 585
R8041 gnd.n6438 gnd.n873 585
R8042 gnd.n6436 gnd.n6435 585
R8043 gnd.n6437 gnd.n6436 585
R8044 gnd.n6434 gnd.n875 585
R8045 gnd.n875 gnd.n874 585
R8046 gnd.n6433 gnd.n6432 585
R8047 gnd.n6432 gnd.n6431 585
R8048 gnd.n881 gnd.n880 585
R8049 gnd.n6430 gnd.n881 585
R8050 gnd.n6428 gnd.n6427 585
R8051 gnd.n6429 gnd.n6428 585
R8052 gnd.n6426 gnd.n883 585
R8053 gnd.n883 gnd.n882 585
R8054 gnd.n6425 gnd.n6424 585
R8055 gnd.n6424 gnd.n6423 585
R8056 gnd.n889 gnd.n888 585
R8057 gnd.n6422 gnd.n889 585
R8058 gnd.n6420 gnd.n6419 585
R8059 gnd.n6421 gnd.n6420 585
R8060 gnd.n6418 gnd.n891 585
R8061 gnd.n891 gnd.n890 585
R8062 gnd.n6417 gnd.n6416 585
R8063 gnd.n6416 gnd.n6415 585
R8064 gnd.n897 gnd.n896 585
R8065 gnd.n6414 gnd.n897 585
R8066 gnd.n6412 gnd.n6411 585
R8067 gnd.n6413 gnd.n6412 585
R8068 gnd.n6410 gnd.n899 585
R8069 gnd.n899 gnd.n898 585
R8070 gnd.n6409 gnd.n6408 585
R8071 gnd.n6408 gnd.n6407 585
R8072 gnd.n905 gnd.n904 585
R8073 gnd.n6406 gnd.n905 585
R8074 gnd.n6404 gnd.n6403 585
R8075 gnd.n6405 gnd.n6404 585
R8076 gnd.n6402 gnd.n907 585
R8077 gnd.n907 gnd.n906 585
R8078 gnd.n6401 gnd.n6400 585
R8079 gnd.n6400 gnd.n6399 585
R8080 gnd.n913 gnd.n912 585
R8081 gnd.n6398 gnd.n913 585
R8082 gnd.n6396 gnd.n6395 585
R8083 gnd.n6397 gnd.n6396 585
R8084 gnd.n6394 gnd.n915 585
R8085 gnd.n915 gnd.n914 585
R8086 gnd.n6393 gnd.n6392 585
R8087 gnd.n6392 gnd.n6391 585
R8088 gnd.n921 gnd.n920 585
R8089 gnd.n6390 gnd.n921 585
R8090 gnd.n6388 gnd.n6387 585
R8091 gnd.n6389 gnd.n6388 585
R8092 gnd.n6386 gnd.n923 585
R8093 gnd.n923 gnd.n922 585
R8094 gnd.n6385 gnd.n6384 585
R8095 gnd.n6384 gnd.n6383 585
R8096 gnd.n929 gnd.n928 585
R8097 gnd.n6382 gnd.n929 585
R8098 gnd.n6380 gnd.n6379 585
R8099 gnd.n6381 gnd.n6380 585
R8100 gnd.n6378 gnd.n931 585
R8101 gnd.n931 gnd.n930 585
R8102 gnd.n6377 gnd.n6376 585
R8103 gnd.n6376 gnd.n6375 585
R8104 gnd.n937 gnd.n936 585
R8105 gnd.n6374 gnd.n937 585
R8106 gnd.n6372 gnd.n6371 585
R8107 gnd.n6373 gnd.n6372 585
R8108 gnd.n6370 gnd.n939 585
R8109 gnd.n939 gnd.n938 585
R8110 gnd.n6369 gnd.n6368 585
R8111 gnd.n6368 gnd.n6367 585
R8112 gnd.n945 gnd.n944 585
R8113 gnd.n6366 gnd.n945 585
R8114 gnd.n6364 gnd.n6363 585
R8115 gnd.n6365 gnd.n6364 585
R8116 gnd.n6362 gnd.n947 585
R8117 gnd.n947 gnd.n946 585
R8118 gnd.n6361 gnd.n6360 585
R8119 gnd.n6360 gnd.n6359 585
R8120 gnd.n953 gnd.n952 585
R8121 gnd.n6358 gnd.n953 585
R8122 gnd.n6356 gnd.n6355 585
R8123 gnd.n6357 gnd.n6356 585
R8124 gnd.n6354 gnd.n955 585
R8125 gnd.n955 gnd.n954 585
R8126 gnd.n6353 gnd.n6352 585
R8127 gnd.n6352 gnd.n6351 585
R8128 gnd.n961 gnd.n960 585
R8129 gnd.n6350 gnd.n961 585
R8130 gnd.n6348 gnd.n6347 585
R8131 gnd.n6349 gnd.n6348 585
R8132 gnd.n6518 gnd.n6517 585
R8133 gnd.n6519 gnd.n6518 585
R8134 gnd.n796 gnd.n795 585
R8135 gnd.n6520 gnd.n796 585
R8136 gnd.n6523 gnd.n6522 585
R8137 gnd.n6522 gnd.n6521 585
R8138 gnd.n793 gnd.n792 585
R8139 gnd.n792 gnd.n791 585
R8140 gnd.n6528 gnd.n6527 585
R8141 gnd.n6529 gnd.n6528 585
R8142 gnd.n790 gnd.n789 585
R8143 gnd.n6530 gnd.n790 585
R8144 gnd.n6533 gnd.n6532 585
R8145 gnd.n6532 gnd.n6531 585
R8146 gnd.n787 gnd.n786 585
R8147 gnd.n786 gnd.n785 585
R8148 gnd.n6538 gnd.n6537 585
R8149 gnd.n6539 gnd.n6538 585
R8150 gnd.n784 gnd.n783 585
R8151 gnd.n6540 gnd.n784 585
R8152 gnd.n6543 gnd.n6542 585
R8153 gnd.n6542 gnd.n6541 585
R8154 gnd.n781 gnd.n780 585
R8155 gnd.n780 gnd.n779 585
R8156 gnd.n6548 gnd.n6547 585
R8157 gnd.n6549 gnd.n6548 585
R8158 gnd.n778 gnd.n777 585
R8159 gnd.n6550 gnd.n778 585
R8160 gnd.n6553 gnd.n6552 585
R8161 gnd.n6552 gnd.n6551 585
R8162 gnd.n775 gnd.n774 585
R8163 gnd.n774 gnd.n773 585
R8164 gnd.n6558 gnd.n6557 585
R8165 gnd.n6559 gnd.n6558 585
R8166 gnd.n772 gnd.n771 585
R8167 gnd.n6560 gnd.n772 585
R8168 gnd.n6563 gnd.n6562 585
R8169 gnd.n6562 gnd.n6561 585
R8170 gnd.n769 gnd.n768 585
R8171 gnd.n768 gnd.n767 585
R8172 gnd.n6568 gnd.n6567 585
R8173 gnd.n6569 gnd.n6568 585
R8174 gnd.n766 gnd.n765 585
R8175 gnd.n6570 gnd.n766 585
R8176 gnd.n6573 gnd.n6572 585
R8177 gnd.n6572 gnd.n6571 585
R8178 gnd.n763 gnd.n762 585
R8179 gnd.n762 gnd.n761 585
R8180 gnd.n6578 gnd.n6577 585
R8181 gnd.n6579 gnd.n6578 585
R8182 gnd.n760 gnd.n759 585
R8183 gnd.n6580 gnd.n760 585
R8184 gnd.n6583 gnd.n6582 585
R8185 gnd.n6582 gnd.n6581 585
R8186 gnd.n757 gnd.n756 585
R8187 gnd.n756 gnd.n755 585
R8188 gnd.n6588 gnd.n6587 585
R8189 gnd.n6589 gnd.n6588 585
R8190 gnd.n754 gnd.n753 585
R8191 gnd.n6590 gnd.n754 585
R8192 gnd.n6593 gnd.n6592 585
R8193 gnd.n6592 gnd.n6591 585
R8194 gnd.n751 gnd.n750 585
R8195 gnd.n750 gnd.n749 585
R8196 gnd.n6598 gnd.n6597 585
R8197 gnd.n6599 gnd.n6598 585
R8198 gnd.n748 gnd.n747 585
R8199 gnd.n6600 gnd.n748 585
R8200 gnd.n6603 gnd.n6602 585
R8201 gnd.n6602 gnd.n6601 585
R8202 gnd.n745 gnd.n744 585
R8203 gnd.n744 gnd.n743 585
R8204 gnd.n6608 gnd.n6607 585
R8205 gnd.n6609 gnd.n6608 585
R8206 gnd.n742 gnd.n741 585
R8207 gnd.n6610 gnd.n742 585
R8208 gnd.n6613 gnd.n6612 585
R8209 gnd.n6612 gnd.n6611 585
R8210 gnd.n739 gnd.n738 585
R8211 gnd.n738 gnd.n737 585
R8212 gnd.n6618 gnd.n6617 585
R8213 gnd.n6619 gnd.n6618 585
R8214 gnd.n736 gnd.n735 585
R8215 gnd.n6620 gnd.n736 585
R8216 gnd.n6623 gnd.n6622 585
R8217 gnd.n6622 gnd.n6621 585
R8218 gnd.n733 gnd.n732 585
R8219 gnd.n732 gnd.n731 585
R8220 gnd.n6628 gnd.n6627 585
R8221 gnd.n6629 gnd.n6628 585
R8222 gnd.n730 gnd.n729 585
R8223 gnd.n6630 gnd.n730 585
R8224 gnd.n6633 gnd.n6632 585
R8225 gnd.n6632 gnd.n6631 585
R8226 gnd.n727 gnd.n726 585
R8227 gnd.n726 gnd.n725 585
R8228 gnd.n6638 gnd.n6637 585
R8229 gnd.n6639 gnd.n6638 585
R8230 gnd.n724 gnd.n723 585
R8231 gnd.n6640 gnd.n724 585
R8232 gnd.n6643 gnd.n6642 585
R8233 gnd.n6642 gnd.n6641 585
R8234 gnd.n721 gnd.n720 585
R8235 gnd.n720 gnd.n719 585
R8236 gnd.n6648 gnd.n6647 585
R8237 gnd.n6649 gnd.n6648 585
R8238 gnd.n718 gnd.n717 585
R8239 gnd.n6650 gnd.n718 585
R8240 gnd.n6653 gnd.n6652 585
R8241 gnd.n6652 gnd.n6651 585
R8242 gnd.n715 gnd.n714 585
R8243 gnd.n714 gnd.n713 585
R8244 gnd.n6658 gnd.n6657 585
R8245 gnd.n6659 gnd.n6658 585
R8246 gnd.n712 gnd.n711 585
R8247 gnd.n6660 gnd.n712 585
R8248 gnd.n6663 gnd.n6662 585
R8249 gnd.n6662 gnd.n6661 585
R8250 gnd.n709 gnd.n708 585
R8251 gnd.n708 gnd.n707 585
R8252 gnd.n6668 gnd.n6667 585
R8253 gnd.n6669 gnd.n6668 585
R8254 gnd.n706 gnd.n705 585
R8255 gnd.n6670 gnd.n706 585
R8256 gnd.n6673 gnd.n6672 585
R8257 gnd.n6672 gnd.n6671 585
R8258 gnd.n703 gnd.n702 585
R8259 gnd.n702 gnd.n701 585
R8260 gnd.n6678 gnd.n6677 585
R8261 gnd.n6679 gnd.n6678 585
R8262 gnd.n700 gnd.n699 585
R8263 gnd.n6680 gnd.n700 585
R8264 gnd.n6683 gnd.n6682 585
R8265 gnd.n6682 gnd.n6681 585
R8266 gnd.n697 gnd.n696 585
R8267 gnd.n696 gnd.n695 585
R8268 gnd.n6688 gnd.n6687 585
R8269 gnd.n6689 gnd.n6688 585
R8270 gnd.n694 gnd.n693 585
R8271 gnd.n6690 gnd.n694 585
R8272 gnd.n6693 gnd.n6692 585
R8273 gnd.n6692 gnd.n6691 585
R8274 gnd.n691 gnd.n690 585
R8275 gnd.n690 gnd.n689 585
R8276 gnd.n6698 gnd.n6697 585
R8277 gnd.n6699 gnd.n6698 585
R8278 gnd.n688 gnd.n687 585
R8279 gnd.n6700 gnd.n688 585
R8280 gnd.n6703 gnd.n6702 585
R8281 gnd.n6702 gnd.n6701 585
R8282 gnd.n685 gnd.n684 585
R8283 gnd.n684 gnd.n683 585
R8284 gnd.n6708 gnd.n6707 585
R8285 gnd.n6709 gnd.n6708 585
R8286 gnd.n682 gnd.n681 585
R8287 gnd.n6710 gnd.n682 585
R8288 gnd.n6713 gnd.n6712 585
R8289 gnd.n6712 gnd.n6711 585
R8290 gnd.n679 gnd.n678 585
R8291 gnd.n678 gnd.n677 585
R8292 gnd.n6718 gnd.n6717 585
R8293 gnd.n6719 gnd.n6718 585
R8294 gnd.n676 gnd.n675 585
R8295 gnd.n6720 gnd.n676 585
R8296 gnd.n6723 gnd.n6722 585
R8297 gnd.n6722 gnd.n6721 585
R8298 gnd.n673 gnd.n672 585
R8299 gnd.n672 gnd.n671 585
R8300 gnd.n6728 gnd.n6727 585
R8301 gnd.n6729 gnd.n6728 585
R8302 gnd.n670 gnd.n669 585
R8303 gnd.n6730 gnd.n670 585
R8304 gnd.n6733 gnd.n6732 585
R8305 gnd.n6732 gnd.n6731 585
R8306 gnd.n667 gnd.n666 585
R8307 gnd.n666 gnd.n665 585
R8308 gnd.n6738 gnd.n6737 585
R8309 gnd.n6739 gnd.n6738 585
R8310 gnd.n664 gnd.n663 585
R8311 gnd.n6740 gnd.n664 585
R8312 gnd.n6743 gnd.n6742 585
R8313 gnd.n6742 gnd.n6741 585
R8314 gnd.n661 gnd.n660 585
R8315 gnd.n660 gnd.n659 585
R8316 gnd.n6748 gnd.n6747 585
R8317 gnd.n6749 gnd.n6748 585
R8318 gnd.n658 gnd.n657 585
R8319 gnd.n6750 gnd.n658 585
R8320 gnd.n6753 gnd.n6752 585
R8321 gnd.n6752 gnd.n6751 585
R8322 gnd.n655 gnd.n654 585
R8323 gnd.n654 gnd.n653 585
R8324 gnd.n6758 gnd.n6757 585
R8325 gnd.n6759 gnd.n6758 585
R8326 gnd.n652 gnd.n651 585
R8327 gnd.n6760 gnd.n652 585
R8328 gnd.n6763 gnd.n6762 585
R8329 gnd.n6762 gnd.n6761 585
R8330 gnd.n649 gnd.n648 585
R8331 gnd.n648 gnd.n647 585
R8332 gnd.n6768 gnd.n6767 585
R8333 gnd.n6769 gnd.n6768 585
R8334 gnd.n646 gnd.n645 585
R8335 gnd.n6770 gnd.n646 585
R8336 gnd.n6773 gnd.n6772 585
R8337 gnd.n6772 gnd.n6771 585
R8338 gnd.n643 gnd.n642 585
R8339 gnd.n642 gnd.n641 585
R8340 gnd.n6778 gnd.n6777 585
R8341 gnd.n6779 gnd.n6778 585
R8342 gnd.n640 gnd.n639 585
R8343 gnd.n6780 gnd.n640 585
R8344 gnd.n6783 gnd.n6782 585
R8345 gnd.n6782 gnd.n6781 585
R8346 gnd.n637 gnd.n636 585
R8347 gnd.n636 gnd.n635 585
R8348 gnd.n6788 gnd.n6787 585
R8349 gnd.n6789 gnd.n6788 585
R8350 gnd.n634 gnd.n633 585
R8351 gnd.n6790 gnd.n634 585
R8352 gnd.n6793 gnd.n6792 585
R8353 gnd.n6792 gnd.n6791 585
R8354 gnd.n631 gnd.n630 585
R8355 gnd.n630 gnd.n629 585
R8356 gnd.n6798 gnd.n6797 585
R8357 gnd.n6799 gnd.n6798 585
R8358 gnd.n628 gnd.n627 585
R8359 gnd.n6800 gnd.n628 585
R8360 gnd.n6803 gnd.n6802 585
R8361 gnd.n6802 gnd.n6801 585
R8362 gnd.n625 gnd.n624 585
R8363 gnd.n624 gnd.n623 585
R8364 gnd.n6808 gnd.n6807 585
R8365 gnd.n6809 gnd.n6808 585
R8366 gnd.n622 gnd.n621 585
R8367 gnd.n6810 gnd.n622 585
R8368 gnd.n6813 gnd.n6812 585
R8369 gnd.n6812 gnd.n6811 585
R8370 gnd.n619 gnd.n618 585
R8371 gnd.n618 gnd.n617 585
R8372 gnd.n6818 gnd.n6817 585
R8373 gnd.n6819 gnd.n6818 585
R8374 gnd.n616 gnd.n615 585
R8375 gnd.n6820 gnd.n616 585
R8376 gnd.n6823 gnd.n6822 585
R8377 gnd.n6822 gnd.n6821 585
R8378 gnd.n613 gnd.n612 585
R8379 gnd.n612 gnd.n611 585
R8380 gnd.n6828 gnd.n6827 585
R8381 gnd.n6829 gnd.n6828 585
R8382 gnd.n610 gnd.n609 585
R8383 gnd.n6830 gnd.n610 585
R8384 gnd.n6833 gnd.n6832 585
R8385 gnd.n6832 gnd.n6831 585
R8386 gnd.n607 gnd.n606 585
R8387 gnd.n606 gnd.n605 585
R8388 gnd.n6838 gnd.n6837 585
R8389 gnd.n6839 gnd.n6838 585
R8390 gnd.n604 gnd.n603 585
R8391 gnd.n6840 gnd.n604 585
R8392 gnd.n6843 gnd.n6842 585
R8393 gnd.n6842 gnd.n6841 585
R8394 gnd.n601 gnd.n600 585
R8395 gnd.n600 gnd.n599 585
R8396 gnd.n6848 gnd.n6847 585
R8397 gnd.n6849 gnd.n6848 585
R8398 gnd.n598 gnd.n597 585
R8399 gnd.n6850 gnd.n598 585
R8400 gnd.n6853 gnd.n6852 585
R8401 gnd.n6852 gnd.n6851 585
R8402 gnd.n595 gnd.n594 585
R8403 gnd.n594 gnd.n593 585
R8404 gnd.n6858 gnd.n6857 585
R8405 gnd.n6859 gnd.n6858 585
R8406 gnd.n592 gnd.n591 585
R8407 gnd.n6860 gnd.n592 585
R8408 gnd.n6863 gnd.n6862 585
R8409 gnd.n6862 gnd.n6861 585
R8410 gnd.n589 gnd.n588 585
R8411 gnd.n588 gnd.n587 585
R8412 gnd.n6868 gnd.n6867 585
R8413 gnd.n6869 gnd.n6868 585
R8414 gnd.n586 gnd.n585 585
R8415 gnd.n6870 gnd.n586 585
R8416 gnd.n6873 gnd.n6872 585
R8417 gnd.n6872 gnd.n6871 585
R8418 gnd.n583 gnd.n582 585
R8419 gnd.n582 gnd.n581 585
R8420 gnd.n6878 gnd.n6877 585
R8421 gnd.n6879 gnd.n6878 585
R8422 gnd.n580 gnd.n579 585
R8423 gnd.n6880 gnd.n580 585
R8424 gnd.n6883 gnd.n6882 585
R8425 gnd.n6882 gnd.n6881 585
R8426 gnd.n577 gnd.n576 585
R8427 gnd.n576 gnd.n575 585
R8428 gnd.n6888 gnd.n6887 585
R8429 gnd.n6889 gnd.n6888 585
R8430 gnd.n574 gnd.n573 585
R8431 gnd.n6890 gnd.n574 585
R8432 gnd.n6893 gnd.n6892 585
R8433 gnd.n6892 gnd.n6891 585
R8434 gnd.n571 gnd.n570 585
R8435 gnd.n570 gnd.n569 585
R8436 gnd.n6898 gnd.n6897 585
R8437 gnd.n6899 gnd.n6898 585
R8438 gnd.n568 gnd.n567 585
R8439 gnd.n6900 gnd.n568 585
R8440 gnd.n6903 gnd.n6902 585
R8441 gnd.n6902 gnd.n6901 585
R8442 gnd.n565 gnd.n564 585
R8443 gnd.n564 gnd.n563 585
R8444 gnd.n6908 gnd.n6907 585
R8445 gnd.n6909 gnd.n6908 585
R8446 gnd.n562 gnd.n561 585
R8447 gnd.n6910 gnd.n562 585
R8448 gnd.n6913 gnd.n6912 585
R8449 gnd.n6912 gnd.n6911 585
R8450 gnd.n559 gnd.n558 585
R8451 gnd.n558 gnd.n557 585
R8452 gnd.n6918 gnd.n6917 585
R8453 gnd.n6919 gnd.n6918 585
R8454 gnd.n556 gnd.n555 585
R8455 gnd.n6920 gnd.n556 585
R8456 gnd.n6923 gnd.n6922 585
R8457 gnd.n6922 gnd.n6921 585
R8458 gnd.n553 gnd.n552 585
R8459 gnd.n552 gnd.n551 585
R8460 gnd.n6929 gnd.n6928 585
R8461 gnd.n6930 gnd.n6929 585
R8462 gnd.n550 gnd.n549 585
R8463 gnd.n6931 gnd.n550 585
R8464 gnd.n6934 gnd.n6933 585
R8465 gnd.n6933 gnd.n6932 585
R8466 gnd.n6935 gnd.n547 585
R8467 gnd.n547 gnd.n546 585
R8468 gnd.n422 gnd.n421 585
R8469 gnd.n7142 gnd.n421 585
R8470 gnd.n7145 gnd.n7144 585
R8471 gnd.n7144 gnd.n7143 585
R8472 gnd.n425 gnd.n424 585
R8473 gnd.n7141 gnd.n425 585
R8474 gnd.n7139 gnd.n7138 585
R8475 gnd.n7140 gnd.n7139 585
R8476 gnd.n428 gnd.n427 585
R8477 gnd.n427 gnd.n426 585
R8478 gnd.n7134 gnd.n7133 585
R8479 gnd.n7133 gnd.n7132 585
R8480 gnd.n431 gnd.n430 585
R8481 gnd.n7131 gnd.n431 585
R8482 gnd.n7129 gnd.n7128 585
R8483 gnd.n7130 gnd.n7129 585
R8484 gnd.n434 gnd.n433 585
R8485 gnd.n433 gnd.n432 585
R8486 gnd.n7124 gnd.n7123 585
R8487 gnd.n7123 gnd.n7122 585
R8488 gnd.n437 gnd.n436 585
R8489 gnd.n7121 gnd.n437 585
R8490 gnd.n7119 gnd.n7118 585
R8491 gnd.n7120 gnd.n7119 585
R8492 gnd.n440 gnd.n439 585
R8493 gnd.n439 gnd.n438 585
R8494 gnd.n7114 gnd.n7113 585
R8495 gnd.n7113 gnd.n7112 585
R8496 gnd.n443 gnd.n442 585
R8497 gnd.n7111 gnd.n443 585
R8498 gnd.n7109 gnd.n7108 585
R8499 gnd.n7110 gnd.n7109 585
R8500 gnd.n446 gnd.n445 585
R8501 gnd.n445 gnd.n444 585
R8502 gnd.n7104 gnd.n7103 585
R8503 gnd.n7103 gnd.n7102 585
R8504 gnd.n449 gnd.n448 585
R8505 gnd.n7101 gnd.n449 585
R8506 gnd.n7099 gnd.n7098 585
R8507 gnd.n7100 gnd.n7099 585
R8508 gnd.n452 gnd.n451 585
R8509 gnd.n451 gnd.n450 585
R8510 gnd.n7094 gnd.n7093 585
R8511 gnd.n7093 gnd.n7092 585
R8512 gnd.n455 gnd.n454 585
R8513 gnd.n7091 gnd.n455 585
R8514 gnd.n7089 gnd.n7088 585
R8515 gnd.n7090 gnd.n7089 585
R8516 gnd.n458 gnd.n457 585
R8517 gnd.n457 gnd.n456 585
R8518 gnd.n7084 gnd.n7083 585
R8519 gnd.n7083 gnd.n7082 585
R8520 gnd.n461 gnd.n460 585
R8521 gnd.n7081 gnd.n461 585
R8522 gnd.n7079 gnd.n7078 585
R8523 gnd.n7080 gnd.n7079 585
R8524 gnd.n464 gnd.n463 585
R8525 gnd.n463 gnd.n462 585
R8526 gnd.n7074 gnd.n7073 585
R8527 gnd.n7073 gnd.n7072 585
R8528 gnd.n467 gnd.n466 585
R8529 gnd.n7071 gnd.n467 585
R8530 gnd.n7069 gnd.n7068 585
R8531 gnd.n7070 gnd.n7069 585
R8532 gnd.n470 gnd.n469 585
R8533 gnd.n469 gnd.n468 585
R8534 gnd.n7064 gnd.n7063 585
R8535 gnd.n7063 gnd.n7062 585
R8536 gnd.n473 gnd.n472 585
R8537 gnd.n7061 gnd.n473 585
R8538 gnd.n7059 gnd.n7058 585
R8539 gnd.n7060 gnd.n7059 585
R8540 gnd.n476 gnd.n475 585
R8541 gnd.n475 gnd.n474 585
R8542 gnd.n7054 gnd.n7053 585
R8543 gnd.n7053 gnd.n7052 585
R8544 gnd.n479 gnd.n478 585
R8545 gnd.n7051 gnd.n479 585
R8546 gnd.n7049 gnd.n7048 585
R8547 gnd.n7050 gnd.n7049 585
R8548 gnd.n482 gnd.n481 585
R8549 gnd.n481 gnd.n480 585
R8550 gnd.n7044 gnd.n7043 585
R8551 gnd.n7043 gnd.n7042 585
R8552 gnd.n485 gnd.n484 585
R8553 gnd.n7041 gnd.n485 585
R8554 gnd.n7039 gnd.n7038 585
R8555 gnd.n7040 gnd.n7039 585
R8556 gnd.n488 gnd.n487 585
R8557 gnd.n487 gnd.n486 585
R8558 gnd.n7034 gnd.n7033 585
R8559 gnd.n7033 gnd.n7032 585
R8560 gnd.n491 gnd.n490 585
R8561 gnd.n7031 gnd.n491 585
R8562 gnd.n7029 gnd.n7028 585
R8563 gnd.n7030 gnd.n7029 585
R8564 gnd.n494 gnd.n493 585
R8565 gnd.n493 gnd.n492 585
R8566 gnd.n7024 gnd.n7023 585
R8567 gnd.n7023 gnd.n7022 585
R8568 gnd.n497 gnd.n496 585
R8569 gnd.n7021 gnd.n497 585
R8570 gnd.n7019 gnd.n7018 585
R8571 gnd.n7020 gnd.n7019 585
R8572 gnd.n500 gnd.n499 585
R8573 gnd.n499 gnd.n498 585
R8574 gnd.n7014 gnd.n7013 585
R8575 gnd.n7013 gnd.n7012 585
R8576 gnd.n503 gnd.n502 585
R8577 gnd.n7011 gnd.n503 585
R8578 gnd.n7009 gnd.n7008 585
R8579 gnd.n7010 gnd.n7009 585
R8580 gnd.n506 gnd.n505 585
R8581 gnd.n505 gnd.n504 585
R8582 gnd.n7004 gnd.n7003 585
R8583 gnd.n7003 gnd.n7002 585
R8584 gnd.n509 gnd.n508 585
R8585 gnd.n7001 gnd.n509 585
R8586 gnd.n6999 gnd.n6998 585
R8587 gnd.n7000 gnd.n6999 585
R8588 gnd.n512 gnd.n511 585
R8589 gnd.n511 gnd.n510 585
R8590 gnd.n6994 gnd.n6993 585
R8591 gnd.n6993 gnd.n6992 585
R8592 gnd.n515 gnd.n514 585
R8593 gnd.n6991 gnd.n515 585
R8594 gnd.n6989 gnd.n6988 585
R8595 gnd.n6990 gnd.n6989 585
R8596 gnd.n518 gnd.n517 585
R8597 gnd.n517 gnd.n516 585
R8598 gnd.n6984 gnd.n6983 585
R8599 gnd.n6983 gnd.n6982 585
R8600 gnd.n521 gnd.n520 585
R8601 gnd.n6981 gnd.n521 585
R8602 gnd.n6979 gnd.n6978 585
R8603 gnd.n6980 gnd.n6979 585
R8604 gnd.n524 gnd.n523 585
R8605 gnd.n523 gnd.n522 585
R8606 gnd.n6974 gnd.n6973 585
R8607 gnd.n6973 gnd.n6972 585
R8608 gnd.n527 gnd.n526 585
R8609 gnd.n6971 gnd.n527 585
R8610 gnd.n6969 gnd.n6968 585
R8611 gnd.n6970 gnd.n6969 585
R8612 gnd.n530 gnd.n529 585
R8613 gnd.n529 gnd.n528 585
R8614 gnd.n6964 gnd.n6963 585
R8615 gnd.n6963 gnd.n6962 585
R8616 gnd.n533 gnd.n532 585
R8617 gnd.n6961 gnd.n533 585
R8618 gnd.n6959 gnd.n6958 585
R8619 gnd.n6960 gnd.n6959 585
R8620 gnd.n536 gnd.n535 585
R8621 gnd.n535 gnd.n534 585
R8622 gnd.n6954 gnd.n6953 585
R8623 gnd.n6953 gnd.n6952 585
R8624 gnd.n539 gnd.n538 585
R8625 gnd.n6951 gnd.n539 585
R8626 gnd.n6949 gnd.n6948 585
R8627 gnd.n6950 gnd.n6949 585
R8628 gnd.n542 gnd.n541 585
R8629 gnd.n541 gnd.n540 585
R8630 gnd.n6944 gnd.n6943 585
R8631 gnd.n6943 gnd.n6942 585
R8632 gnd.n545 gnd.n544 585
R8633 gnd.n6941 gnd.n545 585
R8634 gnd.n6939 gnd.n6938 585
R8635 gnd.n6940 gnd.n6939 585
R8636 gnd.n6260 gnd.n6259 585
R8637 gnd.n6261 gnd.n6260 585
R8638 gnd.n1099 gnd.n1098 585
R8639 gnd.n4553 gnd.n1099 585
R8640 gnd.n6269 gnd.n6268 585
R8641 gnd.n6268 gnd.n6267 585
R8642 gnd.n6270 gnd.n1093 585
R8643 gnd.n4513 gnd.n1093 585
R8644 gnd.n6272 gnd.n6271 585
R8645 gnd.n6273 gnd.n6272 585
R8646 gnd.n1078 gnd.n1077 585
R8647 gnd.n4504 gnd.n1078 585
R8648 gnd.n6281 gnd.n6280 585
R8649 gnd.n6280 gnd.n6279 585
R8650 gnd.n6282 gnd.n1072 585
R8651 gnd.n4496 gnd.n1072 585
R8652 gnd.n6284 gnd.n6283 585
R8653 gnd.n6285 gnd.n6284 585
R8654 gnd.n1056 gnd.n1055 585
R8655 gnd.n4431 gnd.n1056 585
R8656 gnd.n6293 gnd.n6292 585
R8657 gnd.n6292 gnd.n6291 585
R8658 gnd.n6294 gnd.n1050 585
R8659 gnd.n4419 gnd.n1050 585
R8660 gnd.n6296 gnd.n6295 585
R8661 gnd.n6297 gnd.n6296 585
R8662 gnd.n1036 gnd.n1035 585
R8663 gnd.n4442 gnd.n1036 585
R8664 gnd.n6305 gnd.n6304 585
R8665 gnd.n6304 gnd.n6303 585
R8666 gnd.n6306 gnd.n1030 585
R8667 gnd.n4411 gnd.n1030 585
R8668 gnd.n6308 gnd.n6307 585
R8669 gnd.n6309 gnd.n6308 585
R8670 gnd.n1014 gnd.n1013 585
R8671 gnd.n4378 gnd.n1014 585
R8672 gnd.n6317 gnd.n6316 585
R8673 gnd.n6316 gnd.n6315 585
R8674 gnd.n6318 gnd.n1008 585
R8675 gnd.n4370 gnd.n1008 585
R8676 gnd.n6320 gnd.n6319 585
R8677 gnd.n6321 gnd.n6320 585
R8678 gnd.n994 gnd.n993 585
R8679 gnd.n4393 gnd.n994 585
R8680 gnd.n6329 gnd.n6328 585
R8681 gnd.n6328 gnd.n6327 585
R8682 gnd.n6330 gnd.n988 585
R8683 gnd.n4362 gnd.n988 585
R8684 gnd.n6332 gnd.n6331 585
R8685 gnd.n6333 gnd.n6332 585
R8686 gnd.n989 gnd.n987 585
R8687 gnd.n4344 gnd.n987 585
R8688 gnd.n4321 gnd.n974 585
R8689 gnd.n6339 gnd.n974 585
R8690 gnd.n4323 gnd.n4322 585
R8691 gnd.n4322 gnd.n970 585
R8692 gnd.n4324 gnd.n2171 585
R8693 gnd.n4335 gnd.n2171 585
R8694 gnd.n4325 gnd.n2180 585
R8695 gnd.n2180 gnd.n2178 585
R8696 gnd.n4327 gnd.n4326 585
R8697 gnd.n4328 gnd.n4327 585
R8698 gnd.n2181 gnd.n2179 585
R8699 gnd.n2196 gnd.n2179 585
R8700 gnd.n2197 gnd.n2183 585
R8701 gnd.n4309 gnd.n2197 585
R8702 gnd.n4298 gnd.n2205 585
R8703 gnd.n2205 gnd.n2194 585
R8704 gnd.n4300 gnd.n4299 585
R8705 gnd.n4301 gnd.n4300 585
R8706 gnd.n2206 gnd.n2204 585
R8707 gnd.n2204 gnd.n2201 585
R8708 gnd.n4294 gnd.n4293 585
R8709 gnd.n4293 gnd.n4292 585
R8710 gnd.n2209 gnd.n2208 585
R8711 gnd.n2210 gnd.n2209 585
R8712 gnd.n4283 gnd.n4282 585
R8713 gnd.n4284 gnd.n4283 585
R8714 gnd.n2220 gnd.n2219 585
R8715 gnd.n2227 gnd.n2219 585
R8716 gnd.n4278 gnd.n4277 585
R8717 gnd.n4277 gnd.n4276 585
R8718 gnd.n2223 gnd.n2222 585
R8719 gnd.n2224 gnd.n2223 585
R8720 gnd.n4266 gnd.n4265 585
R8721 gnd.n4267 gnd.n4266 585
R8722 gnd.n2237 gnd.n2236 585
R8723 gnd.n2236 gnd.n2233 585
R8724 gnd.n4261 gnd.n4260 585
R8725 gnd.n4260 gnd.n4259 585
R8726 gnd.n2240 gnd.n2239 585
R8727 gnd.n2241 gnd.n2240 585
R8728 gnd.n4250 gnd.n4249 585
R8729 gnd.n4251 gnd.n4250 585
R8730 gnd.n2252 gnd.n2251 585
R8731 gnd.n2259 gnd.n2251 585
R8732 gnd.n4245 gnd.n4244 585
R8733 gnd.n4244 gnd.n4243 585
R8734 gnd.n2255 gnd.n2254 585
R8735 gnd.n2256 gnd.n2255 585
R8736 gnd.n4234 gnd.n4233 585
R8737 gnd.n4235 gnd.n4234 585
R8738 gnd.n2269 gnd.n2268 585
R8739 gnd.n2268 gnd.n2265 585
R8740 gnd.n4229 gnd.n4228 585
R8741 gnd.n4228 gnd.n4227 585
R8742 gnd.n2272 gnd.n2271 585
R8743 gnd.n2273 gnd.n2272 585
R8744 gnd.n4218 gnd.n4217 585
R8745 gnd.n4219 gnd.n4218 585
R8746 gnd.n2284 gnd.n2283 585
R8747 gnd.n2291 gnd.n2283 585
R8748 gnd.n4213 gnd.n4212 585
R8749 gnd.n4212 gnd.n4211 585
R8750 gnd.n2287 gnd.n2286 585
R8751 gnd.n2288 gnd.n2287 585
R8752 gnd.n4202 gnd.n4201 585
R8753 gnd.n4203 gnd.n4202 585
R8754 gnd.n2301 gnd.n2300 585
R8755 gnd.n2300 gnd.n2297 585
R8756 gnd.n4197 gnd.n4196 585
R8757 gnd.n4196 gnd.n4195 585
R8758 gnd.n2304 gnd.n2303 585
R8759 gnd.n2305 gnd.n2304 585
R8760 gnd.n4186 gnd.n4185 585
R8761 gnd.n4187 gnd.n4186 585
R8762 gnd.n2316 gnd.n2315 585
R8763 gnd.n3957 gnd.n2315 585
R8764 gnd.n4181 gnd.n4180 585
R8765 gnd.n4180 gnd.n4179 585
R8766 gnd.n3816 gnd.n2318 585
R8767 gnd.n3819 gnd.n3817 585
R8768 gnd.n3822 gnd.n3821 585
R8769 gnd.n3814 gnd.n3813 585
R8770 gnd.n3827 gnd.n3826 585
R8771 gnd.n3829 gnd.n3812 585
R8772 gnd.n3832 gnd.n3831 585
R8773 gnd.n3810 gnd.n3809 585
R8774 gnd.n3837 gnd.n3836 585
R8775 gnd.n3839 gnd.n3808 585
R8776 gnd.n3842 gnd.n3841 585
R8777 gnd.n3806 gnd.n3805 585
R8778 gnd.n3847 gnd.n3846 585
R8779 gnd.n3849 gnd.n3804 585
R8780 gnd.n3852 gnd.n3851 585
R8781 gnd.n3802 gnd.n3801 585
R8782 gnd.n3857 gnd.n3856 585
R8783 gnd.n3859 gnd.n3800 585
R8784 gnd.n3861 gnd.n3860 585
R8785 gnd.n3860 gnd.n3793 585
R8786 gnd.n5357 gnd.n5356 585
R8787 gnd.n2026 gnd.n2018 585
R8788 gnd.n5364 gnd.n2015 585
R8789 gnd.n5365 gnd.n2014 585
R8790 gnd.n2040 gnd.n2008 585
R8791 gnd.n5372 gnd.n2007 585
R8792 gnd.n5373 gnd.n2006 585
R8793 gnd.n2038 gnd.n1998 585
R8794 gnd.n5380 gnd.n1997 585
R8795 gnd.n5381 gnd.n1996 585
R8796 gnd.n2035 gnd.n1990 585
R8797 gnd.n5388 gnd.n1989 585
R8798 gnd.n5389 gnd.n1988 585
R8799 gnd.n2033 gnd.n1981 585
R8800 gnd.n5396 gnd.n1980 585
R8801 gnd.n5397 gnd.n1979 585
R8802 gnd.n2030 gnd.n1978 585
R8803 gnd.n2029 gnd.n2028 585
R8804 gnd.n1115 gnd.n1113 585
R8805 gnd.n5354 gnd.n1113 585
R8806 gnd.n2111 gnd.n1111 585
R8807 gnd.n6261 gnd.n1111 585
R8808 gnd.n4552 gnd.n4551 585
R8809 gnd.n4553 gnd.n4552 585
R8810 gnd.n2110 gnd.n1102 585
R8811 gnd.n6267 gnd.n1102 585
R8812 gnd.n4515 gnd.n4514 585
R8813 gnd.n4514 gnd.n4513 585
R8814 gnd.n2113 gnd.n1091 585
R8815 gnd.n6273 gnd.n1091 585
R8816 gnd.n4503 gnd.n4502 585
R8817 gnd.n4504 gnd.n4503 585
R8818 gnd.n2117 gnd.n1080 585
R8819 gnd.n6279 gnd.n1080 585
R8820 gnd.n4498 gnd.n4497 585
R8821 gnd.n4497 gnd.n4496 585
R8822 gnd.n2119 gnd.n1070 585
R8823 gnd.n6285 gnd.n1070 585
R8824 gnd.n4434 gnd.n4432 585
R8825 gnd.n4432 gnd.n4431 585
R8826 gnd.n4435 gnd.n1059 585
R8827 gnd.n6291 gnd.n1059 585
R8828 gnd.n4436 gnd.n2136 585
R8829 gnd.n4419 gnd.n2136 585
R8830 gnd.n2133 gnd.n1048 585
R8831 gnd.n6297 gnd.n1048 585
R8832 gnd.n4441 gnd.n4440 585
R8833 gnd.n4442 gnd.n4441 585
R8834 gnd.n2132 gnd.n1038 585
R8835 gnd.n6303 gnd.n1038 585
R8836 gnd.n4381 gnd.n2142 585
R8837 gnd.n4411 gnd.n2142 585
R8838 gnd.n4380 gnd.n1028 585
R8839 gnd.n6309 gnd.n1028 585
R8840 gnd.n4385 gnd.n4379 585
R8841 gnd.n4379 gnd.n4378 585
R8842 gnd.n4386 gnd.n1017 585
R8843 gnd.n6315 gnd.n1017 585
R8844 gnd.n4387 gnd.n2157 585
R8845 gnd.n4370 gnd.n2157 585
R8846 gnd.n2154 gnd.n1006 585
R8847 gnd.n6321 gnd.n1006 585
R8848 gnd.n4392 gnd.n4391 585
R8849 gnd.n4393 gnd.n4392 585
R8850 gnd.n2153 gnd.n996 585
R8851 gnd.n6327 gnd.n996 585
R8852 gnd.n4351 gnd.n4350 585
R8853 gnd.n4362 gnd.n4351 585
R8854 gnd.n2163 gnd.n985 585
R8855 gnd.n6333 gnd.n985 585
R8856 gnd.n4346 gnd.n4345 585
R8857 gnd.n4345 gnd.n4344 585
R8858 gnd.n2165 gnd.n972 585
R8859 gnd.n6339 gnd.n972 585
R8860 gnd.n3900 gnd.n3899 585
R8861 gnd.n3899 gnd.n970 585
R8862 gnd.n3903 gnd.n2170 585
R8863 gnd.n4335 gnd.n2170 585
R8864 gnd.n3904 gnd.n3898 585
R8865 gnd.n3898 gnd.n2178 585
R8866 gnd.n3905 gnd.n2176 585
R8867 gnd.n4328 gnd.n2176 585
R8868 gnd.n3896 gnd.n3895 585
R8869 gnd.n3895 gnd.n2196 585
R8870 gnd.n3909 gnd.n2195 585
R8871 gnd.n4309 gnd.n2195 585
R8872 gnd.n3911 gnd.n3910 585
R8873 gnd.n3910 gnd.n2194 585
R8874 gnd.n3912 gnd.n2203 585
R8875 gnd.n4301 gnd.n2203 585
R8876 gnd.n3914 gnd.n3913 585
R8877 gnd.n3913 gnd.n2201 585
R8878 gnd.n3915 gnd.n2212 585
R8879 gnd.n4292 gnd.n2212 585
R8880 gnd.n3917 gnd.n3916 585
R8881 gnd.n3916 gnd.n2210 585
R8882 gnd.n3918 gnd.n2218 585
R8883 gnd.n4284 gnd.n2218 585
R8884 gnd.n3920 gnd.n3919 585
R8885 gnd.n3919 gnd.n2227 585
R8886 gnd.n3921 gnd.n2226 585
R8887 gnd.n4276 gnd.n2226 585
R8888 gnd.n3923 gnd.n3922 585
R8889 gnd.n3922 gnd.n2224 585
R8890 gnd.n3924 gnd.n2235 585
R8891 gnd.n4267 gnd.n2235 585
R8892 gnd.n3926 gnd.n3925 585
R8893 gnd.n3925 gnd.n2233 585
R8894 gnd.n3927 gnd.n2243 585
R8895 gnd.n4259 gnd.n2243 585
R8896 gnd.n3929 gnd.n3928 585
R8897 gnd.n3928 gnd.n2241 585
R8898 gnd.n3930 gnd.n2250 585
R8899 gnd.n4251 gnd.n2250 585
R8900 gnd.n3932 gnd.n3931 585
R8901 gnd.n3931 gnd.n2259 585
R8902 gnd.n3933 gnd.n2258 585
R8903 gnd.n4243 gnd.n2258 585
R8904 gnd.n3935 gnd.n3934 585
R8905 gnd.n3934 gnd.n2256 585
R8906 gnd.n3936 gnd.n2267 585
R8907 gnd.n4235 gnd.n2267 585
R8908 gnd.n3938 gnd.n3937 585
R8909 gnd.n3937 gnd.n2265 585
R8910 gnd.n3939 gnd.n2275 585
R8911 gnd.n4227 gnd.n2275 585
R8912 gnd.n3941 gnd.n3940 585
R8913 gnd.n3940 gnd.n2273 585
R8914 gnd.n3942 gnd.n2282 585
R8915 gnd.n4219 gnd.n2282 585
R8916 gnd.n3944 gnd.n3943 585
R8917 gnd.n3943 gnd.n2291 585
R8918 gnd.n3945 gnd.n2290 585
R8919 gnd.n4211 gnd.n2290 585
R8920 gnd.n3947 gnd.n3946 585
R8921 gnd.n3946 gnd.n2288 585
R8922 gnd.n3948 gnd.n2299 585
R8923 gnd.n4203 gnd.n2299 585
R8924 gnd.n3950 gnd.n3949 585
R8925 gnd.n3949 gnd.n2297 585
R8926 gnd.n3951 gnd.n2307 585
R8927 gnd.n4195 gnd.n2307 585
R8928 gnd.n3953 gnd.n3952 585
R8929 gnd.n3952 gnd.n2305 585
R8930 gnd.n3954 gnd.n2314 585
R8931 gnd.n4187 gnd.n2314 585
R8932 gnd.n3956 gnd.n3955 585
R8933 gnd.n3957 gnd.n3956 585
R8934 gnd.n3796 gnd.n3795 585
R8935 gnd.n4179 gnd.n3795 585
R8936 gnd.n7506 gnd.n129 585
R8937 gnd.n7602 gnd.n129 585
R8938 gnd.n7507 gnd.n7444 585
R8939 gnd.n7444 gnd.n126 585
R8940 gnd.n7508 gnd.n207 585
R8941 gnd.n7522 gnd.n207 585
R8942 gnd.n219 gnd.n217 585
R8943 gnd.n217 gnd.n206 585
R8944 gnd.n7513 gnd.n7512 585
R8945 gnd.n7514 gnd.n7513 585
R8946 gnd.n218 gnd.n216 585
R8947 gnd.n216 gnd.n213 585
R8948 gnd.n7440 gnd.n7439 585
R8949 gnd.n7439 gnd.n7438 585
R8950 gnd.n222 gnd.n221 585
R8951 gnd.n232 gnd.n222 585
R8952 gnd.n7429 gnd.n7428 585
R8953 gnd.n7430 gnd.n7429 585
R8954 gnd.n234 gnd.n233 585
R8955 gnd.n233 gnd.n229 585
R8956 gnd.n7424 gnd.n7423 585
R8957 gnd.n7423 gnd.n7422 585
R8958 gnd.n237 gnd.n236 585
R8959 gnd.n247 gnd.n237 585
R8960 gnd.n7413 gnd.n7412 585
R8961 gnd.n7414 gnd.n7413 585
R8962 gnd.n249 gnd.n248 585
R8963 gnd.n254 gnd.n248 585
R8964 gnd.n7408 gnd.n7407 585
R8965 gnd.n7407 gnd.n7406 585
R8966 gnd.n252 gnd.n251 585
R8967 gnd.n263 gnd.n252 585
R8968 gnd.n7397 gnd.n7396 585
R8969 gnd.n7398 gnd.n7397 585
R8970 gnd.n265 gnd.n264 585
R8971 gnd.n264 gnd.n260 585
R8972 gnd.n7392 gnd.n7391 585
R8973 gnd.n7391 gnd.n7390 585
R8974 gnd.n268 gnd.n267 585
R8975 gnd.n269 gnd.n268 585
R8976 gnd.n7381 gnd.n7380 585
R8977 gnd.n7382 gnd.n7381 585
R8978 gnd.n279 gnd.n278 585
R8979 gnd.n284 gnd.n278 585
R8980 gnd.n7376 gnd.n7375 585
R8981 gnd.n7375 gnd.n7374 585
R8982 gnd.n282 gnd.n281 585
R8983 gnd.n293 gnd.n282 585
R8984 gnd.n7365 gnd.n7364 585
R8985 gnd.n7366 gnd.n7365 585
R8986 gnd.n295 gnd.n294 585
R8987 gnd.n294 gnd.n290 585
R8988 gnd.n7360 gnd.n7359 585
R8989 gnd.n7359 gnd.n7358 585
R8990 gnd.n298 gnd.n297 585
R8991 gnd.n299 gnd.n298 585
R8992 gnd.n7336 gnd.n7335 585
R8993 gnd.n7335 gnd.n7334 585
R8994 gnd.n7337 gnd.n327 585
R8995 gnd.n7330 gnd.n327 585
R8996 gnd.n333 gnd.n325 585
R8997 gnd.n334 gnd.n333 585
R8998 gnd.n7341 gnd.n324 585
R8999 gnd.n7257 gnd.n324 585
R9000 gnd.n7342 gnd.n323 585
R9001 gnd.n340 gnd.n323 585
R9002 gnd.n7343 gnd.n322 585
R9003 gnd.n7251 gnd.n322 585
R9004 gnd.n319 gnd.n317 585
R9005 gnd.n317 gnd.n315 585
R9006 gnd.n7348 gnd.n7347 585
R9007 gnd.n7349 gnd.n7348 585
R9008 gnd.n318 gnd.n316 585
R9009 gnd.n7242 gnd.n316 585
R9010 gnd.n7210 gnd.n7208 585
R9011 gnd.n7208 gnd.n350 585
R9012 gnd.n7211 gnd.n359 585
R9013 gnd.n7227 gnd.n359 585
R9014 gnd.n7212 gnd.n7207 585
R9015 gnd.n7207 gnd.n7206 585
R9016 gnd.n374 gnd.n372 585
R9017 gnd.n7190 gnd.n372 585
R9018 gnd.n7217 gnd.n7216 585
R9019 gnd.n7218 gnd.n7217 585
R9020 gnd.n373 gnd.n371 585
R9021 gnd.n7196 gnd.n371 585
R9022 gnd.n7165 gnd.n7164 585
R9023 gnd.n7164 gnd.n7163 585
R9024 gnd.n7166 gnd.n392 585
R9025 gnd.n7182 gnd.n392 585
R9026 gnd.n406 gnd.n404 585
R9027 gnd.n5941 gnd.n404 585
R9028 gnd.n7171 gnd.n7170 585
R9029 gnd.n7172 gnd.n7171 585
R9030 gnd.n405 gnd.n403 585
R9031 gnd.n5936 gnd.n403 585
R9032 gnd.n5990 gnd.n5988 585
R9033 gnd.n5988 gnd.n5987 585
R9034 gnd.n5991 gnd.n1360 585
R9035 gnd.n1373 gnd.n1360 585
R9036 gnd.n5992 gnd.n1359 585
R9037 gnd.n5979 gnd.n1359 585
R9038 gnd.n5956 gnd.n1357 585
R9039 gnd.n5957 gnd.n5956 585
R9040 gnd.n5996 gnd.n1356 585
R9041 gnd.n1398 gnd.n1356 585
R9042 gnd.n5997 gnd.n1355 585
R9043 gnd.n5919 gnd.n1355 585
R9044 gnd.n5998 gnd.n1354 585
R9045 gnd.n1407 gnd.n1354 585
R9046 gnd.n5908 gnd.n1352 585
R9047 gnd.n5909 gnd.n5908 585
R9048 gnd.n6002 gnd.n1351 585
R9049 gnd.n5896 gnd.n1351 585
R9050 gnd.n6003 gnd.n1350 585
R9051 gnd.n1414 gnd.n1350 585
R9052 gnd.n6004 gnd.n1349 585
R9053 gnd.n5882 gnd.n1349 585
R9054 gnd.n1434 gnd.n1347 585
R9055 gnd.n1435 gnd.n1434 585
R9056 gnd.n6008 gnd.n1346 585
R9057 gnd.n5872 gnd.n1346 585
R9058 gnd.n6009 gnd.n1345 585
R9059 gnd.n5860 gnd.n1345 585
R9060 gnd.n6010 gnd.n1344 585
R9061 gnd.n1452 gnd.n1344 585
R9062 gnd.n1341 gnd.n1340 585
R9063 gnd.n5851 gnd.n1340 585
R9064 gnd.n6015 gnd.n6014 585
R9065 gnd.n6016 gnd.n6015 585
R9066 gnd.n1517 gnd.n1339 585
R9067 gnd.n1522 gnd.n1521 585
R9068 gnd.n1524 gnd.n1523 585
R9069 gnd.n1527 gnd.n1526 585
R9070 gnd.n1525 gnd.n1510 585
R9071 gnd.n1541 gnd.n1540 585
R9072 gnd.n1543 gnd.n1542 585
R9073 gnd.n1546 gnd.n1545 585
R9074 gnd.n1544 gnd.n1503 585
R9075 gnd.n1560 gnd.n1559 585
R9076 gnd.n1562 gnd.n1561 585
R9077 gnd.n1565 gnd.n1564 585
R9078 gnd.n1563 gnd.n1496 585
R9079 gnd.n1578 gnd.n1577 585
R9080 gnd.n1580 gnd.n1579 585
R9081 gnd.n1489 gnd.n1488 585
R9082 gnd.n1593 gnd.n1490 585
R9083 gnd.n1594 gnd.n1485 585
R9084 gnd.n1595 gnd.n1284 585
R9085 gnd.n6092 gnd.n1284 585
R9086 gnd.n7605 gnd.n7604 585
R9087 gnd.n7477 gnd.n124 585
R9088 gnd.n7479 gnd.n7478 585
R9089 gnd.n7475 gnd.n7474 585
R9090 gnd.n7483 gnd.n7473 585
R9091 gnd.n7484 gnd.n7471 585
R9092 gnd.n7485 gnd.n7470 585
R9093 gnd.n7468 gnd.n7466 585
R9094 gnd.n7489 gnd.n7465 585
R9095 gnd.n7490 gnd.n7463 585
R9096 gnd.n7491 gnd.n7462 585
R9097 gnd.n7460 gnd.n7458 585
R9098 gnd.n7495 gnd.n7457 585
R9099 gnd.n7496 gnd.n7455 585
R9100 gnd.n7497 gnd.n7454 585
R9101 gnd.n7452 gnd.n7450 585
R9102 gnd.n7501 gnd.n7449 585
R9103 gnd.n7502 gnd.n7447 585
R9104 gnd.n7503 gnd.n7446 585
R9105 gnd.n7446 gnd.n128 585
R9106 gnd.n7603 gnd.n120 585
R9107 gnd.n7603 gnd.n7602 585
R9108 gnd.n7609 gnd.n119 585
R9109 gnd.n126 gnd.n119 585
R9110 gnd.n7610 gnd.n118 585
R9111 gnd.n7522 gnd.n118 585
R9112 gnd.n7611 gnd.n117 585
R9113 gnd.n206 gnd.n117 585
R9114 gnd.n215 gnd.n115 585
R9115 gnd.n7514 gnd.n215 585
R9116 gnd.n7615 gnd.n114 585
R9117 gnd.n213 gnd.n114 585
R9118 gnd.n7616 gnd.n113 585
R9119 gnd.n7438 gnd.n113 585
R9120 gnd.n7617 gnd.n112 585
R9121 gnd.n232 gnd.n112 585
R9122 gnd.n231 gnd.n110 585
R9123 gnd.n7430 gnd.n231 585
R9124 gnd.n7621 gnd.n109 585
R9125 gnd.n229 gnd.n109 585
R9126 gnd.n7622 gnd.n108 585
R9127 gnd.n7422 gnd.n108 585
R9128 gnd.n7623 gnd.n107 585
R9129 gnd.n247 gnd.n107 585
R9130 gnd.n246 gnd.n105 585
R9131 gnd.n7414 gnd.n246 585
R9132 gnd.n7627 gnd.n104 585
R9133 gnd.n254 gnd.n104 585
R9134 gnd.n7628 gnd.n103 585
R9135 gnd.n7406 gnd.n103 585
R9136 gnd.n7629 gnd.n102 585
R9137 gnd.n263 gnd.n102 585
R9138 gnd.n262 gnd.n100 585
R9139 gnd.n7398 gnd.n262 585
R9140 gnd.n7633 gnd.n99 585
R9141 gnd.n260 gnd.n99 585
R9142 gnd.n7634 gnd.n98 585
R9143 gnd.n7390 gnd.n98 585
R9144 gnd.n7635 gnd.n97 585
R9145 gnd.n269 gnd.n97 585
R9146 gnd.n277 gnd.n95 585
R9147 gnd.n7382 gnd.n277 585
R9148 gnd.n7639 gnd.n94 585
R9149 gnd.n284 gnd.n94 585
R9150 gnd.n7640 gnd.n93 585
R9151 gnd.n7374 gnd.n93 585
R9152 gnd.n7641 gnd.n92 585
R9153 gnd.n293 gnd.n92 585
R9154 gnd.n292 gnd.n90 585
R9155 gnd.n7366 gnd.n292 585
R9156 gnd.n7645 gnd.n89 585
R9157 gnd.n290 gnd.n89 585
R9158 gnd.n7646 gnd.n88 585
R9159 gnd.n7358 gnd.n88 585
R9160 gnd.n7647 gnd.n87 585
R9161 gnd.n299 gnd.n87 585
R9162 gnd.n329 gnd.n85 585
R9163 gnd.n7334 gnd.n329 585
R9164 gnd.n7651 gnd.n84 585
R9165 gnd.n7330 gnd.n84 585
R9166 gnd.n7652 gnd.n83 585
R9167 gnd.n334 gnd.n83 585
R9168 gnd.n7653 gnd.n82 585
R9169 gnd.n7257 gnd.n82 585
R9170 gnd.n345 gnd.n80 585
R9171 gnd.n345 gnd.n340 585
R9172 gnd.n7250 gnd.n7249 585
R9173 gnd.n7251 gnd.n7250 585
R9174 gnd.n7248 gnd.n344 585
R9175 gnd.n344 gnd.n315 585
R9176 gnd.n346 gnd.n314 585
R9177 gnd.n7349 gnd.n314 585
R9178 gnd.n7244 gnd.n7243 585
R9179 gnd.n7243 gnd.n7242 585
R9180 gnd.n349 gnd.n348 585
R9181 gnd.n350 gnd.n349 585
R9182 gnd.n380 gnd.n357 585
R9183 gnd.n7227 gnd.n357 585
R9184 gnd.n7205 gnd.n7204 585
R9185 gnd.n7206 gnd.n7205 585
R9186 gnd.n379 gnd.n378 585
R9187 gnd.n7190 gnd.n378 585
R9188 gnd.n7199 gnd.n369 585
R9189 gnd.n7218 gnd.n369 585
R9190 gnd.n7198 gnd.n7197 585
R9191 gnd.n7197 gnd.n7196 585
R9192 gnd.n383 gnd.n382 585
R9193 gnd.n7163 gnd.n383 585
R9194 gnd.n5943 gnd.n391 585
R9195 gnd.n7182 gnd.n391 585
R9196 gnd.n5944 gnd.n5942 585
R9197 gnd.n5942 gnd.n5941 585
R9198 gnd.n5938 gnd.n401 585
R9199 gnd.n7172 gnd.n401 585
R9200 gnd.n5948 gnd.n5937 585
R9201 gnd.n5937 gnd.n5936 585
R9202 gnd.n5949 gnd.n1363 585
R9203 gnd.n5987 gnd.n1363 585
R9204 gnd.n5950 gnd.n1386 585
R9205 gnd.n1386 gnd.n1373 585
R9206 gnd.n1383 gnd.n1372 585
R9207 gnd.n5979 gnd.n1372 585
R9208 gnd.n5955 gnd.n5954 585
R9209 gnd.n5957 gnd.n5955 585
R9210 gnd.n1382 gnd.n1381 585
R9211 gnd.n1398 gnd.n1381 585
R9212 gnd.n5889 gnd.n1395 585
R9213 gnd.n5919 gnd.n1395 585
R9214 gnd.n5890 gnd.n5888 585
R9215 gnd.n5888 gnd.n1407 585
R9216 gnd.n1418 gnd.n1406 585
R9217 gnd.n5909 gnd.n1406 585
R9218 gnd.n5895 gnd.n5894 585
R9219 gnd.n5896 gnd.n5895 585
R9220 gnd.n1417 gnd.n1416 585
R9221 gnd.n1416 gnd.n1414 585
R9222 gnd.n5884 gnd.n5883 585
R9223 gnd.n5883 gnd.n5882 585
R9224 gnd.n1421 gnd.n1420 585
R9225 gnd.n1435 gnd.n1421 585
R9226 gnd.n1477 gnd.n1433 585
R9227 gnd.n5872 gnd.n1433 585
R9228 gnd.n5859 gnd.n5858 585
R9229 gnd.n5860 gnd.n5859 585
R9230 gnd.n1476 gnd.n1475 585
R9231 gnd.n1475 gnd.n1452 585
R9232 gnd.n5853 gnd.n5852 585
R9233 gnd.n5852 gnd.n5851 585
R9234 gnd.n5841 gnd.n1337 585
R9235 gnd.n6016 gnd.n1337 585
R9236 gnd.n3700 gnd.n3699 585
R9237 gnd.n3701 gnd.n3700 585
R9238 gnd.n2395 gnd.n2394 585
R9239 gnd.n2401 gnd.n2394 585
R9240 gnd.n3675 gnd.n2413 585
R9241 gnd.n2413 gnd.n2400 585
R9242 gnd.n3677 gnd.n3676 585
R9243 gnd.n3678 gnd.n3677 585
R9244 gnd.n2414 gnd.n2412 585
R9245 gnd.n2412 gnd.n2408 585
R9246 gnd.n3409 gnd.n3408 585
R9247 gnd.n3408 gnd.n3407 585
R9248 gnd.n2419 gnd.n2418 585
R9249 gnd.n3378 gnd.n2419 585
R9250 gnd.n3398 gnd.n3397 585
R9251 gnd.n3397 gnd.n3396 585
R9252 gnd.n2426 gnd.n2425 585
R9253 gnd.n3384 gnd.n2426 585
R9254 gnd.n3354 gnd.n2446 585
R9255 gnd.n2446 gnd.n2445 585
R9256 gnd.n3356 gnd.n3355 585
R9257 gnd.n3357 gnd.n3356 585
R9258 gnd.n2447 gnd.n2444 585
R9259 gnd.n2455 gnd.n2444 585
R9260 gnd.n3332 gnd.n2467 585
R9261 gnd.n2467 gnd.n2454 585
R9262 gnd.n3334 gnd.n3333 585
R9263 gnd.n3335 gnd.n3334 585
R9264 gnd.n2468 gnd.n2466 585
R9265 gnd.n2466 gnd.n2462 585
R9266 gnd.n3320 gnd.n3319 585
R9267 gnd.n3319 gnd.n3318 585
R9268 gnd.n2473 gnd.n2472 585
R9269 gnd.n2483 gnd.n2473 585
R9270 gnd.n3309 gnd.n3308 585
R9271 gnd.n3308 gnd.n3307 585
R9272 gnd.n2480 gnd.n2479 585
R9273 gnd.n3295 gnd.n2480 585
R9274 gnd.n3269 gnd.n2501 585
R9275 gnd.n2501 gnd.n2490 585
R9276 gnd.n3271 gnd.n3270 585
R9277 gnd.n3272 gnd.n3271 585
R9278 gnd.n2502 gnd.n2500 585
R9279 gnd.n2510 gnd.n2500 585
R9280 gnd.n3247 gnd.n2522 585
R9281 gnd.n2522 gnd.n2509 585
R9282 gnd.n3249 gnd.n3248 585
R9283 gnd.n3250 gnd.n3249 585
R9284 gnd.n2523 gnd.n2521 585
R9285 gnd.n2521 gnd.n2517 585
R9286 gnd.n3235 gnd.n3234 585
R9287 gnd.n3234 gnd.n3233 585
R9288 gnd.n2528 gnd.n2527 585
R9289 gnd.n2537 gnd.n2528 585
R9290 gnd.n3224 gnd.n3223 585
R9291 gnd.n3223 gnd.n3222 585
R9292 gnd.n2535 gnd.n2534 585
R9293 gnd.n3210 gnd.n2535 585
R9294 gnd.n2648 gnd.n2647 585
R9295 gnd.n2648 gnd.n2544 585
R9296 gnd.n3167 gnd.n3166 585
R9297 gnd.n3166 gnd.n3165 585
R9298 gnd.n3168 gnd.n2642 585
R9299 gnd.n2653 gnd.n2642 585
R9300 gnd.n3170 gnd.n3169 585
R9301 gnd.n3171 gnd.n3170 585
R9302 gnd.n2643 gnd.n2641 585
R9303 gnd.n2666 gnd.n2641 585
R9304 gnd.n2626 gnd.n2625 585
R9305 gnd.n2629 gnd.n2626 585
R9306 gnd.n3181 gnd.n3180 585
R9307 gnd.n3180 gnd.n3179 585
R9308 gnd.n3182 gnd.n2620 585
R9309 gnd.n3141 gnd.n2620 585
R9310 gnd.n3184 gnd.n3183 585
R9311 gnd.n3185 gnd.n3184 585
R9312 gnd.n2621 gnd.n2619 585
R9313 gnd.n2680 gnd.n2619 585
R9314 gnd.n3133 gnd.n3132 585
R9315 gnd.n3132 gnd.n3131 585
R9316 gnd.n2677 gnd.n2676 585
R9317 gnd.n3115 gnd.n2677 585
R9318 gnd.n3102 gnd.n2696 585
R9319 gnd.n2696 gnd.n2695 585
R9320 gnd.n3104 gnd.n3103 585
R9321 gnd.n3105 gnd.n3104 585
R9322 gnd.n2697 gnd.n2694 585
R9323 gnd.n2703 gnd.n2694 585
R9324 gnd.n3083 gnd.n3082 585
R9325 gnd.n3084 gnd.n3083 585
R9326 gnd.n2714 gnd.n2713 585
R9327 gnd.n2713 gnd.n2709 585
R9328 gnd.n3073 gnd.n3072 585
R9329 gnd.n3074 gnd.n3073 585
R9330 gnd.n2724 gnd.n2723 585
R9331 gnd.n2729 gnd.n2723 585
R9332 gnd.n3051 gnd.n2742 585
R9333 gnd.n2742 gnd.n2728 585
R9334 gnd.n3053 gnd.n3052 585
R9335 gnd.n3054 gnd.n3053 585
R9336 gnd.n2743 gnd.n2741 585
R9337 gnd.n2741 gnd.n2737 585
R9338 gnd.n3042 gnd.n3041 585
R9339 gnd.n3043 gnd.n3042 585
R9340 gnd.n2750 gnd.n2749 585
R9341 gnd.n2754 gnd.n2749 585
R9342 gnd.n3019 gnd.n2771 585
R9343 gnd.n2771 gnd.n2753 585
R9344 gnd.n3021 gnd.n3020 585
R9345 gnd.n3022 gnd.n3021 585
R9346 gnd.n2772 gnd.n2770 585
R9347 gnd.n2770 gnd.n2761 585
R9348 gnd.n3014 gnd.n3013 585
R9349 gnd.n3013 gnd.n3012 585
R9350 gnd.n2819 gnd.n2818 585
R9351 gnd.n2820 gnd.n2819 585
R9352 gnd.n2973 gnd.n2972 585
R9353 gnd.n2974 gnd.n2973 585
R9354 gnd.n2829 gnd.n2828 585
R9355 gnd.n2828 gnd.n2827 585
R9356 gnd.n2968 gnd.n2967 585
R9357 gnd.n2967 gnd.n2966 585
R9358 gnd.n2832 gnd.n2831 585
R9359 gnd.n2833 gnd.n2832 585
R9360 gnd.n2957 gnd.n2956 585
R9361 gnd.n2958 gnd.n2957 585
R9362 gnd.n2840 gnd.n2839 585
R9363 gnd.n2949 gnd.n2839 585
R9364 gnd.n2952 gnd.n2951 585
R9365 gnd.n2951 gnd.n2950 585
R9366 gnd.n2843 gnd.n2842 585
R9367 gnd.n2844 gnd.n2843 585
R9368 gnd.n2938 gnd.n2937 585
R9369 gnd.n2936 gnd.n2862 585
R9370 gnd.n2935 gnd.n2861 585
R9371 gnd.n2940 gnd.n2861 585
R9372 gnd.n2934 gnd.n2933 585
R9373 gnd.n2932 gnd.n2931 585
R9374 gnd.n2930 gnd.n2929 585
R9375 gnd.n2928 gnd.n2927 585
R9376 gnd.n2926 gnd.n2925 585
R9377 gnd.n2924 gnd.n2923 585
R9378 gnd.n2922 gnd.n2921 585
R9379 gnd.n2920 gnd.n2919 585
R9380 gnd.n2918 gnd.n2917 585
R9381 gnd.n2916 gnd.n2915 585
R9382 gnd.n2914 gnd.n2913 585
R9383 gnd.n2912 gnd.n2911 585
R9384 gnd.n2910 gnd.n2909 585
R9385 gnd.n2908 gnd.n2907 585
R9386 gnd.n2906 gnd.n2905 585
R9387 gnd.n2904 gnd.n2903 585
R9388 gnd.n2902 gnd.n2901 585
R9389 gnd.n2900 gnd.n2899 585
R9390 gnd.n2898 gnd.n2897 585
R9391 gnd.n2896 gnd.n2895 585
R9392 gnd.n2894 gnd.n2893 585
R9393 gnd.n2892 gnd.n2891 585
R9394 gnd.n2849 gnd.n2848 585
R9395 gnd.n2943 gnd.n2942 585
R9396 gnd.n3704 gnd.n3703 585
R9397 gnd.n3706 gnd.n3705 585
R9398 gnd.n3708 gnd.n3707 585
R9399 gnd.n3710 gnd.n3709 585
R9400 gnd.n3712 gnd.n3711 585
R9401 gnd.n3714 gnd.n3713 585
R9402 gnd.n3716 gnd.n3715 585
R9403 gnd.n3718 gnd.n3717 585
R9404 gnd.n3720 gnd.n3719 585
R9405 gnd.n3722 gnd.n3721 585
R9406 gnd.n3724 gnd.n3723 585
R9407 gnd.n3726 gnd.n3725 585
R9408 gnd.n3728 gnd.n3727 585
R9409 gnd.n3730 gnd.n3729 585
R9410 gnd.n3732 gnd.n3731 585
R9411 gnd.n3734 gnd.n3733 585
R9412 gnd.n3736 gnd.n3735 585
R9413 gnd.n3738 gnd.n3737 585
R9414 gnd.n3740 gnd.n3739 585
R9415 gnd.n3742 gnd.n3741 585
R9416 gnd.n3744 gnd.n3743 585
R9417 gnd.n3746 gnd.n3745 585
R9418 gnd.n3748 gnd.n3747 585
R9419 gnd.n3750 gnd.n3749 585
R9420 gnd.n3752 gnd.n3751 585
R9421 gnd.n3753 gnd.n2361 585
R9422 gnd.n3754 gnd.n2319 585
R9423 gnd.n3792 gnd.n2319 585
R9424 gnd.n3702 gnd.n2391 585
R9425 gnd.n3702 gnd.n3701 585
R9426 gnd.n3371 gnd.n2390 585
R9427 gnd.n2401 gnd.n2390 585
R9428 gnd.n3373 gnd.n3372 585
R9429 gnd.n3372 gnd.n2400 585
R9430 gnd.n3374 gnd.n2410 585
R9431 gnd.n3678 gnd.n2410 585
R9432 gnd.n3376 gnd.n3375 585
R9433 gnd.n3375 gnd.n2408 585
R9434 gnd.n3377 gnd.n2421 585
R9435 gnd.n3407 gnd.n2421 585
R9436 gnd.n3380 gnd.n3379 585
R9437 gnd.n3379 gnd.n3378 585
R9438 gnd.n3381 gnd.n2428 585
R9439 gnd.n3396 gnd.n2428 585
R9440 gnd.n3383 gnd.n3382 585
R9441 gnd.n3384 gnd.n3383 585
R9442 gnd.n2438 gnd.n2437 585
R9443 gnd.n2445 gnd.n2437 585
R9444 gnd.n3359 gnd.n3358 585
R9445 gnd.n3358 gnd.n3357 585
R9446 gnd.n2441 gnd.n2440 585
R9447 gnd.n2455 gnd.n2441 585
R9448 gnd.n3285 gnd.n3284 585
R9449 gnd.n3284 gnd.n2454 585
R9450 gnd.n3286 gnd.n2464 585
R9451 gnd.n3335 gnd.n2464 585
R9452 gnd.n3288 gnd.n3287 585
R9453 gnd.n3287 gnd.n2462 585
R9454 gnd.n3289 gnd.n2475 585
R9455 gnd.n3318 gnd.n2475 585
R9456 gnd.n3291 gnd.n3290 585
R9457 gnd.n3290 gnd.n2483 585
R9458 gnd.n3292 gnd.n2482 585
R9459 gnd.n3307 gnd.n2482 585
R9460 gnd.n3294 gnd.n3293 585
R9461 gnd.n3295 gnd.n3294 585
R9462 gnd.n2494 gnd.n2493 585
R9463 gnd.n2493 gnd.n2490 585
R9464 gnd.n3274 gnd.n3273 585
R9465 gnd.n3273 gnd.n3272 585
R9466 gnd.n2497 gnd.n2496 585
R9467 gnd.n2510 gnd.n2497 585
R9468 gnd.n3198 gnd.n3197 585
R9469 gnd.n3197 gnd.n2509 585
R9470 gnd.n3199 gnd.n2519 585
R9471 gnd.n3250 gnd.n2519 585
R9472 gnd.n3201 gnd.n3200 585
R9473 gnd.n3200 gnd.n2517 585
R9474 gnd.n3202 gnd.n2530 585
R9475 gnd.n3233 gnd.n2530 585
R9476 gnd.n3204 gnd.n3203 585
R9477 gnd.n3203 gnd.n2537 585
R9478 gnd.n3205 gnd.n2536 585
R9479 gnd.n3222 gnd.n2536 585
R9480 gnd.n3207 gnd.n3206 585
R9481 gnd.n3210 gnd.n3207 585
R9482 gnd.n2547 gnd.n2546 585
R9483 gnd.n2546 gnd.n2544 585
R9484 gnd.n2650 gnd.n2649 585
R9485 gnd.n3165 gnd.n2649 585
R9486 gnd.n2652 gnd.n2651 585
R9487 gnd.n2653 gnd.n2652 585
R9488 gnd.n2663 gnd.n2639 585
R9489 gnd.n3171 gnd.n2639 585
R9490 gnd.n2665 gnd.n2664 585
R9491 gnd.n2666 gnd.n2665 585
R9492 gnd.n2662 gnd.n2661 585
R9493 gnd.n2662 gnd.n2629 585
R9494 gnd.n2660 gnd.n2627 585
R9495 gnd.n3179 gnd.n2627 585
R9496 gnd.n2616 gnd.n2614 585
R9497 gnd.n3141 gnd.n2616 585
R9498 gnd.n3187 gnd.n3186 585
R9499 gnd.n3186 gnd.n3185 585
R9500 gnd.n2615 gnd.n2613 585
R9501 gnd.n2680 gnd.n2615 585
R9502 gnd.n3112 gnd.n2679 585
R9503 gnd.n3131 gnd.n2679 585
R9504 gnd.n3114 gnd.n3113 585
R9505 gnd.n3115 gnd.n3114 585
R9506 gnd.n2689 gnd.n2688 585
R9507 gnd.n2695 gnd.n2688 585
R9508 gnd.n3107 gnd.n3106 585
R9509 gnd.n3106 gnd.n3105 585
R9510 gnd.n2692 gnd.n2691 585
R9511 gnd.n2703 gnd.n2692 585
R9512 gnd.n2992 gnd.n2711 585
R9513 gnd.n3084 gnd.n2711 585
R9514 gnd.n2994 gnd.n2993 585
R9515 gnd.n2993 gnd.n2709 585
R9516 gnd.n2995 gnd.n2722 585
R9517 gnd.n3074 gnd.n2722 585
R9518 gnd.n2997 gnd.n2996 585
R9519 gnd.n2997 gnd.n2729 585
R9520 gnd.n2999 gnd.n2998 585
R9521 gnd.n2998 gnd.n2728 585
R9522 gnd.n3000 gnd.n2739 585
R9523 gnd.n3054 gnd.n2739 585
R9524 gnd.n3002 gnd.n3001 585
R9525 gnd.n3001 gnd.n2737 585
R9526 gnd.n3003 gnd.n2748 585
R9527 gnd.n3043 gnd.n2748 585
R9528 gnd.n3005 gnd.n3004 585
R9529 gnd.n3005 gnd.n2754 585
R9530 gnd.n3007 gnd.n3006 585
R9531 gnd.n3006 gnd.n2753 585
R9532 gnd.n3008 gnd.n2769 585
R9533 gnd.n3022 gnd.n2769 585
R9534 gnd.n3009 gnd.n2822 585
R9535 gnd.n2822 gnd.n2761 585
R9536 gnd.n3011 gnd.n3010 585
R9537 gnd.n3012 gnd.n3011 585
R9538 gnd.n2823 gnd.n2821 585
R9539 gnd.n2821 gnd.n2820 585
R9540 gnd.n2976 gnd.n2975 585
R9541 gnd.n2975 gnd.n2974 585
R9542 gnd.n2826 gnd.n2825 585
R9543 gnd.n2827 gnd.n2826 585
R9544 gnd.n2965 gnd.n2964 585
R9545 gnd.n2966 gnd.n2965 585
R9546 gnd.n2835 gnd.n2834 585
R9547 gnd.n2834 gnd.n2833 585
R9548 gnd.n2960 gnd.n2959 585
R9549 gnd.n2959 gnd.n2958 585
R9550 gnd.n2838 gnd.n2837 585
R9551 gnd.n2949 gnd.n2838 585
R9552 gnd.n2948 gnd.n2947 585
R9553 gnd.n2950 gnd.n2948 585
R9554 gnd.n2846 gnd.n2845 585
R9555 gnd.n2845 gnd.n2844 585
R9556 gnd.n3687 gnd.n2341 585
R9557 gnd.n2393 gnd.n2341 585
R9558 gnd.n3688 gnd.n2403 585
R9559 gnd.n2403 gnd.n2392 585
R9560 gnd.n3690 gnd.n3689 585
R9561 gnd.n3691 gnd.n3690 585
R9562 gnd.n2404 gnd.n2402 585
R9563 gnd.n2411 gnd.n2402 585
R9564 gnd.n3681 gnd.n3680 585
R9565 gnd.n3680 gnd.n3679 585
R9566 gnd.n2407 gnd.n2406 585
R9567 gnd.n3406 gnd.n2407 585
R9568 gnd.n3392 gnd.n2430 585
R9569 gnd.n2430 gnd.n2420 585
R9570 gnd.n3394 gnd.n3393 585
R9571 gnd.n3395 gnd.n3394 585
R9572 gnd.n2431 gnd.n2429 585
R9573 gnd.n2429 gnd.n2427 585
R9574 gnd.n3387 gnd.n3386 585
R9575 gnd.n3386 gnd.n3385 585
R9576 gnd.n2434 gnd.n2433 585
R9577 gnd.n2443 gnd.n2434 585
R9578 gnd.n3343 gnd.n2457 585
R9579 gnd.n2457 gnd.n2442 585
R9580 gnd.n3345 gnd.n3344 585
R9581 gnd.n3346 gnd.n3345 585
R9582 gnd.n2458 gnd.n2456 585
R9583 gnd.n2465 gnd.n2456 585
R9584 gnd.n3338 gnd.n3337 585
R9585 gnd.n3337 gnd.n3336 585
R9586 gnd.n2461 gnd.n2460 585
R9587 gnd.n3317 gnd.n2461 585
R9588 gnd.n3303 gnd.n2485 585
R9589 gnd.n2485 gnd.n2474 585
R9590 gnd.n3305 gnd.n3304 585
R9591 gnd.n3306 gnd.n3305 585
R9592 gnd.n2486 gnd.n2484 585
R9593 gnd.n2484 gnd.n2481 585
R9594 gnd.n3298 gnd.n3297 585
R9595 gnd.n3297 gnd.n3296 585
R9596 gnd.n2489 gnd.n2488 585
R9597 gnd.n2499 gnd.n2489 585
R9598 gnd.n3258 gnd.n2512 585
R9599 gnd.n2512 gnd.n2498 585
R9600 gnd.n3260 gnd.n3259 585
R9601 gnd.n3261 gnd.n3260 585
R9602 gnd.n2513 gnd.n2511 585
R9603 gnd.n2520 gnd.n2511 585
R9604 gnd.n3253 gnd.n3252 585
R9605 gnd.n3252 gnd.n3251 585
R9606 gnd.n2516 gnd.n2515 585
R9607 gnd.n3232 gnd.n2516 585
R9608 gnd.n3218 gnd.n2539 585
R9609 gnd.n2539 gnd.n2529 585
R9610 gnd.n3220 gnd.n3219 585
R9611 gnd.n3221 gnd.n3220 585
R9612 gnd.n2540 gnd.n2538 585
R9613 gnd.n3209 gnd.n2538 585
R9614 gnd.n3213 gnd.n3212 585
R9615 gnd.n3212 gnd.n3211 585
R9616 gnd.n2543 gnd.n2542 585
R9617 gnd.n3164 gnd.n2543 585
R9618 gnd.n2657 gnd.n2656 585
R9619 gnd.n2658 gnd.n2657 585
R9620 gnd.n2637 gnd.n2636 585
R9621 gnd.n2640 gnd.n2637 585
R9622 gnd.n3174 gnd.n3173 585
R9623 gnd.n3173 gnd.n3172 585
R9624 gnd.n3175 gnd.n2631 585
R9625 gnd.n2667 gnd.n2631 585
R9626 gnd.n3177 gnd.n3176 585
R9627 gnd.n3178 gnd.n3177 585
R9628 gnd.n2632 gnd.n2630 585
R9629 gnd.n3142 gnd.n2630 585
R9630 gnd.n3126 gnd.n3125 585
R9631 gnd.n3125 gnd.n2618 585
R9632 gnd.n3127 gnd.n2682 585
R9633 gnd.n2682 gnd.n2617 585
R9634 gnd.n3129 gnd.n3128 585
R9635 gnd.n3130 gnd.n3129 585
R9636 gnd.n2683 gnd.n2681 585
R9637 gnd.n2681 gnd.n2678 585
R9638 gnd.n3118 gnd.n3117 585
R9639 gnd.n3117 gnd.n3116 585
R9640 gnd.n2686 gnd.n2685 585
R9641 gnd.n2693 gnd.n2686 585
R9642 gnd.n3092 gnd.n3091 585
R9643 gnd.n3093 gnd.n3092 585
R9644 gnd.n2705 gnd.n2704 585
R9645 gnd.n2712 gnd.n2704 585
R9646 gnd.n3087 gnd.n3086 585
R9647 gnd.n3086 gnd.n3085 585
R9648 gnd.n2708 gnd.n2707 585
R9649 gnd.n3075 gnd.n2708 585
R9650 gnd.n3062 gnd.n2732 585
R9651 gnd.n2732 gnd.n2731 585
R9652 gnd.n3064 gnd.n3063 585
R9653 gnd.n3065 gnd.n3064 585
R9654 gnd.n2733 gnd.n2730 585
R9655 gnd.n2740 gnd.n2730 585
R9656 gnd.n3057 gnd.n3056 585
R9657 gnd.n3056 gnd.n3055 585
R9658 gnd.n2736 gnd.n2735 585
R9659 gnd.n3044 gnd.n2736 585
R9660 gnd.n3031 gnd.n2757 585
R9661 gnd.n2757 gnd.n2756 585
R9662 gnd.n3033 gnd.n3032 585
R9663 gnd.n3034 gnd.n3033 585
R9664 gnd.n3027 gnd.n2755 585
R9665 gnd.n3026 gnd.n3025 585
R9666 gnd.n2760 gnd.n2759 585
R9667 gnd.n3023 gnd.n2760 585
R9668 gnd.n2782 gnd.n2781 585
R9669 gnd.n2785 gnd.n2784 585
R9670 gnd.n2783 gnd.n2778 585
R9671 gnd.n2790 gnd.n2789 585
R9672 gnd.n2792 gnd.n2791 585
R9673 gnd.n2795 gnd.n2794 585
R9674 gnd.n2793 gnd.n2776 585
R9675 gnd.n2800 gnd.n2799 585
R9676 gnd.n2802 gnd.n2801 585
R9677 gnd.n2805 gnd.n2804 585
R9678 gnd.n2803 gnd.n2774 585
R9679 gnd.n2810 gnd.n2809 585
R9680 gnd.n2814 gnd.n2811 585
R9681 gnd.n2815 gnd.n2752 585
R9682 gnd.n3693 gnd.n2356 585
R9683 gnd.n3760 gnd.n3759 585
R9684 gnd.n3762 gnd.n3761 585
R9685 gnd.n3764 gnd.n3763 585
R9686 gnd.n3766 gnd.n3765 585
R9687 gnd.n3768 gnd.n3767 585
R9688 gnd.n3770 gnd.n3769 585
R9689 gnd.n3772 gnd.n3771 585
R9690 gnd.n3774 gnd.n3773 585
R9691 gnd.n3776 gnd.n3775 585
R9692 gnd.n3778 gnd.n3777 585
R9693 gnd.n3780 gnd.n3779 585
R9694 gnd.n3782 gnd.n3781 585
R9695 gnd.n3785 gnd.n3784 585
R9696 gnd.n3783 gnd.n2344 585
R9697 gnd.n3789 gnd.n2342 585
R9698 gnd.n3791 gnd.n3790 585
R9699 gnd.n3792 gnd.n3791 585
R9700 gnd.n3694 gnd.n2398 585
R9701 gnd.n3694 gnd.n2393 585
R9702 gnd.n3696 gnd.n3695 585
R9703 gnd.n3695 gnd.n2392 585
R9704 gnd.n3692 gnd.n2397 585
R9705 gnd.n3692 gnd.n3691 585
R9706 gnd.n3671 gnd.n2399 585
R9707 gnd.n2411 gnd.n2399 585
R9708 gnd.n3670 gnd.n2409 585
R9709 gnd.n3679 gnd.n2409 585
R9710 gnd.n3405 gnd.n2416 585
R9711 gnd.n3406 gnd.n3405 585
R9712 gnd.n3404 gnd.n3403 585
R9713 gnd.n3404 gnd.n2420 585
R9714 gnd.n3402 gnd.n2422 585
R9715 gnd.n3395 gnd.n2422 585
R9716 gnd.n2435 gnd.n2423 585
R9717 gnd.n2435 gnd.n2427 585
R9718 gnd.n3351 gnd.n2436 585
R9719 gnd.n3385 gnd.n2436 585
R9720 gnd.n3350 gnd.n3349 585
R9721 gnd.n3349 gnd.n2443 585
R9722 gnd.n3348 gnd.n2451 585
R9723 gnd.n3348 gnd.n2442 585
R9724 gnd.n3347 gnd.n2453 585
R9725 gnd.n3347 gnd.n3346 585
R9726 gnd.n3326 gnd.n2452 585
R9727 gnd.n2465 gnd.n2452 585
R9728 gnd.n3325 gnd.n2463 585
R9729 gnd.n3336 gnd.n2463 585
R9730 gnd.n3316 gnd.n2470 585
R9731 gnd.n3317 gnd.n3316 585
R9732 gnd.n3315 gnd.n3314 585
R9733 gnd.n3315 gnd.n2474 585
R9734 gnd.n3313 gnd.n2476 585
R9735 gnd.n3306 gnd.n2476 585
R9736 gnd.n2491 gnd.n2477 585
R9737 gnd.n2491 gnd.n2481 585
R9738 gnd.n3266 gnd.n2492 585
R9739 gnd.n3296 gnd.n2492 585
R9740 gnd.n3265 gnd.n3264 585
R9741 gnd.n3264 gnd.n2499 585
R9742 gnd.n3263 gnd.n2506 585
R9743 gnd.n3263 gnd.n2498 585
R9744 gnd.n3262 gnd.n2508 585
R9745 gnd.n3262 gnd.n3261 585
R9746 gnd.n3241 gnd.n2507 585
R9747 gnd.n2520 gnd.n2507 585
R9748 gnd.n3240 gnd.n2518 585
R9749 gnd.n3251 gnd.n2518 585
R9750 gnd.n3231 gnd.n2525 585
R9751 gnd.n3232 gnd.n3231 585
R9752 gnd.n3230 gnd.n3229 585
R9753 gnd.n3230 gnd.n2529 585
R9754 gnd.n3228 gnd.n2531 585
R9755 gnd.n3221 gnd.n2531 585
R9756 gnd.n3208 gnd.n2532 585
R9757 gnd.n3209 gnd.n3208 585
R9758 gnd.n3161 gnd.n2545 585
R9759 gnd.n3211 gnd.n2545 585
R9760 gnd.n3163 gnd.n3162 585
R9761 gnd.n3164 gnd.n3163 585
R9762 gnd.n3156 gnd.n2659 585
R9763 gnd.n2659 gnd.n2658 585
R9764 gnd.n3154 gnd.n3153 585
R9765 gnd.n3153 gnd.n2640 585
R9766 gnd.n3151 gnd.n2638 585
R9767 gnd.n3172 gnd.n2638 585
R9768 gnd.n2669 gnd.n2668 585
R9769 gnd.n2668 gnd.n2667 585
R9770 gnd.n3145 gnd.n2628 585
R9771 gnd.n3178 gnd.n2628 585
R9772 gnd.n3144 gnd.n3143 585
R9773 gnd.n3143 gnd.n3142 585
R9774 gnd.n3140 gnd.n2671 585
R9775 gnd.n3140 gnd.n2618 585
R9776 gnd.n3139 gnd.n3138 585
R9777 gnd.n3139 gnd.n2617 585
R9778 gnd.n2674 gnd.n2673 585
R9779 gnd.n3130 gnd.n2673 585
R9780 gnd.n3098 gnd.n3097 585
R9781 gnd.n3097 gnd.n2678 585
R9782 gnd.n3099 gnd.n2687 585
R9783 gnd.n3116 gnd.n2687 585
R9784 gnd.n3096 gnd.n3095 585
R9785 gnd.n3095 gnd.n2693 585
R9786 gnd.n3094 gnd.n2701 585
R9787 gnd.n3094 gnd.n3093 585
R9788 gnd.n3079 gnd.n2702 585
R9789 gnd.n2712 gnd.n2702 585
R9790 gnd.n3078 gnd.n2710 585
R9791 gnd.n3085 gnd.n2710 585
R9792 gnd.n3077 gnd.n3076 585
R9793 gnd.n3076 gnd.n3075 585
R9794 gnd.n2721 gnd.n2718 585
R9795 gnd.n2731 gnd.n2721 585
R9796 gnd.n3067 gnd.n3066 585
R9797 gnd.n3066 gnd.n3065 585
R9798 gnd.n2727 gnd.n2726 585
R9799 gnd.n2740 gnd.n2727 585
R9800 gnd.n3047 gnd.n2738 585
R9801 gnd.n3055 gnd.n2738 585
R9802 gnd.n3046 gnd.n3045 585
R9803 gnd.n3045 gnd.n3044 585
R9804 gnd.n2747 gnd.n2745 585
R9805 gnd.n2756 gnd.n2747 585
R9806 gnd.n3036 gnd.n3035 585
R9807 gnd.n3035 gnd.n3034 585
R9808 gnd.n6263 gnd.n6262 585
R9809 gnd.n6262 gnd.n6261 585
R9810 gnd.n6264 gnd.n1103 585
R9811 gnd.n4553 gnd.n1103 585
R9812 gnd.n6266 gnd.n6265 585
R9813 gnd.n6267 gnd.n6266 585
R9814 gnd.n1088 gnd.n1087 585
R9815 gnd.n4513 gnd.n1088 585
R9816 gnd.n6275 gnd.n6274 585
R9817 gnd.n6274 gnd.n6273 585
R9818 gnd.n6276 gnd.n1082 585
R9819 gnd.n4504 gnd.n1082 585
R9820 gnd.n6278 gnd.n6277 585
R9821 gnd.n6279 gnd.n6278 585
R9822 gnd.n1067 gnd.n1066 585
R9823 gnd.n4496 gnd.n1067 585
R9824 gnd.n6287 gnd.n6286 585
R9825 gnd.n6286 gnd.n6285 585
R9826 gnd.n6288 gnd.n1061 585
R9827 gnd.n4431 gnd.n1061 585
R9828 gnd.n6290 gnd.n6289 585
R9829 gnd.n6291 gnd.n6290 585
R9830 gnd.n1046 gnd.n1045 585
R9831 gnd.n4419 gnd.n1046 585
R9832 gnd.n6299 gnd.n6298 585
R9833 gnd.n6298 gnd.n6297 585
R9834 gnd.n6300 gnd.n1040 585
R9835 gnd.n4442 gnd.n1040 585
R9836 gnd.n6302 gnd.n6301 585
R9837 gnd.n6303 gnd.n6302 585
R9838 gnd.n1025 gnd.n1024 585
R9839 gnd.n4411 gnd.n1025 585
R9840 gnd.n6311 gnd.n6310 585
R9841 gnd.n6310 gnd.n6309 585
R9842 gnd.n6312 gnd.n1019 585
R9843 gnd.n4378 gnd.n1019 585
R9844 gnd.n6314 gnd.n6313 585
R9845 gnd.n6315 gnd.n6314 585
R9846 gnd.n1004 gnd.n1003 585
R9847 gnd.n4370 gnd.n1004 585
R9848 gnd.n6323 gnd.n6322 585
R9849 gnd.n6322 gnd.n6321 585
R9850 gnd.n6324 gnd.n998 585
R9851 gnd.n4393 gnd.n998 585
R9852 gnd.n6326 gnd.n6325 585
R9853 gnd.n6327 gnd.n6326 585
R9854 gnd.n982 gnd.n981 585
R9855 gnd.n4362 gnd.n982 585
R9856 gnd.n6335 gnd.n6334 585
R9857 gnd.n6334 gnd.n6333 585
R9858 gnd.n6336 gnd.n976 585
R9859 gnd.n4344 gnd.n976 585
R9860 gnd.n6338 gnd.n6337 585
R9861 gnd.n6339 gnd.n6338 585
R9862 gnd.n977 gnd.n975 585
R9863 gnd.n975 gnd.n970 585
R9864 gnd.n4334 gnd.n4333 585
R9865 gnd.n4335 gnd.n4334 585
R9866 gnd.n4331 gnd.n2172 585
R9867 gnd.n2178 gnd.n2172 585
R9868 gnd.n4330 gnd.n4329 585
R9869 gnd.n4329 gnd.n4328 585
R9870 gnd.n4306 gnd.n2174 585
R9871 gnd.n2196 gnd.n2174 585
R9872 gnd.n4308 gnd.n4307 585
R9873 gnd.n4309 gnd.n4308 585
R9874 gnd.n4304 gnd.n2198 585
R9875 gnd.n2198 gnd.n2194 585
R9876 gnd.n4303 gnd.n4302 585
R9877 gnd.n4302 gnd.n4301 585
R9878 gnd.n4289 gnd.n2200 585
R9879 gnd.n2201 gnd.n2200 585
R9880 gnd.n4291 gnd.n4290 585
R9881 gnd.n4292 gnd.n4291 585
R9882 gnd.n4287 gnd.n2213 585
R9883 gnd.n2213 gnd.n2210 585
R9884 gnd.n4286 gnd.n4285 585
R9885 gnd.n4285 gnd.n4284 585
R9886 gnd.n2216 gnd.n2214 585
R9887 gnd.n2227 gnd.n2216 585
R9888 gnd.n4275 gnd.n4274 585
R9889 gnd.n4276 gnd.n4275 585
R9890 gnd.n2229 gnd.n2228 585
R9891 gnd.n2228 gnd.n2224 585
R9892 gnd.n4269 gnd.n4268 585
R9893 gnd.n4268 gnd.n4267 585
R9894 gnd.n2232 gnd.n2231 585
R9895 gnd.n2233 gnd.n2232 585
R9896 gnd.n4258 gnd.n4257 585
R9897 gnd.n4259 gnd.n4258 585
R9898 gnd.n2245 gnd.n2244 585
R9899 gnd.n2244 gnd.n2241 585
R9900 gnd.n4253 gnd.n4252 585
R9901 gnd.n4252 gnd.n4251 585
R9902 gnd.n2248 gnd.n2247 585
R9903 gnd.n2259 gnd.n2248 585
R9904 gnd.n4242 gnd.n4241 585
R9905 gnd.n4243 gnd.n4242 585
R9906 gnd.n2261 gnd.n2260 585
R9907 gnd.n2260 gnd.n2256 585
R9908 gnd.n4237 gnd.n4236 585
R9909 gnd.n4236 gnd.n4235 585
R9910 gnd.n2264 gnd.n2263 585
R9911 gnd.n2265 gnd.n2264 585
R9912 gnd.n4226 gnd.n4225 585
R9913 gnd.n4227 gnd.n4226 585
R9914 gnd.n2277 gnd.n2276 585
R9915 gnd.n2276 gnd.n2273 585
R9916 gnd.n4221 gnd.n4220 585
R9917 gnd.n4220 gnd.n4219 585
R9918 gnd.n2280 gnd.n2279 585
R9919 gnd.n2291 gnd.n2280 585
R9920 gnd.n4210 gnd.n4209 585
R9921 gnd.n4211 gnd.n4210 585
R9922 gnd.n2293 gnd.n2292 585
R9923 gnd.n2292 gnd.n2288 585
R9924 gnd.n4205 gnd.n4204 585
R9925 gnd.n4204 gnd.n4203 585
R9926 gnd.n2296 gnd.n2295 585
R9927 gnd.n2297 gnd.n2296 585
R9928 gnd.n4194 gnd.n4193 585
R9929 gnd.n4195 gnd.n4194 585
R9930 gnd.n2309 gnd.n2308 585
R9931 gnd.n2308 gnd.n2305 585
R9932 gnd.n4189 gnd.n4188 585
R9933 gnd.n4188 gnd.n4187 585
R9934 gnd.n2312 gnd.n2311 585
R9935 gnd.n3957 gnd.n2312 585
R9936 gnd.n4178 gnd.n4177 585
R9937 gnd.n4179 gnd.n4178 585
R9938 gnd.n4174 gnd.n3958 585
R9939 gnd.n4173 gnd.n4172 585
R9940 gnd.n4170 gnd.n3960 585
R9941 gnd.n4170 gnd.n3793 585
R9942 gnd.n4169 gnd.n4168 585
R9943 gnd.n4167 gnd.n4166 585
R9944 gnd.n4165 gnd.n3965 585
R9945 gnd.n4163 gnd.n4162 585
R9946 gnd.n4161 gnd.n3966 585
R9947 gnd.n4160 gnd.n4159 585
R9948 gnd.n4157 gnd.n3971 585
R9949 gnd.n4155 gnd.n4154 585
R9950 gnd.n4153 gnd.n3972 585
R9951 gnd.n4152 gnd.n4151 585
R9952 gnd.n4149 gnd.n3977 585
R9953 gnd.n4147 gnd.n4146 585
R9954 gnd.n4145 gnd.n3978 585
R9955 gnd.n4144 gnd.n4143 585
R9956 gnd.n4141 gnd.n3983 585
R9957 gnd.n4139 gnd.n4138 585
R9958 gnd.n4137 gnd.n3984 585
R9959 gnd.n4136 gnd.n4135 585
R9960 gnd.n4133 gnd.n3992 585
R9961 gnd.n4131 gnd.n4130 585
R9962 gnd.n4129 gnd.n3993 585
R9963 gnd.n4128 gnd.n4127 585
R9964 gnd.n4125 gnd.n3998 585
R9965 gnd.n4123 gnd.n4122 585
R9966 gnd.n4121 gnd.n3999 585
R9967 gnd.n4120 gnd.n4119 585
R9968 gnd.n4117 gnd.n4004 585
R9969 gnd.n4115 gnd.n4114 585
R9970 gnd.n4113 gnd.n4005 585
R9971 gnd.n4112 gnd.n4111 585
R9972 gnd.n4109 gnd.n4010 585
R9973 gnd.n4107 gnd.n4106 585
R9974 gnd.n4105 gnd.n4011 585
R9975 gnd.n4104 gnd.n4016 585
R9976 gnd.n4097 gnd.n4019 585
R9977 gnd.n4100 gnd.n4099 585
R9978 gnd.n2104 gnd.n2103 585
R9979 gnd.n4561 gnd.n4560 585
R9980 gnd.n4563 gnd.n4562 585
R9981 gnd.n4565 gnd.n4564 585
R9982 gnd.n4567 gnd.n4566 585
R9983 gnd.n4569 gnd.n4568 585
R9984 gnd.n4571 gnd.n4570 585
R9985 gnd.n4573 gnd.n4572 585
R9986 gnd.n4575 gnd.n4574 585
R9987 gnd.n4577 gnd.n4576 585
R9988 gnd.n4579 gnd.n4578 585
R9989 gnd.n4581 gnd.n4580 585
R9990 gnd.n4583 gnd.n4582 585
R9991 gnd.n4585 gnd.n4584 585
R9992 gnd.n4587 gnd.n4586 585
R9993 gnd.n4589 gnd.n4588 585
R9994 gnd.n4591 gnd.n4590 585
R9995 gnd.n4593 gnd.n4592 585
R9996 gnd.n4595 gnd.n4594 585
R9997 gnd.n4598 gnd.n4597 585
R9998 gnd.n4596 gnd.n2082 585
R9999 gnd.n5327 gnd.n5326 585
R10000 gnd.n5329 gnd.n5328 585
R10001 gnd.n5331 gnd.n5330 585
R10002 gnd.n5333 gnd.n5332 585
R10003 gnd.n5335 gnd.n5334 585
R10004 gnd.n5337 gnd.n5336 585
R10005 gnd.n5339 gnd.n5338 585
R10006 gnd.n5341 gnd.n5340 585
R10007 gnd.n5343 gnd.n5342 585
R10008 gnd.n5345 gnd.n5344 585
R10009 gnd.n5347 gnd.n5346 585
R10010 gnd.n5349 gnd.n5348 585
R10011 gnd.n5350 gnd.n2063 585
R10012 gnd.n5352 gnd.n5351 585
R10013 gnd.n2064 gnd.n2062 585
R10014 gnd.n2065 gnd.n1108 585
R10015 gnd.n5354 gnd.n1108 585
R10016 gnd.n4556 gnd.n1110 585
R10017 gnd.n6261 gnd.n1110 585
R10018 gnd.n4555 gnd.n4554 585
R10019 gnd.n4554 gnd.n4553 585
R10020 gnd.n2108 gnd.n1101 585
R10021 gnd.n6267 gnd.n1101 585
R10022 gnd.n4512 gnd.n4511 585
R10023 gnd.n4513 gnd.n4512 585
R10024 gnd.n2114 gnd.n1090 585
R10025 gnd.n6273 gnd.n1090 585
R10026 gnd.n4506 gnd.n4505 585
R10027 gnd.n4505 gnd.n4504 585
R10028 gnd.n2116 gnd.n1079 585
R10029 gnd.n6279 gnd.n1079 585
R10030 gnd.n4427 gnd.n2120 585
R10031 gnd.n4496 gnd.n2120 585
R10032 gnd.n4428 gnd.n1069 585
R10033 gnd.n6285 gnd.n1069 585
R10034 gnd.n4430 gnd.n4429 585
R10035 gnd.n4431 gnd.n4430 585
R10036 gnd.n2137 gnd.n1058 585
R10037 gnd.n6291 gnd.n1058 585
R10038 gnd.n4421 gnd.n4420 585
R10039 gnd.n4420 gnd.n4419 585
R10040 gnd.n4418 gnd.n1047 585
R10041 gnd.n6297 gnd.n1047 585
R10042 gnd.n4417 gnd.n2131 585
R10043 gnd.n4442 gnd.n2131 585
R10044 gnd.n2139 gnd.n1037 585
R10045 gnd.n6303 gnd.n1037 585
R10046 gnd.n4413 gnd.n4412 585
R10047 gnd.n4412 gnd.n4411 585
R10048 gnd.n2141 gnd.n1027 585
R10049 gnd.n6309 gnd.n1027 585
R10050 gnd.n4377 gnd.n4376 585
R10051 gnd.n4378 gnd.n4377 585
R10052 gnd.n2158 gnd.n1016 585
R10053 gnd.n6315 gnd.n1016 585
R10054 gnd.n4372 gnd.n4371 585
R10055 gnd.n4371 gnd.n4370 585
R10056 gnd.n4369 gnd.n1005 585
R10057 gnd.n6321 gnd.n1005 585
R10058 gnd.n4368 gnd.n2152 585
R10059 gnd.n4393 gnd.n2152 585
R10060 gnd.n2160 gnd.n995 585
R10061 gnd.n6327 gnd.n995 585
R10062 gnd.n4364 gnd.n4363 585
R10063 gnd.n4363 gnd.n4362 585
R10064 gnd.n2162 gnd.n984 585
R10065 gnd.n6333 gnd.n984 585
R10066 gnd.n4343 gnd.n4342 585
R10067 gnd.n4344 gnd.n4343 585
R10068 gnd.n2166 gnd.n971 585
R10069 gnd.n6339 gnd.n971 585
R10070 gnd.n4338 gnd.n4337 585
R10071 gnd.n4337 gnd.n970 585
R10072 gnd.n4336 gnd.n2168 585
R10073 gnd.n4336 gnd.n4335 585
R10074 gnd.n2189 gnd.n2169 585
R10075 gnd.n2178 gnd.n2169 585
R10076 gnd.n2190 gnd.n2175 585
R10077 gnd.n4328 gnd.n2175 585
R10078 gnd.n2193 gnd.n2191 585
R10079 gnd.n2196 gnd.n2193 585
R10080 gnd.n4311 gnd.n4310 585
R10081 gnd.n4310 gnd.n4309 585
R10082 gnd.n2192 gnd.n2186 585
R10083 gnd.n2194 gnd.n2192 585
R10084 gnd.n4051 gnd.n2202 585
R10085 gnd.n4301 gnd.n2202 585
R10086 gnd.n4053 gnd.n4052 585
R10087 gnd.n4052 gnd.n2201 585
R10088 gnd.n4054 gnd.n2211 585
R10089 gnd.n4292 gnd.n2211 585
R10090 gnd.n4056 gnd.n4055 585
R10091 gnd.n4055 gnd.n2210 585
R10092 gnd.n4057 gnd.n2217 585
R10093 gnd.n4284 gnd.n2217 585
R10094 gnd.n4059 gnd.n4058 585
R10095 gnd.n4058 gnd.n2227 585
R10096 gnd.n4060 gnd.n2225 585
R10097 gnd.n4276 gnd.n2225 585
R10098 gnd.n4062 gnd.n4061 585
R10099 gnd.n4061 gnd.n2224 585
R10100 gnd.n4063 gnd.n2234 585
R10101 gnd.n4267 gnd.n2234 585
R10102 gnd.n4065 gnd.n4064 585
R10103 gnd.n4064 gnd.n2233 585
R10104 gnd.n4066 gnd.n2242 585
R10105 gnd.n4259 gnd.n2242 585
R10106 gnd.n4068 gnd.n4067 585
R10107 gnd.n4067 gnd.n2241 585
R10108 gnd.n4069 gnd.n2249 585
R10109 gnd.n4251 gnd.n2249 585
R10110 gnd.n4071 gnd.n4070 585
R10111 gnd.n4070 gnd.n2259 585
R10112 gnd.n4072 gnd.n2257 585
R10113 gnd.n4243 gnd.n2257 585
R10114 gnd.n4074 gnd.n4073 585
R10115 gnd.n4073 gnd.n2256 585
R10116 gnd.n4075 gnd.n2266 585
R10117 gnd.n4235 gnd.n2266 585
R10118 gnd.n4077 gnd.n4076 585
R10119 gnd.n4076 gnd.n2265 585
R10120 gnd.n4078 gnd.n2274 585
R10121 gnd.n4227 gnd.n2274 585
R10122 gnd.n4080 gnd.n4079 585
R10123 gnd.n4079 gnd.n2273 585
R10124 gnd.n4081 gnd.n2281 585
R10125 gnd.n4219 gnd.n2281 585
R10126 gnd.n4083 gnd.n4082 585
R10127 gnd.n4082 gnd.n2291 585
R10128 gnd.n4084 gnd.n2289 585
R10129 gnd.n4211 gnd.n2289 585
R10130 gnd.n4086 gnd.n4085 585
R10131 gnd.n4085 gnd.n2288 585
R10132 gnd.n4087 gnd.n2298 585
R10133 gnd.n4203 gnd.n2298 585
R10134 gnd.n4089 gnd.n4088 585
R10135 gnd.n4088 gnd.n2297 585
R10136 gnd.n4090 gnd.n2306 585
R10137 gnd.n4195 gnd.n2306 585
R10138 gnd.n4092 gnd.n4091 585
R10139 gnd.n4091 gnd.n2305 585
R10140 gnd.n4093 gnd.n2313 585
R10141 gnd.n4187 gnd.n2313 585
R10142 gnd.n4094 gnd.n4021 585
R10143 gnd.n4021 gnd.n3957 585
R10144 gnd.n4095 gnd.n3794 585
R10145 gnd.n4179 gnd.n3794 585
R10146 gnd.n7601 gnd.n7600 585
R10147 gnd.n7602 gnd.n7601 585
R10148 gnd.n132 gnd.n130 585
R10149 gnd.n130 gnd.n126 585
R10150 gnd.n7521 gnd.n7520 585
R10151 gnd.n7522 gnd.n7521 585
R10152 gnd.n209 gnd.n208 585
R10153 gnd.n208 gnd.n206 585
R10154 gnd.n7516 gnd.n7515 585
R10155 gnd.n7515 gnd.n7514 585
R10156 gnd.n212 gnd.n211 585
R10157 gnd.n213 gnd.n212 585
R10158 gnd.n7437 gnd.n7436 585
R10159 gnd.n7438 gnd.n7437 585
R10160 gnd.n225 gnd.n224 585
R10161 gnd.n232 gnd.n224 585
R10162 gnd.n7432 gnd.n7431 585
R10163 gnd.n7431 gnd.n7430 585
R10164 gnd.n228 gnd.n227 585
R10165 gnd.n229 gnd.n228 585
R10166 gnd.n7421 gnd.n7420 585
R10167 gnd.n7422 gnd.n7421 585
R10168 gnd.n241 gnd.n240 585
R10169 gnd.n247 gnd.n240 585
R10170 gnd.n7416 gnd.n7415 585
R10171 gnd.n7415 gnd.n7414 585
R10172 gnd.n244 gnd.n243 585
R10173 gnd.n254 gnd.n244 585
R10174 gnd.n7405 gnd.n7404 585
R10175 gnd.n7406 gnd.n7405 585
R10176 gnd.n256 gnd.n255 585
R10177 gnd.n263 gnd.n255 585
R10178 gnd.n7400 gnd.n7399 585
R10179 gnd.n7399 gnd.n7398 585
R10180 gnd.n259 gnd.n258 585
R10181 gnd.n260 gnd.n259 585
R10182 gnd.n7389 gnd.n7388 585
R10183 gnd.n7390 gnd.n7389 585
R10184 gnd.n272 gnd.n271 585
R10185 gnd.n271 gnd.n269 585
R10186 gnd.n7384 gnd.n7383 585
R10187 gnd.n7383 gnd.n7382 585
R10188 gnd.n275 gnd.n274 585
R10189 gnd.n284 gnd.n275 585
R10190 gnd.n7373 gnd.n7372 585
R10191 gnd.n7374 gnd.n7373 585
R10192 gnd.n286 gnd.n285 585
R10193 gnd.n293 gnd.n285 585
R10194 gnd.n7368 gnd.n7367 585
R10195 gnd.n7367 gnd.n7366 585
R10196 gnd.n289 gnd.n288 585
R10197 gnd.n290 gnd.n289 585
R10198 gnd.n7357 gnd.n7356 585
R10199 gnd.n7358 gnd.n7357 585
R10200 gnd.n302 gnd.n301 585
R10201 gnd.n301 gnd.n299 585
R10202 gnd.n7333 gnd.n7332 585
R10203 gnd.n7334 gnd.n7333 585
R10204 gnd.n7331 gnd.n332 585
R10205 gnd.n7331 gnd.n7330 585
R10206 gnd.n331 gnd.n330 585
R10207 gnd.n334 gnd.n330 585
R10208 gnd.n7256 gnd.n7255 585
R10209 gnd.n7257 gnd.n7256 585
R10210 gnd.n7254 gnd.n7253 585
R10211 gnd.n7253 gnd.n340 585
R10212 gnd.n7252 gnd.n342 585
R10213 gnd.n7252 gnd.n7251 585
R10214 gnd.n341 gnd.n311 585
R10215 gnd.n315 gnd.n311 585
R10216 gnd.n7351 gnd.n7350 585
R10217 gnd.n7350 gnd.n7349 585
R10218 gnd.n7352 gnd.n310 585
R10219 gnd.n7242 gnd.n310 585
R10220 gnd.n361 gnd.n309 585
R10221 gnd.n361 gnd.n350 585
R10222 gnd.n7226 gnd.n7225 585
R10223 gnd.n7227 gnd.n7226 585
R10224 gnd.n7224 gnd.n360 585
R10225 gnd.n7206 gnd.n360 585
R10226 gnd.n366 gnd.n362 585
R10227 gnd.n7190 gnd.n366 585
R10228 gnd.n7220 gnd.n7219 585
R10229 gnd.n7219 gnd.n7218 585
R10230 gnd.n365 gnd.n364 585
R10231 gnd.n7196 gnd.n365 585
R10232 gnd.n7179 gnd.n394 585
R10233 gnd.n7163 gnd.n394 585
R10234 gnd.n7181 gnd.n7180 585
R10235 gnd.n7182 gnd.n7181 585
R10236 gnd.n395 gnd.n393 585
R10237 gnd.n5941 gnd.n393 585
R10238 gnd.n7174 gnd.n7173 585
R10239 gnd.n7173 gnd.n7172 585
R10240 gnd.n398 gnd.n397 585
R10241 gnd.n5936 gnd.n398 585
R10242 gnd.n5986 gnd.n5985 585
R10243 gnd.n5987 gnd.n5986 585
R10244 gnd.n1366 gnd.n1365 585
R10245 gnd.n1373 gnd.n1365 585
R10246 gnd.n5981 gnd.n5980 585
R10247 gnd.n5980 gnd.n5979 585
R10248 gnd.n1369 gnd.n1368 585
R10249 gnd.n5957 gnd.n1369 585
R10250 gnd.n5916 gnd.n1399 585
R10251 gnd.n1399 gnd.n1398 585
R10252 gnd.n5918 gnd.n5917 585
R10253 gnd.n5919 gnd.n5918 585
R10254 gnd.n1400 gnd.n1397 585
R10255 gnd.n1407 gnd.n1397 585
R10256 gnd.n5911 gnd.n5910 585
R10257 gnd.n5910 gnd.n5909 585
R10258 gnd.n1403 gnd.n1402 585
R10259 gnd.n5896 gnd.n1403 585
R10260 gnd.n5879 gnd.n1426 585
R10261 gnd.n1426 gnd.n1414 585
R10262 gnd.n5881 gnd.n5880 585
R10263 gnd.n5882 gnd.n5881 585
R10264 gnd.n1427 gnd.n1425 585
R10265 gnd.n1435 gnd.n1425 585
R10266 gnd.n5874 gnd.n5873 585
R10267 gnd.n5873 gnd.n5872 585
R10268 gnd.n1430 gnd.n1429 585
R10269 gnd.n5860 gnd.n1430 585
R10270 gnd.n5848 gnd.n5843 585
R10271 gnd.n5843 gnd.n1452 585
R10272 gnd.n5850 gnd.n5849 585
R10273 gnd.n5851 gnd.n5850 585
R10274 gnd.n5844 gnd.n1288 585
R10275 gnd.n6016 gnd.n1288 585
R10276 gnd.n6090 gnd.n6089 585
R10277 gnd.n6088 gnd.n1287 585
R10278 gnd.n6087 gnd.n1286 585
R10279 gnd.n6092 gnd.n1286 585
R10280 gnd.n6086 gnd.n6085 585
R10281 gnd.n6084 gnd.n6083 585
R10282 gnd.n6082 gnd.n6081 585
R10283 gnd.n6080 gnd.n6079 585
R10284 gnd.n6078 gnd.n6077 585
R10285 gnd.n6076 gnd.n6075 585
R10286 gnd.n6074 gnd.n6073 585
R10287 gnd.n6072 gnd.n6071 585
R10288 gnd.n6070 gnd.n6069 585
R10289 gnd.n6068 gnd.n6067 585
R10290 gnd.n6066 gnd.n6065 585
R10291 gnd.n6064 gnd.n6063 585
R10292 gnd.n6062 gnd.n6061 585
R10293 gnd.n6059 gnd.n6058 585
R10294 gnd.n6057 gnd.n6056 585
R10295 gnd.n6055 gnd.n6054 585
R10296 gnd.n6053 gnd.n6052 585
R10297 gnd.n6051 gnd.n6050 585
R10298 gnd.n6049 gnd.n6048 585
R10299 gnd.n6047 gnd.n6046 585
R10300 gnd.n6045 gnd.n6044 585
R10301 gnd.n6043 gnd.n6042 585
R10302 gnd.n6041 gnd.n6040 585
R10303 gnd.n6039 gnd.n6038 585
R10304 gnd.n6037 gnd.n6036 585
R10305 gnd.n6035 gnd.n6034 585
R10306 gnd.n6033 gnd.n6032 585
R10307 gnd.n6031 gnd.n6030 585
R10308 gnd.n6029 gnd.n6028 585
R10309 gnd.n6027 gnd.n6026 585
R10310 gnd.n6025 gnd.n6024 585
R10311 gnd.n6023 gnd.n1328 585
R10312 gnd.n1332 gnd.n1329 585
R10313 gnd.n6019 gnd.n6018 585
R10314 gnd.n200 gnd.n199 585
R10315 gnd.n7530 gnd.n195 585
R10316 gnd.n7532 gnd.n7531 585
R10317 gnd.n7534 gnd.n193 585
R10318 gnd.n7536 gnd.n7535 585
R10319 gnd.n7537 gnd.n188 585
R10320 gnd.n7539 gnd.n7538 585
R10321 gnd.n7541 gnd.n186 585
R10322 gnd.n7543 gnd.n7542 585
R10323 gnd.n7544 gnd.n181 585
R10324 gnd.n7546 gnd.n7545 585
R10325 gnd.n7548 gnd.n179 585
R10326 gnd.n7550 gnd.n7549 585
R10327 gnd.n7551 gnd.n174 585
R10328 gnd.n7553 gnd.n7552 585
R10329 gnd.n7555 gnd.n172 585
R10330 gnd.n7557 gnd.n7556 585
R10331 gnd.n7558 gnd.n167 585
R10332 gnd.n7560 gnd.n7559 585
R10333 gnd.n7562 gnd.n165 585
R10334 gnd.n7564 gnd.n7563 585
R10335 gnd.n7568 gnd.n160 585
R10336 gnd.n7570 gnd.n7569 585
R10337 gnd.n7572 gnd.n158 585
R10338 gnd.n7574 gnd.n7573 585
R10339 gnd.n7575 gnd.n153 585
R10340 gnd.n7577 gnd.n7576 585
R10341 gnd.n7579 gnd.n151 585
R10342 gnd.n7581 gnd.n7580 585
R10343 gnd.n7582 gnd.n146 585
R10344 gnd.n7584 gnd.n7583 585
R10345 gnd.n7586 gnd.n144 585
R10346 gnd.n7588 gnd.n7587 585
R10347 gnd.n7589 gnd.n139 585
R10348 gnd.n7591 gnd.n7590 585
R10349 gnd.n7593 gnd.n137 585
R10350 gnd.n7595 gnd.n7594 585
R10351 gnd.n7596 gnd.n135 585
R10352 gnd.n7597 gnd.n131 585
R10353 gnd.n131 gnd.n128 585
R10354 gnd.n7526 gnd.n127 585
R10355 gnd.n7602 gnd.n127 585
R10356 gnd.n7525 gnd.n7524 585
R10357 gnd.n7524 gnd.n126 585
R10358 gnd.n7523 gnd.n204 585
R10359 gnd.n7523 gnd.n7522 585
R10360 gnd.n7290 gnd.n205 585
R10361 gnd.n206 gnd.n205 585
R10362 gnd.n7291 gnd.n214 585
R10363 gnd.n7514 gnd.n214 585
R10364 gnd.n7293 gnd.n7292 585
R10365 gnd.n7292 gnd.n213 585
R10366 gnd.n7294 gnd.n223 585
R10367 gnd.n7438 gnd.n223 585
R10368 gnd.n7296 gnd.n7295 585
R10369 gnd.n7295 gnd.n232 585
R10370 gnd.n7297 gnd.n230 585
R10371 gnd.n7430 gnd.n230 585
R10372 gnd.n7299 gnd.n7298 585
R10373 gnd.n7298 gnd.n229 585
R10374 gnd.n7300 gnd.n239 585
R10375 gnd.n7422 gnd.n239 585
R10376 gnd.n7302 gnd.n7301 585
R10377 gnd.n7301 gnd.n247 585
R10378 gnd.n7303 gnd.n245 585
R10379 gnd.n7414 gnd.n245 585
R10380 gnd.n7305 gnd.n7304 585
R10381 gnd.n7304 gnd.n254 585
R10382 gnd.n7306 gnd.n253 585
R10383 gnd.n7406 gnd.n253 585
R10384 gnd.n7308 gnd.n7307 585
R10385 gnd.n7307 gnd.n263 585
R10386 gnd.n7309 gnd.n261 585
R10387 gnd.n7398 gnd.n261 585
R10388 gnd.n7311 gnd.n7310 585
R10389 gnd.n7310 gnd.n260 585
R10390 gnd.n7312 gnd.n270 585
R10391 gnd.n7390 gnd.n270 585
R10392 gnd.n7314 gnd.n7313 585
R10393 gnd.n7313 gnd.n269 585
R10394 gnd.n7315 gnd.n276 585
R10395 gnd.n7382 gnd.n276 585
R10396 gnd.n7317 gnd.n7316 585
R10397 gnd.n7316 gnd.n284 585
R10398 gnd.n7318 gnd.n283 585
R10399 gnd.n7374 gnd.n283 585
R10400 gnd.n7320 gnd.n7319 585
R10401 gnd.n7319 gnd.n293 585
R10402 gnd.n7321 gnd.n291 585
R10403 gnd.n7366 gnd.n291 585
R10404 gnd.n7323 gnd.n7322 585
R10405 gnd.n7322 gnd.n290 585
R10406 gnd.n7324 gnd.n300 585
R10407 gnd.n7358 gnd.n300 585
R10408 gnd.n7326 gnd.n7325 585
R10409 gnd.n7325 gnd.n299 585
R10410 gnd.n7327 gnd.n328 585
R10411 gnd.n7334 gnd.n328 585
R10412 gnd.n7329 gnd.n7328 585
R10413 gnd.n7330 gnd.n7329 585
R10414 gnd.n336 gnd.n335 585
R10415 gnd.n335 gnd.n334 585
R10416 gnd.n7259 gnd.n7258 585
R10417 gnd.n7258 gnd.n7257 585
R10418 gnd.n339 gnd.n338 585
R10419 gnd.n340 gnd.n339 585
R10420 gnd.n7236 gnd.n343 585
R10421 gnd.n7251 gnd.n343 585
R10422 gnd.n7238 gnd.n7237 585
R10423 gnd.n7237 gnd.n315 585
R10424 gnd.n7239 gnd.n313 585
R10425 gnd.n7349 gnd.n313 585
R10426 gnd.n7241 gnd.n7240 585
R10427 gnd.n7242 gnd.n7241 585
R10428 gnd.n352 gnd.n351 585
R10429 gnd.n351 gnd.n350 585
R10430 gnd.n7229 gnd.n7228 585
R10431 gnd.n7228 gnd.n7227 585
R10432 gnd.n355 gnd.n354 585
R10433 gnd.n7206 gnd.n355 585
R10434 gnd.n7192 gnd.n7191 585
R10435 gnd.n7191 gnd.n7190 585
R10436 gnd.n7193 gnd.n368 585
R10437 gnd.n7218 gnd.n368 585
R10438 gnd.n7195 gnd.n7194 585
R10439 gnd.n7196 gnd.n7195 585
R10440 gnd.n386 gnd.n385 585
R10441 gnd.n7163 gnd.n385 585
R10442 gnd.n7184 gnd.n7183 585
R10443 gnd.n7183 gnd.n7182 585
R10444 gnd.n389 gnd.n388 585
R10445 gnd.n5941 gnd.n389 585
R10446 gnd.n5933 gnd.n400 585
R10447 gnd.n7172 gnd.n400 585
R10448 gnd.n5935 gnd.n5934 585
R10449 gnd.n5936 gnd.n5935 585
R10450 gnd.n1387 gnd.n1362 585
R10451 gnd.n5987 gnd.n1362 585
R10452 gnd.n5928 gnd.n5927 585
R10453 gnd.n5927 gnd.n1373 585
R10454 gnd.n5926 gnd.n1371 585
R10455 gnd.n5979 gnd.n1371 585
R10456 gnd.n5925 gnd.n1380 585
R10457 gnd.n5957 gnd.n1380 585
R10458 gnd.n1393 gnd.n1389 585
R10459 gnd.n1398 gnd.n1393 585
R10460 gnd.n5921 gnd.n5920 585
R10461 gnd.n5920 gnd.n5919 585
R10462 gnd.n1392 gnd.n1391 585
R10463 gnd.n1407 gnd.n1392 585
R10464 gnd.n1465 gnd.n1405 585
R10465 gnd.n5909 gnd.n1405 585
R10466 gnd.n1466 gnd.n1415 585
R10467 gnd.n5896 gnd.n1415 585
R10468 gnd.n1468 gnd.n1467 585
R10469 gnd.n1467 gnd.n1414 585
R10470 gnd.n1469 gnd.n1423 585
R10471 gnd.n5882 gnd.n1423 585
R10472 gnd.n1471 gnd.n1470 585
R10473 gnd.n1470 gnd.n1435 585
R10474 gnd.n1472 gnd.n1432 585
R10475 gnd.n5872 gnd.n1432 585
R10476 gnd.n1474 gnd.n1473 585
R10477 gnd.n5860 gnd.n1474 585
R10478 gnd.n1454 gnd.n1453 585
R10479 gnd.n1453 gnd.n1452 585
R10480 gnd.n1455 gnd.n1334 585
R10481 gnd.n5851 gnd.n1334 585
R10482 gnd.n6017 gnd.n1335 585
R10483 gnd.n6017 gnd.n6016 585
R10484 gnd.n4948 gnd.n4923 585
R10485 gnd.n4923 gnd.n1698 585
R10486 gnd.n4947 gnd.n4946 585
R10487 gnd.n4946 gnd.n1707 585
R10488 gnd.n4945 gnd.n4944 585
R10489 gnd.n4945 gnd.n1706 585
R10490 gnd.n4943 gnd.n4882 585
R10491 gnd.n5092 gnd.n4882 585
R10492 gnd.n5095 gnd.n4881 585
R10493 gnd.n5095 gnd.n5094 585
R10494 gnd.n5097 gnd.n5096 585
R10495 gnd.n5096 gnd.n1713 585
R10496 gnd.n5098 gnd.n4879 585
R10497 gnd.n4879 gnd.n4878 585
R10498 gnd.n5100 gnd.n5099 585
R10499 gnd.n5101 gnd.n5100 585
R10500 gnd.n4880 gnd.n4877 585
R10501 gnd.n4877 gnd.n1720 585
R10502 gnd.n4869 gnd.n4868 585
R10503 gnd.n5107 gnd.n4869 585
R10504 gnd.n5111 gnd.n5110 585
R10505 gnd.n5110 gnd.n5109 585
R10506 gnd.n5112 gnd.n4865 585
R10507 gnd.n4865 gnd.n1726 585
R10508 gnd.n5114 gnd.n5113 585
R10509 gnd.n5115 gnd.n5114 585
R10510 gnd.n4867 gnd.n4864 585
R10511 gnd.n4864 gnd.n1734 585
R10512 gnd.n4866 gnd.n4856 585
R10513 gnd.n4856 gnd.n1733 585
R10514 gnd.n5123 gnd.n4855 585
R10515 gnd.n5123 gnd.n5122 585
R10516 gnd.n5125 gnd.n5124 585
R10517 gnd.n5124 gnd.n1742 585
R10518 gnd.n5126 gnd.n4854 585
R10519 gnd.n4854 gnd.n1740 585
R10520 gnd.n5128 gnd.n5127 585
R10521 gnd.n5129 gnd.n5128 585
R10522 gnd.n4848 gnd.n4847 585
R10523 gnd.n4848 gnd.n1748 585
R10524 gnd.n5137 gnd.n5136 585
R10525 gnd.n5136 gnd.n5135 585
R10526 gnd.n5138 gnd.n4845 585
R10527 gnd.n4849 gnd.n4845 585
R10528 gnd.n5140 gnd.n5139 585
R10529 gnd.n5141 gnd.n5140 585
R10530 gnd.n4846 gnd.n4837 585
R10531 gnd.n4837 gnd.n1754 585
R10532 gnd.n5149 gnd.n4836 585
R10533 gnd.n5149 gnd.n5148 585
R10534 gnd.n5151 gnd.n5150 585
R10535 gnd.n5150 gnd.n1762 585
R10536 gnd.n5152 gnd.n4833 585
R10537 gnd.n4833 gnd.n1761 585
R10538 gnd.n5154 gnd.n5153 585
R10539 gnd.n5155 gnd.n5154 585
R10540 gnd.n4835 gnd.n4832 585
R10541 gnd.n4832 gnd.n1770 585
R10542 gnd.n4834 gnd.n4824 585
R10543 gnd.n4824 gnd.n1768 585
R10544 gnd.n5164 gnd.n4823 585
R10545 gnd.n5164 gnd.n5163 585
R10546 gnd.n5166 gnd.n5165 585
R10547 gnd.n5165 gnd.n1776 585
R10548 gnd.n5167 gnd.n4820 585
R10549 gnd.n4820 gnd.n4819 585
R10550 gnd.n5169 gnd.n5168 585
R10551 gnd.n5170 gnd.n5169 585
R10552 gnd.n4822 gnd.n4818 585
R10553 gnd.n4818 gnd.n1784 585
R10554 gnd.n4821 gnd.n4811 585
R10555 gnd.n4811 gnd.n1782 585
R10556 gnd.n5179 gnd.n4810 585
R10557 gnd.n5179 gnd.n5178 585
R10558 gnd.n5181 gnd.n5180 585
R10559 gnd.n5180 gnd.n1790 585
R10560 gnd.n5182 gnd.n4807 585
R10561 gnd.n4807 gnd.n4806 585
R10562 gnd.n5184 gnd.n5183 585
R10563 gnd.n5185 gnd.n5184 585
R10564 gnd.n4809 gnd.n4805 585
R10565 gnd.n4805 gnd.n1797 585
R10566 gnd.n4808 gnd.n4783 585
R10567 gnd.n5191 gnd.n4783 585
R10568 gnd.n5194 gnd.n4784 585
R10569 gnd.n5194 gnd.n5193 585
R10570 gnd.n5195 gnd.n4782 585
R10571 gnd.n5195 gnd.n1804 585
R10572 gnd.n5197 gnd.n5196 585
R10573 gnd.n5196 gnd.n1803 585
R10574 gnd.n5198 gnd.n4781 585
R10575 gnd.n4796 gnd.n4781 585
R10576 gnd.n5200 gnd.n5199 585
R10577 gnd.n5200 gnd.n1812 585
R10578 gnd.n5201 gnd.n4780 585
R10579 gnd.n5201 gnd.n1810 585
R10580 gnd.n5203 gnd.n5202 585
R10581 gnd.n5202 gnd.n1820 585
R10582 gnd.n5204 gnd.n4778 585
R10583 gnd.n4778 gnd.n1818 585
R10584 gnd.n5206 gnd.n5205 585
R10585 gnd.n5207 gnd.n5206 585
R10586 gnd.n4779 gnd.n4777 585
R10587 gnd.n4777 gnd.n1827 585
R10588 gnd.n4762 gnd.n4761 585
R10589 gnd.n5213 gnd.n4762 585
R10590 gnd.n5216 gnd.n5215 585
R10591 gnd.n5215 gnd.n5214 585
R10592 gnd.n5217 gnd.n4759 585
R10593 gnd.n4759 gnd.n1833 585
R10594 gnd.n5219 gnd.n5218 585
R10595 gnd.n5220 gnd.n5219 585
R10596 gnd.n4760 gnd.n4755 585
R10597 gnd.n5221 gnd.n4755 585
R10598 gnd.n5224 gnd.n4754 585
R10599 gnd.n5224 gnd.n5223 585
R10600 gnd.n5226 gnd.n5225 585
R10601 gnd.n5225 gnd.n1839 585
R10602 gnd.n5227 gnd.n4752 585
R10603 gnd.n4752 gnd.n4751 585
R10604 gnd.n5229 gnd.n5228 585
R10605 gnd.n5230 gnd.n5229 585
R10606 gnd.n4753 gnd.n4742 585
R10607 gnd.n4742 gnd.n1846 585
R10608 gnd.n5237 gnd.n4741 585
R10609 gnd.n5237 gnd.n5236 585
R10610 gnd.n5239 gnd.n5238 585
R10611 gnd.n5238 gnd.t304 585
R10612 gnd.n5240 gnd.n4738 585
R10613 gnd.n4738 gnd.n1852 585
R10614 gnd.n5242 gnd.n5241 585
R10615 gnd.n5243 gnd.n5242 585
R10616 gnd.n4740 gnd.n4737 585
R10617 gnd.n4737 gnd.n1860 585
R10618 gnd.n4739 gnd.n4662 585
R10619 gnd.n4662 gnd.n1859 585
R10620 gnd.n5251 gnd.n4661 585
R10621 gnd.n5251 gnd.n5250 585
R10622 gnd.n5253 gnd.n5252 585
R10623 gnd.n5252 gnd.n1868 585
R10624 gnd.n5254 gnd.n4640 585
R10625 gnd.n4640 gnd.n1866 585
R10626 gnd.n5319 gnd.n5318 585
R10627 gnd.n5317 gnd.n4639 585
R10628 gnd.n5316 gnd.n4638 585
R10629 gnd.n5321 gnd.n4638 585
R10630 gnd.n5315 gnd.n5314 585
R10631 gnd.n5313 gnd.n5312 585
R10632 gnd.n5311 gnd.n5310 585
R10633 gnd.n5309 gnd.n5308 585
R10634 gnd.n5307 gnd.n5306 585
R10635 gnd.n5305 gnd.n5304 585
R10636 gnd.n5303 gnd.n5302 585
R10637 gnd.n5301 gnd.n5300 585
R10638 gnd.n5299 gnd.n5298 585
R10639 gnd.n5297 gnd.n5296 585
R10640 gnd.n5295 gnd.n5294 585
R10641 gnd.n5293 gnd.n5292 585
R10642 gnd.n5291 gnd.n5290 585
R10643 gnd.n5289 gnd.n5288 585
R10644 gnd.n5287 gnd.n5286 585
R10645 gnd.n5285 gnd.n5284 585
R10646 gnd.n5283 gnd.n5282 585
R10647 gnd.n5281 gnd.n5280 585
R10648 gnd.n5279 gnd.n5278 585
R10649 gnd.n5277 gnd.n5276 585
R10650 gnd.n5275 gnd.n5274 585
R10651 gnd.n5273 gnd.n5272 585
R10652 gnd.n5271 gnd.n5270 585
R10653 gnd.n5269 gnd.n5268 585
R10654 gnd.n5267 gnd.n5266 585
R10655 gnd.n5265 gnd.n5264 585
R10656 gnd.n5263 gnd.n5262 585
R10657 gnd.n5261 gnd.n5260 585
R10658 gnd.n5259 gnd.n4603 585
R10659 gnd.n5324 gnd.n5323 585
R10660 gnd.n4605 gnd.n4602 585
R10661 gnd.n4669 gnd.n4668 585
R10662 gnd.n4671 gnd.n4670 585
R10663 gnd.n4674 gnd.n4673 585
R10664 gnd.n4676 gnd.n4675 585
R10665 gnd.n4678 gnd.n4677 585
R10666 gnd.n4680 gnd.n4679 585
R10667 gnd.n4682 gnd.n4681 585
R10668 gnd.n4684 gnd.n4683 585
R10669 gnd.n4686 gnd.n4685 585
R10670 gnd.n4688 gnd.n4687 585
R10671 gnd.n4690 gnd.n4689 585
R10672 gnd.n4692 gnd.n4691 585
R10673 gnd.n4694 gnd.n4693 585
R10674 gnd.n4696 gnd.n4695 585
R10675 gnd.n4698 gnd.n4697 585
R10676 gnd.n4700 gnd.n4699 585
R10677 gnd.n4702 gnd.n4701 585
R10678 gnd.n4704 gnd.n4703 585
R10679 gnd.n4706 gnd.n4705 585
R10680 gnd.n4708 gnd.n4707 585
R10681 gnd.n4710 gnd.n4709 585
R10682 gnd.n4712 gnd.n4711 585
R10683 gnd.n4714 gnd.n4713 585
R10684 gnd.n4716 gnd.n4715 585
R10685 gnd.n4718 gnd.n4717 585
R10686 gnd.n4720 gnd.n4719 585
R10687 gnd.n4722 gnd.n4721 585
R10688 gnd.n4724 gnd.n4723 585
R10689 gnd.n4726 gnd.n4725 585
R10690 gnd.n4728 gnd.n4727 585
R10691 gnd.n4730 gnd.n4729 585
R10692 gnd.n5085 gnd.n5084 585
R10693 gnd.n5083 gnd.n5082 585
R10694 gnd.n5081 gnd.n4890 585
R10695 gnd.n5079 gnd.n5078 585
R10696 gnd.n5077 gnd.n4891 585
R10697 gnd.n5076 gnd.n5075 585
R10698 gnd.n5073 gnd.n4892 585
R10699 gnd.n5071 gnd.n5070 585
R10700 gnd.n5069 gnd.n4893 585
R10701 gnd.n5068 gnd.n5067 585
R10702 gnd.n5065 gnd.n4894 585
R10703 gnd.n5063 gnd.n5062 585
R10704 gnd.n5061 gnd.n4895 585
R10705 gnd.n5060 gnd.n5059 585
R10706 gnd.n5057 gnd.n4896 585
R10707 gnd.n5055 gnd.n5054 585
R10708 gnd.n5053 gnd.n4897 585
R10709 gnd.n5052 gnd.n5051 585
R10710 gnd.n5049 gnd.n4898 585
R10711 gnd.n5047 gnd.n5046 585
R10712 gnd.n5045 gnd.n4899 585
R10713 gnd.n5044 gnd.n5043 585
R10714 gnd.n5041 gnd.n4900 585
R10715 gnd.n5039 gnd.n5038 585
R10716 gnd.n5037 gnd.n4901 585
R10717 gnd.n5036 gnd.n5035 585
R10718 gnd.n5033 gnd.n4902 585
R10719 gnd.n5031 gnd.n5030 585
R10720 gnd.n5029 gnd.n4903 585
R10721 gnd.n5027 gnd.n5026 585
R10722 gnd.n5024 gnd.n4906 585
R10723 gnd.n5022 gnd.n5021 585
R10724 gnd.n5020 gnd.n1700 585
R10725 gnd.n5017 gnd.n1305 585
R10726 gnd.n5016 gnd.n5015 585
R10727 gnd.n5014 gnd.n5013 585
R10728 gnd.n5012 gnd.n4908 585
R10729 gnd.n5010 gnd.n5009 585
R10730 gnd.n5005 gnd.n4909 585
R10731 gnd.n5004 gnd.n5003 585
R10732 gnd.n5001 gnd.n4910 585
R10733 gnd.n4999 gnd.n4998 585
R10734 gnd.n4997 gnd.n4911 585
R10735 gnd.n4996 gnd.n4995 585
R10736 gnd.n4993 gnd.n4912 585
R10737 gnd.n4991 gnd.n4990 585
R10738 gnd.n4989 gnd.n4913 585
R10739 gnd.n4988 gnd.n4987 585
R10740 gnd.n4985 gnd.n4914 585
R10741 gnd.n4983 gnd.n4982 585
R10742 gnd.n4981 gnd.n4915 585
R10743 gnd.n4980 gnd.n4979 585
R10744 gnd.n4977 gnd.n4916 585
R10745 gnd.n4975 gnd.n4974 585
R10746 gnd.n4973 gnd.n4917 585
R10747 gnd.n4972 gnd.n4971 585
R10748 gnd.n4969 gnd.n4918 585
R10749 gnd.n4967 gnd.n4966 585
R10750 gnd.n4965 gnd.n4919 585
R10751 gnd.n4964 gnd.n4963 585
R10752 gnd.n4961 gnd.n4920 585
R10753 gnd.n4959 gnd.n4958 585
R10754 gnd.n4957 gnd.n4921 585
R10755 gnd.n4956 gnd.n4955 585
R10756 gnd.n4953 gnd.n4922 585
R10757 gnd.n4951 gnd.n4950 585
R10758 gnd.n5086 gnd.n4888 585
R10759 gnd.n5086 gnd.n1698 585
R10760 gnd.n5088 gnd.n5087 585
R10761 gnd.n5087 gnd.n1707 585
R10762 gnd.n5089 gnd.n4884 585
R10763 gnd.n4884 gnd.n1706 585
R10764 gnd.n5091 gnd.n5090 585
R10765 gnd.n5092 gnd.n5091 585
R10766 gnd.n4887 gnd.n4883 585
R10767 gnd.n5094 gnd.n4883 585
R10768 gnd.n4886 gnd.n4885 585
R10769 gnd.n4885 gnd.n1713 585
R10770 gnd.n4875 gnd.n4874 585
R10771 gnd.n4878 gnd.n4875 585
R10772 gnd.n5103 gnd.n5102 585
R10773 gnd.n5102 gnd.n5101 585
R10774 gnd.n5104 gnd.n4871 585
R10775 gnd.n4871 gnd.n1720 585
R10776 gnd.n5106 gnd.n5105 585
R10777 gnd.n5107 gnd.n5106 585
R10778 gnd.n4873 gnd.n4870 585
R10779 gnd.n5109 gnd.n4870 585
R10780 gnd.n4872 gnd.n4862 585
R10781 gnd.n4862 gnd.n1726 585
R10782 gnd.n5116 gnd.n4861 585
R10783 gnd.n5116 gnd.n5115 585
R10784 gnd.n5118 gnd.n5117 585
R10785 gnd.n5117 gnd.n1734 585
R10786 gnd.n5119 gnd.n4859 585
R10787 gnd.n4859 gnd.n1733 585
R10788 gnd.n5121 gnd.n5120 585
R10789 gnd.n5122 gnd.n5121 585
R10790 gnd.n4860 gnd.n4858 585
R10791 gnd.n4858 gnd.n1742 585
R10792 gnd.n4852 gnd.n4851 585
R10793 gnd.n4852 gnd.n1740 585
R10794 gnd.n5131 gnd.n5130 585
R10795 gnd.n5130 gnd.n5129 585
R10796 gnd.n5132 gnd.n4850 585
R10797 gnd.n4850 gnd.n1748 585
R10798 gnd.n5134 gnd.n5133 585
R10799 gnd.n5135 gnd.n5134 585
R10800 gnd.n4843 gnd.n4842 585
R10801 gnd.n4849 gnd.n4843 585
R10802 gnd.n5143 gnd.n5142 585
R10803 gnd.n5142 gnd.n5141 585
R10804 gnd.n5144 gnd.n4839 585
R10805 gnd.n4839 gnd.n1754 585
R10806 gnd.n5146 gnd.n5145 585
R10807 gnd.n5148 gnd.n5146 585
R10808 gnd.n4841 gnd.n4838 585
R10809 gnd.n4838 gnd.n1762 585
R10810 gnd.n4840 gnd.n4830 585
R10811 gnd.n4830 gnd.n1761 585
R10812 gnd.n5156 gnd.n4829 585
R10813 gnd.n5156 gnd.n5155 585
R10814 gnd.n5158 gnd.n5157 585
R10815 gnd.n5157 gnd.n1770 585
R10816 gnd.n5159 gnd.n4826 585
R10817 gnd.n4826 gnd.n1768 585
R10818 gnd.n5161 gnd.n5160 585
R10819 gnd.n5163 gnd.n5161 585
R10820 gnd.n4828 gnd.n4825 585
R10821 gnd.n4825 gnd.n1776 585
R10822 gnd.n4827 gnd.n4816 585
R10823 gnd.n4819 gnd.n4816 585
R10824 gnd.n5171 gnd.n4815 585
R10825 gnd.n5171 gnd.n5170 585
R10826 gnd.n5173 gnd.n5172 585
R10827 gnd.n5172 gnd.n1784 585
R10828 gnd.n5174 gnd.n4813 585
R10829 gnd.n4813 gnd.n1782 585
R10830 gnd.n5176 gnd.n5175 585
R10831 gnd.n5178 gnd.n5176 585
R10832 gnd.n4814 gnd.n4812 585
R10833 gnd.n4812 gnd.n1790 585
R10834 gnd.n4803 gnd.n4802 585
R10835 gnd.n4806 gnd.n4803 585
R10836 gnd.n5187 gnd.n5186 585
R10837 gnd.n5186 gnd.n5185 585
R10838 gnd.n5188 gnd.n4786 585
R10839 gnd.n4786 gnd.n1797 585
R10840 gnd.n5190 gnd.n5189 585
R10841 gnd.n5191 gnd.n5190 585
R10842 gnd.n4801 gnd.n4785 585
R10843 gnd.n5193 gnd.n4785 585
R10844 gnd.n4800 gnd.n4799 585
R10845 gnd.n4799 gnd.n1804 585
R10846 gnd.n4798 gnd.n4787 585
R10847 gnd.n4798 gnd.n1803 585
R10848 gnd.n4797 gnd.n4794 585
R10849 gnd.n4797 gnd.n4796 585
R10850 gnd.n4793 gnd.n4788 585
R10851 gnd.n4788 gnd.n1812 585
R10852 gnd.n4792 gnd.n4791 585
R10853 gnd.n4791 gnd.n1810 585
R10854 gnd.n4790 gnd.n4789 585
R10855 gnd.n4790 gnd.n1820 585
R10856 gnd.n4775 gnd.n4774 585
R10857 gnd.n4775 gnd.n1818 585
R10858 gnd.n5209 gnd.n5208 585
R10859 gnd.n5208 gnd.n5207 585
R10860 gnd.n5210 gnd.n4765 585
R10861 gnd.n4765 gnd.n1827 585
R10862 gnd.n5212 gnd.n5211 585
R10863 gnd.n5213 gnd.n5212 585
R10864 gnd.n4773 gnd.n4764 585
R10865 gnd.n5214 gnd.n4764 585
R10866 gnd.n4772 gnd.n4771 585
R10867 gnd.n4771 gnd.n1833 585
R10868 gnd.n4770 gnd.n4758 585
R10869 gnd.n5220 gnd.n4758 585
R10870 gnd.n4769 gnd.n4757 585
R10871 gnd.n5221 gnd.n4757 585
R10872 gnd.n4768 gnd.n4756 585
R10873 gnd.n5223 gnd.n4756 585
R10874 gnd.n4767 gnd.n4766 585
R10875 gnd.n4766 gnd.n1839 585
R10876 gnd.n4749 gnd.n4748 585
R10877 gnd.n4751 gnd.n4749 585
R10878 gnd.n5232 gnd.n5231 585
R10879 gnd.n5231 gnd.n5230 585
R10880 gnd.n5233 gnd.n4745 585
R10881 gnd.n4745 gnd.n1846 585
R10882 gnd.n5235 gnd.n5234 585
R10883 gnd.n5236 gnd.n5235 585
R10884 gnd.n4747 gnd.n4744 585
R10885 gnd.n4744 gnd.t304 585
R10886 gnd.n4746 gnd.n4735 585
R10887 gnd.n4735 gnd.n1852 585
R10888 gnd.n5244 gnd.n4734 585
R10889 gnd.n5244 gnd.n5243 585
R10890 gnd.n5246 gnd.n5245 585
R10891 gnd.n5245 gnd.n1860 585
R10892 gnd.n5247 gnd.n4665 585
R10893 gnd.n4665 gnd.n1859 585
R10894 gnd.n5249 gnd.n5248 585
R10895 gnd.n5250 gnd.n5249 585
R10896 gnd.n4733 gnd.n4664 585
R10897 gnd.n4664 gnd.n1868 585
R10898 gnd.n4732 gnd.n4731 585
R10899 gnd.n4731 gnd.n1866 585
R10900 gnd.n6346 gnd.n963 585
R10901 gnd.n2177 gnd.n963 585
R10902 gnd.n7150 gnd.n7149 585
R10903 gnd.n7150 gnd.n312 585
R10904 gnd.n7152 gnd.n7151 585
R10905 gnd.n7151 gnd.n358 585
R10906 gnd.n7153 gnd.n416 585
R10907 gnd.n416 gnd.n356 585
R10908 gnd.n7155 gnd.n7154 585
R10909 gnd.n7155 gnd.n377 585
R10910 gnd.n7156 gnd.n415 585
R10911 gnd.n7156 gnd.n370 585
R10912 gnd.n7158 gnd.n7157 585
R10913 gnd.n7157 gnd.n367 585
R10914 gnd.n7159 gnd.n410 585
R10915 gnd.n410 gnd.n384 585
R10916 gnd.n7161 gnd.n7160 585
R10917 gnd.n7162 gnd.n7161 585
R10918 gnd.n411 gnd.n409 585
R10919 gnd.n409 gnd.n390 585
R10920 gnd.n5971 gnd.n5970 585
R10921 gnd.n5971 gnd.n402 585
R10922 gnd.n5972 gnd.n5966 585
R10923 gnd.n5972 gnd.n399 585
R10924 gnd.n5974 gnd.n5973 585
R10925 gnd.n5973 gnd.n1364 585
R10926 gnd.n5975 gnd.n1375 585
R10927 gnd.n1375 gnd.n1361 585
R10928 gnd.n5977 gnd.n5976 585
R10929 gnd.n5978 gnd.n5977 585
R10930 gnd.n1376 gnd.n1374 585
R10931 gnd.n1374 gnd.n1370 585
R10932 gnd.n5960 gnd.n5959 585
R10933 gnd.n5959 gnd.n5958 585
R10934 gnd.n1379 gnd.n1378 585
R10935 gnd.n1396 gnd.n1379 585
R10936 gnd.n5904 gnd.n1409 585
R10937 gnd.n1409 gnd.n1394 585
R10938 gnd.n5906 gnd.n5905 585
R10939 gnd.n5907 gnd.n5906 585
R10940 gnd.n1410 gnd.n1408 585
R10941 gnd.n1408 gnd.n1404 585
R10942 gnd.n5899 gnd.n5898 585
R10943 gnd.n5898 gnd.n5897 585
R10944 gnd.n1413 gnd.n1412 585
R10945 gnd.n1424 gnd.n1413 585
R10946 gnd.n5868 gnd.n1437 585
R10947 gnd.n1437 gnd.n1422 585
R10948 gnd.n5870 gnd.n5869 585
R10949 gnd.n5871 gnd.n5870 585
R10950 gnd.n1438 gnd.n1436 585
R10951 gnd.n1436 gnd.n1431 585
R10952 gnd.n5863 gnd.n5862 585
R10953 gnd.n5862 gnd.n5861 585
R10954 gnd.n1451 gnd.n1440 585
R10955 gnd.n5842 gnd.n1451 585
R10956 gnd.n1450 gnd.n1449 585
R10957 gnd.n1450 gnd.n1338 585
R10958 gnd.n1442 gnd.n1441 585
R10959 gnd.n1441 gnd.n1336 585
R10960 gnd.n1445 gnd.n1444 585
R10961 gnd.n1444 gnd.n1285 585
R10962 gnd.n1255 gnd.n1254 585
R10963 gnd.n6093 gnd.n1255 585
R10964 gnd.n6096 gnd.n6095 585
R10965 gnd.n6095 gnd.n6094 585
R10966 gnd.n6097 gnd.n1249 585
R10967 gnd.n1256 gnd.n1249 585
R10968 gnd.n6099 gnd.n6098 585
R10969 gnd.n6100 gnd.n6099 585
R10970 gnd.n1250 gnd.n1246 585
R10971 gnd.n6101 gnd.n1246 585
R10972 gnd.n5807 gnd.n1621 585
R10973 gnd.n1621 gnd.n1245 585
R10974 gnd.n5809 gnd.n5808 585
R10975 gnd.n5810 gnd.n5809 585
R10976 gnd.n1622 gnd.n1620 585
R10977 gnd.n1620 gnd.n1618 585
R10978 gnd.n5801 gnd.n5800 585
R10979 gnd.n5800 gnd.n5799 585
R10980 gnd.n1625 gnd.n1624 585
R10981 gnd.n1626 gnd.n1625 585
R10982 gnd.n5788 gnd.n5787 585
R10983 gnd.n5789 gnd.n5788 585
R10984 gnd.n1635 gnd.n1634 585
R10985 gnd.n1640 gnd.n1634 585
R10986 gnd.n5783 gnd.n5782 585
R10987 gnd.n5782 gnd.n5781 585
R10988 gnd.n1638 gnd.n1637 585
R10989 gnd.n1639 gnd.n1638 585
R10990 gnd.n5772 gnd.n5771 585
R10991 gnd.n5773 gnd.n5772 585
R10992 gnd.n1649 gnd.n1648 585
R10993 gnd.n1648 gnd.n1646 585
R10994 gnd.n5767 gnd.n5766 585
R10995 gnd.n5766 gnd.n5765 585
R10996 gnd.n1652 gnd.n1651 585
R10997 gnd.n1653 gnd.n1652 585
R10998 gnd.n5756 gnd.n5755 585
R10999 gnd.n5757 gnd.n5756 585
R11000 gnd.n1662 gnd.n1661 585
R11001 gnd.n1661 gnd.n1659 585
R11002 gnd.n5751 gnd.n5750 585
R11003 gnd.n5750 gnd.n5749 585
R11004 gnd.n1665 gnd.n1664 585
R11005 gnd.n1666 gnd.n1665 585
R11006 gnd.n5740 gnd.n5739 585
R11007 gnd.n5741 gnd.n5740 585
R11008 gnd.n1675 gnd.n1674 585
R11009 gnd.n1674 gnd.n1672 585
R11010 gnd.n5735 gnd.n5734 585
R11011 gnd.n5734 gnd.n5733 585
R11012 gnd.n1678 gnd.n1677 585
R11013 gnd.n1686 gnd.n1678 585
R11014 gnd.n5724 gnd.n5723 585
R11015 gnd.n5725 gnd.n5724 585
R11016 gnd.n1688 gnd.n1687 585
R11017 gnd.n1687 gnd.n1684 585
R11018 gnd.n5719 gnd.n5718 585
R11019 gnd.n5718 gnd.n5717 585
R11020 gnd.n1691 gnd.n1690 585
R11021 gnd.n1692 gnd.n1691 585
R11022 gnd.n5708 gnd.n5707 585
R11023 gnd.n5709 gnd.n5708 585
R11024 gnd.n1702 gnd.n1701 585
R11025 gnd.t333 gnd.n1701 585
R11026 gnd.n5703 gnd.n5702 585
R11027 gnd.n5702 gnd.n5701 585
R11028 gnd.n1705 gnd.n1704 585
R11029 gnd.n5093 gnd.n1705 585
R11030 gnd.n5692 gnd.n5691 585
R11031 gnd.n5693 gnd.n5692 585
R11032 gnd.n1716 gnd.n1715 585
R11033 gnd.n4876 gnd.n1715 585
R11034 gnd.n5687 gnd.n5686 585
R11035 gnd.n5686 gnd.n5685 585
R11036 gnd.n1719 gnd.n1718 585
R11037 gnd.n5108 gnd.n1719 585
R11038 gnd.n5676 gnd.n5675 585
R11039 gnd.n5677 gnd.n5676 585
R11040 gnd.n1729 gnd.n1728 585
R11041 gnd.n4863 gnd.n1728 585
R11042 gnd.n5671 gnd.n5670 585
R11043 gnd.n5670 gnd.n5669 585
R11044 gnd.n1732 gnd.n1731 585
R11045 gnd.n4857 gnd.n1732 585
R11046 gnd.n5660 gnd.n5659 585
R11047 gnd.n5661 gnd.n5660 585
R11048 gnd.n1744 gnd.n1743 585
R11049 gnd.n4853 gnd.n1743 585
R11050 gnd.n5655 gnd.n5654 585
R11051 gnd.n5654 gnd.n5653 585
R11052 gnd.n1747 gnd.n1746 585
R11053 gnd.n4844 gnd.n1747 585
R11054 gnd.n5644 gnd.n5643 585
R11055 gnd.n5645 gnd.n5644 585
R11056 gnd.n1757 gnd.n1756 585
R11057 gnd.n5147 gnd.n1756 585
R11058 gnd.n5639 gnd.n5638 585
R11059 gnd.n5638 gnd.n5637 585
R11060 gnd.n1760 gnd.n1759 585
R11061 gnd.n4831 gnd.n1760 585
R11062 gnd.n5628 gnd.n5627 585
R11063 gnd.n5629 gnd.n5628 585
R11064 gnd.n1772 gnd.n1771 585
R11065 gnd.n5162 gnd.n1771 585
R11066 gnd.n5623 gnd.n5622 585
R11067 gnd.n5622 gnd.n5621 585
R11068 gnd.n1775 gnd.n1774 585
R11069 gnd.n4817 gnd.n1775 585
R11070 gnd.n5612 gnd.n5611 585
R11071 gnd.n5613 gnd.n5612 585
R11072 gnd.n1786 gnd.n1785 585
R11073 gnd.n5177 gnd.n1785 585
R11074 gnd.n5607 gnd.n5606 585
R11075 gnd.n5606 gnd.n5605 585
R11076 gnd.n1789 gnd.n1788 585
R11077 gnd.n4804 gnd.n1789 585
R11078 gnd.n5596 gnd.n5595 585
R11079 gnd.n5597 gnd.n5596 585
R11080 gnd.n1799 gnd.n1798 585
R11081 gnd.n5192 gnd.n1798 585
R11082 gnd.n5591 gnd.n5590 585
R11083 gnd.n5590 gnd.n5589 585
R11084 gnd.n1802 gnd.n1801 585
R11085 gnd.n4795 gnd.n1802 585
R11086 gnd.n5580 gnd.n5579 585
R11087 gnd.n5581 gnd.n5580 585
R11088 gnd.n1814 gnd.n1813 585
R11089 gnd.n1819 gnd.n1813 585
R11090 gnd.n5575 gnd.n5574 585
R11091 gnd.n5574 gnd.n5573 585
R11092 gnd.n1817 gnd.n1816 585
R11093 gnd.n4776 gnd.n1817 585
R11094 gnd.n5564 gnd.n5563 585
R11095 gnd.n5565 gnd.n5564 585
R11096 gnd.n1829 gnd.n1828 585
R11097 gnd.n4763 gnd.n1828 585
R11098 gnd.n5559 gnd.n5558 585
R11099 gnd.n5558 gnd.n5557 585
R11100 gnd.n1832 gnd.n1831 585
R11101 gnd.n5222 gnd.n1832 585
R11102 gnd.n5548 gnd.n5547 585
R11103 gnd.n5549 gnd.n5548 585
R11104 gnd.n1842 gnd.n1841 585
R11105 gnd.n4750 gnd.n1841 585
R11106 gnd.n5543 gnd.n5542 585
R11107 gnd.n5542 gnd.n5541 585
R11108 gnd.n1845 gnd.n1844 585
R11109 gnd.n4743 gnd.n1845 585
R11110 gnd.n5532 gnd.n5531 585
R11111 gnd.n5533 gnd.n5532 585
R11112 gnd.n1855 gnd.n1854 585
R11113 gnd.n4736 gnd.n1854 585
R11114 gnd.n5527 gnd.n5526 585
R11115 gnd.n5526 gnd.n5525 585
R11116 gnd.n1858 gnd.n1857 585
R11117 gnd.n4663 gnd.n1858 585
R11118 gnd.n5516 gnd.n5515 585
R11119 gnd.n5517 gnd.n5516 585
R11120 gnd.n1870 gnd.n1869 585
R11121 gnd.n4637 gnd.n1869 585
R11122 gnd.n5511 gnd.n5510 585
R11123 gnd.n5510 gnd.n5509 585
R11124 gnd.n1873 gnd.n1872 585
R11125 gnd.n1874 gnd.n1873 585
R11126 gnd.n5500 gnd.n5499 585
R11127 gnd.n5501 gnd.n5500 585
R11128 gnd.n1883 gnd.n1882 585
R11129 gnd.n1882 gnd.n1880 585
R11130 gnd.n5495 gnd.n5494 585
R11131 gnd.n5494 gnd.n5493 585
R11132 gnd.n1886 gnd.n1885 585
R11133 gnd.n1894 gnd.n1886 585
R11134 gnd.n5484 gnd.n5483 585
R11135 gnd.n5485 gnd.n5484 585
R11136 gnd.n1896 gnd.n1895 585
R11137 gnd.n1895 gnd.n1892 585
R11138 gnd.n5479 gnd.n5478 585
R11139 gnd.n5478 gnd.n5477 585
R11140 gnd.n1899 gnd.n1898 585
R11141 gnd.n1900 gnd.n1899 585
R11142 gnd.n5468 gnd.n5467 585
R11143 gnd.n5469 gnd.n5468 585
R11144 gnd.n1909 gnd.n1908 585
R11145 gnd.n1908 gnd.n1906 585
R11146 gnd.n5463 gnd.n5462 585
R11147 gnd.n5462 gnd.n5461 585
R11148 gnd.n1912 gnd.n1911 585
R11149 gnd.n1913 gnd.n1912 585
R11150 gnd.n5452 gnd.n5451 585
R11151 gnd.n5453 gnd.n5452 585
R11152 gnd.n1922 gnd.n1921 585
R11153 gnd.n1921 gnd.n1919 585
R11154 gnd.n5447 gnd.n5446 585
R11155 gnd.n5446 gnd.n5445 585
R11156 gnd.n1925 gnd.n1924 585
R11157 gnd.n1926 gnd.n1925 585
R11158 gnd.n5436 gnd.n5435 585
R11159 gnd.n5437 gnd.n5436 585
R11160 gnd.n1934 gnd.n1933 585
R11161 gnd.n1939 gnd.n1933 585
R11162 gnd.n5431 gnd.n5430 585
R11163 gnd.n5430 gnd.n5429 585
R11164 gnd.n1937 gnd.n1936 585
R11165 gnd.n1938 gnd.n1937 585
R11166 gnd.n5420 gnd.n5419 585
R11167 gnd.n5421 gnd.n5420 585
R11168 gnd.n1948 gnd.n1947 585
R11169 gnd.n1947 gnd.n1945 585
R11170 gnd.n5415 gnd.n5414 585
R11171 gnd.n5414 gnd.n5413 585
R11172 gnd.n1951 gnd.n1950 585
R11173 gnd.n1952 gnd.n1951 585
R11174 gnd.n4475 gnd.n4474 585
R11175 gnd.n4475 gnd.n1971 585
R11176 gnd.n4476 gnd.n4471 585
R11177 gnd.n4476 gnd.n1958 585
R11178 gnd.n4479 gnd.n4478 585
R11179 gnd.n4478 gnd.n4477 585
R11180 gnd.n4480 gnd.n4466 585
R11181 gnd.n4466 gnd.n2043 585
R11182 gnd.n4482 gnd.n4481 585
R11183 gnd.n4482 gnd.n2027 585
R11184 gnd.n4483 gnd.n4465 585
R11185 gnd.n4483 gnd.n1112 585
R11186 gnd.n4485 gnd.n4484 585
R11187 gnd.n4484 gnd.n1109 585
R11188 gnd.n4486 gnd.n4460 585
R11189 gnd.n4460 gnd.n2109 585
R11190 gnd.n4488 gnd.n4487 585
R11191 gnd.n4488 gnd.n1100 585
R11192 gnd.n4489 gnd.n4459 585
R11193 gnd.n4489 gnd.n1092 585
R11194 gnd.n4491 gnd.n4490 585
R11195 gnd.n4490 gnd.n1089 585
R11196 gnd.n4492 gnd.n2122 585
R11197 gnd.n2122 gnd.n1081 585
R11198 gnd.n4494 gnd.n4493 585
R11199 gnd.n4495 gnd.n4494 585
R11200 gnd.n2123 gnd.n2121 585
R11201 gnd.n2121 gnd.n1071 585
R11202 gnd.n4453 gnd.n4452 585
R11203 gnd.n4452 gnd.n1068 585
R11204 gnd.n4451 gnd.n2125 585
R11205 gnd.n4451 gnd.n1060 585
R11206 gnd.n4450 gnd.n4449 585
R11207 gnd.n4450 gnd.n1057 585
R11208 gnd.n2127 gnd.n2126 585
R11209 gnd.n2126 gnd.n1049 585
R11210 gnd.n4445 gnd.n4444 585
R11211 gnd.n4444 gnd.n4443 585
R11212 gnd.n2130 gnd.n2129 585
R11213 gnd.n2130 gnd.n1039 585
R11214 gnd.n4409 gnd.n4408 585
R11215 gnd.n4410 gnd.n4409 585
R11216 gnd.n2144 gnd.n2143 585
R11217 gnd.n2143 gnd.n1029 585
R11218 gnd.n4404 gnd.n4403 585
R11219 gnd.n4403 gnd.n1026 585
R11220 gnd.n4402 gnd.n2146 585
R11221 gnd.n4402 gnd.n1018 585
R11222 gnd.n4401 gnd.n4400 585
R11223 gnd.n4401 gnd.n1015 585
R11224 gnd.n2148 gnd.n2147 585
R11225 gnd.n2147 gnd.n1007 585
R11226 gnd.n4396 gnd.n4395 585
R11227 gnd.n4395 gnd.n4394 585
R11228 gnd.n2151 gnd.n2150 585
R11229 gnd.n2151 gnd.n997 585
R11230 gnd.n4360 gnd.n4359 585
R11231 gnd.n4361 gnd.n4360 585
R11232 gnd.n4353 gnd.n4352 585
R11233 gnd.n4352 gnd.n986 585
R11234 gnd.n4355 gnd.n4354 585
R11235 gnd.n4354 gnd.n983 585
R11236 gnd.n969 gnd.n968 585
R11237 gnd.n973 gnd.n969 585
R11238 gnd.n6342 gnd.n6341 585
R11239 gnd.n6341 gnd.n6340 585
R11240 gnd.n6103 gnd.n6102 585
R11241 gnd.n6102 gnd.n6101 585
R11242 gnd.n6104 gnd.n1243 585
R11243 gnd.n1245 gnd.n1243 585
R11244 gnd.n1619 gnd.n1241 585
R11245 gnd.n5810 gnd.n1619 585
R11246 gnd.n6108 gnd.n1240 585
R11247 gnd.n1618 gnd.n1240 585
R11248 gnd.n6109 gnd.n1239 585
R11249 gnd.n5799 gnd.n1239 585
R11250 gnd.n6110 gnd.n1238 585
R11251 gnd.n1626 gnd.n1238 585
R11252 gnd.n1633 gnd.n1236 585
R11253 gnd.n5789 gnd.n1633 585
R11254 gnd.n6114 gnd.n1235 585
R11255 gnd.n1640 gnd.n1235 585
R11256 gnd.n6115 gnd.n1234 585
R11257 gnd.n5781 gnd.n1234 585
R11258 gnd.n6116 gnd.n1233 585
R11259 gnd.n1639 gnd.n1233 585
R11260 gnd.n1647 gnd.n1231 585
R11261 gnd.n5773 gnd.n1647 585
R11262 gnd.n6120 gnd.n1230 585
R11263 gnd.n1646 gnd.n1230 585
R11264 gnd.n6121 gnd.n1229 585
R11265 gnd.n5765 gnd.n1229 585
R11266 gnd.n6122 gnd.n1228 585
R11267 gnd.n1653 gnd.n1228 585
R11268 gnd.n1660 gnd.n1226 585
R11269 gnd.n5757 gnd.n1660 585
R11270 gnd.n6126 gnd.n1225 585
R11271 gnd.n1659 gnd.n1225 585
R11272 gnd.n6127 gnd.n1224 585
R11273 gnd.n5749 gnd.n1224 585
R11274 gnd.n6128 gnd.n1223 585
R11275 gnd.n1666 gnd.n1223 585
R11276 gnd.n1673 gnd.n1221 585
R11277 gnd.n5741 gnd.n1673 585
R11278 gnd.n6132 gnd.n1220 585
R11279 gnd.n1672 gnd.n1220 585
R11280 gnd.n6133 gnd.n1219 585
R11281 gnd.n5733 gnd.n1219 585
R11282 gnd.n6134 gnd.n1218 585
R11283 gnd.n1686 gnd.n1218 585
R11284 gnd.n1685 gnd.n1216 585
R11285 gnd.n5725 gnd.n1685 585
R11286 gnd.n6138 gnd.n1215 585
R11287 gnd.n1684 gnd.n1215 585
R11288 gnd.n6139 gnd.n1214 585
R11289 gnd.n5717 gnd.n1214 585
R11290 gnd.n6140 gnd.n1213 585
R11291 gnd.n1692 gnd.n1213 585
R11292 gnd.n1699 gnd.n1211 585
R11293 gnd.n5709 gnd.n1699 585
R11294 gnd.n6144 gnd.n1210 585
R11295 gnd.t333 gnd.n1210 585
R11296 gnd.n6145 gnd.n1209 585
R11297 gnd.n5701 gnd.n1209 585
R11298 gnd.n6146 gnd.n1208 585
R11299 gnd.n5093 gnd.n1208 585
R11300 gnd.n1714 gnd.n1206 585
R11301 gnd.n5693 gnd.n1714 585
R11302 gnd.n6150 gnd.n1205 585
R11303 gnd.n4876 gnd.n1205 585
R11304 gnd.n6151 gnd.n1204 585
R11305 gnd.n5685 gnd.n1204 585
R11306 gnd.n6152 gnd.n1203 585
R11307 gnd.n5108 gnd.n1203 585
R11308 gnd.n1727 gnd.n1201 585
R11309 gnd.n5677 gnd.n1727 585
R11310 gnd.n6156 gnd.n1200 585
R11311 gnd.n4863 gnd.n1200 585
R11312 gnd.n6157 gnd.n1199 585
R11313 gnd.n5669 gnd.n1199 585
R11314 gnd.n6158 gnd.n1198 585
R11315 gnd.n4857 gnd.n1198 585
R11316 gnd.n1741 gnd.n1196 585
R11317 gnd.n5661 gnd.n1741 585
R11318 gnd.n6162 gnd.n1195 585
R11319 gnd.n4853 gnd.n1195 585
R11320 gnd.n6163 gnd.n1194 585
R11321 gnd.n5653 gnd.n1194 585
R11322 gnd.n6164 gnd.n1193 585
R11323 gnd.n4844 gnd.n1193 585
R11324 gnd.n1755 gnd.n1191 585
R11325 gnd.n5645 gnd.n1755 585
R11326 gnd.n6168 gnd.n1190 585
R11327 gnd.n5147 gnd.n1190 585
R11328 gnd.n6169 gnd.n1189 585
R11329 gnd.n5637 gnd.n1189 585
R11330 gnd.n6170 gnd.n1188 585
R11331 gnd.n4831 gnd.n1188 585
R11332 gnd.n1769 gnd.n1186 585
R11333 gnd.n5629 gnd.n1769 585
R11334 gnd.n6174 gnd.n1185 585
R11335 gnd.n5162 gnd.n1185 585
R11336 gnd.n6175 gnd.n1184 585
R11337 gnd.n5621 gnd.n1184 585
R11338 gnd.n6176 gnd.n1183 585
R11339 gnd.n4817 gnd.n1183 585
R11340 gnd.n1783 gnd.n1181 585
R11341 gnd.n5613 gnd.n1783 585
R11342 gnd.n6180 gnd.n1180 585
R11343 gnd.n5177 gnd.n1180 585
R11344 gnd.n6181 gnd.n1179 585
R11345 gnd.n5605 gnd.n1179 585
R11346 gnd.n6182 gnd.n1178 585
R11347 gnd.n4804 gnd.n1178 585
R11348 gnd.n1796 gnd.n1176 585
R11349 gnd.n5597 gnd.n1796 585
R11350 gnd.n6186 gnd.n1175 585
R11351 gnd.n5192 gnd.n1175 585
R11352 gnd.n6187 gnd.n1174 585
R11353 gnd.n5589 gnd.n1174 585
R11354 gnd.n6188 gnd.n1173 585
R11355 gnd.n4795 gnd.n1173 585
R11356 gnd.n1811 gnd.n1171 585
R11357 gnd.n5581 gnd.n1811 585
R11358 gnd.n6192 gnd.n1170 585
R11359 gnd.n1819 gnd.n1170 585
R11360 gnd.n6193 gnd.n1169 585
R11361 gnd.n5573 gnd.n1169 585
R11362 gnd.n6194 gnd.n1168 585
R11363 gnd.n4776 gnd.n1168 585
R11364 gnd.n1826 gnd.n1166 585
R11365 gnd.n5565 gnd.n1826 585
R11366 gnd.n6198 gnd.n1165 585
R11367 gnd.n4763 gnd.n1165 585
R11368 gnd.n6199 gnd.n1164 585
R11369 gnd.n5557 gnd.n1164 585
R11370 gnd.n6200 gnd.n1163 585
R11371 gnd.n5222 gnd.n1163 585
R11372 gnd.n1840 gnd.n1161 585
R11373 gnd.n5549 gnd.n1840 585
R11374 gnd.n6204 gnd.n1160 585
R11375 gnd.n4750 gnd.n1160 585
R11376 gnd.n6205 gnd.n1159 585
R11377 gnd.n5541 gnd.n1159 585
R11378 gnd.n6206 gnd.n1158 585
R11379 gnd.n4743 gnd.n1158 585
R11380 gnd.n1853 gnd.n1156 585
R11381 gnd.n5533 gnd.n1853 585
R11382 gnd.n6210 gnd.n1155 585
R11383 gnd.n4736 gnd.n1155 585
R11384 gnd.n6211 gnd.n1154 585
R11385 gnd.n5525 gnd.n1154 585
R11386 gnd.n6212 gnd.n1153 585
R11387 gnd.n4663 gnd.n1153 585
R11388 gnd.n1867 gnd.n1151 585
R11389 gnd.n5517 gnd.n1867 585
R11390 gnd.n6216 gnd.n1150 585
R11391 gnd.n4637 gnd.n1150 585
R11392 gnd.n6217 gnd.n1149 585
R11393 gnd.n5509 gnd.n1149 585
R11394 gnd.n6218 gnd.n1148 585
R11395 gnd.n1874 gnd.n1148 585
R11396 gnd.n1881 gnd.n1146 585
R11397 gnd.n5501 gnd.n1881 585
R11398 gnd.n6222 gnd.n1145 585
R11399 gnd.n1880 gnd.n1145 585
R11400 gnd.n6223 gnd.n1144 585
R11401 gnd.n5493 gnd.n1144 585
R11402 gnd.n6224 gnd.n1143 585
R11403 gnd.n1894 gnd.n1143 585
R11404 gnd.n1893 gnd.n1141 585
R11405 gnd.n5485 gnd.n1893 585
R11406 gnd.n6228 gnd.n1140 585
R11407 gnd.n1892 gnd.n1140 585
R11408 gnd.n6229 gnd.n1139 585
R11409 gnd.n5477 gnd.n1139 585
R11410 gnd.n6230 gnd.n1138 585
R11411 gnd.n1900 gnd.n1138 585
R11412 gnd.n1907 gnd.n1136 585
R11413 gnd.n5469 gnd.n1907 585
R11414 gnd.n6234 gnd.n1135 585
R11415 gnd.n1906 gnd.n1135 585
R11416 gnd.n6235 gnd.n1134 585
R11417 gnd.n5461 gnd.n1134 585
R11418 gnd.n6236 gnd.n1133 585
R11419 gnd.n1913 gnd.n1133 585
R11420 gnd.n1920 gnd.n1131 585
R11421 gnd.n5453 gnd.n1920 585
R11422 gnd.n6240 gnd.n1130 585
R11423 gnd.n1919 gnd.n1130 585
R11424 gnd.n6241 gnd.n1129 585
R11425 gnd.n5445 gnd.n1129 585
R11426 gnd.n6242 gnd.n1128 585
R11427 gnd.n1926 gnd.n1128 585
R11428 gnd.n1932 gnd.n1126 585
R11429 gnd.n5437 gnd.n1932 585
R11430 gnd.n6246 gnd.n1125 585
R11431 gnd.n1939 gnd.n1125 585
R11432 gnd.n6247 gnd.n1124 585
R11433 gnd.n5429 gnd.n1124 585
R11434 gnd.n6248 gnd.n1123 585
R11435 gnd.n1938 gnd.n1123 585
R11436 gnd.n1946 gnd.n1121 585
R11437 gnd.n5421 gnd.n1946 585
R11438 gnd.n6252 gnd.n1120 585
R11439 gnd.n1945 gnd.n1120 585
R11440 gnd.n6253 gnd.n1119 585
R11441 gnd.n5413 gnd.n1119 585
R11442 gnd.n6254 gnd.n1118 585
R11443 gnd.n1952 gnd.n1118 585
R11444 gnd.n5402 gnd.n5401 585
R11445 gnd.n5400 gnd.n1973 585
R11446 gnd.n1975 gnd.n1972 585
R11447 gnd.n5404 gnd.n1972 585
R11448 gnd.n5393 gnd.n1983 585
R11449 gnd.n5392 gnd.n1984 585
R11450 gnd.n1986 gnd.n1985 585
R11451 gnd.n5385 gnd.n1992 585
R11452 gnd.n5384 gnd.n1993 585
R11453 gnd.n2000 gnd.n1994 585
R11454 gnd.n5377 gnd.n2001 585
R11455 gnd.n5376 gnd.n2002 585
R11456 gnd.n2004 gnd.n2003 585
R11457 gnd.n5369 gnd.n2010 585
R11458 gnd.n5368 gnd.n2011 585
R11459 gnd.n2020 gnd.n2012 585
R11460 gnd.n5361 gnd.n2021 585
R11461 gnd.n5360 gnd.n2022 585
R11462 gnd.n2024 gnd.n2023 585
R11463 gnd.n4546 gnd.n4519 585
R11464 gnd.n4545 gnd.n4520 585
R11465 gnd.n4544 gnd.n4521 585
R11466 gnd.n4523 gnd.n4522 585
R11467 gnd.n4540 gnd.n4525 585
R11468 gnd.n4539 gnd.n4526 585
R11469 gnd.n4538 gnd.n4527 585
R11470 gnd.n4535 gnd.n4532 585
R11471 gnd.n4534 gnd.n4533 585
R11472 gnd.n1957 gnd.n1956 585
R11473 gnd.n5407 gnd.n5406 585
R11474 gnd.n5814 gnd.n1247 585
R11475 gnd.n6101 gnd.n1247 585
R11476 gnd.n5813 gnd.n5812 585
R11477 gnd.n5812 gnd.n1245 585
R11478 gnd.n5811 gnd.n1616 585
R11479 gnd.n5811 gnd.n5810 585
R11480 gnd.n1629 gnd.n1617 585
R11481 gnd.n1618 gnd.n1617 585
R11482 gnd.n5798 gnd.n5797 585
R11483 gnd.n5799 gnd.n5798 585
R11484 gnd.n1628 gnd.n1627 585
R11485 gnd.n1627 gnd.n1626 585
R11486 gnd.n5791 gnd.n5790 585
R11487 gnd.n5790 gnd.n5789 585
R11488 gnd.n1632 gnd.n1631 585
R11489 gnd.n1640 gnd.n1632 585
R11490 gnd.n5780 gnd.n5779 585
R11491 gnd.n5781 gnd.n5780 585
R11492 gnd.n1642 gnd.n1641 585
R11493 gnd.n1641 gnd.n1639 585
R11494 gnd.n5775 gnd.n5774 585
R11495 gnd.n5774 gnd.n5773 585
R11496 gnd.n1645 gnd.n1644 585
R11497 gnd.n1646 gnd.n1645 585
R11498 gnd.n5764 gnd.n5763 585
R11499 gnd.n5765 gnd.n5764 585
R11500 gnd.n1655 gnd.n1654 585
R11501 gnd.n1654 gnd.n1653 585
R11502 gnd.n5759 gnd.n5758 585
R11503 gnd.n5758 gnd.n5757 585
R11504 gnd.n1658 gnd.n1657 585
R11505 gnd.n1659 gnd.n1658 585
R11506 gnd.n5748 gnd.n5747 585
R11507 gnd.n5749 gnd.n5748 585
R11508 gnd.n1668 gnd.n1667 585
R11509 gnd.n1667 gnd.n1666 585
R11510 gnd.n5743 gnd.n5742 585
R11511 gnd.n5742 gnd.n5741 585
R11512 gnd.n1671 gnd.n1670 585
R11513 gnd.n1672 gnd.n1671 585
R11514 gnd.n5732 gnd.n5731 585
R11515 gnd.n5733 gnd.n5732 585
R11516 gnd.n1680 gnd.n1679 585
R11517 gnd.n1686 gnd.n1679 585
R11518 gnd.n5727 gnd.n5726 585
R11519 gnd.n5726 gnd.n5725 585
R11520 gnd.n1683 gnd.n1682 585
R11521 gnd.n1684 gnd.n1683 585
R11522 gnd.n5716 gnd.n5715 585
R11523 gnd.n5717 gnd.n5716 585
R11524 gnd.n1694 gnd.n1693 585
R11525 gnd.n1693 gnd.n1692 585
R11526 gnd.n5711 gnd.n5710 585
R11527 gnd.n5710 gnd.n5709 585
R11528 gnd.n1697 gnd.n1696 585
R11529 gnd.t333 gnd.n1697 585
R11530 gnd.n5700 gnd.n5699 585
R11531 gnd.n5701 gnd.n5700 585
R11532 gnd.n1709 gnd.n1708 585
R11533 gnd.n5093 gnd.n1708 585
R11534 gnd.n5695 gnd.n5694 585
R11535 gnd.n5694 gnd.n5693 585
R11536 gnd.n1712 gnd.n1711 585
R11537 gnd.n4876 gnd.n1712 585
R11538 gnd.n5684 gnd.n5683 585
R11539 gnd.n5685 gnd.n5684 585
R11540 gnd.n1722 gnd.n1721 585
R11541 gnd.n5108 gnd.n1721 585
R11542 gnd.n5679 gnd.n5678 585
R11543 gnd.n5678 gnd.n5677 585
R11544 gnd.n1725 gnd.n1724 585
R11545 gnd.n4863 gnd.n1725 585
R11546 gnd.n5668 gnd.n5667 585
R11547 gnd.n5669 gnd.n5668 585
R11548 gnd.n1736 gnd.n1735 585
R11549 gnd.n4857 gnd.n1735 585
R11550 gnd.n5663 gnd.n5662 585
R11551 gnd.n5662 gnd.n5661 585
R11552 gnd.n1739 gnd.n1738 585
R11553 gnd.n4853 gnd.n1739 585
R11554 gnd.n5652 gnd.n5651 585
R11555 gnd.n5653 gnd.n5652 585
R11556 gnd.n1750 gnd.n1749 585
R11557 gnd.n4844 gnd.n1749 585
R11558 gnd.n5647 gnd.n5646 585
R11559 gnd.n5646 gnd.n5645 585
R11560 gnd.n1753 gnd.n1752 585
R11561 gnd.n5147 gnd.n1753 585
R11562 gnd.n5636 gnd.n5635 585
R11563 gnd.n5637 gnd.n5636 585
R11564 gnd.n1764 gnd.n1763 585
R11565 gnd.n4831 gnd.n1763 585
R11566 gnd.n5631 gnd.n5630 585
R11567 gnd.n5630 gnd.n5629 585
R11568 gnd.n1767 gnd.n1766 585
R11569 gnd.n5162 gnd.n1767 585
R11570 gnd.n5620 gnd.n5619 585
R11571 gnd.n5621 gnd.n5620 585
R11572 gnd.n1778 gnd.n1777 585
R11573 gnd.n4817 gnd.n1777 585
R11574 gnd.n5615 gnd.n5614 585
R11575 gnd.n5614 gnd.n5613 585
R11576 gnd.n1781 gnd.n1780 585
R11577 gnd.n5177 gnd.n1781 585
R11578 gnd.n5604 gnd.n5603 585
R11579 gnd.n5605 gnd.n5604 585
R11580 gnd.n1792 gnd.n1791 585
R11581 gnd.n4804 gnd.n1791 585
R11582 gnd.n5599 gnd.n5598 585
R11583 gnd.n5598 gnd.n5597 585
R11584 gnd.n1795 gnd.n1794 585
R11585 gnd.n5192 gnd.n1795 585
R11586 gnd.n5588 gnd.n5587 585
R11587 gnd.n5589 gnd.n5588 585
R11588 gnd.n1806 gnd.n1805 585
R11589 gnd.n4795 gnd.n1805 585
R11590 gnd.n5583 gnd.n5582 585
R11591 gnd.n5582 gnd.n5581 585
R11592 gnd.n1809 gnd.n1808 585
R11593 gnd.n1819 gnd.n1809 585
R11594 gnd.n5572 gnd.n5571 585
R11595 gnd.n5573 gnd.n5572 585
R11596 gnd.n1822 gnd.n1821 585
R11597 gnd.n4776 gnd.n1821 585
R11598 gnd.n5567 gnd.n5566 585
R11599 gnd.n5566 gnd.n5565 585
R11600 gnd.n1825 gnd.n1824 585
R11601 gnd.n4763 gnd.n1825 585
R11602 gnd.n5556 gnd.n5555 585
R11603 gnd.n5557 gnd.n5556 585
R11604 gnd.n1835 gnd.n1834 585
R11605 gnd.n5222 gnd.n1834 585
R11606 gnd.n5551 gnd.n5550 585
R11607 gnd.n5550 gnd.n5549 585
R11608 gnd.n1838 gnd.n1837 585
R11609 gnd.n4750 gnd.n1838 585
R11610 gnd.n5540 gnd.n5539 585
R11611 gnd.n5541 gnd.n5540 585
R11612 gnd.n1848 gnd.n1847 585
R11613 gnd.n4743 gnd.n1847 585
R11614 gnd.n5535 gnd.n5534 585
R11615 gnd.n5534 gnd.n5533 585
R11616 gnd.n1851 gnd.n1850 585
R11617 gnd.n4736 gnd.n1851 585
R11618 gnd.n5524 gnd.n5523 585
R11619 gnd.n5525 gnd.n5524 585
R11620 gnd.n1862 gnd.n1861 585
R11621 gnd.n4663 gnd.n1861 585
R11622 gnd.n5519 gnd.n5518 585
R11623 gnd.n5518 gnd.n5517 585
R11624 gnd.n1865 gnd.n1864 585
R11625 gnd.n4637 gnd.n1865 585
R11626 gnd.n5508 gnd.n5507 585
R11627 gnd.n5509 gnd.n5508 585
R11628 gnd.n1876 gnd.n1875 585
R11629 gnd.n1875 gnd.n1874 585
R11630 gnd.n5503 gnd.n5502 585
R11631 gnd.n5502 gnd.n5501 585
R11632 gnd.n1879 gnd.n1878 585
R11633 gnd.n1880 gnd.n1879 585
R11634 gnd.n5492 gnd.n5491 585
R11635 gnd.n5493 gnd.n5492 585
R11636 gnd.n1888 gnd.n1887 585
R11637 gnd.n1894 gnd.n1887 585
R11638 gnd.n5487 gnd.n5486 585
R11639 gnd.n5486 gnd.n5485 585
R11640 gnd.n1891 gnd.n1890 585
R11641 gnd.n1892 gnd.n1891 585
R11642 gnd.n5476 gnd.n5475 585
R11643 gnd.n5477 gnd.n5476 585
R11644 gnd.n1902 gnd.n1901 585
R11645 gnd.n1901 gnd.n1900 585
R11646 gnd.n5471 gnd.n5470 585
R11647 gnd.n5470 gnd.n5469 585
R11648 gnd.n1905 gnd.n1904 585
R11649 gnd.n1906 gnd.n1905 585
R11650 gnd.n5460 gnd.n5459 585
R11651 gnd.n5461 gnd.n5460 585
R11652 gnd.n1915 gnd.n1914 585
R11653 gnd.n1914 gnd.n1913 585
R11654 gnd.n5455 gnd.n5454 585
R11655 gnd.n5454 gnd.n5453 585
R11656 gnd.n1918 gnd.n1917 585
R11657 gnd.n1919 gnd.n1918 585
R11658 gnd.n5444 gnd.n5443 585
R11659 gnd.n5445 gnd.n5444 585
R11660 gnd.n1928 gnd.n1927 585
R11661 gnd.n1927 gnd.n1926 585
R11662 gnd.n5439 gnd.n5438 585
R11663 gnd.n5438 gnd.n5437 585
R11664 gnd.n1931 gnd.n1930 585
R11665 gnd.n1939 gnd.n1931 585
R11666 gnd.n5428 gnd.n5427 585
R11667 gnd.n5429 gnd.n5428 585
R11668 gnd.n1941 gnd.n1940 585
R11669 gnd.n1940 gnd.n1938 585
R11670 gnd.n5423 gnd.n5422 585
R11671 gnd.n5422 gnd.n5421 585
R11672 gnd.n1944 gnd.n1943 585
R11673 gnd.n1945 gnd.n1944 585
R11674 gnd.n5412 gnd.n5411 585
R11675 gnd.n5413 gnd.n5412 585
R11676 gnd.n1954 gnd.n1953 585
R11677 gnd.n1953 gnd.n1952 585
R11678 gnd.n5821 gnd.n5820 585
R11679 gnd.n5820 gnd.n1248 585
R11680 gnd.n5822 gnd.n5819 585
R11681 gnd.n5817 gnd.n1614 585
R11682 gnd.n5826 gnd.n1613 585
R11683 gnd.n5830 gnd.n1611 585
R11684 gnd.n5831 gnd.n1610 585
R11685 gnd.n1608 gnd.n1606 585
R11686 gnd.n5835 gnd.n1605 585
R11687 gnd.n5836 gnd.n1603 585
R11688 gnd.n5837 gnd.n1602 585
R11689 gnd.n1600 gnd.n1480 585
R11690 gnd.n1599 gnd.n1598 585
R11691 gnd.n1588 gnd.n1482 585
R11692 gnd.n1590 gnd.n1589 585
R11693 gnd.n1586 gnd.n1492 585
R11694 gnd.n1585 gnd.n1584 585
R11695 gnd.n1572 gnd.n1494 585
R11696 gnd.n1574 gnd.n1573 585
R11697 gnd.n1570 gnd.n1498 585
R11698 gnd.n1569 gnd.n1568 585
R11699 gnd.n1553 gnd.n1500 585
R11700 gnd.n1555 gnd.n1554 585
R11701 gnd.n1551 gnd.n1505 585
R11702 gnd.n1550 gnd.n1549 585
R11703 gnd.n1534 gnd.n1507 585
R11704 gnd.n1536 gnd.n1535 585
R11705 gnd.n1532 gnd.n1512 585
R11706 gnd.n1531 gnd.n1530 585
R11707 gnd.n1514 gnd.n1244 585
R11708 gnd.n4666 gnd.t322 543.808
R11709 gnd.n4904 gnd.t250 543.808
R11710 gnd.n5256 gnd.t266 543.808
R11711 gnd.n5006 gnd.t294 543.808
R11712 gnd.n4951 gnd.n4923 478.086
R11713 gnd.n5086 gnd.n5085 478.086
R11714 gnd.n4731 gnd.n4730 478.086
R11715 gnd.n5319 gnd.n4640 478.086
R11716 gnd.n6519 gnd.n797 440.005
R11717 gnd.n4528 gnd.t283 371.625
R11718 gnd.n122 gnd.t291 371.625
R11719 gnd.n1486 gnd.t306 371.625
R11720 gnd.n2016 gnd.t335 371.625
R11721 gnd.n1308 gnd.t274 371.625
R11722 gnd.n1330 gnd.t262 371.625
R11723 gnd.n201 gnd.t325 371.625
R11724 gnd.n7565 gnd.t246 371.625
R11725 gnd.n3985 gnd.t347 371.625
R11726 gnd.n4017 gnd.t313 371.625
R11727 gnd.n3798 gnd.t344 371.625
R11728 gnd.n2105 gnd.t341 371.625
R11729 gnd.n2083 gnd.t258 371.625
R11730 gnd.n5827 gnd.t254 371.625
R11731 gnd.n2812 gnd.t328 323.425
R11732 gnd.n2357 gnd.t270 323.425
R11733 gnd.n3660 gnd.n3634 289.615
R11734 gnd.n3628 gnd.n3602 289.615
R11735 gnd.n3596 gnd.n3570 289.615
R11736 gnd.n3565 gnd.n3539 289.615
R11737 gnd.n3533 gnd.n3507 289.615
R11738 gnd.n3501 gnd.n3475 289.615
R11739 gnd.n3469 gnd.n3443 289.615
R11740 gnd.n3438 gnd.n3412 289.615
R11741 gnd.n2886 gnd.t309 279.217
R11742 gnd.n2383 gnd.t287 279.217
R11743 gnd.n4647 gnd.t340 260.649
R11744 gnd.n4935 gnd.t302 260.649
R11745 gnd.n5321 gnd.n5320 256.663
R11746 gnd.n5321 gnd.n4606 256.663
R11747 gnd.n5321 gnd.n4607 256.663
R11748 gnd.n5321 gnd.n4608 256.663
R11749 gnd.n5321 gnd.n4609 256.663
R11750 gnd.n5321 gnd.n4610 256.663
R11751 gnd.n5321 gnd.n4611 256.663
R11752 gnd.n5321 gnd.n4612 256.663
R11753 gnd.n5321 gnd.n4613 256.663
R11754 gnd.n5321 gnd.n4614 256.663
R11755 gnd.n5321 gnd.n4615 256.663
R11756 gnd.n5321 gnd.n4616 256.663
R11757 gnd.n5321 gnd.n4617 256.663
R11758 gnd.n5321 gnd.n4618 256.663
R11759 gnd.n5321 gnd.n4619 256.663
R11760 gnd.n5321 gnd.n4620 256.663
R11761 gnd.n5324 gnd.n4604 256.663
R11762 gnd.n5322 gnd.n5321 256.663
R11763 gnd.n5321 gnd.n4621 256.663
R11764 gnd.n5321 gnd.n4622 256.663
R11765 gnd.n5321 gnd.n4623 256.663
R11766 gnd.n5321 gnd.n4624 256.663
R11767 gnd.n5321 gnd.n4625 256.663
R11768 gnd.n5321 gnd.n4626 256.663
R11769 gnd.n5321 gnd.n4627 256.663
R11770 gnd.n5321 gnd.n4628 256.663
R11771 gnd.n5321 gnd.n4629 256.663
R11772 gnd.n5321 gnd.n4630 256.663
R11773 gnd.n5321 gnd.n4631 256.663
R11774 gnd.n5321 gnd.n4632 256.663
R11775 gnd.n5321 gnd.n4633 256.663
R11776 gnd.n5321 gnd.n4634 256.663
R11777 gnd.n5321 gnd.n4635 256.663
R11778 gnd.n5321 gnd.n4636 256.663
R11779 gnd.n4889 gnd.n1700 256.663
R11780 gnd.n5080 gnd.n1700 256.663
R11781 gnd.n5074 gnd.n1700 256.663
R11782 gnd.n5072 gnd.n1700 256.663
R11783 gnd.n5066 gnd.n1700 256.663
R11784 gnd.n5064 gnd.n1700 256.663
R11785 gnd.n5058 gnd.n1700 256.663
R11786 gnd.n5056 gnd.n1700 256.663
R11787 gnd.n5050 gnd.n1700 256.663
R11788 gnd.n5048 gnd.n1700 256.663
R11789 gnd.n5042 gnd.n1700 256.663
R11790 gnd.n5040 gnd.n1700 256.663
R11791 gnd.n5034 gnd.n1700 256.663
R11792 gnd.n5032 gnd.n1700 256.663
R11793 gnd.n5025 gnd.n1700 256.663
R11794 gnd.n5023 gnd.n1700 256.663
R11795 gnd.n5019 gnd.n1305 256.663
R11796 gnd.n5018 gnd.n1700 256.663
R11797 gnd.n4907 gnd.n1700 256.663
R11798 gnd.n5011 gnd.n1700 256.663
R11799 gnd.n5002 gnd.n1700 256.663
R11800 gnd.n5000 gnd.n1700 256.663
R11801 gnd.n4994 gnd.n1700 256.663
R11802 gnd.n4992 gnd.n1700 256.663
R11803 gnd.n4986 gnd.n1700 256.663
R11804 gnd.n4984 gnd.n1700 256.663
R11805 gnd.n4978 gnd.n1700 256.663
R11806 gnd.n4976 gnd.n1700 256.663
R11807 gnd.n4970 gnd.n1700 256.663
R11808 gnd.n4968 gnd.n1700 256.663
R11809 gnd.n4962 gnd.n1700 256.663
R11810 gnd.n4960 gnd.n1700 256.663
R11811 gnd.n4954 gnd.n1700 256.663
R11812 gnd.n4952 gnd.n1700 256.663
R11813 gnd.n3818 gnd.n3793 242.672
R11814 gnd.n3820 gnd.n3793 242.672
R11815 gnd.n3828 gnd.n3793 242.672
R11816 gnd.n3830 gnd.n3793 242.672
R11817 gnd.n3838 gnd.n3793 242.672
R11818 gnd.n3840 gnd.n3793 242.672
R11819 gnd.n3848 gnd.n3793 242.672
R11820 gnd.n3850 gnd.n3793 242.672
R11821 gnd.n3858 gnd.n3793 242.672
R11822 gnd.n5355 gnd.n5354 242.672
R11823 gnd.n5354 gnd.n2042 242.672
R11824 gnd.n5354 gnd.n2041 242.672
R11825 gnd.n5354 gnd.n2039 242.672
R11826 gnd.n5354 gnd.n2037 242.672
R11827 gnd.n5354 gnd.n2036 242.672
R11828 gnd.n5354 gnd.n2034 242.672
R11829 gnd.n5354 gnd.n2032 242.672
R11830 gnd.n5354 gnd.n2031 242.672
R11831 gnd.n6092 gnd.n1275 242.672
R11832 gnd.n6092 gnd.n1276 242.672
R11833 gnd.n6092 gnd.n1277 242.672
R11834 gnd.n6092 gnd.n1278 242.672
R11835 gnd.n6092 gnd.n1279 242.672
R11836 gnd.n6092 gnd.n1280 242.672
R11837 gnd.n6092 gnd.n1281 242.672
R11838 gnd.n6092 gnd.n1282 242.672
R11839 gnd.n6092 gnd.n1283 242.672
R11840 gnd.n128 gnd.n125 242.672
R11841 gnd.n7476 gnd.n128 242.672
R11842 gnd.n7472 gnd.n128 242.672
R11843 gnd.n7469 gnd.n128 242.672
R11844 gnd.n7464 gnd.n128 242.672
R11845 gnd.n7461 gnd.n128 242.672
R11846 gnd.n7456 gnd.n128 242.672
R11847 gnd.n7453 gnd.n128 242.672
R11848 gnd.n7448 gnd.n128 242.672
R11849 gnd.n2940 gnd.n2939 242.672
R11850 gnd.n2940 gnd.n2850 242.672
R11851 gnd.n2940 gnd.n2851 242.672
R11852 gnd.n2940 gnd.n2852 242.672
R11853 gnd.n2940 gnd.n2853 242.672
R11854 gnd.n2940 gnd.n2854 242.672
R11855 gnd.n2940 gnd.n2855 242.672
R11856 gnd.n2940 gnd.n2856 242.672
R11857 gnd.n2940 gnd.n2857 242.672
R11858 gnd.n2940 gnd.n2858 242.672
R11859 gnd.n2940 gnd.n2859 242.672
R11860 gnd.n2940 gnd.n2860 242.672
R11861 gnd.n2941 gnd.n2940 242.672
R11862 gnd.n3792 gnd.n2332 242.672
R11863 gnd.n3792 gnd.n2331 242.672
R11864 gnd.n3792 gnd.n2330 242.672
R11865 gnd.n3792 gnd.n2329 242.672
R11866 gnd.n3792 gnd.n2328 242.672
R11867 gnd.n3792 gnd.n2327 242.672
R11868 gnd.n3792 gnd.n2326 242.672
R11869 gnd.n3792 gnd.n2325 242.672
R11870 gnd.n3792 gnd.n2324 242.672
R11871 gnd.n3792 gnd.n2323 242.672
R11872 gnd.n3792 gnd.n2322 242.672
R11873 gnd.n3792 gnd.n2321 242.672
R11874 gnd.n3792 gnd.n2320 242.672
R11875 gnd.n3024 gnd.n3023 242.672
R11876 gnd.n3023 gnd.n2762 242.672
R11877 gnd.n3023 gnd.n2763 242.672
R11878 gnd.n3023 gnd.n2764 242.672
R11879 gnd.n3023 gnd.n2765 242.672
R11880 gnd.n3023 gnd.n2766 242.672
R11881 gnd.n3023 gnd.n2767 242.672
R11882 gnd.n3023 gnd.n2768 242.672
R11883 gnd.n3792 gnd.n2333 242.672
R11884 gnd.n3792 gnd.n2334 242.672
R11885 gnd.n3792 gnd.n2335 242.672
R11886 gnd.n3792 gnd.n2336 242.672
R11887 gnd.n3792 gnd.n2337 242.672
R11888 gnd.n3792 gnd.n2338 242.672
R11889 gnd.n3792 gnd.n2339 242.672
R11890 gnd.n3792 gnd.n2340 242.672
R11891 gnd.n4171 gnd.n3793 242.672
R11892 gnd.n3961 gnd.n3793 242.672
R11893 gnd.n4164 gnd.n3793 242.672
R11894 gnd.n4158 gnd.n3793 242.672
R11895 gnd.n4156 gnd.n3793 242.672
R11896 gnd.n4150 gnd.n3793 242.672
R11897 gnd.n4148 gnd.n3793 242.672
R11898 gnd.n4142 gnd.n3793 242.672
R11899 gnd.n4140 gnd.n3793 242.672
R11900 gnd.n4134 gnd.n3793 242.672
R11901 gnd.n4132 gnd.n3793 242.672
R11902 gnd.n4126 gnd.n3793 242.672
R11903 gnd.n4124 gnd.n3793 242.672
R11904 gnd.n4118 gnd.n3793 242.672
R11905 gnd.n4116 gnd.n3793 242.672
R11906 gnd.n4110 gnd.n3793 242.672
R11907 gnd.n4108 gnd.n3793 242.672
R11908 gnd.n4015 gnd.n3793 242.672
R11909 gnd.n4098 gnd.n3793 242.672
R11910 gnd.n5354 gnd.n2044 242.672
R11911 gnd.n5354 gnd.n2045 242.672
R11912 gnd.n5354 gnd.n2046 242.672
R11913 gnd.n5354 gnd.n2047 242.672
R11914 gnd.n5354 gnd.n2048 242.672
R11915 gnd.n5354 gnd.n2049 242.672
R11916 gnd.n5354 gnd.n2050 242.672
R11917 gnd.n5354 gnd.n2051 242.672
R11918 gnd.n5354 gnd.n2052 242.672
R11919 gnd.n5354 gnd.n2053 242.672
R11920 gnd.n5354 gnd.n2054 242.672
R11921 gnd.n5325 gnd.n2085 242.672
R11922 gnd.n5354 gnd.n2055 242.672
R11923 gnd.n5354 gnd.n2056 242.672
R11924 gnd.n5354 gnd.n2057 242.672
R11925 gnd.n5354 gnd.n2058 242.672
R11926 gnd.n5354 gnd.n2059 242.672
R11927 gnd.n5354 gnd.n2060 242.672
R11928 gnd.n5354 gnd.n2061 242.672
R11929 gnd.n5354 gnd.n5353 242.672
R11930 gnd.n6092 gnd.n6091 242.672
R11931 gnd.n6092 gnd.n1257 242.672
R11932 gnd.n6092 gnd.n1258 242.672
R11933 gnd.n6092 gnd.n1259 242.672
R11934 gnd.n6092 gnd.n1260 242.672
R11935 gnd.n6092 gnd.n1261 242.672
R11936 gnd.n6092 gnd.n1262 242.672
R11937 gnd.n6092 gnd.n1263 242.672
R11938 gnd.n6060 gnd.n1306 242.672
R11939 gnd.n6092 gnd.n1264 242.672
R11940 gnd.n6092 gnd.n1265 242.672
R11941 gnd.n6092 gnd.n1266 242.672
R11942 gnd.n6092 gnd.n1267 242.672
R11943 gnd.n6092 gnd.n1268 242.672
R11944 gnd.n6092 gnd.n1269 242.672
R11945 gnd.n6092 gnd.n1270 242.672
R11946 gnd.n6092 gnd.n1271 242.672
R11947 gnd.n6092 gnd.n1272 242.672
R11948 gnd.n6092 gnd.n1273 242.672
R11949 gnd.n6092 gnd.n1274 242.672
R11950 gnd.n198 gnd.n128 242.672
R11951 gnd.n7533 gnd.n128 242.672
R11952 gnd.n194 gnd.n128 242.672
R11953 gnd.n7540 gnd.n128 242.672
R11954 gnd.n187 gnd.n128 242.672
R11955 gnd.n7547 gnd.n128 242.672
R11956 gnd.n180 gnd.n128 242.672
R11957 gnd.n7554 gnd.n128 242.672
R11958 gnd.n173 gnd.n128 242.672
R11959 gnd.n7561 gnd.n128 242.672
R11960 gnd.n166 gnd.n128 242.672
R11961 gnd.n7571 gnd.n128 242.672
R11962 gnd.n159 gnd.n128 242.672
R11963 gnd.n7578 gnd.n128 242.672
R11964 gnd.n152 gnd.n128 242.672
R11965 gnd.n7585 gnd.n128 242.672
R11966 gnd.n145 gnd.n128 242.672
R11967 gnd.n7592 gnd.n128 242.672
R11968 gnd.n138 gnd.n128 242.672
R11969 gnd.n5404 gnd.n5403 242.672
R11970 gnd.n5404 gnd.n1959 242.672
R11971 gnd.n5404 gnd.n1960 242.672
R11972 gnd.n5404 gnd.n1961 242.672
R11973 gnd.n5404 gnd.n1962 242.672
R11974 gnd.n5404 gnd.n1963 242.672
R11975 gnd.n5404 gnd.n1964 242.672
R11976 gnd.n5404 gnd.n1965 242.672
R11977 gnd.n5404 gnd.n1966 242.672
R11978 gnd.n5404 gnd.n1967 242.672
R11979 gnd.n5404 gnd.n1968 242.672
R11980 gnd.n5404 gnd.n1969 242.672
R11981 gnd.n5404 gnd.n1970 242.672
R11982 gnd.n5405 gnd.n5404 242.672
R11983 gnd.n5818 gnd.n1248 242.672
R11984 gnd.n1612 gnd.n1248 242.672
R11985 gnd.n1609 gnd.n1248 242.672
R11986 gnd.n1604 gnd.n1248 242.672
R11987 gnd.n1601 gnd.n1248 242.672
R11988 gnd.n1481 gnd.n1248 242.672
R11989 gnd.n1587 gnd.n1248 242.672
R11990 gnd.n1493 gnd.n1248 242.672
R11991 gnd.n1571 gnd.n1248 242.672
R11992 gnd.n1499 gnd.n1248 242.672
R11993 gnd.n1552 gnd.n1248 242.672
R11994 gnd.n1506 gnd.n1248 242.672
R11995 gnd.n1533 gnd.n1248 242.672
R11996 gnd.n1513 gnd.n1248 242.672
R11997 gnd.n135 gnd.n131 240.244
R11998 gnd.n7594 gnd.n7593 240.244
R11999 gnd.n7591 gnd.n139 240.244
R12000 gnd.n7587 gnd.n7586 240.244
R12001 gnd.n7584 gnd.n146 240.244
R12002 gnd.n7580 gnd.n7579 240.244
R12003 gnd.n7577 gnd.n153 240.244
R12004 gnd.n7573 gnd.n7572 240.244
R12005 gnd.n7570 gnd.n160 240.244
R12006 gnd.n7563 gnd.n7562 240.244
R12007 gnd.n7560 gnd.n167 240.244
R12008 gnd.n7556 gnd.n7555 240.244
R12009 gnd.n7553 gnd.n174 240.244
R12010 gnd.n7549 gnd.n7548 240.244
R12011 gnd.n7546 gnd.n181 240.244
R12012 gnd.n7542 gnd.n7541 240.244
R12013 gnd.n7539 gnd.n188 240.244
R12014 gnd.n7535 gnd.n7534 240.244
R12015 gnd.n7532 gnd.n195 240.244
R12016 gnd.n6017 gnd.n1334 240.244
R12017 gnd.n1453 gnd.n1334 240.244
R12018 gnd.n1474 gnd.n1453 240.244
R12019 gnd.n1474 gnd.n1432 240.244
R12020 gnd.n1470 gnd.n1432 240.244
R12021 gnd.n1470 gnd.n1423 240.244
R12022 gnd.n1467 gnd.n1423 240.244
R12023 gnd.n1467 gnd.n1415 240.244
R12024 gnd.n1415 gnd.n1405 240.244
R12025 gnd.n1405 gnd.n1392 240.244
R12026 gnd.n5920 gnd.n1392 240.244
R12027 gnd.n5920 gnd.n1393 240.244
R12028 gnd.n1393 gnd.n1380 240.244
R12029 gnd.n1380 gnd.n1371 240.244
R12030 gnd.n5927 gnd.n1371 240.244
R12031 gnd.n5927 gnd.n1362 240.244
R12032 gnd.n5935 gnd.n1362 240.244
R12033 gnd.n5935 gnd.n400 240.244
R12034 gnd.n400 gnd.n389 240.244
R12035 gnd.n7183 gnd.n389 240.244
R12036 gnd.n7183 gnd.n385 240.244
R12037 gnd.n7195 gnd.n385 240.244
R12038 gnd.n7195 gnd.n368 240.244
R12039 gnd.n7191 gnd.n368 240.244
R12040 gnd.n7191 gnd.n355 240.244
R12041 gnd.n7228 gnd.n355 240.244
R12042 gnd.n7228 gnd.n351 240.244
R12043 gnd.n7241 gnd.n351 240.244
R12044 gnd.n7241 gnd.n313 240.244
R12045 gnd.n7237 gnd.n313 240.244
R12046 gnd.n7237 gnd.n343 240.244
R12047 gnd.n343 gnd.n339 240.244
R12048 gnd.n7258 gnd.n339 240.244
R12049 gnd.n7258 gnd.n335 240.244
R12050 gnd.n7329 gnd.n335 240.244
R12051 gnd.n7329 gnd.n328 240.244
R12052 gnd.n7325 gnd.n328 240.244
R12053 gnd.n7325 gnd.n300 240.244
R12054 gnd.n7322 gnd.n300 240.244
R12055 gnd.n7322 gnd.n291 240.244
R12056 gnd.n7319 gnd.n291 240.244
R12057 gnd.n7319 gnd.n283 240.244
R12058 gnd.n7316 gnd.n283 240.244
R12059 gnd.n7316 gnd.n276 240.244
R12060 gnd.n7313 gnd.n276 240.244
R12061 gnd.n7313 gnd.n270 240.244
R12062 gnd.n7310 gnd.n270 240.244
R12063 gnd.n7310 gnd.n261 240.244
R12064 gnd.n7307 gnd.n261 240.244
R12065 gnd.n7307 gnd.n253 240.244
R12066 gnd.n7304 gnd.n253 240.244
R12067 gnd.n7304 gnd.n245 240.244
R12068 gnd.n7301 gnd.n245 240.244
R12069 gnd.n7301 gnd.n239 240.244
R12070 gnd.n7298 gnd.n239 240.244
R12071 gnd.n7298 gnd.n230 240.244
R12072 gnd.n7295 gnd.n230 240.244
R12073 gnd.n7295 gnd.n223 240.244
R12074 gnd.n7292 gnd.n223 240.244
R12075 gnd.n7292 gnd.n214 240.244
R12076 gnd.n214 gnd.n205 240.244
R12077 gnd.n7523 gnd.n205 240.244
R12078 gnd.n7524 gnd.n7523 240.244
R12079 gnd.n7524 gnd.n127 240.244
R12080 gnd.n1287 gnd.n1286 240.244
R12081 gnd.n6085 gnd.n1286 240.244
R12082 gnd.n6083 gnd.n6082 240.244
R12083 gnd.n6079 gnd.n6078 240.244
R12084 gnd.n6075 gnd.n6074 240.244
R12085 gnd.n6071 gnd.n6070 240.244
R12086 gnd.n6067 gnd.n6066 240.244
R12087 gnd.n6063 gnd.n6062 240.244
R12088 gnd.n6058 gnd.n6057 240.244
R12089 gnd.n6054 gnd.n6053 240.244
R12090 gnd.n6050 gnd.n6049 240.244
R12091 gnd.n6046 gnd.n6045 240.244
R12092 gnd.n6042 gnd.n6041 240.244
R12093 gnd.n6038 gnd.n6037 240.244
R12094 gnd.n6034 gnd.n6033 240.244
R12095 gnd.n6030 gnd.n6029 240.244
R12096 gnd.n6026 gnd.n6025 240.244
R12097 gnd.n1329 gnd.n1328 240.244
R12098 gnd.n5850 gnd.n1288 240.244
R12099 gnd.n5850 gnd.n5843 240.244
R12100 gnd.n5843 gnd.n1430 240.244
R12101 gnd.n5873 gnd.n1430 240.244
R12102 gnd.n5873 gnd.n1425 240.244
R12103 gnd.n5881 gnd.n1425 240.244
R12104 gnd.n5881 gnd.n1426 240.244
R12105 gnd.n1426 gnd.n1403 240.244
R12106 gnd.n5910 gnd.n1403 240.244
R12107 gnd.n5910 gnd.n1397 240.244
R12108 gnd.n5918 gnd.n1397 240.244
R12109 gnd.n5918 gnd.n1399 240.244
R12110 gnd.n1399 gnd.n1369 240.244
R12111 gnd.n5980 gnd.n1369 240.244
R12112 gnd.n5980 gnd.n1365 240.244
R12113 gnd.n5986 gnd.n1365 240.244
R12114 gnd.n5986 gnd.n398 240.244
R12115 gnd.n7173 gnd.n398 240.244
R12116 gnd.n7173 gnd.n393 240.244
R12117 gnd.n7181 gnd.n393 240.244
R12118 gnd.n7181 gnd.n394 240.244
R12119 gnd.n394 gnd.n365 240.244
R12120 gnd.n7219 gnd.n365 240.244
R12121 gnd.n7219 gnd.n366 240.244
R12122 gnd.n366 gnd.n360 240.244
R12123 gnd.n7226 gnd.n360 240.244
R12124 gnd.n7226 gnd.n361 240.244
R12125 gnd.n361 gnd.n310 240.244
R12126 gnd.n7350 gnd.n310 240.244
R12127 gnd.n7350 gnd.n311 240.244
R12128 gnd.n7252 gnd.n311 240.244
R12129 gnd.n7253 gnd.n7252 240.244
R12130 gnd.n7256 gnd.n7253 240.244
R12131 gnd.n7256 gnd.n330 240.244
R12132 gnd.n7331 gnd.n330 240.244
R12133 gnd.n7333 gnd.n7331 240.244
R12134 gnd.n7333 gnd.n301 240.244
R12135 gnd.n7357 gnd.n301 240.244
R12136 gnd.n7357 gnd.n289 240.244
R12137 gnd.n7367 gnd.n289 240.244
R12138 gnd.n7367 gnd.n285 240.244
R12139 gnd.n7373 gnd.n285 240.244
R12140 gnd.n7373 gnd.n275 240.244
R12141 gnd.n7383 gnd.n275 240.244
R12142 gnd.n7383 gnd.n271 240.244
R12143 gnd.n7389 gnd.n271 240.244
R12144 gnd.n7389 gnd.n259 240.244
R12145 gnd.n7399 gnd.n259 240.244
R12146 gnd.n7399 gnd.n255 240.244
R12147 gnd.n7405 gnd.n255 240.244
R12148 gnd.n7405 gnd.n244 240.244
R12149 gnd.n7415 gnd.n244 240.244
R12150 gnd.n7415 gnd.n240 240.244
R12151 gnd.n7421 gnd.n240 240.244
R12152 gnd.n7421 gnd.n228 240.244
R12153 gnd.n7431 gnd.n228 240.244
R12154 gnd.n7431 gnd.n224 240.244
R12155 gnd.n7437 gnd.n224 240.244
R12156 gnd.n7437 gnd.n212 240.244
R12157 gnd.n7515 gnd.n212 240.244
R12158 gnd.n7515 gnd.n208 240.244
R12159 gnd.n7521 gnd.n208 240.244
R12160 gnd.n7521 gnd.n130 240.244
R12161 gnd.n7601 gnd.n130 240.244
R12162 gnd.n2062 gnd.n1108 240.244
R12163 gnd.n5352 gnd.n2063 240.244
R12164 gnd.n5348 gnd.n5347 240.244
R12165 gnd.n5344 gnd.n5343 240.244
R12166 gnd.n5340 gnd.n5339 240.244
R12167 gnd.n5336 gnd.n5335 240.244
R12168 gnd.n5332 gnd.n5331 240.244
R12169 gnd.n5328 gnd.n5327 240.244
R12170 gnd.n4597 gnd.n4596 240.244
R12171 gnd.n4594 gnd.n4593 240.244
R12172 gnd.n4590 gnd.n4589 240.244
R12173 gnd.n4586 gnd.n4585 240.244
R12174 gnd.n4582 gnd.n4581 240.244
R12175 gnd.n4578 gnd.n4577 240.244
R12176 gnd.n4574 gnd.n4573 240.244
R12177 gnd.n4570 gnd.n4569 240.244
R12178 gnd.n4566 gnd.n4565 240.244
R12179 gnd.n4562 gnd.n4561 240.244
R12180 gnd.n4021 gnd.n3794 240.244
R12181 gnd.n4021 gnd.n2313 240.244
R12182 gnd.n4091 gnd.n2313 240.244
R12183 gnd.n4091 gnd.n2306 240.244
R12184 gnd.n4088 gnd.n2306 240.244
R12185 gnd.n4088 gnd.n2298 240.244
R12186 gnd.n4085 gnd.n2298 240.244
R12187 gnd.n4085 gnd.n2289 240.244
R12188 gnd.n4082 gnd.n2289 240.244
R12189 gnd.n4082 gnd.n2281 240.244
R12190 gnd.n4079 gnd.n2281 240.244
R12191 gnd.n4079 gnd.n2274 240.244
R12192 gnd.n4076 gnd.n2274 240.244
R12193 gnd.n4076 gnd.n2266 240.244
R12194 gnd.n4073 gnd.n2266 240.244
R12195 gnd.n4073 gnd.n2257 240.244
R12196 gnd.n4070 gnd.n2257 240.244
R12197 gnd.n4070 gnd.n2249 240.244
R12198 gnd.n4067 gnd.n2249 240.244
R12199 gnd.n4067 gnd.n2242 240.244
R12200 gnd.n4064 gnd.n2242 240.244
R12201 gnd.n4064 gnd.n2234 240.244
R12202 gnd.n4061 gnd.n2234 240.244
R12203 gnd.n4061 gnd.n2225 240.244
R12204 gnd.n4058 gnd.n2225 240.244
R12205 gnd.n4058 gnd.n2217 240.244
R12206 gnd.n4055 gnd.n2217 240.244
R12207 gnd.n4055 gnd.n2211 240.244
R12208 gnd.n4052 gnd.n2211 240.244
R12209 gnd.n4052 gnd.n2202 240.244
R12210 gnd.n2202 gnd.n2192 240.244
R12211 gnd.n4310 gnd.n2192 240.244
R12212 gnd.n4310 gnd.n2193 240.244
R12213 gnd.n2193 gnd.n2175 240.244
R12214 gnd.n2175 gnd.n2169 240.244
R12215 gnd.n4336 gnd.n2169 240.244
R12216 gnd.n4337 gnd.n4336 240.244
R12217 gnd.n4337 gnd.n971 240.244
R12218 gnd.n4343 gnd.n971 240.244
R12219 gnd.n4343 gnd.n984 240.244
R12220 gnd.n4363 gnd.n984 240.244
R12221 gnd.n4363 gnd.n995 240.244
R12222 gnd.n2152 gnd.n995 240.244
R12223 gnd.n2152 gnd.n1005 240.244
R12224 gnd.n4371 gnd.n1005 240.244
R12225 gnd.n4371 gnd.n1016 240.244
R12226 gnd.n4377 gnd.n1016 240.244
R12227 gnd.n4377 gnd.n1027 240.244
R12228 gnd.n4412 gnd.n1027 240.244
R12229 gnd.n4412 gnd.n1037 240.244
R12230 gnd.n2131 gnd.n1037 240.244
R12231 gnd.n2131 gnd.n1047 240.244
R12232 gnd.n4420 gnd.n1047 240.244
R12233 gnd.n4420 gnd.n1058 240.244
R12234 gnd.n4430 gnd.n1058 240.244
R12235 gnd.n4430 gnd.n1069 240.244
R12236 gnd.n2120 gnd.n1069 240.244
R12237 gnd.n2120 gnd.n1079 240.244
R12238 gnd.n4505 gnd.n1079 240.244
R12239 gnd.n4505 gnd.n1090 240.244
R12240 gnd.n4512 gnd.n1090 240.244
R12241 gnd.n4512 gnd.n1101 240.244
R12242 gnd.n4554 gnd.n1101 240.244
R12243 gnd.n4554 gnd.n1110 240.244
R12244 gnd.n4172 gnd.n4170 240.244
R12245 gnd.n4170 gnd.n4169 240.244
R12246 gnd.n4166 gnd.n4165 240.244
R12247 gnd.n4163 gnd.n3966 240.244
R12248 gnd.n4159 gnd.n4157 240.244
R12249 gnd.n4155 gnd.n3972 240.244
R12250 gnd.n4151 gnd.n4149 240.244
R12251 gnd.n4147 gnd.n3978 240.244
R12252 gnd.n4143 gnd.n4141 240.244
R12253 gnd.n4139 gnd.n3984 240.244
R12254 gnd.n4135 gnd.n4133 240.244
R12255 gnd.n4131 gnd.n3993 240.244
R12256 gnd.n4127 gnd.n4125 240.244
R12257 gnd.n4123 gnd.n3999 240.244
R12258 gnd.n4119 gnd.n4117 240.244
R12259 gnd.n4115 gnd.n4005 240.244
R12260 gnd.n4111 gnd.n4109 240.244
R12261 gnd.n4107 gnd.n4011 240.244
R12262 gnd.n4097 gnd.n4016 240.244
R12263 gnd.n4178 gnd.n2312 240.244
R12264 gnd.n4188 gnd.n2312 240.244
R12265 gnd.n4188 gnd.n2308 240.244
R12266 gnd.n4194 gnd.n2308 240.244
R12267 gnd.n4194 gnd.n2296 240.244
R12268 gnd.n4204 gnd.n2296 240.244
R12269 gnd.n4204 gnd.n2292 240.244
R12270 gnd.n4210 gnd.n2292 240.244
R12271 gnd.n4210 gnd.n2280 240.244
R12272 gnd.n4220 gnd.n2280 240.244
R12273 gnd.n4220 gnd.n2276 240.244
R12274 gnd.n4226 gnd.n2276 240.244
R12275 gnd.n4226 gnd.n2264 240.244
R12276 gnd.n4236 gnd.n2264 240.244
R12277 gnd.n4236 gnd.n2260 240.244
R12278 gnd.n4242 gnd.n2260 240.244
R12279 gnd.n4242 gnd.n2248 240.244
R12280 gnd.n4252 gnd.n2248 240.244
R12281 gnd.n4252 gnd.n2244 240.244
R12282 gnd.n4258 gnd.n2244 240.244
R12283 gnd.n4258 gnd.n2232 240.244
R12284 gnd.n4268 gnd.n2232 240.244
R12285 gnd.n4268 gnd.n2228 240.244
R12286 gnd.n4275 gnd.n2228 240.244
R12287 gnd.n4275 gnd.n2216 240.244
R12288 gnd.n4285 gnd.n2216 240.244
R12289 gnd.n4285 gnd.n2213 240.244
R12290 gnd.n4291 gnd.n2213 240.244
R12291 gnd.n4291 gnd.n2200 240.244
R12292 gnd.n4302 gnd.n2200 240.244
R12293 gnd.n4302 gnd.n2198 240.244
R12294 gnd.n4308 gnd.n2198 240.244
R12295 gnd.n4308 gnd.n2174 240.244
R12296 gnd.n4329 gnd.n2174 240.244
R12297 gnd.n4329 gnd.n2172 240.244
R12298 gnd.n4334 gnd.n2172 240.244
R12299 gnd.n4334 gnd.n975 240.244
R12300 gnd.n6338 gnd.n975 240.244
R12301 gnd.n6338 gnd.n976 240.244
R12302 gnd.n6334 gnd.n976 240.244
R12303 gnd.n6334 gnd.n982 240.244
R12304 gnd.n6326 gnd.n982 240.244
R12305 gnd.n6326 gnd.n998 240.244
R12306 gnd.n6322 gnd.n998 240.244
R12307 gnd.n6322 gnd.n1004 240.244
R12308 gnd.n6314 gnd.n1004 240.244
R12309 gnd.n6314 gnd.n1019 240.244
R12310 gnd.n6310 gnd.n1019 240.244
R12311 gnd.n6310 gnd.n1025 240.244
R12312 gnd.n6302 gnd.n1025 240.244
R12313 gnd.n6302 gnd.n1040 240.244
R12314 gnd.n6298 gnd.n1040 240.244
R12315 gnd.n6298 gnd.n1046 240.244
R12316 gnd.n6290 gnd.n1046 240.244
R12317 gnd.n6290 gnd.n1061 240.244
R12318 gnd.n6286 gnd.n1061 240.244
R12319 gnd.n6286 gnd.n1067 240.244
R12320 gnd.n6278 gnd.n1067 240.244
R12321 gnd.n6278 gnd.n1082 240.244
R12322 gnd.n6274 gnd.n1082 240.244
R12323 gnd.n6274 gnd.n1088 240.244
R12324 gnd.n6266 gnd.n1088 240.244
R12325 gnd.n6266 gnd.n1103 240.244
R12326 gnd.n6262 gnd.n1103 240.244
R12327 gnd.n3791 gnd.n2342 240.244
R12328 gnd.n3784 gnd.n3783 240.244
R12329 gnd.n3781 gnd.n3780 240.244
R12330 gnd.n3777 gnd.n3776 240.244
R12331 gnd.n3773 gnd.n3772 240.244
R12332 gnd.n3769 gnd.n3768 240.244
R12333 gnd.n3765 gnd.n3764 240.244
R12334 gnd.n3761 gnd.n3760 240.244
R12335 gnd.n3035 gnd.n2747 240.244
R12336 gnd.n3045 gnd.n2747 240.244
R12337 gnd.n3045 gnd.n2738 240.244
R12338 gnd.n2738 gnd.n2727 240.244
R12339 gnd.n3066 gnd.n2727 240.244
R12340 gnd.n3066 gnd.n2721 240.244
R12341 gnd.n3076 gnd.n2721 240.244
R12342 gnd.n3076 gnd.n2710 240.244
R12343 gnd.n2710 gnd.n2702 240.244
R12344 gnd.n3094 gnd.n2702 240.244
R12345 gnd.n3095 gnd.n3094 240.244
R12346 gnd.n3095 gnd.n2687 240.244
R12347 gnd.n3097 gnd.n2687 240.244
R12348 gnd.n3097 gnd.n2673 240.244
R12349 gnd.n3139 gnd.n2673 240.244
R12350 gnd.n3140 gnd.n3139 240.244
R12351 gnd.n3143 gnd.n3140 240.244
R12352 gnd.n3143 gnd.n2628 240.244
R12353 gnd.n2668 gnd.n2628 240.244
R12354 gnd.n2668 gnd.n2638 240.244
R12355 gnd.n3153 gnd.n2638 240.244
R12356 gnd.n3153 gnd.n2659 240.244
R12357 gnd.n3163 gnd.n2659 240.244
R12358 gnd.n3163 gnd.n2545 240.244
R12359 gnd.n3208 gnd.n2545 240.244
R12360 gnd.n3208 gnd.n2531 240.244
R12361 gnd.n3230 gnd.n2531 240.244
R12362 gnd.n3231 gnd.n3230 240.244
R12363 gnd.n3231 gnd.n2518 240.244
R12364 gnd.n2518 gnd.n2507 240.244
R12365 gnd.n3262 gnd.n2507 240.244
R12366 gnd.n3263 gnd.n3262 240.244
R12367 gnd.n3264 gnd.n3263 240.244
R12368 gnd.n3264 gnd.n2492 240.244
R12369 gnd.n2492 gnd.n2491 240.244
R12370 gnd.n2491 gnd.n2476 240.244
R12371 gnd.n3315 gnd.n2476 240.244
R12372 gnd.n3316 gnd.n3315 240.244
R12373 gnd.n3316 gnd.n2463 240.244
R12374 gnd.n2463 gnd.n2452 240.244
R12375 gnd.n3347 gnd.n2452 240.244
R12376 gnd.n3348 gnd.n3347 240.244
R12377 gnd.n3349 gnd.n3348 240.244
R12378 gnd.n3349 gnd.n2436 240.244
R12379 gnd.n2436 gnd.n2435 240.244
R12380 gnd.n2435 gnd.n2422 240.244
R12381 gnd.n3404 gnd.n2422 240.244
R12382 gnd.n3405 gnd.n3404 240.244
R12383 gnd.n3405 gnd.n2409 240.244
R12384 gnd.n2409 gnd.n2399 240.244
R12385 gnd.n3692 gnd.n2399 240.244
R12386 gnd.n3695 gnd.n3692 240.244
R12387 gnd.n3695 gnd.n3694 240.244
R12388 gnd.n3025 gnd.n2760 240.244
R12389 gnd.n2781 gnd.n2760 240.244
R12390 gnd.n2784 gnd.n2783 240.244
R12391 gnd.n2791 gnd.n2790 240.244
R12392 gnd.n2794 gnd.n2793 240.244
R12393 gnd.n2801 gnd.n2800 240.244
R12394 gnd.n2804 gnd.n2803 240.244
R12395 gnd.n2811 gnd.n2810 240.244
R12396 gnd.n3033 gnd.n2757 240.244
R12397 gnd.n2757 gnd.n2736 240.244
R12398 gnd.n3056 gnd.n2736 240.244
R12399 gnd.n3056 gnd.n2730 240.244
R12400 gnd.n3064 gnd.n2730 240.244
R12401 gnd.n3064 gnd.n2732 240.244
R12402 gnd.n2732 gnd.n2708 240.244
R12403 gnd.n3086 gnd.n2708 240.244
R12404 gnd.n3086 gnd.n2704 240.244
R12405 gnd.n3092 gnd.n2704 240.244
R12406 gnd.n3092 gnd.n2686 240.244
R12407 gnd.n3117 gnd.n2686 240.244
R12408 gnd.n3117 gnd.n2681 240.244
R12409 gnd.n3129 gnd.n2681 240.244
R12410 gnd.n3129 gnd.n2682 240.244
R12411 gnd.n3125 gnd.n2682 240.244
R12412 gnd.n3125 gnd.n2630 240.244
R12413 gnd.n3177 gnd.n2630 240.244
R12414 gnd.n3177 gnd.n2631 240.244
R12415 gnd.n3173 gnd.n2631 240.244
R12416 gnd.n3173 gnd.n2637 240.244
R12417 gnd.n2657 gnd.n2637 240.244
R12418 gnd.n2657 gnd.n2543 240.244
R12419 gnd.n3212 gnd.n2543 240.244
R12420 gnd.n3212 gnd.n2538 240.244
R12421 gnd.n3220 gnd.n2538 240.244
R12422 gnd.n3220 gnd.n2539 240.244
R12423 gnd.n2539 gnd.n2516 240.244
R12424 gnd.n3252 gnd.n2516 240.244
R12425 gnd.n3252 gnd.n2511 240.244
R12426 gnd.n3260 gnd.n2511 240.244
R12427 gnd.n3260 gnd.n2512 240.244
R12428 gnd.n2512 gnd.n2489 240.244
R12429 gnd.n3297 gnd.n2489 240.244
R12430 gnd.n3297 gnd.n2484 240.244
R12431 gnd.n3305 gnd.n2484 240.244
R12432 gnd.n3305 gnd.n2485 240.244
R12433 gnd.n2485 gnd.n2461 240.244
R12434 gnd.n3337 gnd.n2461 240.244
R12435 gnd.n3337 gnd.n2456 240.244
R12436 gnd.n3345 gnd.n2456 240.244
R12437 gnd.n3345 gnd.n2457 240.244
R12438 gnd.n2457 gnd.n2434 240.244
R12439 gnd.n3386 gnd.n2434 240.244
R12440 gnd.n3386 gnd.n2429 240.244
R12441 gnd.n3394 gnd.n2429 240.244
R12442 gnd.n3394 gnd.n2430 240.244
R12443 gnd.n2430 gnd.n2407 240.244
R12444 gnd.n3680 gnd.n2407 240.244
R12445 gnd.n3680 gnd.n2402 240.244
R12446 gnd.n3690 gnd.n2402 240.244
R12447 gnd.n3690 gnd.n2403 240.244
R12448 gnd.n2403 gnd.n2341 240.244
R12449 gnd.n2361 gnd.n2319 240.244
R12450 gnd.n3751 gnd.n3750 240.244
R12451 gnd.n3747 gnd.n3746 240.244
R12452 gnd.n3743 gnd.n3742 240.244
R12453 gnd.n3739 gnd.n3738 240.244
R12454 gnd.n3735 gnd.n3734 240.244
R12455 gnd.n3731 gnd.n3730 240.244
R12456 gnd.n3727 gnd.n3726 240.244
R12457 gnd.n3723 gnd.n3722 240.244
R12458 gnd.n3719 gnd.n3718 240.244
R12459 gnd.n3715 gnd.n3714 240.244
R12460 gnd.n3711 gnd.n3710 240.244
R12461 gnd.n3707 gnd.n3706 240.244
R12462 gnd.n2948 gnd.n2845 240.244
R12463 gnd.n2948 gnd.n2838 240.244
R12464 gnd.n2959 gnd.n2838 240.244
R12465 gnd.n2959 gnd.n2834 240.244
R12466 gnd.n2965 gnd.n2834 240.244
R12467 gnd.n2965 gnd.n2826 240.244
R12468 gnd.n2975 gnd.n2826 240.244
R12469 gnd.n2975 gnd.n2821 240.244
R12470 gnd.n3011 gnd.n2821 240.244
R12471 gnd.n3011 gnd.n2822 240.244
R12472 gnd.n2822 gnd.n2769 240.244
R12473 gnd.n3006 gnd.n2769 240.244
R12474 gnd.n3006 gnd.n3005 240.244
R12475 gnd.n3005 gnd.n2748 240.244
R12476 gnd.n3001 gnd.n2748 240.244
R12477 gnd.n3001 gnd.n2739 240.244
R12478 gnd.n2998 gnd.n2739 240.244
R12479 gnd.n2998 gnd.n2997 240.244
R12480 gnd.n2997 gnd.n2722 240.244
R12481 gnd.n2993 gnd.n2722 240.244
R12482 gnd.n2993 gnd.n2711 240.244
R12483 gnd.n2711 gnd.n2692 240.244
R12484 gnd.n3106 gnd.n2692 240.244
R12485 gnd.n3106 gnd.n2688 240.244
R12486 gnd.n3114 gnd.n2688 240.244
R12487 gnd.n3114 gnd.n2679 240.244
R12488 gnd.n2679 gnd.n2615 240.244
R12489 gnd.n3186 gnd.n2615 240.244
R12490 gnd.n3186 gnd.n2616 240.244
R12491 gnd.n2627 gnd.n2616 240.244
R12492 gnd.n2662 gnd.n2627 240.244
R12493 gnd.n2665 gnd.n2662 240.244
R12494 gnd.n2665 gnd.n2639 240.244
R12495 gnd.n2652 gnd.n2639 240.244
R12496 gnd.n2652 gnd.n2649 240.244
R12497 gnd.n2649 gnd.n2546 240.244
R12498 gnd.n3207 gnd.n2546 240.244
R12499 gnd.n3207 gnd.n2536 240.244
R12500 gnd.n3203 gnd.n2536 240.244
R12501 gnd.n3203 gnd.n2530 240.244
R12502 gnd.n3200 gnd.n2530 240.244
R12503 gnd.n3200 gnd.n2519 240.244
R12504 gnd.n3197 gnd.n2519 240.244
R12505 gnd.n3197 gnd.n2497 240.244
R12506 gnd.n3273 gnd.n2497 240.244
R12507 gnd.n3273 gnd.n2493 240.244
R12508 gnd.n3294 gnd.n2493 240.244
R12509 gnd.n3294 gnd.n2482 240.244
R12510 gnd.n3290 gnd.n2482 240.244
R12511 gnd.n3290 gnd.n2475 240.244
R12512 gnd.n3287 gnd.n2475 240.244
R12513 gnd.n3287 gnd.n2464 240.244
R12514 gnd.n3284 gnd.n2464 240.244
R12515 gnd.n3284 gnd.n2441 240.244
R12516 gnd.n3358 gnd.n2441 240.244
R12517 gnd.n3358 gnd.n2437 240.244
R12518 gnd.n3383 gnd.n2437 240.244
R12519 gnd.n3383 gnd.n2428 240.244
R12520 gnd.n3379 gnd.n2428 240.244
R12521 gnd.n3379 gnd.n2421 240.244
R12522 gnd.n3375 gnd.n2421 240.244
R12523 gnd.n3375 gnd.n2410 240.244
R12524 gnd.n3372 gnd.n2410 240.244
R12525 gnd.n3372 gnd.n2390 240.244
R12526 gnd.n3702 gnd.n2390 240.244
R12527 gnd.n2862 gnd.n2861 240.244
R12528 gnd.n2933 gnd.n2861 240.244
R12529 gnd.n2931 gnd.n2930 240.244
R12530 gnd.n2927 gnd.n2926 240.244
R12531 gnd.n2923 gnd.n2922 240.244
R12532 gnd.n2919 gnd.n2918 240.244
R12533 gnd.n2915 gnd.n2914 240.244
R12534 gnd.n2911 gnd.n2910 240.244
R12535 gnd.n2907 gnd.n2906 240.244
R12536 gnd.n2903 gnd.n2902 240.244
R12537 gnd.n2899 gnd.n2898 240.244
R12538 gnd.n2895 gnd.n2894 240.244
R12539 gnd.n2891 gnd.n2849 240.244
R12540 gnd.n2951 gnd.n2843 240.244
R12541 gnd.n2951 gnd.n2839 240.244
R12542 gnd.n2957 gnd.n2839 240.244
R12543 gnd.n2957 gnd.n2832 240.244
R12544 gnd.n2967 gnd.n2832 240.244
R12545 gnd.n2967 gnd.n2828 240.244
R12546 gnd.n2973 gnd.n2828 240.244
R12547 gnd.n2973 gnd.n2819 240.244
R12548 gnd.n3013 gnd.n2819 240.244
R12549 gnd.n3013 gnd.n2770 240.244
R12550 gnd.n3021 gnd.n2770 240.244
R12551 gnd.n3021 gnd.n2771 240.244
R12552 gnd.n2771 gnd.n2749 240.244
R12553 gnd.n3042 gnd.n2749 240.244
R12554 gnd.n3042 gnd.n2741 240.244
R12555 gnd.n3053 gnd.n2741 240.244
R12556 gnd.n3053 gnd.n2742 240.244
R12557 gnd.n2742 gnd.n2723 240.244
R12558 gnd.n3073 gnd.n2723 240.244
R12559 gnd.n3073 gnd.n2713 240.244
R12560 gnd.n3083 gnd.n2713 240.244
R12561 gnd.n3083 gnd.n2694 240.244
R12562 gnd.n3104 gnd.n2694 240.244
R12563 gnd.n3104 gnd.n2696 240.244
R12564 gnd.n2696 gnd.n2677 240.244
R12565 gnd.n3132 gnd.n2677 240.244
R12566 gnd.n3132 gnd.n2619 240.244
R12567 gnd.n3184 gnd.n2619 240.244
R12568 gnd.n3184 gnd.n2620 240.244
R12569 gnd.n3180 gnd.n2620 240.244
R12570 gnd.n3180 gnd.n2626 240.244
R12571 gnd.n2641 gnd.n2626 240.244
R12572 gnd.n3170 gnd.n2641 240.244
R12573 gnd.n3170 gnd.n2642 240.244
R12574 gnd.n3166 gnd.n2642 240.244
R12575 gnd.n3166 gnd.n2648 240.244
R12576 gnd.n2648 gnd.n2535 240.244
R12577 gnd.n3223 gnd.n2535 240.244
R12578 gnd.n3223 gnd.n2528 240.244
R12579 gnd.n3234 gnd.n2528 240.244
R12580 gnd.n3234 gnd.n2521 240.244
R12581 gnd.n3249 gnd.n2521 240.244
R12582 gnd.n3249 gnd.n2522 240.244
R12583 gnd.n2522 gnd.n2500 240.244
R12584 gnd.n3271 gnd.n2500 240.244
R12585 gnd.n3271 gnd.n2501 240.244
R12586 gnd.n2501 gnd.n2480 240.244
R12587 gnd.n3308 gnd.n2480 240.244
R12588 gnd.n3308 gnd.n2473 240.244
R12589 gnd.n3319 gnd.n2473 240.244
R12590 gnd.n3319 gnd.n2466 240.244
R12591 gnd.n3334 gnd.n2466 240.244
R12592 gnd.n3334 gnd.n2467 240.244
R12593 gnd.n2467 gnd.n2444 240.244
R12594 gnd.n3356 gnd.n2444 240.244
R12595 gnd.n3356 gnd.n2446 240.244
R12596 gnd.n2446 gnd.n2426 240.244
R12597 gnd.n3397 gnd.n2426 240.244
R12598 gnd.n3397 gnd.n2419 240.244
R12599 gnd.n3408 gnd.n2419 240.244
R12600 gnd.n3408 gnd.n2412 240.244
R12601 gnd.n3677 gnd.n2412 240.244
R12602 gnd.n3677 gnd.n2413 240.244
R12603 gnd.n2413 gnd.n2394 240.244
R12604 gnd.n3700 gnd.n2394 240.244
R12605 gnd.n7447 gnd.n7446 240.244
R12606 gnd.n7452 gnd.n7449 240.244
R12607 gnd.n7455 gnd.n7454 240.244
R12608 gnd.n7460 gnd.n7457 240.244
R12609 gnd.n7463 gnd.n7462 240.244
R12610 gnd.n7468 gnd.n7465 240.244
R12611 gnd.n7471 gnd.n7470 240.244
R12612 gnd.n7475 gnd.n7473 240.244
R12613 gnd.n7478 gnd.n7477 240.244
R12614 gnd.n5852 gnd.n1337 240.244
R12615 gnd.n5852 gnd.n1475 240.244
R12616 gnd.n5859 gnd.n1475 240.244
R12617 gnd.n5859 gnd.n1433 240.244
R12618 gnd.n1433 gnd.n1421 240.244
R12619 gnd.n5883 gnd.n1421 240.244
R12620 gnd.n5883 gnd.n1416 240.244
R12621 gnd.n5895 gnd.n1416 240.244
R12622 gnd.n5895 gnd.n1406 240.244
R12623 gnd.n5888 gnd.n1406 240.244
R12624 gnd.n5888 gnd.n1395 240.244
R12625 gnd.n1395 gnd.n1381 240.244
R12626 gnd.n5955 gnd.n1381 240.244
R12627 gnd.n5955 gnd.n1372 240.244
R12628 gnd.n1386 gnd.n1372 240.244
R12629 gnd.n1386 gnd.n1363 240.244
R12630 gnd.n5937 gnd.n1363 240.244
R12631 gnd.n5937 gnd.n401 240.244
R12632 gnd.n5942 gnd.n401 240.244
R12633 gnd.n5942 gnd.n391 240.244
R12634 gnd.n391 gnd.n383 240.244
R12635 gnd.n7197 gnd.n383 240.244
R12636 gnd.n7197 gnd.n369 240.244
R12637 gnd.n378 gnd.n369 240.244
R12638 gnd.n7205 gnd.n378 240.244
R12639 gnd.n7205 gnd.n357 240.244
R12640 gnd.n357 gnd.n349 240.244
R12641 gnd.n7243 gnd.n349 240.244
R12642 gnd.n7243 gnd.n314 240.244
R12643 gnd.n344 gnd.n314 240.244
R12644 gnd.n7250 gnd.n344 240.244
R12645 gnd.n7250 gnd.n345 240.244
R12646 gnd.n345 gnd.n82 240.244
R12647 gnd.n83 gnd.n82 240.244
R12648 gnd.n84 gnd.n83 240.244
R12649 gnd.n329 gnd.n84 240.244
R12650 gnd.n329 gnd.n87 240.244
R12651 gnd.n88 gnd.n87 240.244
R12652 gnd.n89 gnd.n88 240.244
R12653 gnd.n292 gnd.n89 240.244
R12654 gnd.n292 gnd.n92 240.244
R12655 gnd.n93 gnd.n92 240.244
R12656 gnd.n94 gnd.n93 240.244
R12657 gnd.n277 gnd.n94 240.244
R12658 gnd.n277 gnd.n97 240.244
R12659 gnd.n98 gnd.n97 240.244
R12660 gnd.n99 gnd.n98 240.244
R12661 gnd.n262 gnd.n99 240.244
R12662 gnd.n262 gnd.n102 240.244
R12663 gnd.n103 gnd.n102 240.244
R12664 gnd.n104 gnd.n103 240.244
R12665 gnd.n246 gnd.n104 240.244
R12666 gnd.n246 gnd.n107 240.244
R12667 gnd.n108 gnd.n107 240.244
R12668 gnd.n109 gnd.n108 240.244
R12669 gnd.n231 gnd.n109 240.244
R12670 gnd.n231 gnd.n112 240.244
R12671 gnd.n113 gnd.n112 240.244
R12672 gnd.n114 gnd.n113 240.244
R12673 gnd.n215 gnd.n114 240.244
R12674 gnd.n215 gnd.n117 240.244
R12675 gnd.n118 gnd.n117 240.244
R12676 gnd.n119 gnd.n118 240.244
R12677 gnd.n7603 gnd.n119 240.244
R12678 gnd.n1523 gnd.n1522 240.244
R12679 gnd.n1526 gnd.n1525 240.244
R12680 gnd.n1542 gnd.n1541 240.244
R12681 gnd.n1545 gnd.n1544 240.244
R12682 gnd.n1561 gnd.n1560 240.244
R12683 gnd.n1564 gnd.n1563 240.244
R12684 gnd.n1579 gnd.n1578 240.244
R12685 gnd.n1490 gnd.n1489 240.244
R12686 gnd.n1485 gnd.n1284 240.244
R12687 gnd.n6015 gnd.n1340 240.244
R12688 gnd.n1344 gnd.n1340 240.244
R12689 gnd.n1345 gnd.n1344 240.244
R12690 gnd.n1346 gnd.n1345 240.244
R12691 gnd.n1434 gnd.n1346 240.244
R12692 gnd.n1434 gnd.n1349 240.244
R12693 gnd.n1350 gnd.n1349 240.244
R12694 gnd.n1351 gnd.n1350 240.244
R12695 gnd.n5908 gnd.n1351 240.244
R12696 gnd.n5908 gnd.n1354 240.244
R12697 gnd.n1355 gnd.n1354 240.244
R12698 gnd.n1356 gnd.n1355 240.244
R12699 gnd.n5956 gnd.n1356 240.244
R12700 gnd.n5956 gnd.n1359 240.244
R12701 gnd.n1360 gnd.n1359 240.244
R12702 gnd.n5988 gnd.n1360 240.244
R12703 gnd.n5988 gnd.n403 240.244
R12704 gnd.n7171 gnd.n403 240.244
R12705 gnd.n7171 gnd.n404 240.244
R12706 gnd.n404 gnd.n392 240.244
R12707 gnd.n7164 gnd.n392 240.244
R12708 gnd.n7164 gnd.n371 240.244
R12709 gnd.n7217 gnd.n371 240.244
R12710 gnd.n7217 gnd.n372 240.244
R12711 gnd.n7207 gnd.n372 240.244
R12712 gnd.n7207 gnd.n359 240.244
R12713 gnd.n7208 gnd.n359 240.244
R12714 gnd.n7208 gnd.n316 240.244
R12715 gnd.n7348 gnd.n316 240.244
R12716 gnd.n7348 gnd.n317 240.244
R12717 gnd.n322 gnd.n317 240.244
R12718 gnd.n323 gnd.n322 240.244
R12719 gnd.n324 gnd.n323 240.244
R12720 gnd.n333 gnd.n324 240.244
R12721 gnd.n333 gnd.n327 240.244
R12722 gnd.n7335 gnd.n327 240.244
R12723 gnd.n7335 gnd.n298 240.244
R12724 gnd.n7359 gnd.n298 240.244
R12725 gnd.n7359 gnd.n294 240.244
R12726 gnd.n7365 gnd.n294 240.244
R12727 gnd.n7365 gnd.n282 240.244
R12728 gnd.n7375 gnd.n282 240.244
R12729 gnd.n7375 gnd.n278 240.244
R12730 gnd.n7381 gnd.n278 240.244
R12731 gnd.n7381 gnd.n268 240.244
R12732 gnd.n7391 gnd.n268 240.244
R12733 gnd.n7391 gnd.n264 240.244
R12734 gnd.n7397 gnd.n264 240.244
R12735 gnd.n7397 gnd.n252 240.244
R12736 gnd.n7407 gnd.n252 240.244
R12737 gnd.n7407 gnd.n248 240.244
R12738 gnd.n7413 gnd.n248 240.244
R12739 gnd.n7413 gnd.n237 240.244
R12740 gnd.n7423 gnd.n237 240.244
R12741 gnd.n7423 gnd.n233 240.244
R12742 gnd.n7429 gnd.n233 240.244
R12743 gnd.n7429 gnd.n222 240.244
R12744 gnd.n7439 gnd.n222 240.244
R12745 gnd.n7439 gnd.n216 240.244
R12746 gnd.n7513 gnd.n216 240.244
R12747 gnd.n7513 gnd.n217 240.244
R12748 gnd.n217 gnd.n207 240.244
R12749 gnd.n7444 gnd.n207 240.244
R12750 gnd.n7444 gnd.n129 240.244
R12751 gnd.n2029 gnd.n1113 240.244
R12752 gnd.n2030 gnd.n1979 240.244
R12753 gnd.n2033 gnd.n1980 240.244
R12754 gnd.n1989 gnd.n1988 240.244
R12755 gnd.n2035 gnd.n1996 240.244
R12756 gnd.n2038 gnd.n1997 240.244
R12757 gnd.n2007 gnd.n2006 240.244
R12758 gnd.n2040 gnd.n2014 240.244
R12759 gnd.n2026 gnd.n2015 240.244
R12760 gnd.n3956 gnd.n3795 240.244
R12761 gnd.n3956 gnd.n2314 240.244
R12762 gnd.n3952 gnd.n2314 240.244
R12763 gnd.n3952 gnd.n2307 240.244
R12764 gnd.n3949 gnd.n2307 240.244
R12765 gnd.n3949 gnd.n2299 240.244
R12766 gnd.n3946 gnd.n2299 240.244
R12767 gnd.n3946 gnd.n2290 240.244
R12768 gnd.n3943 gnd.n2290 240.244
R12769 gnd.n3943 gnd.n2282 240.244
R12770 gnd.n3940 gnd.n2282 240.244
R12771 gnd.n3940 gnd.n2275 240.244
R12772 gnd.n3937 gnd.n2275 240.244
R12773 gnd.n3937 gnd.n2267 240.244
R12774 gnd.n3934 gnd.n2267 240.244
R12775 gnd.n3934 gnd.n2258 240.244
R12776 gnd.n3931 gnd.n2258 240.244
R12777 gnd.n3931 gnd.n2250 240.244
R12778 gnd.n3928 gnd.n2250 240.244
R12779 gnd.n3928 gnd.n2243 240.244
R12780 gnd.n3925 gnd.n2243 240.244
R12781 gnd.n3925 gnd.n2235 240.244
R12782 gnd.n3922 gnd.n2235 240.244
R12783 gnd.n3922 gnd.n2226 240.244
R12784 gnd.n3919 gnd.n2226 240.244
R12785 gnd.n3919 gnd.n2218 240.244
R12786 gnd.n3916 gnd.n2218 240.244
R12787 gnd.n3916 gnd.n2212 240.244
R12788 gnd.n3913 gnd.n2212 240.244
R12789 gnd.n3913 gnd.n2203 240.244
R12790 gnd.n3910 gnd.n2203 240.244
R12791 gnd.n3910 gnd.n2195 240.244
R12792 gnd.n3895 gnd.n2195 240.244
R12793 gnd.n3895 gnd.n2176 240.244
R12794 gnd.n3898 gnd.n2176 240.244
R12795 gnd.n3898 gnd.n2170 240.244
R12796 gnd.n3899 gnd.n2170 240.244
R12797 gnd.n3899 gnd.n972 240.244
R12798 gnd.n4345 gnd.n972 240.244
R12799 gnd.n4345 gnd.n985 240.244
R12800 gnd.n4351 gnd.n985 240.244
R12801 gnd.n4351 gnd.n996 240.244
R12802 gnd.n4392 gnd.n996 240.244
R12803 gnd.n4392 gnd.n1006 240.244
R12804 gnd.n2157 gnd.n1006 240.244
R12805 gnd.n2157 gnd.n1017 240.244
R12806 gnd.n4379 gnd.n1017 240.244
R12807 gnd.n4379 gnd.n1028 240.244
R12808 gnd.n2142 gnd.n1028 240.244
R12809 gnd.n2142 gnd.n1038 240.244
R12810 gnd.n4441 gnd.n1038 240.244
R12811 gnd.n4441 gnd.n1048 240.244
R12812 gnd.n2136 gnd.n1048 240.244
R12813 gnd.n2136 gnd.n1059 240.244
R12814 gnd.n4432 gnd.n1059 240.244
R12815 gnd.n4432 gnd.n1070 240.244
R12816 gnd.n4497 gnd.n1070 240.244
R12817 gnd.n4497 gnd.n1080 240.244
R12818 gnd.n4503 gnd.n1080 240.244
R12819 gnd.n4503 gnd.n1091 240.244
R12820 gnd.n4514 gnd.n1091 240.244
R12821 gnd.n4514 gnd.n1102 240.244
R12822 gnd.n4552 gnd.n1102 240.244
R12823 gnd.n4552 gnd.n1111 240.244
R12824 gnd.n3821 gnd.n3819 240.244
R12825 gnd.n3827 gnd.n3813 240.244
R12826 gnd.n3831 gnd.n3829 240.244
R12827 gnd.n3837 gnd.n3809 240.244
R12828 gnd.n3841 gnd.n3839 240.244
R12829 gnd.n3847 gnd.n3805 240.244
R12830 gnd.n3851 gnd.n3849 240.244
R12831 gnd.n3857 gnd.n3801 240.244
R12832 gnd.n3860 gnd.n3859 240.244
R12833 gnd.n4180 gnd.n2315 240.244
R12834 gnd.n4186 gnd.n2315 240.244
R12835 gnd.n4186 gnd.n2304 240.244
R12836 gnd.n4196 gnd.n2304 240.244
R12837 gnd.n4196 gnd.n2300 240.244
R12838 gnd.n4202 gnd.n2300 240.244
R12839 gnd.n4202 gnd.n2287 240.244
R12840 gnd.n4212 gnd.n2287 240.244
R12841 gnd.n4212 gnd.n2283 240.244
R12842 gnd.n4218 gnd.n2283 240.244
R12843 gnd.n4218 gnd.n2272 240.244
R12844 gnd.n4228 gnd.n2272 240.244
R12845 gnd.n4228 gnd.n2268 240.244
R12846 gnd.n4234 gnd.n2268 240.244
R12847 gnd.n4234 gnd.n2255 240.244
R12848 gnd.n4244 gnd.n2255 240.244
R12849 gnd.n4244 gnd.n2251 240.244
R12850 gnd.n4250 gnd.n2251 240.244
R12851 gnd.n4250 gnd.n2240 240.244
R12852 gnd.n4260 gnd.n2240 240.244
R12853 gnd.n4260 gnd.n2236 240.244
R12854 gnd.n4266 gnd.n2236 240.244
R12855 gnd.n4266 gnd.n2223 240.244
R12856 gnd.n4277 gnd.n2223 240.244
R12857 gnd.n4277 gnd.n2219 240.244
R12858 gnd.n4283 gnd.n2219 240.244
R12859 gnd.n4283 gnd.n2209 240.244
R12860 gnd.n4293 gnd.n2209 240.244
R12861 gnd.n4293 gnd.n2204 240.244
R12862 gnd.n4300 gnd.n2204 240.244
R12863 gnd.n4300 gnd.n2205 240.244
R12864 gnd.n2205 gnd.n2197 240.244
R12865 gnd.n2197 gnd.n2179 240.244
R12866 gnd.n4327 gnd.n2179 240.244
R12867 gnd.n4327 gnd.n2180 240.244
R12868 gnd.n2180 gnd.n2171 240.244
R12869 gnd.n4322 gnd.n2171 240.244
R12870 gnd.n4322 gnd.n974 240.244
R12871 gnd.n987 gnd.n974 240.244
R12872 gnd.n6332 gnd.n987 240.244
R12873 gnd.n6332 gnd.n988 240.244
R12874 gnd.n6328 gnd.n988 240.244
R12875 gnd.n6328 gnd.n994 240.244
R12876 gnd.n6320 gnd.n994 240.244
R12877 gnd.n6320 gnd.n1008 240.244
R12878 gnd.n6316 gnd.n1008 240.244
R12879 gnd.n6316 gnd.n1014 240.244
R12880 gnd.n6308 gnd.n1014 240.244
R12881 gnd.n6308 gnd.n1030 240.244
R12882 gnd.n6304 gnd.n1030 240.244
R12883 gnd.n6304 gnd.n1036 240.244
R12884 gnd.n6296 gnd.n1036 240.244
R12885 gnd.n6296 gnd.n1050 240.244
R12886 gnd.n6292 gnd.n1050 240.244
R12887 gnd.n6292 gnd.n1056 240.244
R12888 gnd.n6284 gnd.n1056 240.244
R12889 gnd.n6284 gnd.n1072 240.244
R12890 gnd.n6280 gnd.n1072 240.244
R12891 gnd.n6280 gnd.n1078 240.244
R12892 gnd.n6272 gnd.n1078 240.244
R12893 gnd.n6272 gnd.n1093 240.244
R12894 gnd.n6268 gnd.n1093 240.244
R12895 gnd.n6268 gnd.n1099 240.244
R12896 gnd.n6260 gnd.n1099 240.244
R12897 gnd.n6518 gnd.n796 240.244
R12898 gnd.n6522 gnd.n796 240.244
R12899 gnd.n6522 gnd.n792 240.244
R12900 gnd.n6528 gnd.n792 240.244
R12901 gnd.n6528 gnd.n790 240.244
R12902 gnd.n6532 gnd.n790 240.244
R12903 gnd.n6532 gnd.n786 240.244
R12904 gnd.n6538 gnd.n786 240.244
R12905 gnd.n6538 gnd.n784 240.244
R12906 gnd.n6542 gnd.n784 240.244
R12907 gnd.n6542 gnd.n780 240.244
R12908 gnd.n6548 gnd.n780 240.244
R12909 gnd.n6548 gnd.n778 240.244
R12910 gnd.n6552 gnd.n778 240.244
R12911 gnd.n6552 gnd.n774 240.244
R12912 gnd.n6558 gnd.n774 240.244
R12913 gnd.n6558 gnd.n772 240.244
R12914 gnd.n6562 gnd.n772 240.244
R12915 gnd.n6562 gnd.n768 240.244
R12916 gnd.n6568 gnd.n768 240.244
R12917 gnd.n6568 gnd.n766 240.244
R12918 gnd.n6572 gnd.n766 240.244
R12919 gnd.n6572 gnd.n762 240.244
R12920 gnd.n6578 gnd.n762 240.244
R12921 gnd.n6578 gnd.n760 240.244
R12922 gnd.n6582 gnd.n760 240.244
R12923 gnd.n6582 gnd.n756 240.244
R12924 gnd.n6588 gnd.n756 240.244
R12925 gnd.n6588 gnd.n754 240.244
R12926 gnd.n6592 gnd.n754 240.244
R12927 gnd.n6592 gnd.n750 240.244
R12928 gnd.n6598 gnd.n750 240.244
R12929 gnd.n6598 gnd.n748 240.244
R12930 gnd.n6602 gnd.n748 240.244
R12931 gnd.n6602 gnd.n744 240.244
R12932 gnd.n6608 gnd.n744 240.244
R12933 gnd.n6608 gnd.n742 240.244
R12934 gnd.n6612 gnd.n742 240.244
R12935 gnd.n6612 gnd.n738 240.244
R12936 gnd.n6618 gnd.n738 240.244
R12937 gnd.n6618 gnd.n736 240.244
R12938 gnd.n6622 gnd.n736 240.244
R12939 gnd.n6622 gnd.n732 240.244
R12940 gnd.n6628 gnd.n732 240.244
R12941 gnd.n6628 gnd.n730 240.244
R12942 gnd.n6632 gnd.n730 240.244
R12943 gnd.n6632 gnd.n726 240.244
R12944 gnd.n6638 gnd.n726 240.244
R12945 gnd.n6638 gnd.n724 240.244
R12946 gnd.n6642 gnd.n724 240.244
R12947 gnd.n6642 gnd.n720 240.244
R12948 gnd.n6648 gnd.n720 240.244
R12949 gnd.n6648 gnd.n718 240.244
R12950 gnd.n6652 gnd.n718 240.244
R12951 gnd.n6652 gnd.n714 240.244
R12952 gnd.n6658 gnd.n714 240.244
R12953 gnd.n6658 gnd.n712 240.244
R12954 gnd.n6662 gnd.n712 240.244
R12955 gnd.n6662 gnd.n708 240.244
R12956 gnd.n6668 gnd.n708 240.244
R12957 gnd.n6668 gnd.n706 240.244
R12958 gnd.n6672 gnd.n706 240.244
R12959 gnd.n6672 gnd.n702 240.244
R12960 gnd.n6678 gnd.n702 240.244
R12961 gnd.n6678 gnd.n700 240.244
R12962 gnd.n6682 gnd.n700 240.244
R12963 gnd.n6682 gnd.n696 240.244
R12964 gnd.n6688 gnd.n696 240.244
R12965 gnd.n6688 gnd.n694 240.244
R12966 gnd.n6692 gnd.n694 240.244
R12967 gnd.n6692 gnd.n690 240.244
R12968 gnd.n6698 gnd.n690 240.244
R12969 gnd.n6698 gnd.n688 240.244
R12970 gnd.n6702 gnd.n688 240.244
R12971 gnd.n6702 gnd.n684 240.244
R12972 gnd.n6708 gnd.n684 240.244
R12973 gnd.n6708 gnd.n682 240.244
R12974 gnd.n6712 gnd.n682 240.244
R12975 gnd.n6712 gnd.n678 240.244
R12976 gnd.n6718 gnd.n678 240.244
R12977 gnd.n6718 gnd.n676 240.244
R12978 gnd.n6722 gnd.n676 240.244
R12979 gnd.n6722 gnd.n672 240.244
R12980 gnd.n6728 gnd.n672 240.244
R12981 gnd.n6728 gnd.n670 240.244
R12982 gnd.n6732 gnd.n670 240.244
R12983 gnd.n6732 gnd.n666 240.244
R12984 gnd.n6738 gnd.n666 240.244
R12985 gnd.n6738 gnd.n664 240.244
R12986 gnd.n6742 gnd.n664 240.244
R12987 gnd.n6742 gnd.n660 240.244
R12988 gnd.n6748 gnd.n660 240.244
R12989 gnd.n6748 gnd.n658 240.244
R12990 gnd.n6752 gnd.n658 240.244
R12991 gnd.n6752 gnd.n654 240.244
R12992 gnd.n6758 gnd.n654 240.244
R12993 gnd.n6758 gnd.n652 240.244
R12994 gnd.n6762 gnd.n652 240.244
R12995 gnd.n6762 gnd.n648 240.244
R12996 gnd.n6768 gnd.n648 240.244
R12997 gnd.n6768 gnd.n646 240.244
R12998 gnd.n6772 gnd.n646 240.244
R12999 gnd.n6772 gnd.n642 240.244
R13000 gnd.n6778 gnd.n642 240.244
R13001 gnd.n6778 gnd.n640 240.244
R13002 gnd.n6782 gnd.n640 240.244
R13003 gnd.n6782 gnd.n636 240.244
R13004 gnd.n6788 gnd.n636 240.244
R13005 gnd.n6788 gnd.n634 240.244
R13006 gnd.n6792 gnd.n634 240.244
R13007 gnd.n6792 gnd.n630 240.244
R13008 gnd.n6798 gnd.n630 240.244
R13009 gnd.n6798 gnd.n628 240.244
R13010 gnd.n6802 gnd.n628 240.244
R13011 gnd.n6802 gnd.n624 240.244
R13012 gnd.n6808 gnd.n624 240.244
R13013 gnd.n6808 gnd.n622 240.244
R13014 gnd.n6812 gnd.n622 240.244
R13015 gnd.n6812 gnd.n618 240.244
R13016 gnd.n6818 gnd.n618 240.244
R13017 gnd.n6818 gnd.n616 240.244
R13018 gnd.n6822 gnd.n616 240.244
R13019 gnd.n6822 gnd.n612 240.244
R13020 gnd.n6828 gnd.n612 240.244
R13021 gnd.n6828 gnd.n610 240.244
R13022 gnd.n6832 gnd.n610 240.244
R13023 gnd.n6832 gnd.n606 240.244
R13024 gnd.n6838 gnd.n606 240.244
R13025 gnd.n6838 gnd.n604 240.244
R13026 gnd.n6842 gnd.n604 240.244
R13027 gnd.n6842 gnd.n600 240.244
R13028 gnd.n6848 gnd.n600 240.244
R13029 gnd.n6848 gnd.n598 240.244
R13030 gnd.n6852 gnd.n598 240.244
R13031 gnd.n6852 gnd.n594 240.244
R13032 gnd.n6858 gnd.n594 240.244
R13033 gnd.n6858 gnd.n592 240.244
R13034 gnd.n6862 gnd.n592 240.244
R13035 gnd.n6862 gnd.n588 240.244
R13036 gnd.n6868 gnd.n588 240.244
R13037 gnd.n6868 gnd.n586 240.244
R13038 gnd.n6872 gnd.n586 240.244
R13039 gnd.n6872 gnd.n582 240.244
R13040 gnd.n6878 gnd.n582 240.244
R13041 gnd.n6878 gnd.n580 240.244
R13042 gnd.n6882 gnd.n580 240.244
R13043 gnd.n6882 gnd.n576 240.244
R13044 gnd.n6888 gnd.n576 240.244
R13045 gnd.n6888 gnd.n574 240.244
R13046 gnd.n6892 gnd.n574 240.244
R13047 gnd.n6892 gnd.n570 240.244
R13048 gnd.n6898 gnd.n570 240.244
R13049 gnd.n6898 gnd.n568 240.244
R13050 gnd.n6902 gnd.n568 240.244
R13051 gnd.n6902 gnd.n564 240.244
R13052 gnd.n6908 gnd.n564 240.244
R13053 gnd.n6908 gnd.n562 240.244
R13054 gnd.n6912 gnd.n562 240.244
R13055 gnd.n6912 gnd.n558 240.244
R13056 gnd.n6918 gnd.n558 240.244
R13057 gnd.n6918 gnd.n556 240.244
R13058 gnd.n6922 gnd.n556 240.244
R13059 gnd.n6922 gnd.n552 240.244
R13060 gnd.n6929 gnd.n552 240.244
R13061 gnd.n6929 gnd.n550 240.244
R13062 gnd.n6933 gnd.n550 240.244
R13063 gnd.n6933 gnd.n547 240.244
R13064 gnd.n6939 gnd.n545 240.244
R13065 gnd.n6943 gnd.n545 240.244
R13066 gnd.n6943 gnd.n541 240.244
R13067 gnd.n6949 gnd.n541 240.244
R13068 gnd.n6949 gnd.n539 240.244
R13069 gnd.n6953 gnd.n539 240.244
R13070 gnd.n6953 gnd.n535 240.244
R13071 gnd.n6959 gnd.n535 240.244
R13072 gnd.n6959 gnd.n533 240.244
R13073 gnd.n6963 gnd.n533 240.244
R13074 gnd.n6963 gnd.n529 240.244
R13075 gnd.n6969 gnd.n529 240.244
R13076 gnd.n6969 gnd.n527 240.244
R13077 gnd.n6973 gnd.n527 240.244
R13078 gnd.n6973 gnd.n523 240.244
R13079 gnd.n6979 gnd.n523 240.244
R13080 gnd.n6979 gnd.n521 240.244
R13081 gnd.n6983 gnd.n521 240.244
R13082 gnd.n6983 gnd.n517 240.244
R13083 gnd.n6989 gnd.n517 240.244
R13084 gnd.n6989 gnd.n515 240.244
R13085 gnd.n6993 gnd.n515 240.244
R13086 gnd.n6993 gnd.n511 240.244
R13087 gnd.n6999 gnd.n511 240.244
R13088 gnd.n6999 gnd.n509 240.244
R13089 gnd.n7003 gnd.n509 240.244
R13090 gnd.n7003 gnd.n505 240.244
R13091 gnd.n7009 gnd.n505 240.244
R13092 gnd.n7009 gnd.n503 240.244
R13093 gnd.n7013 gnd.n503 240.244
R13094 gnd.n7013 gnd.n499 240.244
R13095 gnd.n7019 gnd.n499 240.244
R13096 gnd.n7019 gnd.n497 240.244
R13097 gnd.n7023 gnd.n497 240.244
R13098 gnd.n7023 gnd.n493 240.244
R13099 gnd.n7029 gnd.n493 240.244
R13100 gnd.n7029 gnd.n491 240.244
R13101 gnd.n7033 gnd.n491 240.244
R13102 gnd.n7033 gnd.n487 240.244
R13103 gnd.n7039 gnd.n487 240.244
R13104 gnd.n7039 gnd.n485 240.244
R13105 gnd.n7043 gnd.n485 240.244
R13106 gnd.n7043 gnd.n481 240.244
R13107 gnd.n7049 gnd.n481 240.244
R13108 gnd.n7049 gnd.n479 240.244
R13109 gnd.n7053 gnd.n479 240.244
R13110 gnd.n7053 gnd.n475 240.244
R13111 gnd.n7059 gnd.n475 240.244
R13112 gnd.n7059 gnd.n473 240.244
R13113 gnd.n7063 gnd.n473 240.244
R13114 gnd.n7063 gnd.n469 240.244
R13115 gnd.n7069 gnd.n469 240.244
R13116 gnd.n7069 gnd.n467 240.244
R13117 gnd.n7073 gnd.n467 240.244
R13118 gnd.n7073 gnd.n463 240.244
R13119 gnd.n7079 gnd.n463 240.244
R13120 gnd.n7079 gnd.n461 240.244
R13121 gnd.n7083 gnd.n461 240.244
R13122 gnd.n7083 gnd.n457 240.244
R13123 gnd.n7089 gnd.n457 240.244
R13124 gnd.n7089 gnd.n455 240.244
R13125 gnd.n7093 gnd.n455 240.244
R13126 gnd.n7093 gnd.n451 240.244
R13127 gnd.n7099 gnd.n451 240.244
R13128 gnd.n7099 gnd.n449 240.244
R13129 gnd.n7103 gnd.n449 240.244
R13130 gnd.n7103 gnd.n445 240.244
R13131 gnd.n7109 gnd.n445 240.244
R13132 gnd.n7109 gnd.n443 240.244
R13133 gnd.n7113 gnd.n443 240.244
R13134 gnd.n7113 gnd.n439 240.244
R13135 gnd.n7119 gnd.n439 240.244
R13136 gnd.n7119 gnd.n437 240.244
R13137 gnd.n7123 gnd.n437 240.244
R13138 gnd.n7123 gnd.n433 240.244
R13139 gnd.n7129 gnd.n433 240.244
R13140 gnd.n7129 gnd.n431 240.244
R13141 gnd.n7133 gnd.n431 240.244
R13142 gnd.n7133 gnd.n427 240.244
R13143 gnd.n7139 gnd.n427 240.244
R13144 gnd.n7139 gnd.n425 240.244
R13145 gnd.n7144 gnd.n425 240.244
R13146 gnd.n7144 gnd.n421 240.244
R13147 gnd.n7150 gnd.n421 240.244
R13148 gnd.n6341 gnd.n969 240.244
R13149 gnd.n4354 gnd.n969 240.244
R13150 gnd.n4354 gnd.n4352 240.244
R13151 gnd.n4360 gnd.n4352 240.244
R13152 gnd.n4360 gnd.n2151 240.244
R13153 gnd.n4395 gnd.n2151 240.244
R13154 gnd.n4395 gnd.n2147 240.244
R13155 gnd.n4401 gnd.n2147 240.244
R13156 gnd.n4402 gnd.n4401 240.244
R13157 gnd.n4403 gnd.n4402 240.244
R13158 gnd.n4403 gnd.n2143 240.244
R13159 gnd.n4409 gnd.n2143 240.244
R13160 gnd.n4409 gnd.n2130 240.244
R13161 gnd.n4444 gnd.n2130 240.244
R13162 gnd.n4444 gnd.n2126 240.244
R13163 gnd.n4450 gnd.n2126 240.244
R13164 gnd.n4451 gnd.n4450 240.244
R13165 gnd.n4452 gnd.n4451 240.244
R13166 gnd.n4452 gnd.n2121 240.244
R13167 gnd.n4494 gnd.n2121 240.244
R13168 gnd.n4494 gnd.n2122 240.244
R13169 gnd.n4490 gnd.n2122 240.244
R13170 gnd.n4490 gnd.n4489 240.244
R13171 gnd.n4489 gnd.n4488 240.244
R13172 gnd.n4488 gnd.n4460 240.244
R13173 gnd.n4484 gnd.n4460 240.244
R13174 gnd.n4484 gnd.n4483 240.244
R13175 gnd.n4483 gnd.n4482 240.244
R13176 gnd.n4482 gnd.n4466 240.244
R13177 gnd.n4478 gnd.n4466 240.244
R13178 gnd.n4478 gnd.n4476 240.244
R13179 gnd.n4476 gnd.n4475 240.244
R13180 gnd.n4475 gnd.n1951 240.244
R13181 gnd.n5414 gnd.n1951 240.244
R13182 gnd.n5414 gnd.n1947 240.244
R13183 gnd.n5420 gnd.n1947 240.244
R13184 gnd.n5420 gnd.n1937 240.244
R13185 gnd.n5430 gnd.n1937 240.244
R13186 gnd.n5430 gnd.n1933 240.244
R13187 gnd.n5436 gnd.n1933 240.244
R13188 gnd.n5436 gnd.n1925 240.244
R13189 gnd.n5446 gnd.n1925 240.244
R13190 gnd.n5446 gnd.n1921 240.244
R13191 gnd.n5452 gnd.n1921 240.244
R13192 gnd.n5452 gnd.n1912 240.244
R13193 gnd.n5462 gnd.n1912 240.244
R13194 gnd.n5462 gnd.n1908 240.244
R13195 gnd.n5468 gnd.n1908 240.244
R13196 gnd.n5468 gnd.n1899 240.244
R13197 gnd.n5478 gnd.n1899 240.244
R13198 gnd.n5478 gnd.n1895 240.244
R13199 gnd.n5484 gnd.n1895 240.244
R13200 gnd.n5484 gnd.n1886 240.244
R13201 gnd.n5494 gnd.n1886 240.244
R13202 gnd.n5494 gnd.n1882 240.244
R13203 gnd.n5500 gnd.n1882 240.244
R13204 gnd.n5500 gnd.n1873 240.244
R13205 gnd.n5510 gnd.n1873 240.244
R13206 gnd.n5510 gnd.n1869 240.244
R13207 gnd.n5516 gnd.n1869 240.244
R13208 gnd.n5516 gnd.n1858 240.244
R13209 gnd.n5526 gnd.n1858 240.244
R13210 gnd.n5526 gnd.n1854 240.244
R13211 gnd.n5532 gnd.n1854 240.244
R13212 gnd.n5532 gnd.n1845 240.244
R13213 gnd.n5542 gnd.n1845 240.244
R13214 gnd.n5542 gnd.n1841 240.244
R13215 gnd.n5548 gnd.n1841 240.244
R13216 gnd.n5548 gnd.n1832 240.244
R13217 gnd.n5558 gnd.n1832 240.244
R13218 gnd.n5558 gnd.n1828 240.244
R13219 gnd.n5564 gnd.n1828 240.244
R13220 gnd.n5564 gnd.n1817 240.244
R13221 gnd.n5574 gnd.n1817 240.244
R13222 gnd.n5574 gnd.n1813 240.244
R13223 gnd.n5580 gnd.n1813 240.244
R13224 gnd.n5580 gnd.n1802 240.244
R13225 gnd.n5590 gnd.n1802 240.244
R13226 gnd.n5590 gnd.n1798 240.244
R13227 gnd.n5596 gnd.n1798 240.244
R13228 gnd.n5596 gnd.n1789 240.244
R13229 gnd.n5606 gnd.n1789 240.244
R13230 gnd.n5606 gnd.n1785 240.244
R13231 gnd.n5612 gnd.n1785 240.244
R13232 gnd.n5612 gnd.n1775 240.244
R13233 gnd.n5622 gnd.n1775 240.244
R13234 gnd.n5622 gnd.n1771 240.244
R13235 gnd.n5628 gnd.n1771 240.244
R13236 gnd.n5628 gnd.n1760 240.244
R13237 gnd.n5638 gnd.n1760 240.244
R13238 gnd.n5638 gnd.n1756 240.244
R13239 gnd.n5644 gnd.n1756 240.244
R13240 gnd.n5644 gnd.n1747 240.244
R13241 gnd.n5654 gnd.n1747 240.244
R13242 gnd.n5654 gnd.n1743 240.244
R13243 gnd.n5660 gnd.n1743 240.244
R13244 gnd.n5660 gnd.n1732 240.244
R13245 gnd.n5670 gnd.n1732 240.244
R13246 gnd.n5670 gnd.n1728 240.244
R13247 gnd.n5676 gnd.n1728 240.244
R13248 gnd.n5676 gnd.n1719 240.244
R13249 gnd.n5686 gnd.n1719 240.244
R13250 gnd.n5686 gnd.n1715 240.244
R13251 gnd.n5692 gnd.n1715 240.244
R13252 gnd.n5692 gnd.n1705 240.244
R13253 gnd.n5702 gnd.n1705 240.244
R13254 gnd.n5702 gnd.n1701 240.244
R13255 gnd.n5708 gnd.n1701 240.244
R13256 gnd.n5708 gnd.n1691 240.244
R13257 gnd.n5718 gnd.n1691 240.244
R13258 gnd.n5718 gnd.n1687 240.244
R13259 gnd.n5724 gnd.n1687 240.244
R13260 gnd.n5724 gnd.n1678 240.244
R13261 gnd.n5734 gnd.n1678 240.244
R13262 gnd.n5734 gnd.n1674 240.244
R13263 gnd.n5740 gnd.n1674 240.244
R13264 gnd.n5740 gnd.n1665 240.244
R13265 gnd.n5750 gnd.n1665 240.244
R13266 gnd.n5750 gnd.n1661 240.244
R13267 gnd.n5756 gnd.n1661 240.244
R13268 gnd.n5756 gnd.n1652 240.244
R13269 gnd.n5766 gnd.n1652 240.244
R13270 gnd.n5766 gnd.n1648 240.244
R13271 gnd.n5772 gnd.n1648 240.244
R13272 gnd.n5772 gnd.n1638 240.244
R13273 gnd.n5782 gnd.n1638 240.244
R13274 gnd.n5782 gnd.n1634 240.244
R13275 gnd.n5788 gnd.n1634 240.244
R13276 gnd.n5788 gnd.n1625 240.244
R13277 gnd.n5800 gnd.n1625 240.244
R13278 gnd.n5800 gnd.n1620 240.244
R13279 gnd.n5809 gnd.n1620 240.244
R13280 gnd.n5809 gnd.n1621 240.244
R13281 gnd.n1621 gnd.n1246 240.244
R13282 gnd.n6099 gnd.n1246 240.244
R13283 gnd.n6099 gnd.n1249 240.244
R13284 gnd.n6095 gnd.n1249 240.244
R13285 gnd.n6095 gnd.n1255 240.244
R13286 gnd.n1444 gnd.n1255 240.244
R13287 gnd.n1444 gnd.n1441 240.244
R13288 gnd.n1450 gnd.n1441 240.244
R13289 gnd.n1451 gnd.n1450 240.244
R13290 gnd.n5862 gnd.n1451 240.244
R13291 gnd.n5862 gnd.n1436 240.244
R13292 gnd.n5870 gnd.n1436 240.244
R13293 gnd.n5870 gnd.n1437 240.244
R13294 gnd.n1437 gnd.n1413 240.244
R13295 gnd.n5898 gnd.n1413 240.244
R13296 gnd.n5898 gnd.n1408 240.244
R13297 gnd.n5906 gnd.n1408 240.244
R13298 gnd.n5906 gnd.n1409 240.244
R13299 gnd.n1409 gnd.n1379 240.244
R13300 gnd.n5959 gnd.n1379 240.244
R13301 gnd.n5959 gnd.n1374 240.244
R13302 gnd.n5977 gnd.n1374 240.244
R13303 gnd.n5977 gnd.n1375 240.244
R13304 gnd.n5973 gnd.n1375 240.244
R13305 gnd.n5973 gnd.n5972 240.244
R13306 gnd.n5972 gnd.n5971 240.244
R13307 gnd.n5971 gnd.n409 240.244
R13308 gnd.n7161 gnd.n409 240.244
R13309 gnd.n7161 gnd.n410 240.244
R13310 gnd.n7157 gnd.n410 240.244
R13311 gnd.n7157 gnd.n7156 240.244
R13312 gnd.n7156 gnd.n7155 240.244
R13313 gnd.n7155 gnd.n416 240.244
R13314 gnd.n7151 gnd.n416 240.244
R13315 gnd.n6512 gnd.n798 240.244
R13316 gnd.n6512 gnd.n801 240.244
R13317 gnd.n6508 gnd.n801 240.244
R13318 gnd.n6508 gnd.n803 240.244
R13319 gnd.n6504 gnd.n803 240.244
R13320 gnd.n6504 gnd.n809 240.244
R13321 gnd.n6500 gnd.n809 240.244
R13322 gnd.n6500 gnd.n811 240.244
R13323 gnd.n6496 gnd.n811 240.244
R13324 gnd.n6496 gnd.n817 240.244
R13325 gnd.n6492 gnd.n817 240.244
R13326 gnd.n6492 gnd.n819 240.244
R13327 gnd.n6488 gnd.n819 240.244
R13328 gnd.n6488 gnd.n825 240.244
R13329 gnd.n6484 gnd.n825 240.244
R13330 gnd.n6484 gnd.n827 240.244
R13331 gnd.n6480 gnd.n827 240.244
R13332 gnd.n6480 gnd.n833 240.244
R13333 gnd.n6476 gnd.n833 240.244
R13334 gnd.n6476 gnd.n835 240.244
R13335 gnd.n6472 gnd.n835 240.244
R13336 gnd.n6472 gnd.n841 240.244
R13337 gnd.n6468 gnd.n841 240.244
R13338 gnd.n6468 gnd.n843 240.244
R13339 gnd.n6464 gnd.n843 240.244
R13340 gnd.n6464 gnd.n849 240.244
R13341 gnd.n6460 gnd.n849 240.244
R13342 gnd.n6460 gnd.n851 240.244
R13343 gnd.n6456 gnd.n851 240.244
R13344 gnd.n6456 gnd.n857 240.244
R13345 gnd.n6452 gnd.n857 240.244
R13346 gnd.n6452 gnd.n859 240.244
R13347 gnd.n6448 gnd.n859 240.244
R13348 gnd.n6448 gnd.n865 240.244
R13349 gnd.n6444 gnd.n865 240.244
R13350 gnd.n6444 gnd.n867 240.244
R13351 gnd.n6440 gnd.n867 240.244
R13352 gnd.n6440 gnd.n873 240.244
R13353 gnd.n6436 gnd.n873 240.244
R13354 gnd.n6436 gnd.n875 240.244
R13355 gnd.n6432 gnd.n875 240.244
R13356 gnd.n6432 gnd.n881 240.244
R13357 gnd.n6428 gnd.n881 240.244
R13358 gnd.n6428 gnd.n883 240.244
R13359 gnd.n6424 gnd.n883 240.244
R13360 gnd.n6424 gnd.n889 240.244
R13361 gnd.n6420 gnd.n889 240.244
R13362 gnd.n6420 gnd.n891 240.244
R13363 gnd.n6416 gnd.n891 240.244
R13364 gnd.n6416 gnd.n897 240.244
R13365 gnd.n6412 gnd.n897 240.244
R13366 gnd.n6412 gnd.n899 240.244
R13367 gnd.n6408 gnd.n899 240.244
R13368 gnd.n6408 gnd.n905 240.244
R13369 gnd.n6404 gnd.n905 240.244
R13370 gnd.n6404 gnd.n907 240.244
R13371 gnd.n6400 gnd.n907 240.244
R13372 gnd.n6400 gnd.n913 240.244
R13373 gnd.n6396 gnd.n913 240.244
R13374 gnd.n6396 gnd.n915 240.244
R13375 gnd.n6392 gnd.n915 240.244
R13376 gnd.n6392 gnd.n921 240.244
R13377 gnd.n6388 gnd.n921 240.244
R13378 gnd.n6388 gnd.n923 240.244
R13379 gnd.n6384 gnd.n923 240.244
R13380 gnd.n6384 gnd.n929 240.244
R13381 gnd.n6380 gnd.n929 240.244
R13382 gnd.n6380 gnd.n931 240.244
R13383 gnd.n6376 gnd.n931 240.244
R13384 gnd.n6376 gnd.n937 240.244
R13385 gnd.n6372 gnd.n937 240.244
R13386 gnd.n6372 gnd.n939 240.244
R13387 gnd.n6368 gnd.n939 240.244
R13388 gnd.n6368 gnd.n945 240.244
R13389 gnd.n6364 gnd.n945 240.244
R13390 gnd.n6364 gnd.n947 240.244
R13391 gnd.n6360 gnd.n947 240.244
R13392 gnd.n6360 gnd.n953 240.244
R13393 gnd.n6356 gnd.n953 240.244
R13394 gnd.n6356 gnd.n955 240.244
R13395 gnd.n6352 gnd.n955 240.244
R13396 gnd.n6352 gnd.n961 240.244
R13397 gnd.n6348 gnd.n961 240.244
R13398 gnd.n6348 gnd.n963 240.244
R13399 gnd.n1119 gnd.n1118 240.244
R13400 gnd.n1120 gnd.n1119 240.244
R13401 gnd.n1946 gnd.n1120 240.244
R13402 gnd.n1946 gnd.n1123 240.244
R13403 gnd.n1124 gnd.n1123 240.244
R13404 gnd.n1125 gnd.n1124 240.244
R13405 gnd.n1932 gnd.n1125 240.244
R13406 gnd.n1932 gnd.n1128 240.244
R13407 gnd.n1129 gnd.n1128 240.244
R13408 gnd.n1130 gnd.n1129 240.244
R13409 gnd.n1920 gnd.n1130 240.244
R13410 gnd.n1920 gnd.n1133 240.244
R13411 gnd.n1134 gnd.n1133 240.244
R13412 gnd.n1135 gnd.n1134 240.244
R13413 gnd.n1907 gnd.n1135 240.244
R13414 gnd.n1907 gnd.n1138 240.244
R13415 gnd.n1139 gnd.n1138 240.244
R13416 gnd.n1140 gnd.n1139 240.244
R13417 gnd.n1893 gnd.n1140 240.244
R13418 gnd.n1893 gnd.n1143 240.244
R13419 gnd.n1144 gnd.n1143 240.244
R13420 gnd.n1145 gnd.n1144 240.244
R13421 gnd.n1881 gnd.n1145 240.244
R13422 gnd.n1881 gnd.n1148 240.244
R13423 gnd.n1149 gnd.n1148 240.244
R13424 gnd.n1150 gnd.n1149 240.244
R13425 gnd.n1867 gnd.n1150 240.244
R13426 gnd.n1867 gnd.n1153 240.244
R13427 gnd.n1154 gnd.n1153 240.244
R13428 gnd.n1155 gnd.n1154 240.244
R13429 gnd.n1853 gnd.n1155 240.244
R13430 gnd.n1853 gnd.n1158 240.244
R13431 gnd.n1159 gnd.n1158 240.244
R13432 gnd.n1160 gnd.n1159 240.244
R13433 gnd.n1840 gnd.n1160 240.244
R13434 gnd.n1840 gnd.n1163 240.244
R13435 gnd.n1164 gnd.n1163 240.244
R13436 gnd.n1165 gnd.n1164 240.244
R13437 gnd.n1826 gnd.n1165 240.244
R13438 gnd.n1826 gnd.n1168 240.244
R13439 gnd.n1169 gnd.n1168 240.244
R13440 gnd.n1170 gnd.n1169 240.244
R13441 gnd.n1811 gnd.n1170 240.244
R13442 gnd.n1811 gnd.n1173 240.244
R13443 gnd.n1174 gnd.n1173 240.244
R13444 gnd.n1175 gnd.n1174 240.244
R13445 gnd.n1796 gnd.n1175 240.244
R13446 gnd.n1796 gnd.n1178 240.244
R13447 gnd.n1179 gnd.n1178 240.244
R13448 gnd.n1180 gnd.n1179 240.244
R13449 gnd.n1783 gnd.n1180 240.244
R13450 gnd.n1783 gnd.n1183 240.244
R13451 gnd.n1184 gnd.n1183 240.244
R13452 gnd.n1185 gnd.n1184 240.244
R13453 gnd.n1769 gnd.n1185 240.244
R13454 gnd.n1769 gnd.n1188 240.244
R13455 gnd.n1189 gnd.n1188 240.244
R13456 gnd.n1190 gnd.n1189 240.244
R13457 gnd.n1755 gnd.n1190 240.244
R13458 gnd.n1755 gnd.n1193 240.244
R13459 gnd.n1194 gnd.n1193 240.244
R13460 gnd.n1195 gnd.n1194 240.244
R13461 gnd.n1741 gnd.n1195 240.244
R13462 gnd.n1741 gnd.n1198 240.244
R13463 gnd.n1199 gnd.n1198 240.244
R13464 gnd.n1200 gnd.n1199 240.244
R13465 gnd.n1727 gnd.n1200 240.244
R13466 gnd.n1727 gnd.n1203 240.244
R13467 gnd.n1204 gnd.n1203 240.244
R13468 gnd.n1205 gnd.n1204 240.244
R13469 gnd.n1714 gnd.n1205 240.244
R13470 gnd.n1714 gnd.n1208 240.244
R13471 gnd.n1209 gnd.n1208 240.244
R13472 gnd.n1210 gnd.n1209 240.244
R13473 gnd.n1699 gnd.n1210 240.244
R13474 gnd.n1699 gnd.n1213 240.244
R13475 gnd.n1214 gnd.n1213 240.244
R13476 gnd.n1215 gnd.n1214 240.244
R13477 gnd.n1685 gnd.n1215 240.244
R13478 gnd.n1685 gnd.n1218 240.244
R13479 gnd.n1219 gnd.n1218 240.244
R13480 gnd.n1220 gnd.n1219 240.244
R13481 gnd.n1673 gnd.n1220 240.244
R13482 gnd.n1673 gnd.n1223 240.244
R13483 gnd.n1224 gnd.n1223 240.244
R13484 gnd.n1225 gnd.n1224 240.244
R13485 gnd.n1660 gnd.n1225 240.244
R13486 gnd.n1660 gnd.n1228 240.244
R13487 gnd.n1229 gnd.n1228 240.244
R13488 gnd.n1230 gnd.n1229 240.244
R13489 gnd.n1647 gnd.n1230 240.244
R13490 gnd.n1647 gnd.n1233 240.244
R13491 gnd.n1234 gnd.n1233 240.244
R13492 gnd.n1235 gnd.n1234 240.244
R13493 gnd.n1633 gnd.n1235 240.244
R13494 gnd.n1633 gnd.n1238 240.244
R13495 gnd.n1239 gnd.n1238 240.244
R13496 gnd.n1240 gnd.n1239 240.244
R13497 gnd.n1619 gnd.n1240 240.244
R13498 gnd.n1619 gnd.n1243 240.244
R13499 gnd.n6102 gnd.n1243 240.244
R13500 gnd.n1973 gnd.n1972 240.244
R13501 gnd.n1983 gnd.n1972 240.244
R13502 gnd.n1985 gnd.n1984 240.244
R13503 gnd.n1993 gnd.n1992 240.244
R13504 gnd.n2001 gnd.n2000 240.244
R13505 gnd.n2003 gnd.n2002 240.244
R13506 gnd.n2011 gnd.n2010 240.244
R13507 gnd.n2021 gnd.n2020 240.244
R13508 gnd.n2023 gnd.n2022 240.244
R13509 gnd.n4520 gnd.n4519 240.244
R13510 gnd.n4522 gnd.n4521 240.244
R13511 gnd.n4526 gnd.n4525 240.244
R13512 gnd.n4532 gnd.n4527 240.244
R13513 gnd.n4533 gnd.n1957 240.244
R13514 gnd.n5412 gnd.n1953 240.244
R13515 gnd.n5412 gnd.n1944 240.244
R13516 gnd.n5422 gnd.n1944 240.244
R13517 gnd.n5422 gnd.n1940 240.244
R13518 gnd.n5428 gnd.n1940 240.244
R13519 gnd.n5428 gnd.n1931 240.244
R13520 gnd.n5438 gnd.n1931 240.244
R13521 gnd.n5438 gnd.n1927 240.244
R13522 gnd.n5444 gnd.n1927 240.244
R13523 gnd.n5444 gnd.n1918 240.244
R13524 gnd.n5454 gnd.n1918 240.244
R13525 gnd.n5454 gnd.n1914 240.244
R13526 gnd.n5460 gnd.n1914 240.244
R13527 gnd.n5460 gnd.n1905 240.244
R13528 gnd.n5470 gnd.n1905 240.244
R13529 gnd.n5470 gnd.n1901 240.244
R13530 gnd.n5476 gnd.n1901 240.244
R13531 gnd.n5476 gnd.n1891 240.244
R13532 gnd.n5486 gnd.n1891 240.244
R13533 gnd.n5486 gnd.n1887 240.244
R13534 gnd.n5492 gnd.n1887 240.244
R13535 gnd.n5492 gnd.n1879 240.244
R13536 gnd.n5502 gnd.n1879 240.244
R13537 gnd.n5502 gnd.n1875 240.244
R13538 gnd.n5508 gnd.n1875 240.244
R13539 gnd.n5508 gnd.n1865 240.244
R13540 gnd.n5518 gnd.n1865 240.244
R13541 gnd.n5518 gnd.n1861 240.244
R13542 gnd.n5524 gnd.n1861 240.244
R13543 gnd.n5524 gnd.n1851 240.244
R13544 gnd.n5534 gnd.n1851 240.244
R13545 gnd.n5534 gnd.n1847 240.244
R13546 gnd.n5540 gnd.n1847 240.244
R13547 gnd.n5540 gnd.n1838 240.244
R13548 gnd.n5550 gnd.n1838 240.244
R13549 gnd.n5550 gnd.n1834 240.244
R13550 gnd.n5556 gnd.n1834 240.244
R13551 gnd.n5556 gnd.n1825 240.244
R13552 gnd.n5566 gnd.n1825 240.244
R13553 gnd.n5566 gnd.n1821 240.244
R13554 gnd.n5572 gnd.n1821 240.244
R13555 gnd.n5572 gnd.n1809 240.244
R13556 gnd.n5582 gnd.n1809 240.244
R13557 gnd.n5582 gnd.n1805 240.244
R13558 gnd.n5588 gnd.n1805 240.244
R13559 gnd.n5588 gnd.n1795 240.244
R13560 gnd.n5598 gnd.n1795 240.244
R13561 gnd.n5598 gnd.n1791 240.244
R13562 gnd.n5604 gnd.n1791 240.244
R13563 gnd.n5604 gnd.n1781 240.244
R13564 gnd.n5614 gnd.n1781 240.244
R13565 gnd.n5614 gnd.n1777 240.244
R13566 gnd.n5620 gnd.n1777 240.244
R13567 gnd.n5620 gnd.n1767 240.244
R13568 gnd.n5630 gnd.n1767 240.244
R13569 gnd.n5630 gnd.n1763 240.244
R13570 gnd.n5636 gnd.n1763 240.244
R13571 gnd.n5636 gnd.n1753 240.244
R13572 gnd.n5646 gnd.n1753 240.244
R13573 gnd.n5646 gnd.n1749 240.244
R13574 gnd.n5652 gnd.n1749 240.244
R13575 gnd.n5652 gnd.n1739 240.244
R13576 gnd.n5662 gnd.n1739 240.244
R13577 gnd.n5662 gnd.n1735 240.244
R13578 gnd.n5668 gnd.n1735 240.244
R13579 gnd.n5668 gnd.n1725 240.244
R13580 gnd.n5678 gnd.n1725 240.244
R13581 gnd.n5678 gnd.n1721 240.244
R13582 gnd.n5684 gnd.n1721 240.244
R13583 gnd.n5684 gnd.n1712 240.244
R13584 gnd.n5694 gnd.n1712 240.244
R13585 gnd.n5694 gnd.n1708 240.244
R13586 gnd.n5700 gnd.n1708 240.244
R13587 gnd.n5700 gnd.n1697 240.244
R13588 gnd.n5710 gnd.n1697 240.244
R13589 gnd.n5710 gnd.n1693 240.244
R13590 gnd.n5716 gnd.n1693 240.244
R13591 gnd.n5716 gnd.n1683 240.244
R13592 gnd.n5726 gnd.n1683 240.244
R13593 gnd.n5726 gnd.n1679 240.244
R13594 gnd.n5732 gnd.n1679 240.244
R13595 gnd.n5732 gnd.n1671 240.244
R13596 gnd.n5742 gnd.n1671 240.244
R13597 gnd.n5742 gnd.n1667 240.244
R13598 gnd.n5748 gnd.n1667 240.244
R13599 gnd.n5748 gnd.n1658 240.244
R13600 gnd.n5758 gnd.n1658 240.244
R13601 gnd.n5758 gnd.n1654 240.244
R13602 gnd.n5764 gnd.n1654 240.244
R13603 gnd.n5764 gnd.n1645 240.244
R13604 gnd.n5774 gnd.n1645 240.244
R13605 gnd.n5774 gnd.n1641 240.244
R13606 gnd.n5780 gnd.n1641 240.244
R13607 gnd.n5780 gnd.n1632 240.244
R13608 gnd.n5790 gnd.n1632 240.244
R13609 gnd.n5790 gnd.n1627 240.244
R13610 gnd.n5798 gnd.n1627 240.244
R13611 gnd.n5798 gnd.n1617 240.244
R13612 gnd.n5811 gnd.n1617 240.244
R13613 gnd.n5812 gnd.n5811 240.244
R13614 gnd.n5812 gnd.n1247 240.244
R13615 gnd.n1532 gnd.n1531 240.244
R13616 gnd.n1535 gnd.n1534 240.244
R13617 gnd.n1551 gnd.n1550 240.244
R13618 gnd.n1554 gnd.n1553 240.244
R13619 gnd.n1570 gnd.n1569 240.244
R13620 gnd.n1573 gnd.n1572 240.244
R13621 gnd.n1586 gnd.n1585 240.244
R13622 gnd.n1589 gnd.n1588 240.244
R13623 gnd.n1600 gnd.n1599 240.244
R13624 gnd.n1603 gnd.n1602 240.244
R13625 gnd.n1608 gnd.n1605 240.244
R13626 gnd.n1611 gnd.n1610 240.244
R13627 gnd.n5817 gnd.n1613 240.244
R13628 gnd.n5820 gnd.n5819 240.244
R13629 gnd.n4647 gnd.n4646 240.132
R13630 gnd.n4935 gnd.n4934 240.132
R13631 gnd.n6520 gnd.n6519 225.874
R13632 gnd.n6521 gnd.n6520 225.874
R13633 gnd.n6521 gnd.n791 225.874
R13634 gnd.n6529 gnd.n791 225.874
R13635 gnd.n6530 gnd.n6529 225.874
R13636 gnd.n6531 gnd.n6530 225.874
R13637 gnd.n6531 gnd.n785 225.874
R13638 gnd.n6539 gnd.n785 225.874
R13639 gnd.n6540 gnd.n6539 225.874
R13640 gnd.n6541 gnd.n6540 225.874
R13641 gnd.n6541 gnd.n779 225.874
R13642 gnd.n6549 gnd.n779 225.874
R13643 gnd.n6550 gnd.n6549 225.874
R13644 gnd.n6551 gnd.n6550 225.874
R13645 gnd.n6551 gnd.n773 225.874
R13646 gnd.n6559 gnd.n773 225.874
R13647 gnd.n6560 gnd.n6559 225.874
R13648 gnd.n6561 gnd.n6560 225.874
R13649 gnd.n6561 gnd.n767 225.874
R13650 gnd.n6569 gnd.n767 225.874
R13651 gnd.n6570 gnd.n6569 225.874
R13652 gnd.n6571 gnd.n6570 225.874
R13653 gnd.n6571 gnd.n761 225.874
R13654 gnd.n6579 gnd.n761 225.874
R13655 gnd.n6580 gnd.n6579 225.874
R13656 gnd.n6581 gnd.n6580 225.874
R13657 gnd.n6581 gnd.n755 225.874
R13658 gnd.n6589 gnd.n755 225.874
R13659 gnd.n6590 gnd.n6589 225.874
R13660 gnd.n6591 gnd.n6590 225.874
R13661 gnd.n6591 gnd.n749 225.874
R13662 gnd.n6599 gnd.n749 225.874
R13663 gnd.n6600 gnd.n6599 225.874
R13664 gnd.n6601 gnd.n6600 225.874
R13665 gnd.n6601 gnd.n743 225.874
R13666 gnd.n6609 gnd.n743 225.874
R13667 gnd.n6610 gnd.n6609 225.874
R13668 gnd.n6611 gnd.n6610 225.874
R13669 gnd.n6611 gnd.n737 225.874
R13670 gnd.n6619 gnd.n737 225.874
R13671 gnd.n6620 gnd.n6619 225.874
R13672 gnd.n6621 gnd.n6620 225.874
R13673 gnd.n6621 gnd.n731 225.874
R13674 gnd.n6629 gnd.n731 225.874
R13675 gnd.n6630 gnd.n6629 225.874
R13676 gnd.n6631 gnd.n6630 225.874
R13677 gnd.n6631 gnd.n725 225.874
R13678 gnd.n6639 gnd.n725 225.874
R13679 gnd.n6640 gnd.n6639 225.874
R13680 gnd.n6641 gnd.n6640 225.874
R13681 gnd.n6641 gnd.n719 225.874
R13682 gnd.n6649 gnd.n719 225.874
R13683 gnd.n6650 gnd.n6649 225.874
R13684 gnd.n6651 gnd.n6650 225.874
R13685 gnd.n6651 gnd.n713 225.874
R13686 gnd.n6659 gnd.n713 225.874
R13687 gnd.n6660 gnd.n6659 225.874
R13688 gnd.n6661 gnd.n6660 225.874
R13689 gnd.n6661 gnd.n707 225.874
R13690 gnd.n6669 gnd.n707 225.874
R13691 gnd.n6670 gnd.n6669 225.874
R13692 gnd.n6671 gnd.n6670 225.874
R13693 gnd.n6671 gnd.n701 225.874
R13694 gnd.n6679 gnd.n701 225.874
R13695 gnd.n6680 gnd.n6679 225.874
R13696 gnd.n6681 gnd.n6680 225.874
R13697 gnd.n6681 gnd.n695 225.874
R13698 gnd.n6689 gnd.n695 225.874
R13699 gnd.n6690 gnd.n6689 225.874
R13700 gnd.n6691 gnd.n6690 225.874
R13701 gnd.n6691 gnd.n689 225.874
R13702 gnd.n6699 gnd.n689 225.874
R13703 gnd.n6700 gnd.n6699 225.874
R13704 gnd.n6701 gnd.n6700 225.874
R13705 gnd.n6701 gnd.n683 225.874
R13706 gnd.n6709 gnd.n683 225.874
R13707 gnd.n6710 gnd.n6709 225.874
R13708 gnd.n6711 gnd.n6710 225.874
R13709 gnd.n6711 gnd.n677 225.874
R13710 gnd.n6719 gnd.n677 225.874
R13711 gnd.n6720 gnd.n6719 225.874
R13712 gnd.n6721 gnd.n6720 225.874
R13713 gnd.n6721 gnd.n671 225.874
R13714 gnd.n6729 gnd.n671 225.874
R13715 gnd.n6730 gnd.n6729 225.874
R13716 gnd.n6731 gnd.n6730 225.874
R13717 gnd.n6731 gnd.n665 225.874
R13718 gnd.n6739 gnd.n665 225.874
R13719 gnd.n6740 gnd.n6739 225.874
R13720 gnd.n6741 gnd.n6740 225.874
R13721 gnd.n6741 gnd.n659 225.874
R13722 gnd.n6749 gnd.n659 225.874
R13723 gnd.n6750 gnd.n6749 225.874
R13724 gnd.n6751 gnd.n6750 225.874
R13725 gnd.n6751 gnd.n653 225.874
R13726 gnd.n6759 gnd.n653 225.874
R13727 gnd.n6760 gnd.n6759 225.874
R13728 gnd.n6761 gnd.n6760 225.874
R13729 gnd.n6761 gnd.n647 225.874
R13730 gnd.n6769 gnd.n647 225.874
R13731 gnd.n6770 gnd.n6769 225.874
R13732 gnd.n6771 gnd.n6770 225.874
R13733 gnd.n6771 gnd.n641 225.874
R13734 gnd.n6779 gnd.n641 225.874
R13735 gnd.n6780 gnd.n6779 225.874
R13736 gnd.n6781 gnd.n6780 225.874
R13737 gnd.n6781 gnd.n635 225.874
R13738 gnd.n6789 gnd.n635 225.874
R13739 gnd.n6790 gnd.n6789 225.874
R13740 gnd.n6791 gnd.n6790 225.874
R13741 gnd.n6791 gnd.n629 225.874
R13742 gnd.n6799 gnd.n629 225.874
R13743 gnd.n6800 gnd.n6799 225.874
R13744 gnd.n6801 gnd.n6800 225.874
R13745 gnd.n6801 gnd.n623 225.874
R13746 gnd.n6809 gnd.n623 225.874
R13747 gnd.n6810 gnd.n6809 225.874
R13748 gnd.n6811 gnd.n6810 225.874
R13749 gnd.n6811 gnd.n617 225.874
R13750 gnd.n6819 gnd.n617 225.874
R13751 gnd.n6820 gnd.n6819 225.874
R13752 gnd.n6821 gnd.n6820 225.874
R13753 gnd.n6821 gnd.n611 225.874
R13754 gnd.n6829 gnd.n611 225.874
R13755 gnd.n6830 gnd.n6829 225.874
R13756 gnd.n6831 gnd.n6830 225.874
R13757 gnd.n6831 gnd.n605 225.874
R13758 gnd.n6839 gnd.n605 225.874
R13759 gnd.n6840 gnd.n6839 225.874
R13760 gnd.n6841 gnd.n6840 225.874
R13761 gnd.n6841 gnd.n599 225.874
R13762 gnd.n6849 gnd.n599 225.874
R13763 gnd.n6850 gnd.n6849 225.874
R13764 gnd.n6851 gnd.n6850 225.874
R13765 gnd.n6851 gnd.n593 225.874
R13766 gnd.n6859 gnd.n593 225.874
R13767 gnd.n6860 gnd.n6859 225.874
R13768 gnd.n6861 gnd.n6860 225.874
R13769 gnd.n6861 gnd.n587 225.874
R13770 gnd.n6869 gnd.n587 225.874
R13771 gnd.n6870 gnd.n6869 225.874
R13772 gnd.n6871 gnd.n6870 225.874
R13773 gnd.n6871 gnd.n581 225.874
R13774 gnd.n6879 gnd.n581 225.874
R13775 gnd.n6880 gnd.n6879 225.874
R13776 gnd.n6881 gnd.n6880 225.874
R13777 gnd.n6881 gnd.n575 225.874
R13778 gnd.n6889 gnd.n575 225.874
R13779 gnd.n6890 gnd.n6889 225.874
R13780 gnd.n6891 gnd.n6890 225.874
R13781 gnd.n6891 gnd.n569 225.874
R13782 gnd.n6899 gnd.n569 225.874
R13783 gnd.n6900 gnd.n6899 225.874
R13784 gnd.n6901 gnd.n6900 225.874
R13785 gnd.n6901 gnd.n563 225.874
R13786 gnd.n6909 gnd.n563 225.874
R13787 gnd.n6910 gnd.n6909 225.874
R13788 gnd.n6911 gnd.n6910 225.874
R13789 gnd.n6911 gnd.n557 225.874
R13790 gnd.n6919 gnd.n557 225.874
R13791 gnd.n6920 gnd.n6919 225.874
R13792 gnd.n6921 gnd.n6920 225.874
R13793 gnd.n6921 gnd.n551 225.874
R13794 gnd.n6930 gnd.n551 225.874
R13795 gnd.n6931 gnd.n6930 225.874
R13796 gnd.n6932 gnd.n6931 225.874
R13797 gnd.n6932 gnd.n546 225.874
R13798 gnd.n2886 gnd.t312 224.174
R13799 gnd.n2383 gnd.t289 224.174
R13800 gnd.n1306 gnd.n1263 199.319
R13801 gnd.n1306 gnd.n1264 199.319
R13802 gnd.n2085 gnd.n2055 199.319
R13803 gnd.n2085 gnd.n2054 199.319
R13804 gnd.n6060 gnd.n1305 192.704
R13805 gnd.n5325 gnd.n5324 192.704
R13806 gnd.n4648 gnd.n4645 186.49
R13807 gnd.n4936 gnd.n4933 186.49
R13808 gnd.n3661 gnd.n3660 185
R13809 gnd.n3659 gnd.n3658 185
R13810 gnd.n3638 gnd.n3637 185
R13811 gnd.n3653 gnd.n3652 185
R13812 gnd.n3651 gnd.n3650 185
R13813 gnd.n3642 gnd.n3641 185
R13814 gnd.n3645 gnd.n3644 185
R13815 gnd.n3629 gnd.n3628 185
R13816 gnd.n3627 gnd.n3626 185
R13817 gnd.n3606 gnd.n3605 185
R13818 gnd.n3621 gnd.n3620 185
R13819 gnd.n3619 gnd.n3618 185
R13820 gnd.n3610 gnd.n3609 185
R13821 gnd.n3613 gnd.n3612 185
R13822 gnd.n3597 gnd.n3596 185
R13823 gnd.n3595 gnd.n3594 185
R13824 gnd.n3574 gnd.n3573 185
R13825 gnd.n3589 gnd.n3588 185
R13826 gnd.n3587 gnd.n3586 185
R13827 gnd.n3578 gnd.n3577 185
R13828 gnd.n3581 gnd.n3580 185
R13829 gnd.n3566 gnd.n3565 185
R13830 gnd.n3564 gnd.n3563 185
R13831 gnd.n3543 gnd.n3542 185
R13832 gnd.n3558 gnd.n3557 185
R13833 gnd.n3556 gnd.n3555 185
R13834 gnd.n3547 gnd.n3546 185
R13835 gnd.n3550 gnd.n3549 185
R13836 gnd.n3534 gnd.n3533 185
R13837 gnd.n3532 gnd.n3531 185
R13838 gnd.n3511 gnd.n3510 185
R13839 gnd.n3526 gnd.n3525 185
R13840 gnd.n3524 gnd.n3523 185
R13841 gnd.n3515 gnd.n3514 185
R13842 gnd.n3518 gnd.n3517 185
R13843 gnd.n3502 gnd.n3501 185
R13844 gnd.n3500 gnd.n3499 185
R13845 gnd.n3479 gnd.n3478 185
R13846 gnd.n3494 gnd.n3493 185
R13847 gnd.n3492 gnd.n3491 185
R13848 gnd.n3483 gnd.n3482 185
R13849 gnd.n3486 gnd.n3485 185
R13850 gnd.n3470 gnd.n3469 185
R13851 gnd.n3468 gnd.n3467 185
R13852 gnd.n3447 gnd.n3446 185
R13853 gnd.n3462 gnd.n3461 185
R13854 gnd.n3460 gnd.n3459 185
R13855 gnd.n3451 gnd.n3450 185
R13856 gnd.n3454 gnd.n3453 185
R13857 gnd.n3439 gnd.n3438 185
R13858 gnd.n3437 gnd.n3436 185
R13859 gnd.n3416 gnd.n3415 185
R13860 gnd.n3431 gnd.n3430 185
R13861 gnd.n3429 gnd.n3428 185
R13862 gnd.n3420 gnd.n3419 185
R13863 gnd.n3423 gnd.n3422 185
R13864 gnd.n2887 gnd.t311 178.987
R13865 gnd.n2384 gnd.t290 178.987
R13866 gnd.n1 gnd.t351 170.774
R13867 gnd.n9 gnd.t237 170.103
R13868 gnd.n8 gnd.t78 170.103
R13869 gnd.n7 gnd.t204 170.103
R13870 gnd.n6 gnd.t353 170.103
R13871 gnd.n5 gnd.t94 170.103
R13872 gnd.n4 gnd.t125 170.103
R13873 gnd.n3 gnd.t192 170.103
R13874 gnd.n2 gnd.t25 170.103
R13875 gnd.n1 gnd.t80 170.103
R13876 gnd.n4955 gnd.n4953 163.367
R13877 gnd.n4959 gnd.n4921 163.367
R13878 gnd.n4963 gnd.n4961 163.367
R13879 gnd.n4967 gnd.n4919 163.367
R13880 gnd.n4971 gnd.n4969 163.367
R13881 gnd.n4975 gnd.n4917 163.367
R13882 gnd.n4979 gnd.n4977 163.367
R13883 gnd.n4983 gnd.n4915 163.367
R13884 gnd.n4987 gnd.n4985 163.367
R13885 gnd.n4991 gnd.n4913 163.367
R13886 gnd.n4995 gnd.n4993 163.367
R13887 gnd.n4999 gnd.n4911 163.367
R13888 gnd.n5003 gnd.n5001 163.367
R13889 gnd.n5010 gnd.n4909 163.367
R13890 gnd.n5013 gnd.n5012 163.367
R13891 gnd.n5017 gnd.n5016 163.367
R13892 gnd.n5022 gnd.n5020 163.367
R13893 gnd.n5026 gnd.n5024 163.367
R13894 gnd.n5031 gnd.n4903 163.367
R13895 gnd.n5035 gnd.n5033 163.367
R13896 gnd.n5039 gnd.n4901 163.367
R13897 gnd.n5043 gnd.n5041 163.367
R13898 gnd.n5047 gnd.n4899 163.367
R13899 gnd.n5051 gnd.n5049 163.367
R13900 gnd.n5055 gnd.n4897 163.367
R13901 gnd.n5059 gnd.n5057 163.367
R13902 gnd.n5063 gnd.n4895 163.367
R13903 gnd.n5067 gnd.n5065 163.367
R13904 gnd.n5071 gnd.n4893 163.367
R13905 gnd.n5075 gnd.n5073 163.367
R13906 gnd.n5079 gnd.n4891 163.367
R13907 gnd.n5082 gnd.n5081 163.367
R13908 gnd.n4731 gnd.n4664 163.367
R13909 gnd.n5249 gnd.n4664 163.367
R13910 gnd.n5249 gnd.n4665 163.367
R13911 gnd.n5245 gnd.n4665 163.367
R13912 gnd.n5245 gnd.n5244 163.367
R13913 gnd.n5244 gnd.n4735 163.367
R13914 gnd.n4744 gnd.n4735 163.367
R13915 gnd.n5235 gnd.n4744 163.367
R13916 gnd.n5235 gnd.n4745 163.367
R13917 gnd.n5231 gnd.n4745 163.367
R13918 gnd.n5231 gnd.n4749 163.367
R13919 gnd.n4766 gnd.n4749 163.367
R13920 gnd.n4766 gnd.n4756 163.367
R13921 gnd.n4757 gnd.n4756 163.367
R13922 gnd.n4758 gnd.n4757 163.367
R13923 gnd.n4771 gnd.n4758 163.367
R13924 gnd.n4771 gnd.n4764 163.367
R13925 gnd.n5212 gnd.n4764 163.367
R13926 gnd.n5212 gnd.n4765 163.367
R13927 gnd.n5208 gnd.n4765 163.367
R13928 gnd.n5208 gnd.n4775 163.367
R13929 gnd.n4790 gnd.n4775 163.367
R13930 gnd.n4791 gnd.n4790 163.367
R13931 gnd.n4791 gnd.n4788 163.367
R13932 gnd.n4797 gnd.n4788 163.367
R13933 gnd.n4798 gnd.n4797 163.367
R13934 gnd.n4799 gnd.n4798 163.367
R13935 gnd.n4799 gnd.n4785 163.367
R13936 gnd.n5190 gnd.n4785 163.367
R13937 gnd.n5190 gnd.n4786 163.367
R13938 gnd.n5186 gnd.n4786 163.367
R13939 gnd.n5186 gnd.n4803 163.367
R13940 gnd.n4812 gnd.n4803 163.367
R13941 gnd.n5176 gnd.n4812 163.367
R13942 gnd.n5176 gnd.n4813 163.367
R13943 gnd.n5172 gnd.n4813 163.367
R13944 gnd.n5172 gnd.n5171 163.367
R13945 gnd.n5171 gnd.n4816 163.367
R13946 gnd.n4825 gnd.n4816 163.367
R13947 gnd.n5161 gnd.n4825 163.367
R13948 gnd.n5161 gnd.n4826 163.367
R13949 gnd.n5157 gnd.n4826 163.367
R13950 gnd.n5157 gnd.n5156 163.367
R13951 gnd.n5156 gnd.n4830 163.367
R13952 gnd.n4838 gnd.n4830 163.367
R13953 gnd.n5146 gnd.n4838 163.367
R13954 gnd.n5146 gnd.n4839 163.367
R13955 gnd.n5142 gnd.n4839 163.367
R13956 gnd.n5142 gnd.n4843 163.367
R13957 gnd.n5134 gnd.n4843 163.367
R13958 gnd.n5134 gnd.n4850 163.367
R13959 gnd.n5130 gnd.n4850 163.367
R13960 gnd.n5130 gnd.n4852 163.367
R13961 gnd.n4858 gnd.n4852 163.367
R13962 gnd.n5121 gnd.n4858 163.367
R13963 gnd.n5121 gnd.n4859 163.367
R13964 gnd.n5117 gnd.n4859 163.367
R13965 gnd.n5117 gnd.n5116 163.367
R13966 gnd.n5116 gnd.n4862 163.367
R13967 gnd.n4870 gnd.n4862 163.367
R13968 gnd.n5106 gnd.n4870 163.367
R13969 gnd.n5106 gnd.n4871 163.367
R13970 gnd.n5102 gnd.n4871 163.367
R13971 gnd.n5102 gnd.n4875 163.367
R13972 gnd.n4885 gnd.n4875 163.367
R13973 gnd.n4885 gnd.n4883 163.367
R13974 gnd.n5091 gnd.n4883 163.367
R13975 gnd.n5091 gnd.n4884 163.367
R13976 gnd.n5087 gnd.n4884 163.367
R13977 gnd.n5087 gnd.n5086 163.367
R13978 gnd.n4639 gnd.n4638 163.367
R13979 gnd.n5314 gnd.n4638 163.367
R13980 gnd.n5312 gnd.n5311 163.367
R13981 gnd.n5308 gnd.n5307 163.367
R13982 gnd.n5304 gnd.n5303 163.367
R13983 gnd.n5300 gnd.n5299 163.367
R13984 gnd.n5296 gnd.n5295 163.367
R13985 gnd.n5292 gnd.n5291 163.367
R13986 gnd.n5288 gnd.n5287 163.367
R13987 gnd.n5284 gnd.n5283 163.367
R13988 gnd.n5280 gnd.n5279 163.367
R13989 gnd.n5276 gnd.n5275 163.367
R13990 gnd.n5272 gnd.n5271 163.367
R13991 gnd.n5268 gnd.n5267 163.367
R13992 gnd.n5264 gnd.n5263 163.367
R13993 gnd.n5260 gnd.n5259 163.367
R13994 gnd.n5323 gnd.n4605 163.367
R13995 gnd.n4670 gnd.n4669 163.367
R13996 gnd.n4675 gnd.n4674 163.367
R13997 gnd.n4679 gnd.n4678 163.367
R13998 gnd.n4683 gnd.n4682 163.367
R13999 gnd.n4687 gnd.n4686 163.367
R14000 gnd.n4691 gnd.n4690 163.367
R14001 gnd.n4695 gnd.n4694 163.367
R14002 gnd.n4699 gnd.n4698 163.367
R14003 gnd.n4703 gnd.n4702 163.367
R14004 gnd.n4707 gnd.n4706 163.367
R14005 gnd.n4711 gnd.n4710 163.367
R14006 gnd.n4715 gnd.n4714 163.367
R14007 gnd.n4719 gnd.n4718 163.367
R14008 gnd.n4723 gnd.n4722 163.367
R14009 gnd.n4727 gnd.n4726 163.367
R14010 gnd.n5252 gnd.n4640 163.367
R14011 gnd.n5252 gnd.n5251 163.367
R14012 gnd.n5251 gnd.n4662 163.367
R14013 gnd.n4737 gnd.n4662 163.367
R14014 gnd.n5242 gnd.n4737 163.367
R14015 gnd.n5242 gnd.n4738 163.367
R14016 gnd.n5238 gnd.n4738 163.367
R14017 gnd.n5238 gnd.n5237 163.367
R14018 gnd.n5237 gnd.n4742 163.367
R14019 gnd.n5229 gnd.n4742 163.367
R14020 gnd.n5229 gnd.n4752 163.367
R14021 gnd.n5225 gnd.n4752 163.367
R14022 gnd.n5225 gnd.n5224 163.367
R14023 gnd.n5224 gnd.n4755 163.367
R14024 gnd.n5219 gnd.n4755 163.367
R14025 gnd.n5219 gnd.n4759 163.367
R14026 gnd.n5215 gnd.n4759 163.367
R14027 gnd.n5215 gnd.n4762 163.367
R14028 gnd.n4777 gnd.n4762 163.367
R14029 gnd.n5206 gnd.n4777 163.367
R14030 gnd.n5206 gnd.n4778 163.367
R14031 gnd.n5202 gnd.n4778 163.367
R14032 gnd.n5202 gnd.n5201 163.367
R14033 gnd.n5201 gnd.n5200 163.367
R14034 gnd.n5200 gnd.n4781 163.367
R14035 gnd.n5196 gnd.n4781 163.367
R14036 gnd.n5196 gnd.n5195 163.367
R14037 gnd.n5195 gnd.n5194 163.367
R14038 gnd.n5194 gnd.n4783 163.367
R14039 gnd.n4805 gnd.n4783 163.367
R14040 gnd.n5184 gnd.n4805 163.367
R14041 gnd.n5184 gnd.n4807 163.367
R14042 gnd.n5180 gnd.n4807 163.367
R14043 gnd.n5180 gnd.n5179 163.367
R14044 gnd.n5179 gnd.n4811 163.367
R14045 gnd.n4818 gnd.n4811 163.367
R14046 gnd.n5169 gnd.n4818 163.367
R14047 gnd.n5169 gnd.n4820 163.367
R14048 gnd.n5165 gnd.n4820 163.367
R14049 gnd.n5165 gnd.n5164 163.367
R14050 gnd.n5164 gnd.n4824 163.367
R14051 gnd.n4832 gnd.n4824 163.367
R14052 gnd.n5154 gnd.n4832 163.367
R14053 gnd.n5154 gnd.n4833 163.367
R14054 gnd.n5150 gnd.n4833 163.367
R14055 gnd.n5150 gnd.n5149 163.367
R14056 gnd.n5149 gnd.n4837 163.367
R14057 gnd.n5140 gnd.n4837 163.367
R14058 gnd.n5140 gnd.n4845 163.367
R14059 gnd.n5136 gnd.n4845 163.367
R14060 gnd.n5136 gnd.n4848 163.367
R14061 gnd.n5128 gnd.n4848 163.367
R14062 gnd.n5128 gnd.n4854 163.367
R14063 gnd.n5124 gnd.n4854 163.367
R14064 gnd.n5124 gnd.n5123 163.367
R14065 gnd.n5123 gnd.n4856 163.367
R14066 gnd.n4864 gnd.n4856 163.367
R14067 gnd.n5114 gnd.n4864 163.367
R14068 gnd.n5114 gnd.n4865 163.367
R14069 gnd.n5110 gnd.n4865 163.367
R14070 gnd.n5110 gnd.n4869 163.367
R14071 gnd.n4877 gnd.n4869 163.367
R14072 gnd.n5100 gnd.n4877 163.367
R14073 gnd.n5100 gnd.n4879 163.367
R14074 gnd.n5096 gnd.n4879 163.367
R14075 gnd.n5096 gnd.n5095 163.367
R14076 gnd.n5095 gnd.n4882 163.367
R14077 gnd.n4945 gnd.n4882 163.367
R14078 gnd.n4946 gnd.n4945 163.367
R14079 gnd.n4946 gnd.n4923 163.367
R14080 gnd.n4942 gnd.n4941 156.462
R14081 gnd.n3601 gnd.n3569 153.042
R14082 gnd.n3665 gnd.n3664 152.079
R14083 gnd.n3633 gnd.n3632 152.079
R14084 gnd.n3601 gnd.n3600 152.079
R14085 gnd.n4653 gnd.n4652 152
R14086 gnd.n4654 gnd.n4643 152
R14087 gnd.n4656 gnd.n4655 152
R14088 gnd.n4658 gnd.n4641 152
R14089 gnd.n4660 gnd.n4659 152
R14090 gnd.n4940 gnd.n4924 152
R14091 gnd.n4932 gnd.n4925 152
R14092 gnd.n4931 gnd.n4930 152
R14093 gnd.n4929 gnd.n4926 152
R14094 gnd.n4927 gnd.t300 150.546
R14095 gnd.t69 gnd.n3643 147.661
R14096 gnd.t65 gnd.n3611 147.661
R14097 gnd.t67 gnd.n3579 147.661
R14098 gnd.t63 gnd.n3548 147.661
R14099 gnd.t61 gnd.n3516 147.661
R14100 gnd.t59 gnd.n3484 147.661
R14101 gnd.t57 gnd.n3452 147.661
R14102 gnd.t71 gnd.n3421 147.661
R14103 gnd.n5019 gnd.n5018 143.351
R14104 gnd.n4620 gnd.n4604 143.351
R14105 gnd.n5322 gnd.n4604 143.351
R14106 gnd.n4650 gnd.t243 130.484
R14107 gnd.n4659 gnd.t338 126.766
R14108 gnd.n4657 gnd.t280 126.766
R14109 gnd.n4643 gnd.t320 126.766
R14110 gnd.n4651 gnd.t303 126.766
R14111 gnd.n4928 gnd.t317 126.766
R14112 gnd.n4930 gnd.t277 126.766
R14113 gnd.n4939 gnd.t332 126.766
R14114 gnd.n4941 gnd.t297 126.766
R14115 gnd.n3660 gnd.n3659 104.615
R14116 gnd.n3659 gnd.n3637 104.615
R14117 gnd.n3652 gnd.n3637 104.615
R14118 gnd.n3652 gnd.n3651 104.615
R14119 gnd.n3651 gnd.n3641 104.615
R14120 gnd.n3644 gnd.n3641 104.615
R14121 gnd.n3628 gnd.n3627 104.615
R14122 gnd.n3627 gnd.n3605 104.615
R14123 gnd.n3620 gnd.n3605 104.615
R14124 gnd.n3620 gnd.n3619 104.615
R14125 gnd.n3619 gnd.n3609 104.615
R14126 gnd.n3612 gnd.n3609 104.615
R14127 gnd.n3596 gnd.n3595 104.615
R14128 gnd.n3595 gnd.n3573 104.615
R14129 gnd.n3588 gnd.n3573 104.615
R14130 gnd.n3588 gnd.n3587 104.615
R14131 gnd.n3587 gnd.n3577 104.615
R14132 gnd.n3580 gnd.n3577 104.615
R14133 gnd.n3565 gnd.n3564 104.615
R14134 gnd.n3564 gnd.n3542 104.615
R14135 gnd.n3557 gnd.n3542 104.615
R14136 gnd.n3557 gnd.n3556 104.615
R14137 gnd.n3556 gnd.n3546 104.615
R14138 gnd.n3549 gnd.n3546 104.615
R14139 gnd.n3533 gnd.n3532 104.615
R14140 gnd.n3532 gnd.n3510 104.615
R14141 gnd.n3525 gnd.n3510 104.615
R14142 gnd.n3525 gnd.n3524 104.615
R14143 gnd.n3524 gnd.n3514 104.615
R14144 gnd.n3517 gnd.n3514 104.615
R14145 gnd.n3501 gnd.n3500 104.615
R14146 gnd.n3500 gnd.n3478 104.615
R14147 gnd.n3493 gnd.n3478 104.615
R14148 gnd.n3493 gnd.n3492 104.615
R14149 gnd.n3492 gnd.n3482 104.615
R14150 gnd.n3485 gnd.n3482 104.615
R14151 gnd.n3469 gnd.n3468 104.615
R14152 gnd.n3468 gnd.n3446 104.615
R14153 gnd.n3461 gnd.n3446 104.615
R14154 gnd.n3461 gnd.n3460 104.615
R14155 gnd.n3460 gnd.n3450 104.615
R14156 gnd.n3453 gnd.n3450 104.615
R14157 gnd.n3438 gnd.n3437 104.615
R14158 gnd.n3437 gnd.n3415 104.615
R14159 gnd.n3430 gnd.n3415 104.615
R14160 gnd.n3430 gnd.n3429 104.615
R14161 gnd.n3429 gnd.n3419 104.615
R14162 gnd.n3422 gnd.n3419 104.615
R14163 gnd.n2812 gnd.t331 100.632
R14164 gnd.n2357 gnd.t272 100.632
R14165 gnd.n7594 gnd.n138 99.6594
R14166 gnd.n7592 gnd.n7591 99.6594
R14167 gnd.n7587 gnd.n145 99.6594
R14168 gnd.n7585 gnd.n7584 99.6594
R14169 gnd.n7580 gnd.n152 99.6594
R14170 gnd.n7578 gnd.n7577 99.6594
R14171 gnd.n7573 gnd.n159 99.6594
R14172 gnd.n7571 gnd.n7570 99.6594
R14173 gnd.n7563 gnd.n166 99.6594
R14174 gnd.n7561 gnd.n7560 99.6594
R14175 gnd.n7556 gnd.n173 99.6594
R14176 gnd.n7554 gnd.n7553 99.6594
R14177 gnd.n7549 gnd.n180 99.6594
R14178 gnd.n7547 gnd.n7546 99.6594
R14179 gnd.n7542 gnd.n187 99.6594
R14180 gnd.n7540 gnd.n7539 99.6594
R14181 gnd.n7535 gnd.n194 99.6594
R14182 gnd.n7533 gnd.n7532 99.6594
R14183 gnd.n199 gnd.n198 99.6594
R14184 gnd.n6091 gnd.n6090 99.6594
R14185 gnd.n6085 gnd.n1257 99.6594
R14186 gnd.n6082 gnd.n1258 99.6594
R14187 gnd.n6078 gnd.n1259 99.6594
R14188 gnd.n6074 gnd.n1260 99.6594
R14189 gnd.n6070 gnd.n1261 99.6594
R14190 gnd.n6066 gnd.n1262 99.6594
R14191 gnd.n6062 gnd.n1263 99.6594
R14192 gnd.n6057 gnd.n1265 99.6594
R14193 gnd.n6053 gnd.n1266 99.6594
R14194 gnd.n6049 gnd.n1267 99.6594
R14195 gnd.n6045 gnd.n1268 99.6594
R14196 gnd.n6041 gnd.n1269 99.6594
R14197 gnd.n6037 gnd.n1270 99.6594
R14198 gnd.n6033 gnd.n1271 99.6594
R14199 gnd.n6029 gnd.n1272 99.6594
R14200 gnd.n6025 gnd.n1273 99.6594
R14201 gnd.n1329 gnd.n1274 99.6594
R14202 gnd.n5353 gnd.n5352 99.6594
R14203 gnd.n5348 gnd.n2061 99.6594
R14204 gnd.n5344 gnd.n2060 99.6594
R14205 gnd.n5340 gnd.n2059 99.6594
R14206 gnd.n5336 gnd.n2058 99.6594
R14207 gnd.n5332 gnd.n2057 99.6594
R14208 gnd.n5328 gnd.n2056 99.6594
R14209 gnd.n4596 gnd.n2054 99.6594
R14210 gnd.n4594 gnd.n2053 99.6594
R14211 gnd.n4590 gnd.n2052 99.6594
R14212 gnd.n4586 gnd.n2051 99.6594
R14213 gnd.n4582 gnd.n2050 99.6594
R14214 gnd.n4578 gnd.n2049 99.6594
R14215 gnd.n4574 gnd.n2048 99.6594
R14216 gnd.n4570 gnd.n2047 99.6594
R14217 gnd.n4566 gnd.n2046 99.6594
R14218 gnd.n4562 gnd.n2045 99.6594
R14219 gnd.n2103 gnd.n2044 99.6594
R14220 gnd.n4171 gnd.n3958 99.6594
R14221 gnd.n4169 gnd.n3961 99.6594
R14222 gnd.n4165 gnd.n4164 99.6594
R14223 gnd.n4158 gnd.n3966 99.6594
R14224 gnd.n4157 gnd.n4156 99.6594
R14225 gnd.n4150 gnd.n3972 99.6594
R14226 gnd.n4149 gnd.n4148 99.6594
R14227 gnd.n4142 gnd.n3978 99.6594
R14228 gnd.n4141 gnd.n4140 99.6594
R14229 gnd.n4134 gnd.n3984 99.6594
R14230 gnd.n4133 gnd.n4132 99.6594
R14231 gnd.n4126 gnd.n3993 99.6594
R14232 gnd.n4125 gnd.n4124 99.6594
R14233 gnd.n4118 gnd.n3999 99.6594
R14234 gnd.n4117 gnd.n4116 99.6594
R14235 gnd.n4110 gnd.n4005 99.6594
R14236 gnd.n4109 gnd.n4108 99.6594
R14237 gnd.n4015 gnd.n4011 99.6594
R14238 gnd.n4098 gnd.n4097 99.6594
R14239 gnd.n3783 gnd.n2340 99.6594
R14240 gnd.n3781 gnd.n2339 99.6594
R14241 gnd.n3777 gnd.n2338 99.6594
R14242 gnd.n3773 gnd.n2337 99.6594
R14243 gnd.n3769 gnd.n2336 99.6594
R14244 gnd.n3765 gnd.n2335 99.6594
R14245 gnd.n3761 gnd.n2334 99.6594
R14246 gnd.n3693 gnd.n2333 99.6594
R14247 gnd.n3024 gnd.n2755 99.6594
R14248 gnd.n2781 gnd.n2762 99.6594
R14249 gnd.n2783 gnd.n2763 99.6594
R14250 gnd.n2791 gnd.n2764 99.6594
R14251 gnd.n2793 gnd.n2765 99.6594
R14252 gnd.n2801 gnd.n2766 99.6594
R14253 gnd.n2803 gnd.n2767 99.6594
R14254 gnd.n2811 gnd.n2768 99.6594
R14255 gnd.n3751 gnd.n2320 99.6594
R14256 gnd.n3747 gnd.n2321 99.6594
R14257 gnd.n3743 gnd.n2322 99.6594
R14258 gnd.n3739 gnd.n2323 99.6594
R14259 gnd.n3735 gnd.n2324 99.6594
R14260 gnd.n3731 gnd.n2325 99.6594
R14261 gnd.n3727 gnd.n2326 99.6594
R14262 gnd.n3723 gnd.n2327 99.6594
R14263 gnd.n3719 gnd.n2328 99.6594
R14264 gnd.n3715 gnd.n2329 99.6594
R14265 gnd.n3711 gnd.n2330 99.6594
R14266 gnd.n3707 gnd.n2331 99.6594
R14267 gnd.n3703 gnd.n2332 99.6594
R14268 gnd.n2939 gnd.n2938 99.6594
R14269 gnd.n2933 gnd.n2850 99.6594
R14270 gnd.n2930 gnd.n2851 99.6594
R14271 gnd.n2926 gnd.n2852 99.6594
R14272 gnd.n2922 gnd.n2853 99.6594
R14273 gnd.n2918 gnd.n2854 99.6594
R14274 gnd.n2914 gnd.n2855 99.6594
R14275 gnd.n2910 gnd.n2856 99.6594
R14276 gnd.n2906 gnd.n2857 99.6594
R14277 gnd.n2902 gnd.n2858 99.6594
R14278 gnd.n2898 gnd.n2859 99.6594
R14279 gnd.n2894 gnd.n2860 99.6594
R14280 gnd.n2941 gnd.n2849 99.6594
R14281 gnd.n7449 gnd.n7448 99.6594
R14282 gnd.n7454 gnd.n7453 99.6594
R14283 gnd.n7457 gnd.n7456 99.6594
R14284 gnd.n7462 gnd.n7461 99.6594
R14285 gnd.n7465 gnd.n7464 99.6594
R14286 gnd.n7470 gnd.n7469 99.6594
R14287 gnd.n7473 gnd.n7472 99.6594
R14288 gnd.n7478 gnd.n7476 99.6594
R14289 gnd.n7604 gnd.n125 99.6594
R14290 gnd.n1339 gnd.n1275 99.6594
R14291 gnd.n1523 gnd.n1276 99.6594
R14292 gnd.n1525 gnd.n1277 99.6594
R14293 gnd.n1542 gnd.n1278 99.6594
R14294 gnd.n1544 gnd.n1279 99.6594
R14295 gnd.n1561 gnd.n1280 99.6594
R14296 gnd.n1563 gnd.n1281 99.6594
R14297 gnd.n1579 gnd.n1282 99.6594
R14298 gnd.n1490 gnd.n1283 99.6594
R14299 gnd.n2031 gnd.n2030 99.6594
R14300 gnd.n2032 gnd.n1980 99.6594
R14301 gnd.n2034 gnd.n1988 99.6594
R14302 gnd.n2036 gnd.n2035 99.6594
R14303 gnd.n2037 gnd.n1997 99.6594
R14304 gnd.n2039 gnd.n2006 99.6594
R14305 gnd.n2041 gnd.n2040 99.6594
R14306 gnd.n2042 gnd.n2015 99.6594
R14307 gnd.n5356 gnd.n5355 99.6594
R14308 gnd.n3818 gnd.n2318 99.6594
R14309 gnd.n3821 gnd.n3820 99.6594
R14310 gnd.n3828 gnd.n3827 99.6594
R14311 gnd.n3831 gnd.n3830 99.6594
R14312 gnd.n3838 gnd.n3837 99.6594
R14313 gnd.n3841 gnd.n3840 99.6594
R14314 gnd.n3848 gnd.n3847 99.6594
R14315 gnd.n3851 gnd.n3850 99.6594
R14316 gnd.n3858 gnd.n3857 99.6594
R14317 gnd.n3819 gnd.n3818 99.6594
R14318 gnd.n3820 gnd.n3813 99.6594
R14319 gnd.n3829 gnd.n3828 99.6594
R14320 gnd.n3830 gnd.n3809 99.6594
R14321 gnd.n3839 gnd.n3838 99.6594
R14322 gnd.n3840 gnd.n3805 99.6594
R14323 gnd.n3849 gnd.n3848 99.6594
R14324 gnd.n3850 gnd.n3801 99.6594
R14325 gnd.n3859 gnd.n3858 99.6594
R14326 gnd.n5355 gnd.n2026 99.6594
R14327 gnd.n2042 gnd.n2014 99.6594
R14328 gnd.n2041 gnd.n2007 99.6594
R14329 gnd.n2039 gnd.n2038 99.6594
R14330 gnd.n2037 gnd.n1996 99.6594
R14331 gnd.n2036 gnd.n1989 99.6594
R14332 gnd.n2034 gnd.n2033 99.6594
R14333 gnd.n2032 gnd.n1979 99.6594
R14334 gnd.n2031 gnd.n2029 99.6594
R14335 gnd.n1522 gnd.n1275 99.6594
R14336 gnd.n1526 gnd.n1276 99.6594
R14337 gnd.n1541 gnd.n1277 99.6594
R14338 gnd.n1545 gnd.n1278 99.6594
R14339 gnd.n1560 gnd.n1279 99.6594
R14340 gnd.n1564 gnd.n1280 99.6594
R14341 gnd.n1578 gnd.n1281 99.6594
R14342 gnd.n1489 gnd.n1282 99.6594
R14343 gnd.n1485 gnd.n1283 99.6594
R14344 gnd.n7477 gnd.n125 99.6594
R14345 gnd.n7476 gnd.n7475 99.6594
R14346 gnd.n7472 gnd.n7471 99.6594
R14347 gnd.n7469 gnd.n7468 99.6594
R14348 gnd.n7464 gnd.n7463 99.6594
R14349 gnd.n7461 gnd.n7460 99.6594
R14350 gnd.n7456 gnd.n7455 99.6594
R14351 gnd.n7453 gnd.n7452 99.6594
R14352 gnd.n7448 gnd.n7447 99.6594
R14353 gnd.n2939 gnd.n2862 99.6594
R14354 gnd.n2931 gnd.n2850 99.6594
R14355 gnd.n2927 gnd.n2851 99.6594
R14356 gnd.n2923 gnd.n2852 99.6594
R14357 gnd.n2919 gnd.n2853 99.6594
R14358 gnd.n2915 gnd.n2854 99.6594
R14359 gnd.n2911 gnd.n2855 99.6594
R14360 gnd.n2907 gnd.n2856 99.6594
R14361 gnd.n2903 gnd.n2857 99.6594
R14362 gnd.n2899 gnd.n2858 99.6594
R14363 gnd.n2895 gnd.n2859 99.6594
R14364 gnd.n2891 gnd.n2860 99.6594
R14365 gnd.n2942 gnd.n2941 99.6594
R14366 gnd.n3706 gnd.n2332 99.6594
R14367 gnd.n3710 gnd.n2331 99.6594
R14368 gnd.n3714 gnd.n2330 99.6594
R14369 gnd.n3718 gnd.n2329 99.6594
R14370 gnd.n3722 gnd.n2328 99.6594
R14371 gnd.n3726 gnd.n2327 99.6594
R14372 gnd.n3730 gnd.n2326 99.6594
R14373 gnd.n3734 gnd.n2325 99.6594
R14374 gnd.n3738 gnd.n2324 99.6594
R14375 gnd.n3742 gnd.n2323 99.6594
R14376 gnd.n3746 gnd.n2322 99.6594
R14377 gnd.n3750 gnd.n2321 99.6594
R14378 gnd.n2361 gnd.n2320 99.6594
R14379 gnd.n3025 gnd.n3024 99.6594
R14380 gnd.n2784 gnd.n2762 99.6594
R14381 gnd.n2790 gnd.n2763 99.6594
R14382 gnd.n2794 gnd.n2764 99.6594
R14383 gnd.n2800 gnd.n2765 99.6594
R14384 gnd.n2804 gnd.n2766 99.6594
R14385 gnd.n2810 gnd.n2767 99.6594
R14386 gnd.n2768 gnd.n2752 99.6594
R14387 gnd.n3760 gnd.n2333 99.6594
R14388 gnd.n3764 gnd.n2334 99.6594
R14389 gnd.n3768 gnd.n2335 99.6594
R14390 gnd.n3772 gnd.n2336 99.6594
R14391 gnd.n3776 gnd.n2337 99.6594
R14392 gnd.n3780 gnd.n2338 99.6594
R14393 gnd.n3784 gnd.n2339 99.6594
R14394 gnd.n2342 gnd.n2340 99.6594
R14395 gnd.n4172 gnd.n4171 99.6594
R14396 gnd.n4166 gnd.n3961 99.6594
R14397 gnd.n4164 gnd.n4163 99.6594
R14398 gnd.n4159 gnd.n4158 99.6594
R14399 gnd.n4156 gnd.n4155 99.6594
R14400 gnd.n4151 gnd.n4150 99.6594
R14401 gnd.n4148 gnd.n4147 99.6594
R14402 gnd.n4143 gnd.n4142 99.6594
R14403 gnd.n4140 gnd.n4139 99.6594
R14404 gnd.n4135 gnd.n4134 99.6594
R14405 gnd.n4132 gnd.n4131 99.6594
R14406 gnd.n4127 gnd.n4126 99.6594
R14407 gnd.n4124 gnd.n4123 99.6594
R14408 gnd.n4119 gnd.n4118 99.6594
R14409 gnd.n4116 gnd.n4115 99.6594
R14410 gnd.n4111 gnd.n4110 99.6594
R14411 gnd.n4108 gnd.n4107 99.6594
R14412 gnd.n4016 gnd.n4015 99.6594
R14413 gnd.n4099 gnd.n4098 99.6594
R14414 gnd.n4561 gnd.n2044 99.6594
R14415 gnd.n4565 gnd.n2045 99.6594
R14416 gnd.n4569 gnd.n2046 99.6594
R14417 gnd.n4573 gnd.n2047 99.6594
R14418 gnd.n4577 gnd.n2048 99.6594
R14419 gnd.n4581 gnd.n2049 99.6594
R14420 gnd.n4585 gnd.n2050 99.6594
R14421 gnd.n4589 gnd.n2051 99.6594
R14422 gnd.n4593 gnd.n2052 99.6594
R14423 gnd.n4597 gnd.n2053 99.6594
R14424 gnd.n5327 gnd.n2055 99.6594
R14425 gnd.n5331 gnd.n2056 99.6594
R14426 gnd.n5335 gnd.n2057 99.6594
R14427 gnd.n5339 gnd.n2058 99.6594
R14428 gnd.n5343 gnd.n2059 99.6594
R14429 gnd.n5347 gnd.n2060 99.6594
R14430 gnd.n2063 gnd.n2061 99.6594
R14431 gnd.n5353 gnd.n2062 99.6594
R14432 gnd.n6091 gnd.n1287 99.6594
R14433 gnd.n6083 gnd.n1257 99.6594
R14434 gnd.n6079 gnd.n1258 99.6594
R14435 gnd.n6075 gnd.n1259 99.6594
R14436 gnd.n6071 gnd.n1260 99.6594
R14437 gnd.n6067 gnd.n1261 99.6594
R14438 gnd.n6063 gnd.n1262 99.6594
R14439 gnd.n6058 gnd.n1264 99.6594
R14440 gnd.n6054 gnd.n1265 99.6594
R14441 gnd.n6050 gnd.n1266 99.6594
R14442 gnd.n6046 gnd.n1267 99.6594
R14443 gnd.n6042 gnd.n1268 99.6594
R14444 gnd.n6038 gnd.n1269 99.6594
R14445 gnd.n6034 gnd.n1270 99.6594
R14446 gnd.n6030 gnd.n1271 99.6594
R14447 gnd.n6026 gnd.n1272 99.6594
R14448 gnd.n1328 gnd.n1273 99.6594
R14449 gnd.n6018 gnd.n1274 99.6594
R14450 gnd.n198 gnd.n195 99.6594
R14451 gnd.n7534 gnd.n7533 99.6594
R14452 gnd.n194 gnd.n188 99.6594
R14453 gnd.n7541 gnd.n7540 99.6594
R14454 gnd.n187 gnd.n181 99.6594
R14455 gnd.n7548 gnd.n7547 99.6594
R14456 gnd.n180 gnd.n174 99.6594
R14457 gnd.n7555 gnd.n7554 99.6594
R14458 gnd.n173 gnd.n167 99.6594
R14459 gnd.n7562 gnd.n7561 99.6594
R14460 gnd.n166 gnd.n160 99.6594
R14461 gnd.n7572 gnd.n7571 99.6594
R14462 gnd.n159 gnd.n153 99.6594
R14463 gnd.n7579 gnd.n7578 99.6594
R14464 gnd.n152 gnd.n146 99.6594
R14465 gnd.n7586 gnd.n7585 99.6594
R14466 gnd.n145 gnd.n139 99.6594
R14467 gnd.n7593 gnd.n7592 99.6594
R14468 gnd.n138 gnd.n135 99.6594
R14469 gnd.n5403 gnd.n5402 99.6594
R14470 gnd.n1983 gnd.n1959 99.6594
R14471 gnd.n1985 gnd.n1960 99.6594
R14472 gnd.n1993 gnd.n1961 99.6594
R14473 gnd.n2001 gnd.n1962 99.6594
R14474 gnd.n2003 gnd.n1963 99.6594
R14475 gnd.n2011 gnd.n1964 99.6594
R14476 gnd.n2021 gnd.n1965 99.6594
R14477 gnd.n2023 gnd.n1966 99.6594
R14478 gnd.n4520 gnd.n1967 99.6594
R14479 gnd.n4522 gnd.n1968 99.6594
R14480 gnd.n4526 gnd.n1969 99.6594
R14481 gnd.n4532 gnd.n1970 99.6594
R14482 gnd.n5405 gnd.n1957 99.6594
R14483 gnd.n5403 gnd.n1973 99.6594
R14484 gnd.n1984 gnd.n1959 99.6594
R14485 gnd.n1992 gnd.n1960 99.6594
R14486 gnd.n2000 gnd.n1961 99.6594
R14487 gnd.n2002 gnd.n1962 99.6594
R14488 gnd.n2010 gnd.n1963 99.6594
R14489 gnd.n2020 gnd.n1964 99.6594
R14490 gnd.n2022 gnd.n1965 99.6594
R14491 gnd.n4519 gnd.n1966 99.6594
R14492 gnd.n4521 gnd.n1967 99.6594
R14493 gnd.n4525 gnd.n1968 99.6594
R14494 gnd.n4527 gnd.n1969 99.6594
R14495 gnd.n4533 gnd.n1970 99.6594
R14496 gnd.n5406 gnd.n5405 99.6594
R14497 gnd.n1531 gnd.n1513 99.6594
R14498 gnd.n1535 gnd.n1533 99.6594
R14499 gnd.n1550 gnd.n1506 99.6594
R14500 gnd.n1554 gnd.n1552 99.6594
R14501 gnd.n1569 gnd.n1499 99.6594
R14502 gnd.n1573 gnd.n1571 99.6594
R14503 gnd.n1585 gnd.n1493 99.6594
R14504 gnd.n1589 gnd.n1587 99.6594
R14505 gnd.n1599 gnd.n1481 99.6594
R14506 gnd.n1602 gnd.n1601 99.6594
R14507 gnd.n1605 gnd.n1604 99.6594
R14508 gnd.n1610 gnd.n1609 99.6594
R14509 gnd.n1613 gnd.n1612 99.6594
R14510 gnd.n5819 gnd.n5818 99.6594
R14511 gnd.n5818 gnd.n5817 99.6594
R14512 gnd.n1612 gnd.n1611 99.6594
R14513 gnd.n1609 gnd.n1608 99.6594
R14514 gnd.n1604 gnd.n1603 99.6594
R14515 gnd.n1601 gnd.n1600 99.6594
R14516 gnd.n1588 gnd.n1481 99.6594
R14517 gnd.n1587 gnd.n1586 99.6594
R14518 gnd.n1572 gnd.n1493 99.6594
R14519 gnd.n1571 gnd.n1570 99.6594
R14520 gnd.n1553 gnd.n1499 99.6594
R14521 gnd.n1552 gnd.n1551 99.6594
R14522 gnd.n1534 gnd.n1506 99.6594
R14523 gnd.n1533 gnd.n1532 99.6594
R14524 gnd.n1513 gnd.n1244 99.6594
R14525 gnd.n4528 gnd.t286 98.63
R14526 gnd.n122 gnd.t292 98.63
R14527 gnd.n1486 gnd.t308 98.63
R14528 gnd.n2016 gnd.t336 98.63
R14529 gnd.n1308 gnd.t276 98.63
R14530 gnd.n1330 gnd.t265 98.63
R14531 gnd.n201 gnd.t326 98.63
R14532 gnd.n7565 gnd.t248 98.63
R14533 gnd.n3985 gnd.t349 98.63
R14534 gnd.n4017 gnd.t316 98.63
R14535 gnd.n3798 gnd.t346 98.63
R14536 gnd.n2105 gnd.t342 98.63
R14537 gnd.n2083 gnd.t260 98.63
R14538 gnd.n5827 gnd.t256 98.63
R14539 gnd.n4666 gnd.t324 88.9408
R14540 gnd.n4904 gnd.t252 88.9408
R14541 gnd.n5256 gnd.t269 88.933
R14542 gnd.n5006 gnd.t295 88.933
R14543 gnd.n6941 gnd.n6940 84.8607
R14544 gnd.n6942 gnd.n6941 84.8607
R14545 gnd.n6942 gnd.n540 84.8607
R14546 gnd.n6950 gnd.n540 84.8607
R14547 gnd.n6951 gnd.n6950 84.8607
R14548 gnd.n6952 gnd.n6951 84.8607
R14549 gnd.n6952 gnd.n534 84.8607
R14550 gnd.n6960 gnd.n534 84.8607
R14551 gnd.n6961 gnd.n6960 84.8607
R14552 gnd.n6962 gnd.n6961 84.8607
R14553 gnd.n6962 gnd.n528 84.8607
R14554 gnd.n6970 gnd.n528 84.8607
R14555 gnd.n6971 gnd.n6970 84.8607
R14556 gnd.n6972 gnd.n6971 84.8607
R14557 gnd.n6972 gnd.n522 84.8607
R14558 gnd.n6980 gnd.n522 84.8607
R14559 gnd.n6981 gnd.n6980 84.8607
R14560 gnd.n6982 gnd.n6981 84.8607
R14561 gnd.n6982 gnd.n516 84.8607
R14562 gnd.n6990 gnd.n516 84.8607
R14563 gnd.n6991 gnd.n6990 84.8607
R14564 gnd.n6992 gnd.n6991 84.8607
R14565 gnd.n6992 gnd.n510 84.8607
R14566 gnd.n7000 gnd.n510 84.8607
R14567 gnd.n7001 gnd.n7000 84.8607
R14568 gnd.n7002 gnd.n7001 84.8607
R14569 gnd.n7002 gnd.n504 84.8607
R14570 gnd.n7010 gnd.n504 84.8607
R14571 gnd.n7011 gnd.n7010 84.8607
R14572 gnd.n7012 gnd.n7011 84.8607
R14573 gnd.n7012 gnd.n498 84.8607
R14574 gnd.n7020 gnd.n498 84.8607
R14575 gnd.n7021 gnd.n7020 84.8607
R14576 gnd.n7022 gnd.n7021 84.8607
R14577 gnd.n7022 gnd.n492 84.8607
R14578 gnd.n7030 gnd.n492 84.8607
R14579 gnd.n7031 gnd.n7030 84.8607
R14580 gnd.n7032 gnd.n7031 84.8607
R14581 gnd.n7032 gnd.n486 84.8607
R14582 gnd.n7040 gnd.n486 84.8607
R14583 gnd.n7041 gnd.n7040 84.8607
R14584 gnd.n7042 gnd.n7041 84.8607
R14585 gnd.n7042 gnd.n480 84.8607
R14586 gnd.n7050 gnd.n480 84.8607
R14587 gnd.n7051 gnd.n7050 84.8607
R14588 gnd.n7052 gnd.n7051 84.8607
R14589 gnd.n7052 gnd.n474 84.8607
R14590 gnd.n7060 gnd.n474 84.8607
R14591 gnd.n7061 gnd.n7060 84.8607
R14592 gnd.n7062 gnd.n7061 84.8607
R14593 gnd.n7062 gnd.n468 84.8607
R14594 gnd.n7070 gnd.n468 84.8607
R14595 gnd.n7071 gnd.n7070 84.8607
R14596 gnd.n7072 gnd.n7071 84.8607
R14597 gnd.n7072 gnd.n462 84.8607
R14598 gnd.n7080 gnd.n462 84.8607
R14599 gnd.n7081 gnd.n7080 84.8607
R14600 gnd.n7082 gnd.n7081 84.8607
R14601 gnd.n7082 gnd.n456 84.8607
R14602 gnd.n7090 gnd.n456 84.8607
R14603 gnd.n7091 gnd.n7090 84.8607
R14604 gnd.n7092 gnd.n7091 84.8607
R14605 gnd.n7092 gnd.n450 84.8607
R14606 gnd.n7100 gnd.n450 84.8607
R14607 gnd.n7101 gnd.n7100 84.8607
R14608 gnd.n7102 gnd.n7101 84.8607
R14609 gnd.n7102 gnd.n444 84.8607
R14610 gnd.n7110 gnd.n444 84.8607
R14611 gnd.n7111 gnd.n7110 84.8607
R14612 gnd.n7112 gnd.n7111 84.8607
R14613 gnd.n7112 gnd.n438 84.8607
R14614 gnd.n7120 gnd.n438 84.8607
R14615 gnd.n7121 gnd.n7120 84.8607
R14616 gnd.n7122 gnd.n7121 84.8607
R14617 gnd.n7122 gnd.n432 84.8607
R14618 gnd.n7130 gnd.n432 84.8607
R14619 gnd.n7131 gnd.n7130 84.8607
R14620 gnd.n7132 gnd.n7131 84.8607
R14621 gnd.n7132 gnd.n426 84.8607
R14622 gnd.n7140 gnd.n426 84.8607
R14623 gnd.n7141 gnd.n7140 84.8607
R14624 gnd.n7143 gnd.n7141 84.8607
R14625 gnd.n7143 gnd.n7142 84.8607
R14626 gnd.n4650 gnd.n4649 81.8399
R14627 gnd.n2813 gnd.t330 74.8376
R14628 gnd.n2358 gnd.t273 74.8376
R14629 gnd.n4667 gnd.t323 72.8438
R14630 gnd.n4905 gnd.t253 72.8438
R14631 gnd.n4651 gnd.n4644 72.8411
R14632 gnd.n4657 gnd.n4642 72.8411
R14633 gnd.n4939 gnd.n4938 72.8411
R14634 gnd.n4529 gnd.t285 72.836
R14635 gnd.n5257 gnd.t268 72.836
R14636 gnd.n5007 gnd.t296 72.836
R14637 gnd.n123 gnd.t293 72.836
R14638 gnd.n1487 gnd.t307 72.836
R14639 gnd.n2017 gnd.t337 72.836
R14640 gnd.n1309 gnd.t275 72.836
R14641 gnd.n1331 gnd.t264 72.836
R14642 gnd.n202 gnd.t327 72.836
R14643 gnd.n7566 gnd.t249 72.836
R14644 gnd.n3986 gnd.t348 72.836
R14645 gnd.n4018 gnd.t315 72.836
R14646 gnd.n3799 gnd.t345 72.836
R14647 gnd.n2106 gnd.t343 72.836
R14648 gnd.n2084 gnd.t261 72.836
R14649 gnd.n5828 gnd.t257 72.836
R14650 gnd.n4953 gnd.n4952 71.676
R14651 gnd.n4954 gnd.n4921 71.676
R14652 gnd.n4961 gnd.n4960 71.676
R14653 gnd.n4962 gnd.n4919 71.676
R14654 gnd.n4969 gnd.n4968 71.676
R14655 gnd.n4970 gnd.n4917 71.676
R14656 gnd.n4977 gnd.n4976 71.676
R14657 gnd.n4978 gnd.n4915 71.676
R14658 gnd.n4985 gnd.n4984 71.676
R14659 gnd.n4986 gnd.n4913 71.676
R14660 gnd.n4993 gnd.n4992 71.676
R14661 gnd.n4994 gnd.n4911 71.676
R14662 gnd.n5001 gnd.n5000 71.676
R14663 gnd.n5002 gnd.n4909 71.676
R14664 gnd.n5012 gnd.n5011 71.676
R14665 gnd.n5016 gnd.n4907 71.676
R14666 gnd.n5020 gnd.n5019 71.676
R14667 gnd.n5024 gnd.n5023 71.676
R14668 gnd.n5025 gnd.n4903 71.676
R14669 gnd.n5033 gnd.n5032 71.676
R14670 gnd.n5034 gnd.n4901 71.676
R14671 gnd.n5041 gnd.n5040 71.676
R14672 gnd.n5042 gnd.n4899 71.676
R14673 gnd.n5049 gnd.n5048 71.676
R14674 gnd.n5050 gnd.n4897 71.676
R14675 gnd.n5057 gnd.n5056 71.676
R14676 gnd.n5058 gnd.n4895 71.676
R14677 gnd.n5065 gnd.n5064 71.676
R14678 gnd.n5066 gnd.n4893 71.676
R14679 gnd.n5073 gnd.n5072 71.676
R14680 gnd.n5074 gnd.n4891 71.676
R14681 gnd.n5081 gnd.n5080 71.676
R14682 gnd.n5085 gnd.n4889 71.676
R14683 gnd.n5320 gnd.n5319 71.676
R14684 gnd.n5314 gnd.n4606 71.676
R14685 gnd.n5311 gnd.n4607 71.676
R14686 gnd.n5307 gnd.n4608 71.676
R14687 gnd.n5303 gnd.n4609 71.676
R14688 gnd.n5299 gnd.n4610 71.676
R14689 gnd.n5295 gnd.n4611 71.676
R14690 gnd.n5291 gnd.n4612 71.676
R14691 gnd.n5287 gnd.n4613 71.676
R14692 gnd.n5283 gnd.n4614 71.676
R14693 gnd.n5279 gnd.n4615 71.676
R14694 gnd.n5275 gnd.n4616 71.676
R14695 gnd.n5271 gnd.n4617 71.676
R14696 gnd.n5267 gnd.n4618 71.676
R14697 gnd.n5263 gnd.n4619 71.676
R14698 gnd.n5259 gnd.n4620 71.676
R14699 gnd.n4621 gnd.n4605 71.676
R14700 gnd.n4670 gnd.n4622 71.676
R14701 gnd.n4675 gnd.n4623 71.676
R14702 gnd.n4679 gnd.n4624 71.676
R14703 gnd.n4683 gnd.n4625 71.676
R14704 gnd.n4687 gnd.n4626 71.676
R14705 gnd.n4691 gnd.n4627 71.676
R14706 gnd.n4695 gnd.n4628 71.676
R14707 gnd.n4699 gnd.n4629 71.676
R14708 gnd.n4703 gnd.n4630 71.676
R14709 gnd.n4707 gnd.n4631 71.676
R14710 gnd.n4711 gnd.n4632 71.676
R14711 gnd.n4715 gnd.n4633 71.676
R14712 gnd.n4719 gnd.n4634 71.676
R14713 gnd.n4723 gnd.n4635 71.676
R14714 gnd.n4727 gnd.n4636 71.676
R14715 gnd.n5320 gnd.n4639 71.676
R14716 gnd.n5312 gnd.n4606 71.676
R14717 gnd.n5308 gnd.n4607 71.676
R14718 gnd.n5304 gnd.n4608 71.676
R14719 gnd.n5300 gnd.n4609 71.676
R14720 gnd.n5296 gnd.n4610 71.676
R14721 gnd.n5292 gnd.n4611 71.676
R14722 gnd.n5288 gnd.n4612 71.676
R14723 gnd.n5284 gnd.n4613 71.676
R14724 gnd.n5280 gnd.n4614 71.676
R14725 gnd.n5276 gnd.n4615 71.676
R14726 gnd.n5272 gnd.n4616 71.676
R14727 gnd.n5268 gnd.n4617 71.676
R14728 gnd.n5264 gnd.n4618 71.676
R14729 gnd.n5260 gnd.n4619 71.676
R14730 gnd.n5323 gnd.n5322 71.676
R14731 gnd.n4669 gnd.n4621 71.676
R14732 gnd.n4674 gnd.n4622 71.676
R14733 gnd.n4678 gnd.n4623 71.676
R14734 gnd.n4682 gnd.n4624 71.676
R14735 gnd.n4686 gnd.n4625 71.676
R14736 gnd.n4690 gnd.n4626 71.676
R14737 gnd.n4694 gnd.n4627 71.676
R14738 gnd.n4698 gnd.n4628 71.676
R14739 gnd.n4702 gnd.n4629 71.676
R14740 gnd.n4706 gnd.n4630 71.676
R14741 gnd.n4710 gnd.n4631 71.676
R14742 gnd.n4714 gnd.n4632 71.676
R14743 gnd.n4718 gnd.n4633 71.676
R14744 gnd.n4722 gnd.n4634 71.676
R14745 gnd.n4726 gnd.n4635 71.676
R14746 gnd.n4730 gnd.n4636 71.676
R14747 gnd.n5082 gnd.n4889 71.676
R14748 gnd.n5080 gnd.n5079 71.676
R14749 gnd.n5075 gnd.n5074 71.676
R14750 gnd.n5072 gnd.n5071 71.676
R14751 gnd.n5067 gnd.n5066 71.676
R14752 gnd.n5064 gnd.n5063 71.676
R14753 gnd.n5059 gnd.n5058 71.676
R14754 gnd.n5056 gnd.n5055 71.676
R14755 gnd.n5051 gnd.n5050 71.676
R14756 gnd.n5048 gnd.n5047 71.676
R14757 gnd.n5043 gnd.n5042 71.676
R14758 gnd.n5040 gnd.n5039 71.676
R14759 gnd.n5035 gnd.n5034 71.676
R14760 gnd.n5032 gnd.n5031 71.676
R14761 gnd.n5026 gnd.n5025 71.676
R14762 gnd.n5023 gnd.n5022 71.676
R14763 gnd.n5018 gnd.n5017 71.676
R14764 gnd.n5013 gnd.n4907 71.676
R14765 gnd.n5011 gnd.n5010 71.676
R14766 gnd.n5003 gnd.n5002 71.676
R14767 gnd.n5000 gnd.n4999 71.676
R14768 gnd.n4995 gnd.n4994 71.676
R14769 gnd.n4992 gnd.n4991 71.676
R14770 gnd.n4987 gnd.n4986 71.676
R14771 gnd.n4984 gnd.n4983 71.676
R14772 gnd.n4979 gnd.n4978 71.676
R14773 gnd.n4976 gnd.n4975 71.676
R14774 gnd.n4971 gnd.n4970 71.676
R14775 gnd.n4968 gnd.n4967 71.676
R14776 gnd.n4963 gnd.n4962 71.676
R14777 gnd.n4960 gnd.n4959 71.676
R14778 gnd.n4955 gnd.n4954 71.676
R14779 gnd.n4952 gnd.n4951 71.676
R14780 gnd.n10 gnd.t155 69.1507
R14781 gnd.n18 gnd.t134 68.4792
R14782 gnd.n17 gnd.t104 68.4792
R14783 gnd.n16 gnd.t355 68.4792
R14784 gnd.n15 gnd.t118 68.4792
R14785 gnd.n14 gnd.t194 68.4792
R14786 gnd.n13 gnd.t235 68.4792
R14787 gnd.n12 gnd.t123 68.4792
R14788 gnd.n11 gnd.t157 68.4792
R14789 gnd.n10 gnd.t131 68.4792
R14790 gnd.n2940 gnd.n2844 64.369
R14791 gnd.n4672 gnd.n4667 59.5399
R14792 gnd.n5028 gnd.n4905 59.5399
R14793 gnd.n5258 gnd.n5257 59.5399
R14794 gnd.n5008 gnd.n5007 59.5399
R14795 gnd.n5255 gnd.n4660 59.1804
R14796 gnd.n2591 gnd.t208 56.607
R14797 gnd.n60 gnd.t75 56.607
R14798 gnd.n2552 gnd.t92 56.407
R14799 gnd.n2571 gnd.t43 56.407
R14800 gnd.n21 gnd.t144 56.407
R14801 gnd.n40 gnd.t30 56.407
R14802 gnd.n2608 gnd.t153 55.8337
R14803 gnd.n2569 gnd.t113 55.8337
R14804 gnd.n2588 gnd.t4 55.8337
R14805 gnd.n77 gnd.t74 55.8337
R14806 gnd.n38 gnd.t145 55.8337
R14807 gnd.n57 gnd.t83 55.8337
R14808 gnd.n4648 gnd.n4647 54.358
R14809 gnd.n4936 gnd.n4935 54.358
R14810 gnd.n2591 gnd.n2590 53.0052
R14811 gnd.n2593 gnd.n2592 53.0052
R14812 gnd.n2595 gnd.n2594 53.0052
R14813 gnd.n2597 gnd.n2596 53.0052
R14814 gnd.n2599 gnd.n2598 53.0052
R14815 gnd.n2601 gnd.n2600 53.0052
R14816 gnd.n2603 gnd.n2602 53.0052
R14817 gnd.n2605 gnd.n2604 53.0052
R14818 gnd.n2607 gnd.n2606 53.0052
R14819 gnd.n2552 gnd.n2551 53.0052
R14820 gnd.n2554 gnd.n2553 53.0052
R14821 gnd.n2556 gnd.n2555 53.0052
R14822 gnd.n2558 gnd.n2557 53.0052
R14823 gnd.n2560 gnd.n2559 53.0052
R14824 gnd.n2562 gnd.n2561 53.0052
R14825 gnd.n2564 gnd.n2563 53.0052
R14826 gnd.n2566 gnd.n2565 53.0052
R14827 gnd.n2568 gnd.n2567 53.0052
R14828 gnd.n2571 gnd.n2570 53.0052
R14829 gnd.n2573 gnd.n2572 53.0052
R14830 gnd.n2575 gnd.n2574 53.0052
R14831 gnd.n2577 gnd.n2576 53.0052
R14832 gnd.n2579 gnd.n2578 53.0052
R14833 gnd.n2581 gnd.n2580 53.0052
R14834 gnd.n2583 gnd.n2582 53.0052
R14835 gnd.n2585 gnd.n2584 53.0052
R14836 gnd.n2587 gnd.n2586 53.0052
R14837 gnd.n76 gnd.n75 53.0052
R14838 gnd.n74 gnd.n73 53.0052
R14839 gnd.n72 gnd.n71 53.0052
R14840 gnd.n70 gnd.n69 53.0052
R14841 gnd.n68 gnd.n67 53.0052
R14842 gnd.n66 gnd.n65 53.0052
R14843 gnd.n64 gnd.n63 53.0052
R14844 gnd.n62 gnd.n61 53.0052
R14845 gnd.n60 gnd.n59 53.0052
R14846 gnd.n37 gnd.n36 53.0052
R14847 gnd.n35 gnd.n34 53.0052
R14848 gnd.n33 gnd.n32 53.0052
R14849 gnd.n31 gnd.n30 53.0052
R14850 gnd.n29 gnd.n28 53.0052
R14851 gnd.n27 gnd.n26 53.0052
R14852 gnd.n25 gnd.n24 53.0052
R14853 gnd.n23 gnd.n22 53.0052
R14854 gnd.n21 gnd.n20 53.0052
R14855 gnd.n56 gnd.n55 53.0052
R14856 gnd.n54 gnd.n53 53.0052
R14857 gnd.n52 gnd.n51 53.0052
R14858 gnd.n50 gnd.n49 53.0052
R14859 gnd.n48 gnd.n47 53.0052
R14860 gnd.n46 gnd.n45 53.0052
R14861 gnd.n44 gnd.n43 53.0052
R14862 gnd.n42 gnd.n41 53.0052
R14863 gnd.n40 gnd.n39 53.0052
R14864 gnd.n4927 gnd.n4926 52.4801
R14865 gnd.n3644 gnd.t69 52.3082
R14866 gnd.n3612 gnd.t65 52.3082
R14867 gnd.n3580 gnd.t67 52.3082
R14868 gnd.n3549 gnd.t63 52.3082
R14869 gnd.n3517 gnd.t61 52.3082
R14870 gnd.n3485 gnd.t59 52.3082
R14871 gnd.n3453 gnd.t57 52.3082
R14872 gnd.n3422 gnd.t71 52.3082
R14873 gnd.n4179 gnd.n3793 51.6227
R14874 gnd.n7602 gnd.n128 51.6227
R14875 gnd.n3474 gnd.n3442 51.4173
R14876 gnd.n7142 gnd.n238 50.9166
R14877 gnd.n3538 gnd.n3537 50.455
R14878 gnd.n3506 gnd.n3505 50.455
R14879 gnd.n3474 gnd.n3473 50.455
R14880 gnd.n2887 gnd.n2886 45.1884
R14881 gnd.n2384 gnd.n2383 45.1884
R14882 gnd.n4949 gnd.n4942 44.3322
R14883 gnd.n4651 gnd.n4650 44.3189
R14884 gnd.n4530 gnd.n4529 42.4732
R14885 gnd.n5829 gnd.n5828 42.4732
R14886 gnd.n2888 gnd.n2887 42.2793
R14887 gnd.n2385 gnd.n2384 42.2793
R14888 gnd.n2814 gnd.n2813 42.2793
R14889 gnd.n3759 gnd.n2358 42.2793
R14890 gnd.n124 gnd.n123 42.2793
R14891 gnd.n1594 gnd.n1487 42.2793
R14892 gnd.n2018 gnd.n2017 42.2793
R14893 gnd.n1332 gnd.n1331 42.2793
R14894 gnd.n7530 gnd.n202 42.2793
R14895 gnd.n7567 gnd.n7566 42.2793
R14896 gnd.n3987 gnd.n3986 42.2793
R14897 gnd.n4019 gnd.n4018 42.2793
R14898 gnd.n3800 gnd.n3799 42.2793
R14899 gnd.n4560 gnd.n2106 42.2793
R14900 gnd.n4649 gnd.n4648 41.6274
R14901 gnd.n4937 gnd.n4936 41.6274
R14902 gnd.n4658 gnd.n4657 40.8975
R14903 gnd.n4940 gnd.n4939 40.8975
R14904 gnd.n6060 gnd.n1309 36.9518
R14905 gnd.n5325 gnd.n2084 36.9518
R14906 gnd.n4657 gnd.n4656 35.055
R14907 gnd.n4652 gnd.n4651 35.055
R14908 gnd.n4929 gnd.n4928 35.055
R14909 gnd.n4939 gnd.n4925 35.055
R14910 gnd.n6511 gnd.n797 31.9958
R14911 gnd.n6511 gnd.n6510 31.9958
R14912 gnd.n6510 gnd.n6509 31.9958
R14913 gnd.n6509 gnd.n802 31.9958
R14914 gnd.n6503 gnd.n802 31.9958
R14915 gnd.n6503 gnd.n6502 31.9958
R14916 gnd.n6502 gnd.n6501 31.9958
R14917 gnd.n6501 gnd.n810 31.9958
R14918 gnd.n6495 gnd.n810 31.9958
R14919 gnd.n6495 gnd.n6494 31.9958
R14920 gnd.n6494 gnd.n6493 31.9958
R14921 gnd.n6493 gnd.n818 31.9958
R14922 gnd.n6487 gnd.n818 31.9958
R14923 gnd.n6487 gnd.n6486 31.9958
R14924 gnd.n6486 gnd.n6485 31.9958
R14925 gnd.n6485 gnd.n826 31.9958
R14926 gnd.n6479 gnd.n826 31.9958
R14927 gnd.n6479 gnd.n6478 31.9958
R14928 gnd.n6478 gnd.n6477 31.9958
R14929 gnd.n6477 gnd.n834 31.9958
R14930 gnd.n6471 gnd.n834 31.9958
R14931 gnd.n6471 gnd.n6470 31.9958
R14932 gnd.n6470 gnd.n6469 31.9958
R14933 gnd.n6469 gnd.n842 31.9958
R14934 gnd.n6463 gnd.n842 31.9958
R14935 gnd.n6463 gnd.n6462 31.9958
R14936 gnd.n6462 gnd.n6461 31.9958
R14937 gnd.n6461 gnd.n850 31.9958
R14938 gnd.n6455 gnd.n850 31.9958
R14939 gnd.n6455 gnd.n6454 31.9958
R14940 gnd.n6454 gnd.n6453 31.9958
R14941 gnd.n6453 gnd.n858 31.9958
R14942 gnd.n6447 gnd.n858 31.9958
R14943 gnd.n6447 gnd.n6446 31.9958
R14944 gnd.n6446 gnd.n6445 31.9958
R14945 gnd.n6445 gnd.n866 31.9958
R14946 gnd.n6439 gnd.n866 31.9958
R14947 gnd.n6439 gnd.n6438 31.9958
R14948 gnd.n6438 gnd.n6437 31.9958
R14949 gnd.n6437 gnd.n874 31.9958
R14950 gnd.n6431 gnd.n874 31.9958
R14951 gnd.n6431 gnd.n6430 31.9958
R14952 gnd.n6430 gnd.n6429 31.9958
R14953 gnd.n6429 gnd.n882 31.9958
R14954 gnd.n6423 gnd.n882 31.9958
R14955 gnd.n6423 gnd.n6422 31.9958
R14956 gnd.n6422 gnd.n6421 31.9958
R14957 gnd.n6421 gnd.n890 31.9958
R14958 gnd.n6415 gnd.n890 31.9958
R14959 gnd.n6415 gnd.n6414 31.9958
R14960 gnd.n6414 gnd.n6413 31.9958
R14961 gnd.n6413 gnd.n898 31.9958
R14962 gnd.n6407 gnd.n898 31.9958
R14963 gnd.n6407 gnd.n6406 31.9958
R14964 gnd.n6406 gnd.n6405 31.9958
R14965 gnd.n6405 gnd.n906 31.9958
R14966 gnd.n6399 gnd.n906 31.9958
R14967 gnd.n6399 gnd.n6398 31.9958
R14968 gnd.n6398 gnd.n6397 31.9958
R14969 gnd.n6397 gnd.n914 31.9958
R14970 gnd.n6391 gnd.n914 31.9958
R14971 gnd.n6391 gnd.n6390 31.9958
R14972 gnd.n6390 gnd.n6389 31.9958
R14973 gnd.n6389 gnd.n922 31.9958
R14974 gnd.n6383 gnd.n922 31.9958
R14975 gnd.n6383 gnd.n6382 31.9958
R14976 gnd.n6382 gnd.n6381 31.9958
R14977 gnd.n6381 gnd.n930 31.9958
R14978 gnd.n6375 gnd.n930 31.9958
R14979 gnd.n6375 gnd.n6374 31.9958
R14980 gnd.n6374 gnd.n6373 31.9958
R14981 gnd.n6373 gnd.n938 31.9958
R14982 gnd.n6367 gnd.n938 31.9958
R14983 gnd.n6367 gnd.n6366 31.9958
R14984 gnd.n6366 gnd.n6365 31.9958
R14985 gnd.n6365 gnd.n946 31.9958
R14986 gnd.n6359 gnd.n946 31.9958
R14987 gnd.n6359 gnd.n6358 31.9958
R14988 gnd.n6358 gnd.n6357 31.9958
R14989 gnd.n6357 gnd.n954 31.9958
R14990 gnd.n6351 gnd.n954 31.9958
R14991 gnd.n6351 gnd.n6350 31.9958
R14992 gnd.n6350 gnd.n6349 31.9958
R14993 gnd.n2950 gnd.n2844 31.8661
R14994 gnd.n2950 gnd.n2949 31.8661
R14995 gnd.n2958 gnd.n2833 31.8661
R14996 gnd.n2966 gnd.n2833 31.8661
R14997 gnd.n2966 gnd.n2827 31.8661
R14998 gnd.n2974 gnd.n2827 31.8661
R14999 gnd.n2974 gnd.n2820 31.8661
R15000 gnd.n3012 gnd.n2820 31.8661
R15001 gnd.n3022 gnd.n2753 31.8661
R15002 gnd.n4179 gnd.n3957 31.8661
R15003 gnd.n4187 gnd.n2305 31.8661
R15004 gnd.n4195 gnd.n2305 31.8661
R15005 gnd.n4195 gnd.n2297 31.8661
R15006 gnd.n4203 gnd.n2297 31.8661
R15007 gnd.n4211 gnd.n2288 31.8661
R15008 gnd.n4211 gnd.n2291 31.8661
R15009 gnd.n4219 gnd.n2273 31.8661
R15010 gnd.n4227 gnd.n2273 31.8661
R15011 gnd.n4235 gnd.n2265 31.8661
R15012 gnd.n4243 gnd.n2256 31.8661
R15013 gnd.n4243 gnd.n2259 31.8661
R15014 gnd.n4251 gnd.n2241 31.8661
R15015 gnd.n4259 gnd.n2241 31.8661
R15016 gnd.n4267 gnd.n2233 31.8661
R15017 gnd.n4276 gnd.n2224 31.8661
R15018 gnd.n4276 gnd.n2227 31.8661
R15019 gnd.n4284 gnd.n2210 31.8661
R15020 gnd.n4292 gnd.n2210 31.8661
R15021 gnd.n4301 gnd.n2201 31.8661
R15022 gnd.n4309 gnd.n2194 31.8661
R15023 gnd.n4309 gnd.n2196 31.8661
R15024 gnd.n4328 gnd.n2178 31.8661
R15025 gnd.n4335 gnd.n970 31.8661
R15026 gnd.n2027 gnd.n1112 31.8661
R15027 gnd.n4477 gnd.n2043 31.8661
R15028 gnd.n4477 gnd.n1958 31.8661
R15029 gnd.n1971 gnd.n1952 31.8661
R15030 gnd.n5413 gnd.n1952 31.8661
R15031 gnd.n5421 gnd.n1945 31.8661
R15032 gnd.n5421 gnd.n1938 31.8661
R15033 gnd.n5429 gnd.n1938 31.8661
R15034 gnd.n5429 gnd.n1939 31.8661
R15035 gnd.n5437 gnd.n1926 31.8661
R15036 gnd.n5445 gnd.n1926 31.8661
R15037 gnd.n5445 gnd.n1919 31.8661
R15038 gnd.n5453 gnd.n1919 31.8661
R15039 gnd.n5461 gnd.n1913 31.8661
R15040 gnd.n5461 gnd.n1906 31.8661
R15041 gnd.n5469 gnd.n1906 31.8661
R15042 gnd.n5477 gnd.n1900 31.8661
R15043 gnd.n5477 gnd.n1892 31.8661
R15044 gnd.n5485 gnd.n1892 31.8661
R15045 gnd.n5485 gnd.n1894 31.8661
R15046 gnd.n5493 gnd.n1880 31.8661
R15047 gnd.n5501 gnd.n1880 31.8661
R15048 gnd.n5501 gnd.n1874 31.8661
R15049 gnd.n5509 gnd.n1874 31.8661
R15050 gnd.n5717 gnd.n1692 31.8661
R15051 gnd.n5717 gnd.n1684 31.8661
R15052 gnd.n5725 gnd.n1684 31.8661
R15053 gnd.n5725 gnd.n1686 31.8661
R15054 gnd.n5733 gnd.n1672 31.8661
R15055 gnd.n5741 gnd.n1672 31.8661
R15056 gnd.n5741 gnd.n1666 31.8661
R15057 gnd.n5749 gnd.n1666 31.8661
R15058 gnd.n5757 gnd.n1659 31.8661
R15059 gnd.n5757 gnd.n1653 31.8661
R15060 gnd.n5765 gnd.n1653 31.8661
R15061 gnd.n5773 gnd.n1646 31.8661
R15062 gnd.n5773 gnd.n1639 31.8661
R15063 gnd.n5781 gnd.n1639 31.8661
R15064 gnd.n5781 gnd.n1640 31.8661
R15065 gnd.n5789 gnd.n1626 31.8661
R15066 gnd.n5799 gnd.n1626 31.8661
R15067 gnd.n5799 gnd.n1618 31.8661
R15068 gnd.n5810 gnd.n1618 31.8661
R15069 gnd.n6101 gnd.n1245 31.8661
R15070 gnd.n6101 gnd.n6100 31.8661
R15071 gnd.n6094 gnd.n1256 31.8661
R15072 gnd.n6094 gnd.n6093 31.8661
R15073 gnd.n1336 gnd.n1285 31.8661
R15074 gnd.n7242 gnd.n350 31.8661
R15075 gnd.n7349 gnd.n315 31.8661
R15076 gnd.n7251 gnd.n340 31.8661
R15077 gnd.n7257 gnd.n340 31.8661
R15078 gnd.n7330 gnd.n334 31.8661
R15079 gnd.n7334 gnd.n299 31.8661
R15080 gnd.n7358 gnd.n299 31.8661
R15081 gnd.n7366 gnd.n290 31.8661
R15082 gnd.n7366 gnd.n293 31.8661
R15083 gnd.n7374 gnd.n284 31.8661
R15084 gnd.n7382 gnd.n269 31.8661
R15085 gnd.n7390 gnd.n269 31.8661
R15086 gnd.n7398 gnd.n260 31.8661
R15087 gnd.n7398 gnd.n263 31.8661
R15088 gnd.n7406 gnd.n254 31.8661
R15089 gnd.n7414 gnd.n247 31.8661
R15090 gnd.n7430 gnd.n229 31.8661
R15091 gnd.n7430 gnd.n232 31.8661
R15092 gnd.n7438 gnd.n213 31.8661
R15093 gnd.n7514 gnd.n213 31.8661
R15094 gnd.n7514 gnd.n206 31.8661
R15095 gnd.n7522 gnd.n206 31.8661
R15096 gnd.n7602 gnd.n126 31.8661
R15097 gnd.t107 gnd.n2201 31.5474
R15098 gnd.n7330 gnd.t13 31.5474
R15099 gnd.n5084 gnd.n4888 31.0639
R15100 gnd.n4732 gnd.n4729 31.0639
R15101 gnd.t141 gnd.n2233 30.9101
R15102 gnd.n284 gnd.t19 30.9101
R15103 gnd.n3792 gnd.n962 30.2728
R15104 gnd.t40 gnd.n2265 30.2728
R15105 gnd.n254 gnd.t89 30.2728
R15106 gnd.n3957 gnd.t314 28.3609
R15107 gnd.t247 gnd.n126 28.3609
R15108 gnd.n2393 gnd.n962 27.0862
R15109 gnd.n5469 gnd.t79 27.0862
R15110 gnd.t103 gnd.n1659 27.0862
R15111 gnd.n4529 gnd.n4528 25.7944
R15112 gnd.n2813 gnd.n2812 25.7944
R15113 gnd.n2358 gnd.n2357 25.7944
R15114 gnd.n123 gnd.n122 25.7944
R15115 gnd.n1487 gnd.n1486 25.7944
R15116 gnd.n2017 gnd.n2016 25.7944
R15117 gnd.n1309 gnd.n1308 25.7944
R15118 gnd.n1331 gnd.n1330 25.7944
R15119 gnd.n202 gnd.n201 25.7944
R15120 gnd.n7566 gnd.n7565 25.7944
R15121 gnd.n3986 gnd.n3985 25.7944
R15122 gnd.n4018 gnd.n4017 25.7944
R15123 gnd.n3799 gnd.n3798 25.7944
R15124 gnd.n2106 gnd.n2105 25.7944
R15125 gnd.n2084 gnd.n2083 25.7944
R15126 gnd.n5828 gnd.n5827 25.7944
R15127 gnd.n3034 gnd.n2754 24.8557
R15128 gnd.n3044 gnd.n2737 24.8557
R15129 gnd.n2740 gnd.n2728 24.8557
R15130 gnd.n3065 gnd.n2729 24.8557
R15131 gnd.n3075 gnd.n2709 24.8557
R15132 gnd.n3085 gnd.n3084 24.8557
R15133 gnd.n2695 gnd.n2693 24.8557
R15134 gnd.n3116 gnd.n3115 24.8557
R15135 gnd.n3131 gnd.n2678 24.8557
R15136 gnd.n3185 gnd.n2617 24.8557
R15137 gnd.n3141 gnd.n2618 24.8557
R15138 gnd.n3178 gnd.n2629 24.8557
R15139 gnd.n2667 gnd.n2666 24.8557
R15140 gnd.n3172 gnd.n3171 24.8557
R15141 gnd.n2653 gnd.n2640 24.8557
R15142 gnd.n3211 gnd.n3210 24.8557
R15143 gnd.n3221 gnd.n2537 24.8557
R15144 gnd.n3233 gnd.n2529 24.8557
R15145 gnd.n3232 gnd.n2517 24.8557
R15146 gnd.n3251 gnd.n3250 24.8557
R15147 gnd.n3261 gnd.n2510 24.8557
R15148 gnd.n3272 gnd.n2498 24.8557
R15149 gnd.n3296 gnd.n3295 24.8557
R15150 gnd.n3307 gnd.n2481 24.8557
R15151 gnd.n3306 gnd.n2483 24.8557
R15152 gnd.n3318 gnd.n2474 24.8557
R15153 gnd.n3336 gnd.n3335 24.8557
R15154 gnd.n2465 gnd.n2454 24.8557
R15155 gnd.n3357 gnd.n2442 24.8557
R15156 gnd.n3385 gnd.n3384 24.8557
R15157 gnd.n3396 gnd.n2427 24.8557
R15158 gnd.n3407 gnd.n2420 24.8557
R15159 gnd.n3406 gnd.n2408 24.8557
R15160 gnd.n3679 gnd.n3678 24.8557
R15161 gnd.n3701 gnd.n2392 24.8557
R15162 gnd.n5413 gnd.t284 24.537
R15163 gnd.t154 gnd.n1913 24.537
R15164 gnd.n5765 gnd.t236 24.537
R15165 gnd.t255 gnd.n1245 24.537
R15166 gnd.n7422 gnd.n238 24.537
R15167 gnd.n6340 gnd.n6339 24.2183
R15168 gnd.n6333 gnd.n983 24.2183
R15169 gnd.n4362 gnd.n986 24.2183
R15170 gnd.n4393 gnd.n997 24.2183
R15171 gnd.n4370 gnd.n1007 24.2183
R15172 gnd.n6315 gnd.n1015 24.2183
R15173 gnd.n6309 gnd.n1026 24.2183
R15174 gnd.n4411 gnd.n1029 24.2183
R15175 gnd.n4442 gnd.n1039 24.2183
R15176 gnd.n4419 gnd.n1049 24.2183
R15177 gnd.n6291 gnd.n1057 24.2183
R15178 gnd.n6285 gnd.n1068 24.2183
R15179 gnd.n4496 gnd.n1071 24.2183
R15180 gnd.n4504 gnd.n1081 24.2183
R15181 gnd.n6273 gnd.n1089 24.2183
R15182 gnd.n4513 gnd.n1092 24.2183
R15183 gnd.n6267 gnd.n1100 24.2183
R15184 gnd.n4553 gnd.n2109 24.2183
R15185 gnd.n6261 gnd.n1109 24.2183
R15186 gnd.n6016 gnd.n1338 24.2183
R15187 gnd.n5851 gnd.n5842 24.2183
R15188 gnd.n5861 gnd.n1452 24.2183
R15189 gnd.n5860 gnd.n1431 24.2183
R15190 gnd.n5872 gnd.n5871 24.2183
R15191 gnd.n1435 gnd.n1422 24.2183
R15192 gnd.n5897 gnd.n1414 24.2183
R15193 gnd.n5896 gnd.n1404 24.2183
R15194 gnd.n1407 gnd.n1394 24.2183
R15195 gnd.n5919 gnd.n1396 24.2183
R15196 gnd.n5957 gnd.n1370 24.2183
R15197 gnd.n1373 gnd.n1361 24.2183
R15198 gnd.n5987 gnd.n1364 24.2183
R15199 gnd.n7172 gnd.n402 24.2183
R15200 gnd.n5941 gnd.n390 24.2183
R15201 gnd.n7163 gnd.n384 24.2183
R15202 gnd.n7218 gnd.n370 24.2183
R15203 gnd.n7190 gnd.n377 24.2183
R15204 gnd.n7227 gnd.n358 24.2183
R15205 gnd.n5404 gnd.n1971 23.8997
R15206 gnd.n6100 gnd.n1248 23.8997
R15207 gnd.n3055 gnd.t70 23.2624
R15208 gnd.n4203 gnd.t3 23.2624
R15209 gnd.n4394 gnd.t17 23.2624
R15210 gnd.n6279 gnd.t42 23.2624
R15211 gnd.n5882 gnd.t29 23.2624
R15212 gnd.n7162 gnd.t84 23.2624
R15213 gnd.n7438 gnd.t73 23.2624
R15214 gnd.n2756 gnd.t329 22.6251
R15215 gnd.n4235 gnd.t81 22.6251
R15216 gnd.n6303 gnd.t52 22.6251
R15217 gnd.n4443 gnd.t37 22.6251
R15218 gnd.n5958 gnd.t44 22.6251
R15219 gnd.n5979 gnd.t33 22.6251
R15220 gnd.n7406 gnd.t50 22.6251
R15221 gnd.n2177 gnd.t31 22.3064
R15222 gnd.n5709 gnd.n1698 22.3064
R15223 gnd.t46 gnd.n312 22.3064
R15224 gnd.n4267 gnd.t169 21.9878
R15225 gnd.n6327 gnd.t150 21.9878
R15226 gnd.n7196 gnd.t5 21.9878
R15227 gnd.n7374 gnd.t11 21.9878
R15228 gnd.n5243 gnd.n1852 21.6691
R15229 gnd.n5236 gnd.n1846 21.6691
R15230 gnd.n5221 gnd.n5220 21.6691
R15231 gnd.n5207 gnd.n1818 21.6691
R15232 gnd.n5185 gnd.n1797 21.6691
R15233 gnd.n5178 gnd.n1790 21.6691
R15234 gnd.n5170 gnd.n1784 21.6691
R15235 gnd.n5163 gnd.n1776 21.6691
R15236 gnd.n5135 gnd.n4849 21.6691
R15237 gnd.n5122 gnd.n1733 21.6691
R15238 gnd.n5107 gnd.n1720 21.6691
R15239 gnd.t62 gnd.n2761 21.3504
R15240 gnd.n4301 gnd.t86 21.3504
R15241 gnd.n4328 gnd.t160 21.3504
R15242 gnd.t101 gnd.n315 21.3504
R15243 gnd.t195 gnd.n334 21.3504
R15244 gnd.n5573 gnd.n1820 21.0318
R15245 gnd.n5581 gnd.n1810 21.0318
R15246 gnd.n5147 gnd.n1754 21.0318
R15247 gnd.n5141 gnd.n4844 21.0318
R15248 gnd.t224 gnd.n2455 20.7131
R15249 gnd.n4284 gnd.t98 20.7131
R15250 gnd.n7358 gnd.t9 20.7131
R15251 gnd.t210 gnd.n2490 20.0758
R15252 gnd.n4251 gnd.t27 20.0758
R15253 gnd.n7390 gnd.t35 20.0758
R15254 gnd.n4645 gnd.t305 19.8005
R15255 gnd.n4645 gnd.t245 19.8005
R15256 gnd.n4646 gnd.t282 19.8005
R15257 gnd.n4646 gnd.t321 19.8005
R15258 gnd.n4933 gnd.t334 19.8005
R15259 gnd.n4933 gnd.t299 19.8005
R15260 gnd.n4934 gnd.t319 19.8005
R15261 gnd.n4934 gnd.t279 19.8005
R15262 gnd.n5354 gnd.n2043 19.7572
R15263 gnd.n4663 gnd.n1868 19.7572
R15264 gnd.n5565 gnd.n1827 19.7572
R15265 gnd.n5589 gnd.n1803 19.7572
R15266 gnd.n4831 gnd.n1761 19.7572
R15267 gnd.n4853 gnd.n1748 19.7572
R15268 gnd.n5701 gnd.n1707 19.7572
R15269 gnd.n6093 gnd.n6092 19.7572
R15270 gnd.n4642 gnd.n4641 19.5087
R15271 gnd.n4655 gnd.n4642 19.5087
R15272 gnd.n4653 gnd.n4644 19.5087
R15273 gnd.n4938 gnd.n4932 19.5087
R15274 gnd.n3222 gnd.t216 19.4385
R15275 gnd.n4219 gnd.t7 19.4385
R15276 gnd.n1939 gnd.t350 19.4385
R15277 gnd.n5789 gnd.t133 19.4385
R15278 gnd.n7422 gnd.t148 19.4385
R15279 gnd.n5411 gnd.n1954 19.3944
R15280 gnd.n5411 gnd.n1943 19.3944
R15281 gnd.n5423 gnd.n1943 19.3944
R15282 gnd.n5423 gnd.n1941 19.3944
R15283 gnd.n5427 gnd.n1941 19.3944
R15284 gnd.n5427 gnd.n1930 19.3944
R15285 gnd.n5439 gnd.n1930 19.3944
R15286 gnd.n5439 gnd.n1928 19.3944
R15287 gnd.n5443 gnd.n1928 19.3944
R15288 gnd.n5443 gnd.n1917 19.3944
R15289 gnd.n5455 gnd.n1917 19.3944
R15290 gnd.n5455 gnd.n1915 19.3944
R15291 gnd.n5459 gnd.n1915 19.3944
R15292 gnd.n5459 gnd.n1904 19.3944
R15293 gnd.n5471 gnd.n1904 19.3944
R15294 gnd.n5471 gnd.n1902 19.3944
R15295 gnd.n5475 gnd.n1902 19.3944
R15296 gnd.n5475 gnd.n1890 19.3944
R15297 gnd.n5487 gnd.n1890 19.3944
R15298 gnd.n5487 gnd.n1888 19.3944
R15299 gnd.n5491 gnd.n1888 19.3944
R15300 gnd.n5491 gnd.n1878 19.3944
R15301 gnd.n5503 gnd.n1878 19.3944
R15302 gnd.n5503 gnd.n1876 19.3944
R15303 gnd.n5507 gnd.n1876 19.3944
R15304 gnd.n5507 gnd.n1864 19.3944
R15305 gnd.n5519 gnd.n1864 19.3944
R15306 gnd.n5519 gnd.n1862 19.3944
R15307 gnd.n5523 gnd.n1862 19.3944
R15308 gnd.n5523 gnd.n1850 19.3944
R15309 gnd.n5535 gnd.n1850 19.3944
R15310 gnd.n5535 gnd.n1848 19.3944
R15311 gnd.n5539 gnd.n1848 19.3944
R15312 gnd.n5539 gnd.n1837 19.3944
R15313 gnd.n5551 gnd.n1837 19.3944
R15314 gnd.n5551 gnd.n1835 19.3944
R15315 gnd.n5555 gnd.n1835 19.3944
R15316 gnd.n5555 gnd.n1824 19.3944
R15317 gnd.n5567 gnd.n1824 19.3944
R15318 gnd.n5567 gnd.n1822 19.3944
R15319 gnd.n5571 gnd.n1822 19.3944
R15320 gnd.n5571 gnd.n1808 19.3944
R15321 gnd.n5583 gnd.n1808 19.3944
R15322 gnd.n5583 gnd.n1806 19.3944
R15323 gnd.n5587 gnd.n1806 19.3944
R15324 gnd.n5587 gnd.n1794 19.3944
R15325 gnd.n5599 gnd.n1794 19.3944
R15326 gnd.n5599 gnd.n1792 19.3944
R15327 gnd.n5603 gnd.n1792 19.3944
R15328 gnd.n5603 gnd.n1780 19.3944
R15329 gnd.n5615 gnd.n1780 19.3944
R15330 gnd.n5615 gnd.n1778 19.3944
R15331 gnd.n5619 gnd.n1778 19.3944
R15332 gnd.n5619 gnd.n1766 19.3944
R15333 gnd.n5631 gnd.n1766 19.3944
R15334 gnd.n5631 gnd.n1764 19.3944
R15335 gnd.n5635 gnd.n1764 19.3944
R15336 gnd.n5635 gnd.n1752 19.3944
R15337 gnd.n5647 gnd.n1752 19.3944
R15338 gnd.n5647 gnd.n1750 19.3944
R15339 gnd.n5651 gnd.n1750 19.3944
R15340 gnd.n5651 gnd.n1738 19.3944
R15341 gnd.n5663 gnd.n1738 19.3944
R15342 gnd.n5663 gnd.n1736 19.3944
R15343 gnd.n5667 gnd.n1736 19.3944
R15344 gnd.n5667 gnd.n1724 19.3944
R15345 gnd.n5679 gnd.n1724 19.3944
R15346 gnd.n5679 gnd.n1722 19.3944
R15347 gnd.n5683 gnd.n1722 19.3944
R15348 gnd.n5683 gnd.n1711 19.3944
R15349 gnd.n5695 gnd.n1711 19.3944
R15350 gnd.n5695 gnd.n1709 19.3944
R15351 gnd.n5699 gnd.n1709 19.3944
R15352 gnd.n5699 gnd.n1696 19.3944
R15353 gnd.n5711 gnd.n1696 19.3944
R15354 gnd.n5711 gnd.n1694 19.3944
R15355 gnd.n5715 gnd.n1694 19.3944
R15356 gnd.n5715 gnd.n1682 19.3944
R15357 gnd.n5727 gnd.n1682 19.3944
R15358 gnd.n5727 gnd.n1680 19.3944
R15359 gnd.n5731 gnd.n1680 19.3944
R15360 gnd.n5731 gnd.n1670 19.3944
R15361 gnd.n5743 gnd.n1670 19.3944
R15362 gnd.n5743 gnd.n1668 19.3944
R15363 gnd.n5747 gnd.n1668 19.3944
R15364 gnd.n5747 gnd.n1657 19.3944
R15365 gnd.n5759 gnd.n1657 19.3944
R15366 gnd.n5759 gnd.n1655 19.3944
R15367 gnd.n5763 gnd.n1655 19.3944
R15368 gnd.n5763 gnd.n1644 19.3944
R15369 gnd.n5775 gnd.n1644 19.3944
R15370 gnd.n5775 gnd.n1642 19.3944
R15371 gnd.n5779 gnd.n1642 19.3944
R15372 gnd.n5779 gnd.n1631 19.3944
R15373 gnd.n5791 gnd.n1631 19.3944
R15374 gnd.n5791 gnd.n1628 19.3944
R15375 gnd.n5797 gnd.n1628 19.3944
R15376 gnd.n5797 gnd.n1629 19.3944
R15377 gnd.n1629 gnd.n1616 19.3944
R15378 gnd.n5813 gnd.n1616 19.3944
R15379 gnd.n5814 gnd.n5813 19.3944
R15380 gnd.n4535 gnd.n4534 19.3944
R15381 gnd.n4534 gnd.n1956 19.3944
R15382 gnd.n5407 gnd.n1956 19.3944
R15383 gnd.n5401 gnd.n5400 19.3944
R15384 gnd.n5400 gnd.n1975 19.3944
R15385 gnd.n5393 gnd.n1975 19.3944
R15386 gnd.n5393 gnd.n5392 19.3944
R15387 gnd.n5392 gnd.n1986 19.3944
R15388 gnd.n5385 gnd.n1986 19.3944
R15389 gnd.n5385 gnd.n5384 19.3944
R15390 gnd.n5384 gnd.n1994 19.3944
R15391 gnd.n5377 gnd.n1994 19.3944
R15392 gnd.n5377 gnd.n5376 19.3944
R15393 gnd.n5376 gnd.n2004 19.3944
R15394 gnd.n5369 gnd.n2004 19.3944
R15395 gnd.n5369 gnd.n5368 19.3944
R15396 gnd.n5368 gnd.n2012 19.3944
R15397 gnd.n5361 gnd.n2012 19.3944
R15398 gnd.n5361 gnd.n5360 19.3944
R15399 gnd.n5360 gnd.n2024 19.3944
R15400 gnd.n4546 gnd.n2024 19.3944
R15401 gnd.n4546 gnd.n4545 19.3944
R15402 gnd.n4545 gnd.n4544 19.3944
R15403 gnd.n4544 gnd.n4523 19.3944
R15404 gnd.n4540 gnd.n4523 19.3944
R15405 gnd.n4540 gnd.n4539 19.3944
R15406 gnd.n4539 gnd.n4538 19.3944
R15407 gnd.n2937 gnd.n2936 19.3944
R15408 gnd.n2936 gnd.n2935 19.3944
R15409 gnd.n2935 gnd.n2934 19.3944
R15410 gnd.n2934 gnd.n2932 19.3944
R15411 gnd.n2932 gnd.n2929 19.3944
R15412 gnd.n2929 gnd.n2928 19.3944
R15413 gnd.n2928 gnd.n2925 19.3944
R15414 gnd.n2925 gnd.n2924 19.3944
R15415 gnd.n2924 gnd.n2921 19.3944
R15416 gnd.n2921 gnd.n2920 19.3944
R15417 gnd.n2920 gnd.n2917 19.3944
R15418 gnd.n2917 gnd.n2916 19.3944
R15419 gnd.n2916 gnd.n2913 19.3944
R15420 gnd.n2913 gnd.n2912 19.3944
R15421 gnd.n2912 gnd.n2909 19.3944
R15422 gnd.n2909 gnd.n2908 19.3944
R15423 gnd.n2908 gnd.n2905 19.3944
R15424 gnd.n2905 gnd.n2904 19.3944
R15425 gnd.n2904 gnd.n2901 19.3944
R15426 gnd.n2901 gnd.n2900 19.3944
R15427 gnd.n2900 gnd.n2897 19.3944
R15428 gnd.n2897 gnd.n2896 19.3944
R15429 gnd.n2893 gnd.n2892 19.3944
R15430 gnd.n2892 gnd.n2848 19.3944
R15431 gnd.n2943 gnd.n2848 19.3944
R15432 gnd.n3709 gnd.n3708 19.3944
R15433 gnd.n3708 gnd.n3705 19.3944
R15434 gnd.n3705 gnd.n3704 19.3944
R15435 gnd.n3754 gnd.n3753 19.3944
R15436 gnd.n3753 gnd.n3752 19.3944
R15437 gnd.n3752 gnd.n3749 19.3944
R15438 gnd.n3749 gnd.n3748 19.3944
R15439 gnd.n3748 gnd.n3745 19.3944
R15440 gnd.n3745 gnd.n3744 19.3944
R15441 gnd.n3744 gnd.n3741 19.3944
R15442 gnd.n3741 gnd.n3740 19.3944
R15443 gnd.n3740 gnd.n3737 19.3944
R15444 gnd.n3737 gnd.n3736 19.3944
R15445 gnd.n3736 gnd.n3733 19.3944
R15446 gnd.n3733 gnd.n3732 19.3944
R15447 gnd.n3732 gnd.n3729 19.3944
R15448 gnd.n3729 gnd.n3728 19.3944
R15449 gnd.n3728 gnd.n3725 19.3944
R15450 gnd.n3725 gnd.n3724 19.3944
R15451 gnd.n3724 gnd.n3721 19.3944
R15452 gnd.n3721 gnd.n3720 19.3944
R15453 gnd.n3720 gnd.n3717 19.3944
R15454 gnd.n3717 gnd.n3716 19.3944
R15455 gnd.n3716 gnd.n3713 19.3944
R15456 gnd.n3713 gnd.n3712 19.3944
R15457 gnd.n3036 gnd.n2745 19.3944
R15458 gnd.n3046 gnd.n2745 19.3944
R15459 gnd.n3047 gnd.n3046 19.3944
R15460 gnd.n3047 gnd.n2726 19.3944
R15461 gnd.n3067 gnd.n2726 19.3944
R15462 gnd.n3067 gnd.n2718 19.3944
R15463 gnd.n3077 gnd.n2718 19.3944
R15464 gnd.n3078 gnd.n3077 19.3944
R15465 gnd.n3079 gnd.n3078 19.3944
R15466 gnd.n3079 gnd.n2701 19.3944
R15467 gnd.n3096 gnd.n2701 19.3944
R15468 gnd.n3099 gnd.n3096 19.3944
R15469 gnd.n3099 gnd.n3098 19.3944
R15470 gnd.n3098 gnd.n2674 19.3944
R15471 gnd.n3138 gnd.n2674 19.3944
R15472 gnd.n3138 gnd.n2671 19.3944
R15473 gnd.n3144 gnd.n2671 19.3944
R15474 gnd.n3145 gnd.n3144 19.3944
R15475 gnd.n3145 gnd.n2669 19.3944
R15476 gnd.n3151 gnd.n2669 19.3944
R15477 gnd.n3154 gnd.n3151 19.3944
R15478 gnd.n3156 gnd.n3154 19.3944
R15479 gnd.n3162 gnd.n3156 19.3944
R15480 gnd.n3162 gnd.n3161 19.3944
R15481 gnd.n3161 gnd.n2532 19.3944
R15482 gnd.n3228 gnd.n2532 19.3944
R15483 gnd.n3229 gnd.n3228 19.3944
R15484 gnd.n3229 gnd.n2525 19.3944
R15485 gnd.n3240 gnd.n2525 19.3944
R15486 gnd.n3241 gnd.n3240 19.3944
R15487 gnd.n3241 gnd.n2508 19.3944
R15488 gnd.n2508 gnd.n2506 19.3944
R15489 gnd.n3265 gnd.n2506 19.3944
R15490 gnd.n3266 gnd.n3265 19.3944
R15491 gnd.n3266 gnd.n2477 19.3944
R15492 gnd.n3313 gnd.n2477 19.3944
R15493 gnd.n3314 gnd.n3313 19.3944
R15494 gnd.n3314 gnd.n2470 19.3944
R15495 gnd.n3325 gnd.n2470 19.3944
R15496 gnd.n3326 gnd.n3325 19.3944
R15497 gnd.n3326 gnd.n2453 19.3944
R15498 gnd.n2453 gnd.n2451 19.3944
R15499 gnd.n3350 gnd.n2451 19.3944
R15500 gnd.n3351 gnd.n3350 19.3944
R15501 gnd.n3351 gnd.n2423 19.3944
R15502 gnd.n3402 gnd.n2423 19.3944
R15503 gnd.n3403 gnd.n3402 19.3944
R15504 gnd.n3403 gnd.n2416 19.3944
R15505 gnd.n3670 gnd.n2416 19.3944
R15506 gnd.n3671 gnd.n3670 19.3944
R15507 gnd.n3671 gnd.n2397 19.3944
R15508 gnd.n3696 gnd.n2397 19.3944
R15509 gnd.n3696 gnd.n2398 19.3944
R15510 gnd.n3027 gnd.n3026 19.3944
R15511 gnd.n3026 gnd.n2759 19.3944
R15512 gnd.n2782 gnd.n2759 19.3944
R15513 gnd.n2785 gnd.n2782 19.3944
R15514 gnd.n2785 gnd.n2778 19.3944
R15515 gnd.n2789 gnd.n2778 19.3944
R15516 gnd.n2792 gnd.n2789 19.3944
R15517 gnd.n2795 gnd.n2792 19.3944
R15518 gnd.n2795 gnd.n2776 19.3944
R15519 gnd.n2799 gnd.n2776 19.3944
R15520 gnd.n2802 gnd.n2799 19.3944
R15521 gnd.n2805 gnd.n2802 19.3944
R15522 gnd.n2805 gnd.n2774 19.3944
R15523 gnd.n2809 gnd.n2774 19.3944
R15524 gnd.n3032 gnd.n3031 19.3944
R15525 gnd.n3031 gnd.n2735 19.3944
R15526 gnd.n3057 gnd.n2735 19.3944
R15527 gnd.n3057 gnd.n2733 19.3944
R15528 gnd.n3063 gnd.n2733 19.3944
R15529 gnd.n3063 gnd.n3062 19.3944
R15530 gnd.n3062 gnd.n2707 19.3944
R15531 gnd.n3087 gnd.n2707 19.3944
R15532 gnd.n3087 gnd.n2705 19.3944
R15533 gnd.n3091 gnd.n2705 19.3944
R15534 gnd.n3091 gnd.n2685 19.3944
R15535 gnd.n3118 gnd.n2685 19.3944
R15536 gnd.n3118 gnd.n2683 19.3944
R15537 gnd.n3128 gnd.n2683 19.3944
R15538 gnd.n3128 gnd.n3127 19.3944
R15539 gnd.n3127 gnd.n3126 19.3944
R15540 gnd.n3126 gnd.n2632 19.3944
R15541 gnd.n3176 gnd.n2632 19.3944
R15542 gnd.n3176 gnd.n3175 19.3944
R15543 gnd.n3175 gnd.n3174 19.3944
R15544 gnd.n3174 gnd.n2636 19.3944
R15545 gnd.n2656 gnd.n2636 19.3944
R15546 gnd.n2656 gnd.n2542 19.3944
R15547 gnd.n3213 gnd.n2542 19.3944
R15548 gnd.n3213 gnd.n2540 19.3944
R15549 gnd.n3219 gnd.n2540 19.3944
R15550 gnd.n3219 gnd.n3218 19.3944
R15551 gnd.n3218 gnd.n2515 19.3944
R15552 gnd.n3253 gnd.n2515 19.3944
R15553 gnd.n3253 gnd.n2513 19.3944
R15554 gnd.n3259 gnd.n2513 19.3944
R15555 gnd.n3259 gnd.n3258 19.3944
R15556 gnd.n3258 gnd.n2488 19.3944
R15557 gnd.n3298 gnd.n2488 19.3944
R15558 gnd.n3298 gnd.n2486 19.3944
R15559 gnd.n3304 gnd.n2486 19.3944
R15560 gnd.n3304 gnd.n3303 19.3944
R15561 gnd.n3303 gnd.n2460 19.3944
R15562 gnd.n3338 gnd.n2460 19.3944
R15563 gnd.n3338 gnd.n2458 19.3944
R15564 gnd.n3344 gnd.n2458 19.3944
R15565 gnd.n3344 gnd.n3343 19.3944
R15566 gnd.n3343 gnd.n2433 19.3944
R15567 gnd.n3387 gnd.n2433 19.3944
R15568 gnd.n3387 gnd.n2431 19.3944
R15569 gnd.n3393 gnd.n2431 19.3944
R15570 gnd.n3393 gnd.n3392 19.3944
R15571 gnd.n3392 gnd.n2406 19.3944
R15572 gnd.n3681 gnd.n2406 19.3944
R15573 gnd.n3681 gnd.n2404 19.3944
R15574 gnd.n3689 gnd.n2404 19.3944
R15575 gnd.n3689 gnd.n3688 19.3944
R15576 gnd.n3688 gnd.n3687 19.3944
R15577 gnd.n3790 gnd.n3789 19.3944
R15578 gnd.n3789 gnd.n2344 19.3944
R15579 gnd.n3785 gnd.n2344 19.3944
R15580 gnd.n3785 gnd.n3782 19.3944
R15581 gnd.n3782 gnd.n3779 19.3944
R15582 gnd.n3779 gnd.n3778 19.3944
R15583 gnd.n3778 gnd.n3775 19.3944
R15584 gnd.n3775 gnd.n3774 19.3944
R15585 gnd.n3774 gnd.n3771 19.3944
R15586 gnd.n3771 gnd.n3770 19.3944
R15587 gnd.n3770 gnd.n3767 19.3944
R15588 gnd.n3767 gnd.n3766 19.3944
R15589 gnd.n3766 gnd.n3763 19.3944
R15590 gnd.n3763 gnd.n3762 19.3944
R15591 gnd.n2947 gnd.n2846 19.3944
R15592 gnd.n2947 gnd.n2837 19.3944
R15593 gnd.n2960 gnd.n2837 19.3944
R15594 gnd.n2960 gnd.n2835 19.3944
R15595 gnd.n2964 gnd.n2835 19.3944
R15596 gnd.n2964 gnd.n2825 19.3944
R15597 gnd.n2976 gnd.n2825 19.3944
R15598 gnd.n2976 gnd.n2823 19.3944
R15599 gnd.n3010 gnd.n2823 19.3944
R15600 gnd.n3010 gnd.n3009 19.3944
R15601 gnd.n3009 gnd.n3008 19.3944
R15602 gnd.n3008 gnd.n3007 19.3944
R15603 gnd.n3007 gnd.n3004 19.3944
R15604 gnd.n3004 gnd.n3003 19.3944
R15605 gnd.n3003 gnd.n3002 19.3944
R15606 gnd.n3002 gnd.n3000 19.3944
R15607 gnd.n3000 gnd.n2999 19.3944
R15608 gnd.n2999 gnd.n2996 19.3944
R15609 gnd.n2996 gnd.n2995 19.3944
R15610 gnd.n2995 gnd.n2994 19.3944
R15611 gnd.n2994 gnd.n2992 19.3944
R15612 gnd.n2992 gnd.n2691 19.3944
R15613 gnd.n3107 gnd.n2691 19.3944
R15614 gnd.n3107 gnd.n2689 19.3944
R15615 gnd.n3113 gnd.n2689 19.3944
R15616 gnd.n3113 gnd.n3112 19.3944
R15617 gnd.n3112 gnd.n2613 19.3944
R15618 gnd.n3187 gnd.n2613 19.3944
R15619 gnd.n3187 gnd.n2614 19.3944
R15620 gnd.n2661 gnd.n2660 19.3944
R15621 gnd.n2664 gnd.n2663 19.3944
R15622 gnd.n2651 gnd.n2650 19.3944
R15623 gnd.n3206 gnd.n2547 19.3944
R15624 gnd.n3206 gnd.n3205 19.3944
R15625 gnd.n3205 gnd.n3204 19.3944
R15626 gnd.n3204 gnd.n3202 19.3944
R15627 gnd.n3202 gnd.n3201 19.3944
R15628 gnd.n3201 gnd.n3199 19.3944
R15629 gnd.n3199 gnd.n3198 19.3944
R15630 gnd.n3198 gnd.n2496 19.3944
R15631 gnd.n3274 gnd.n2496 19.3944
R15632 gnd.n3274 gnd.n2494 19.3944
R15633 gnd.n3293 gnd.n2494 19.3944
R15634 gnd.n3293 gnd.n3292 19.3944
R15635 gnd.n3292 gnd.n3291 19.3944
R15636 gnd.n3291 gnd.n3289 19.3944
R15637 gnd.n3289 gnd.n3288 19.3944
R15638 gnd.n3288 gnd.n3286 19.3944
R15639 gnd.n3286 gnd.n3285 19.3944
R15640 gnd.n3285 gnd.n2440 19.3944
R15641 gnd.n3359 gnd.n2440 19.3944
R15642 gnd.n3359 gnd.n2438 19.3944
R15643 gnd.n3382 gnd.n2438 19.3944
R15644 gnd.n3382 gnd.n3381 19.3944
R15645 gnd.n3381 gnd.n3380 19.3944
R15646 gnd.n3380 gnd.n3377 19.3944
R15647 gnd.n3377 gnd.n3376 19.3944
R15648 gnd.n3376 gnd.n3374 19.3944
R15649 gnd.n3374 gnd.n3373 19.3944
R15650 gnd.n3373 gnd.n3371 19.3944
R15651 gnd.n3371 gnd.n2391 19.3944
R15652 gnd.n2952 gnd.n2842 19.3944
R15653 gnd.n2952 gnd.n2840 19.3944
R15654 gnd.n2956 gnd.n2840 19.3944
R15655 gnd.n2956 gnd.n2831 19.3944
R15656 gnd.n2968 gnd.n2831 19.3944
R15657 gnd.n2968 gnd.n2829 19.3944
R15658 gnd.n2972 gnd.n2829 19.3944
R15659 gnd.n2972 gnd.n2818 19.3944
R15660 gnd.n3014 gnd.n2818 19.3944
R15661 gnd.n3014 gnd.n2772 19.3944
R15662 gnd.n3020 gnd.n2772 19.3944
R15663 gnd.n3020 gnd.n3019 19.3944
R15664 gnd.n3019 gnd.n2750 19.3944
R15665 gnd.n3041 gnd.n2750 19.3944
R15666 gnd.n3041 gnd.n2743 19.3944
R15667 gnd.n3052 gnd.n2743 19.3944
R15668 gnd.n3052 gnd.n3051 19.3944
R15669 gnd.n3051 gnd.n2724 19.3944
R15670 gnd.n3072 gnd.n2724 19.3944
R15671 gnd.n3072 gnd.n2714 19.3944
R15672 gnd.n3082 gnd.n2714 19.3944
R15673 gnd.n3082 gnd.n2697 19.3944
R15674 gnd.n3103 gnd.n2697 19.3944
R15675 gnd.n3103 gnd.n3102 19.3944
R15676 gnd.n3102 gnd.n2676 19.3944
R15677 gnd.n3133 gnd.n2676 19.3944
R15678 gnd.n3133 gnd.n2621 19.3944
R15679 gnd.n3183 gnd.n2621 19.3944
R15680 gnd.n3183 gnd.n3182 19.3944
R15681 gnd.n3182 gnd.n3181 19.3944
R15682 gnd.n3181 gnd.n2625 19.3944
R15683 gnd.n2643 gnd.n2625 19.3944
R15684 gnd.n3169 gnd.n2643 19.3944
R15685 gnd.n3169 gnd.n3168 19.3944
R15686 gnd.n3168 gnd.n3167 19.3944
R15687 gnd.n3167 gnd.n2647 19.3944
R15688 gnd.n2647 gnd.n2534 19.3944
R15689 gnd.n3224 gnd.n2534 19.3944
R15690 gnd.n3224 gnd.n2527 19.3944
R15691 gnd.n3235 gnd.n2527 19.3944
R15692 gnd.n3235 gnd.n2523 19.3944
R15693 gnd.n3248 gnd.n2523 19.3944
R15694 gnd.n3248 gnd.n3247 19.3944
R15695 gnd.n3247 gnd.n2502 19.3944
R15696 gnd.n3270 gnd.n2502 19.3944
R15697 gnd.n3270 gnd.n3269 19.3944
R15698 gnd.n3269 gnd.n2479 19.3944
R15699 gnd.n3309 gnd.n2479 19.3944
R15700 gnd.n3309 gnd.n2472 19.3944
R15701 gnd.n3320 gnd.n2472 19.3944
R15702 gnd.n3320 gnd.n2468 19.3944
R15703 gnd.n3333 gnd.n2468 19.3944
R15704 gnd.n3333 gnd.n3332 19.3944
R15705 gnd.n3332 gnd.n2447 19.3944
R15706 gnd.n3355 gnd.n2447 19.3944
R15707 gnd.n3355 gnd.n3354 19.3944
R15708 gnd.n3354 gnd.n2425 19.3944
R15709 gnd.n3398 gnd.n2425 19.3944
R15710 gnd.n3398 gnd.n2418 19.3944
R15711 gnd.n3409 gnd.n2418 19.3944
R15712 gnd.n3409 gnd.n2414 19.3944
R15713 gnd.n3676 gnd.n2414 19.3944
R15714 gnd.n3676 gnd.n3675 19.3944
R15715 gnd.n3675 gnd.n2395 19.3944
R15716 gnd.n3699 gnd.n2395 19.3944
R15717 gnd.n5853 gnd.n5841 19.3944
R15718 gnd.n5853 gnd.n1476 19.3944
R15719 gnd.n5858 gnd.n1476 19.3944
R15720 gnd.n5858 gnd.n1477 19.3944
R15721 gnd.n1477 gnd.n1420 19.3944
R15722 gnd.n5884 gnd.n1420 19.3944
R15723 gnd.n5884 gnd.n1417 19.3944
R15724 gnd.n5894 gnd.n1417 19.3944
R15725 gnd.n5894 gnd.n1418 19.3944
R15726 gnd.n5890 gnd.n1418 19.3944
R15727 gnd.n5890 gnd.n5889 19.3944
R15728 gnd.n5889 gnd.n1382 19.3944
R15729 gnd.n5954 gnd.n1382 19.3944
R15730 gnd.n5954 gnd.n1383 19.3944
R15731 gnd.n5950 gnd.n1383 19.3944
R15732 gnd.n5950 gnd.n5949 19.3944
R15733 gnd.n5949 gnd.n5948 19.3944
R15734 gnd.n5948 gnd.n5938 19.3944
R15735 gnd.n5944 gnd.n5938 19.3944
R15736 gnd.n5944 gnd.n5943 19.3944
R15737 gnd.n5943 gnd.n382 19.3944
R15738 gnd.n7198 gnd.n382 19.3944
R15739 gnd.n7199 gnd.n7198 19.3944
R15740 gnd.n7199 gnd.n379 19.3944
R15741 gnd.n7204 gnd.n379 19.3944
R15742 gnd.n7204 gnd.n380 19.3944
R15743 gnd.n380 gnd.n348 19.3944
R15744 gnd.n7244 gnd.n348 19.3944
R15745 gnd.n7244 gnd.n346 19.3944
R15746 gnd.n7248 gnd.n346 19.3944
R15747 gnd.n7249 gnd.n7248 19.3944
R15748 gnd.n7249 gnd.n80 19.3944
R15749 gnd.n7653 gnd.n80 19.3944
R15750 gnd.n7653 gnd.n7652 19.3944
R15751 gnd.n7652 gnd.n7651 19.3944
R15752 gnd.n7651 gnd.n85 19.3944
R15753 gnd.n7647 gnd.n85 19.3944
R15754 gnd.n7647 gnd.n7646 19.3944
R15755 gnd.n7646 gnd.n7645 19.3944
R15756 gnd.n7645 gnd.n90 19.3944
R15757 gnd.n7641 gnd.n90 19.3944
R15758 gnd.n7641 gnd.n7640 19.3944
R15759 gnd.n7640 gnd.n7639 19.3944
R15760 gnd.n7639 gnd.n95 19.3944
R15761 gnd.n7635 gnd.n95 19.3944
R15762 gnd.n7635 gnd.n7634 19.3944
R15763 gnd.n7634 gnd.n7633 19.3944
R15764 gnd.n7633 gnd.n100 19.3944
R15765 gnd.n7629 gnd.n100 19.3944
R15766 gnd.n7629 gnd.n7628 19.3944
R15767 gnd.n7628 gnd.n7627 19.3944
R15768 gnd.n7627 gnd.n105 19.3944
R15769 gnd.n7623 gnd.n105 19.3944
R15770 gnd.n7623 gnd.n7622 19.3944
R15771 gnd.n7622 gnd.n7621 19.3944
R15772 gnd.n7621 gnd.n110 19.3944
R15773 gnd.n7617 gnd.n110 19.3944
R15774 gnd.n7617 gnd.n7616 19.3944
R15775 gnd.n7616 gnd.n7615 19.3944
R15776 gnd.n7615 gnd.n115 19.3944
R15777 gnd.n7611 gnd.n115 19.3944
R15778 gnd.n7611 gnd.n7610 19.3944
R15779 gnd.n7610 gnd.n7609 19.3944
R15780 gnd.n7609 gnd.n120 19.3944
R15781 gnd.n7503 gnd.n7502 19.3944
R15782 gnd.n7502 gnd.n7501 19.3944
R15783 gnd.n7501 gnd.n7450 19.3944
R15784 gnd.n7497 gnd.n7450 19.3944
R15785 gnd.n7497 gnd.n7496 19.3944
R15786 gnd.n7496 gnd.n7495 19.3944
R15787 gnd.n7495 gnd.n7458 19.3944
R15788 gnd.n7491 gnd.n7458 19.3944
R15789 gnd.n7491 gnd.n7490 19.3944
R15790 gnd.n7490 gnd.n7489 19.3944
R15791 gnd.n7489 gnd.n7466 19.3944
R15792 gnd.n7485 gnd.n7466 19.3944
R15793 gnd.n7485 gnd.n7484 19.3944
R15794 gnd.n7484 gnd.n7483 19.3944
R15795 gnd.n7483 gnd.n7474 19.3944
R15796 gnd.n7479 gnd.n7474 19.3944
R15797 gnd.n1521 gnd.n1517 19.3944
R15798 gnd.n1524 gnd.n1521 19.3944
R15799 gnd.n1527 gnd.n1524 19.3944
R15800 gnd.n1527 gnd.n1510 19.3944
R15801 gnd.n1540 gnd.n1510 19.3944
R15802 gnd.n1543 gnd.n1540 19.3944
R15803 gnd.n1546 gnd.n1543 19.3944
R15804 gnd.n1546 gnd.n1503 19.3944
R15805 gnd.n1559 gnd.n1503 19.3944
R15806 gnd.n1562 gnd.n1559 19.3944
R15807 gnd.n1565 gnd.n1562 19.3944
R15808 gnd.n1565 gnd.n1496 19.3944
R15809 gnd.n1577 gnd.n1496 19.3944
R15810 gnd.n1580 gnd.n1577 19.3944
R15811 gnd.n1580 gnd.n1488 19.3944
R15812 gnd.n1593 gnd.n1488 19.3944
R15813 gnd.n6014 gnd.n1341 19.3944
R15814 gnd.n6010 gnd.n1341 19.3944
R15815 gnd.n6010 gnd.n6009 19.3944
R15816 gnd.n6009 gnd.n6008 19.3944
R15817 gnd.n6008 gnd.n1347 19.3944
R15818 gnd.n6004 gnd.n1347 19.3944
R15819 gnd.n6004 gnd.n6003 19.3944
R15820 gnd.n6003 gnd.n6002 19.3944
R15821 gnd.n6002 gnd.n1352 19.3944
R15822 gnd.n5998 gnd.n1352 19.3944
R15823 gnd.n5998 gnd.n5997 19.3944
R15824 gnd.n5997 gnd.n5996 19.3944
R15825 gnd.n5996 gnd.n1357 19.3944
R15826 gnd.n5992 gnd.n1357 19.3944
R15827 gnd.n5992 gnd.n5991 19.3944
R15828 gnd.n5991 gnd.n5990 19.3944
R15829 gnd.n5990 gnd.n405 19.3944
R15830 gnd.n7170 gnd.n405 19.3944
R15831 gnd.n7170 gnd.n406 19.3944
R15832 gnd.n7166 gnd.n406 19.3944
R15833 gnd.n7166 gnd.n7165 19.3944
R15834 gnd.n7165 gnd.n373 19.3944
R15835 gnd.n7216 gnd.n373 19.3944
R15836 gnd.n7216 gnd.n374 19.3944
R15837 gnd.n7212 gnd.n374 19.3944
R15838 gnd.n7212 gnd.n7211 19.3944
R15839 gnd.n7211 gnd.n7210 19.3944
R15840 gnd.n7210 gnd.n318 19.3944
R15841 gnd.n7347 gnd.n318 19.3944
R15842 gnd.n7347 gnd.n319 19.3944
R15843 gnd.n7343 gnd.n319 19.3944
R15844 gnd.n7343 gnd.n7342 19.3944
R15845 gnd.n7342 gnd.n7341 19.3944
R15846 gnd.n7341 gnd.n325 19.3944
R15847 gnd.n7337 gnd.n325 19.3944
R15848 gnd.n7337 gnd.n7336 19.3944
R15849 gnd.n7336 gnd.n297 19.3944
R15850 gnd.n7360 gnd.n297 19.3944
R15851 gnd.n7360 gnd.n295 19.3944
R15852 gnd.n7364 gnd.n295 19.3944
R15853 gnd.n7364 gnd.n281 19.3944
R15854 gnd.n7376 gnd.n281 19.3944
R15855 gnd.n7376 gnd.n279 19.3944
R15856 gnd.n7380 gnd.n279 19.3944
R15857 gnd.n7380 gnd.n267 19.3944
R15858 gnd.n7392 gnd.n267 19.3944
R15859 gnd.n7392 gnd.n265 19.3944
R15860 gnd.n7396 gnd.n265 19.3944
R15861 gnd.n7396 gnd.n251 19.3944
R15862 gnd.n7408 gnd.n251 19.3944
R15863 gnd.n7408 gnd.n249 19.3944
R15864 gnd.n7412 gnd.n249 19.3944
R15865 gnd.n7412 gnd.n236 19.3944
R15866 gnd.n7424 gnd.n236 19.3944
R15867 gnd.n7424 gnd.n234 19.3944
R15868 gnd.n7428 gnd.n234 19.3944
R15869 gnd.n7428 gnd.n221 19.3944
R15870 gnd.n7440 gnd.n221 19.3944
R15871 gnd.n7440 gnd.n218 19.3944
R15872 gnd.n7512 gnd.n218 19.3944
R15873 gnd.n7512 gnd.n219 19.3944
R15874 gnd.n7508 gnd.n219 19.3944
R15875 gnd.n7508 gnd.n7507 19.3944
R15876 gnd.n7507 gnd.n7506 19.3944
R15877 gnd.n2028 gnd.n1115 19.3944
R15878 gnd.n2028 gnd.n1978 19.3944
R15879 gnd.n5397 gnd.n1978 19.3944
R15880 gnd.n5397 gnd.n5396 19.3944
R15881 gnd.n5396 gnd.n1981 19.3944
R15882 gnd.n5389 gnd.n1981 19.3944
R15883 gnd.n5389 gnd.n5388 19.3944
R15884 gnd.n5388 gnd.n1990 19.3944
R15885 gnd.n5381 gnd.n1990 19.3944
R15886 gnd.n5381 gnd.n5380 19.3944
R15887 gnd.n5380 gnd.n1998 19.3944
R15888 gnd.n5373 gnd.n1998 19.3944
R15889 gnd.n5373 gnd.n5372 19.3944
R15890 gnd.n5372 gnd.n2008 19.3944
R15891 gnd.n5365 gnd.n2008 19.3944
R15892 gnd.n5365 gnd.n5364 19.3944
R15893 gnd.n6342 gnd.n968 19.3944
R15894 gnd.n4355 gnd.n968 19.3944
R15895 gnd.n4355 gnd.n4353 19.3944
R15896 gnd.n4359 gnd.n4353 19.3944
R15897 gnd.n4359 gnd.n2150 19.3944
R15898 gnd.n4396 gnd.n2150 19.3944
R15899 gnd.n4396 gnd.n2148 19.3944
R15900 gnd.n4400 gnd.n2148 19.3944
R15901 gnd.n4400 gnd.n2146 19.3944
R15902 gnd.n4404 gnd.n2146 19.3944
R15903 gnd.n4404 gnd.n2144 19.3944
R15904 gnd.n4408 gnd.n2144 19.3944
R15905 gnd.n4408 gnd.n2129 19.3944
R15906 gnd.n4445 gnd.n2129 19.3944
R15907 gnd.n4445 gnd.n2127 19.3944
R15908 gnd.n4449 gnd.n2127 19.3944
R15909 gnd.n4449 gnd.n2125 19.3944
R15910 gnd.n4453 gnd.n2125 19.3944
R15911 gnd.n4453 gnd.n2123 19.3944
R15912 gnd.n4493 gnd.n2123 19.3944
R15913 gnd.n4493 gnd.n4492 19.3944
R15914 gnd.n4492 gnd.n4491 19.3944
R15915 gnd.n4491 gnd.n4459 19.3944
R15916 gnd.n4487 gnd.n4459 19.3944
R15917 gnd.n4487 gnd.n4486 19.3944
R15918 gnd.n4486 gnd.n4485 19.3944
R15919 gnd.n4485 gnd.n4465 19.3944
R15920 gnd.n4481 gnd.n4465 19.3944
R15921 gnd.n4481 gnd.n4480 19.3944
R15922 gnd.n4480 gnd.n4479 19.3944
R15923 gnd.n4479 gnd.n4471 19.3944
R15924 gnd.n4474 gnd.n4471 19.3944
R15925 gnd.n4474 gnd.n1950 19.3944
R15926 gnd.n5415 gnd.n1950 19.3944
R15927 gnd.n5415 gnd.n1948 19.3944
R15928 gnd.n5419 gnd.n1948 19.3944
R15929 gnd.n5419 gnd.n1936 19.3944
R15930 gnd.n5431 gnd.n1936 19.3944
R15931 gnd.n5431 gnd.n1934 19.3944
R15932 gnd.n5435 gnd.n1934 19.3944
R15933 gnd.n5435 gnd.n1924 19.3944
R15934 gnd.n5447 gnd.n1924 19.3944
R15935 gnd.n5447 gnd.n1922 19.3944
R15936 gnd.n5451 gnd.n1922 19.3944
R15937 gnd.n5451 gnd.n1911 19.3944
R15938 gnd.n5463 gnd.n1911 19.3944
R15939 gnd.n5463 gnd.n1909 19.3944
R15940 gnd.n5467 gnd.n1909 19.3944
R15941 gnd.n5467 gnd.n1898 19.3944
R15942 gnd.n5479 gnd.n1898 19.3944
R15943 gnd.n5479 gnd.n1896 19.3944
R15944 gnd.n5483 gnd.n1896 19.3944
R15945 gnd.n5483 gnd.n1885 19.3944
R15946 gnd.n5495 gnd.n1885 19.3944
R15947 gnd.n5495 gnd.n1883 19.3944
R15948 gnd.n5499 gnd.n1883 19.3944
R15949 gnd.n5499 gnd.n1872 19.3944
R15950 gnd.n5511 gnd.n1872 19.3944
R15951 gnd.n5511 gnd.n1870 19.3944
R15952 gnd.n5515 gnd.n1870 19.3944
R15953 gnd.n5515 gnd.n1857 19.3944
R15954 gnd.n5527 gnd.n1857 19.3944
R15955 gnd.n5527 gnd.n1855 19.3944
R15956 gnd.n5531 gnd.n1855 19.3944
R15957 gnd.n5531 gnd.n1844 19.3944
R15958 gnd.n5543 gnd.n1844 19.3944
R15959 gnd.n5543 gnd.n1842 19.3944
R15960 gnd.n5547 gnd.n1842 19.3944
R15961 gnd.n5547 gnd.n1831 19.3944
R15962 gnd.n5559 gnd.n1831 19.3944
R15963 gnd.n5559 gnd.n1829 19.3944
R15964 gnd.n5563 gnd.n1829 19.3944
R15965 gnd.n5563 gnd.n1816 19.3944
R15966 gnd.n5575 gnd.n1816 19.3944
R15967 gnd.n5575 gnd.n1814 19.3944
R15968 gnd.n5579 gnd.n1814 19.3944
R15969 gnd.n5579 gnd.n1801 19.3944
R15970 gnd.n5591 gnd.n1801 19.3944
R15971 gnd.n5591 gnd.n1799 19.3944
R15972 gnd.n5595 gnd.n1799 19.3944
R15973 gnd.n5595 gnd.n1788 19.3944
R15974 gnd.n5607 gnd.n1788 19.3944
R15975 gnd.n5607 gnd.n1786 19.3944
R15976 gnd.n5611 gnd.n1786 19.3944
R15977 gnd.n5611 gnd.n1774 19.3944
R15978 gnd.n5623 gnd.n1774 19.3944
R15979 gnd.n5623 gnd.n1772 19.3944
R15980 gnd.n5627 gnd.n1772 19.3944
R15981 gnd.n5627 gnd.n1759 19.3944
R15982 gnd.n5639 gnd.n1759 19.3944
R15983 gnd.n5639 gnd.n1757 19.3944
R15984 gnd.n5643 gnd.n1757 19.3944
R15985 gnd.n5643 gnd.n1746 19.3944
R15986 gnd.n5655 gnd.n1746 19.3944
R15987 gnd.n5655 gnd.n1744 19.3944
R15988 gnd.n5659 gnd.n1744 19.3944
R15989 gnd.n5659 gnd.n1731 19.3944
R15990 gnd.n5671 gnd.n1731 19.3944
R15991 gnd.n5671 gnd.n1729 19.3944
R15992 gnd.n5675 gnd.n1729 19.3944
R15993 gnd.n5675 gnd.n1718 19.3944
R15994 gnd.n5687 gnd.n1718 19.3944
R15995 gnd.n5687 gnd.n1716 19.3944
R15996 gnd.n5691 gnd.n1716 19.3944
R15997 gnd.n5691 gnd.n1704 19.3944
R15998 gnd.n5703 gnd.n1704 19.3944
R15999 gnd.n5703 gnd.n1702 19.3944
R16000 gnd.n5707 gnd.n1702 19.3944
R16001 gnd.n5707 gnd.n1690 19.3944
R16002 gnd.n5719 gnd.n1690 19.3944
R16003 gnd.n5719 gnd.n1688 19.3944
R16004 gnd.n5723 gnd.n1688 19.3944
R16005 gnd.n5723 gnd.n1677 19.3944
R16006 gnd.n5735 gnd.n1677 19.3944
R16007 gnd.n5735 gnd.n1675 19.3944
R16008 gnd.n5739 gnd.n1675 19.3944
R16009 gnd.n5739 gnd.n1664 19.3944
R16010 gnd.n5751 gnd.n1664 19.3944
R16011 gnd.n5751 gnd.n1662 19.3944
R16012 gnd.n5755 gnd.n1662 19.3944
R16013 gnd.n5755 gnd.n1651 19.3944
R16014 gnd.n5767 gnd.n1651 19.3944
R16015 gnd.n5767 gnd.n1649 19.3944
R16016 gnd.n5771 gnd.n1649 19.3944
R16017 gnd.n5771 gnd.n1637 19.3944
R16018 gnd.n5783 gnd.n1637 19.3944
R16019 gnd.n5783 gnd.n1635 19.3944
R16020 gnd.n5787 gnd.n1635 19.3944
R16021 gnd.n5787 gnd.n1624 19.3944
R16022 gnd.n5801 gnd.n1624 19.3944
R16023 gnd.n5801 gnd.n1622 19.3944
R16024 gnd.n5808 gnd.n1622 19.3944
R16025 gnd.n5808 gnd.n5807 19.3944
R16026 gnd.n5807 gnd.n1250 19.3944
R16027 gnd.n6098 gnd.n1250 19.3944
R16028 gnd.n6098 gnd.n6097 19.3944
R16029 gnd.n6097 gnd.n6096 19.3944
R16030 gnd.n6096 gnd.n1254 19.3944
R16031 gnd.n1445 gnd.n1254 19.3944
R16032 gnd.n1445 gnd.n1442 19.3944
R16033 gnd.n1449 gnd.n1442 19.3944
R16034 gnd.n1449 gnd.n1440 19.3944
R16035 gnd.n5863 gnd.n1440 19.3944
R16036 gnd.n5863 gnd.n1438 19.3944
R16037 gnd.n5869 gnd.n1438 19.3944
R16038 gnd.n5869 gnd.n5868 19.3944
R16039 gnd.n5868 gnd.n1412 19.3944
R16040 gnd.n5899 gnd.n1412 19.3944
R16041 gnd.n5899 gnd.n1410 19.3944
R16042 gnd.n5905 gnd.n1410 19.3944
R16043 gnd.n5905 gnd.n5904 19.3944
R16044 gnd.n5904 gnd.n1378 19.3944
R16045 gnd.n5960 gnd.n1378 19.3944
R16046 gnd.n5960 gnd.n1376 19.3944
R16047 gnd.n5976 gnd.n1376 19.3944
R16048 gnd.n5976 gnd.n5975 19.3944
R16049 gnd.n5975 gnd.n5974 19.3944
R16050 gnd.n5974 gnd.n5966 19.3944
R16051 gnd.n5970 gnd.n5966 19.3944
R16052 gnd.n5970 gnd.n411 19.3944
R16053 gnd.n7160 gnd.n411 19.3944
R16054 gnd.n7160 gnd.n7159 19.3944
R16055 gnd.n7159 gnd.n7158 19.3944
R16056 gnd.n7158 gnd.n415 19.3944
R16057 gnd.n7154 gnd.n415 19.3944
R16058 gnd.n7154 gnd.n7153 19.3944
R16059 gnd.n7153 gnd.n7152 19.3944
R16060 gnd.n6938 gnd.n544 19.3944
R16061 gnd.n6944 gnd.n544 19.3944
R16062 gnd.n6944 gnd.n542 19.3944
R16063 gnd.n6948 gnd.n542 19.3944
R16064 gnd.n6948 gnd.n538 19.3944
R16065 gnd.n6954 gnd.n538 19.3944
R16066 gnd.n6954 gnd.n536 19.3944
R16067 gnd.n6958 gnd.n536 19.3944
R16068 gnd.n6958 gnd.n532 19.3944
R16069 gnd.n6964 gnd.n532 19.3944
R16070 gnd.n6964 gnd.n530 19.3944
R16071 gnd.n6968 gnd.n530 19.3944
R16072 gnd.n6968 gnd.n526 19.3944
R16073 gnd.n6974 gnd.n526 19.3944
R16074 gnd.n6974 gnd.n524 19.3944
R16075 gnd.n6978 gnd.n524 19.3944
R16076 gnd.n6978 gnd.n520 19.3944
R16077 gnd.n6984 gnd.n520 19.3944
R16078 gnd.n6984 gnd.n518 19.3944
R16079 gnd.n6988 gnd.n518 19.3944
R16080 gnd.n6988 gnd.n514 19.3944
R16081 gnd.n6994 gnd.n514 19.3944
R16082 gnd.n6994 gnd.n512 19.3944
R16083 gnd.n6998 gnd.n512 19.3944
R16084 gnd.n6998 gnd.n508 19.3944
R16085 gnd.n7004 gnd.n508 19.3944
R16086 gnd.n7004 gnd.n506 19.3944
R16087 gnd.n7008 gnd.n506 19.3944
R16088 gnd.n7008 gnd.n502 19.3944
R16089 gnd.n7014 gnd.n502 19.3944
R16090 gnd.n7014 gnd.n500 19.3944
R16091 gnd.n7018 gnd.n500 19.3944
R16092 gnd.n7018 gnd.n496 19.3944
R16093 gnd.n7024 gnd.n496 19.3944
R16094 gnd.n7024 gnd.n494 19.3944
R16095 gnd.n7028 gnd.n494 19.3944
R16096 gnd.n7028 gnd.n490 19.3944
R16097 gnd.n7034 gnd.n490 19.3944
R16098 gnd.n7034 gnd.n488 19.3944
R16099 gnd.n7038 gnd.n488 19.3944
R16100 gnd.n7038 gnd.n484 19.3944
R16101 gnd.n7044 gnd.n484 19.3944
R16102 gnd.n7044 gnd.n482 19.3944
R16103 gnd.n7048 gnd.n482 19.3944
R16104 gnd.n7048 gnd.n478 19.3944
R16105 gnd.n7054 gnd.n478 19.3944
R16106 gnd.n7054 gnd.n476 19.3944
R16107 gnd.n7058 gnd.n476 19.3944
R16108 gnd.n7058 gnd.n472 19.3944
R16109 gnd.n7064 gnd.n472 19.3944
R16110 gnd.n7064 gnd.n470 19.3944
R16111 gnd.n7068 gnd.n470 19.3944
R16112 gnd.n7068 gnd.n466 19.3944
R16113 gnd.n7074 gnd.n466 19.3944
R16114 gnd.n7074 gnd.n464 19.3944
R16115 gnd.n7078 gnd.n464 19.3944
R16116 gnd.n7078 gnd.n460 19.3944
R16117 gnd.n7084 gnd.n460 19.3944
R16118 gnd.n7084 gnd.n458 19.3944
R16119 gnd.n7088 gnd.n458 19.3944
R16120 gnd.n7088 gnd.n454 19.3944
R16121 gnd.n7094 gnd.n454 19.3944
R16122 gnd.n7094 gnd.n452 19.3944
R16123 gnd.n7098 gnd.n452 19.3944
R16124 gnd.n7098 gnd.n448 19.3944
R16125 gnd.n7104 gnd.n448 19.3944
R16126 gnd.n7104 gnd.n446 19.3944
R16127 gnd.n7108 gnd.n446 19.3944
R16128 gnd.n7108 gnd.n442 19.3944
R16129 gnd.n7114 gnd.n442 19.3944
R16130 gnd.n7114 gnd.n440 19.3944
R16131 gnd.n7118 gnd.n440 19.3944
R16132 gnd.n7118 gnd.n436 19.3944
R16133 gnd.n7124 gnd.n436 19.3944
R16134 gnd.n7124 gnd.n434 19.3944
R16135 gnd.n7128 gnd.n434 19.3944
R16136 gnd.n7128 gnd.n430 19.3944
R16137 gnd.n7134 gnd.n430 19.3944
R16138 gnd.n7134 gnd.n428 19.3944
R16139 gnd.n7138 gnd.n428 19.3944
R16140 gnd.n7138 gnd.n424 19.3944
R16141 gnd.n7145 gnd.n424 19.3944
R16142 gnd.n7145 gnd.n422 19.3944
R16143 gnd.n7149 gnd.n422 19.3944
R16144 gnd.n6517 gnd.n795 19.3944
R16145 gnd.n6523 gnd.n795 19.3944
R16146 gnd.n6523 gnd.n793 19.3944
R16147 gnd.n6527 gnd.n793 19.3944
R16148 gnd.n6527 gnd.n789 19.3944
R16149 gnd.n6533 gnd.n789 19.3944
R16150 gnd.n6533 gnd.n787 19.3944
R16151 gnd.n6537 gnd.n787 19.3944
R16152 gnd.n6537 gnd.n783 19.3944
R16153 gnd.n6543 gnd.n783 19.3944
R16154 gnd.n6543 gnd.n781 19.3944
R16155 gnd.n6547 gnd.n781 19.3944
R16156 gnd.n6547 gnd.n777 19.3944
R16157 gnd.n6553 gnd.n777 19.3944
R16158 gnd.n6553 gnd.n775 19.3944
R16159 gnd.n6557 gnd.n775 19.3944
R16160 gnd.n6557 gnd.n771 19.3944
R16161 gnd.n6563 gnd.n771 19.3944
R16162 gnd.n6563 gnd.n769 19.3944
R16163 gnd.n6567 gnd.n769 19.3944
R16164 gnd.n6567 gnd.n765 19.3944
R16165 gnd.n6573 gnd.n765 19.3944
R16166 gnd.n6573 gnd.n763 19.3944
R16167 gnd.n6577 gnd.n763 19.3944
R16168 gnd.n6577 gnd.n759 19.3944
R16169 gnd.n6583 gnd.n759 19.3944
R16170 gnd.n6583 gnd.n757 19.3944
R16171 gnd.n6587 gnd.n757 19.3944
R16172 gnd.n6587 gnd.n753 19.3944
R16173 gnd.n6593 gnd.n753 19.3944
R16174 gnd.n6593 gnd.n751 19.3944
R16175 gnd.n6597 gnd.n751 19.3944
R16176 gnd.n6597 gnd.n747 19.3944
R16177 gnd.n6603 gnd.n747 19.3944
R16178 gnd.n6603 gnd.n745 19.3944
R16179 gnd.n6607 gnd.n745 19.3944
R16180 gnd.n6607 gnd.n741 19.3944
R16181 gnd.n6613 gnd.n741 19.3944
R16182 gnd.n6613 gnd.n739 19.3944
R16183 gnd.n6617 gnd.n739 19.3944
R16184 gnd.n6617 gnd.n735 19.3944
R16185 gnd.n6623 gnd.n735 19.3944
R16186 gnd.n6623 gnd.n733 19.3944
R16187 gnd.n6627 gnd.n733 19.3944
R16188 gnd.n6627 gnd.n729 19.3944
R16189 gnd.n6633 gnd.n729 19.3944
R16190 gnd.n6633 gnd.n727 19.3944
R16191 gnd.n6637 gnd.n727 19.3944
R16192 gnd.n6637 gnd.n723 19.3944
R16193 gnd.n6643 gnd.n723 19.3944
R16194 gnd.n6643 gnd.n721 19.3944
R16195 gnd.n6647 gnd.n721 19.3944
R16196 gnd.n6647 gnd.n717 19.3944
R16197 gnd.n6653 gnd.n717 19.3944
R16198 gnd.n6653 gnd.n715 19.3944
R16199 gnd.n6657 gnd.n715 19.3944
R16200 gnd.n6657 gnd.n711 19.3944
R16201 gnd.n6663 gnd.n711 19.3944
R16202 gnd.n6663 gnd.n709 19.3944
R16203 gnd.n6667 gnd.n709 19.3944
R16204 gnd.n6667 gnd.n705 19.3944
R16205 gnd.n6673 gnd.n705 19.3944
R16206 gnd.n6673 gnd.n703 19.3944
R16207 gnd.n6677 gnd.n703 19.3944
R16208 gnd.n6677 gnd.n699 19.3944
R16209 gnd.n6683 gnd.n699 19.3944
R16210 gnd.n6683 gnd.n697 19.3944
R16211 gnd.n6687 gnd.n697 19.3944
R16212 gnd.n6687 gnd.n693 19.3944
R16213 gnd.n6693 gnd.n693 19.3944
R16214 gnd.n6693 gnd.n691 19.3944
R16215 gnd.n6697 gnd.n691 19.3944
R16216 gnd.n6697 gnd.n687 19.3944
R16217 gnd.n6703 gnd.n687 19.3944
R16218 gnd.n6703 gnd.n685 19.3944
R16219 gnd.n6707 gnd.n685 19.3944
R16220 gnd.n6707 gnd.n681 19.3944
R16221 gnd.n6713 gnd.n681 19.3944
R16222 gnd.n6713 gnd.n679 19.3944
R16223 gnd.n6717 gnd.n679 19.3944
R16224 gnd.n6717 gnd.n675 19.3944
R16225 gnd.n6723 gnd.n675 19.3944
R16226 gnd.n6723 gnd.n673 19.3944
R16227 gnd.n6727 gnd.n673 19.3944
R16228 gnd.n6727 gnd.n669 19.3944
R16229 gnd.n6733 gnd.n669 19.3944
R16230 gnd.n6733 gnd.n667 19.3944
R16231 gnd.n6737 gnd.n667 19.3944
R16232 gnd.n6737 gnd.n663 19.3944
R16233 gnd.n6743 gnd.n663 19.3944
R16234 gnd.n6743 gnd.n661 19.3944
R16235 gnd.n6747 gnd.n661 19.3944
R16236 gnd.n6747 gnd.n657 19.3944
R16237 gnd.n6753 gnd.n657 19.3944
R16238 gnd.n6753 gnd.n655 19.3944
R16239 gnd.n6757 gnd.n655 19.3944
R16240 gnd.n6757 gnd.n651 19.3944
R16241 gnd.n6763 gnd.n651 19.3944
R16242 gnd.n6763 gnd.n649 19.3944
R16243 gnd.n6767 gnd.n649 19.3944
R16244 gnd.n6767 gnd.n645 19.3944
R16245 gnd.n6773 gnd.n645 19.3944
R16246 gnd.n6773 gnd.n643 19.3944
R16247 gnd.n6777 gnd.n643 19.3944
R16248 gnd.n6777 gnd.n639 19.3944
R16249 gnd.n6783 gnd.n639 19.3944
R16250 gnd.n6783 gnd.n637 19.3944
R16251 gnd.n6787 gnd.n637 19.3944
R16252 gnd.n6787 gnd.n633 19.3944
R16253 gnd.n6793 gnd.n633 19.3944
R16254 gnd.n6793 gnd.n631 19.3944
R16255 gnd.n6797 gnd.n631 19.3944
R16256 gnd.n6797 gnd.n627 19.3944
R16257 gnd.n6803 gnd.n627 19.3944
R16258 gnd.n6803 gnd.n625 19.3944
R16259 gnd.n6807 gnd.n625 19.3944
R16260 gnd.n6807 gnd.n621 19.3944
R16261 gnd.n6813 gnd.n621 19.3944
R16262 gnd.n6813 gnd.n619 19.3944
R16263 gnd.n6817 gnd.n619 19.3944
R16264 gnd.n6817 gnd.n615 19.3944
R16265 gnd.n6823 gnd.n615 19.3944
R16266 gnd.n6823 gnd.n613 19.3944
R16267 gnd.n6827 gnd.n613 19.3944
R16268 gnd.n6827 gnd.n609 19.3944
R16269 gnd.n6833 gnd.n609 19.3944
R16270 gnd.n6833 gnd.n607 19.3944
R16271 gnd.n6837 gnd.n607 19.3944
R16272 gnd.n6837 gnd.n603 19.3944
R16273 gnd.n6843 gnd.n603 19.3944
R16274 gnd.n6843 gnd.n601 19.3944
R16275 gnd.n6847 gnd.n601 19.3944
R16276 gnd.n6847 gnd.n597 19.3944
R16277 gnd.n6853 gnd.n597 19.3944
R16278 gnd.n6853 gnd.n595 19.3944
R16279 gnd.n6857 gnd.n595 19.3944
R16280 gnd.n6857 gnd.n591 19.3944
R16281 gnd.n6863 gnd.n591 19.3944
R16282 gnd.n6863 gnd.n589 19.3944
R16283 gnd.n6867 gnd.n589 19.3944
R16284 gnd.n6867 gnd.n585 19.3944
R16285 gnd.n6873 gnd.n585 19.3944
R16286 gnd.n6873 gnd.n583 19.3944
R16287 gnd.n6877 gnd.n583 19.3944
R16288 gnd.n6877 gnd.n579 19.3944
R16289 gnd.n6883 gnd.n579 19.3944
R16290 gnd.n6883 gnd.n577 19.3944
R16291 gnd.n6887 gnd.n577 19.3944
R16292 gnd.n6887 gnd.n573 19.3944
R16293 gnd.n6893 gnd.n573 19.3944
R16294 gnd.n6893 gnd.n571 19.3944
R16295 gnd.n6897 gnd.n571 19.3944
R16296 gnd.n6897 gnd.n567 19.3944
R16297 gnd.n6903 gnd.n567 19.3944
R16298 gnd.n6903 gnd.n565 19.3944
R16299 gnd.n6907 gnd.n565 19.3944
R16300 gnd.n6907 gnd.n561 19.3944
R16301 gnd.n6913 gnd.n561 19.3944
R16302 gnd.n6913 gnd.n559 19.3944
R16303 gnd.n6917 gnd.n559 19.3944
R16304 gnd.n6917 gnd.n555 19.3944
R16305 gnd.n6923 gnd.n555 19.3944
R16306 gnd.n6923 gnd.n553 19.3944
R16307 gnd.n6928 gnd.n553 19.3944
R16308 gnd.n6928 gnd.n549 19.3944
R16309 gnd.n6934 gnd.n549 19.3944
R16310 gnd.n6935 gnd.n6934 19.3944
R16311 gnd.n6089 gnd.n6088 19.3944
R16312 gnd.n6088 gnd.n6087 19.3944
R16313 gnd.n6087 gnd.n6086 19.3944
R16314 gnd.n6086 gnd.n6084 19.3944
R16315 gnd.n6084 gnd.n6081 19.3944
R16316 gnd.n6081 gnd.n6080 19.3944
R16317 gnd.n6080 gnd.n6077 19.3944
R16318 gnd.n6077 gnd.n6076 19.3944
R16319 gnd.n6076 gnd.n6073 19.3944
R16320 gnd.n6073 gnd.n6072 19.3944
R16321 gnd.n6072 gnd.n6069 19.3944
R16322 gnd.n6069 gnd.n6068 19.3944
R16323 gnd.n6068 gnd.n6065 19.3944
R16324 gnd.n6065 gnd.n6064 19.3944
R16325 gnd.n6064 gnd.n6061 19.3944
R16326 gnd.n6059 gnd.n6056 19.3944
R16327 gnd.n6056 gnd.n6055 19.3944
R16328 gnd.n6055 gnd.n6052 19.3944
R16329 gnd.n6052 gnd.n6051 19.3944
R16330 gnd.n6051 gnd.n6048 19.3944
R16331 gnd.n6048 gnd.n6047 19.3944
R16332 gnd.n6047 gnd.n6044 19.3944
R16333 gnd.n6044 gnd.n6043 19.3944
R16334 gnd.n6043 gnd.n6040 19.3944
R16335 gnd.n6040 gnd.n6039 19.3944
R16336 gnd.n6039 gnd.n6036 19.3944
R16337 gnd.n6036 gnd.n6035 19.3944
R16338 gnd.n6035 gnd.n6032 19.3944
R16339 gnd.n6032 gnd.n6031 19.3944
R16340 gnd.n6031 gnd.n6028 19.3944
R16341 gnd.n6028 gnd.n6027 19.3944
R16342 gnd.n6027 gnd.n6024 19.3944
R16343 gnd.n6024 gnd.n6023 19.3944
R16344 gnd.n1455 gnd.n1335 19.3944
R16345 gnd.n1455 gnd.n1454 19.3944
R16346 gnd.n1473 gnd.n1454 19.3944
R16347 gnd.n1473 gnd.n1472 19.3944
R16348 gnd.n1472 gnd.n1471 19.3944
R16349 gnd.n1471 gnd.n1469 19.3944
R16350 gnd.n1469 gnd.n1468 19.3944
R16351 gnd.n1468 gnd.n1466 19.3944
R16352 gnd.n1466 gnd.n1465 19.3944
R16353 gnd.n1465 gnd.n1391 19.3944
R16354 gnd.n5921 gnd.n1391 19.3944
R16355 gnd.n5921 gnd.n1389 19.3944
R16356 gnd.n5925 gnd.n1389 19.3944
R16357 gnd.n5926 gnd.n5925 19.3944
R16358 gnd.n5928 gnd.n5926 19.3944
R16359 gnd.n5928 gnd.n1387 19.3944
R16360 gnd.n5934 gnd.n1387 19.3944
R16361 gnd.n5934 gnd.n5933 19.3944
R16362 gnd.n5933 gnd.n388 19.3944
R16363 gnd.n7184 gnd.n388 19.3944
R16364 gnd.n7184 gnd.n386 19.3944
R16365 gnd.n7194 gnd.n386 19.3944
R16366 gnd.n7194 gnd.n7193 19.3944
R16367 gnd.n7193 gnd.n7192 19.3944
R16368 gnd.n7192 gnd.n354 19.3944
R16369 gnd.n7229 gnd.n354 19.3944
R16370 gnd.n7229 gnd.n352 19.3944
R16371 gnd.n7240 gnd.n352 19.3944
R16372 gnd.n7240 gnd.n7239 19.3944
R16373 gnd.n7239 gnd.n7238 19.3944
R16374 gnd.n7238 gnd.n7236 19.3944
R16375 gnd.n7236 gnd.n338 19.3944
R16376 gnd.n7259 gnd.n338 19.3944
R16377 gnd.n7259 gnd.n336 19.3944
R16378 gnd.n7328 gnd.n336 19.3944
R16379 gnd.n7328 gnd.n7327 19.3944
R16380 gnd.n7327 gnd.n7326 19.3944
R16381 gnd.n7326 gnd.n7324 19.3944
R16382 gnd.n7324 gnd.n7323 19.3944
R16383 gnd.n7323 gnd.n7321 19.3944
R16384 gnd.n7321 gnd.n7320 19.3944
R16385 gnd.n7320 gnd.n7318 19.3944
R16386 gnd.n7318 gnd.n7317 19.3944
R16387 gnd.n7317 gnd.n7315 19.3944
R16388 gnd.n7315 gnd.n7314 19.3944
R16389 gnd.n7314 gnd.n7312 19.3944
R16390 gnd.n7312 gnd.n7311 19.3944
R16391 gnd.n7311 gnd.n7309 19.3944
R16392 gnd.n7309 gnd.n7308 19.3944
R16393 gnd.n7308 gnd.n7306 19.3944
R16394 gnd.n7306 gnd.n7305 19.3944
R16395 gnd.n7305 gnd.n7303 19.3944
R16396 gnd.n7303 gnd.n7302 19.3944
R16397 gnd.n7302 gnd.n7300 19.3944
R16398 gnd.n7300 gnd.n7299 19.3944
R16399 gnd.n7299 gnd.n7297 19.3944
R16400 gnd.n7297 gnd.n7296 19.3944
R16401 gnd.n7296 gnd.n7294 19.3944
R16402 gnd.n7294 gnd.n7293 19.3944
R16403 gnd.n7293 gnd.n7291 19.3944
R16404 gnd.n7291 gnd.n7290 19.3944
R16405 gnd.n7290 gnd.n204 19.3944
R16406 gnd.n7525 gnd.n204 19.3944
R16407 gnd.n7526 gnd.n7525 19.3944
R16408 gnd.n7564 gnd.n165 19.3944
R16409 gnd.n7559 gnd.n165 19.3944
R16410 gnd.n7559 gnd.n7558 19.3944
R16411 gnd.n7558 gnd.n7557 19.3944
R16412 gnd.n7557 gnd.n172 19.3944
R16413 gnd.n7552 gnd.n172 19.3944
R16414 gnd.n7552 gnd.n7551 19.3944
R16415 gnd.n7551 gnd.n7550 19.3944
R16416 gnd.n7550 gnd.n179 19.3944
R16417 gnd.n7545 gnd.n179 19.3944
R16418 gnd.n7545 gnd.n7544 19.3944
R16419 gnd.n7544 gnd.n7543 19.3944
R16420 gnd.n7543 gnd.n186 19.3944
R16421 gnd.n7538 gnd.n186 19.3944
R16422 gnd.n7538 gnd.n7537 19.3944
R16423 gnd.n7537 gnd.n7536 19.3944
R16424 gnd.n7536 gnd.n193 19.3944
R16425 gnd.n7531 gnd.n193 19.3944
R16426 gnd.n7597 gnd.n7596 19.3944
R16427 gnd.n7596 gnd.n7595 19.3944
R16428 gnd.n7595 gnd.n137 19.3944
R16429 gnd.n7590 gnd.n137 19.3944
R16430 gnd.n7590 gnd.n7589 19.3944
R16431 gnd.n7589 gnd.n7588 19.3944
R16432 gnd.n7588 gnd.n144 19.3944
R16433 gnd.n7583 gnd.n144 19.3944
R16434 gnd.n7583 gnd.n7582 19.3944
R16435 gnd.n7582 gnd.n7581 19.3944
R16436 gnd.n7581 gnd.n151 19.3944
R16437 gnd.n7576 gnd.n151 19.3944
R16438 gnd.n7576 gnd.n7575 19.3944
R16439 gnd.n7575 gnd.n7574 19.3944
R16440 gnd.n7574 gnd.n158 19.3944
R16441 gnd.n7569 gnd.n158 19.3944
R16442 gnd.n7569 gnd.n7568 19.3944
R16443 gnd.n5849 gnd.n5844 19.3944
R16444 gnd.n5849 gnd.n5848 19.3944
R16445 gnd.n5848 gnd.n1429 19.3944
R16446 gnd.n5874 gnd.n1429 19.3944
R16447 gnd.n5874 gnd.n1427 19.3944
R16448 gnd.n5880 gnd.n1427 19.3944
R16449 gnd.n5880 gnd.n5879 19.3944
R16450 gnd.n5879 gnd.n1402 19.3944
R16451 gnd.n5911 gnd.n1402 19.3944
R16452 gnd.n5911 gnd.n1400 19.3944
R16453 gnd.n5917 gnd.n1400 19.3944
R16454 gnd.n5917 gnd.n5916 19.3944
R16455 gnd.n5916 gnd.n1368 19.3944
R16456 gnd.n5981 gnd.n1368 19.3944
R16457 gnd.n5981 gnd.n1366 19.3944
R16458 gnd.n5985 gnd.n1366 19.3944
R16459 gnd.n5985 gnd.n397 19.3944
R16460 gnd.n7174 gnd.n397 19.3944
R16461 gnd.n7174 gnd.n395 19.3944
R16462 gnd.n7180 gnd.n395 19.3944
R16463 gnd.n7180 gnd.n7179 19.3944
R16464 gnd.n7179 gnd.n364 19.3944
R16465 gnd.n7220 gnd.n364 19.3944
R16466 gnd.n7220 gnd.n362 19.3944
R16467 gnd.n7224 gnd.n362 19.3944
R16468 gnd.n7225 gnd.n7224 19.3944
R16469 gnd.n7225 gnd.n309 19.3944
R16470 gnd.n7352 gnd.n7351 19.3944
R16471 gnd.n342 gnd.n341 19.3944
R16472 gnd.n7255 gnd.n7254 19.3944
R16473 gnd.n332 gnd.n331 19.3944
R16474 gnd.n7332 gnd.n302 19.3944
R16475 gnd.n7356 gnd.n302 19.3944
R16476 gnd.n7356 gnd.n288 19.3944
R16477 gnd.n7368 gnd.n288 19.3944
R16478 gnd.n7368 gnd.n286 19.3944
R16479 gnd.n7372 gnd.n286 19.3944
R16480 gnd.n7372 gnd.n274 19.3944
R16481 gnd.n7384 gnd.n274 19.3944
R16482 gnd.n7384 gnd.n272 19.3944
R16483 gnd.n7388 gnd.n272 19.3944
R16484 gnd.n7388 gnd.n258 19.3944
R16485 gnd.n7400 gnd.n258 19.3944
R16486 gnd.n7400 gnd.n256 19.3944
R16487 gnd.n7404 gnd.n256 19.3944
R16488 gnd.n7404 gnd.n243 19.3944
R16489 gnd.n7416 gnd.n243 19.3944
R16490 gnd.n7416 gnd.n241 19.3944
R16491 gnd.n7420 gnd.n241 19.3944
R16492 gnd.n7420 gnd.n227 19.3944
R16493 gnd.n7432 gnd.n227 19.3944
R16494 gnd.n7432 gnd.n225 19.3944
R16495 gnd.n7436 gnd.n225 19.3944
R16496 gnd.n7436 gnd.n211 19.3944
R16497 gnd.n7516 gnd.n211 19.3944
R16498 gnd.n7516 gnd.n209 19.3944
R16499 gnd.n7520 gnd.n209 19.3944
R16500 gnd.n7520 gnd.n132 19.3944
R16501 gnd.n7600 gnd.n132 19.3944
R16502 gnd.n4174 gnd.n4173 19.3944
R16503 gnd.n4173 gnd.n3960 19.3944
R16504 gnd.n4168 gnd.n3960 19.3944
R16505 gnd.n4168 gnd.n4167 19.3944
R16506 gnd.n4167 gnd.n3965 19.3944
R16507 gnd.n4162 gnd.n3965 19.3944
R16508 gnd.n4162 gnd.n4161 19.3944
R16509 gnd.n4161 gnd.n4160 19.3944
R16510 gnd.n4160 gnd.n3971 19.3944
R16511 gnd.n4154 gnd.n3971 19.3944
R16512 gnd.n4154 gnd.n4153 19.3944
R16513 gnd.n4153 gnd.n4152 19.3944
R16514 gnd.n4152 gnd.n3977 19.3944
R16515 gnd.n4146 gnd.n3977 19.3944
R16516 gnd.n4146 gnd.n4145 19.3944
R16517 gnd.n4145 gnd.n4144 19.3944
R16518 gnd.n4144 gnd.n3983 19.3944
R16519 gnd.n4138 gnd.n4137 19.3944
R16520 gnd.n4137 gnd.n4136 19.3944
R16521 gnd.n4136 gnd.n3992 19.3944
R16522 gnd.n4130 gnd.n3992 19.3944
R16523 gnd.n4130 gnd.n4129 19.3944
R16524 gnd.n4129 gnd.n4128 19.3944
R16525 gnd.n4128 gnd.n3998 19.3944
R16526 gnd.n4122 gnd.n3998 19.3944
R16527 gnd.n4122 gnd.n4121 19.3944
R16528 gnd.n4121 gnd.n4120 19.3944
R16529 gnd.n4120 gnd.n4004 19.3944
R16530 gnd.n4114 gnd.n4004 19.3944
R16531 gnd.n4114 gnd.n4113 19.3944
R16532 gnd.n4113 gnd.n4112 19.3944
R16533 gnd.n4112 gnd.n4010 19.3944
R16534 gnd.n4106 gnd.n4010 19.3944
R16535 gnd.n4106 gnd.n4105 19.3944
R16536 gnd.n4105 gnd.n4104 19.3944
R16537 gnd.n4181 gnd.n2316 19.3944
R16538 gnd.n4185 gnd.n2316 19.3944
R16539 gnd.n4185 gnd.n2303 19.3944
R16540 gnd.n4197 gnd.n2303 19.3944
R16541 gnd.n4197 gnd.n2301 19.3944
R16542 gnd.n4201 gnd.n2301 19.3944
R16543 gnd.n4201 gnd.n2286 19.3944
R16544 gnd.n4213 gnd.n2286 19.3944
R16545 gnd.n4213 gnd.n2284 19.3944
R16546 gnd.n4217 gnd.n2284 19.3944
R16547 gnd.n4217 gnd.n2271 19.3944
R16548 gnd.n4229 gnd.n2271 19.3944
R16549 gnd.n4229 gnd.n2269 19.3944
R16550 gnd.n4233 gnd.n2269 19.3944
R16551 gnd.n4233 gnd.n2254 19.3944
R16552 gnd.n4245 gnd.n2254 19.3944
R16553 gnd.n4245 gnd.n2252 19.3944
R16554 gnd.n4249 gnd.n2252 19.3944
R16555 gnd.n4249 gnd.n2239 19.3944
R16556 gnd.n4261 gnd.n2239 19.3944
R16557 gnd.n4261 gnd.n2237 19.3944
R16558 gnd.n4265 gnd.n2237 19.3944
R16559 gnd.n4265 gnd.n2222 19.3944
R16560 gnd.n4278 gnd.n2222 19.3944
R16561 gnd.n4278 gnd.n2220 19.3944
R16562 gnd.n4282 gnd.n2220 19.3944
R16563 gnd.n4282 gnd.n2208 19.3944
R16564 gnd.n4294 gnd.n2208 19.3944
R16565 gnd.n4294 gnd.n2206 19.3944
R16566 gnd.n4299 gnd.n2206 19.3944
R16567 gnd.n4299 gnd.n4298 19.3944
R16568 gnd.n4298 gnd.n2183 19.3944
R16569 gnd.n2183 gnd.n2181 19.3944
R16570 gnd.n4326 gnd.n2181 19.3944
R16571 gnd.n4326 gnd.n4325 19.3944
R16572 gnd.n4325 gnd.n4324 19.3944
R16573 gnd.n4324 gnd.n4323 19.3944
R16574 gnd.n4323 gnd.n4321 19.3944
R16575 gnd.n4321 gnd.n989 19.3944
R16576 gnd.n6331 gnd.n989 19.3944
R16577 gnd.n6331 gnd.n6330 19.3944
R16578 gnd.n6330 gnd.n6329 19.3944
R16579 gnd.n6329 gnd.n993 19.3944
R16580 gnd.n6319 gnd.n993 19.3944
R16581 gnd.n6319 gnd.n6318 19.3944
R16582 gnd.n6318 gnd.n6317 19.3944
R16583 gnd.n6317 gnd.n1013 19.3944
R16584 gnd.n6307 gnd.n1013 19.3944
R16585 gnd.n6307 gnd.n6306 19.3944
R16586 gnd.n6306 gnd.n6305 19.3944
R16587 gnd.n6305 gnd.n1035 19.3944
R16588 gnd.n6295 gnd.n1035 19.3944
R16589 gnd.n6295 gnd.n6294 19.3944
R16590 gnd.n6294 gnd.n6293 19.3944
R16591 gnd.n6293 gnd.n1055 19.3944
R16592 gnd.n6283 gnd.n1055 19.3944
R16593 gnd.n6283 gnd.n6282 19.3944
R16594 gnd.n6282 gnd.n6281 19.3944
R16595 gnd.n6281 gnd.n1077 19.3944
R16596 gnd.n6271 gnd.n1077 19.3944
R16597 gnd.n6271 gnd.n6270 19.3944
R16598 gnd.n6270 gnd.n6269 19.3944
R16599 gnd.n6269 gnd.n1098 19.3944
R16600 gnd.n6259 gnd.n1098 19.3944
R16601 gnd.n3817 gnd.n3816 19.3944
R16602 gnd.n3822 gnd.n3817 19.3944
R16603 gnd.n3822 gnd.n3814 19.3944
R16604 gnd.n3826 gnd.n3814 19.3944
R16605 gnd.n3826 gnd.n3812 19.3944
R16606 gnd.n3832 gnd.n3812 19.3944
R16607 gnd.n3832 gnd.n3810 19.3944
R16608 gnd.n3836 gnd.n3810 19.3944
R16609 gnd.n3836 gnd.n3808 19.3944
R16610 gnd.n3842 gnd.n3808 19.3944
R16611 gnd.n3842 gnd.n3806 19.3944
R16612 gnd.n3846 gnd.n3806 19.3944
R16613 gnd.n3846 gnd.n3804 19.3944
R16614 gnd.n3852 gnd.n3804 19.3944
R16615 gnd.n3852 gnd.n3802 19.3944
R16616 gnd.n3856 gnd.n3802 19.3944
R16617 gnd.n3955 gnd.n3796 19.3944
R16618 gnd.n3955 gnd.n3954 19.3944
R16619 gnd.n3954 gnd.n3953 19.3944
R16620 gnd.n3953 gnd.n3951 19.3944
R16621 gnd.n3951 gnd.n3950 19.3944
R16622 gnd.n3950 gnd.n3948 19.3944
R16623 gnd.n3948 gnd.n3947 19.3944
R16624 gnd.n3947 gnd.n3945 19.3944
R16625 gnd.n3945 gnd.n3944 19.3944
R16626 gnd.n3944 gnd.n3942 19.3944
R16627 gnd.n3942 gnd.n3941 19.3944
R16628 gnd.n3941 gnd.n3939 19.3944
R16629 gnd.n3939 gnd.n3938 19.3944
R16630 gnd.n3938 gnd.n3936 19.3944
R16631 gnd.n3936 gnd.n3935 19.3944
R16632 gnd.n3935 gnd.n3933 19.3944
R16633 gnd.n3933 gnd.n3932 19.3944
R16634 gnd.n3932 gnd.n3930 19.3944
R16635 gnd.n3930 gnd.n3929 19.3944
R16636 gnd.n3929 gnd.n3927 19.3944
R16637 gnd.n3927 gnd.n3926 19.3944
R16638 gnd.n3926 gnd.n3924 19.3944
R16639 gnd.n3924 gnd.n3923 19.3944
R16640 gnd.n3923 gnd.n3921 19.3944
R16641 gnd.n3921 gnd.n3920 19.3944
R16642 gnd.n3920 gnd.n3918 19.3944
R16643 gnd.n3918 gnd.n3917 19.3944
R16644 gnd.n3917 gnd.n3915 19.3944
R16645 gnd.n3915 gnd.n3914 19.3944
R16646 gnd.n3914 gnd.n3912 19.3944
R16647 gnd.n3912 gnd.n3911 19.3944
R16648 gnd.n3911 gnd.n3909 19.3944
R16649 gnd.n3909 gnd.n3896 19.3944
R16650 gnd.n3905 gnd.n3896 19.3944
R16651 gnd.n3905 gnd.n3904 19.3944
R16652 gnd.n3904 gnd.n3903 19.3944
R16653 gnd.n3903 gnd.n3900 19.3944
R16654 gnd.n3900 gnd.n2165 19.3944
R16655 gnd.n4346 gnd.n2165 19.3944
R16656 gnd.n4346 gnd.n2163 19.3944
R16657 gnd.n4350 gnd.n2163 19.3944
R16658 gnd.n4350 gnd.n2153 19.3944
R16659 gnd.n4391 gnd.n2153 19.3944
R16660 gnd.n4391 gnd.n2154 19.3944
R16661 gnd.n4387 gnd.n2154 19.3944
R16662 gnd.n4387 gnd.n4386 19.3944
R16663 gnd.n4386 gnd.n4385 19.3944
R16664 gnd.n4385 gnd.n4380 19.3944
R16665 gnd.n4381 gnd.n4380 19.3944
R16666 gnd.n4381 gnd.n2132 19.3944
R16667 gnd.n4440 gnd.n2132 19.3944
R16668 gnd.n4440 gnd.n2133 19.3944
R16669 gnd.n4436 gnd.n2133 19.3944
R16670 gnd.n4436 gnd.n4435 19.3944
R16671 gnd.n4435 gnd.n4434 19.3944
R16672 gnd.n4434 gnd.n2119 19.3944
R16673 gnd.n4498 gnd.n2119 19.3944
R16674 gnd.n4498 gnd.n2117 19.3944
R16675 gnd.n4502 gnd.n2117 19.3944
R16676 gnd.n4502 gnd.n2113 19.3944
R16677 gnd.n4515 gnd.n2113 19.3944
R16678 gnd.n4515 gnd.n2110 19.3944
R16679 gnd.n4551 gnd.n2110 19.3944
R16680 gnd.n4551 gnd.n2111 19.3944
R16681 gnd.n4095 gnd.n4094 19.3944
R16682 gnd.n4094 gnd.n4093 19.3944
R16683 gnd.n4093 gnd.n4092 19.3944
R16684 gnd.n4092 gnd.n4090 19.3944
R16685 gnd.n4090 gnd.n4089 19.3944
R16686 gnd.n4089 gnd.n4087 19.3944
R16687 gnd.n4087 gnd.n4086 19.3944
R16688 gnd.n4086 gnd.n4084 19.3944
R16689 gnd.n4084 gnd.n4083 19.3944
R16690 gnd.n4083 gnd.n4081 19.3944
R16691 gnd.n4081 gnd.n4080 19.3944
R16692 gnd.n4080 gnd.n4078 19.3944
R16693 gnd.n4078 gnd.n4077 19.3944
R16694 gnd.n4077 gnd.n4075 19.3944
R16695 gnd.n4075 gnd.n4074 19.3944
R16696 gnd.n4074 gnd.n4072 19.3944
R16697 gnd.n4072 gnd.n4071 19.3944
R16698 gnd.n4071 gnd.n4069 19.3944
R16699 gnd.n4069 gnd.n4068 19.3944
R16700 gnd.n4068 gnd.n4066 19.3944
R16701 gnd.n4066 gnd.n4065 19.3944
R16702 gnd.n4065 gnd.n4063 19.3944
R16703 gnd.n4063 gnd.n4062 19.3944
R16704 gnd.n4062 gnd.n4060 19.3944
R16705 gnd.n4060 gnd.n4059 19.3944
R16706 gnd.n4059 gnd.n4057 19.3944
R16707 gnd.n4057 gnd.n4056 19.3944
R16708 gnd.n4056 gnd.n4054 19.3944
R16709 gnd.n4054 gnd.n4053 19.3944
R16710 gnd.n4053 gnd.n4051 19.3944
R16711 gnd.n4051 gnd.n2186 19.3944
R16712 gnd.n4311 gnd.n2186 19.3944
R16713 gnd.n4311 gnd.n2191 19.3944
R16714 gnd.n2191 gnd.n2190 19.3944
R16715 gnd.n2190 gnd.n2189 19.3944
R16716 gnd.n2189 gnd.n2168 19.3944
R16717 gnd.n4338 gnd.n2168 19.3944
R16718 gnd.n4338 gnd.n2166 19.3944
R16719 gnd.n4342 gnd.n2166 19.3944
R16720 gnd.n4342 gnd.n2162 19.3944
R16721 gnd.n4364 gnd.n2162 19.3944
R16722 gnd.n4364 gnd.n2160 19.3944
R16723 gnd.n4368 gnd.n2160 19.3944
R16724 gnd.n4369 gnd.n4368 19.3944
R16725 gnd.n4372 gnd.n4369 19.3944
R16726 gnd.n4372 gnd.n2158 19.3944
R16727 gnd.n4376 gnd.n2158 19.3944
R16728 gnd.n4376 gnd.n2141 19.3944
R16729 gnd.n4413 gnd.n2141 19.3944
R16730 gnd.n4413 gnd.n2139 19.3944
R16731 gnd.n4417 gnd.n2139 19.3944
R16732 gnd.n4418 gnd.n4417 19.3944
R16733 gnd.n4421 gnd.n4418 19.3944
R16734 gnd.n4421 gnd.n2137 19.3944
R16735 gnd.n4429 gnd.n2137 19.3944
R16736 gnd.n4429 gnd.n4428 19.3944
R16737 gnd.n4428 gnd.n4427 19.3944
R16738 gnd.n4427 gnd.n2116 19.3944
R16739 gnd.n4506 gnd.n2116 19.3944
R16740 gnd.n4506 gnd.n2114 19.3944
R16741 gnd.n4511 gnd.n2114 19.3944
R16742 gnd.n4511 gnd.n2108 19.3944
R16743 gnd.n4555 gnd.n2108 19.3944
R16744 gnd.n4556 gnd.n4555 19.3944
R16745 gnd.n4598 gnd.n2082 19.3944
R16746 gnd.n4598 gnd.n4595 19.3944
R16747 gnd.n4595 gnd.n4592 19.3944
R16748 gnd.n4592 gnd.n4591 19.3944
R16749 gnd.n4591 gnd.n4588 19.3944
R16750 gnd.n4588 gnd.n4587 19.3944
R16751 gnd.n4587 gnd.n4584 19.3944
R16752 gnd.n4584 gnd.n4583 19.3944
R16753 gnd.n4583 gnd.n4580 19.3944
R16754 gnd.n4580 gnd.n4579 19.3944
R16755 gnd.n4579 gnd.n4576 19.3944
R16756 gnd.n4576 gnd.n4575 19.3944
R16757 gnd.n4575 gnd.n4572 19.3944
R16758 gnd.n4572 gnd.n4571 19.3944
R16759 gnd.n4571 gnd.n4568 19.3944
R16760 gnd.n4568 gnd.n4567 19.3944
R16761 gnd.n4567 gnd.n4564 19.3944
R16762 gnd.n4564 gnd.n4563 19.3944
R16763 gnd.n2065 gnd.n2064 19.3944
R16764 gnd.n5351 gnd.n2064 19.3944
R16765 gnd.n5351 gnd.n5350 19.3944
R16766 gnd.n5350 gnd.n5349 19.3944
R16767 gnd.n5349 gnd.n5346 19.3944
R16768 gnd.n5346 gnd.n5345 19.3944
R16769 gnd.n5345 gnd.n5342 19.3944
R16770 gnd.n5342 gnd.n5341 19.3944
R16771 gnd.n5341 gnd.n5338 19.3944
R16772 gnd.n5338 gnd.n5337 19.3944
R16773 gnd.n5337 gnd.n5334 19.3944
R16774 gnd.n5334 gnd.n5333 19.3944
R16775 gnd.n5333 gnd.n5330 19.3944
R16776 gnd.n5330 gnd.n5329 19.3944
R16777 gnd.n5329 gnd.n5326 19.3944
R16778 gnd.n4177 gnd.n2311 19.3944
R16779 gnd.n4189 gnd.n2311 19.3944
R16780 gnd.n4189 gnd.n2309 19.3944
R16781 gnd.n4193 gnd.n2309 19.3944
R16782 gnd.n4193 gnd.n2295 19.3944
R16783 gnd.n4205 gnd.n2295 19.3944
R16784 gnd.n4205 gnd.n2293 19.3944
R16785 gnd.n4209 gnd.n2293 19.3944
R16786 gnd.n4209 gnd.n2279 19.3944
R16787 gnd.n4221 gnd.n2279 19.3944
R16788 gnd.n4221 gnd.n2277 19.3944
R16789 gnd.n4225 gnd.n2277 19.3944
R16790 gnd.n4225 gnd.n2263 19.3944
R16791 gnd.n4237 gnd.n2263 19.3944
R16792 gnd.n4237 gnd.n2261 19.3944
R16793 gnd.n4241 gnd.n2261 19.3944
R16794 gnd.n4241 gnd.n2247 19.3944
R16795 gnd.n4253 gnd.n2247 19.3944
R16796 gnd.n4253 gnd.n2245 19.3944
R16797 gnd.n4257 gnd.n2245 19.3944
R16798 gnd.n4257 gnd.n2231 19.3944
R16799 gnd.n4269 gnd.n2231 19.3944
R16800 gnd.n4269 gnd.n2229 19.3944
R16801 gnd.n4274 gnd.n2229 19.3944
R16802 gnd.n4274 gnd.n2214 19.3944
R16803 gnd.n4286 gnd.n2214 19.3944
R16804 gnd.n4287 gnd.n4286 19.3944
R16805 gnd.n4290 gnd.n4289 19.3944
R16806 gnd.n4304 gnd.n4303 19.3944
R16807 gnd.n4307 gnd.n4306 19.3944
R16808 gnd.n4331 gnd.n4330 19.3944
R16809 gnd.n4333 gnd.n977 19.3944
R16810 gnd.n6337 gnd.n977 19.3944
R16811 gnd.n6337 gnd.n6336 19.3944
R16812 gnd.n6336 gnd.n6335 19.3944
R16813 gnd.n6335 gnd.n981 19.3944
R16814 gnd.n6325 gnd.n981 19.3944
R16815 gnd.n6325 gnd.n6324 19.3944
R16816 gnd.n6324 gnd.n6323 19.3944
R16817 gnd.n6323 gnd.n1003 19.3944
R16818 gnd.n6313 gnd.n1003 19.3944
R16819 gnd.n6313 gnd.n6312 19.3944
R16820 gnd.n6312 gnd.n6311 19.3944
R16821 gnd.n6311 gnd.n1024 19.3944
R16822 gnd.n6301 gnd.n1024 19.3944
R16823 gnd.n6301 gnd.n6300 19.3944
R16824 gnd.n6300 gnd.n6299 19.3944
R16825 gnd.n6299 gnd.n1045 19.3944
R16826 gnd.n6289 gnd.n1045 19.3944
R16827 gnd.n6289 gnd.n6288 19.3944
R16828 gnd.n6288 gnd.n6287 19.3944
R16829 gnd.n6287 gnd.n1066 19.3944
R16830 gnd.n6277 gnd.n1066 19.3944
R16831 gnd.n6277 gnd.n6276 19.3944
R16832 gnd.n6276 gnd.n6275 19.3944
R16833 gnd.n6275 gnd.n1087 19.3944
R16834 gnd.n6265 gnd.n1087 19.3944
R16835 gnd.n6265 gnd.n6264 19.3944
R16836 gnd.n6264 gnd.n6263 19.3944
R16837 gnd.n6514 gnd.n6513 19.3944
R16838 gnd.n6513 gnd.n800 19.3944
R16839 gnd.n6507 gnd.n800 19.3944
R16840 gnd.n6507 gnd.n6506 19.3944
R16841 gnd.n6506 gnd.n6505 19.3944
R16842 gnd.n6505 gnd.n808 19.3944
R16843 gnd.n6499 gnd.n808 19.3944
R16844 gnd.n6499 gnd.n6498 19.3944
R16845 gnd.n6498 gnd.n6497 19.3944
R16846 gnd.n6497 gnd.n816 19.3944
R16847 gnd.n6491 gnd.n816 19.3944
R16848 gnd.n6491 gnd.n6490 19.3944
R16849 gnd.n6490 gnd.n6489 19.3944
R16850 gnd.n6489 gnd.n824 19.3944
R16851 gnd.n6483 gnd.n824 19.3944
R16852 gnd.n6483 gnd.n6482 19.3944
R16853 gnd.n6482 gnd.n6481 19.3944
R16854 gnd.n6481 gnd.n832 19.3944
R16855 gnd.n6475 gnd.n832 19.3944
R16856 gnd.n6475 gnd.n6474 19.3944
R16857 gnd.n6474 gnd.n6473 19.3944
R16858 gnd.n6473 gnd.n840 19.3944
R16859 gnd.n6467 gnd.n840 19.3944
R16860 gnd.n6467 gnd.n6466 19.3944
R16861 gnd.n6466 gnd.n6465 19.3944
R16862 gnd.n6465 gnd.n848 19.3944
R16863 gnd.n6459 gnd.n848 19.3944
R16864 gnd.n6459 gnd.n6458 19.3944
R16865 gnd.n6458 gnd.n6457 19.3944
R16866 gnd.n6457 gnd.n856 19.3944
R16867 gnd.n6451 gnd.n856 19.3944
R16868 gnd.n6451 gnd.n6450 19.3944
R16869 gnd.n6450 gnd.n6449 19.3944
R16870 gnd.n6449 gnd.n864 19.3944
R16871 gnd.n6443 gnd.n864 19.3944
R16872 gnd.n6443 gnd.n6442 19.3944
R16873 gnd.n6442 gnd.n6441 19.3944
R16874 gnd.n6441 gnd.n872 19.3944
R16875 gnd.n6435 gnd.n872 19.3944
R16876 gnd.n6435 gnd.n6434 19.3944
R16877 gnd.n6434 gnd.n6433 19.3944
R16878 gnd.n6433 gnd.n880 19.3944
R16879 gnd.n6427 gnd.n880 19.3944
R16880 gnd.n6427 gnd.n6426 19.3944
R16881 gnd.n6426 gnd.n6425 19.3944
R16882 gnd.n6425 gnd.n888 19.3944
R16883 gnd.n6419 gnd.n888 19.3944
R16884 gnd.n6419 gnd.n6418 19.3944
R16885 gnd.n6418 gnd.n6417 19.3944
R16886 gnd.n6417 gnd.n896 19.3944
R16887 gnd.n6411 gnd.n896 19.3944
R16888 gnd.n6411 gnd.n6410 19.3944
R16889 gnd.n6410 gnd.n6409 19.3944
R16890 gnd.n6409 gnd.n904 19.3944
R16891 gnd.n6403 gnd.n904 19.3944
R16892 gnd.n6403 gnd.n6402 19.3944
R16893 gnd.n6402 gnd.n6401 19.3944
R16894 gnd.n6401 gnd.n912 19.3944
R16895 gnd.n6395 gnd.n912 19.3944
R16896 gnd.n6395 gnd.n6394 19.3944
R16897 gnd.n6394 gnd.n6393 19.3944
R16898 gnd.n6393 gnd.n920 19.3944
R16899 gnd.n6387 gnd.n920 19.3944
R16900 gnd.n6387 gnd.n6386 19.3944
R16901 gnd.n6386 gnd.n6385 19.3944
R16902 gnd.n6385 gnd.n928 19.3944
R16903 gnd.n6379 gnd.n928 19.3944
R16904 gnd.n6379 gnd.n6378 19.3944
R16905 gnd.n6378 gnd.n6377 19.3944
R16906 gnd.n6377 gnd.n936 19.3944
R16907 gnd.n6371 gnd.n936 19.3944
R16908 gnd.n6371 gnd.n6370 19.3944
R16909 gnd.n6370 gnd.n6369 19.3944
R16910 gnd.n6369 gnd.n944 19.3944
R16911 gnd.n6363 gnd.n944 19.3944
R16912 gnd.n6363 gnd.n6362 19.3944
R16913 gnd.n6362 gnd.n6361 19.3944
R16914 gnd.n6361 gnd.n952 19.3944
R16915 gnd.n6355 gnd.n952 19.3944
R16916 gnd.n6355 gnd.n6354 19.3944
R16917 gnd.n6354 gnd.n6353 19.3944
R16918 gnd.n6353 gnd.n960 19.3944
R16919 gnd.n6347 gnd.n960 19.3944
R16920 gnd.n6347 gnd.n6346 19.3944
R16921 gnd.n6254 gnd.n6253 19.3944
R16922 gnd.n6253 gnd.n6252 19.3944
R16923 gnd.n6252 gnd.n1121 19.3944
R16924 gnd.n6248 gnd.n1121 19.3944
R16925 gnd.n6248 gnd.n6247 19.3944
R16926 gnd.n6247 gnd.n6246 19.3944
R16927 gnd.n6246 gnd.n1126 19.3944
R16928 gnd.n6242 gnd.n1126 19.3944
R16929 gnd.n6242 gnd.n6241 19.3944
R16930 gnd.n6241 gnd.n6240 19.3944
R16931 gnd.n6240 gnd.n1131 19.3944
R16932 gnd.n6236 gnd.n1131 19.3944
R16933 gnd.n6236 gnd.n6235 19.3944
R16934 gnd.n6235 gnd.n6234 19.3944
R16935 gnd.n6234 gnd.n1136 19.3944
R16936 gnd.n6230 gnd.n1136 19.3944
R16937 gnd.n6230 gnd.n6229 19.3944
R16938 gnd.n6229 gnd.n6228 19.3944
R16939 gnd.n6228 gnd.n1141 19.3944
R16940 gnd.n6224 gnd.n1141 19.3944
R16941 gnd.n6224 gnd.n6223 19.3944
R16942 gnd.n6223 gnd.n6222 19.3944
R16943 gnd.n6222 gnd.n1146 19.3944
R16944 gnd.n6218 gnd.n1146 19.3944
R16945 gnd.n6218 gnd.n6217 19.3944
R16946 gnd.n6217 gnd.n6216 19.3944
R16947 gnd.n6216 gnd.n1151 19.3944
R16948 gnd.n6212 gnd.n1151 19.3944
R16949 gnd.n6212 gnd.n6211 19.3944
R16950 gnd.n6211 gnd.n6210 19.3944
R16951 gnd.n6210 gnd.n1156 19.3944
R16952 gnd.n6206 gnd.n1156 19.3944
R16953 gnd.n6206 gnd.n6205 19.3944
R16954 gnd.n6205 gnd.n6204 19.3944
R16955 gnd.n6204 gnd.n1161 19.3944
R16956 gnd.n6200 gnd.n1161 19.3944
R16957 gnd.n6200 gnd.n6199 19.3944
R16958 gnd.n6199 gnd.n6198 19.3944
R16959 gnd.n6198 gnd.n1166 19.3944
R16960 gnd.n6194 gnd.n1166 19.3944
R16961 gnd.n6194 gnd.n6193 19.3944
R16962 gnd.n6193 gnd.n6192 19.3944
R16963 gnd.n6192 gnd.n1171 19.3944
R16964 gnd.n6188 gnd.n1171 19.3944
R16965 gnd.n6188 gnd.n6187 19.3944
R16966 gnd.n6187 gnd.n6186 19.3944
R16967 gnd.n6186 gnd.n1176 19.3944
R16968 gnd.n6182 gnd.n1176 19.3944
R16969 gnd.n6182 gnd.n6181 19.3944
R16970 gnd.n6181 gnd.n6180 19.3944
R16971 gnd.n6180 gnd.n1181 19.3944
R16972 gnd.n6176 gnd.n1181 19.3944
R16973 gnd.n6176 gnd.n6175 19.3944
R16974 gnd.n6175 gnd.n6174 19.3944
R16975 gnd.n6174 gnd.n1186 19.3944
R16976 gnd.n6170 gnd.n1186 19.3944
R16977 gnd.n6170 gnd.n6169 19.3944
R16978 gnd.n6169 gnd.n6168 19.3944
R16979 gnd.n6168 gnd.n1191 19.3944
R16980 gnd.n6164 gnd.n1191 19.3944
R16981 gnd.n6164 gnd.n6163 19.3944
R16982 gnd.n6163 gnd.n6162 19.3944
R16983 gnd.n6162 gnd.n1196 19.3944
R16984 gnd.n6158 gnd.n1196 19.3944
R16985 gnd.n6158 gnd.n6157 19.3944
R16986 gnd.n6157 gnd.n6156 19.3944
R16987 gnd.n6156 gnd.n1201 19.3944
R16988 gnd.n6152 gnd.n1201 19.3944
R16989 gnd.n6152 gnd.n6151 19.3944
R16990 gnd.n6151 gnd.n6150 19.3944
R16991 gnd.n6150 gnd.n1206 19.3944
R16992 gnd.n6146 gnd.n1206 19.3944
R16993 gnd.n6146 gnd.n6145 19.3944
R16994 gnd.n6145 gnd.n6144 19.3944
R16995 gnd.n6144 gnd.n1211 19.3944
R16996 gnd.n6140 gnd.n1211 19.3944
R16997 gnd.n6140 gnd.n6139 19.3944
R16998 gnd.n6139 gnd.n6138 19.3944
R16999 gnd.n6138 gnd.n1216 19.3944
R17000 gnd.n6134 gnd.n1216 19.3944
R17001 gnd.n6134 gnd.n6133 19.3944
R17002 gnd.n6133 gnd.n6132 19.3944
R17003 gnd.n6132 gnd.n1221 19.3944
R17004 gnd.n6128 gnd.n1221 19.3944
R17005 gnd.n6128 gnd.n6127 19.3944
R17006 gnd.n6127 gnd.n6126 19.3944
R17007 gnd.n6126 gnd.n1226 19.3944
R17008 gnd.n6122 gnd.n1226 19.3944
R17009 gnd.n6122 gnd.n6121 19.3944
R17010 gnd.n6121 gnd.n6120 19.3944
R17011 gnd.n6120 gnd.n1231 19.3944
R17012 gnd.n6116 gnd.n1231 19.3944
R17013 gnd.n6116 gnd.n6115 19.3944
R17014 gnd.n6115 gnd.n6114 19.3944
R17015 gnd.n6114 gnd.n1236 19.3944
R17016 gnd.n6110 gnd.n1236 19.3944
R17017 gnd.n6110 gnd.n6109 19.3944
R17018 gnd.n6109 gnd.n6108 19.3944
R17019 gnd.n6108 gnd.n1241 19.3944
R17020 gnd.n6104 gnd.n1241 19.3944
R17021 gnd.n6104 gnd.n6103 19.3944
R17022 gnd.n5826 gnd.n1614 19.3944
R17023 gnd.n5822 gnd.n1614 19.3944
R17024 gnd.n5822 gnd.n5821 19.3944
R17025 gnd.n1530 gnd.n1514 19.3944
R17026 gnd.n1530 gnd.n1512 19.3944
R17027 gnd.n1536 gnd.n1512 19.3944
R17028 gnd.n1536 gnd.n1507 19.3944
R17029 gnd.n1549 gnd.n1507 19.3944
R17030 gnd.n1549 gnd.n1505 19.3944
R17031 gnd.n1555 gnd.n1505 19.3944
R17032 gnd.n1555 gnd.n1500 19.3944
R17033 gnd.n1568 gnd.n1500 19.3944
R17034 gnd.n1568 gnd.n1498 19.3944
R17035 gnd.n1574 gnd.n1498 19.3944
R17036 gnd.n1574 gnd.n1494 19.3944
R17037 gnd.n1584 gnd.n1494 19.3944
R17038 gnd.n1584 gnd.n1492 19.3944
R17039 gnd.n1590 gnd.n1492 19.3944
R17040 gnd.n1590 gnd.n1482 19.3944
R17041 gnd.n1598 gnd.n1482 19.3944
R17042 gnd.n1598 gnd.n1480 19.3944
R17043 gnd.n5837 gnd.n1480 19.3944
R17044 gnd.n5837 gnd.n5836 19.3944
R17045 gnd.n5836 gnd.n5835 19.3944
R17046 gnd.n5835 gnd.n1606 19.3944
R17047 gnd.n5831 gnd.n1606 19.3944
R17048 gnd.n5831 gnd.n5830 19.3944
R17049 gnd.n6349 gnd.n962 19.1977
R17050 gnd.t281 gnd.n1859 19.1199
R17051 gnd.t278 gnd.n1706 19.1199
R17052 gnd.n5255 gnd.n5254 18.8883
R17053 gnd.n4949 gnd.n4948 18.8883
R17054 gnd.n3179 gnd.t222 18.8012
R17055 gnd.n3164 gnd.t64 18.8012
R17056 gnd.n3023 gnd.n3022 18.4825
R17057 gnd.n5557 gnd.n1833 18.4825
R17058 gnd.n4857 gnd.n1742 18.4825
R17059 gnd.n6061 gnd.n6060 18.4247
R17060 gnd.n5326 gnd.n5325 18.4247
R17061 gnd.n7479 gnd.n124 18.2308
R17062 gnd.n1594 gnd.n1593 18.2308
R17063 gnd.n5364 gnd.n2018 18.2308
R17064 gnd.n3856 gnd.n3800 18.2308
R17065 gnd.t223 gnd.n2703 18.1639
R17066 gnd.n2731 gnd.t220 17.5266
R17067 gnd.t124 gnd.n1812 17.5266
R17068 gnd.n5148 gnd.t193 17.5266
R17069 gnd.n4743 gnd.t304 17.2079
R17070 gnd.n3130 gnd.t215 16.8893
R17071 gnd.n5493 gnd.t130 16.8893
R17072 gnd.t191 gnd.n1839 16.8893
R17073 gnd.n5115 gnd.t117 16.8893
R17074 gnd.n1686 gnd.t77 16.8893
R17075 gnd.n5101 gnd.t301 16.5706
R17076 gnd.n2958 gnd.t310 16.2519
R17077 gnd.n2658 gnd.t214 16.2519
R17078 gnd.n5321 gnd.n4637 16.2519
R17079 gnd.n5709 gnd.n1700 16.2519
R17080 gnd.n4667 gnd.n4666 16.0975
R17081 gnd.n4905 gnd.n4904 16.0975
R17082 gnd.n5257 gnd.n5256 16.0975
R17083 gnd.n5007 gnd.n5006 16.0975
R17084 gnd.n5191 gnd.t129 15.9333
R17085 gnd.n5177 gnd.n1782 15.9333
R17086 gnd.n5613 gnd.n1782 15.9333
R17087 gnd.t23 gnd.n1768 15.9333
R17088 gnd.n5109 gnd.n5108 15.9333
R17089 gnd.n3645 gnd.n3643 15.6674
R17090 gnd.n3613 gnd.n3611 15.6674
R17091 gnd.n3581 gnd.n3579 15.6674
R17092 gnd.n3550 gnd.n3548 15.6674
R17093 gnd.n3518 gnd.n3516 15.6674
R17094 gnd.n3486 gnd.n3484 15.6674
R17095 gnd.n3454 gnd.n3452 15.6674
R17096 gnd.n3423 gnd.n3421 15.6674
R17097 gnd.n2949 gnd.t310 15.6146
R17098 gnd.t288 gnd.n2400 15.6146
R17099 gnd.t271 gnd.n2401 15.6146
R17100 gnd.n4637 gnd.t339 15.296
R17101 gnd.n5193 gnd.t21 15.296
R17102 gnd.t1 gnd.n1770 15.296
R17103 gnd.n4928 gnd.n4927 15.0827
R17104 gnd.n4649 gnd.n4644 15.0481
R17105 gnd.n4938 gnd.n4937 15.0481
R17106 gnd.n3317 gnd.t209 14.9773
R17107 gnd.n1894 gnd.t130 14.9773
R17108 gnd.n5733 gnd.t77 14.9773
R17109 gnd.n5533 gnd.t304 14.6587
R17110 gnd.n5223 gnd.n5222 14.6587
R17111 gnd.n5669 gnd.n1734 14.6587
R17112 gnd.n5101 gnd.n4876 14.6587
R17113 gnd.n4878 gnd.t318 14.6587
R17114 gnd.t60 gnd.n2443 14.34
R17115 gnd.n3395 gnd.t218 14.34
R17116 gnd.n3105 gnd.t66 13.7027
R17117 gnd.n2815 gnd.n2814 13.5763
R17118 gnd.n3759 gnd.n2356 13.5763
R17119 gnd.n6023 gnd.n1332 13.5763
R17120 gnd.n7531 gnd.n7530 13.5763
R17121 gnd.n4104 gnd.n4019 13.5763
R17122 gnd.n4563 gnd.n4560 13.5763
R17123 gnd.n3023 gnd.n2761 13.384
R17124 gnd.n5525 gnd.n1860 13.384
R17125 gnd.n4763 gnd.n1833 13.384
R17126 gnd.n5192 gnd.n5191 13.384
R17127 gnd.n5605 gnd.t174 13.384
R17128 gnd.t116 gnd.n4817 13.384
R17129 gnd.n5629 gnd.n1768 13.384
R17130 gnd.n5661 gnd.n1742 13.384
R17131 gnd.n5094 gnd.n5093 13.384
R17132 gnd.n4660 gnd.n4641 13.1884
R17133 gnd.n4655 gnd.n4654 13.1884
R17134 gnd.n4654 gnd.n4653 13.1884
R17135 gnd.n4931 gnd.n4926 13.1884
R17136 gnd.n4932 gnd.n4931 13.1884
R17137 gnd.n4656 gnd.n4643 13.146
R17138 gnd.n4652 gnd.n4643 13.146
R17139 gnd.n4930 gnd.n4929 13.146
R17140 gnd.n4930 gnd.n4925 13.146
R17141 gnd.t111 gnd.n973 13.0654
R17142 gnd.t172 gnd.n356 13.0654
R17143 gnd.n3646 gnd.n3642 12.8005
R17144 gnd.n3614 gnd.n3610 12.8005
R17145 gnd.n3582 gnd.n3578 12.8005
R17146 gnd.n3551 gnd.n3547 12.8005
R17147 gnd.n3519 gnd.n3515 12.8005
R17148 gnd.n3487 gnd.n3483 12.8005
R17149 gnd.n3455 gnd.n3451 12.8005
R17150 gnd.n3424 gnd.n3420 12.8005
R17151 gnd.n5321 gnd.t24 12.7467
R17152 gnd.n2291 gnd.t7 12.4281
R17153 gnd.t137 gnd.n1018 12.4281
R17154 gnd.n4431 gnd.t183 12.4281
R17155 gnd.n5437 gnd.t350 12.4281
R17156 gnd.n1640 gnd.t133 12.4281
R17157 gnd.n5909 gnd.t48 12.4281
R17158 gnd.t15 gnd.n399 12.4281
R17159 gnd.t148 gnd.n229 12.4281
R17160 gnd.n2814 gnd.n2809 12.4126
R17161 gnd.n3762 gnd.n3759 12.4126
R17162 gnd.n6019 gnd.n1332 12.4126
R17163 gnd.n7530 gnd.n200 12.4126
R17164 gnd.n4100 gnd.n4019 12.4126
R17165 gnd.n4560 gnd.n2104 12.4126
R17166 gnd.n5318 gnd.n5255 12.1761
R17167 gnd.n4950 gnd.n4949 12.1761
R17168 gnd.n5354 gnd.n2027 12.1094
R17169 gnd.n5517 gnd.n1868 12.1094
R17170 gnd.n5230 gnd.t244 12.1094
R17171 gnd.n4776 gnd.n1827 12.1094
R17172 gnd.n4795 gnd.n1803 12.1094
R17173 gnd.n5637 gnd.n1761 12.1094
R17174 gnd.n5653 gnd.n1748 12.1094
R17175 gnd.n1707 gnd.t333 12.1094
R17176 gnd.n6092 gnd.n1285 12.1094
R17177 gnd.n3650 gnd.n3649 12.0247
R17178 gnd.n3618 gnd.n3617 12.0247
R17179 gnd.n3586 gnd.n3585 12.0247
R17180 gnd.n3555 gnd.n3554 12.0247
R17181 gnd.n3523 gnd.n3522 12.0247
R17182 gnd.n3491 gnd.n3490 12.0247
R17183 gnd.n3459 gnd.n3458 12.0247
R17184 gnd.n3428 gnd.n3427 12.0247
R17185 gnd.n2259 gnd.t27 11.7908
R17186 gnd.n4378 gnd.t137 11.7908
R17187 gnd.t183 gnd.n1060 11.7908
R17188 gnd.t48 gnd.n5907 11.7908
R17189 gnd.n5936 gnd.t15 11.7908
R17190 gnd.t35 gnd.n260 11.7908
R17191 gnd.n4750 gnd.t95 11.4721
R17192 gnd.n5214 gnd.t190 11.4721
R17193 gnd.t26 gnd.n1740 11.4721
R17194 gnd.n5677 gnd.t22 11.4721
R17195 gnd.n3653 gnd.n3640 11.249
R17196 gnd.n3621 gnd.n3608 11.249
R17197 gnd.n3589 gnd.n3576 11.249
R17198 gnd.n3558 gnd.n3545 11.249
R17199 gnd.n3526 gnd.n3513 11.249
R17200 gnd.n3494 gnd.n3481 11.249
R17201 gnd.n3462 gnd.n3449 11.249
R17202 gnd.n3431 gnd.n3418 11.249
R17203 gnd.n3093 gnd.t66 11.1535
R17204 gnd.n2227 gnd.t98 11.1535
R17205 gnd.n4344 gnd.t111 11.1535
R17206 gnd.n7206 gnd.t172 11.1535
R17207 gnd.t9 gnd.n290 11.1535
R17208 gnd.n1819 gnd.n1810 10.8348
R17209 gnd.n5645 gnd.n1754 10.8348
R17210 gnd.n5021 gnd.n4906 10.6151
R17211 gnd.n5027 gnd.n4906 10.6151
R17212 gnd.n5030 gnd.n5029 10.6151
R17213 gnd.n5030 gnd.n4902 10.6151
R17214 gnd.n5036 gnd.n4902 10.6151
R17215 gnd.n5037 gnd.n5036 10.6151
R17216 gnd.n5038 gnd.n5037 10.6151
R17217 gnd.n5038 gnd.n4900 10.6151
R17218 gnd.n5044 gnd.n4900 10.6151
R17219 gnd.n5045 gnd.n5044 10.6151
R17220 gnd.n5046 gnd.n5045 10.6151
R17221 gnd.n5046 gnd.n4898 10.6151
R17222 gnd.n5052 gnd.n4898 10.6151
R17223 gnd.n5053 gnd.n5052 10.6151
R17224 gnd.n5054 gnd.n5053 10.6151
R17225 gnd.n5054 gnd.n4896 10.6151
R17226 gnd.n5060 gnd.n4896 10.6151
R17227 gnd.n5061 gnd.n5060 10.6151
R17228 gnd.n5062 gnd.n5061 10.6151
R17229 gnd.n5062 gnd.n4894 10.6151
R17230 gnd.n5068 gnd.n4894 10.6151
R17231 gnd.n5069 gnd.n5068 10.6151
R17232 gnd.n5070 gnd.n5069 10.6151
R17233 gnd.n5070 gnd.n4892 10.6151
R17234 gnd.n5076 gnd.n4892 10.6151
R17235 gnd.n5077 gnd.n5076 10.6151
R17236 gnd.n5078 gnd.n5077 10.6151
R17237 gnd.n5078 gnd.n4890 10.6151
R17238 gnd.n5083 gnd.n4890 10.6151
R17239 gnd.n5084 gnd.n5083 10.6151
R17240 gnd.n4733 gnd.n4732 10.6151
R17241 gnd.n5248 gnd.n4733 10.6151
R17242 gnd.n5248 gnd.n5247 10.6151
R17243 gnd.n5247 gnd.n5246 10.6151
R17244 gnd.n5246 gnd.n4734 10.6151
R17245 gnd.n4746 gnd.n4734 10.6151
R17246 gnd.n4747 gnd.n4746 10.6151
R17247 gnd.n5234 gnd.n4747 10.6151
R17248 gnd.n5234 gnd.n5233 10.6151
R17249 gnd.n5233 gnd.n5232 10.6151
R17250 gnd.n5232 gnd.n4748 10.6151
R17251 gnd.n4767 gnd.n4748 10.6151
R17252 gnd.n4768 gnd.n4767 10.6151
R17253 gnd.n4769 gnd.n4768 10.6151
R17254 gnd.n4770 gnd.n4769 10.6151
R17255 gnd.n4772 gnd.n4770 10.6151
R17256 gnd.n4773 gnd.n4772 10.6151
R17257 gnd.n5211 gnd.n4773 10.6151
R17258 gnd.n5211 gnd.n5210 10.6151
R17259 gnd.n5210 gnd.n5209 10.6151
R17260 gnd.n5209 gnd.n4774 10.6151
R17261 gnd.n4789 gnd.n4774 10.6151
R17262 gnd.n4792 gnd.n4789 10.6151
R17263 gnd.n4793 gnd.n4792 10.6151
R17264 gnd.n4794 gnd.n4793 10.6151
R17265 gnd.n4794 gnd.n4787 10.6151
R17266 gnd.n4800 gnd.n4787 10.6151
R17267 gnd.n4801 gnd.n4800 10.6151
R17268 gnd.n5189 gnd.n4801 10.6151
R17269 gnd.n5189 gnd.n5188 10.6151
R17270 gnd.n5188 gnd.n5187 10.6151
R17271 gnd.n5187 gnd.n4802 10.6151
R17272 gnd.n4814 gnd.n4802 10.6151
R17273 gnd.n5175 gnd.n4814 10.6151
R17274 gnd.n5175 gnd.n5174 10.6151
R17275 gnd.n5174 gnd.n5173 10.6151
R17276 gnd.n5173 gnd.n4815 10.6151
R17277 gnd.n4827 gnd.n4815 10.6151
R17278 gnd.n4828 gnd.n4827 10.6151
R17279 gnd.n5160 gnd.n4828 10.6151
R17280 gnd.n5160 gnd.n5159 10.6151
R17281 gnd.n5159 gnd.n5158 10.6151
R17282 gnd.n5158 gnd.n4829 10.6151
R17283 gnd.n4840 gnd.n4829 10.6151
R17284 gnd.n4841 gnd.n4840 10.6151
R17285 gnd.n5145 gnd.n4841 10.6151
R17286 gnd.n5145 gnd.n5144 10.6151
R17287 gnd.n5144 gnd.n5143 10.6151
R17288 gnd.n5143 gnd.n4842 10.6151
R17289 gnd.n5133 gnd.n4842 10.6151
R17290 gnd.n5133 gnd.n5132 10.6151
R17291 gnd.n5132 gnd.n5131 10.6151
R17292 gnd.n5131 gnd.n4851 10.6151
R17293 gnd.n4860 gnd.n4851 10.6151
R17294 gnd.n5120 gnd.n4860 10.6151
R17295 gnd.n5120 gnd.n5119 10.6151
R17296 gnd.n5119 gnd.n5118 10.6151
R17297 gnd.n5118 gnd.n4861 10.6151
R17298 gnd.n4872 gnd.n4861 10.6151
R17299 gnd.n4873 gnd.n4872 10.6151
R17300 gnd.n5105 gnd.n4873 10.6151
R17301 gnd.n5105 gnd.n5104 10.6151
R17302 gnd.n5104 gnd.n5103 10.6151
R17303 gnd.n5103 gnd.n4874 10.6151
R17304 gnd.n4886 gnd.n4874 10.6151
R17305 gnd.n4887 gnd.n4886 10.6151
R17306 gnd.n5090 gnd.n4887 10.6151
R17307 gnd.n5090 gnd.n5089 10.6151
R17308 gnd.n5089 gnd.n5088 10.6151
R17309 gnd.n5088 gnd.n4888 10.6151
R17310 gnd.n4668 gnd.n4602 10.6151
R17311 gnd.n4671 gnd.n4668 10.6151
R17312 gnd.n4676 gnd.n4673 10.6151
R17313 gnd.n4677 gnd.n4676 10.6151
R17314 gnd.n4680 gnd.n4677 10.6151
R17315 gnd.n4681 gnd.n4680 10.6151
R17316 gnd.n4684 gnd.n4681 10.6151
R17317 gnd.n4685 gnd.n4684 10.6151
R17318 gnd.n4688 gnd.n4685 10.6151
R17319 gnd.n4689 gnd.n4688 10.6151
R17320 gnd.n4692 gnd.n4689 10.6151
R17321 gnd.n4693 gnd.n4692 10.6151
R17322 gnd.n4696 gnd.n4693 10.6151
R17323 gnd.n4697 gnd.n4696 10.6151
R17324 gnd.n4700 gnd.n4697 10.6151
R17325 gnd.n4701 gnd.n4700 10.6151
R17326 gnd.n4704 gnd.n4701 10.6151
R17327 gnd.n4705 gnd.n4704 10.6151
R17328 gnd.n4708 gnd.n4705 10.6151
R17329 gnd.n4709 gnd.n4708 10.6151
R17330 gnd.n4712 gnd.n4709 10.6151
R17331 gnd.n4713 gnd.n4712 10.6151
R17332 gnd.n4716 gnd.n4713 10.6151
R17333 gnd.n4717 gnd.n4716 10.6151
R17334 gnd.n4720 gnd.n4717 10.6151
R17335 gnd.n4721 gnd.n4720 10.6151
R17336 gnd.n4724 gnd.n4721 10.6151
R17337 gnd.n4725 gnd.n4724 10.6151
R17338 gnd.n4728 gnd.n4725 10.6151
R17339 gnd.n4729 gnd.n4728 10.6151
R17340 gnd.n5318 gnd.n5317 10.6151
R17341 gnd.n5317 gnd.n5316 10.6151
R17342 gnd.n5316 gnd.n5315 10.6151
R17343 gnd.n5315 gnd.n5313 10.6151
R17344 gnd.n5313 gnd.n5310 10.6151
R17345 gnd.n5310 gnd.n5309 10.6151
R17346 gnd.n5309 gnd.n5306 10.6151
R17347 gnd.n5306 gnd.n5305 10.6151
R17348 gnd.n5305 gnd.n5302 10.6151
R17349 gnd.n5302 gnd.n5301 10.6151
R17350 gnd.n5301 gnd.n5298 10.6151
R17351 gnd.n5298 gnd.n5297 10.6151
R17352 gnd.n5297 gnd.n5294 10.6151
R17353 gnd.n5294 gnd.n5293 10.6151
R17354 gnd.n5293 gnd.n5290 10.6151
R17355 gnd.n5290 gnd.n5289 10.6151
R17356 gnd.n5289 gnd.n5286 10.6151
R17357 gnd.n5286 gnd.n5285 10.6151
R17358 gnd.n5285 gnd.n5282 10.6151
R17359 gnd.n5282 gnd.n5281 10.6151
R17360 gnd.n5281 gnd.n5278 10.6151
R17361 gnd.n5278 gnd.n5277 10.6151
R17362 gnd.n5277 gnd.n5274 10.6151
R17363 gnd.n5274 gnd.n5273 10.6151
R17364 gnd.n5273 gnd.n5270 10.6151
R17365 gnd.n5270 gnd.n5269 10.6151
R17366 gnd.n5269 gnd.n5266 10.6151
R17367 gnd.n5266 gnd.n5265 10.6151
R17368 gnd.n5262 gnd.n5261 10.6151
R17369 gnd.n5261 gnd.n4603 10.6151
R17370 gnd.n4950 gnd.n4922 10.6151
R17371 gnd.n4956 gnd.n4922 10.6151
R17372 gnd.n4957 gnd.n4956 10.6151
R17373 gnd.n4958 gnd.n4957 10.6151
R17374 gnd.n4958 gnd.n4920 10.6151
R17375 gnd.n4964 gnd.n4920 10.6151
R17376 gnd.n4965 gnd.n4964 10.6151
R17377 gnd.n4966 gnd.n4965 10.6151
R17378 gnd.n4966 gnd.n4918 10.6151
R17379 gnd.n4972 gnd.n4918 10.6151
R17380 gnd.n4973 gnd.n4972 10.6151
R17381 gnd.n4974 gnd.n4973 10.6151
R17382 gnd.n4974 gnd.n4916 10.6151
R17383 gnd.n4980 gnd.n4916 10.6151
R17384 gnd.n4981 gnd.n4980 10.6151
R17385 gnd.n4982 gnd.n4981 10.6151
R17386 gnd.n4982 gnd.n4914 10.6151
R17387 gnd.n4988 gnd.n4914 10.6151
R17388 gnd.n4989 gnd.n4988 10.6151
R17389 gnd.n4990 gnd.n4989 10.6151
R17390 gnd.n4990 gnd.n4912 10.6151
R17391 gnd.n4996 gnd.n4912 10.6151
R17392 gnd.n4997 gnd.n4996 10.6151
R17393 gnd.n4998 gnd.n4997 10.6151
R17394 gnd.n4998 gnd.n4910 10.6151
R17395 gnd.n5004 gnd.n4910 10.6151
R17396 gnd.n5005 gnd.n5004 10.6151
R17397 gnd.n5009 gnd.n5005 10.6151
R17398 gnd.n5014 gnd.n4908 10.6151
R17399 gnd.n5015 gnd.n5014 10.6151
R17400 gnd.n5254 gnd.n5253 10.6151
R17401 gnd.n5253 gnd.n4661 10.6151
R17402 gnd.n4739 gnd.n4661 10.6151
R17403 gnd.n4740 gnd.n4739 10.6151
R17404 gnd.n5241 gnd.n4740 10.6151
R17405 gnd.n5241 gnd.n5240 10.6151
R17406 gnd.n5240 gnd.n5239 10.6151
R17407 gnd.n5239 gnd.n4741 10.6151
R17408 gnd.n4753 gnd.n4741 10.6151
R17409 gnd.n5228 gnd.n4753 10.6151
R17410 gnd.n5228 gnd.n5227 10.6151
R17411 gnd.n5227 gnd.n5226 10.6151
R17412 gnd.n5226 gnd.n4754 10.6151
R17413 gnd.n4760 gnd.n4754 10.6151
R17414 gnd.n5218 gnd.n4760 10.6151
R17415 gnd.n5218 gnd.n5217 10.6151
R17416 gnd.n5217 gnd.n5216 10.6151
R17417 gnd.n5216 gnd.n4761 10.6151
R17418 gnd.n4779 gnd.n4761 10.6151
R17419 gnd.n5205 gnd.n4779 10.6151
R17420 gnd.n5205 gnd.n5204 10.6151
R17421 gnd.n5204 gnd.n5203 10.6151
R17422 gnd.n5203 gnd.n4780 10.6151
R17423 gnd.n5199 gnd.n4780 10.6151
R17424 gnd.n5199 gnd.n5198 10.6151
R17425 gnd.n5198 gnd.n5197 10.6151
R17426 gnd.n5197 gnd.n4782 10.6151
R17427 gnd.n4784 gnd.n4782 10.6151
R17428 gnd.n4808 gnd.n4784 10.6151
R17429 gnd.n4809 gnd.n4808 10.6151
R17430 gnd.n5183 gnd.n4809 10.6151
R17431 gnd.n5183 gnd.n5182 10.6151
R17432 gnd.n5182 gnd.n5181 10.6151
R17433 gnd.n5181 gnd.n4810 10.6151
R17434 gnd.n4821 gnd.n4810 10.6151
R17435 gnd.n4822 gnd.n4821 10.6151
R17436 gnd.n5168 gnd.n4822 10.6151
R17437 gnd.n5168 gnd.n5167 10.6151
R17438 gnd.n5167 gnd.n5166 10.6151
R17439 gnd.n5166 gnd.n4823 10.6151
R17440 gnd.n4834 gnd.n4823 10.6151
R17441 gnd.n4835 gnd.n4834 10.6151
R17442 gnd.n5153 gnd.n4835 10.6151
R17443 gnd.n5153 gnd.n5152 10.6151
R17444 gnd.n5152 gnd.n5151 10.6151
R17445 gnd.n5151 gnd.n4836 10.6151
R17446 gnd.n4846 gnd.n4836 10.6151
R17447 gnd.n5139 gnd.n4846 10.6151
R17448 gnd.n5139 gnd.n5138 10.6151
R17449 gnd.n5138 gnd.n5137 10.6151
R17450 gnd.n5137 gnd.n4847 10.6151
R17451 gnd.n5127 gnd.n4847 10.6151
R17452 gnd.n5127 gnd.n5126 10.6151
R17453 gnd.n5126 gnd.n5125 10.6151
R17454 gnd.n5125 gnd.n4855 10.6151
R17455 gnd.n4866 gnd.n4855 10.6151
R17456 gnd.n4867 gnd.n4866 10.6151
R17457 gnd.n5113 gnd.n4867 10.6151
R17458 gnd.n5113 gnd.n5112 10.6151
R17459 gnd.n5112 gnd.n5111 10.6151
R17460 gnd.n5111 gnd.n4868 10.6151
R17461 gnd.n4880 gnd.n4868 10.6151
R17462 gnd.n5099 gnd.n4880 10.6151
R17463 gnd.n5099 gnd.n5098 10.6151
R17464 gnd.n5098 gnd.n5097 10.6151
R17465 gnd.n5097 gnd.n4881 10.6151
R17466 gnd.n4943 gnd.n4881 10.6151
R17467 gnd.n4944 gnd.n4943 10.6151
R17468 gnd.n4947 gnd.n4944 10.6151
R17469 gnd.n4948 gnd.n4947 10.6151
R17470 gnd.n3012 gnd.t62 10.5161
R17471 gnd.n2445 gnd.t60 10.5161
R17472 gnd.n3378 gnd.t218 10.5161
R17473 gnd.t86 gnd.n2194 10.5161
R17474 gnd.n2196 gnd.t160 10.5161
R17475 gnd.n7251 gnd.t101 10.5161
R17476 gnd.n7257 gnd.t195 10.5161
R17477 gnd.n3654 gnd.n3638 10.4732
R17478 gnd.n3622 gnd.n3606 10.4732
R17479 gnd.n3590 gnd.n3574 10.4732
R17480 gnd.n3559 gnd.n3543 10.4732
R17481 gnd.n3527 gnd.n3511 10.4732
R17482 gnd.n3495 gnd.n3479 10.4732
R17483 gnd.n3463 gnd.n3447 10.4732
R17484 gnd.n3432 gnd.n3416 10.4732
R17485 gnd.t190 gnd.n5213 10.1975
R17486 gnd.n5129 gnd.t26 10.1975
R17487 gnd.t209 gnd.n2462 9.87883
R17488 gnd.t169 gnd.n2224 9.87883
R17489 gnd.n293 gnd.t11 9.87883
R17490 gnd.n7656 gnd.n78 9.81789
R17491 gnd.n3658 gnd.n3657 9.69747
R17492 gnd.n3626 gnd.n3625 9.69747
R17493 gnd.n3594 gnd.n3593 9.69747
R17494 gnd.n3563 gnd.n3562 9.69747
R17495 gnd.n3531 gnd.n3530 9.69747
R17496 gnd.n3499 gnd.n3498 9.69747
R17497 gnd.n3467 gnd.n3466 9.69747
R17498 gnd.n3436 gnd.n3435 9.69747
R17499 gnd.n5517 gnd.n1866 9.56018
R17500 gnd.n5549 gnd.t132 9.56018
R17501 gnd.n4796 gnd.n4795 9.56018
R17502 gnd.n5637 gnd.n1762 9.56018
R17503 gnd.n4863 gnd.t119 9.56018
R17504 gnd.t333 gnd.n1698 9.56018
R17505 gnd.n6257 gnd.n1115 9.45751
R17506 gnd.n1517 gnd.n1342 9.45599
R17507 gnd.n3664 gnd.n3663 9.45567
R17508 gnd.n3632 gnd.n3631 9.45567
R17509 gnd.n3600 gnd.n3599 9.45567
R17510 gnd.n3569 gnd.n3568 9.45567
R17511 gnd.n3537 gnd.n3536 9.45567
R17512 gnd.n3505 gnd.n3504 9.45567
R17513 gnd.n3473 gnd.n3472 9.45567
R17514 gnd.n3442 gnd.n3441 9.45567
R17515 gnd.n2610 gnd.n2609 9.39724
R17516 gnd.n3663 gnd.n3662 9.3005
R17517 gnd.n3636 gnd.n3635 9.3005
R17518 gnd.n3657 gnd.n3656 9.3005
R17519 gnd.n3655 gnd.n3654 9.3005
R17520 gnd.n3640 gnd.n3639 9.3005
R17521 gnd.n3649 gnd.n3648 9.3005
R17522 gnd.n3647 gnd.n3646 9.3005
R17523 gnd.n3631 gnd.n3630 9.3005
R17524 gnd.n3604 gnd.n3603 9.3005
R17525 gnd.n3625 gnd.n3624 9.3005
R17526 gnd.n3623 gnd.n3622 9.3005
R17527 gnd.n3608 gnd.n3607 9.3005
R17528 gnd.n3617 gnd.n3616 9.3005
R17529 gnd.n3615 gnd.n3614 9.3005
R17530 gnd.n3599 gnd.n3598 9.3005
R17531 gnd.n3572 gnd.n3571 9.3005
R17532 gnd.n3593 gnd.n3592 9.3005
R17533 gnd.n3591 gnd.n3590 9.3005
R17534 gnd.n3576 gnd.n3575 9.3005
R17535 gnd.n3585 gnd.n3584 9.3005
R17536 gnd.n3583 gnd.n3582 9.3005
R17537 gnd.n3568 gnd.n3567 9.3005
R17538 gnd.n3541 gnd.n3540 9.3005
R17539 gnd.n3562 gnd.n3561 9.3005
R17540 gnd.n3560 gnd.n3559 9.3005
R17541 gnd.n3545 gnd.n3544 9.3005
R17542 gnd.n3554 gnd.n3553 9.3005
R17543 gnd.n3552 gnd.n3551 9.3005
R17544 gnd.n3536 gnd.n3535 9.3005
R17545 gnd.n3509 gnd.n3508 9.3005
R17546 gnd.n3530 gnd.n3529 9.3005
R17547 gnd.n3528 gnd.n3527 9.3005
R17548 gnd.n3513 gnd.n3512 9.3005
R17549 gnd.n3522 gnd.n3521 9.3005
R17550 gnd.n3520 gnd.n3519 9.3005
R17551 gnd.n3504 gnd.n3503 9.3005
R17552 gnd.n3477 gnd.n3476 9.3005
R17553 gnd.n3498 gnd.n3497 9.3005
R17554 gnd.n3496 gnd.n3495 9.3005
R17555 gnd.n3481 gnd.n3480 9.3005
R17556 gnd.n3490 gnd.n3489 9.3005
R17557 gnd.n3488 gnd.n3487 9.3005
R17558 gnd.n3472 gnd.n3471 9.3005
R17559 gnd.n3445 gnd.n3444 9.3005
R17560 gnd.n3466 gnd.n3465 9.3005
R17561 gnd.n3464 gnd.n3463 9.3005
R17562 gnd.n3449 gnd.n3448 9.3005
R17563 gnd.n3458 gnd.n3457 9.3005
R17564 gnd.n3456 gnd.n3455 9.3005
R17565 gnd.n3441 gnd.n3440 9.3005
R17566 gnd.n3414 gnd.n3413 9.3005
R17567 gnd.n3435 gnd.n3434 9.3005
R17568 gnd.n3433 gnd.n3432 9.3005
R17569 gnd.n3418 gnd.n3417 9.3005
R17570 gnd.n3427 gnd.n3426 9.3005
R17571 gnd.n3425 gnd.n3424 9.3005
R17572 gnd.n3789 gnd.n3788 9.3005
R17573 gnd.n3787 gnd.n2344 9.3005
R17574 gnd.n3786 gnd.n3785 9.3005
R17575 gnd.n3782 gnd.n2345 9.3005
R17576 gnd.n3779 gnd.n2346 9.3005
R17577 gnd.n3778 gnd.n2347 9.3005
R17578 gnd.n3775 gnd.n2348 9.3005
R17579 gnd.n3774 gnd.n2349 9.3005
R17580 gnd.n3771 gnd.n2350 9.3005
R17581 gnd.n3770 gnd.n2351 9.3005
R17582 gnd.n3767 gnd.n2352 9.3005
R17583 gnd.n3766 gnd.n2353 9.3005
R17584 gnd.n3763 gnd.n2354 9.3005
R17585 gnd.n3762 gnd.n2355 9.3005
R17586 gnd.n3759 gnd.n3758 9.3005
R17587 gnd.n3757 gnd.n2356 9.3005
R17588 gnd.n3790 gnd.n2343 9.3005
R17589 gnd.n3031 gnd.n3030 9.3005
R17590 gnd.n2735 gnd.n2734 9.3005
R17591 gnd.n3058 gnd.n3057 9.3005
R17592 gnd.n3059 gnd.n2733 9.3005
R17593 gnd.n3063 gnd.n3060 9.3005
R17594 gnd.n3062 gnd.n3061 9.3005
R17595 gnd.n2707 gnd.n2706 9.3005
R17596 gnd.n3088 gnd.n3087 9.3005
R17597 gnd.n3089 gnd.n2705 9.3005
R17598 gnd.n3091 gnd.n3090 9.3005
R17599 gnd.n2685 gnd.n2684 9.3005
R17600 gnd.n3119 gnd.n3118 9.3005
R17601 gnd.n3120 gnd.n2683 9.3005
R17602 gnd.n3128 gnd.n3121 9.3005
R17603 gnd.n3127 gnd.n3122 9.3005
R17604 gnd.n3126 gnd.n3124 9.3005
R17605 gnd.n3123 gnd.n2632 9.3005
R17606 gnd.n3176 gnd.n2633 9.3005
R17607 gnd.n3175 gnd.n2634 9.3005
R17608 gnd.n3174 gnd.n2635 9.3005
R17609 gnd.n2654 gnd.n2636 9.3005
R17610 gnd.n2656 gnd.n2655 9.3005
R17611 gnd.n2542 gnd.n2541 9.3005
R17612 gnd.n3214 gnd.n3213 9.3005
R17613 gnd.n3215 gnd.n2540 9.3005
R17614 gnd.n3219 gnd.n3216 9.3005
R17615 gnd.n3218 gnd.n3217 9.3005
R17616 gnd.n2515 gnd.n2514 9.3005
R17617 gnd.n3254 gnd.n3253 9.3005
R17618 gnd.n3255 gnd.n2513 9.3005
R17619 gnd.n3259 gnd.n3256 9.3005
R17620 gnd.n3258 gnd.n3257 9.3005
R17621 gnd.n2488 gnd.n2487 9.3005
R17622 gnd.n3299 gnd.n3298 9.3005
R17623 gnd.n3300 gnd.n2486 9.3005
R17624 gnd.n3304 gnd.n3301 9.3005
R17625 gnd.n3303 gnd.n3302 9.3005
R17626 gnd.n2460 gnd.n2459 9.3005
R17627 gnd.n3339 gnd.n3338 9.3005
R17628 gnd.n3340 gnd.n2458 9.3005
R17629 gnd.n3344 gnd.n3341 9.3005
R17630 gnd.n3343 gnd.n3342 9.3005
R17631 gnd.n2433 gnd.n2432 9.3005
R17632 gnd.n3388 gnd.n3387 9.3005
R17633 gnd.n3389 gnd.n2431 9.3005
R17634 gnd.n3393 gnd.n3390 9.3005
R17635 gnd.n3392 gnd.n3391 9.3005
R17636 gnd.n2406 gnd.n2405 9.3005
R17637 gnd.n3682 gnd.n3681 9.3005
R17638 gnd.n3683 gnd.n2404 9.3005
R17639 gnd.n3689 gnd.n3684 9.3005
R17640 gnd.n3688 gnd.n3685 9.3005
R17641 gnd.n3687 gnd.n3686 9.3005
R17642 gnd.n3032 gnd.n3029 9.3005
R17643 gnd.n2814 gnd.n2773 9.3005
R17644 gnd.n2809 gnd.n2808 9.3005
R17645 gnd.n2807 gnd.n2774 9.3005
R17646 gnd.n2806 gnd.n2805 9.3005
R17647 gnd.n2802 gnd.n2775 9.3005
R17648 gnd.n2799 gnd.n2798 9.3005
R17649 gnd.n2797 gnd.n2776 9.3005
R17650 gnd.n2796 gnd.n2795 9.3005
R17651 gnd.n2792 gnd.n2777 9.3005
R17652 gnd.n2789 gnd.n2788 9.3005
R17653 gnd.n2787 gnd.n2778 9.3005
R17654 gnd.n2786 gnd.n2785 9.3005
R17655 gnd.n2782 gnd.n2780 9.3005
R17656 gnd.n2779 gnd.n2759 9.3005
R17657 gnd.n3026 gnd.n2758 9.3005
R17658 gnd.n3028 gnd.n3027 9.3005
R17659 gnd.n2816 gnd.n2815 9.3005
R17660 gnd.n3039 gnd.n2745 9.3005
R17661 gnd.n3046 gnd.n2746 9.3005
R17662 gnd.n3048 gnd.n3047 9.3005
R17663 gnd.n3049 gnd.n2726 9.3005
R17664 gnd.n3068 gnd.n3067 9.3005
R17665 gnd.n3070 gnd.n2718 9.3005
R17666 gnd.n3077 gnd.n2720 9.3005
R17667 gnd.n3078 gnd.n2715 9.3005
R17668 gnd.n3080 gnd.n3079 9.3005
R17669 gnd.n2716 gnd.n2701 9.3005
R17670 gnd.n3096 gnd.n2699 9.3005
R17671 gnd.n3100 gnd.n3099 9.3005
R17672 gnd.n3098 gnd.n2675 9.3005
R17673 gnd.n3135 gnd.n2674 9.3005
R17674 gnd.n3138 gnd.n3137 9.3005
R17675 gnd.n2671 gnd.n2670 9.3005
R17676 gnd.n3144 gnd.n2672 9.3005
R17677 gnd.n3146 gnd.n3145 9.3005
R17678 gnd.n3148 gnd.n2669 9.3005
R17679 gnd.n3151 gnd.n3150 9.3005
R17680 gnd.n3154 gnd.n3152 9.3005
R17681 gnd.n3156 gnd.n3155 9.3005
R17682 gnd.n3162 gnd.n3157 9.3005
R17683 gnd.n3161 gnd.n3160 9.3005
R17684 gnd.n2533 gnd.n2532 9.3005
R17685 gnd.n3228 gnd.n3227 9.3005
R17686 gnd.n3229 gnd.n2526 9.3005
R17687 gnd.n3237 gnd.n2525 9.3005
R17688 gnd.n3240 gnd.n3239 9.3005
R17689 gnd.n3242 gnd.n3241 9.3005
R17690 gnd.n3245 gnd.n2508 9.3005
R17691 gnd.n3243 gnd.n2506 9.3005
R17692 gnd.n3265 gnd.n2504 9.3005
R17693 gnd.n3267 gnd.n3266 9.3005
R17694 gnd.n2478 gnd.n2477 9.3005
R17695 gnd.n3313 gnd.n3312 9.3005
R17696 gnd.n3314 gnd.n2471 9.3005
R17697 gnd.n3322 gnd.n2470 9.3005
R17698 gnd.n3325 gnd.n3324 9.3005
R17699 gnd.n3327 gnd.n3326 9.3005
R17700 gnd.n3330 gnd.n2453 9.3005
R17701 gnd.n3328 gnd.n2451 9.3005
R17702 gnd.n3350 gnd.n2449 9.3005
R17703 gnd.n3352 gnd.n3351 9.3005
R17704 gnd.n2424 gnd.n2423 9.3005
R17705 gnd.n3402 gnd.n3401 9.3005
R17706 gnd.n3403 gnd.n2417 9.3005
R17707 gnd.n3411 gnd.n2416 9.3005
R17708 gnd.n3670 gnd.n3669 9.3005
R17709 gnd.n3672 gnd.n3671 9.3005
R17710 gnd.n3673 gnd.n2397 9.3005
R17711 gnd.n3697 gnd.n3696 9.3005
R17712 gnd.n2398 gnd.n2359 9.3005
R17713 gnd.n3037 gnd.n3036 9.3005
R17714 gnd.n3753 gnd.n2360 9.3005
R17715 gnd.n3752 gnd.n2362 9.3005
R17716 gnd.n3749 gnd.n2363 9.3005
R17717 gnd.n3748 gnd.n2364 9.3005
R17718 gnd.n3745 gnd.n2365 9.3005
R17719 gnd.n3744 gnd.n2366 9.3005
R17720 gnd.n3741 gnd.n2367 9.3005
R17721 gnd.n3740 gnd.n2368 9.3005
R17722 gnd.n3737 gnd.n2369 9.3005
R17723 gnd.n3736 gnd.n2370 9.3005
R17724 gnd.n3733 gnd.n2371 9.3005
R17725 gnd.n3732 gnd.n2372 9.3005
R17726 gnd.n3729 gnd.n2373 9.3005
R17727 gnd.n3728 gnd.n2374 9.3005
R17728 gnd.n3725 gnd.n2375 9.3005
R17729 gnd.n3724 gnd.n2376 9.3005
R17730 gnd.n3721 gnd.n2377 9.3005
R17731 gnd.n3720 gnd.n2378 9.3005
R17732 gnd.n3717 gnd.n2379 9.3005
R17733 gnd.n3716 gnd.n2380 9.3005
R17734 gnd.n3713 gnd.n2381 9.3005
R17735 gnd.n3712 gnd.n2382 9.3005
R17736 gnd.n3709 gnd.n2386 9.3005
R17737 gnd.n3708 gnd.n2387 9.3005
R17738 gnd.n3705 gnd.n2388 9.3005
R17739 gnd.n3704 gnd.n2389 9.3005
R17740 gnd.n3755 gnd.n3754 9.3005
R17741 gnd.n3206 gnd.n3190 9.3005
R17742 gnd.n3205 gnd.n3191 9.3005
R17743 gnd.n3204 gnd.n3192 9.3005
R17744 gnd.n3202 gnd.n3193 9.3005
R17745 gnd.n3201 gnd.n3194 9.3005
R17746 gnd.n3199 gnd.n3195 9.3005
R17747 gnd.n3198 gnd.n3196 9.3005
R17748 gnd.n2496 gnd.n2495 9.3005
R17749 gnd.n3275 gnd.n3274 9.3005
R17750 gnd.n3276 gnd.n2494 9.3005
R17751 gnd.n3293 gnd.n3277 9.3005
R17752 gnd.n3292 gnd.n3278 9.3005
R17753 gnd.n3291 gnd.n3279 9.3005
R17754 gnd.n3289 gnd.n3280 9.3005
R17755 gnd.n3288 gnd.n3281 9.3005
R17756 gnd.n3286 gnd.n3282 9.3005
R17757 gnd.n3285 gnd.n3283 9.3005
R17758 gnd.n2440 gnd.n2439 9.3005
R17759 gnd.n3360 gnd.n3359 9.3005
R17760 gnd.n3361 gnd.n2438 9.3005
R17761 gnd.n3382 gnd.n3362 9.3005
R17762 gnd.n3381 gnd.n3363 9.3005
R17763 gnd.n3380 gnd.n3364 9.3005
R17764 gnd.n3377 gnd.n3365 9.3005
R17765 gnd.n3376 gnd.n3366 9.3005
R17766 gnd.n3374 gnd.n3367 9.3005
R17767 gnd.n3373 gnd.n3368 9.3005
R17768 gnd.n3371 gnd.n3370 9.3005
R17769 gnd.n3369 gnd.n2391 9.3005
R17770 gnd.n2947 gnd.n2946 9.3005
R17771 gnd.n2837 gnd.n2836 9.3005
R17772 gnd.n2961 gnd.n2960 9.3005
R17773 gnd.n2962 gnd.n2835 9.3005
R17774 gnd.n2964 gnd.n2963 9.3005
R17775 gnd.n2825 gnd.n2824 9.3005
R17776 gnd.n2977 gnd.n2976 9.3005
R17777 gnd.n2978 gnd.n2823 9.3005
R17778 gnd.n3010 gnd.n2979 9.3005
R17779 gnd.n3009 gnd.n2980 9.3005
R17780 gnd.n3008 gnd.n2981 9.3005
R17781 gnd.n3007 gnd.n2982 9.3005
R17782 gnd.n3004 gnd.n2983 9.3005
R17783 gnd.n3003 gnd.n2984 9.3005
R17784 gnd.n3002 gnd.n2985 9.3005
R17785 gnd.n3000 gnd.n2986 9.3005
R17786 gnd.n2999 gnd.n2987 9.3005
R17787 gnd.n2996 gnd.n2988 9.3005
R17788 gnd.n2995 gnd.n2989 9.3005
R17789 gnd.n2994 gnd.n2990 9.3005
R17790 gnd.n2992 gnd.n2991 9.3005
R17791 gnd.n2691 gnd.n2690 9.3005
R17792 gnd.n3108 gnd.n3107 9.3005
R17793 gnd.n3109 gnd.n2689 9.3005
R17794 gnd.n3113 gnd.n3110 9.3005
R17795 gnd.n3112 gnd.n3111 9.3005
R17796 gnd.n2613 gnd.n2612 9.3005
R17797 gnd.n3188 gnd.n3187 9.3005
R17798 gnd.n2945 gnd.n2846 9.3005
R17799 gnd.n2848 gnd.n2847 9.3005
R17800 gnd.n2892 gnd.n2890 9.3005
R17801 gnd.n2893 gnd.n2889 9.3005
R17802 gnd.n2896 gnd.n2885 9.3005
R17803 gnd.n2897 gnd.n2884 9.3005
R17804 gnd.n2900 gnd.n2883 9.3005
R17805 gnd.n2901 gnd.n2882 9.3005
R17806 gnd.n2904 gnd.n2881 9.3005
R17807 gnd.n2905 gnd.n2880 9.3005
R17808 gnd.n2908 gnd.n2879 9.3005
R17809 gnd.n2909 gnd.n2878 9.3005
R17810 gnd.n2912 gnd.n2877 9.3005
R17811 gnd.n2913 gnd.n2876 9.3005
R17812 gnd.n2916 gnd.n2875 9.3005
R17813 gnd.n2917 gnd.n2874 9.3005
R17814 gnd.n2920 gnd.n2873 9.3005
R17815 gnd.n2921 gnd.n2872 9.3005
R17816 gnd.n2924 gnd.n2871 9.3005
R17817 gnd.n2925 gnd.n2870 9.3005
R17818 gnd.n2928 gnd.n2869 9.3005
R17819 gnd.n2929 gnd.n2868 9.3005
R17820 gnd.n2932 gnd.n2867 9.3005
R17821 gnd.n2934 gnd.n2866 9.3005
R17822 gnd.n2935 gnd.n2865 9.3005
R17823 gnd.n2936 gnd.n2864 9.3005
R17824 gnd.n2937 gnd.n2863 9.3005
R17825 gnd.n2944 gnd.n2943 9.3005
R17826 gnd.n2953 gnd.n2952 9.3005
R17827 gnd.n2954 gnd.n2840 9.3005
R17828 gnd.n2956 gnd.n2955 9.3005
R17829 gnd.n2831 gnd.n2830 9.3005
R17830 gnd.n2969 gnd.n2968 9.3005
R17831 gnd.n2970 gnd.n2829 9.3005
R17832 gnd.n2972 gnd.n2971 9.3005
R17833 gnd.n2818 gnd.n2817 9.3005
R17834 gnd.n3015 gnd.n3014 9.3005
R17835 gnd.n3016 gnd.n2772 9.3005
R17836 gnd.n3020 gnd.n3018 9.3005
R17837 gnd.n3019 gnd.n2751 9.3005
R17838 gnd.n3038 gnd.n2750 9.3005
R17839 gnd.n3041 gnd.n3040 9.3005
R17840 gnd.n2744 gnd.n2743 9.3005
R17841 gnd.n3052 gnd.n3050 9.3005
R17842 gnd.n3051 gnd.n2725 9.3005
R17843 gnd.n3069 gnd.n2724 9.3005
R17844 gnd.n3072 gnd.n3071 9.3005
R17845 gnd.n2719 gnd.n2714 9.3005
R17846 gnd.n3082 gnd.n3081 9.3005
R17847 gnd.n2717 gnd.n2697 9.3005
R17848 gnd.n3103 gnd.n2698 9.3005
R17849 gnd.n3102 gnd.n3101 9.3005
R17850 gnd.n2700 gnd.n2676 9.3005
R17851 gnd.n3134 gnd.n3133 9.3005
R17852 gnd.n3136 gnd.n2621 9.3005
R17853 gnd.n3183 gnd.n2622 9.3005
R17854 gnd.n3182 gnd.n2623 9.3005
R17855 gnd.n3181 gnd.n2624 9.3005
R17856 gnd.n3147 gnd.n2625 9.3005
R17857 gnd.n3149 gnd.n2643 9.3005
R17858 gnd.n3169 gnd.n2644 9.3005
R17859 gnd.n3168 gnd.n2645 9.3005
R17860 gnd.n3167 gnd.n2646 9.3005
R17861 gnd.n3158 gnd.n2647 9.3005
R17862 gnd.n3159 gnd.n2534 9.3005
R17863 gnd.n3225 gnd.n3224 9.3005
R17864 gnd.n3226 gnd.n2527 9.3005
R17865 gnd.n3236 gnd.n3235 9.3005
R17866 gnd.n3238 gnd.n2523 9.3005
R17867 gnd.n3248 gnd.n2524 9.3005
R17868 gnd.n3247 gnd.n3246 9.3005
R17869 gnd.n3244 gnd.n2502 9.3005
R17870 gnd.n3270 gnd.n2503 9.3005
R17871 gnd.n3269 gnd.n3268 9.3005
R17872 gnd.n2505 gnd.n2479 9.3005
R17873 gnd.n3310 gnd.n3309 9.3005
R17874 gnd.n3311 gnd.n2472 9.3005
R17875 gnd.n3321 gnd.n3320 9.3005
R17876 gnd.n3323 gnd.n2468 9.3005
R17877 gnd.n3333 gnd.n2469 9.3005
R17878 gnd.n3332 gnd.n3331 9.3005
R17879 gnd.n3329 gnd.n2447 9.3005
R17880 gnd.n3355 gnd.n2448 9.3005
R17881 gnd.n3354 gnd.n3353 9.3005
R17882 gnd.n2450 gnd.n2425 9.3005
R17883 gnd.n3399 gnd.n3398 9.3005
R17884 gnd.n3400 gnd.n2418 9.3005
R17885 gnd.n3410 gnd.n3409 9.3005
R17886 gnd.n3668 gnd.n2414 9.3005
R17887 gnd.n3676 gnd.n2415 9.3005
R17888 gnd.n3675 gnd.n3674 9.3005
R17889 gnd.n2396 gnd.n2395 9.3005
R17890 gnd.n3699 gnd.n3698 9.3005
R17891 gnd.n2842 gnd.n2841 9.3005
R17892 gnd.n6517 gnd.n6516 9.3005
R17893 gnd.n795 gnd.n794 9.3005
R17894 gnd.n6524 gnd.n6523 9.3005
R17895 gnd.n6525 gnd.n793 9.3005
R17896 gnd.n6527 gnd.n6526 9.3005
R17897 gnd.n789 gnd.n788 9.3005
R17898 gnd.n6534 gnd.n6533 9.3005
R17899 gnd.n6535 gnd.n787 9.3005
R17900 gnd.n6537 gnd.n6536 9.3005
R17901 gnd.n783 gnd.n782 9.3005
R17902 gnd.n6544 gnd.n6543 9.3005
R17903 gnd.n6545 gnd.n781 9.3005
R17904 gnd.n6547 gnd.n6546 9.3005
R17905 gnd.n777 gnd.n776 9.3005
R17906 gnd.n6554 gnd.n6553 9.3005
R17907 gnd.n6555 gnd.n775 9.3005
R17908 gnd.n6557 gnd.n6556 9.3005
R17909 gnd.n771 gnd.n770 9.3005
R17910 gnd.n6564 gnd.n6563 9.3005
R17911 gnd.n6565 gnd.n769 9.3005
R17912 gnd.n6567 gnd.n6566 9.3005
R17913 gnd.n765 gnd.n764 9.3005
R17914 gnd.n6574 gnd.n6573 9.3005
R17915 gnd.n6575 gnd.n763 9.3005
R17916 gnd.n6577 gnd.n6576 9.3005
R17917 gnd.n759 gnd.n758 9.3005
R17918 gnd.n6584 gnd.n6583 9.3005
R17919 gnd.n6585 gnd.n757 9.3005
R17920 gnd.n6587 gnd.n6586 9.3005
R17921 gnd.n753 gnd.n752 9.3005
R17922 gnd.n6594 gnd.n6593 9.3005
R17923 gnd.n6595 gnd.n751 9.3005
R17924 gnd.n6597 gnd.n6596 9.3005
R17925 gnd.n747 gnd.n746 9.3005
R17926 gnd.n6604 gnd.n6603 9.3005
R17927 gnd.n6605 gnd.n745 9.3005
R17928 gnd.n6607 gnd.n6606 9.3005
R17929 gnd.n741 gnd.n740 9.3005
R17930 gnd.n6614 gnd.n6613 9.3005
R17931 gnd.n6615 gnd.n739 9.3005
R17932 gnd.n6617 gnd.n6616 9.3005
R17933 gnd.n735 gnd.n734 9.3005
R17934 gnd.n6624 gnd.n6623 9.3005
R17935 gnd.n6625 gnd.n733 9.3005
R17936 gnd.n6627 gnd.n6626 9.3005
R17937 gnd.n729 gnd.n728 9.3005
R17938 gnd.n6634 gnd.n6633 9.3005
R17939 gnd.n6635 gnd.n727 9.3005
R17940 gnd.n6637 gnd.n6636 9.3005
R17941 gnd.n723 gnd.n722 9.3005
R17942 gnd.n6644 gnd.n6643 9.3005
R17943 gnd.n6645 gnd.n721 9.3005
R17944 gnd.n6647 gnd.n6646 9.3005
R17945 gnd.n717 gnd.n716 9.3005
R17946 gnd.n6654 gnd.n6653 9.3005
R17947 gnd.n6655 gnd.n715 9.3005
R17948 gnd.n6657 gnd.n6656 9.3005
R17949 gnd.n711 gnd.n710 9.3005
R17950 gnd.n6664 gnd.n6663 9.3005
R17951 gnd.n6665 gnd.n709 9.3005
R17952 gnd.n6667 gnd.n6666 9.3005
R17953 gnd.n705 gnd.n704 9.3005
R17954 gnd.n6674 gnd.n6673 9.3005
R17955 gnd.n6675 gnd.n703 9.3005
R17956 gnd.n6677 gnd.n6676 9.3005
R17957 gnd.n699 gnd.n698 9.3005
R17958 gnd.n6684 gnd.n6683 9.3005
R17959 gnd.n6685 gnd.n697 9.3005
R17960 gnd.n6687 gnd.n6686 9.3005
R17961 gnd.n693 gnd.n692 9.3005
R17962 gnd.n6694 gnd.n6693 9.3005
R17963 gnd.n6695 gnd.n691 9.3005
R17964 gnd.n6697 gnd.n6696 9.3005
R17965 gnd.n687 gnd.n686 9.3005
R17966 gnd.n6704 gnd.n6703 9.3005
R17967 gnd.n6705 gnd.n685 9.3005
R17968 gnd.n6707 gnd.n6706 9.3005
R17969 gnd.n681 gnd.n680 9.3005
R17970 gnd.n6714 gnd.n6713 9.3005
R17971 gnd.n6715 gnd.n679 9.3005
R17972 gnd.n6717 gnd.n6716 9.3005
R17973 gnd.n675 gnd.n674 9.3005
R17974 gnd.n6724 gnd.n6723 9.3005
R17975 gnd.n6725 gnd.n673 9.3005
R17976 gnd.n6727 gnd.n6726 9.3005
R17977 gnd.n669 gnd.n668 9.3005
R17978 gnd.n6734 gnd.n6733 9.3005
R17979 gnd.n6735 gnd.n667 9.3005
R17980 gnd.n6737 gnd.n6736 9.3005
R17981 gnd.n663 gnd.n662 9.3005
R17982 gnd.n6744 gnd.n6743 9.3005
R17983 gnd.n6745 gnd.n661 9.3005
R17984 gnd.n6747 gnd.n6746 9.3005
R17985 gnd.n657 gnd.n656 9.3005
R17986 gnd.n6754 gnd.n6753 9.3005
R17987 gnd.n6755 gnd.n655 9.3005
R17988 gnd.n6757 gnd.n6756 9.3005
R17989 gnd.n651 gnd.n650 9.3005
R17990 gnd.n6764 gnd.n6763 9.3005
R17991 gnd.n6765 gnd.n649 9.3005
R17992 gnd.n6767 gnd.n6766 9.3005
R17993 gnd.n645 gnd.n644 9.3005
R17994 gnd.n6774 gnd.n6773 9.3005
R17995 gnd.n6775 gnd.n643 9.3005
R17996 gnd.n6777 gnd.n6776 9.3005
R17997 gnd.n639 gnd.n638 9.3005
R17998 gnd.n6784 gnd.n6783 9.3005
R17999 gnd.n6785 gnd.n637 9.3005
R18000 gnd.n6787 gnd.n6786 9.3005
R18001 gnd.n633 gnd.n632 9.3005
R18002 gnd.n6794 gnd.n6793 9.3005
R18003 gnd.n6795 gnd.n631 9.3005
R18004 gnd.n6797 gnd.n6796 9.3005
R18005 gnd.n627 gnd.n626 9.3005
R18006 gnd.n6804 gnd.n6803 9.3005
R18007 gnd.n6805 gnd.n625 9.3005
R18008 gnd.n6807 gnd.n6806 9.3005
R18009 gnd.n621 gnd.n620 9.3005
R18010 gnd.n6814 gnd.n6813 9.3005
R18011 gnd.n6815 gnd.n619 9.3005
R18012 gnd.n6817 gnd.n6816 9.3005
R18013 gnd.n615 gnd.n614 9.3005
R18014 gnd.n6824 gnd.n6823 9.3005
R18015 gnd.n6825 gnd.n613 9.3005
R18016 gnd.n6827 gnd.n6826 9.3005
R18017 gnd.n609 gnd.n608 9.3005
R18018 gnd.n6834 gnd.n6833 9.3005
R18019 gnd.n6835 gnd.n607 9.3005
R18020 gnd.n6837 gnd.n6836 9.3005
R18021 gnd.n603 gnd.n602 9.3005
R18022 gnd.n6844 gnd.n6843 9.3005
R18023 gnd.n6845 gnd.n601 9.3005
R18024 gnd.n6847 gnd.n6846 9.3005
R18025 gnd.n597 gnd.n596 9.3005
R18026 gnd.n6854 gnd.n6853 9.3005
R18027 gnd.n6855 gnd.n595 9.3005
R18028 gnd.n6857 gnd.n6856 9.3005
R18029 gnd.n591 gnd.n590 9.3005
R18030 gnd.n6864 gnd.n6863 9.3005
R18031 gnd.n6865 gnd.n589 9.3005
R18032 gnd.n6867 gnd.n6866 9.3005
R18033 gnd.n585 gnd.n584 9.3005
R18034 gnd.n6874 gnd.n6873 9.3005
R18035 gnd.n6875 gnd.n583 9.3005
R18036 gnd.n6877 gnd.n6876 9.3005
R18037 gnd.n579 gnd.n578 9.3005
R18038 gnd.n6884 gnd.n6883 9.3005
R18039 gnd.n6885 gnd.n577 9.3005
R18040 gnd.n6887 gnd.n6886 9.3005
R18041 gnd.n573 gnd.n572 9.3005
R18042 gnd.n6894 gnd.n6893 9.3005
R18043 gnd.n6895 gnd.n571 9.3005
R18044 gnd.n6897 gnd.n6896 9.3005
R18045 gnd.n567 gnd.n566 9.3005
R18046 gnd.n6904 gnd.n6903 9.3005
R18047 gnd.n6905 gnd.n565 9.3005
R18048 gnd.n6907 gnd.n6906 9.3005
R18049 gnd.n561 gnd.n560 9.3005
R18050 gnd.n6914 gnd.n6913 9.3005
R18051 gnd.n6915 gnd.n559 9.3005
R18052 gnd.n6917 gnd.n6916 9.3005
R18053 gnd.n555 gnd.n554 9.3005
R18054 gnd.n6924 gnd.n6923 9.3005
R18055 gnd.n6925 gnd.n553 9.3005
R18056 gnd.n6928 gnd.n6927 9.3005
R18057 gnd.n6926 gnd.n549 9.3005
R18058 gnd.n6934 gnd.n548 9.3005
R18059 gnd.n6936 gnd.n6935 9.3005
R18060 gnd.n544 gnd.n543 9.3005
R18061 gnd.n6945 gnd.n6944 9.3005
R18062 gnd.n6946 gnd.n542 9.3005
R18063 gnd.n6948 gnd.n6947 9.3005
R18064 gnd.n538 gnd.n537 9.3005
R18065 gnd.n6955 gnd.n6954 9.3005
R18066 gnd.n6956 gnd.n536 9.3005
R18067 gnd.n6958 gnd.n6957 9.3005
R18068 gnd.n532 gnd.n531 9.3005
R18069 gnd.n6965 gnd.n6964 9.3005
R18070 gnd.n6966 gnd.n530 9.3005
R18071 gnd.n6968 gnd.n6967 9.3005
R18072 gnd.n526 gnd.n525 9.3005
R18073 gnd.n6975 gnd.n6974 9.3005
R18074 gnd.n6976 gnd.n524 9.3005
R18075 gnd.n6978 gnd.n6977 9.3005
R18076 gnd.n520 gnd.n519 9.3005
R18077 gnd.n6985 gnd.n6984 9.3005
R18078 gnd.n6986 gnd.n518 9.3005
R18079 gnd.n6988 gnd.n6987 9.3005
R18080 gnd.n514 gnd.n513 9.3005
R18081 gnd.n6995 gnd.n6994 9.3005
R18082 gnd.n6996 gnd.n512 9.3005
R18083 gnd.n6998 gnd.n6997 9.3005
R18084 gnd.n508 gnd.n507 9.3005
R18085 gnd.n7005 gnd.n7004 9.3005
R18086 gnd.n7006 gnd.n506 9.3005
R18087 gnd.n7008 gnd.n7007 9.3005
R18088 gnd.n502 gnd.n501 9.3005
R18089 gnd.n7015 gnd.n7014 9.3005
R18090 gnd.n7016 gnd.n500 9.3005
R18091 gnd.n7018 gnd.n7017 9.3005
R18092 gnd.n496 gnd.n495 9.3005
R18093 gnd.n7025 gnd.n7024 9.3005
R18094 gnd.n7026 gnd.n494 9.3005
R18095 gnd.n7028 gnd.n7027 9.3005
R18096 gnd.n490 gnd.n489 9.3005
R18097 gnd.n7035 gnd.n7034 9.3005
R18098 gnd.n7036 gnd.n488 9.3005
R18099 gnd.n7038 gnd.n7037 9.3005
R18100 gnd.n484 gnd.n483 9.3005
R18101 gnd.n7045 gnd.n7044 9.3005
R18102 gnd.n7046 gnd.n482 9.3005
R18103 gnd.n7048 gnd.n7047 9.3005
R18104 gnd.n478 gnd.n477 9.3005
R18105 gnd.n7055 gnd.n7054 9.3005
R18106 gnd.n7056 gnd.n476 9.3005
R18107 gnd.n7058 gnd.n7057 9.3005
R18108 gnd.n472 gnd.n471 9.3005
R18109 gnd.n7065 gnd.n7064 9.3005
R18110 gnd.n7066 gnd.n470 9.3005
R18111 gnd.n7068 gnd.n7067 9.3005
R18112 gnd.n466 gnd.n465 9.3005
R18113 gnd.n7075 gnd.n7074 9.3005
R18114 gnd.n7076 gnd.n464 9.3005
R18115 gnd.n7078 gnd.n7077 9.3005
R18116 gnd.n460 gnd.n459 9.3005
R18117 gnd.n7085 gnd.n7084 9.3005
R18118 gnd.n7086 gnd.n458 9.3005
R18119 gnd.n7088 gnd.n7087 9.3005
R18120 gnd.n454 gnd.n453 9.3005
R18121 gnd.n7095 gnd.n7094 9.3005
R18122 gnd.n7096 gnd.n452 9.3005
R18123 gnd.n7098 gnd.n7097 9.3005
R18124 gnd.n448 gnd.n447 9.3005
R18125 gnd.n7105 gnd.n7104 9.3005
R18126 gnd.n7106 gnd.n446 9.3005
R18127 gnd.n7108 gnd.n7107 9.3005
R18128 gnd.n442 gnd.n441 9.3005
R18129 gnd.n7115 gnd.n7114 9.3005
R18130 gnd.n7116 gnd.n440 9.3005
R18131 gnd.n7118 gnd.n7117 9.3005
R18132 gnd.n436 gnd.n435 9.3005
R18133 gnd.n7125 gnd.n7124 9.3005
R18134 gnd.n7126 gnd.n434 9.3005
R18135 gnd.n7128 gnd.n7127 9.3005
R18136 gnd.n430 gnd.n429 9.3005
R18137 gnd.n7135 gnd.n7134 9.3005
R18138 gnd.n7136 gnd.n428 9.3005
R18139 gnd.n7138 gnd.n7137 9.3005
R18140 gnd.n424 gnd.n423 9.3005
R18141 gnd.n7146 gnd.n7145 9.3005
R18142 gnd.n7147 gnd.n422 9.3005
R18143 gnd.n7149 gnd.n7148 9.3005
R18144 gnd.n6938 gnd.n6937 9.3005
R18145 gnd.n7596 gnd.n134 9.3005
R18146 gnd.n7595 gnd.n136 9.3005
R18147 gnd.n140 gnd.n137 9.3005
R18148 gnd.n7590 gnd.n141 9.3005
R18149 gnd.n7589 gnd.n142 9.3005
R18150 gnd.n7588 gnd.n143 9.3005
R18151 gnd.n147 gnd.n144 9.3005
R18152 gnd.n7583 gnd.n148 9.3005
R18153 gnd.n7582 gnd.n149 9.3005
R18154 gnd.n7581 gnd.n150 9.3005
R18155 gnd.n154 gnd.n151 9.3005
R18156 gnd.n7576 gnd.n155 9.3005
R18157 gnd.n7575 gnd.n156 9.3005
R18158 gnd.n7574 gnd.n157 9.3005
R18159 gnd.n161 gnd.n158 9.3005
R18160 gnd.n7569 gnd.n162 9.3005
R18161 gnd.n7568 gnd.n163 9.3005
R18162 gnd.n7564 gnd.n164 9.3005
R18163 gnd.n168 gnd.n165 9.3005
R18164 gnd.n7559 gnd.n169 9.3005
R18165 gnd.n7558 gnd.n170 9.3005
R18166 gnd.n7557 gnd.n171 9.3005
R18167 gnd.n175 gnd.n172 9.3005
R18168 gnd.n7552 gnd.n176 9.3005
R18169 gnd.n7551 gnd.n177 9.3005
R18170 gnd.n7550 gnd.n178 9.3005
R18171 gnd.n182 gnd.n179 9.3005
R18172 gnd.n7545 gnd.n183 9.3005
R18173 gnd.n7544 gnd.n184 9.3005
R18174 gnd.n7543 gnd.n185 9.3005
R18175 gnd.n189 gnd.n186 9.3005
R18176 gnd.n7538 gnd.n190 9.3005
R18177 gnd.n7537 gnd.n191 9.3005
R18178 gnd.n7536 gnd.n192 9.3005
R18179 gnd.n196 gnd.n193 9.3005
R18180 gnd.n7531 gnd.n197 9.3005
R18181 gnd.n7530 gnd.n7529 9.3005
R18182 gnd.n7528 gnd.n200 9.3005
R18183 gnd.n7598 gnd.n7597 9.3005
R18184 gnd.n1456 gnd.n1455 9.3005
R18185 gnd.n1457 gnd.n1454 9.3005
R18186 gnd.n1473 gnd.n1458 9.3005
R18187 gnd.n1472 gnd.n1459 9.3005
R18188 gnd.n1471 gnd.n1460 9.3005
R18189 gnd.n1469 gnd.n1461 9.3005
R18190 gnd.n1468 gnd.n1462 9.3005
R18191 gnd.n1466 gnd.n1463 9.3005
R18192 gnd.n1465 gnd.n1464 9.3005
R18193 gnd.n1391 gnd.n1390 9.3005
R18194 gnd.n5922 gnd.n5921 9.3005
R18195 gnd.n5923 gnd.n1389 9.3005
R18196 gnd.n5925 gnd.n5924 9.3005
R18197 gnd.n5926 gnd.n1388 9.3005
R18198 gnd.n5929 gnd.n5928 9.3005
R18199 gnd.n5930 gnd.n1387 9.3005
R18200 gnd.n5934 gnd.n5931 9.3005
R18201 gnd.n5933 gnd.n5932 9.3005
R18202 gnd.n388 gnd.n387 9.3005
R18203 gnd.n7185 gnd.n7184 9.3005
R18204 gnd.n7186 gnd.n386 9.3005
R18205 gnd.n7194 gnd.n7187 9.3005
R18206 gnd.n7193 gnd.n7188 9.3005
R18207 gnd.n7192 gnd.n7189 9.3005
R18208 gnd.n354 gnd.n353 9.3005
R18209 gnd.n7230 gnd.n7229 9.3005
R18210 gnd.n7231 gnd.n352 9.3005
R18211 gnd.n7240 gnd.n7232 9.3005
R18212 gnd.n7239 gnd.n7233 9.3005
R18213 gnd.n7238 gnd.n7234 9.3005
R18214 gnd.n7236 gnd.n7235 9.3005
R18215 gnd.n338 gnd.n337 9.3005
R18216 gnd.n7260 gnd.n7259 9.3005
R18217 gnd.n7261 gnd.n336 9.3005
R18218 gnd.n7328 gnd.n7262 9.3005
R18219 gnd.n7327 gnd.n7263 9.3005
R18220 gnd.n7326 gnd.n7264 9.3005
R18221 gnd.n7324 gnd.n7265 9.3005
R18222 gnd.n7323 gnd.n7266 9.3005
R18223 gnd.n7321 gnd.n7267 9.3005
R18224 gnd.n7320 gnd.n7268 9.3005
R18225 gnd.n7318 gnd.n7269 9.3005
R18226 gnd.n7317 gnd.n7270 9.3005
R18227 gnd.n7315 gnd.n7271 9.3005
R18228 gnd.n7314 gnd.n7272 9.3005
R18229 gnd.n7312 gnd.n7273 9.3005
R18230 gnd.n7311 gnd.n7274 9.3005
R18231 gnd.n7309 gnd.n7275 9.3005
R18232 gnd.n7308 gnd.n7276 9.3005
R18233 gnd.n7306 gnd.n7277 9.3005
R18234 gnd.n7305 gnd.n7278 9.3005
R18235 gnd.n7303 gnd.n7279 9.3005
R18236 gnd.n7302 gnd.n7280 9.3005
R18237 gnd.n7300 gnd.n7281 9.3005
R18238 gnd.n7299 gnd.n7282 9.3005
R18239 gnd.n7297 gnd.n7283 9.3005
R18240 gnd.n7296 gnd.n7284 9.3005
R18241 gnd.n7294 gnd.n7285 9.3005
R18242 gnd.n7293 gnd.n7286 9.3005
R18243 gnd.n7291 gnd.n7287 9.3005
R18244 gnd.n7290 gnd.n7289 9.3005
R18245 gnd.n7288 gnd.n204 9.3005
R18246 gnd.n7525 gnd.n203 9.3005
R18247 gnd.n7527 gnd.n7526 9.3005
R18248 gnd.n1335 gnd.n1333 9.3005
R18249 gnd.n6023 gnd.n6022 9.3005
R18250 gnd.n6024 gnd.n1327 9.3005
R18251 gnd.n6027 gnd.n1326 9.3005
R18252 gnd.n6028 gnd.n1325 9.3005
R18253 gnd.n6031 gnd.n1324 9.3005
R18254 gnd.n6032 gnd.n1323 9.3005
R18255 gnd.n6035 gnd.n1322 9.3005
R18256 gnd.n6036 gnd.n1321 9.3005
R18257 gnd.n6039 gnd.n1320 9.3005
R18258 gnd.n6040 gnd.n1319 9.3005
R18259 gnd.n6043 gnd.n1318 9.3005
R18260 gnd.n6044 gnd.n1317 9.3005
R18261 gnd.n6047 gnd.n1316 9.3005
R18262 gnd.n6048 gnd.n1315 9.3005
R18263 gnd.n6051 gnd.n1314 9.3005
R18264 gnd.n6052 gnd.n1313 9.3005
R18265 gnd.n6055 gnd.n1312 9.3005
R18266 gnd.n6056 gnd.n1311 9.3005
R18267 gnd.n6059 gnd.n1310 9.3005
R18268 gnd.n6061 gnd.n1304 9.3005
R18269 gnd.n6064 gnd.n1303 9.3005
R18270 gnd.n6065 gnd.n1302 9.3005
R18271 gnd.n6068 gnd.n1301 9.3005
R18272 gnd.n6069 gnd.n1300 9.3005
R18273 gnd.n6072 gnd.n1299 9.3005
R18274 gnd.n6073 gnd.n1298 9.3005
R18275 gnd.n6076 gnd.n1297 9.3005
R18276 gnd.n6077 gnd.n1296 9.3005
R18277 gnd.n6080 gnd.n1295 9.3005
R18278 gnd.n6081 gnd.n1294 9.3005
R18279 gnd.n6084 gnd.n1293 9.3005
R18280 gnd.n6086 gnd.n1292 9.3005
R18281 gnd.n6087 gnd.n1291 9.3005
R18282 gnd.n6088 gnd.n1290 9.3005
R18283 gnd.n6089 gnd.n1289 9.3005
R18284 gnd.n6021 gnd.n1332 9.3005
R18285 gnd.n6020 gnd.n6019 9.3005
R18286 gnd.n5849 gnd.n5846 9.3005
R18287 gnd.n5848 gnd.n5847 9.3005
R18288 gnd.n1429 gnd.n1428 9.3005
R18289 gnd.n5875 gnd.n5874 9.3005
R18290 gnd.n5876 gnd.n1427 9.3005
R18291 gnd.n5880 gnd.n5877 9.3005
R18292 gnd.n5879 gnd.n5878 9.3005
R18293 gnd.n1402 gnd.n1401 9.3005
R18294 gnd.n5912 gnd.n5911 9.3005
R18295 gnd.n5913 gnd.n1400 9.3005
R18296 gnd.n5917 gnd.n5914 9.3005
R18297 gnd.n5916 gnd.n5915 9.3005
R18298 gnd.n1368 gnd.n1367 9.3005
R18299 gnd.n5982 gnd.n5981 9.3005
R18300 gnd.n5983 gnd.n1366 9.3005
R18301 gnd.n5985 gnd.n5984 9.3005
R18302 gnd.n397 gnd.n396 9.3005
R18303 gnd.n7175 gnd.n7174 9.3005
R18304 gnd.n7176 gnd.n395 9.3005
R18305 gnd.n7180 gnd.n7177 9.3005
R18306 gnd.n7179 gnd.n7178 9.3005
R18307 gnd.n364 gnd.n363 9.3005
R18308 gnd.n7221 gnd.n7220 9.3005
R18309 gnd.n7222 gnd.n362 9.3005
R18310 gnd.n7224 gnd.n7223 9.3005
R18311 gnd.n7225 gnd.n303 9.3005
R18312 gnd.n7356 gnd.n7355 9.3005
R18313 gnd.n288 gnd.n287 9.3005
R18314 gnd.n7369 gnd.n7368 9.3005
R18315 gnd.n7370 gnd.n286 9.3005
R18316 gnd.n7372 gnd.n7371 9.3005
R18317 gnd.n274 gnd.n273 9.3005
R18318 gnd.n7385 gnd.n7384 9.3005
R18319 gnd.n7386 gnd.n272 9.3005
R18320 gnd.n7388 gnd.n7387 9.3005
R18321 gnd.n258 gnd.n257 9.3005
R18322 gnd.n7401 gnd.n7400 9.3005
R18323 gnd.n7402 gnd.n256 9.3005
R18324 gnd.n7404 gnd.n7403 9.3005
R18325 gnd.n243 gnd.n242 9.3005
R18326 gnd.n7417 gnd.n7416 9.3005
R18327 gnd.n7418 gnd.n241 9.3005
R18328 gnd.n7420 gnd.n7419 9.3005
R18329 gnd.n227 gnd.n226 9.3005
R18330 gnd.n7433 gnd.n7432 9.3005
R18331 gnd.n7434 gnd.n225 9.3005
R18332 gnd.n7436 gnd.n7435 9.3005
R18333 gnd.n211 gnd.n210 9.3005
R18334 gnd.n7517 gnd.n7516 9.3005
R18335 gnd.n7518 gnd.n209 9.3005
R18336 gnd.n7520 gnd.n7519 9.3005
R18337 gnd.n133 gnd.n132 9.3005
R18338 gnd.n7600 gnd.n7599 9.3005
R18339 gnd.n5845 gnd.n5844 9.3005
R18340 gnd.n7354 gnd.n302 9.3005
R18341 gnd.n968 gnd.n967 9.3005
R18342 gnd.n4356 gnd.n4355 9.3005
R18343 gnd.n4357 gnd.n4353 9.3005
R18344 gnd.n4359 gnd.n4358 9.3005
R18345 gnd.n2150 gnd.n2149 9.3005
R18346 gnd.n4397 gnd.n4396 9.3005
R18347 gnd.n4398 gnd.n2148 9.3005
R18348 gnd.n4400 gnd.n4399 9.3005
R18349 gnd.n2146 gnd.n2145 9.3005
R18350 gnd.n4405 gnd.n4404 9.3005
R18351 gnd.n4406 gnd.n2144 9.3005
R18352 gnd.n4408 gnd.n4407 9.3005
R18353 gnd.n2129 gnd.n2128 9.3005
R18354 gnd.n4446 gnd.n4445 9.3005
R18355 gnd.n4447 gnd.n2127 9.3005
R18356 gnd.n4449 gnd.n4448 9.3005
R18357 gnd.n2125 gnd.n2124 9.3005
R18358 gnd.n4454 gnd.n4453 9.3005
R18359 gnd.n4455 gnd.n2123 9.3005
R18360 gnd.n4493 gnd.n4456 9.3005
R18361 gnd.n4492 gnd.n4457 9.3005
R18362 gnd.n4491 gnd.n4458 9.3005
R18363 gnd.n4461 gnd.n4459 9.3005
R18364 gnd.n4487 gnd.n4462 9.3005
R18365 gnd.n4486 gnd.n4463 9.3005
R18366 gnd.n4485 gnd.n4464 9.3005
R18367 gnd.n4467 gnd.n4465 9.3005
R18368 gnd.n4481 gnd.n4468 9.3005
R18369 gnd.n4480 gnd.n4469 9.3005
R18370 gnd.n4479 gnd.n4470 9.3005
R18371 gnd.n4472 gnd.n4471 9.3005
R18372 gnd.n4474 gnd.n4473 9.3005
R18373 gnd.n1950 gnd.n1949 9.3005
R18374 gnd.n5416 gnd.n5415 9.3005
R18375 gnd.n5417 gnd.n1948 9.3005
R18376 gnd.n5419 gnd.n5418 9.3005
R18377 gnd.n1936 gnd.n1935 9.3005
R18378 gnd.n5432 gnd.n5431 9.3005
R18379 gnd.n5433 gnd.n1934 9.3005
R18380 gnd.n5435 gnd.n5434 9.3005
R18381 gnd.n1924 gnd.n1923 9.3005
R18382 gnd.n5448 gnd.n5447 9.3005
R18383 gnd.n5449 gnd.n1922 9.3005
R18384 gnd.n5451 gnd.n5450 9.3005
R18385 gnd.n1911 gnd.n1910 9.3005
R18386 gnd.n5464 gnd.n5463 9.3005
R18387 gnd.n5465 gnd.n1909 9.3005
R18388 gnd.n5467 gnd.n5466 9.3005
R18389 gnd.n1898 gnd.n1897 9.3005
R18390 gnd.n5480 gnd.n5479 9.3005
R18391 gnd.n5481 gnd.n1896 9.3005
R18392 gnd.n5483 gnd.n5482 9.3005
R18393 gnd.n1885 gnd.n1884 9.3005
R18394 gnd.n5496 gnd.n5495 9.3005
R18395 gnd.n5497 gnd.n1883 9.3005
R18396 gnd.n5499 gnd.n5498 9.3005
R18397 gnd.n1872 gnd.n1871 9.3005
R18398 gnd.n5512 gnd.n5511 9.3005
R18399 gnd.n5513 gnd.n1870 9.3005
R18400 gnd.n5515 gnd.n5514 9.3005
R18401 gnd.n1857 gnd.n1856 9.3005
R18402 gnd.n5528 gnd.n5527 9.3005
R18403 gnd.n5529 gnd.n1855 9.3005
R18404 gnd.n5531 gnd.n5530 9.3005
R18405 gnd.n1844 gnd.n1843 9.3005
R18406 gnd.n5544 gnd.n5543 9.3005
R18407 gnd.n5545 gnd.n1842 9.3005
R18408 gnd.n5547 gnd.n5546 9.3005
R18409 gnd.n1831 gnd.n1830 9.3005
R18410 gnd.n5560 gnd.n5559 9.3005
R18411 gnd.n5561 gnd.n1829 9.3005
R18412 gnd.n5563 gnd.n5562 9.3005
R18413 gnd.n1816 gnd.n1815 9.3005
R18414 gnd.n5576 gnd.n5575 9.3005
R18415 gnd.n5577 gnd.n1814 9.3005
R18416 gnd.n5579 gnd.n5578 9.3005
R18417 gnd.n1801 gnd.n1800 9.3005
R18418 gnd.n5592 gnd.n5591 9.3005
R18419 gnd.n5593 gnd.n1799 9.3005
R18420 gnd.n5595 gnd.n5594 9.3005
R18421 gnd.n1788 gnd.n1787 9.3005
R18422 gnd.n5608 gnd.n5607 9.3005
R18423 gnd.n5609 gnd.n1786 9.3005
R18424 gnd.n5611 gnd.n5610 9.3005
R18425 gnd.n1774 gnd.n1773 9.3005
R18426 gnd.n5624 gnd.n5623 9.3005
R18427 gnd.n5625 gnd.n1772 9.3005
R18428 gnd.n5627 gnd.n5626 9.3005
R18429 gnd.n1759 gnd.n1758 9.3005
R18430 gnd.n5640 gnd.n5639 9.3005
R18431 gnd.n5641 gnd.n1757 9.3005
R18432 gnd.n5643 gnd.n5642 9.3005
R18433 gnd.n1746 gnd.n1745 9.3005
R18434 gnd.n5656 gnd.n5655 9.3005
R18435 gnd.n5657 gnd.n1744 9.3005
R18436 gnd.n5659 gnd.n5658 9.3005
R18437 gnd.n1731 gnd.n1730 9.3005
R18438 gnd.n5672 gnd.n5671 9.3005
R18439 gnd.n5673 gnd.n1729 9.3005
R18440 gnd.n5675 gnd.n5674 9.3005
R18441 gnd.n1718 gnd.n1717 9.3005
R18442 gnd.n5688 gnd.n5687 9.3005
R18443 gnd.n5689 gnd.n1716 9.3005
R18444 gnd.n5691 gnd.n5690 9.3005
R18445 gnd.n1704 gnd.n1703 9.3005
R18446 gnd.n5704 gnd.n5703 9.3005
R18447 gnd.n5705 gnd.n1702 9.3005
R18448 gnd.n5707 gnd.n5706 9.3005
R18449 gnd.n1690 gnd.n1689 9.3005
R18450 gnd.n5720 gnd.n5719 9.3005
R18451 gnd.n5721 gnd.n1688 9.3005
R18452 gnd.n5723 gnd.n5722 9.3005
R18453 gnd.n1677 gnd.n1676 9.3005
R18454 gnd.n5736 gnd.n5735 9.3005
R18455 gnd.n5737 gnd.n1675 9.3005
R18456 gnd.n5739 gnd.n5738 9.3005
R18457 gnd.n1664 gnd.n1663 9.3005
R18458 gnd.n5752 gnd.n5751 9.3005
R18459 gnd.n5753 gnd.n1662 9.3005
R18460 gnd.n5755 gnd.n5754 9.3005
R18461 gnd.n1651 gnd.n1650 9.3005
R18462 gnd.n5768 gnd.n5767 9.3005
R18463 gnd.n5769 gnd.n1649 9.3005
R18464 gnd.n5771 gnd.n5770 9.3005
R18465 gnd.n1637 gnd.n1636 9.3005
R18466 gnd.n5784 gnd.n5783 9.3005
R18467 gnd.n5785 gnd.n1635 9.3005
R18468 gnd.n5787 gnd.n5786 9.3005
R18469 gnd.n1624 gnd.n1623 9.3005
R18470 gnd.n5802 gnd.n5801 9.3005
R18471 gnd.n5803 gnd.n1622 9.3005
R18472 gnd.n5808 gnd.n5804 9.3005
R18473 gnd.n5807 gnd.n5806 9.3005
R18474 gnd.n5805 gnd.n1250 9.3005
R18475 gnd.n6098 gnd.n1251 9.3005
R18476 gnd.n6097 gnd.n1252 9.3005
R18477 gnd.n6096 gnd.n1253 9.3005
R18478 gnd.n1443 gnd.n1254 9.3005
R18479 gnd.n1446 gnd.n1445 9.3005
R18480 gnd.n1447 gnd.n1442 9.3005
R18481 gnd.n1449 gnd.n1448 9.3005
R18482 gnd.n1440 gnd.n1439 9.3005
R18483 gnd.n5864 gnd.n5863 9.3005
R18484 gnd.n5865 gnd.n1438 9.3005
R18485 gnd.n5869 gnd.n5866 9.3005
R18486 gnd.n5868 gnd.n5867 9.3005
R18487 gnd.n1412 gnd.n1411 9.3005
R18488 gnd.n5900 gnd.n5899 9.3005
R18489 gnd.n5901 gnd.n1410 9.3005
R18490 gnd.n5905 gnd.n5902 9.3005
R18491 gnd.n5904 gnd.n5903 9.3005
R18492 gnd.n1378 gnd.n1377 9.3005
R18493 gnd.n5961 gnd.n5960 9.3005
R18494 gnd.n5962 gnd.n1376 9.3005
R18495 gnd.n5976 gnd.n5963 9.3005
R18496 gnd.n5975 gnd.n5964 9.3005
R18497 gnd.n5974 gnd.n5965 9.3005
R18498 gnd.n5967 gnd.n5966 9.3005
R18499 gnd.n5970 gnd.n5969 9.3005
R18500 gnd.n5968 gnd.n411 9.3005
R18501 gnd.n7160 gnd.n412 9.3005
R18502 gnd.n7159 gnd.n413 9.3005
R18503 gnd.n7158 gnd.n414 9.3005
R18504 gnd.n417 gnd.n415 9.3005
R18505 gnd.n7154 gnd.n418 9.3005
R18506 gnd.n7153 gnd.n419 9.3005
R18507 gnd.n7152 gnd.n420 9.3005
R18508 gnd.n6343 gnd.n6342 9.3005
R18509 gnd.n3909 gnd.n3908 9.3005
R18510 gnd.n3955 gnd.n3864 9.3005
R18511 gnd.n3954 gnd.n3865 9.3005
R18512 gnd.n3953 gnd.n3866 9.3005
R18513 gnd.n3951 gnd.n3867 9.3005
R18514 gnd.n3950 gnd.n3868 9.3005
R18515 gnd.n3948 gnd.n3869 9.3005
R18516 gnd.n3947 gnd.n3870 9.3005
R18517 gnd.n3945 gnd.n3871 9.3005
R18518 gnd.n3944 gnd.n3872 9.3005
R18519 gnd.n3942 gnd.n3873 9.3005
R18520 gnd.n3941 gnd.n3874 9.3005
R18521 gnd.n3939 gnd.n3875 9.3005
R18522 gnd.n3938 gnd.n3876 9.3005
R18523 gnd.n3936 gnd.n3877 9.3005
R18524 gnd.n3935 gnd.n3878 9.3005
R18525 gnd.n3933 gnd.n3879 9.3005
R18526 gnd.n3932 gnd.n3880 9.3005
R18527 gnd.n3930 gnd.n3881 9.3005
R18528 gnd.n3929 gnd.n3882 9.3005
R18529 gnd.n3927 gnd.n3883 9.3005
R18530 gnd.n3926 gnd.n3884 9.3005
R18531 gnd.n3924 gnd.n3885 9.3005
R18532 gnd.n3923 gnd.n3886 9.3005
R18533 gnd.n3921 gnd.n3887 9.3005
R18534 gnd.n3920 gnd.n3888 9.3005
R18535 gnd.n3918 gnd.n3889 9.3005
R18536 gnd.n3917 gnd.n3890 9.3005
R18537 gnd.n3915 gnd.n3891 9.3005
R18538 gnd.n3914 gnd.n3892 9.3005
R18539 gnd.n3912 gnd.n3893 9.3005
R18540 gnd.n3911 gnd.n3894 9.3005
R18541 gnd.n3863 gnd.n3796 9.3005
R18542 gnd.n3856 gnd.n3855 9.3005
R18543 gnd.n3854 gnd.n3802 9.3005
R18544 gnd.n3853 gnd.n3852 9.3005
R18545 gnd.n3804 gnd.n3803 9.3005
R18546 gnd.n3846 gnd.n3845 9.3005
R18547 gnd.n3844 gnd.n3806 9.3005
R18548 gnd.n3843 gnd.n3842 9.3005
R18549 gnd.n3808 gnd.n3807 9.3005
R18550 gnd.n3836 gnd.n3835 9.3005
R18551 gnd.n3834 gnd.n3810 9.3005
R18552 gnd.n3833 gnd.n3832 9.3005
R18553 gnd.n3812 gnd.n3811 9.3005
R18554 gnd.n3826 gnd.n3825 9.3005
R18555 gnd.n3824 gnd.n3814 9.3005
R18556 gnd.n3823 gnd.n3822 9.3005
R18557 gnd.n3817 gnd.n3815 9.3005
R18558 gnd.n3816 gnd.n2317 9.3005
R18559 gnd.n3800 gnd.n3797 9.3005
R18560 gnd.n3862 gnd.n3861 9.3005
R18561 gnd.n4183 gnd.n2316 9.3005
R18562 gnd.n4185 gnd.n4184 9.3005
R18563 gnd.n2303 gnd.n2302 9.3005
R18564 gnd.n4198 gnd.n4197 9.3005
R18565 gnd.n4199 gnd.n2301 9.3005
R18566 gnd.n4201 gnd.n4200 9.3005
R18567 gnd.n2286 gnd.n2285 9.3005
R18568 gnd.n4214 gnd.n4213 9.3005
R18569 gnd.n4215 gnd.n2284 9.3005
R18570 gnd.n4217 gnd.n4216 9.3005
R18571 gnd.n2271 gnd.n2270 9.3005
R18572 gnd.n4230 gnd.n4229 9.3005
R18573 gnd.n4231 gnd.n2269 9.3005
R18574 gnd.n4233 gnd.n4232 9.3005
R18575 gnd.n2254 gnd.n2253 9.3005
R18576 gnd.n4246 gnd.n4245 9.3005
R18577 gnd.n4247 gnd.n2252 9.3005
R18578 gnd.n4249 gnd.n4248 9.3005
R18579 gnd.n2239 gnd.n2238 9.3005
R18580 gnd.n4262 gnd.n4261 9.3005
R18581 gnd.n4263 gnd.n2237 9.3005
R18582 gnd.n4265 gnd.n4264 9.3005
R18583 gnd.n2222 gnd.n2221 9.3005
R18584 gnd.n4279 gnd.n4278 9.3005
R18585 gnd.n4280 gnd.n2220 9.3005
R18586 gnd.n4282 gnd.n4281 9.3005
R18587 gnd.n2208 gnd.n2207 9.3005
R18588 gnd.n4295 gnd.n4294 9.3005
R18589 gnd.n4296 gnd.n2206 9.3005
R18590 gnd.n4299 gnd.n4297 9.3005
R18591 gnd.n4298 gnd.n2182 9.3005
R18592 gnd.n4313 gnd.n2183 9.3005
R18593 gnd.n4314 gnd.n2181 9.3005
R18594 gnd.n4326 gnd.n4315 9.3005
R18595 gnd.n4325 gnd.n4316 9.3005
R18596 gnd.n4324 gnd.n4317 9.3005
R18597 gnd.n4323 gnd.n4318 9.3005
R18598 gnd.n4321 gnd.n4320 9.3005
R18599 gnd.n4319 gnd.n989 9.3005
R18600 gnd.n6331 gnd.n990 9.3005
R18601 gnd.n6330 gnd.n991 9.3005
R18602 gnd.n6329 gnd.n992 9.3005
R18603 gnd.n1009 gnd.n993 9.3005
R18604 gnd.n6319 gnd.n1010 9.3005
R18605 gnd.n6318 gnd.n1011 9.3005
R18606 gnd.n6317 gnd.n1012 9.3005
R18607 gnd.n1031 gnd.n1013 9.3005
R18608 gnd.n6307 gnd.n1032 9.3005
R18609 gnd.n6306 gnd.n1033 9.3005
R18610 gnd.n6305 gnd.n1034 9.3005
R18611 gnd.n1051 gnd.n1035 9.3005
R18612 gnd.n6295 gnd.n1052 9.3005
R18613 gnd.n6294 gnd.n1053 9.3005
R18614 gnd.n6293 gnd.n1054 9.3005
R18615 gnd.n1073 gnd.n1055 9.3005
R18616 gnd.n6283 gnd.n1074 9.3005
R18617 gnd.n6282 gnd.n1075 9.3005
R18618 gnd.n6281 gnd.n1076 9.3005
R18619 gnd.n1094 gnd.n1077 9.3005
R18620 gnd.n6271 gnd.n1095 9.3005
R18621 gnd.n6270 gnd.n1096 9.3005
R18622 gnd.n6269 gnd.n1097 9.3005
R18623 gnd.n1114 gnd.n1098 9.3005
R18624 gnd.n6259 gnd.n6258 9.3005
R18625 gnd.n4182 gnd.n4181 9.3005
R18626 gnd.n5326 gnd.n2081 9.3005
R18627 gnd.n5329 gnd.n2080 9.3005
R18628 gnd.n5330 gnd.n2079 9.3005
R18629 gnd.n5333 gnd.n2078 9.3005
R18630 gnd.n5334 gnd.n2077 9.3005
R18631 gnd.n5337 gnd.n2076 9.3005
R18632 gnd.n5338 gnd.n2075 9.3005
R18633 gnd.n5341 gnd.n2074 9.3005
R18634 gnd.n5342 gnd.n2073 9.3005
R18635 gnd.n5345 gnd.n2072 9.3005
R18636 gnd.n5346 gnd.n2071 9.3005
R18637 gnd.n5349 gnd.n2070 9.3005
R18638 gnd.n5350 gnd.n2069 9.3005
R18639 gnd.n5351 gnd.n2068 9.3005
R18640 gnd.n2067 gnd.n2064 9.3005
R18641 gnd.n2066 gnd.n2065 9.3005
R18642 gnd.n4599 gnd.n4598 9.3005
R18643 gnd.n4595 gnd.n2086 9.3005
R18644 gnd.n4592 gnd.n2087 9.3005
R18645 gnd.n4591 gnd.n2088 9.3005
R18646 gnd.n4588 gnd.n2089 9.3005
R18647 gnd.n4587 gnd.n2090 9.3005
R18648 gnd.n4584 gnd.n2091 9.3005
R18649 gnd.n4583 gnd.n2092 9.3005
R18650 gnd.n4580 gnd.n2093 9.3005
R18651 gnd.n4579 gnd.n2094 9.3005
R18652 gnd.n4576 gnd.n2095 9.3005
R18653 gnd.n4575 gnd.n2096 9.3005
R18654 gnd.n4572 gnd.n2097 9.3005
R18655 gnd.n4571 gnd.n2098 9.3005
R18656 gnd.n4568 gnd.n2099 9.3005
R18657 gnd.n4567 gnd.n2100 9.3005
R18658 gnd.n4564 gnd.n2101 9.3005
R18659 gnd.n4563 gnd.n2102 9.3005
R18660 gnd.n4560 gnd.n4559 9.3005
R18661 gnd.n4558 gnd.n2104 9.3005
R18662 gnd.n4600 gnd.n2082 9.3005
R18663 gnd.n4094 gnd.n4020 9.3005
R18664 gnd.n4093 gnd.n4022 9.3005
R18665 gnd.n4092 gnd.n4023 9.3005
R18666 gnd.n4090 gnd.n4024 9.3005
R18667 gnd.n4089 gnd.n4025 9.3005
R18668 gnd.n4087 gnd.n4026 9.3005
R18669 gnd.n4086 gnd.n4027 9.3005
R18670 gnd.n4084 gnd.n4028 9.3005
R18671 gnd.n4083 gnd.n4029 9.3005
R18672 gnd.n4081 gnd.n4030 9.3005
R18673 gnd.n4080 gnd.n4031 9.3005
R18674 gnd.n4078 gnd.n4032 9.3005
R18675 gnd.n4077 gnd.n4033 9.3005
R18676 gnd.n4075 gnd.n4034 9.3005
R18677 gnd.n4074 gnd.n4035 9.3005
R18678 gnd.n4072 gnd.n4036 9.3005
R18679 gnd.n4071 gnd.n4037 9.3005
R18680 gnd.n4069 gnd.n4038 9.3005
R18681 gnd.n4068 gnd.n4039 9.3005
R18682 gnd.n4066 gnd.n4040 9.3005
R18683 gnd.n4065 gnd.n4041 9.3005
R18684 gnd.n4063 gnd.n4042 9.3005
R18685 gnd.n4062 gnd.n4043 9.3005
R18686 gnd.n4060 gnd.n4044 9.3005
R18687 gnd.n4059 gnd.n4045 9.3005
R18688 gnd.n4057 gnd.n4046 9.3005
R18689 gnd.n4056 gnd.n4047 9.3005
R18690 gnd.n4054 gnd.n4048 9.3005
R18691 gnd.n4053 gnd.n4049 9.3005
R18692 gnd.n4051 gnd.n4050 9.3005
R18693 gnd.n2186 gnd.n2184 9.3005
R18694 gnd.n4312 gnd.n4311 9.3005
R18695 gnd.n2191 gnd.n2185 9.3005
R18696 gnd.n2190 gnd.n2187 9.3005
R18697 gnd.n2189 gnd.n2188 9.3005
R18698 gnd.n2168 gnd.n2167 9.3005
R18699 gnd.n4339 gnd.n4338 9.3005
R18700 gnd.n4340 gnd.n2166 9.3005
R18701 gnd.n4342 gnd.n4341 9.3005
R18702 gnd.n2162 gnd.n2161 9.3005
R18703 gnd.n4365 gnd.n4364 9.3005
R18704 gnd.n4366 gnd.n2160 9.3005
R18705 gnd.n4368 gnd.n4367 9.3005
R18706 gnd.n4369 gnd.n2159 9.3005
R18707 gnd.n4373 gnd.n4372 9.3005
R18708 gnd.n4374 gnd.n2158 9.3005
R18709 gnd.n4376 gnd.n4375 9.3005
R18710 gnd.n2141 gnd.n2140 9.3005
R18711 gnd.n4414 gnd.n4413 9.3005
R18712 gnd.n4415 gnd.n2139 9.3005
R18713 gnd.n4417 gnd.n4416 9.3005
R18714 gnd.n4418 gnd.n2138 9.3005
R18715 gnd.n4422 gnd.n4421 9.3005
R18716 gnd.n4423 gnd.n2137 9.3005
R18717 gnd.n4429 gnd.n4424 9.3005
R18718 gnd.n4428 gnd.n4425 9.3005
R18719 gnd.n4427 gnd.n4426 9.3005
R18720 gnd.n2116 gnd.n2115 9.3005
R18721 gnd.n4507 gnd.n4506 9.3005
R18722 gnd.n4508 gnd.n2114 9.3005
R18723 gnd.n4511 gnd.n4510 9.3005
R18724 gnd.n4509 gnd.n2108 9.3005
R18725 gnd.n4555 gnd.n2107 9.3005
R18726 gnd.n4557 gnd.n4556 9.3005
R18727 gnd.n4096 gnd.n4095 9.3005
R18728 gnd.n4104 gnd.n4103 9.3005
R18729 gnd.n4105 gnd.n4014 9.3005
R18730 gnd.n4106 gnd.n4013 9.3005
R18731 gnd.n4012 gnd.n4010 9.3005
R18732 gnd.n4112 gnd.n4009 9.3005
R18733 gnd.n4113 gnd.n4008 9.3005
R18734 gnd.n4114 gnd.n4007 9.3005
R18735 gnd.n4006 gnd.n4004 9.3005
R18736 gnd.n4120 gnd.n4003 9.3005
R18737 gnd.n4121 gnd.n4002 9.3005
R18738 gnd.n4122 gnd.n4001 9.3005
R18739 gnd.n4000 gnd.n3998 9.3005
R18740 gnd.n4128 gnd.n3997 9.3005
R18741 gnd.n4129 gnd.n3996 9.3005
R18742 gnd.n4130 gnd.n3995 9.3005
R18743 gnd.n3994 gnd.n3992 9.3005
R18744 gnd.n4136 gnd.n3991 9.3005
R18745 gnd.n4137 gnd.n3990 9.3005
R18746 gnd.n4138 gnd.n3989 9.3005
R18747 gnd.n3988 gnd.n3983 9.3005
R18748 gnd.n4144 gnd.n3982 9.3005
R18749 gnd.n4145 gnd.n3981 9.3005
R18750 gnd.n4146 gnd.n3980 9.3005
R18751 gnd.n3979 gnd.n3977 9.3005
R18752 gnd.n4152 gnd.n3976 9.3005
R18753 gnd.n4153 gnd.n3975 9.3005
R18754 gnd.n4154 gnd.n3974 9.3005
R18755 gnd.n3973 gnd.n3971 9.3005
R18756 gnd.n4160 gnd.n3970 9.3005
R18757 gnd.n4161 gnd.n3969 9.3005
R18758 gnd.n4162 gnd.n3968 9.3005
R18759 gnd.n3967 gnd.n3965 9.3005
R18760 gnd.n4167 gnd.n3964 9.3005
R18761 gnd.n4168 gnd.n3963 9.3005
R18762 gnd.n3962 gnd.n3960 9.3005
R18763 gnd.n4173 gnd.n3959 9.3005
R18764 gnd.n4175 gnd.n4174 9.3005
R18765 gnd.n4102 gnd.n4019 9.3005
R18766 gnd.n4101 gnd.n4100 9.3005
R18767 gnd.n2311 gnd.n2310 9.3005
R18768 gnd.n4190 gnd.n4189 9.3005
R18769 gnd.n4191 gnd.n2309 9.3005
R18770 gnd.n4193 gnd.n4192 9.3005
R18771 gnd.n2295 gnd.n2294 9.3005
R18772 gnd.n4206 gnd.n4205 9.3005
R18773 gnd.n4207 gnd.n2293 9.3005
R18774 gnd.n4209 gnd.n4208 9.3005
R18775 gnd.n2279 gnd.n2278 9.3005
R18776 gnd.n4222 gnd.n4221 9.3005
R18777 gnd.n4223 gnd.n2277 9.3005
R18778 gnd.n4225 gnd.n4224 9.3005
R18779 gnd.n2263 gnd.n2262 9.3005
R18780 gnd.n4238 gnd.n4237 9.3005
R18781 gnd.n4239 gnd.n2261 9.3005
R18782 gnd.n4241 gnd.n4240 9.3005
R18783 gnd.n2247 gnd.n2246 9.3005
R18784 gnd.n4254 gnd.n4253 9.3005
R18785 gnd.n4255 gnd.n2245 9.3005
R18786 gnd.n4257 gnd.n4256 9.3005
R18787 gnd.n2231 gnd.n2230 9.3005
R18788 gnd.n4270 gnd.n4269 9.3005
R18789 gnd.n4271 gnd.n2229 9.3005
R18790 gnd.n4274 gnd.n4273 9.3005
R18791 gnd.n4272 gnd.n2214 9.3005
R18792 gnd.n4286 gnd.n2215 9.3005
R18793 gnd.n6337 gnd.n978 9.3005
R18794 gnd.n6336 gnd.n979 9.3005
R18795 gnd.n6335 gnd.n980 9.3005
R18796 gnd.n999 gnd.n981 9.3005
R18797 gnd.n6325 gnd.n1000 9.3005
R18798 gnd.n6324 gnd.n1001 9.3005
R18799 gnd.n6323 gnd.n1002 9.3005
R18800 gnd.n1020 gnd.n1003 9.3005
R18801 gnd.n6313 gnd.n1021 9.3005
R18802 gnd.n6312 gnd.n1022 9.3005
R18803 gnd.n6311 gnd.n1023 9.3005
R18804 gnd.n1041 gnd.n1024 9.3005
R18805 gnd.n6301 gnd.n1042 9.3005
R18806 gnd.n6300 gnd.n1043 9.3005
R18807 gnd.n6299 gnd.n1044 9.3005
R18808 gnd.n1062 gnd.n1045 9.3005
R18809 gnd.n6289 gnd.n1063 9.3005
R18810 gnd.n6288 gnd.n1064 9.3005
R18811 gnd.n6287 gnd.n1065 9.3005
R18812 gnd.n1083 gnd.n1066 9.3005
R18813 gnd.n6277 gnd.n1084 9.3005
R18814 gnd.n6276 gnd.n1085 9.3005
R18815 gnd.n6275 gnd.n1086 9.3005
R18816 gnd.n1104 gnd.n1087 9.3005
R18817 gnd.n6265 gnd.n1105 9.3005
R18818 gnd.n6264 gnd.n1106 9.3005
R18819 gnd.n6263 gnd.n1107 9.3005
R18820 gnd.n4177 gnd.n4176 9.3005
R18821 gnd.n977 gnd.n966 9.3005
R18822 gnd.n6347 gnd.n965 9.3005
R18823 gnd.n964 gnd.n960 9.3005
R18824 gnd.n6353 gnd.n959 9.3005
R18825 gnd.n6354 gnd.n958 9.3005
R18826 gnd.n6355 gnd.n957 9.3005
R18827 gnd.n956 gnd.n952 9.3005
R18828 gnd.n6361 gnd.n951 9.3005
R18829 gnd.n6362 gnd.n950 9.3005
R18830 gnd.n6363 gnd.n949 9.3005
R18831 gnd.n948 gnd.n944 9.3005
R18832 gnd.n6369 gnd.n943 9.3005
R18833 gnd.n6370 gnd.n942 9.3005
R18834 gnd.n6371 gnd.n941 9.3005
R18835 gnd.n940 gnd.n936 9.3005
R18836 gnd.n6377 gnd.n935 9.3005
R18837 gnd.n6378 gnd.n934 9.3005
R18838 gnd.n6379 gnd.n933 9.3005
R18839 gnd.n932 gnd.n928 9.3005
R18840 gnd.n6385 gnd.n927 9.3005
R18841 gnd.n6386 gnd.n926 9.3005
R18842 gnd.n6387 gnd.n925 9.3005
R18843 gnd.n924 gnd.n920 9.3005
R18844 gnd.n6393 gnd.n919 9.3005
R18845 gnd.n6394 gnd.n918 9.3005
R18846 gnd.n6395 gnd.n917 9.3005
R18847 gnd.n916 gnd.n912 9.3005
R18848 gnd.n6401 gnd.n911 9.3005
R18849 gnd.n6402 gnd.n910 9.3005
R18850 gnd.n6403 gnd.n909 9.3005
R18851 gnd.n908 gnd.n904 9.3005
R18852 gnd.n6409 gnd.n903 9.3005
R18853 gnd.n6410 gnd.n902 9.3005
R18854 gnd.n6411 gnd.n901 9.3005
R18855 gnd.n900 gnd.n896 9.3005
R18856 gnd.n6417 gnd.n895 9.3005
R18857 gnd.n6418 gnd.n894 9.3005
R18858 gnd.n6419 gnd.n893 9.3005
R18859 gnd.n892 gnd.n888 9.3005
R18860 gnd.n6425 gnd.n887 9.3005
R18861 gnd.n6426 gnd.n886 9.3005
R18862 gnd.n6427 gnd.n885 9.3005
R18863 gnd.n884 gnd.n880 9.3005
R18864 gnd.n6433 gnd.n879 9.3005
R18865 gnd.n6434 gnd.n878 9.3005
R18866 gnd.n6435 gnd.n877 9.3005
R18867 gnd.n876 gnd.n872 9.3005
R18868 gnd.n6441 gnd.n871 9.3005
R18869 gnd.n6442 gnd.n870 9.3005
R18870 gnd.n6443 gnd.n869 9.3005
R18871 gnd.n868 gnd.n864 9.3005
R18872 gnd.n6449 gnd.n863 9.3005
R18873 gnd.n6450 gnd.n862 9.3005
R18874 gnd.n6451 gnd.n861 9.3005
R18875 gnd.n860 gnd.n856 9.3005
R18876 gnd.n6457 gnd.n855 9.3005
R18877 gnd.n6458 gnd.n854 9.3005
R18878 gnd.n6459 gnd.n853 9.3005
R18879 gnd.n852 gnd.n848 9.3005
R18880 gnd.n6465 gnd.n847 9.3005
R18881 gnd.n6466 gnd.n846 9.3005
R18882 gnd.n6467 gnd.n845 9.3005
R18883 gnd.n844 gnd.n840 9.3005
R18884 gnd.n6473 gnd.n839 9.3005
R18885 gnd.n6474 gnd.n838 9.3005
R18886 gnd.n6475 gnd.n837 9.3005
R18887 gnd.n836 gnd.n832 9.3005
R18888 gnd.n6481 gnd.n831 9.3005
R18889 gnd.n6482 gnd.n830 9.3005
R18890 gnd.n6483 gnd.n829 9.3005
R18891 gnd.n828 gnd.n824 9.3005
R18892 gnd.n6489 gnd.n823 9.3005
R18893 gnd.n6490 gnd.n822 9.3005
R18894 gnd.n6491 gnd.n821 9.3005
R18895 gnd.n820 gnd.n816 9.3005
R18896 gnd.n6497 gnd.n815 9.3005
R18897 gnd.n6498 gnd.n814 9.3005
R18898 gnd.n6499 gnd.n813 9.3005
R18899 gnd.n812 gnd.n808 9.3005
R18900 gnd.n6505 gnd.n807 9.3005
R18901 gnd.n6506 gnd.n806 9.3005
R18902 gnd.n6507 gnd.n805 9.3005
R18903 gnd.n804 gnd.n800 9.3005
R18904 gnd.n6513 gnd.n799 9.3005
R18905 gnd.n6515 gnd.n6514 9.3005
R18906 gnd.n6346 gnd.n6345 9.3005
R18907 gnd.n1530 gnd.n1529 9.3005
R18908 gnd.n1516 gnd.n1512 9.3005
R18909 gnd.n1537 gnd.n1536 9.3005
R18910 gnd.n1538 gnd.n1507 9.3005
R18911 gnd.n1549 gnd.n1548 9.3005
R18912 gnd.n1509 gnd.n1505 9.3005
R18913 gnd.n1556 gnd.n1555 9.3005
R18914 gnd.n1557 gnd.n1500 9.3005
R18915 gnd.n1568 gnd.n1567 9.3005
R18916 gnd.n1502 gnd.n1498 9.3005
R18917 gnd.n1575 gnd.n1574 9.3005
R18918 gnd.n1495 gnd.n1494 9.3005
R18919 gnd.n1584 gnd.n1583 9.3005
R18920 gnd.n1492 gnd.n1491 9.3005
R18921 gnd.n1591 gnd.n1590 9.3005
R18922 gnd.n1483 gnd.n1482 9.3005
R18923 gnd.n1598 gnd.n1597 9.3005
R18924 gnd.n1480 gnd.n1478 9.3005
R18925 gnd.n1519 gnd.n1514 9.3005
R18926 gnd.n1593 gnd.n1592 9.3005
R18927 gnd.n1582 gnd.n1488 9.3005
R18928 gnd.n1581 gnd.n1580 9.3005
R18929 gnd.n1577 gnd.n1576 9.3005
R18930 gnd.n1497 gnd.n1496 9.3005
R18931 gnd.n1566 gnd.n1565 9.3005
R18932 gnd.n1562 gnd.n1501 9.3005
R18933 gnd.n1559 gnd.n1558 9.3005
R18934 gnd.n1504 gnd.n1503 9.3005
R18935 gnd.n1547 gnd.n1546 9.3005
R18936 gnd.n1543 gnd.n1508 9.3005
R18937 gnd.n1540 gnd.n1539 9.3005
R18938 gnd.n1511 gnd.n1510 9.3005
R18939 gnd.n1528 gnd.n1527 9.3005
R18940 gnd.n1524 gnd.n1515 9.3005
R18941 gnd.n1521 gnd.n1520 9.3005
R18942 gnd.n1594 gnd.n1484 9.3005
R18943 gnd.n1596 gnd.n1595 9.3005
R18944 gnd.n5838 gnd.n5837 9.3005
R18945 gnd.n5836 gnd.n1479 9.3005
R18946 gnd.n5835 gnd.n5834 9.3005
R18947 gnd.n5833 gnd.n1606 9.3005
R18948 gnd.n5832 gnd.n5831 9.3005
R18949 gnd.n5830 gnd.n1607 9.3005
R18950 gnd.n5826 gnd.n5825 9.3005
R18951 gnd.n5824 gnd.n1614 9.3005
R18952 gnd.n5823 gnd.n5822 9.3005
R18953 gnd.n5821 gnd.n5816 9.3005
R18954 gnd.n5411 gnd.n5410 9.3005
R18955 gnd.n1943 gnd.n1942 9.3005
R18956 gnd.n5424 gnd.n5423 9.3005
R18957 gnd.n5425 gnd.n1941 9.3005
R18958 gnd.n5427 gnd.n5426 9.3005
R18959 gnd.n1930 gnd.n1929 9.3005
R18960 gnd.n5440 gnd.n5439 9.3005
R18961 gnd.n5441 gnd.n1928 9.3005
R18962 gnd.n5443 gnd.n5442 9.3005
R18963 gnd.n1917 gnd.n1916 9.3005
R18964 gnd.n5456 gnd.n5455 9.3005
R18965 gnd.n5457 gnd.n1915 9.3005
R18966 gnd.n5459 gnd.n5458 9.3005
R18967 gnd.n1904 gnd.n1903 9.3005
R18968 gnd.n5472 gnd.n5471 9.3005
R18969 gnd.n5473 gnd.n1902 9.3005
R18970 gnd.n5475 gnd.n5474 9.3005
R18971 gnd.n1890 gnd.n1889 9.3005
R18972 gnd.n5488 gnd.n5487 9.3005
R18973 gnd.n5489 gnd.n1888 9.3005
R18974 gnd.n5491 gnd.n5490 9.3005
R18975 gnd.n1878 gnd.n1877 9.3005
R18976 gnd.n5504 gnd.n5503 9.3005
R18977 gnd.n5505 gnd.n1876 9.3005
R18978 gnd.n5507 gnd.n5506 9.3005
R18979 gnd.n1864 gnd.n1863 9.3005
R18980 gnd.n5520 gnd.n5519 9.3005
R18981 gnd.n5521 gnd.n1862 9.3005
R18982 gnd.n5523 gnd.n5522 9.3005
R18983 gnd.n1850 gnd.n1849 9.3005
R18984 gnd.n5536 gnd.n5535 9.3005
R18985 gnd.n5537 gnd.n1848 9.3005
R18986 gnd.n5539 gnd.n5538 9.3005
R18987 gnd.n1837 gnd.n1836 9.3005
R18988 gnd.n5552 gnd.n5551 9.3005
R18989 gnd.n5553 gnd.n1835 9.3005
R18990 gnd.n5555 gnd.n5554 9.3005
R18991 gnd.n1824 gnd.n1823 9.3005
R18992 gnd.n5568 gnd.n5567 9.3005
R18993 gnd.n5569 gnd.n1822 9.3005
R18994 gnd.n5571 gnd.n5570 9.3005
R18995 gnd.n1808 gnd.n1807 9.3005
R18996 gnd.n5584 gnd.n5583 9.3005
R18997 gnd.n5585 gnd.n1806 9.3005
R18998 gnd.n5587 gnd.n5586 9.3005
R18999 gnd.n1794 gnd.n1793 9.3005
R19000 gnd.n5600 gnd.n5599 9.3005
R19001 gnd.n5601 gnd.n1792 9.3005
R19002 gnd.n5603 gnd.n5602 9.3005
R19003 gnd.n1780 gnd.n1779 9.3005
R19004 gnd.n5616 gnd.n5615 9.3005
R19005 gnd.n5617 gnd.n1778 9.3005
R19006 gnd.n5619 gnd.n5618 9.3005
R19007 gnd.n1766 gnd.n1765 9.3005
R19008 gnd.n5632 gnd.n5631 9.3005
R19009 gnd.n5633 gnd.n1764 9.3005
R19010 gnd.n5635 gnd.n5634 9.3005
R19011 gnd.n1752 gnd.n1751 9.3005
R19012 gnd.n5648 gnd.n5647 9.3005
R19013 gnd.n5649 gnd.n1750 9.3005
R19014 gnd.n5651 gnd.n5650 9.3005
R19015 gnd.n1738 gnd.n1737 9.3005
R19016 gnd.n5664 gnd.n5663 9.3005
R19017 gnd.n5665 gnd.n1736 9.3005
R19018 gnd.n5667 gnd.n5666 9.3005
R19019 gnd.n1724 gnd.n1723 9.3005
R19020 gnd.n5680 gnd.n5679 9.3005
R19021 gnd.n5681 gnd.n1722 9.3005
R19022 gnd.n5683 gnd.n5682 9.3005
R19023 gnd.n1711 gnd.n1710 9.3005
R19024 gnd.n5696 gnd.n5695 9.3005
R19025 gnd.n5697 gnd.n1709 9.3005
R19026 gnd.n5699 gnd.n5698 9.3005
R19027 gnd.n1696 gnd.n1695 9.3005
R19028 gnd.n5712 gnd.n5711 9.3005
R19029 gnd.n5713 gnd.n1694 9.3005
R19030 gnd.n5715 gnd.n5714 9.3005
R19031 gnd.n1682 gnd.n1681 9.3005
R19032 gnd.n5728 gnd.n5727 9.3005
R19033 gnd.n5729 gnd.n1680 9.3005
R19034 gnd.n5731 gnd.n5730 9.3005
R19035 gnd.n1670 gnd.n1669 9.3005
R19036 gnd.n5744 gnd.n5743 9.3005
R19037 gnd.n5745 gnd.n1668 9.3005
R19038 gnd.n5747 gnd.n5746 9.3005
R19039 gnd.n1657 gnd.n1656 9.3005
R19040 gnd.n5760 gnd.n5759 9.3005
R19041 gnd.n5761 gnd.n1655 9.3005
R19042 gnd.n5763 gnd.n5762 9.3005
R19043 gnd.n1644 gnd.n1643 9.3005
R19044 gnd.n5776 gnd.n5775 9.3005
R19045 gnd.n5777 gnd.n1642 9.3005
R19046 gnd.n5779 gnd.n5778 9.3005
R19047 gnd.n1631 gnd.n1630 9.3005
R19048 gnd.n5792 gnd.n5791 9.3005
R19049 gnd.n5793 gnd.n1628 9.3005
R19050 gnd.n5797 gnd.n5796 9.3005
R19051 gnd.n5795 gnd.n1629 9.3005
R19052 gnd.n5794 gnd.n1616 9.3005
R19053 gnd.n5813 gnd.n1615 9.3005
R19054 gnd.n5815 gnd.n5814 9.3005
R19055 gnd.n5409 gnd.n1954 9.3005
R19056 gnd.n1956 gnd.n1955 9.3005
R19057 gnd.n4534 gnd.n4531 9.3005
R19058 gnd.n4536 gnd.n4535 9.3005
R19059 gnd.n4538 gnd.n4537 9.3005
R19060 gnd.n4539 gnd.n4524 9.3005
R19061 gnd.n4541 gnd.n4540 9.3005
R19062 gnd.n4542 gnd.n4523 9.3005
R19063 gnd.n4544 gnd.n4543 9.3005
R19064 gnd.n4545 gnd.n4518 9.3005
R19065 gnd.n5408 gnd.n5407 9.3005
R19066 gnd.n3907 gnd.n3896 9.3005
R19067 gnd.n3906 gnd.n3905 9.3005
R19068 gnd.n3904 gnd.n3897 9.3005
R19069 gnd.n3903 gnd.n3902 9.3005
R19070 gnd.n3901 gnd.n3900 9.3005
R19071 gnd.n2165 gnd.n2164 9.3005
R19072 gnd.n4347 gnd.n4346 9.3005
R19073 gnd.n4348 gnd.n2163 9.3005
R19074 gnd.n4350 gnd.n4349 9.3005
R19075 gnd.n2155 gnd.n2153 9.3005
R19076 gnd.n4391 gnd.n4390 9.3005
R19077 gnd.n4389 gnd.n2154 9.3005
R19078 gnd.n4388 gnd.n4387 9.3005
R19079 gnd.n4386 gnd.n2156 9.3005
R19080 gnd.n4385 gnd.n4384 9.3005
R19081 gnd.n4383 gnd.n4380 9.3005
R19082 gnd.n4382 gnd.n4381 9.3005
R19083 gnd.n2134 gnd.n2132 9.3005
R19084 gnd.n4440 gnd.n4439 9.3005
R19085 gnd.n4438 gnd.n2133 9.3005
R19086 gnd.n4437 gnd.n4436 9.3005
R19087 gnd.n4435 gnd.n2135 9.3005
R19088 gnd.n4434 gnd.n4433 9.3005
R19089 gnd.n2119 gnd.n2118 9.3005
R19090 gnd.n4499 gnd.n4498 9.3005
R19091 gnd.n4500 gnd.n2117 9.3005
R19092 gnd.n4502 gnd.n4501 9.3005
R19093 gnd.n2113 gnd.n2112 9.3005
R19094 gnd.n4516 gnd.n4515 9.3005
R19095 gnd.n4517 gnd.n2110 9.3005
R19096 gnd.n4551 gnd.n4550 9.3005
R19097 gnd.n4549 gnd.n2111 9.3005
R19098 gnd.n4547 gnd.n4546 9.3005
R19099 gnd.n2025 gnd.n2024 9.3005
R19100 gnd.n5360 gnd.n5359 9.3005
R19101 gnd.n5362 gnd.n5361 9.3005
R19102 gnd.n2013 gnd.n2012 9.3005
R19103 gnd.n5368 gnd.n5367 9.3005
R19104 gnd.n5370 gnd.n5369 9.3005
R19105 gnd.n2005 gnd.n2004 9.3005
R19106 gnd.n5376 gnd.n5375 9.3005
R19107 gnd.n5378 gnd.n5377 9.3005
R19108 gnd.n1995 gnd.n1994 9.3005
R19109 gnd.n5384 gnd.n5383 9.3005
R19110 gnd.n5386 gnd.n5385 9.3005
R19111 gnd.n1987 gnd.n1986 9.3005
R19112 gnd.n5392 gnd.n5391 9.3005
R19113 gnd.n5394 gnd.n5393 9.3005
R19114 gnd.n1977 gnd.n1975 9.3005
R19115 gnd.n5400 gnd.n5399 9.3005
R19116 gnd.n5401 gnd.n1974 9.3005
R19117 gnd.n2028 gnd.n1116 9.3005
R19118 gnd.n1978 gnd.n1976 9.3005
R19119 gnd.n5398 gnd.n5397 9.3005
R19120 gnd.n5396 gnd.n5395 9.3005
R19121 gnd.n1982 gnd.n1981 9.3005
R19122 gnd.n5390 gnd.n5389 9.3005
R19123 gnd.n5388 gnd.n5387 9.3005
R19124 gnd.n1991 gnd.n1990 9.3005
R19125 gnd.n5382 gnd.n5381 9.3005
R19126 gnd.n5380 gnd.n5379 9.3005
R19127 gnd.n1999 gnd.n1998 9.3005
R19128 gnd.n5374 gnd.n5373 9.3005
R19129 gnd.n5372 gnd.n5371 9.3005
R19130 gnd.n2009 gnd.n2008 9.3005
R19131 gnd.n5366 gnd.n5365 9.3005
R19132 gnd.n5364 gnd.n5363 9.3005
R19133 gnd.n2019 gnd.n2018 9.3005
R19134 gnd.n5358 gnd.n5357 9.3005
R19135 gnd.n6253 gnd.n1117 9.3005
R19136 gnd.n6252 gnd.n6251 9.3005
R19137 gnd.n6250 gnd.n1121 9.3005
R19138 gnd.n6249 gnd.n6248 9.3005
R19139 gnd.n6247 gnd.n1122 9.3005
R19140 gnd.n6246 gnd.n6245 9.3005
R19141 gnd.n6244 gnd.n1126 9.3005
R19142 gnd.n6243 gnd.n6242 9.3005
R19143 gnd.n6241 gnd.n1127 9.3005
R19144 gnd.n6240 gnd.n6239 9.3005
R19145 gnd.n6238 gnd.n1131 9.3005
R19146 gnd.n6237 gnd.n6236 9.3005
R19147 gnd.n6235 gnd.n1132 9.3005
R19148 gnd.n6234 gnd.n6233 9.3005
R19149 gnd.n6232 gnd.n1136 9.3005
R19150 gnd.n6231 gnd.n6230 9.3005
R19151 gnd.n6229 gnd.n1137 9.3005
R19152 gnd.n6228 gnd.n6227 9.3005
R19153 gnd.n6226 gnd.n1141 9.3005
R19154 gnd.n6225 gnd.n6224 9.3005
R19155 gnd.n6223 gnd.n1142 9.3005
R19156 gnd.n6222 gnd.n6221 9.3005
R19157 gnd.n6220 gnd.n1146 9.3005
R19158 gnd.n6219 gnd.n6218 9.3005
R19159 gnd.n6217 gnd.n1147 9.3005
R19160 gnd.n6216 gnd.n6215 9.3005
R19161 gnd.n6214 gnd.n1151 9.3005
R19162 gnd.n6213 gnd.n6212 9.3005
R19163 gnd.n6211 gnd.n1152 9.3005
R19164 gnd.n6210 gnd.n6209 9.3005
R19165 gnd.n6208 gnd.n1156 9.3005
R19166 gnd.n6207 gnd.n6206 9.3005
R19167 gnd.n6205 gnd.n1157 9.3005
R19168 gnd.n6204 gnd.n6203 9.3005
R19169 gnd.n6202 gnd.n1161 9.3005
R19170 gnd.n6201 gnd.n6200 9.3005
R19171 gnd.n6199 gnd.n1162 9.3005
R19172 gnd.n6198 gnd.n6197 9.3005
R19173 gnd.n6196 gnd.n1166 9.3005
R19174 gnd.n6195 gnd.n6194 9.3005
R19175 gnd.n6193 gnd.n1167 9.3005
R19176 gnd.n6192 gnd.n6191 9.3005
R19177 gnd.n6190 gnd.n1171 9.3005
R19178 gnd.n6189 gnd.n6188 9.3005
R19179 gnd.n6187 gnd.n1172 9.3005
R19180 gnd.n6186 gnd.n6185 9.3005
R19181 gnd.n6184 gnd.n1176 9.3005
R19182 gnd.n6183 gnd.n6182 9.3005
R19183 gnd.n6181 gnd.n1177 9.3005
R19184 gnd.n6180 gnd.n6179 9.3005
R19185 gnd.n6178 gnd.n1181 9.3005
R19186 gnd.n6177 gnd.n6176 9.3005
R19187 gnd.n6175 gnd.n1182 9.3005
R19188 gnd.n6174 gnd.n6173 9.3005
R19189 gnd.n6172 gnd.n1186 9.3005
R19190 gnd.n6171 gnd.n6170 9.3005
R19191 gnd.n6169 gnd.n1187 9.3005
R19192 gnd.n6168 gnd.n6167 9.3005
R19193 gnd.n6166 gnd.n1191 9.3005
R19194 gnd.n6165 gnd.n6164 9.3005
R19195 gnd.n6163 gnd.n1192 9.3005
R19196 gnd.n6162 gnd.n6161 9.3005
R19197 gnd.n6160 gnd.n1196 9.3005
R19198 gnd.n6159 gnd.n6158 9.3005
R19199 gnd.n6157 gnd.n1197 9.3005
R19200 gnd.n6156 gnd.n6155 9.3005
R19201 gnd.n6154 gnd.n1201 9.3005
R19202 gnd.n6153 gnd.n6152 9.3005
R19203 gnd.n6151 gnd.n1202 9.3005
R19204 gnd.n6150 gnd.n6149 9.3005
R19205 gnd.n6148 gnd.n1206 9.3005
R19206 gnd.n6147 gnd.n6146 9.3005
R19207 gnd.n6145 gnd.n1207 9.3005
R19208 gnd.n6144 gnd.n6143 9.3005
R19209 gnd.n6142 gnd.n1211 9.3005
R19210 gnd.n6141 gnd.n6140 9.3005
R19211 gnd.n6139 gnd.n1212 9.3005
R19212 gnd.n6138 gnd.n6137 9.3005
R19213 gnd.n6136 gnd.n1216 9.3005
R19214 gnd.n6135 gnd.n6134 9.3005
R19215 gnd.n6133 gnd.n1217 9.3005
R19216 gnd.n6132 gnd.n6131 9.3005
R19217 gnd.n6130 gnd.n1221 9.3005
R19218 gnd.n6129 gnd.n6128 9.3005
R19219 gnd.n6127 gnd.n1222 9.3005
R19220 gnd.n6126 gnd.n6125 9.3005
R19221 gnd.n6124 gnd.n1226 9.3005
R19222 gnd.n6123 gnd.n6122 9.3005
R19223 gnd.n6121 gnd.n1227 9.3005
R19224 gnd.n6120 gnd.n6119 9.3005
R19225 gnd.n6118 gnd.n1231 9.3005
R19226 gnd.n6117 gnd.n6116 9.3005
R19227 gnd.n6115 gnd.n1232 9.3005
R19228 gnd.n6114 gnd.n6113 9.3005
R19229 gnd.n6112 gnd.n1236 9.3005
R19230 gnd.n6111 gnd.n6110 9.3005
R19231 gnd.n6109 gnd.n1237 9.3005
R19232 gnd.n6108 gnd.n6107 9.3005
R19233 gnd.n6106 gnd.n1241 9.3005
R19234 gnd.n6105 gnd.n6104 9.3005
R19235 gnd.n6103 gnd.n1242 9.3005
R19236 gnd.n6255 gnd.n6254 9.3005
R19237 gnd.n6012 gnd.n1341 9.3005
R19238 gnd.n6011 gnd.n6010 9.3005
R19239 gnd.n6009 gnd.n1343 9.3005
R19240 gnd.n6008 gnd.n6007 9.3005
R19241 gnd.n6006 gnd.n1347 9.3005
R19242 gnd.n6005 gnd.n6004 9.3005
R19243 gnd.n6003 gnd.n1348 9.3005
R19244 gnd.n6002 gnd.n6001 9.3005
R19245 gnd.n6000 gnd.n1352 9.3005
R19246 gnd.n5999 gnd.n5998 9.3005
R19247 gnd.n5997 gnd.n1353 9.3005
R19248 gnd.n5996 gnd.n5995 9.3005
R19249 gnd.n5994 gnd.n1357 9.3005
R19250 gnd.n5993 gnd.n5992 9.3005
R19251 gnd.n5991 gnd.n1358 9.3005
R19252 gnd.n5990 gnd.n5989 9.3005
R19253 gnd.n407 gnd.n405 9.3005
R19254 gnd.n7170 gnd.n7169 9.3005
R19255 gnd.n7168 gnd.n406 9.3005
R19256 gnd.n7167 gnd.n7166 9.3005
R19257 gnd.n7165 gnd.n408 9.3005
R19258 gnd.n375 gnd.n373 9.3005
R19259 gnd.n7216 gnd.n7215 9.3005
R19260 gnd.n7214 gnd.n374 9.3005
R19261 gnd.n7213 gnd.n7212 9.3005
R19262 gnd.n7211 gnd.n376 9.3005
R19263 gnd.n7210 gnd.n7209 9.3005
R19264 gnd.n320 gnd.n318 9.3005
R19265 gnd.n7347 gnd.n7346 9.3005
R19266 gnd.n7345 gnd.n319 9.3005
R19267 gnd.n7344 gnd.n7343 9.3005
R19268 gnd.n7342 gnd.n321 9.3005
R19269 gnd.n7341 gnd.n7340 9.3005
R19270 gnd.n7339 gnd.n325 9.3005
R19271 gnd.n7338 gnd.n7337 9.3005
R19272 gnd.n7336 gnd.n326 9.3005
R19273 gnd.n297 gnd.n296 9.3005
R19274 gnd.n7361 gnd.n7360 9.3005
R19275 gnd.n7362 gnd.n295 9.3005
R19276 gnd.n7364 gnd.n7363 9.3005
R19277 gnd.n281 gnd.n280 9.3005
R19278 gnd.n7377 gnd.n7376 9.3005
R19279 gnd.n7378 gnd.n279 9.3005
R19280 gnd.n7380 gnd.n7379 9.3005
R19281 gnd.n267 gnd.n266 9.3005
R19282 gnd.n7393 gnd.n7392 9.3005
R19283 gnd.n7394 gnd.n265 9.3005
R19284 gnd.n7396 gnd.n7395 9.3005
R19285 gnd.n251 gnd.n250 9.3005
R19286 gnd.n7409 gnd.n7408 9.3005
R19287 gnd.n7410 gnd.n249 9.3005
R19288 gnd.n7412 gnd.n7411 9.3005
R19289 gnd.n236 gnd.n235 9.3005
R19290 gnd.n7425 gnd.n7424 9.3005
R19291 gnd.n7426 gnd.n234 9.3005
R19292 gnd.n7428 gnd.n7427 9.3005
R19293 gnd.n221 gnd.n220 9.3005
R19294 gnd.n7441 gnd.n7440 9.3005
R19295 gnd.n7442 gnd.n218 9.3005
R19296 gnd.n7512 gnd.n7511 9.3005
R19297 gnd.n7510 gnd.n219 9.3005
R19298 gnd.n7509 gnd.n7508 9.3005
R19299 gnd.n7507 gnd.n7443 9.3005
R19300 gnd.n7506 gnd.n7505 9.3005
R19301 gnd.n6014 gnd.n6013 9.3005
R19302 gnd.n7502 gnd.n7445 9.3005
R19303 gnd.n7501 gnd.n7500 9.3005
R19304 gnd.n7499 gnd.n7450 9.3005
R19305 gnd.n7498 gnd.n7497 9.3005
R19306 gnd.n7496 gnd.n7451 9.3005
R19307 gnd.n7495 gnd.n7494 9.3005
R19308 gnd.n7493 gnd.n7458 9.3005
R19309 gnd.n7492 gnd.n7491 9.3005
R19310 gnd.n7490 gnd.n7459 9.3005
R19311 gnd.n7489 gnd.n7488 9.3005
R19312 gnd.n7487 gnd.n7466 9.3005
R19313 gnd.n7486 gnd.n7485 9.3005
R19314 gnd.n7484 gnd.n7467 9.3005
R19315 gnd.n7483 gnd.n7482 9.3005
R19316 gnd.n7481 gnd.n7474 9.3005
R19317 gnd.n7480 gnd.n7479 9.3005
R19318 gnd.n124 gnd.n121 9.3005
R19319 gnd.n7606 gnd.n7605 9.3005
R19320 gnd.n7504 gnd.n7503 9.3005
R19321 gnd.n5854 gnd.n5853 9.3005
R19322 gnd.n5855 gnd.n1476 9.3005
R19323 gnd.n5858 gnd.n5857 9.3005
R19324 gnd.n5856 gnd.n1477 9.3005
R19325 gnd.n1420 gnd.n1419 9.3005
R19326 gnd.n5885 gnd.n5884 9.3005
R19327 gnd.n5886 gnd.n1417 9.3005
R19328 gnd.n5894 gnd.n5893 9.3005
R19329 gnd.n5892 gnd.n1418 9.3005
R19330 gnd.n5891 gnd.n5890 9.3005
R19331 gnd.n5889 gnd.n5887 9.3005
R19332 gnd.n1384 gnd.n1382 9.3005
R19333 gnd.n5954 gnd.n5953 9.3005
R19334 gnd.n5952 gnd.n1383 9.3005
R19335 gnd.n5951 gnd.n5950 9.3005
R19336 gnd.n5949 gnd.n1385 9.3005
R19337 gnd.n5948 gnd.n5947 9.3005
R19338 gnd.n5946 gnd.n5938 9.3005
R19339 gnd.n5945 gnd.n5944 9.3005
R19340 gnd.n5943 gnd.n5940 9.3005
R19341 gnd.n5939 gnd.n382 9.3005
R19342 gnd.n7198 gnd.n381 9.3005
R19343 gnd.n7200 gnd.n7199 9.3005
R19344 gnd.n7201 gnd.n379 9.3005
R19345 gnd.n7204 gnd.n7203 9.3005
R19346 gnd.n7202 gnd.n380 9.3005
R19347 gnd.n348 gnd.n347 9.3005
R19348 gnd.n7245 gnd.n7244 9.3005
R19349 gnd.n7246 gnd.n346 9.3005
R19350 gnd.n7248 gnd.n7247 9.3005
R19351 gnd.n7249 gnd.n79 9.3005
R19352 gnd.n7655 gnd.n80 9.3005
R19353 gnd.n7654 gnd.n7653 9.3005
R19354 gnd.n7652 gnd.n81 9.3005
R19355 gnd.n7651 gnd.n7650 9.3005
R19356 gnd.n7649 gnd.n85 9.3005
R19357 gnd.n7648 gnd.n7647 9.3005
R19358 gnd.n7646 gnd.n86 9.3005
R19359 gnd.n7645 gnd.n7644 9.3005
R19360 gnd.n7643 gnd.n90 9.3005
R19361 gnd.n7642 gnd.n7641 9.3005
R19362 gnd.n7640 gnd.n91 9.3005
R19363 gnd.n7639 gnd.n7638 9.3005
R19364 gnd.n7637 gnd.n95 9.3005
R19365 gnd.n7636 gnd.n7635 9.3005
R19366 gnd.n7634 gnd.n96 9.3005
R19367 gnd.n7633 gnd.n7632 9.3005
R19368 gnd.n7631 gnd.n100 9.3005
R19369 gnd.n7630 gnd.n7629 9.3005
R19370 gnd.n7628 gnd.n101 9.3005
R19371 gnd.n7627 gnd.n7626 9.3005
R19372 gnd.n7625 gnd.n105 9.3005
R19373 gnd.n7624 gnd.n7623 9.3005
R19374 gnd.n7622 gnd.n106 9.3005
R19375 gnd.n7621 gnd.n7620 9.3005
R19376 gnd.n7619 gnd.n110 9.3005
R19377 gnd.n7618 gnd.n7617 9.3005
R19378 gnd.n7616 gnd.n111 9.3005
R19379 gnd.n7615 gnd.n7614 9.3005
R19380 gnd.n7613 gnd.n115 9.3005
R19381 gnd.n7612 gnd.n7611 9.3005
R19382 gnd.n7610 gnd.n116 9.3005
R19383 gnd.n7609 gnd.n7608 9.3005
R19384 gnd.n7607 gnd.n120 9.3005
R19385 gnd.n5841 gnd.n5840 9.3005
R19386 gnd.t211 gnd.n2509 9.24152
R19387 gnd.n2411 gnd.t288 9.24152
R19388 gnd.n3691 gnd.t271 9.24152
R19389 gnd.t81 gnd.n2256 9.24152
R19390 gnd.n2178 gnd.n2177 9.24152
R19391 gnd.t156 gnd.n1860 9.24152
R19392 gnd.n5094 gnd.t203 9.24152
R19393 gnd.n7349 gnd.n312 9.24152
R19394 gnd.n263 gnd.t50 9.24152
R19395 gnd.t58 gnd.t211 8.92286
R19396 gnd.t189 gnd.n4776 8.92286
R19397 gnd.n1820 gnd.t2 8.92286
R19398 gnd.n5141 gnd.t96 8.92286
R19399 gnd.n5653 gnd.t127 8.92286
R19400 gnd.n3661 gnd.n3636 8.92171
R19401 gnd.n3629 gnd.n3604 8.92171
R19402 gnd.n3597 gnd.n3572 8.92171
R19403 gnd.n3566 gnd.n3541 8.92171
R19404 gnd.n3534 gnd.n3509 8.92171
R19405 gnd.n3502 gnd.n3477 8.92171
R19406 gnd.n3470 gnd.n3445 8.92171
R19407 gnd.n3439 gnd.n3414 8.92171
R19408 gnd.n4942 gnd.n4924 8.72777
R19409 gnd.n3165 gnd.t214 8.60421
R19410 gnd.t3 gnd.n2288 8.60421
R19411 gnd.n4806 gnd.t234 8.60421
R19412 gnd.n4819 gnd.t93 8.60421
R19413 gnd.n232 gnd.t73 8.60421
R19414 gnd.n2589 gnd.n2569 8.43467
R19415 gnd.n58 gnd.n38 8.43467
R19416 gnd.n3908 gnd.n0 8.41456
R19417 gnd.n7656 gnd.n7655 8.41456
R19418 gnd.n5525 gnd.n1859 8.28555
R19419 gnd.n5214 gnd.n4763 8.28555
R19420 gnd.n5193 gnd.n5192 8.28555
R19421 gnd.n5629 gnd.n1770 8.28555
R19422 gnd.n5661 gnd.n1740 8.28555
R19423 gnd.n5093 gnd.n5092 8.28555
R19424 gnd.n3662 gnd.n3634 8.14595
R19425 gnd.n3630 gnd.n3602 8.14595
R19426 gnd.n3598 gnd.n3570 8.14595
R19427 gnd.n3567 gnd.n3539 8.14595
R19428 gnd.n3535 gnd.n3507 8.14595
R19429 gnd.n3503 gnd.n3475 8.14595
R19430 gnd.n3471 gnd.n3443 8.14595
R19431 gnd.n3440 gnd.n3412 8.14595
R19432 gnd.n3667 gnd.n3666 7.97301
R19433 gnd.t215 gnd.n2680 7.9669
R19434 gnd.n5404 gnd.n1958 7.9669
R19435 gnd.t298 gnd.t354 7.9669
R19436 gnd.n1256 gnd.n1248 7.9669
R19437 gnd.n7605 gnd.n124 7.75808
R19438 gnd.n1595 gnd.n1594 7.75808
R19439 gnd.n5357 gnd.n2018 7.75808
R19440 gnd.n3861 gnd.n3800 7.75808
R19441 gnd.n6340 gnd.n970 7.64824
R19442 gnd.n6339 gnd.n973 7.64824
R19443 gnd.n4344 gnd.n983 7.64824
R19444 gnd.n6333 gnd.n986 7.64824
R19445 gnd.n4362 gnd.n4361 7.64824
R19446 gnd.n6327 gnd.n997 7.64824
R19447 gnd.n4394 gnd.n4393 7.64824
R19448 gnd.n6321 gnd.n1007 7.64824
R19449 gnd.n4370 gnd.n1015 7.64824
R19450 gnd.n6315 gnd.n1018 7.64824
R19451 gnd.n4378 gnd.n1026 7.64824
R19452 gnd.n6309 gnd.n1029 7.64824
R19453 gnd.n4411 gnd.n4410 7.64824
R19454 gnd.n6303 gnd.n1039 7.64824
R19455 gnd.n4443 gnd.n4442 7.64824
R19456 gnd.n6297 gnd.n1049 7.64824
R19457 gnd.n4419 gnd.n1057 7.64824
R19458 gnd.n6291 gnd.n1060 7.64824
R19459 gnd.n4431 gnd.n1068 7.64824
R19460 gnd.n6285 gnd.n1071 7.64824
R19461 gnd.n4496 gnd.n4495 7.64824
R19462 gnd.n6279 gnd.n1081 7.64824
R19463 gnd.n4504 gnd.n1089 7.64824
R19464 gnd.n6273 gnd.n1092 7.64824
R19465 gnd.n4513 gnd.n1100 7.64824
R19466 gnd.n4553 gnd.n1109 7.64824
R19467 gnd.n6261 gnd.n1112 7.64824
R19468 gnd.n5223 gnd.t132 7.64824
R19469 gnd.t119 gnd.n1734 7.64824
R19470 gnd.n6016 gnd.n1336 7.64824
R19471 gnd.n5851 gnd.n1338 7.64824
R19472 gnd.n5861 gnd.n5860 7.64824
R19473 gnd.n5872 gnd.n1431 7.64824
R19474 gnd.n5871 gnd.n1435 7.64824
R19475 gnd.n5882 gnd.n1422 7.64824
R19476 gnd.n1424 gnd.n1414 7.64824
R19477 gnd.n5897 gnd.n5896 7.64824
R19478 gnd.n5909 gnd.n1404 7.64824
R19479 gnd.n5907 gnd.n1407 7.64824
R19480 gnd.n5919 gnd.n1394 7.64824
R19481 gnd.n1398 gnd.n1396 7.64824
R19482 gnd.n5958 gnd.n5957 7.64824
R19483 gnd.n5979 gnd.n1370 7.64824
R19484 gnd.n5978 gnd.n1373 7.64824
R19485 gnd.n5987 gnd.n1361 7.64824
R19486 gnd.n5936 gnd.n1364 7.64824
R19487 gnd.n7172 gnd.n399 7.64824
R19488 gnd.n5941 gnd.n402 7.64824
R19489 gnd.n7182 gnd.n390 7.64824
R19490 gnd.n7163 gnd.n7162 7.64824
R19491 gnd.n7196 gnd.n384 7.64824
R19492 gnd.n7218 gnd.n367 7.64824
R19493 gnd.n7190 gnd.n370 7.64824
R19494 gnd.n7206 gnd.n377 7.64824
R19495 gnd.n7227 gnd.n356 7.64824
R19496 gnd.n358 gnd.n350 7.64824
R19497 gnd.n3074 gnd.t220 7.32958
R19498 gnd.t284 gnd.n1945 7.32958
R19499 gnd.n5453 gnd.t154 7.32958
R19500 gnd.t236 gnd.n1646 7.32958
R19501 gnd.n5810 gnd.t255 7.32958
R19502 gnd.n247 gnd.n238 7.32958
R19503 gnd.n4659 gnd.n4658 7.30353
R19504 gnd.n4941 gnd.n4940 7.30353
R19505 gnd.n3034 gnd.n2753 7.01093
R19506 gnd.n2756 gnd.n2754 7.01093
R19507 gnd.n3044 gnd.n3043 7.01093
R19508 gnd.n3055 gnd.n2737 7.01093
R19509 gnd.n3054 gnd.n2740 7.01093
R19510 gnd.n3065 gnd.n2728 7.01093
R19511 gnd.n2731 gnd.n2729 7.01093
R19512 gnd.n3075 gnd.n3074 7.01093
R19513 gnd.n3085 gnd.n2709 7.01093
R19514 gnd.n3084 gnd.n2712 7.01093
R19515 gnd.n3093 gnd.n2703 7.01093
R19516 gnd.n3105 gnd.n2693 7.01093
R19517 gnd.n3115 gnd.n2678 7.01093
R19518 gnd.n3131 gnd.n3130 7.01093
R19519 gnd.n2680 gnd.n2617 7.01093
R19520 gnd.n3185 gnd.n2618 7.01093
R19521 gnd.n3179 gnd.n3178 7.01093
R19522 gnd.n2667 gnd.n2629 7.01093
R19523 gnd.n3171 gnd.n2640 7.01093
R19524 gnd.n2658 gnd.n2653 7.01093
R19525 gnd.n3165 gnd.n3164 7.01093
R19526 gnd.n3211 gnd.n2544 7.01093
R19527 gnd.n3210 gnd.n3209 7.01093
R19528 gnd.n3222 gnd.n3221 7.01093
R19529 gnd.n2537 gnd.n2529 7.01093
R19530 gnd.n3251 gnd.n2517 7.01093
R19531 gnd.n3250 gnd.n2520 7.01093
R19532 gnd.n3261 gnd.n2509 7.01093
R19533 gnd.n2510 gnd.n2498 7.01093
R19534 gnd.n3272 gnd.n2499 7.01093
R19535 gnd.n3296 gnd.n2490 7.01093
R19536 gnd.n3295 gnd.n2481 7.01093
R19537 gnd.n3318 gnd.n3317 7.01093
R19538 gnd.n3336 gnd.n2462 7.01093
R19539 gnd.n3335 gnd.n2465 7.01093
R19540 gnd.n3346 gnd.n2454 7.01093
R19541 gnd.n2455 gnd.n2442 7.01093
R19542 gnd.n3357 gnd.n2443 7.01093
R19543 gnd.n3384 gnd.n2427 7.01093
R19544 gnd.n3396 gnd.n3395 7.01093
R19545 gnd.n3378 gnd.n2420 7.01093
R19546 gnd.n3407 gnd.n3406 7.01093
R19547 gnd.n3679 gnd.n2408 7.01093
R19548 gnd.n3678 gnd.n2411 7.01093
R19549 gnd.n3691 gnd.n2400 7.01093
R19550 gnd.n2401 gnd.n2392 7.01093
R19551 gnd.n3701 gnd.n2393 7.01093
R19552 gnd.t339 gnd.n1866 7.01093
R19553 gnd.n5533 gnd.n1852 7.01093
R19554 gnd.n5222 gnd.n5221 7.01093
R19555 gnd.n5185 gnd.n4804 7.01093
R19556 gnd.n5621 gnd.n1776 7.01093
R19557 gnd.n5669 gnd.n1733 7.01093
R19558 gnd.n4878 gnd.n4876 7.01093
R19559 gnd.t318 gnd.n1713 7.01093
R19560 gnd.n2712 gnd.t223 6.69227
R19561 gnd.n2520 gnd.t58 6.69227
R19562 gnd.n3385 gnd.t213 6.69227
R19563 gnd.n5028 gnd.n5027 6.5566
R19564 gnd.n4672 gnd.n4671 6.5566
R19565 gnd.n5262 gnd.n5258 6.5566
R19566 gnd.n5008 gnd.n4908 6.5566
R19567 gnd.n4736 gnd.t267 6.37362
R19568 gnd.t21 gnd.n1804 6.37362
R19569 gnd.n5155 gnd.t1 6.37362
R19570 gnd.n5693 gnd.t251 6.37362
R19571 gnd.n4535 gnd.n4530 6.20656
R19572 gnd.n7567 gnd.n7564 6.20656
R19573 gnd.n4138 gnd.n3987 6.20656
R19574 gnd.n5829 gnd.n5826 6.20656
R19575 gnd.t56 gnd.n3141 6.05496
R19576 gnd.n3142 gnd.t222 6.05496
R19577 gnd.t64 gnd.n2544 6.05496
R19578 gnd.t217 gnd.n3306 6.05496
R19579 gnd.t234 gnd.n4804 6.05496
R19580 gnd.n5621 gnd.t93 6.05496
R19581 gnd.n3664 gnd.n3634 5.81868
R19582 gnd.n3632 gnd.n3602 5.81868
R19583 gnd.n3600 gnd.n3570 5.81868
R19584 gnd.n3569 gnd.n3539 5.81868
R19585 gnd.n3537 gnd.n3507 5.81868
R19586 gnd.n3505 gnd.n3475 5.81868
R19587 gnd.n3473 gnd.n3443 5.81868
R19588 gnd.n3442 gnd.n3412 5.81868
R19589 gnd.n5541 gnd.n1846 5.73631
R19590 gnd.n4751 gnd.n4750 5.73631
R19591 gnd.n5178 gnd.n5177 5.73631
R19592 gnd.n5613 gnd.n1784 5.73631
R19593 gnd.n5677 gnd.n1726 5.73631
R19594 gnd.n5108 gnd.n5107 5.73631
R19595 gnd.n5021 gnd.n1305 5.62001
R19596 gnd.n5324 gnd.n4602 5.62001
R19597 gnd.n5324 gnd.n4603 5.62001
R19598 gnd.n5015 gnd.n1305 5.62001
R19599 gnd.n2893 gnd.n2888 5.4308
R19600 gnd.n3709 gnd.n2385 5.4308
R19601 gnd.n3209 gnd.t216 5.41765
R19602 gnd.t219 gnd.n3232 5.41765
R19603 gnd.t68 gnd.n2474 5.41765
R19604 gnd.n3662 gnd.n3661 5.04292
R19605 gnd.n3630 gnd.n3629 5.04292
R19606 gnd.n3598 gnd.n3597 5.04292
R19607 gnd.n3567 gnd.n3566 5.04292
R19608 gnd.n3535 gnd.n3534 5.04292
R19609 gnd.n3503 gnd.n3502 5.04292
R19610 gnd.n3471 gnd.n3470 5.04292
R19611 gnd.n3440 gnd.n3439 5.04292
R19612 gnd.n2609 gnd.n2608 4.82753
R19613 gnd.n78 gnd.n77 4.82753
R19614 gnd.n3172 gnd.t221 4.78034
R19615 gnd.n2499 gnd.t210 4.78034
R19616 gnd.t79 gnd.n1900 4.78034
R19617 gnd.n4751 gnd.t191 4.78034
R19618 gnd.t117 gnd.n1726 4.78034
R19619 gnd.n1700 gnd.t298 4.78034
R19620 gnd.n5749 gnd.t103 4.78034
R19621 gnd.n2614 gnd.n2611 4.74817
R19622 gnd.n2664 gnd.n2550 4.74817
R19623 gnd.n2651 gnd.n2549 4.74817
R19624 gnd.n2548 gnd.n2547 4.74817
R19625 gnd.n2660 gnd.n2611 4.74817
R19626 gnd.n2661 gnd.n2550 4.74817
R19627 gnd.n2663 gnd.n2549 4.74817
R19628 gnd.n2650 gnd.n2548 4.74817
R19629 gnd.n7353 gnd.n7352 4.74817
R19630 gnd.n341 gnd.n308 4.74817
R19631 gnd.n7254 gnd.n307 4.74817
R19632 gnd.n331 gnd.n306 4.74817
R19633 gnd.n7332 gnd.n305 4.74817
R19634 gnd.n7353 gnd.n309 4.74817
R19635 gnd.n7351 gnd.n308 4.74817
R19636 gnd.n342 gnd.n307 4.74817
R19637 gnd.n7255 gnd.n306 4.74817
R19638 gnd.n332 gnd.n305 4.74817
R19639 gnd.n4290 gnd.n4288 4.74817
R19640 gnd.n4303 gnd.n2199 4.74817
R19641 gnd.n4307 gnd.n4305 4.74817
R19642 gnd.n4330 gnd.n2173 4.74817
R19643 gnd.n4333 gnd.n4332 4.74817
R19644 gnd.n4288 gnd.n4287 4.74817
R19645 gnd.n4289 gnd.n2199 4.74817
R19646 gnd.n4305 gnd.n4304 4.74817
R19647 gnd.n4306 gnd.n2173 4.74817
R19648 gnd.n4332 gnd.n4331 4.74817
R19649 gnd.n2589 gnd.n2588 4.7074
R19650 gnd.n58 gnd.n57 4.7074
R19651 gnd.n2609 gnd.n2589 4.65959
R19652 gnd.n78 gnd.n58 4.65959
R19653 gnd.n6060 gnd.n1307 4.6132
R19654 gnd.n5325 gnd.n4601 4.6132
R19655 gnd.n5236 gnd.n4743 4.46168
R19656 gnd.n5230 gnd.t95 4.46168
R19657 gnd.n5549 gnd.n1839 4.46168
R19658 gnd.n5605 gnd.n1790 4.46168
R19659 gnd.n5170 gnd.n4817 4.46168
R19660 gnd.n5115 gnd.n4863 4.46168
R19661 gnd.n5109 gnd.t22 4.46168
R19662 gnd.n5685 gnd.n1720 4.46168
R19663 gnd.n4937 gnd.n4924 4.46111
R19664 gnd.n3647 gnd.n3643 4.38594
R19665 gnd.n3615 gnd.n3611 4.38594
R19666 gnd.n3583 gnd.n3579 4.38594
R19667 gnd.n3552 gnd.n3548 4.38594
R19668 gnd.n3520 gnd.n3516 4.38594
R19669 gnd.n3488 gnd.n3484 4.38594
R19670 gnd.n3456 gnd.n3452 4.38594
R19671 gnd.n3425 gnd.n3421 4.38594
R19672 gnd.n3658 gnd.n3636 4.26717
R19673 gnd.n3626 gnd.n3604 4.26717
R19674 gnd.n3594 gnd.n3572 4.26717
R19675 gnd.n3563 gnd.n3541 4.26717
R19676 gnd.n3531 gnd.n3509 4.26717
R19677 gnd.n3499 gnd.n3477 4.26717
R19678 gnd.n3467 gnd.n3445 4.26717
R19679 gnd.n3436 gnd.n3414 4.26717
R19680 gnd.n3116 gnd.t212 4.14303
R19681 gnd.n3346 gnd.t224 4.14303
R19682 gnd.n2109 gnd.t259 4.14303
R19683 gnd.n5842 gnd.t263 4.14303
R19684 gnd.n3666 gnd.n3665 4.08274
R19685 gnd.n5029 gnd.n5028 4.05904
R19686 gnd.n4673 gnd.n4672 4.05904
R19687 gnd.n5265 gnd.n5258 4.05904
R19688 gnd.n5009 gnd.n5008 4.05904
R19689 gnd.n19 gnd.n9 3.99943
R19690 gnd.n5541 gnd.t244 3.82437
R19691 gnd.n4806 gnd.t174 3.82437
R19692 gnd.n4819 gnd.t116 3.82437
R19693 gnd.n3666 gnd.n3538 3.70378
R19694 gnd.n3189 gnd.n2610 3.65935
R19695 gnd.n19 gnd.n18 3.60163
R19696 gnd.n4187 gnd.t314 3.50571
R19697 gnd.n6267 gnd.t259 3.50571
R19698 gnd.t263 gnd.n1452 3.50571
R19699 gnd.n7522 gnd.t247 3.50571
R19700 gnd.n3657 gnd.n3638 3.49141
R19701 gnd.n3625 gnd.n3606 3.49141
R19702 gnd.n3593 gnd.n3574 3.49141
R19703 gnd.n3562 gnd.n3543 3.49141
R19704 gnd.n3530 gnd.n3511 3.49141
R19705 gnd.n3498 gnd.n3479 3.49141
R19706 gnd.n3466 gnd.n3447 3.49141
R19707 gnd.n3435 gnd.n3416 3.49141
R19708 gnd.n5243 gnd.n4736 3.18706
R19709 gnd.n4796 gnd.t0 3.18706
R19710 gnd.n5597 gnd.n1797 3.18706
R19711 gnd.n5163 gnd.n5162 3.18706
R19712 gnd.t135 gnd.n1762 3.18706
R19713 gnd.n5693 gnd.n1713 3.18706
R19714 gnd.n2695 gnd.t212 2.8684
R19715 gnd.n5509 gnd.t24 2.8684
R19716 gnd.t267 gnd.t156 2.8684
R19717 gnd.t203 gnd.t251 2.8684
R19718 gnd.t354 gnd.n1692 2.8684
R19719 gnd.n2590 gnd.t38 2.82907
R19720 gnd.n2590 gnd.t185 2.82907
R19721 gnd.n2592 gnd.t228 2.82907
R19722 gnd.n2592 gnd.t241 2.82907
R19723 gnd.n2594 gnd.t151 2.82907
R19724 gnd.n2594 gnd.t188 2.82907
R19725 gnd.n2596 gnd.t32 2.82907
R19726 gnd.n2596 gnd.t225 2.82907
R19727 gnd.n2598 gnd.t87 2.82907
R19728 gnd.n2598 gnd.t165 2.82907
R19729 gnd.n2600 gnd.t227 2.82907
R19730 gnd.n2600 gnd.t231 2.82907
R19731 gnd.n2602 gnd.t226 2.82907
R19732 gnd.n2602 gnd.t242 2.82907
R19733 gnd.n2604 gnd.t121 2.82907
R19734 gnd.n2604 gnd.t88 2.82907
R19735 gnd.n2606 gnd.t8 2.82907
R19736 gnd.n2606 gnd.t147 2.82907
R19737 gnd.n2551 gnd.t97 2.82907
R19738 gnd.n2551 gnd.t184 2.82907
R19739 gnd.n2553 gnd.t138 2.82907
R19740 gnd.n2553 gnd.t53 2.82907
R19741 gnd.n2555 gnd.t168 2.82907
R19742 gnd.n2555 gnd.t18 2.82907
R19743 gnd.n2557 gnd.t100 2.82907
R19744 gnd.n2557 gnd.t177 2.82907
R19745 gnd.n2559 gnd.t233 2.82907
R19746 gnd.n2559 gnd.t181 2.82907
R19747 gnd.n2561 gnd.t238 2.82907
R19748 gnd.n2561 gnd.t108 2.82907
R19749 gnd.n2563 gnd.t198 2.82907
R19750 gnd.n2563 gnd.t170 2.82907
R19751 gnd.n2565 gnd.t82 2.82907
R19752 gnd.n2565 gnd.t176 2.82907
R19753 gnd.n2567 gnd.t197 2.82907
R19754 gnd.n2567 gnd.t136 2.82907
R19755 gnd.n2570 gnd.t159 2.82907
R19756 gnd.n2570 gnd.t206 2.82907
R19757 gnd.n2572 gnd.t158 2.82907
R19758 gnd.n2572 gnd.t128 2.82907
R19759 gnd.n2574 gnd.t200 2.82907
R19760 gnd.n2574 gnd.t167 2.82907
R19761 gnd.n2576 gnd.t39 2.82907
R19762 gnd.n2576 gnd.t112 2.82907
R19763 gnd.n2578 gnd.t171 2.82907
R19764 gnd.n2578 gnd.t161 2.82907
R19765 gnd.n2580 gnd.t99 2.82907
R19766 gnd.n2580 gnd.t162 2.82907
R19767 gnd.n2582 gnd.t142 2.82907
R19768 gnd.n2582 gnd.t180 2.82907
R19769 gnd.n2584 gnd.t106 2.82907
R19770 gnd.n2584 gnd.t28 2.82907
R19771 gnd.n2586 gnd.t55 2.82907
R19772 gnd.n2586 gnd.t41 2.82907
R19773 gnd.n75 gnd.t90 2.82907
R19774 gnd.n75 gnd.t149 2.82907
R19775 gnd.n73 gnd.t36 2.82907
R19776 gnd.n73 gnd.t230 2.82907
R19777 gnd.n71 gnd.t76 2.82907
R19778 gnd.n71 gnd.t20 2.82907
R19779 gnd.n69 gnd.t205 2.82907
R19780 gnd.n69 gnd.t152 2.82907
R19781 gnd.n67 gnd.t186 2.82907
R19782 gnd.n67 gnd.t229 2.82907
R19783 gnd.n65 gnd.t178 2.82907
R19784 gnd.n65 gnd.t179 2.82907
R19785 gnd.n63 gnd.t85 2.82907
R19786 gnd.n63 gnd.t6 2.82907
R19787 gnd.n61 gnd.t34 2.82907
R19788 gnd.n61 gnd.t120 2.82907
R19789 gnd.n59 gnd.t187 2.82907
R19790 gnd.n59 gnd.t146 2.82907
R19791 gnd.n36 gnd.t109 2.82907
R19792 gnd.n36 gnd.t202 2.82907
R19793 gnd.n34 gnd.t240 2.82907
R19794 gnd.n34 gnd.t51 2.82907
R19795 gnd.n32 gnd.t12 2.82907
R19796 gnd.n32 gnd.t358 2.82907
R19797 gnd.n30 gnd.t14 2.82907
R19798 gnd.n30 gnd.t54 2.82907
R19799 gnd.n28 gnd.t102 2.82907
R19800 gnd.n28 gnd.t196 2.82907
R19801 gnd.n26 gnd.t173 2.82907
R19802 gnd.n26 gnd.t47 2.82907
R19803 gnd.n24 gnd.t139 2.82907
R19804 gnd.n24 gnd.t201 2.82907
R19805 gnd.n22 gnd.t239 2.82907
R19806 gnd.n22 gnd.t16 2.82907
R19807 gnd.n20 gnd.t49 2.82907
R19808 gnd.n20 gnd.t45 2.82907
R19809 gnd.n55 gnd.t166 2.82907
R19810 gnd.n55 gnd.t164 2.82907
R19811 gnd.n53 gnd.t114 2.82907
R19812 gnd.n53 gnd.t140 2.82907
R19813 gnd.n51 gnd.t91 2.82907
R19814 gnd.n51 gnd.t110 2.82907
R19815 gnd.n49 gnd.t356 2.82907
R19816 gnd.n49 gnd.t10 2.82907
R19817 gnd.n47 gnd.t207 2.82907
R19818 gnd.n47 gnd.t199 2.82907
R19819 gnd.n45 gnd.t357 2.82907
R19820 gnd.n45 gnd.t105 2.82907
R19821 gnd.n43 gnd.t182 2.82907
R19822 gnd.n43 gnd.t163 2.82907
R19823 gnd.n41 gnd.t143 2.82907
R19824 gnd.n41 gnd.t175 2.82907
R19825 gnd.n39 gnd.t72 2.82907
R19826 gnd.n39 gnd.t232 2.82907
R19827 gnd.n3654 gnd.n3653 2.71565
R19828 gnd.n3622 gnd.n3621 2.71565
R19829 gnd.n3590 gnd.n3589 2.71565
R19830 gnd.n3559 gnd.n3558 2.71565
R19831 gnd.n3527 gnd.n3526 2.71565
R19832 gnd.n3495 gnd.n3494 2.71565
R19833 gnd.n3463 gnd.n3462 2.71565
R19834 gnd.n3432 gnd.n3431 2.71565
R19835 gnd.n5250 gnd.t281 2.54975
R19836 gnd.n5597 gnd.t129 2.54975
R19837 gnd.n5162 gnd.t23 2.54975
R19838 gnd.n5092 gnd.t278 2.54975
R19839 gnd.n3189 gnd.n2611 2.27742
R19840 gnd.n3189 gnd.n2550 2.27742
R19841 gnd.n3189 gnd.n2549 2.27742
R19842 gnd.n3189 gnd.n2548 2.27742
R19843 gnd.n7354 gnd.n7353 2.27742
R19844 gnd.n7354 gnd.n308 2.27742
R19845 gnd.n7354 gnd.n307 2.27742
R19846 gnd.n7354 gnd.n306 2.27742
R19847 gnd.n7354 gnd.n305 2.27742
R19848 gnd.n4288 gnd.n966 2.27742
R19849 gnd.n2199 gnd.n966 2.27742
R19850 gnd.n4305 gnd.n966 2.27742
R19851 gnd.n2173 gnd.n966 2.27742
R19852 gnd.n4332 gnd.n966 2.27742
R19853 gnd.n3043 gnd.t329 2.23109
R19854 gnd.n2666 gnd.t221 2.23109
R19855 gnd.n4361 gnd.t150 2.23109
R19856 gnd.t5 gnd.n367 2.23109
R19857 gnd.n3650 gnd.n3640 1.93989
R19858 gnd.n3618 gnd.n3608 1.93989
R19859 gnd.n3586 gnd.n3576 1.93989
R19860 gnd.n3555 gnd.n3545 1.93989
R19861 gnd.n3523 gnd.n3513 1.93989
R19862 gnd.n3491 gnd.n3481 1.93989
R19863 gnd.n3459 gnd.n3449 1.93989
R19864 gnd.n3428 gnd.n3418 1.93989
R19865 gnd.n5250 gnd.n4663 1.91244
R19866 gnd.n5220 gnd.t126 1.91244
R19867 gnd.t2 gnd.n1819 1.91244
R19868 gnd.n5589 gnd.n1804 1.91244
R19869 gnd.n5155 gnd.n4831 1.91244
R19870 gnd.n5645 gnd.t96 1.91244
R19871 gnd.n5122 gnd.t115 1.91244
R19872 gnd.n5701 gnd.n1706 1.91244
R19873 gnd.t70 gnd.n3054 1.59378
R19874 gnd.n3233 gnd.t219 1.59378
R19875 gnd.n2483 gnd.t68 1.59378
R19876 gnd.n4227 gnd.t40 1.59378
R19877 gnd.n4410 gnd.t52 1.59378
R19878 gnd.n6297 gnd.t37 1.59378
R19879 gnd.n5565 gnd.t122 1.59378
R19880 gnd.t352 gnd.n4853 1.59378
R19881 gnd.n1398 gnd.t44 1.59378
R19882 gnd.t33 gnd.n5978 1.59378
R19883 gnd.n7414 gnd.t89 1.59378
R19884 gnd.n5557 gnd.t126 1.27512
R19885 gnd.t115 gnd.n4857 1.27512
R19886 gnd.n2896 gnd.n2888 1.16414
R19887 gnd.n3712 gnd.n2385 1.16414
R19888 gnd.n3649 gnd.n3642 1.16414
R19889 gnd.n3617 gnd.n3610 1.16414
R19890 gnd.n3585 gnd.n3578 1.16414
R19891 gnd.n3554 gnd.n3547 1.16414
R19892 gnd.n3522 gnd.n3515 1.16414
R19893 gnd.n3490 gnd.n3483 1.16414
R19894 gnd.n3458 gnd.n3451 1.16414
R19895 gnd.n3427 gnd.n3420 1.16414
R19896 gnd.n6060 gnd.n6059 0.970197
R19897 gnd.n5325 gnd.n2082 0.970197
R19898 gnd.n3633 gnd.n3601 0.962709
R19899 gnd.n3665 gnd.n3633 0.962709
R19900 gnd.n3506 gnd.n3474 0.962709
R19901 gnd.n3538 gnd.n3506 0.962709
R19902 gnd.n3142 gnd.t56 0.956468
R19903 gnd.n3307 gnd.t217 0.956468
R19904 gnd.n4259 gnd.t141 0.956468
R19905 gnd.n6321 gnd.t17 0.956468
R19906 gnd.n4495 gnd.t42 0.956468
R19907 gnd.t0 gnd.t124 0.956468
R19908 gnd.t193 gnd.t135 0.956468
R19909 gnd.t29 gnd.n1424 0.956468
R19910 gnd.n7182 gnd.t84 0.956468
R19911 gnd.n7382 gnd.t19 0.956468
R19912 gnd.n2601 gnd.n2599 0.773756
R19913 gnd.n70 gnd.n68 0.773756
R19914 gnd.n2608 gnd.n2607 0.773756
R19915 gnd.n2607 gnd.n2605 0.773756
R19916 gnd.n2605 gnd.n2603 0.773756
R19917 gnd.n2603 gnd.n2601 0.773756
R19918 gnd.n2599 gnd.n2597 0.773756
R19919 gnd.n2597 gnd.n2595 0.773756
R19920 gnd.n2595 gnd.n2593 0.773756
R19921 gnd.n2593 gnd.n2591 0.773756
R19922 gnd.n62 gnd.n60 0.773756
R19923 gnd.n64 gnd.n62 0.773756
R19924 gnd.n66 gnd.n64 0.773756
R19925 gnd.n68 gnd.n66 0.773756
R19926 gnd.n72 gnd.n70 0.773756
R19927 gnd.n74 gnd.n72 0.773756
R19928 gnd.n76 gnd.n74 0.773756
R19929 gnd.n77 gnd.n76 0.773756
R19930 gnd gnd.n0 0.70738
R19931 gnd.n2 gnd.n1 0.672012
R19932 gnd.n3 gnd.n2 0.672012
R19933 gnd.n4 gnd.n3 0.672012
R19934 gnd.n5 gnd.n4 0.672012
R19935 gnd.n6 gnd.n5 0.672012
R19936 gnd.n7 gnd.n6 0.672012
R19937 gnd.n8 gnd.n7 0.672012
R19938 gnd.n9 gnd.n8 0.672012
R19939 gnd.n11 gnd.n10 0.672012
R19940 gnd.n12 gnd.n11 0.672012
R19941 gnd.n13 gnd.n12 0.672012
R19942 gnd.n14 gnd.n13 0.672012
R19943 gnd.n15 gnd.n14 0.672012
R19944 gnd.n16 gnd.n15 0.672012
R19945 gnd.n17 gnd.n16 0.672012
R19946 gnd.n18 gnd.n17 0.672012
R19947 gnd.n5207 gnd.t189 0.637812
R19948 gnd.n5573 gnd.n1818 0.637812
R19949 gnd.n5581 gnd.n1812 0.637812
R19950 gnd.n5148 gnd.n5147 0.637812
R19951 gnd.n4849 gnd.n4844 0.637812
R19952 gnd.n5135 gnd.t127 0.637812
R19953 gnd.n5685 gnd.t301 0.637812
R19954 gnd.n7657 gnd.n7656 0.637193
R19955 gnd.n2569 gnd.n2568 0.573776
R19956 gnd.n2568 gnd.n2566 0.573776
R19957 gnd.n2566 gnd.n2564 0.573776
R19958 gnd.n2564 gnd.n2562 0.573776
R19959 gnd.n2562 gnd.n2560 0.573776
R19960 gnd.n2560 gnd.n2558 0.573776
R19961 gnd.n2558 gnd.n2556 0.573776
R19962 gnd.n2556 gnd.n2554 0.573776
R19963 gnd.n2554 gnd.n2552 0.573776
R19964 gnd.n2588 gnd.n2587 0.573776
R19965 gnd.n2587 gnd.n2585 0.573776
R19966 gnd.n2585 gnd.n2583 0.573776
R19967 gnd.n2583 gnd.n2581 0.573776
R19968 gnd.n2581 gnd.n2579 0.573776
R19969 gnd.n2579 gnd.n2577 0.573776
R19970 gnd.n2577 gnd.n2575 0.573776
R19971 gnd.n2575 gnd.n2573 0.573776
R19972 gnd.n2573 gnd.n2571 0.573776
R19973 gnd.n23 gnd.n21 0.573776
R19974 gnd.n25 gnd.n23 0.573776
R19975 gnd.n27 gnd.n25 0.573776
R19976 gnd.n29 gnd.n27 0.573776
R19977 gnd.n31 gnd.n29 0.573776
R19978 gnd.n33 gnd.n31 0.573776
R19979 gnd.n35 gnd.n33 0.573776
R19980 gnd.n37 gnd.n35 0.573776
R19981 gnd.n38 gnd.n37 0.573776
R19982 gnd.n42 gnd.n40 0.573776
R19983 gnd.n44 gnd.n42 0.573776
R19984 gnd.n46 gnd.n44 0.573776
R19985 gnd.n48 gnd.n46 0.573776
R19986 gnd.n50 gnd.n48 0.573776
R19987 gnd.n52 gnd.n50 0.573776
R19988 gnd.n54 gnd.n52 0.573776
R19989 gnd.n56 gnd.n54 0.573776
R19990 gnd.n57 gnd.n56 0.573776
R19991 gnd.n7354 gnd.n304 0.5435
R19992 gnd.n6344 gnd.n966 0.5435
R19993 gnd.n3369 gnd.n2389 0.486781
R19994 gnd.n1518 gnd.n1242 0.486781
R19995 gnd.n2945 gnd.n2944 0.48678
R19996 gnd.n6256 gnd.n6255 0.485256
R19997 gnd.n3686 gnd.n2343 0.480683
R19998 gnd.n3029 gnd.n3028 0.480683
R19999 gnd.n6516 gnd.n6515 0.480683
R20000 gnd.n6937 gnd.n6936 0.480683
R20001 gnd.n3863 gnd.n3862 0.477634
R20002 gnd.n4182 gnd.n2317 0.477634
R20003 gnd.n7505 gnd.n7504 0.477634
R20004 gnd.n7607 gnd.n7606 0.477634
R20005 gnd.n7599 gnd.n7598 0.465439
R20006 gnd.n7528 gnd.n7527 0.465439
R20007 gnd.n6020 gnd.n1333 0.465439
R20008 gnd.n5845 gnd.n1289 0.465439
R20009 gnd.n2066 gnd.n1107 0.465439
R20010 gnd.n4558 gnd.n4557 0.465439
R20011 gnd.n4101 gnd.n4096 0.465439
R20012 gnd.n4176 gnd.n4175 0.465439
R20013 gnd.n5816 gnd.n5815 0.451719
R20014 gnd.n5409 gnd.n5408 0.451719
R20015 gnd.n4538 gnd.n4530 0.388379
R20016 gnd.n3646 gnd.n3645 0.388379
R20017 gnd.n3614 gnd.n3613 0.388379
R20018 gnd.n3582 gnd.n3581 0.388379
R20019 gnd.n3551 gnd.n3550 0.388379
R20020 gnd.n3519 gnd.n3518 0.388379
R20021 gnd.n3487 gnd.n3486 0.388379
R20022 gnd.n3455 gnd.n3454 0.388379
R20023 gnd.n3424 gnd.n3423 0.388379
R20024 gnd.n7568 gnd.n7567 0.388379
R20025 gnd.n3987 gnd.n3983 0.388379
R20026 gnd.n5830 gnd.n5829 0.388379
R20027 gnd.n6258 gnd.n6257 0.378829
R20028 gnd.n6013 gnd.n1342 0.377553
R20029 gnd.n7657 gnd.n19 0.374463
R20030 gnd gnd.n7657 0.367492
R20031 gnd.n2445 gnd.t213 0.319156
R20032 gnd.n4292 gnd.t107 0.319156
R20033 gnd.n4335 gnd.t31 0.319156
R20034 gnd.n5213 gnd.t122 0.319156
R20035 gnd.n5129 gnd.t352 0.319156
R20036 gnd.n7242 gnd.t46 0.319156
R20037 gnd.n7334 gnd.t13 0.319156
R20038 gnd.n2863 gnd.n2841 0.311721
R20039 gnd.n7148 gnd.n304 0.282512
R20040 gnd.n6345 gnd.n6344 0.282512
R20041 gnd.n3757 gnd.n3756 0.268793
R20042 gnd.n4549 gnd.n4548 0.247451
R20043 gnd.n5840 gnd.n5839 0.247451
R20044 gnd.n3756 gnd.n3755 0.241354
R20045 gnd.n1307 gnd.n1304 0.229039
R20046 gnd.n1310 gnd.n1307 0.229039
R20047 gnd.n4601 gnd.n2081 0.229039
R20048 gnd.n4601 gnd.n4600 0.229039
R20049 gnd.n2610 gnd.n0 0.210825
R20050 gnd.n3017 gnd.n2816 0.206293
R20051 gnd.n420 gnd.n304 0.198671
R20052 gnd.n6344 gnd.n6343 0.198671
R20053 gnd.n3663 gnd.n3635 0.155672
R20054 gnd.n3656 gnd.n3635 0.155672
R20055 gnd.n3656 gnd.n3655 0.155672
R20056 gnd.n3655 gnd.n3639 0.155672
R20057 gnd.n3648 gnd.n3639 0.155672
R20058 gnd.n3648 gnd.n3647 0.155672
R20059 gnd.n3631 gnd.n3603 0.155672
R20060 gnd.n3624 gnd.n3603 0.155672
R20061 gnd.n3624 gnd.n3623 0.155672
R20062 gnd.n3623 gnd.n3607 0.155672
R20063 gnd.n3616 gnd.n3607 0.155672
R20064 gnd.n3616 gnd.n3615 0.155672
R20065 gnd.n3599 gnd.n3571 0.155672
R20066 gnd.n3592 gnd.n3571 0.155672
R20067 gnd.n3592 gnd.n3591 0.155672
R20068 gnd.n3591 gnd.n3575 0.155672
R20069 gnd.n3584 gnd.n3575 0.155672
R20070 gnd.n3584 gnd.n3583 0.155672
R20071 gnd.n3568 gnd.n3540 0.155672
R20072 gnd.n3561 gnd.n3540 0.155672
R20073 gnd.n3561 gnd.n3560 0.155672
R20074 gnd.n3560 gnd.n3544 0.155672
R20075 gnd.n3553 gnd.n3544 0.155672
R20076 gnd.n3553 gnd.n3552 0.155672
R20077 gnd.n3536 gnd.n3508 0.155672
R20078 gnd.n3529 gnd.n3508 0.155672
R20079 gnd.n3529 gnd.n3528 0.155672
R20080 gnd.n3528 gnd.n3512 0.155672
R20081 gnd.n3521 gnd.n3512 0.155672
R20082 gnd.n3521 gnd.n3520 0.155672
R20083 gnd.n3504 gnd.n3476 0.155672
R20084 gnd.n3497 gnd.n3476 0.155672
R20085 gnd.n3497 gnd.n3496 0.155672
R20086 gnd.n3496 gnd.n3480 0.155672
R20087 gnd.n3489 gnd.n3480 0.155672
R20088 gnd.n3489 gnd.n3488 0.155672
R20089 gnd.n3472 gnd.n3444 0.155672
R20090 gnd.n3465 gnd.n3444 0.155672
R20091 gnd.n3465 gnd.n3464 0.155672
R20092 gnd.n3464 gnd.n3448 0.155672
R20093 gnd.n3457 gnd.n3448 0.155672
R20094 gnd.n3457 gnd.n3456 0.155672
R20095 gnd.n3441 gnd.n3413 0.155672
R20096 gnd.n3434 gnd.n3413 0.155672
R20097 gnd.n3434 gnd.n3433 0.155672
R20098 gnd.n3433 gnd.n3417 0.155672
R20099 gnd.n3426 gnd.n3417 0.155672
R20100 gnd.n3426 gnd.n3425 0.155672
R20101 gnd.n3788 gnd.n2343 0.152939
R20102 gnd.n3788 gnd.n3787 0.152939
R20103 gnd.n3787 gnd.n3786 0.152939
R20104 gnd.n3786 gnd.n2345 0.152939
R20105 gnd.n2346 gnd.n2345 0.152939
R20106 gnd.n2347 gnd.n2346 0.152939
R20107 gnd.n2348 gnd.n2347 0.152939
R20108 gnd.n2349 gnd.n2348 0.152939
R20109 gnd.n2350 gnd.n2349 0.152939
R20110 gnd.n2351 gnd.n2350 0.152939
R20111 gnd.n2352 gnd.n2351 0.152939
R20112 gnd.n2353 gnd.n2352 0.152939
R20113 gnd.n2354 gnd.n2353 0.152939
R20114 gnd.n2355 gnd.n2354 0.152939
R20115 gnd.n3758 gnd.n2355 0.152939
R20116 gnd.n3758 gnd.n3757 0.152939
R20117 gnd.n3030 gnd.n3029 0.152939
R20118 gnd.n3030 gnd.n2734 0.152939
R20119 gnd.n3058 gnd.n2734 0.152939
R20120 gnd.n3059 gnd.n3058 0.152939
R20121 gnd.n3060 gnd.n3059 0.152939
R20122 gnd.n3061 gnd.n3060 0.152939
R20123 gnd.n3061 gnd.n2706 0.152939
R20124 gnd.n3088 gnd.n2706 0.152939
R20125 gnd.n3089 gnd.n3088 0.152939
R20126 gnd.n3090 gnd.n3089 0.152939
R20127 gnd.n3090 gnd.n2684 0.152939
R20128 gnd.n3119 gnd.n2684 0.152939
R20129 gnd.n3120 gnd.n3119 0.152939
R20130 gnd.n3121 gnd.n3120 0.152939
R20131 gnd.n3122 gnd.n3121 0.152939
R20132 gnd.n3124 gnd.n3122 0.152939
R20133 gnd.n3124 gnd.n3123 0.152939
R20134 gnd.n3123 gnd.n2633 0.152939
R20135 gnd.n2634 gnd.n2633 0.152939
R20136 gnd.n2635 gnd.n2634 0.152939
R20137 gnd.n2654 gnd.n2635 0.152939
R20138 gnd.n2655 gnd.n2654 0.152939
R20139 gnd.n2655 gnd.n2541 0.152939
R20140 gnd.n3214 gnd.n2541 0.152939
R20141 gnd.n3215 gnd.n3214 0.152939
R20142 gnd.n3216 gnd.n3215 0.152939
R20143 gnd.n3217 gnd.n3216 0.152939
R20144 gnd.n3217 gnd.n2514 0.152939
R20145 gnd.n3254 gnd.n2514 0.152939
R20146 gnd.n3255 gnd.n3254 0.152939
R20147 gnd.n3256 gnd.n3255 0.152939
R20148 gnd.n3257 gnd.n3256 0.152939
R20149 gnd.n3257 gnd.n2487 0.152939
R20150 gnd.n3299 gnd.n2487 0.152939
R20151 gnd.n3300 gnd.n3299 0.152939
R20152 gnd.n3301 gnd.n3300 0.152939
R20153 gnd.n3302 gnd.n3301 0.152939
R20154 gnd.n3302 gnd.n2459 0.152939
R20155 gnd.n3339 gnd.n2459 0.152939
R20156 gnd.n3340 gnd.n3339 0.152939
R20157 gnd.n3341 gnd.n3340 0.152939
R20158 gnd.n3342 gnd.n3341 0.152939
R20159 gnd.n3342 gnd.n2432 0.152939
R20160 gnd.n3388 gnd.n2432 0.152939
R20161 gnd.n3389 gnd.n3388 0.152939
R20162 gnd.n3390 gnd.n3389 0.152939
R20163 gnd.n3391 gnd.n3390 0.152939
R20164 gnd.n3391 gnd.n2405 0.152939
R20165 gnd.n3682 gnd.n2405 0.152939
R20166 gnd.n3683 gnd.n3682 0.152939
R20167 gnd.n3684 gnd.n3683 0.152939
R20168 gnd.n3685 gnd.n3684 0.152939
R20169 gnd.n3686 gnd.n3685 0.152939
R20170 gnd.n3028 gnd.n2758 0.152939
R20171 gnd.n2779 gnd.n2758 0.152939
R20172 gnd.n2780 gnd.n2779 0.152939
R20173 gnd.n2786 gnd.n2780 0.152939
R20174 gnd.n2787 gnd.n2786 0.152939
R20175 gnd.n2788 gnd.n2787 0.152939
R20176 gnd.n2788 gnd.n2777 0.152939
R20177 gnd.n2796 gnd.n2777 0.152939
R20178 gnd.n2797 gnd.n2796 0.152939
R20179 gnd.n2798 gnd.n2797 0.152939
R20180 gnd.n2798 gnd.n2775 0.152939
R20181 gnd.n2806 gnd.n2775 0.152939
R20182 gnd.n2807 gnd.n2806 0.152939
R20183 gnd.n2808 gnd.n2807 0.152939
R20184 gnd.n2808 gnd.n2773 0.152939
R20185 gnd.n2816 gnd.n2773 0.152939
R20186 gnd.n3755 gnd.n2360 0.152939
R20187 gnd.n2362 gnd.n2360 0.152939
R20188 gnd.n2363 gnd.n2362 0.152939
R20189 gnd.n2364 gnd.n2363 0.152939
R20190 gnd.n2365 gnd.n2364 0.152939
R20191 gnd.n2366 gnd.n2365 0.152939
R20192 gnd.n2367 gnd.n2366 0.152939
R20193 gnd.n2368 gnd.n2367 0.152939
R20194 gnd.n2369 gnd.n2368 0.152939
R20195 gnd.n2370 gnd.n2369 0.152939
R20196 gnd.n2371 gnd.n2370 0.152939
R20197 gnd.n2372 gnd.n2371 0.152939
R20198 gnd.n2373 gnd.n2372 0.152939
R20199 gnd.n2374 gnd.n2373 0.152939
R20200 gnd.n2375 gnd.n2374 0.152939
R20201 gnd.n2376 gnd.n2375 0.152939
R20202 gnd.n2377 gnd.n2376 0.152939
R20203 gnd.n2378 gnd.n2377 0.152939
R20204 gnd.n2379 gnd.n2378 0.152939
R20205 gnd.n2380 gnd.n2379 0.152939
R20206 gnd.n2381 gnd.n2380 0.152939
R20207 gnd.n2382 gnd.n2381 0.152939
R20208 gnd.n2386 gnd.n2382 0.152939
R20209 gnd.n2387 gnd.n2386 0.152939
R20210 gnd.n2388 gnd.n2387 0.152939
R20211 gnd.n2389 gnd.n2388 0.152939
R20212 gnd.n3191 gnd.n3190 0.152939
R20213 gnd.n3192 gnd.n3191 0.152939
R20214 gnd.n3193 gnd.n3192 0.152939
R20215 gnd.n3194 gnd.n3193 0.152939
R20216 gnd.n3195 gnd.n3194 0.152939
R20217 gnd.n3196 gnd.n3195 0.152939
R20218 gnd.n3196 gnd.n2495 0.152939
R20219 gnd.n3275 gnd.n2495 0.152939
R20220 gnd.n3276 gnd.n3275 0.152939
R20221 gnd.n3277 gnd.n3276 0.152939
R20222 gnd.n3278 gnd.n3277 0.152939
R20223 gnd.n3279 gnd.n3278 0.152939
R20224 gnd.n3280 gnd.n3279 0.152939
R20225 gnd.n3281 gnd.n3280 0.152939
R20226 gnd.n3282 gnd.n3281 0.152939
R20227 gnd.n3283 gnd.n3282 0.152939
R20228 gnd.n3283 gnd.n2439 0.152939
R20229 gnd.n3360 gnd.n2439 0.152939
R20230 gnd.n3361 gnd.n3360 0.152939
R20231 gnd.n3362 gnd.n3361 0.152939
R20232 gnd.n3363 gnd.n3362 0.152939
R20233 gnd.n3364 gnd.n3363 0.152939
R20234 gnd.n3365 gnd.n3364 0.152939
R20235 gnd.n3366 gnd.n3365 0.152939
R20236 gnd.n3367 gnd.n3366 0.152939
R20237 gnd.n3368 gnd.n3367 0.152939
R20238 gnd.n3370 gnd.n3368 0.152939
R20239 gnd.n3370 gnd.n3369 0.152939
R20240 gnd.n2946 gnd.n2945 0.152939
R20241 gnd.n2946 gnd.n2836 0.152939
R20242 gnd.n2961 gnd.n2836 0.152939
R20243 gnd.n2962 gnd.n2961 0.152939
R20244 gnd.n2963 gnd.n2962 0.152939
R20245 gnd.n2963 gnd.n2824 0.152939
R20246 gnd.n2977 gnd.n2824 0.152939
R20247 gnd.n2978 gnd.n2977 0.152939
R20248 gnd.n2979 gnd.n2978 0.152939
R20249 gnd.n2980 gnd.n2979 0.152939
R20250 gnd.n2981 gnd.n2980 0.152939
R20251 gnd.n2982 gnd.n2981 0.152939
R20252 gnd.n2983 gnd.n2982 0.152939
R20253 gnd.n2984 gnd.n2983 0.152939
R20254 gnd.n2985 gnd.n2984 0.152939
R20255 gnd.n2986 gnd.n2985 0.152939
R20256 gnd.n2987 gnd.n2986 0.152939
R20257 gnd.n2988 gnd.n2987 0.152939
R20258 gnd.n2989 gnd.n2988 0.152939
R20259 gnd.n2990 gnd.n2989 0.152939
R20260 gnd.n2991 gnd.n2990 0.152939
R20261 gnd.n2991 gnd.n2690 0.152939
R20262 gnd.n3108 gnd.n2690 0.152939
R20263 gnd.n3109 gnd.n3108 0.152939
R20264 gnd.n3110 gnd.n3109 0.152939
R20265 gnd.n3111 gnd.n3110 0.152939
R20266 gnd.n3111 gnd.n2612 0.152939
R20267 gnd.n3188 gnd.n2612 0.152939
R20268 gnd.n2864 gnd.n2863 0.152939
R20269 gnd.n2865 gnd.n2864 0.152939
R20270 gnd.n2866 gnd.n2865 0.152939
R20271 gnd.n2867 gnd.n2866 0.152939
R20272 gnd.n2868 gnd.n2867 0.152939
R20273 gnd.n2869 gnd.n2868 0.152939
R20274 gnd.n2870 gnd.n2869 0.152939
R20275 gnd.n2871 gnd.n2870 0.152939
R20276 gnd.n2872 gnd.n2871 0.152939
R20277 gnd.n2873 gnd.n2872 0.152939
R20278 gnd.n2874 gnd.n2873 0.152939
R20279 gnd.n2875 gnd.n2874 0.152939
R20280 gnd.n2876 gnd.n2875 0.152939
R20281 gnd.n2877 gnd.n2876 0.152939
R20282 gnd.n2878 gnd.n2877 0.152939
R20283 gnd.n2879 gnd.n2878 0.152939
R20284 gnd.n2880 gnd.n2879 0.152939
R20285 gnd.n2881 gnd.n2880 0.152939
R20286 gnd.n2882 gnd.n2881 0.152939
R20287 gnd.n2883 gnd.n2882 0.152939
R20288 gnd.n2884 gnd.n2883 0.152939
R20289 gnd.n2885 gnd.n2884 0.152939
R20290 gnd.n2889 gnd.n2885 0.152939
R20291 gnd.n2890 gnd.n2889 0.152939
R20292 gnd.n2890 gnd.n2847 0.152939
R20293 gnd.n2944 gnd.n2847 0.152939
R20294 gnd.n6516 gnd.n794 0.152939
R20295 gnd.n6524 gnd.n794 0.152939
R20296 gnd.n6525 gnd.n6524 0.152939
R20297 gnd.n6526 gnd.n6525 0.152939
R20298 gnd.n6526 gnd.n788 0.152939
R20299 gnd.n6534 gnd.n788 0.152939
R20300 gnd.n6535 gnd.n6534 0.152939
R20301 gnd.n6536 gnd.n6535 0.152939
R20302 gnd.n6536 gnd.n782 0.152939
R20303 gnd.n6544 gnd.n782 0.152939
R20304 gnd.n6545 gnd.n6544 0.152939
R20305 gnd.n6546 gnd.n6545 0.152939
R20306 gnd.n6546 gnd.n776 0.152939
R20307 gnd.n6554 gnd.n776 0.152939
R20308 gnd.n6555 gnd.n6554 0.152939
R20309 gnd.n6556 gnd.n6555 0.152939
R20310 gnd.n6556 gnd.n770 0.152939
R20311 gnd.n6564 gnd.n770 0.152939
R20312 gnd.n6565 gnd.n6564 0.152939
R20313 gnd.n6566 gnd.n6565 0.152939
R20314 gnd.n6566 gnd.n764 0.152939
R20315 gnd.n6574 gnd.n764 0.152939
R20316 gnd.n6575 gnd.n6574 0.152939
R20317 gnd.n6576 gnd.n6575 0.152939
R20318 gnd.n6576 gnd.n758 0.152939
R20319 gnd.n6584 gnd.n758 0.152939
R20320 gnd.n6585 gnd.n6584 0.152939
R20321 gnd.n6586 gnd.n6585 0.152939
R20322 gnd.n6586 gnd.n752 0.152939
R20323 gnd.n6594 gnd.n752 0.152939
R20324 gnd.n6595 gnd.n6594 0.152939
R20325 gnd.n6596 gnd.n6595 0.152939
R20326 gnd.n6596 gnd.n746 0.152939
R20327 gnd.n6604 gnd.n746 0.152939
R20328 gnd.n6605 gnd.n6604 0.152939
R20329 gnd.n6606 gnd.n6605 0.152939
R20330 gnd.n6606 gnd.n740 0.152939
R20331 gnd.n6614 gnd.n740 0.152939
R20332 gnd.n6615 gnd.n6614 0.152939
R20333 gnd.n6616 gnd.n6615 0.152939
R20334 gnd.n6616 gnd.n734 0.152939
R20335 gnd.n6624 gnd.n734 0.152939
R20336 gnd.n6625 gnd.n6624 0.152939
R20337 gnd.n6626 gnd.n6625 0.152939
R20338 gnd.n6626 gnd.n728 0.152939
R20339 gnd.n6634 gnd.n728 0.152939
R20340 gnd.n6635 gnd.n6634 0.152939
R20341 gnd.n6636 gnd.n6635 0.152939
R20342 gnd.n6636 gnd.n722 0.152939
R20343 gnd.n6644 gnd.n722 0.152939
R20344 gnd.n6645 gnd.n6644 0.152939
R20345 gnd.n6646 gnd.n6645 0.152939
R20346 gnd.n6646 gnd.n716 0.152939
R20347 gnd.n6654 gnd.n716 0.152939
R20348 gnd.n6655 gnd.n6654 0.152939
R20349 gnd.n6656 gnd.n6655 0.152939
R20350 gnd.n6656 gnd.n710 0.152939
R20351 gnd.n6664 gnd.n710 0.152939
R20352 gnd.n6665 gnd.n6664 0.152939
R20353 gnd.n6666 gnd.n6665 0.152939
R20354 gnd.n6666 gnd.n704 0.152939
R20355 gnd.n6674 gnd.n704 0.152939
R20356 gnd.n6675 gnd.n6674 0.152939
R20357 gnd.n6676 gnd.n6675 0.152939
R20358 gnd.n6676 gnd.n698 0.152939
R20359 gnd.n6684 gnd.n698 0.152939
R20360 gnd.n6685 gnd.n6684 0.152939
R20361 gnd.n6686 gnd.n6685 0.152939
R20362 gnd.n6686 gnd.n692 0.152939
R20363 gnd.n6694 gnd.n692 0.152939
R20364 gnd.n6695 gnd.n6694 0.152939
R20365 gnd.n6696 gnd.n6695 0.152939
R20366 gnd.n6696 gnd.n686 0.152939
R20367 gnd.n6704 gnd.n686 0.152939
R20368 gnd.n6705 gnd.n6704 0.152939
R20369 gnd.n6706 gnd.n6705 0.152939
R20370 gnd.n6706 gnd.n680 0.152939
R20371 gnd.n6714 gnd.n680 0.152939
R20372 gnd.n6715 gnd.n6714 0.152939
R20373 gnd.n6716 gnd.n6715 0.152939
R20374 gnd.n6716 gnd.n674 0.152939
R20375 gnd.n6724 gnd.n674 0.152939
R20376 gnd.n6725 gnd.n6724 0.152939
R20377 gnd.n6726 gnd.n6725 0.152939
R20378 gnd.n6726 gnd.n668 0.152939
R20379 gnd.n6734 gnd.n668 0.152939
R20380 gnd.n6735 gnd.n6734 0.152939
R20381 gnd.n6736 gnd.n6735 0.152939
R20382 gnd.n6736 gnd.n662 0.152939
R20383 gnd.n6744 gnd.n662 0.152939
R20384 gnd.n6745 gnd.n6744 0.152939
R20385 gnd.n6746 gnd.n6745 0.152939
R20386 gnd.n6746 gnd.n656 0.152939
R20387 gnd.n6754 gnd.n656 0.152939
R20388 gnd.n6755 gnd.n6754 0.152939
R20389 gnd.n6756 gnd.n6755 0.152939
R20390 gnd.n6756 gnd.n650 0.152939
R20391 gnd.n6764 gnd.n650 0.152939
R20392 gnd.n6765 gnd.n6764 0.152939
R20393 gnd.n6766 gnd.n6765 0.152939
R20394 gnd.n6766 gnd.n644 0.152939
R20395 gnd.n6774 gnd.n644 0.152939
R20396 gnd.n6775 gnd.n6774 0.152939
R20397 gnd.n6776 gnd.n6775 0.152939
R20398 gnd.n6776 gnd.n638 0.152939
R20399 gnd.n6784 gnd.n638 0.152939
R20400 gnd.n6785 gnd.n6784 0.152939
R20401 gnd.n6786 gnd.n6785 0.152939
R20402 gnd.n6786 gnd.n632 0.152939
R20403 gnd.n6794 gnd.n632 0.152939
R20404 gnd.n6795 gnd.n6794 0.152939
R20405 gnd.n6796 gnd.n6795 0.152939
R20406 gnd.n6796 gnd.n626 0.152939
R20407 gnd.n6804 gnd.n626 0.152939
R20408 gnd.n6805 gnd.n6804 0.152939
R20409 gnd.n6806 gnd.n6805 0.152939
R20410 gnd.n6806 gnd.n620 0.152939
R20411 gnd.n6814 gnd.n620 0.152939
R20412 gnd.n6815 gnd.n6814 0.152939
R20413 gnd.n6816 gnd.n6815 0.152939
R20414 gnd.n6816 gnd.n614 0.152939
R20415 gnd.n6824 gnd.n614 0.152939
R20416 gnd.n6825 gnd.n6824 0.152939
R20417 gnd.n6826 gnd.n6825 0.152939
R20418 gnd.n6826 gnd.n608 0.152939
R20419 gnd.n6834 gnd.n608 0.152939
R20420 gnd.n6835 gnd.n6834 0.152939
R20421 gnd.n6836 gnd.n6835 0.152939
R20422 gnd.n6836 gnd.n602 0.152939
R20423 gnd.n6844 gnd.n602 0.152939
R20424 gnd.n6845 gnd.n6844 0.152939
R20425 gnd.n6846 gnd.n6845 0.152939
R20426 gnd.n6846 gnd.n596 0.152939
R20427 gnd.n6854 gnd.n596 0.152939
R20428 gnd.n6855 gnd.n6854 0.152939
R20429 gnd.n6856 gnd.n6855 0.152939
R20430 gnd.n6856 gnd.n590 0.152939
R20431 gnd.n6864 gnd.n590 0.152939
R20432 gnd.n6865 gnd.n6864 0.152939
R20433 gnd.n6866 gnd.n6865 0.152939
R20434 gnd.n6866 gnd.n584 0.152939
R20435 gnd.n6874 gnd.n584 0.152939
R20436 gnd.n6875 gnd.n6874 0.152939
R20437 gnd.n6876 gnd.n6875 0.152939
R20438 gnd.n6876 gnd.n578 0.152939
R20439 gnd.n6884 gnd.n578 0.152939
R20440 gnd.n6885 gnd.n6884 0.152939
R20441 gnd.n6886 gnd.n6885 0.152939
R20442 gnd.n6886 gnd.n572 0.152939
R20443 gnd.n6894 gnd.n572 0.152939
R20444 gnd.n6895 gnd.n6894 0.152939
R20445 gnd.n6896 gnd.n6895 0.152939
R20446 gnd.n6896 gnd.n566 0.152939
R20447 gnd.n6904 gnd.n566 0.152939
R20448 gnd.n6905 gnd.n6904 0.152939
R20449 gnd.n6906 gnd.n6905 0.152939
R20450 gnd.n6906 gnd.n560 0.152939
R20451 gnd.n6914 gnd.n560 0.152939
R20452 gnd.n6915 gnd.n6914 0.152939
R20453 gnd.n6916 gnd.n6915 0.152939
R20454 gnd.n6916 gnd.n554 0.152939
R20455 gnd.n6924 gnd.n554 0.152939
R20456 gnd.n6925 gnd.n6924 0.152939
R20457 gnd.n6927 gnd.n6925 0.152939
R20458 gnd.n6927 gnd.n6926 0.152939
R20459 gnd.n6926 gnd.n548 0.152939
R20460 gnd.n6936 gnd.n548 0.152939
R20461 gnd.n6937 gnd.n543 0.152939
R20462 gnd.n6945 gnd.n543 0.152939
R20463 gnd.n6946 gnd.n6945 0.152939
R20464 gnd.n6947 gnd.n6946 0.152939
R20465 gnd.n6947 gnd.n537 0.152939
R20466 gnd.n6955 gnd.n537 0.152939
R20467 gnd.n6956 gnd.n6955 0.152939
R20468 gnd.n6957 gnd.n6956 0.152939
R20469 gnd.n6957 gnd.n531 0.152939
R20470 gnd.n6965 gnd.n531 0.152939
R20471 gnd.n6966 gnd.n6965 0.152939
R20472 gnd.n6967 gnd.n6966 0.152939
R20473 gnd.n6967 gnd.n525 0.152939
R20474 gnd.n6975 gnd.n525 0.152939
R20475 gnd.n6976 gnd.n6975 0.152939
R20476 gnd.n6977 gnd.n6976 0.152939
R20477 gnd.n6977 gnd.n519 0.152939
R20478 gnd.n6985 gnd.n519 0.152939
R20479 gnd.n6986 gnd.n6985 0.152939
R20480 gnd.n6987 gnd.n6986 0.152939
R20481 gnd.n6987 gnd.n513 0.152939
R20482 gnd.n6995 gnd.n513 0.152939
R20483 gnd.n6996 gnd.n6995 0.152939
R20484 gnd.n6997 gnd.n6996 0.152939
R20485 gnd.n6997 gnd.n507 0.152939
R20486 gnd.n7005 gnd.n507 0.152939
R20487 gnd.n7006 gnd.n7005 0.152939
R20488 gnd.n7007 gnd.n7006 0.152939
R20489 gnd.n7007 gnd.n501 0.152939
R20490 gnd.n7015 gnd.n501 0.152939
R20491 gnd.n7016 gnd.n7015 0.152939
R20492 gnd.n7017 gnd.n7016 0.152939
R20493 gnd.n7017 gnd.n495 0.152939
R20494 gnd.n7025 gnd.n495 0.152939
R20495 gnd.n7026 gnd.n7025 0.152939
R20496 gnd.n7027 gnd.n7026 0.152939
R20497 gnd.n7027 gnd.n489 0.152939
R20498 gnd.n7035 gnd.n489 0.152939
R20499 gnd.n7036 gnd.n7035 0.152939
R20500 gnd.n7037 gnd.n7036 0.152939
R20501 gnd.n7037 gnd.n483 0.152939
R20502 gnd.n7045 gnd.n483 0.152939
R20503 gnd.n7046 gnd.n7045 0.152939
R20504 gnd.n7047 gnd.n7046 0.152939
R20505 gnd.n7047 gnd.n477 0.152939
R20506 gnd.n7055 gnd.n477 0.152939
R20507 gnd.n7056 gnd.n7055 0.152939
R20508 gnd.n7057 gnd.n7056 0.152939
R20509 gnd.n7057 gnd.n471 0.152939
R20510 gnd.n7065 gnd.n471 0.152939
R20511 gnd.n7066 gnd.n7065 0.152939
R20512 gnd.n7067 gnd.n7066 0.152939
R20513 gnd.n7067 gnd.n465 0.152939
R20514 gnd.n7075 gnd.n465 0.152939
R20515 gnd.n7076 gnd.n7075 0.152939
R20516 gnd.n7077 gnd.n7076 0.152939
R20517 gnd.n7077 gnd.n459 0.152939
R20518 gnd.n7085 gnd.n459 0.152939
R20519 gnd.n7086 gnd.n7085 0.152939
R20520 gnd.n7087 gnd.n7086 0.152939
R20521 gnd.n7087 gnd.n453 0.152939
R20522 gnd.n7095 gnd.n453 0.152939
R20523 gnd.n7096 gnd.n7095 0.152939
R20524 gnd.n7097 gnd.n7096 0.152939
R20525 gnd.n7097 gnd.n447 0.152939
R20526 gnd.n7105 gnd.n447 0.152939
R20527 gnd.n7106 gnd.n7105 0.152939
R20528 gnd.n7107 gnd.n7106 0.152939
R20529 gnd.n7107 gnd.n441 0.152939
R20530 gnd.n7115 gnd.n441 0.152939
R20531 gnd.n7116 gnd.n7115 0.152939
R20532 gnd.n7117 gnd.n7116 0.152939
R20533 gnd.n7117 gnd.n435 0.152939
R20534 gnd.n7125 gnd.n435 0.152939
R20535 gnd.n7126 gnd.n7125 0.152939
R20536 gnd.n7127 gnd.n7126 0.152939
R20537 gnd.n7127 gnd.n429 0.152939
R20538 gnd.n7135 gnd.n429 0.152939
R20539 gnd.n7136 gnd.n7135 0.152939
R20540 gnd.n7137 gnd.n7136 0.152939
R20541 gnd.n7137 gnd.n423 0.152939
R20542 gnd.n7146 gnd.n423 0.152939
R20543 gnd.n7147 gnd.n7146 0.152939
R20544 gnd.n7148 gnd.n7147 0.152939
R20545 gnd.n7355 gnd.n7354 0.152939
R20546 gnd.n7355 gnd.n287 0.152939
R20547 gnd.n7369 gnd.n287 0.152939
R20548 gnd.n7370 gnd.n7369 0.152939
R20549 gnd.n7371 gnd.n7370 0.152939
R20550 gnd.n7371 gnd.n273 0.152939
R20551 gnd.n7385 gnd.n273 0.152939
R20552 gnd.n7386 gnd.n7385 0.152939
R20553 gnd.n7387 gnd.n7386 0.152939
R20554 gnd.n7387 gnd.n257 0.152939
R20555 gnd.n7401 gnd.n257 0.152939
R20556 gnd.n7402 gnd.n7401 0.152939
R20557 gnd.n7403 gnd.n7402 0.152939
R20558 gnd.n7403 gnd.n242 0.152939
R20559 gnd.n7417 gnd.n242 0.152939
R20560 gnd.n7418 gnd.n7417 0.152939
R20561 gnd.n7419 gnd.n7418 0.152939
R20562 gnd.n7419 gnd.n226 0.152939
R20563 gnd.n7433 gnd.n226 0.152939
R20564 gnd.n7434 gnd.n7433 0.152939
R20565 gnd.n7435 gnd.n7434 0.152939
R20566 gnd.n7435 gnd.n210 0.152939
R20567 gnd.n7517 gnd.n210 0.152939
R20568 gnd.n7518 gnd.n7517 0.152939
R20569 gnd.n7519 gnd.n7518 0.152939
R20570 gnd.n7519 gnd.n133 0.152939
R20571 gnd.n7599 gnd.n133 0.152939
R20572 gnd.n7598 gnd.n134 0.152939
R20573 gnd.n136 gnd.n134 0.152939
R20574 gnd.n140 gnd.n136 0.152939
R20575 gnd.n141 gnd.n140 0.152939
R20576 gnd.n142 gnd.n141 0.152939
R20577 gnd.n143 gnd.n142 0.152939
R20578 gnd.n147 gnd.n143 0.152939
R20579 gnd.n148 gnd.n147 0.152939
R20580 gnd.n149 gnd.n148 0.152939
R20581 gnd.n150 gnd.n149 0.152939
R20582 gnd.n154 gnd.n150 0.152939
R20583 gnd.n155 gnd.n154 0.152939
R20584 gnd.n156 gnd.n155 0.152939
R20585 gnd.n157 gnd.n156 0.152939
R20586 gnd.n161 gnd.n157 0.152939
R20587 gnd.n162 gnd.n161 0.152939
R20588 gnd.n163 gnd.n162 0.152939
R20589 gnd.n164 gnd.n163 0.152939
R20590 gnd.n168 gnd.n164 0.152939
R20591 gnd.n169 gnd.n168 0.152939
R20592 gnd.n170 gnd.n169 0.152939
R20593 gnd.n171 gnd.n170 0.152939
R20594 gnd.n175 gnd.n171 0.152939
R20595 gnd.n176 gnd.n175 0.152939
R20596 gnd.n177 gnd.n176 0.152939
R20597 gnd.n178 gnd.n177 0.152939
R20598 gnd.n182 gnd.n178 0.152939
R20599 gnd.n183 gnd.n182 0.152939
R20600 gnd.n184 gnd.n183 0.152939
R20601 gnd.n185 gnd.n184 0.152939
R20602 gnd.n189 gnd.n185 0.152939
R20603 gnd.n190 gnd.n189 0.152939
R20604 gnd.n191 gnd.n190 0.152939
R20605 gnd.n192 gnd.n191 0.152939
R20606 gnd.n196 gnd.n192 0.152939
R20607 gnd.n197 gnd.n196 0.152939
R20608 gnd.n7529 gnd.n197 0.152939
R20609 gnd.n7529 gnd.n7528 0.152939
R20610 gnd.n1456 gnd.n1333 0.152939
R20611 gnd.n1457 gnd.n1456 0.152939
R20612 gnd.n1458 gnd.n1457 0.152939
R20613 gnd.n1459 gnd.n1458 0.152939
R20614 gnd.n1460 gnd.n1459 0.152939
R20615 gnd.n1461 gnd.n1460 0.152939
R20616 gnd.n1462 gnd.n1461 0.152939
R20617 gnd.n1463 gnd.n1462 0.152939
R20618 gnd.n1464 gnd.n1463 0.152939
R20619 gnd.n1464 gnd.n1390 0.152939
R20620 gnd.n5922 gnd.n1390 0.152939
R20621 gnd.n5923 gnd.n5922 0.152939
R20622 gnd.n5924 gnd.n5923 0.152939
R20623 gnd.n5924 gnd.n1388 0.152939
R20624 gnd.n5929 gnd.n1388 0.152939
R20625 gnd.n5930 gnd.n5929 0.152939
R20626 gnd.n5931 gnd.n5930 0.152939
R20627 gnd.n5932 gnd.n5931 0.152939
R20628 gnd.n5932 gnd.n387 0.152939
R20629 gnd.n7185 gnd.n387 0.152939
R20630 gnd.n7186 gnd.n7185 0.152939
R20631 gnd.n7187 gnd.n7186 0.152939
R20632 gnd.n7188 gnd.n7187 0.152939
R20633 gnd.n7189 gnd.n7188 0.152939
R20634 gnd.n7189 gnd.n353 0.152939
R20635 gnd.n7230 gnd.n353 0.152939
R20636 gnd.n7231 gnd.n7230 0.152939
R20637 gnd.n7232 gnd.n7231 0.152939
R20638 gnd.n7233 gnd.n7232 0.152939
R20639 gnd.n7234 gnd.n7233 0.152939
R20640 gnd.n7235 gnd.n7234 0.152939
R20641 gnd.n7235 gnd.n337 0.152939
R20642 gnd.n7260 gnd.n337 0.152939
R20643 gnd.n7261 gnd.n7260 0.152939
R20644 gnd.n7262 gnd.n7261 0.152939
R20645 gnd.n7263 gnd.n7262 0.152939
R20646 gnd.n7264 gnd.n7263 0.152939
R20647 gnd.n7265 gnd.n7264 0.152939
R20648 gnd.n7266 gnd.n7265 0.152939
R20649 gnd.n7267 gnd.n7266 0.152939
R20650 gnd.n7268 gnd.n7267 0.152939
R20651 gnd.n7269 gnd.n7268 0.152939
R20652 gnd.n7270 gnd.n7269 0.152939
R20653 gnd.n7271 gnd.n7270 0.152939
R20654 gnd.n7272 gnd.n7271 0.152939
R20655 gnd.n7273 gnd.n7272 0.152939
R20656 gnd.n7274 gnd.n7273 0.152939
R20657 gnd.n7275 gnd.n7274 0.152939
R20658 gnd.n7276 gnd.n7275 0.152939
R20659 gnd.n7277 gnd.n7276 0.152939
R20660 gnd.n7278 gnd.n7277 0.152939
R20661 gnd.n7279 gnd.n7278 0.152939
R20662 gnd.n7280 gnd.n7279 0.152939
R20663 gnd.n7281 gnd.n7280 0.152939
R20664 gnd.n7282 gnd.n7281 0.152939
R20665 gnd.n7283 gnd.n7282 0.152939
R20666 gnd.n7284 gnd.n7283 0.152939
R20667 gnd.n7285 gnd.n7284 0.152939
R20668 gnd.n7286 gnd.n7285 0.152939
R20669 gnd.n7287 gnd.n7286 0.152939
R20670 gnd.n7289 gnd.n7287 0.152939
R20671 gnd.n7289 gnd.n7288 0.152939
R20672 gnd.n7288 gnd.n203 0.152939
R20673 gnd.n7527 gnd.n203 0.152939
R20674 gnd.n1290 gnd.n1289 0.152939
R20675 gnd.n1291 gnd.n1290 0.152939
R20676 gnd.n1292 gnd.n1291 0.152939
R20677 gnd.n1293 gnd.n1292 0.152939
R20678 gnd.n1294 gnd.n1293 0.152939
R20679 gnd.n1295 gnd.n1294 0.152939
R20680 gnd.n1296 gnd.n1295 0.152939
R20681 gnd.n1297 gnd.n1296 0.152939
R20682 gnd.n1298 gnd.n1297 0.152939
R20683 gnd.n1299 gnd.n1298 0.152939
R20684 gnd.n1300 gnd.n1299 0.152939
R20685 gnd.n1301 gnd.n1300 0.152939
R20686 gnd.n1302 gnd.n1301 0.152939
R20687 gnd.n1303 gnd.n1302 0.152939
R20688 gnd.n1304 gnd.n1303 0.152939
R20689 gnd.n1311 gnd.n1310 0.152939
R20690 gnd.n1312 gnd.n1311 0.152939
R20691 gnd.n1313 gnd.n1312 0.152939
R20692 gnd.n1314 gnd.n1313 0.152939
R20693 gnd.n1315 gnd.n1314 0.152939
R20694 gnd.n1316 gnd.n1315 0.152939
R20695 gnd.n1317 gnd.n1316 0.152939
R20696 gnd.n1318 gnd.n1317 0.152939
R20697 gnd.n1319 gnd.n1318 0.152939
R20698 gnd.n1320 gnd.n1319 0.152939
R20699 gnd.n1321 gnd.n1320 0.152939
R20700 gnd.n1322 gnd.n1321 0.152939
R20701 gnd.n1323 gnd.n1322 0.152939
R20702 gnd.n1324 gnd.n1323 0.152939
R20703 gnd.n1325 gnd.n1324 0.152939
R20704 gnd.n1326 gnd.n1325 0.152939
R20705 gnd.n1327 gnd.n1326 0.152939
R20706 gnd.n6022 gnd.n1327 0.152939
R20707 gnd.n6022 gnd.n6021 0.152939
R20708 gnd.n6021 gnd.n6020 0.152939
R20709 gnd.n5846 gnd.n5845 0.152939
R20710 gnd.n5847 gnd.n5846 0.152939
R20711 gnd.n5847 gnd.n1428 0.152939
R20712 gnd.n5875 gnd.n1428 0.152939
R20713 gnd.n5876 gnd.n5875 0.152939
R20714 gnd.n5877 gnd.n5876 0.152939
R20715 gnd.n5878 gnd.n5877 0.152939
R20716 gnd.n5878 gnd.n1401 0.152939
R20717 gnd.n5912 gnd.n1401 0.152939
R20718 gnd.n5913 gnd.n5912 0.152939
R20719 gnd.n5914 gnd.n5913 0.152939
R20720 gnd.n5915 gnd.n5914 0.152939
R20721 gnd.n5915 gnd.n1367 0.152939
R20722 gnd.n5982 gnd.n1367 0.152939
R20723 gnd.n5983 gnd.n5982 0.152939
R20724 gnd.n5984 gnd.n5983 0.152939
R20725 gnd.n5984 gnd.n396 0.152939
R20726 gnd.n7175 gnd.n396 0.152939
R20727 gnd.n7176 gnd.n7175 0.152939
R20728 gnd.n7177 gnd.n7176 0.152939
R20729 gnd.n7178 gnd.n7177 0.152939
R20730 gnd.n7178 gnd.n363 0.152939
R20731 gnd.n7221 gnd.n363 0.152939
R20732 gnd.n7222 gnd.n7221 0.152939
R20733 gnd.n7223 gnd.n7222 0.152939
R20734 gnd.n7223 gnd.n303 0.152939
R20735 gnd.n7354 gnd.n303 0.152939
R20736 gnd.n6343 gnd.n967 0.152939
R20737 gnd.n4356 gnd.n967 0.152939
R20738 gnd.n4357 gnd.n4356 0.152939
R20739 gnd.n4358 gnd.n4357 0.152939
R20740 gnd.n4358 gnd.n2149 0.152939
R20741 gnd.n4397 gnd.n2149 0.152939
R20742 gnd.n4398 gnd.n4397 0.152939
R20743 gnd.n4399 gnd.n4398 0.152939
R20744 gnd.n4399 gnd.n2145 0.152939
R20745 gnd.n4405 gnd.n2145 0.152939
R20746 gnd.n4406 gnd.n4405 0.152939
R20747 gnd.n4407 gnd.n4406 0.152939
R20748 gnd.n4407 gnd.n2128 0.152939
R20749 gnd.n4446 gnd.n2128 0.152939
R20750 gnd.n4447 gnd.n4446 0.152939
R20751 gnd.n4448 gnd.n4447 0.152939
R20752 gnd.n4448 gnd.n2124 0.152939
R20753 gnd.n4454 gnd.n2124 0.152939
R20754 gnd.n4455 gnd.n4454 0.152939
R20755 gnd.n4456 gnd.n4455 0.152939
R20756 gnd.n4457 gnd.n4456 0.152939
R20757 gnd.n4458 gnd.n4457 0.152939
R20758 gnd.n4461 gnd.n4458 0.152939
R20759 gnd.n4462 gnd.n4461 0.152939
R20760 gnd.n4463 gnd.n4462 0.152939
R20761 gnd.n4464 gnd.n4463 0.152939
R20762 gnd.n4467 gnd.n4464 0.152939
R20763 gnd.n4468 gnd.n4467 0.152939
R20764 gnd.n4469 gnd.n4468 0.152939
R20765 gnd.n4470 gnd.n4469 0.152939
R20766 gnd.n4472 gnd.n4470 0.152939
R20767 gnd.n4473 gnd.n4472 0.152939
R20768 gnd.n4473 gnd.n1949 0.152939
R20769 gnd.n5416 gnd.n1949 0.152939
R20770 gnd.n5417 gnd.n5416 0.152939
R20771 gnd.n5418 gnd.n5417 0.152939
R20772 gnd.n5418 gnd.n1935 0.152939
R20773 gnd.n5432 gnd.n1935 0.152939
R20774 gnd.n5433 gnd.n5432 0.152939
R20775 gnd.n5434 gnd.n5433 0.152939
R20776 gnd.n5434 gnd.n1923 0.152939
R20777 gnd.n5448 gnd.n1923 0.152939
R20778 gnd.n5449 gnd.n5448 0.152939
R20779 gnd.n5450 gnd.n5449 0.152939
R20780 gnd.n5450 gnd.n1910 0.152939
R20781 gnd.n5464 gnd.n1910 0.152939
R20782 gnd.n5465 gnd.n5464 0.152939
R20783 gnd.n5466 gnd.n5465 0.152939
R20784 gnd.n5466 gnd.n1897 0.152939
R20785 gnd.n5480 gnd.n1897 0.152939
R20786 gnd.n5481 gnd.n5480 0.152939
R20787 gnd.n5482 gnd.n5481 0.152939
R20788 gnd.n5482 gnd.n1884 0.152939
R20789 gnd.n5496 gnd.n1884 0.152939
R20790 gnd.n5497 gnd.n5496 0.152939
R20791 gnd.n5498 gnd.n5497 0.152939
R20792 gnd.n5498 gnd.n1871 0.152939
R20793 gnd.n5512 gnd.n1871 0.152939
R20794 gnd.n5513 gnd.n5512 0.152939
R20795 gnd.n5514 gnd.n5513 0.152939
R20796 gnd.n5514 gnd.n1856 0.152939
R20797 gnd.n5528 gnd.n1856 0.152939
R20798 gnd.n5529 gnd.n5528 0.152939
R20799 gnd.n5530 gnd.n5529 0.152939
R20800 gnd.n5530 gnd.n1843 0.152939
R20801 gnd.n5544 gnd.n1843 0.152939
R20802 gnd.n5545 gnd.n5544 0.152939
R20803 gnd.n5546 gnd.n5545 0.152939
R20804 gnd.n5546 gnd.n1830 0.152939
R20805 gnd.n5560 gnd.n1830 0.152939
R20806 gnd.n5561 gnd.n5560 0.152939
R20807 gnd.n5562 gnd.n5561 0.152939
R20808 gnd.n5562 gnd.n1815 0.152939
R20809 gnd.n5576 gnd.n1815 0.152939
R20810 gnd.n5577 gnd.n5576 0.152939
R20811 gnd.n5578 gnd.n5577 0.152939
R20812 gnd.n5578 gnd.n1800 0.152939
R20813 gnd.n5592 gnd.n1800 0.152939
R20814 gnd.n5593 gnd.n5592 0.152939
R20815 gnd.n5594 gnd.n5593 0.152939
R20816 gnd.n5594 gnd.n1787 0.152939
R20817 gnd.n5608 gnd.n1787 0.152939
R20818 gnd.n5609 gnd.n5608 0.152939
R20819 gnd.n5610 gnd.n5609 0.152939
R20820 gnd.n5610 gnd.n1773 0.152939
R20821 gnd.n5624 gnd.n1773 0.152939
R20822 gnd.n5625 gnd.n5624 0.152939
R20823 gnd.n5626 gnd.n5625 0.152939
R20824 gnd.n5626 gnd.n1758 0.152939
R20825 gnd.n5640 gnd.n1758 0.152939
R20826 gnd.n5641 gnd.n5640 0.152939
R20827 gnd.n5642 gnd.n5641 0.152939
R20828 gnd.n5642 gnd.n1745 0.152939
R20829 gnd.n5656 gnd.n1745 0.152939
R20830 gnd.n5657 gnd.n5656 0.152939
R20831 gnd.n5658 gnd.n5657 0.152939
R20832 gnd.n5658 gnd.n1730 0.152939
R20833 gnd.n5672 gnd.n1730 0.152939
R20834 gnd.n5673 gnd.n5672 0.152939
R20835 gnd.n5674 gnd.n5673 0.152939
R20836 gnd.n5674 gnd.n1717 0.152939
R20837 gnd.n5688 gnd.n1717 0.152939
R20838 gnd.n5689 gnd.n5688 0.152939
R20839 gnd.n5690 gnd.n5689 0.152939
R20840 gnd.n5690 gnd.n1703 0.152939
R20841 gnd.n5704 gnd.n1703 0.152939
R20842 gnd.n5705 gnd.n5704 0.152939
R20843 gnd.n5706 gnd.n5705 0.152939
R20844 gnd.n5706 gnd.n1689 0.152939
R20845 gnd.n5720 gnd.n1689 0.152939
R20846 gnd.n5721 gnd.n5720 0.152939
R20847 gnd.n5722 gnd.n5721 0.152939
R20848 gnd.n5722 gnd.n1676 0.152939
R20849 gnd.n5736 gnd.n1676 0.152939
R20850 gnd.n5737 gnd.n5736 0.152939
R20851 gnd.n5738 gnd.n5737 0.152939
R20852 gnd.n5738 gnd.n1663 0.152939
R20853 gnd.n5752 gnd.n1663 0.152939
R20854 gnd.n5753 gnd.n5752 0.152939
R20855 gnd.n5754 gnd.n5753 0.152939
R20856 gnd.n5754 gnd.n1650 0.152939
R20857 gnd.n5768 gnd.n1650 0.152939
R20858 gnd.n5769 gnd.n5768 0.152939
R20859 gnd.n5770 gnd.n5769 0.152939
R20860 gnd.n5770 gnd.n1636 0.152939
R20861 gnd.n5784 gnd.n1636 0.152939
R20862 gnd.n5785 gnd.n5784 0.152939
R20863 gnd.n5786 gnd.n5785 0.152939
R20864 gnd.n5786 gnd.n1623 0.152939
R20865 gnd.n5802 gnd.n1623 0.152939
R20866 gnd.n5803 gnd.n5802 0.152939
R20867 gnd.n5804 gnd.n5803 0.152939
R20868 gnd.n5806 gnd.n5804 0.152939
R20869 gnd.n5806 gnd.n5805 0.152939
R20870 gnd.n5805 gnd.n1251 0.152939
R20871 gnd.n1252 gnd.n1251 0.152939
R20872 gnd.n1253 gnd.n1252 0.152939
R20873 gnd.n1443 gnd.n1253 0.152939
R20874 gnd.n1446 gnd.n1443 0.152939
R20875 gnd.n1447 gnd.n1446 0.152939
R20876 gnd.n1448 gnd.n1447 0.152939
R20877 gnd.n1448 gnd.n1439 0.152939
R20878 gnd.n5864 gnd.n1439 0.152939
R20879 gnd.n5865 gnd.n5864 0.152939
R20880 gnd.n5866 gnd.n5865 0.152939
R20881 gnd.n5867 gnd.n5866 0.152939
R20882 gnd.n5867 gnd.n1411 0.152939
R20883 gnd.n5900 gnd.n1411 0.152939
R20884 gnd.n5901 gnd.n5900 0.152939
R20885 gnd.n5902 gnd.n5901 0.152939
R20886 gnd.n5903 gnd.n5902 0.152939
R20887 gnd.n5903 gnd.n1377 0.152939
R20888 gnd.n5961 gnd.n1377 0.152939
R20889 gnd.n5962 gnd.n5961 0.152939
R20890 gnd.n5963 gnd.n5962 0.152939
R20891 gnd.n5964 gnd.n5963 0.152939
R20892 gnd.n5965 gnd.n5964 0.152939
R20893 gnd.n5967 gnd.n5965 0.152939
R20894 gnd.n5969 gnd.n5967 0.152939
R20895 gnd.n5969 gnd.n5968 0.152939
R20896 gnd.n5968 gnd.n412 0.152939
R20897 gnd.n413 gnd.n412 0.152939
R20898 gnd.n414 gnd.n413 0.152939
R20899 gnd.n417 gnd.n414 0.152939
R20900 gnd.n418 gnd.n417 0.152939
R20901 gnd.n419 gnd.n418 0.152939
R20902 gnd.n420 gnd.n419 0.152939
R20903 gnd.n3864 gnd.n3863 0.152939
R20904 gnd.n3865 gnd.n3864 0.152939
R20905 gnd.n3866 gnd.n3865 0.152939
R20906 gnd.n3867 gnd.n3866 0.152939
R20907 gnd.n3868 gnd.n3867 0.152939
R20908 gnd.n3869 gnd.n3868 0.152939
R20909 gnd.n3870 gnd.n3869 0.152939
R20910 gnd.n3871 gnd.n3870 0.152939
R20911 gnd.n3872 gnd.n3871 0.152939
R20912 gnd.n3873 gnd.n3872 0.152939
R20913 gnd.n3874 gnd.n3873 0.152939
R20914 gnd.n3875 gnd.n3874 0.152939
R20915 gnd.n3876 gnd.n3875 0.152939
R20916 gnd.n3877 gnd.n3876 0.152939
R20917 gnd.n3878 gnd.n3877 0.152939
R20918 gnd.n3879 gnd.n3878 0.152939
R20919 gnd.n3880 gnd.n3879 0.152939
R20920 gnd.n3881 gnd.n3880 0.152939
R20921 gnd.n3882 gnd.n3881 0.152939
R20922 gnd.n3883 gnd.n3882 0.152939
R20923 gnd.n3884 gnd.n3883 0.152939
R20924 gnd.n3885 gnd.n3884 0.152939
R20925 gnd.n3886 gnd.n3885 0.152939
R20926 gnd.n3887 gnd.n3886 0.152939
R20927 gnd.n3888 gnd.n3887 0.152939
R20928 gnd.n3889 gnd.n3888 0.152939
R20929 gnd.n3890 gnd.n3889 0.152939
R20930 gnd.n3891 gnd.n3890 0.152939
R20931 gnd.n3892 gnd.n3891 0.152939
R20932 gnd.n3893 gnd.n3892 0.152939
R20933 gnd.n3894 gnd.n3893 0.152939
R20934 gnd.n3815 gnd.n2317 0.152939
R20935 gnd.n3823 gnd.n3815 0.152939
R20936 gnd.n3824 gnd.n3823 0.152939
R20937 gnd.n3825 gnd.n3824 0.152939
R20938 gnd.n3825 gnd.n3811 0.152939
R20939 gnd.n3833 gnd.n3811 0.152939
R20940 gnd.n3834 gnd.n3833 0.152939
R20941 gnd.n3835 gnd.n3834 0.152939
R20942 gnd.n3835 gnd.n3807 0.152939
R20943 gnd.n3843 gnd.n3807 0.152939
R20944 gnd.n3844 gnd.n3843 0.152939
R20945 gnd.n3845 gnd.n3844 0.152939
R20946 gnd.n3845 gnd.n3803 0.152939
R20947 gnd.n3853 gnd.n3803 0.152939
R20948 gnd.n3854 gnd.n3853 0.152939
R20949 gnd.n3855 gnd.n3854 0.152939
R20950 gnd.n3855 gnd.n3797 0.152939
R20951 gnd.n3862 gnd.n3797 0.152939
R20952 gnd.n4183 gnd.n4182 0.152939
R20953 gnd.n4184 gnd.n4183 0.152939
R20954 gnd.n4184 gnd.n2302 0.152939
R20955 gnd.n4198 gnd.n2302 0.152939
R20956 gnd.n4199 gnd.n4198 0.152939
R20957 gnd.n4200 gnd.n4199 0.152939
R20958 gnd.n4200 gnd.n2285 0.152939
R20959 gnd.n4214 gnd.n2285 0.152939
R20960 gnd.n4215 gnd.n4214 0.152939
R20961 gnd.n4216 gnd.n4215 0.152939
R20962 gnd.n4216 gnd.n2270 0.152939
R20963 gnd.n4230 gnd.n2270 0.152939
R20964 gnd.n4231 gnd.n4230 0.152939
R20965 gnd.n4232 gnd.n4231 0.152939
R20966 gnd.n4232 gnd.n2253 0.152939
R20967 gnd.n4246 gnd.n2253 0.152939
R20968 gnd.n4247 gnd.n4246 0.152939
R20969 gnd.n4248 gnd.n4247 0.152939
R20970 gnd.n4248 gnd.n2238 0.152939
R20971 gnd.n4262 gnd.n2238 0.152939
R20972 gnd.n4263 gnd.n4262 0.152939
R20973 gnd.n4264 gnd.n4263 0.152939
R20974 gnd.n4264 gnd.n2221 0.152939
R20975 gnd.n4279 gnd.n2221 0.152939
R20976 gnd.n4280 gnd.n4279 0.152939
R20977 gnd.n4281 gnd.n4280 0.152939
R20978 gnd.n4281 gnd.n2207 0.152939
R20979 gnd.n4295 gnd.n2207 0.152939
R20980 gnd.n4296 gnd.n4295 0.152939
R20981 gnd.n4297 gnd.n4296 0.152939
R20982 gnd.n4297 gnd.n2182 0.152939
R20983 gnd.n4313 gnd.n2182 0.152939
R20984 gnd.n4314 gnd.n4313 0.152939
R20985 gnd.n4315 gnd.n4314 0.152939
R20986 gnd.n4316 gnd.n4315 0.152939
R20987 gnd.n4317 gnd.n4316 0.152939
R20988 gnd.n4318 gnd.n4317 0.152939
R20989 gnd.n4320 gnd.n4318 0.152939
R20990 gnd.n4320 gnd.n4319 0.152939
R20991 gnd.n4319 gnd.n990 0.152939
R20992 gnd.n991 gnd.n990 0.152939
R20993 gnd.n992 gnd.n991 0.152939
R20994 gnd.n1009 gnd.n992 0.152939
R20995 gnd.n1010 gnd.n1009 0.152939
R20996 gnd.n1011 gnd.n1010 0.152939
R20997 gnd.n1012 gnd.n1011 0.152939
R20998 gnd.n1031 gnd.n1012 0.152939
R20999 gnd.n1032 gnd.n1031 0.152939
R21000 gnd.n1033 gnd.n1032 0.152939
R21001 gnd.n1034 gnd.n1033 0.152939
R21002 gnd.n1051 gnd.n1034 0.152939
R21003 gnd.n1052 gnd.n1051 0.152939
R21004 gnd.n1053 gnd.n1052 0.152939
R21005 gnd.n1054 gnd.n1053 0.152939
R21006 gnd.n1073 gnd.n1054 0.152939
R21007 gnd.n1074 gnd.n1073 0.152939
R21008 gnd.n1075 gnd.n1074 0.152939
R21009 gnd.n1076 gnd.n1075 0.152939
R21010 gnd.n1094 gnd.n1076 0.152939
R21011 gnd.n1095 gnd.n1094 0.152939
R21012 gnd.n1096 gnd.n1095 0.152939
R21013 gnd.n1097 gnd.n1096 0.152939
R21014 gnd.n1114 gnd.n1097 0.152939
R21015 gnd.n6258 gnd.n1114 0.152939
R21016 gnd.n978 gnd.n966 0.152939
R21017 gnd.n979 gnd.n978 0.152939
R21018 gnd.n980 gnd.n979 0.152939
R21019 gnd.n999 gnd.n980 0.152939
R21020 gnd.n1000 gnd.n999 0.152939
R21021 gnd.n1001 gnd.n1000 0.152939
R21022 gnd.n1002 gnd.n1001 0.152939
R21023 gnd.n1020 gnd.n1002 0.152939
R21024 gnd.n1021 gnd.n1020 0.152939
R21025 gnd.n1022 gnd.n1021 0.152939
R21026 gnd.n1023 gnd.n1022 0.152939
R21027 gnd.n1041 gnd.n1023 0.152939
R21028 gnd.n1042 gnd.n1041 0.152939
R21029 gnd.n1043 gnd.n1042 0.152939
R21030 gnd.n1044 gnd.n1043 0.152939
R21031 gnd.n1062 gnd.n1044 0.152939
R21032 gnd.n1063 gnd.n1062 0.152939
R21033 gnd.n1064 gnd.n1063 0.152939
R21034 gnd.n1065 gnd.n1064 0.152939
R21035 gnd.n1083 gnd.n1065 0.152939
R21036 gnd.n1084 gnd.n1083 0.152939
R21037 gnd.n1085 gnd.n1084 0.152939
R21038 gnd.n1086 gnd.n1085 0.152939
R21039 gnd.n1104 gnd.n1086 0.152939
R21040 gnd.n1105 gnd.n1104 0.152939
R21041 gnd.n1106 gnd.n1105 0.152939
R21042 gnd.n1107 gnd.n1106 0.152939
R21043 gnd.n2067 gnd.n2066 0.152939
R21044 gnd.n2068 gnd.n2067 0.152939
R21045 gnd.n2069 gnd.n2068 0.152939
R21046 gnd.n2070 gnd.n2069 0.152939
R21047 gnd.n2071 gnd.n2070 0.152939
R21048 gnd.n2072 gnd.n2071 0.152939
R21049 gnd.n2073 gnd.n2072 0.152939
R21050 gnd.n2074 gnd.n2073 0.152939
R21051 gnd.n2075 gnd.n2074 0.152939
R21052 gnd.n2076 gnd.n2075 0.152939
R21053 gnd.n2077 gnd.n2076 0.152939
R21054 gnd.n2078 gnd.n2077 0.152939
R21055 gnd.n2079 gnd.n2078 0.152939
R21056 gnd.n2080 gnd.n2079 0.152939
R21057 gnd.n2081 gnd.n2080 0.152939
R21058 gnd.n4600 gnd.n4599 0.152939
R21059 gnd.n4599 gnd.n2086 0.152939
R21060 gnd.n2087 gnd.n2086 0.152939
R21061 gnd.n2088 gnd.n2087 0.152939
R21062 gnd.n2089 gnd.n2088 0.152939
R21063 gnd.n2090 gnd.n2089 0.152939
R21064 gnd.n2091 gnd.n2090 0.152939
R21065 gnd.n2092 gnd.n2091 0.152939
R21066 gnd.n2093 gnd.n2092 0.152939
R21067 gnd.n2094 gnd.n2093 0.152939
R21068 gnd.n2095 gnd.n2094 0.152939
R21069 gnd.n2096 gnd.n2095 0.152939
R21070 gnd.n2097 gnd.n2096 0.152939
R21071 gnd.n2098 gnd.n2097 0.152939
R21072 gnd.n2099 gnd.n2098 0.152939
R21073 gnd.n2100 gnd.n2099 0.152939
R21074 gnd.n2101 gnd.n2100 0.152939
R21075 gnd.n2102 gnd.n2101 0.152939
R21076 gnd.n4559 gnd.n2102 0.152939
R21077 gnd.n4559 gnd.n4558 0.152939
R21078 gnd.n4096 gnd.n4020 0.152939
R21079 gnd.n4022 gnd.n4020 0.152939
R21080 gnd.n4023 gnd.n4022 0.152939
R21081 gnd.n4024 gnd.n4023 0.152939
R21082 gnd.n4025 gnd.n4024 0.152939
R21083 gnd.n4026 gnd.n4025 0.152939
R21084 gnd.n4027 gnd.n4026 0.152939
R21085 gnd.n4028 gnd.n4027 0.152939
R21086 gnd.n4029 gnd.n4028 0.152939
R21087 gnd.n4030 gnd.n4029 0.152939
R21088 gnd.n4031 gnd.n4030 0.152939
R21089 gnd.n4032 gnd.n4031 0.152939
R21090 gnd.n4033 gnd.n4032 0.152939
R21091 gnd.n4034 gnd.n4033 0.152939
R21092 gnd.n4035 gnd.n4034 0.152939
R21093 gnd.n4036 gnd.n4035 0.152939
R21094 gnd.n4037 gnd.n4036 0.152939
R21095 gnd.n4038 gnd.n4037 0.152939
R21096 gnd.n4039 gnd.n4038 0.152939
R21097 gnd.n4040 gnd.n4039 0.152939
R21098 gnd.n4041 gnd.n4040 0.152939
R21099 gnd.n4042 gnd.n4041 0.152939
R21100 gnd.n4043 gnd.n4042 0.152939
R21101 gnd.n4044 gnd.n4043 0.152939
R21102 gnd.n4045 gnd.n4044 0.152939
R21103 gnd.n4046 gnd.n4045 0.152939
R21104 gnd.n4047 gnd.n4046 0.152939
R21105 gnd.n4048 gnd.n4047 0.152939
R21106 gnd.n4049 gnd.n4048 0.152939
R21107 gnd.n4050 gnd.n4049 0.152939
R21108 gnd.n4050 gnd.n2184 0.152939
R21109 gnd.n4312 gnd.n2184 0.152939
R21110 gnd.n4312 gnd.n2185 0.152939
R21111 gnd.n2187 gnd.n2185 0.152939
R21112 gnd.n2188 gnd.n2187 0.152939
R21113 gnd.n2188 gnd.n2167 0.152939
R21114 gnd.n4339 gnd.n2167 0.152939
R21115 gnd.n4340 gnd.n4339 0.152939
R21116 gnd.n4341 gnd.n4340 0.152939
R21117 gnd.n4341 gnd.n2161 0.152939
R21118 gnd.n4365 gnd.n2161 0.152939
R21119 gnd.n4366 gnd.n4365 0.152939
R21120 gnd.n4367 gnd.n4366 0.152939
R21121 gnd.n4367 gnd.n2159 0.152939
R21122 gnd.n4373 gnd.n2159 0.152939
R21123 gnd.n4374 gnd.n4373 0.152939
R21124 gnd.n4375 gnd.n4374 0.152939
R21125 gnd.n4375 gnd.n2140 0.152939
R21126 gnd.n4414 gnd.n2140 0.152939
R21127 gnd.n4415 gnd.n4414 0.152939
R21128 gnd.n4416 gnd.n4415 0.152939
R21129 gnd.n4416 gnd.n2138 0.152939
R21130 gnd.n4422 gnd.n2138 0.152939
R21131 gnd.n4423 gnd.n4422 0.152939
R21132 gnd.n4424 gnd.n4423 0.152939
R21133 gnd.n4425 gnd.n4424 0.152939
R21134 gnd.n4426 gnd.n4425 0.152939
R21135 gnd.n4426 gnd.n2115 0.152939
R21136 gnd.n4507 gnd.n2115 0.152939
R21137 gnd.n4508 gnd.n4507 0.152939
R21138 gnd.n4510 gnd.n4508 0.152939
R21139 gnd.n4510 gnd.n4509 0.152939
R21140 gnd.n4509 gnd.n2107 0.152939
R21141 gnd.n4557 gnd.n2107 0.152939
R21142 gnd.n4175 gnd.n3959 0.152939
R21143 gnd.n3962 gnd.n3959 0.152939
R21144 gnd.n3963 gnd.n3962 0.152939
R21145 gnd.n3964 gnd.n3963 0.152939
R21146 gnd.n3967 gnd.n3964 0.152939
R21147 gnd.n3968 gnd.n3967 0.152939
R21148 gnd.n3969 gnd.n3968 0.152939
R21149 gnd.n3970 gnd.n3969 0.152939
R21150 gnd.n3973 gnd.n3970 0.152939
R21151 gnd.n3974 gnd.n3973 0.152939
R21152 gnd.n3975 gnd.n3974 0.152939
R21153 gnd.n3976 gnd.n3975 0.152939
R21154 gnd.n3979 gnd.n3976 0.152939
R21155 gnd.n3980 gnd.n3979 0.152939
R21156 gnd.n3981 gnd.n3980 0.152939
R21157 gnd.n3982 gnd.n3981 0.152939
R21158 gnd.n3988 gnd.n3982 0.152939
R21159 gnd.n3989 gnd.n3988 0.152939
R21160 gnd.n3990 gnd.n3989 0.152939
R21161 gnd.n3991 gnd.n3990 0.152939
R21162 gnd.n3994 gnd.n3991 0.152939
R21163 gnd.n3995 gnd.n3994 0.152939
R21164 gnd.n3996 gnd.n3995 0.152939
R21165 gnd.n3997 gnd.n3996 0.152939
R21166 gnd.n4000 gnd.n3997 0.152939
R21167 gnd.n4001 gnd.n4000 0.152939
R21168 gnd.n4002 gnd.n4001 0.152939
R21169 gnd.n4003 gnd.n4002 0.152939
R21170 gnd.n4006 gnd.n4003 0.152939
R21171 gnd.n4007 gnd.n4006 0.152939
R21172 gnd.n4008 gnd.n4007 0.152939
R21173 gnd.n4009 gnd.n4008 0.152939
R21174 gnd.n4012 gnd.n4009 0.152939
R21175 gnd.n4013 gnd.n4012 0.152939
R21176 gnd.n4014 gnd.n4013 0.152939
R21177 gnd.n4103 gnd.n4014 0.152939
R21178 gnd.n4103 gnd.n4102 0.152939
R21179 gnd.n4102 gnd.n4101 0.152939
R21180 gnd.n4176 gnd.n2310 0.152939
R21181 gnd.n4190 gnd.n2310 0.152939
R21182 gnd.n4191 gnd.n4190 0.152939
R21183 gnd.n4192 gnd.n4191 0.152939
R21184 gnd.n4192 gnd.n2294 0.152939
R21185 gnd.n4206 gnd.n2294 0.152939
R21186 gnd.n4207 gnd.n4206 0.152939
R21187 gnd.n4208 gnd.n4207 0.152939
R21188 gnd.n4208 gnd.n2278 0.152939
R21189 gnd.n4222 gnd.n2278 0.152939
R21190 gnd.n4223 gnd.n4222 0.152939
R21191 gnd.n4224 gnd.n4223 0.152939
R21192 gnd.n4224 gnd.n2262 0.152939
R21193 gnd.n4238 gnd.n2262 0.152939
R21194 gnd.n4239 gnd.n4238 0.152939
R21195 gnd.n4240 gnd.n4239 0.152939
R21196 gnd.n4240 gnd.n2246 0.152939
R21197 gnd.n4254 gnd.n2246 0.152939
R21198 gnd.n4255 gnd.n4254 0.152939
R21199 gnd.n4256 gnd.n4255 0.152939
R21200 gnd.n4256 gnd.n2230 0.152939
R21201 gnd.n4270 gnd.n2230 0.152939
R21202 gnd.n4271 gnd.n4270 0.152939
R21203 gnd.n4273 gnd.n4271 0.152939
R21204 gnd.n4273 gnd.n4272 0.152939
R21205 gnd.n4272 gnd.n2215 0.152939
R21206 gnd.n2215 gnd.n966 0.152939
R21207 gnd.n6515 gnd.n799 0.152939
R21208 gnd.n804 gnd.n799 0.152939
R21209 gnd.n805 gnd.n804 0.152939
R21210 gnd.n806 gnd.n805 0.152939
R21211 gnd.n807 gnd.n806 0.152939
R21212 gnd.n812 gnd.n807 0.152939
R21213 gnd.n813 gnd.n812 0.152939
R21214 gnd.n814 gnd.n813 0.152939
R21215 gnd.n815 gnd.n814 0.152939
R21216 gnd.n820 gnd.n815 0.152939
R21217 gnd.n821 gnd.n820 0.152939
R21218 gnd.n822 gnd.n821 0.152939
R21219 gnd.n823 gnd.n822 0.152939
R21220 gnd.n828 gnd.n823 0.152939
R21221 gnd.n829 gnd.n828 0.152939
R21222 gnd.n830 gnd.n829 0.152939
R21223 gnd.n831 gnd.n830 0.152939
R21224 gnd.n836 gnd.n831 0.152939
R21225 gnd.n837 gnd.n836 0.152939
R21226 gnd.n838 gnd.n837 0.152939
R21227 gnd.n839 gnd.n838 0.152939
R21228 gnd.n844 gnd.n839 0.152939
R21229 gnd.n845 gnd.n844 0.152939
R21230 gnd.n846 gnd.n845 0.152939
R21231 gnd.n847 gnd.n846 0.152939
R21232 gnd.n852 gnd.n847 0.152939
R21233 gnd.n853 gnd.n852 0.152939
R21234 gnd.n854 gnd.n853 0.152939
R21235 gnd.n855 gnd.n854 0.152939
R21236 gnd.n860 gnd.n855 0.152939
R21237 gnd.n861 gnd.n860 0.152939
R21238 gnd.n862 gnd.n861 0.152939
R21239 gnd.n863 gnd.n862 0.152939
R21240 gnd.n868 gnd.n863 0.152939
R21241 gnd.n869 gnd.n868 0.152939
R21242 gnd.n870 gnd.n869 0.152939
R21243 gnd.n871 gnd.n870 0.152939
R21244 gnd.n876 gnd.n871 0.152939
R21245 gnd.n877 gnd.n876 0.152939
R21246 gnd.n878 gnd.n877 0.152939
R21247 gnd.n879 gnd.n878 0.152939
R21248 gnd.n884 gnd.n879 0.152939
R21249 gnd.n885 gnd.n884 0.152939
R21250 gnd.n886 gnd.n885 0.152939
R21251 gnd.n887 gnd.n886 0.152939
R21252 gnd.n892 gnd.n887 0.152939
R21253 gnd.n893 gnd.n892 0.152939
R21254 gnd.n894 gnd.n893 0.152939
R21255 gnd.n895 gnd.n894 0.152939
R21256 gnd.n900 gnd.n895 0.152939
R21257 gnd.n901 gnd.n900 0.152939
R21258 gnd.n902 gnd.n901 0.152939
R21259 gnd.n903 gnd.n902 0.152939
R21260 gnd.n908 gnd.n903 0.152939
R21261 gnd.n909 gnd.n908 0.152939
R21262 gnd.n910 gnd.n909 0.152939
R21263 gnd.n911 gnd.n910 0.152939
R21264 gnd.n916 gnd.n911 0.152939
R21265 gnd.n917 gnd.n916 0.152939
R21266 gnd.n918 gnd.n917 0.152939
R21267 gnd.n919 gnd.n918 0.152939
R21268 gnd.n924 gnd.n919 0.152939
R21269 gnd.n925 gnd.n924 0.152939
R21270 gnd.n926 gnd.n925 0.152939
R21271 gnd.n927 gnd.n926 0.152939
R21272 gnd.n932 gnd.n927 0.152939
R21273 gnd.n933 gnd.n932 0.152939
R21274 gnd.n934 gnd.n933 0.152939
R21275 gnd.n935 gnd.n934 0.152939
R21276 gnd.n940 gnd.n935 0.152939
R21277 gnd.n941 gnd.n940 0.152939
R21278 gnd.n942 gnd.n941 0.152939
R21279 gnd.n943 gnd.n942 0.152939
R21280 gnd.n948 gnd.n943 0.152939
R21281 gnd.n949 gnd.n948 0.152939
R21282 gnd.n950 gnd.n949 0.152939
R21283 gnd.n951 gnd.n950 0.152939
R21284 gnd.n956 gnd.n951 0.152939
R21285 gnd.n957 gnd.n956 0.152939
R21286 gnd.n958 gnd.n957 0.152939
R21287 gnd.n959 gnd.n958 0.152939
R21288 gnd.n964 gnd.n959 0.152939
R21289 gnd.n965 gnd.n964 0.152939
R21290 gnd.n6345 gnd.n965 0.152939
R21291 gnd.n5838 gnd.n1479 0.152939
R21292 gnd.n5834 gnd.n1479 0.152939
R21293 gnd.n5834 gnd.n5833 0.152939
R21294 gnd.n5833 gnd.n5832 0.152939
R21295 gnd.n5832 gnd.n1607 0.152939
R21296 gnd.n5825 gnd.n1607 0.152939
R21297 gnd.n5825 gnd.n5824 0.152939
R21298 gnd.n5824 gnd.n5823 0.152939
R21299 gnd.n5823 gnd.n5816 0.152939
R21300 gnd.n5410 gnd.n5409 0.152939
R21301 gnd.n5410 gnd.n1942 0.152939
R21302 gnd.n5424 gnd.n1942 0.152939
R21303 gnd.n5425 gnd.n5424 0.152939
R21304 gnd.n5426 gnd.n5425 0.152939
R21305 gnd.n5426 gnd.n1929 0.152939
R21306 gnd.n5440 gnd.n1929 0.152939
R21307 gnd.n5441 gnd.n5440 0.152939
R21308 gnd.n5442 gnd.n5441 0.152939
R21309 gnd.n5442 gnd.n1916 0.152939
R21310 gnd.n5456 gnd.n1916 0.152939
R21311 gnd.n5457 gnd.n5456 0.152939
R21312 gnd.n5458 gnd.n5457 0.152939
R21313 gnd.n5458 gnd.n1903 0.152939
R21314 gnd.n5472 gnd.n1903 0.152939
R21315 gnd.n5473 gnd.n5472 0.152939
R21316 gnd.n5474 gnd.n5473 0.152939
R21317 gnd.n5474 gnd.n1889 0.152939
R21318 gnd.n5488 gnd.n1889 0.152939
R21319 gnd.n5489 gnd.n5488 0.152939
R21320 gnd.n5490 gnd.n5489 0.152939
R21321 gnd.n5490 gnd.n1877 0.152939
R21322 gnd.n5504 gnd.n1877 0.152939
R21323 gnd.n5505 gnd.n5504 0.152939
R21324 gnd.n5506 gnd.n5505 0.152939
R21325 gnd.n5506 gnd.n1863 0.152939
R21326 gnd.n5520 gnd.n1863 0.152939
R21327 gnd.n5521 gnd.n5520 0.152939
R21328 gnd.n5522 gnd.n5521 0.152939
R21329 gnd.n5522 gnd.n1849 0.152939
R21330 gnd.n5536 gnd.n1849 0.152939
R21331 gnd.n5537 gnd.n5536 0.152939
R21332 gnd.n5538 gnd.n5537 0.152939
R21333 gnd.n5538 gnd.n1836 0.152939
R21334 gnd.n5552 gnd.n1836 0.152939
R21335 gnd.n5553 gnd.n5552 0.152939
R21336 gnd.n5554 gnd.n5553 0.152939
R21337 gnd.n5554 gnd.n1823 0.152939
R21338 gnd.n5568 gnd.n1823 0.152939
R21339 gnd.n5569 gnd.n5568 0.152939
R21340 gnd.n5570 gnd.n5569 0.152939
R21341 gnd.n5570 gnd.n1807 0.152939
R21342 gnd.n5584 gnd.n1807 0.152939
R21343 gnd.n5585 gnd.n5584 0.152939
R21344 gnd.n5586 gnd.n5585 0.152939
R21345 gnd.n5586 gnd.n1793 0.152939
R21346 gnd.n5600 gnd.n1793 0.152939
R21347 gnd.n5601 gnd.n5600 0.152939
R21348 gnd.n5602 gnd.n5601 0.152939
R21349 gnd.n5602 gnd.n1779 0.152939
R21350 gnd.n5616 gnd.n1779 0.152939
R21351 gnd.n5617 gnd.n5616 0.152939
R21352 gnd.n5618 gnd.n5617 0.152939
R21353 gnd.n5618 gnd.n1765 0.152939
R21354 gnd.n5632 gnd.n1765 0.152939
R21355 gnd.n5633 gnd.n5632 0.152939
R21356 gnd.n5634 gnd.n5633 0.152939
R21357 gnd.n5634 gnd.n1751 0.152939
R21358 gnd.n5648 gnd.n1751 0.152939
R21359 gnd.n5649 gnd.n5648 0.152939
R21360 gnd.n5650 gnd.n5649 0.152939
R21361 gnd.n5650 gnd.n1737 0.152939
R21362 gnd.n5664 gnd.n1737 0.152939
R21363 gnd.n5665 gnd.n5664 0.152939
R21364 gnd.n5666 gnd.n5665 0.152939
R21365 gnd.n5666 gnd.n1723 0.152939
R21366 gnd.n5680 gnd.n1723 0.152939
R21367 gnd.n5681 gnd.n5680 0.152939
R21368 gnd.n5682 gnd.n5681 0.152939
R21369 gnd.n5682 gnd.n1710 0.152939
R21370 gnd.n5696 gnd.n1710 0.152939
R21371 gnd.n5697 gnd.n5696 0.152939
R21372 gnd.n5698 gnd.n5697 0.152939
R21373 gnd.n5698 gnd.n1695 0.152939
R21374 gnd.n5712 gnd.n1695 0.152939
R21375 gnd.n5713 gnd.n5712 0.152939
R21376 gnd.n5714 gnd.n5713 0.152939
R21377 gnd.n5714 gnd.n1681 0.152939
R21378 gnd.n5728 gnd.n1681 0.152939
R21379 gnd.n5729 gnd.n5728 0.152939
R21380 gnd.n5730 gnd.n5729 0.152939
R21381 gnd.n5730 gnd.n1669 0.152939
R21382 gnd.n5744 gnd.n1669 0.152939
R21383 gnd.n5745 gnd.n5744 0.152939
R21384 gnd.n5746 gnd.n5745 0.152939
R21385 gnd.n5746 gnd.n1656 0.152939
R21386 gnd.n5760 gnd.n1656 0.152939
R21387 gnd.n5761 gnd.n5760 0.152939
R21388 gnd.n5762 gnd.n5761 0.152939
R21389 gnd.n5762 gnd.n1643 0.152939
R21390 gnd.n5776 gnd.n1643 0.152939
R21391 gnd.n5777 gnd.n5776 0.152939
R21392 gnd.n5778 gnd.n5777 0.152939
R21393 gnd.n5778 gnd.n1630 0.152939
R21394 gnd.n5792 gnd.n1630 0.152939
R21395 gnd.n5793 gnd.n5792 0.152939
R21396 gnd.n5796 gnd.n5793 0.152939
R21397 gnd.n5796 gnd.n5795 0.152939
R21398 gnd.n5795 gnd.n5794 0.152939
R21399 gnd.n5794 gnd.n1615 0.152939
R21400 gnd.n5815 gnd.n1615 0.152939
R21401 gnd.n4543 gnd.n4518 0.152939
R21402 gnd.n4543 gnd.n4542 0.152939
R21403 gnd.n4542 gnd.n4541 0.152939
R21404 gnd.n4541 gnd.n4524 0.152939
R21405 gnd.n4537 gnd.n4524 0.152939
R21406 gnd.n4537 gnd.n4536 0.152939
R21407 gnd.n4536 gnd.n4531 0.152939
R21408 gnd.n4531 gnd.n1955 0.152939
R21409 gnd.n5408 gnd.n1955 0.152939
R21410 gnd.n3907 gnd.n3906 0.152939
R21411 gnd.n3906 gnd.n3897 0.152939
R21412 gnd.n3902 gnd.n3897 0.152939
R21413 gnd.n3902 gnd.n3901 0.152939
R21414 gnd.n3901 gnd.n2164 0.152939
R21415 gnd.n4347 gnd.n2164 0.152939
R21416 gnd.n4348 gnd.n4347 0.152939
R21417 gnd.n4349 gnd.n4348 0.152939
R21418 gnd.n4349 gnd.n2155 0.152939
R21419 gnd.n4390 gnd.n2155 0.152939
R21420 gnd.n4390 gnd.n4389 0.152939
R21421 gnd.n4389 gnd.n4388 0.152939
R21422 gnd.n4388 gnd.n2156 0.152939
R21423 gnd.n4384 gnd.n2156 0.152939
R21424 gnd.n4384 gnd.n4383 0.152939
R21425 gnd.n4383 gnd.n4382 0.152939
R21426 gnd.n4382 gnd.n2134 0.152939
R21427 gnd.n4439 gnd.n2134 0.152939
R21428 gnd.n4439 gnd.n4438 0.152939
R21429 gnd.n4438 gnd.n4437 0.152939
R21430 gnd.n4437 gnd.n2135 0.152939
R21431 gnd.n4433 gnd.n2135 0.152939
R21432 gnd.n4433 gnd.n2118 0.152939
R21433 gnd.n4499 gnd.n2118 0.152939
R21434 gnd.n4500 gnd.n4499 0.152939
R21435 gnd.n4501 gnd.n4500 0.152939
R21436 gnd.n4501 gnd.n2112 0.152939
R21437 gnd.n4516 gnd.n2112 0.152939
R21438 gnd.n4517 gnd.n4516 0.152939
R21439 gnd.n4550 gnd.n4517 0.152939
R21440 gnd.n4550 gnd.n4549 0.152939
R21441 gnd.n6255 gnd.n1117 0.152939
R21442 gnd.n6251 gnd.n1117 0.152939
R21443 gnd.n6251 gnd.n6250 0.152939
R21444 gnd.n6250 gnd.n6249 0.152939
R21445 gnd.n6249 gnd.n1122 0.152939
R21446 gnd.n6245 gnd.n1122 0.152939
R21447 gnd.n6245 gnd.n6244 0.152939
R21448 gnd.n6244 gnd.n6243 0.152939
R21449 gnd.n6243 gnd.n1127 0.152939
R21450 gnd.n6239 gnd.n1127 0.152939
R21451 gnd.n6239 gnd.n6238 0.152939
R21452 gnd.n6238 gnd.n6237 0.152939
R21453 gnd.n6237 gnd.n1132 0.152939
R21454 gnd.n6233 gnd.n1132 0.152939
R21455 gnd.n6233 gnd.n6232 0.152939
R21456 gnd.n6232 gnd.n6231 0.152939
R21457 gnd.n6231 gnd.n1137 0.152939
R21458 gnd.n6227 gnd.n1137 0.152939
R21459 gnd.n6227 gnd.n6226 0.152939
R21460 gnd.n6226 gnd.n6225 0.152939
R21461 gnd.n6225 gnd.n1142 0.152939
R21462 gnd.n6221 gnd.n1142 0.152939
R21463 gnd.n6221 gnd.n6220 0.152939
R21464 gnd.n6220 gnd.n6219 0.152939
R21465 gnd.n6219 gnd.n1147 0.152939
R21466 gnd.n6215 gnd.n1147 0.152939
R21467 gnd.n6215 gnd.n6214 0.152939
R21468 gnd.n6214 gnd.n6213 0.152939
R21469 gnd.n6213 gnd.n1152 0.152939
R21470 gnd.n6209 gnd.n1152 0.152939
R21471 gnd.n6209 gnd.n6208 0.152939
R21472 gnd.n6208 gnd.n6207 0.152939
R21473 gnd.n6207 gnd.n1157 0.152939
R21474 gnd.n6203 gnd.n1157 0.152939
R21475 gnd.n6203 gnd.n6202 0.152939
R21476 gnd.n6202 gnd.n6201 0.152939
R21477 gnd.n6201 gnd.n1162 0.152939
R21478 gnd.n6197 gnd.n1162 0.152939
R21479 gnd.n6197 gnd.n6196 0.152939
R21480 gnd.n6196 gnd.n6195 0.152939
R21481 gnd.n6195 gnd.n1167 0.152939
R21482 gnd.n6191 gnd.n1167 0.152939
R21483 gnd.n6191 gnd.n6190 0.152939
R21484 gnd.n6190 gnd.n6189 0.152939
R21485 gnd.n6189 gnd.n1172 0.152939
R21486 gnd.n6185 gnd.n1172 0.152939
R21487 gnd.n6185 gnd.n6184 0.152939
R21488 gnd.n6184 gnd.n6183 0.152939
R21489 gnd.n6183 gnd.n1177 0.152939
R21490 gnd.n6179 gnd.n1177 0.152939
R21491 gnd.n6179 gnd.n6178 0.152939
R21492 gnd.n6178 gnd.n6177 0.152939
R21493 gnd.n6177 gnd.n1182 0.152939
R21494 gnd.n6173 gnd.n1182 0.152939
R21495 gnd.n6173 gnd.n6172 0.152939
R21496 gnd.n6172 gnd.n6171 0.152939
R21497 gnd.n6171 gnd.n1187 0.152939
R21498 gnd.n6167 gnd.n1187 0.152939
R21499 gnd.n6167 gnd.n6166 0.152939
R21500 gnd.n6166 gnd.n6165 0.152939
R21501 gnd.n6165 gnd.n1192 0.152939
R21502 gnd.n6161 gnd.n1192 0.152939
R21503 gnd.n6161 gnd.n6160 0.152939
R21504 gnd.n6160 gnd.n6159 0.152939
R21505 gnd.n6159 gnd.n1197 0.152939
R21506 gnd.n6155 gnd.n1197 0.152939
R21507 gnd.n6155 gnd.n6154 0.152939
R21508 gnd.n6154 gnd.n6153 0.152939
R21509 gnd.n6153 gnd.n1202 0.152939
R21510 gnd.n6149 gnd.n1202 0.152939
R21511 gnd.n6149 gnd.n6148 0.152939
R21512 gnd.n6148 gnd.n6147 0.152939
R21513 gnd.n6147 gnd.n1207 0.152939
R21514 gnd.n6143 gnd.n1207 0.152939
R21515 gnd.n6143 gnd.n6142 0.152939
R21516 gnd.n6142 gnd.n6141 0.152939
R21517 gnd.n6141 gnd.n1212 0.152939
R21518 gnd.n6137 gnd.n1212 0.152939
R21519 gnd.n6137 gnd.n6136 0.152939
R21520 gnd.n6136 gnd.n6135 0.152939
R21521 gnd.n6135 gnd.n1217 0.152939
R21522 gnd.n6131 gnd.n1217 0.152939
R21523 gnd.n6131 gnd.n6130 0.152939
R21524 gnd.n6130 gnd.n6129 0.152939
R21525 gnd.n6129 gnd.n1222 0.152939
R21526 gnd.n6125 gnd.n1222 0.152939
R21527 gnd.n6125 gnd.n6124 0.152939
R21528 gnd.n6124 gnd.n6123 0.152939
R21529 gnd.n6123 gnd.n1227 0.152939
R21530 gnd.n6119 gnd.n1227 0.152939
R21531 gnd.n6119 gnd.n6118 0.152939
R21532 gnd.n6118 gnd.n6117 0.152939
R21533 gnd.n6117 gnd.n1232 0.152939
R21534 gnd.n6113 gnd.n1232 0.152939
R21535 gnd.n6113 gnd.n6112 0.152939
R21536 gnd.n6112 gnd.n6111 0.152939
R21537 gnd.n6111 gnd.n1237 0.152939
R21538 gnd.n6107 gnd.n1237 0.152939
R21539 gnd.n6107 gnd.n6106 0.152939
R21540 gnd.n6106 gnd.n6105 0.152939
R21541 gnd.n6105 gnd.n1242 0.152939
R21542 gnd.n6013 gnd.n6012 0.152939
R21543 gnd.n6012 gnd.n6011 0.152939
R21544 gnd.n6011 gnd.n1343 0.152939
R21545 gnd.n6007 gnd.n1343 0.152939
R21546 gnd.n6007 gnd.n6006 0.152939
R21547 gnd.n6006 gnd.n6005 0.152939
R21548 gnd.n6005 gnd.n1348 0.152939
R21549 gnd.n6001 gnd.n1348 0.152939
R21550 gnd.n6001 gnd.n6000 0.152939
R21551 gnd.n6000 gnd.n5999 0.152939
R21552 gnd.n5999 gnd.n1353 0.152939
R21553 gnd.n5995 gnd.n1353 0.152939
R21554 gnd.n5995 gnd.n5994 0.152939
R21555 gnd.n5994 gnd.n5993 0.152939
R21556 gnd.n5993 gnd.n1358 0.152939
R21557 gnd.n5989 gnd.n1358 0.152939
R21558 gnd.n5989 gnd.n407 0.152939
R21559 gnd.n7169 gnd.n407 0.152939
R21560 gnd.n7169 gnd.n7168 0.152939
R21561 gnd.n7168 gnd.n7167 0.152939
R21562 gnd.n7167 gnd.n408 0.152939
R21563 gnd.n408 gnd.n375 0.152939
R21564 gnd.n7215 gnd.n375 0.152939
R21565 gnd.n7215 gnd.n7214 0.152939
R21566 gnd.n7214 gnd.n7213 0.152939
R21567 gnd.n7213 gnd.n376 0.152939
R21568 gnd.n7209 gnd.n376 0.152939
R21569 gnd.n7209 gnd.n320 0.152939
R21570 gnd.n7346 gnd.n320 0.152939
R21571 gnd.n7346 gnd.n7345 0.152939
R21572 gnd.n7345 gnd.n7344 0.152939
R21573 gnd.n7344 gnd.n321 0.152939
R21574 gnd.n7340 gnd.n321 0.152939
R21575 gnd.n7340 gnd.n7339 0.152939
R21576 gnd.n7339 gnd.n7338 0.152939
R21577 gnd.n7338 gnd.n326 0.152939
R21578 gnd.n326 gnd.n296 0.152939
R21579 gnd.n7361 gnd.n296 0.152939
R21580 gnd.n7362 gnd.n7361 0.152939
R21581 gnd.n7363 gnd.n7362 0.152939
R21582 gnd.n7363 gnd.n280 0.152939
R21583 gnd.n7377 gnd.n280 0.152939
R21584 gnd.n7378 gnd.n7377 0.152939
R21585 gnd.n7379 gnd.n7378 0.152939
R21586 gnd.n7379 gnd.n266 0.152939
R21587 gnd.n7393 gnd.n266 0.152939
R21588 gnd.n7394 gnd.n7393 0.152939
R21589 gnd.n7395 gnd.n7394 0.152939
R21590 gnd.n7395 gnd.n250 0.152939
R21591 gnd.n7409 gnd.n250 0.152939
R21592 gnd.n7410 gnd.n7409 0.152939
R21593 gnd.n7411 gnd.n7410 0.152939
R21594 gnd.n7411 gnd.n235 0.152939
R21595 gnd.n7425 gnd.n235 0.152939
R21596 gnd.n7426 gnd.n7425 0.152939
R21597 gnd.n7427 gnd.n7426 0.152939
R21598 gnd.n7427 gnd.n220 0.152939
R21599 gnd.n7441 gnd.n220 0.152939
R21600 gnd.n7442 gnd.n7441 0.152939
R21601 gnd.n7511 gnd.n7442 0.152939
R21602 gnd.n7511 gnd.n7510 0.152939
R21603 gnd.n7510 gnd.n7509 0.152939
R21604 gnd.n7509 gnd.n7443 0.152939
R21605 gnd.n7505 gnd.n7443 0.152939
R21606 gnd.n7504 gnd.n7445 0.152939
R21607 gnd.n7500 gnd.n7445 0.152939
R21608 gnd.n7500 gnd.n7499 0.152939
R21609 gnd.n7499 gnd.n7498 0.152939
R21610 gnd.n7498 gnd.n7451 0.152939
R21611 gnd.n7494 gnd.n7451 0.152939
R21612 gnd.n7494 gnd.n7493 0.152939
R21613 gnd.n7493 gnd.n7492 0.152939
R21614 gnd.n7492 gnd.n7459 0.152939
R21615 gnd.n7488 gnd.n7459 0.152939
R21616 gnd.n7488 gnd.n7487 0.152939
R21617 gnd.n7487 gnd.n7486 0.152939
R21618 gnd.n7486 gnd.n7467 0.152939
R21619 gnd.n7482 gnd.n7467 0.152939
R21620 gnd.n7482 gnd.n7481 0.152939
R21621 gnd.n7481 gnd.n7480 0.152939
R21622 gnd.n7480 gnd.n121 0.152939
R21623 gnd.n7606 gnd.n121 0.152939
R21624 gnd.n5854 gnd.n5840 0.152939
R21625 gnd.n5855 gnd.n5854 0.152939
R21626 gnd.n5857 gnd.n5855 0.152939
R21627 gnd.n5857 gnd.n5856 0.152939
R21628 gnd.n5856 gnd.n1419 0.152939
R21629 gnd.n5885 gnd.n1419 0.152939
R21630 gnd.n5886 gnd.n5885 0.152939
R21631 gnd.n5893 gnd.n5886 0.152939
R21632 gnd.n5893 gnd.n5892 0.152939
R21633 gnd.n5892 gnd.n5891 0.152939
R21634 gnd.n5891 gnd.n5887 0.152939
R21635 gnd.n5887 gnd.n1384 0.152939
R21636 gnd.n5953 gnd.n1384 0.152939
R21637 gnd.n5953 gnd.n5952 0.152939
R21638 gnd.n5952 gnd.n5951 0.152939
R21639 gnd.n5951 gnd.n1385 0.152939
R21640 gnd.n5947 gnd.n1385 0.152939
R21641 gnd.n5947 gnd.n5946 0.152939
R21642 gnd.n5946 gnd.n5945 0.152939
R21643 gnd.n5945 gnd.n5940 0.152939
R21644 gnd.n5940 gnd.n5939 0.152939
R21645 gnd.n5939 gnd.n381 0.152939
R21646 gnd.n7200 gnd.n381 0.152939
R21647 gnd.n7201 gnd.n7200 0.152939
R21648 gnd.n7203 gnd.n7201 0.152939
R21649 gnd.n7203 gnd.n7202 0.152939
R21650 gnd.n7202 gnd.n347 0.152939
R21651 gnd.n7245 gnd.n347 0.152939
R21652 gnd.n7246 gnd.n7245 0.152939
R21653 gnd.n7247 gnd.n7246 0.152939
R21654 gnd.n7247 gnd.n79 0.152939
R21655 gnd.n7655 gnd.n79 0.152939
R21656 gnd.n7655 gnd.n7654 0.152939
R21657 gnd.n7654 gnd.n81 0.152939
R21658 gnd.n7650 gnd.n81 0.152939
R21659 gnd.n7650 gnd.n7649 0.152939
R21660 gnd.n7649 gnd.n7648 0.152939
R21661 gnd.n7648 gnd.n86 0.152939
R21662 gnd.n7644 gnd.n86 0.152939
R21663 gnd.n7644 gnd.n7643 0.152939
R21664 gnd.n7643 gnd.n7642 0.152939
R21665 gnd.n7642 gnd.n91 0.152939
R21666 gnd.n7638 gnd.n91 0.152939
R21667 gnd.n7638 gnd.n7637 0.152939
R21668 gnd.n7637 gnd.n7636 0.152939
R21669 gnd.n7636 gnd.n96 0.152939
R21670 gnd.n7632 gnd.n96 0.152939
R21671 gnd.n7632 gnd.n7631 0.152939
R21672 gnd.n7631 gnd.n7630 0.152939
R21673 gnd.n7630 gnd.n101 0.152939
R21674 gnd.n7626 gnd.n101 0.152939
R21675 gnd.n7626 gnd.n7625 0.152939
R21676 gnd.n7625 gnd.n7624 0.152939
R21677 gnd.n7624 gnd.n106 0.152939
R21678 gnd.n7620 gnd.n106 0.152939
R21679 gnd.n7620 gnd.n7619 0.152939
R21680 gnd.n7619 gnd.n7618 0.152939
R21681 gnd.n7618 gnd.n111 0.152939
R21682 gnd.n7614 gnd.n111 0.152939
R21683 gnd.n7614 gnd.n7613 0.152939
R21684 gnd.n7613 gnd.n7612 0.152939
R21685 gnd.n7612 gnd.n116 0.152939
R21686 gnd.n7608 gnd.n116 0.152939
R21687 gnd.n7608 gnd.n7607 0.152939
R21688 gnd.n5839 gnd.n5838 0.151415
R21689 gnd.n4548 gnd.n4518 0.151415
R21690 gnd.n3908 gnd.n3894 0.145814
R21691 gnd.n3908 gnd.n3907 0.145814
R21692 gnd.n3190 gnd.n3189 0.0767195
R21693 gnd.n3189 gnd.n3188 0.0767195
R21694 gnd.n6257 gnd.n6256 0.063
R21695 gnd.n1518 gnd.n1342 0.063
R21696 gnd.n3756 gnd.n2359 0.0477147
R21697 gnd.n2953 gnd.n2841 0.0442063
R21698 gnd.n2954 gnd.n2953 0.0442063
R21699 gnd.n2955 gnd.n2954 0.0442063
R21700 gnd.n2955 gnd.n2830 0.0442063
R21701 gnd.n2969 gnd.n2830 0.0442063
R21702 gnd.n2970 gnd.n2969 0.0442063
R21703 gnd.n2971 gnd.n2970 0.0442063
R21704 gnd.n2971 gnd.n2817 0.0442063
R21705 gnd.n3015 gnd.n2817 0.0442063
R21706 gnd.n3016 gnd.n3015 0.0442063
R21707 gnd.n3018 gnd.n2751 0.0344674
R21708 gnd.n1597 gnd.n1478 0.0343753
R21709 gnd.n4547 gnd.n2025 0.0343753
R21710 gnd.n3038 gnd.n3037 0.0269946
R21711 gnd.n3040 gnd.n3039 0.0269946
R21712 gnd.n2746 gnd.n2744 0.0269946
R21713 gnd.n3050 gnd.n3048 0.0269946
R21714 gnd.n3049 gnd.n2725 0.0269946
R21715 gnd.n3069 gnd.n3068 0.0269946
R21716 gnd.n3071 gnd.n3070 0.0269946
R21717 gnd.n2720 gnd.n2719 0.0269946
R21718 gnd.n3081 gnd.n2715 0.0269946
R21719 gnd.n3080 gnd.n2717 0.0269946
R21720 gnd.n2716 gnd.n2698 0.0269946
R21721 gnd.n3101 gnd.n2699 0.0269946
R21722 gnd.n3100 gnd.n2700 0.0269946
R21723 gnd.n3134 gnd.n2675 0.0269946
R21724 gnd.n3136 gnd.n3135 0.0269946
R21725 gnd.n3137 gnd.n2622 0.0269946
R21726 gnd.n2670 gnd.n2623 0.0269946
R21727 gnd.n2672 gnd.n2624 0.0269946
R21728 gnd.n3147 gnd.n3146 0.0269946
R21729 gnd.n3149 gnd.n3148 0.0269946
R21730 gnd.n3150 gnd.n2644 0.0269946
R21731 gnd.n3152 gnd.n2645 0.0269946
R21732 gnd.n3155 gnd.n2646 0.0269946
R21733 gnd.n3158 gnd.n3157 0.0269946
R21734 gnd.n3160 gnd.n3159 0.0269946
R21735 gnd.n3225 gnd.n2533 0.0269946
R21736 gnd.n3227 gnd.n3226 0.0269946
R21737 gnd.n3236 gnd.n2526 0.0269946
R21738 gnd.n3238 gnd.n3237 0.0269946
R21739 gnd.n3239 gnd.n2524 0.0269946
R21740 gnd.n3246 gnd.n3242 0.0269946
R21741 gnd.n3245 gnd.n3244 0.0269946
R21742 gnd.n3243 gnd.n2503 0.0269946
R21743 gnd.n3268 gnd.n2504 0.0269946
R21744 gnd.n3267 gnd.n2505 0.0269946
R21745 gnd.n3310 gnd.n2478 0.0269946
R21746 gnd.n3312 gnd.n3311 0.0269946
R21747 gnd.n3321 gnd.n2471 0.0269946
R21748 gnd.n3323 gnd.n3322 0.0269946
R21749 gnd.n3324 gnd.n2469 0.0269946
R21750 gnd.n3331 gnd.n3327 0.0269946
R21751 gnd.n3330 gnd.n3329 0.0269946
R21752 gnd.n3328 gnd.n2448 0.0269946
R21753 gnd.n3353 gnd.n2449 0.0269946
R21754 gnd.n3352 gnd.n2450 0.0269946
R21755 gnd.n3399 gnd.n2424 0.0269946
R21756 gnd.n3401 gnd.n3400 0.0269946
R21757 gnd.n3410 gnd.n2417 0.0269946
R21758 gnd.n3669 gnd.n2415 0.0269946
R21759 gnd.n3674 gnd.n3672 0.0269946
R21760 gnd.n3673 gnd.n2396 0.0269946
R21761 gnd.n3698 gnd.n3697 0.0269946
R21762 gnd.n1520 gnd.n1518 0.0245515
R21763 gnd.n6256 gnd.n1116 0.0245515
R21764 gnd.n3018 gnd.n3017 0.0202011
R21765 gnd.n1520 gnd.n1519 0.0174377
R21766 gnd.n1519 gnd.n1515 0.0174377
R21767 gnd.n1529 gnd.n1515 0.0174377
R21768 gnd.n1529 gnd.n1528 0.0174377
R21769 gnd.n1528 gnd.n1516 0.0174377
R21770 gnd.n1516 gnd.n1511 0.0174377
R21771 gnd.n1537 gnd.n1511 0.0174377
R21772 gnd.n1539 gnd.n1537 0.0174377
R21773 gnd.n1539 gnd.n1538 0.0174377
R21774 gnd.n1538 gnd.n1508 0.0174377
R21775 gnd.n1548 gnd.n1508 0.0174377
R21776 gnd.n1548 gnd.n1547 0.0174377
R21777 gnd.n1547 gnd.n1509 0.0174377
R21778 gnd.n1509 gnd.n1504 0.0174377
R21779 gnd.n1556 gnd.n1504 0.0174377
R21780 gnd.n1558 gnd.n1556 0.0174377
R21781 gnd.n1558 gnd.n1557 0.0174377
R21782 gnd.n1557 gnd.n1501 0.0174377
R21783 gnd.n1567 gnd.n1501 0.0174377
R21784 gnd.n1567 gnd.n1566 0.0174377
R21785 gnd.n1566 gnd.n1502 0.0174377
R21786 gnd.n1502 gnd.n1497 0.0174377
R21787 gnd.n1575 gnd.n1497 0.0174377
R21788 gnd.n1576 gnd.n1575 0.0174377
R21789 gnd.n1576 gnd.n1495 0.0174377
R21790 gnd.n1581 gnd.n1495 0.0174377
R21791 gnd.n1583 gnd.n1581 0.0174377
R21792 gnd.n1583 gnd.n1582 0.0174377
R21793 gnd.n1582 gnd.n1491 0.0174377
R21794 gnd.n1592 gnd.n1491 0.0174377
R21795 gnd.n1592 gnd.n1591 0.0174377
R21796 gnd.n1591 gnd.n1484 0.0174377
R21797 gnd.n1484 gnd.n1483 0.0174377
R21798 gnd.n1596 gnd.n1483 0.0174377
R21799 gnd.n1597 gnd.n1596 0.0174377
R21800 gnd.n1974 gnd.n1116 0.0174377
R21801 gnd.n1976 gnd.n1974 0.0174377
R21802 gnd.n5399 gnd.n1976 0.0174377
R21803 gnd.n5399 gnd.n5398 0.0174377
R21804 gnd.n5398 gnd.n1977 0.0174377
R21805 gnd.n5395 gnd.n1977 0.0174377
R21806 gnd.n5395 gnd.n5394 0.0174377
R21807 gnd.n5394 gnd.n1982 0.0174377
R21808 gnd.n5391 gnd.n1982 0.0174377
R21809 gnd.n5391 gnd.n5390 0.0174377
R21810 gnd.n5390 gnd.n1987 0.0174377
R21811 gnd.n5387 gnd.n1987 0.0174377
R21812 gnd.n5387 gnd.n5386 0.0174377
R21813 gnd.n5386 gnd.n1991 0.0174377
R21814 gnd.n5383 gnd.n1991 0.0174377
R21815 gnd.n5383 gnd.n5382 0.0174377
R21816 gnd.n5382 gnd.n1995 0.0174377
R21817 gnd.n5379 gnd.n1995 0.0174377
R21818 gnd.n5379 gnd.n5378 0.0174377
R21819 gnd.n5378 gnd.n1999 0.0174377
R21820 gnd.n5375 gnd.n1999 0.0174377
R21821 gnd.n5375 gnd.n5374 0.0174377
R21822 gnd.n5374 gnd.n2005 0.0174377
R21823 gnd.n5371 gnd.n2005 0.0174377
R21824 gnd.n5371 gnd.n5370 0.0174377
R21825 gnd.n5370 gnd.n2009 0.0174377
R21826 gnd.n5367 gnd.n2009 0.0174377
R21827 gnd.n5367 gnd.n5366 0.0174377
R21828 gnd.n5366 gnd.n2013 0.0174377
R21829 gnd.n5363 gnd.n2013 0.0174377
R21830 gnd.n5363 gnd.n5362 0.0174377
R21831 gnd.n5362 gnd.n2019 0.0174377
R21832 gnd.n5359 gnd.n2019 0.0174377
R21833 gnd.n5359 gnd.n5358 0.0174377
R21834 gnd.n5358 gnd.n2025 0.0174377
R21835 gnd.n3017 gnd.n3016 0.0148637
R21836 gnd.n3667 gnd.n3411 0.0144266
R21837 gnd.n3668 gnd.n3667 0.0130679
R21838 gnd.n3037 gnd.n2751 0.00797283
R21839 gnd.n3039 gnd.n3038 0.00797283
R21840 gnd.n3040 gnd.n2746 0.00797283
R21841 gnd.n3048 gnd.n2744 0.00797283
R21842 gnd.n3050 gnd.n3049 0.00797283
R21843 gnd.n3068 gnd.n2725 0.00797283
R21844 gnd.n3070 gnd.n3069 0.00797283
R21845 gnd.n3071 gnd.n2720 0.00797283
R21846 gnd.n2719 gnd.n2715 0.00797283
R21847 gnd.n3081 gnd.n3080 0.00797283
R21848 gnd.n2717 gnd.n2716 0.00797283
R21849 gnd.n2699 gnd.n2698 0.00797283
R21850 gnd.n3101 gnd.n3100 0.00797283
R21851 gnd.n2700 gnd.n2675 0.00797283
R21852 gnd.n3135 gnd.n3134 0.00797283
R21853 gnd.n3137 gnd.n3136 0.00797283
R21854 gnd.n2670 gnd.n2622 0.00797283
R21855 gnd.n2672 gnd.n2623 0.00797283
R21856 gnd.n3146 gnd.n2624 0.00797283
R21857 gnd.n3148 gnd.n3147 0.00797283
R21858 gnd.n3150 gnd.n3149 0.00797283
R21859 gnd.n3152 gnd.n2644 0.00797283
R21860 gnd.n3155 gnd.n2645 0.00797283
R21861 gnd.n3157 gnd.n2646 0.00797283
R21862 gnd.n3160 gnd.n3158 0.00797283
R21863 gnd.n3159 gnd.n2533 0.00797283
R21864 gnd.n3227 gnd.n3225 0.00797283
R21865 gnd.n3226 gnd.n2526 0.00797283
R21866 gnd.n3237 gnd.n3236 0.00797283
R21867 gnd.n3239 gnd.n3238 0.00797283
R21868 gnd.n3242 gnd.n2524 0.00797283
R21869 gnd.n3246 gnd.n3245 0.00797283
R21870 gnd.n3244 gnd.n3243 0.00797283
R21871 gnd.n2504 gnd.n2503 0.00797283
R21872 gnd.n3268 gnd.n3267 0.00797283
R21873 gnd.n2505 gnd.n2478 0.00797283
R21874 gnd.n3312 gnd.n3310 0.00797283
R21875 gnd.n3311 gnd.n2471 0.00797283
R21876 gnd.n3322 gnd.n3321 0.00797283
R21877 gnd.n3324 gnd.n3323 0.00797283
R21878 gnd.n3327 gnd.n2469 0.00797283
R21879 gnd.n3331 gnd.n3330 0.00797283
R21880 gnd.n3329 gnd.n3328 0.00797283
R21881 gnd.n2449 gnd.n2448 0.00797283
R21882 gnd.n3353 gnd.n3352 0.00797283
R21883 gnd.n2450 gnd.n2424 0.00797283
R21884 gnd.n3401 gnd.n3399 0.00797283
R21885 gnd.n3400 gnd.n2417 0.00797283
R21886 gnd.n3411 gnd.n3410 0.00797283
R21887 gnd.n3669 gnd.n3668 0.00797283
R21888 gnd.n3672 gnd.n2415 0.00797283
R21889 gnd.n3674 gnd.n3673 0.00797283
R21890 gnd.n3697 gnd.n2396 0.00797283
R21891 gnd.n3698 gnd.n2359 0.00797283
R21892 gnd.n337 gnd.n321 0.00433921
R21893 gnd.n4313 gnd.n4312 0.00433921
R21894 gnd.n5839 gnd.n1478 0.000838753
R21895 gnd.n4548 gnd.n4547 0.000838753
R21896 diffpairibias.n0 diffpairibias.t27 436.822
R21897 diffpairibias.n27 diffpairibias.t24 435.479
R21898 diffpairibias.n26 diffpairibias.t21 435.479
R21899 diffpairibias.n25 diffpairibias.t22 435.479
R21900 diffpairibias.n24 diffpairibias.t26 435.479
R21901 diffpairibias.n23 diffpairibias.t20 435.479
R21902 diffpairibias.n0 diffpairibias.t23 435.479
R21903 diffpairibias.n1 diffpairibias.t28 435.479
R21904 diffpairibias.n2 diffpairibias.t25 435.479
R21905 diffpairibias.n3 diffpairibias.t29 435.479
R21906 diffpairibias.n13 diffpairibias.t14 377.536
R21907 diffpairibias.n13 diffpairibias.t0 376.193
R21908 diffpairibias.n14 diffpairibias.t10 376.193
R21909 diffpairibias.n15 diffpairibias.t12 376.193
R21910 diffpairibias.n16 diffpairibias.t6 376.193
R21911 diffpairibias.n17 diffpairibias.t2 376.193
R21912 diffpairibias.n18 diffpairibias.t16 376.193
R21913 diffpairibias.n19 diffpairibias.t4 376.193
R21914 diffpairibias.n20 diffpairibias.t18 376.193
R21915 diffpairibias.n21 diffpairibias.t8 376.193
R21916 diffpairibias.n4 diffpairibias.t15 113.368
R21917 diffpairibias.n4 diffpairibias.t1 112.698
R21918 diffpairibias.n5 diffpairibias.t11 112.698
R21919 diffpairibias.n6 diffpairibias.t13 112.698
R21920 diffpairibias.n7 diffpairibias.t7 112.698
R21921 diffpairibias.n8 diffpairibias.t3 112.698
R21922 diffpairibias.n9 diffpairibias.t17 112.698
R21923 diffpairibias.n10 diffpairibias.t5 112.698
R21924 diffpairibias.n11 diffpairibias.t19 112.698
R21925 diffpairibias.n12 diffpairibias.t9 112.698
R21926 diffpairibias.n22 diffpairibias.n21 4.77242
R21927 diffpairibias.n22 diffpairibias.n12 4.30807
R21928 diffpairibias.n23 diffpairibias.n22 4.13945
R21929 diffpairibias.n21 diffpairibias.n20 1.34352
R21930 diffpairibias.n20 diffpairibias.n19 1.34352
R21931 diffpairibias.n19 diffpairibias.n18 1.34352
R21932 diffpairibias.n18 diffpairibias.n17 1.34352
R21933 diffpairibias.n17 diffpairibias.n16 1.34352
R21934 diffpairibias.n16 diffpairibias.n15 1.34352
R21935 diffpairibias.n15 diffpairibias.n14 1.34352
R21936 diffpairibias.n14 diffpairibias.n13 1.34352
R21937 diffpairibias.n3 diffpairibias.n2 1.34352
R21938 diffpairibias.n2 diffpairibias.n1 1.34352
R21939 diffpairibias.n1 diffpairibias.n0 1.34352
R21940 diffpairibias.n24 diffpairibias.n23 1.34352
R21941 diffpairibias.n25 diffpairibias.n24 1.34352
R21942 diffpairibias.n26 diffpairibias.n25 1.34352
R21943 diffpairibias.n27 diffpairibias.n26 1.34352
R21944 diffpairibias.n28 diffpairibias.n27 0.862419
R21945 diffpairibias diffpairibias.n28 0.684875
R21946 diffpairibias.n12 diffpairibias.n11 0.672012
R21947 diffpairibias.n11 diffpairibias.n10 0.672012
R21948 diffpairibias.n10 diffpairibias.n9 0.672012
R21949 diffpairibias.n9 diffpairibias.n8 0.672012
R21950 diffpairibias.n8 diffpairibias.n7 0.672012
R21951 diffpairibias.n7 diffpairibias.n6 0.672012
R21952 diffpairibias.n6 diffpairibias.n5 0.672012
R21953 diffpairibias.n5 diffpairibias.n4 0.672012
R21954 diffpairibias.n28 diffpairibias.n3 0.190907
R21955 a_n3827_n3924.n42 a_n3827_n3924.t10 214.994
R21956 a_n3827_n3924.t17 a_n3827_n3924.n51 214.994
R21957 a_n3827_n3924.n42 a_n3827_n3924.t14 214.321
R21958 a_n3827_n3924.n44 a_n3827_n3924.t9 214.321
R21959 a_n3827_n3924.n45 a_n3827_n3924.t12 214.321
R21960 a_n3827_n3924.n46 a_n3827_n3924.t8 214.321
R21961 a_n3827_n3924.n47 a_n3827_n3924.t13 214.321
R21962 a_n3827_n3924.n48 a_n3827_n3924.t16 214.321
R21963 a_n3827_n3924.n50 a_n3827_n3924.t15 214.321
R21964 a_n3827_n3924.n51 a_n3827_n3924.t11 214.321
R21965 a_n3827_n3924.n11 a_n3827_n3924.t22 55.8337
R21966 a_n3827_n3924.n10 a_n3827_n3924.t45 55.8337
R21967 a_n3827_n3924.n1 a_n3827_n3924.t47 55.8337
R21968 a_n3827_n3924.n20 a_n3827_n3924.t6 55.8335
R21969 a_n3827_n3924.n40 a_n3827_n3924.t4 55.8335
R21970 a_n3827_n3924.n31 a_n3827_n3924.t37 55.8335
R21971 a_n3827_n3924.n30 a_n3827_n3924.t34 55.8335
R21972 a_n3827_n3924.n21 a_n3827_n3924.t19 55.8335
R21973 a_n3827_n3924.n19 a_n3827_n3924.n18 53.0052
R21974 a_n3827_n3924.n17 a_n3827_n3924.n16 53.0052
R21975 a_n3827_n3924.n15 a_n3827_n3924.n14 53.0052
R21976 a_n3827_n3924.n13 a_n3827_n3924.n12 53.0052
R21977 a_n3827_n3924.n9 a_n3827_n3924.n8 53.0052
R21978 a_n3827_n3924.n7 a_n3827_n3924.n6 53.0052
R21979 a_n3827_n3924.n5 a_n3827_n3924.n4 53.0052
R21980 a_n3827_n3924.n3 a_n3827_n3924.n2 53.0052
R21981 a_n3827_n3924.n39 a_n3827_n3924.n38 53.0051
R21982 a_n3827_n3924.n37 a_n3827_n3924.n36 53.0051
R21983 a_n3827_n3924.n35 a_n3827_n3924.n34 53.0051
R21984 a_n3827_n3924.n33 a_n3827_n3924.n32 53.0051
R21985 a_n3827_n3924.n29 a_n3827_n3924.n28 53.0051
R21986 a_n3827_n3924.n27 a_n3827_n3924.n26 53.0051
R21987 a_n3827_n3924.n25 a_n3827_n3924.n24 53.0051
R21988 a_n3827_n3924.n23 a_n3827_n3924.n22 53.0051
R21989 a_n3827_n3924.n1 a_n3827_n3924.n0 12.1555
R21990 a_n3827_n3924.n41 a_n3827_n3924.n20 12.1555
R21991 a_n3827_n3924.n21 a_n3827_n3924.n0 5.07593
R21992 a_n3827_n3924.n41 a_n3827_n3924.n40 5.07593
R21993 a_n3827_n3924.n38 a_n3827_n3924.t41 2.82907
R21994 a_n3827_n3924.n38 a_n3827_n3924.t24 2.82907
R21995 a_n3827_n3924.n36 a_n3827_n3924.t26 2.82907
R21996 a_n3827_n3924.n36 a_n3827_n3924.t30 2.82907
R21997 a_n3827_n3924.n34 a_n3827_n3924.t48 2.82907
R21998 a_n3827_n3924.n34 a_n3827_n3924.t23 2.82907
R21999 a_n3827_n3924.n32 a_n3827_n3924.t5 2.82907
R22000 a_n3827_n3924.n32 a_n3827_n3924.t1 2.82907
R22001 a_n3827_n3924.n28 a_n3827_n3924.t3 2.82907
R22002 a_n3827_n3924.n28 a_n3827_n3924.t40 2.82907
R22003 a_n3827_n3924.n26 a_n3827_n3924.t18 2.82907
R22004 a_n3827_n3924.n26 a_n3827_n3924.t0 2.82907
R22005 a_n3827_n3924.n24 a_n3827_n3924.t39 2.82907
R22006 a_n3827_n3924.n24 a_n3827_n3924.t35 2.82907
R22007 a_n3827_n3924.n22 a_n3827_n3924.t36 2.82907
R22008 a_n3827_n3924.n22 a_n3827_n3924.t49 2.82907
R22009 a_n3827_n3924.n18 a_n3827_n3924.t21 2.82907
R22010 a_n3827_n3924.n18 a_n3827_n3924.t33 2.82907
R22011 a_n3827_n3924.n16 a_n3827_n3924.t44 2.82907
R22012 a_n3827_n3924.n16 a_n3827_n3924.t7 2.82907
R22013 a_n3827_n3924.n14 a_n3827_n3924.t32 2.82907
R22014 a_n3827_n3924.n14 a_n3827_n3924.t20 2.82907
R22015 a_n3827_n3924.n12 a_n3827_n3924.t43 2.82907
R22016 a_n3827_n3924.n12 a_n3827_n3924.t27 2.82907
R22017 a_n3827_n3924.n8 a_n3827_n3924.t46 2.82907
R22018 a_n3827_n3924.n8 a_n3827_n3924.t29 2.82907
R22019 a_n3827_n3924.n6 a_n3827_n3924.t2 2.82907
R22020 a_n3827_n3924.n6 a_n3827_n3924.t28 2.82907
R22021 a_n3827_n3924.n4 a_n3827_n3924.t38 2.82907
R22022 a_n3827_n3924.n4 a_n3827_n3924.t42 2.82907
R22023 a_n3827_n3924.n2 a_n3827_n3924.t31 2.82907
R22024 a_n3827_n3924.n2 a_n3827_n3924.t25 2.82907
R22025 a_n3827_n3924.n49 a_n3827_n3924.n0 1.95694
R22026 a_n3827_n3924.n43 a_n3827_n3924.n41 1.95694
R22027 a_n3827_n3924.n51 a_n3827_n3924.n50 0.672012
R22028 a_n3827_n3924.n48 a_n3827_n3924.n47 0.672012
R22029 a_n3827_n3924.n47 a_n3827_n3924.n46 0.672012
R22030 a_n3827_n3924.n46 a_n3827_n3924.n45 0.672012
R22031 a_n3827_n3924.n45 a_n3827_n3924.n44 0.672012
R22032 a_n3827_n3924.n43 a_n3827_n3924.n42 0.412564
R22033 a_n3827_n3924.n49 a_n3827_n3924.n48 0.40239
R22034 a_n3827_n3924.n3 a_n3827_n3924.n1 0.358259
R22035 a_n3827_n3924.n5 a_n3827_n3924.n3 0.358259
R22036 a_n3827_n3924.n7 a_n3827_n3924.n5 0.358259
R22037 a_n3827_n3924.n9 a_n3827_n3924.n7 0.358259
R22038 a_n3827_n3924.n10 a_n3827_n3924.n9 0.358259
R22039 a_n3827_n3924.n13 a_n3827_n3924.n11 0.358259
R22040 a_n3827_n3924.n15 a_n3827_n3924.n13 0.358259
R22041 a_n3827_n3924.n17 a_n3827_n3924.n15 0.358259
R22042 a_n3827_n3924.n19 a_n3827_n3924.n17 0.358259
R22043 a_n3827_n3924.n20 a_n3827_n3924.n19 0.358259
R22044 a_n3827_n3924.n23 a_n3827_n3924.n21 0.358259
R22045 a_n3827_n3924.n25 a_n3827_n3924.n23 0.358259
R22046 a_n3827_n3924.n27 a_n3827_n3924.n25 0.358259
R22047 a_n3827_n3924.n29 a_n3827_n3924.n27 0.358259
R22048 a_n3827_n3924.n30 a_n3827_n3924.n29 0.358259
R22049 a_n3827_n3924.n33 a_n3827_n3924.n31 0.358259
R22050 a_n3827_n3924.n35 a_n3827_n3924.n33 0.358259
R22051 a_n3827_n3924.n37 a_n3827_n3924.n35 0.358259
R22052 a_n3827_n3924.n39 a_n3827_n3924.n37 0.358259
R22053 a_n3827_n3924.n40 a_n3827_n3924.n39 0.358259
R22054 a_n3827_n3924.n50 a_n3827_n3924.n49 0.270122
R22055 a_n3827_n3924.n44 a_n3827_n3924.n43 0.259948
R22056 a_n3827_n3924.n11 a_n3827_n3924.n10 0.235414
R22057 a_n3827_n3924.n31 a_n3827_n3924.n30 0.235414
R22058 commonsourceibias.n281 commonsourceibias.t101 222.032
R22059 commonsourceibias.n44 commonsourceibias.t78 222.032
R22060 commonsourceibias.n166 commonsourceibias.t117 222.032
R22061 commonsourceibias.n643 commonsourceibias.t106 222.032
R22062 commonsourceibias.n413 commonsourceibias.t28 222.032
R22063 commonsourceibias.n529 commonsourceibias.t123 222.032
R22064 commonsourceibias.n364 commonsourceibias.t100 207.983
R22065 commonsourceibias.n127 commonsourceibias.t74 207.983
R22066 commonsourceibias.n249 commonsourceibias.t115 207.983
R22067 commonsourceibias.n731 commonsourceibias.t122 207.983
R22068 commonsourceibias.n501 commonsourceibias.t14 207.983
R22069 commonsourceibias.n616 commonsourceibias.t140 207.983
R22070 commonsourceibias.n280 commonsourceibias.t87 168.701
R22071 commonsourceibias.n286 commonsourceibias.t129 168.701
R22072 commonsourceibias.n292 commonsourceibias.t110 168.701
R22073 commonsourceibias.n276 commonsourceibias.t93 168.701
R22074 commonsourceibias.n300 commonsourceibias.t95 168.701
R22075 commonsourceibias.n306 commonsourceibias.t121 168.701
R22076 commonsourceibias.n271 commonsourceibias.t102 168.701
R22077 commonsourceibias.n314 commonsourceibias.t108 168.701
R22078 commonsourceibias.n320 commonsourceibias.t159 168.701
R22079 commonsourceibias.n266 commonsourceibias.t138 168.701
R22080 commonsourceibias.n328 commonsourceibias.t118 168.701
R22081 commonsourceibias.n334 commonsourceibias.t83 168.701
R22082 commonsourceibias.n261 commonsourceibias.t86 168.701
R22083 commonsourceibias.n342 commonsourceibias.t128 168.701
R22084 commonsourceibias.n348 commonsourceibias.t109 168.701
R22085 commonsourceibias.n256 commonsourceibias.t92 168.701
R22086 commonsourceibias.n356 commonsourceibias.t137 168.701
R22087 commonsourceibias.n362 commonsourceibias.t119 168.701
R22088 commonsourceibias.n125 commonsourceibias.t20 168.701
R22089 commonsourceibias.n119 commonsourceibias.t50 168.701
R22090 commonsourceibias.n19 commonsourceibias.t8 168.701
R22091 commonsourceibias.n111 commonsourceibias.t36 168.701
R22092 commonsourceibias.n105 commonsourceibias.t76 168.701
R22093 commonsourceibias.n24 commonsourceibias.t24 168.701
R22094 commonsourceibias.n97 commonsourceibias.t34 168.701
R22095 commonsourceibias.n91 commonsourceibias.t10 168.701
R22096 commonsourceibias.n29 commonsourceibias.t40 168.701
R22097 commonsourceibias.n83 commonsourceibias.t56 168.701
R22098 commonsourceibias.n77 commonsourceibias.t26 168.701
R22099 commonsourceibias.n34 commonsourceibias.t38 168.701
R22100 commonsourceibias.n69 commonsourceibias.t70 168.701
R22101 commonsourceibias.n63 commonsourceibias.t18 168.701
R22102 commonsourceibias.n39 commonsourceibias.t22 168.701
R22103 commonsourceibias.n55 commonsourceibias.t54 168.701
R22104 commonsourceibias.n49 commonsourceibias.t4 168.701
R22105 commonsourceibias.n43 commonsourceibias.t46 168.701
R22106 commonsourceibias.n247 commonsourceibias.t136 168.701
R22107 commonsourceibias.n241 commonsourceibias.t151 168.701
R22108 commonsourceibias.n5 commonsourceibias.t105 168.701
R22109 commonsourceibias.n233 commonsourceibias.t126 168.701
R22110 commonsourceibias.n227 commonsourceibias.t144 168.701
R22111 commonsourceibias.n10 commonsourceibias.t98 168.701
R22112 commonsourceibias.n219 commonsourceibias.t94 168.701
R22113 commonsourceibias.n213 commonsourceibias.t135 168.701
R22114 commonsourceibias.n150 commonsourceibias.t153 168.701
R22115 commonsourceibias.n151 commonsourceibias.t88 168.701
R22116 commonsourceibias.n153 commonsourceibias.t125 168.701
R22117 commonsourceibias.n155 commonsourceibias.t120 168.701
R22118 commonsourceibias.n191 commonsourceibias.t139 168.701
R22119 commonsourceibias.n185 commonsourceibias.t112 168.701
R22120 commonsourceibias.n161 commonsourceibias.t107 168.701
R22121 commonsourceibias.n177 commonsourceibias.t127 168.701
R22122 commonsourceibias.n171 commonsourceibias.t146 168.701
R22123 commonsourceibias.n165 commonsourceibias.t99 168.701
R22124 commonsourceibias.n642 commonsourceibias.t90 168.701
R22125 commonsourceibias.n648 commonsourceibias.t134 168.701
R22126 commonsourceibias.n654 commonsourceibias.t116 168.701
R22127 commonsourceibias.n656 commonsourceibias.t96 168.701
R22128 commonsourceibias.n663 commonsourceibias.t91 168.701
R22129 commonsourceibias.n669 commonsourceibias.t145 168.701
R22130 commonsourceibias.n671 commonsourceibias.t124 168.701
R22131 commonsourceibias.n678 commonsourceibias.t131 168.701
R22132 commonsourceibias.n684 commonsourceibias.t152 168.701
R22133 commonsourceibias.n686 commonsourceibias.t157 168.701
R22134 commonsourceibias.n693 commonsourceibias.t141 168.701
R22135 commonsourceibias.n699 commonsourceibias.t97 168.701
R22136 commonsourceibias.n701 commonsourceibias.t81 168.701
R22137 commonsourceibias.n708 commonsourceibias.t149 168.701
R22138 commonsourceibias.n714 commonsourceibias.t132 168.701
R22139 commonsourceibias.n716 commonsourceibias.t111 168.701
R22140 commonsourceibias.n723 commonsourceibias.t156 168.701
R22141 commonsourceibias.n729 commonsourceibias.t142 168.701
R22142 commonsourceibias.n412 commonsourceibias.t2 168.701
R22143 commonsourceibias.n418 commonsourceibias.t48 168.701
R22144 commonsourceibias.n424 commonsourceibias.t12 168.701
R22145 commonsourceibias.n426 commonsourceibias.t68 168.701
R22146 commonsourceibias.n433 commonsourceibias.t66 168.701
R22147 commonsourceibias.n439 commonsourceibias.t6 168.701
R22148 commonsourceibias.n441 commonsourceibias.t62 168.701
R22149 commonsourceibias.n448 commonsourceibias.t52 168.701
R22150 commonsourceibias.n454 commonsourceibias.t72 168.701
R22151 commonsourceibias.n456 commonsourceibias.t64 168.701
R22152 commonsourceibias.n463 commonsourceibias.t32 168.701
R22153 commonsourceibias.n469 commonsourceibias.t58 168.701
R22154 commonsourceibias.n471 commonsourceibias.t44 168.701
R22155 commonsourceibias.n478 commonsourceibias.t16 168.701
R22156 commonsourceibias.n484 commonsourceibias.t60 168.701
R22157 commonsourceibias.n486 commonsourceibias.t30 168.701
R22158 commonsourceibias.n493 commonsourceibias.t0 168.701
R22159 commonsourceibias.n499 commonsourceibias.t42 168.701
R22160 commonsourceibias.n614 commonsourceibias.t155 168.701
R22161 commonsourceibias.n608 commonsourceibias.t84 168.701
R22162 commonsourceibias.n601 commonsourceibias.t130 168.701
R22163 commonsourceibias.n599 commonsourceibias.t148 168.701
R22164 commonsourceibias.n593 commonsourceibias.t80 168.701
R22165 commonsourceibias.n586 commonsourceibias.t89 168.701
R22166 commonsourceibias.n584 commonsourceibias.t113 168.701
R22167 commonsourceibias.n578 commonsourceibias.t154 168.701
R22168 commonsourceibias.n571 commonsourceibias.t85 168.701
R22169 commonsourceibias.n528 commonsourceibias.t103 168.701
R22170 commonsourceibias.n534 commonsourceibias.t150 168.701
R22171 commonsourceibias.n540 commonsourceibias.t133 168.701
R22172 commonsourceibias.n542 commonsourceibias.t114 168.701
R22173 commonsourceibias.n549 commonsourceibias.t104 168.701
R22174 commonsourceibias.n555 commonsourceibias.t158 168.701
R22175 commonsourceibias.n519 commonsourceibias.t143 168.701
R22176 commonsourceibias.n517 commonsourceibias.t147 168.701
R22177 commonsourceibias.n515 commonsourceibias.t82 168.701
R22178 commonsourceibias.n363 commonsourceibias.n251 161.3
R22179 commonsourceibias.n361 commonsourceibias.n360 161.3
R22180 commonsourceibias.n359 commonsourceibias.n252 161.3
R22181 commonsourceibias.n358 commonsourceibias.n357 161.3
R22182 commonsourceibias.n355 commonsourceibias.n253 161.3
R22183 commonsourceibias.n354 commonsourceibias.n353 161.3
R22184 commonsourceibias.n352 commonsourceibias.n254 161.3
R22185 commonsourceibias.n351 commonsourceibias.n350 161.3
R22186 commonsourceibias.n349 commonsourceibias.n255 161.3
R22187 commonsourceibias.n347 commonsourceibias.n346 161.3
R22188 commonsourceibias.n345 commonsourceibias.n257 161.3
R22189 commonsourceibias.n344 commonsourceibias.n343 161.3
R22190 commonsourceibias.n341 commonsourceibias.n258 161.3
R22191 commonsourceibias.n340 commonsourceibias.n339 161.3
R22192 commonsourceibias.n338 commonsourceibias.n259 161.3
R22193 commonsourceibias.n337 commonsourceibias.n336 161.3
R22194 commonsourceibias.n335 commonsourceibias.n260 161.3
R22195 commonsourceibias.n333 commonsourceibias.n332 161.3
R22196 commonsourceibias.n331 commonsourceibias.n262 161.3
R22197 commonsourceibias.n330 commonsourceibias.n329 161.3
R22198 commonsourceibias.n327 commonsourceibias.n263 161.3
R22199 commonsourceibias.n326 commonsourceibias.n325 161.3
R22200 commonsourceibias.n324 commonsourceibias.n264 161.3
R22201 commonsourceibias.n323 commonsourceibias.n322 161.3
R22202 commonsourceibias.n321 commonsourceibias.n265 161.3
R22203 commonsourceibias.n319 commonsourceibias.n318 161.3
R22204 commonsourceibias.n317 commonsourceibias.n267 161.3
R22205 commonsourceibias.n316 commonsourceibias.n315 161.3
R22206 commonsourceibias.n313 commonsourceibias.n268 161.3
R22207 commonsourceibias.n312 commonsourceibias.n311 161.3
R22208 commonsourceibias.n310 commonsourceibias.n269 161.3
R22209 commonsourceibias.n309 commonsourceibias.n308 161.3
R22210 commonsourceibias.n307 commonsourceibias.n270 161.3
R22211 commonsourceibias.n305 commonsourceibias.n304 161.3
R22212 commonsourceibias.n303 commonsourceibias.n272 161.3
R22213 commonsourceibias.n302 commonsourceibias.n301 161.3
R22214 commonsourceibias.n299 commonsourceibias.n273 161.3
R22215 commonsourceibias.n298 commonsourceibias.n297 161.3
R22216 commonsourceibias.n296 commonsourceibias.n274 161.3
R22217 commonsourceibias.n295 commonsourceibias.n294 161.3
R22218 commonsourceibias.n293 commonsourceibias.n275 161.3
R22219 commonsourceibias.n291 commonsourceibias.n290 161.3
R22220 commonsourceibias.n289 commonsourceibias.n277 161.3
R22221 commonsourceibias.n288 commonsourceibias.n287 161.3
R22222 commonsourceibias.n285 commonsourceibias.n278 161.3
R22223 commonsourceibias.n284 commonsourceibias.n283 161.3
R22224 commonsourceibias.n282 commonsourceibias.n279 161.3
R22225 commonsourceibias.n45 commonsourceibias.n42 161.3
R22226 commonsourceibias.n47 commonsourceibias.n46 161.3
R22227 commonsourceibias.n48 commonsourceibias.n41 161.3
R22228 commonsourceibias.n51 commonsourceibias.n50 161.3
R22229 commonsourceibias.n52 commonsourceibias.n40 161.3
R22230 commonsourceibias.n54 commonsourceibias.n53 161.3
R22231 commonsourceibias.n56 commonsourceibias.n38 161.3
R22232 commonsourceibias.n58 commonsourceibias.n57 161.3
R22233 commonsourceibias.n59 commonsourceibias.n37 161.3
R22234 commonsourceibias.n61 commonsourceibias.n60 161.3
R22235 commonsourceibias.n62 commonsourceibias.n36 161.3
R22236 commonsourceibias.n65 commonsourceibias.n64 161.3
R22237 commonsourceibias.n66 commonsourceibias.n35 161.3
R22238 commonsourceibias.n68 commonsourceibias.n67 161.3
R22239 commonsourceibias.n70 commonsourceibias.n33 161.3
R22240 commonsourceibias.n72 commonsourceibias.n71 161.3
R22241 commonsourceibias.n73 commonsourceibias.n32 161.3
R22242 commonsourceibias.n75 commonsourceibias.n74 161.3
R22243 commonsourceibias.n76 commonsourceibias.n31 161.3
R22244 commonsourceibias.n79 commonsourceibias.n78 161.3
R22245 commonsourceibias.n80 commonsourceibias.n30 161.3
R22246 commonsourceibias.n82 commonsourceibias.n81 161.3
R22247 commonsourceibias.n84 commonsourceibias.n28 161.3
R22248 commonsourceibias.n86 commonsourceibias.n85 161.3
R22249 commonsourceibias.n87 commonsourceibias.n27 161.3
R22250 commonsourceibias.n89 commonsourceibias.n88 161.3
R22251 commonsourceibias.n90 commonsourceibias.n26 161.3
R22252 commonsourceibias.n93 commonsourceibias.n92 161.3
R22253 commonsourceibias.n94 commonsourceibias.n25 161.3
R22254 commonsourceibias.n96 commonsourceibias.n95 161.3
R22255 commonsourceibias.n98 commonsourceibias.n23 161.3
R22256 commonsourceibias.n100 commonsourceibias.n99 161.3
R22257 commonsourceibias.n101 commonsourceibias.n22 161.3
R22258 commonsourceibias.n103 commonsourceibias.n102 161.3
R22259 commonsourceibias.n104 commonsourceibias.n21 161.3
R22260 commonsourceibias.n107 commonsourceibias.n106 161.3
R22261 commonsourceibias.n108 commonsourceibias.n20 161.3
R22262 commonsourceibias.n110 commonsourceibias.n109 161.3
R22263 commonsourceibias.n112 commonsourceibias.n18 161.3
R22264 commonsourceibias.n114 commonsourceibias.n113 161.3
R22265 commonsourceibias.n115 commonsourceibias.n17 161.3
R22266 commonsourceibias.n117 commonsourceibias.n116 161.3
R22267 commonsourceibias.n118 commonsourceibias.n16 161.3
R22268 commonsourceibias.n121 commonsourceibias.n120 161.3
R22269 commonsourceibias.n122 commonsourceibias.n15 161.3
R22270 commonsourceibias.n124 commonsourceibias.n123 161.3
R22271 commonsourceibias.n126 commonsourceibias.n14 161.3
R22272 commonsourceibias.n167 commonsourceibias.n164 161.3
R22273 commonsourceibias.n169 commonsourceibias.n168 161.3
R22274 commonsourceibias.n170 commonsourceibias.n163 161.3
R22275 commonsourceibias.n173 commonsourceibias.n172 161.3
R22276 commonsourceibias.n174 commonsourceibias.n162 161.3
R22277 commonsourceibias.n176 commonsourceibias.n175 161.3
R22278 commonsourceibias.n178 commonsourceibias.n160 161.3
R22279 commonsourceibias.n180 commonsourceibias.n179 161.3
R22280 commonsourceibias.n181 commonsourceibias.n159 161.3
R22281 commonsourceibias.n183 commonsourceibias.n182 161.3
R22282 commonsourceibias.n184 commonsourceibias.n158 161.3
R22283 commonsourceibias.n187 commonsourceibias.n186 161.3
R22284 commonsourceibias.n188 commonsourceibias.n157 161.3
R22285 commonsourceibias.n190 commonsourceibias.n189 161.3
R22286 commonsourceibias.n192 commonsourceibias.n156 161.3
R22287 commonsourceibias.n194 commonsourceibias.n193 161.3
R22288 commonsourceibias.n196 commonsourceibias.n195 161.3
R22289 commonsourceibias.n197 commonsourceibias.n154 161.3
R22290 commonsourceibias.n199 commonsourceibias.n198 161.3
R22291 commonsourceibias.n201 commonsourceibias.n200 161.3
R22292 commonsourceibias.n202 commonsourceibias.n152 161.3
R22293 commonsourceibias.n204 commonsourceibias.n203 161.3
R22294 commonsourceibias.n206 commonsourceibias.n205 161.3
R22295 commonsourceibias.n208 commonsourceibias.n207 161.3
R22296 commonsourceibias.n209 commonsourceibias.n13 161.3
R22297 commonsourceibias.n211 commonsourceibias.n210 161.3
R22298 commonsourceibias.n212 commonsourceibias.n12 161.3
R22299 commonsourceibias.n215 commonsourceibias.n214 161.3
R22300 commonsourceibias.n216 commonsourceibias.n11 161.3
R22301 commonsourceibias.n218 commonsourceibias.n217 161.3
R22302 commonsourceibias.n220 commonsourceibias.n9 161.3
R22303 commonsourceibias.n222 commonsourceibias.n221 161.3
R22304 commonsourceibias.n223 commonsourceibias.n8 161.3
R22305 commonsourceibias.n225 commonsourceibias.n224 161.3
R22306 commonsourceibias.n226 commonsourceibias.n7 161.3
R22307 commonsourceibias.n229 commonsourceibias.n228 161.3
R22308 commonsourceibias.n230 commonsourceibias.n6 161.3
R22309 commonsourceibias.n232 commonsourceibias.n231 161.3
R22310 commonsourceibias.n234 commonsourceibias.n4 161.3
R22311 commonsourceibias.n236 commonsourceibias.n235 161.3
R22312 commonsourceibias.n237 commonsourceibias.n3 161.3
R22313 commonsourceibias.n239 commonsourceibias.n238 161.3
R22314 commonsourceibias.n240 commonsourceibias.n2 161.3
R22315 commonsourceibias.n243 commonsourceibias.n242 161.3
R22316 commonsourceibias.n244 commonsourceibias.n1 161.3
R22317 commonsourceibias.n246 commonsourceibias.n245 161.3
R22318 commonsourceibias.n248 commonsourceibias.n0 161.3
R22319 commonsourceibias.n730 commonsourceibias.n618 161.3
R22320 commonsourceibias.n728 commonsourceibias.n727 161.3
R22321 commonsourceibias.n726 commonsourceibias.n619 161.3
R22322 commonsourceibias.n725 commonsourceibias.n724 161.3
R22323 commonsourceibias.n722 commonsourceibias.n620 161.3
R22324 commonsourceibias.n721 commonsourceibias.n720 161.3
R22325 commonsourceibias.n719 commonsourceibias.n621 161.3
R22326 commonsourceibias.n718 commonsourceibias.n717 161.3
R22327 commonsourceibias.n715 commonsourceibias.n622 161.3
R22328 commonsourceibias.n713 commonsourceibias.n712 161.3
R22329 commonsourceibias.n711 commonsourceibias.n623 161.3
R22330 commonsourceibias.n710 commonsourceibias.n709 161.3
R22331 commonsourceibias.n707 commonsourceibias.n624 161.3
R22332 commonsourceibias.n706 commonsourceibias.n705 161.3
R22333 commonsourceibias.n704 commonsourceibias.n625 161.3
R22334 commonsourceibias.n703 commonsourceibias.n702 161.3
R22335 commonsourceibias.n700 commonsourceibias.n626 161.3
R22336 commonsourceibias.n698 commonsourceibias.n697 161.3
R22337 commonsourceibias.n696 commonsourceibias.n627 161.3
R22338 commonsourceibias.n695 commonsourceibias.n694 161.3
R22339 commonsourceibias.n692 commonsourceibias.n628 161.3
R22340 commonsourceibias.n691 commonsourceibias.n690 161.3
R22341 commonsourceibias.n689 commonsourceibias.n629 161.3
R22342 commonsourceibias.n688 commonsourceibias.n687 161.3
R22343 commonsourceibias.n685 commonsourceibias.n630 161.3
R22344 commonsourceibias.n683 commonsourceibias.n682 161.3
R22345 commonsourceibias.n681 commonsourceibias.n631 161.3
R22346 commonsourceibias.n680 commonsourceibias.n679 161.3
R22347 commonsourceibias.n677 commonsourceibias.n632 161.3
R22348 commonsourceibias.n676 commonsourceibias.n675 161.3
R22349 commonsourceibias.n674 commonsourceibias.n633 161.3
R22350 commonsourceibias.n673 commonsourceibias.n672 161.3
R22351 commonsourceibias.n670 commonsourceibias.n634 161.3
R22352 commonsourceibias.n668 commonsourceibias.n667 161.3
R22353 commonsourceibias.n666 commonsourceibias.n635 161.3
R22354 commonsourceibias.n665 commonsourceibias.n664 161.3
R22355 commonsourceibias.n662 commonsourceibias.n636 161.3
R22356 commonsourceibias.n661 commonsourceibias.n660 161.3
R22357 commonsourceibias.n659 commonsourceibias.n637 161.3
R22358 commonsourceibias.n658 commonsourceibias.n657 161.3
R22359 commonsourceibias.n655 commonsourceibias.n638 161.3
R22360 commonsourceibias.n653 commonsourceibias.n652 161.3
R22361 commonsourceibias.n651 commonsourceibias.n639 161.3
R22362 commonsourceibias.n650 commonsourceibias.n649 161.3
R22363 commonsourceibias.n647 commonsourceibias.n640 161.3
R22364 commonsourceibias.n646 commonsourceibias.n645 161.3
R22365 commonsourceibias.n644 commonsourceibias.n641 161.3
R22366 commonsourceibias.n500 commonsourceibias.n388 161.3
R22367 commonsourceibias.n498 commonsourceibias.n497 161.3
R22368 commonsourceibias.n496 commonsourceibias.n389 161.3
R22369 commonsourceibias.n495 commonsourceibias.n494 161.3
R22370 commonsourceibias.n492 commonsourceibias.n390 161.3
R22371 commonsourceibias.n491 commonsourceibias.n490 161.3
R22372 commonsourceibias.n489 commonsourceibias.n391 161.3
R22373 commonsourceibias.n488 commonsourceibias.n487 161.3
R22374 commonsourceibias.n485 commonsourceibias.n392 161.3
R22375 commonsourceibias.n483 commonsourceibias.n482 161.3
R22376 commonsourceibias.n481 commonsourceibias.n393 161.3
R22377 commonsourceibias.n480 commonsourceibias.n479 161.3
R22378 commonsourceibias.n477 commonsourceibias.n394 161.3
R22379 commonsourceibias.n476 commonsourceibias.n475 161.3
R22380 commonsourceibias.n474 commonsourceibias.n395 161.3
R22381 commonsourceibias.n473 commonsourceibias.n472 161.3
R22382 commonsourceibias.n470 commonsourceibias.n396 161.3
R22383 commonsourceibias.n468 commonsourceibias.n467 161.3
R22384 commonsourceibias.n466 commonsourceibias.n397 161.3
R22385 commonsourceibias.n465 commonsourceibias.n464 161.3
R22386 commonsourceibias.n462 commonsourceibias.n398 161.3
R22387 commonsourceibias.n461 commonsourceibias.n460 161.3
R22388 commonsourceibias.n459 commonsourceibias.n399 161.3
R22389 commonsourceibias.n458 commonsourceibias.n457 161.3
R22390 commonsourceibias.n455 commonsourceibias.n400 161.3
R22391 commonsourceibias.n453 commonsourceibias.n452 161.3
R22392 commonsourceibias.n451 commonsourceibias.n401 161.3
R22393 commonsourceibias.n450 commonsourceibias.n449 161.3
R22394 commonsourceibias.n447 commonsourceibias.n402 161.3
R22395 commonsourceibias.n446 commonsourceibias.n445 161.3
R22396 commonsourceibias.n444 commonsourceibias.n403 161.3
R22397 commonsourceibias.n443 commonsourceibias.n442 161.3
R22398 commonsourceibias.n440 commonsourceibias.n404 161.3
R22399 commonsourceibias.n438 commonsourceibias.n437 161.3
R22400 commonsourceibias.n436 commonsourceibias.n405 161.3
R22401 commonsourceibias.n435 commonsourceibias.n434 161.3
R22402 commonsourceibias.n432 commonsourceibias.n406 161.3
R22403 commonsourceibias.n431 commonsourceibias.n430 161.3
R22404 commonsourceibias.n429 commonsourceibias.n407 161.3
R22405 commonsourceibias.n428 commonsourceibias.n427 161.3
R22406 commonsourceibias.n425 commonsourceibias.n408 161.3
R22407 commonsourceibias.n423 commonsourceibias.n422 161.3
R22408 commonsourceibias.n421 commonsourceibias.n409 161.3
R22409 commonsourceibias.n420 commonsourceibias.n419 161.3
R22410 commonsourceibias.n417 commonsourceibias.n410 161.3
R22411 commonsourceibias.n416 commonsourceibias.n415 161.3
R22412 commonsourceibias.n414 commonsourceibias.n411 161.3
R22413 commonsourceibias.n570 commonsourceibias.n569 161.3
R22414 commonsourceibias.n568 commonsourceibias.n567 161.3
R22415 commonsourceibias.n566 commonsourceibias.n516 161.3
R22416 commonsourceibias.n565 commonsourceibias.n564 161.3
R22417 commonsourceibias.n563 commonsourceibias.n562 161.3
R22418 commonsourceibias.n561 commonsourceibias.n518 161.3
R22419 commonsourceibias.n560 commonsourceibias.n559 161.3
R22420 commonsourceibias.n558 commonsourceibias.n557 161.3
R22421 commonsourceibias.n556 commonsourceibias.n520 161.3
R22422 commonsourceibias.n554 commonsourceibias.n553 161.3
R22423 commonsourceibias.n552 commonsourceibias.n521 161.3
R22424 commonsourceibias.n551 commonsourceibias.n550 161.3
R22425 commonsourceibias.n548 commonsourceibias.n522 161.3
R22426 commonsourceibias.n547 commonsourceibias.n546 161.3
R22427 commonsourceibias.n545 commonsourceibias.n523 161.3
R22428 commonsourceibias.n544 commonsourceibias.n543 161.3
R22429 commonsourceibias.n541 commonsourceibias.n524 161.3
R22430 commonsourceibias.n539 commonsourceibias.n538 161.3
R22431 commonsourceibias.n537 commonsourceibias.n525 161.3
R22432 commonsourceibias.n536 commonsourceibias.n535 161.3
R22433 commonsourceibias.n533 commonsourceibias.n526 161.3
R22434 commonsourceibias.n532 commonsourceibias.n531 161.3
R22435 commonsourceibias.n530 commonsourceibias.n527 161.3
R22436 commonsourceibias.n615 commonsourceibias.n367 161.3
R22437 commonsourceibias.n613 commonsourceibias.n612 161.3
R22438 commonsourceibias.n611 commonsourceibias.n368 161.3
R22439 commonsourceibias.n610 commonsourceibias.n609 161.3
R22440 commonsourceibias.n607 commonsourceibias.n369 161.3
R22441 commonsourceibias.n606 commonsourceibias.n605 161.3
R22442 commonsourceibias.n604 commonsourceibias.n370 161.3
R22443 commonsourceibias.n603 commonsourceibias.n602 161.3
R22444 commonsourceibias.n600 commonsourceibias.n371 161.3
R22445 commonsourceibias.n598 commonsourceibias.n597 161.3
R22446 commonsourceibias.n596 commonsourceibias.n372 161.3
R22447 commonsourceibias.n595 commonsourceibias.n594 161.3
R22448 commonsourceibias.n592 commonsourceibias.n373 161.3
R22449 commonsourceibias.n591 commonsourceibias.n590 161.3
R22450 commonsourceibias.n589 commonsourceibias.n374 161.3
R22451 commonsourceibias.n588 commonsourceibias.n587 161.3
R22452 commonsourceibias.n585 commonsourceibias.n375 161.3
R22453 commonsourceibias.n583 commonsourceibias.n582 161.3
R22454 commonsourceibias.n581 commonsourceibias.n376 161.3
R22455 commonsourceibias.n580 commonsourceibias.n579 161.3
R22456 commonsourceibias.n577 commonsourceibias.n377 161.3
R22457 commonsourceibias.n576 commonsourceibias.n575 161.3
R22458 commonsourceibias.n574 commonsourceibias.n378 161.3
R22459 commonsourceibias.n573 commonsourceibias.n572 161.3
R22460 commonsourceibias.n141 commonsourceibias.n139 81.5057
R22461 commonsourceibias.n381 commonsourceibias.n379 81.5057
R22462 commonsourceibias.n141 commonsourceibias.n140 80.9324
R22463 commonsourceibias.n143 commonsourceibias.n142 80.9324
R22464 commonsourceibias.n145 commonsourceibias.n144 80.9324
R22465 commonsourceibias.n147 commonsourceibias.n146 80.9324
R22466 commonsourceibias.n138 commonsourceibias.n137 80.9324
R22467 commonsourceibias.n136 commonsourceibias.n135 80.9324
R22468 commonsourceibias.n134 commonsourceibias.n133 80.9324
R22469 commonsourceibias.n132 commonsourceibias.n131 80.9324
R22470 commonsourceibias.n130 commonsourceibias.n129 80.9324
R22471 commonsourceibias.n504 commonsourceibias.n503 80.9324
R22472 commonsourceibias.n506 commonsourceibias.n505 80.9324
R22473 commonsourceibias.n508 commonsourceibias.n507 80.9324
R22474 commonsourceibias.n510 commonsourceibias.n509 80.9324
R22475 commonsourceibias.n512 commonsourceibias.n511 80.9324
R22476 commonsourceibias.n387 commonsourceibias.n386 80.9324
R22477 commonsourceibias.n385 commonsourceibias.n384 80.9324
R22478 commonsourceibias.n383 commonsourceibias.n382 80.9324
R22479 commonsourceibias.n381 commonsourceibias.n380 80.9324
R22480 commonsourceibias.n365 commonsourceibias.n364 80.6037
R22481 commonsourceibias.n128 commonsourceibias.n127 80.6037
R22482 commonsourceibias.n250 commonsourceibias.n249 80.6037
R22483 commonsourceibias.n732 commonsourceibias.n731 80.6037
R22484 commonsourceibias.n502 commonsourceibias.n501 80.6037
R22485 commonsourceibias.n617 commonsourceibias.n616 80.6037
R22486 commonsourceibias.n322 commonsourceibias.n321 56.5617
R22487 commonsourceibias.n336 commonsourceibias.n335 56.5617
R22488 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22489 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22490 commonsourceibias.n207 commonsourceibias.n206 56.5617
R22491 commonsourceibias.n193 commonsourceibias.n192 56.5617
R22492 commonsourceibias.n687 commonsourceibias.n685 56.5617
R22493 commonsourceibias.n702 commonsourceibias.n700 56.5617
R22494 commonsourceibias.n457 commonsourceibias.n455 56.5617
R22495 commonsourceibias.n472 commonsourceibias.n470 56.5617
R22496 commonsourceibias.n572 commonsourceibias.n570 56.5617
R22497 commonsourceibias.n294 commonsourceibias.n293 56.5617
R22498 commonsourceibias.n308 commonsourceibias.n307 56.5617
R22499 commonsourceibias.n350 commonsourceibias.n349 56.5617
R22500 commonsourceibias.n113 commonsourceibias.n112 56.5617
R22501 commonsourceibias.n99 commonsourceibias.n98 56.5617
R22502 commonsourceibias.n57 commonsourceibias.n56 56.5617
R22503 commonsourceibias.n235 commonsourceibias.n234 56.5617
R22504 commonsourceibias.n221 commonsourceibias.n220 56.5617
R22505 commonsourceibias.n179 commonsourceibias.n178 56.5617
R22506 commonsourceibias.n657 commonsourceibias.n655 56.5617
R22507 commonsourceibias.n672 commonsourceibias.n670 56.5617
R22508 commonsourceibias.n717 commonsourceibias.n715 56.5617
R22509 commonsourceibias.n427 commonsourceibias.n425 56.5617
R22510 commonsourceibias.n442 commonsourceibias.n440 56.5617
R22511 commonsourceibias.n487 commonsourceibias.n485 56.5617
R22512 commonsourceibias.n602 commonsourceibias.n600 56.5617
R22513 commonsourceibias.n587 commonsourceibias.n585 56.5617
R22514 commonsourceibias.n543 commonsourceibias.n541 56.5617
R22515 commonsourceibias.n557 commonsourceibias.n556 56.5617
R22516 commonsourceibias.n285 commonsourceibias.n284 51.2335
R22517 commonsourceibias.n357 commonsourceibias.n252 51.2335
R22518 commonsourceibias.n120 commonsourceibias.n15 51.2335
R22519 commonsourceibias.n48 commonsourceibias.n47 51.2335
R22520 commonsourceibias.n242 commonsourceibias.n1 51.2335
R22521 commonsourceibias.n170 commonsourceibias.n169 51.2335
R22522 commonsourceibias.n647 commonsourceibias.n646 51.2335
R22523 commonsourceibias.n724 commonsourceibias.n619 51.2335
R22524 commonsourceibias.n417 commonsourceibias.n416 51.2335
R22525 commonsourceibias.n494 commonsourceibias.n389 51.2335
R22526 commonsourceibias.n609 commonsourceibias.n368 51.2335
R22527 commonsourceibias.n533 commonsourceibias.n532 51.2335
R22528 commonsourceibias.n364 commonsourceibias.n363 50.9056
R22529 commonsourceibias.n127 commonsourceibias.n126 50.9056
R22530 commonsourceibias.n249 commonsourceibias.n248 50.9056
R22531 commonsourceibias.n731 commonsourceibias.n730 50.9056
R22532 commonsourceibias.n501 commonsourceibias.n500 50.9056
R22533 commonsourceibias.n616 commonsourceibias.n615 50.9056
R22534 commonsourceibias.n299 commonsourceibias.n298 50.2647
R22535 commonsourceibias.n343 commonsourceibias.n257 50.2647
R22536 commonsourceibias.n106 commonsourceibias.n20 50.2647
R22537 commonsourceibias.n62 commonsourceibias.n61 50.2647
R22538 commonsourceibias.n228 commonsourceibias.n6 50.2647
R22539 commonsourceibias.n184 commonsourceibias.n183 50.2647
R22540 commonsourceibias.n662 commonsourceibias.n661 50.2647
R22541 commonsourceibias.n709 commonsourceibias.n623 50.2647
R22542 commonsourceibias.n432 commonsourceibias.n431 50.2647
R22543 commonsourceibias.n479 commonsourceibias.n393 50.2647
R22544 commonsourceibias.n594 commonsourceibias.n372 50.2647
R22545 commonsourceibias.n548 commonsourceibias.n547 50.2647
R22546 commonsourceibias.n281 commonsourceibias.n280 49.9027
R22547 commonsourceibias.n44 commonsourceibias.n43 49.9027
R22548 commonsourceibias.n166 commonsourceibias.n165 49.9027
R22549 commonsourceibias.n643 commonsourceibias.n642 49.9027
R22550 commonsourceibias.n413 commonsourceibias.n412 49.9027
R22551 commonsourceibias.n529 commonsourceibias.n528 49.9027
R22552 commonsourceibias.n313 commonsourceibias.n312 49.296
R22553 commonsourceibias.n329 commonsourceibias.n262 49.296
R22554 commonsourceibias.n92 commonsourceibias.n25 49.296
R22555 commonsourceibias.n76 commonsourceibias.n75 49.296
R22556 commonsourceibias.n214 commonsourceibias.n11 49.296
R22557 commonsourceibias.n198 commonsourceibias.n197 49.296
R22558 commonsourceibias.n677 commonsourceibias.n676 49.296
R22559 commonsourceibias.n694 commonsourceibias.n627 49.296
R22560 commonsourceibias.n447 commonsourceibias.n446 49.296
R22561 commonsourceibias.n464 commonsourceibias.n397 49.296
R22562 commonsourceibias.n579 commonsourceibias.n376 49.296
R22563 commonsourceibias.n562 commonsourceibias.n561 49.296
R22564 commonsourceibias.n315 commonsourceibias.n267 48.3272
R22565 commonsourceibias.n327 commonsourceibias.n326 48.3272
R22566 commonsourceibias.n90 commonsourceibias.n89 48.3272
R22567 commonsourceibias.n78 commonsourceibias.n30 48.3272
R22568 commonsourceibias.n212 commonsourceibias.n211 48.3272
R22569 commonsourceibias.n202 commonsourceibias.n201 48.3272
R22570 commonsourceibias.n679 commonsourceibias.n631 48.3272
R22571 commonsourceibias.n692 commonsourceibias.n691 48.3272
R22572 commonsourceibias.n449 commonsourceibias.n401 48.3272
R22573 commonsourceibias.n462 commonsourceibias.n461 48.3272
R22574 commonsourceibias.n577 commonsourceibias.n576 48.3272
R22575 commonsourceibias.n566 commonsourceibias.n565 48.3272
R22576 commonsourceibias.n301 commonsourceibias.n272 47.3584
R22577 commonsourceibias.n341 commonsourceibias.n340 47.3584
R22578 commonsourceibias.n104 commonsourceibias.n103 47.3584
R22579 commonsourceibias.n64 commonsourceibias.n35 47.3584
R22580 commonsourceibias.n226 commonsourceibias.n225 47.3584
R22581 commonsourceibias.n186 commonsourceibias.n157 47.3584
R22582 commonsourceibias.n664 commonsourceibias.n635 47.3584
R22583 commonsourceibias.n707 commonsourceibias.n706 47.3584
R22584 commonsourceibias.n434 commonsourceibias.n405 47.3584
R22585 commonsourceibias.n477 commonsourceibias.n476 47.3584
R22586 commonsourceibias.n592 commonsourceibias.n591 47.3584
R22587 commonsourceibias.n550 commonsourceibias.n521 47.3584
R22588 commonsourceibias.n287 commonsourceibias.n277 46.3896
R22589 commonsourceibias.n355 commonsourceibias.n354 46.3896
R22590 commonsourceibias.n118 commonsourceibias.n117 46.3896
R22591 commonsourceibias.n50 commonsourceibias.n40 46.3896
R22592 commonsourceibias.n240 commonsourceibias.n239 46.3896
R22593 commonsourceibias.n172 commonsourceibias.n162 46.3896
R22594 commonsourceibias.n649 commonsourceibias.n639 46.3896
R22595 commonsourceibias.n722 commonsourceibias.n721 46.3896
R22596 commonsourceibias.n419 commonsourceibias.n409 46.3896
R22597 commonsourceibias.n492 commonsourceibias.n491 46.3896
R22598 commonsourceibias.n607 commonsourceibias.n606 46.3896
R22599 commonsourceibias.n535 commonsourceibias.n525 46.3896
R22600 commonsourceibias.n282 commonsourceibias.n281 44.7059
R22601 commonsourceibias.n644 commonsourceibias.n643 44.7059
R22602 commonsourceibias.n414 commonsourceibias.n413 44.7059
R22603 commonsourceibias.n530 commonsourceibias.n529 44.7059
R22604 commonsourceibias.n45 commonsourceibias.n44 44.7059
R22605 commonsourceibias.n167 commonsourceibias.n166 44.7059
R22606 commonsourceibias.n291 commonsourceibias.n277 34.7644
R22607 commonsourceibias.n354 commonsourceibias.n254 34.7644
R22608 commonsourceibias.n117 commonsourceibias.n17 34.7644
R22609 commonsourceibias.n54 commonsourceibias.n40 34.7644
R22610 commonsourceibias.n239 commonsourceibias.n3 34.7644
R22611 commonsourceibias.n176 commonsourceibias.n162 34.7644
R22612 commonsourceibias.n653 commonsourceibias.n639 34.7644
R22613 commonsourceibias.n721 commonsourceibias.n621 34.7644
R22614 commonsourceibias.n423 commonsourceibias.n409 34.7644
R22615 commonsourceibias.n491 commonsourceibias.n391 34.7644
R22616 commonsourceibias.n606 commonsourceibias.n370 34.7644
R22617 commonsourceibias.n539 commonsourceibias.n525 34.7644
R22618 commonsourceibias.n305 commonsourceibias.n272 33.7956
R22619 commonsourceibias.n340 commonsourceibias.n259 33.7956
R22620 commonsourceibias.n103 commonsourceibias.n22 33.7956
R22621 commonsourceibias.n68 commonsourceibias.n35 33.7956
R22622 commonsourceibias.n225 commonsourceibias.n8 33.7956
R22623 commonsourceibias.n190 commonsourceibias.n157 33.7956
R22624 commonsourceibias.n668 commonsourceibias.n635 33.7956
R22625 commonsourceibias.n706 commonsourceibias.n625 33.7956
R22626 commonsourceibias.n438 commonsourceibias.n405 33.7956
R22627 commonsourceibias.n476 commonsourceibias.n395 33.7956
R22628 commonsourceibias.n591 commonsourceibias.n374 33.7956
R22629 commonsourceibias.n554 commonsourceibias.n521 33.7956
R22630 commonsourceibias.n319 commonsourceibias.n267 32.8269
R22631 commonsourceibias.n326 commonsourceibias.n264 32.8269
R22632 commonsourceibias.n89 commonsourceibias.n27 32.8269
R22633 commonsourceibias.n82 commonsourceibias.n30 32.8269
R22634 commonsourceibias.n211 commonsourceibias.n13 32.8269
R22635 commonsourceibias.n203 commonsourceibias.n202 32.8269
R22636 commonsourceibias.n683 commonsourceibias.n631 32.8269
R22637 commonsourceibias.n691 commonsourceibias.n629 32.8269
R22638 commonsourceibias.n453 commonsourceibias.n401 32.8269
R22639 commonsourceibias.n461 commonsourceibias.n399 32.8269
R22640 commonsourceibias.n576 commonsourceibias.n378 32.8269
R22641 commonsourceibias.n567 commonsourceibias.n566 32.8269
R22642 commonsourceibias.n312 commonsourceibias.n269 31.8581
R22643 commonsourceibias.n333 commonsourceibias.n262 31.8581
R22644 commonsourceibias.n96 commonsourceibias.n25 31.8581
R22645 commonsourceibias.n75 commonsourceibias.n32 31.8581
R22646 commonsourceibias.n218 commonsourceibias.n11 31.8581
R22647 commonsourceibias.n197 commonsourceibias.n196 31.8581
R22648 commonsourceibias.n676 commonsourceibias.n633 31.8581
R22649 commonsourceibias.n698 commonsourceibias.n627 31.8581
R22650 commonsourceibias.n446 commonsourceibias.n403 31.8581
R22651 commonsourceibias.n468 commonsourceibias.n397 31.8581
R22652 commonsourceibias.n583 commonsourceibias.n376 31.8581
R22653 commonsourceibias.n561 commonsourceibias.n560 31.8581
R22654 commonsourceibias.n298 commonsourceibias.n274 30.8893
R22655 commonsourceibias.n347 commonsourceibias.n257 30.8893
R22656 commonsourceibias.n110 commonsourceibias.n20 30.8893
R22657 commonsourceibias.n61 commonsourceibias.n37 30.8893
R22658 commonsourceibias.n232 commonsourceibias.n6 30.8893
R22659 commonsourceibias.n183 commonsourceibias.n159 30.8893
R22660 commonsourceibias.n661 commonsourceibias.n637 30.8893
R22661 commonsourceibias.n713 commonsourceibias.n623 30.8893
R22662 commonsourceibias.n431 commonsourceibias.n407 30.8893
R22663 commonsourceibias.n483 commonsourceibias.n393 30.8893
R22664 commonsourceibias.n598 commonsourceibias.n372 30.8893
R22665 commonsourceibias.n547 commonsourceibias.n523 30.8893
R22666 commonsourceibias.n284 commonsourceibias.n279 29.9206
R22667 commonsourceibias.n361 commonsourceibias.n252 29.9206
R22668 commonsourceibias.n124 commonsourceibias.n15 29.9206
R22669 commonsourceibias.n47 commonsourceibias.n42 29.9206
R22670 commonsourceibias.n246 commonsourceibias.n1 29.9206
R22671 commonsourceibias.n169 commonsourceibias.n164 29.9206
R22672 commonsourceibias.n646 commonsourceibias.n641 29.9206
R22673 commonsourceibias.n728 commonsourceibias.n619 29.9206
R22674 commonsourceibias.n416 commonsourceibias.n411 29.9206
R22675 commonsourceibias.n498 commonsourceibias.n389 29.9206
R22676 commonsourceibias.n613 commonsourceibias.n368 29.9206
R22677 commonsourceibias.n532 commonsourceibias.n527 29.9206
R22678 commonsourceibias.n363 commonsourceibias.n362 21.8872
R22679 commonsourceibias.n126 commonsourceibias.n125 21.8872
R22680 commonsourceibias.n248 commonsourceibias.n247 21.8872
R22681 commonsourceibias.n730 commonsourceibias.n729 21.8872
R22682 commonsourceibias.n500 commonsourceibias.n499 21.8872
R22683 commonsourceibias.n615 commonsourceibias.n614 21.8872
R22684 commonsourceibias.n294 commonsourceibias.n276 21.3954
R22685 commonsourceibias.n349 commonsourceibias.n348 21.3954
R22686 commonsourceibias.n112 commonsourceibias.n111 21.3954
R22687 commonsourceibias.n57 commonsourceibias.n39 21.3954
R22688 commonsourceibias.n234 commonsourceibias.n233 21.3954
R22689 commonsourceibias.n179 commonsourceibias.n161 21.3954
R22690 commonsourceibias.n657 commonsourceibias.n656 21.3954
R22691 commonsourceibias.n715 commonsourceibias.n714 21.3954
R22692 commonsourceibias.n427 commonsourceibias.n426 21.3954
R22693 commonsourceibias.n485 commonsourceibias.n484 21.3954
R22694 commonsourceibias.n600 commonsourceibias.n599 21.3954
R22695 commonsourceibias.n543 commonsourceibias.n542 21.3954
R22696 commonsourceibias.n308 commonsourceibias.n271 20.9036
R22697 commonsourceibias.n335 commonsourceibias.n334 20.9036
R22698 commonsourceibias.n98 commonsourceibias.n97 20.9036
R22699 commonsourceibias.n71 commonsourceibias.n34 20.9036
R22700 commonsourceibias.n220 commonsourceibias.n219 20.9036
R22701 commonsourceibias.n193 commonsourceibias.n155 20.9036
R22702 commonsourceibias.n672 commonsourceibias.n671 20.9036
R22703 commonsourceibias.n700 commonsourceibias.n699 20.9036
R22704 commonsourceibias.n442 commonsourceibias.n441 20.9036
R22705 commonsourceibias.n470 commonsourceibias.n469 20.9036
R22706 commonsourceibias.n585 commonsourceibias.n584 20.9036
R22707 commonsourceibias.n557 commonsourceibias.n519 20.9036
R22708 commonsourceibias.n321 commonsourceibias.n320 20.4117
R22709 commonsourceibias.n322 commonsourceibias.n266 20.4117
R22710 commonsourceibias.n85 commonsourceibias.n29 20.4117
R22711 commonsourceibias.n84 commonsourceibias.n83 20.4117
R22712 commonsourceibias.n207 commonsourceibias.n150 20.4117
R22713 commonsourceibias.n206 commonsourceibias.n151 20.4117
R22714 commonsourceibias.n685 commonsourceibias.n684 20.4117
R22715 commonsourceibias.n687 commonsourceibias.n686 20.4117
R22716 commonsourceibias.n455 commonsourceibias.n454 20.4117
R22717 commonsourceibias.n457 commonsourceibias.n456 20.4117
R22718 commonsourceibias.n572 commonsourceibias.n571 20.4117
R22719 commonsourceibias.n570 commonsourceibias.n515 20.4117
R22720 commonsourceibias.n307 commonsourceibias.n306 19.9199
R22721 commonsourceibias.n336 commonsourceibias.n261 19.9199
R22722 commonsourceibias.n99 commonsourceibias.n24 19.9199
R22723 commonsourceibias.n70 commonsourceibias.n69 19.9199
R22724 commonsourceibias.n221 commonsourceibias.n10 19.9199
R22725 commonsourceibias.n192 commonsourceibias.n191 19.9199
R22726 commonsourceibias.n670 commonsourceibias.n669 19.9199
R22727 commonsourceibias.n702 commonsourceibias.n701 19.9199
R22728 commonsourceibias.n440 commonsourceibias.n439 19.9199
R22729 commonsourceibias.n472 commonsourceibias.n471 19.9199
R22730 commonsourceibias.n587 commonsourceibias.n586 19.9199
R22731 commonsourceibias.n556 commonsourceibias.n555 19.9199
R22732 commonsourceibias.n293 commonsourceibias.n292 19.4281
R22733 commonsourceibias.n350 commonsourceibias.n256 19.4281
R22734 commonsourceibias.n113 commonsourceibias.n19 19.4281
R22735 commonsourceibias.n56 commonsourceibias.n55 19.4281
R22736 commonsourceibias.n235 commonsourceibias.n5 19.4281
R22737 commonsourceibias.n178 commonsourceibias.n177 19.4281
R22738 commonsourceibias.n655 commonsourceibias.n654 19.4281
R22739 commonsourceibias.n717 commonsourceibias.n716 19.4281
R22740 commonsourceibias.n425 commonsourceibias.n424 19.4281
R22741 commonsourceibias.n487 commonsourceibias.n486 19.4281
R22742 commonsourceibias.n602 commonsourceibias.n601 19.4281
R22743 commonsourceibias.n541 commonsourceibias.n540 19.4281
R22744 commonsourceibias.n286 commonsourceibias.n285 13.526
R22745 commonsourceibias.n357 commonsourceibias.n356 13.526
R22746 commonsourceibias.n120 commonsourceibias.n119 13.526
R22747 commonsourceibias.n49 commonsourceibias.n48 13.526
R22748 commonsourceibias.n242 commonsourceibias.n241 13.526
R22749 commonsourceibias.n171 commonsourceibias.n170 13.526
R22750 commonsourceibias.n648 commonsourceibias.n647 13.526
R22751 commonsourceibias.n724 commonsourceibias.n723 13.526
R22752 commonsourceibias.n418 commonsourceibias.n417 13.526
R22753 commonsourceibias.n494 commonsourceibias.n493 13.526
R22754 commonsourceibias.n609 commonsourceibias.n608 13.526
R22755 commonsourceibias.n534 commonsourceibias.n533 13.526
R22756 commonsourceibias.n130 commonsourceibias.n128 13.2322
R22757 commonsourceibias.n504 commonsourceibias.n502 13.2322
R22758 commonsourceibias.n300 commonsourceibias.n299 13.0342
R22759 commonsourceibias.n343 commonsourceibias.n342 13.0342
R22760 commonsourceibias.n106 commonsourceibias.n105 13.0342
R22761 commonsourceibias.n63 commonsourceibias.n62 13.0342
R22762 commonsourceibias.n228 commonsourceibias.n227 13.0342
R22763 commonsourceibias.n185 commonsourceibias.n184 13.0342
R22764 commonsourceibias.n663 commonsourceibias.n662 13.0342
R22765 commonsourceibias.n709 commonsourceibias.n708 13.0342
R22766 commonsourceibias.n433 commonsourceibias.n432 13.0342
R22767 commonsourceibias.n479 commonsourceibias.n478 13.0342
R22768 commonsourceibias.n594 commonsourceibias.n593 13.0342
R22769 commonsourceibias.n549 commonsourceibias.n548 13.0342
R22770 commonsourceibias.n314 commonsourceibias.n313 12.5423
R22771 commonsourceibias.n329 commonsourceibias.n328 12.5423
R22772 commonsourceibias.n92 commonsourceibias.n91 12.5423
R22773 commonsourceibias.n77 commonsourceibias.n76 12.5423
R22774 commonsourceibias.n214 commonsourceibias.n213 12.5423
R22775 commonsourceibias.n198 commonsourceibias.n153 12.5423
R22776 commonsourceibias.n678 commonsourceibias.n677 12.5423
R22777 commonsourceibias.n694 commonsourceibias.n693 12.5423
R22778 commonsourceibias.n448 commonsourceibias.n447 12.5423
R22779 commonsourceibias.n464 commonsourceibias.n463 12.5423
R22780 commonsourceibias.n579 commonsourceibias.n578 12.5423
R22781 commonsourceibias.n562 commonsourceibias.n517 12.5423
R22782 commonsourceibias.n734 commonsourceibias.n366 12.2777
R22783 commonsourceibias.n315 commonsourceibias.n314 12.0505
R22784 commonsourceibias.n328 commonsourceibias.n327 12.0505
R22785 commonsourceibias.n91 commonsourceibias.n90 12.0505
R22786 commonsourceibias.n78 commonsourceibias.n77 12.0505
R22787 commonsourceibias.n213 commonsourceibias.n212 12.0505
R22788 commonsourceibias.n201 commonsourceibias.n153 12.0505
R22789 commonsourceibias.n679 commonsourceibias.n678 12.0505
R22790 commonsourceibias.n693 commonsourceibias.n692 12.0505
R22791 commonsourceibias.n449 commonsourceibias.n448 12.0505
R22792 commonsourceibias.n463 commonsourceibias.n462 12.0505
R22793 commonsourceibias.n578 commonsourceibias.n577 12.0505
R22794 commonsourceibias.n565 commonsourceibias.n517 12.0505
R22795 commonsourceibias.n301 commonsourceibias.n300 11.5587
R22796 commonsourceibias.n342 commonsourceibias.n341 11.5587
R22797 commonsourceibias.n105 commonsourceibias.n104 11.5587
R22798 commonsourceibias.n64 commonsourceibias.n63 11.5587
R22799 commonsourceibias.n227 commonsourceibias.n226 11.5587
R22800 commonsourceibias.n186 commonsourceibias.n185 11.5587
R22801 commonsourceibias.n664 commonsourceibias.n663 11.5587
R22802 commonsourceibias.n708 commonsourceibias.n707 11.5587
R22803 commonsourceibias.n434 commonsourceibias.n433 11.5587
R22804 commonsourceibias.n478 commonsourceibias.n477 11.5587
R22805 commonsourceibias.n593 commonsourceibias.n592 11.5587
R22806 commonsourceibias.n550 commonsourceibias.n549 11.5587
R22807 commonsourceibias.n287 commonsourceibias.n286 11.0668
R22808 commonsourceibias.n356 commonsourceibias.n355 11.0668
R22809 commonsourceibias.n119 commonsourceibias.n118 11.0668
R22810 commonsourceibias.n50 commonsourceibias.n49 11.0668
R22811 commonsourceibias.n241 commonsourceibias.n240 11.0668
R22812 commonsourceibias.n172 commonsourceibias.n171 11.0668
R22813 commonsourceibias.n649 commonsourceibias.n648 11.0668
R22814 commonsourceibias.n723 commonsourceibias.n722 11.0668
R22815 commonsourceibias.n419 commonsourceibias.n418 11.0668
R22816 commonsourceibias.n493 commonsourceibias.n492 11.0668
R22817 commonsourceibias.n608 commonsourceibias.n607 11.0668
R22818 commonsourceibias.n535 commonsourceibias.n534 11.0668
R22819 commonsourceibias.n734 commonsourceibias.n733 10.3347
R22820 commonsourceibias.n149 commonsourceibias.n148 9.50363
R22821 commonsourceibias.n514 commonsourceibias.n513 9.50363
R22822 commonsourceibias.n366 commonsourceibias.n250 8.75852
R22823 commonsourceibias.n733 commonsourceibias.n617 8.75852
R22824 commonsourceibias.n292 commonsourceibias.n291 5.16479
R22825 commonsourceibias.n256 commonsourceibias.n254 5.16479
R22826 commonsourceibias.n19 commonsourceibias.n17 5.16479
R22827 commonsourceibias.n55 commonsourceibias.n54 5.16479
R22828 commonsourceibias.n5 commonsourceibias.n3 5.16479
R22829 commonsourceibias.n177 commonsourceibias.n176 5.16479
R22830 commonsourceibias.n654 commonsourceibias.n653 5.16479
R22831 commonsourceibias.n716 commonsourceibias.n621 5.16479
R22832 commonsourceibias.n424 commonsourceibias.n423 5.16479
R22833 commonsourceibias.n486 commonsourceibias.n391 5.16479
R22834 commonsourceibias.n601 commonsourceibias.n370 5.16479
R22835 commonsourceibias.n540 commonsourceibias.n539 5.16479
R22836 commonsourceibias.n366 commonsourceibias.n365 5.03125
R22837 commonsourceibias.n733 commonsourceibias.n732 5.03125
R22838 commonsourceibias.n306 commonsourceibias.n305 4.67295
R22839 commonsourceibias.n261 commonsourceibias.n259 4.67295
R22840 commonsourceibias.n24 commonsourceibias.n22 4.67295
R22841 commonsourceibias.n69 commonsourceibias.n68 4.67295
R22842 commonsourceibias.n10 commonsourceibias.n8 4.67295
R22843 commonsourceibias.n191 commonsourceibias.n190 4.67295
R22844 commonsourceibias.n669 commonsourceibias.n668 4.67295
R22845 commonsourceibias.n701 commonsourceibias.n625 4.67295
R22846 commonsourceibias.n439 commonsourceibias.n438 4.67295
R22847 commonsourceibias.n471 commonsourceibias.n395 4.67295
R22848 commonsourceibias.n586 commonsourceibias.n374 4.67295
R22849 commonsourceibias.n555 commonsourceibias.n554 4.67295
R22850 commonsourceibias commonsourceibias.n734 4.20978
R22851 commonsourceibias.n320 commonsourceibias.n319 4.18111
R22852 commonsourceibias.n266 commonsourceibias.n264 4.18111
R22853 commonsourceibias.n29 commonsourceibias.n27 4.18111
R22854 commonsourceibias.n83 commonsourceibias.n82 4.18111
R22855 commonsourceibias.n150 commonsourceibias.n13 4.18111
R22856 commonsourceibias.n203 commonsourceibias.n151 4.18111
R22857 commonsourceibias.n684 commonsourceibias.n683 4.18111
R22858 commonsourceibias.n686 commonsourceibias.n629 4.18111
R22859 commonsourceibias.n454 commonsourceibias.n453 4.18111
R22860 commonsourceibias.n456 commonsourceibias.n399 4.18111
R22861 commonsourceibias.n571 commonsourceibias.n378 4.18111
R22862 commonsourceibias.n567 commonsourceibias.n515 4.18111
R22863 commonsourceibias.n271 commonsourceibias.n269 3.68928
R22864 commonsourceibias.n334 commonsourceibias.n333 3.68928
R22865 commonsourceibias.n97 commonsourceibias.n96 3.68928
R22866 commonsourceibias.n34 commonsourceibias.n32 3.68928
R22867 commonsourceibias.n219 commonsourceibias.n218 3.68928
R22868 commonsourceibias.n196 commonsourceibias.n155 3.68928
R22869 commonsourceibias.n671 commonsourceibias.n633 3.68928
R22870 commonsourceibias.n699 commonsourceibias.n698 3.68928
R22871 commonsourceibias.n441 commonsourceibias.n403 3.68928
R22872 commonsourceibias.n469 commonsourceibias.n468 3.68928
R22873 commonsourceibias.n584 commonsourceibias.n583 3.68928
R22874 commonsourceibias.n560 commonsourceibias.n519 3.68928
R22875 commonsourceibias.n276 commonsourceibias.n274 3.19744
R22876 commonsourceibias.n348 commonsourceibias.n347 3.19744
R22877 commonsourceibias.n111 commonsourceibias.n110 3.19744
R22878 commonsourceibias.n39 commonsourceibias.n37 3.19744
R22879 commonsourceibias.n233 commonsourceibias.n232 3.19744
R22880 commonsourceibias.n161 commonsourceibias.n159 3.19744
R22881 commonsourceibias.n656 commonsourceibias.n637 3.19744
R22882 commonsourceibias.n714 commonsourceibias.n713 3.19744
R22883 commonsourceibias.n426 commonsourceibias.n407 3.19744
R22884 commonsourceibias.n484 commonsourceibias.n483 3.19744
R22885 commonsourceibias.n599 commonsourceibias.n598 3.19744
R22886 commonsourceibias.n542 commonsourceibias.n523 3.19744
R22887 commonsourceibias.n139 commonsourceibias.t47 2.82907
R22888 commonsourceibias.n139 commonsourceibias.t79 2.82907
R22889 commonsourceibias.n140 commonsourceibias.t55 2.82907
R22890 commonsourceibias.n140 commonsourceibias.t5 2.82907
R22891 commonsourceibias.n142 commonsourceibias.t19 2.82907
R22892 commonsourceibias.n142 commonsourceibias.t23 2.82907
R22893 commonsourceibias.n144 commonsourceibias.t39 2.82907
R22894 commonsourceibias.n144 commonsourceibias.t71 2.82907
R22895 commonsourceibias.n146 commonsourceibias.t57 2.82907
R22896 commonsourceibias.n146 commonsourceibias.t27 2.82907
R22897 commonsourceibias.n137 commonsourceibias.t11 2.82907
R22898 commonsourceibias.n137 commonsourceibias.t41 2.82907
R22899 commonsourceibias.n135 commonsourceibias.t25 2.82907
R22900 commonsourceibias.n135 commonsourceibias.t35 2.82907
R22901 commonsourceibias.n133 commonsourceibias.t37 2.82907
R22902 commonsourceibias.n133 commonsourceibias.t77 2.82907
R22903 commonsourceibias.n131 commonsourceibias.t51 2.82907
R22904 commonsourceibias.n131 commonsourceibias.t9 2.82907
R22905 commonsourceibias.n129 commonsourceibias.t75 2.82907
R22906 commonsourceibias.n129 commonsourceibias.t21 2.82907
R22907 commonsourceibias.n503 commonsourceibias.t43 2.82907
R22908 commonsourceibias.n503 commonsourceibias.t15 2.82907
R22909 commonsourceibias.n505 commonsourceibias.t31 2.82907
R22910 commonsourceibias.n505 commonsourceibias.t1 2.82907
R22911 commonsourceibias.n507 commonsourceibias.t17 2.82907
R22912 commonsourceibias.n507 commonsourceibias.t61 2.82907
R22913 commonsourceibias.n509 commonsourceibias.t59 2.82907
R22914 commonsourceibias.n509 commonsourceibias.t45 2.82907
R22915 commonsourceibias.n511 commonsourceibias.t65 2.82907
R22916 commonsourceibias.n511 commonsourceibias.t33 2.82907
R22917 commonsourceibias.n386 commonsourceibias.t53 2.82907
R22918 commonsourceibias.n386 commonsourceibias.t73 2.82907
R22919 commonsourceibias.n384 commonsourceibias.t7 2.82907
R22920 commonsourceibias.n384 commonsourceibias.t63 2.82907
R22921 commonsourceibias.n382 commonsourceibias.t69 2.82907
R22922 commonsourceibias.n382 commonsourceibias.t67 2.82907
R22923 commonsourceibias.n380 commonsourceibias.t49 2.82907
R22924 commonsourceibias.n380 commonsourceibias.t13 2.82907
R22925 commonsourceibias.n379 commonsourceibias.t29 2.82907
R22926 commonsourceibias.n379 commonsourceibias.t3 2.82907
R22927 commonsourceibias.n280 commonsourceibias.n279 2.7056
R22928 commonsourceibias.n362 commonsourceibias.n361 2.7056
R22929 commonsourceibias.n125 commonsourceibias.n124 2.7056
R22930 commonsourceibias.n43 commonsourceibias.n42 2.7056
R22931 commonsourceibias.n247 commonsourceibias.n246 2.7056
R22932 commonsourceibias.n165 commonsourceibias.n164 2.7056
R22933 commonsourceibias.n642 commonsourceibias.n641 2.7056
R22934 commonsourceibias.n729 commonsourceibias.n728 2.7056
R22935 commonsourceibias.n412 commonsourceibias.n411 2.7056
R22936 commonsourceibias.n499 commonsourceibias.n498 2.7056
R22937 commonsourceibias.n614 commonsourceibias.n613 2.7056
R22938 commonsourceibias.n528 commonsourceibias.n527 2.7056
R22939 commonsourceibias.n132 commonsourceibias.n130 0.573776
R22940 commonsourceibias.n134 commonsourceibias.n132 0.573776
R22941 commonsourceibias.n136 commonsourceibias.n134 0.573776
R22942 commonsourceibias.n138 commonsourceibias.n136 0.573776
R22943 commonsourceibias.n147 commonsourceibias.n145 0.573776
R22944 commonsourceibias.n145 commonsourceibias.n143 0.573776
R22945 commonsourceibias.n143 commonsourceibias.n141 0.573776
R22946 commonsourceibias.n383 commonsourceibias.n381 0.573776
R22947 commonsourceibias.n385 commonsourceibias.n383 0.573776
R22948 commonsourceibias.n387 commonsourceibias.n385 0.573776
R22949 commonsourceibias.n512 commonsourceibias.n510 0.573776
R22950 commonsourceibias.n510 commonsourceibias.n508 0.573776
R22951 commonsourceibias.n508 commonsourceibias.n506 0.573776
R22952 commonsourceibias.n506 commonsourceibias.n504 0.573776
R22953 commonsourceibias.n148 commonsourceibias.n138 0.287138
R22954 commonsourceibias.n148 commonsourceibias.n147 0.287138
R22955 commonsourceibias.n513 commonsourceibias.n387 0.287138
R22956 commonsourceibias.n513 commonsourceibias.n512 0.287138
R22957 commonsourceibias.n365 commonsourceibias.n251 0.285035
R22958 commonsourceibias.n128 commonsourceibias.n14 0.285035
R22959 commonsourceibias.n250 commonsourceibias.n0 0.285035
R22960 commonsourceibias.n732 commonsourceibias.n618 0.285035
R22961 commonsourceibias.n502 commonsourceibias.n388 0.285035
R22962 commonsourceibias.n617 commonsourceibias.n367 0.285035
R22963 commonsourceibias.n360 commonsourceibias.n251 0.189894
R22964 commonsourceibias.n360 commonsourceibias.n359 0.189894
R22965 commonsourceibias.n359 commonsourceibias.n358 0.189894
R22966 commonsourceibias.n358 commonsourceibias.n253 0.189894
R22967 commonsourceibias.n353 commonsourceibias.n253 0.189894
R22968 commonsourceibias.n353 commonsourceibias.n352 0.189894
R22969 commonsourceibias.n352 commonsourceibias.n351 0.189894
R22970 commonsourceibias.n351 commonsourceibias.n255 0.189894
R22971 commonsourceibias.n346 commonsourceibias.n255 0.189894
R22972 commonsourceibias.n346 commonsourceibias.n345 0.189894
R22973 commonsourceibias.n345 commonsourceibias.n344 0.189894
R22974 commonsourceibias.n344 commonsourceibias.n258 0.189894
R22975 commonsourceibias.n339 commonsourceibias.n258 0.189894
R22976 commonsourceibias.n339 commonsourceibias.n338 0.189894
R22977 commonsourceibias.n338 commonsourceibias.n337 0.189894
R22978 commonsourceibias.n337 commonsourceibias.n260 0.189894
R22979 commonsourceibias.n332 commonsourceibias.n260 0.189894
R22980 commonsourceibias.n332 commonsourceibias.n331 0.189894
R22981 commonsourceibias.n331 commonsourceibias.n330 0.189894
R22982 commonsourceibias.n330 commonsourceibias.n263 0.189894
R22983 commonsourceibias.n325 commonsourceibias.n263 0.189894
R22984 commonsourceibias.n325 commonsourceibias.n324 0.189894
R22985 commonsourceibias.n324 commonsourceibias.n323 0.189894
R22986 commonsourceibias.n323 commonsourceibias.n265 0.189894
R22987 commonsourceibias.n318 commonsourceibias.n265 0.189894
R22988 commonsourceibias.n318 commonsourceibias.n317 0.189894
R22989 commonsourceibias.n317 commonsourceibias.n316 0.189894
R22990 commonsourceibias.n316 commonsourceibias.n268 0.189894
R22991 commonsourceibias.n311 commonsourceibias.n268 0.189894
R22992 commonsourceibias.n311 commonsourceibias.n310 0.189894
R22993 commonsourceibias.n310 commonsourceibias.n309 0.189894
R22994 commonsourceibias.n309 commonsourceibias.n270 0.189894
R22995 commonsourceibias.n304 commonsourceibias.n270 0.189894
R22996 commonsourceibias.n304 commonsourceibias.n303 0.189894
R22997 commonsourceibias.n303 commonsourceibias.n302 0.189894
R22998 commonsourceibias.n302 commonsourceibias.n273 0.189894
R22999 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23000 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23001 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23002 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23003 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23004 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23005 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23006 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23007 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23008 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23009 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23010 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23011 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23012 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23013 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23014 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23015 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23016 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23017 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23018 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23019 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23020 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23021 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23022 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23023 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23024 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23025 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23026 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23027 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23028 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23029 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23030 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23031 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23032 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23033 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23034 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23035 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23036 commonsourceibias.n79 commonsourceibias.n31 0.189894
R23037 commonsourceibias.n74 commonsourceibias.n31 0.189894
R23038 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23039 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23040 commonsourceibias.n72 commonsourceibias.n33 0.189894
R23041 commonsourceibias.n67 commonsourceibias.n33 0.189894
R23042 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23043 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23044 commonsourceibias.n65 commonsourceibias.n36 0.189894
R23045 commonsourceibias.n60 commonsourceibias.n36 0.189894
R23046 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23047 commonsourceibias.n59 commonsourceibias.n58 0.189894
R23048 commonsourceibias.n58 commonsourceibias.n38 0.189894
R23049 commonsourceibias.n53 commonsourceibias.n38 0.189894
R23050 commonsourceibias.n53 commonsourceibias.n52 0.189894
R23051 commonsourceibias.n52 commonsourceibias.n51 0.189894
R23052 commonsourceibias.n51 commonsourceibias.n41 0.189894
R23053 commonsourceibias.n46 commonsourceibias.n41 0.189894
R23054 commonsourceibias.n46 commonsourceibias.n45 0.189894
R23055 commonsourceibias.n205 commonsourceibias.n204 0.189894
R23056 commonsourceibias.n204 commonsourceibias.n152 0.189894
R23057 commonsourceibias.n200 commonsourceibias.n152 0.189894
R23058 commonsourceibias.n200 commonsourceibias.n199 0.189894
R23059 commonsourceibias.n199 commonsourceibias.n154 0.189894
R23060 commonsourceibias.n195 commonsourceibias.n154 0.189894
R23061 commonsourceibias.n195 commonsourceibias.n194 0.189894
R23062 commonsourceibias.n194 commonsourceibias.n156 0.189894
R23063 commonsourceibias.n189 commonsourceibias.n156 0.189894
R23064 commonsourceibias.n189 commonsourceibias.n188 0.189894
R23065 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23066 commonsourceibias.n187 commonsourceibias.n158 0.189894
R23067 commonsourceibias.n182 commonsourceibias.n158 0.189894
R23068 commonsourceibias.n182 commonsourceibias.n181 0.189894
R23069 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23070 commonsourceibias.n180 commonsourceibias.n160 0.189894
R23071 commonsourceibias.n175 commonsourceibias.n160 0.189894
R23072 commonsourceibias.n175 commonsourceibias.n174 0.189894
R23073 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23074 commonsourceibias.n173 commonsourceibias.n163 0.189894
R23075 commonsourceibias.n168 commonsourceibias.n163 0.189894
R23076 commonsourceibias.n168 commonsourceibias.n167 0.189894
R23077 commonsourceibias.n245 commonsourceibias.n0 0.189894
R23078 commonsourceibias.n245 commonsourceibias.n244 0.189894
R23079 commonsourceibias.n244 commonsourceibias.n243 0.189894
R23080 commonsourceibias.n243 commonsourceibias.n2 0.189894
R23081 commonsourceibias.n238 commonsourceibias.n2 0.189894
R23082 commonsourceibias.n238 commonsourceibias.n237 0.189894
R23083 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23084 commonsourceibias.n236 commonsourceibias.n4 0.189894
R23085 commonsourceibias.n231 commonsourceibias.n4 0.189894
R23086 commonsourceibias.n231 commonsourceibias.n230 0.189894
R23087 commonsourceibias.n230 commonsourceibias.n229 0.189894
R23088 commonsourceibias.n229 commonsourceibias.n7 0.189894
R23089 commonsourceibias.n224 commonsourceibias.n7 0.189894
R23090 commonsourceibias.n224 commonsourceibias.n223 0.189894
R23091 commonsourceibias.n223 commonsourceibias.n222 0.189894
R23092 commonsourceibias.n222 commonsourceibias.n9 0.189894
R23093 commonsourceibias.n217 commonsourceibias.n9 0.189894
R23094 commonsourceibias.n217 commonsourceibias.n216 0.189894
R23095 commonsourceibias.n216 commonsourceibias.n215 0.189894
R23096 commonsourceibias.n215 commonsourceibias.n12 0.189894
R23097 commonsourceibias.n210 commonsourceibias.n12 0.189894
R23098 commonsourceibias.n210 commonsourceibias.n209 0.189894
R23099 commonsourceibias.n209 commonsourceibias.n208 0.189894
R23100 commonsourceibias.n645 commonsourceibias.n644 0.189894
R23101 commonsourceibias.n645 commonsourceibias.n640 0.189894
R23102 commonsourceibias.n650 commonsourceibias.n640 0.189894
R23103 commonsourceibias.n651 commonsourceibias.n650 0.189894
R23104 commonsourceibias.n652 commonsourceibias.n651 0.189894
R23105 commonsourceibias.n652 commonsourceibias.n638 0.189894
R23106 commonsourceibias.n658 commonsourceibias.n638 0.189894
R23107 commonsourceibias.n659 commonsourceibias.n658 0.189894
R23108 commonsourceibias.n660 commonsourceibias.n659 0.189894
R23109 commonsourceibias.n660 commonsourceibias.n636 0.189894
R23110 commonsourceibias.n665 commonsourceibias.n636 0.189894
R23111 commonsourceibias.n666 commonsourceibias.n665 0.189894
R23112 commonsourceibias.n667 commonsourceibias.n666 0.189894
R23113 commonsourceibias.n667 commonsourceibias.n634 0.189894
R23114 commonsourceibias.n673 commonsourceibias.n634 0.189894
R23115 commonsourceibias.n674 commonsourceibias.n673 0.189894
R23116 commonsourceibias.n675 commonsourceibias.n674 0.189894
R23117 commonsourceibias.n675 commonsourceibias.n632 0.189894
R23118 commonsourceibias.n680 commonsourceibias.n632 0.189894
R23119 commonsourceibias.n681 commonsourceibias.n680 0.189894
R23120 commonsourceibias.n682 commonsourceibias.n681 0.189894
R23121 commonsourceibias.n682 commonsourceibias.n630 0.189894
R23122 commonsourceibias.n688 commonsourceibias.n630 0.189894
R23123 commonsourceibias.n689 commonsourceibias.n688 0.189894
R23124 commonsourceibias.n690 commonsourceibias.n689 0.189894
R23125 commonsourceibias.n690 commonsourceibias.n628 0.189894
R23126 commonsourceibias.n695 commonsourceibias.n628 0.189894
R23127 commonsourceibias.n696 commonsourceibias.n695 0.189894
R23128 commonsourceibias.n697 commonsourceibias.n696 0.189894
R23129 commonsourceibias.n697 commonsourceibias.n626 0.189894
R23130 commonsourceibias.n703 commonsourceibias.n626 0.189894
R23131 commonsourceibias.n704 commonsourceibias.n703 0.189894
R23132 commonsourceibias.n705 commonsourceibias.n704 0.189894
R23133 commonsourceibias.n705 commonsourceibias.n624 0.189894
R23134 commonsourceibias.n710 commonsourceibias.n624 0.189894
R23135 commonsourceibias.n711 commonsourceibias.n710 0.189894
R23136 commonsourceibias.n712 commonsourceibias.n711 0.189894
R23137 commonsourceibias.n712 commonsourceibias.n622 0.189894
R23138 commonsourceibias.n718 commonsourceibias.n622 0.189894
R23139 commonsourceibias.n719 commonsourceibias.n718 0.189894
R23140 commonsourceibias.n720 commonsourceibias.n719 0.189894
R23141 commonsourceibias.n720 commonsourceibias.n620 0.189894
R23142 commonsourceibias.n725 commonsourceibias.n620 0.189894
R23143 commonsourceibias.n726 commonsourceibias.n725 0.189894
R23144 commonsourceibias.n727 commonsourceibias.n726 0.189894
R23145 commonsourceibias.n727 commonsourceibias.n618 0.189894
R23146 commonsourceibias.n415 commonsourceibias.n414 0.189894
R23147 commonsourceibias.n415 commonsourceibias.n410 0.189894
R23148 commonsourceibias.n420 commonsourceibias.n410 0.189894
R23149 commonsourceibias.n421 commonsourceibias.n420 0.189894
R23150 commonsourceibias.n422 commonsourceibias.n421 0.189894
R23151 commonsourceibias.n422 commonsourceibias.n408 0.189894
R23152 commonsourceibias.n428 commonsourceibias.n408 0.189894
R23153 commonsourceibias.n429 commonsourceibias.n428 0.189894
R23154 commonsourceibias.n430 commonsourceibias.n429 0.189894
R23155 commonsourceibias.n430 commonsourceibias.n406 0.189894
R23156 commonsourceibias.n435 commonsourceibias.n406 0.189894
R23157 commonsourceibias.n436 commonsourceibias.n435 0.189894
R23158 commonsourceibias.n437 commonsourceibias.n436 0.189894
R23159 commonsourceibias.n437 commonsourceibias.n404 0.189894
R23160 commonsourceibias.n443 commonsourceibias.n404 0.189894
R23161 commonsourceibias.n444 commonsourceibias.n443 0.189894
R23162 commonsourceibias.n445 commonsourceibias.n444 0.189894
R23163 commonsourceibias.n445 commonsourceibias.n402 0.189894
R23164 commonsourceibias.n450 commonsourceibias.n402 0.189894
R23165 commonsourceibias.n451 commonsourceibias.n450 0.189894
R23166 commonsourceibias.n452 commonsourceibias.n451 0.189894
R23167 commonsourceibias.n452 commonsourceibias.n400 0.189894
R23168 commonsourceibias.n458 commonsourceibias.n400 0.189894
R23169 commonsourceibias.n459 commonsourceibias.n458 0.189894
R23170 commonsourceibias.n460 commonsourceibias.n459 0.189894
R23171 commonsourceibias.n460 commonsourceibias.n398 0.189894
R23172 commonsourceibias.n465 commonsourceibias.n398 0.189894
R23173 commonsourceibias.n466 commonsourceibias.n465 0.189894
R23174 commonsourceibias.n467 commonsourceibias.n466 0.189894
R23175 commonsourceibias.n467 commonsourceibias.n396 0.189894
R23176 commonsourceibias.n473 commonsourceibias.n396 0.189894
R23177 commonsourceibias.n474 commonsourceibias.n473 0.189894
R23178 commonsourceibias.n475 commonsourceibias.n474 0.189894
R23179 commonsourceibias.n475 commonsourceibias.n394 0.189894
R23180 commonsourceibias.n480 commonsourceibias.n394 0.189894
R23181 commonsourceibias.n481 commonsourceibias.n480 0.189894
R23182 commonsourceibias.n482 commonsourceibias.n481 0.189894
R23183 commonsourceibias.n482 commonsourceibias.n392 0.189894
R23184 commonsourceibias.n488 commonsourceibias.n392 0.189894
R23185 commonsourceibias.n489 commonsourceibias.n488 0.189894
R23186 commonsourceibias.n490 commonsourceibias.n489 0.189894
R23187 commonsourceibias.n490 commonsourceibias.n390 0.189894
R23188 commonsourceibias.n495 commonsourceibias.n390 0.189894
R23189 commonsourceibias.n496 commonsourceibias.n495 0.189894
R23190 commonsourceibias.n497 commonsourceibias.n496 0.189894
R23191 commonsourceibias.n497 commonsourceibias.n388 0.189894
R23192 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23193 commonsourceibias.n531 commonsourceibias.n526 0.189894
R23194 commonsourceibias.n536 commonsourceibias.n526 0.189894
R23195 commonsourceibias.n537 commonsourceibias.n536 0.189894
R23196 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23197 commonsourceibias.n538 commonsourceibias.n524 0.189894
R23198 commonsourceibias.n544 commonsourceibias.n524 0.189894
R23199 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23200 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23201 commonsourceibias.n546 commonsourceibias.n522 0.189894
R23202 commonsourceibias.n551 commonsourceibias.n522 0.189894
R23203 commonsourceibias.n552 commonsourceibias.n551 0.189894
R23204 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23205 commonsourceibias.n553 commonsourceibias.n520 0.189894
R23206 commonsourceibias.n558 commonsourceibias.n520 0.189894
R23207 commonsourceibias.n559 commonsourceibias.n558 0.189894
R23208 commonsourceibias.n559 commonsourceibias.n518 0.189894
R23209 commonsourceibias.n563 commonsourceibias.n518 0.189894
R23210 commonsourceibias.n564 commonsourceibias.n563 0.189894
R23211 commonsourceibias.n564 commonsourceibias.n516 0.189894
R23212 commonsourceibias.n568 commonsourceibias.n516 0.189894
R23213 commonsourceibias.n569 commonsourceibias.n568 0.189894
R23214 commonsourceibias.n574 commonsourceibias.n573 0.189894
R23215 commonsourceibias.n575 commonsourceibias.n574 0.189894
R23216 commonsourceibias.n575 commonsourceibias.n377 0.189894
R23217 commonsourceibias.n580 commonsourceibias.n377 0.189894
R23218 commonsourceibias.n581 commonsourceibias.n580 0.189894
R23219 commonsourceibias.n582 commonsourceibias.n581 0.189894
R23220 commonsourceibias.n582 commonsourceibias.n375 0.189894
R23221 commonsourceibias.n588 commonsourceibias.n375 0.189894
R23222 commonsourceibias.n589 commonsourceibias.n588 0.189894
R23223 commonsourceibias.n590 commonsourceibias.n589 0.189894
R23224 commonsourceibias.n590 commonsourceibias.n373 0.189894
R23225 commonsourceibias.n595 commonsourceibias.n373 0.189894
R23226 commonsourceibias.n596 commonsourceibias.n595 0.189894
R23227 commonsourceibias.n597 commonsourceibias.n596 0.189894
R23228 commonsourceibias.n597 commonsourceibias.n371 0.189894
R23229 commonsourceibias.n603 commonsourceibias.n371 0.189894
R23230 commonsourceibias.n604 commonsourceibias.n603 0.189894
R23231 commonsourceibias.n605 commonsourceibias.n604 0.189894
R23232 commonsourceibias.n605 commonsourceibias.n369 0.189894
R23233 commonsourceibias.n610 commonsourceibias.n369 0.189894
R23234 commonsourceibias.n611 commonsourceibias.n610 0.189894
R23235 commonsourceibias.n612 commonsourceibias.n611 0.189894
R23236 commonsourceibias.n612 commonsourceibias.n367 0.189894
R23237 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R23238 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R23239 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R23240 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R23241 output.n41 output.n15 289.615
R23242 output.n72 output.n46 289.615
R23243 output.n104 output.n78 289.615
R23244 output.n136 output.n110 289.615
R23245 output.n77 output.n45 197.26
R23246 output.n77 output.n76 196.298
R23247 output.n109 output.n108 196.298
R23248 output.n141 output.n140 196.298
R23249 output.n42 output.n41 185
R23250 output.n40 output.n39 185
R23251 output.n19 output.n18 185
R23252 output.n34 output.n33 185
R23253 output.n32 output.n31 185
R23254 output.n23 output.n22 185
R23255 output.n26 output.n25 185
R23256 output.n73 output.n72 185
R23257 output.n71 output.n70 185
R23258 output.n50 output.n49 185
R23259 output.n65 output.n64 185
R23260 output.n63 output.n62 185
R23261 output.n54 output.n53 185
R23262 output.n57 output.n56 185
R23263 output.n105 output.n104 185
R23264 output.n103 output.n102 185
R23265 output.n82 output.n81 185
R23266 output.n97 output.n96 185
R23267 output.n95 output.n94 185
R23268 output.n86 output.n85 185
R23269 output.n89 output.n88 185
R23270 output.n137 output.n136 185
R23271 output.n135 output.n134 185
R23272 output.n114 output.n113 185
R23273 output.n129 output.n128 185
R23274 output.n127 output.n126 185
R23275 output.n118 output.n117 185
R23276 output.n121 output.n120 185
R23277 output.t3 output.n24 147.661
R23278 output.t1 output.n55 147.661
R23279 output.t2 output.n87 147.661
R23280 output.t0 output.n119 147.661
R23281 output.n41 output.n40 104.615
R23282 output.n40 output.n18 104.615
R23283 output.n33 output.n18 104.615
R23284 output.n33 output.n32 104.615
R23285 output.n32 output.n22 104.615
R23286 output.n25 output.n22 104.615
R23287 output.n72 output.n71 104.615
R23288 output.n71 output.n49 104.615
R23289 output.n64 output.n49 104.615
R23290 output.n64 output.n63 104.615
R23291 output.n63 output.n53 104.615
R23292 output.n56 output.n53 104.615
R23293 output.n104 output.n103 104.615
R23294 output.n103 output.n81 104.615
R23295 output.n96 output.n81 104.615
R23296 output.n96 output.n95 104.615
R23297 output.n95 output.n85 104.615
R23298 output.n88 output.n85 104.615
R23299 output.n136 output.n135 104.615
R23300 output.n135 output.n113 104.615
R23301 output.n128 output.n113 104.615
R23302 output.n128 output.n127 104.615
R23303 output.n127 output.n117 104.615
R23304 output.n120 output.n117 104.615
R23305 output.n1 output.t13 77.056
R23306 output.n14 output.t15 76.6694
R23307 output.n1 output.n0 72.7095
R23308 output.n3 output.n2 72.7095
R23309 output.n5 output.n4 72.7095
R23310 output.n7 output.n6 72.7095
R23311 output.n9 output.n8 72.7095
R23312 output.n11 output.n10 72.7095
R23313 output.n13 output.n12 72.7095
R23314 output.n25 output.t3 52.3082
R23315 output.n56 output.t1 52.3082
R23316 output.n88 output.t2 52.3082
R23317 output.n120 output.t0 52.3082
R23318 output.n26 output.n24 15.6674
R23319 output.n57 output.n55 15.6674
R23320 output.n89 output.n87 15.6674
R23321 output.n121 output.n119 15.6674
R23322 output.n27 output.n23 12.8005
R23323 output.n58 output.n54 12.8005
R23324 output.n90 output.n86 12.8005
R23325 output.n122 output.n118 12.8005
R23326 output.n31 output.n30 12.0247
R23327 output.n62 output.n61 12.0247
R23328 output.n94 output.n93 12.0247
R23329 output.n126 output.n125 12.0247
R23330 output.n34 output.n21 11.249
R23331 output.n65 output.n52 11.249
R23332 output.n97 output.n84 11.249
R23333 output.n129 output.n116 11.249
R23334 output.n35 output.n19 10.4732
R23335 output.n66 output.n50 10.4732
R23336 output.n98 output.n82 10.4732
R23337 output.n130 output.n114 10.4732
R23338 output.n39 output.n38 9.69747
R23339 output.n70 output.n69 9.69747
R23340 output.n102 output.n101 9.69747
R23341 output.n134 output.n133 9.69747
R23342 output.n45 output.n44 9.45567
R23343 output.n76 output.n75 9.45567
R23344 output.n108 output.n107 9.45567
R23345 output.n140 output.n139 9.45567
R23346 output.n44 output.n43 9.3005
R23347 output.n17 output.n16 9.3005
R23348 output.n38 output.n37 9.3005
R23349 output.n36 output.n35 9.3005
R23350 output.n21 output.n20 9.3005
R23351 output.n30 output.n29 9.3005
R23352 output.n28 output.n27 9.3005
R23353 output.n75 output.n74 9.3005
R23354 output.n48 output.n47 9.3005
R23355 output.n69 output.n68 9.3005
R23356 output.n67 output.n66 9.3005
R23357 output.n52 output.n51 9.3005
R23358 output.n61 output.n60 9.3005
R23359 output.n59 output.n58 9.3005
R23360 output.n107 output.n106 9.3005
R23361 output.n80 output.n79 9.3005
R23362 output.n101 output.n100 9.3005
R23363 output.n99 output.n98 9.3005
R23364 output.n84 output.n83 9.3005
R23365 output.n93 output.n92 9.3005
R23366 output.n91 output.n90 9.3005
R23367 output.n139 output.n138 9.3005
R23368 output.n112 output.n111 9.3005
R23369 output.n133 output.n132 9.3005
R23370 output.n131 output.n130 9.3005
R23371 output.n116 output.n115 9.3005
R23372 output.n125 output.n124 9.3005
R23373 output.n123 output.n122 9.3005
R23374 output.n42 output.n17 8.92171
R23375 output.n73 output.n48 8.92171
R23376 output.n105 output.n80 8.92171
R23377 output.n137 output.n112 8.92171
R23378 output output.n141 8.15037
R23379 output.n43 output.n15 8.14595
R23380 output.n74 output.n46 8.14595
R23381 output.n106 output.n78 8.14595
R23382 output.n138 output.n110 8.14595
R23383 output.n45 output.n15 5.81868
R23384 output.n76 output.n46 5.81868
R23385 output.n108 output.n78 5.81868
R23386 output.n140 output.n110 5.81868
R23387 output.n43 output.n42 5.04292
R23388 output.n74 output.n73 5.04292
R23389 output.n106 output.n105 5.04292
R23390 output.n138 output.n137 5.04292
R23391 output.n28 output.n24 4.38594
R23392 output.n59 output.n55 4.38594
R23393 output.n91 output.n87 4.38594
R23394 output.n123 output.n119 4.38594
R23395 output.n39 output.n17 4.26717
R23396 output.n70 output.n48 4.26717
R23397 output.n102 output.n80 4.26717
R23398 output.n134 output.n112 4.26717
R23399 output.n0 output.t19 3.9605
R23400 output.n0 output.t8 3.9605
R23401 output.n2 output.t12 3.9605
R23402 output.n2 output.t4 3.9605
R23403 output.n4 output.t6 3.9605
R23404 output.n4 output.t5 3.9605
R23405 output.n6 output.t11 3.9605
R23406 output.n6 output.t14 3.9605
R23407 output.n8 output.t16 3.9605
R23408 output.n8 output.t9 3.9605
R23409 output.n10 output.t10 3.9605
R23410 output.n10 output.t17 3.9605
R23411 output.n12 output.t18 3.9605
R23412 output.n12 output.t7 3.9605
R23413 output.n38 output.n19 3.49141
R23414 output.n69 output.n50 3.49141
R23415 output.n101 output.n82 3.49141
R23416 output.n133 output.n114 3.49141
R23417 output.n35 output.n34 2.71565
R23418 output.n66 output.n65 2.71565
R23419 output.n98 output.n97 2.71565
R23420 output.n130 output.n129 2.71565
R23421 output.n31 output.n21 1.93989
R23422 output.n62 output.n52 1.93989
R23423 output.n94 output.n84 1.93989
R23424 output.n126 output.n116 1.93989
R23425 output.n30 output.n23 1.16414
R23426 output.n61 output.n54 1.16414
R23427 output.n93 output.n86 1.16414
R23428 output.n125 output.n118 1.16414
R23429 output.n141 output.n109 0.962709
R23430 output.n109 output.n77 0.962709
R23431 output.n27 output.n26 0.388379
R23432 output.n58 output.n57 0.388379
R23433 output.n90 output.n89 0.388379
R23434 output.n122 output.n121 0.388379
R23435 output.n14 output.n13 0.387128
R23436 output.n13 output.n11 0.387128
R23437 output.n11 output.n9 0.387128
R23438 output.n9 output.n7 0.387128
R23439 output.n7 output.n5 0.387128
R23440 output.n5 output.n3 0.387128
R23441 output.n3 output.n1 0.387128
R23442 output.n44 output.n16 0.155672
R23443 output.n37 output.n16 0.155672
R23444 output.n37 output.n36 0.155672
R23445 output.n36 output.n20 0.155672
R23446 output.n29 output.n20 0.155672
R23447 output.n29 output.n28 0.155672
R23448 output.n75 output.n47 0.155672
R23449 output.n68 output.n47 0.155672
R23450 output.n68 output.n67 0.155672
R23451 output.n67 output.n51 0.155672
R23452 output.n60 output.n51 0.155672
R23453 output.n60 output.n59 0.155672
R23454 output.n107 output.n79 0.155672
R23455 output.n100 output.n79 0.155672
R23456 output.n100 output.n99 0.155672
R23457 output.n99 output.n83 0.155672
R23458 output.n92 output.n83 0.155672
R23459 output.n92 output.n91 0.155672
R23460 output.n139 output.n111 0.155672
R23461 output.n132 output.n111 0.155672
R23462 output.n132 output.n131 0.155672
R23463 output.n131 output.n115 0.155672
R23464 output.n124 output.n115 0.155672
R23465 output.n124 output.n123 0.155672
R23466 output output.n14 0.126227
R23467 a_n2318_8322.n8 a_n2318_8322.t3 74.6477
R23468 a_n2318_8322.n1 a_n2318_8322.t22 74.6477
R23469 a_n2318_8322.n20 a_n2318_8322.t21 74.6474
R23470 a_n2318_8322.n16 a_n2318_8322.t11 74.2899
R23471 a_n2318_8322.n9 a_n2318_8322.t1 74.2899
R23472 a_n2318_8322.n10 a_n2318_8322.t4 74.2899
R23473 a_n2318_8322.n13 a_n2318_8322.t5 74.2899
R23474 a_n2318_8322.n6 a_n2318_8322.t8 74.2899
R23475 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23476 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23477 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R23478 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R23479 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23480 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23481 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23482 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R23483 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R23484 a_n2318_8322.n15 a_n2318_8322.t24 10.1716
R23485 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R23486 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R23487 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R23488 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R23489 a_n2318_8322.n19 a_n2318_8322.t15 3.61217
R23490 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R23491 a_n2318_8322.n17 a_n2318_8322.t13 3.61217
R23492 a_n2318_8322.n7 a_n2318_8322.t7 3.61217
R23493 a_n2318_8322.n7 a_n2318_8322.t6 3.61217
R23494 a_n2318_8322.n11 a_n2318_8322.t2 3.61217
R23495 a_n2318_8322.n11 a_n2318_8322.t0 3.61217
R23496 a_n2318_8322.n0 a_n2318_8322.t10 3.61217
R23497 a_n2318_8322.n0 a_n2318_8322.t9 3.61217
R23498 a_n2318_8322.n2 a_n2318_8322.t19 3.61217
R23499 a_n2318_8322.n2 a_n2318_8322.t14 3.61217
R23500 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R23501 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R23502 a_n2318_8322.n22 a_n2318_8322.t12 3.61217
R23503 a_n2318_8322.t23 a_n2318_8322.n22 3.61217
R23504 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R23505 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R23506 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R23507 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23508 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23509 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23510 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23511 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R23512 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R23513 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R23514 a_n2318_8322.t27 a_n2318_8322.t26 0.0788333
R23515 a_n2318_8322.t25 a_n2318_8322.t27 0.0631667
R23516 a_n2318_8322.t24 a_n2318_8322.t25 0.0471944
R23517 a_n2318_8322.t24 a_n2318_8322.t26 0.0453889
R23518 plus.n34 plus.t22 436.949
R23519 plus.n8 plus.t12 436.949
R23520 plus.n35 plus.t5 415.966
R23521 plus.n33 plus.t19 415.966
R23522 plus.n41 plus.t23 415.966
R23523 plus.n42 plus.t11 415.966
R23524 plus.n46 plus.t6 415.966
R23525 plus.n47 plus.t10 415.966
R23526 plus.n29 plus.t18 415.966
R23527 plus.n53 plus.t8 415.966
R23528 plus.n54 plus.t15 415.966
R23529 plus.n26 plus.t24 415.966
R23530 plus.n25 plus.t20 415.966
R23531 plus.n1 plus.t7 415.966
R23532 plus.n19 plus.t17 415.966
R23533 plus.n18 plus.t13 415.966
R23534 plus.n4 plus.t21 415.966
R23535 plus.n13 plus.t16 415.966
R23536 plus.n11 plus.t9 415.966
R23537 plus.n7 plus.t14 415.966
R23538 plus.n58 plus.t0 243.97
R23539 plus.n58 plus.n57 223.454
R23540 plus.n60 plus.n59 223.454
R23541 plus.n55 plus.n54 161.3
R23542 plus.n53 plus.n28 161.3
R23543 plus.n52 plus.n51 161.3
R23544 plus.n50 plus.n29 161.3
R23545 plus.n49 plus.n48 161.3
R23546 plus.n47 plus.n30 161.3
R23547 plus.n46 plus.n45 161.3
R23548 plus.n44 plus.n31 161.3
R23549 plus.n43 plus.n42 161.3
R23550 plus.n41 plus.n32 161.3
R23551 plus.n40 plus.n39 161.3
R23552 plus.n38 plus.n33 161.3
R23553 plus.n37 plus.n36 161.3
R23554 plus.n10 plus.n9 161.3
R23555 plus.n11 plus.n6 161.3
R23556 plus.n12 plus.n5 161.3
R23557 plus.n14 plus.n13 161.3
R23558 plus.n15 plus.n4 161.3
R23559 plus.n17 plus.n16 161.3
R23560 plus.n18 plus.n3 161.3
R23561 plus.n19 plus.n2 161.3
R23562 plus.n21 plus.n20 161.3
R23563 plus.n22 plus.n1 161.3
R23564 plus.n24 plus.n23 161.3
R23565 plus.n25 plus.n0 161.3
R23566 plus.n27 plus.n26 161.3
R23567 plus.n37 plus.n34 70.4033
R23568 plus.n9 plus.n8 70.4033
R23569 plus.n42 plus.n41 48.2005
R23570 plus.n47 plus.n46 48.2005
R23571 plus.n54 plus.n53 48.2005
R23572 plus.n26 plus.n25 48.2005
R23573 plus.n19 plus.n18 48.2005
R23574 plus.n13 plus.n4 48.2005
R23575 plus.n40 plus.n33 47.4702
R23576 plus.n48 plus.n29 47.4702
R23577 plus.n20 plus.n1 47.4702
R23578 plus.n12 plus.n11 47.4702
R23579 plus.n56 plus.n55 29.8622
R23580 plus.n36 plus.n33 25.5611
R23581 plus.n52 plus.n29 25.5611
R23582 plus.n24 plus.n1 25.5611
R23583 plus.n11 plus.n10 25.5611
R23584 plus.n42 plus.n31 24.1005
R23585 plus.n46 plus.n31 24.1005
R23586 plus.n18 plus.n17 24.1005
R23587 plus.n17 plus.n4 24.1005
R23588 plus.n36 plus.n35 22.6399
R23589 plus.n53 plus.n52 22.6399
R23590 plus.n25 plus.n24 22.6399
R23591 plus.n10 plus.n7 22.6399
R23592 plus.n35 plus.n34 20.9576
R23593 plus.n8 plus.n7 20.9576
R23594 plus.n57 plus.t3 19.8005
R23595 plus.n57 plus.t2 19.8005
R23596 plus.n59 plus.t4 19.8005
R23597 plus.n59 plus.t1 19.8005
R23598 plus plus.n61 14.929
R23599 plus.n56 plus.n27 11.7903
R23600 plus.n61 plus.n60 5.40567
R23601 plus.n61 plus.n56 1.188
R23602 plus.n41 plus.n40 0.730803
R23603 plus.n48 plus.n47 0.730803
R23604 plus.n20 plus.n19 0.730803
R23605 plus.n13 plus.n12 0.730803
R23606 plus.n60 plus.n58 0.716017
R23607 plus.n38 plus.n37 0.189894
R23608 plus.n39 plus.n38 0.189894
R23609 plus.n39 plus.n32 0.189894
R23610 plus.n43 plus.n32 0.189894
R23611 plus.n44 plus.n43 0.189894
R23612 plus.n45 plus.n44 0.189894
R23613 plus.n45 plus.n30 0.189894
R23614 plus.n49 plus.n30 0.189894
R23615 plus.n50 plus.n49 0.189894
R23616 plus.n51 plus.n50 0.189894
R23617 plus.n51 plus.n28 0.189894
R23618 plus.n55 plus.n28 0.189894
R23619 plus.n27 plus.n0 0.189894
R23620 plus.n23 plus.n0 0.189894
R23621 plus.n23 plus.n22 0.189894
R23622 plus.n22 plus.n21 0.189894
R23623 plus.n21 plus.n2 0.189894
R23624 plus.n3 plus.n2 0.189894
R23625 plus.n16 plus.n3 0.189894
R23626 plus.n16 plus.n15 0.189894
R23627 plus.n15 plus.n14 0.189894
R23628 plus.n14 plus.n5 0.189894
R23629 plus.n6 plus.n5 0.189894
R23630 plus.n9 plus.n6 0.189894
R23631 minus.n36 minus.t23 436.949
R23632 minus.n6 minus.t11 436.949
R23633 minus.n54 minus.t18 415.966
R23634 minus.n53 minus.t13 415.966
R23635 minus.n29 minus.t20 415.966
R23636 minus.n47 minus.t10 415.966
R23637 minus.n46 minus.t5 415.966
R23638 minus.n32 minus.t14 415.966
R23639 minus.n41 minus.t9 415.966
R23640 minus.n39 minus.t22 415.966
R23641 minus.n35 minus.t7 415.966
R23642 minus.n7 minus.t15 415.966
R23643 minus.n5 minus.t8 415.966
R23644 minus.n13 minus.t12 415.966
R23645 minus.n14 minus.t21 415.966
R23646 minus.n18 minus.t16 415.966
R23647 minus.n19 minus.t19 415.966
R23648 minus.n1 minus.t6 415.966
R23649 minus.n25 minus.t17 415.966
R23650 minus.n26 minus.t24 415.966
R23651 minus.n60 minus.t1 243.255
R23652 minus.n59 minus.n57 224.169
R23653 minus.n59 minus.n58 223.454
R23654 minus.n38 minus.n37 161.3
R23655 minus.n39 minus.n34 161.3
R23656 minus.n40 minus.n33 161.3
R23657 minus.n42 minus.n41 161.3
R23658 minus.n43 minus.n32 161.3
R23659 minus.n45 minus.n44 161.3
R23660 minus.n46 minus.n31 161.3
R23661 minus.n47 minus.n30 161.3
R23662 minus.n49 minus.n48 161.3
R23663 minus.n50 minus.n29 161.3
R23664 minus.n52 minus.n51 161.3
R23665 minus.n53 minus.n28 161.3
R23666 minus.n55 minus.n54 161.3
R23667 minus.n27 minus.n26 161.3
R23668 minus.n25 minus.n0 161.3
R23669 minus.n24 minus.n23 161.3
R23670 minus.n22 minus.n1 161.3
R23671 minus.n21 minus.n20 161.3
R23672 minus.n19 minus.n2 161.3
R23673 minus.n18 minus.n17 161.3
R23674 minus.n16 minus.n3 161.3
R23675 minus.n15 minus.n14 161.3
R23676 minus.n13 minus.n4 161.3
R23677 minus.n12 minus.n11 161.3
R23678 minus.n10 minus.n5 161.3
R23679 minus.n9 minus.n8 161.3
R23680 minus.n37 minus.n36 70.4033
R23681 minus.n9 minus.n6 70.4033
R23682 minus.n54 minus.n53 48.2005
R23683 minus.n47 minus.n46 48.2005
R23684 minus.n41 minus.n32 48.2005
R23685 minus.n14 minus.n13 48.2005
R23686 minus.n19 minus.n18 48.2005
R23687 minus.n26 minus.n25 48.2005
R23688 minus.n48 minus.n29 47.4702
R23689 minus.n40 minus.n39 47.4702
R23690 minus.n12 minus.n5 47.4702
R23691 minus.n20 minus.n1 47.4702
R23692 minus.n56 minus.n55 30.0782
R23693 minus.n52 minus.n29 25.5611
R23694 minus.n39 minus.n38 25.5611
R23695 minus.n8 minus.n5 25.5611
R23696 minus.n24 minus.n1 25.5611
R23697 minus.n46 minus.n45 24.1005
R23698 minus.n45 minus.n32 24.1005
R23699 minus.n14 minus.n3 24.1005
R23700 minus.n18 minus.n3 24.1005
R23701 minus.n53 minus.n52 22.6399
R23702 minus.n38 minus.n35 22.6399
R23703 minus.n8 minus.n7 22.6399
R23704 minus.n25 minus.n24 22.6399
R23705 minus.n36 minus.n35 20.9576
R23706 minus.n7 minus.n6 20.9576
R23707 minus.n58 minus.t0 19.8005
R23708 minus.n58 minus.t4 19.8005
R23709 minus.n57 minus.t2 19.8005
R23710 minus.n57 minus.t3 19.8005
R23711 minus minus.n61 12.2993
R23712 minus.n56 minus.n27 12.0062
R23713 minus.n61 minus.n60 4.80222
R23714 minus.n61 minus.n56 0.972091
R23715 minus.n48 minus.n47 0.730803
R23716 minus.n41 minus.n40 0.730803
R23717 minus.n13 minus.n12 0.730803
R23718 minus.n20 minus.n19 0.730803
R23719 minus.n60 minus.n59 0.716017
R23720 minus.n55 minus.n28 0.189894
R23721 minus.n51 minus.n28 0.189894
R23722 minus.n51 minus.n50 0.189894
R23723 minus.n50 minus.n49 0.189894
R23724 minus.n49 minus.n30 0.189894
R23725 minus.n31 minus.n30 0.189894
R23726 minus.n44 minus.n31 0.189894
R23727 minus.n44 minus.n43 0.189894
R23728 minus.n43 minus.n42 0.189894
R23729 minus.n42 minus.n33 0.189894
R23730 minus.n34 minus.n33 0.189894
R23731 minus.n37 minus.n34 0.189894
R23732 minus.n10 minus.n9 0.189894
R23733 minus.n11 minus.n10 0.189894
R23734 minus.n11 minus.n4 0.189894
R23735 minus.n15 minus.n4 0.189894
R23736 minus.n16 minus.n15 0.189894
R23737 minus.n17 minus.n16 0.189894
R23738 minus.n17 minus.n2 0.189894
R23739 minus.n21 minus.n2 0.189894
R23740 minus.n22 minus.n21 0.189894
R23741 minus.n23 minus.n22 0.189894
R23742 minus.n23 minus.n0 0.189894
R23743 minus.n27 minus.n0 0.189894
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.116614p
C5 minus diffpairibias 2.77e-19
C6 commonsourceibias output 0.006808f
C7 vdd plus 0.082936f
C8 CSoutput minus 3.3847f
C9 plus diffpairibias 2.54e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.87913f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 45.462303f
C15 minus plus 9.54777f
C16 minus commonsourceibias 0.327318f
C17 plus commonsourceibias 0.272687f
C18 diffpairibias gnd 59.991035f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.182016p
C22 plus gnd 32.634003f
C23 minus gnd 28.6196f
C24 CSoutput gnd 0.115659p
C25 vdd gnd 0.443442p
C26 minus.n0 gnd 0.030606f
C27 minus.t6 gnd 0.309209f
C28 minus.n1 gnd 0.142957f
C29 minus.n2 gnd 0.030606f
C30 minus.n3 gnd 0.006945f
C31 minus.n4 gnd 0.030606f
C32 minus.t8 gnd 0.309209f
C33 minus.n5 gnd 0.142957f
C34 minus.t11 gnd 0.315922f
C35 minus.n6 gnd 0.133271f
C36 minus.t15 gnd 0.309209f
C37 minus.n7 gnd 0.142674f
C38 minus.n8 gnd 0.006945f
C39 minus.n9 gnd 0.100452f
C40 minus.n10 gnd 0.030606f
C41 minus.n11 gnd 0.030606f
C42 minus.n12 gnd 0.006945f
C43 minus.t12 gnd 0.309209f
C44 minus.n13 gnd 0.139844f
C45 minus.t21 gnd 0.309209f
C46 minus.n14 gnd 0.142863f
C47 minus.n15 gnd 0.030606f
C48 minus.n16 gnd 0.030606f
C49 minus.n17 gnd 0.030606f
C50 minus.t16 gnd 0.309209f
C51 minus.n18 gnd 0.142863f
C52 minus.t19 gnd 0.309209f
C53 minus.n19 gnd 0.139844f
C54 minus.n20 gnd 0.006945f
C55 minus.n21 gnd 0.030606f
C56 minus.n22 gnd 0.030606f
C57 minus.n23 gnd 0.030606f
C58 minus.n24 gnd 0.006945f
C59 minus.t17 gnd 0.309209f
C60 minus.n25 gnd 0.142674f
C61 minus.t24 gnd 0.309209f
C62 minus.n26 gnd 0.139749f
C63 minus.n27 gnd 0.348154f
C64 minus.n28 gnd 0.030606f
C65 minus.t18 gnd 0.309209f
C66 minus.t13 gnd 0.309209f
C67 minus.t20 gnd 0.309209f
C68 minus.n29 gnd 0.142957f
C69 minus.n30 gnd 0.030606f
C70 minus.t10 gnd 0.309209f
C71 minus.t5 gnd 0.309209f
C72 minus.n31 gnd 0.030606f
C73 minus.t14 gnd 0.309209f
C74 minus.n32 gnd 0.142863f
C75 minus.n33 gnd 0.030606f
C76 minus.t9 gnd 0.309209f
C77 minus.t22 gnd 0.309209f
C78 minus.n34 gnd 0.030606f
C79 minus.t7 gnd 0.309209f
C80 minus.n35 gnd 0.142674f
C81 minus.t23 gnd 0.315922f
C82 minus.n36 gnd 0.133271f
C83 minus.n37 gnd 0.100452f
C84 minus.n38 gnd 0.006945f
C85 minus.n39 gnd 0.142957f
C86 minus.n40 gnd 0.006945f
C87 minus.n41 gnd 0.139844f
C88 minus.n42 gnd 0.030606f
C89 minus.n43 gnd 0.030606f
C90 minus.n44 gnd 0.030606f
C91 minus.n45 gnd 0.006945f
C92 minus.n46 gnd 0.142863f
C93 minus.n47 gnd 0.139844f
C94 minus.n48 gnd 0.006945f
C95 minus.n49 gnd 0.030606f
C96 minus.n50 gnd 0.030606f
C97 minus.n51 gnd 0.030606f
C98 minus.n52 gnd 0.006945f
C99 minus.n53 gnd 0.142674f
C100 minus.n54 gnd 0.139749f
C101 minus.n55 gnd 0.879238f
C102 minus.n56 gnd 1.34121f
C103 minus.t2 gnd 0.009435f
C104 minus.t3 gnd 0.009435f
C105 minus.n57 gnd 0.031024f
C106 minus.t0 gnd 0.009435f
C107 minus.t4 gnd 0.009435f
C108 minus.n58 gnd 0.030599f
C109 minus.n59 gnd 0.26115f
C110 minus.t1 gnd 0.052514f
C111 minus.n60 gnd 0.142507f
C112 minus.n61 gnd 2.47488f
C113 plus.n0 gnd 0.022157f
C114 plus.t24 gnd 0.22385f
C115 plus.t20 gnd 0.22385f
C116 plus.t7 gnd 0.22385f
C117 plus.n1 gnd 0.103493f
C118 plus.n2 gnd 0.022157f
C119 plus.t17 gnd 0.22385f
C120 plus.n3 gnd 0.022157f
C121 plus.t13 gnd 0.22385f
C122 plus.t21 gnd 0.22385f
C123 plus.n4 gnd 0.103425f
C124 plus.n5 gnd 0.022157f
C125 plus.t16 gnd 0.22385f
C126 plus.n6 gnd 0.022157f
C127 plus.t9 gnd 0.22385f
C128 plus.t14 gnd 0.22385f
C129 plus.n7 gnd 0.103288f
C130 plus.t12 gnd 0.22871f
C131 plus.n8 gnd 0.096481f
C132 plus.n9 gnd 0.072722f
C133 plus.n10 gnd 0.005028f
C134 plus.n11 gnd 0.103493f
C135 plus.n12 gnd 0.005028f
C136 plus.n13 gnd 0.101239f
C137 plus.n14 gnd 0.022157f
C138 plus.n15 gnd 0.022157f
C139 plus.n16 gnd 0.022157f
C140 plus.n17 gnd 0.005028f
C141 plus.n18 gnd 0.103425f
C142 plus.n19 gnd 0.101239f
C143 plus.n20 gnd 0.005028f
C144 plus.n21 gnd 0.022157f
C145 plus.n22 gnd 0.022157f
C146 plus.n23 gnd 0.022157f
C147 plus.n24 gnd 0.005028f
C148 plus.n25 gnd 0.103288f
C149 plus.n26 gnd 0.101171f
C150 plus.n27 gnd 0.246327f
C151 plus.n28 gnd 0.022157f
C152 plus.t18 gnd 0.22385f
C153 plus.n29 gnd 0.103493f
C154 plus.n30 gnd 0.022157f
C155 plus.n31 gnd 0.005028f
C156 plus.t6 gnd 0.22385f
C157 plus.n32 gnd 0.022157f
C158 plus.t19 gnd 0.22385f
C159 plus.n33 gnd 0.103493f
C160 plus.t22 gnd 0.22871f
C161 plus.n34 gnd 0.096481f
C162 plus.t5 gnd 0.22385f
C163 plus.n35 gnd 0.103288f
C164 plus.n36 gnd 0.005028f
C165 plus.n37 gnd 0.072722f
C166 plus.n38 gnd 0.022157f
C167 plus.n39 gnd 0.022157f
C168 plus.n40 gnd 0.005028f
C169 plus.t23 gnd 0.22385f
C170 plus.n41 gnd 0.101239f
C171 plus.t11 gnd 0.22385f
C172 plus.n42 gnd 0.103425f
C173 plus.n43 gnd 0.022157f
C174 plus.n44 gnd 0.022157f
C175 plus.n45 gnd 0.022157f
C176 plus.n46 gnd 0.103425f
C177 plus.t10 gnd 0.22385f
C178 plus.n47 gnd 0.101239f
C179 plus.n48 gnd 0.005028f
C180 plus.n49 gnd 0.022157f
C181 plus.n50 gnd 0.022157f
C182 plus.n51 gnd 0.022157f
C183 plus.n52 gnd 0.005028f
C184 plus.t8 gnd 0.22385f
C185 plus.n53 gnd 0.103288f
C186 plus.t15 gnd 0.22385f
C187 plus.n54 gnd 0.101171f
C188 plus.n55 gnd 0.627617f
C189 plus.n56 gnd 0.962217f
C190 plus.t0 gnd 0.038249f
C191 plus.t3 gnd 0.00683f
C192 plus.t2 gnd 0.00683f
C193 plus.n57 gnd 0.022152f
C194 plus.n58 gnd 0.171968f
C195 plus.t4 gnd 0.00683f
C196 plus.t1 gnd 0.00683f
C197 plus.n59 gnd 0.022152f
C198 plus.n60 gnd 0.129083f
C199 plus.n61 gnd 2.84006f
C200 a_n2318_8322.t26 gnd 39.5788f
C201 a_n2318_8322.t24 gnd 29.8018f
C202 a_n2318_8322.t27 gnd 19.7198f
C203 a_n2318_8322.t25 gnd 39.5788f
C204 a_n2318_8322.t12 gnd 0.095725f
C205 a_n2318_8322.t22 gnd 0.89632f
C206 a_n2318_8322.t10 gnd 0.095725f
C207 a_n2318_8322.t9 gnd 0.095725f
C208 a_n2318_8322.n0 gnd 0.674286f
C209 a_n2318_8322.n1 gnd 0.753416f
C210 a_n2318_8322.t19 gnd 0.095725f
C211 a_n2318_8322.t14 gnd 0.095725f
C212 a_n2318_8322.n2 gnd 0.674286f
C213 a_n2318_8322.n3 gnd 0.382801f
C214 a_n2318_8322.t17 gnd 0.095725f
C215 a_n2318_8322.t16 gnd 0.095725f
C216 a_n2318_8322.n4 gnd 0.674286f
C217 a_n2318_8322.n5 gnd 0.382801f
C218 a_n2318_8322.t8 gnd 0.894535f
C219 a_n2318_8322.n6 gnd 1.55036f
C220 a_n2318_8322.t3 gnd 0.89632f
C221 a_n2318_8322.t7 gnd 0.095725f
C222 a_n2318_8322.t6 gnd 0.095725f
C223 a_n2318_8322.n7 gnd 0.674286f
C224 a_n2318_8322.n8 gnd 0.753416f
C225 a_n2318_8322.t1 gnd 0.894535f
C226 a_n2318_8322.n9 gnd 0.379129f
C227 a_n2318_8322.t4 gnd 0.894535f
C228 a_n2318_8322.n10 gnd 0.379129f
C229 a_n2318_8322.t2 gnd 0.095725f
C230 a_n2318_8322.t0 gnd 0.095725f
C231 a_n2318_8322.n11 gnd 0.674286f
C232 a_n2318_8322.n12 gnd 0.382801f
C233 a_n2318_8322.t5 gnd 0.894535f
C234 a_n2318_8322.n13 gnd 1.07361f
C235 a_n2318_8322.n14 gnd 1.82505f
C236 a_n2318_8322.n15 gnd 3.97113f
C237 a_n2318_8322.t11 gnd 0.894535f
C238 a_n2318_8322.n16 gnd 0.880601f
C239 a_n2318_8322.t20 gnd 0.095725f
C240 a_n2318_8322.t13 gnd 0.095725f
C241 a_n2318_8322.n17 gnd 0.674286f
C242 a_n2318_8322.n18 gnd 0.382801f
C243 a_n2318_8322.t21 gnd 0.896317f
C244 a_n2318_8322.t18 gnd 0.095725f
C245 a_n2318_8322.t15 gnd 0.095725f
C246 a_n2318_8322.n19 gnd 0.674286f
C247 a_n2318_8322.n20 gnd 0.753418f
C248 a_n2318_8322.n21 gnd 0.382799f
C249 a_n2318_8322.n22 gnd 0.674288f
C250 a_n2318_8322.t23 gnd 0.095725f
C251 output.t13 gnd 0.464308f
C252 output.t19 gnd 0.044422f
C253 output.t8 gnd 0.044422f
C254 output.n0 gnd 0.364624f
C255 output.n1 gnd 0.614102f
C256 output.t12 gnd 0.044422f
C257 output.t4 gnd 0.044422f
C258 output.n2 gnd 0.364624f
C259 output.n3 gnd 0.350265f
C260 output.t6 gnd 0.044422f
C261 output.t5 gnd 0.044422f
C262 output.n4 gnd 0.364624f
C263 output.n5 gnd 0.350265f
C264 output.t11 gnd 0.044422f
C265 output.t14 gnd 0.044422f
C266 output.n6 gnd 0.364624f
C267 output.n7 gnd 0.350265f
C268 output.t16 gnd 0.044422f
C269 output.t9 gnd 0.044422f
C270 output.n8 gnd 0.364624f
C271 output.n9 gnd 0.350265f
C272 output.t10 gnd 0.044422f
C273 output.t17 gnd 0.044422f
C274 output.n10 gnd 0.364624f
C275 output.n11 gnd 0.350265f
C276 output.t18 gnd 0.044422f
C277 output.t7 gnd 0.044422f
C278 output.n12 gnd 0.364624f
C279 output.n13 gnd 0.350265f
C280 output.t15 gnd 0.462979f
C281 output.n14 gnd 0.28994f
C282 output.n15 gnd 0.015803f
C283 output.n16 gnd 0.011243f
C284 output.n17 gnd 0.006041f
C285 output.n18 gnd 0.01428f
C286 output.n19 gnd 0.006397f
C287 output.n20 gnd 0.011243f
C288 output.n21 gnd 0.006041f
C289 output.n22 gnd 0.01428f
C290 output.n23 gnd 0.006397f
C291 output.n24 gnd 0.048111f
C292 output.t3 gnd 0.023274f
C293 output.n25 gnd 0.01071f
C294 output.n26 gnd 0.008435f
C295 output.n27 gnd 0.006041f
C296 output.n28 gnd 0.267512f
C297 output.n29 gnd 0.011243f
C298 output.n30 gnd 0.006041f
C299 output.n31 gnd 0.006397f
C300 output.n32 gnd 0.01428f
C301 output.n33 gnd 0.01428f
C302 output.n34 gnd 0.006397f
C303 output.n35 gnd 0.006041f
C304 output.n36 gnd 0.011243f
C305 output.n37 gnd 0.011243f
C306 output.n38 gnd 0.006041f
C307 output.n39 gnd 0.006397f
C308 output.n40 gnd 0.01428f
C309 output.n41 gnd 0.030913f
C310 output.n42 gnd 0.006397f
C311 output.n43 gnd 0.006041f
C312 output.n44 gnd 0.025987f
C313 output.n45 gnd 0.097665f
C314 output.n46 gnd 0.015803f
C315 output.n47 gnd 0.011243f
C316 output.n48 gnd 0.006041f
C317 output.n49 gnd 0.01428f
C318 output.n50 gnd 0.006397f
C319 output.n51 gnd 0.011243f
C320 output.n52 gnd 0.006041f
C321 output.n53 gnd 0.01428f
C322 output.n54 gnd 0.006397f
C323 output.n55 gnd 0.048111f
C324 output.t1 gnd 0.023274f
C325 output.n56 gnd 0.01071f
C326 output.n57 gnd 0.008435f
C327 output.n58 gnd 0.006041f
C328 output.n59 gnd 0.267512f
C329 output.n60 gnd 0.011243f
C330 output.n61 gnd 0.006041f
C331 output.n62 gnd 0.006397f
C332 output.n63 gnd 0.01428f
C333 output.n64 gnd 0.01428f
C334 output.n65 gnd 0.006397f
C335 output.n66 gnd 0.006041f
C336 output.n67 gnd 0.011243f
C337 output.n68 gnd 0.011243f
C338 output.n69 gnd 0.006041f
C339 output.n70 gnd 0.006397f
C340 output.n71 gnd 0.01428f
C341 output.n72 gnd 0.030913f
C342 output.n73 gnd 0.006397f
C343 output.n74 gnd 0.006041f
C344 output.n75 gnd 0.025987f
C345 output.n76 gnd 0.09306f
C346 output.n77 gnd 1.65264f
C347 output.n78 gnd 0.015803f
C348 output.n79 gnd 0.011243f
C349 output.n80 gnd 0.006041f
C350 output.n81 gnd 0.01428f
C351 output.n82 gnd 0.006397f
C352 output.n83 gnd 0.011243f
C353 output.n84 gnd 0.006041f
C354 output.n85 gnd 0.01428f
C355 output.n86 gnd 0.006397f
C356 output.n87 gnd 0.048111f
C357 output.t2 gnd 0.023274f
C358 output.n88 gnd 0.01071f
C359 output.n89 gnd 0.008435f
C360 output.n90 gnd 0.006041f
C361 output.n91 gnd 0.267512f
C362 output.n92 gnd 0.011243f
C363 output.n93 gnd 0.006041f
C364 output.n94 gnd 0.006397f
C365 output.n95 gnd 0.01428f
C366 output.n96 gnd 0.01428f
C367 output.n97 gnd 0.006397f
C368 output.n98 gnd 0.006041f
C369 output.n99 gnd 0.011243f
C370 output.n100 gnd 0.011243f
C371 output.n101 gnd 0.006041f
C372 output.n102 gnd 0.006397f
C373 output.n103 gnd 0.01428f
C374 output.n104 gnd 0.030913f
C375 output.n105 gnd 0.006397f
C376 output.n106 gnd 0.006041f
C377 output.n107 gnd 0.025987f
C378 output.n108 gnd 0.09306f
C379 output.n109 gnd 0.713089f
C380 output.n110 gnd 0.015803f
C381 output.n111 gnd 0.011243f
C382 output.n112 gnd 0.006041f
C383 output.n113 gnd 0.01428f
C384 output.n114 gnd 0.006397f
C385 output.n115 gnd 0.011243f
C386 output.n116 gnd 0.006041f
C387 output.n117 gnd 0.01428f
C388 output.n118 gnd 0.006397f
C389 output.n119 gnd 0.048111f
C390 output.t0 gnd 0.023274f
C391 output.n120 gnd 0.01071f
C392 output.n121 gnd 0.008435f
C393 output.n122 gnd 0.006041f
C394 output.n123 gnd 0.267512f
C395 output.n124 gnd 0.011243f
C396 output.n125 gnd 0.006041f
C397 output.n126 gnd 0.006397f
C398 output.n127 gnd 0.01428f
C399 output.n128 gnd 0.01428f
C400 output.n129 gnd 0.006397f
C401 output.n130 gnd 0.006041f
C402 output.n131 gnd 0.011243f
C403 output.n132 gnd 0.011243f
C404 output.n133 gnd 0.006041f
C405 output.n134 gnd 0.006397f
C406 output.n135 gnd 0.01428f
C407 output.n136 gnd 0.030913f
C408 output.n137 gnd 0.006397f
C409 output.n138 gnd 0.006041f
C410 output.n139 gnd 0.025987f
C411 output.n140 gnd 0.09306f
C412 output.n141 gnd 1.67353f
C413 commonsourceibias.n0 gnd 0.010724f
C414 commonsourceibias.t115 gnd 0.162395f
C415 commonsourceibias.t136 gnd 0.150157f
C416 commonsourceibias.n1 gnd 0.007823f
C417 commonsourceibias.n2 gnd 0.008037f
C418 commonsourceibias.t151 gnd 0.150157f
C419 commonsourceibias.n3 gnd 0.01034f
C420 commonsourceibias.n4 gnd 0.008037f
C421 commonsourceibias.t105 gnd 0.150157f
C422 commonsourceibias.n5 gnd 0.059912f
C423 commonsourceibias.t126 gnd 0.150157f
C424 commonsourceibias.n6 gnd 0.007578f
C425 commonsourceibias.n7 gnd 0.008037f
C426 commonsourceibias.t144 gnd 0.150157f
C427 commonsourceibias.n8 gnd 0.010186f
C428 commonsourceibias.n9 gnd 0.008037f
C429 commonsourceibias.t98 gnd 0.150157f
C430 commonsourceibias.n10 gnd 0.059912f
C431 commonsourceibias.t94 gnd 0.150157f
C432 commonsourceibias.n11 gnd 0.007361f
C433 commonsourceibias.n12 gnd 0.008037f
C434 commonsourceibias.t135 gnd 0.150157f
C435 commonsourceibias.n13 gnd 0.010015f
C436 commonsourceibias.n14 gnd 0.010724f
C437 commonsourceibias.t74 gnd 0.162395f
C438 commonsourceibias.t20 gnd 0.150157f
C439 commonsourceibias.n15 gnd 0.007823f
C440 commonsourceibias.n16 gnd 0.008037f
C441 commonsourceibias.t50 gnd 0.150157f
C442 commonsourceibias.n17 gnd 0.01034f
C443 commonsourceibias.n18 gnd 0.008037f
C444 commonsourceibias.t8 gnd 0.150157f
C445 commonsourceibias.n19 gnd 0.059912f
C446 commonsourceibias.t36 gnd 0.150157f
C447 commonsourceibias.n20 gnd 0.007578f
C448 commonsourceibias.n21 gnd 0.008037f
C449 commonsourceibias.t76 gnd 0.150157f
C450 commonsourceibias.n22 gnd 0.010186f
C451 commonsourceibias.n23 gnd 0.008037f
C452 commonsourceibias.t24 gnd 0.150157f
C453 commonsourceibias.n24 gnd 0.059912f
C454 commonsourceibias.t34 gnd 0.150157f
C455 commonsourceibias.n25 gnd 0.007361f
C456 commonsourceibias.n26 gnd 0.008037f
C457 commonsourceibias.t10 gnd 0.150157f
C458 commonsourceibias.n27 gnd 0.010015f
C459 commonsourceibias.n28 gnd 0.008037f
C460 commonsourceibias.t40 gnd 0.150157f
C461 commonsourceibias.n29 gnd 0.059912f
C462 commonsourceibias.t56 gnd 0.150157f
C463 commonsourceibias.n30 gnd 0.007172f
C464 commonsourceibias.n31 gnd 0.008037f
C465 commonsourceibias.t26 gnd 0.150157f
C466 commonsourceibias.n32 gnd 0.009825f
C467 commonsourceibias.n33 gnd 0.008037f
C468 commonsourceibias.t38 gnd 0.150157f
C469 commonsourceibias.n34 gnd 0.059912f
C470 commonsourceibias.t70 gnd 0.150157f
C471 commonsourceibias.n35 gnd 0.007008f
C472 commonsourceibias.n36 gnd 0.008037f
C473 commonsourceibias.t18 gnd 0.150157f
C474 commonsourceibias.n37 gnd 0.009613f
C475 commonsourceibias.n38 gnd 0.008037f
C476 commonsourceibias.t22 gnd 0.150157f
C477 commonsourceibias.n39 gnd 0.059912f
C478 commonsourceibias.t54 gnd 0.150157f
C479 commonsourceibias.n40 gnd 0.006868f
C480 commonsourceibias.n41 gnd 0.008037f
C481 commonsourceibias.t4 gnd 0.150157f
C482 commonsourceibias.n42 gnd 0.009378f
C483 commonsourceibias.t78 gnd 0.166947f
C484 commonsourceibias.t46 gnd 0.150157f
C485 commonsourceibias.n43 gnd 0.065449f
C486 commonsourceibias.n44 gnd 0.071822f
C487 commonsourceibias.n45 gnd 0.033327f
C488 commonsourceibias.n46 gnd 0.008037f
C489 commonsourceibias.n47 gnd 0.007823f
C490 commonsourceibias.n48 gnd 0.01121f
C491 commonsourceibias.n49 gnd 0.059912f
C492 commonsourceibias.n50 gnd 0.011203f
C493 commonsourceibias.n51 gnd 0.008037f
C494 commonsourceibias.n52 gnd 0.008037f
C495 commonsourceibias.n53 gnd 0.008037f
C496 commonsourceibias.n54 gnd 0.01034f
C497 commonsourceibias.n55 gnd 0.059912f
C498 commonsourceibias.n56 gnd 0.010583f
C499 commonsourceibias.n57 gnd 0.010282f
C500 commonsourceibias.n58 gnd 0.008037f
C501 commonsourceibias.n59 gnd 0.008037f
C502 commonsourceibias.n60 gnd 0.008037f
C503 commonsourceibias.n61 gnd 0.007578f
C504 commonsourceibias.n62 gnd 0.01122f
C505 commonsourceibias.n63 gnd 0.059912f
C506 commonsourceibias.n64 gnd 0.011217f
C507 commonsourceibias.n65 gnd 0.008037f
C508 commonsourceibias.n66 gnd 0.008037f
C509 commonsourceibias.n67 gnd 0.008037f
C510 commonsourceibias.n68 gnd 0.010186f
C511 commonsourceibias.n69 gnd 0.059912f
C512 commonsourceibias.n70 gnd 0.010507f
C513 commonsourceibias.n71 gnd 0.010357f
C514 commonsourceibias.n72 gnd 0.008037f
C515 commonsourceibias.n73 gnd 0.008037f
C516 commonsourceibias.n74 gnd 0.008037f
C517 commonsourceibias.n75 gnd 0.007361f
C518 commonsourceibias.n76 gnd 0.011225f
C519 commonsourceibias.n77 gnd 0.059912f
C520 commonsourceibias.n78 gnd 0.011224f
C521 commonsourceibias.n79 gnd 0.008037f
C522 commonsourceibias.n80 gnd 0.008037f
C523 commonsourceibias.n81 gnd 0.008037f
C524 commonsourceibias.n82 gnd 0.010015f
C525 commonsourceibias.n83 gnd 0.059912f
C526 commonsourceibias.n84 gnd 0.010432f
C527 commonsourceibias.n85 gnd 0.010432f
C528 commonsourceibias.n86 gnd 0.008037f
C529 commonsourceibias.n87 gnd 0.008037f
C530 commonsourceibias.n88 gnd 0.008037f
C531 commonsourceibias.n89 gnd 0.007172f
C532 commonsourceibias.n90 gnd 0.011224f
C533 commonsourceibias.n91 gnd 0.059912f
C534 commonsourceibias.n92 gnd 0.011225f
C535 commonsourceibias.n93 gnd 0.008037f
C536 commonsourceibias.n94 gnd 0.008037f
C537 commonsourceibias.n95 gnd 0.008037f
C538 commonsourceibias.n96 gnd 0.009825f
C539 commonsourceibias.n97 gnd 0.059912f
C540 commonsourceibias.n98 gnd 0.010357f
C541 commonsourceibias.n99 gnd 0.010507f
C542 commonsourceibias.n100 gnd 0.008037f
C543 commonsourceibias.n101 gnd 0.008037f
C544 commonsourceibias.n102 gnd 0.008037f
C545 commonsourceibias.n103 gnd 0.007008f
C546 commonsourceibias.n104 gnd 0.011217f
C547 commonsourceibias.n105 gnd 0.059912f
C548 commonsourceibias.n106 gnd 0.01122f
C549 commonsourceibias.n107 gnd 0.008037f
C550 commonsourceibias.n108 gnd 0.008037f
C551 commonsourceibias.n109 gnd 0.008037f
C552 commonsourceibias.n110 gnd 0.009613f
C553 commonsourceibias.n111 gnd 0.059912f
C554 commonsourceibias.n112 gnd 0.010282f
C555 commonsourceibias.n113 gnd 0.010583f
C556 commonsourceibias.n114 gnd 0.008037f
C557 commonsourceibias.n115 gnd 0.008037f
C558 commonsourceibias.n116 gnd 0.008037f
C559 commonsourceibias.n117 gnd 0.006868f
C560 commonsourceibias.n118 gnd 0.011203f
C561 commonsourceibias.n119 gnd 0.059912f
C562 commonsourceibias.n120 gnd 0.01121f
C563 commonsourceibias.n121 gnd 0.008037f
C564 commonsourceibias.n122 gnd 0.008037f
C565 commonsourceibias.n123 gnd 0.008037f
C566 commonsourceibias.n124 gnd 0.009378f
C567 commonsourceibias.n125 gnd 0.059912f
C568 commonsourceibias.n126 gnd 0.009861f
C569 commonsourceibias.n127 gnd 0.07189f
C570 commonsourceibias.n128 gnd 0.080075f
C571 commonsourceibias.t75 gnd 0.017343f
C572 commonsourceibias.t21 gnd 0.017343f
C573 commonsourceibias.n129 gnd 0.15325f
C574 commonsourceibias.n130 gnd 0.132562f
C575 commonsourceibias.t51 gnd 0.017343f
C576 commonsourceibias.t9 gnd 0.017343f
C577 commonsourceibias.n131 gnd 0.15325f
C578 commonsourceibias.n132 gnd 0.070394f
C579 commonsourceibias.t37 gnd 0.017343f
C580 commonsourceibias.t77 gnd 0.017343f
C581 commonsourceibias.n133 gnd 0.15325f
C582 commonsourceibias.n134 gnd 0.070394f
C583 commonsourceibias.t25 gnd 0.017343f
C584 commonsourceibias.t35 gnd 0.017343f
C585 commonsourceibias.n135 gnd 0.15325f
C586 commonsourceibias.n136 gnd 0.070394f
C587 commonsourceibias.t11 gnd 0.017343f
C588 commonsourceibias.t41 gnd 0.017343f
C589 commonsourceibias.n137 gnd 0.15325f
C590 commonsourceibias.n138 gnd 0.058811f
C591 commonsourceibias.t47 gnd 0.017343f
C592 commonsourceibias.t79 gnd 0.017343f
C593 commonsourceibias.n139 gnd 0.153763f
C594 commonsourceibias.t55 gnd 0.017343f
C595 commonsourceibias.t5 gnd 0.017343f
C596 commonsourceibias.n140 gnd 0.15325f
C597 commonsourceibias.n141 gnd 0.1428f
C598 commonsourceibias.t19 gnd 0.017343f
C599 commonsourceibias.t23 gnd 0.017343f
C600 commonsourceibias.n142 gnd 0.15325f
C601 commonsourceibias.n143 gnd 0.070394f
C602 commonsourceibias.t39 gnd 0.017343f
C603 commonsourceibias.t71 gnd 0.017343f
C604 commonsourceibias.n144 gnd 0.15325f
C605 commonsourceibias.n145 gnd 0.070394f
C606 commonsourceibias.t57 gnd 0.017343f
C607 commonsourceibias.t27 gnd 0.017343f
C608 commonsourceibias.n146 gnd 0.15325f
C609 commonsourceibias.n147 gnd 0.058811f
C610 commonsourceibias.n148 gnd 0.071213f
C611 commonsourceibias.n149 gnd 0.052016f
C612 commonsourceibias.t153 gnd 0.150157f
C613 commonsourceibias.n150 gnd 0.059912f
C614 commonsourceibias.t88 gnd 0.150157f
C615 commonsourceibias.n151 gnd 0.059912f
C616 commonsourceibias.n152 gnd 0.008037f
C617 commonsourceibias.t125 gnd 0.150157f
C618 commonsourceibias.n153 gnd 0.059912f
C619 commonsourceibias.n154 gnd 0.008037f
C620 commonsourceibias.t120 gnd 0.150157f
C621 commonsourceibias.n155 gnd 0.059912f
C622 commonsourceibias.n156 gnd 0.008037f
C623 commonsourceibias.t139 gnd 0.150157f
C624 commonsourceibias.n157 gnd 0.007008f
C625 commonsourceibias.n158 gnd 0.008037f
C626 commonsourceibias.t112 gnd 0.150157f
C627 commonsourceibias.n159 gnd 0.009613f
C628 commonsourceibias.n160 gnd 0.008037f
C629 commonsourceibias.t107 gnd 0.150157f
C630 commonsourceibias.n161 gnd 0.059912f
C631 commonsourceibias.t127 gnd 0.150157f
C632 commonsourceibias.n162 gnd 0.006868f
C633 commonsourceibias.n163 gnd 0.008037f
C634 commonsourceibias.t146 gnd 0.150157f
C635 commonsourceibias.n164 gnd 0.009378f
C636 commonsourceibias.t117 gnd 0.166947f
C637 commonsourceibias.t99 gnd 0.150157f
C638 commonsourceibias.n165 gnd 0.065449f
C639 commonsourceibias.n166 gnd 0.071822f
C640 commonsourceibias.n167 gnd 0.033327f
C641 commonsourceibias.n168 gnd 0.008037f
C642 commonsourceibias.n169 gnd 0.007823f
C643 commonsourceibias.n170 gnd 0.01121f
C644 commonsourceibias.n171 gnd 0.059912f
C645 commonsourceibias.n172 gnd 0.011203f
C646 commonsourceibias.n173 gnd 0.008037f
C647 commonsourceibias.n174 gnd 0.008037f
C648 commonsourceibias.n175 gnd 0.008037f
C649 commonsourceibias.n176 gnd 0.01034f
C650 commonsourceibias.n177 gnd 0.059912f
C651 commonsourceibias.n178 gnd 0.010583f
C652 commonsourceibias.n179 gnd 0.010282f
C653 commonsourceibias.n180 gnd 0.008037f
C654 commonsourceibias.n181 gnd 0.008037f
C655 commonsourceibias.n182 gnd 0.008037f
C656 commonsourceibias.n183 gnd 0.007578f
C657 commonsourceibias.n184 gnd 0.01122f
C658 commonsourceibias.n185 gnd 0.059912f
C659 commonsourceibias.n186 gnd 0.011217f
C660 commonsourceibias.n187 gnd 0.008037f
C661 commonsourceibias.n188 gnd 0.008037f
C662 commonsourceibias.n189 gnd 0.008037f
C663 commonsourceibias.n190 gnd 0.010186f
C664 commonsourceibias.n191 gnd 0.059912f
C665 commonsourceibias.n192 gnd 0.010507f
C666 commonsourceibias.n193 gnd 0.010357f
C667 commonsourceibias.n194 gnd 0.008037f
C668 commonsourceibias.n195 gnd 0.008037f
C669 commonsourceibias.n196 gnd 0.009825f
C670 commonsourceibias.n197 gnd 0.007361f
C671 commonsourceibias.n198 gnd 0.011225f
C672 commonsourceibias.n199 gnd 0.008037f
C673 commonsourceibias.n200 gnd 0.008037f
C674 commonsourceibias.n201 gnd 0.011224f
C675 commonsourceibias.n202 gnd 0.007172f
C676 commonsourceibias.n203 gnd 0.010015f
C677 commonsourceibias.n204 gnd 0.008037f
C678 commonsourceibias.n205 gnd 0.007021f
C679 commonsourceibias.n206 gnd 0.010432f
C680 commonsourceibias.n207 gnd 0.010432f
C681 commonsourceibias.n208 gnd 0.007021f
C682 commonsourceibias.n209 gnd 0.008037f
C683 commonsourceibias.n210 gnd 0.008037f
C684 commonsourceibias.n211 gnd 0.007172f
C685 commonsourceibias.n212 gnd 0.011224f
C686 commonsourceibias.n213 gnd 0.059912f
C687 commonsourceibias.n214 gnd 0.011225f
C688 commonsourceibias.n215 gnd 0.008037f
C689 commonsourceibias.n216 gnd 0.008037f
C690 commonsourceibias.n217 gnd 0.008037f
C691 commonsourceibias.n218 gnd 0.009825f
C692 commonsourceibias.n219 gnd 0.059912f
C693 commonsourceibias.n220 gnd 0.010357f
C694 commonsourceibias.n221 gnd 0.010507f
C695 commonsourceibias.n222 gnd 0.008037f
C696 commonsourceibias.n223 gnd 0.008037f
C697 commonsourceibias.n224 gnd 0.008037f
C698 commonsourceibias.n225 gnd 0.007008f
C699 commonsourceibias.n226 gnd 0.011217f
C700 commonsourceibias.n227 gnd 0.059912f
C701 commonsourceibias.n228 gnd 0.01122f
C702 commonsourceibias.n229 gnd 0.008037f
C703 commonsourceibias.n230 gnd 0.008037f
C704 commonsourceibias.n231 gnd 0.008037f
C705 commonsourceibias.n232 gnd 0.009613f
C706 commonsourceibias.n233 gnd 0.059912f
C707 commonsourceibias.n234 gnd 0.010282f
C708 commonsourceibias.n235 gnd 0.010583f
C709 commonsourceibias.n236 gnd 0.008037f
C710 commonsourceibias.n237 gnd 0.008037f
C711 commonsourceibias.n238 gnd 0.008037f
C712 commonsourceibias.n239 gnd 0.006868f
C713 commonsourceibias.n240 gnd 0.011203f
C714 commonsourceibias.n241 gnd 0.059912f
C715 commonsourceibias.n242 gnd 0.01121f
C716 commonsourceibias.n243 gnd 0.008037f
C717 commonsourceibias.n244 gnd 0.008037f
C718 commonsourceibias.n245 gnd 0.008037f
C719 commonsourceibias.n246 gnd 0.009378f
C720 commonsourceibias.n247 gnd 0.059912f
C721 commonsourceibias.n248 gnd 0.009861f
C722 commonsourceibias.n249 gnd 0.07189f
C723 commonsourceibias.n250 gnd 0.04697f
C724 commonsourceibias.n251 gnd 0.010724f
C725 commonsourceibias.t119 gnd 0.150157f
C726 commonsourceibias.n252 gnd 0.007823f
C727 commonsourceibias.n253 gnd 0.008037f
C728 commonsourceibias.t137 gnd 0.150157f
C729 commonsourceibias.n254 gnd 0.01034f
C730 commonsourceibias.n255 gnd 0.008037f
C731 commonsourceibias.t92 gnd 0.150157f
C732 commonsourceibias.n256 gnd 0.059912f
C733 commonsourceibias.t109 gnd 0.150157f
C734 commonsourceibias.n257 gnd 0.007578f
C735 commonsourceibias.n258 gnd 0.008037f
C736 commonsourceibias.t128 gnd 0.150157f
C737 commonsourceibias.n259 gnd 0.010186f
C738 commonsourceibias.n260 gnd 0.008037f
C739 commonsourceibias.t86 gnd 0.150157f
C740 commonsourceibias.n261 gnd 0.059912f
C741 commonsourceibias.t83 gnd 0.150157f
C742 commonsourceibias.n262 gnd 0.007361f
C743 commonsourceibias.n263 gnd 0.008037f
C744 commonsourceibias.t118 gnd 0.150157f
C745 commonsourceibias.n264 gnd 0.010015f
C746 commonsourceibias.n265 gnd 0.008037f
C747 commonsourceibias.t138 gnd 0.150157f
C748 commonsourceibias.n266 gnd 0.059912f
C749 commonsourceibias.t159 gnd 0.150157f
C750 commonsourceibias.n267 gnd 0.007172f
C751 commonsourceibias.n268 gnd 0.008037f
C752 commonsourceibias.t108 gnd 0.150157f
C753 commonsourceibias.n269 gnd 0.009825f
C754 commonsourceibias.n270 gnd 0.008037f
C755 commonsourceibias.t102 gnd 0.150157f
C756 commonsourceibias.n271 gnd 0.059912f
C757 commonsourceibias.t121 gnd 0.150157f
C758 commonsourceibias.n272 gnd 0.007008f
C759 commonsourceibias.n273 gnd 0.008037f
C760 commonsourceibias.t95 gnd 0.150157f
C761 commonsourceibias.n274 gnd 0.009613f
C762 commonsourceibias.n275 gnd 0.008037f
C763 commonsourceibias.t93 gnd 0.150157f
C764 commonsourceibias.n276 gnd 0.059912f
C765 commonsourceibias.t110 gnd 0.150157f
C766 commonsourceibias.n277 gnd 0.006868f
C767 commonsourceibias.n278 gnd 0.008037f
C768 commonsourceibias.t129 gnd 0.150157f
C769 commonsourceibias.n279 gnd 0.009378f
C770 commonsourceibias.t101 gnd 0.166947f
C771 commonsourceibias.t87 gnd 0.150157f
C772 commonsourceibias.n280 gnd 0.065449f
C773 commonsourceibias.n281 gnd 0.071822f
C774 commonsourceibias.n282 gnd 0.033327f
C775 commonsourceibias.n283 gnd 0.008037f
C776 commonsourceibias.n284 gnd 0.007823f
C777 commonsourceibias.n285 gnd 0.01121f
C778 commonsourceibias.n286 gnd 0.059912f
C779 commonsourceibias.n287 gnd 0.011203f
C780 commonsourceibias.n288 gnd 0.008037f
C781 commonsourceibias.n289 gnd 0.008037f
C782 commonsourceibias.n290 gnd 0.008037f
C783 commonsourceibias.n291 gnd 0.01034f
C784 commonsourceibias.n292 gnd 0.059912f
C785 commonsourceibias.n293 gnd 0.010583f
C786 commonsourceibias.n294 gnd 0.010282f
C787 commonsourceibias.n295 gnd 0.008037f
C788 commonsourceibias.n296 gnd 0.008037f
C789 commonsourceibias.n297 gnd 0.008037f
C790 commonsourceibias.n298 gnd 0.007578f
C791 commonsourceibias.n299 gnd 0.01122f
C792 commonsourceibias.n300 gnd 0.059912f
C793 commonsourceibias.n301 gnd 0.011217f
C794 commonsourceibias.n302 gnd 0.008037f
C795 commonsourceibias.n303 gnd 0.008037f
C796 commonsourceibias.n304 gnd 0.008037f
C797 commonsourceibias.n305 gnd 0.010186f
C798 commonsourceibias.n306 gnd 0.059912f
C799 commonsourceibias.n307 gnd 0.010507f
C800 commonsourceibias.n308 gnd 0.010357f
C801 commonsourceibias.n309 gnd 0.008037f
C802 commonsourceibias.n310 gnd 0.008037f
C803 commonsourceibias.n311 gnd 0.008037f
C804 commonsourceibias.n312 gnd 0.007361f
C805 commonsourceibias.n313 gnd 0.011225f
C806 commonsourceibias.n314 gnd 0.059912f
C807 commonsourceibias.n315 gnd 0.011224f
C808 commonsourceibias.n316 gnd 0.008037f
C809 commonsourceibias.n317 gnd 0.008037f
C810 commonsourceibias.n318 gnd 0.008037f
C811 commonsourceibias.n319 gnd 0.010015f
C812 commonsourceibias.n320 gnd 0.059912f
C813 commonsourceibias.n321 gnd 0.010432f
C814 commonsourceibias.n322 gnd 0.010432f
C815 commonsourceibias.n323 gnd 0.008037f
C816 commonsourceibias.n324 gnd 0.008037f
C817 commonsourceibias.n325 gnd 0.008037f
C818 commonsourceibias.n326 gnd 0.007172f
C819 commonsourceibias.n327 gnd 0.011224f
C820 commonsourceibias.n328 gnd 0.059912f
C821 commonsourceibias.n329 gnd 0.011225f
C822 commonsourceibias.n330 gnd 0.008037f
C823 commonsourceibias.n331 gnd 0.008037f
C824 commonsourceibias.n332 gnd 0.008037f
C825 commonsourceibias.n333 gnd 0.009825f
C826 commonsourceibias.n334 gnd 0.059912f
C827 commonsourceibias.n335 gnd 0.010357f
C828 commonsourceibias.n336 gnd 0.010507f
C829 commonsourceibias.n337 gnd 0.008037f
C830 commonsourceibias.n338 gnd 0.008037f
C831 commonsourceibias.n339 gnd 0.008037f
C832 commonsourceibias.n340 gnd 0.007008f
C833 commonsourceibias.n341 gnd 0.011217f
C834 commonsourceibias.n342 gnd 0.059912f
C835 commonsourceibias.n343 gnd 0.01122f
C836 commonsourceibias.n344 gnd 0.008037f
C837 commonsourceibias.n345 gnd 0.008037f
C838 commonsourceibias.n346 gnd 0.008037f
C839 commonsourceibias.n347 gnd 0.009613f
C840 commonsourceibias.n348 gnd 0.059912f
C841 commonsourceibias.n349 gnd 0.010282f
C842 commonsourceibias.n350 gnd 0.010583f
C843 commonsourceibias.n351 gnd 0.008037f
C844 commonsourceibias.n352 gnd 0.008037f
C845 commonsourceibias.n353 gnd 0.008037f
C846 commonsourceibias.n354 gnd 0.006868f
C847 commonsourceibias.n355 gnd 0.011203f
C848 commonsourceibias.n356 gnd 0.059912f
C849 commonsourceibias.n357 gnd 0.01121f
C850 commonsourceibias.n358 gnd 0.008037f
C851 commonsourceibias.n359 gnd 0.008037f
C852 commonsourceibias.n360 gnd 0.008037f
C853 commonsourceibias.n361 gnd 0.009378f
C854 commonsourceibias.n362 gnd 0.059912f
C855 commonsourceibias.n363 gnd 0.009861f
C856 commonsourceibias.t100 gnd 0.162395f
C857 commonsourceibias.n364 gnd 0.07189f
C858 commonsourceibias.n365 gnd 0.025003f
C859 commonsourceibias.n366 gnd 0.464917f
C860 commonsourceibias.n367 gnd 0.010724f
C861 commonsourceibias.t140 gnd 0.162395f
C862 commonsourceibias.t155 gnd 0.150157f
C863 commonsourceibias.n368 gnd 0.007823f
C864 commonsourceibias.n369 gnd 0.008037f
C865 commonsourceibias.t84 gnd 0.150157f
C866 commonsourceibias.n370 gnd 0.01034f
C867 commonsourceibias.n371 gnd 0.008037f
C868 commonsourceibias.t148 gnd 0.150157f
C869 commonsourceibias.n372 gnd 0.007578f
C870 commonsourceibias.n373 gnd 0.008037f
C871 commonsourceibias.t80 gnd 0.150157f
C872 commonsourceibias.n374 gnd 0.010186f
C873 commonsourceibias.n375 gnd 0.008037f
C874 commonsourceibias.t113 gnd 0.150157f
C875 commonsourceibias.n376 gnd 0.007361f
C876 commonsourceibias.n377 gnd 0.008037f
C877 commonsourceibias.t154 gnd 0.150157f
C878 commonsourceibias.n378 gnd 0.010015f
C879 commonsourceibias.t29 gnd 0.017343f
C880 commonsourceibias.t3 gnd 0.017343f
C881 commonsourceibias.n379 gnd 0.153763f
C882 commonsourceibias.t49 gnd 0.017343f
C883 commonsourceibias.t13 gnd 0.017343f
C884 commonsourceibias.n380 gnd 0.15325f
C885 commonsourceibias.n381 gnd 0.1428f
C886 commonsourceibias.t69 gnd 0.017343f
C887 commonsourceibias.t67 gnd 0.017343f
C888 commonsourceibias.n382 gnd 0.15325f
C889 commonsourceibias.n383 gnd 0.070394f
C890 commonsourceibias.t7 gnd 0.017343f
C891 commonsourceibias.t63 gnd 0.017343f
C892 commonsourceibias.n384 gnd 0.15325f
C893 commonsourceibias.n385 gnd 0.070394f
C894 commonsourceibias.t53 gnd 0.017343f
C895 commonsourceibias.t73 gnd 0.017343f
C896 commonsourceibias.n386 gnd 0.15325f
C897 commonsourceibias.n387 gnd 0.058811f
C898 commonsourceibias.n388 gnd 0.010724f
C899 commonsourceibias.t42 gnd 0.150157f
C900 commonsourceibias.n389 gnd 0.007823f
C901 commonsourceibias.n390 gnd 0.008037f
C902 commonsourceibias.t0 gnd 0.150157f
C903 commonsourceibias.n391 gnd 0.01034f
C904 commonsourceibias.n392 gnd 0.008037f
C905 commonsourceibias.t60 gnd 0.150157f
C906 commonsourceibias.n393 gnd 0.007578f
C907 commonsourceibias.n394 gnd 0.008037f
C908 commonsourceibias.t16 gnd 0.150157f
C909 commonsourceibias.n395 gnd 0.010186f
C910 commonsourceibias.n396 gnd 0.008037f
C911 commonsourceibias.t58 gnd 0.150157f
C912 commonsourceibias.n397 gnd 0.007361f
C913 commonsourceibias.n398 gnd 0.008037f
C914 commonsourceibias.t32 gnd 0.150157f
C915 commonsourceibias.n399 gnd 0.010015f
C916 commonsourceibias.n400 gnd 0.008037f
C917 commonsourceibias.t72 gnd 0.150157f
C918 commonsourceibias.n401 gnd 0.007172f
C919 commonsourceibias.n402 gnd 0.008037f
C920 commonsourceibias.t52 gnd 0.150157f
C921 commonsourceibias.n403 gnd 0.009825f
C922 commonsourceibias.n404 gnd 0.008037f
C923 commonsourceibias.t6 gnd 0.150157f
C924 commonsourceibias.n405 gnd 0.007008f
C925 commonsourceibias.n406 gnd 0.008037f
C926 commonsourceibias.t66 gnd 0.150157f
C927 commonsourceibias.n407 gnd 0.009613f
C928 commonsourceibias.n408 gnd 0.008037f
C929 commonsourceibias.t12 gnd 0.150157f
C930 commonsourceibias.n409 gnd 0.006868f
C931 commonsourceibias.n410 gnd 0.008037f
C932 commonsourceibias.t48 gnd 0.150157f
C933 commonsourceibias.n411 gnd 0.009378f
C934 commonsourceibias.t28 gnd 0.166947f
C935 commonsourceibias.t2 gnd 0.150157f
C936 commonsourceibias.n412 gnd 0.065449f
C937 commonsourceibias.n413 gnd 0.071822f
C938 commonsourceibias.n414 gnd 0.033327f
C939 commonsourceibias.n415 gnd 0.008037f
C940 commonsourceibias.n416 gnd 0.007823f
C941 commonsourceibias.n417 gnd 0.01121f
C942 commonsourceibias.n418 gnd 0.059912f
C943 commonsourceibias.n419 gnd 0.011203f
C944 commonsourceibias.n420 gnd 0.008037f
C945 commonsourceibias.n421 gnd 0.008037f
C946 commonsourceibias.n422 gnd 0.008037f
C947 commonsourceibias.n423 gnd 0.01034f
C948 commonsourceibias.n424 gnd 0.059912f
C949 commonsourceibias.n425 gnd 0.010583f
C950 commonsourceibias.t68 gnd 0.150157f
C951 commonsourceibias.n426 gnd 0.059912f
C952 commonsourceibias.n427 gnd 0.010282f
C953 commonsourceibias.n428 gnd 0.008037f
C954 commonsourceibias.n429 gnd 0.008037f
C955 commonsourceibias.n430 gnd 0.008037f
C956 commonsourceibias.n431 gnd 0.007578f
C957 commonsourceibias.n432 gnd 0.01122f
C958 commonsourceibias.n433 gnd 0.059912f
C959 commonsourceibias.n434 gnd 0.011217f
C960 commonsourceibias.n435 gnd 0.008037f
C961 commonsourceibias.n436 gnd 0.008037f
C962 commonsourceibias.n437 gnd 0.008037f
C963 commonsourceibias.n438 gnd 0.010186f
C964 commonsourceibias.n439 gnd 0.059912f
C965 commonsourceibias.n440 gnd 0.010507f
C966 commonsourceibias.t62 gnd 0.150157f
C967 commonsourceibias.n441 gnd 0.059912f
C968 commonsourceibias.n442 gnd 0.010357f
C969 commonsourceibias.n443 gnd 0.008037f
C970 commonsourceibias.n444 gnd 0.008037f
C971 commonsourceibias.n445 gnd 0.008037f
C972 commonsourceibias.n446 gnd 0.007361f
C973 commonsourceibias.n447 gnd 0.011225f
C974 commonsourceibias.n448 gnd 0.059912f
C975 commonsourceibias.n449 gnd 0.011224f
C976 commonsourceibias.n450 gnd 0.008037f
C977 commonsourceibias.n451 gnd 0.008037f
C978 commonsourceibias.n452 gnd 0.008037f
C979 commonsourceibias.n453 gnd 0.010015f
C980 commonsourceibias.n454 gnd 0.059912f
C981 commonsourceibias.n455 gnd 0.010432f
C982 commonsourceibias.t64 gnd 0.150157f
C983 commonsourceibias.n456 gnd 0.059912f
C984 commonsourceibias.n457 gnd 0.010432f
C985 commonsourceibias.n458 gnd 0.008037f
C986 commonsourceibias.n459 gnd 0.008037f
C987 commonsourceibias.n460 gnd 0.008037f
C988 commonsourceibias.n461 gnd 0.007172f
C989 commonsourceibias.n462 gnd 0.011224f
C990 commonsourceibias.n463 gnd 0.059912f
C991 commonsourceibias.n464 gnd 0.011225f
C992 commonsourceibias.n465 gnd 0.008037f
C993 commonsourceibias.n466 gnd 0.008037f
C994 commonsourceibias.n467 gnd 0.008037f
C995 commonsourceibias.n468 gnd 0.009825f
C996 commonsourceibias.n469 gnd 0.059912f
C997 commonsourceibias.n470 gnd 0.010357f
C998 commonsourceibias.t44 gnd 0.150157f
C999 commonsourceibias.n471 gnd 0.059912f
C1000 commonsourceibias.n472 gnd 0.010507f
C1001 commonsourceibias.n473 gnd 0.008037f
C1002 commonsourceibias.n474 gnd 0.008037f
C1003 commonsourceibias.n475 gnd 0.008037f
C1004 commonsourceibias.n476 gnd 0.007008f
C1005 commonsourceibias.n477 gnd 0.011217f
C1006 commonsourceibias.n478 gnd 0.059912f
C1007 commonsourceibias.n479 gnd 0.01122f
C1008 commonsourceibias.n480 gnd 0.008037f
C1009 commonsourceibias.n481 gnd 0.008037f
C1010 commonsourceibias.n482 gnd 0.008037f
C1011 commonsourceibias.n483 gnd 0.009613f
C1012 commonsourceibias.n484 gnd 0.059912f
C1013 commonsourceibias.n485 gnd 0.010282f
C1014 commonsourceibias.t30 gnd 0.150157f
C1015 commonsourceibias.n486 gnd 0.059912f
C1016 commonsourceibias.n487 gnd 0.010583f
C1017 commonsourceibias.n488 gnd 0.008037f
C1018 commonsourceibias.n489 gnd 0.008037f
C1019 commonsourceibias.n490 gnd 0.008037f
C1020 commonsourceibias.n491 gnd 0.006868f
C1021 commonsourceibias.n492 gnd 0.011203f
C1022 commonsourceibias.n493 gnd 0.059912f
C1023 commonsourceibias.n494 gnd 0.01121f
C1024 commonsourceibias.n495 gnd 0.008037f
C1025 commonsourceibias.n496 gnd 0.008037f
C1026 commonsourceibias.n497 gnd 0.008037f
C1027 commonsourceibias.n498 gnd 0.009378f
C1028 commonsourceibias.n499 gnd 0.059912f
C1029 commonsourceibias.n500 gnd 0.009861f
C1030 commonsourceibias.t14 gnd 0.162395f
C1031 commonsourceibias.n501 gnd 0.07189f
C1032 commonsourceibias.n502 gnd 0.080075f
C1033 commonsourceibias.t43 gnd 0.017343f
C1034 commonsourceibias.t15 gnd 0.017343f
C1035 commonsourceibias.n503 gnd 0.15325f
C1036 commonsourceibias.n504 gnd 0.132562f
C1037 commonsourceibias.t31 gnd 0.017343f
C1038 commonsourceibias.t1 gnd 0.017343f
C1039 commonsourceibias.n505 gnd 0.15325f
C1040 commonsourceibias.n506 gnd 0.070394f
C1041 commonsourceibias.t17 gnd 0.017343f
C1042 commonsourceibias.t61 gnd 0.017343f
C1043 commonsourceibias.n507 gnd 0.15325f
C1044 commonsourceibias.n508 gnd 0.070394f
C1045 commonsourceibias.t59 gnd 0.017343f
C1046 commonsourceibias.t45 gnd 0.017343f
C1047 commonsourceibias.n509 gnd 0.15325f
C1048 commonsourceibias.n510 gnd 0.070394f
C1049 commonsourceibias.t65 gnd 0.017343f
C1050 commonsourceibias.t33 gnd 0.017343f
C1051 commonsourceibias.n511 gnd 0.15325f
C1052 commonsourceibias.n512 gnd 0.058811f
C1053 commonsourceibias.n513 gnd 0.071213f
C1054 commonsourceibias.n514 gnd 0.052016f
C1055 commonsourceibias.t82 gnd 0.150157f
C1056 commonsourceibias.n515 gnd 0.059912f
C1057 commonsourceibias.n516 gnd 0.008037f
C1058 commonsourceibias.t147 gnd 0.150157f
C1059 commonsourceibias.n517 gnd 0.059912f
C1060 commonsourceibias.n518 gnd 0.008037f
C1061 commonsourceibias.t143 gnd 0.150157f
C1062 commonsourceibias.n519 gnd 0.059912f
C1063 commonsourceibias.n520 gnd 0.008037f
C1064 commonsourceibias.t158 gnd 0.150157f
C1065 commonsourceibias.n521 gnd 0.007008f
C1066 commonsourceibias.n522 gnd 0.008037f
C1067 commonsourceibias.t104 gnd 0.150157f
C1068 commonsourceibias.n523 gnd 0.009613f
C1069 commonsourceibias.n524 gnd 0.008037f
C1070 commonsourceibias.t133 gnd 0.150157f
C1071 commonsourceibias.n525 gnd 0.006868f
C1072 commonsourceibias.n526 gnd 0.008037f
C1073 commonsourceibias.t150 gnd 0.150157f
C1074 commonsourceibias.n527 gnd 0.009378f
C1075 commonsourceibias.t123 gnd 0.166947f
C1076 commonsourceibias.t103 gnd 0.150157f
C1077 commonsourceibias.n528 gnd 0.065449f
C1078 commonsourceibias.n529 gnd 0.071822f
C1079 commonsourceibias.n530 gnd 0.033327f
C1080 commonsourceibias.n531 gnd 0.008037f
C1081 commonsourceibias.n532 gnd 0.007823f
C1082 commonsourceibias.n533 gnd 0.01121f
C1083 commonsourceibias.n534 gnd 0.059912f
C1084 commonsourceibias.n535 gnd 0.011203f
C1085 commonsourceibias.n536 gnd 0.008037f
C1086 commonsourceibias.n537 gnd 0.008037f
C1087 commonsourceibias.n538 gnd 0.008037f
C1088 commonsourceibias.n539 gnd 0.01034f
C1089 commonsourceibias.n540 gnd 0.059912f
C1090 commonsourceibias.n541 gnd 0.010583f
C1091 commonsourceibias.t114 gnd 0.150157f
C1092 commonsourceibias.n542 gnd 0.059912f
C1093 commonsourceibias.n543 gnd 0.010282f
C1094 commonsourceibias.n544 gnd 0.008037f
C1095 commonsourceibias.n545 gnd 0.008037f
C1096 commonsourceibias.n546 gnd 0.008037f
C1097 commonsourceibias.n547 gnd 0.007578f
C1098 commonsourceibias.n548 gnd 0.01122f
C1099 commonsourceibias.n549 gnd 0.059912f
C1100 commonsourceibias.n550 gnd 0.011217f
C1101 commonsourceibias.n551 gnd 0.008037f
C1102 commonsourceibias.n552 gnd 0.008037f
C1103 commonsourceibias.n553 gnd 0.008037f
C1104 commonsourceibias.n554 gnd 0.010186f
C1105 commonsourceibias.n555 gnd 0.059912f
C1106 commonsourceibias.n556 gnd 0.010507f
C1107 commonsourceibias.n557 gnd 0.010357f
C1108 commonsourceibias.n558 gnd 0.008037f
C1109 commonsourceibias.n559 gnd 0.008037f
C1110 commonsourceibias.n560 gnd 0.009825f
C1111 commonsourceibias.n561 gnd 0.007361f
C1112 commonsourceibias.n562 gnd 0.011225f
C1113 commonsourceibias.n563 gnd 0.008037f
C1114 commonsourceibias.n564 gnd 0.008037f
C1115 commonsourceibias.n565 gnd 0.011224f
C1116 commonsourceibias.n566 gnd 0.007172f
C1117 commonsourceibias.n567 gnd 0.010015f
C1118 commonsourceibias.n568 gnd 0.008037f
C1119 commonsourceibias.n569 gnd 0.007021f
C1120 commonsourceibias.n570 gnd 0.010432f
C1121 commonsourceibias.t85 gnd 0.150157f
C1122 commonsourceibias.n571 gnd 0.059912f
C1123 commonsourceibias.n572 gnd 0.010432f
C1124 commonsourceibias.n573 gnd 0.007021f
C1125 commonsourceibias.n574 gnd 0.008037f
C1126 commonsourceibias.n575 gnd 0.008037f
C1127 commonsourceibias.n576 gnd 0.007172f
C1128 commonsourceibias.n577 gnd 0.011224f
C1129 commonsourceibias.n578 gnd 0.059912f
C1130 commonsourceibias.n579 gnd 0.011225f
C1131 commonsourceibias.n580 gnd 0.008037f
C1132 commonsourceibias.n581 gnd 0.008037f
C1133 commonsourceibias.n582 gnd 0.008037f
C1134 commonsourceibias.n583 gnd 0.009825f
C1135 commonsourceibias.n584 gnd 0.059912f
C1136 commonsourceibias.n585 gnd 0.010357f
C1137 commonsourceibias.t89 gnd 0.150157f
C1138 commonsourceibias.n586 gnd 0.059912f
C1139 commonsourceibias.n587 gnd 0.010507f
C1140 commonsourceibias.n588 gnd 0.008037f
C1141 commonsourceibias.n589 gnd 0.008037f
C1142 commonsourceibias.n590 gnd 0.008037f
C1143 commonsourceibias.n591 gnd 0.007008f
C1144 commonsourceibias.n592 gnd 0.011217f
C1145 commonsourceibias.n593 gnd 0.059912f
C1146 commonsourceibias.n594 gnd 0.01122f
C1147 commonsourceibias.n595 gnd 0.008037f
C1148 commonsourceibias.n596 gnd 0.008037f
C1149 commonsourceibias.n597 gnd 0.008037f
C1150 commonsourceibias.n598 gnd 0.009613f
C1151 commonsourceibias.n599 gnd 0.059912f
C1152 commonsourceibias.n600 gnd 0.010282f
C1153 commonsourceibias.t130 gnd 0.150157f
C1154 commonsourceibias.n601 gnd 0.059912f
C1155 commonsourceibias.n602 gnd 0.010583f
C1156 commonsourceibias.n603 gnd 0.008037f
C1157 commonsourceibias.n604 gnd 0.008037f
C1158 commonsourceibias.n605 gnd 0.008037f
C1159 commonsourceibias.n606 gnd 0.006868f
C1160 commonsourceibias.n607 gnd 0.011203f
C1161 commonsourceibias.n608 gnd 0.059912f
C1162 commonsourceibias.n609 gnd 0.01121f
C1163 commonsourceibias.n610 gnd 0.008037f
C1164 commonsourceibias.n611 gnd 0.008037f
C1165 commonsourceibias.n612 gnd 0.008037f
C1166 commonsourceibias.n613 gnd 0.009378f
C1167 commonsourceibias.n614 gnd 0.059912f
C1168 commonsourceibias.n615 gnd 0.009861f
C1169 commonsourceibias.n616 gnd 0.07189f
C1170 commonsourceibias.n617 gnd 0.04697f
C1171 commonsourceibias.n618 gnd 0.010724f
C1172 commonsourceibias.t142 gnd 0.150157f
C1173 commonsourceibias.n619 gnd 0.007823f
C1174 commonsourceibias.n620 gnd 0.008037f
C1175 commonsourceibias.t156 gnd 0.150157f
C1176 commonsourceibias.n621 gnd 0.01034f
C1177 commonsourceibias.n622 gnd 0.008037f
C1178 commonsourceibias.t132 gnd 0.150157f
C1179 commonsourceibias.n623 gnd 0.007578f
C1180 commonsourceibias.n624 gnd 0.008037f
C1181 commonsourceibias.t149 gnd 0.150157f
C1182 commonsourceibias.n625 gnd 0.010186f
C1183 commonsourceibias.n626 gnd 0.008037f
C1184 commonsourceibias.t97 gnd 0.150157f
C1185 commonsourceibias.n627 gnd 0.007361f
C1186 commonsourceibias.n628 gnd 0.008037f
C1187 commonsourceibias.t141 gnd 0.150157f
C1188 commonsourceibias.n629 gnd 0.010015f
C1189 commonsourceibias.n630 gnd 0.008037f
C1190 commonsourceibias.t152 gnd 0.150157f
C1191 commonsourceibias.n631 gnd 0.007172f
C1192 commonsourceibias.n632 gnd 0.008037f
C1193 commonsourceibias.t131 gnd 0.150157f
C1194 commonsourceibias.n633 gnd 0.009825f
C1195 commonsourceibias.n634 gnd 0.008037f
C1196 commonsourceibias.t145 gnd 0.150157f
C1197 commonsourceibias.n635 gnd 0.007008f
C1198 commonsourceibias.n636 gnd 0.008037f
C1199 commonsourceibias.t91 gnd 0.150157f
C1200 commonsourceibias.n637 gnd 0.009613f
C1201 commonsourceibias.n638 gnd 0.008037f
C1202 commonsourceibias.t116 gnd 0.150157f
C1203 commonsourceibias.n639 gnd 0.006868f
C1204 commonsourceibias.n640 gnd 0.008037f
C1205 commonsourceibias.t134 gnd 0.150157f
C1206 commonsourceibias.n641 gnd 0.009378f
C1207 commonsourceibias.t106 gnd 0.166947f
C1208 commonsourceibias.t90 gnd 0.150157f
C1209 commonsourceibias.n642 gnd 0.065449f
C1210 commonsourceibias.n643 gnd 0.071822f
C1211 commonsourceibias.n644 gnd 0.033327f
C1212 commonsourceibias.n645 gnd 0.008037f
C1213 commonsourceibias.n646 gnd 0.007823f
C1214 commonsourceibias.n647 gnd 0.01121f
C1215 commonsourceibias.n648 gnd 0.059912f
C1216 commonsourceibias.n649 gnd 0.011203f
C1217 commonsourceibias.n650 gnd 0.008037f
C1218 commonsourceibias.n651 gnd 0.008037f
C1219 commonsourceibias.n652 gnd 0.008037f
C1220 commonsourceibias.n653 gnd 0.01034f
C1221 commonsourceibias.n654 gnd 0.059912f
C1222 commonsourceibias.n655 gnd 0.010583f
C1223 commonsourceibias.t96 gnd 0.150157f
C1224 commonsourceibias.n656 gnd 0.059912f
C1225 commonsourceibias.n657 gnd 0.010282f
C1226 commonsourceibias.n658 gnd 0.008037f
C1227 commonsourceibias.n659 gnd 0.008037f
C1228 commonsourceibias.n660 gnd 0.008037f
C1229 commonsourceibias.n661 gnd 0.007578f
C1230 commonsourceibias.n662 gnd 0.01122f
C1231 commonsourceibias.n663 gnd 0.059912f
C1232 commonsourceibias.n664 gnd 0.011217f
C1233 commonsourceibias.n665 gnd 0.008037f
C1234 commonsourceibias.n666 gnd 0.008037f
C1235 commonsourceibias.n667 gnd 0.008037f
C1236 commonsourceibias.n668 gnd 0.010186f
C1237 commonsourceibias.n669 gnd 0.059912f
C1238 commonsourceibias.n670 gnd 0.010507f
C1239 commonsourceibias.t124 gnd 0.150157f
C1240 commonsourceibias.n671 gnd 0.059912f
C1241 commonsourceibias.n672 gnd 0.010357f
C1242 commonsourceibias.n673 gnd 0.008037f
C1243 commonsourceibias.n674 gnd 0.008037f
C1244 commonsourceibias.n675 gnd 0.008037f
C1245 commonsourceibias.n676 gnd 0.007361f
C1246 commonsourceibias.n677 gnd 0.011225f
C1247 commonsourceibias.n678 gnd 0.059912f
C1248 commonsourceibias.n679 gnd 0.011224f
C1249 commonsourceibias.n680 gnd 0.008037f
C1250 commonsourceibias.n681 gnd 0.008037f
C1251 commonsourceibias.n682 gnd 0.008037f
C1252 commonsourceibias.n683 gnd 0.010015f
C1253 commonsourceibias.n684 gnd 0.059912f
C1254 commonsourceibias.n685 gnd 0.010432f
C1255 commonsourceibias.t157 gnd 0.150157f
C1256 commonsourceibias.n686 gnd 0.059912f
C1257 commonsourceibias.n687 gnd 0.010432f
C1258 commonsourceibias.n688 gnd 0.008037f
C1259 commonsourceibias.n689 gnd 0.008037f
C1260 commonsourceibias.n690 gnd 0.008037f
C1261 commonsourceibias.n691 gnd 0.007172f
C1262 commonsourceibias.n692 gnd 0.011224f
C1263 commonsourceibias.n693 gnd 0.059912f
C1264 commonsourceibias.n694 gnd 0.011225f
C1265 commonsourceibias.n695 gnd 0.008037f
C1266 commonsourceibias.n696 gnd 0.008037f
C1267 commonsourceibias.n697 gnd 0.008037f
C1268 commonsourceibias.n698 gnd 0.009825f
C1269 commonsourceibias.n699 gnd 0.059912f
C1270 commonsourceibias.n700 gnd 0.010357f
C1271 commonsourceibias.t81 gnd 0.150157f
C1272 commonsourceibias.n701 gnd 0.059912f
C1273 commonsourceibias.n702 gnd 0.010507f
C1274 commonsourceibias.n703 gnd 0.008037f
C1275 commonsourceibias.n704 gnd 0.008037f
C1276 commonsourceibias.n705 gnd 0.008037f
C1277 commonsourceibias.n706 gnd 0.007008f
C1278 commonsourceibias.n707 gnd 0.011217f
C1279 commonsourceibias.n708 gnd 0.059912f
C1280 commonsourceibias.n709 gnd 0.01122f
C1281 commonsourceibias.n710 gnd 0.008037f
C1282 commonsourceibias.n711 gnd 0.008037f
C1283 commonsourceibias.n712 gnd 0.008037f
C1284 commonsourceibias.n713 gnd 0.009613f
C1285 commonsourceibias.n714 gnd 0.059912f
C1286 commonsourceibias.n715 gnd 0.010282f
C1287 commonsourceibias.t111 gnd 0.150157f
C1288 commonsourceibias.n716 gnd 0.059912f
C1289 commonsourceibias.n717 gnd 0.010583f
C1290 commonsourceibias.n718 gnd 0.008037f
C1291 commonsourceibias.n719 gnd 0.008037f
C1292 commonsourceibias.n720 gnd 0.008037f
C1293 commonsourceibias.n721 gnd 0.006868f
C1294 commonsourceibias.n722 gnd 0.011203f
C1295 commonsourceibias.n723 gnd 0.059912f
C1296 commonsourceibias.n724 gnd 0.01121f
C1297 commonsourceibias.n725 gnd 0.008037f
C1298 commonsourceibias.n726 gnd 0.008037f
C1299 commonsourceibias.n727 gnd 0.008037f
C1300 commonsourceibias.n728 gnd 0.009378f
C1301 commonsourceibias.n729 gnd 0.059912f
C1302 commonsourceibias.n730 gnd 0.009861f
C1303 commonsourceibias.t122 gnd 0.162395f
C1304 commonsourceibias.n731 gnd 0.07189f
C1305 commonsourceibias.n732 gnd 0.025003f
C1306 commonsourceibias.n733 gnd 0.221951f
C1307 commonsourceibias.n734 gnd 4.85761f
C1308 a_n3827_n3924.n0 gnd 0.899874f
C1309 a_n3827_n3924.t47 gnd 1.00187f
C1310 a_n3827_n3924.n1 gnd 0.864582f
C1311 a_n3827_n3924.t31 gnd 0.096397f
C1312 a_n3827_n3924.t25 gnd 0.096397f
C1313 a_n3827_n3924.n2 gnd 0.787293f
C1314 a_n3827_n3924.n3 gnd 0.319299f
C1315 a_n3827_n3924.t38 gnd 0.096397f
C1316 a_n3827_n3924.t42 gnd 0.096397f
C1317 a_n3827_n3924.n4 gnd 0.787293f
C1318 a_n3827_n3924.n5 gnd 0.319299f
C1319 a_n3827_n3924.t2 gnd 0.096397f
C1320 a_n3827_n3924.t28 gnd 0.096397f
C1321 a_n3827_n3924.n6 gnd 0.787293f
C1322 a_n3827_n3924.n7 gnd 0.319299f
C1323 a_n3827_n3924.t46 gnd 0.096397f
C1324 a_n3827_n3924.t29 gnd 0.096397f
C1325 a_n3827_n3924.n8 gnd 0.787293f
C1326 a_n3827_n3924.n9 gnd 0.319299f
C1327 a_n3827_n3924.t45 gnd 1.00187f
C1328 a_n3827_n3924.n10 gnd 0.340028f
C1329 a_n3827_n3924.t22 gnd 1.00187f
C1330 a_n3827_n3924.n11 gnd 0.340028f
C1331 a_n3827_n3924.t43 gnd 0.096397f
C1332 a_n3827_n3924.t27 gnd 0.096397f
C1333 a_n3827_n3924.n12 gnd 0.787293f
C1334 a_n3827_n3924.n13 gnd 0.319299f
C1335 a_n3827_n3924.t32 gnd 0.096397f
C1336 a_n3827_n3924.t20 gnd 0.096397f
C1337 a_n3827_n3924.n14 gnd 0.787293f
C1338 a_n3827_n3924.n15 gnd 0.319299f
C1339 a_n3827_n3924.t44 gnd 0.096397f
C1340 a_n3827_n3924.t7 gnd 0.096397f
C1341 a_n3827_n3924.n16 gnd 0.787293f
C1342 a_n3827_n3924.n17 gnd 0.319299f
C1343 a_n3827_n3924.t21 gnd 0.096397f
C1344 a_n3827_n3924.t33 gnd 0.096397f
C1345 a_n3827_n3924.n18 gnd 0.787293f
C1346 a_n3827_n3924.n19 gnd 0.319299f
C1347 a_n3827_n3924.t6 gnd 1.00187f
C1348 a_n3827_n3924.n20 gnd 0.864586f
C1349 a_n3827_n3924.t19 gnd 1.00187f
C1350 a_n3827_n3924.n21 gnd 0.549564f
C1351 a_n3827_n3924.t36 gnd 0.096397f
C1352 a_n3827_n3924.t49 gnd 0.096397f
C1353 a_n3827_n3924.n22 gnd 0.787292f
C1354 a_n3827_n3924.n23 gnd 0.319301f
C1355 a_n3827_n3924.t39 gnd 0.096397f
C1356 a_n3827_n3924.t35 gnd 0.096397f
C1357 a_n3827_n3924.n24 gnd 0.787292f
C1358 a_n3827_n3924.n25 gnd 0.319301f
C1359 a_n3827_n3924.t18 gnd 0.096397f
C1360 a_n3827_n3924.t0 gnd 0.096397f
C1361 a_n3827_n3924.n26 gnd 0.787292f
C1362 a_n3827_n3924.n27 gnd 0.319301f
C1363 a_n3827_n3924.t3 gnd 0.096397f
C1364 a_n3827_n3924.t40 gnd 0.096397f
C1365 a_n3827_n3924.n28 gnd 0.787292f
C1366 a_n3827_n3924.n29 gnd 0.319301f
C1367 a_n3827_n3924.t34 gnd 1.00187f
C1368 a_n3827_n3924.n30 gnd 0.340031f
C1369 a_n3827_n3924.t37 gnd 1.00187f
C1370 a_n3827_n3924.n31 gnd 0.340031f
C1371 a_n3827_n3924.t5 gnd 0.096397f
C1372 a_n3827_n3924.t1 gnd 0.096397f
C1373 a_n3827_n3924.n32 gnd 0.787292f
C1374 a_n3827_n3924.n33 gnd 0.319301f
C1375 a_n3827_n3924.t48 gnd 0.096397f
C1376 a_n3827_n3924.t23 gnd 0.096397f
C1377 a_n3827_n3924.n34 gnd 0.787292f
C1378 a_n3827_n3924.n35 gnd 0.319301f
C1379 a_n3827_n3924.t26 gnd 0.096397f
C1380 a_n3827_n3924.t30 gnd 0.096397f
C1381 a_n3827_n3924.n36 gnd 0.787292f
C1382 a_n3827_n3924.n37 gnd 0.319301f
C1383 a_n3827_n3924.t41 gnd 0.096397f
C1384 a_n3827_n3924.t24 gnd 0.096397f
C1385 a_n3827_n3924.n38 gnd 0.787292f
C1386 a_n3827_n3924.n39 gnd 0.319301f
C1387 a_n3827_n3924.t4 gnd 1.00187f
C1388 a_n3827_n3924.n40 gnd 0.549564f
C1389 a_n3827_n3924.n41 gnd 0.899874f
C1390 a_n3827_n3924.t10 gnd 1.24822f
C1391 a_n3827_n3924.t14 gnd 1.24481f
C1392 a_n3827_n3924.n42 gnd 1.83656f
C1393 a_n3827_n3924.n43 gnd 0.473862f
C1394 a_n3827_n3924.t9 gnd 1.24481f
C1395 a_n3827_n3924.n44 gnd 0.673252f
C1396 a_n3827_n3924.t12 gnd 1.24481f
C1397 a_n3827_n3924.n45 gnd 0.876738f
C1398 a_n3827_n3924.t8 gnd 1.24481f
C1399 a_n3827_n3924.n46 gnd 0.876738f
C1400 a_n3827_n3924.t13 gnd 1.24481f
C1401 a_n3827_n3924.n47 gnd 0.876738f
C1402 a_n3827_n3924.t16 gnd 1.24481f
C1403 a_n3827_n3924.n48 gnd 0.743593f
C1404 a_n3827_n3924.n49 gnd 0.473862f
C1405 a_n3827_n3924.t15 gnd 1.24481f
C1406 a_n3827_n3924.n50 gnd 0.678276f
C1407 a_n3827_n3924.t11 gnd 1.24481f
C1408 a_n3827_n3924.n51 gnd 1.44378f
C1409 a_n3827_n3924.t17 gnd 1.24658f
C1410 diffpairibias.t27 gnd 0.090128f
C1411 diffpairibias.t23 gnd 0.08996f
C1412 diffpairibias.n0 gnd 0.105991f
C1413 diffpairibias.t28 gnd 0.08996f
C1414 diffpairibias.n1 gnd 0.051736f
C1415 diffpairibias.t25 gnd 0.08996f
C1416 diffpairibias.n2 gnd 0.051736f
C1417 diffpairibias.t29 gnd 0.08996f
C1418 diffpairibias.n3 gnd 0.041084f
C1419 diffpairibias.t15 gnd 0.086371f
C1420 diffpairibias.t1 gnd 0.085993f
C1421 diffpairibias.n4 gnd 0.13579f
C1422 diffpairibias.t11 gnd 0.085993f
C1423 diffpairibias.n5 gnd 0.072463f
C1424 diffpairibias.t13 gnd 0.085993f
C1425 diffpairibias.n6 gnd 0.072463f
C1426 diffpairibias.t7 gnd 0.085993f
C1427 diffpairibias.n7 gnd 0.072463f
C1428 diffpairibias.t3 gnd 0.085993f
C1429 diffpairibias.n8 gnd 0.072463f
C1430 diffpairibias.t17 gnd 0.085993f
C1431 diffpairibias.n9 gnd 0.072463f
C1432 diffpairibias.t5 gnd 0.085993f
C1433 diffpairibias.n10 gnd 0.072463f
C1434 diffpairibias.t19 gnd 0.085993f
C1435 diffpairibias.n11 gnd 0.072463f
C1436 diffpairibias.t9 gnd 0.085993f
C1437 diffpairibias.n12 gnd 0.102883f
C1438 diffpairibias.t14 gnd 0.086899f
C1439 diffpairibias.t0 gnd 0.086748f
C1440 diffpairibias.n13 gnd 0.094648f
C1441 diffpairibias.t10 gnd 0.086748f
C1442 diffpairibias.n14 gnd 0.052262f
C1443 diffpairibias.t12 gnd 0.086748f
C1444 diffpairibias.n15 gnd 0.052262f
C1445 diffpairibias.t6 gnd 0.086748f
C1446 diffpairibias.n16 gnd 0.052262f
C1447 diffpairibias.t2 gnd 0.086748f
C1448 diffpairibias.n17 gnd 0.052262f
C1449 diffpairibias.t16 gnd 0.086748f
C1450 diffpairibias.n18 gnd 0.052262f
C1451 diffpairibias.t4 gnd 0.086748f
C1452 diffpairibias.n19 gnd 0.052262f
C1453 diffpairibias.t18 gnd 0.086748f
C1454 diffpairibias.n20 gnd 0.052262f
C1455 diffpairibias.t8 gnd 0.086748f
C1456 diffpairibias.n21 gnd 0.061849f
C1457 diffpairibias.n22 gnd 0.233513f
C1458 diffpairibias.t20 gnd 0.08996f
C1459 diffpairibias.n23 gnd 0.051747f
C1460 diffpairibias.t26 gnd 0.08996f
C1461 diffpairibias.n24 gnd 0.051736f
C1462 diffpairibias.t22 gnd 0.08996f
C1463 diffpairibias.n25 gnd 0.051736f
C1464 diffpairibias.t21 gnd 0.08996f
C1465 diffpairibias.n26 gnd 0.051736f
C1466 diffpairibias.t24 gnd 0.08996f
C1467 diffpairibias.n27 gnd 0.04729f
C1468 diffpairibias.n28 gnd 0.047711f
C1469 outputibias.t10 gnd 0.11477f
C1470 outputibias.t8 gnd 0.115567f
C1471 outputibias.n0 gnd 0.130108f
C1472 outputibias.n1 gnd 0.001372f
C1473 outputibias.n2 gnd 9.76e-19
C1474 outputibias.n3 gnd 5.24e-19
C1475 outputibias.n4 gnd 0.001239f
C1476 outputibias.n5 gnd 5.55e-19
C1477 outputibias.n6 gnd 9.76e-19
C1478 outputibias.n7 gnd 5.24e-19
C1479 outputibias.n8 gnd 0.001239f
C1480 outputibias.n9 gnd 5.55e-19
C1481 outputibias.n10 gnd 0.004176f
C1482 outputibias.t7 gnd 0.00202f
C1483 outputibias.n11 gnd 9.3e-19
C1484 outputibias.n12 gnd 7.32e-19
C1485 outputibias.n13 gnd 5.24e-19
C1486 outputibias.n14 gnd 0.02322f
C1487 outputibias.n15 gnd 9.76e-19
C1488 outputibias.n16 gnd 5.24e-19
C1489 outputibias.n17 gnd 5.55e-19
C1490 outputibias.n18 gnd 0.001239f
C1491 outputibias.n19 gnd 0.001239f
C1492 outputibias.n20 gnd 5.55e-19
C1493 outputibias.n21 gnd 5.24e-19
C1494 outputibias.n22 gnd 9.76e-19
C1495 outputibias.n23 gnd 9.76e-19
C1496 outputibias.n24 gnd 5.24e-19
C1497 outputibias.n25 gnd 5.55e-19
C1498 outputibias.n26 gnd 0.001239f
C1499 outputibias.n27 gnd 0.002683f
C1500 outputibias.n28 gnd 5.55e-19
C1501 outputibias.n29 gnd 5.24e-19
C1502 outputibias.n30 gnd 0.002256f
C1503 outputibias.n31 gnd 0.005781f
C1504 outputibias.n32 gnd 0.001372f
C1505 outputibias.n33 gnd 9.76e-19
C1506 outputibias.n34 gnd 5.24e-19
C1507 outputibias.n35 gnd 0.001239f
C1508 outputibias.n36 gnd 5.55e-19
C1509 outputibias.n37 gnd 9.76e-19
C1510 outputibias.n38 gnd 5.24e-19
C1511 outputibias.n39 gnd 0.001239f
C1512 outputibias.n40 gnd 5.55e-19
C1513 outputibias.n41 gnd 0.004176f
C1514 outputibias.t5 gnd 0.00202f
C1515 outputibias.n42 gnd 9.3e-19
C1516 outputibias.n43 gnd 7.32e-19
C1517 outputibias.n44 gnd 5.24e-19
C1518 outputibias.n45 gnd 0.02322f
C1519 outputibias.n46 gnd 9.76e-19
C1520 outputibias.n47 gnd 5.24e-19
C1521 outputibias.n48 gnd 5.55e-19
C1522 outputibias.n49 gnd 0.001239f
C1523 outputibias.n50 gnd 0.001239f
C1524 outputibias.n51 gnd 5.55e-19
C1525 outputibias.n52 gnd 5.24e-19
C1526 outputibias.n53 gnd 9.76e-19
C1527 outputibias.n54 gnd 9.76e-19
C1528 outputibias.n55 gnd 5.24e-19
C1529 outputibias.n56 gnd 5.55e-19
C1530 outputibias.n57 gnd 0.001239f
C1531 outputibias.n58 gnd 0.002683f
C1532 outputibias.n59 gnd 5.55e-19
C1533 outputibias.n60 gnd 5.24e-19
C1534 outputibias.n61 gnd 0.002256f
C1535 outputibias.n62 gnd 0.005197f
C1536 outputibias.n63 gnd 0.121892f
C1537 outputibias.n64 gnd 0.001372f
C1538 outputibias.n65 gnd 9.76e-19
C1539 outputibias.n66 gnd 5.24e-19
C1540 outputibias.n67 gnd 0.001239f
C1541 outputibias.n68 gnd 5.55e-19
C1542 outputibias.n69 gnd 9.76e-19
C1543 outputibias.n70 gnd 5.24e-19
C1544 outputibias.n71 gnd 0.001239f
C1545 outputibias.n72 gnd 5.55e-19
C1546 outputibias.n73 gnd 0.004176f
C1547 outputibias.t3 gnd 0.00202f
C1548 outputibias.n74 gnd 9.3e-19
C1549 outputibias.n75 gnd 7.32e-19
C1550 outputibias.n76 gnd 5.24e-19
C1551 outputibias.n77 gnd 0.02322f
C1552 outputibias.n78 gnd 9.76e-19
C1553 outputibias.n79 gnd 5.24e-19
C1554 outputibias.n80 gnd 5.55e-19
C1555 outputibias.n81 gnd 0.001239f
C1556 outputibias.n82 gnd 0.001239f
C1557 outputibias.n83 gnd 5.55e-19
C1558 outputibias.n84 gnd 5.24e-19
C1559 outputibias.n85 gnd 9.76e-19
C1560 outputibias.n86 gnd 9.76e-19
C1561 outputibias.n87 gnd 5.24e-19
C1562 outputibias.n88 gnd 5.55e-19
C1563 outputibias.n89 gnd 0.001239f
C1564 outputibias.n90 gnd 0.002683f
C1565 outputibias.n91 gnd 5.55e-19
C1566 outputibias.n92 gnd 5.24e-19
C1567 outputibias.n93 gnd 0.002256f
C1568 outputibias.n94 gnd 0.005197f
C1569 outputibias.n95 gnd 0.064513f
C1570 outputibias.n96 gnd 0.001372f
C1571 outputibias.n97 gnd 9.76e-19
C1572 outputibias.n98 gnd 5.24e-19
C1573 outputibias.n99 gnd 0.001239f
C1574 outputibias.n100 gnd 5.55e-19
C1575 outputibias.n101 gnd 9.76e-19
C1576 outputibias.n102 gnd 5.24e-19
C1577 outputibias.n103 gnd 0.001239f
C1578 outputibias.n104 gnd 5.55e-19
C1579 outputibias.n105 gnd 0.004176f
C1580 outputibias.t1 gnd 0.00202f
C1581 outputibias.n106 gnd 9.3e-19
C1582 outputibias.n107 gnd 7.32e-19
C1583 outputibias.n108 gnd 5.24e-19
C1584 outputibias.n109 gnd 0.02322f
C1585 outputibias.n110 gnd 9.76e-19
C1586 outputibias.n111 gnd 5.24e-19
C1587 outputibias.n112 gnd 5.55e-19
C1588 outputibias.n113 gnd 0.001239f
C1589 outputibias.n114 gnd 0.001239f
C1590 outputibias.n115 gnd 5.55e-19
C1591 outputibias.n116 gnd 5.24e-19
C1592 outputibias.n117 gnd 9.76e-19
C1593 outputibias.n118 gnd 9.76e-19
C1594 outputibias.n119 gnd 5.24e-19
C1595 outputibias.n120 gnd 5.55e-19
C1596 outputibias.n121 gnd 0.001239f
C1597 outputibias.n122 gnd 0.002683f
C1598 outputibias.n123 gnd 5.55e-19
C1599 outputibias.n124 gnd 5.24e-19
C1600 outputibias.n125 gnd 0.002256f
C1601 outputibias.n126 gnd 0.005197f
C1602 outputibias.n127 gnd 0.084814f
C1603 outputibias.t0 gnd 0.108319f
C1604 outputibias.t2 gnd 0.108319f
C1605 outputibias.t4 gnd 0.108319f
C1606 outputibias.t6 gnd 0.109238f
C1607 outputibias.n128 gnd 0.134674f
C1608 outputibias.n129 gnd 0.07244f
C1609 outputibias.n130 gnd 0.079818f
C1610 outputibias.n131 gnd 0.164901f
C1611 outputibias.t11 gnd 0.11477f
C1612 outputibias.n132 gnd 0.067481f
C1613 outputibias.t9 gnd 0.11477f
C1614 outputibias.n133 gnd 0.065115f
C1615 outputibias.n134 gnd 0.029159f
C1616 a_n2140_13878.t11 gnd 0.186452f
C1617 a_n2140_13878.t10 gnd 0.186452f
C1618 a_n2140_13878.t5 gnd 0.186452f
C1619 a_n2140_13878.n0 gnd 1.46971f
C1620 a_n2140_13878.t2 gnd 0.186452f
C1621 a_n2140_13878.t4 gnd 0.186452f
C1622 a_n2140_13878.n1 gnd 1.46815f
C1623 a_n2140_13878.n2 gnd 2.05145f
C1624 a_n2140_13878.t12 gnd 0.186452f
C1625 a_n2140_13878.t3 gnd 0.186452f
C1626 a_n2140_13878.n3 gnd 1.46815f
C1627 a_n2140_13878.n4 gnd 1.00065f
C1628 a_n2140_13878.t9 gnd 0.186452f
C1629 a_n2140_13878.t1 gnd 0.186452f
C1630 a_n2140_13878.n5 gnd 1.46815f
C1631 a_n2140_13878.n6 gnd 4.05307f
C1632 a_n2140_13878.t17 gnd 1.74584f
C1633 a_n2140_13878.t20 gnd 0.186452f
C1634 a_n2140_13878.t21 gnd 0.186452f
C1635 a_n2140_13878.n7 gnd 1.31337f
C1636 a_n2140_13878.n8 gnd 1.4675f
C1637 a_n2140_13878.t16 gnd 1.74237f
C1638 a_n2140_13878.n9 gnd 0.738464f
C1639 a_n2140_13878.t19 gnd 1.74237f
C1640 a_n2140_13878.n10 gnd 0.738464f
C1641 a_n2140_13878.t22 gnd 0.186452f
C1642 a_n2140_13878.t23 gnd 0.186452f
C1643 a_n2140_13878.n11 gnd 1.31337f
C1644 a_n2140_13878.n12 gnd 0.745616f
C1645 a_n2140_13878.t18 gnd 1.74237f
C1646 a_n2140_13878.n13 gnd 2.09116f
C1647 a_n2140_13878.n14 gnd 2.85337f
C1648 a_n2140_13878.t6 gnd 0.186452f
C1649 a_n2140_13878.t7 gnd 0.186452f
C1650 a_n2140_13878.n15 gnd 1.46815f
C1651 a_n2140_13878.n16 gnd 2.01216f
C1652 a_n2140_13878.t13 gnd 0.186452f
C1653 a_n2140_13878.t14 gnd 0.186452f
C1654 a_n2140_13878.n17 gnd 1.46815f
C1655 a_n2140_13878.n18 gnd 0.650499f
C1656 a_n2140_13878.t0 gnd 0.186452f
C1657 a_n2140_13878.t8 gnd 0.186452f
C1658 a_n2140_13878.n19 gnd 1.46815f
C1659 a_n2140_13878.n20 gnd 1.31969f
C1660 a_n2140_13878.n21 gnd 1.47058f
C1661 a_n2140_13878.t15 gnd 0.186452f
C1662 a_n2318_13878.n0 gnd 0.217886f
C1663 a_n2318_13878.n1 gnd 3.16141f
C1664 a_n2318_13878.n2 gnd 0.217886f
C1665 a_n2318_13878.n3 gnd 0.674574f
C1666 a_n2318_13878.n4 gnd 0.217886f
C1667 a_n2318_13878.n5 gnd 0.753716f
C1668 a_n2318_13878.n6 gnd 0.217886f
C1669 a_n2318_13878.n7 gnd 0.42604f
C1670 a_n2318_13878.n8 gnd 0.674551f
C1671 a_n2318_13878.n9 gnd 0.206738f
C1672 a_n2318_13878.n10 gnd 0.152266f
C1673 a_n2318_13878.n11 gnd 0.239314f
C1674 a_n2318_13878.n12 gnd 0.184843f
C1675 a_n2318_13878.n13 gnd 0.206738f
C1676 a_n2318_13878.n14 gnd 1.12829f
C1677 a_n2318_13878.n15 gnd 0.152266f
C1678 a_n2318_13878.n16 gnd 0.729022f
C1679 a_n2318_13878.n17 gnd 0.51701f
C1680 a_n2318_13878.n18 gnd 0.217886f
C1681 a_n2318_13878.n19 gnd 0.217886f
C1682 a_n2318_13878.n20 gnd 0.447806f
C1683 a_n2318_13878.n21 gnd 0.217886f
C1684 a_n2318_13878.n22 gnd 0.217886f
C1685 a_n2318_13878.n23 gnd 0.733554f
C1686 a_n2318_13878.n24 gnd 2.98994f
C1687 a_n2318_13878.n25 gnd 2.92523f
C1688 a_n2318_13878.n26 gnd 3.7969f
C1689 a_n2318_13878.n27 gnd 1.79383f
C1690 a_n2318_13878.n28 gnd 2.09784f
C1691 a_n2318_13878.n29 gnd 1.91464f
C1692 a_n2318_13878.n30 gnd 1.79383f
C1693 a_n2318_13878.n31 gnd 0.287827f
C1694 a_n2318_13878.n32 gnd 0.766802f
C1695 a_n2318_13878.n33 gnd 0.004897f
C1696 a_n2318_13878.n34 gnd 0.010591f
C1697 a_n2318_13878.n35 gnd 0.010591f
C1698 a_n2318_13878.n36 gnd 0.004897f
C1699 a_n2318_13878.n37 gnd 0.287827f
C1700 a_n2318_13878.n38 gnd 0.287827f
C1701 a_n2318_13878.n39 gnd 0.447806f
C1702 a_n2318_13878.n40 gnd 0.004897f
C1703 a_n2318_13878.n41 gnd 0.010591f
C1704 a_n2318_13878.n42 gnd 0.010591f
C1705 a_n2318_13878.n43 gnd 0.004897f
C1706 a_n2318_13878.n44 gnd 0.287827f
C1707 a_n2318_13878.n45 gnd 0.008436f
C1708 a_n2318_13878.n46 gnd 0.287827f
C1709 a_n2318_13878.n47 gnd 0.008436f
C1710 a_n2318_13878.n48 gnd 0.287827f
C1711 a_n2318_13878.n49 gnd 0.008436f
C1712 a_n2318_13878.n50 gnd 0.287827f
C1713 a_n2318_13878.n51 gnd 0.008436f
C1714 a_n2318_13878.n52 gnd 0.287827f
C1715 a_n2318_13878.n53 gnd 0.287827f
C1716 a_n2318_13878.n54 gnd 0.004897f
C1717 a_n2318_13878.n55 gnd 0.010591f
C1718 a_n2318_13878.n56 gnd 0.010591f
C1719 a_n2318_13878.n57 gnd 0.004897f
C1720 a_n2318_13878.n58 gnd 0.287827f
C1721 a_n2318_13878.n59 gnd 0.287827f
C1722 a_n2318_13878.n60 gnd 0.004897f
C1723 a_n2318_13878.n61 gnd 0.010591f
C1724 a_n2318_13878.n62 gnd 0.010591f
C1725 a_n2318_13878.n63 gnd 0.004897f
C1726 a_n2318_13878.n64 gnd 0.287827f
C1727 a_n2318_13878.t15 gnd 0.151128f
C1728 a_n2318_13878.t28 gnd 0.714753f
C1729 a_n2318_13878.t22 gnd 0.702974f
C1730 a_n2318_13878.t26 gnd 0.702974f
C1731 a_n2318_13878.n65 gnd 0.307084f
C1732 a_n2318_13878.t4 gnd 0.702974f
C1733 a_n2318_13878.t14 gnd 0.702974f
C1734 a_n2318_13878.t32 gnd 0.702974f
C1735 a_n2318_13878.n66 gnd 0.307084f
C1736 a_n2318_13878.t24 gnd 0.702974f
C1737 a_n2318_13878.t16 gnd 0.714753f
C1738 a_n2318_13878.t82 gnd 0.714753f
C1739 a_n2318_13878.t63 gnd 0.702974f
C1740 a_n2318_13878.t67 gnd 0.702974f
C1741 a_n2318_13878.n67 gnd 0.307084f
C1742 a_n2318_13878.t57 gnd 0.702974f
C1743 a_n2318_13878.t72 gnd 0.702974f
C1744 a_n2318_13878.t79 gnd 0.702974f
C1745 a_n2318_13878.n68 gnd 0.307084f
C1746 a_n2318_13878.t80 gnd 0.702974f
C1747 a_n2318_13878.t54 gnd 0.714753f
C1748 a_n2318_13878.t9 gnd 1.41509f
C1749 a_n2318_13878.t21 gnd 0.151128f
C1750 a_n2318_13878.t31 gnd 0.151128f
C1751 a_n2318_13878.n69 gnd 1.06455f
C1752 a_n2318_13878.t11 gnd 0.151128f
C1753 a_n2318_13878.t7 gnd 0.151128f
C1754 a_n2318_13878.n70 gnd 1.06455f
C1755 a_n2318_13878.t13 gnd 0.151128f
C1756 a_n2318_13878.t35 gnd 0.151128f
C1757 a_n2318_13878.n71 gnd 1.06455f
C1758 a_n2318_13878.t19 gnd 1.41226f
C1759 a_n2318_13878.t12 gnd 0.702974f
C1760 a_n2318_13878.n72 gnd 0.307084f
C1761 a_n2318_13878.t10 gnd 0.702974f
C1762 a_n2318_13878.t8 gnd 0.714753f
C1763 a_n2318_13878.t20 gnd 0.702974f
C1764 a_n2318_13878.t62 gnd 0.702974f
C1765 a_n2318_13878.n73 gnd 0.307084f
C1766 a_n2318_13878.t76 gnd 0.702974f
C1767 a_n2318_13878.t78 gnd 0.714753f
C1768 a_n2318_13878.t56 gnd 0.702974f
C1769 a_n2318_13878.n74 gnd 0.309588f
C1770 a_n2318_13878.t75 gnd 0.702974f
C1771 a_n2318_13878.n75 gnd 0.307084f
C1772 a_n2318_13878.n76 gnd 0.30246f
C1773 a_n2318_13878.t53 gnd 0.702974f
C1774 a_n2318_13878.n77 gnd 0.30246f
C1775 a_n2318_13878.t71 gnd 0.702974f
C1776 a_n2318_13878.n78 gnd 0.309588f
C1777 a_n2318_13878.t55 gnd 0.714753f
C1778 a_n2318_13878.n79 gnd 0.309588f
C1779 a_n2318_13878.t30 gnd 0.702974f
C1780 a_n2318_13878.n80 gnd 0.307084f
C1781 a_n2318_13878.n81 gnd 0.30246f
C1782 a_n2318_13878.t6 gnd 0.702974f
C1783 a_n2318_13878.n82 gnd 0.30246f
C1784 a_n2318_13878.t34 gnd 0.702974f
C1785 a_n2318_13878.n83 gnd 0.309588f
C1786 a_n2318_13878.t18 gnd 0.714753f
C1787 a_n2318_13878.n84 gnd 1.20932f
C1788 a_n2318_13878.t60 gnd 0.702974f
C1789 a_n2318_13878.n85 gnd 0.305147f
C1790 a_n2318_13878.t66 gnd 0.702974f
C1791 a_n2318_13878.n86 gnd 0.305147f
C1792 a_n2318_13878.t58 gnd 0.702974f
C1793 a_n2318_13878.n87 gnd 0.305147f
C1794 a_n2318_13878.t70 gnd 0.702974f
C1795 a_n2318_13878.n88 gnd 0.305147f
C1796 a_n2318_13878.t61 gnd 0.702974f
C1797 a_n2318_13878.n89 gnd 0.299606f
C1798 a_n2318_13878.t83 gnd 0.702974f
C1799 a_n2318_13878.n90 gnd 0.309072f
C1800 a_n2318_13878.t64 gnd 0.714753f
C1801 a_n2318_13878.t73 gnd 0.702974f
C1802 a_n2318_13878.n91 gnd 0.299606f
C1803 a_n2318_13878.t59 gnd 0.702974f
C1804 a_n2318_13878.n92 gnd 0.309072f
C1805 a_n2318_13878.t68 gnd 0.714753f
C1806 a_n2318_13878.t77 gnd 0.702974f
C1807 a_n2318_13878.n93 gnd 0.299606f
C1808 a_n2318_13878.t65 gnd 0.702974f
C1809 a_n2318_13878.n94 gnd 0.309072f
C1810 a_n2318_13878.t81 gnd 0.714753f
C1811 a_n2318_13878.t69 gnd 0.702974f
C1812 a_n2318_13878.n95 gnd 0.299606f
C1813 a_n2318_13878.t52 gnd 0.702974f
C1814 a_n2318_13878.n96 gnd 0.309072f
C1815 a_n2318_13878.t74 gnd 0.714753f
C1816 a_n2318_13878.n97 gnd 1.46328f
C1817 a_n2318_13878.n98 gnd 0.309588f
C1818 a_n2318_13878.n99 gnd 0.30246f
C1819 a_n2318_13878.n100 gnd 0.30246f
C1820 a_n2318_13878.n101 gnd 0.309588f
C1821 a_n2318_13878.t44 gnd 0.117544f
C1822 a_n2318_13878.t3 gnd 0.117544f
C1823 a_n2318_13878.n102 gnd 1.04031f
C1824 a_n2318_13878.t0 gnd 0.117544f
C1825 a_n2318_13878.t51 gnd 0.117544f
C1826 a_n2318_13878.n103 gnd 1.03866f
C1827 a_n2318_13878.t36 gnd 0.117544f
C1828 a_n2318_13878.t39 gnd 0.117544f
C1829 a_n2318_13878.n104 gnd 1.03866f
C1830 a_n2318_13878.t37 gnd 0.117544f
C1831 a_n2318_13878.t2 gnd 0.117544f
C1832 a_n2318_13878.n105 gnd 1.04031f
C1833 a_n2318_13878.t42 gnd 0.117544f
C1834 a_n2318_13878.t46 gnd 0.117544f
C1835 a_n2318_13878.n106 gnd 1.03866f
C1836 a_n2318_13878.t50 gnd 0.117544f
C1837 a_n2318_13878.t43 gnd 0.117544f
C1838 a_n2318_13878.n107 gnd 1.03866f
C1839 a_n2318_13878.t38 gnd 0.117544f
C1840 a_n2318_13878.t45 gnd 0.117544f
C1841 a_n2318_13878.n108 gnd 1.03866f
C1842 a_n2318_13878.t47 gnd 0.117544f
C1843 a_n2318_13878.t1 gnd 0.117544f
C1844 a_n2318_13878.n109 gnd 1.03866f
C1845 a_n2318_13878.t41 gnd 0.117544f
C1846 a_n2318_13878.t48 gnd 0.117544f
C1847 a_n2318_13878.n110 gnd 1.04032f
C1848 a_n2318_13878.t40 gnd 0.117544f
C1849 a_n2318_13878.t49 gnd 0.117544f
C1850 a_n2318_13878.n111 gnd 1.03866f
C1851 a_n2318_13878.n112 gnd 0.309588f
C1852 a_n2318_13878.n113 gnd 0.30246f
C1853 a_n2318_13878.n114 gnd 0.30246f
C1854 a_n2318_13878.n115 gnd 0.309588f
C1855 a_n2318_13878.n116 gnd 0.867362f
C1856 a_n2318_13878.t29 gnd 1.41227f
C1857 a_n2318_13878.t23 gnd 0.151128f
C1858 a_n2318_13878.t27 gnd 0.151128f
C1859 a_n2318_13878.n117 gnd 1.06455f
C1860 a_n2318_13878.t17 gnd 1.41509f
C1861 a_n2318_13878.t33 gnd 0.151128f
C1862 a_n2318_13878.t25 gnd 0.151128f
C1863 a_n2318_13878.n118 gnd 1.06455f
C1864 a_n2318_13878.n119 gnd 1.06455f
C1865 a_n2318_13878.t5 gnd 0.151128f
C1866 CSoutput.n0 gnd 0.044648f
C1867 CSoutput.t193 gnd 0.295337f
C1868 CSoutput.n1 gnd 0.13336f
C1869 CSoutput.n2 gnd 0.044648f
C1870 CSoutput.t176 gnd 0.295337f
C1871 CSoutput.n3 gnd 0.035387f
C1872 CSoutput.n4 gnd 0.044648f
C1873 CSoutput.t185 gnd 0.295337f
C1874 CSoutput.n5 gnd 0.030515f
C1875 CSoutput.n6 gnd 0.044648f
C1876 CSoutput.t196 gnd 0.295337f
C1877 CSoutput.t195 gnd 0.295337f
C1878 CSoutput.n7 gnd 0.131906f
C1879 CSoutput.n8 gnd 0.044648f
C1880 CSoutput.t182 gnd 0.295337f
C1881 CSoutput.n9 gnd 0.029094f
C1882 CSoutput.n10 gnd 0.044648f
C1883 CSoutput.t188 gnd 0.295337f
C1884 CSoutput.t191 gnd 0.295337f
C1885 CSoutput.n11 gnd 0.131906f
C1886 CSoutput.n12 gnd 0.044648f
C1887 CSoutput.t179 gnd 0.295337f
C1888 CSoutput.n13 gnd 0.030515f
C1889 CSoutput.n14 gnd 0.044648f
C1890 CSoutput.t178 gnd 0.295337f
C1891 CSoutput.t189 gnd 0.295337f
C1892 CSoutput.n15 gnd 0.131906f
C1893 CSoutput.n16 gnd 0.044648f
C1894 CSoutput.t194 gnd 0.295337f
C1895 CSoutput.n17 gnd 0.032591f
C1896 CSoutput.t180 gnd 0.352936f
C1897 CSoutput.t177 gnd 0.295337f
C1898 CSoutput.n18 gnd 0.168393f
C1899 CSoutput.n19 gnd 0.163399f
C1900 CSoutput.n20 gnd 0.189563f
C1901 CSoutput.n21 gnd 0.044648f
C1902 CSoutput.n22 gnd 0.037264f
C1903 CSoutput.n23 gnd 0.131906f
C1904 CSoutput.n24 gnd 0.035921f
C1905 CSoutput.n25 gnd 0.035387f
C1906 CSoutput.n26 gnd 0.044648f
C1907 CSoutput.n27 gnd 0.044648f
C1908 CSoutput.n28 gnd 0.036977f
C1909 CSoutput.n29 gnd 0.031395f
C1910 CSoutput.n30 gnd 0.134843f
C1911 CSoutput.n31 gnd 0.031827f
C1912 CSoutput.n32 gnd 0.044648f
C1913 CSoutput.n33 gnd 0.044648f
C1914 CSoutput.n34 gnd 0.044648f
C1915 CSoutput.n35 gnd 0.036583f
C1916 CSoutput.n36 gnd 0.131906f
C1917 CSoutput.n37 gnd 0.034987f
C1918 CSoutput.n38 gnd 0.036322f
C1919 CSoutput.n39 gnd 0.044648f
C1920 CSoutput.n40 gnd 0.044648f
C1921 CSoutput.n41 gnd 0.037256f
C1922 CSoutput.n42 gnd 0.034052f
C1923 CSoutput.n43 gnd 0.131906f
C1924 CSoutput.n44 gnd 0.034916f
C1925 CSoutput.n45 gnd 0.044648f
C1926 CSoutput.n46 gnd 0.044648f
C1927 CSoutput.n47 gnd 0.044648f
C1928 CSoutput.n48 gnd 0.034916f
C1929 CSoutput.n49 gnd 0.131906f
C1930 CSoutput.n50 gnd 0.034052f
C1931 CSoutput.n51 gnd 0.037256f
C1932 CSoutput.n52 gnd 0.044648f
C1933 CSoutput.n53 gnd 0.044648f
C1934 CSoutput.n54 gnd 0.036322f
C1935 CSoutput.n55 gnd 0.034987f
C1936 CSoutput.n56 gnd 0.131906f
C1937 CSoutput.n57 gnd 0.036583f
C1938 CSoutput.n58 gnd 0.044648f
C1939 CSoutput.n59 gnd 0.044648f
C1940 CSoutput.n60 gnd 0.044648f
C1941 CSoutput.n61 gnd 0.031827f
C1942 CSoutput.n62 gnd 0.134843f
C1943 CSoutput.n63 gnd 0.031395f
C1944 CSoutput.t197 gnd 0.295337f
C1945 CSoutput.n64 gnd 0.131906f
C1946 CSoutput.n65 gnd 0.036977f
C1947 CSoutput.n66 gnd 0.044648f
C1948 CSoutput.n67 gnd 0.044648f
C1949 CSoutput.n68 gnd 0.044648f
C1950 CSoutput.n69 gnd 0.035921f
C1951 CSoutput.n70 gnd 0.131906f
C1952 CSoutput.n71 gnd 0.037264f
C1953 CSoutput.n72 gnd 0.032591f
C1954 CSoutput.n73 gnd 0.044648f
C1955 CSoutput.n74 gnd 0.044648f
C1956 CSoutput.n75 gnd 0.033799f
C1957 CSoutput.n76 gnd 0.020073f
C1958 CSoutput.t183 gnd 0.331833f
C1959 CSoutput.n77 gnd 0.164841f
C1960 CSoutput.n78 gnd 0.70534f
C1961 CSoutput.t150 gnd 0.055692f
C1962 CSoutput.t97 gnd 0.055692f
C1963 CSoutput.n79 gnd 0.431188f
C1964 CSoutput.t162 gnd 0.055692f
C1965 CSoutput.t114 gnd 0.055692f
C1966 CSoutput.n80 gnd 0.430419f
C1967 CSoutput.n81 gnd 0.436874f
C1968 CSoutput.t78 gnd 0.055692f
C1969 CSoutput.t126 gnd 0.055692f
C1970 CSoutput.n82 gnd 0.430419f
C1971 CSoutput.n83 gnd 0.215273f
C1972 CSoutput.t82 gnd 0.055692f
C1973 CSoutput.t106 gnd 0.055692f
C1974 CSoutput.n84 gnd 0.430419f
C1975 CSoutput.n85 gnd 0.215273f
C1976 CSoutput.t166 gnd 0.055692f
C1977 CSoutput.t121 gnd 0.055692f
C1978 CSoutput.n86 gnd 0.430419f
C1979 CSoutput.n87 gnd 0.215273f
C1980 CSoutput.t85 gnd 0.055692f
C1981 CSoutput.t154 gnd 0.055692f
C1982 CSoutput.n88 gnd 0.430419f
C1983 CSoutput.n89 gnd 0.215273f
C1984 CSoutput.t93 gnd 0.055692f
C1985 CSoutput.t136 gnd 0.055692f
C1986 CSoutput.n90 gnd 0.430419f
C1987 CSoutput.n91 gnd 0.215273f
C1988 CSoutput.t109 gnd 0.055692f
C1989 CSoutput.t127 gnd 0.055692f
C1990 CSoutput.n92 gnd 0.430419f
C1991 CSoutput.n93 gnd 0.394762f
C1992 CSoutput.t74 gnd 0.055692f
C1993 CSoutput.t148 gnd 0.055692f
C1994 CSoutput.n94 gnd 0.431188f
C1995 CSoutput.t137 gnd 0.055692f
C1996 CSoutput.t116 gnd 0.055692f
C1997 CSoutput.n95 gnd 0.430419f
C1998 CSoutput.n96 gnd 0.436874f
C1999 CSoutput.t98 gnd 0.055692f
C2000 CSoutput.t159 gnd 0.055692f
C2001 CSoutput.n97 gnd 0.430419f
C2002 CSoutput.n98 gnd 0.215273f
C2003 CSoutput.t134 gnd 0.055692f
C2004 CSoutput.t133 gnd 0.055692f
C2005 CSoutput.n99 gnd 0.430419f
C2006 CSoutput.n100 gnd 0.215273f
C2007 CSoutput.t123 gnd 0.055692f
C2008 CSoutput.t94 gnd 0.055692f
C2009 CSoutput.n101 gnd 0.430419f
C2010 CSoutput.n102 gnd 0.215273f
C2011 CSoutput.t77 gnd 0.055692f
C2012 CSoutput.t124 gnd 0.055692f
C2013 CSoutput.n103 gnd 0.430419f
C2014 CSoutput.n104 gnd 0.215273f
C2015 CSoutput.t122 gnd 0.055692f
C2016 CSoutput.t92 gnd 0.055692f
C2017 CSoutput.n105 gnd 0.430419f
C2018 CSoutput.n106 gnd 0.215273f
C2019 CSoutput.t75 gnd 0.055692f
C2020 CSoutput.t73 gnd 0.055692f
C2021 CSoutput.n107 gnd 0.430419f
C2022 CSoutput.n108 gnd 0.321027f
C2023 CSoutput.n109 gnd 0.404813f
C2024 CSoutput.t87 gnd 0.055692f
C2025 CSoutput.t158 gnd 0.055692f
C2026 CSoutput.n110 gnd 0.431188f
C2027 CSoutput.t143 gnd 0.055692f
C2028 CSoutput.t125 gnd 0.055692f
C2029 CSoutput.n111 gnd 0.430419f
C2030 CSoutput.n112 gnd 0.436874f
C2031 CSoutput.t110 gnd 0.055692f
C2032 CSoutput.t167 gnd 0.055692f
C2033 CSoutput.n113 gnd 0.430419f
C2034 CSoutput.n114 gnd 0.215273f
C2035 CSoutput.t142 gnd 0.055692f
C2036 CSoutput.t141 gnd 0.055692f
C2037 CSoutput.n115 gnd 0.430419f
C2038 CSoutput.n116 gnd 0.215273f
C2039 CSoutput.t131 gnd 0.055692f
C2040 CSoutput.t107 gnd 0.055692f
C2041 CSoutput.n117 gnd 0.430419f
C2042 CSoutput.n118 gnd 0.215273f
C2043 CSoutput.t89 gnd 0.055692f
C2044 CSoutput.t132 gnd 0.055692f
C2045 CSoutput.n119 gnd 0.430419f
C2046 CSoutput.n120 gnd 0.215273f
C2047 CSoutput.t130 gnd 0.055692f
C2048 CSoutput.t105 gnd 0.055692f
C2049 CSoutput.n121 gnd 0.430419f
C2050 CSoutput.n122 gnd 0.215273f
C2051 CSoutput.t88 gnd 0.055692f
C2052 CSoutput.t86 gnd 0.055692f
C2053 CSoutput.n123 gnd 0.430419f
C2054 CSoutput.n124 gnd 0.321027f
C2055 CSoutput.n125 gnd 0.452477f
C2056 CSoutput.n126 gnd 9.424299f
C2057 CSoutput.n128 gnd 0.789817f
C2058 CSoutput.n129 gnd 0.592363f
C2059 CSoutput.n130 gnd 0.789817f
C2060 CSoutput.n131 gnd 0.789817f
C2061 CSoutput.n132 gnd 2.12643f
C2062 CSoutput.n133 gnd 0.789817f
C2063 CSoutput.n134 gnd 0.789817f
C2064 CSoutput.t187 gnd 0.987271f
C2065 CSoutput.n135 gnd 0.789817f
C2066 CSoutput.n136 gnd 0.789817f
C2067 CSoutput.n140 gnd 0.789817f
C2068 CSoutput.n144 gnd 0.789817f
C2069 CSoutput.n145 gnd 0.789817f
C2070 CSoutput.n147 gnd 0.789817f
C2071 CSoutput.n152 gnd 0.789817f
C2072 CSoutput.n154 gnd 0.789817f
C2073 CSoutput.n155 gnd 0.789817f
C2074 CSoutput.n157 gnd 0.789817f
C2075 CSoutput.n158 gnd 0.789817f
C2076 CSoutput.n160 gnd 0.789817f
C2077 CSoutput.t181 gnd 13.1978f
C2078 CSoutput.n162 gnd 0.789817f
C2079 CSoutput.n163 gnd 0.592363f
C2080 CSoutput.n164 gnd 0.789817f
C2081 CSoutput.n165 gnd 0.789817f
C2082 CSoutput.n166 gnd 2.12643f
C2083 CSoutput.n167 gnd 0.789817f
C2084 CSoutput.n168 gnd 0.789817f
C2085 CSoutput.t184 gnd 0.987271f
C2086 CSoutput.n169 gnd 0.789817f
C2087 CSoutput.n170 gnd 0.789817f
C2088 CSoutput.n174 gnd 0.789817f
C2089 CSoutput.n178 gnd 0.789817f
C2090 CSoutput.n179 gnd 0.789817f
C2091 CSoutput.n181 gnd 0.789817f
C2092 CSoutput.n186 gnd 0.789817f
C2093 CSoutput.n188 gnd 0.789817f
C2094 CSoutput.n189 gnd 0.789817f
C2095 CSoutput.n191 gnd 0.789817f
C2096 CSoutput.n192 gnd 0.789817f
C2097 CSoutput.n194 gnd 0.789817f
C2098 CSoutput.n195 gnd 0.592363f
C2099 CSoutput.n197 gnd 0.789817f
C2100 CSoutput.n198 gnd 0.592363f
C2101 CSoutput.n199 gnd 0.789817f
C2102 CSoutput.n200 gnd 0.789817f
C2103 CSoutput.n201 gnd 2.12643f
C2104 CSoutput.n202 gnd 0.789817f
C2105 CSoutput.n203 gnd 0.789817f
C2106 CSoutput.t186 gnd 0.987271f
C2107 CSoutput.n204 gnd 0.789817f
C2108 CSoutput.n205 gnd 2.12643f
C2109 CSoutput.n207 gnd 0.789817f
C2110 CSoutput.n208 gnd 0.789817f
C2111 CSoutput.n210 gnd 0.789817f
C2112 CSoutput.n211 gnd 0.789817f
C2113 CSoutput.t192 gnd 12.9827f
C2114 CSoutput.t190 gnd 13.1978f
C2115 CSoutput.n217 gnd 2.47777f
C2116 CSoutput.n218 gnd 10.0935f
C2117 CSoutput.n219 gnd 10.515901f
C2118 CSoutput.n224 gnd 2.68409f
C2119 CSoutput.n230 gnd 0.789817f
C2120 CSoutput.n232 gnd 0.789817f
C2121 CSoutput.n234 gnd 0.789817f
C2122 CSoutput.n236 gnd 0.789817f
C2123 CSoutput.n238 gnd 0.789817f
C2124 CSoutput.n244 gnd 0.789817f
C2125 CSoutput.n251 gnd 1.44901f
C2126 CSoutput.n252 gnd 1.44901f
C2127 CSoutput.n253 gnd 0.789817f
C2128 CSoutput.n254 gnd 0.789817f
C2129 CSoutput.n256 gnd 0.592363f
C2130 CSoutput.n257 gnd 0.507305f
C2131 CSoutput.n259 gnd 0.592363f
C2132 CSoutput.n260 gnd 0.507305f
C2133 CSoutput.n261 gnd 0.592363f
C2134 CSoutput.n263 gnd 0.789817f
C2135 CSoutput.n265 gnd 2.12643f
C2136 CSoutput.n266 gnd 2.47777f
C2137 CSoutput.n267 gnd 9.28346f
C2138 CSoutput.n269 gnd 0.592363f
C2139 CSoutput.n270 gnd 1.52419f
C2140 CSoutput.n271 gnd 0.592363f
C2141 CSoutput.n273 gnd 0.789817f
C2142 CSoutput.n275 gnd 2.12643f
C2143 CSoutput.n276 gnd 4.63171f
C2144 CSoutput.t96 gnd 0.055692f
C2145 CSoutput.t149 gnd 0.055692f
C2146 CSoutput.n277 gnd 0.431188f
C2147 CSoutput.t113 gnd 0.055692f
C2148 CSoutput.t161 gnd 0.055692f
C2149 CSoutput.n278 gnd 0.430419f
C2150 CSoutput.n279 gnd 0.436874f
C2151 CSoutput.t144 gnd 0.055692f
C2152 CSoutput.t76 gnd 0.055692f
C2153 CSoutput.n280 gnd 0.430419f
C2154 CSoutput.n281 gnd 0.215273f
C2155 CSoutput.t104 gnd 0.055692f
C2156 CSoutput.t81 gnd 0.055692f
C2157 CSoutput.n282 gnd 0.430419f
C2158 CSoutput.n283 gnd 0.215273f
C2159 CSoutput.t120 gnd 0.055692f
C2160 CSoutput.t101 gnd 0.055692f
C2161 CSoutput.n284 gnd 0.430419f
C2162 CSoutput.n285 gnd 0.215273f
C2163 CSoutput.t153 gnd 0.055692f
C2164 CSoutput.t84 gnd 0.055692f
C2165 CSoutput.n286 gnd 0.430419f
C2166 CSoutput.n287 gnd 0.215273f
C2167 CSoutput.t135 gnd 0.055692f
C2168 CSoutput.t90 gnd 0.055692f
C2169 CSoutput.n288 gnd 0.430419f
C2170 CSoutput.n289 gnd 0.215273f
C2171 CSoutput.t145 gnd 0.055692f
C2172 CSoutput.t108 gnd 0.055692f
C2173 CSoutput.n290 gnd 0.430419f
C2174 CSoutput.n291 gnd 0.394762f
C2175 CSoutput.t119 gnd 0.055692f
C2176 CSoutput.t139 gnd 0.055692f
C2177 CSoutput.n292 gnd 0.431188f
C2178 CSoutput.t72 gnd 0.055692f
C2179 CSoutput.t102 gnd 0.055692f
C2180 CSoutput.n293 gnd 0.430419f
C2181 CSoutput.n294 gnd 0.436874f
C2182 CSoutput.t103 gnd 0.055692f
C2183 CSoutput.t157 gnd 0.055692f
C2184 CSoutput.n295 gnd 0.430419f
C2185 CSoutput.n296 gnd 0.215273f
C2186 CSoutput.t99 gnd 0.055692f
C2187 CSoutput.t100 gnd 0.055692f
C2188 CSoutput.n297 gnd 0.430419f
C2189 CSoutput.n298 gnd 0.215273f
C2190 CSoutput.t155 gnd 0.055692f
C2191 CSoutput.t156 gnd 0.055692f
C2192 CSoutput.n299 gnd 0.430419f
C2193 CSoutput.n300 gnd 0.215273f
C2194 CSoutput.t80 gnd 0.055692f
C2195 CSoutput.t140 gnd 0.055692f
C2196 CSoutput.n301 gnd 0.430419f
C2197 CSoutput.n302 gnd 0.215273f
C2198 CSoutput.t152 gnd 0.055692f
C2199 CSoutput.t79 gnd 0.055692f
C2200 CSoutput.n303 gnd 0.430419f
C2201 CSoutput.n304 gnd 0.215273f
C2202 CSoutput.t118 gnd 0.055692f
C2203 CSoutput.t138 gnd 0.055692f
C2204 CSoutput.n305 gnd 0.430419f
C2205 CSoutput.n306 gnd 0.321027f
C2206 CSoutput.n307 gnd 0.404813f
C2207 CSoutput.t128 gnd 0.055692f
C2208 CSoutput.t146 gnd 0.055692f
C2209 CSoutput.n308 gnd 0.431188f
C2210 CSoutput.t83 gnd 0.055692f
C2211 CSoutput.t115 gnd 0.055692f
C2212 CSoutput.n309 gnd 0.430419f
C2213 CSoutput.n310 gnd 0.436874f
C2214 CSoutput.t117 gnd 0.055692f
C2215 CSoutput.t165 gnd 0.055692f
C2216 CSoutput.n311 gnd 0.430419f
C2217 CSoutput.n312 gnd 0.215273f
C2218 CSoutput.t111 gnd 0.055692f
C2219 CSoutput.t112 gnd 0.055692f
C2220 CSoutput.n313 gnd 0.430419f
C2221 CSoutput.n314 gnd 0.215273f
C2222 CSoutput.t163 gnd 0.055692f
C2223 CSoutput.t164 gnd 0.055692f
C2224 CSoutput.n315 gnd 0.430419f
C2225 CSoutput.n316 gnd 0.215273f
C2226 CSoutput.t95 gnd 0.055692f
C2227 CSoutput.t151 gnd 0.055692f
C2228 CSoutput.n317 gnd 0.430419f
C2229 CSoutput.n318 gnd 0.215273f
C2230 CSoutput.t160 gnd 0.055692f
C2231 CSoutput.t91 gnd 0.055692f
C2232 CSoutput.n319 gnd 0.430419f
C2233 CSoutput.n320 gnd 0.215273f
C2234 CSoutput.t129 gnd 0.055692f
C2235 CSoutput.t147 gnd 0.055692f
C2236 CSoutput.n321 gnd 0.430417f
C2237 CSoutput.n322 gnd 0.321028f
C2238 CSoutput.n323 gnd 0.452477f
C2239 CSoutput.n324 gnd 12.9707f
C2240 CSoutput.t7 gnd 0.048731f
C2241 CSoutput.t18 gnd 0.048731f
C2242 CSoutput.n325 gnd 0.432043f
C2243 CSoutput.t168 gnd 0.048731f
C2244 CSoutput.t41 gnd 0.048731f
C2245 CSoutput.n326 gnd 0.430601f
C2246 CSoutput.n327 gnd 0.40124f
C2247 CSoutput.t56 gnd 0.048731f
C2248 CSoutput.t61 gnd 0.048731f
C2249 CSoutput.n328 gnd 0.430601f
C2250 CSoutput.n329 gnd 0.197792f
C2251 CSoutput.t48 gnd 0.048731f
C2252 CSoutput.t174 gnd 0.048731f
C2253 CSoutput.n330 gnd 0.430601f
C2254 CSoutput.n331 gnd 0.197792f
C2255 CSoutput.t27 gnd 0.048731f
C2256 CSoutput.t71 gnd 0.048731f
C2257 CSoutput.n332 gnd 0.430601f
C2258 CSoutput.n333 gnd 0.197792f
C2259 CSoutput.t66 gnd 0.048731f
C2260 CSoutput.t173 gnd 0.048731f
C2261 CSoutput.n334 gnd 0.430601f
C2262 CSoutput.n335 gnd 0.197792f
C2263 CSoutput.t1 gnd 0.048731f
C2264 CSoutput.t21 gnd 0.048731f
C2265 CSoutput.n336 gnd 0.430601f
C2266 CSoutput.n337 gnd 0.197792f
C2267 CSoutput.t31 gnd 0.048731f
C2268 CSoutput.t34 gnd 0.048731f
C2269 CSoutput.n338 gnd 0.430601f
C2270 CSoutput.n339 gnd 0.197792f
C2271 CSoutput.t39 gnd 0.048731f
C2272 CSoutput.t50 gnd 0.048731f
C2273 CSoutput.n340 gnd 0.430601f
C2274 CSoutput.n341 gnd 0.197792f
C2275 CSoutput.t49 gnd 0.048731f
C2276 CSoutput.t20 gnd 0.048731f
C2277 CSoutput.n342 gnd 0.430601f
C2278 CSoutput.n343 gnd 0.364769f
C2279 CSoutput.t42 gnd 0.048731f
C2280 CSoutput.t13 gnd 0.048731f
C2281 CSoutput.n344 gnd 0.432043f
C2282 CSoutput.t11 gnd 0.048731f
C2283 CSoutput.t171 gnd 0.048731f
C2284 CSoutput.n345 gnd 0.430601f
C2285 CSoutput.n346 gnd 0.40124f
C2286 CSoutput.t4 gnd 0.048731f
C2287 CSoutput.t38 gnd 0.048731f
C2288 CSoutput.n347 gnd 0.430601f
C2289 CSoutput.n348 gnd 0.197792f
C2290 CSoutput.t68 gnd 0.048731f
C2291 CSoutput.t55 gnd 0.048731f
C2292 CSoutput.n349 gnd 0.430601f
C2293 CSoutput.n350 gnd 0.197792f
C2294 CSoutput.t12 gnd 0.048731f
C2295 CSoutput.t26 gnd 0.048731f
C2296 CSoutput.n351 gnd 0.430601f
C2297 CSoutput.n352 gnd 0.197792f
C2298 CSoutput.t63 gnd 0.048731f
C2299 CSoutput.t3 gnd 0.048731f
C2300 CSoutput.n353 gnd 0.430601f
C2301 CSoutput.n354 gnd 0.197792f
C2302 CSoutput.t16 gnd 0.048731f
C2303 CSoutput.t2 gnd 0.048731f
C2304 CSoutput.n355 gnd 0.430601f
C2305 CSoutput.n356 gnd 0.197792f
C2306 CSoutput.t175 gnd 0.048731f
C2307 CSoutput.t172 gnd 0.048731f
C2308 CSoutput.n357 gnd 0.430601f
C2309 CSoutput.n358 gnd 0.197792f
C2310 CSoutput.t14 gnd 0.048731f
C2311 CSoutput.t30 gnd 0.048731f
C2312 CSoutput.n359 gnd 0.430601f
C2313 CSoutput.n360 gnd 0.197792f
C2314 CSoutput.t69 gnd 0.048731f
C2315 CSoutput.t43 gnd 0.048731f
C2316 CSoutput.n361 gnd 0.430601f
C2317 CSoutput.n362 gnd 0.300291f
C2318 CSoutput.n363 gnd 0.557964f
C2319 CSoutput.n364 gnd 13.862901f
C2320 CSoutput.t70 gnd 0.048731f
C2321 CSoutput.t10 gnd 0.048731f
C2322 CSoutput.n365 gnd 0.432043f
C2323 CSoutput.t35 gnd 0.048731f
C2324 CSoutput.t45 gnd 0.048731f
C2325 CSoutput.n366 gnd 0.430601f
C2326 CSoutput.n367 gnd 0.40124f
C2327 CSoutput.t51 gnd 0.048731f
C2328 CSoutput.t44 gnd 0.048731f
C2329 CSoutput.n368 gnd 0.430601f
C2330 CSoutput.n369 gnd 0.197792f
C2331 CSoutput.t32 gnd 0.048731f
C2332 CSoutput.t67 gnd 0.048731f
C2333 CSoutput.n370 gnd 0.430601f
C2334 CSoutput.n371 gnd 0.197792f
C2335 CSoutput.t46 gnd 0.048731f
C2336 CSoutput.t8 gnd 0.048731f
C2337 CSoutput.n372 gnd 0.430601f
C2338 CSoutput.n373 gnd 0.197792f
C2339 CSoutput.t47 gnd 0.048731f
C2340 CSoutput.t54 gnd 0.048731f
C2341 CSoutput.n374 gnd 0.430601f
C2342 CSoutput.n375 gnd 0.197792f
C2343 CSoutput.t59 gnd 0.048731f
C2344 CSoutput.t24 gnd 0.048731f
C2345 CSoutput.n376 gnd 0.430601f
C2346 CSoutput.n377 gnd 0.197792f
C2347 CSoutput.t6 gnd 0.048731f
C2348 CSoutput.t40 gnd 0.048731f
C2349 CSoutput.n378 gnd 0.430601f
C2350 CSoutput.n379 gnd 0.197792f
C2351 CSoutput.t9 gnd 0.048731f
C2352 CSoutput.t28 gnd 0.048731f
C2353 CSoutput.n380 gnd 0.430601f
C2354 CSoutput.n381 gnd 0.197792f
C2355 CSoutput.t0 gnd 0.048731f
C2356 CSoutput.t17 gnd 0.048731f
C2357 CSoutput.n382 gnd 0.430601f
C2358 CSoutput.n383 gnd 0.364769f
C2359 CSoutput.t62 gnd 0.048731f
C2360 CSoutput.t22 gnd 0.048731f
C2361 CSoutput.n384 gnd 0.432043f
C2362 CSoutput.t15 gnd 0.048731f
C2363 CSoutput.t23 gnd 0.048731f
C2364 CSoutput.n385 gnd 0.430601f
C2365 CSoutput.n386 gnd 0.40124f
C2366 CSoutput.t5 gnd 0.048731f
C2367 CSoutput.t37 gnd 0.048731f
C2368 CSoutput.n387 gnd 0.430601f
C2369 CSoutput.n388 gnd 0.197792f
C2370 CSoutput.t58 gnd 0.048731f
C2371 CSoutput.t52 gnd 0.048731f
C2372 CSoutput.n389 gnd 0.430601f
C2373 CSoutput.n390 gnd 0.197792f
C2374 CSoutput.t60 gnd 0.048731f
C2375 CSoutput.t25 gnd 0.048731f
C2376 CSoutput.n391 gnd 0.430601f
C2377 CSoutput.n392 gnd 0.197792f
C2378 CSoutput.t29 gnd 0.048731f
C2379 CSoutput.t169 gnd 0.048731f
C2380 CSoutput.n393 gnd 0.430601f
C2381 CSoutput.n394 gnd 0.197792f
C2382 CSoutput.t53 gnd 0.048731f
C2383 CSoutput.t170 gnd 0.048731f
C2384 CSoutput.n395 gnd 0.430601f
C2385 CSoutput.n396 gnd 0.197792f
C2386 CSoutput.t57 gnd 0.048731f
C2387 CSoutput.t65 gnd 0.048731f
C2388 CSoutput.n397 gnd 0.430601f
C2389 CSoutput.n398 gnd 0.197792f
C2390 CSoutput.t36 gnd 0.048731f
C2391 CSoutput.t19 gnd 0.048731f
C2392 CSoutput.n399 gnd 0.430601f
C2393 CSoutput.n400 gnd 0.197792f
C2394 CSoutput.t33 gnd 0.048731f
C2395 CSoutput.t64 gnd 0.048731f
C2396 CSoutput.n401 gnd 0.430601f
C2397 CSoutput.n402 gnd 0.300291f
C2398 CSoutput.n403 gnd 0.557964f
C2399 CSoutput.n404 gnd 8.431059f
C2400 CSoutput.n405 gnd 14.554401f
C2401 vdd.t25 gnd 0.037051f
C2402 vdd.t127 gnd 0.037051f
C2403 vdd.n0 gnd 0.29223f
C2404 vdd.t3 gnd 0.037051f
C2405 vdd.t38 gnd 0.037051f
C2406 vdd.n1 gnd 0.291748f
C2407 vdd.n2 gnd 0.269047f
C2408 vdd.t47 gnd 0.037051f
C2409 vdd.t6 gnd 0.037051f
C2410 vdd.n3 gnd 0.291748f
C2411 vdd.n4 gnd 0.136067f
C2412 vdd.t267 gnd 0.037051f
C2413 vdd.t27 gnd 0.037051f
C2414 vdd.n5 gnd 0.291748f
C2415 vdd.n6 gnd 0.127674f
C2416 vdd.t21 gnd 0.037051f
C2417 vdd.t49 gnd 0.037051f
C2418 vdd.n7 gnd 0.29223f
C2419 vdd.t13 gnd 0.037051f
C2420 vdd.t35 gnd 0.037051f
C2421 vdd.n8 gnd 0.291748f
C2422 vdd.n9 gnd 0.269047f
C2423 vdd.t32 gnd 0.037051f
C2424 vdd.t30 gnd 0.037051f
C2425 vdd.n10 gnd 0.291748f
C2426 vdd.n11 gnd 0.136067f
C2427 vdd.t15 gnd 0.037051f
C2428 vdd.t18 gnd 0.037051f
C2429 vdd.n12 gnd 0.291748f
C2430 vdd.n13 gnd 0.127674f
C2431 vdd.n14 gnd 0.090263f
C2432 vdd.t130 gnd 0.020584f
C2433 vdd.t43 gnd 0.020584f
C2434 vdd.n15 gnd 0.189468f
C2435 vdd.t134 gnd 0.020584f
C2436 vdd.t39 gnd 0.020584f
C2437 vdd.n16 gnd 0.188913f
C2438 vdd.n17 gnd 0.328768f
C2439 vdd.t133 gnd 0.020584f
C2440 vdd.t44 gnd 0.020584f
C2441 vdd.n18 gnd 0.188913f
C2442 vdd.n19 gnd 0.136016f
C2443 vdd.t135 gnd 0.020584f
C2444 vdd.t40 gnd 0.020584f
C2445 vdd.n20 gnd 0.189468f
C2446 vdd.t131 gnd 0.020584f
C2447 vdd.t128 gnd 0.020584f
C2448 vdd.n21 gnd 0.188913f
C2449 vdd.n22 gnd 0.328768f
C2450 vdd.t41 gnd 0.020584f
C2451 vdd.t42 gnd 0.020584f
C2452 vdd.n23 gnd 0.188913f
C2453 vdd.n24 gnd 0.136016f
C2454 vdd.t129 gnd 0.020584f
C2455 vdd.t137 gnd 0.020584f
C2456 vdd.n25 gnd 0.188913f
C2457 vdd.t136 gnd 0.020584f
C2458 vdd.t132 gnd 0.020584f
C2459 vdd.n26 gnd 0.188913f
C2460 vdd.n27 gnd 22.1869f
C2461 vdd.n28 gnd 8.48422f
C2462 vdd.n29 gnd 0.005614f
C2463 vdd.n30 gnd 0.00521f
C2464 vdd.n31 gnd 0.002882f
C2465 vdd.n32 gnd 0.006617f
C2466 vdd.n33 gnd 0.002799f
C2467 vdd.n34 gnd 0.002964f
C2468 vdd.n35 gnd 0.00521f
C2469 vdd.n36 gnd 0.002799f
C2470 vdd.n37 gnd 0.006617f
C2471 vdd.n38 gnd 0.002964f
C2472 vdd.n39 gnd 0.00521f
C2473 vdd.n40 gnd 0.002799f
C2474 vdd.n41 gnd 0.004963f
C2475 vdd.n42 gnd 0.004977f
C2476 vdd.t178 gnd 0.014216f
C2477 vdd.n43 gnd 0.03163f
C2478 vdd.n44 gnd 0.164609f
C2479 vdd.n45 gnd 0.002799f
C2480 vdd.n46 gnd 0.002964f
C2481 vdd.n47 gnd 0.006617f
C2482 vdd.n48 gnd 0.006617f
C2483 vdd.n49 gnd 0.002964f
C2484 vdd.n50 gnd 0.002799f
C2485 vdd.n51 gnd 0.00521f
C2486 vdd.n52 gnd 0.00521f
C2487 vdd.n53 gnd 0.002799f
C2488 vdd.n54 gnd 0.002964f
C2489 vdd.n55 gnd 0.006617f
C2490 vdd.n56 gnd 0.006617f
C2491 vdd.n57 gnd 0.002964f
C2492 vdd.n58 gnd 0.002799f
C2493 vdd.n59 gnd 0.00521f
C2494 vdd.n60 gnd 0.00521f
C2495 vdd.n61 gnd 0.002799f
C2496 vdd.n62 gnd 0.002964f
C2497 vdd.n63 gnd 0.006617f
C2498 vdd.n64 gnd 0.006617f
C2499 vdd.n65 gnd 0.015644f
C2500 vdd.n66 gnd 0.002882f
C2501 vdd.n67 gnd 0.002799f
C2502 vdd.n68 gnd 0.013465f
C2503 vdd.n69 gnd 0.009401f
C2504 vdd.t247 gnd 0.032935f
C2505 vdd.t202 gnd 0.032935f
C2506 vdd.n70 gnd 0.226349f
C2507 vdd.n71 gnd 0.177989f
C2508 vdd.t259 gnd 0.032935f
C2509 vdd.t242 gnd 0.032935f
C2510 vdd.n72 gnd 0.226349f
C2511 vdd.n73 gnd 0.143636f
C2512 vdd.t147 gnd 0.032935f
C2513 vdd.t193 gnd 0.032935f
C2514 vdd.n74 gnd 0.226349f
C2515 vdd.n75 gnd 0.143636f
C2516 vdd.t157 gnd 0.032935f
C2517 vdd.t212 gnd 0.032935f
C2518 vdd.n76 gnd 0.226349f
C2519 vdd.n77 gnd 0.143636f
C2520 vdd.t183 gnd 0.032935f
C2521 vdd.t251 gnd 0.032935f
C2522 vdd.n78 gnd 0.226349f
C2523 vdd.n79 gnd 0.143636f
C2524 vdd.t162 gnd 0.032935f
C2525 vdd.t231 gnd 0.032935f
C2526 vdd.n80 gnd 0.226349f
C2527 vdd.n81 gnd 0.143636f
C2528 vdd.t168 gnd 0.032935f
C2529 vdd.t243 gnd 0.032935f
C2530 vdd.n82 gnd 0.226349f
C2531 vdd.n83 gnd 0.143636f
C2532 vdd.n84 gnd 0.005614f
C2533 vdd.n85 gnd 0.00521f
C2534 vdd.n86 gnd 0.002882f
C2535 vdd.n87 gnd 0.006617f
C2536 vdd.n88 gnd 0.002799f
C2537 vdd.n89 gnd 0.002964f
C2538 vdd.n90 gnd 0.00521f
C2539 vdd.n91 gnd 0.002799f
C2540 vdd.n92 gnd 0.006617f
C2541 vdd.n93 gnd 0.002964f
C2542 vdd.n94 gnd 0.00521f
C2543 vdd.n95 gnd 0.002799f
C2544 vdd.n96 gnd 0.004963f
C2545 vdd.n97 gnd 0.004977f
C2546 vdd.t197 gnd 0.014216f
C2547 vdd.n98 gnd 0.03163f
C2548 vdd.n99 gnd 0.164609f
C2549 vdd.n100 gnd 0.002799f
C2550 vdd.n101 gnd 0.002964f
C2551 vdd.n102 gnd 0.006617f
C2552 vdd.n103 gnd 0.006617f
C2553 vdd.n104 gnd 0.002964f
C2554 vdd.n105 gnd 0.002799f
C2555 vdd.n106 gnd 0.00521f
C2556 vdd.n107 gnd 0.00521f
C2557 vdd.n108 gnd 0.002799f
C2558 vdd.n109 gnd 0.002964f
C2559 vdd.n110 gnd 0.006617f
C2560 vdd.n111 gnd 0.006617f
C2561 vdd.n112 gnd 0.002964f
C2562 vdd.n113 gnd 0.002799f
C2563 vdd.n114 gnd 0.00521f
C2564 vdd.n115 gnd 0.00521f
C2565 vdd.n116 gnd 0.002799f
C2566 vdd.n117 gnd 0.002964f
C2567 vdd.n118 gnd 0.006617f
C2568 vdd.n119 gnd 0.006617f
C2569 vdd.n120 gnd 0.015644f
C2570 vdd.n121 gnd 0.002882f
C2571 vdd.n122 gnd 0.002799f
C2572 vdd.n123 gnd 0.013465f
C2573 vdd.n124 gnd 0.009106f
C2574 vdd.n125 gnd 0.106866f
C2575 vdd.n126 gnd 0.005614f
C2576 vdd.n127 gnd 0.00521f
C2577 vdd.n128 gnd 0.002882f
C2578 vdd.n129 gnd 0.006617f
C2579 vdd.n130 gnd 0.002799f
C2580 vdd.n131 gnd 0.002964f
C2581 vdd.n132 gnd 0.00521f
C2582 vdd.n133 gnd 0.002799f
C2583 vdd.n134 gnd 0.006617f
C2584 vdd.n135 gnd 0.002964f
C2585 vdd.n136 gnd 0.00521f
C2586 vdd.n137 gnd 0.002799f
C2587 vdd.n138 gnd 0.004963f
C2588 vdd.n139 gnd 0.004977f
C2589 vdd.t210 gnd 0.014216f
C2590 vdd.n140 gnd 0.03163f
C2591 vdd.n141 gnd 0.164609f
C2592 vdd.n142 gnd 0.002799f
C2593 vdd.n143 gnd 0.002964f
C2594 vdd.n144 gnd 0.006617f
C2595 vdd.n145 gnd 0.006617f
C2596 vdd.n146 gnd 0.002964f
C2597 vdd.n147 gnd 0.002799f
C2598 vdd.n148 gnd 0.00521f
C2599 vdd.n149 gnd 0.00521f
C2600 vdd.n150 gnd 0.002799f
C2601 vdd.n151 gnd 0.002964f
C2602 vdd.n152 gnd 0.006617f
C2603 vdd.n153 gnd 0.006617f
C2604 vdd.n154 gnd 0.002964f
C2605 vdd.n155 gnd 0.002799f
C2606 vdd.n156 gnd 0.00521f
C2607 vdd.n157 gnd 0.00521f
C2608 vdd.n158 gnd 0.002799f
C2609 vdd.n159 gnd 0.002964f
C2610 vdd.n160 gnd 0.006617f
C2611 vdd.n161 gnd 0.006617f
C2612 vdd.n162 gnd 0.015644f
C2613 vdd.n163 gnd 0.002882f
C2614 vdd.n164 gnd 0.002799f
C2615 vdd.n165 gnd 0.013465f
C2616 vdd.n166 gnd 0.009401f
C2617 vdd.t237 gnd 0.032935f
C2618 vdd.t139 gnd 0.032935f
C2619 vdd.n167 gnd 0.226349f
C2620 vdd.n168 gnd 0.177989f
C2621 vdd.t188 gnd 0.032935f
C2622 vdd.t190 gnd 0.032935f
C2623 vdd.n169 gnd 0.226349f
C2624 vdd.n170 gnd 0.143636f
C2625 vdd.t255 gnd 0.032935f
C2626 vdd.t185 gnd 0.032935f
C2627 vdd.n171 gnd 0.226349f
C2628 vdd.n172 gnd 0.143636f
C2629 vdd.t186 gnd 0.032935f
C2630 vdd.t253 gnd 0.032935f
C2631 vdd.n173 gnd 0.226349f
C2632 vdd.n174 gnd 0.143636f
C2633 vdd.t254 gnd 0.032935f
C2634 vdd.t155 gnd 0.032935f
C2635 vdd.n175 gnd 0.226349f
C2636 vdd.n176 gnd 0.143636f
C2637 vdd.t238 gnd 0.032935f
C2638 vdd.t250 gnd 0.032935f
C2639 vdd.n177 gnd 0.226349f
C2640 vdd.n178 gnd 0.143636f
C2641 vdd.t153 gnd 0.032935f
C2642 vdd.t207 gnd 0.032935f
C2643 vdd.n179 gnd 0.226349f
C2644 vdd.n180 gnd 0.143636f
C2645 vdd.n181 gnd 0.005614f
C2646 vdd.n182 gnd 0.00521f
C2647 vdd.n183 gnd 0.002882f
C2648 vdd.n184 gnd 0.006617f
C2649 vdd.n185 gnd 0.002799f
C2650 vdd.n186 gnd 0.002964f
C2651 vdd.n187 gnd 0.00521f
C2652 vdd.n188 gnd 0.002799f
C2653 vdd.n189 gnd 0.006617f
C2654 vdd.n190 gnd 0.002964f
C2655 vdd.n191 gnd 0.00521f
C2656 vdd.n192 gnd 0.002799f
C2657 vdd.n193 gnd 0.004963f
C2658 vdd.n194 gnd 0.004977f
C2659 vdd.t235 gnd 0.014216f
C2660 vdd.n195 gnd 0.03163f
C2661 vdd.n196 gnd 0.164609f
C2662 vdd.n197 gnd 0.002799f
C2663 vdd.n198 gnd 0.002964f
C2664 vdd.n199 gnd 0.006617f
C2665 vdd.n200 gnd 0.006617f
C2666 vdd.n201 gnd 0.002964f
C2667 vdd.n202 gnd 0.002799f
C2668 vdd.n203 gnd 0.00521f
C2669 vdd.n204 gnd 0.00521f
C2670 vdd.n205 gnd 0.002799f
C2671 vdd.n206 gnd 0.002964f
C2672 vdd.n207 gnd 0.006617f
C2673 vdd.n208 gnd 0.006617f
C2674 vdd.n209 gnd 0.002964f
C2675 vdd.n210 gnd 0.002799f
C2676 vdd.n211 gnd 0.00521f
C2677 vdd.n212 gnd 0.00521f
C2678 vdd.n213 gnd 0.002799f
C2679 vdd.n214 gnd 0.002964f
C2680 vdd.n215 gnd 0.006617f
C2681 vdd.n216 gnd 0.006617f
C2682 vdd.n217 gnd 0.015644f
C2683 vdd.n218 gnd 0.002882f
C2684 vdd.n219 gnd 0.002799f
C2685 vdd.n220 gnd 0.013465f
C2686 vdd.n221 gnd 0.009106f
C2687 vdd.n222 gnd 0.063574f
C2688 vdd.n223 gnd 0.229075f
C2689 vdd.n224 gnd 0.005614f
C2690 vdd.n225 gnd 0.00521f
C2691 vdd.n226 gnd 0.002882f
C2692 vdd.n227 gnd 0.006617f
C2693 vdd.n228 gnd 0.002799f
C2694 vdd.n229 gnd 0.002964f
C2695 vdd.n230 gnd 0.00521f
C2696 vdd.n231 gnd 0.002799f
C2697 vdd.n232 gnd 0.006617f
C2698 vdd.n233 gnd 0.002964f
C2699 vdd.n234 gnd 0.00521f
C2700 vdd.n235 gnd 0.002799f
C2701 vdd.n236 gnd 0.004963f
C2702 vdd.n237 gnd 0.004977f
C2703 vdd.t223 gnd 0.014216f
C2704 vdd.n238 gnd 0.03163f
C2705 vdd.n239 gnd 0.164609f
C2706 vdd.n240 gnd 0.002799f
C2707 vdd.n241 gnd 0.002964f
C2708 vdd.n242 gnd 0.006617f
C2709 vdd.n243 gnd 0.006617f
C2710 vdd.n244 gnd 0.002964f
C2711 vdd.n245 gnd 0.002799f
C2712 vdd.n246 gnd 0.00521f
C2713 vdd.n247 gnd 0.00521f
C2714 vdd.n248 gnd 0.002799f
C2715 vdd.n249 gnd 0.002964f
C2716 vdd.n250 gnd 0.006617f
C2717 vdd.n251 gnd 0.006617f
C2718 vdd.n252 gnd 0.002964f
C2719 vdd.n253 gnd 0.002799f
C2720 vdd.n254 gnd 0.00521f
C2721 vdd.n255 gnd 0.00521f
C2722 vdd.n256 gnd 0.002799f
C2723 vdd.n257 gnd 0.002964f
C2724 vdd.n258 gnd 0.006617f
C2725 vdd.n259 gnd 0.006617f
C2726 vdd.n260 gnd 0.015644f
C2727 vdd.n261 gnd 0.002882f
C2728 vdd.n262 gnd 0.002799f
C2729 vdd.n263 gnd 0.013465f
C2730 vdd.n264 gnd 0.009401f
C2731 vdd.t244 gnd 0.032935f
C2732 vdd.t160 gnd 0.032935f
C2733 vdd.n265 gnd 0.226349f
C2734 vdd.n266 gnd 0.177989f
C2735 vdd.t205 gnd 0.032935f
C2736 vdd.t209 gnd 0.032935f
C2737 vdd.n267 gnd 0.226349f
C2738 vdd.n268 gnd 0.143636f
C2739 vdd.t263 gnd 0.032935f
C2740 vdd.t200 gnd 0.032935f
C2741 vdd.n269 gnd 0.226349f
C2742 vdd.n270 gnd 0.143636f
C2743 vdd.t201 gnd 0.032935f
C2744 vdd.t261 gnd 0.032935f
C2745 vdd.n271 gnd 0.226349f
C2746 vdd.n272 gnd 0.143636f
C2747 vdd.t262 gnd 0.032935f
C2748 vdd.t176 gnd 0.032935f
C2749 vdd.n273 gnd 0.226349f
C2750 vdd.n274 gnd 0.143636f
C2751 vdd.t249 gnd 0.032935f
C2752 vdd.t258 gnd 0.032935f
C2753 vdd.n275 gnd 0.226349f
C2754 vdd.n276 gnd 0.143636f
C2755 vdd.t169 gnd 0.032935f
C2756 vdd.t224 gnd 0.032935f
C2757 vdd.n277 gnd 0.226349f
C2758 vdd.n278 gnd 0.143636f
C2759 vdd.n279 gnd 0.005614f
C2760 vdd.n280 gnd 0.00521f
C2761 vdd.n281 gnd 0.002882f
C2762 vdd.n282 gnd 0.006617f
C2763 vdd.n283 gnd 0.002799f
C2764 vdd.n284 gnd 0.002964f
C2765 vdd.n285 gnd 0.00521f
C2766 vdd.n286 gnd 0.002799f
C2767 vdd.n287 gnd 0.006617f
C2768 vdd.n288 gnd 0.002964f
C2769 vdd.n289 gnd 0.00521f
C2770 vdd.n290 gnd 0.002799f
C2771 vdd.n291 gnd 0.004963f
C2772 vdd.n292 gnd 0.004977f
C2773 vdd.t245 gnd 0.014216f
C2774 vdd.n293 gnd 0.03163f
C2775 vdd.n294 gnd 0.164609f
C2776 vdd.n295 gnd 0.002799f
C2777 vdd.n296 gnd 0.002964f
C2778 vdd.n297 gnd 0.006617f
C2779 vdd.n298 gnd 0.006617f
C2780 vdd.n299 gnd 0.002964f
C2781 vdd.n300 gnd 0.002799f
C2782 vdd.n301 gnd 0.00521f
C2783 vdd.n302 gnd 0.00521f
C2784 vdd.n303 gnd 0.002799f
C2785 vdd.n304 gnd 0.002964f
C2786 vdd.n305 gnd 0.006617f
C2787 vdd.n306 gnd 0.006617f
C2788 vdd.n307 gnd 0.002964f
C2789 vdd.n308 gnd 0.002799f
C2790 vdd.n309 gnd 0.00521f
C2791 vdd.n310 gnd 0.00521f
C2792 vdd.n311 gnd 0.002799f
C2793 vdd.n312 gnd 0.002964f
C2794 vdd.n313 gnd 0.006617f
C2795 vdd.n314 gnd 0.006617f
C2796 vdd.n315 gnd 0.015644f
C2797 vdd.n316 gnd 0.002882f
C2798 vdd.n317 gnd 0.002799f
C2799 vdd.n318 gnd 0.013465f
C2800 vdd.n319 gnd 0.009106f
C2801 vdd.n320 gnd 0.063574f
C2802 vdd.n321 gnd 0.256534f
C2803 vdd.n322 gnd 0.007862f
C2804 vdd.n323 gnd 0.01023f
C2805 vdd.n324 gnd 0.008234f
C2806 vdd.n325 gnd 0.008234f
C2807 vdd.n326 gnd 0.01023f
C2808 vdd.n327 gnd 0.01023f
C2809 vdd.n328 gnd 0.747477f
C2810 vdd.n329 gnd 0.01023f
C2811 vdd.n330 gnd 0.01023f
C2812 vdd.n331 gnd 0.01023f
C2813 vdd.n332 gnd 0.810202f
C2814 vdd.n333 gnd 0.01023f
C2815 vdd.n334 gnd 0.01023f
C2816 vdd.n335 gnd 0.01023f
C2817 vdd.n336 gnd 0.01023f
C2818 vdd.n337 gnd 0.008234f
C2819 vdd.n338 gnd 0.01023f
C2820 vdd.t154 gnd 0.522711f
C2821 vdd.n339 gnd 0.01023f
C2822 vdd.n340 gnd 0.01023f
C2823 vdd.n341 gnd 0.01023f
C2824 vdd.t230 gnd 0.522711f
C2825 vdd.n342 gnd 0.01023f
C2826 vdd.n343 gnd 0.01023f
C2827 vdd.n344 gnd 0.01023f
C2828 vdd.n345 gnd 0.01023f
C2829 vdd.n346 gnd 0.01023f
C2830 vdd.n347 gnd 0.008234f
C2831 vdd.n348 gnd 0.01023f
C2832 vdd.n349 gnd 0.590664f
C2833 vdd.n350 gnd 0.01023f
C2834 vdd.n351 gnd 0.01023f
C2835 vdd.n352 gnd 0.01023f
C2836 vdd.t206 gnd 0.522711f
C2837 vdd.n353 gnd 0.01023f
C2838 vdd.n354 gnd 0.01023f
C2839 vdd.n355 gnd 0.01023f
C2840 vdd.n356 gnd 0.01023f
C2841 vdd.n357 gnd 0.01023f
C2842 vdd.n358 gnd 0.008234f
C2843 vdd.n359 gnd 0.01023f
C2844 vdd.t196 gnd 0.522711f
C2845 vdd.n360 gnd 0.01023f
C2846 vdd.n361 gnd 0.01023f
C2847 vdd.n362 gnd 0.01023f
C2848 vdd.n363 gnd 0.883382f
C2849 vdd.n364 gnd 0.01023f
C2850 vdd.n365 gnd 0.01023f
C2851 vdd.n366 gnd 0.01023f
C2852 vdd.n367 gnd 0.01023f
C2853 vdd.n368 gnd 0.01023f
C2854 vdd.n369 gnd 0.006834f
C2855 vdd.n370 gnd 0.023295f
C2856 vdd.t84 gnd 0.522711f
C2857 vdd.n371 gnd 0.01023f
C2858 vdd.n372 gnd 0.023295f
C2859 vdd.n404 gnd 0.01023f
C2860 vdd.t86 gnd 0.125851f
C2861 vdd.t85 gnd 0.134501f
C2862 vdd.t83 gnd 0.164361f
C2863 vdd.n405 gnd 0.210687f
C2864 vdd.n406 gnd 0.177839f
C2865 vdd.n407 gnd 0.013503f
C2866 vdd.n408 gnd 0.01023f
C2867 vdd.n409 gnd 0.008234f
C2868 vdd.n410 gnd 0.01023f
C2869 vdd.n411 gnd 0.008234f
C2870 vdd.n412 gnd 0.01023f
C2871 vdd.n413 gnd 0.008234f
C2872 vdd.n414 gnd 0.01023f
C2873 vdd.n415 gnd 0.008234f
C2874 vdd.n416 gnd 0.01023f
C2875 vdd.n417 gnd 0.008234f
C2876 vdd.n418 gnd 0.01023f
C2877 vdd.t119 gnd 0.125851f
C2878 vdd.t118 gnd 0.134501f
C2879 vdd.t117 gnd 0.164361f
C2880 vdd.n419 gnd 0.210687f
C2881 vdd.n420 gnd 0.177839f
C2882 vdd.n421 gnd 0.008234f
C2883 vdd.n422 gnd 0.01023f
C2884 vdd.n423 gnd 0.008234f
C2885 vdd.n424 gnd 0.01023f
C2886 vdd.n425 gnd 0.008234f
C2887 vdd.n426 gnd 0.01023f
C2888 vdd.n427 gnd 0.008234f
C2889 vdd.n428 gnd 0.01023f
C2890 vdd.n429 gnd 0.008234f
C2891 vdd.n430 gnd 0.01023f
C2892 vdd.t125 gnd 0.125851f
C2893 vdd.t124 gnd 0.134501f
C2894 vdd.t123 gnd 0.164361f
C2895 vdd.n431 gnd 0.210687f
C2896 vdd.n432 gnd 0.177839f
C2897 vdd.n433 gnd 0.01762f
C2898 vdd.n434 gnd 0.01023f
C2899 vdd.n435 gnd 0.008234f
C2900 vdd.n436 gnd 0.01023f
C2901 vdd.n437 gnd 0.008234f
C2902 vdd.n438 gnd 0.01023f
C2903 vdd.n439 gnd 0.008234f
C2904 vdd.n440 gnd 0.01023f
C2905 vdd.n441 gnd 0.008234f
C2906 vdd.n442 gnd 0.01023f
C2907 vdd.n443 gnd 0.023295f
C2908 vdd.n444 gnd 0.023454f
C2909 vdd.n445 gnd 0.023454f
C2910 vdd.n446 gnd 0.006834f
C2911 vdd.n447 gnd 0.008234f
C2912 vdd.n448 gnd 0.01023f
C2913 vdd.n449 gnd 0.01023f
C2914 vdd.n450 gnd 0.008234f
C2915 vdd.n451 gnd 0.01023f
C2916 vdd.n452 gnd 0.01023f
C2917 vdd.n453 gnd 0.01023f
C2918 vdd.n454 gnd 0.01023f
C2919 vdd.n455 gnd 0.01023f
C2920 vdd.n456 gnd 0.008234f
C2921 vdd.n457 gnd 0.008234f
C2922 vdd.n458 gnd 0.01023f
C2923 vdd.n459 gnd 0.01023f
C2924 vdd.n460 gnd 0.008234f
C2925 vdd.n461 gnd 0.01023f
C2926 vdd.n462 gnd 0.01023f
C2927 vdd.n463 gnd 0.01023f
C2928 vdd.n464 gnd 0.01023f
C2929 vdd.n465 gnd 0.01023f
C2930 vdd.n466 gnd 0.008234f
C2931 vdd.n467 gnd 0.008234f
C2932 vdd.n468 gnd 0.01023f
C2933 vdd.n469 gnd 0.01023f
C2934 vdd.n470 gnd 0.008234f
C2935 vdd.n471 gnd 0.01023f
C2936 vdd.n472 gnd 0.01023f
C2937 vdd.n473 gnd 0.01023f
C2938 vdd.n474 gnd 0.01023f
C2939 vdd.n475 gnd 0.01023f
C2940 vdd.n476 gnd 0.008234f
C2941 vdd.n477 gnd 0.008234f
C2942 vdd.n478 gnd 0.01023f
C2943 vdd.n479 gnd 0.01023f
C2944 vdd.n480 gnd 0.008234f
C2945 vdd.n481 gnd 0.01023f
C2946 vdd.n482 gnd 0.01023f
C2947 vdd.n483 gnd 0.01023f
C2948 vdd.n484 gnd 0.01023f
C2949 vdd.n485 gnd 0.01023f
C2950 vdd.n486 gnd 0.008234f
C2951 vdd.n487 gnd 0.008234f
C2952 vdd.n488 gnd 0.01023f
C2953 vdd.n489 gnd 0.01023f
C2954 vdd.n490 gnd 0.006875f
C2955 vdd.n491 gnd 0.01023f
C2956 vdd.n492 gnd 0.01023f
C2957 vdd.n493 gnd 0.01023f
C2958 vdd.n494 gnd 0.01023f
C2959 vdd.n495 gnd 0.01023f
C2960 vdd.n496 gnd 0.006875f
C2961 vdd.n497 gnd 0.008234f
C2962 vdd.n498 gnd 0.01023f
C2963 vdd.n499 gnd 0.01023f
C2964 vdd.n500 gnd 0.008234f
C2965 vdd.n501 gnd 0.01023f
C2966 vdd.n502 gnd 0.01023f
C2967 vdd.n503 gnd 0.01023f
C2968 vdd.n504 gnd 0.01023f
C2969 vdd.n505 gnd 0.01023f
C2970 vdd.n506 gnd 0.008234f
C2971 vdd.n507 gnd 0.008234f
C2972 vdd.n508 gnd 0.01023f
C2973 vdd.n509 gnd 0.01023f
C2974 vdd.n510 gnd 0.008234f
C2975 vdd.n511 gnd 0.01023f
C2976 vdd.n512 gnd 0.01023f
C2977 vdd.n513 gnd 0.01023f
C2978 vdd.n514 gnd 0.01023f
C2979 vdd.n515 gnd 0.01023f
C2980 vdd.n516 gnd 0.008234f
C2981 vdd.n517 gnd 0.008234f
C2982 vdd.n518 gnd 0.01023f
C2983 vdd.n519 gnd 0.01023f
C2984 vdd.n520 gnd 0.008234f
C2985 vdd.n521 gnd 0.01023f
C2986 vdd.n522 gnd 0.01023f
C2987 vdd.n523 gnd 0.01023f
C2988 vdd.n524 gnd 0.01023f
C2989 vdd.n525 gnd 0.01023f
C2990 vdd.n526 gnd 0.008234f
C2991 vdd.n527 gnd 0.008234f
C2992 vdd.n528 gnd 0.01023f
C2993 vdd.n529 gnd 0.01023f
C2994 vdd.n530 gnd 0.008234f
C2995 vdd.n531 gnd 0.01023f
C2996 vdd.n532 gnd 0.01023f
C2997 vdd.n533 gnd 0.01023f
C2998 vdd.n534 gnd 0.01023f
C2999 vdd.n535 gnd 0.01023f
C3000 vdd.n536 gnd 0.008234f
C3001 vdd.n537 gnd 0.008234f
C3002 vdd.n538 gnd 0.01023f
C3003 vdd.n539 gnd 0.01023f
C3004 vdd.n540 gnd 0.008234f
C3005 vdd.n541 gnd 0.01023f
C3006 vdd.n542 gnd 0.01023f
C3007 vdd.n543 gnd 0.01023f
C3008 vdd.n544 gnd 0.01023f
C3009 vdd.n545 gnd 0.01023f
C3010 vdd.n546 gnd 0.005599f
C3011 vdd.n547 gnd 0.01762f
C3012 vdd.n548 gnd 0.01023f
C3013 vdd.n549 gnd 0.01023f
C3014 vdd.n550 gnd 0.008151f
C3015 vdd.n551 gnd 0.01023f
C3016 vdd.n552 gnd 0.01023f
C3017 vdd.n553 gnd 0.01023f
C3018 vdd.n554 gnd 0.01023f
C3019 vdd.n555 gnd 0.01023f
C3020 vdd.n556 gnd 0.008234f
C3021 vdd.n557 gnd 0.008234f
C3022 vdd.n558 gnd 0.01023f
C3023 vdd.n559 gnd 0.01023f
C3024 vdd.n560 gnd 0.008234f
C3025 vdd.n561 gnd 0.01023f
C3026 vdd.n562 gnd 0.01023f
C3027 vdd.n563 gnd 0.01023f
C3028 vdd.n564 gnd 0.01023f
C3029 vdd.n565 gnd 0.01023f
C3030 vdd.n566 gnd 0.008234f
C3031 vdd.n567 gnd 0.008234f
C3032 vdd.n568 gnd 0.01023f
C3033 vdd.n569 gnd 0.01023f
C3034 vdd.n570 gnd 0.008234f
C3035 vdd.n571 gnd 0.01023f
C3036 vdd.n572 gnd 0.01023f
C3037 vdd.n573 gnd 0.01023f
C3038 vdd.n574 gnd 0.01023f
C3039 vdd.n575 gnd 0.01023f
C3040 vdd.n576 gnd 0.008234f
C3041 vdd.n577 gnd 0.008234f
C3042 vdd.n578 gnd 0.01023f
C3043 vdd.n579 gnd 0.01023f
C3044 vdd.n580 gnd 0.008234f
C3045 vdd.n581 gnd 0.01023f
C3046 vdd.n582 gnd 0.01023f
C3047 vdd.n583 gnd 0.01023f
C3048 vdd.n584 gnd 0.01023f
C3049 vdd.n585 gnd 0.01023f
C3050 vdd.n586 gnd 0.008234f
C3051 vdd.n587 gnd 0.008234f
C3052 vdd.n588 gnd 0.01023f
C3053 vdd.n589 gnd 0.01023f
C3054 vdd.n590 gnd 0.008234f
C3055 vdd.n591 gnd 0.01023f
C3056 vdd.n592 gnd 0.01023f
C3057 vdd.n593 gnd 0.01023f
C3058 vdd.n594 gnd 0.01023f
C3059 vdd.n595 gnd 0.01023f
C3060 vdd.n596 gnd 0.008234f
C3061 vdd.n597 gnd 0.01023f
C3062 vdd.n598 gnd 0.008234f
C3063 vdd.n599 gnd 0.004323f
C3064 vdd.n600 gnd 0.01023f
C3065 vdd.n601 gnd 0.01023f
C3066 vdd.n602 gnd 0.008234f
C3067 vdd.n603 gnd 0.01023f
C3068 vdd.n604 gnd 0.008234f
C3069 vdd.n605 gnd 0.01023f
C3070 vdd.n606 gnd 0.008234f
C3071 vdd.n607 gnd 0.01023f
C3072 vdd.n608 gnd 0.008234f
C3073 vdd.n609 gnd 0.01023f
C3074 vdd.n610 gnd 0.008234f
C3075 vdd.n611 gnd 0.01023f
C3076 vdd.n612 gnd 0.01023f
C3077 vdd.n613 gnd 0.569755f
C3078 vdd.t156 gnd 0.522711f
C3079 vdd.n614 gnd 0.01023f
C3080 vdd.n615 gnd 0.008234f
C3081 vdd.n616 gnd 0.01023f
C3082 vdd.n617 gnd 0.008234f
C3083 vdd.n618 gnd 0.01023f
C3084 vdd.t146 gnd 0.522711f
C3085 vdd.n619 gnd 0.01023f
C3086 vdd.n620 gnd 0.008234f
C3087 vdd.n621 gnd 0.01023f
C3088 vdd.n622 gnd 0.008234f
C3089 vdd.n623 gnd 0.01023f
C3090 vdd.t189 gnd 0.522711f
C3091 vdd.n624 gnd 0.653389f
C3092 vdd.n625 gnd 0.01023f
C3093 vdd.n626 gnd 0.008234f
C3094 vdd.n627 gnd 0.01023f
C3095 vdd.n628 gnd 0.008234f
C3096 vdd.n629 gnd 0.01023f
C3097 vdd.t187 gnd 0.522711f
C3098 vdd.n630 gnd 0.01023f
C3099 vdd.n631 gnd 0.008234f
C3100 vdd.n632 gnd 0.01023f
C3101 vdd.n633 gnd 0.008234f
C3102 vdd.n634 gnd 0.01023f
C3103 vdd.n635 gnd 0.726568f
C3104 vdd.n636 gnd 0.8677f
C3105 vdd.t138 gnd 0.522711f
C3106 vdd.n637 gnd 0.01023f
C3107 vdd.n638 gnd 0.008234f
C3108 vdd.n639 gnd 0.01023f
C3109 vdd.n640 gnd 0.008234f
C3110 vdd.n641 gnd 0.01023f
C3111 vdd.n642 gnd 0.548847f
C3112 vdd.n643 gnd 0.01023f
C3113 vdd.n644 gnd 0.008234f
C3114 vdd.n645 gnd 0.01023f
C3115 vdd.n646 gnd 0.008234f
C3116 vdd.n647 gnd 0.01023f
C3117 vdd.n648 gnd 1.04542f
C3118 vdd.t177 gnd 0.522711f
C3119 vdd.n649 gnd 0.01023f
C3120 vdd.n650 gnd 0.008234f
C3121 vdd.n651 gnd 0.01023f
C3122 vdd.n652 gnd 0.008234f
C3123 vdd.n653 gnd 0.01023f
C3124 vdd.t59 gnd 0.522711f
C3125 vdd.n654 gnd 0.01023f
C3126 vdd.n655 gnd 0.008234f
C3127 vdd.n656 gnd 0.023454f
C3128 vdd.n657 gnd 0.023454f
C3129 vdd.n658 gnd 9.12654f
C3130 vdd.n659 gnd 0.580209f
C3131 vdd.n660 gnd 0.023454f
C3132 vdd.n661 gnd 0.008798f
C3133 vdd.n662 gnd 0.008234f
C3134 vdd.n667 gnd 0.006547f
C3135 vdd.n668 gnd 0.008234f
C3136 vdd.n669 gnd 0.01023f
C3137 vdd.n670 gnd 0.01023f
C3138 vdd.n671 gnd 0.01023f
C3139 vdd.n672 gnd 0.01023f
C3140 vdd.n673 gnd 0.01023f
C3141 vdd.n674 gnd 0.008234f
C3142 vdd.n675 gnd 0.01023f
C3143 vdd.n676 gnd 0.01023f
C3144 vdd.n677 gnd 0.01023f
C3145 vdd.n678 gnd 0.01023f
C3146 vdd.n679 gnd 0.01023f
C3147 vdd.n680 gnd 0.008234f
C3148 vdd.n681 gnd 0.01023f
C3149 vdd.n682 gnd 0.01023f
C3150 vdd.n683 gnd 0.01023f
C3151 vdd.n684 gnd 0.01023f
C3152 vdd.n685 gnd 0.01023f
C3153 vdd.t77 gnd 0.125851f
C3154 vdd.t78 gnd 0.134501f
C3155 vdd.t76 gnd 0.164361f
C3156 vdd.n686 gnd 0.210687f
C3157 vdd.n687 gnd 0.177015f
C3158 vdd.n688 gnd 0.016797f
C3159 vdd.n689 gnd 0.01023f
C3160 vdd.n690 gnd 0.01023f
C3161 vdd.n691 gnd 0.01023f
C3162 vdd.n692 gnd 0.01023f
C3163 vdd.n693 gnd 0.01023f
C3164 vdd.n694 gnd 0.008234f
C3165 vdd.n695 gnd 0.01023f
C3166 vdd.n696 gnd 0.01023f
C3167 vdd.n697 gnd 0.01023f
C3168 vdd.n698 gnd 0.01023f
C3169 vdd.n699 gnd 0.01023f
C3170 vdd.n700 gnd 0.008234f
C3171 vdd.n701 gnd 0.01023f
C3172 vdd.n702 gnd 0.01023f
C3173 vdd.n703 gnd 0.01023f
C3174 vdd.n704 gnd 0.01023f
C3175 vdd.n705 gnd 0.01023f
C3176 vdd.n706 gnd 0.008234f
C3177 vdd.n707 gnd 0.01023f
C3178 vdd.n708 gnd 0.01023f
C3179 vdd.n709 gnd 0.01023f
C3180 vdd.n710 gnd 0.01023f
C3181 vdd.n711 gnd 0.01023f
C3182 vdd.n712 gnd 0.008234f
C3183 vdd.n713 gnd 0.01023f
C3184 vdd.n714 gnd 0.01023f
C3185 vdd.n715 gnd 0.01023f
C3186 vdd.n716 gnd 0.01023f
C3187 vdd.n717 gnd 0.01023f
C3188 vdd.n718 gnd 0.008234f
C3189 vdd.n719 gnd 0.01023f
C3190 vdd.n720 gnd 0.01023f
C3191 vdd.n721 gnd 0.01023f
C3192 vdd.n722 gnd 0.008151f
C3193 vdd.t67 gnd 0.125851f
C3194 vdd.t68 gnd 0.134501f
C3195 vdd.t66 gnd 0.164361f
C3196 vdd.n723 gnd 0.210687f
C3197 vdd.n724 gnd 0.177015f
C3198 vdd.n725 gnd 0.01023f
C3199 vdd.n726 gnd 0.008234f
C3200 vdd.n728 gnd 0.01023f
C3201 vdd.n730 gnd 0.01023f
C3202 vdd.n731 gnd 0.01023f
C3203 vdd.n732 gnd 0.008234f
C3204 vdd.n733 gnd 0.01023f
C3205 vdd.n734 gnd 0.01023f
C3206 vdd.n735 gnd 0.01023f
C3207 vdd.n736 gnd 0.01023f
C3208 vdd.n737 gnd 0.01023f
C3209 vdd.n738 gnd 0.008234f
C3210 vdd.n739 gnd 0.01023f
C3211 vdd.n740 gnd 0.01023f
C3212 vdd.n741 gnd 0.01023f
C3213 vdd.n742 gnd 0.01023f
C3214 vdd.n743 gnd 0.01023f
C3215 vdd.n744 gnd 0.008234f
C3216 vdd.n745 gnd 0.01023f
C3217 vdd.n746 gnd 0.01023f
C3218 vdd.n747 gnd 0.01023f
C3219 vdd.n748 gnd 0.006547f
C3220 vdd.n753 gnd 0.006956f
C3221 vdd.n754 gnd 0.006956f
C3222 vdd.n755 gnd 0.006956f
C3223 vdd.n756 gnd 8.91745f
C3224 vdd.n757 gnd 0.006956f
C3225 vdd.n758 gnd 0.006956f
C3226 vdd.n759 gnd 0.006956f
C3227 vdd.n761 gnd 0.006956f
C3228 vdd.n762 gnd 0.006956f
C3229 vdd.n764 gnd 0.006956f
C3230 vdd.n765 gnd 0.005064f
C3231 vdd.n767 gnd 0.006956f
C3232 vdd.t53 gnd 0.281098f
C3233 vdd.t52 gnd 0.287738f
C3234 vdd.t50 gnd 0.183511f
C3235 vdd.n768 gnd 0.099178f
C3236 vdd.n769 gnd 0.056257f
C3237 vdd.n770 gnd 0.009941f
C3238 vdd.n771 gnd 0.016101f
C3239 vdd.n773 gnd 0.006956f
C3240 vdd.n774 gnd 0.710887f
C3241 vdd.n775 gnd 0.015237f
C3242 vdd.n776 gnd 0.015237f
C3243 vdd.n777 gnd 0.006956f
C3244 vdd.n778 gnd 0.01627f
C3245 vdd.n779 gnd 0.006956f
C3246 vdd.n780 gnd 0.006956f
C3247 vdd.n781 gnd 0.006956f
C3248 vdd.n782 gnd 0.006956f
C3249 vdd.n783 gnd 0.006956f
C3250 vdd.n785 gnd 0.006956f
C3251 vdd.n786 gnd 0.006956f
C3252 vdd.n788 gnd 0.006956f
C3253 vdd.n789 gnd 0.006956f
C3254 vdd.n791 gnd 0.006956f
C3255 vdd.n792 gnd 0.006956f
C3256 vdd.n794 gnd 0.006956f
C3257 vdd.n795 gnd 0.006956f
C3258 vdd.n797 gnd 0.006956f
C3259 vdd.n798 gnd 0.006956f
C3260 vdd.n800 gnd 0.006956f
C3261 vdd.n801 gnd 0.005064f
C3262 vdd.n803 gnd 0.006956f
C3263 vdd.t122 gnd 0.281098f
C3264 vdd.t121 gnd 0.287738f
C3265 vdd.t120 gnd 0.183511f
C3266 vdd.n804 gnd 0.099178f
C3267 vdd.n805 gnd 0.056257f
C3268 vdd.n806 gnd 0.009941f
C3269 vdd.n807 gnd 0.006956f
C3270 vdd.n808 gnd 0.006956f
C3271 vdd.t51 gnd 0.355444f
C3272 vdd.n809 gnd 0.006956f
C3273 vdd.n810 gnd 0.006956f
C3274 vdd.n811 gnd 0.006956f
C3275 vdd.n812 gnd 0.006956f
C3276 vdd.n813 gnd 0.006956f
C3277 vdd.n814 gnd 0.710887f
C3278 vdd.n815 gnd 0.006956f
C3279 vdd.n816 gnd 0.006956f
C3280 vdd.n817 gnd 0.601118f
C3281 vdd.n818 gnd 0.006956f
C3282 vdd.n819 gnd 0.006956f
C3283 vdd.n820 gnd 0.006956f
C3284 vdd.n821 gnd 0.006956f
C3285 vdd.n822 gnd 0.695206f
C3286 vdd.n823 gnd 0.006956f
C3287 vdd.n824 gnd 0.006956f
C3288 vdd.n825 gnd 0.006956f
C3289 vdd.n826 gnd 0.006956f
C3290 vdd.n827 gnd 0.006956f
C3291 vdd.n828 gnd 0.710887f
C3292 vdd.n829 gnd 0.006956f
C3293 vdd.n830 gnd 0.006956f
C3294 vdd.t10 gnd 0.355444f
C3295 vdd.n831 gnd 0.006956f
C3296 vdd.n832 gnd 0.006956f
C3297 vdd.n833 gnd 0.006956f
C3298 vdd.t7 gnd 0.355444f
C3299 vdd.n834 gnd 0.006956f
C3300 vdd.n835 gnd 0.006956f
C3301 vdd.n836 gnd 0.006956f
C3302 vdd.n837 gnd 0.006956f
C3303 vdd.n838 gnd 0.006956f
C3304 vdd.t73 gnd 0.297945f
C3305 vdd.n839 gnd 0.006956f
C3306 vdd.n840 gnd 0.006956f
C3307 vdd.n841 gnd 0.569755f
C3308 vdd.n842 gnd 0.006956f
C3309 vdd.t74 gnd 0.287738f
C3310 vdd.t72 gnd 0.183511f
C3311 vdd.t75 gnd 0.287738f
C3312 vdd.n843 gnd 0.161721f
C3313 vdd.n844 gnd 0.006956f
C3314 vdd.n845 gnd 0.006956f
C3315 vdd.n846 gnd 0.454759f
C3316 vdd.n847 gnd 0.006956f
C3317 vdd.n848 gnd 0.006956f
C3318 vdd.t19 gnd 0.104542f
C3319 vdd.n849 gnd 0.412942f
C3320 vdd.n850 gnd 0.006956f
C3321 vdd.n851 gnd 0.006956f
C3322 vdd.n852 gnd 0.006956f
C3323 vdd.n853 gnd 0.611572f
C3324 vdd.n854 gnd 0.006956f
C3325 vdd.n855 gnd 0.006956f
C3326 vdd.t36 gnd 0.355444f
C3327 vdd.n856 gnd 0.006956f
C3328 vdd.n857 gnd 0.006956f
C3329 vdd.n858 gnd 0.006956f
C3330 vdd.t48 gnd 0.355444f
C3331 vdd.n859 gnd 0.006956f
C3332 vdd.n860 gnd 0.006956f
C3333 vdd.t1 gnd 0.355444f
C3334 vdd.n861 gnd 0.006956f
C3335 vdd.n862 gnd 0.006956f
C3336 vdd.n863 gnd 0.006956f
C3337 vdd.t33 gnd 0.282264f
C3338 vdd.n864 gnd 0.006956f
C3339 vdd.n865 gnd 0.006956f
C3340 vdd.n866 gnd 0.585436f
C3341 vdd.n867 gnd 0.006956f
C3342 vdd.n868 gnd 0.006956f
C3343 vdd.n869 gnd 0.006956f
C3344 vdd.t45 gnd 0.355444f
C3345 vdd.n870 gnd 0.006956f
C3346 vdd.n871 gnd 0.006956f
C3347 vdd.t20 gnd 0.297945f
C3348 vdd.n872 gnd 0.428623f
C3349 vdd.n873 gnd 0.006956f
C3350 vdd.n874 gnd 0.006956f
C3351 vdd.n875 gnd 0.006956f
C3352 vdd.n876 gnd 0.371125f
C3353 vdd.n877 gnd 0.006956f
C3354 vdd.n878 gnd 0.006956f
C3355 vdd.t34 gnd 0.355444f
C3356 vdd.n879 gnd 0.006956f
C3357 vdd.n880 gnd 0.006956f
C3358 vdd.n881 gnd 0.006956f
C3359 vdd.n882 gnd 0.710887f
C3360 vdd.n883 gnd 0.006956f
C3361 vdd.n884 gnd 0.006956f
C3362 vdd.t11 gnd 0.240447f
C3363 vdd.t12 gnd 0.339762f
C3364 vdd.n885 gnd 0.006956f
C3365 vdd.n886 gnd 0.006956f
C3366 vdd.n887 gnd 0.006956f
C3367 vdd.n888 gnd 0.533165f
C3368 vdd.n889 gnd 0.006956f
C3369 vdd.n890 gnd 0.006956f
C3370 vdd.n891 gnd 0.006956f
C3371 vdd.n892 gnd 0.006956f
C3372 vdd.n893 gnd 0.006956f
C3373 vdd.t101 gnd 0.355444f
C3374 vdd.n894 gnd 0.006956f
C3375 vdd.n895 gnd 0.006956f
C3376 vdd.t29 gnd 0.355444f
C3377 vdd.n896 gnd 0.006956f
C3378 vdd.n897 gnd 0.015237f
C3379 vdd.n898 gnd 0.015237f
C3380 vdd.n899 gnd 0.846792f
C3381 vdd.n900 gnd 0.006956f
C3382 vdd.n901 gnd 0.006956f
C3383 vdd.t31 gnd 0.355444f
C3384 vdd.n902 gnd 0.015237f
C3385 vdd.n903 gnd 0.006956f
C3386 vdd.n904 gnd 0.006956f
C3387 vdd.t266 gnd 0.648162f
C3388 vdd.n922 gnd 0.01627f
C3389 vdd.n940 gnd 0.015237f
C3390 vdd.n941 gnd 0.006956f
C3391 vdd.n942 gnd 0.015237f
C3392 vdd.t116 gnd 0.281098f
C3393 vdd.t115 gnd 0.287738f
C3394 vdd.t114 gnd 0.183511f
C3395 vdd.n943 gnd 0.099178f
C3396 vdd.n944 gnd 0.056257f
C3397 vdd.n945 gnd 0.016101f
C3398 vdd.n946 gnd 0.006956f
C3399 vdd.n947 gnd 0.376352f
C3400 vdd.n948 gnd 0.015237f
C3401 vdd.n949 gnd 0.006956f
C3402 vdd.n950 gnd 0.01627f
C3403 vdd.n951 gnd 0.006956f
C3404 vdd.t99 gnd 0.281098f
C3405 vdd.t98 gnd 0.287738f
C3406 vdd.t96 gnd 0.183511f
C3407 vdd.n952 gnd 0.099178f
C3408 vdd.n953 gnd 0.056257f
C3409 vdd.n954 gnd 0.009941f
C3410 vdd.n955 gnd 0.006956f
C3411 vdd.n956 gnd 0.006956f
C3412 vdd.t97 gnd 0.355444f
C3413 vdd.n957 gnd 0.006956f
C3414 vdd.t5 gnd 0.355444f
C3415 vdd.n958 gnd 0.006956f
C3416 vdd.n959 gnd 0.006956f
C3417 vdd.n960 gnd 0.006956f
C3418 vdd.n961 gnd 0.006956f
C3419 vdd.n962 gnd 0.006956f
C3420 vdd.n963 gnd 0.710887f
C3421 vdd.n964 gnd 0.006956f
C3422 vdd.n965 gnd 0.006956f
C3423 vdd.t46 gnd 0.355444f
C3424 vdd.n966 gnd 0.006956f
C3425 vdd.n967 gnd 0.006956f
C3426 vdd.n968 gnd 0.006956f
C3427 vdd.n969 gnd 0.006956f
C3428 vdd.n970 gnd 0.47044f
C3429 vdd.n971 gnd 0.006956f
C3430 vdd.n972 gnd 0.006956f
C3431 vdd.n973 gnd 0.006956f
C3432 vdd.n974 gnd 0.006956f
C3433 vdd.n975 gnd 0.006956f
C3434 vdd.n976 gnd 0.627253f
C3435 vdd.n977 gnd 0.006956f
C3436 vdd.n978 gnd 0.006956f
C3437 vdd.t37 gnd 0.339762f
C3438 vdd.t9 gnd 0.240447f
C3439 vdd.n979 gnd 0.006956f
C3440 vdd.n980 gnd 0.006956f
C3441 vdd.n981 gnd 0.006956f
C3442 vdd.t8 gnd 0.355444f
C3443 vdd.n982 gnd 0.006956f
C3444 vdd.n983 gnd 0.006956f
C3445 vdd.t2 gnd 0.355444f
C3446 vdd.n984 gnd 0.006956f
C3447 vdd.n985 gnd 0.006956f
C3448 vdd.n986 gnd 0.006956f
C3449 vdd.t126 gnd 0.297945f
C3450 vdd.n987 gnd 0.006956f
C3451 vdd.n988 gnd 0.006956f
C3452 vdd.n989 gnd 0.569755f
C3453 vdd.n990 gnd 0.006956f
C3454 vdd.n991 gnd 0.006956f
C3455 vdd.n992 gnd 0.006956f
C3456 vdd.t24 gnd 0.355444f
C3457 vdd.n993 gnd 0.006956f
C3458 vdd.n994 gnd 0.006956f
C3459 vdd.t4 gnd 0.282264f
C3460 vdd.n995 gnd 0.412942f
C3461 vdd.n996 gnd 0.006956f
C3462 vdd.n997 gnd 0.006956f
C3463 vdd.n998 gnd 0.006956f
C3464 vdd.n999 gnd 0.611572f
C3465 vdd.n1000 gnd 0.006956f
C3466 vdd.n1001 gnd 0.006956f
C3467 vdd.t0 gnd 0.355444f
C3468 vdd.n1002 gnd 0.006956f
C3469 vdd.n1003 gnd 0.006956f
C3470 vdd.n1004 gnd 0.006956f
C3471 vdd.n1005 gnd 0.710887f
C3472 vdd.n1006 gnd 0.006956f
C3473 vdd.n1007 gnd 0.006956f
C3474 vdd.t23 gnd 0.355444f
C3475 vdd.n1008 gnd 0.006956f
C3476 vdd.n1009 gnd 0.006956f
C3477 vdd.n1010 gnd 0.006956f
C3478 vdd.t22 gnd 0.104542f
C3479 vdd.n1011 gnd 0.006956f
C3480 vdd.n1012 gnd 0.006956f
C3481 vdd.n1013 gnd 0.006956f
C3482 vdd.t106 gnd 0.287738f
C3483 vdd.t104 gnd 0.183511f
C3484 vdd.t107 gnd 0.287738f
C3485 vdd.n1014 gnd 0.161721f
C3486 vdd.n1015 gnd 0.006956f
C3487 vdd.n1016 gnd 0.006956f
C3488 vdd.t16 gnd 0.355444f
C3489 vdd.n1017 gnd 0.006956f
C3490 vdd.n1018 gnd 0.006956f
C3491 vdd.t105 gnd 0.297945f
C3492 vdd.n1019 gnd 0.606345f
C3493 vdd.n1020 gnd 0.006956f
C3494 vdd.n1021 gnd 0.006956f
C3495 vdd.n1022 gnd 0.006956f
C3496 vdd.n1023 gnd 0.371125f
C3497 vdd.n1024 gnd 0.006956f
C3498 vdd.n1025 gnd 0.006956f
C3499 vdd.n1026 gnd 0.496576f
C3500 vdd.n1027 gnd 0.006956f
C3501 vdd.n1028 gnd 0.006956f
C3502 vdd.n1029 gnd 0.006956f
C3503 vdd.n1030 gnd 0.710887f
C3504 vdd.n1031 gnd 0.006956f
C3505 vdd.n1032 gnd 0.006956f
C3506 vdd.t28 gnd 0.355444f
C3507 vdd.n1033 gnd 0.006956f
C3508 vdd.n1034 gnd 0.006956f
C3509 vdd.n1035 gnd 0.006956f
C3510 vdd.n1036 gnd 0.710887f
C3511 vdd.n1037 gnd 0.006956f
C3512 vdd.n1038 gnd 0.006956f
C3513 vdd.n1039 gnd 0.006956f
C3514 vdd.n1040 gnd 0.006956f
C3515 vdd.n1041 gnd 0.006956f
C3516 vdd.t55 gnd 0.355444f
C3517 vdd.n1042 gnd 0.006956f
C3518 vdd.n1043 gnd 0.006956f
C3519 vdd.n1044 gnd 0.006956f
C3520 vdd.n1045 gnd 0.015237f
C3521 vdd.n1046 gnd 0.015237f
C3522 vdd.n1047 gnd 1.00361f
C3523 vdd.n1048 gnd 0.006956f
C3524 vdd.n1049 gnd 0.006956f
C3525 vdd.n1050 gnd 0.465213f
C3526 vdd.n1051 gnd 0.015237f
C3527 vdd.n1052 gnd 0.006956f
C3528 vdd.n1053 gnd 0.006956f
C3529 vdd.n1054 gnd 9.12654f
C3530 vdd.n1087 gnd 0.01627f
C3531 vdd.n1088 gnd 0.006956f
C3532 vdd.n1089 gnd 0.006956f
C3533 vdd.n1090 gnd 0.006956f
C3534 vdd.n1091 gnd 0.006547f
C3535 vdd.n1094 gnd 0.023454f
C3536 vdd.n1095 gnd 0.006834f
C3537 vdd.n1096 gnd 0.008234f
C3538 vdd.n1098 gnd 0.01023f
C3539 vdd.n1099 gnd 0.01023f
C3540 vdd.n1100 gnd 0.008234f
C3541 vdd.n1102 gnd 0.01023f
C3542 vdd.n1103 gnd 0.01023f
C3543 vdd.n1104 gnd 0.01023f
C3544 vdd.n1105 gnd 0.01023f
C3545 vdd.n1106 gnd 0.01023f
C3546 vdd.n1107 gnd 0.008234f
C3547 vdd.n1109 gnd 0.01023f
C3548 vdd.n1110 gnd 0.01023f
C3549 vdd.n1111 gnd 0.01023f
C3550 vdd.n1112 gnd 0.01023f
C3551 vdd.n1113 gnd 0.01023f
C3552 vdd.n1114 gnd 0.008234f
C3553 vdd.n1116 gnd 0.01023f
C3554 vdd.n1117 gnd 0.01023f
C3555 vdd.n1118 gnd 0.01023f
C3556 vdd.n1119 gnd 0.01023f
C3557 vdd.n1120 gnd 0.006875f
C3558 vdd.t110 gnd 0.125851f
C3559 vdd.t109 gnd 0.134501f
C3560 vdd.t108 gnd 0.164361f
C3561 vdd.n1121 gnd 0.210687f
C3562 vdd.n1122 gnd 0.177015f
C3563 vdd.n1124 gnd 0.01023f
C3564 vdd.n1125 gnd 0.01023f
C3565 vdd.n1126 gnd 0.008234f
C3566 vdd.n1127 gnd 0.01023f
C3567 vdd.n1129 gnd 0.01023f
C3568 vdd.n1130 gnd 0.01023f
C3569 vdd.n1131 gnd 0.01023f
C3570 vdd.n1132 gnd 0.01023f
C3571 vdd.n1133 gnd 0.008234f
C3572 vdd.n1135 gnd 0.01023f
C3573 vdd.n1136 gnd 0.01023f
C3574 vdd.n1137 gnd 0.01023f
C3575 vdd.n1138 gnd 0.01023f
C3576 vdd.n1139 gnd 0.01023f
C3577 vdd.n1140 gnd 0.008234f
C3578 vdd.n1142 gnd 0.01023f
C3579 vdd.n1143 gnd 0.01023f
C3580 vdd.n1144 gnd 0.01023f
C3581 vdd.n1145 gnd 0.01023f
C3582 vdd.n1146 gnd 0.01023f
C3583 vdd.n1147 gnd 0.008234f
C3584 vdd.n1149 gnd 0.01023f
C3585 vdd.n1150 gnd 0.01023f
C3586 vdd.n1151 gnd 0.01023f
C3587 vdd.n1152 gnd 0.01023f
C3588 vdd.n1153 gnd 0.01023f
C3589 vdd.n1154 gnd 0.008234f
C3590 vdd.n1156 gnd 0.01023f
C3591 vdd.n1157 gnd 0.01023f
C3592 vdd.n1158 gnd 0.01023f
C3593 vdd.n1159 gnd 0.01023f
C3594 vdd.n1160 gnd 0.008151f
C3595 vdd.t95 gnd 0.125851f
C3596 vdd.t94 gnd 0.134501f
C3597 vdd.t93 gnd 0.164361f
C3598 vdd.n1161 gnd 0.210687f
C3599 vdd.n1162 gnd 0.177015f
C3600 vdd.n1164 gnd 0.01023f
C3601 vdd.n1165 gnd 0.01023f
C3602 vdd.n1166 gnd 0.008234f
C3603 vdd.n1167 gnd 0.01023f
C3604 vdd.n1169 gnd 0.01023f
C3605 vdd.n1170 gnd 0.01023f
C3606 vdd.n1171 gnd 0.01023f
C3607 vdd.n1172 gnd 0.01023f
C3608 vdd.n1173 gnd 0.008234f
C3609 vdd.n1175 gnd 0.01023f
C3610 vdd.n1176 gnd 0.01023f
C3611 vdd.n1177 gnd 0.01023f
C3612 vdd.n1178 gnd 0.01023f
C3613 vdd.n1179 gnd 0.01023f
C3614 vdd.n1180 gnd 0.008234f
C3615 vdd.n1182 gnd 0.01023f
C3616 vdd.n1183 gnd 0.01023f
C3617 vdd.n1184 gnd 0.01023f
C3618 vdd.n1185 gnd 0.01023f
C3619 vdd.n1186 gnd 0.01023f
C3620 vdd.n1187 gnd 0.008234f
C3621 vdd.n1189 gnd 0.01023f
C3622 vdd.n1190 gnd 0.01023f
C3623 vdd.n1191 gnd 0.006547f
C3624 vdd.n1192 gnd 0.008234f
C3625 vdd.n1193 gnd 0.006956f
C3626 vdd.n1194 gnd 0.006956f
C3627 vdd.n1195 gnd 0.006956f
C3628 vdd.n1196 gnd 0.006956f
C3629 vdd.n1197 gnd 0.006956f
C3630 vdd.n1198 gnd 0.006956f
C3631 vdd.n1199 gnd 0.006956f
C3632 vdd.n1200 gnd 0.006956f
C3633 vdd.n1201 gnd 0.006956f
C3634 vdd.n1202 gnd 0.006956f
C3635 vdd.n1203 gnd 0.006956f
C3636 vdd.n1204 gnd 0.006956f
C3637 vdd.n1205 gnd 0.006956f
C3638 vdd.n1206 gnd 0.006956f
C3639 vdd.n1207 gnd 0.006956f
C3640 vdd.n1208 gnd 0.006956f
C3641 vdd.n1209 gnd 0.006956f
C3642 vdd.n1210 gnd 0.006956f
C3643 vdd.n1211 gnd 0.006956f
C3644 vdd.n1212 gnd 0.006956f
C3645 vdd.n1213 gnd 0.006956f
C3646 vdd.n1214 gnd 0.006956f
C3647 vdd.n1215 gnd 0.006956f
C3648 vdd.n1216 gnd 0.006956f
C3649 vdd.n1217 gnd 0.006956f
C3650 vdd.n1218 gnd 0.006956f
C3651 vdd.n1219 gnd 0.006956f
C3652 vdd.n1220 gnd 0.006956f
C3653 vdd.n1221 gnd 0.006956f
C3654 vdd.n1222 gnd 0.006956f
C3655 vdd.n1223 gnd 0.006956f
C3656 vdd.t56 gnd 0.281098f
C3657 vdd.t57 gnd 0.287738f
C3658 vdd.t54 gnd 0.183511f
C3659 vdd.n1224 gnd 0.099178f
C3660 vdd.n1225 gnd 0.056257f
C3661 vdd.n1226 gnd 0.009941f
C3662 vdd.n1227 gnd 0.006956f
C3663 vdd.n1228 gnd 0.006956f
C3664 vdd.n1229 gnd 0.006956f
C3665 vdd.n1230 gnd 0.006956f
C3666 vdd.n1231 gnd 0.006956f
C3667 vdd.n1232 gnd 0.006956f
C3668 vdd.n1233 gnd 0.006956f
C3669 vdd.n1234 gnd 0.006956f
C3670 vdd.n1235 gnd 0.006956f
C3671 vdd.n1236 gnd 0.006956f
C3672 vdd.n1237 gnd 0.006956f
C3673 vdd.n1238 gnd 0.006956f
C3674 vdd.n1239 gnd 0.006956f
C3675 vdd.n1240 gnd 0.006956f
C3676 vdd.n1241 gnd 0.006956f
C3677 vdd.n1242 gnd 0.006956f
C3678 vdd.n1243 gnd 0.006956f
C3679 vdd.t70 gnd 0.281098f
C3680 vdd.t71 gnd 0.287738f
C3681 vdd.t69 gnd 0.183511f
C3682 vdd.n1244 gnd 0.099178f
C3683 vdd.n1245 gnd 0.056257f
C3684 vdd.n1246 gnd 0.006956f
C3685 vdd.n1247 gnd 0.006956f
C3686 vdd.n1248 gnd 0.006956f
C3687 vdd.n1249 gnd 0.006956f
C3688 vdd.n1250 gnd 0.006956f
C3689 vdd.n1251 gnd 0.006956f
C3690 vdd.n1252 gnd 0.006956f
C3691 vdd.n1253 gnd 0.006956f
C3692 vdd.n1254 gnd 0.006956f
C3693 vdd.n1255 gnd 0.006956f
C3694 vdd.n1256 gnd 0.006956f
C3695 vdd.n1257 gnd 0.006956f
C3696 vdd.n1258 gnd 0.006956f
C3697 vdd.n1259 gnd 0.006956f
C3698 vdd.n1260 gnd 0.006956f
C3699 vdd.n1261 gnd 0.006956f
C3700 vdd.n1262 gnd 0.006956f
C3701 vdd.n1263 gnd 0.006956f
C3702 vdd.n1264 gnd 0.006956f
C3703 vdd.n1265 gnd 0.006956f
C3704 vdd.n1266 gnd 0.006956f
C3705 vdd.n1267 gnd 0.006956f
C3706 vdd.n1268 gnd 0.006956f
C3707 vdd.n1269 gnd 0.006956f
C3708 vdd.n1270 gnd 0.006956f
C3709 vdd.n1271 gnd 0.006956f
C3710 vdd.n1272 gnd 0.005064f
C3711 vdd.n1273 gnd 0.009941f
C3712 vdd.n1274 gnd 0.005371f
C3713 vdd.n1275 gnd 0.006956f
C3714 vdd.n1276 gnd 0.006956f
C3715 vdd.n1277 gnd 0.006956f
C3716 vdd.n1278 gnd 0.01627f
C3717 vdd.n1279 gnd 0.01627f
C3718 vdd.n1280 gnd 0.015237f
C3719 vdd.n1281 gnd 0.015237f
C3720 vdd.n1282 gnd 0.006956f
C3721 vdd.n1283 gnd 0.006956f
C3722 vdd.n1284 gnd 0.006956f
C3723 vdd.n1285 gnd 0.006956f
C3724 vdd.n1286 gnd 0.006956f
C3725 vdd.n1287 gnd 0.006956f
C3726 vdd.n1288 gnd 0.006956f
C3727 vdd.n1289 gnd 0.006956f
C3728 vdd.n1290 gnd 0.006956f
C3729 vdd.n1291 gnd 0.006956f
C3730 vdd.n1292 gnd 0.006956f
C3731 vdd.n1293 gnd 0.006956f
C3732 vdd.n1294 gnd 0.006956f
C3733 vdd.n1295 gnd 0.006956f
C3734 vdd.n1296 gnd 0.006956f
C3735 vdd.n1297 gnd 0.006956f
C3736 vdd.n1298 gnd 0.006956f
C3737 vdd.n1299 gnd 0.006956f
C3738 vdd.n1300 gnd 0.006956f
C3739 vdd.n1301 gnd 0.006956f
C3740 vdd.n1302 gnd 0.006956f
C3741 vdd.n1303 gnd 0.006956f
C3742 vdd.n1304 gnd 0.006956f
C3743 vdd.n1305 gnd 0.006956f
C3744 vdd.n1306 gnd 0.006956f
C3745 vdd.n1307 gnd 0.006956f
C3746 vdd.n1308 gnd 0.006956f
C3747 vdd.n1309 gnd 0.423396f
C3748 vdd.n1310 gnd 0.006956f
C3749 vdd.n1311 gnd 0.006956f
C3750 vdd.n1312 gnd 0.006956f
C3751 vdd.n1313 gnd 0.006956f
C3752 vdd.n1314 gnd 0.006956f
C3753 vdd.n1315 gnd 0.006956f
C3754 vdd.n1316 gnd 0.006956f
C3755 vdd.n1317 gnd 0.006956f
C3756 vdd.n1318 gnd 0.006956f
C3757 vdd.n1319 gnd 0.006956f
C3758 vdd.n1320 gnd 0.006956f
C3759 vdd.n1321 gnd 0.006956f
C3760 vdd.n1322 gnd 0.006956f
C3761 vdd.n1323 gnd 0.006956f
C3762 vdd.n1324 gnd 0.006956f
C3763 vdd.n1325 gnd 0.006956f
C3764 vdd.n1326 gnd 0.006956f
C3765 vdd.n1327 gnd 0.006956f
C3766 vdd.n1328 gnd 0.006956f
C3767 vdd.n1329 gnd 0.006956f
C3768 vdd.n1330 gnd 0.224766f
C3769 vdd.n1331 gnd 0.006956f
C3770 vdd.n1332 gnd 0.006956f
C3771 vdd.n1333 gnd 0.006956f
C3772 vdd.n1334 gnd 0.006956f
C3773 vdd.n1335 gnd 0.006956f
C3774 vdd.n1336 gnd 0.006956f
C3775 vdd.n1337 gnd 0.006956f
C3776 vdd.n1338 gnd 0.006956f
C3777 vdd.n1339 gnd 0.006956f
C3778 vdd.n1340 gnd 0.006956f
C3779 vdd.n1341 gnd 0.006956f
C3780 vdd.n1342 gnd 0.006956f
C3781 vdd.n1343 gnd 0.006956f
C3782 vdd.n1344 gnd 0.006956f
C3783 vdd.n1345 gnd 0.006956f
C3784 vdd.n1346 gnd 0.006956f
C3785 vdd.n1347 gnd 0.006956f
C3786 vdd.n1348 gnd 0.006956f
C3787 vdd.n1349 gnd 0.006956f
C3788 vdd.n1350 gnd 0.006956f
C3789 vdd.n1351 gnd 0.006956f
C3790 vdd.n1352 gnd 0.006956f
C3791 vdd.n1353 gnd 0.006956f
C3792 vdd.n1354 gnd 0.006956f
C3793 vdd.n1355 gnd 0.006956f
C3794 vdd.n1356 gnd 0.006956f
C3795 vdd.n1357 gnd 0.006956f
C3796 vdd.n1358 gnd 0.015237f
C3797 vdd.n1359 gnd 0.015237f
C3798 vdd.n1360 gnd 0.01627f
C3799 vdd.n1361 gnd 0.006956f
C3800 vdd.n1362 gnd 0.006956f
C3801 vdd.n1363 gnd 0.005371f
C3802 vdd.n1364 gnd 0.006956f
C3803 vdd.n1365 gnd 0.006956f
C3804 vdd.n1366 gnd 0.005064f
C3805 vdd.n1367 gnd 0.006956f
C3806 vdd.n1368 gnd 0.006956f
C3807 vdd.n1369 gnd 0.006956f
C3808 vdd.n1370 gnd 0.006956f
C3809 vdd.n1371 gnd 0.006956f
C3810 vdd.n1372 gnd 0.006956f
C3811 vdd.n1373 gnd 0.006956f
C3812 vdd.n1374 gnd 0.006956f
C3813 vdd.n1375 gnd 0.006956f
C3814 vdd.n1376 gnd 0.006956f
C3815 vdd.n1377 gnd 0.006956f
C3816 vdd.n1378 gnd 0.006956f
C3817 vdd.n1379 gnd 0.006956f
C3818 vdd.n1380 gnd 0.006956f
C3819 vdd.n1381 gnd 0.006956f
C3820 vdd.n1382 gnd 0.006956f
C3821 vdd.n1383 gnd 0.006956f
C3822 vdd.n1384 gnd 0.006956f
C3823 vdd.n1385 gnd 0.006956f
C3824 vdd.n1386 gnd 0.006956f
C3825 vdd.n1387 gnd 0.006956f
C3826 vdd.n1388 gnd 0.006956f
C3827 vdd.n1389 gnd 0.006956f
C3828 vdd.n1390 gnd 0.006956f
C3829 vdd.n1391 gnd 0.006956f
C3830 vdd.n1392 gnd 0.006956f
C3831 vdd.n1393 gnd 0.02788f
C3832 vdd.n1395 gnd 0.023454f
C3833 vdd.n1396 gnd 0.008234f
C3834 vdd.n1398 gnd 0.01023f
C3835 vdd.n1399 gnd 0.008234f
C3836 vdd.n1400 gnd 0.01023f
C3837 vdd.n1402 gnd 0.01023f
C3838 vdd.n1403 gnd 0.01023f
C3839 vdd.n1405 gnd 0.01023f
C3840 vdd.n1406 gnd 0.006834f
C3841 vdd.n1407 gnd 0.580209f
C3842 vdd.n1408 gnd 0.01023f
C3843 vdd.n1409 gnd 0.023454f
C3844 vdd.n1410 gnd 0.008234f
C3845 vdd.n1411 gnd 0.01023f
C3846 vdd.n1412 gnd 0.008234f
C3847 vdd.n1413 gnd 0.01023f
C3848 vdd.n1414 gnd 1.04542f
C3849 vdd.n1415 gnd 0.01023f
C3850 vdd.n1416 gnd 0.008234f
C3851 vdd.n1417 gnd 0.008234f
C3852 vdd.n1418 gnd 0.01023f
C3853 vdd.n1419 gnd 0.008234f
C3854 vdd.n1420 gnd 0.01023f
C3855 vdd.t179 gnd 0.522711f
C3856 vdd.n1421 gnd 0.01023f
C3857 vdd.n1422 gnd 0.008234f
C3858 vdd.n1423 gnd 0.01023f
C3859 vdd.n1424 gnd 0.008234f
C3860 vdd.n1425 gnd 0.01023f
C3861 vdd.t142 gnd 0.522711f
C3862 vdd.n1426 gnd 0.01023f
C3863 vdd.n1427 gnd 0.008234f
C3864 vdd.n1428 gnd 0.01023f
C3865 vdd.n1429 gnd 0.008234f
C3866 vdd.n1430 gnd 0.01023f
C3867 vdd.t203 gnd 0.522711f
C3868 vdd.n1431 gnd 0.726568f
C3869 vdd.n1432 gnd 0.01023f
C3870 vdd.n1433 gnd 0.008234f
C3871 vdd.n1434 gnd 0.01023f
C3872 vdd.n1435 gnd 0.008234f
C3873 vdd.n1436 gnd 0.01023f
C3874 vdd.n1437 gnd 0.831111f
C3875 vdd.n1438 gnd 0.01023f
C3876 vdd.n1439 gnd 0.008234f
C3877 vdd.n1440 gnd 0.01023f
C3878 vdd.n1441 gnd 0.008234f
C3879 vdd.n1442 gnd 0.01023f
C3880 vdd.n1443 gnd 0.653389f
C3881 vdd.t220 gnd 0.522711f
C3882 vdd.n1444 gnd 0.01023f
C3883 vdd.n1445 gnd 0.008234f
C3884 vdd.n1446 gnd 0.01023f
C3885 vdd.n1447 gnd 0.008234f
C3886 vdd.n1448 gnd 0.01023f
C3887 vdd.t194 gnd 0.522711f
C3888 vdd.n1449 gnd 0.01023f
C3889 vdd.n1450 gnd 0.008234f
C3890 vdd.n1451 gnd 0.01023f
C3891 vdd.n1452 gnd 0.008234f
C3892 vdd.n1453 gnd 0.01023f
C3893 vdd.t158 gnd 0.522711f
C3894 vdd.n1454 gnd 0.569755f
C3895 vdd.n1455 gnd 0.01023f
C3896 vdd.n1456 gnd 0.008234f
C3897 vdd.n1457 gnd 0.01023f
C3898 vdd.n1458 gnd 0.008234f
C3899 vdd.n1459 gnd 0.01023f
C3900 vdd.t174 gnd 0.522711f
C3901 vdd.n1460 gnd 0.01023f
C3902 vdd.n1461 gnd 0.008234f
C3903 vdd.n1462 gnd 0.01023f
C3904 vdd.n1463 gnd 0.008234f
C3905 vdd.n1464 gnd 0.01023f
C3906 vdd.n1465 gnd 0.810202f
C3907 vdd.n1466 gnd 0.8677f
C3908 vdd.t215 gnd 0.522711f
C3909 vdd.n1467 gnd 0.01023f
C3910 vdd.n1468 gnd 0.008234f
C3911 vdd.n1469 gnd 0.01023f
C3912 vdd.n1470 gnd 0.008234f
C3913 vdd.n1471 gnd 0.01023f
C3914 vdd.n1472 gnd 0.63248f
C3915 vdd.n1473 gnd 0.01023f
C3916 vdd.n1474 gnd 0.008234f
C3917 vdd.n1475 gnd 0.01023f
C3918 vdd.n1476 gnd 0.008234f
C3919 vdd.n1477 gnd 0.01023f
C3920 vdd.t170 gnd 0.522711f
C3921 vdd.t148 gnd 0.522711f
C3922 vdd.n1478 gnd 0.01023f
C3923 vdd.n1479 gnd 0.008234f
C3924 vdd.n1480 gnd 0.01023f
C3925 vdd.n1481 gnd 0.008234f
C3926 vdd.n1482 gnd 0.01023f
C3927 vdd.t172 gnd 0.522711f
C3928 vdd.n1483 gnd 0.01023f
C3929 vdd.n1484 gnd 0.008234f
C3930 vdd.n1485 gnd 0.01023f
C3931 vdd.n1486 gnd 0.008234f
C3932 vdd.n1487 gnd 0.01023f
C3933 vdd.t140 gnd 0.522711f
C3934 vdd.n1488 gnd 0.768385f
C3935 vdd.n1489 gnd 0.01023f
C3936 vdd.n1490 gnd 0.008234f
C3937 vdd.n1491 gnd 0.01023f
C3938 vdd.n1492 gnd 0.008234f
C3939 vdd.n1493 gnd 0.01023f
C3940 vdd.n1494 gnd 1.04542f
C3941 vdd.n1495 gnd 0.01023f
C3942 vdd.n1496 gnd 0.008234f
C3943 vdd.n1497 gnd 0.01023f
C3944 vdd.n1498 gnd 0.008234f
C3945 vdd.n1499 gnd 0.01023f
C3946 vdd.n1500 gnd 0.883382f
C3947 vdd.n1501 gnd 0.01023f
C3948 vdd.n1502 gnd 0.008234f
C3949 vdd.n1503 gnd 0.023295f
C3950 vdd.n1504 gnd 0.006834f
C3951 vdd.n1505 gnd 0.023295f
C3952 vdd.n1506 gnd 1.37996f
C3953 vdd.n1507 gnd 0.023295f
C3954 vdd.n1508 gnd 0.006834f
C3955 vdd.n1509 gnd 0.01023f
C3956 vdd.t88 gnd 0.125851f
C3957 vdd.t89 gnd 0.134501f
C3958 vdd.t87 gnd 0.164361f
C3959 vdd.n1510 gnd 0.210687f
C3960 vdd.n1511 gnd 0.177839f
C3961 vdd.n1512 gnd 0.013503f
C3962 vdd.n1513 gnd 0.01023f
C3963 vdd.n1544 gnd 0.01023f
C3964 vdd.n1545 gnd 0.01023f
C3965 vdd.n1546 gnd 0.023454f
C3966 vdd.n1547 gnd 0.008234f
C3967 vdd.n1548 gnd 0.01023f
C3968 vdd.n1549 gnd 0.01023f
C3969 vdd.n1550 gnd 0.01023f
C3970 vdd.n1551 gnd 0.01023f
C3971 vdd.n1552 gnd 0.008234f
C3972 vdd.n1553 gnd 0.01023f
C3973 vdd.n1554 gnd 0.01023f
C3974 vdd.n1555 gnd 0.01023f
C3975 vdd.n1556 gnd 0.01023f
C3976 vdd.n1557 gnd 0.01023f
C3977 vdd.n1558 gnd 0.008234f
C3978 vdd.n1559 gnd 0.01023f
C3979 vdd.n1560 gnd 0.01023f
C3980 vdd.n1561 gnd 0.01023f
C3981 vdd.n1562 gnd 0.01023f
C3982 vdd.n1563 gnd 0.01023f
C3983 vdd.n1564 gnd 0.008234f
C3984 vdd.n1565 gnd 0.01023f
C3985 vdd.n1566 gnd 0.01023f
C3986 vdd.n1567 gnd 0.01023f
C3987 vdd.n1568 gnd 0.01023f
C3988 vdd.n1569 gnd 0.01023f
C3989 vdd.n1570 gnd 0.006875f
C3990 vdd.n1571 gnd 0.01023f
C3991 vdd.n1572 gnd 0.01023f
C3992 vdd.n1573 gnd 0.01023f
C3993 vdd.n1574 gnd 0.008234f
C3994 vdd.n1575 gnd 0.01023f
C3995 vdd.n1576 gnd 0.01023f
C3996 vdd.n1577 gnd 0.01023f
C3997 vdd.n1578 gnd 0.01023f
C3998 vdd.n1579 gnd 0.01023f
C3999 vdd.n1580 gnd 0.008234f
C4000 vdd.n1581 gnd 0.01023f
C4001 vdd.n1582 gnd 0.01023f
C4002 vdd.n1583 gnd 0.01023f
C4003 vdd.n1584 gnd 0.01023f
C4004 vdd.n1585 gnd 0.01023f
C4005 vdd.n1586 gnd 0.008234f
C4006 vdd.n1587 gnd 0.01023f
C4007 vdd.n1588 gnd 0.01023f
C4008 vdd.n1589 gnd 0.01023f
C4009 vdd.n1590 gnd 0.01023f
C4010 vdd.n1591 gnd 0.01023f
C4011 vdd.n1592 gnd 0.008234f
C4012 vdd.n1593 gnd 0.01023f
C4013 vdd.n1594 gnd 0.01023f
C4014 vdd.n1595 gnd 0.01023f
C4015 vdd.n1596 gnd 0.01023f
C4016 vdd.n1597 gnd 0.01023f
C4017 vdd.n1598 gnd 0.008234f
C4018 vdd.n1599 gnd 0.01023f
C4019 vdd.n1600 gnd 0.01023f
C4020 vdd.n1601 gnd 0.01023f
C4021 vdd.n1602 gnd 0.01023f
C4022 vdd.n1603 gnd 0.008151f
C4023 vdd.n1604 gnd 0.01023f
C4024 vdd.n1605 gnd 0.01023f
C4025 vdd.n1606 gnd 0.01023f
C4026 vdd.n1607 gnd 0.01023f
C4027 vdd.n1608 gnd 0.01023f
C4028 vdd.n1609 gnd 0.008234f
C4029 vdd.n1610 gnd 0.01023f
C4030 vdd.n1611 gnd 0.01023f
C4031 vdd.n1612 gnd 0.01023f
C4032 vdd.n1613 gnd 0.01023f
C4033 vdd.n1614 gnd 0.01023f
C4034 vdd.n1615 gnd 0.008234f
C4035 vdd.n1616 gnd 0.01023f
C4036 vdd.n1617 gnd 0.01023f
C4037 vdd.n1618 gnd 0.01023f
C4038 vdd.n1619 gnd 0.01023f
C4039 vdd.n1620 gnd 0.01023f
C4040 vdd.n1621 gnd 0.008234f
C4041 vdd.n1622 gnd 0.01023f
C4042 vdd.n1623 gnd 0.01023f
C4043 vdd.n1624 gnd 0.01023f
C4044 vdd.n1625 gnd 0.01023f
C4045 vdd.n1626 gnd 0.01023f
C4046 vdd.n1627 gnd 0.008234f
C4047 vdd.n1628 gnd 0.01023f
C4048 vdd.n1629 gnd 0.01023f
C4049 vdd.n1630 gnd 0.01023f
C4050 vdd.n1631 gnd 0.01023f
C4051 vdd.n1632 gnd 0.01023f
C4052 vdd.n1633 gnd 0.004323f
C4053 vdd.n1634 gnd 0.01023f
C4054 vdd.n1635 gnd 0.008234f
C4055 vdd.n1636 gnd 0.008234f
C4056 vdd.n1637 gnd 0.008234f
C4057 vdd.n1638 gnd 0.01023f
C4058 vdd.n1639 gnd 0.01023f
C4059 vdd.n1640 gnd 0.01023f
C4060 vdd.n1641 gnd 0.008234f
C4061 vdd.n1642 gnd 0.008234f
C4062 vdd.n1643 gnd 0.008234f
C4063 vdd.n1644 gnd 0.01023f
C4064 vdd.n1645 gnd 0.01023f
C4065 vdd.n1646 gnd 0.01023f
C4066 vdd.n1647 gnd 0.008234f
C4067 vdd.n1648 gnd 0.008234f
C4068 vdd.n1649 gnd 0.008234f
C4069 vdd.n1650 gnd 0.01023f
C4070 vdd.n1651 gnd 0.01023f
C4071 vdd.n1652 gnd 0.01023f
C4072 vdd.n1653 gnd 0.008234f
C4073 vdd.n1654 gnd 0.008234f
C4074 vdd.n1655 gnd 0.008234f
C4075 vdd.n1656 gnd 0.01023f
C4076 vdd.n1657 gnd 0.01023f
C4077 vdd.n1658 gnd 0.01023f
C4078 vdd.n1659 gnd 0.008234f
C4079 vdd.n1660 gnd 0.008234f
C4080 vdd.n1661 gnd 0.008234f
C4081 vdd.n1662 gnd 0.01023f
C4082 vdd.n1663 gnd 0.01023f
C4083 vdd.n1664 gnd 0.01023f
C4084 vdd.n1665 gnd 0.01023f
C4085 vdd.t81 gnd 0.125851f
C4086 vdd.t82 gnd 0.134501f
C4087 vdd.t79 gnd 0.164361f
C4088 vdd.n1666 gnd 0.210687f
C4089 vdd.n1667 gnd 0.177839f
C4090 vdd.n1668 gnd 0.01762f
C4091 vdd.n1669 gnd 0.005599f
C4092 vdd.n1670 gnd 0.008234f
C4093 vdd.n1671 gnd 0.01023f
C4094 vdd.n1672 gnd 0.01023f
C4095 vdd.n1673 gnd 0.01023f
C4096 vdd.n1674 gnd 0.008234f
C4097 vdd.n1675 gnd 0.008234f
C4098 vdd.n1676 gnd 0.008234f
C4099 vdd.n1677 gnd 0.01023f
C4100 vdd.n1678 gnd 0.01023f
C4101 vdd.n1679 gnd 0.01023f
C4102 vdd.n1680 gnd 0.008234f
C4103 vdd.n1681 gnd 0.008234f
C4104 vdd.n1682 gnd 0.008234f
C4105 vdd.n1683 gnd 0.01023f
C4106 vdd.n1684 gnd 0.01023f
C4107 vdd.n1685 gnd 0.01023f
C4108 vdd.n1686 gnd 0.008234f
C4109 vdd.n1687 gnd 0.008234f
C4110 vdd.n1688 gnd 0.008234f
C4111 vdd.n1689 gnd 0.01023f
C4112 vdd.n1690 gnd 0.01023f
C4113 vdd.n1691 gnd 0.01023f
C4114 vdd.n1692 gnd 0.008234f
C4115 vdd.n1693 gnd 0.008234f
C4116 vdd.n1694 gnd 0.008234f
C4117 vdd.n1695 gnd 0.01023f
C4118 vdd.n1696 gnd 0.01023f
C4119 vdd.n1697 gnd 0.01023f
C4120 vdd.n1698 gnd 0.008234f
C4121 vdd.n1699 gnd 0.006875f
C4122 vdd.n1700 gnd 0.01023f
C4123 vdd.n1701 gnd 0.01023f
C4124 vdd.t91 gnd 0.125851f
C4125 vdd.t92 gnd 0.134501f
C4126 vdd.t90 gnd 0.164361f
C4127 vdd.n1702 gnd 0.210687f
C4128 vdd.n1703 gnd 0.177839f
C4129 vdd.n1704 gnd 0.01762f
C4130 vdd.n1705 gnd 0.01023f
C4131 vdd.n1706 gnd 0.01023f
C4132 vdd.n1707 gnd 0.01023f
C4133 vdd.n1708 gnd 0.008234f
C4134 vdd.n1709 gnd 0.008234f
C4135 vdd.n1710 gnd 0.008234f
C4136 vdd.n1711 gnd 0.01023f
C4137 vdd.n1712 gnd 0.01023f
C4138 vdd.n1713 gnd 0.01023f
C4139 vdd.n1714 gnd 0.008234f
C4140 vdd.n1715 gnd 0.008234f
C4141 vdd.n1716 gnd 0.008234f
C4142 vdd.n1717 gnd 0.01023f
C4143 vdd.n1718 gnd 0.01023f
C4144 vdd.n1719 gnd 0.01023f
C4145 vdd.n1720 gnd 0.008234f
C4146 vdd.n1721 gnd 0.008234f
C4147 vdd.n1722 gnd 0.008234f
C4148 vdd.n1723 gnd 0.01023f
C4149 vdd.n1724 gnd 0.01023f
C4150 vdd.n1725 gnd 0.01023f
C4151 vdd.n1726 gnd 0.008234f
C4152 vdd.n1727 gnd 0.008234f
C4153 vdd.n1728 gnd 0.008234f
C4154 vdd.n1729 gnd 0.01023f
C4155 vdd.n1730 gnd 0.01023f
C4156 vdd.n1731 gnd 0.01023f
C4157 vdd.n1732 gnd 0.008234f
C4158 vdd.n1733 gnd 0.006834f
C4159 vdd.n1734 gnd 0.023454f
C4160 vdd.n1736 gnd 2.31038f
C4161 vdd.n1737 gnd 0.023454f
C4162 vdd.n1738 gnd 0.003911f
C4163 vdd.n1739 gnd 0.023454f
C4164 vdd.n1740 gnd 0.023295f
C4165 vdd.n1741 gnd 0.01023f
C4166 vdd.n1742 gnd 0.008234f
C4167 vdd.n1743 gnd 0.01023f
C4168 vdd.t80 gnd 0.522711f
C4169 vdd.n1744 gnd 0.684752f
C4170 vdd.n1745 gnd 0.01023f
C4171 vdd.n1746 gnd 0.008234f
C4172 vdd.n1747 gnd 0.01023f
C4173 vdd.n1748 gnd 0.01023f
C4174 vdd.n1749 gnd 0.01023f
C4175 vdd.n1750 gnd 0.008234f
C4176 vdd.n1751 gnd 0.01023f
C4177 vdd.n1752 gnd 1.04542f
C4178 vdd.n1753 gnd 0.01023f
C4179 vdd.n1754 gnd 0.008234f
C4180 vdd.n1755 gnd 0.01023f
C4181 vdd.n1756 gnd 0.01023f
C4182 vdd.n1757 gnd 0.01023f
C4183 vdd.n1758 gnd 0.008234f
C4184 vdd.n1759 gnd 0.01023f
C4185 vdd.n1760 gnd 0.8677f
C4186 vdd.t144 gnd 0.522711f
C4187 vdd.n1761 gnd 0.601118f
C4188 vdd.n1762 gnd 0.01023f
C4189 vdd.n1763 gnd 0.008234f
C4190 vdd.n1764 gnd 0.01023f
C4191 vdd.n1765 gnd 0.01023f
C4192 vdd.n1766 gnd 0.01023f
C4193 vdd.n1767 gnd 0.008234f
C4194 vdd.n1768 gnd 0.01023f
C4195 vdd.n1769 gnd 0.622026f
C4196 vdd.n1770 gnd 0.01023f
C4197 vdd.n1771 gnd 0.008234f
C4198 vdd.n1772 gnd 0.01023f
C4199 vdd.n1773 gnd 0.01023f
C4200 vdd.n1774 gnd 0.01023f
C4201 vdd.n1775 gnd 0.008234f
C4202 vdd.n1776 gnd 0.01023f
C4203 vdd.n1777 gnd 0.590664f
C4204 vdd.n1778 gnd 0.799748f
C4205 vdd.n1779 gnd 0.01023f
C4206 vdd.n1780 gnd 0.008234f
C4207 vdd.n1781 gnd 0.01023f
C4208 vdd.n1782 gnd 0.01023f
C4209 vdd.n1783 gnd 0.01023f
C4210 vdd.n1784 gnd 0.008234f
C4211 vdd.n1785 gnd 0.01023f
C4212 vdd.n1786 gnd 0.8677f
C4213 vdd.n1787 gnd 0.01023f
C4214 vdd.n1788 gnd 0.008234f
C4215 vdd.n1789 gnd 0.01023f
C4216 vdd.n1790 gnd 0.01023f
C4217 vdd.n1791 gnd 0.01023f
C4218 vdd.n1792 gnd 0.008234f
C4219 vdd.n1793 gnd 0.01023f
C4220 vdd.t217 gnd 0.522711f
C4221 vdd.n1794 gnd 0.757931f
C4222 vdd.n1795 gnd 0.01023f
C4223 vdd.n1796 gnd 0.008234f
C4224 vdd.n1797 gnd 0.01023f
C4225 vdd.n1798 gnd 0.01023f
C4226 vdd.n1799 gnd 0.01023f
C4227 vdd.n1800 gnd 0.008234f
C4228 vdd.n1801 gnd 0.01023f
C4229 vdd.n1802 gnd 0.580209f
C4230 vdd.n1803 gnd 0.01023f
C4231 vdd.n1804 gnd 0.008234f
C4232 vdd.n1805 gnd 0.01023f
C4233 vdd.n1806 gnd 0.01023f
C4234 vdd.n1807 gnd 0.01023f
C4235 vdd.n1808 gnd 0.008234f
C4236 vdd.n1809 gnd 0.01023f
C4237 vdd.n1810 gnd 0.747477f
C4238 vdd.n1811 gnd 0.642935f
C4239 vdd.n1812 gnd 0.01023f
C4240 vdd.n1813 gnd 0.008234f
C4241 vdd.n1814 gnd 0.007862f
C4242 vdd.n1815 gnd 0.005614f
C4243 vdd.n1816 gnd 0.00521f
C4244 vdd.n1817 gnd 0.002882f
C4245 vdd.n1818 gnd 0.006617f
C4246 vdd.n1819 gnd 0.002799f
C4247 vdd.n1820 gnd 0.002964f
C4248 vdd.n1821 gnd 0.00521f
C4249 vdd.n1822 gnd 0.002799f
C4250 vdd.n1823 gnd 0.006617f
C4251 vdd.n1824 gnd 0.002964f
C4252 vdd.n1825 gnd 0.00521f
C4253 vdd.n1826 gnd 0.002799f
C4254 vdd.n1827 gnd 0.004963f
C4255 vdd.n1828 gnd 0.004977f
C4256 vdd.t180 gnd 0.014216f
C4257 vdd.n1829 gnd 0.03163f
C4258 vdd.n1830 gnd 0.164609f
C4259 vdd.n1831 gnd 0.002799f
C4260 vdd.n1832 gnd 0.002964f
C4261 vdd.n1833 gnd 0.006617f
C4262 vdd.n1834 gnd 0.006617f
C4263 vdd.n1835 gnd 0.002964f
C4264 vdd.n1836 gnd 0.002799f
C4265 vdd.n1837 gnd 0.00521f
C4266 vdd.n1838 gnd 0.00521f
C4267 vdd.n1839 gnd 0.002799f
C4268 vdd.n1840 gnd 0.002964f
C4269 vdd.n1841 gnd 0.006617f
C4270 vdd.n1842 gnd 0.006617f
C4271 vdd.n1843 gnd 0.002964f
C4272 vdd.n1844 gnd 0.002799f
C4273 vdd.n1845 gnd 0.00521f
C4274 vdd.n1846 gnd 0.00521f
C4275 vdd.n1847 gnd 0.002799f
C4276 vdd.n1848 gnd 0.002964f
C4277 vdd.n1849 gnd 0.006617f
C4278 vdd.n1850 gnd 0.006617f
C4279 vdd.n1851 gnd 0.015644f
C4280 vdd.n1852 gnd 0.002882f
C4281 vdd.n1853 gnd 0.002799f
C4282 vdd.n1854 gnd 0.013465f
C4283 vdd.n1855 gnd 0.009401f
C4284 vdd.t204 gnd 0.032935f
C4285 vdd.t248 gnd 0.032935f
C4286 vdd.n1856 gnd 0.226349f
C4287 vdd.n1857 gnd 0.177989f
C4288 vdd.t221 gnd 0.032935f
C4289 vdd.t260 gnd 0.032935f
C4290 vdd.n1858 gnd 0.226349f
C4291 vdd.n1859 gnd 0.143636f
C4292 vdd.t195 gnd 0.032935f
C4293 vdd.t151 gnd 0.032935f
C4294 vdd.n1860 gnd 0.226349f
C4295 vdd.n1861 gnd 0.143636f
C4296 vdd.t213 gnd 0.032935f
C4297 vdd.t159 gnd 0.032935f
C4298 vdd.n1862 gnd 0.226349f
C4299 vdd.n1863 gnd 0.143636f
C4300 vdd.t252 gnd 0.032935f
C4301 vdd.t264 gnd 0.032935f
C4302 vdd.n1864 gnd 0.226349f
C4303 vdd.n1865 gnd 0.143636f
C4304 vdd.t232 gnd 0.032935f
C4305 vdd.t163 gnd 0.032935f
C4306 vdd.n1866 gnd 0.226349f
C4307 vdd.n1867 gnd 0.143636f
C4308 vdd.t222 gnd 0.032935f
C4309 vdd.t173 gnd 0.032935f
C4310 vdd.n1868 gnd 0.226349f
C4311 vdd.n1869 gnd 0.143636f
C4312 vdd.n1870 gnd 0.005614f
C4313 vdd.n1871 gnd 0.00521f
C4314 vdd.n1872 gnd 0.002882f
C4315 vdd.n1873 gnd 0.006617f
C4316 vdd.n1874 gnd 0.002799f
C4317 vdd.n1875 gnd 0.002964f
C4318 vdd.n1876 gnd 0.00521f
C4319 vdd.n1877 gnd 0.002799f
C4320 vdd.n1878 gnd 0.006617f
C4321 vdd.n1879 gnd 0.002964f
C4322 vdd.n1880 gnd 0.00521f
C4323 vdd.n1881 gnd 0.002799f
C4324 vdd.n1882 gnd 0.004963f
C4325 vdd.n1883 gnd 0.004977f
C4326 vdd.t198 gnd 0.014216f
C4327 vdd.n1884 gnd 0.03163f
C4328 vdd.n1885 gnd 0.164609f
C4329 vdd.n1886 gnd 0.002799f
C4330 vdd.n1887 gnd 0.002964f
C4331 vdd.n1888 gnd 0.006617f
C4332 vdd.n1889 gnd 0.006617f
C4333 vdd.n1890 gnd 0.002964f
C4334 vdd.n1891 gnd 0.002799f
C4335 vdd.n1892 gnd 0.00521f
C4336 vdd.n1893 gnd 0.00521f
C4337 vdd.n1894 gnd 0.002799f
C4338 vdd.n1895 gnd 0.002964f
C4339 vdd.n1896 gnd 0.006617f
C4340 vdd.n1897 gnd 0.006617f
C4341 vdd.n1898 gnd 0.002964f
C4342 vdd.n1899 gnd 0.002799f
C4343 vdd.n1900 gnd 0.00521f
C4344 vdd.n1901 gnd 0.00521f
C4345 vdd.n1902 gnd 0.002799f
C4346 vdd.n1903 gnd 0.002964f
C4347 vdd.n1904 gnd 0.006617f
C4348 vdd.n1905 gnd 0.006617f
C4349 vdd.n1906 gnd 0.015644f
C4350 vdd.n1907 gnd 0.002882f
C4351 vdd.n1908 gnd 0.002799f
C4352 vdd.n1909 gnd 0.013465f
C4353 vdd.n1910 gnd 0.009106f
C4354 vdd.n1911 gnd 0.106866f
C4355 vdd.n1912 gnd 0.005614f
C4356 vdd.n1913 gnd 0.00521f
C4357 vdd.n1914 gnd 0.002882f
C4358 vdd.n1915 gnd 0.006617f
C4359 vdd.n1916 gnd 0.002799f
C4360 vdd.n1917 gnd 0.002964f
C4361 vdd.n1918 gnd 0.00521f
C4362 vdd.n1919 gnd 0.002799f
C4363 vdd.n1920 gnd 0.006617f
C4364 vdd.n1921 gnd 0.002964f
C4365 vdd.n1922 gnd 0.00521f
C4366 vdd.n1923 gnd 0.002799f
C4367 vdd.n1924 gnd 0.004963f
C4368 vdd.n1925 gnd 0.004977f
C4369 vdd.t246 gnd 0.014216f
C4370 vdd.n1926 gnd 0.03163f
C4371 vdd.n1927 gnd 0.164609f
C4372 vdd.n1928 gnd 0.002799f
C4373 vdd.n1929 gnd 0.002964f
C4374 vdd.n1930 gnd 0.006617f
C4375 vdd.n1931 gnd 0.006617f
C4376 vdd.n1932 gnd 0.002964f
C4377 vdd.n1933 gnd 0.002799f
C4378 vdd.n1934 gnd 0.00521f
C4379 vdd.n1935 gnd 0.00521f
C4380 vdd.n1936 gnd 0.002799f
C4381 vdd.n1937 gnd 0.002964f
C4382 vdd.n1938 gnd 0.006617f
C4383 vdd.n1939 gnd 0.006617f
C4384 vdd.n1940 gnd 0.002964f
C4385 vdd.n1941 gnd 0.002799f
C4386 vdd.n1942 gnd 0.00521f
C4387 vdd.n1943 gnd 0.00521f
C4388 vdd.n1944 gnd 0.002799f
C4389 vdd.n1945 gnd 0.002964f
C4390 vdd.n1946 gnd 0.006617f
C4391 vdd.n1947 gnd 0.006617f
C4392 vdd.n1948 gnd 0.015644f
C4393 vdd.n1949 gnd 0.002882f
C4394 vdd.n1950 gnd 0.002799f
C4395 vdd.n1951 gnd 0.013465f
C4396 vdd.n1952 gnd 0.009401f
C4397 vdd.t208 gnd 0.032935f
C4398 vdd.t143 gnd 0.032935f
C4399 vdd.n1953 gnd 0.226349f
C4400 vdd.n1954 gnd 0.177989f
C4401 vdd.t257 gnd 0.032935f
C4402 vdd.t234 gnd 0.032935f
C4403 vdd.n1955 gnd 0.226349f
C4404 vdd.n1956 gnd 0.143636f
C4405 vdd.t228 gnd 0.032935f
C4406 vdd.t181 gnd 0.032935f
C4407 vdd.n1957 gnd 0.226349f
C4408 vdd.n1958 gnd 0.143636f
C4409 vdd.t175 gnd 0.032935f
C4410 vdd.t229 gnd 0.032935f
C4411 vdd.n1959 gnd 0.226349f
C4412 vdd.n1960 gnd 0.143636f
C4413 vdd.t218 gnd 0.032935f
C4414 vdd.t216 gnd 0.032935f
C4415 vdd.n1961 gnd 0.226349f
C4416 vdd.n1962 gnd 0.143636f
C4417 vdd.t171 gnd 0.032935f
C4418 vdd.t149 gnd 0.032935f
C4419 vdd.n1963 gnd 0.226349f
C4420 vdd.n1964 gnd 0.143636f
C4421 vdd.t141 gnd 0.032935f
C4422 vdd.t214 gnd 0.032935f
C4423 vdd.n1965 gnd 0.226349f
C4424 vdd.n1966 gnd 0.143636f
C4425 vdd.n1967 gnd 0.005614f
C4426 vdd.n1968 gnd 0.00521f
C4427 vdd.n1969 gnd 0.002882f
C4428 vdd.n1970 gnd 0.006617f
C4429 vdd.n1971 gnd 0.002799f
C4430 vdd.n1972 gnd 0.002964f
C4431 vdd.n1973 gnd 0.00521f
C4432 vdd.n1974 gnd 0.002799f
C4433 vdd.n1975 gnd 0.006617f
C4434 vdd.n1976 gnd 0.002964f
C4435 vdd.n1977 gnd 0.00521f
C4436 vdd.n1978 gnd 0.002799f
C4437 vdd.n1979 gnd 0.004963f
C4438 vdd.n1980 gnd 0.004977f
C4439 vdd.t145 gnd 0.014216f
C4440 vdd.n1981 gnd 0.03163f
C4441 vdd.n1982 gnd 0.164609f
C4442 vdd.n1983 gnd 0.002799f
C4443 vdd.n1984 gnd 0.002964f
C4444 vdd.n1985 gnd 0.006617f
C4445 vdd.n1986 gnd 0.006617f
C4446 vdd.n1987 gnd 0.002964f
C4447 vdd.n1988 gnd 0.002799f
C4448 vdd.n1989 gnd 0.00521f
C4449 vdd.n1990 gnd 0.00521f
C4450 vdd.n1991 gnd 0.002799f
C4451 vdd.n1992 gnd 0.002964f
C4452 vdd.n1993 gnd 0.006617f
C4453 vdd.n1994 gnd 0.006617f
C4454 vdd.n1995 gnd 0.002964f
C4455 vdd.n1996 gnd 0.002799f
C4456 vdd.n1997 gnd 0.00521f
C4457 vdd.n1998 gnd 0.00521f
C4458 vdd.n1999 gnd 0.002799f
C4459 vdd.n2000 gnd 0.002964f
C4460 vdd.n2001 gnd 0.006617f
C4461 vdd.n2002 gnd 0.006617f
C4462 vdd.n2003 gnd 0.015644f
C4463 vdd.n2004 gnd 0.002882f
C4464 vdd.n2005 gnd 0.002799f
C4465 vdd.n2006 gnd 0.013465f
C4466 vdd.n2007 gnd 0.009106f
C4467 vdd.n2008 gnd 0.063574f
C4468 vdd.n2009 gnd 0.229075f
C4469 vdd.n2010 gnd 0.005614f
C4470 vdd.n2011 gnd 0.00521f
C4471 vdd.n2012 gnd 0.002882f
C4472 vdd.n2013 gnd 0.006617f
C4473 vdd.n2014 gnd 0.002799f
C4474 vdd.n2015 gnd 0.002964f
C4475 vdd.n2016 gnd 0.00521f
C4476 vdd.n2017 gnd 0.002799f
C4477 vdd.n2018 gnd 0.006617f
C4478 vdd.n2019 gnd 0.002964f
C4479 vdd.n2020 gnd 0.00521f
C4480 vdd.n2021 gnd 0.002799f
C4481 vdd.n2022 gnd 0.004963f
C4482 vdd.n2023 gnd 0.004977f
C4483 vdd.t256 gnd 0.014216f
C4484 vdd.n2024 gnd 0.03163f
C4485 vdd.n2025 gnd 0.164609f
C4486 vdd.n2026 gnd 0.002799f
C4487 vdd.n2027 gnd 0.002964f
C4488 vdd.n2028 gnd 0.006617f
C4489 vdd.n2029 gnd 0.006617f
C4490 vdd.n2030 gnd 0.002964f
C4491 vdd.n2031 gnd 0.002799f
C4492 vdd.n2032 gnd 0.00521f
C4493 vdd.n2033 gnd 0.00521f
C4494 vdd.n2034 gnd 0.002799f
C4495 vdd.n2035 gnd 0.002964f
C4496 vdd.n2036 gnd 0.006617f
C4497 vdd.n2037 gnd 0.006617f
C4498 vdd.n2038 gnd 0.002964f
C4499 vdd.n2039 gnd 0.002799f
C4500 vdd.n2040 gnd 0.00521f
C4501 vdd.n2041 gnd 0.00521f
C4502 vdd.n2042 gnd 0.002799f
C4503 vdd.n2043 gnd 0.002964f
C4504 vdd.n2044 gnd 0.006617f
C4505 vdd.n2045 gnd 0.006617f
C4506 vdd.n2046 gnd 0.015644f
C4507 vdd.n2047 gnd 0.002882f
C4508 vdd.n2048 gnd 0.002799f
C4509 vdd.n2049 gnd 0.013465f
C4510 vdd.n2050 gnd 0.009401f
C4511 vdd.t219 gnd 0.032935f
C4512 vdd.t165 gnd 0.032935f
C4513 vdd.n2051 gnd 0.226349f
C4514 vdd.n2052 gnd 0.177989f
C4515 vdd.t265 gnd 0.032935f
C4516 vdd.t241 gnd 0.032935f
C4517 vdd.n2053 gnd 0.226349f
C4518 vdd.n2054 gnd 0.143636f
C4519 vdd.t239 gnd 0.032935f
C4520 vdd.t199 gnd 0.032935f
C4521 vdd.n2055 gnd 0.226349f
C4522 vdd.n2056 gnd 0.143636f
C4523 vdd.t192 gnd 0.032935f
C4524 vdd.t240 gnd 0.032935f
C4525 vdd.n2057 gnd 0.226349f
C4526 vdd.n2058 gnd 0.143636f
C4527 vdd.t227 gnd 0.032935f
C4528 vdd.t226 gnd 0.032935f
C4529 vdd.n2059 gnd 0.226349f
C4530 vdd.n2060 gnd 0.143636f
C4531 vdd.t191 gnd 0.032935f
C4532 vdd.t167 gnd 0.032935f
C4533 vdd.n2061 gnd 0.226349f
C4534 vdd.n2062 gnd 0.143636f
C4535 vdd.t164 gnd 0.032935f
C4536 vdd.t225 gnd 0.032935f
C4537 vdd.n2063 gnd 0.226349f
C4538 vdd.n2064 gnd 0.143636f
C4539 vdd.n2065 gnd 0.005614f
C4540 vdd.n2066 gnd 0.00521f
C4541 vdd.n2067 gnd 0.002882f
C4542 vdd.n2068 gnd 0.006617f
C4543 vdd.n2069 gnd 0.002799f
C4544 vdd.n2070 gnd 0.002964f
C4545 vdd.n2071 gnd 0.00521f
C4546 vdd.n2072 gnd 0.002799f
C4547 vdd.n2073 gnd 0.006617f
C4548 vdd.n2074 gnd 0.002964f
C4549 vdd.n2075 gnd 0.00521f
C4550 vdd.n2076 gnd 0.002799f
C4551 vdd.n2077 gnd 0.004963f
C4552 vdd.n2078 gnd 0.004977f
C4553 vdd.t166 gnd 0.014216f
C4554 vdd.n2079 gnd 0.03163f
C4555 vdd.n2080 gnd 0.164609f
C4556 vdd.n2081 gnd 0.002799f
C4557 vdd.n2082 gnd 0.002964f
C4558 vdd.n2083 gnd 0.006617f
C4559 vdd.n2084 gnd 0.006617f
C4560 vdd.n2085 gnd 0.002964f
C4561 vdd.n2086 gnd 0.002799f
C4562 vdd.n2087 gnd 0.00521f
C4563 vdd.n2088 gnd 0.00521f
C4564 vdd.n2089 gnd 0.002799f
C4565 vdd.n2090 gnd 0.002964f
C4566 vdd.n2091 gnd 0.006617f
C4567 vdd.n2092 gnd 0.006617f
C4568 vdd.n2093 gnd 0.002964f
C4569 vdd.n2094 gnd 0.002799f
C4570 vdd.n2095 gnd 0.00521f
C4571 vdd.n2096 gnd 0.00521f
C4572 vdd.n2097 gnd 0.002799f
C4573 vdd.n2098 gnd 0.002964f
C4574 vdd.n2099 gnd 0.006617f
C4575 vdd.n2100 gnd 0.006617f
C4576 vdd.n2101 gnd 0.015644f
C4577 vdd.n2102 gnd 0.002882f
C4578 vdd.n2103 gnd 0.002799f
C4579 vdd.n2104 gnd 0.013465f
C4580 vdd.n2105 gnd 0.009106f
C4581 vdd.n2106 gnd 0.063574f
C4582 vdd.n2107 gnd 0.256534f
C4583 vdd.n2108 gnd 2.57063f
C4584 vdd.n2109 gnd 0.603384f
C4585 vdd.n2110 gnd 0.007862f
C4586 vdd.n2111 gnd 0.01023f
C4587 vdd.n2112 gnd 0.008234f
C4588 vdd.n2113 gnd 0.01023f
C4589 vdd.n2114 gnd 0.820656f
C4590 vdd.n2115 gnd 0.01023f
C4591 vdd.n2116 gnd 0.008234f
C4592 vdd.n2117 gnd 0.01023f
C4593 vdd.n2118 gnd 0.01023f
C4594 vdd.n2119 gnd 0.01023f
C4595 vdd.n2120 gnd 0.008234f
C4596 vdd.n2121 gnd 0.01023f
C4597 vdd.t150 gnd 0.522711f
C4598 vdd.n2122 gnd 0.8677f
C4599 vdd.n2123 gnd 0.01023f
C4600 vdd.n2124 gnd 0.008234f
C4601 vdd.n2125 gnd 0.01023f
C4602 vdd.n2126 gnd 0.01023f
C4603 vdd.n2127 gnd 0.01023f
C4604 vdd.n2128 gnd 0.008234f
C4605 vdd.n2129 gnd 0.01023f
C4606 vdd.n2130 gnd 0.737023f
C4607 vdd.n2131 gnd 0.01023f
C4608 vdd.n2132 gnd 0.008234f
C4609 vdd.n2133 gnd 0.01023f
C4610 vdd.n2134 gnd 0.01023f
C4611 vdd.n2135 gnd 0.01023f
C4612 vdd.n2136 gnd 0.008234f
C4613 vdd.n2137 gnd 0.01023f
C4614 vdd.n2138 gnd 0.8677f
C4615 vdd.t233 gnd 0.522711f
C4616 vdd.n2139 gnd 0.559301f
C4617 vdd.n2140 gnd 0.01023f
C4618 vdd.n2141 gnd 0.008234f
C4619 vdd.n2142 gnd 0.01023f
C4620 vdd.n2143 gnd 0.01023f
C4621 vdd.n2144 gnd 0.01023f
C4622 vdd.n2145 gnd 0.008234f
C4623 vdd.n2146 gnd 0.01023f
C4624 vdd.n2147 gnd 0.663843f
C4625 vdd.n2148 gnd 0.01023f
C4626 vdd.n2149 gnd 0.008234f
C4627 vdd.n2150 gnd 0.01023f
C4628 vdd.n2151 gnd 0.01023f
C4629 vdd.n2152 gnd 0.01023f
C4630 vdd.n2153 gnd 0.008234f
C4631 vdd.n2154 gnd 0.01023f
C4632 vdd.n2155 gnd 0.548847f
C4633 vdd.n2156 gnd 0.841565f
C4634 vdd.n2157 gnd 0.01023f
C4635 vdd.n2158 gnd 0.008234f
C4636 vdd.n2159 gnd 0.01023f
C4637 vdd.n2160 gnd 0.01023f
C4638 vdd.n2161 gnd 0.01023f
C4639 vdd.n2162 gnd 0.008234f
C4640 vdd.n2163 gnd 0.01023f
C4641 vdd.n2164 gnd 1.01929f
C4642 vdd.n2165 gnd 0.01023f
C4643 vdd.n2166 gnd 0.008234f
C4644 vdd.n2167 gnd 0.01023f
C4645 vdd.n2168 gnd 0.01023f
C4646 vdd.n2169 gnd 0.023295f
C4647 vdd.n2170 gnd 0.01023f
C4648 vdd.n2171 gnd 0.01023f
C4649 vdd.n2172 gnd 0.008234f
C4650 vdd.n2173 gnd 0.01023f
C4651 vdd.t63 gnd 0.522711f
C4652 vdd.n2174 gnd 0.987924f
C4653 vdd.n2175 gnd 0.01023f
C4654 vdd.n2176 gnd 0.008234f
C4655 vdd.n2177 gnd 0.01023f
C4656 vdd.n2178 gnd 0.01023f
C4657 vdd.n2179 gnd 0.023295f
C4658 vdd.n2180 gnd 0.006834f
C4659 vdd.n2181 gnd 0.023295f
C4660 vdd.n2182 gnd 1.37996f
C4661 vdd.n2183 gnd 0.023295f
C4662 vdd.n2184 gnd 0.023454f
C4663 vdd.n2185 gnd 0.003911f
C4664 vdd.t65 gnd 0.125851f
C4665 vdd.t64 gnd 0.134501f
C4666 vdd.t62 gnd 0.164361f
C4667 vdd.n2186 gnd 0.210687f
C4668 vdd.n2187 gnd 0.177015f
C4669 vdd.n2188 gnd 0.01268f
C4670 vdd.n2189 gnd 0.004323f
C4671 vdd.n2190 gnd 0.008798f
C4672 vdd.n2191 gnd 0.773622f
C4673 vdd.n2193 gnd 0.008234f
C4674 vdd.n2194 gnd 0.008234f
C4675 vdd.n2195 gnd 0.01023f
C4676 vdd.n2197 gnd 0.01023f
C4677 vdd.n2198 gnd 0.01023f
C4678 vdd.n2199 gnd 0.008234f
C4679 vdd.n2200 gnd 0.008234f
C4680 vdd.n2201 gnd 0.008234f
C4681 vdd.n2202 gnd 0.01023f
C4682 vdd.n2204 gnd 0.01023f
C4683 vdd.n2205 gnd 0.01023f
C4684 vdd.n2206 gnd 0.008234f
C4685 vdd.n2207 gnd 0.008234f
C4686 vdd.n2208 gnd 0.008234f
C4687 vdd.n2209 gnd 0.01023f
C4688 vdd.n2211 gnd 0.01023f
C4689 vdd.n2212 gnd 0.01023f
C4690 vdd.n2213 gnd 0.008234f
C4691 vdd.n2214 gnd 0.008234f
C4692 vdd.n2215 gnd 0.008234f
C4693 vdd.n2216 gnd 0.01023f
C4694 vdd.n2218 gnd 0.01023f
C4695 vdd.n2219 gnd 0.01023f
C4696 vdd.n2220 gnd 0.008234f
C4697 vdd.n2221 gnd 0.01023f
C4698 vdd.n2222 gnd 0.01023f
C4699 vdd.n2223 gnd 0.01023f
C4700 vdd.n2224 gnd 0.016797f
C4701 vdd.n2225 gnd 0.005599f
C4702 vdd.n2226 gnd 0.008234f
C4703 vdd.n2227 gnd 0.01023f
C4704 vdd.n2229 gnd 0.01023f
C4705 vdd.n2230 gnd 0.01023f
C4706 vdd.n2231 gnd 0.008234f
C4707 vdd.n2232 gnd 0.008234f
C4708 vdd.n2233 gnd 0.008234f
C4709 vdd.n2234 gnd 0.01023f
C4710 vdd.n2236 gnd 0.01023f
C4711 vdd.n2237 gnd 0.01023f
C4712 vdd.n2238 gnd 0.008234f
C4713 vdd.n2239 gnd 0.008234f
C4714 vdd.n2240 gnd 0.008234f
C4715 vdd.n2241 gnd 0.01023f
C4716 vdd.n2243 gnd 0.01023f
C4717 vdd.n2244 gnd 0.01023f
C4718 vdd.n2245 gnd 0.008234f
C4719 vdd.n2246 gnd 0.008234f
C4720 vdd.n2247 gnd 0.008234f
C4721 vdd.n2248 gnd 0.01023f
C4722 vdd.n2250 gnd 0.01023f
C4723 vdd.n2251 gnd 0.01023f
C4724 vdd.n2252 gnd 0.008234f
C4725 vdd.n2253 gnd 0.008234f
C4726 vdd.n2254 gnd 0.008234f
C4727 vdd.n2255 gnd 0.01023f
C4728 vdd.n2257 gnd 0.01023f
C4729 vdd.n2258 gnd 0.01023f
C4730 vdd.n2259 gnd 0.008234f
C4731 vdd.n2260 gnd 0.01023f
C4732 vdd.n2261 gnd 0.01023f
C4733 vdd.n2262 gnd 0.01023f
C4734 vdd.n2263 gnd 0.016797f
C4735 vdd.n2264 gnd 0.006875f
C4736 vdd.n2265 gnd 0.008234f
C4737 vdd.n2266 gnd 0.01023f
C4738 vdd.n2268 gnd 0.01023f
C4739 vdd.n2269 gnd 0.01023f
C4740 vdd.n2270 gnd 0.008234f
C4741 vdd.n2271 gnd 0.008234f
C4742 vdd.n2272 gnd 0.008234f
C4743 vdd.n2273 gnd 0.01023f
C4744 vdd.n2275 gnd 0.01023f
C4745 vdd.n2276 gnd 0.01023f
C4746 vdd.n2277 gnd 0.008234f
C4747 vdd.n2278 gnd 0.008234f
C4748 vdd.n2279 gnd 0.008234f
C4749 vdd.n2280 gnd 0.01023f
C4750 vdd.n2282 gnd 0.01023f
C4751 vdd.n2283 gnd 0.01023f
C4752 vdd.n2284 gnd 0.008234f
C4753 vdd.n2285 gnd 0.008234f
C4754 vdd.n2286 gnd 0.008234f
C4755 vdd.n2287 gnd 0.01023f
C4756 vdd.n2289 gnd 0.01023f
C4757 vdd.n2290 gnd 0.008234f
C4758 vdd.n2291 gnd 0.008234f
C4759 vdd.n2292 gnd 0.01023f
C4760 vdd.n2294 gnd 0.01023f
C4761 vdd.n2295 gnd 0.01023f
C4762 vdd.n2296 gnd 0.008234f
C4763 vdd.n2297 gnd 0.008798f
C4764 vdd.n2298 gnd 0.773622f
C4765 vdd.n2299 gnd 0.02788f
C4766 vdd.n2300 gnd 0.006956f
C4767 vdd.n2301 gnd 0.006956f
C4768 vdd.n2302 gnd 0.006956f
C4769 vdd.n2303 gnd 0.006956f
C4770 vdd.n2304 gnd 0.006956f
C4771 vdd.n2305 gnd 0.006956f
C4772 vdd.n2306 gnd 0.006956f
C4773 vdd.n2307 gnd 0.006956f
C4774 vdd.n2308 gnd 0.006956f
C4775 vdd.n2309 gnd 0.006956f
C4776 vdd.n2310 gnd 0.006956f
C4777 vdd.n2311 gnd 0.006956f
C4778 vdd.n2312 gnd 0.006956f
C4779 vdd.n2313 gnd 0.006956f
C4780 vdd.n2314 gnd 0.006956f
C4781 vdd.n2315 gnd 0.006956f
C4782 vdd.n2316 gnd 0.006956f
C4783 vdd.n2317 gnd 0.006956f
C4784 vdd.n2318 gnd 0.006956f
C4785 vdd.n2319 gnd 0.006956f
C4786 vdd.n2320 gnd 0.006956f
C4787 vdd.n2321 gnd 0.006956f
C4788 vdd.n2322 gnd 0.006956f
C4789 vdd.n2323 gnd 0.006956f
C4790 vdd.n2324 gnd 0.006956f
C4791 vdd.n2325 gnd 0.006956f
C4792 vdd.n2326 gnd 0.006956f
C4793 vdd.n2327 gnd 0.006956f
C4794 vdd.n2328 gnd 0.006956f
C4795 vdd.n2329 gnd 0.006956f
C4796 vdd.n2330 gnd 0.006956f
C4797 vdd.n2331 gnd 0.01627f
C4798 vdd.n2332 gnd 0.01627f
C4799 vdd.n2334 gnd 8.91745f
C4800 vdd.n2336 gnd 0.01627f
C4801 vdd.n2337 gnd 0.01627f
C4802 vdd.n2338 gnd 0.015237f
C4803 vdd.n2339 gnd 0.006956f
C4804 vdd.n2340 gnd 0.006956f
C4805 vdd.n2341 gnd 0.710887f
C4806 vdd.n2342 gnd 0.006956f
C4807 vdd.n2343 gnd 0.006956f
C4808 vdd.n2344 gnd 0.006956f
C4809 vdd.n2345 gnd 0.006956f
C4810 vdd.n2346 gnd 0.006956f
C4811 vdd.n2347 gnd 0.601118f
C4812 vdd.n2348 gnd 0.006956f
C4813 vdd.n2349 gnd 0.006956f
C4814 vdd.n2350 gnd 0.006956f
C4815 vdd.n2351 gnd 0.006956f
C4816 vdd.n2352 gnd 0.006956f
C4817 vdd.n2353 gnd 0.710887f
C4818 vdd.n2354 gnd 0.006956f
C4819 vdd.n2355 gnd 0.006956f
C4820 vdd.n2356 gnd 0.006956f
C4821 vdd.n2357 gnd 0.006956f
C4822 vdd.n2358 gnd 0.006956f
C4823 vdd.n2359 gnd 0.695206f
C4824 vdd.n2360 gnd 0.006956f
C4825 vdd.n2361 gnd 0.006956f
C4826 vdd.n2362 gnd 0.006956f
C4827 vdd.n2363 gnd 0.006956f
C4828 vdd.n2364 gnd 0.006956f
C4829 vdd.n2365 gnd 0.710887f
C4830 vdd.n2366 gnd 0.006956f
C4831 vdd.n2367 gnd 0.006956f
C4832 vdd.n2368 gnd 0.006956f
C4833 vdd.n2369 gnd 0.006956f
C4834 vdd.n2370 gnd 0.006956f
C4835 vdd.n2371 gnd 0.569755f
C4836 vdd.n2372 gnd 0.006956f
C4837 vdd.n2373 gnd 0.006956f
C4838 vdd.n2374 gnd 0.005933f
C4839 vdd.n2375 gnd 0.020151f
C4840 vdd.n2376 gnd 0.004501f
C4841 vdd.n2377 gnd 0.006956f
C4842 vdd.n2378 gnd 0.412942f
C4843 vdd.n2379 gnd 0.006956f
C4844 vdd.n2380 gnd 0.006956f
C4845 vdd.n2381 gnd 0.006956f
C4846 vdd.n2382 gnd 0.006956f
C4847 vdd.n2383 gnd 0.006956f
C4848 vdd.n2384 gnd 0.454759f
C4849 vdd.n2385 gnd 0.006956f
C4850 vdd.n2386 gnd 0.006956f
C4851 vdd.n2387 gnd 0.006956f
C4852 vdd.n2388 gnd 0.006956f
C4853 vdd.n2389 gnd 0.006956f
C4854 vdd.n2390 gnd 0.611572f
C4855 vdd.n2391 gnd 0.006956f
C4856 vdd.n2392 gnd 0.006956f
C4857 vdd.n2393 gnd 0.006956f
C4858 vdd.n2394 gnd 0.006956f
C4859 vdd.n2395 gnd 0.006956f
C4860 vdd.n2396 gnd 0.585436f
C4861 vdd.n2397 gnd 0.006956f
C4862 vdd.n2398 gnd 0.006956f
C4863 vdd.n2399 gnd 0.006956f
C4864 vdd.n2400 gnd 0.006956f
C4865 vdd.n2401 gnd 0.006956f
C4866 vdd.n2402 gnd 0.428623f
C4867 vdd.n2403 gnd 0.006956f
C4868 vdd.n2404 gnd 0.006956f
C4869 vdd.n2405 gnd 0.006956f
C4870 vdd.n2406 gnd 0.006956f
C4871 vdd.n2407 gnd 0.006956f
C4872 vdd.n2408 gnd 0.224766f
C4873 vdd.n2409 gnd 0.006956f
C4874 vdd.n2410 gnd 0.006956f
C4875 vdd.n2411 gnd 0.006956f
C4876 vdd.n2412 gnd 0.006956f
C4877 vdd.n2413 gnd 0.006956f
C4878 vdd.n2414 gnd 0.371125f
C4879 vdd.n2415 gnd 0.006956f
C4880 vdd.n2416 gnd 0.006956f
C4881 vdd.n2417 gnd 0.006956f
C4882 vdd.n2418 gnd 0.006956f
C4883 vdd.n2419 gnd 0.006956f
C4884 vdd.n2420 gnd 0.710887f
C4885 vdd.n2421 gnd 0.006956f
C4886 vdd.n2422 gnd 0.006956f
C4887 vdd.n2423 gnd 0.006956f
C4888 vdd.n2424 gnd 0.006956f
C4889 vdd.n2425 gnd 0.006956f
C4890 vdd.n2426 gnd 0.006956f
C4891 vdd.n2427 gnd 0.006956f
C4892 vdd.n2428 gnd 0.533165f
C4893 vdd.n2429 gnd 0.006956f
C4894 vdd.n2430 gnd 0.006956f
C4895 vdd.n2431 gnd 0.006956f
C4896 vdd.n2432 gnd 0.006956f
C4897 vdd.n2433 gnd 0.006956f
C4898 vdd.n2434 gnd 0.006956f
C4899 vdd.n2435 gnd 0.444304f
C4900 vdd.n2436 gnd 0.006956f
C4901 vdd.n2437 gnd 0.006956f
C4902 vdd.n2438 gnd 0.006956f
C4903 vdd.n2439 gnd 0.016101f
C4904 vdd.n2440 gnd 0.015406f
C4905 vdd.n2441 gnd 0.006956f
C4906 vdd.n2442 gnd 0.006956f
C4907 vdd.n2443 gnd 0.005371f
C4908 vdd.n2444 gnd 0.006956f
C4909 vdd.n2445 gnd 0.006956f
C4910 vdd.n2446 gnd 0.005064f
C4911 vdd.n2447 gnd 0.006956f
C4912 vdd.n2448 gnd 0.006956f
C4913 vdd.n2449 gnd 0.006956f
C4914 vdd.n2450 gnd 0.006956f
C4915 vdd.n2451 gnd 0.006956f
C4916 vdd.n2452 gnd 0.006956f
C4917 vdd.n2453 gnd 0.006956f
C4918 vdd.n2454 gnd 0.006956f
C4919 vdd.n2455 gnd 0.006956f
C4920 vdd.n2456 gnd 0.006956f
C4921 vdd.n2457 gnd 0.006956f
C4922 vdd.n2458 gnd 0.006956f
C4923 vdd.n2459 gnd 0.006956f
C4924 vdd.n2460 gnd 0.006956f
C4925 vdd.n2461 gnd 0.006956f
C4926 vdd.n2462 gnd 0.006956f
C4927 vdd.n2463 gnd 0.006956f
C4928 vdd.n2464 gnd 0.006956f
C4929 vdd.n2465 gnd 0.006956f
C4930 vdd.n2466 gnd 0.006956f
C4931 vdd.n2467 gnd 0.006956f
C4932 vdd.n2468 gnd 0.006956f
C4933 vdd.n2469 gnd 0.006956f
C4934 vdd.n2470 gnd 0.006956f
C4935 vdd.n2471 gnd 0.006956f
C4936 vdd.n2472 gnd 0.006956f
C4937 vdd.n2473 gnd 0.006956f
C4938 vdd.n2474 gnd 0.006956f
C4939 vdd.n2475 gnd 0.006956f
C4940 vdd.n2476 gnd 0.006956f
C4941 vdd.n2477 gnd 0.006956f
C4942 vdd.n2478 gnd 0.006956f
C4943 vdd.n2479 gnd 0.006956f
C4944 vdd.n2480 gnd 0.006956f
C4945 vdd.n2481 gnd 0.006956f
C4946 vdd.n2482 gnd 0.006956f
C4947 vdd.n2483 gnd 0.006956f
C4948 vdd.n2484 gnd 0.006956f
C4949 vdd.n2485 gnd 0.006956f
C4950 vdd.n2486 gnd 0.006956f
C4951 vdd.n2487 gnd 0.006956f
C4952 vdd.n2488 gnd 0.006956f
C4953 vdd.n2489 gnd 0.006956f
C4954 vdd.n2490 gnd 0.006956f
C4955 vdd.n2491 gnd 0.006956f
C4956 vdd.n2492 gnd 0.006956f
C4957 vdd.n2493 gnd 0.006956f
C4958 vdd.n2494 gnd 0.006956f
C4959 vdd.n2495 gnd 0.006956f
C4960 vdd.n2496 gnd 0.006956f
C4961 vdd.n2497 gnd 0.006956f
C4962 vdd.n2498 gnd 0.006956f
C4963 vdd.n2499 gnd 0.006956f
C4964 vdd.n2500 gnd 0.006956f
C4965 vdd.n2501 gnd 0.006956f
C4966 vdd.n2502 gnd 0.006956f
C4967 vdd.n2503 gnd 0.006956f
C4968 vdd.n2504 gnd 0.006956f
C4969 vdd.n2505 gnd 0.006956f
C4970 vdd.n2506 gnd 0.006956f
C4971 vdd.n2507 gnd 0.01627f
C4972 vdd.n2508 gnd 0.015237f
C4973 vdd.n2509 gnd 0.015237f
C4974 vdd.n2510 gnd 0.846792f
C4975 vdd.n2511 gnd 0.015237f
C4976 vdd.n2512 gnd 0.01627f
C4977 vdd.n2513 gnd 0.015406f
C4978 vdd.n2514 gnd 0.006956f
C4979 vdd.n2515 gnd 0.006956f
C4980 vdd.n2516 gnd 0.006956f
C4981 vdd.n2517 gnd 0.005371f
C4982 vdd.n2518 gnd 0.009941f
C4983 vdd.n2519 gnd 0.005064f
C4984 vdd.n2520 gnd 0.006956f
C4985 vdd.n2521 gnd 0.006956f
C4986 vdd.n2522 gnd 0.006956f
C4987 vdd.n2523 gnd 0.006956f
C4988 vdd.n2524 gnd 0.006956f
C4989 vdd.n2525 gnd 0.006956f
C4990 vdd.n2526 gnd 0.006956f
C4991 vdd.n2527 gnd 0.006956f
C4992 vdd.n2528 gnd 0.006956f
C4993 vdd.n2529 gnd 0.006956f
C4994 vdd.n2530 gnd 0.006956f
C4995 vdd.n2531 gnd 0.006956f
C4996 vdd.n2532 gnd 0.006956f
C4997 vdd.n2533 gnd 0.006956f
C4998 vdd.n2534 gnd 0.006956f
C4999 vdd.n2535 gnd 0.006956f
C5000 vdd.n2536 gnd 0.006956f
C5001 vdd.n2537 gnd 0.006956f
C5002 vdd.n2538 gnd 0.006956f
C5003 vdd.n2539 gnd 0.006956f
C5004 vdd.n2540 gnd 0.006956f
C5005 vdd.n2541 gnd 0.006956f
C5006 vdd.n2542 gnd 0.006956f
C5007 vdd.n2543 gnd 0.006956f
C5008 vdd.n2544 gnd 0.006956f
C5009 vdd.n2545 gnd 0.006956f
C5010 vdd.n2546 gnd 0.006956f
C5011 vdd.n2547 gnd 0.006956f
C5012 vdd.n2548 gnd 0.006956f
C5013 vdd.n2549 gnd 0.006956f
C5014 vdd.n2550 gnd 0.006956f
C5015 vdd.n2551 gnd 0.006956f
C5016 vdd.n2552 gnd 0.006956f
C5017 vdd.n2553 gnd 0.006956f
C5018 vdd.n2554 gnd 0.006956f
C5019 vdd.n2555 gnd 0.006956f
C5020 vdd.n2556 gnd 0.006956f
C5021 vdd.n2557 gnd 0.006956f
C5022 vdd.n2558 gnd 0.006956f
C5023 vdd.n2559 gnd 0.006956f
C5024 vdd.n2560 gnd 0.006956f
C5025 vdd.n2561 gnd 0.006956f
C5026 vdd.n2562 gnd 0.006956f
C5027 vdd.n2563 gnd 0.006956f
C5028 vdd.n2564 gnd 0.006956f
C5029 vdd.n2565 gnd 0.006956f
C5030 vdd.n2566 gnd 0.006956f
C5031 vdd.n2567 gnd 0.006956f
C5032 vdd.n2568 gnd 0.006956f
C5033 vdd.n2569 gnd 0.006956f
C5034 vdd.n2570 gnd 0.006956f
C5035 vdd.n2571 gnd 0.006956f
C5036 vdd.n2572 gnd 0.006956f
C5037 vdd.n2573 gnd 0.006956f
C5038 vdd.n2574 gnd 0.006956f
C5039 vdd.n2575 gnd 0.006956f
C5040 vdd.n2576 gnd 0.006956f
C5041 vdd.n2577 gnd 0.006956f
C5042 vdd.n2578 gnd 0.006956f
C5043 vdd.n2579 gnd 0.006956f
C5044 vdd.n2580 gnd 0.01627f
C5045 vdd.n2581 gnd 0.01627f
C5046 vdd.n2582 gnd 0.8677f
C5047 vdd.t26 gnd 3.084f
C5048 vdd.t14 gnd 3.084f
C5049 vdd.n2615 gnd 0.01627f
C5050 vdd.t17 gnd 0.648162f
C5051 vdd.n2616 gnd 0.006956f
C5052 vdd.n2617 gnd 0.006956f
C5053 vdd.t102 gnd 0.281098f
C5054 vdd.t103 gnd 0.287738f
C5055 vdd.t100 gnd 0.183511f
C5056 vdd.n2618 gnd 0.099178f
C5057 vdd.n2619 gnd 0.056257f
C5058 vdd.n2620 gnd 0.006956f
C5059 vdd.t112 gnd 0.281098f
C5060 vdd.t113 gnd 0.287738f
C5061 vdd.t111 gnd 0.183511f
C5062 vdd.n2621 gnd 0.099178f
C5063 vdd.n2622 gnd 0.056257f
C5064 vdd.n2623 gnd 0.009941f
C5065 vdd.n2624 gnd 0.006956f
C5066 vdd.n2625 gnd 0.006956f
C5067 vdd.n2626 gnd 0.006956f
C5068 vdd.n2627 gnd 0.006956f
C5069 vdd.n2628 gnd 0.006956f
C5070 vdd.n2629 gnd 0.006956f
C5071 vdd.n2630 gnd 0.006956f
C5072 vdd.n2631 gnd 0.006956f
C5073 vdd.n2632 gnd 0.006956f
C5074 vdd.n2633 gnd 0.006956f
C5075 vdd.n2634 gnd 0.006956f
C5076 vdd.n2635 gnd 0.006956f
C5077 vdd.n2636 gnd 0.006956f
C5078 vdd.n2637 gnd 0.006956f
C5079 vdd.n2638 gnd 0.006956f
C5080 vdd.n2639 gnd 0.006956f
C5081 vdd.n2640 gnd 0.006956f
C5082 vdd.n2641 gnd 0.006956f
C5083 vdd.n2642 gnd 0.006956f
C5084 vdd.n2643 gnd 0.006956f
C5085 vdd.n2644 gnd 0.006956f
C5086 vdd.n2645 gnd 0.006956f
C5087 vdd.n2646 gnd 0.006956f
C5088 vdd.n2647 gnd 0.006956f
C5089 vdd.n2648 gnd 0.006956f
C5090 vdd.n2649 gnd 0.006956f
C5091 vdd.n2650 gnd 0.006956f
C5092 vdd.n2651 gnd 0.006956f
C5093 vdd.n2652 gnd 0.006956f
C5094 vdd.n2653 gnd 0.006956f
C5095 vdd.n2654 gnd 0.006956f
C5096 vdd.n2655 gnd 0.006956f
C5097 vdd.n2656 gnd 0.006956f
C5098 vdd.n2657 gnd 0.006956f
C5099 vdd.n2658 gnd 0.006956f
C5100 vdd.n2659 gnd 0.006956f
C5101 vdd.n2660 gnd 0.006956f
C5102 vdd.n2661 gnd 0.006956f
C5103 vdd.n2662 gnd 0.006956f
C5104 vdd.n2663 gnd 0.006956f
C5105 vdd.n2664 gnd 0.006956f
C5106 vdd.n2665 gnd 0.006956f
C5107 vdd.n2666 gnd 0.006956f
C5108 vdd.n2667 gnd 0.006956f
C5109 vdd.n2668 gnd 0.006956f
C5110 vdd.n2669 gnd 0.006956f
C5111 vdd.n2670 gnd 0.006956f
C5112 vdd.n2671 gnd 0.006956f
C5113 vdd.n2672 gnd 0.006956f
C5114 vdd.n2673 gnd 0.006956f
C5115 vdd.n2674 gnd 0.006956f
C5116 vdd.n2675 gnd 0.006956f
C5117 vdd.n2676 gnd 0.006956f
C5118 vdd.n2677 gnd 0.006956f
C5119 vdd.n2678 gnd 0.006956f
C5120 vdd.n2679 gnd 0.006956f
C5121 vdd.n2680 gnd 0.006956f
C5122 vdd.n2681 gnd 0.006956f
C5123 vdd.n2682 gnd 0.005064f
C5124 vdd.n2683 gnd 0.006956f
C5125 vdd.n2684 gnd 0.006956f
C5126 vdd.n2685 gnd 0.005371f
C5127 vdd.n2686 gnd 0.006956f
C5128 vdd.n2687 gnd 0.006956f
C5129 vdd.n2688 gnd 0.01627f
C5130 vdd.n2689 gnd 0.015237f
C5131 vdd.n2690 gnd 0.015237f
C5132 vdd.n2691 gnd 0.006956f
C5133 vdd.n2692 gnd 0.006956f
C5134 vdd.n2693 gnd 0.006956f
C5135 vdd.n2694 gnd 0.006956f
C5136 vdd.n2695 gnd 0.006956f
C5137 vdd.n2696 gnd 0.006956f
C5138 vdd.n2697 gnd 0.006956f
C5139 vdd.n2698 gnd 0.006956f
C5140 vdd.n2699 gnd 0.006956f
C5141 vdd.n2700 gnd 0.006956f
C5142 vdd.n2701 gnd 0.006956f
C5143 vdd.n2702 gnd 0.006956f
C5144 vdd.n2703 gnd 0.006956f
C5145 vdd.n2704 gnd 0.006956f
C5146 vdd.n2705 gnd 0.006956f
C5147 vdd.n2706 gnd 0.006956f
C5148 vdd.n2707 gnd 0.006956f
C5149 vdd.n2708 gnd 0.006956f
C5150 vdd.n2709 gnd 0.006956f
C5151 vdd.n2710 gnd 0.006956f
C5152 vdd.n2711 gnd 0.006956f
C5153 vdd.n2712 gnd 0.006956f
C5154 vdd.n2713 gnd 0.006956f
C5155 vdd.n2714 gnd 0.006956f
C5156 vdd.n2715 gnd 0.006956f
C5157 vdd.n2716 gnd 0.006956f
C5158 vdd.n2717 gnd 0.006956f
C5159 vdd.n2718 gnd 0.006956f
C5160 vdd.n2719 gnd 0.006956f
C5161 vdd.n2720 gnd 0.006956f
C5162 vdd.n2721 gnd 0.006956f
C5163 vdd.n2722 gnd 0.006956f
C5164 vdd.n2723 gnd 0.006956f
C5165 vdd.n2724 gnd 0.006956f
C5166 vdd.n2725 gnd 0.006956f
C5167 vdd.n2726 gnd 0.006956f
C5168 vdd.n2727 gnd 0.006956f
C5169 vdd.n2728 gnd 0.006956f
C5170 vdd.n2729 gnd 0.006956f
C5171 vdd.n2730 gnd 0.006956f
C5172 vdd.n2731 gnd 0.006956f
C5173 vdd.n2732 gnd 0.006956f
C5174 vdd.n2733 gnd 0.006956f
C5175 vdd.n2734 gnd 0.006956f
C5176 vdd.n2735 gnd 0.006956f
C5177 vdd.n2736 gnd 0.006956f
C5178 vdd.n2737 gnd 0.006956f
C5179 vdd.n2738 gnd 0.006956f
C5180 vdd.n2739 gnd 0.006956f
C5181 vdd.n2740 gnd 0.006956f
C5182 vdd.n2741 gnd 0.006956f
C5183 vdd.n2742 gnd 0.006956f
C5184 vdd.n2743 gnd 0.006956f
C5185 vdd.n2744 gnd 0.006956f
C5186 vdd.n2745 gnd 0.006956f
C5187 vdd.n2746 gnd 0.006956f
C5188 vdd.n2747 gnd 0.006956f
C5189 vdd.n2748 gnd 0.006956f
C5190 vdd.n2749 gnd 0.006956f
C5191 vdd.n2750 gnd 0.006956f
C5192 vdd.n2751 gnd 0.006956f
C5193 vdd.n2752 gnd 0.006956f
C5194 vdd.n2753 gnd 0.006956f
C5195 vdd.n2754 gnd 0.006956f
C5196 vdd.n2755 gnd 0.006956f
C5197 vdd.n2756 gnd 0.006956f
C5198 vdd.n2757 gnd 0.006956f
C5199 vdd.n2758 gnd 0.006956f
C5200 vdd.n2759 gnd 0.006956f
C5201 vdd.n2760 gnd 0.006956f
C5202 vdd.n2761 gnd 0.006956f
C5203 vdd.n2762 gnd 0.006956f
C5204 vdd.n2763 gnd 0.006956f
C5205 vdd.n2764 gnd 0.224766f
C5206 vdd.n2765 gnd 0.006956f
C5207 vdd.n2766 gnd 0.006956f
C5208 vdd.n2767 gnd 0.006956f
C5209 vdd.n2768 gnd 0.006956f
C5210 vdd.n2769 gnd 0.006956f
C5211 vdd.n2770 gnd 0.006956f
C5212 vdd.n2771 gnd 0.006956f
C5213 vdd.n2772 gnd 0.006956f
C5214 vdd.n2773 gnd 0.006956f
C5215 vdd.n2774 gnd 0.006956f
C5216 vdd.n2775 gnd 0.006956f
C5217 vdd.n2776 gnd 0.006956f
C5218 vdd.n2777 gnd 0.006956f
C5219 vdd.n2778 gnd 0.006956f
C5220 vdd.n2779 gnd 0.444304f
C5221 vdd.n2780 gnd 0.006956f
C5222 vdd.n2781 gnd 0.006956f
C5223 vdd.n2782 gnd 0.006956f
C5224 vdd.n2783 gnd 0.015237f
C5225 vdd.n2784 gnd 0.015237f
C5226 vdd.n2785 gnd 0.01627f
C5227 vdd.n2786 gnd 0.01627f
C5228 vdd.n2787 gnd 0.006956f
C5229 vdd.n2788 gnd 0.006956f
C5230 vdd.n2789 gnd 0.006956f
C5231 vdd.n2790 gnd 0.005371f
C5232 vdd.n2791 gnd 0.009941f
C5233 vdd.n2792 gnd 0.005064f
C5234 vdd.n2793 gnd 0.006956f
C5235 vdd.n2794 gnd 0.006956f
C5236 vdd.n2795 gnd 0.006956f
C5237 vdd.n2796 gnd 0.006956f
C5238 vdd.n2797 gnd 0.006956f
C5239 vdd.n2798 gnd 0.006956f
C5240 vdd.n2799 gnd 0.006956f
C5241 vdd.n2800 gnd 0.006956f
C5242 vdd.n2801 gnd 0.006956f
C5243 vdd.n2802 gnd 0.006956f
C5244 vdd.n2803 gnd 0.006956f
C5245 vdd.n2804 gnd 0.006956f
C5246 vdd.n2805 gnd 0.006956f
C5247 vdd.n2806 gnd 0.006956f
C5248 vdd.n2807 gnd 0.006956f
C5249 vdd.n2808 gnd 0.006956f
C5250 vdd.n2809 gnd 0.006956f
C5251 vdd.n2810 gnd 0.006956f
C5252 vdd.n2811 gnd 0.006956f
C5253 vdd.n2812 gnd 0.006956f
C5254 vdd.n2813 gnd 0.006956f
C5255 vdd.n2814 gnd 0.006956f
C5256 vdd.n2815 gnd 0.006956f
C5257 vdd.n2816 gnd 0.006956f
C5258 vdd.n2817 gnd 0.006956f
C5259 vdd.n2818 gnd 0.006956f
C5260 vdd.n2819 gnd 0.006956f
C5261 vdd.n2820 gnd 0.006956f
C5262 vdd.n2821 gnd 0.006956f
C5263 vdd.n2822 gnd 0.006956f
C5264 vdd.n2823 gnd 0.006956f
C5265 vdd.n2824 gnd 0.006956f
C5266 vdd.n2825 gnd 0.006956f
C5267 vdd.n2826 gnd 0.006956f
C5268 vdd.n2827 gnd 0.006956f
C5269 vdd.n2828 gnd 0.006956f
C5270 vdd.n2829 gnd 0.006956f
C5271 vdd.n2830 gnd 0.006956f
C5272 vdd.n2831 gnd 0.006956f
C5273 vdd.n2832 gnd 0.006956f
C5274 vdd.n2833 gnd 0.006956f
C5275 vdd.n2834 gnd 0.006956f
C5276 vdd.n2835 gnd 0.006956f
C5277 vdd.n2836 gnd 0.006956f
C5278 vdd.n2837 gnd 0.006956f
C5279 vdd.n2838 gnd 0.006956f
C5280 vdd.n2839 gnd 0.006956f
C5281 vdd.n2840 gnd 0.006956f
C5282 vdd.n2841 gnd 0.006956f
C5283 vdd.n2842 gnd 0.006956f
C5284 vdd.n2843 gnd 0.006956f
C5285 vdd.n2844 gnd 0.006956f
C5286 vdd.n2845 gnd 0.006956f
C5287 vdd.n2846 gnd 0.006956f
C5288 vdd.n2847 gnd 0.006956f
C5289 vdd.n2848 gnd 0.006956f
C5290 vdd.n2849 gnd 0.006956f
C5291 vdd.n2850 gnd 0.006956f
C5292 vdd.n2851 gnd 0.006956f
C5293 vdd.n2852 gnd 0.01627f
C5294 vdd.n2853 gnd 0.01627f
C5295 vdd.n2855 gnd 0.8677f
C5296 vdd.n2857 gnd 0.01627f
C5297 vdd.n2858 gnd 0.01627f
C5298 vdd.n2859 gnd 0.015237f
C5299 vdd.n2860 gnd 0.006956f
C5300 vdd.n2861 gnd 0.006956f
C5301 vdd.n2862 gnd 0.376352f
C5302 vdd.n2863 gnd 0.006956f
C5303 vdd.n2864 gnd 0.006956f
C5304 vdd.n2865 gnd 0.006956f
C5305 vdd.n2866 gnd 0.006956f
C5306 vdd.n2867 gnd 0.006956f
C5307 vdd.n2868 gnd 0.423396f
C5308 vdd.n2869 gnd 0.006956f
C5309 vdd.n2870 gnd 0.006956f
C5310 vdd.n2871 gnd 0.006956f
C5311 vdd.n2872 gnd 0.006956f
C5312 vdd.n2873 gnd 0.006956f
C5313 vdd.n2874 gnd 0.710887f
C5314 vdd.n2875 gnd 0.006956f
C5315 vdd.n2876 gnd 0.006956f
C5316 vdd.n2877 gnd 0.006956f
C5317 vdd.n2878 gnd 0.006956f
C5318 vdd.n2879 gnd 0.006956f
C5319 vdd.n2880 gnd 0.47044f
C5320 vdd.n2881 gnd 0.006956f
C5321 vdd.n2882 gnd 0.006956f
C5322 vdd.n2883 gnd 0.006956f
C5323 vdd.n2884 gnd 0.006956f
C5324 vdd.n2885 gnd 0.006956f
C5325 vdd.n2886 gnd 0.627253f
C5326 vdd.n2887 gnd 0.006956f
C5327 vdd.n2888 gnd 0.006956f
C5328 vdd.n2889 gnd 0.006956f
C5329 vdd.n2890 gnd 0.006956f
C5330 vdd.n2891 gnd 0.006956f
C5331 vdd.n2892 gnd 0.569755f
C5332 vdd.n2893 gnd 0.006956f
C5333 vdd.n2894 gnd 0.006956f
C5334 vdd.n2895 gnd 0.006956f
C5335 vdd.n2896 gnd 0.006956f
C5336 vdd.n2897 gnd 0.006956f
C5337 vdd.n2898 gnd 0.412942f
C5338 vdd.n2899 gnd 0.006956f
C5339 vdd.n2900 gnd 0.006956f
C5340 vdd.n2901 gnd 0.006956f
C5341 vdd.n2902 gnd 0.006956f
C5342 vdd.n2903 gnd 0.006956f
C5343 vdd.n2904 gnd 0.224766f
C5344 vdd.n2905 gnd 0.006956f
C5345 vdd.n2906 gnd 0.006956f
C5346 vdd.n2907 gnd 0.006956f
C5347 vdd.n2908 gnd 0.006956f
C5348 vdd.n2909 gnd 0.006956f
C5349 vdd.n2910 gnd 0.611572f
C5350 vdd.n2911 gnd 0.006956f
C5351 vdd.n2912 gnd 0.006956f
C5352 vdd.n2913 gnd 0.006956f
C5353 vdd.n2914 gnd 0.006956f
C5354 vdd.n2915 gnd 0.006956f
C5355 vdd.n2916 gnd 0.710887f
C5356 vdd.n2917 gnd 0.006956f
C5357 vdd.n2918 gnd 0.006956f
C5358 vdd.n2919 gnd 0.004501f
C5359 vdd.n2920 gnd 0.020151f
C5360 vdd.n2921 gnd 0.005933f
C5361 vdd.n2922 gnd 0.006956f
C5362 vdd.n2923 gnd 0.606345f
C5363 vdd.n2924 gnd 0.006956f
C5364 vdd.n2925 gnd 0.006956f
C5365 vdd.n2926 gnd 0.006956f
C5366 vdd.n2927 gnd 0.006956f
C5367 vdd.n2928 gnd 0.006956f
C5368 vdd.n2929 gnd 0.496576f
C5369 vdd.n2930 gnd 0.006956f
C5370 vdd.n2931 gnd 0.006956f
C5371 vdd.n2932 gnd 0.006956f
C5372 vdd.n2933 gnd 0.006956f
C5373 vdd.n2934 gnd 0.006956f
C5374 vdd.n2935 gnd 0.371125f
C5375 vdd.n2936 gnd 0.006956f
C5376 vdd.n2937 gnd 0.006956f
C5377 vdd.n2938 gnd 0.006956f
C5378 vdd.n2939 gnd 0.006956f
C5379 vdd.n2940 gnd 0.006956f
C5380 vdd.n2941 gnd 0.710887f
C5381 vdd.n2942 gnd 0.006956f
C5382 vdd.n2943 gnd 0.006956f
C5383 vdd.n2944 gnd 0.006956f
C5384 vdd.n2945 gnd 0.006956f
C5385 vdd.n2946 gnd 0.006956f
C5386 vdd.n2947 gnd 0.006956f
C5387 vdd.n2949 gnd 0.006956f
C5388 vdd.n2950 gnd 0.006956f
C5389 vdd.n2952 gnd 0.006956f
C5390 vdd.n2953 gnd 0.006956f
C5391 vdd.n2956 gnd 0.006956f
C5392 vdd.n2957 gnd 0.006956f
C5393 vdd.n2958 gnd 0.006956f
C5394 vdd.n2959 gnd 0.006956f
C5395 vdd.n2961 gnd 0.006956f
C5396 vdd.n2962 gnd 0.006956f
C5397 vdd.n2963 gnd 0.006956f
C5398 vdd.n2964 gnd 0.006956f
C5399 vdd.n2965 gnd 0.006956f
C5400 vdd.n2966 gnd 0.006956f
C5401 vdd.n2968 gnd 0.006956f
C5402 vdd.n2969 gnd 0.006956f
C5403 vdd.n2970 gnd 0.006956f
C5404 vdd.n2971 gnd 0.006956f
C5405 vdd.n2972 gnd 0.006956f
C5406 vdd.n2973 gnd 0.006956f
C5407 vdd.n2975 gnd 0.006956f
C5408 vdd.n2976 gnd 0.006956f
C5409 vdd.n2977 gnd 0.006956f
C5410 vdd.n2978 gnd 0.006956f
C5411 vdd.n2979 gnd 0.006956f
C5412 vdd.n2980 gnd 0.006956f
C5413 vdd.n2982 gnd 0.006956f
C5414 vdd.n2983 gnd 0.01627f
C5415 vdd.n2984 gnd 0.01627f
C5416 vdd.n2985 gnd 0.015237f
C5417 vdd.n2986 gnd 0.006956f
C5418 vdd.n2987 gnd 0.006956f
C5419 vdd.n2988 gnd 0.006956f
C5420 vdd.n2989 gnd 0.006956f
C5421 vdd.n2990 gnd 0.006956f
C5422 vdd.n2991 gnd 0.006956f
C5423 vdd.n2992 gnd 0.710887f
C5424 vdd.n2993 gnd 0.006956f
C5425 vdd.n2994 gnd 0.006956f
C5426 vdd.n2995 gnd 0.006956f
C5427 vdd.n2996 gnd 0.006956f
C5428 vdd.n2997 gnd 0.006956f
C5429 vdd.n2998 gnd 0.465213f
C5430 vdd.n2999 gnd 0.006956f
C5431 vdd.n3000 gnd 0.006956f
C5432 vdd.n3001 gnd 0.006956f
C5433 vdd.n3002 gnd 0.016101f
C5434 vdd.n3004 gnd 0.01627f
C5435 vdd.n3005 gnd 0.015406f
C5436 vdd.n3006 gnd 0.006956f
C5437 vdd.n3007 gnd 0.005371f
C5438 vdd.n3008 gnd 0.006956f
C5439 vdd.n3010 gnd 0.006956f
C5440 vdd.n3011 gnd 0.006956f
C5441 vdd.n3012 gnd 0.006956f
C5442 vdd.n3013 gnd 0.006956f
C5443 vdd.n3014 gnd 0.006956f
C5444 vdd.n3015 gnd 0.006956f
C5445 vdd.n3017 gnd 0.006956f
C5446 vdd.n3018 gnd 0.006956f
C5447 vdd.n3019 gnd 0.006956f
C5448 vdd.n3020 gnd 0.006956f
C5449 vdd.n3021 gnd 0.006956f
C5450 vdd.n3022 gnd 0.006956f
C5451 vdd.n3024 gnd 0.006956f
C5452 vdd.n3025 gnd 0.006956f
C5453 vdd.n3026 gnd 0.006956f
C5454 vdd.n3027 gnd 0.006956f
C5455 vdd.n3028 gnd 0.006956f
C5456 vdd.n3029 gnd 0.006956f
C5457 vdd.n3031 gnd 0.006956f
C5458 vdd.n3032 gnd 0.006956f
C5459 vdd.n3033 gnd 0.006956f
C5460 vdd.n3034 gnd 0.777612f
C5461 vdd.n3035 gnd 0.02389f
C5462 vdd.n3036 gnd 0.006956f
C5463 vdd.n3037 gnd 0.006956f
C5464 vdd.n3039 gnd 0.006956f
C5465 vdd.n3040 gnd 0.006956f
C5466 vdd.n3041 gnd 0.006956f
C5467 vdd.n3042 gnd 0.006956f
C5468 vdd.n3043 gnd 0.006956f
C5469 vdd.n3044 gnd 0.006956f
C5470 vdd.n3046 gnd 0.006956f
C5471 vdd.n3047 gnd 0.006956f
C5472 vdd.n3048 gnd 0.006956f
C5473 vdd.n3049 gnd 0.006956f
C5474 vdd.n3050 gnd 0.006956f
C5475 vdd.n3051 gnd 0.006956f
C5476 vdd.n3053 gnd 0.006956f
C5477 vdd.n3054 gnd 0.006956f
C5478 vdd.n3055 gnd 0.006956f
C5479 vdd.n3056 gnd 0.006956f
C5480 vdd.n3057 gnd 0.006956f
C5481 vdd.n3058 gnd 0.006956f
C5482 vdd.n3060 gnd 0.006956f
C5483 vdd.n3061 gnd 0.006956f
C5484 vdd.n3063 gnd 0.006956f
C5485 vdd.n3064 gnd 0.006956f
C5486 vdd.n3065 gnd 0.01627f
C5487 vdd.n3066 gnd 0.015237f
C5488 vdd.n3067 gnd 0.015237f
C5489 vdd.n3068 gnd 1.00361f
C5490 vdd.n3069 gnd 0.015237f
C5491 vdd.n3070 gnd 0.01627f
C5492 vdd.n3071 gnd 0.015406f
C5493 vdd.n3072 gnd 0.006956f
C5494 vdd.n3073 gnd 0.005371f
C5495 vdd.n3074 gnd 0.006956f
C5496 vdd.n3076 gnd 0.006956f
C5497 vdd.n3077 gnd 0.006956f
C5498 vdd.n3078 gnd 0.006956f
C5499 vdd.n3079 gnd 0.006956f
C5500 vdd.n3080 gnd 0.006956f
C5501 vdd.n3081 gnd 0.006956f
C5502 vdd.n3083 gnd 0.006956f
C5503 vdd.n3084 gnd 0.006956f
C5504 vdd.n3085 gnd 0.006956f
C5505 vdd.n3086 gnd 0.006956f
C5506 vdd.n3087 gnd 0.006956f
C5507 vdd.n3088 gnd 0.006956f
C5508 vdd.n3090 gnd 0.006956f
C5509 vdd.n3091 gnd 0.006956f
C5510 vdd.n3092 gnd 0.006956f
C5511 vdd.n3093 gnd 0.006956f
C5512 vdd.n3094 gnd 0.006956f
C5513 vdd.n3095 gnd 0.006956f
C5514 vdd.n3097 gnd 0.006956f
C5515 vdd.n3098 gnd 0.006956f
C5516 vdd.n3100 gnd 0.006956f
C5517 vdd.n3101 gnd 0.02389f
C5518 vdd.n3102 gnd 0.777612f
C5519 vdd.n3103 gnd 0.008798f
C5520 vdd.n3104 gnd 0.003911f
C5521 vdd.t60 gnd 0.125851f
C5522 vdd.t61 gnd 0.134501f
C5523 vdd.t58 gnd 0.164361f
C5524 vdd.n3105 gnd 0.210687f
C5525 vdd.n3106 gnd 0.177015f
C5526 vdd.n3107 gnd 0.01268f
C5527 vdd.n3108 gnd 0.01023f
C5528 vdd.n3109 gnd 0.004323f
C5529 vdd.n3110 gnd 0.008234f
C5530 vdd.n3111 gnd 0.01023f
C5531 vdd.n3112 gnd 0.01023f
C5532 vdd.n3113 gnd 0.008234f
C5533 vdd.n3114 gnd 0.008234f
C5534 vdd.n3115 gnd 0.01023f
C5535 vdd.n3117 gnd 0.01023f
C5536 vdd.n3118 gnd 0.008234f
C5537 vdd.n3119 gnd 0.008234f
C5538 vdd.n3120 gnd 0.008234f
C5539 vdd.n3121 gnd 0.01023f
C5540 vdd.n3123 gnd 0.01023f
C5541 vdd.n3125 gnd 0.01023f
C5542 vdd.n3126 gnd 0.008234f
C5543 vdd.n3127 gnd 0.008234f
C5544 vdd.n3128 gnd 0.008234f
C5545 vdd.n3129 gnd 0.01023f
C5546 vdd.n3131 gnd 0.01023f
C5547 vdd.n3133 gnd 0.01023f
C5548 vdd.n3134 gnd 0.008234f
C5549 vdd.n3135 gnd 0.008234f
C5550 vdd.n3136 gnd 0.008234f
C5551 vdd.n3137 gnd 0.01023f
C5552 vdd.n3139 gnd 0.01023f
C5553 vdd.n3140 gnd 0.01023f
C5554 vdd.n3141 gnd 0.008234f
C5555 vdd.n3142 gnd 0.008234f
C5556 vdd.n3143 gnd 0.01023f
C5557 vdd.n3144 gnd 0.01023f
C5558 vdd.n3146 gnd 0.01023f
C5559 vdd.n3147 gnd 0.008234f
C5560 vdd.n3148 gnd 0.01023f
C5561 vdd.n3149 gnd 0.01023f
C5562 vdd.n3150 gnd 0.01023f
C5563 vdd.n3151 gnd 0.016797f
C5564 vdd.n3152 gnd 0.005599f
C5565 vdd.n3153 gnd 0.01023f
C5566 vdd.n3155 gnd 0.01023f
C5567 vdd.n3157 gnd 0.01023f
C5568 vdd.n3158 gnd 0.008234f
C5569 vdd.n3159 gnd 0.008234f
C5570 vdd.n3160 gnd 0.008234f
C5571 vdd.n3161 gnd 0.01023f
C5572 vdd.n3163 gnd 0.01023f
C5573 vdd.n3165 gnd 0.01023f
C5574 vdd.n3166 gnd 0.008234f
C5575 vdd.n3167 gnd 0.008234f
C5576 vdd.n3168 gnd 0.008234f
C5577 vdd.n3169 gnd 0.01023f
C5578 vdd.n3171 gnd 0.01023f
C5579 vdd.n3173 gnd 0.01023f
C5580 vdd.n3174 gnd 0.008234f
C5581 vdd.n3175 gnd 0.008234f
C5582 vdd.n3176 gnd 0.008234f
C5583 vdd.n3177 gnd 0.01023f
C5584 vdd.n3179 gnd 0.01023f
C5585 vdd.n3181 gnd 0.01023f
C5586 vdd.n3182 gnd 0.008234f
C5587 vdd.n3183 gnd 0.008234f
C5588 vdd.n3184 gnd 0.008234f
C5589 vdd.n3185 gnd 0.01023f
C5590 vdd.n3187 gnd 0.01023f
C5591 vdd.n3189 gnd 0.01023f
C5592 vdd.n3190 gnd 0.008234f
C5593 vdd.n3191 gnd 0.008234f
C5594 vdd.n3192 gnd 0.006875f
C5595 vdd.n3193 gnd 0.01023f
C5596 vdd.n3195 gnd 0.01023f
C5597 vdd.n3197 gnd 0.01023f
C5598 vdd.n3198 gnd 0.006875f
C5599 vdd.n3199 gnd 0.008234f
C5600 vdd.n3200 gnd 0.008234f
C5601 vdd.n3201 gnd 0.01023f
C5602 vdd.n3203 gnd 0.01023f
C5603 vdd.n3205 gnd 0.01023f
C5604 vdd.n3206 gnd 0.008234f
C5605 vdd.n3207 gnd 0.008234f
C5606 vdd.n3208 gnd 0.008234f
C5607 vdd.n3209 gnd 0.01023f
C5608 vdd.n3211 gnd 0.01023f
C5609 vdd.n3213 gnd 0.01023f
C5610 vdd.n3214 gnd 0.008234f
C5611 vdd.n3215 gnd 0.008234f
C5612 vdd.n3216 gnd 0.008234f
C5613 vdd.n3217 gnd 0.01023f
C5614 vdd.n3219 gnd 0.01023f
C5615 vdd.n3220 gnd 0.01023f
C5616 vdd.n3221 gnd 0.008234f
C5617 vdd.n3222 gnd 0.008234f
C5618 vdd.n3223 gnd 0.01023f
C5619 vdd.n3224 gnd 0.01023f
C5620 vdd.n3225 gnd 0.008234f
C5621 vdd.n3226 gnd 0.008234f
C5622 vdd.n3227 gnd 0.01023f
C5623 vdd.n3228 gnd 0.01023f
C5624 vdd.n3230 gnd 0.01023f
C5625 vdd.n3231 gnd 0.008234f
C5626 vdd.n3232 gnd 0.006834f
C5627 vdd.n3233 gnd 0.023454f
C5628 vdd.n3234 gnd 0.023295f
C5629 vdd.n3235 gnd 0.006834f
C5630 vdd.n3236 gnd 0.023295f
C5631 vdd.n3237 gnd 1.37996f
C5632 vdd.n3238 gnd 0.023295f
C5633 vdd.n3239 gnd 0.006834f
C5634 vdd.n3240 gnd 0.023295f
C5635 vdd.n3241 gnd 0.01023f
C5636 vdd.n3242 gnd 0.01023f
C5637 vdd.n3243 gnd 0.008234f
C5638 vdd.n3244 gnd 0.01023f
C5639 vdd.n3245 gnd 0.987924f
C5640 vdd.n3246 gnd 0.01023f
C5641 vdd.n3247 gnd 0.008234f
C5642 vdd.n3248 gnd 0.01023f
C5643 vdd.n3249 gnd 0.01023f
C5644 vdd.n3250 gnd 0.01023f
C5645 vdd.n3251 gnd 0.008234f
C5646 vdd.n3252 gnd 0.01023f
C5647 vdd.n3253 gnd 1.01929f
C5648 vdd.n3254 gnd 0.01023f
C5649 vdd.n3255 gnd 0.008234f
C5650 vdd.n3256 gnd 0.01023f
C5651 vdd.n3257 gnd 0.01023f
C5652 vdd.n3258 gnd 0.01023f
C5653 vdd.n3259 gnd 0.008234f
C5654 vdd.n3260 gnd 0.01023f
C5655 vdd.t236 gnd 0.522711f
C5656 vdd.n3261 gnd 0.841565f
C5657 vdd.n3262 gnd 0.01023f
C5658 vdd.n3263 gnd 0.008234f
C5659 vdd.n3264 gnd 0.01023f
C5660 vdd.n3265 gnd 0.01023f
C5661 vdd.n3266 gnd 0.01023f
C5662 vdd.n3267 gnd 0.008234f
C5663 vdd.n3268 gnd 0.01023f
C5664 vdd.n3269 gnd 0.663843f
C5665 vdd.n3270 gnd 0.01023f
C5666 vdd.n3271 gnd 0.008234f
C5667 vdd.n3272 gnd 0.01023f
C5668 vdd.n3273 gnd 0.01023f
C5669 vdd.n3274 gnd 0.01023f
C5670 vdd.n3275 gnd 0.008234f
C5671 vdd.n3276 gnd 0.01023f
C5672 vdd.n3277 gnd 0.831111f
C5673 vdd.n3278 gnd 0.559301f
C5674 vdd.n3279 gnd 0.01023f
C5675 vdd.n3280 gnd 0.008234f
C5676 vdd.n3281 gnd 0.01023f
C5677 vdd.n3282 gnd 0.01023f
C5678 vdd.n3283 gnd 0.01023f
C5679 vdd.n3284 gnd 0.008234f
C5680 vdd.n3285 gnd 0.01023f
C5681 vdd.n3286 gnd 0.737023f
C5682 vdd.n3287 gnd 0.01023f
C5683 vdd.n3288 gnd 0.008234f
C5684 vdd.n3289 gnd 0.01023f
C5685 vdd.n3290 gnd 0.01023f
C5686 vdd.n3291 gnd 0.01023f
C5687 vdd.n3292 gnd 0.01023f
C5688 vdd.n3293 gnd 0.01023f
C5689 vdd.n3294 gnd 0.008234f
C5690 vdd.n3295 gnd 0.008234f
C5691 vdd.n3296 gnd 0.01023f
C5692 vdd.t184 gnd 0.522711f
C5693 vdd.n3297 gnd 0.8677f
C5694 vdd.n3298 gnd 0.01023f
C5695 vdd.n3299 gnd 0.008234f
C5696 vdd.n3300 gnd 0.01023f
C5697 vdd.n3301 gnd 0.01023f
C5698 vdd.n3302 gnd 0.01023f
C5699 vdd.n3303 gnd 0.008234f
C5700 vdd.n3304 gnd 0.01023f
C5701 vdd.n3305 gnd 0.820656f
C5702 vdd.n3306 gnd 0.01023f
C5703 vdd.n3307 gnd 0.01023f
C5704 vdd.n3308 gnd 0.008234f
C5705 vdd.n3309 gnd 0.008234f
C5706 vdd.n3310 gnd 0.008234f
C5707 vdd.n3311 gnd 0.01023f
C5708 vdd.n3312 gnd 0.01023f
C5709 vdd.n3313 gnd 0.01023f
C5710 vdd.n3314 gnd 0.01023f
C5711 vdd.n3315 gnd 0.008234f
C5712 vdd.n3316 gnd 0.008234f
C5713 vdd.n3317 gnd 0.008234f
C5714 vdd.n3318 gnd 0.01023f
C5715 vdd.n3319 gnd 0.01023f
C5716 vdd.n3320 gnd 0.01023f
C5717 vdd.n3321 gnd 0.01023f
C5718 vdd.n3322 gnd 0.008234f
C5719 vdd.n3323 gnd 0.008234f
C5720 vdd.n3324 gnd 0.008234f
C5721 vdd.n3325 gnd 0.01023f
C5722 vdd.n3326 gnd 0.01023f
C5723 vdd.n3327 gnd 0.01023f
C5724 vdd.n3328 gnd 0.8677f
C5725 vdd.n3329 gnd 0.01023f
C5726 vdd.n3330 gnd 0.008234f
C5727 vdd.n3331 gnd 0.008234f
C5728 vdd.n3332 gnd 0.008234f
C5729 vdd.n3333 gnd 0.01023f
C5730 vdd.n3334 gnd 0.01023f
C5731 vdd.n3335 gnd 0.01023f
C5732 vdd.n3336 gnd 0.01023f
C5733 vdd.n3337 gnd 0.008234f
C5734 vdd.n3338 gnd 0.008234f
C5735 vdd.n3339 gnd 0.006834f
C5736 vdd.n3340 gnd 0.023295f
C5737 vdd.n3341 gnd 0.023454f
C5738 vdd.n3342 gnd 0.003911f
C5739 vdd.n3343 gnd 0.023454f
C5740 vdd.n3345 gnd 2.31038f
C5741 vdd.n3346 gnd 1.37996f
C5742 vdd.n3347 gnd 0.684752f
C5743 vdd.n3348 gnd 0.01023f
C5744 vdd.n3349 gnd 0.008234f
C5745 vdd.n3350 gnd 0.008234f
C5746 vdd.n3351 gnd 0.008234f
C5747 vdd.n3352 gnd 0.01023f
C5748 vdd.n3353 gnd 1.04542f
C5749 vdd.n3354 gnd 1.04542f
C5750 vdd.n3355 gnd 0.601118f
C5751 vdd.n3356 gnd 0.01023f
C5752 vdd.n3357 gnd 0.008234f
C5753 vdd.n3358 gnd 0.008234f
C5754 vdd.n3359 gnd 0.008234f
C5755 vdd.n3360 gnd 0.01023f
C5756 vdd.n3361 gnd 0.622026f
C5757 vdd.n3362 gnd 0.768385f
C5758 vdd.t152 gnd 0.522711f
C5759 vdd.n3363 gnd 0.799748f
C5760 vdd.n3364 gnd 0.01023f
C5761 vdd.n3365 gnd 0.008234f
C5762 vdd.n3366 gnd 0.008234f
C5763 vdd.n3367 gnd 0.008234f
C5764 vdd.n3368 gnd 0.01023f
C5765 vdd.n3369 gnd 0.8677f
C5766 vdd.t161 gnd 0.522711f
C5767 vdd.n3370 gnd 0.63248f
C5768 vdd.n3371 gnd 0.757931f
C5769 vdd.n3372 gnd 0.01023f
C5770 vdd.n3373 gnd 0.008234f
C5771 vdd.n3374 gnd 0.008234f
C5772 vdd.n3375 gnd 0.008234f
C5773 vdd.n3376 gnd 0.01023f
C5774 vdd.n3377 gnd 0.580209f
C5775 vdd.t182 gnd 0.522711f
C5776 vdd.n3378 gnd 0.8677f
C5777 vdd.t211 gnd 0.522711f
C5778 vdd.n3379 gnd 0.642935f
C5779 vdd.n3380 gnd 0.01023f
C5780 vdd.n3381 gnd 0.008234f
C5781 vdd.n3382 gnd 0.007862f
C5782 vdd.n3383 gnd 0.603384f
C5783 vdd.n3384 gnd 2.55924f
C5784 a_n7636_8799.n0 gnd 0.21002f
C5785 a_n7636_8799.n1 gnd 0.293544f
C5786 a_n7636_8799.n2 gnd 0.21002f
C5787 a_n7636_8799.n3 gnd 0.21002f
C5788 a_n7636_8799.n4 gnd 0.21002f
C5789 a_n7636_8799.n5 gnd 0.276692f
C5790 a_n7636_8799.n6 gnd 0.21002f
C5791 a_n7636_8799.n7 gnd 0.293544f
C5792 a_n7636_8799.n8 gnd 0.21002f
C5793 a_n7636_8799.n9 gnd 0.21002f
C5794 a_n7636_8799.n10 gnd 0.21002f
C5795 a_n7636_8799.n11 gnd 0.276692f
C5796 a_n7636_8799.n12 gnd 0.21002f
C5797 a_n7636_8799.n13 gnd 0.46004f
C5798 a_n7636_8799.n14 gnd 0.21002f
C5799 a_n7636_8799.n15 gnd 0.21002f
C5800 a_n7636_8799.n16 gnd 0.21002f
C5801 a_n7636_8799.n17 gnd 0.276692f
C5802 a_n7636_8799.n18 gnd 0.329198f
C5803 a_n7636_8799.n19 gnd 0.21002f
C5804 a_n7636_8799.n20 gnd 0.21002f
C5805 a_n7636_8799.n21 gnd 0.21002f
C5806 a_n7636_8799.n22 gnd 0.21002f
C5807 a_n7636_8799.n23 gnd 0.241039f
C5808 a_n7636_8799.n24 gnd 0.329198f
C5809 a_n7636_8799.n25 gnd 0.21002f
C5810 a_n7636_8799.n26 gnd 0.21002f
C5811 a_n7636_8799.n27 gnd 0.21002f
C5812 a_n7636_8799.n28 gnd 0.21002f
C5813 a_n7636_8799.n29 gnd 0.241039f
C5814 a_n7636_8799.n30 gnd 0.329198f
C5815 a_n7636_8799.n31 gnd 0.21002f
C5816 a_n7636_8799.n32 gnd 0.21002f
C5817 a_n7636_8799.n33 gnd 0.21002f
C5818 a_n7636_8799.n34 gnd 0.21002f
C5819 a_n7636_8799.n35 gnd 0.407535f
C5820 a_n7636_8799.n36 gnd 0.707073f
C5821 a_n7636_8799.n37 gnd 2.93241f
C5822 a_n7636_8799.n38 gnd 2.87509f
C5823 a_n7636_8799.n39 gnd 1.41136f
C5824 a_n7636_8799.n40 gnd 1.53928f
C5825 a_n7636_8799.n41 gnd 2.59195f
C5826 a_n7636_8799.n42 gnd 0.008711f
C5827 a_n7636_8799.n43 gnd 0.001169f
C5828 a_n7636_8799.n45 gnd 0.007823f
C5829 a_n7636_8799.n46 gnd 0.011824f
C5830 a_n7636_8799.n47 gnd 0.008131f
C5831 a_n7636_8799.n49 gnd 4.06e-19
C5832 a_n7636_8799.n50 gnd 0.008427f
C5833 a_n7636_8799.n51 gnd 0.011639f
C5834 a_n7636_8799.n52 gnd 0.0075f
C5835 a_n7636_8799.n53 gnd 0.008711f
C5836 a_n7636_8799.n54 gnd 0.001169f
C5837 a_n7636_8799.n56 gnd 0.007823f
C5838 a_n7636_8799.n57 gnd 0.011824f
C5839 a_n7636_8799.n58 gnd 0.008131f
C5840 a_n7636_8799.n60 gnd 4.06e-19
C5841 a_n7636_8799.n61 gnd 0.008427f
C5842 a_n7636_8799.n62 gnd 0.011639f
C5843 a_n7636_8799.n63 gnd 0.0075f
C5844 a_n7636_8799.n64 gnd 0.008711f
C5845 a_n7636_8799.n65 gnd 0.001169f
C5846 a_n7636_8799.n67 gnd 0.007823f
C5847 a_n7636_8799.n68 gnd 0.011824f
C5848 a_n7636_8799.n69 gnd 0.008131f
C5849 a_n7636_8799.n71 gnd 4.06e-19
C5850 a_n7636_8799.n72 gnd 0.008427f
C5851 a_n7636_8799.n73 gnd 0.011639f
C5852 a_n7636_8799.n74 gnd 0.0075f
C5853 a_n7636_8799.n75 gnd 0.001169f
C5854 a_n7636_8799.n77 gnd 0.007823f
C5855 a_n7636_8799.n78 gnd 0.011824f
C5856 a_n7636_8799.n79 gnd 0.008131f
C5857 a_n7636_8799.n81 gnd 4.06e-19
C5858 a_n7636_8799.n82 gnd 0.008427f
C5859 a_n7636_8799.n83 gnd 0.011639f
C5860 a_n7636_8799.n84 gnd 0.0075f
C5861 a_n7636_8799.n85 gnd 0.252844f
C5862 a_n7636_8799.n86 gnd 0.001169f
C5863 a_n7636_8799.n88 gnd 0.007823f
C5864 a_n7636_8799.n89 gnd 0.011824f
C5865 a_n7636_8799.n90 gnd 0.008131f
C5866 a_n7636_8799.n92 gnd 4.06e-19
C5867 a_n7636_8799.n93 gnd 0.008427f
C5868 a_n7636_8799.n94 gnd 0.011639f
C5869 a_n7636_8799.n95 gnd 0.0075f
C5870 a_n7636_8799.n96 gnd 0.252844f
C5871 a_n7636_8799.n97 gnd 0.001169f
C5872 a_n7636_8799.n99 gnd 0.007823f
C5873 a_n7636_8799.n100 gnd 0.011824f
C5874 a_n7636_8799.n101 gnd 0.008131f
C5875 a_n7636_8799.n103 gnd 4.06e-19
C5876 a_n7636_8799.n104 gnd 0.008427f
C5877 a_n7636_8799.n105 gnd 0.011639f
C5878 a_n7636_8799.n106 gnd 0.0075f
C5879 a_n7636_8799.n107 gnd 0.252844f
C5880 a_n7636_8799.t19 gnd 0.145672f
C5881 a_n7636_8799.t12 gnd 0.145672f
C5882 a_n7636_8799.t29 gnd 0.145672f
C5883 a_n7636_8799.n108 gnd 1.14894f
C5884 a_n7636_8799.t23 gnd 0.145672f
C5885 a_n7636_8799.t7 gnd 0.145672f
C5886 a_n7636_8799.n109 gnd 1.14894f
C5887 a_n7636_8799.t32 gnd 0.145672f
C5888 a_n7636_8799.t6 gnd 0.145672f
C5889 a_n7636_8799.n110 gnd 1.14704f
C5890 a_n7636_8799.t31 gnd 0.145672f
C5891 a_n7636_8799.t28 gnd 0.145672f
C5892 a_n7636_8799.n111 gnd 1.14704f
C5893 a_n7636_8799.t18 gnd 0.145672f
C5894 a_n7636_8799.t21 gnd 0.145672f
C5895 a_n7636_8799.n112 gnd 1.14704f
C5896 a_n7636_8799.n113 gnd 3.20169f
C5897 a_n7636_8799.t14 gnd 0.113301f
C5898 a_n7636_8799.t33 gnd 0.113301f
C5899 a_n7636_8799.n114 gnd 1.00276f
C5900 a_n7636_8799.t15 gnd 0.113301f
C5901 a_n7636_8799.t17 gnd 0.113301f
C5902 a_n7636_8799.n115 gnd 1.00117f
C5903 a_n7636_8799.t11 gnd 0.113301f
C5904 a_n7636_8799.t34 gnd 0.113301f
C5905 a_n7636_8799.n116 gnd 1.00117f
C5906 a_n7636_8799.t10 gnd 0.113301f
C5907 a_n7636_8799.t25 gnd 0.113301f
C5908 a_n7636_8799.n117 gnd 1.00276f
C5909 a_n7636_8799.t35 gnd 0.113301f
C5910 a_n7636_8799.t26 gnd 0.113301f
C5911 a_n7636_8799.n118 gnd 1.00116f
C5912 a_n7636_8799.t24 gnd 0.113301f
C5913 a_n7636_8799.t9 gnd 0.113301f
C5914 a_n7636_8799.n119 gnd 1.00116f
C5915 a_n7636_8799.t27 gnd 0.113301f
C5916 a_n7636_8799.t22 gnd 0.113301f
C5917 a_n7636_8799.n120 gnd 1.00276f
C5918 a_n7636_8799.t0 gnd 0.113301f
C5919 a_n7636_8799.t2 gnd 0.113301f
C5920 a_n7636_8799.n121 gnd 1.00116f
C5921 a_n7636_8799.t20 gnd 0.113301f
C5922 a_n7636_8799.t4 gnd 0.113301f
C5923 a_n7636_8799.n122 gnd 1.00117f
C5924 a_n7636_8799.t5 gnd 0.113301f
C5925 a_n7636_8799.t13 gnd 0.113301f
C5926 a_n7636_8799.n123 gnd 1.00117f
C5927 a_n7636_8799.t78 gnd 0.604025f
C5928 a_n7636_8799.n124 gnd 0.270045f
C5929 a_n7636_8799.t36 gnd 0.604025f
C5930 a_n7636_8799.t61 gnd 0.604025f
C5931 a_n7636_8799.n125 gnd 0.273391f
C5932 a_n7636_8799.t62 gnd 0.604025f
C5933 a_n7636_8799.t72 gnd 0.604025f
C5934 a_n7636_8799.t98 gnd 0.604025f
C5935 a_n7636_8799.n126 gnd 0.275497f
C5936 a_n7636_8799.t114 gnd 0.604025f
C5937 a_n7636_8799.t117 gnd 0.604025f
C5938 a_n7636_8799.n127 gnd 0.26896f
C5939 a_n7636_8799.t115 gnd 0.615458f
C5940 a_n7636_8799.n128 gnd 0.253234f
C5941 a_n7636_8799.n129 gnd 0.011915f
C5942 a_n7636_8799.t73 gnd 0.604025f
C5943 a_n7636_8799.n130 gnd 0.269769f
C5944 a_n7636_8799.n131 gnd 0.273376f
C5945 a_n7636_8799.t71 gnd 0.604025f
C5946 a_n7636_8799.n132 gnd 0.26986f
C5947 a_n7636_8799.n133 gnd 0.264428f
C5948 a_n7636_8799.t96 gnd 0.604025f
C5949 a_n7636_8799.n134 gnd 0.269607f
C5950 a_n7636_8799.n135 gnd 0.275936f
C5951 a_n7636_8799.t93 gnd 0.604025f
C5952 a_n7636_8799.n136 gnd 0.273257f
C5953 a_n7636_8799.n137 gnd 0.269284f
C5954 a_n7636_8799.t60 gnd 0.604025f
C5955 a_n7636_8799.n138 gnd 0.264752f
C5956 a_n7636_8799.t116 gnd 0.604025f
C5957 a_n7636_8799.n139 gnd 0.273375f
C5958 a_n7636_8799.t45 gnd 0.615447f
C5959 a_n7636_8799.t87 gnd 0.604025f
C5960 a_n7636_8799.n140 gnd 0.270045f
C5961 a_n7636_8799.t44 gnd 0.604025f
C5962 a_n7636_8799.t69 gnd 0.604025f
C5963 a_n7636_8799.n141 gnd 0.273391f
C5964 a_n7636_8799.t70 gnd 0.604025f
C5965 a_n7636_8799.t80 gnd 0.604025f
C5966 a_n7636_8799.t111 gnd 0.604025f
C5967 a_n7636_8799.n142 gnd 0.275497f
C5968 a_n7636_8799.t126 gnd 0.604025f
C5969 a_n7636_8799.t130 gnd 0.604025f
C5970 a_n7636_8799.n143 gnd 0.26896f
C5971 a_n7636_8799.t128 gnd 0.615458f
C5972 a_n7636_8799.n144 gnd 0.253234f
C5973 a_n7636_8799.n145 gnd 0.011915f
C5974 a_n7636_8799.t81 gnd 0.604025f
C5975 a_n7636_8799.n146 gnd 0.269769f
C5976 a_n7636_8799.n147 gnd 0.273376f
C5977 a_n7636_8799.t79 gnd 0.604025f
C5978 a_n7636_8799.n148 gnd 0.26986f
C5979 a_n7636_8799.n149 gnd 0.264428f
C5980 a_n7636_8799.t109 gnd 0.604025f
C5981 a_n7636_8799.n150 gnd 0.269607f
C5982 a_n7636_8799.n151 gnd 0.275936f
C5983 a_n7636_8799.t105 gnd 0.604025f
C5984 a_n7636_8799.n152 gnd 0.273257f
C5985 a_n7636_8799.n153 gnd 0.269284f
C5986 a_n7636_8799.t66 gnd 0.604025f
C5987 a_n7636_8799.n154 gnd 0.264752f
C5988 a_n7636_8799.t129 gnd 0.604025f
C5989 a_n7636_8799.n155 gnd 0.273375f
C5990 a_n7636_8799.t55 gnd 0.615447f
C5991 a_n7636_8799.n156 gnd 0.909729f
C5992 a_n7636_8799.t89 gnd 0.604025f
C5993 a_n7636_8799.n157 gnd 0.270045f
C5994 a_n7636_8799.t77 gnd 0.604025f
C5995 a_n7636_8799.t121 gnd 0.604025f
C5996 a_n7636_8799.n158 gnd 0.273391f
C5997 a_n7636_8799.t97 gnd 0.604025f
C5998 a_n7636_8799.t37 gnd 0.604025f
C5999 a_n7636_8799.t67 gnd 0.604025f
C6000 a_n7636_8799.n159 gnd 0.275497f
C6001 a_n7636_8799.t118 gnd 0.604025f
C6002 a_n7636_8799.t76 gnd 0.604025f
C6003 a_n7636_8799.n160 gnd 0.26896f
C6004 a_n7636_8799.t94 gnd 0.615458f
C6005 a_n7636_8799.n161 gnd 0.253234f
C6006 a_n7636_8799.n162 gnd 0.011915f
C6007 a_n7636_8799.t110 gnd 0.604025f
C6008 a_n7636_8799.n163 gnd 0.269769f
C6009 a_n7636_8799.n164 gnd 0.273376f
C6010 a_n7636_8799.t49 gnd 0.604025f
C6011 a_n7636_8799.n165 gnd 0.26986f
C6012 a_n7636_8799.n166 gnd 0.264428f
C6013 a_n7636_8799.t82 gnd 0.604025f
C6014 a_n7636_8799.n167 gnd 0.269607f
C6015 a_n7636_8799.n168 gnd 0.275936f
C6016 a_n7636_8799.t125 gnd 0.604025f
C6017 a_n7636_8799.n169 gnd 0.273257f
C6018 a_n7636_8799.n170 gnd 0.269284f
C6019 a_n7636_8799.t41 gnd 0.604025f
C6020 a_n7636_8799.n171 gnd 0.264752f
C6021 a_n7636_8799.t53 gnd 0.604025f
C6022 a_n7636_8799.n172 gnd 0.273375f
C6023 a_n7636_8799.t106 gnd 0.615447f
C6024 a_n7636_8799.n173 gnd 1.55929f
C6025 a_n7636_8799.t75 gnd 0.604025f
C6026 a_n7636_8799.t57 gnd 0.604025f
C6027 a_n7636_8799.t120 gnd 0.604025f
C6028 a_n7636_8799.n174 gnd 0.272973f
C6029 a_n7636_8799.t88 gnd 0.604025f
C6030 a_n7636_8799.t86 gnd 0.604025f
C6031 a_n7636_8799.t38 gnd 0.604025f
C6032 a_n7636_8799.n175 gnd 0.26986f
C6033 a_n7636_8799.t92 gnd 0.604025f
C6034 a_n7636_8799.t91 gnd 0.604025f
C6035 a_n7636_8799.t40 gnd 0.604025f
C6036 a_n7636_8799.n176 gnd 0.273391f
C6037 a_n7636_8799.t39 gnd 0.604025f
C6038 a_n7636_8799.t108 gnd 0.604025f
C6039 a_n7636_8799.t52 gnd 0.604025f
C6040 a_n7636_8799.n177 gnd 0.269284f
C6041 a_n7636_8799.t43 gnd 0.604025f
C6042 a_n7636_8799.t112 gnd 0.604025f
C6043 a_n7636_8799.t74 gnd 0.604025f
C6044 a_n7636_8799.n178 gnd 0.273375f
C6045 a_n7636_8799.t56 gnd 0.615458f
C6046 a_n7636_8799.n179 gnd 0.253234f
C6047 a_n7636_8799.n180 gnd 0.270045f
C6048 a_n7636_8799.n181 gnd 0.264752f
C6049 a_n7636_8799.n182 gnd 0.273257f
C6050 a_n7636_8799.n183 gnd 0.275936f
C6051 a_n7636_8799.n184 gnd 0.269607f
C6052 a_n7636_8799.n185 gnd 0.264428f
C6053 a_n7636_8799.n186 gnd 0.273376f
C6054 a_n7636_8799.n187 gnd 0.275497f
C6055 a_n7636_8799.n188 gnd 0.26896f
C6056 a_n7636_8799.n189 gnd 0.264266f
C6057 a_n7636_8799.t84 gnd 0.604025f
C6058 a_n7636_8799.t64 gnd 0.604025f
C6059 a_n7636_8799.t131 gnd 0.604025f
C6060 a_n7636_8799.n190 gnd 0.272973f
C6061 a_n7636_8799.t101 gnd 0.604025f
C6062 a_n7636_8799.t100 gnd 0.604025f
C6063 a_n7636_8799.t46 gnd 0.604025f
C6064 a_n7636_8799.n191 gnd 0.26986f
C6065 a_n7636_8799.t104 gnd 0.604025f
C6066 a_n7636_8799.t103 gnd 0.604025f
C6067 a_n7636_8799.t48 gnd 0.604025f
C6068 a_n7636_8799.n192 gnd 0.273391f
C6069 a_n7636_8799.t47 gnd 0.604025f
C6070 a_n7636_8799.t123 gnd 0.604025f
C6071 a_n7636_8799.t63 gnd 0.604025f
C6072 a_n7636_8799.n193 gnd 0.269284f
C6073 a_n7636_8799.t51 gnd 0.604025f
C6074 a_n7636_8799.t124 gnd 0.604025f
C6075 a_n7636_8799.t85 gnd 0.604025f
C6076 a_n7636_8799.n194 gnd 0.273375f
C6077 a_n7636_8799.t65 gnd 0.615458f
C6078 a_n7636_8799.n195 gnd 0.253234f
C6079 a_n7636_8799.n196 gnd 0.270045f
C6080 a_n7636_8799.n197 gnd 0.264752f
C6081 a_n7636_8799.n198 gnd 0.273257f
C6082 a_n7636_8799.n199 gnd 0.275936f
C6083 a_n7636_8799.n200 gnd 0.269607f
C6084 a_n7636_8799.n201 gnd 0.264428f
C6085 a_n7636_8799.n202 gnd 0.273376f
C6086 a_n7636_8799.n203 gnd 0.275497f
C6087 a_n7636_8799.n204 gnd 0.26896f
C6088 a_n7636_8799.n205 gnd 0.264266f
C6089 a_n7636_8799.n206 gnd 0.909729f
C6090 a_n7636_8799.t107 gnd 0.604025f
C6091 a_n7636_8799.t54 gnd 0.604025f
C6092 a_n7636_8799.t90 gnd 0.604025f
C6093 a_n7636_8799.n207 gnd 0.272973f
C6094 a_n7636_8799.t42 gnd 0.604025f
C6095 a_n7636_8799.t59 gnd 0.604025f
C6096 a_n7636_8799.t127 gnd 0.604025f
C6097 a_n7636_8799.n208 gnd 0.26986f
C6098 a_n7636_8799.t99 gnd 0.604025f
C6099 a_n7636_8799.t122 gnd 0.604025f
C6100 a_n7636_8799.t83 gnd 0.604025f
C6101 a_n7636_8799.n209 gnd 0.273391f
C6102 a_n7636_8799.t102 gnd 0.604025f
C6103 a_n7636_8799.t50 gnd 0.604025f
C6104 a_n7636_8799.t119 gnd 0.604025f
C6105 a_n7636_8799.n210 gnd 0.269284f
C6106 a_n7636_8799.t68 gnd 0.604025f
C6107 a_n7636_8799.t113 gnd 0.604025f
C6108 a_n7636_8799.t58 gnd 0.604025f
C6109 a_n7636_8799.n211 gnd 0.273375f
C6110 a_n7636_8799.t95 gnd 0.615458f
C6111 a_n7636_8799.n212 gnd 0.253234f
C6112 a_n7636_8799.n213 gnd 0.270045f
C6113 a_n7636_8799.n214 gnd 0.264752f
C6114 a_n7636_8799.n215 gnd 0.273257f
C6115 a_n7636_8799.n216 gnd 0.275936f
C6116 a_n7636_8799.n217 gnd 0.269607f
C6117 a_n7636_8799.n218 gnd 0.264428f
C6118 a_n7636_8799.n219 gnd 0.273376f
C6119 a_n7636_8799.n220 gnd 0.275497f
C6120 a_n7636_8799.n221 gnd 0.26896f
C6121 a_n7636_8799.n222 gnd 0.264266f
C6122 a_n7636_8799.n223 gnd 1.25333f
C6123 a_n7636_8799.n224 gnd 14.1324f
C6124 a_n7636_8799.n225 gnd 4.42059f
C6125 a_n7636_8799.n226 gnd 6.41463f
C6126 a_n7636_8799.t3 gnd 0.145672f
C6127 a_n7636_8799.t8 gnd 0.145672f
C6128 a_n7636_8799.n227 gnd 1.14704f
C6129 a_n7636_8799.t30 gnd 0.145672f
C6130 a_n7636_8799.t16 gnd 0.145672f
C6131 a_n7636_8799.n228 gnd 1.14704f
C6132 a_n7636_8799.n229 gnd 1.03105f
C6133 a_n7636_8799.n230 gnd 1.14705f
C6134 a_n7636_8799.t1 gnd 0.145672f
.ends

