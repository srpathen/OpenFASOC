* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t160 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X1 commonsourceibias.t63 commonsourceibias.t62 gnd.t284 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 gnd.t283 commonsourceibias.t64 CSoutput.t89 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 vdd.t146 a_n6972_8799.t36 CSoutput.t69 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 a_n1986_8322.t13 a_n2848_n452.t48 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 a_n1808_13878.t11 a_n2848_n452.t15 a_n2848_n452.t16 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X6 a_n6972_8799.t27 plus.t5 a_n3106_n452.t52 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X7 gnd.t282 commonsourceibias.t65 CSoutput.t49 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n3106_n452.t51 plus.t6 a_n6972_8799.t6 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 a_n2848_n452.t36 a_n2848_n452.t35 a_n1808_13878.t10 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 a_n1808_13878.t9 a_n2848_n452.t27 a_n2848_n452.t28 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 vdd.t239 vdd.t237 vdd.t238 vdd.t215 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X12 CSoutput.t147 a_n6972_8799.t37 vdd.t145 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 a_n1808_13878.t19 a_n2848_n452.t49 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 gnd.t126 gnd.t124 gnd.t125 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X15 gnd.t281 commonsourceibias.t60 commonsourceibias.t61 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 vdd.t253 CSoutput.t161 output.t17 gnd.t315 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X17 vdd.t236 vdd.t234 vdd.t235 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X18 CSoutput.t109 a_n6972_8799.t38 vdd.t144 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 vdd.t143 a_n6972_8799.t39 CSoutput.t143 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t280 commonsourceibias.t66 CSoutput.t48 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t62 a_n6972_8799.t40 vdd.t142 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t279 commonsourceibias.t67 CSoutput.t46 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 output.t16 CSoutput.t162 vdd.t252 gnd.t314 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X24 a_n1986_8322.t9 a_n2848_n452.t50 a_n6972_8799.t8 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 a_n2848_n452.t47 minus.t5 a_n3106_n452.t53 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 a_n6972_8799.t26 plus.t7 a_n3106_n452.t50 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 gnd.t278 commonsourceibias.t58 commonsourceibias.t59 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 CSoutput.t150 a_n6972_8799.t41 vdd.t141 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 plus.t4 gnd.t121 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X30 a_n2848_n452.t10 minus.t6 a_n3106_n452.t11 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 vdd.t140 a_n6972_8799.t42 CSoutput.t151 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 CSoutput.t163 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 output.t18 outputibias.t8 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X34 gnd.t120 gnd.t118 gnd.t119 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X35 CSoutput.t117 commonsourceibias.t68 gnd.t277 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t276 commonsourceibias.t56 commonsourceibias.t57 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t149 a_n6972_8799.t43 vdd.t139 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 vdd.t138 a_n6972_8799.t44 CSoutput.t14 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 a_n3106_n452.t49 plus.t8 a_n6972_8799.t17 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 output.t19 outputibias.t9 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X41 a_n6972_8799.t9 a_n2848_n452.t51 a_n1986_8322.t10 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X42 CSoutput.t118 a_n6972_8799.t45 vdd.t137 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X43 vdd.t136 a_n6972_8799.t46 CSoutput.t65 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 a_n3106_n452.t8 minus.t7 a_n2848_n452.t7 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 CSoutput.t144 commonsourceibias.t69 gnd.t275 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 a_n3106_n452.t54 diffpairibias.t16 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X47 vdd.t255 CSoutput.t164 output.t15 gnd.t313 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X48 output.t14 CSoutput.t165 vdd.t249 gnd.t312 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X49 output.t0 outputibias.t10 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 CSoutput.t120 commonsourceibias.t70 gnd.t274 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t99 a_n6972_8799.t47 vdd.t135 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 CSoutput.t43 a_n6972_8799.t48 vdd.t134 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t233 vdd.t231 vdd.t232 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X54 gnd.t227 commonsourceibias.t30 commonsourceibias.t31 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X55 vdd.t230 vdd.t228 vdd.t229 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X56 CSoutput.t76 commonsourceibias.t71 gnd.t273 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t117 gnd.t115 gnd.t116 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X58 CSoutput.t36 a_n6972_8799.t49 vdd.t133 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 a_n3106_n452.t48 plus.t9 a_n6972_8799.t16 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X60 a_n1808_13878.t8 a_n2848_n452.t31 a_n2848_n452.t32 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X61 vdd.t132 a_n6972_8799.t50 CSoutput.t146 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 a_n3106_n452.t47 plus.t10 a_n6972_8799.t19 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X63 a_n3106_n452.t24 minus.t8 a_n2848_n452.t43 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X64 diffpairibias.t15 diffpairibias.t14 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X65 a_n2848_n452.t22 a_n2848_n452.t21 a_n1808_13878.t7 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t125 a_n6972_8799.t51 vdd.t131 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 vdd.t227 vdd.t225 vdd.t226 vdd.t200 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X68 CSoutput.t87 a_n6972_8799.t52 vdd.t130 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 vdd.t129 a_n6972_8799.t53 CSoutput.t131 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 gnd.t272 commonsourceibias.t72 CSoutput.t115 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 gnd.t271 commonsourceibias.t73 CSoutput.t54 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 diffpairibias.t13 diffpairibias.t12 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X73 CSoutput.t41 a_n6972_8799.t54 vdd.t128 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 gnd.t270 commonsourceibias.t74 CSoutput.t0 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 commonsourceibias.t55 commonsourceibias.t54 gnd.t269 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t127 a_n6972_8799.t55 CSoutput.t155 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 vdd.t125 a_n6972_8799.t56 CSoutput.t10 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 vdd.t250 CSoutput.t166 output.t13 gnd.t311 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X79 CSoutput.t16 a_n6972_8799.t57 vdd.t124 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X80 vdd.t123 a_n6972_8799.t58 CSoutput.t159 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t153 a_n6972_8799.t59 vdd.t122 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X82 gnd.t268 commonsourceibias.t75 CSoutput.t6 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 a_n3106_n452.t10 minus.t9 a_n2848_n452.t9 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X84 CSoutput.t167 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X85 commonsourceibias.t29 commonsourceibias.t28 gnd.t226 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 a_n3106_n452.t46 plus.t11 a_n6972_8799.t22 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X87 vdd.t121 a_n6972_8799.t60 CSoutput.t44 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 gnd.t267 commonsourceibias.t76 CSoutput.t40 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n6972_8799.t21 plus.t12 a_n3106_n452.t45 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X90 commonsourceibias.t53 commonsourceibias.t52 gnd.t266 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 CSoutput.t61 a_n6972_8799.t61 vdd.t120 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 CSoutput.t17 a_n6972_8799.t62 vdd.t119 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 CSoutput.t74 commonsourceibias.t77 gnd.t265 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X94 a_n3106_n452.t55 diffpairibias.t17 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 gnd.t264 commonsourceibias.t50 commonsourceibias.t51 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 CSoutput.t57 a_n6972_8799.t63 vdd.t118 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n3106_n452.t44 plus.t13 a_n6972_8799.t30 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X98 vdd.t117 a_n6972_8799.t64 CSoutput.t137 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 gnd.t263 commonsourceibias.t48 commonsourceibias.t49 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X100 gnd.t114 gnd.t112 gnd.t113 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X101 commonsourceibias.t47 commonsourceibias.t46 gnd.t262 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 a_n2848_n452.t20 a_n2848_n452.t19 a_n1808_13878.t6 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X103 a_n2848_n452.t30 a_n2848_n452.t29 a_n1808_13878.t5 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X104 vdd.t116 a_n6972_8799.t65 CSoutput.t94 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 vdd.t115 a_n6972_8799.t66 CSoutput.t60 vdd.t65 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 a_n6972_8799.t5 a_n2848_n452.t52 a_n1986_8322.t6 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X107 CSoutput.t8 commonsourceibias.t78 gnd.t261 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t114 a_n6972_8799.t67 CSoutput.t105 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 a_n2848_n452.t8 minus.t10 a_n3106_n452.t9 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X110 CSoutput.t79 commonsourceibias.t79 gnd.t260 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 CSoutput.t119 commonsourceibias.t80 gnd.t259 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 vdd.t113 a_n6972_8799.t68 CSoutput.t107 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 gnd.t258 commonsourceibias.t81 CSoutput.t22 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X114 commonsourceibias.t17 commonsourceibias.t16 gnd.t257 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 CSoutput.t82 a_n6972_8799.t69 vdd.t112 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 CSoutput.t112 commonsourceibias.t82 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 CSoutput.t168 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X118 vdd.t111 a_n6972_8799.t70 CSoutput.t111 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 vdd.t224 vdd.t222 vdd.t223 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 CSoutput.t18 a_n6972_8799.t71 vdd.t110 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X121 vdd.t221 vdd.t218 vdd.t220 vdd.t219 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 gnd.t254 commonsourceibias.t83 CSoutput.t122 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 output.t1 outputibias.t11 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X124 a_n3106_n452.t22 diffpairibias.t18 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X125 vdd.t217 vdd.t214 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 gnd.t111 gnd.t109 minus.t4 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X127 gnd.t108 gnd.t106 gnd.t107 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X128 CSoutput.t169 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X129 commonsourceibias.t15 commonsourceibias.t14 gnd.t253 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t16 a_n2848_n452.t53 a_n1986_8322.t7 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 vdd.t213 vdd.t211 vdd.t212 vdd.t204 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X132 CSoutput.t63 a_n6972_8799.t72 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 a_n1986_8322.t4 a_n2848_n452.t54 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 vdd.t107 a_n6972_8799.t73 CSoutput.t157 vdd.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 gnd.t252 commonsourceibias.t12 commonsourceibias.t13 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 gnd.t250 commonsourceibias.t84 CSoutput.t27 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 vdd.t9 a_n2848_n452.t55 a_n1808_13878.t18 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 gnd.t105 gnd.t103 plus.t3 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X139 gnd.t249 commonsourceibias.t85 CSoutput.t134 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n2848_n452.t11 minus.t11 a_n3106_n452.t12 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X141 a_n6972_8799.t14 plus.t14 a_n3106_n452.t43 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X142 gnd.t247 commonsourceibias.t86 CSoutput.t58 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 commonsourceibias.t37 commonsourceibias.t36 gnd.t246 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 vdd.t210 vdd.t207 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X145 a_n6972_8799.t29 plus.t15 a_n3106_n452.t42 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X146 a_n2848_n452.t45 minus.t12 a_n3106_n452.t27 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X147 vdd.t243 CSoutput.t170 output.t12 gnd.t310 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X148 diffpairibias.t11 diffpairibias.t10 gnd.t295 gnd.t294 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X149 vdd.t206 vdd.t203 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 vdd.t105 a_n6972_8799.t74 CSoutput.t19 vdd.t104 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 gnd.t245 commonsourceibias.t87 CSoutput.t59 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 gnd.t102 gnd.t99 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X153 a_n6972_8799.t2 a_n2848_n452.t56 a_n1986_8322.t2 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 a_n1986_8322.t3 a_n2848_n452.t57 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X155 vdd.t202 vdd.t199 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X156 CSoutput.t148 commonsourceibias.t88 gnd.t244 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X157 gnd.t243 commonsourceibias.t89 CSoutput.t136 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 vdd.t103 a_n6972_8799.t75 CSoutput.t34 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n2848_n452.t34 a_n2848_n452.t33 a_n1808_13878.t4 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 a_n3106_n452.t6 minus.t13 a_n2848_n452.t5 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 commonsourceibias.t35 commonsourceibias.t34 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X162 CSoutput.t66 a_n6972_8799.t76 vdd.t102 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 a_n6972_8799.t34 a_n2848_n452.t58 a_n1986_8322.t19 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 CSoutput.t78 commonsourceibias.t90 gnd.t239 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n1808_13878.t3 a_n2848_n452.t17 a_n2848_n452.t18 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X166 a_n3106_n452.t41 plus.t16 a_n6972_8799.t20 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X167 a_n2848_n452.t44 minus.t14 a_n3106_n452.t26 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X168 vdd.t101 a_n6972_8799.t77 CSoutput.t83 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 CSoutput.t158 a_n6972_8799.t78 vdd.t100 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 vdd.t263 a_n2848_n452.t59 a_n1986_8322.t20 vdd.t262 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X171 gnd.t98 gnd.t95 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X172 a_n3106_n452.t20 diffpairibias.t19 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X173 CSoutput.t121 commonsourceibias.t91 gnd.t238 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 CSoutput.t141 a_n6972_8799.t79 vdd.t99 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 CSoutput.t96 commonsourceibias.t92 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 a_n6972_8799.t18 plus.t17 a_n3106_n452.t40 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X177 CSoutput.t3 commonsourceibias.t93 gnd.t235 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n3106_n452.t0 diffpairibias.t20 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X179 vdd.t98 a_n6972_8799.t80 CSoutput.t5 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X180 gnd.t234 commonsourceibias.t94 CSoutput.t9 gnd.t233 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X181 gnd.t232 commonsourceibias.t95 CSoutput.t39 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X182 CSoutput.t33 commonsourceibias.t96 gnd.t231 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 commonsourceibias.t33 commonsourceibias.t32 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 vdd.t244 CSoutput.t171 output.t11 gnd.t309 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X185 a_n6972_8799.t23 plus.t18 a_n3106_n452.t39 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X186 vdd.t97 a_n6972_8799.t81 CSoutput.t101 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 gnd.t228 commonsourceibias.t97 CSoutput.t64 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 gnd.t94 gnd.t91 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X189 minus.t3 gnd.t88 gnd.t90 gnd.t89 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X190 CSoutput.t26 commonsourceibias.t98 gnd.t225 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 gnd.t87 gnd.t85 gnd.t86 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X192 diffpairibias.t9 diffpairibias.t8 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 a_n2848_n452.t13 minus.t15 a_n3106_n452.t15 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 CSoutput.t127 a_n6972_8799.t82 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 a_n3106_n452.t38 plus.t19 a_n6972_8799.t31 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X196 CSoutput.t116 a_n6972_8799.t83 vdd.t94 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t45 commonsourceibias.t99 gnd.t224 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X198 gnd.t223 commonsourceibias.t100 CSoutput.t21 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 vdd.t198 vdd.t196 vdd.t197 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 a_n1808_13878.t17 a_n2848_n452.t60 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 vdd.t160 a_n2848_n452.t61 a_n1808_13878.t16 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 gnd.t222 commonsourceibias.t26 commonsourceibias.t27 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 gnd.t221 commonsourceibias.t101 CSoutput.t20 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 CSoutput.t130 a_n6972_8799.t84 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 vdd.t91 a_n6972_8799.t85 CSoutput.t98 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 gnd.t220 commonsourceibias.t102 CSoutput.t114 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 a_n3106_n452.t19 minus.t16 a_n2848_n452.t41 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X208 CSoutput.t37 commonsourceibias.t103 gnd.t219 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 diffpairibias.t7 diffpairibias.t6 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X210 CSoutput.t140 a_n6972_8799.t86 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 gnd.t218 commonsourceibias.t24 commonsourceibias.t25 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 output.t10 CSoutput.t172 vdd.t241 gnd.t308 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X213 vdd.t87 a_n6972_8799.t87 CSoutput.t126 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X214 CSoutput.t32 commonsourceibias.t104 gnd.t216 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n3106_n452.t28 minus.t17 a_n2848_n452.t46 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X216 a_n3106_n452.t37 plus.t20 a_n6972_8799.t15 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X217 gnd.t84 gnd.t82 gnd.t83 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X218 a_n1986_8322.t11 a_n2848_n452.t62 a_n6972_8799.t10 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 CSoutput.t73 a_n6972_8799.t88 vdd.t86 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 CSoutput.t138 commonsourceibias.t105 gnd.t215 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 a_n3106_n452.t7 minus.t18 a_n2848_n452.t6 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X222 vdd.t85 a_n6972_8799.t89 CSoutput.t4 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 vdd.t83 a_n6972_8799.t90 CSoutput.t2 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 CSoutput.t30 a_n6972_8799.t91 vdd.t81 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 vdd.t80 a_n6972_8799.t92 CSoutput.t51 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 vdd.t152 a_n2848_n452.t63 a_n1986_8322.t12 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X227 gnd.t214 commonsourceibias.t22 commonsourceibias.t23 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 a_n1808_13878.t15 a_n2848_n452.t64 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X229 gnd.t81 gnd.t78 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 minus.t2 gnd.t75 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X231 CSoutput.t11 commonsourceibias.t106 gnd.t213 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 gnd.t74 gnd.t71 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X233 a_n3106_n452.t25 diffpairibias.t21 gnd.t297 gnd.t296 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 vdd.t79 a_n6972_8799.t93 CSoutput.t97 vdd.t65 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 CSoutput.t53 a_n6972_8799.t94 vdd.t78 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 a_n6972_8799.t13 plus.t21 a_n3106_n452.t36 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X237 a_n2848_n452.t1 minus.t19 a_n3106_n452.t2 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X238 output.t9 CSoutput.t173 vdd.t251 gnd.t307 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X239 CSoutput.t25 commonsourceibias.t107 gnd.t212 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 CSoutput.t12 a_n6972_8799.t95 vdd.t77 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 a_n3106_n452.t5 minus.t20 a_n2848_n452.t4 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X242 gnd.t211 commonsourceibias.t108 CSoutput.t38 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t195 vdd.t193 vdd.t194 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 CSoutput.t31 commonsourceibias.t109 gnd.t209 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 gnd.t70 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X246 gnd.t208 commonsourceibias.t10 commonsourceibias.t11 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 a_n1986_8322.t8 a_n2848_n452.t65 a_n6972_8799.t7 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 vdd.t192 vdd.t190 vdd.t191 vdd.t169 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 vdd.t1 a_n2848_n452.t66 a_n1986_8322.t0 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 vdd.t76 a_n6972_8799.t96 CSoutput.t29 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t56 a_n6972_8799.t97 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 gnd.t206 commonsourceibias.t110 CSoutput.t110 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t88 a_n6972_8799.t98 vdd.t73 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 a_n3106_n452.t1 minus.t21 a_n2848_n452.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X255 vdd.t247 CSoutput.t174 output.t8 gnd.t306 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X256 gnd.t66 gnd.t64 gnd.t65 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X257 output.t7 CSoutput.t175 vdd.t246 gnd.t305 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X258 vdd.t72 a_n6972_8799.t99 CSoutput.t28 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 vdd.t71 a_n6972_8799.t100 CSoutput.t13 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 a_n3106_n452.t18 minus.t22 a_n2848_n452.t40 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X261 outputibias.t7 outputibias.t6 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X262 gnd.t63 gnd.t61 gnd.t62 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X263 CSoutput.t123 commonsourceibias.t111 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 diffpairibias.t5 diffpairibias.t4 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X265 vdd.t189 vdd.t186 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X266 outputibias.t5 outputibias.t4 gnd.t293 gnd.t292 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X267 CSoutput.t85 a_n6972_8799.t101 vdd.t70 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 a_n1808_13878.t2 a_n2848_n452.t25 a_n2848_n452.t26 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X269 gnd.t203 commonsourceibias.t112 CSoutput.t102 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 CSoutput.t92 commonsourceibias.t113 gnd.t201 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X271 a_n1986_8322.t1 a_n2848_n452.t67 a_n6972_8799.t0 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 outputibias.t3 outputibias.t2 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X273 gnd.t60 gnd.t57 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X274 gnd.t200 commonsourceibias.t114 CSoutput.t84 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 outputibias.t1 outputibias.t0 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X276 gnd.t199 commonsourceibias.t8 commonsourceibias.t9 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 vdd.t69 a_n6972_8799.t102 CSoutput.t100 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 CSoutput.t70 a_n6972_8799.t103 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 a_n3106_n452.t17 minus.t23 a_n2848_n452.t39 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X280 output.t6 CSoutput.t176 vdd.t245 gnd.t304 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X281 CSoutput.t47 commonsourceibias.t115 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 vdd.t66 a_n6972_8799.t104 CSoutput.t35 vdd.t65 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 CSoutput.t86 a_n6972_8799.t105 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 a_n1986_8322.t18 a_n2848_n452.t68 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X285 gnd.t25 gnd.t22 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X286 gnd.t56 gnd.t54 plus.t2 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X287 CSoutput.t142 commonsourceibias.t116 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 gnd.t53 gnd.t50 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X289 CSoutput.t113 commonsourceibias.t117 gnd.t193 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t192 commonsourceibias.t118 CSoutput.t81 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 gnd.t191 commonsourceibias.t20 commonsourceibias.t21 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 gnd.t49 gnd.t46 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X293 output.t5 CSoutput.t177 vdd.t254 gnd.t303 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X294 vdd.t261 a_n2848_n452.t69 a_n1808_13878.t14 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X295 vdd.t185 vdd.t183 vdd.t184 vdd.t169 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X296 CSoutput.t106 a_n6972_8799.t106 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 CSoutput.t67 a_n6972_8799.t107 vdd.t60 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t59 a_n6972_8799.t108 CSoutput.t156 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 vdd.t57 a_n6972_8799.t109 CSoutput.t72 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t182 vdd.t179 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X301 a_n1986_8322.t14 a_n2848_n452.t70 a_n6972_8799.t11 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X302 a_n3106_n452.t35 plus.t22 a_n6972_8799.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X303 vdd.t178 vdd.t176 vdd.t177 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 a_n6972_8799.t12 a_n2848_n452.t71 a_n1986_8322.t15 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X305 a_n1808_13878.t13 a_n2848_n452.t72 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X306 vdd.t56 a_n6972_8799.t110 CSoutput.t108 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 CSoutput.t95 a_n6972_8799.t111 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 gnd.t45 gnd.t43 minus.t1 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X309 a_n2848_n452.t12 minus.t24 a_n3106_n452.t14 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X310 a_n6972_8799.t3 plus.t23 a_n3106_n452.t34 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X311 CSoutput.t24 commonsourceibias.t119 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 vdd.t52 a_n6972_8799.t112 CSoutput.t145 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 a_n2848_n452.t2 minus.t25 a_n3106_n452.t3 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X314 CSoutput.t52 a_n6972_8799.t113 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 commonsourceibias.t19 commonsourceibias.t18 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 gnd.t185 commonsourceibias.t120 CSoutput.t23 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 vdd.t240 CSoutput.t178 output.t4 gnd.t302 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X318 vdd.t175 vdd.t172 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X319 vdd.t171 vdd.t168 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X320 gnd.t184 commonsourceibias.t121 CSoutput.t75 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t104 a_n6972_8799.t114 vdd.t49 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t48 a_n6972_8799.t115 CSoutput.t103 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X323 a_n1808_13878.t1 a_n2848_n452.t37 a_n2848_n452.t38 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X324 gnd.t42 gnd.t40 gnd.t41 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X325 gnd.t39 gnd.t36 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X326 a_n3106_n452.t16 minus.t26 a_n2848_n452.t14 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X327 a_n3106_n452.t21 diffpairibias.t22 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X328 gnd.t182 commonsourceibias.t122 CSoutput.t80 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 commonsourceibias.t45 commonsourceibias.t44 gnd.t180 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 vdd.t242 CSoutput.t179 output.t3 gnd.t301 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X331 a_n6972_8799.t25 plus.t24 a_n3106_n452.t33 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X332 CSoutput.t124 a_n6972_8799.t116 vdd.t47 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 vdd.t46 a_n6972_8799.t117 CSoutput.t71 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 CSoutput.t180 a_n1986_8322.t16 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X335 diffpairibias.t3 diffpairibias.t2 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X336 a_n6972_8799.t4 a_n2848_n452.t73 a_n1986_8322.t5 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X337 a_n2848_n452.t24 a_n2848_n452.t23 a_n1808_13878.t0 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X338 vdd.t45 a_n6972_8799.t118 CSoutput.t135 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X339 gnd.t35 gnd.t33 plus.t1 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X340 a_n2848_n452.t3 minus.t27 a_n3106_n452.t4 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X341 vdd.t44 a_n6972_8799.t119 CSoutput.t77 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t1 a_n6972_8799.t120 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X343 commonsourceibias.t43 commonsourceibias.t42 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t177 commonsourceibias.t123 CSoutput.t91 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 vdd.t167 vdd.t164 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X346 vdd.t40 a_n6972_8799.t121 CSoutput.t7 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 diffpairibias.t1 diffpairibias.t0 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X348 gnd.t32 gnd.t29 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X349 CSoutput.t42 a_n6972_8799.t122 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 CSoutput.t50 commonsourceibias.t124 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 vdd.t36 a_n6972_8799.t123 CSoutput.t15 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 plus.t0 gnd.t26 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X353 gnd.t173 commonsourceibias.t125 CSoutput.t129 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 CSoutput.t128 commonsourceibias.t126 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 commonsourceibias.t41 commonsourceibias.t40 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 gnd.t21 gnd.t19 minus.t0 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X357 a_n6972_8799.t24 plus.t25 a_n3106_n452.t32 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X358 gnd.t168 commonsourceibias.t38 commonsourceibias.t39 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 vdd.t257 a_n2848_n452.t74 a_n1808_13878.t12 vdd.t256 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X360 CSoutput.t152 a_n6972_8799.t124 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 CSoutput.t133 commonsourceibias.t127 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 a_n6972_8799.t28 plus.t26 a_n3106_n452.t31 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X363 a_n2848_n452.t42 minus.t28 a_n3106_n452.t23 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X364 output.t2 CSoutput.t181 vdd.t248 gnd.t300 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X365 vdd.t32 a_n6972_8799.t125 CSoutput.t132 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X366 CSoutput.t154 a_n6972_8799.t126 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 vdd.t28 a_n6972_8799.t127 CSoutput.t68 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t164 commonsourceibias.t6 commonsourceibias.t7 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 commonsourceibias.t5 commonsourceibias.t4 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t139 a_n6972_8799.t128 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 vdd.t24 a_n6972_8799.t129 CSoutput.t93 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 a_n1986_8322.t17 a_n2848_n452.t75 a_n6972_8799.t33 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X373 a_n3106_n452.t30 plus.t27 a_n6972_8799.t32 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X374 commonsourceibias.t3 commonsourceibias.t2 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X375 vdd.t22 a_n6972_8799.t130 CSoutput.t90 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t55 a_n6972_8799.t131 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 a_n3106_n452.t29 plus.t28 a_n6972_8799.t35 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X378 gnd.t158 commonsourceibias.t0 commonsourceibias.t1 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 a_n3106_n452.t13 diffpairibias.t23 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 CSoutput.n19 CSoutput.t162 184.661
R1 CSoutput.n78 CSoutput.n77 165.8
R2 CSoutput.n76 CSoutput.n0 165.8
R3 CSoutput.n75 CSoutput.n74 165.8
R4 CSoutput.n73 CSoutput.n72 165.8
R5 CSoutput.n71 CSoutput.n2 165.8
R6 CSoutput.n69 CSoutput.n68 165.8
R7 CSoutput.n67 CSoutput.n3 165.8
R8 CSoutput.n66 CSoutput.n65 165.8
R9 CSoutput.n63 CSoutput.n4 165.8
R10 CSoutput.n61 CSoutput.n60 165.8
R11 CSoutput.n59 CSoutput.n5 165.8
R12 CSoutput.n58 CSoutput.n57 165.8
R13 CSoutput.n55 CSoutput.n6 165.8
R14 CSoutput.n54 CSoutput.n53 165.8
R15 CSoutput.n52 CSoutput.n51 165.8
R16 CSoutput.n50 CSoutput.n8 165.8
R17 CSoutput.n48 CSoutput.n47 165.8
R18 CSoutput.n46 CSoutput.n9 165.8
R19 CSoutput.n45 CSoutput.n44 165.8
R20 CSoutput.n42 CSoutput.n10 165.8
R21 CSoutput.n41 CSoutput.n40 165.8
R22 CSoutput.n39 CSoutput.n38 165.8
R23 CSoutput.n37 CSoutput.n12 165.8
R24 CSoutput.n35 CSoutput.n34 165.8
R25 CSoutput.n33 CSoutput.n13 165.8
R26 CSoutput.n32 CSoutput.n31 165.8
R27 CSoutput.n29 CSoutput.n14 165.8
R28 CSoutput.n28 CSoutput.n27 165.8
R29 CSoutput.n26 CSoutput.n25 165.8
R30 CSoutput.n24 CSoutput.n16 165.8
R31 CSoutput.n22 CSoutput.n21 165.8
R32 CSoutput.n20 CSoutput.n17 165.8
R33 CSoutput.n77 CSoutput.t164 162.194
R34 CSoutput.n18 CSoutput.t179 120.501
R35 CSoutput.n23 CSoutput.t175 120.501
R36 CSoutput.n15 CSoutput.t171 120.501
R37 CSoutput.n30 CSoutput.t181 120.501
R38 CSoutput.n36 CSoutput.t161 120.501
R39 CSoutput.n11 CSoutput.t172 120.501
R40 CSoutput.n43 CSoutput.t170 120.501
R41 CSoutput.n49 CSoutput.t165 120.501
R42 CSoutput.n7 CSoutput.t174 120.501
R43 CSoutput.n56 CSoutput.t176 120.501
R44 CSoutput.n62 CSoutput.t166 120.501
R45 CSoutput.n64 CSoutput.t177 120.501
R46 CSoutput.n70 CSoutput.t178 120.501
R47 CSoutput.n1 CSoutput.t173 120.501
R48 CSoutput.n310 CSoutput.n308 103.469
R49 CSoutput.n294 CSoutput.n292 103.469
R50 CSoutput.n279 CSoutput.n277 103.469
R51 CSoutput.n112 CSoutput.n110 103.469
R52 CSoutput.n96 CSoutput.n94 103.469
R53 CSoutput.n81 CSoutput.n79 103.469
R54 CSoutput.n320 CSoutput.n319 103.111
R55 CSoutput.n318 CSoutput.n317 103.111
R56 CSoutput.n316 CSoutput.n315 103.111
R57 CSoutput.n314 CSoutput.n313 103.111
R58 CSoutput.n312 CSoutput.n311 103.111
R59 CSoutput.n310 CSoutput.n309 103.111
R60 CSoutput.n306 CSoutput.n305 103.111
R61 CSoutput.n304 CSoutput.n303 103.111
R62 CSoutput.n302 CSoutput.n301 103.111
R63 CSoutput.n300 CSoutput.n299 103.111
R64 CSoutput.n298 CSoutput.n297 103.111
R65 CSoutput.n296 CSoutput.n295 103.111
R66 CSoutput.n294 CSoutput.n293 103.111
R67 CSoutput.n291 CSoutput.n290 103.111
R68 CSoutput.n289 CSoutput.n288 103.111
R69 CSoutput.n287 CSoutput.n286 103.111
R70 CSoutput.n285 CSoutput.n284 103.111
R71 CSoutput.n283 CSoutput.n282 103.111
R72 CSoutput.n281 CSoutput.n280 103.111
R73 CSoutput.n279 CSoutput.n278 103.111
R74 CSoutput.n112 CSoutput.n111 103.111
R75 CSoutput.n114 CSoutput.n113 103.111
R76 CSoutput.n116 CSoutput.n115 103.111
R77 CSoutput.n118 CSoutput.n117 103.111
R78 CSoutput.n120 CSoutput.n119 103.111
R79 CSoutput.n122 CSoutput.n121 103.111
R80 CSoutput.n124 CSoutput.n123 103.111
R81 CSoutput.n96 CSoutput.n95 103.111
R82 CSoutput.n98 CSoutput.n97 103.111
R83 CSoutput.n100 CSoutput.n99 103.111
R84 CSoutput.n102 CSoutput.n101 103.111
R85 CSoutput.n104 CSoutput.n103 103.111
R86 CSoutput.n106 CSoutput.n105 103.111
R87 CSoutput.n108 CSoutput.n107 103.111
R88 CSoutput.n81 CSoutput.n80 103.111
R89 CSoutput.n83 CSoutput.n82 103.111
R90 CSoutput.n85 CSoutput.n84 103.111
R91 CSoutput.n87 CSoutput.n86 103.111
R92 CSoutput.n89 CSoutput.n88 103.111
R93 CSoutput.n91 CSoutput.n90 103.111
R94 CSoutput.n93 CSoutput.n92 103.111
R95 CSoutput.n322 CSoutput.n321 103.111
R96 CSoutput.n342 CSoutput.n340 81.5057
R97 CSoutput.n327 CSoutput.n325 81.5057
R98 CSoutput.n374 CSoutput.n372 81.5057
R99 CSoutput.n359 CSoutput.n357 81.5057
R100 CSoutput.n354 CSoutput.n353 80.9324
R101 CSoutput.n352 CSoutput.n351 80.9324
R102 CSoutput.n350 CSoutput.n349 80.9324
R103 CSoutput.n348 CSoutput.n347 80.9324
R104 CSoutput.n346 CSoutput.n345 80.9324
R105 CSoutput.n344 CSoutput.n343 80.9324
R106 CSoutput.n342 CSoutput.n341 80.9324
R107 CSoutput.n339 CSoutput.n338 80.9324
R108 CSoutput.n337 CSoutput.n336 80.9324
R109 CSoutput.n335 CSoutput.n334 80.9324
R110 CSoutput.n333 CSoutput.n332 80.9324
R111 CSoutput.n331 CSoutput.n330 80.9324
R112 CSoutput.n329 CSoutput.n328 80.9324
R113 CSoutput.n327 CSoutput.n326 80.9324
R114 CSoutput.n374 CSoutput.n373 80.9324
R115 CSoutput.n376 CSoutput.n375 80.9324
R116 CSoutput.n378 CSoutput.n377 80.9324
R117 CSoutput.n380 CSoutput.n379 80.9324
R118 CSoutput.n382 CSoutput.n381 80.9324
R119 CSoutput.n384 CSoutput.n383 80.9324
R120 CSoutput.n386 CSoutput.n385 80.9324
R121 CSoutput.n359 CSoutput.n358 80.9324
R122 CSoutput.n361 CSoutput.n360 80.9324
R123 CSoutput.n363 CSoutput.n362 80.9324
R124 CSoutput.n365 CSoutput.n364 80.9324
R125 CSoutput.n367 CSoutput.n366 80.9324
R126 CSoutput.n369 CSoutput.n368 80.9324
R127 CSoutput.n371 CSoutput.n370 80.9324
R128 CSoutput.n25 CSoutput.n24 48.1486
R129 CSoutput.n69 CSoutput.n3 48.1486
R130 CSoutput.n38 CSoutput.n37 48.1486
R131 CSoutput.n42 CSoutput.n41 48.1486
R132 CSoutput.n51 CSoutput.n50 48.1486
R133 CSoutput.n55 CSoutput.n54 48.1486
R134 CSoutput.n22 CSoutput.n17 46.462
R135 CSoutput.n72 CSoutput.n71 46.462
R136 CSoutput.n20 CSoutput.n19 44.9055
R137 CSoutput.n29 CSoutput.n28 43.7635
R138 CSoutput.n65 CSoutput.n63 43.7635
R139 CSoutput.n35 CSoutput.n13 41.7396
R140 CSoutput.n57 CSoutput.n5 41.7396
R141 CSoutput.n44 CSoutput.n9 37.0171
R142 CSoutput.n48 CSoutput.n9 37.0171
R143 CSoutput.n76 CSoutput.n75 34.9932
R144 CSoutput.n31 CSoutput.n13 32.2947
R145 CSoutput.n61 CSoutput.n5 32.2947
R146 CSoutput.n30 CSoutput.n29 29.6014
R147 CSoutput.n63 CSoutput.n62 29.6014
R148 CSoutput.n19 CSoutput.n18 28.4085
R149 CSoutput.n18 CSoutput.n17 25.1176
R150 CSoutput.n72 CSoutput.n1 25.1176
R151 CSoutput.n43 CSoutput.n42 22.0922
R152 CSoutput.n50 CSoutput.n49 22.0922
R153 CSoutput.n77 CSoutput.n76 21.8586
R154 CSoutput.n37 CSoutput.n36 18.9681
R155 CSoutput.n56 CSoutput.n55 18.9681
R156 CSoutput.n25 CSoutput.n15 17.6292
R157 CSoutput.n64 CSoutput.n3 17.6292
R158 CSoutput.n24 CSoutput.n23 15.844
R159 CSoutput.n70 CSoutput.n69 15.844
R160 CSoutput.n38 CSoutput.n11 14.5051
R161 CSoutput.n54 CSoutput.n7 14.5051
R162 CSoutput.n389 CSoutput.n78 11.6139
R163 CSoutput.n41 CSoutput.n11 11.3811
R164 CSoutput.n51 CSoutput.n7 11.3811
R165 CSoutput.n23 CSoutput.n22 10.0422
R166 CSoutput.n71 CSoutput.n70 10.0422
R167 CSoutput.n307 CSoutput.n291 9.25285
R168 CSoutput.n109 CSoutput.n93 9.25285
R169 CSoutput.n355 CSoutput.n339 8.97993
R170 CSoutput.n387 CSoutput.n371 8.97993
R171 CSoutput.n356 CSoutput.n324 8.88693
R172 CSoutput.n28 CSoutput.n15 8.25698
R173 CSoutput.n65 CSoutput.n64 8.25698
R174 CSoutput.n356 CSoutput.n355 7.89345
R175 CSoutput.n388 CSoutput.n387 7.89345
R176 CSoutput.n324 CSoutput.n323 7.12641
R177 CSoutput.n126 CSoutput.n125 7.12641
R178 CSoutput.n36 CSoutput.n35 6.91809
R179 CSoutput.n57 CSoutput.n56 6.91809
R180 CSoutput.n389 CSoutput.n126 5.29449
R181 CSoutput.n355 CSoutput.n354 5.25266
R182 CSoutput.n387 CSoutput.n386 5.25266
R183 CSoutput.n323 CSoutput.n322 5.1449
R184 CSoutput.n307 CSoutput.n306 5.1449
R185 CSoutput.n125 CSoutput.n124 5.1449
R186 CSoutput.n109 CSoutput.n108 5.1449
R187 CSoutput.n217 CSoutput.n170 4.5005
R188 CSoutput.n186 CSoutput.n170 4.5005
R189 CSoutput.n181 CSoutput.n165 4.5005
R190 CSoutput.n181 CSoutput.n167 4.5005
R191 CSoutput.n181 CSoutput.n164 4.5005
R192 CSoutput.n181 CSoutput.n168 4.5005
R193 CSoutput.n181 CSoutput.n163 4.5005
R194 CSoutput.n181 CSoutput.t180 4.5005
R195 CSoutput.n181 CSoutput.n162 4.5005
R196 CSoutput.n181 CSoutput.n169 4.5005
R197 CSoutput.n181 CSoutput.n170 4.5005
R198 CSoutput.n179 CSoutput.n165 4.5005
R199 CSoutput.n179 CSoutput.n167 4.5005
R200 CSoutput.n179 CSoutput.n164 4.5005
R201 CSoutput.n179 CSoutput.n168 4.5005
R202 CSoutput.n179 CSoutput.n163 4.5005
R203 CSoutput.n179 CSoutput.t180 4.5005
R204 CSoutput.n179 CSoutput.n162 4.5005
R205 CSoutput.n179 CSoutput.n169 4.5005
R206 CSoutput.n179 CSoutput.n170 4.5005
R207 CSoutput.n178 CSoutput.n165 4.5005
R208 CSoutput.n178 CSoutput.n167 4.5005
R209 CSoutput.n178 CSoutput.n164 4.5005
R210 CSoutput.n178 CSoutput.n168 4.5005
R211 CSoutput.n178 CSoutput.n163 4.5005
R212 CSoutput.n178 CSoutput.t180 4.5005
R213 CSoutput.n178 CSoutput.n162 4.5005
R214 CSoutput.n178 CSoutput.n169 4.5005
R215 CSoutput.n178 CSoutput.n170 4.5005
R216 CSoutput.n263 CSoutput.n165 4.5005
R217 CSoutput.n263 CSoutput.n167 4.5005
R218 CSoutput.n263 CSoutput.n164 4.5005
R219 CSoutput.n263 CSoutput.n168 4.5005
R220 CSoutput.n263 CSoutput.n163 4.5005
R221 CSoutput.n263 CSoutput.t180 4.5005
R222 CSoutput.n263 CSoutput.n162 4.5005
R223 CSoutput.n263 CSoutput.n169 4.5005
R224 CSoutput.n263 CSoutput.n170 4.5005
R225 CSoutput.n261 CSoutput.n165 4.5005
R226 CSoutput.n261 CSoutput.n167 4.5005
R227 CSoutput.n261 CSoutput.n164 4.5005
R228 CSoutput.n261 CSoutput.n168 4.5005
R229 CSoutput.n261 CSoutput.n163 4.5005
R230 CSoutput.n261 CSoutput.t180 4.5005
R231 CSoutput.n261 CSoutput.n162 4.5005
R232 CSoutput.n261 CSoutput.n169 4.5005
R233 CSoutput.n259 CSoutput.n165 4.5005
R234 CSoutput.n259 CSoutput.n167 4.5005
R235 CSoutput.n259 CSoutput.n164 4.5005
R236 CSoutput.n259 CSoutput.n168 4.5005
R237 CSoutput.n259 CSoutput.n163 4.5005
R238 CSoutput.n259 CSoutput.t180 4.5005
R239 CSoutput.n259 CSoutput.n162 4.5005
R240 CSoutput.n259 CSoutput.n169 4.5005
R241 CSoutput.n189 CSoutput.n165 4.5005
R242 CSoutput.n189 CSoutput.n167 4.5005
R243 CSoutput.n189 CSoutput.n164 4.5005
R244 CSoutput.n189 CSoutput.n168 4.5005
R245 CSoutput.n189 CSoutput.n163 4.5005
R246 CSoutput.n189 CSoutput.t180 4.5005
R247 CSoutput.n189 CSoutput.n162 4.5005
R248 CSoutput.n189 CSoutput.n169 4.5005
R249 CSoutput.n189 CSoutput.n170 4.5005
R250 CSoutput.n188 CSoutput.n165 4.5005
R251 CSoutput.n188 CSoutput.n167 4.5005
R252 CSoutput.n188 CSoutput.n164 4.5005
R253 CSoutput.n188 CSoutput.n168 4.5005
R254 CSoutput.n188 CSoutput.n163 4.5005
R255 CSoutput.n188 CSoutput.t180 4.5005
R256 CSoutput.n188 CSoutput.n162 4.5005
R257 CSoutput.n188 CSoutput.n169 4.5005
R258 CSoutput.n188 CSoutput.n170 4.5005
R259 CSoutput.n192 CSoutput.n165 4.5005
R260 CSoutput.n192 CSoutput.n167 4.5005
R261 CSoutput.n192 CSoutput.n164 4.5005
R262 CSoutput.n192 CSoutput.n168 4.5005
R263 CSoutput.n192 CSoutput.n163 4.5005
R264 CSoutput.n192 CSoutput.t180 4.5005
R265 CSoutput.n192 CSoutput.n162 4.5005
R266 CSoutput.n192 CSoutput.n169 4.5005
R267 CSoutput.n192 CSoutput.n170 4.5005
R268 CSoutput.n191 CSoutput.n165 4.5005
R269 CSoutput.n191 CSoutput.n167 4.5005
R270 CSoutput.n191 CSoutput.n164 4.5005
R271 CSoutput.n191 CSoutput.n168 4.5005
R272 CSoutput.n191 CSoutput.n163 4.5005
R273 CSoutput.n191 CSoutput.t180 4.5005
R274 CSoutput.n191 CSoutput.n162 4.5005
R275 CSoutput.n191 CSoutput.n169 4.5005
R276 CSoutput.n191 CSoutput.n170 4.5005
R277 CSoutput.n174 CSoutput.n165 4.5005
R278 CSoutput.n174 CSoutput.n167 4.5005
R279 CSoutput.n174 CSoutput.n164 4.5005
R280 CSoutput.n174 CSoutput.n168 4.5005
R281 CSoutput.n174 CSoutput.n163 4.5005
R282 CSoutput.n174 CSoutput.t180 4.5005
R283 CSoutput.n174 CSoutput.n162 4.5005
R284 CSoutput.n174 CSoutput.n169 4.5005
R285 CSoutput.n174 CSoutput.n170 4.5005
R286 CSoutput.n266 CSoutput.n165 4.5005
R287 CSoutput.n266 CSoutput.n167 4.5005
R288 CSoutput.n266 CSoutput.n164 4.5005
R289 CSoutput.n266 CSoutput.n168 4.5005
R290 CSoutput.n266 CSoutput.n163 4.5005
R291 CSoutput.n266 CSoutput.t180 4.5005
R292 CSoutput.n266 CSoutput.n162 4.5005
R293 CSoutput.n266 CSoutput.n169 4.5005
R294 CSoutput.n266 CSoutput.n170 4.5005
R295 CSoutput.n253 CSoutput.n224 4.5005
R296 CSoutput.n253 CSoutput.n230 4.5005
R297 CSoutput.n211 CSoutput.n200 4.5005
R298 CSoutput.n211 CSoutput.n202 4.5005
R299 CSoutput.n211 CSoutput.n199 4.5005
R300 CSoutput.n211 CSoutput.n203 4.5005
R301 CSoutput.n211 CSoutput.n198 4.5005
R302 CSoutput.n211 CSoutput.t160 4.5005
R303 CSoutput.n211 CSoutput.n197 4.5005
R304 CSoutput.n211 CSoutput.n204 4.5005
R305 CSoutput.n253 CSoutput.n211 4.5005
R306 CSoutput.n232 CSoutput.n200 4.5005
R307 CSoutput.n232 CSoutput.n202 4.5005
R308 CSoutput.n232 CSoutput.n199 4.5005
R309 CSoutput.n232 CSoutput.n203 4.5005
R310 CSoutput.n232 CSoutput.n198 4.5005
R311 CSoutput.n232 CSoutput.t160 4.5005
R312 CSoutput.n232 CSoutput.n197 4.5005
R313 CSoutput.n232 CSoutput.n204 4.5005
R314 CSoutput.n253 CSoutput.n232 4.5005
R315 CSoutput.n210 CSoutput.n200 4.5005
R316 CSoutput.n210 CSoutput.n202 4.5005
R317 CSoutput.n210 CSoutput.n199 4.5005
R318 CSoutput.n210 CSoutput.n203 4.5005
R319 CSoutput.n210 CSoutput.n198 4.5005
R320 CSoutput.n210 CSoutput.t160 4.5005
R321 CSoutput.n210 CSoutput.n197 4.5005
R322 CSoutput.n210 CSoutput.n204 4.5005
R323 CSoutput.n253 CSoutput.n210 4.5005
R324 CSoutput.n234 CSoutput.n200 4.5005
R325 CSoutput.n234 CSoutput.n202 4.5005
R326 CSoutput.n234 CSoutput.n199 4.5005
R327 CSoutput.n234 CSoutput.n203 4.5005
R328 CSoutput.n234 CSoutput.n198 4.5005
R329 CSoutput.n234 CSoutput.t160 4.5005
R330 CSoutput.n234 CSoutput.n197 4.5005
R331 CSoutput.n234 CSoutput.n204 4.5005
R332 CSoutput.n253 CSoutput.n234 4.5005
R333 CSoutput.n200 CSoutput.n195 4.5005
R334 CSoutput.n202 CSoutput.n195 4.5005
R335 CSoutput.n199 CSoutput.n195 4.5005
R336 CSoutput.n203 CSoutput.n195 4.5005
R337 CSoutput.n198 CSoutput.n195 4.5005
R338 CSoutput.t160 CSoutput.n195 4.5005
R339 CSoutput.n197 CSoutput.n195 4.5005
R340 CSoutput.n204 CSoutput.n195 4.5005
R341 CSoutput.n256 CSoutput.n200 4.5005
R342 CSoutput.n256 CSoutput.n202 4.5005
R343 CSoutput.n256 CSoutput.n199 4.5005
R344 CSoutput.n256 CSoutput.n203 4.5005
R345 CSoutput.n256 CSoutput.n198 4.5005
R346 CSoutput.n256 CSoutput.t160 4.5005
R347 CSoutput.n256 CSoutput.n197 4.5005
R348 CSoutput.n256 CSoutput.n204 4.5005
R349 CSoutput.n254 CSoutput.n200 4.5005
R350 CSoutput.n254 CSoutput.n202 4.5005
R351 CSoutput.n254 CSoutput.n199 4.5005
R352 CSoutput.n254 CSoutput.n203 4.5005
R353 CSoutput.n254 CSoutput.n198 4.5005
R354 CSoutput.n254 CSoutput.t160 4.5005
R355 CSoutput.n254 CSoutput.n197 4.5005
R356 CSoutput.n254 CSoutput.n204 4.5005
R357 CSoutput.n254 CSoutput.n253 4.5005
R358 CSoutput.n236 CSoutput.n200 4.5005
R359 CSoutput.n236 CSoutput.n202 4.5005
R360 CSoutput.n236 CSoutput.n199 4.5005
R361 CSoutput.n236 CSoutput.n203 4.5005
R362 CSoutput.n236 CSoutput.n198 4.5005
R363 CSoutput.n236 CSoutput.t160 4.5005
R364 CSoutput.n236 CSoutput.n197 4.5005
R365 CSoutput.n236 CSoutput.n204 4.5005
R366 CSoutput.n253 CSoutput.n236 4.5005
R367 CSoutput.n208 CSoutput.n200 4.5005
R368 CSoutput.n208 CSoutput.n202 4.5005
R369 CSoutput.n208 CSoutput.n199 4.5005
R370 CSoutput.n208 CSoutput.n203 4.5005
R371 CSoutput.n208 CSoutput.n198 4.5005
R372 CSoutput.n208 CSoutput.t160 4.5005
R373 CSoutput.n208 CSoutput.n197 4.5005
R374 CSoutput.n208 CSoutput.n204 4.5005
R375 CSoutput.n253 CSoutput.n208 4.5005
R376 CSoutput.n238 CSoutput.n200 4.5005
R377 CSoutput.n238 CSoutput.n202 4.5005
R378 CSoutput.n238 CSoutput.n199 4.5005
R379 CSoutput.n238 CSoutput.n203 4.5005
R380 CSoutput.n238 CSoutput.n198 4.5005
R381 CSoutput.n238 CSoutput.t160 4.5005
R382 CSoutput.n238 CSoutput.n197 4.5005
R383 CSoutput.n238 CSoutput.n204 4.5005
R384 CSoutput.n253 CSoutput.n238 4.5005
R385 CSoutput.n207 CSoutput.n200 4.5005
R386 CSoutput.n207 CSoutput.n202 4.5005
R387 CSoutput.n207 CSoutput.n199 4.5005
R388 CSoutput.n207 CSoutput.n203 4.5005
R389 CSoutput.n207 CSoutput.n198 4.5005
R390 CSoutput.n207 CSoutput.t160 4.5005
R391 CSoutput.n207 CSoutput.n197 4.5005
R392 CSoutput.n207 CSoutput.n204 4.5005
R393 CSoutput.n253 CSoutput.n207 4.5005
R394 CSoutput.n252 CSoutput.n200 4.5005
R395 CSoutput.n252 CSoutput.n202 4.5005
R396 CSoutput.n252 CSoutput.n199 4.5005
R397 CSoutput.n252 CSoutput.n203 4.5005
R398 CSoutput.n252 CSoutput.n198 4.5005
R399 CSoutput.n252 CSoutput.t160 4.5005
R400 CSoutput.n252 CSoutput.n197 4.5005
R401 CSoutput.n252 CSoutput.n204 4.5005
R402 CSoutput.n253 CSoutput.n252 4.5005
R403 CSoutput.n251 CSoutput.n136 4.5005
R404 CSoutput.n152 CSoutput.n136 4.5005
R405 CSoutput.n147 CSoutput.n131 4.5005
R406 CSoutput.n147 CSoutput.n133 4.5005
R407 CSoutput.n147 CSoutput.n130 4.5005
R408 CSoutput.n147 CSoutput.n134 4.5005
R409 CSoutput.n147 CSoutput.n129 4.5005
R410 CSoutput.n147 CSoutput.t168 4.5005
R411 CSoutput.n147 CSoutput.n128 4.5005
R412 CSoutput.n147 CSoutput.n135 4.5005
R413 CSoutput.n147 CSoutput.n136 4.5005
R414 CSoutput.n145 CSoutput.n131 4.5005
R415 CSoutput.n145 CSoutput.n133 4.5005
R416 CSoutput.n145 CSoutput.n130 4.5005
R417 CSoutput.n145 CSoutput.n134 4.5005
R418 CSoutput.n145 CSoutput.n129 4.5005
R419 CSoutput.n145 CSoutput.t168 4.5005
R420 CSoutput.n145 CSoutput.n128 4.5005
R421 CSoutput.n145 CSoutput.n135 4.5005
R422 CSoutput.n145 CSoutput.n136 4.5005
R423 CSoutput.n144 CSoutput.n131 4.5005
R424 CSoutput.n144 CSoutput.n133 4.5005
R425 CSoutput.n144 CSoutput.n130 4.5005
R426 CSoutput.n144 CSoutput.n134 4.5005
R427 CSoutput.n144 CSoutput.n129 4.5005
R428 CSoutput.n144 CSoutput.t168 4.5005
R429 CSoutput.n144 CSoutput.n128 4.5005
R430 CSoutput.n144 CSoutput.n135 4.5005
R431 CSoutput.n144 CSoutput.n136 4.5005
R432 CSoutput.n273 CSoutput.n131 4.5005
R433 CSoutput.n273 CSoutput.n133 4.5005
R434 CSoutput.n273 CSoutput.n130 4.5005
R435 CSoutput.n273 CSoutput.n134 4.5005
R436 CSoutput.n273 CSoutput.n129 4.5005
R437 CSoutput.n273 CSoutput.t168 4.5005
R438 CSoutput.n273 CSoutput.n128 4.5005
R439 CSoutput.n273 CSoutput.n135 4.5005
R440 CSoutput.n273 CSoutput.n136 4.5005
R441 CSoutput.n271 CSoutput.n131 4.5005
R442 CSoutput.n271 CSoutput.n133 4.5005
R443 CSoutput.n271 CSoutput.n130 4.5005
R444 CSoutput.n271 CSoutput.n134 4.5005
R445 CSoutput.n271 CSoutput.n129 4.5005
R446 CSoutput.n271 CSoutput.t168 4.5005
R447 CSoutput.n271 CSoutput.n128 4.5005
R448 CSoutput.n271 CSoutput.n135 4.5005
R449 CSoutput.n269 CSoutput.n131 4.5005
R450 CSoutput.n269 CSoutput.n133 4.5005
R451 CSoutput.n269 CSoutput.n130 4.5005
R452 CSoutput.n269 CSoutput.n134 4.5005
R453 CSoutput.n269 CSoutput.n129 4.5005
R454 CSoutput.n269 CSoutput.t168 4.5005
R455 CSoutput.n269 CSoutput.n128 4.5005
R456 CSoutput.n269 CSoutput.n135 4.5005
R457 CSoutput.n155 CSoutput.n131 4.5005
R458 CSoutput.n155 CSoutput.n133 4.5005
R459 CSoutput.n155 CSoutput.n130 4.5005
R460 CSoutput.n155 CSoutput.n134 4.5005
R461 CSoutput.n155 CSoutput.n129 4.5005
R462 CSoutput.n155 CSoutput.t168 4.5005
R463 CSoutput.n155 CSoutput.n128 4.5005
R464 CSoutput.n155 CSoutput.n135 4.5005
R465 CSoutput.n155 CSoutput.n136 4.5005
R466 CSoutput.n154 CSoutput.n131 4.5005
R467 CSoutput.n154 CSoutput.n133 4.5005
R468 CSoutput.n154 CSoutput.n130 4.5005
R469 CSoutput.n154 CSoutput.n134 4.5005
R470 CSoutput.n154 CSoutput.n129 4.5005
R471 CSoutput.n154 CSoutput.t168 4.5005
R472 CSoutput.n154 CSoutput.n128 4.5005
R473 CSoutput.n154 CSoutput.n135 4.5005
R474 CSoutput.n154 CSoutput.n136 4.5005
R475 CSoutput.n158 CSoutput.n131 4.5005
R476 CSoutput.n158 CSoutput.n133 4.5005
R477 CSoutput.n158 CSoutput.n130 4.5005
R478 CSoutput.n158 CSoutput.n134 4.5005
R479 CSoutput.n158 CSoutput.n129 4.5005
R480 CSoutput.n158 CSoutput.t168 4.5005
R481 CSoutput.n158 CSoutput.n128 4.5005
R482 CSoutput.n158 CSoutput.n135 4.5005
R483 CSoutput.n158 CSoutput.n136 4.5005
R484 CSoutput.n157 CSoutput.n131 4.5005
R485 CSoutput.n157 CSoutput.n133 4.5005
R486 CSoutput.n157 CSoutput.n130 4.5005
R487 CSoutput.n157 CSoutput.n134 4.5005
R488 CSoutput.n157 CSoutput.n129 4.5005
R489 CSoutput.n157 CSoutput.t168 4.5005
R490 CSoutput.n157 CSoutput.n128 4.5005
R491 CSoutput.n157 CSoutput.n135 4.5005
R492 CSoutput.n157 CSoutput.n136 4.5005
R493 CSoutput.n140 CSoutput.n131 4.5005
R494 CSoutput.n140 CSoutput.n133 4.5005
R495 CSoutput.n140 CSoutput.n130 4.5005
R496 CSoutput.n140 CSoutput.n134 4.5005
R497 CSoutput.n140 CSoutput.n129 4.5005
R498 CSoutput.n140 CSoutput.t168 4.5005
R499 CSoutput.n140 CSoutput.n128 4.5005
R500 CSoutput.n140 CSoutput.n135 4.5005
R501 CSoutput.n140 CSoutput.n136 4.5005
R502 CSoutput.n276 CSoutput.n131 4.5005
R503 CSoutput.n276 CSoutput.n133 4.5005
R504 CSoutput.n276 CSoutput.n130 4.5005
R505 CSoutput.n276 CSoutput.n134 4.5005
R506 CSoutput.n276 CSoutput.n129 4.5005
R507 CSoutput.n276 CSoutput.t168 4.5005
R508 CSoutput.n276 CSoutput.n128 4.5005
R509 CSoutput.n276 CSoutput.n135 4.5005
R510 CSoutput.n276 CSoutput.n136 4.5005
R511 CSoutput.n323 CSoutput.n307 4.10845
R512 CSoutput.n125 CSoutput.n109 4.10845
R513 CSoutput.n321 CSoutput.t145 4.06363
R514 CSoutput.n321 CSoutput.t16 4.06363
R515 CSoutput.n319 CSoutput.t151 4.06363
R516 CSoutput.n319 CSoutput.t150 4.06363
R517 CSoutput.n317 CSoutput.t28 4.06363
R518 CSoutput.n317 CSoutput.t88 4.06363
R519 CSoutput.n315 CSoutput.t97 4.06363
R520 CSoutput.n315 CSoutput.t62 4.06363
R521 CSoutput.n313 CSoutput.t77 4.06363
R522 CSoutput.n313 CSoutput.t12 4.06363
R523 CSoutput.n311 CSoutput.t101 4.06363
R524 CSoutput.n311 CSoutput.t57 4.06363
R525 CSoutput.n309 CSoutput.t159 4.06363
R526 CSoutput.n309 CSoutput.t124 4.06363
R527 CSoutput.n308 CSoutput.t5 4.06363
R528 CSoutput.n308 CSoutput.t141 4.06363
R529 CSoutput.n305 CSoutput.t15 4.06363
R530 CSoutput.n305 CSoutput.t18 4.06363
R531 CSoutput.n303 CSoutput.t131 4.06363
R532 CSoutput.n303 CSoutput.t87 4.06363
R533 CSoutput.n301 CSoutput.t156 4.06363
R534 CSoutput.n301 CSoutput.t67 4.06363
R535 CSoutput.n299 CSoutput.t35 4.06363
R536 CSoutput.n299 CSoutput.t36 4.06363
R537 CSoutput.n297 CSoutput.t69 4.06363
R538 CSoutput.n297 CSoutput.t86 4.06363
R539 CSoutput.n295 CSoutput.t51 4.06363
R540 CSoutput.n295 CSoutput.t63 4.06363
R541 CSoutput.n293 CSoutput.t111 4.06363
R542 CSoutput.n293 CSoutput.t139 4.06363
R543 CSoutput.n292 CSoutput.t126 4.06363
R544 CSoutput.n292 CSoutput.t140 4.06363
R545 CSoutput.n290 CSoutput.t10 4.06363
R546 CSoutput.n290 CSoutput.t1 4.06363
R547 CSoutput.n288 CSoutput.t4 4.06363
R548 CSoutput.n288 CSoutput.t106 4.06363
R549 CSoutput.n286 CSoutput.t100 4.06363
R550 CSoutput.n286 CSoutput.t42 4.06363
R551 CSoutput.n284 CSoutput.t60 4.06363
R552 CSoutput.n284 CSoutput.t154 4.06363
R553 CSoutput.n282 CSoutput.t29 4.06363
R554 CSoutput.n282 CSoutput.t149 4.06363
R555 CSoutput.n280 CSoutput.t108 4.06363
R556 CSoutput.n280 CSoutput.t17 4.06363
R557 CSoutput.n278 CSoutput.t2 4.06363
R558 CSoutput.n278 CSoutput.t109 4.06363
R559 CSoutput.n277 CSoutput.t90 4.06363
R560 CSoutput.n277 CSoutput.t125 4.06363
R561 CSoutput.n110 CSoutput.t65 4.06363
R562 CSoutput.n110 CSoutput.t118 4.06363
R563 CSoutput.n111 CSoutput.t137 4.06363
R564 CSoutput.n111 CSoutput.t104 4.06363
R565 CSoutput.n113 CSoutput.t71 4.06363
R566 CSoutput.n113 CSoutput.t99 4.06363
R567 CSoutput.n115 CSoutput.t94 4.06363
R568 CSoutput.n115 CSoutput.t116 4.06363
R569 CSoutput.n117 CSoutput.t13 4.06363
R570 CSoutput.n117 CSoutput.t147 4.06363
R571 CSoutput.n119 CSoutput.t107 4.06363
R572 CSoutput.n119 CSoutput.t82 4.06363
R573 CSoutput.n121 CSoutput.t83 4.06363
R574 CSoutput.n121 CSoutput.t85 4.06363
R575 CSoutput.n123 CSoutput.t103 4.06363
R576 CSoutput.n123 CSoutput.t158 4.06363
R577 CSoutput.n94 CSoutput.t155 4.06363
R578 CSoutput.n94 CSoutput.t153 4.06363
R579 CSoutput.n95 CSoutput.t157 4.06363
R580 CSoutput.n95 CSoutput.t152 4.06363
R581 CSoutput.n97 CSoutput.t93 4.06363
R582 CSoutput.n97 CSoutput.t61 4.06363
R583 CSoutput.n99 CSoutput.t19 4.06363
R584 CSoutput.n99 CSoutput.t53 4.06363
R585 CSoutput.n101 CSoutput.t72 4.06363
R586 CSoutput.n101 CSoutput.t43 4.06363
R587 CSoutput.n103 CSoutput.t34 4.06363
R588 CSoutput.n103 CSoutput.t66 4.06363
R589 CSoutput.n105 CSoutput.t98 4.06363
R590 CSoutput.n105 CSoutput.t52 4.06363
R591 CSoutput.n107 CSoutput.t132 4.06363
R592 CSoutput.n107 CSoutput.t130 4.06363
R593 CSoutput.n79 CSoutput.t146 4.06363
R594 CSoutput.n79 CSoutput.t55 4.06363
R595 CSoutput.n80 CSoutput.t105 4.06363
R596 CSoutput.n80 CSoutput.t30 4.06363
R597 CSoutput.n82 CSoutput.t44 4.06363
R598 CSoutput.n82 CSoutput.t95 4.06363
R599 CSoutput.n84 CSoutput.t14 4.06363
R600 CSoutput.n84 CSoutput.t56 4.06363
R601 CSoutput.n86 CSoutput.t68 4.06363
R602 CSoutput.n86 CSoutput.t127 4.06363
R603 CSoutput.n88 CSoutput.t7 4.06363
R604 CSoutput.n88 CSoutput.t70 4.06363
R605 CSoutput.n90 CSoutput.t143 4.06363
R606 CSoutput.n90 CSoutput.t73 4.06363
R607 CSoutput.n92 CSoutput.t135 4.06363
R608 CSoutput.n92 CSoutput.t41 4.06363
R609 CSoutput.n44 CSoutput.n43 3.79402
R610 CSoutput.n49 CSoutput.n48 3.79402
R611 CSoutput.n389 CSoutput.n388 3.57343
R612 CSoutput.n388 CSoutput.n356 3.08965
R613 CSoutput.n353 CSoutput.t46 2.82907
R614 CSoutput.n353 CSoutput.t74 2.82907
R615 CSoutput.n351 CSoutput.t122 2.82907
R616 CSoutput.n351 CSoutput.t26 2.82907
R617 CSoutput.n349 CSoutput.t0 2.82907
R618 CSoutput.n349 CSoutput.t76 2.82907
R619 CSoutput.n347 CSoutput.t40 2.82907
R620 CSoutput.n347 CSoutput.t78 2.82907
R621 CSoutput.n345 CSoutput.t80 2.82907
R622 CSoutput.n345 CSoutput.t119 2.82907
R623 CSoutput.n343 CSoutput.t59 2.82907
R624 CSoutput.n343 CSoutput.t32 2.82907
R625 CSoutput.n341 CSoutput.t49 2.82907
R626 CSoutput.n341 CSoutput.t133 2.82907
R627 CSoutput.n340 CSoutput.t22 2.82907
R628 CSoutput.n340 CSoutput.t33 2.82907
R629 CSoutput.n338 CSoutput.t6 2.82907
R630 CSoutput.n338 CSoutput.t148 2.82907
R631 CSoutput.n336 CSoutput.t64 2.82907
R632 CSoutput.n336 CSoutput.t123 2.82907
R633 CSoutput.n334 CSoutput.t134 2.82907
R634 CSoutput.n334 CSoutput.t112 2.82907
R635 CSoutput.n332 CSoutput.t136 2.82907
R636 CSoutput.n332 CSoutput.t138 2.82907
R637 CSoutput.n330 CSoutput.t48 2.82907
R638 CSoutput.n330 CSoutput.t96 2.82907
R639 CSoutput.n328 CSoutput.t114 2.82907
R640 CSoutput.n328 CSoutput.t142 2.82907
R641 CSoutput.n326 CSoutput.t115 2.82907
R642 CSoutput.n326 CSoutput.t120 2.82907
R643 CSoutput.n325 CSoutput.t9 2.82907
R644 CSoutput.n325 CSoutput.t31 2.82907
R645 CSoutput.n372 CSoutput.t84 2.82907
R646 CSoutput.n372 CSoutput.t45 2.82907
R647 CSoutput.n373 CSoutput.t54 2.82907
R648 CSoutput.n373 CSoutput.t50 2.82907
R649 CSoutput.n375 CSoutput.t23 2.82907
R650 CSoutput.n375 CSoutput.t11 2.82907
R651 CSoutput.n377 CSoutput.t21 2.82907
R652 CSoutput.n377 CSoutput.t113 2.82907
R653 CSoutput.n379 CSoutput.t110 2.82907
R654 CSoutput.n379 CSoutput.t3 2.82907
R655 CSoutput.n381 CSoutput.t58 2.82907
R656 CSoutput.n381 CSoutput.t144 2.82907
R657 CSoutput.n383 CSoutput.t81 2.82907
R658 CSoutput.n383 CSoutput.t37 2.82907
R659 CSoutput.n385 CSoutput.t39 2.82907
R660 CSoutput.n385 CSoutput.t79 2.82907
R661 CSoutput.n357 CSoutput.t91 2.82907
R662 CSoutput.n357 CSoutput.t92 2.82907
R663 CSoutput.n358 CSoutput.t27 2.82907
R664 CSoutput.n358 CSoutput.t117 2.82907
R665 CSoutput.n360 CSoutput.t89 2.82907
R666 CSoutput.n360 CSoutput.t24 2.82907
R667 CSoutput.n362 CSoutput.t102 2.82907
R668 CSoutput.n362 CSoutput.t128 2.82907
R669 CSoutput.n364 CSoutput.t75 2.82907
R670 CSoutput.n364 CSoutput.t25 2.82907
R671 CSoutput.n366 CSoutput.t20 2.82907
R672 CSoutput.n366 CSoutput.t8 2.82907
R673 CSoutput.n368 CSoutput.t129 2.82907
R674 CSoutput.n368 CSoutput.t47 2.82907
R675 CSoutput.n370 CSoutput.t38 2.82907
R676 CSoutput.n370 CSoutput.t121 2.82907
R677 CSoutput.n75 CSoutput.n1 2.45513
R678 CSoutput.n324 CSoutput.n126 2.36742
R679 CSoutput.n217 CSoutput.n215 2.251
R680 CSoutput.n217 CSoutput.n214 2.251
R681 CSoutput.n217 CSoutput.n213 2.251
R682 CSoutput.n217 CSoutput.n212 2.251
R683 CSoutput.n186 CSoutput.n185 2.251
R684 CSoutput.n186 CSoutput.n184 2.251
R685 CSoutput.n186 CSoutput.n183 2.251
R686 CSoutput.n186 CSoutput.n182 2.251
R687 CSoutput.n259 CSoutput.n258 2.251
R688 CSoutput.n224 CSoutput.n222 2.251
R689 CSoutput.n224 CSoutput.n221 2.251
R690 CSoutput.n224 CSoutput.n220 2.251
R691 CSoutput.n242 CSoutput.n224 2.251
R692 CSoutput.n230 CSoutput.n229 2.251
R693 CSoutput.n230 CSoutput.n228 2.251
R694 CSoutput.n230 CSoutput.n227 2.251
R695 CSoutput.n230 CSoutput.n226 2.251
R696 CSoutput.n256 CSoutput.n196 2.251
R697 CSoutput.n251 CSoutput.n249 2.251
R698 CSoutput.n251 CSoutput.n248 2.251
R699 CSoutput.n251 CSoutput.n247 2.251
R700 CSoutput.n251 CSoutput.n246 2.251
R701 CSoutput.n152 CSoutput.n151 2.251
R702 CSoutput.n152 CSoutput.n150 2.251
R703 CSoutput.n152 CSoutput.n149 2.251
R704 CSoutput.n152 CSoutput.n148 2.251
R705 CSoutput.n269 CSoutput.n268 2.251
R706 CSoutput.n186 CSoutput.n166 2.2505
R707 CSoutput.n181 CSoutput.n166 2.2505
R708 CSoutput.n179 CSoutput.n166 2.2505
R709 CSoutput.n178 CSoutput.n166 2.2505
R710 CSoutput.n263 CSoutput.n166 2.2505
R711 CSoutput.n261 CSoutput.n166 2.2505
R712 CSoutput.n259 CSoutput.n166 2.2505
R713 CSoutput.n189 CSoutput.n166 2.2505
R714 CSoutput.n188 CSoutput.n166 2.2505
R715 CSoutput.n192 CSoutput.n166 2.2505
R716 CSoutput.n191 CSoutput.n166 2.2505
R717 CSoutput.n174 CSoutput.n166 2.2505
R718 CSoutput.n266 CSoutput.n166 2.2505
R719 CSoutput.n266 CSoutput.n265 2.2505
R720 CSoutput.n230 CSoutput.n201 2.2505
R721 CSoutput.n211 CSoutput.n201 2.2505
R722 CSoutput.n232 CSoutput.n201 2.2505
R723 CSoutput.n210 CSoutput.n201 2.2505
R724 CSoutput.n234 CSoutput.n201 2.2505
R725 CSoutput.n201 CSoutput.n195 2.2505
R726 CSoutput.n256 CSoutput.n201 2.2505
R727 CSoutput.n254 CSoutput.n201 2.2505
R728 CSoutput.n236 CSoutput.n201 2.2505
R729 CSoutput.n208 CSoutput.n201 2.2505
R730 CSoutput.n238 CSoutput.n201 2.2505
R731 CSoutput.n207 CSoutput.n201 2.2505
R732 CSoutput.n252 CSoutput.n201 2.2505
R733 CSoutput.n252 CSoutput.n205 2.2505
R734 CSoutput.n152 CSoutput.n132 2.2505
R735 CSoutput.n147 CSoutput.n132 2.2505
R736 CSoutput.n145 CSoutput.n132 2.2505
R737 CSoutput.n144 CSoutput.n132 2.2505
R738 CSoutput.n273 CSoutput.n132 2.2505
R739 CSoutput.n271 CSoutput.n132 2.2505
R740 CSoutput.n269 CSoutput.n132 2.2505
R741 CSoutput.n155 CSoutput.n132 2.2505
R742 CSoutput.n154 CSoutput.n132 2.2505
R743 CSoutput.n158 CSoutput.n132 2.2505
R744 CSoutput.n157 CSoutput.n132 2.2505
R745 CSoutput.n140 CSoutput.n132 2.2505
R746 CSoutput.n276 CSoutput.n132 2.2505
R747 CSoutput.n276 CSoutput.n275 2.2505
R748 CSoutput.n194 CSoutput.n187 2.25024
R749 CSoutput.n194 CSoutput.n180 2.25024
R750 CSoutput.n262 CSoutput.n194 2.25024
R751 CSoutput.n194 CSoutput.n190 2.25024
R752 CSoutput.n194 CSoutput.n193 2.25024
R753 CSoutput.n194 CSoutput.n161 2.25024
R754 CSoutput.n244 CSoutput.n241 2.25024
R755 CSoutput.n244 CSoutput.n240 2.25024
R756 CSoutput.n244 CSoutput.n239 2.25024
R757 CSoutput.n244 CSoutput.n206 2.25024
R758 CSoutput.n244 CSoutput.n243 2.25024
R759 CSoutput.n245 CSoutput.n244 2.25024
R760 CSoutput.n160 CSoutput.n153 2.25024
R761 CSoutput.n160 CSoutput.n146 2.25024
R762 CSoutput.n272 CSoutput.n160 2.25024
R763 CSoutput.n160 CSoutput.n156 2.25024
R764 CSoutput.n160 CSoutput.n159 2.25024
R765 CSoutput.n160 CSoutput.n127 2.25024
R766 CSoutput.n261 CSoutput.n171 1.50111
R767 CSoutput.n209 CSoutput.n195 1.50111
R768 CSoutput.n271 CSoutput.n137 1.50111
R769 CSoutput.n217 CSoutput.n216 1.501
R770 CSoutput.n224 CSoutput.n223 1.501
R771 CSoutput.n251 CSoutput.n250 1.501
R772 CSoutput.n265 CSoutput.n176 1.12536
R773 CSoutput.n265 CSoutput.n177 1.12536
R774 CSoutput.n265 CSoutput.n264 1.12536
R775 CSoutput.n225 CSoutput.n205 1.12536
R776 CSoutput.n231 CSoutput.n205 1.12536
R777 CSoutput.n233 CSoutput.n205 1.12536
R778 CSoutput.n275 CSoutput.n142 1.12536
R779 CSoutput.n275 CSoutput.n143 1.12536
R780 CSoutput.n275 CSoutput.n274 1.12536
R781 CSoutput.n265 CSoutput.n172 1.12536
R782 CSoutput.n265 CSoutput.n173 1.12536
R783 CSoutput.n265 CSoutput.n175 1.12536
R784 CSoutput.n255 CSoutput.n205 1.12536
R785 CSoutput.n235 CSoutput.n205 1.12536
R786 CSoutput.n237 CSoutput.n205 1.12536
R787 CSoutput.n275 CSoutput.n138 1.12536
R788 CSoutput.n275 CSoutput.n139 1.12536
R789 CSoutput.n275 CSoutput.n141 1.12536
R790 CSoutput.n31 CSoutput.n30 0.669944
R791 CSoutput.n62 CSoutput.n61 0.669944
R792 CSoutput.n344 CSoutput.n342 0.573776
R793 CSoutput.n346 CSoutput.n344 0.573776
R794 CSoutput.n348 CSoutput.n346 0.573776
R795 CSoutput.n350 CSoutput.n348 0.573776
R796 CSoutput.n352 CSoutput.n350 0.573776
R797 CSoutput.n354 CSoutput.n352 0.573776
R798 CSoutput.n329 CSoutput.n327 0.573776
R799 CSoutput.n331 CSoutput.n329 0.573776
R800 CSoutput.n333 CSoutput.n331 0.573776
R801 CSoutput.n335 CSoutput.n333 0.573776
R802 CSoutput.n337 CSoutput.n335 0.573776
R803 CSoutput.n339 CSoutput.n337 0.573776
R804 CSoutput.n386 CSoutput.n384 0.573776
R805 CSoutput.n384 CSoutput.n382 0.573776
R806 CSoutput.n382 CSoutput.n380 0.573776
R807 CSoutput.n380 CSoutput.n378 0.573776
R808 CSoutput.n378 CSoutput.n376 0.573776
R809 CSoutput.n376 CSoutput.n374 0.573776
R810 CSoutput.n371 CSoutput.n369 0.573776
R811 CSoutput.n369 CSoutput.n367 0.573776
R812 CSoutput.n367 CSoutput.n365 0.573776
R813 CSoutput.n365 CSoutput.n363 0.573776
R814 CSoutput.n363 CSoutput.n361 0.573776
R815 CSoutput.n361 CSoutput.n359 0.573776
R816 CSoutput.n389 CSoutput.n276 0.53442
R817 CSoutput.n312 CSoutput.n310 0.358259
R818 CSoutput.n314 CSoutput.n312 0.358259
R819 CSoutput.n316 CSoutput.n314 0.358259
R820 CSoutput.n318 CSoutput.n316 0.358259
R821 CSoutput.n320 CSoutput.n318 0.358259
R822 CSoutput.n322 CSoutput.n320 0.358259
R823 CSoutput.n296 CSoutput.n294 0.358259
R824 CSoutput.n298 CSoutput.n296 0.358259
R825 CSoutput.n300 CSoutput.n298 0.358259
R826 CSoutput.n302 CSoutput.n300 0.358259
R827 CSoutput.n304 CSoutput.n302 0.358259
R828 CSoutput.n306 CSoutput.n304 0.358259
R829 CSoutput.n281 CSoutput.n279 0.358259
R830 CSoutput.n283 CSoutput.n281 0.358259
R831 CSoutput.n285 CSoutput.n283 0.358259
R832 CSoutput.n287 CSoutput.n285 0.358259
R833 CSoutput.n289 CSoutput.n287 0.358259
R834 CSoutput.n291 CSoutput.n289 0.358259
R835 CSoutput.n124 CSoutput.n122 0.358259
R836 CSoutput.n122 CSoutput.n120 0.358259
R837 CSoutput.n120 CSoutput.n118 0.358259
R838 CSoutput.n118 CSoutput.n116 0.358259
R839 CSoutput.n116 CSoutput.n114 0.358259
R840 CSoutput.n114 CSoutput.n112 0.358259
R841 CSoutput.n108 CSoutput.n106 0.358259
R842 CSoutput.n106 CSoutput.n104 0.358259
R843 CSoutput.n104 CSoutput.n102 0.358259
R844 CSoutput.n102 CSoutput.n100 0.358259
R845 CSoutput.n100 CSoutput.n98 0.358259
R846 CSoutput.n98 CSoutput.n96 0.358259
R847 CSoutput.n93 CSoutput.n91 0.358259
R848 CSoutput.n91 CSoutput.n89 0.358259
R849 CSoutput.n89 CSoutput.n87 0.358259
R850 CSoutput.n87 CSoutput.n85 0.358259
R851 CSoutput.n85 CSoutput.n83 0.358259
R852 CSoutput.n83 CSoutput.n81 0.358259
R853 CSoutput.n21 CSoutput.n20 0.169105
R854 CSoutput.n21 CSoutput.n16 0.169105
R855 CSoutput.n26 CSoutput.n16 0.169105
R856 CSoutput.n27 CSoutput.n26 0.169105
R857 CSoutput.n27 CSoutput.n14 0.169105
R858 CSoutput.n32 CSoutput.n14 0.169105
R859 CSoutput.n33 CSoutput.n32 0.169105
R860 CSoutput.n34 CSoutput.n33 0.169105
R861 CSoutput.n34 CSoutput.n12 0.169105
R862 CSoutput.n39 CSoutput.n12 0.169105
R863 CSoutput.n40 CSoutput.n39 0.169105
R864 CSoutput.n40 CSoutput.n10 0.169105
R865 CSoutput.n45 CSoutput.n10 0.169105
R866 CSoutput.n46 CSoutput.n45 0.169105
R867 CSoutput.n47 CSoutput.n46 0.169105
R868 CSoutput.n47 CSoutput.n8 0.169105
R869 CSoutput.n52 CSoutput.n8 0.169105
R870 CSoutput.n53 CSoutput.n52 0.169105
R871 CSoutput.n53 CSoutput.n6 0.169105
R872 CSoutput.n58 CSoutput.n6 0.169105
R873 CSoutput.n59 CSoutput.n58 0.169105
R874 CSoutput.n60 CSoutput.n59 0.169105
R875 CSoutput.n60 CSoutput.n4 0.169105
R876 CSoutput.n66 CSoutput.n4 0.169105
R877 CSoutput.n67 CSoutput.n66 0.169105
R878 CSoutput.n68 CSoutput.n67 0.169105
R879 CSoutput.n68 CSoutput.n2 0.169105
R880 CSoutput.n73 CSoutput.n2 0.169105
R881 CSoutput.n74 CSoutput.n73 0.169105
R882 CSoutput.n74 CSoutput.n0 0.169105
R883 CSoutput.n78 CSoutput.n0 0.169105
R884 CSoutput.n219 CSoutput.n218 0.0910737
R885 CSoutput.n270 CSoutput.n267 0.0723685
R886 CSoutput.n224 CSoutput.n219 0.0522944
R887 CSoutput.n267 CSoutput.n266 0.0499135
R888 CSoutput.n218 CSoutput.n217 0.0499135
R889 CSoutput.n252 CSoutput.n251 0.0464294
R890 CSoutput.n260 CSoutput.n257 0.0391444
R891 CSoutput.n219 CSoutput.t169 0.023435
R892 CSoutput.n267 CSoutput.t163 0.02262
R893 CSoutput.n218 CSoutput.t167 0.02262
R894 CSoutput CSoutput.n389 0.0052
R895 CSoutput.n189 CSoutput.n172 0.00365111
R896 CSoutput.n192 CSoutput.n173 0.00365111
R897 CSoutput.n175 CSoutput.n174 0.00365111
R898 CSoutput.n217 CSoutput.n176 0.00365111
R899 CSoutput.n181 CSoutput.n177 0.00365111
R900 CSoutput.n264 CSoutput.n178 0.00365111
R901 CSoutput.n255 CSoutput.n254 0.00365111
R902 CSoutput.n235 CSoutput.n208 0.00365111
R903 CSoutput.n237 CSoutput.n207 0.00365111
R904 CSoutput.n225 CSoutput.n224 0.00365111
R905 CSoutput.n231 CSoutput.n211 0.00365111
R906 CSoutput.n233 CSoutput.n210 0.00365111
R907 CSoutput.n155 CSoutput.n138 0.00365111
R908 CSoutput.n158 CSoutput.n139 0.00365111
R909 CSoutput.n141 CSoutput.n140 0.00365111
R910 CSoutput.n251 CSoutput.n142 0.00365111
R911 CSoutput.n147 CSoutput.n143 0.00365111
R912 CSoutput.n274 CSoutput.n144 0.00365111
R913 CSoutput.n186 CSoutput.n176 0.00340054
R914 CSoutput.n179 CSoutput.n177 0.00340054
R915 CSoutput.n264 CSoutput.n263 0.00340054
R916 CSoutput.n259 CSoutput.n172 0.00340054
R917 CSoutput.n188 CSoutput.n173 0.00340054
R918 CSoutput.n191 CSoutput.n175 0.00340054
R919 CSoutput.n230 CSoutput.n225 0.00340054
R920 CSoutput.n232 CSoutput.n231 0.00340054
R921 CSoutput.n234 CSoutput.n233 0.00340054
R922 CSoutput.n256 CSoutput.n255 0.00340054
R923 CSoutput.n236 CSoutput.n235 0.00340054
R924 CSoutput.n238 CSoutput.n237 0.00340054
R925 CSoutput.n152 CSoutput.n142 0.00340054
R926 CSoutput.n145 CSoutput.n143 0.00340054
R927 CSoutput.n274 CSoutput.n273 0.00340054
R928 CSoutput.n269 CSoutput.n138 0.00340054
R929 CSoutput.n154 CSoutput.n139 0.00340054
R930 CSoutput.n157 CSoutput.n141 0.00340054
R931 CSoutput.n187 CSoutput.n181 0.00252698
R932 CSoutput.n180 CSoutput.n178 0.00252698
R933 CSoutput.n262 CSoutput.n261 0.00252698
R934 CSoutput.n190 CSoutput.n188 0.00252698
R935 CSoutput.n193 CSoutput.n191 0.00252698
R936 CSoutput.n266 CSoutput.n161 0.00252698
R937 CSoutput.n187 CSoutput.n186 0.00252698
R938 CSoutput.n180 CSoutput.n179 0.00252698
R939 CSoutput.n263 CSoutput.n262 0.00252698
R940 CSoutput.n190 CSoutput.n189 0.00252698
R941 CSoutput.n193 CSoutput.n192 0.00252698
R942 CSoutput.n174 CSoutput.n161 0.00252698
R943 CSoutput.n241 CSoutput.n211 0.00252698
R944 CSoutput.n240 CSoutput.n210 0.00252698
R945 CSoutput.n239 CSoutput.n195 0.00252698
R946 CSoutput.n236 CSoutput.n206 0.00252698
R947 CSoutput.n243 CSoutput.n238 0.00252698
R948 CSoutput.n252 CSoutput.n245 0.00252698
R949 CSoutput.n241 CSoutput.n230 0.00252698
R950 CSoutput.n240 CSoutput.n232 0.00252698
R951 CSoutput.n239 CSoutput.n234 0.00252698
R952 CSoutput.n254 CSoutput.n206 0.00252698
R953 CSoutput.n243 CSoutput.n208 0.00252698
R954 CSoutput.n245 CSoutput.n207 0.00252698
R955 CSoutput.n153 CSoutput.n147 0.00252698
R956 CSoutput.n146 CSoutput.n144 0.00252698
R957 CSoutput.n272 CSoutput.n271 0.00252698
R958 CSoutput.n156 CSoutput.n154 0.00252698
R959 CSoutput.n159 CSoutput.n157 0.00252698
R960 CSoutput.n276 CSoutput.n127 0.00252698
R961 CSoutput.n153 CSoutput.n152 0.00252698
R962 CSoutput.n146 CSoutput.n145 0.00252698
R963 CSoutput.n273 CSoutput.n272 0.00252698
R964 CSoutput.n156 CSoutput.n155 0.00252698
R965 CSoutput.n159 CSoutput.n158 0.00252698
R966 CSoutput.n140 CSoutput.n127 0.00252698
R967 CSoutput.n261 CSoutput.n260 0.0020275
R968 CSoutput.n260 CSoutput.n259 0.0020275
R969 CSoutput.n257 CSoutput.n195 0.0020275
R970 CSoutput.n257 CSoutput.n256 0.0020275
R971 CSoutput.n271 CSoutput.n270 0.0020275
R972 CSoutput.n270 CSoutput.n269 0.0020275
R973 CSoutput.n171 CSoutput.n170 0.00166668
R974 CSoutput.n253 CSoutput.n209 0.00166668
R975 CSoutput.n137 CSoutput.n136 0.00166668
R976 CSoutput.n275 CSoutput.n137 0.00133328
R977 CSoutput.n209 CSoutput.n205 0.00133328
R978 CSoutput.n265 CSoutput.n171 0.00133328
R979 CSoutput.n268 CSoutput.n160 0.001
R980 CSoutput.n246 CSoutput.n160 0.001
R981 CSoutput.n148 CSoutput.n128 0.001
R982 CSoutput.n247 CSoutput.n128 0.001
R983 CSoutput.n149 CSoutput.n129 0.001
R984 CSoutput.n248 CSoutput.n129 0.001
R985 CSoutput.n150 CSoutput.n130 0.001
R986 CSoutput.n249 CSoutput.n130 0.001
R987 CSoutput.n151 CSoutput.n131 0.001
R988 CSoutput.n250 CSoutput.n131 0.001
R989 CSoutput.n244 CSoutput.n196 0.001
R990 CSoutput.n244 CSoutput.n242 0.001
R991 CSoutput.n226 CSoutput.n197 0.001
R992 CSoutput.n220 CSoutput.n197 0.001
R993 CSoutput.n227 CSoutput.n198 0.001
R994 CSoutput.n221 CSoutput.n198 0.001
R995 CSoutput.n228 CSoutput.n199 0.001
R996 CSoutput.n222 CSoutput.n199 0.001
R997 CSoutput.n229 CSoutput.n200 0.001
R998 CSoutput.n223 CSoutput.n200 0.001
R999 CSoutput.n258 CSoutput.n194 0.001
R1000 CSoutput.n212 CSoutput.n194 0.001
R1001 CSoutput.n182 CSoutput.n162 0.001
R1002 CSoutput.n213 CSoutput.n162 0.001
R1003 CSoutput.n183 CSoutput.n163 0.001
R1004 CSoutput.n214 CSoutput.n163 0.001
R1005 CSoutput.n184 CSoutput.n164 0.001
R1006 CSoutput.n215 CSoutput.n164 0.001
R1007 CSoutput.n185 CSoutput.n165 0.001
R1008 CSoutput.n216 CSoutput.n165 0.001
R1009 CSoutput.n216 CSoutput.n166 0.001
R1010 CSoutput.n215 CSoutput.n167 0.001
R1011 CSoutput.n214 CSoutput.n168 0.001
R1012 CSoutput.n213 CSoutput.t180 0.001
R1013 CSoutput.n212 CSoutput.n169 0.001
R1014 CSoutput.n185 CSoutput.n167 0.001
R1015 CSoutput.n184 CSoutput.n168 0.001
R1016 CSoutput.n183 CSoutput.t180 0.001
R1017 CSoutput.n182 CSoutput.n169 0.001
R1018 CSoutput.n258 CSoutput.n170 0.001
R1019 CSoutput.n223 CSoutput.n201 0.001
R1020 CSoutput.n222 CSoutput.n202 0.001
R1021 CSoutput.n221 CSoutput.n203 0.001
R1022 CSoutput.n220 CSoutput.t160 0.001
R1023 CSoutput.n242 CSoutput.n204 0.001
R1024 CSoutput.n229 CSoutput.n202 0.001
R1025 CSoutput.n228 CSoutput.n203 0.001
R1026 CSoutput.n227 CSoutput.t160 0.001
R1027 CSoutput.n226 CSoutput.n204 0.001
R1028 CSoutput.n253 CSoutput.n196 0.001
R1029 CSoutput.n250 CSoutput.n132 0.001
R1030 CSoutput.n249 CSoutput.n133 0.001
R1031 CSoutput.n248 CSoutput.n134 0.001
R1032 CSoutput.n247 CSoutput.t168 0.001
R1033 CSoutput.n246 CSoutput.n135 0.001
R1034 CSoutput.n151 CSoutput.n133 0.001
R1035 CSoutput.n150 CSoutput.n134 0.001
R1036 CSoutput.n149 CSoutput.t168 0.001
R1037 CSoutput.n148 CSoutput.n135 0.001
R1038 CSoutput.n268 CSoutput.n136 0.001
R1039 a_n1986_8322.n2 a_n1986_8322.t12 74.6477
R1040 a_n1986_8322.n1 a_n1986_8322.t5 74.6477
R1041 a_n1986_8322.n0 a_n1986_8322.t10 74.6474
R1042 a_n1986_8322.n2 a_n1986_8322.t18 74.2899
R1043 a_n1986_8322.n2 a_n1986_8322.t20 74.2899
R1044 a_n1986_8322.n3 a_n1986_8322.t3 74.2899
R1045 a_n1986_8322.n6 a_n1986_8322.t14 74.2899
R1046 a_n1986_8322.n10 a_n1986_8322.t17 74.2899
R1047 a_n1986_8322.n2 a_n1986_8322.n12 70.6783
R1048 a_n1986_8322.n0 a_n1986_8322.n4 70.6783
R1049 a_n1986_8322.n0 a_n1986_8322.n5 70.6783
R1050 a_n1986_8322.n1 a_n1986_8322.n8 70.6783
R1051 a_n1986_8322.n1 a_n1986_8322.n9 70.6783
R1052 a_n1986_8322.n13 a_n1986_8322.n3 70.6782
R1053 a_n1986_8322.n11 a_n1986_8322.n10 22.7556
R1054 a_n1986_8322.n7 a_n1986_8322.t16 9.96389
R1055 a_n1986_8322.n3 a_n1986_8322.n11 6.2408
R1056 a_n1986_8322.n7 a_n1986_8322.n6 5.83671
R1057 a_n1986_8322.n11 a_n1986_8322.n7 5.3452
R1058 a_n1986_8322.n12 a_n1986_8322.t7 3.61217
R1059 a_n1986_8322.n12 a_n1986_8322.t4 3.61217
R1060 a_n1986_8322.n4 a_n1986_8322.t2 3.61217
R1061 a_n1986_8322.n4 a_n1986_8322.t8 3.61217
R1062 a_n1986_8322.n5 a_n1986_8322.t15 3.61217
R1063 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R1064 a_n1986_8322.n8 a_n1986_8322.t6 3.61217
R1065 a_n1986_8322.n8 a_n1986_8322.t1 3.61217
R1066 a_n1986_8322.n9 a_n1986_8322.t19 3.61217
R1067 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R1068 a_n1986_8322.t0 a_n1986_8322.n13 3.61217
R1069 a_n1986_8322.n13 a_n1986_8322.t13 3.61217
R1070 a_n1986_8322.n3 a_n1986_8322.n2 1.17507
R1071 a_n1986_8322.n10 a_n1986_8322.n1 0.716017
R1072 a_n1986_8322.n6 a_n1986_8322.n0 0.716017
R1073 commonsourceibias.n35 commonsourceibias.t34 223.028
R1074 commonsourceibias.n128 commonsourceibias.t88 223.028
R1075 commonsourceibias.n217 commonsourceibias.t77 223.028
R1076 commonsourceibias.n364 commonsourceibias.t30 223.028
R1077 commonsourceibias.n305 commonsourceibias.t108 223.028
R1078 commonsourceibias.n499 commonsourceibias.t95 223.028
R1079 commonsourceibias.n99 commonsourceibias.t48 207.983
R1080 commonsourceibias.n192 commonsourceibias.t94 207.983
R1081 commonsourceibias.n281 commonsourceibias.t81 207.983
R1082 commonsourceibias.n430 commonsourceibias.t2 207.983
R1083 commonsourceibias.n476 commonsourceibias.t113 207.983
R1084 commonsourceibias.n565 commonsourceibias.t99 207.983
R1085 commonsourceibias.n97 commonsourceibias.t18 168.701
R1086 commonsourceibias.n91 commonsourceibias.t12 168.701
R1087 commonsourceibias.n17 commonsourceibias.t46 168.701
R1088 commonsourceibias.n83 commonsourceibias.t24 168.701
R1089 commonsourceibias.n77 commonsourceibias.t52 168.701
R1090 commonsourceibias.n22 commonsourceibias.t60 168.701
R1091 commonsourceibias.n69 commonsourceibias.t14 168.701
R1092 commonsourceibias.n63 commonsourceibias.t50 168.701
R1093 commonsourceibias.n25 commonsourceibias.t42 168.701
R1094 commonsourceibias.n27 commonsourceibias.t56 168.701
R1095 commonsourceibias.n29 commonsourceibias.t62 168.701
R1096 commonsourceibias.n46 commonsourceibias.t10 168.701
R1097 commonsourceibias.n40 commonsourceibias.t28 168.701
R1098 commonsourceibias.n34 commonsourceibias.t20 168.701
R1099 commonsourceibias.n190 commonsourceibias.t109 168.701
R1100 commonsourceibias.n184 commonsourceibias.t72 168.701
R1101 commonsourceibias.n5 commonsourceibias.t70 168.701
R1102 commonsourceibias.n176 commonsourceibias.t102 168.701
R1103 commonsourceibias.n170 commonsourceibias.t116 168.701
R1104 commonsourceibias.n10 commonsourceibias.t66 168.701
R1105 commonsourceibias.n162 commonsourceibias.t92 168.701
R1106 commonsourceibias.n156 commonsourceibias.t89 168.701
R1107 commonsourceibias.n118 commonsourceibias.t105 168.701
R1108 commonsourceibias.n120 commonsourceibias.t85 168.701
R1109 commonsourceibias.n122 commonsourceibias.t82 168.701
R1110 commonsourceibias.n139 commonsourceibias.t97 168.701
R1111 commonsourceibias.n133 commonsourceibias.t111 168.701
R1112 commonsourceibias.n127 commonsourceibias.t75 168.701
R1113 commonsourceibias.n216 commonsourceibias.t67 168.701
R1114 commonsourceibias.n222 commonsourceibias.t98 168.701
R1115 commonsourceibias.n228 commonsourceibias.t83 168.701
R1116 commonsourceibias.n211 commonsourceibias.t71 168.701
R1117 commonsourceibias.n209 commonsourceibias.t74 168.701
R1118 commonsourceibias.n207 commonsourceibias.t90 168.701
R1119 commonsourceibias.n245 commonsourceibias.t76 168.701
R1120 commonsourceibias.n251 commonsourceibias.t80 168.701
R1121 commonsourceibias.n204 commonsourceibias.t122 168.701
R1122 commonsourceibias.n259 commonsourceibias.t104 168.701
R1123 commonsourceibias.n265 commonsourceibias.t87 168.701
R1124 commonsourceibias.n199 commonsourceibias.t127 168.701
R1125 commonsourceibias.n273 commonsourceibias.t65 168.701
R1126 commonsourceibias.n279 commonsourceibias.t96 168.701
R1127 commonsourceibias.n363 commonsourceibias.t32 168.701
R1128 commonsourceibias.n369 commonsourceibias.t38 168.701
R1129 commonsourceibias.n375 commonsourceibias.t36 168.701
R1130 commonsourceibias.n358 commonsourceibias.t8 168.701
R1131 commonsourceibias.n356 commonsourceibias.t40 168.701
R1132 commonsourceibias.n354 commonsourceibias.t22 168.701
R1133 commonsourceibias.n392 commonsourceibias.t4 168.701
R1134 commonsourceibias.n398 commonsourceibias.t58 168.701
R1135 commonsourceibias.n400 commonsourceibias.t44 168.701
R1136 commonsourceibias.n407 commonsourceibias.t6 168.701
R1137 commonsourceibias.n413 commonsourceibias.t16 168.701
R1138 commonsourceibias.n415 commonsourceibias.t0 168.701
R1139 commonsourceibias.n422 commonsourceibias.t54 168.701
R1140 commonsourceibias.n428 commonsourceibias.t26 168.701
R1141 commonsourceibias.n474 commonsourceibias.t123 168.701
R1142 commonsourceibias.n468 commonsourceibias.t68 168.701
R1143 commonsourceibias.n461 commonsourceibias.t84 168.701
R1144 commonsourceibias.n459 commonsourceibias.t119 168.701
R1145 commonsourceibias.n453 commonsourceibias.t64 168.701
R1146 commonsourceibias.n446 commonsourceibias.t126 168.701
R1147 commonsourceibias.n444 commonsourceibias.t112 168.701
R1148 commonsourceibias.n304 commonsourceibias.t91 168.701
R1149 commonsourceibias.n310 commonsourceibias.t125 168.701
R1150 commonsourceibias.n316 commonsourceibias.t115 168.701
R1151 commonsourceibias.n299 commonsourceibias.t101 168.701
R1152 commonsourceibias.n297 commonsourceibias.t78 168.701
R1153 commonsourceibias.n295 commonsourceibias.t121 168.701
R1154 commonsourceibias.n333 commonsourceibias.t107 168.701
R1155 commonsourceibias.n498 commonsourceibias.t79 168.701
R1156 commonsourceibias.n504 commonsourceibias.t118 168.701
R1157 commonsourceibias.n510 commonsourceibias.t103 168.701
R1158 commonsourceibias.n493 commonsourceibias.t86 168.701
R1159 commonsourceibias.n491 commonsourceibias.t69 168.701
R1160 commonsourceibias.n489 commonsourceibias.t110 168.701
R1161 commonsourceibias.n527 commonsourceibias.t93 168.701
R1162 commonsourceibias.n533 commonsourceibias.t100 168.701
R1163 commonsourceibias.n535 commonsourceibias.t117 168.701
R1164 commonsourceibias.n542 commonsourceibias.t120 168.701
R1165 commonsourceibias.n548 commonsourceibias.t106 168.701
R1166 commonsourceibias.n550 commonsourceibias.t73 168.701
R1167 commonsourceibias.n557 commonsourceibias.t124 168.701
R1168 commonsourceibias.n563 commonsourceibias.t114 168.701
R1169 commonsourceibias.n36 commonsourceibias.n33 161.3
R1170 commonsourceibias.n38 commonsourceibias.n37 161.3
R1171 commonsourceibias.n39 commonsourceibias.n32 161.3
R1172 commonsourceibias.n42 commonsourceibias.n41 161.3
R1173 commonsourceibias.n43 commonsourceibias.n31 161.3
R1174 commonsourceibias.n45 commonsourceibias.n44 161.3
R1175 commonsourceibias.n47 commonsourceibias.n30 161.3
R1176 commonsourceibias.n49 commonsourceibias.n48 161.3
R1177 commonsourceibias.n51 commonsourceibias.n50 161.3
R1178 commonsourceibias.n52 commonsourceibias.n28 161.3
R1179 commonsourceibias.n54 commonsourceibias.n53 161.3
R1180 commonsourceibias.n56 commonsourceibias.n55 161.3
R1181 commonsourceibias.n57 commonsourceibias.n26 161.3
R1182 commonsourceibias.n59 commonsourceibias.n58 161.3
R1183 commonsourceibias.n61 commonsourceibias.n60 161.3
R1184 commonsourceibias.n62 commonsourceibias.n24 161.3
R1185 commonsourceibias.n65 commonsourceibias.n64 161.3
R1186 commonsourceibias.n66 commonsourceibias.n23 161.3
R1187 commonsourceibias.n68 commonsourceibias.n67 161.3
R1188 commonsourceibias.n70 commonsourceibias.n21 161.3
R1189 commonsourceibias.n72 commonsourceibias.n71 161.3
R1190 commonsourceibias.n73 commonsourceibias.n20 161.3
R1191 commonsourceibias.n75 commonsourceibias.n74 161.3
R1192 commonsourceibias.n76 commonsourceibias.n19 161.3
R1193 commonsourceibias.n79 commonsourceibias.n78 161.3
R1194 commonsourceibias.n80 commonsourceibias.n18 161.3
R1195 commonsourceibias.n82 commonsourceibias.n81 161.3
R1196 commonsourceibias.n84 commonsourceibias.n16 161.3
R1197 commonsourceibias.n86 commonsourceibias.n85 161.3
R1198 commonsourceibias.n87 commonsourceibias.n15 161.3
R1199 commonsourceibias.n89 commonsourceibias.n88 161.3
R1200 commonsourceibias.n90 commonsourceibias.n14 161.3
R1201 commonsourceibias.n93 commonsourceibias.n92 161.3
R1202 commonsourceibias.n94 commonsourceibias.n13 161.3
R1203 commonsourceibias.n96 commonsourceibias.n95 161.3
R1204 commonsourceibias.n98 commonsourceibias.n12 161.3
R1205 commonsourceibias.n129 commonsourceibias.n126 161.3
R1206 commonsourceibias.n131 commonsourceibias.n130 161.3
R1207 commonsourceibias.n132 commonsourceibias.n125 161.3
R1208 commonsourceibias.n135 commonsourceibias.n134 161.3
R1209 commonsourceibias.n136 commonsourceibias.n124 161.3
R1210 commonsourceibias.n138 commonsourceibias.n137 161.3
R1211 commonsourceibias.n140 commonsourceibias.n123 161.3
R1212 commonsourceibias.n142 commonsourceibias.n141 161.3
R1213 commonsourceibias.n144 commonsourceibias.n143 161.3
R1214 commonsourceibias.n145 commonsourceibias.n121 161.3
R1215 commonsourceibias.n147 commonsourceibias.n146 161.3
R1216 commonsourceibias.n149 commonsourceibias.n148 161.3
R1217 commonsourceibias.n150 commonsourceibias.n119 161.3
R1218 commonsourceibias.n152 commonsourceibias.n151 161.3
R1219 commonsourceibias.n154 commonsourceibias.n153 161.3
R1220 commonsourceibias.n155 commonsourceibias.n117 161.3
R1221 commonsourceibias.n158 commonsourceibias.n157 161.3
R1222 commonsourceibias.n159 commonsourceibias.n11 161.3
R1223 commonsourceibias.n161 commonsourceibias.n160 161.3
R1224 commonsourceibias.n163 commonsourceibias.n9 161.3
R1225 commonsourceibias.n165 commonsourceibias.n164 161.3
R1226 commonsourceibias.n166 commonsourceibias.n8 161.3
R1227 commonsourceibias.n168 commonsourceibias.n167 161.3
R1228 commonsourceibias.n169 commonsourceibias.n7 161.3
R1229 commonsourceibias.n172 commonsourceibias.n171 161.3
R1230 commonsourceibias.n173 commonsourceibias.n6 161.3
R1231 commonsourceibias.n175 commonsourceibias.n174 161.3
R1232 commonsourceibias.n177 commonsourceibias.n4 161.3
R1233 commonsourceibias.n179 commonsourceibias.n178 161.3
R1234 commonsourceibias.n180 commonsourceibias.n3 161.3
R1235 commonsourceibias.n182 commonsourceibias.n181 161.3
R1236 commonsourceibias.n183 commonsourceibias.n2 161.3
R1237 commonsourceibias.n186 commonsourceibias.n185 161.3
R1238 commonsourceibias.n187 commonsourceibias.n1 161.3
R1239 commonsourceibias.n189 commonsourceibias.n188 161.3
R1240 commonsourceibias.n191 commonsourceibias.n0 161.3
R1241 commonsourceibias.n280 commonsourceibias.n194 161.3
R1242 commonsourceibias.n278 commonsourceibias.n277 161.3
R1243 commonsourceibias.n276 commonsourceibias.n195 161.3
R1244 commonsourceibias.n275 commonsourceibias.n274 161.3
R1245 commonsourceibias.n272 commonsourceibias.n196 161.3
R1246 commonsourceibias.n271 commonsourceibias.n270 161.3
R1247 commonsourceibias.n269 commonsourceibias.n197 161.3
R1248 commonsourceibias.n268 commonsourceibias.n267 161.3
R1249 commonsourceibias.n266 commonsourceibias.n198 161.3
R1250 commonsourceibias.n264 commonsourceibias.n263 161.3
R1251 commonsourceibias.n262 commonsourceibias.n200 161.3
R1252 commonsourceibias.n261 commonsourceibias.n260 161.3
R1253 commonsourceibias.n258 commonsourceibias.n201 161.3
R1254 commonsourceibias.n257 commonsourceibias.n256 161.3
R1255 commonsourceibias.n255 commonsourceibias.n202 161.3
R1256 commonsourceibias.n254 commonsourceibias.n253 161.3
R1257 commonsourceibias.n252 commonsourceibias.n203 161.3
R1258 commonsourceibias.n250 commonsourceibias.n249 161.3
R1259 commonsourceibias.n248 commonsourceibias.n205 161.3
R1260 commonsourceibias.n247 commonsourceibias.n246 161.3
R1261 commonsourceibias.n244 commonsourceibias.n206 161.3
R1262 commonsourceibias.n243 commonsourceibias.n242 161.3
R1263 commonsourceibias.n241 commonsourceibias.n240 161.3
R1264 commonsourceibias.n239 commonsourceibias.n208 161.3
R1265 commonsourceibias.n238 commonsourceibias.n237 161.3
R1266 commonsourceibias.n236 commonsourceibias.n235 161.3
R1267 commonsourceibias.n234 commonsourceibias.n210 161.3
R1268 commonsourceibias.n233 commonsourceibias.n232 161.3
R1269 commonsourceibias.n231 commonsourceibias.n230 161.3
R1270 commonsourceibias.n229 commonsourceibias.n212 161.3
R1271 commonsourceibias.n227 commonsourceibias.n226 161.3
R1272 commonsourceibias.n225 commonsourceibias.n213 161.3
R1273 commonsourceibias.n224 commonsourceibias.n223 161.3
R1274 commonsourceibias.n221 commonsourceibias.n214 161.3
R1275 commonsourceibias.n220 commonsourceibias.n219 161.3
R1276 commonsourceibias.n218 commonsourceibias.n215 161.3
R1277 commonsourceibias.n429 commonsourceibias.n343 161.3
R1278 commonsourceibias.n427 commonsourceibias.n426 161.3
R1279 commonsourceibias.n425 commonsourceibias.n344 161.3
R1280 commonsourceibias.n424 commonsourceibias.n423 161.3
R1281 commonsourceibias.n421 commonsourceibias.n345 161.3
R1282 commonsourceibias.n420 commonsourceibias.n419 161.3
R1283 commonsourceibias.n418 commonsourceibias.n346 161.3
R1284 commonsourceibias.n417 commonsourceibias.n416 161.3
R1285 commonsourceibias.n414 commonsourceibias.n347 161.3
R1286 commonsourceibias.n412 commonsourceibias.n411 161.3
R1287 commonsourceibias.n410 commonsourceibias.n348 161.3
R1288 commonsourceibias.n409 commonsourceibias.n408 161.3
R1289 commonsourceibias.n406 commonsourceibias.n349 161.3
R1290 commonsourceibias.n405 commonsourceibias.n404 161.3
R1291 commonsourceibias.n403 commonsourceibias.n350 161.3
R1292 commonsourceibias.n402 commonsourceibias.n401 161.3
R1293 commonsourceibias.n399 commonsourceibias.n351 161.3
R1294 commonsourceibias.n397 commonsourceibias.n396 161.3
R1295 commonsourceibias.n395 commonsourceibias.n352 161.3
R1296 commonsourceibias.n394 commonsourceibias.n393 161.3
R1297 commonsourceibias.n391 commonsourceibias.n353 161.3
R1298 commonsourceibias.n390 commonsourceibias.n389 161.3
R1299 commonsourceibias.n388 commonsourceibias.n387 161.3
R1300 commonsourceibias.n386 commonsourceibias.n355 161.3
R1301 commonsourceibias.n385 commonsourceibias.n384 161.3
R1302 commonsourceibias.n383 commonsourceibias.n382 161.3
R1303 commonsourceibias.n381 commonsourceibias.n357 161.3
R1304 commonsourceibias.n380 commonsourceibias.n379 161.3
R1305 commonsourceibias.n378 commonsourceibias.n377 161.3
R1306 commonsourceibias.n376 commonsourceibias.n359 161.3
R1307 commonsourceibias.n374 commonsourceibias.n373 161.3
R1308 commonsourceibias.n372 commonsourceibias.n360 161.3
R1309 commonsourceibias.n371 commonsourceibias.n370 161.3
R1310 commonsourceibias.n368 commonsourceibias.n361 161.3
R1311 commonsourceibias.n367 commonsourceibias.n366 161.3
R1312 commonsourceibias.n365 commonsourceibias.n362 161.3
R1313 commonsourceibias.n335 commonsourceibias.n334 161.3
R1314 commonsourceibias.n332 commonsourceibias.n294 161.3
R1315 commonsourceibias.n331 commonsourceibias.n330 161.3
R1316 commonsourceibias.n329 commonsourceibias.n328 161.3
R1317 commonsourceibias.n327 commonsourceibias.n296 161.3
R1318 commonsourceibias.n326 commonsourceibias.n325 161.3
R1319 commonsourceibias.n324 commonsourceibias.n323 161.3
R1320 commonsourceibias.n322 commonsourceibias.n298 161.3
R1321 commonsourceibias.n321 commonsourceibias.n320 161.3
R1322 commonsourceibias.n319 commonsourceibias.n318 161.3
R1323 commonsourceibias.n317 commonsourceibias.n300 161.3
R1324 commonsourceibias.n315 commonsourceibias.n314 161.3
R1325 commonsourceibias.n313 commonsourceibias.n301 161.3
R1326 commonsourceibias.n312 commonsourceibias.n311 161.3
R1327 commonsourceibias.n309 commonsourceibias.n302 161.3
R1328 commonsourceibias.n308 commonsourceibias.n307 161.3
R1329 commonsourceibias.n306 commonsourceibias.n303 161.3
R1330 commonsourceibias.n441 commonsourceibias.n293 161.3
R1331 commonsourceibias.n475 commonsourceibias.n284 161.3
R1332 commonsourceibias.n473 commonsourceibias.n472 161.3
R1333 commonsourceibias.n471 commonsourceibias.n285 161.3
R1334 commonsourceibias.n470 commonsourceibias.n469 161.3
R1335 commonsourceibias.n467 commonsourceibias.n286 161.3
R1336 commonsourceibias.n466 commonsourceibias.n465 161.3
R1337 commonsourceibias.n464 commonsourceibias.n287 161.3
R1338 commonsourceibias.n463 commonsourceibias.n462 161.3
R1339 commonsourceibias.n460 commonsourceibias.n288 161.3
R1340 commonsourceibias.n458 commonsourceibias.n457 161.3
R1341 commonsourceibias.n456 commonsourceibias.n289 161.3
R1342 commonsourceibias.n455 commonsourceibias.n454 161.3
R1343 commonsourceibias.n452 commonsourceibias.n290 161.3
R1344 commonsourceibias.n451 commonsourceibias.n450 161.3
R1345 commonsourceibias.n449 commonsourceibias.n291 161.3
R1346 commonsourceibias.n448 commonsourceibias.n447 161.3
R1347 commonsourceibias.n445 commonsourceibias.n292 161.3
R1348 commonsourceibias.n443 commonsourceibias.n442 161.3
R1349 commonsourceibias.n564 commonsourceibias.n478 161.3
R1350 commonsourceibias.n562 commonsourceibias.n561 161.3
R1351 commonsourceibias.n560 commonsourceibias.n479 161.3
R1352 commonsourceibias.n559 commonsourceibias.n558 161.3
R1353 commonsourceibias.n556 commonsourceibias.n480 161.3
R1354 commonsourceibias.n555 commonsourceibias.n554 161.3
R1355 commonsourceibias.n553 commonsourceibias.n481 161.3
R1356 commonsourceibias.n552 commonsourceibias.n551 161.3
R1357 commonsourceibias.n549 commonsourceibias.n482 161.3
R1358 commonsourceibias.n547 commonsourceibias.n546 161.3
R1359 commonsourceibias.n545 commonsourceibias.n483 161.3
R1360 commonsourceibias.n544 commonsourceibias.n543 161.3
R1361 commonsourceibias.n541 commonsourceibias.n484 161.3
R1362 commonsourceibias.n540 commonsourceibias.n539 161.3
R1363 commonsourceibias.n538 commonsourceibias.n485 161.3
R1364 commonsourceibias.n537 commonsourceibias.n536 161.3
R1365 commonsourceibias.n534 commonsourceibias.n486 161.3
R1366 commonsourceibias.n532 commonsourceibias.n531 161.3
R1367 commonsourceibias.n530 commonsourceibias.n487 161.3
R1368 commonsourceibias.n529 commonsourceibias.n528 161.3
R1369 commonsourceibias.n526 commonsourceibias.n488 161.3
R1370 commonsourceibias.n525 commonsourceibias.n524 161.3
R1371 commonsourceibias.n523 commonsourceibias.n522 161.3
R1372 commonsourceibias.n521 commonsourceibias.n490 161.3
R1373 commonsourceibias.n520 commonsourceibias.n519 161.3
R1374 commonsourceibias.n518 commonsourceibias.n517 161.3
R1375 commonsourceibias.n516 commonsourceibias.n492 161.3
R1376 commonsourceibias.n515 commonsourceibias.n514 161.3
R1377 commonsourceibias.n513 commonsourceibias.n512 161.3
R1378 commonsourceibias.n511 commonsourceibias.n494 161.3
R1379 commonsourceibias.n509 commonsourceibias.n508 161.3
R1380 commonsourceibias.n507 commonsourceibias.n495 161.3
R1381 commonsourceibias.n506 commonsourceibias.n505 161.3
R1382 commonsourceibias.n503 commonsourceibias.n496 161.3
R1383 commonsourceibias.n502 commonsourceibias.n501 161.3
R1384 commonsourceibias.n500 commonsourceibias.n497 161.3
R1385 commonsourceibias.n111 commonsourceibias.n109 81.5057
R1386 commonsourceibias.n338 commonsourceibias.n336 81.5057
R1387 commonsourceibias.n111 commonsourceibias.n110 80.9324
R1388 commonsourceibias.n113 commonsourceibias.n112 80.9324
R1389 commonsourceibias.n115 commonsourceibias.n114 80.9324
R1390 commonsourceibias.n108 commonsourceibias.n107 80.9324
R1391 commonsourceibias.n106 commonsourceibias.n105 80.9324
R1392 commonsourceibias.n104 commonsourceibias.n103 80.9324
R1393 commonsourceibias.n102 commonsourceibias.n101 80.9324
R1394 commonsourceibias.n433 commonsourceibias.n432 80.9324
R1395 commonsourceibias.n435 commonsourceibias.n434 80.9324
R1396 commonsourceibias.n437 commonsourceibias.n436 80.9324
R1397 commonsourceibias.n439 commonsourceibias.n438 80.9324
R1398 commonsourceibias.n342 commonsourceibias.n341 80.9324
R1399 commonsourceibias.n340 commonsourceibias.n339 80.9324
R1400 commonsourceibias.n338 commonsourceibias.n337 80.9324
R1401 commonsourceibias.n100 commonsourceibias.n99 80.6037
R1402 commonsourceibias.n193 commonsourceibias.n192 80.6037
R1403 commonsourceibias.n282 commonsourceibias.n281 80.6037
R1404 commonsourceibias.n431 commonsourceibias.n430 80.6037
R1405 commonsourceibias.n477 commonsourceibias.n476 80.6037
R1406 commonsourceibias.n566 commonsourceibias.n565 80.6037
R1407 commonsourceibias.n85 commonsourceibias.n84 56.5617
R1408 commonsourceibias.n71 commonsourceibias.n70 56.5617
R1409 commonsourceibias.n62 commonsourceibias.n61 56.5617
R1410 commonsourceibias.n48 commonsourceibias.n47 56.5617
R1411 commonsourceibias.n178 commonsourceibias.n177 56.5617
R1412 commonsourceibias.n164 commonsourceibias.n163 56.5617
R1413 commonsourceibias.n155 commonsourceibias.n154 56.5617
R1414 commonsourceibias.n141 commonsourceibias.n140 56.5617
R1415 commonsourceibias.n230 commonsourceibias.n229 56.5617
R1416 commonsourceibias.n244 commonsourceibias.n243 56.5617
R1417 commonsourceibias.n253 commonsourceibias.n252 56.5617
R1418 commonsourceibias.n267 commonsourceibias.n266 56.5617
R1419 commonsourceibias.n377 commonsourceibias.n376 56.5617
R1420 commonsourceibias.n391 commonsourceibias.n390 56.5617
R1421 commonsourceibias.n401 commonsourceibias.n399 56.5617
R1422 commonsourceibias.n416 commonsourceibias.n414 56.5617
R1423 commonsourceibias.n462 commonsourceibias.n460 56.5617
R1424 commonsourceibias.n447 commonsourceibias.n445 56.5617
R1425 commonsourceibias.n318 commonsourceibias.n317 56.5617
R1426 commonsourceibias.n332 commonsourceibias.n331 56.5617
R1427 commonsourceibias.n512 commonsourceibias.n511 56.5617
R1428 commonsourceibias.n526 commonsourceibias.n525 56.5617
R1429 commonsourceibias.n536 commonsourceibias.n534 56.5617
R1430 commonsourceibias.n551 commonsourceibias.n549 56.5617
R1431 commonsourceibias.n76 commonsourceibias.n75 56.0773
R1432 commonsourceibias.n57 commonsourceibias.n56 56.0773
R1433 commonsourceibias.n169 commonsourceibias.n168 56.0773
R1434 commonsourceibias.n150 commonsourceibias.n149 56.0773
R1435 commonsourceibias.n239 commonsourceibias.n238 56.0773
R1436 commonsourceibias.n258 commonsourceibias.n257 56.0773
R1437 commonsourceibias.n386 commonsourceibias.n385 56.0773
R1438 commonsourceibias.n406 commonsourceibias.n405 56.0773
R1439 commonsourceibias.n452 commonsourceibias.n451 56.0773
R1440 commonsourceibias.n327 commonsourceibias.n326 56.0773
R1441 commonsourceibias.n521 commonsourceibias.n520 56.0773
R1442 commonsourceibias.n541 commonsourceibias.n540 56.0773
R1443 commonsourceibias.n99 commonsourceibias.n98 55.3321
R1444 commonsourceibias.n192 commonsourceibias.n191 55.3321
R1445 commonsourceibias.n281 commonsourceibias.n280 55.3321
R1446 commonsourceibias.n430 commonsourceibias.n429 55.3321
R1447 commonsourceibias.n476 commonsourceibias.n475 55.3321
R1448 commonsourceibias.n565 commonsourceibias.n564 55.3321
R1449 commonsourceibias.n90 commonsourceibias.n89 55.1086
R1450 commonsourceibias.n41 commonsourceibias.n31 55.1086
R1451 commonsourceibias.n183 commonsourceibias.n182 55.1086
R1452 commonsourceibias.n134 commonsourceibias.n124 55.1086
R1453 commonsourceibias.n223 commonsourceibias.n213 55.1086
R1454 commonsourceibias.n272 commonsourceibias.n271 55.1086
R1455 commonsourceibias.n370 commonsourceibias.n360 55.1086
R1456 commonsourceibias.n421 commonsourceibias.n420 55.1086
R1457 commonsourceibias.n467 commonsourceibias.n466 55.1086
R1458 commonsourceibias.n311 commonsourceibias.n301 55.1086
R1459 commonsourceibias.n505 commonsourceibias.n495 55.1086
R1460 commonsourceibias.n556 commonsourceibias.n555 55.1086
R1461 commonsourceibias.n35 commonsourceibias.n34 47.4592
R1462 commonsourceibias.n128 commonsourceibias.n127 47.4592
R1463 commonsourceibias.n217 commonsourceibias.n216 47.4592
R1464 commonsourceibias.n364 commonsourceibias.n363 47.4592
R1465 commonsourceibias.n305 commonsourceibias.n304 47.4592
R1466 commonsourceibias.n499 commonsourceibias.n498 47.4592
R1467 commonsourceibias.n218 commonsourceibias.n217 44.0436
R1468 commonsourceibias.n365 commonsourceibias.n364 44.0436
R1469 commonsourceibias.n306 commonsourceibias.n305 44.0436
R1470 commonsourceibias.n500 commonsourceibias.n499 44.0436
R1471 commonsourceibias.n36 commonsourceibias.n35 44.0436
R1472 commonsourceibias.n129 commonsourceibias.n128 44.0436
R1473 commonsourceibias.n92 commonsourceibias.n13 42.5146
R1474 commonsourceibias.n39 commonsourceibias.n38 42.5146
R1475 commonsourceibias.n185 commonsourceibias.n1 42.5146
R1476 commonsourceibias.n132 commonsourceibias.n131 42.5146
R1477 commonsourceibias.n221 commonsourceibias.n220 42.5146
R1478 commonsourceibias.n274 commonsourceibias.n195 42.5146
R1479 commonsourceibias.n368 commonsourceibias.n367 42.5146
R1480 commonsourceibias.n423 commonsourceibias.n344 42.5146
R1481 commonsourceibias.n469 commonsourceibias.n285 42.5146
R1482 commonsourceibias.n309 commonsourceibias.n308 42.5146
R1483 commonsourceibias.n503 commonsourceibias.n502 42.5146
R1484 commonsourceibias.n558 commonsourceibias.n479 42.5146
R1485 commonsourceibias.n78 commonsourceibias.n18 41.5458
R1486 commonsourceibias.n53 commonsourceibias.n52 41.5458
R1487 commonsourceibias.n171 commonsourceibias.n6 41.5458
R1488 commonsourceibias.n146 commonsourceibias.n145 41.5458
R1489 commonsourceibias.n235 commonsourceibias.n234 41.5458
R1490 commonsourceibias.n260 commonsourceibias.n200 41.5458
R1491 commonsourceibias.n382 commonsourceibias.n381 41.5458
R1492 commonsourceibias.n408 commonsourceibias.n348 41.5458
R1493 commonsourceibias.n454 commonsourceibias.n289 41.5458
R1494 commonsourceibias.n323 commonsourceibias.n322 41.5458
R1495 commonsourceibias.n517 commonsourceibias.n516 41.5458
R1496 commonsourceibias.n543 commonsourceibias.n483 41.5458
R1497 commonsourceibias.n68 commonsourceibias.n23 40.577
R1498 commonsourceibias.n64 commonsourceibias.n23 40.577
R1499 commonsourceibias.n161 commonsourceibias.n11 40.577
R1500 commonsourceibias.n157 commonsourceibias.n11 40.577
R1501 commonsourceibias.n246 commonsourceibias.n205 40.577
R1502 commonsourceibias.n250 commonsourceibias.n205 40.577
R1503 commonsourceibias.n393 commonsourceibias.n352 40.577
R1504 commonsourceibias.n397 commonsourceibias.n352 40.577
R1505 commonsourceibias.n443 commonsourceibias.n293 40.577
R1506 commonsourceibias.n334 commonsourceibias.n293 40.577
R1507 commonsourceibias.n528 commonsourceibias.n487 40.577
R1508 commonsourceibias.n532 commonsourceibias.n487 40.577
R1509 commonsourceibias.n82 commonsourceibias.n18 39.6083
R1510 commonsourceibias.n52 commonsourceibias.n51 39.6083
R1511 commonsourceibias.n175 commonsourceibias.n6 39.6083
R1512 commonsourceibias.n145 commonsourceibias.n144 39.6083
R1513 commonsourceibias.n234 commonsourceibias.n233 39.6083
R1514 commonsourceibias.n264 commonsourceibias.n200 39.6083
R1515 commonsourceibias.n381 commonsourceibias.n380 39.6083
R1516 commonsourceibias.n412 commonsourceibias.n348 39.6083
R1517 commonsourceibias.n458 commonsourceibias.n289 39.6083
R1518 commonsourceibias.n322 commonsourceibias.n321 39.6083
R1519 commonsourceibias.n516 commonsourceibias.n515 39.6083
R1520 commonsourceibias.n547 commonsourceibias.n483 39.6083
R1521 commonsourceibias.n96 commonsourceibias.n13 38.6395
R1522 commonsourceibias.n38 commonsourceibias.n33 38.6395
R1523 commonsourceibias.n189 commonsourceibias.n1 38.6395
R1524 commonsourceibias.n131 commonsourceibias.n126 38.6395
R1525 commonsourceibias.n220 commonsourceibias.n215 38.6395
R1526 commonsourceibias.n278 commonsourceibias.n195 38.6395
R1527 commonsourceibias.n367 commonsourceibias.n362 38.6395
R1528 commonsourceibias.n427 commonsourceibias.n344 38.6395
R1529 commonsourceibias.n473 commonsourceibias.n285 38.6395
R1530 commonsourceibias.n308 commonsourceibias.n303 38.6395
R1531 commonsourceibias.n502 commonsourceibias.n497 38.6395
R1532 commonsourceibias.n562 commonsourceibias.n479 38.6395
R1533 commonsourceibias.n89 commonsourceibias.n15 26.0455
R1534 commonsourceibias.n45 commonsourceibias.n31 26.0455
R1535 commonsourceibias.n182 commonsourceibias.n3 26.0455
R1536 commonsourceibias.n138 commonsourceibias.n124 26.0455
R1537 commonsourceibias.n227 commonsourceibias.n213 26.0455
R1538 commonsourceibias.n271 commonsourceibias.n197 26.0455
R1539 commonsourceibias.n374 commonsourceibias.n360 26.0455
R1540 commonsourceibias.n420 commonsourceibias.n346 26.0455
R1541 commonsourceibias.n466 commonsourceibias.n287 26.0455
R1542 commonsourceibias.n315 commonsourceibias.n301 26.0455
R1543 commonsourceibias.n509 commonsourceibias.n495 26.0455
R1544 commonsourceibias.n555 commonsourceibias.n481 26.0455
R1545 commonsourceibias.n75 commonsourceibias.n20 25.0767
R1546 commonsourceibias.n58 commonsourceibias.n57 25.0767
R1547 commonsourceibias.n168 commonsourceibias.n8 25.0767
R1548 commonsourceibias.n151 commonsourceibias.n150 25.0767
R1549 commonsourceibias.n240 commonsourceibias.n239 25.0767
R1550 commonsourceibias.n257 commonsourceibias.n202 25.0767
R1551 commonsourceibias.n387 commonsourceibias.n386 25.0767
R1552 commonsourceibias.n405 commonsourceibias.n350 25.0767
R1553 commonsourceibias.n451 commonsourceibias.n291 25.0767
R1554 commonsourceibias.n328 commonsourceibias.n327 25.0767
R1555 commonsourceibias.n522 commonsourceibias.n521 25.0767
R1556 commonsourceibias.n540 commonsourceibias.n485 25.0767
R1557 commonsourceibias.n71 commonsourceibias.n22 24.3464
R1558 commonsourceibias.n61 commonsourceibias.n25 24.3464
R1559 commonsourceibias.n164 commonsourceibias.n10 24.3464
R1560 commonsourceibias.n154 commonsourceibias.n118 24.3464
R1561 commonsourceibias.n243 commonsourceibias.n207 24.3464
R1562 commonsourceibias.n253 commonsourceibias.n204 24.3464
R1563 commonsourceibias.n390 commonsourceibias.n354 24.3464
R1564 commonsourceibias.n401 commonsourceibias.n400 24.3464
R1565 commonsourceibias.n447 commonsourceibias.n446 24.3464
R1566 commonsourceibias.n331 commonsourceibias.n295 24.3464
R1567 commonsourceibias.n525 commonsourceibias.n489 24.3464
R1568 commonsourceibias.n536 commonsourceibias.n535 24.3464
R1569 commonsourceibias.n85 commonsourceibias.n17 23.8546
R1570 commonsourceibias.n47 commonsourceibias.n46 23.8546
R1571 commonsourceibias.n178 commonsourceibias.n5 23.8546
R1572 commonsourceibias.n140 commonsourceibias.n139 23.8546
R1573 commonsourceibias.n229 commonsourceibias.n228 23.8546
R1574 commonsourceibias.n267 commonsourceibias.n199 23.8546
R1575 commonsourceibias.n376 commonsourceibias.n375 23.8546
R1576 commonsourceibias.n416 commonsourceibias.n415 23.8546
R1577 commonsourceibias.n462 commonsourceibias.n461 23.8546
R1578 commonsourceibias.n317 commonsourceibias.n316 23.8546
R1579 commonsourceibias.n511 commonsourceibias.n510 23.8546
R1580 commonsourceibias.n551 commonsourceibias.n550 23.8546
R1581 commonsourceibias.n98 commonsourceibias.n97 17.4607
R1582 commonsourceibias.n191 commonsourceibias.n190 17.4607
R1583 commonsourceibias.n280 commonsourceibias.n279 17.4607
R1584 commonsourceibias.n429 commonsourceibias.n428 17.4607
R1585 commonsourceibias.n475 commonsourceibias.n474 17.4607
R1586 commonsourceibias.n564 commonsourceibias.n563 17.4607
R1587 commonsourceibias.n84 commonsourceibias.n83 16.9689
R1588 commonsourceibias.n48 commonsourceibias.n29 16.9689
R1589 commonsourceibias.n177 commonsourceibias.n176 16.9689
R1590 commonsourceibias.n141 commonsourceibias.n122 16.9689
R1591 commonsourceibias.n230 commonsourceibias.n211 16.9689
R1592 commonsourceibias.n266 commonsourceibias.n265 16.9689
R1593 commonsourceibias.n377 commonsourceibias.n358 16.9689
R1594 commonsourceibias.n414 commonsourceibias.n413 16.9689
R1595 commonsourceibias.n460 commonsourceibias.n459 16.9689
R1596 commonsourceibias.n318 commonsourceibias.n299 16.9689
R1597 commonsourceibias.n512 commonsourceibias.n493 16.9689
R1598 commonsourceibias.n549 commonsourceibias.n548 16.9689
R1599 commonsourceibias.n70 commonsourceibias.n69 16.477
R1600 commonsourceibias.n63 commonsourceibias.n62 16.477
R1601 commonsourceibias.n163 commonsourceibias.n162 16.477
R1602 commonsourceibias.n156 commonsourceibias.n155 16.477
R1603 commonsourceibias.n245 commonsourceibias.n244 16.477
R1604 commonsourceibias.n252 commonsourceibias.n251 16.477
R1605 commonsourceibias.n392 commonsourceibias.n391 16.477
R1606 commonsourceibias.n399 commonsourceibias.n398 16.477
R1607 commonsourceibias.n445 commonsourceibias.n444 16.477
R1608 commonsourceibias.n333 commonsourceibias.n332 16.477
R1609 commonsourceibias.n527 commonsourceibias.n526 16.477
R1610 commonsourceibias.n534 commonsourceibias.n533 16.477
R1611 commonsourceibias.n77 commonsourceibias.n76 15.9852
R1612 commonsourceibias.n56 commonsourceibias.n27 15.9852
R1613 commonsourceibias.n170 commonsourceibias.n169 15.9852
R1614 commonsourceibias.n149 commonsourceibias.n120 15.9852
R1615 commonsourceibias.n238 commonsourceibias.n209 15.9852
R1616 commonsourceibias.n259 commonsourceibias.n258 15.9852
R1617 commonsourceibias.n385 commonsourceibias.n356 15.9852
R1618 commonsourceibias.n407 commonsourceibias.n406 15.9852
R1619 commonsourceibias.n453 commonsourceibias.n452 15.9852
R1620 commonsourceibias.n326 commonsourceibias.n297 15.9852
R1621 commonsourceibias.n520 commonsourceibias.n491 15.9852
R1622 commonsourceibias.n542 commonsourceibias.n541 15.9852
R1623 commonsourceibias.n91 commonsourceibias.n90 15.4934
R1624 commonsourceibias.n41 commonsourceibias.n40 15.4934
R1625 commonsourceibias.n184 commonsourceibias.n183 15.4934
R1626 commonsourceibias.n134 commonsourceibias.n133 15.4934
R1627 commonsourceibias.n223 commonsourceibias.n222 15.4934
R1628 commonsourceibias.n273 commonsourceibias.n272 15.4934
R1629 commonsourceibias.n370 commonsourceibias.n369 15.4934
R1630 commonsourceibias.n422 commonsourceibias.n421 15.4934
R1631 commonsourceibias.n468 commonsourceibias.n467 15.4934
R1632 commonsourceibias.n311 commonsourceibias.n310 15.4934
R1633 commonsourceibias.n505 commonsourceibias.n504 15.4934
R1634 commonsourceibias.n557 commonsourceibias.n556 15.4934
R1635 commonsourceibias.n102 commonsourceibias.n100 13.2663
R1636 commonsourceibias.n433 commonsourceibias.n431 13.2663
R1637 commonsourceibias.n568 commonsourceibias.n283 11.9876
R1638 commonsourceibias.n568 commonsourceibias.n567 10.3347
R1639 commonsourceibias.n159 commonsourceibias.n116 9.50363
R1640 commonsourceibias.n441 commonsourceibias.n440 9.50363
R1641 commonsourceibias.n92 commonsourceibias.n91 9.09948
R1642 commonsourceibias.n40 commonsourceibias.n39 9.09948
R1643 commonsourceibias.n185 commonsourceibias.n184 9.09948
R1644 commonsourceibias.n133 commonsourceibias.n132 9.09948
R1645 commonsourceibias.n222 commonsourceibias.n221 9.09948
R1646 commonsourceibias.n274 commonsourceibias.n273 9.09948
R1647 commonsourceibias.n369 commonsourceibias.n368 9.09948
R1648 commonsourceibias.n423 commonsourceibias.n422 9.09948
R1649 commonsourceibias.n469 commonsourceibias.n468 9.09948
R1650 commonsourceibias.n310 commonsourceibias.n309 9.09948
R1651 commonsourceibias.n504 commonsourceibias.n503 9.09948
R1652 commonsourceibias.n558 commonsourceibias.n557 9.09948
R1653 commonsourceibias.n283 commonsourceibias.n193 8.79261
R1654 commonsourceibias.n567 commonsourceibias.n477 8.79261
R1655 commonsourceibias.n78 commonsourceibias.n77 8.60764
R1656 commonsourceibias.n53 commonsourceibias.n27 8.60764
R1657 commonsourceibias.n171 commonsourceibias.n170 8.60764
R1658 commonsourceibias.n146 commonsourceibias.n120 8.60764
R1659 commonsourceibias.n235 commonsourceibias.n209 8.60764
R1660 commonsourceibias.n260 commonsourceibias.n259 8.60764
R1661 commonsourceibias.n382 commonsourceibias.n356 8.60764
R1662 commonsourceibias.n408 commonsourceibias.n407 8.60764
R1663 commonsourceibias.n454 commonsourceibias.n453 8.60764
R1664 commonsourceibias.n323 commonsourceibias.n297 8.60764
R1665 commonsourceibias.n517 commonsourceibias.n491 8.60764
R1666 commonsourceibias.n543 commonsourceibias.n542 8.60764
R1667 commonsourceibias.n69 commonsourceibias.n68 8.11581
R1668 commonsourceibias.n64 commonsourceibias.n63 8.11581
R1669 commonsourceibias.n162 commonsourceibias.n161 8.11581
R1670 commonsourceibias.n157 commonsourceibias.n156 8.11581
R1671 commonsourceibias.n246 commonsourceibias.n245 8.11581
R1672 commonsourceibias.n251 commonsourceibias.n250 8.11581
R1673 commonsourceibias.n393 commonsourceibias.n392 8.11581
R1674 commonsourceibias.n398 commonsourceibias.n397 8.11581
R1675 commonsourceibias.n444 commonsourceibias.n443 8.11581
R1676 commonsourceibias.n334 commonsourceibias.n333 8.11581
R1677 commonsourceibias.n528 commonsourceibias.n527 8.11581
R1678 commonsourceibias.n533 commonsourceibias.n532 8.11581
R1679 commonsourceibias.n83 commonsourceibias.n82 7.62397
R1680 commonsourceibias.n51 commonsourceibias.n29 7.62397
R1681 commonsourceibias.n176 commonsourceibias.n175 7.62397
R1682 commonsourceibias.n144 commonsourceibias.n122 7.62397
R1683 commonsourceibias.n233 commonsourceibias.n211 7.62397
R1684 commonsourceibias.n265 commonsourceibias.n264 7.62397
R1685 commonsourceibias.n380 commonsourceibias.n358 7.62397
R1686 commonsourceibias.n413 commonsourceibias.n412 7.62397
R1687 commonsourceibias.n459 commonsourceibias.n458 7.62397
R1688 commonsourceibias.n321 commonsourceibias.n299 7.62397
R1689 commonsourceibias.n515 commonsourceibias.n493 7.62397
R1690 commonsourceibias.n548 commonsourceibias.n547 7.62397
R1691 commonsourceibias.n97 commonsourceibias.n96 7.13213
R1692 commonsourceibias.n34 commonsourceibias.n33 7.13213
R1693 commonsourceibias.n190 commonsourceibias.n189 7.13213
R1694 commonsourceibias.n127 commonsourceibias.n126 7.13213
R1695 commonsourceibias.n216 commonsourceibias.n215 7.13213
R1696 commonsourceibias.n279 commonsourceibias.n278 7.13213
R1697 commonsourceibias.n363 commonsourceibias.n362 7.13213
R1698 commonsourceibias.n428 commonsourceibias.n427 7.13213
R1699 commonsourceibias.n474 commonsourceibias.n473 7.13213
R1700 commonsourceibias.n304 commonsourceibias.n303 7.13213
R1701 commonsourceibias.n498 commonsourceibias.n497 7.13213
R1702 commonsourceibias.n563 commonsourceibias.n562 7.13213
R1703 commonsourceibias.n283 commonsourceibias.n282 5.06534
R1704 commonsourceibias.n567 commonsourceibias.n566 5.06534
R1705 commonsourceibias commonsourceibias.n568 4.04308
R1706 commonsourceibias.n109 commonsourceibias.t21 2.82907
R1707 commonsourceibias.n109 commonsourceibias.t35 2.82907
R1708 commonsourceibias.n110 commonsourceibias.t11 2.82907
R1709 commonsourceibias.n110 commonsourceibias.t29 2.82907
R1710 commonsourceibias.n112 commonsourceibias.t57 2.82907
R1711 commonsourceibias.n112 commonsourceibias.t63 2.82907
R1712 commonsourceibias.n114 commonsourceibias.t51 2.82907
R1713 commonsourceibias.n114 commonsourceibias.t43 2.82907
R1714 commonsourceibias.n107 commonsourceibias.t61 2.82907
R1715 commonsourceibias.n107 commonsourceibias.t15 2.82907
R1716 commonsourceibias.n105 commonsourceibias.t25 2.82907
R1717 commonsourceibias.n105 commonsourceibias.t53 2.82907
R1718 commonsourceibias.n103 commonsourceibias.t13 2.82907
R1719 commonsourceibias.n103 commonsourceibias.t47 2.82907
R1720 commonsourceibias.n101 commonsourceibias.t49 2.82907
R1721 commonsourceibias.n101 commonsourceibias.t19 2.82907
R1722 commonsourceibias.n432 commonsourceibias.t27 2.82907
R1723 commonsourceibias.n432 commonsourceibias.t3 2.82907
R1724 commonsourceibias.n434 commonsourceibias.t1 2.82907
R1725 commonsourceibias.n434 commonsourceibias.t55 2.82907
R1726 commonsourceibias.n436 commonsourceibias.t7 2.82907
R1727 commonsourceibias.n436 commonsourceibias.t17 2.82907
R1728 commonsourceibias.n438 commonsourceibias.t59 2.82907
R1729 commonsourceibias.n438 commonsourceibias.t45 2.82907
R1730 commonsourceibias.n341 commonsourceibias.t23 2.82907
R1731 commonsourceibias.n341 commonsourceibias.t5 2.82907
R1732 commonsourceibias.n339 commonsourceibias.t9 2.82907
R1733 commonsourceibias.n339 commonsourceibias.t41 2.82907
R1734 commonsourceibias.n337 commonsourceibias.t39 2.82907
R1735 commonsourceibias.n337 commonsourceibias.t37 2.82907
R1736 commonsourceibias.n336 commonsourceibias.t31 2.82907
R1737 commonsourceibias.n336 commonsourceibias.t33 2.82907
R1738 commonsourceibias.n17 commonsourceibias.n15 0.738255
R1739 commonsourceibias.n46 commonsourceibias.n45 0.738255
R1740 commonsourceibias.n5 commonsourceibias.n3 0.738255
R1741 commonsourceibias.n139 commonsourceibias.n138 0.738255
R1742 commonsourceibias.n228 commonsourceibias.n227 0.738255
R1743 commonsourceibias.n199 commonsourceibias.n197 0.738255
R1744 commonsourceibias.n375 commonsourceibias.n374 0.738255
R1745 commonsourceibias.n415 commonsourceibias.n346 0.738255
R1746 commonsourceibias.n461 commonsourceibias.n287 0.738255
R1747 commonsourceibias.n316 commonsourceibias.n315 0.738255
R1748 commonsourceibias.n510 commonsourceibias.n509 0.738255
R1749 commonsourceibias.n550 commonsourceibias.n481 0.738255
R1750 commonsourceibias.n104 commonsourceibias.n102 0.573776
R1751 commonsourceibias.n106 commonsourceibias.n104 0.573776
R1752 commonsourceibias.n108 commonsourceibias.n106 0.573776
R1753 commonsourceibias.n115 commonsourceibias.n113 0.573776
R1754 commonsourceibias.n113 commonsourceibias.n111 0.573776
R1755 commonsourceibias.n340 commonsourceibias.n338 0.573776
R1756 commonsourceibias.n342 commonsourceibias.n340 0.573776
R1757 commonsourceibias.n439 commonsourceibias.n437 0.573776
R1758 commonsourceibias.n437 commonsourceibias.n435 0.573776
R1759 commonsourceibias.n435 commonsourceibias.n433 0.573776
R1760 commonsourceibias.n116 commonsourceibias.n108 0.287138
R1761 commonsourceibias.n116 commonsourceibias.n115 0.287138
R1762 commonsourceibias.n440 commonsourceibias.n342 0.287138
R1763 commonsourceibias.n440 commonsourceibias.n439 0.287138
R1764 commonsourceibias.n100 commonsourceibias.n12 0.285035
R1765 commonsourceibias.n193 commonsourceibias.n0 0.285035
R1766 commonsourceibias.n282 commonsourceibias.n194 0.285035
R1767 commonsourceibias.n431 commonsourceibias.n343 0.285035
R1768 commonsourceibias.n477 commonsourceibias.n284 0.285035
R1769 commonsourceibias.n566 commonsourceibias.n478 0.285035
R1770 commonsourceibias.n22 commonsourceibias.n20 0.246418
R1771 commonsourceibias.n58 commonsourceibias.n25 0.246418
R1772 commonsourceibias.n10 commonsourceibias.n8 0.246418
R1773 commonsourceibias.n151 commonsourceibias.n118 0.246418
R1774 commonsourceibias.n240 commonsourceibias.n207 0.246418
R1775 commonsourceibias.n204 commonsourceibias.n202 0.246418
R1776 commonsourceibias.n387 commonsourceibias.n354 0.246418
R1777 commonsourceibias.n400 commonsourceibias.n350 0.246418
R1778 commonsourceibias.n446 commonsourceibias.n291 0.246418
R1779 commonsourceibias.n328 commonsourceibias.n295 0.246418
R1780 commonsourceibias.n522 commonsourceibias.n489 0.246418
R1781 commonsourceibias.n535 commonsourceibias.n485 0.246418
R1782 commonsourceibias.n95 commonsourceibias.n12 0.189894
R1783 commonsourceibias.n95 commonsourceibias.n94 0.189894
R1784 commonsourceibias.n94 commonsourceibias.n93 0.189894
R1785 commonsourceibias.n93 commonsourceibias.n14 0.189894
R1786 commonsourceibias.n88 commonsourceibias.n14 0.189894
R1787 commonsourceibias.n88 commonsourceibias.n87 0.189894
R1788 commonsourceibias.n87 commonsourceibias.n86 0.189894
R1789 commonsourceibias.n86 commonsourceibias.n16 0.189894
R1790 commonsourceibias.n81 commonsourceibias.n16 0.189894
R1791 commonsourceibias.n81 commonsourceibias.n80 0.189894
R1792 commonsourceibias.n80 commonsourceibias.n79 0.189894
R1793 commonsourceibias.n79 commonsourceibias.n19 0.189894
R1794 commonsourceibias.n74 commonsourceibias.n19 0.189894
R1795 commonsourceibias.n74 commonsourceibias.n73 0.189894
R1796 commonsourceibias.n73 commonsourceibias.n72 0.189894
R1797 commonsourceibias.n72 commonsourceibias.n21 0.189894
R1798 commonsourceibias.n67 commonsourceibias.n21 0.189894
R1799 commonsourceibias.n67 commonsourceibias.n66 0.189894
R1800 commonsourceibias.n66 commonsourceibias.n65 0.189894
R1801 commonsourceibias.n65 commonsourceibias.n24 0.189894
R1802 commonsourceibias.n60 commonsourceibias.n24 0.189894
R1803 commonsourceibias.n60 commonsourceibias.n59 0.189894
R1804 commonsourceibias.n59 commonsourceibias.n26 0.189894
R1805 commonsourceibias.n55 commonsourceibias.n26 0.189894
R1806 commonsourceibias.n55 commonsourceibias.n54 0.189894
R1807 commonsourceibias.n54 commonsourceibias.n28 0.189894
R1808 commonsourceibias.n50 commonsourceibias.n28 0.189894
R1809 commonsourceibias.n50 commonsourceibias.n49 0.189894
R1810 commonsourceibias.n49 commonsourceibias.n30 0.189894
R1811 commonsourceibias.n44 commonsourceibias.n30 0.189894
R1812 commonsourceibias.n44 commonsourceibias.n43 0.189894
R1813 commonsourceibias.n43 commonsourceibias.n42 0.189894
R1814 commonsourceibias.n42 commonsourceibias.n32 0.189894
R1815 commonsourceibias.n37 commonsourceibias.n32 0.189894
R1816 commonsourceibias.n37 commonsourceibias.n36 0.189894
R1817 commonsourceibias.n158 commonsourceibias.n117 0.189894
R1818 commonsourceibias.n153 commonsourceibias.n117 0.189894
R1819 commonsourceibias.n153 commonsourceibias.n152 0.189894
R1820 commonsourceibias.n152 commonsourceibias.n119 0.189894
R1821 commonsourceibias.n148 commonsourceibias.n119 0.189894
R1822 commonsourceibias.n148 commonsourceibias.n147 0.189894
R1823 commonsourceibias.n147 commonsourceibias.n121 0.189894
R1824 commonsourceibias.n143 commonsourceibias.n121 0.189894
R1825 commonsourceibias.n143 commonsourceibias.n142 0.189894
R1826 commonsourceibias.n142 commonsourceibias.n123 0.189894
R1827 commonsourceibias.n137 commonsourceibias.n123 0.189894
R1828 commonsourceibias.n137 commonsourceibias.n136 0.189894
R1829 commonsourceibias.n136 commonsourceibias.n135 0.189894
R1830 commonsourceibias.n135 commonsourceibias.n125 0.189894
R1831 commonsourceibias.n130 commonsourceibias.n125 0.189894
R1832 commonsourceibias.n130 commonsourceibias.n129 0.189894
R1833 commonsourceibias.n188 commonsourceibias.n0 0.189894
R1834 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1835 commonsourceibias.n187 commonsourceibias.n186 0.189894
R1836 commonsourceibias.n186 commonsourceibias.n2 0.189894
R1837 commonsourceibias.n181 commonsourceibias.n2 0.189894
R1838 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1839 commonsourceibias.n180 commonsourceibias.n179 0.189894
R1840 commonsourceibias.n179 commonsourceibias.n4 0.189894
R1841 commonsourceibias.n174 commonsourceibias.n4 0.189894
R1842 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1843 commonsourceibias.n173 commonsourceibias.n172 0.189894
R1844 commonsourceibias.n172 commonsourceibias.n7 0.189894
R1845 commonsourceibias.n167 commonsourceibias.n7 0.189894
R1846 commonsourceibias.n167 commonsourceibias.n166 0.189894
R1847 commonsourceibias.n166 commonsourceibias.n165 0.189894
R1848 commonsourceibias.n165 commonsourceibias.n9 0.189894
R1849 commonsourceibias.n160 commonsourceibias.n9 0.189894
R1850 commonsourceibias.n277 commonsourceibias.n194 0.189894
R1851 commonsourceibias.n277 commonsourceibias.n276 0.189894
R1852 commonsourceibias.n276 commonsourceibias.n275 0.189894
R1853 commonsourceibias.n275 commonsourceibias.n196 0.189894
R1854 commonsourceibias.n270 commonsourceibias.n196 0.189894
R1855 commonsourceibias.n270 commonsourceibias.n269 0.189894
R1856 commonsourceibias.n269 commonsourceibias.n268 0.189894
R1857 commonsourceibias.n268 commonsourceibias.n198 0.189894
R1858 commonsourceibias.n263 commonsourceibias.n198 0.189894
R1859 commonsourceibias.n263 commonsourceibias.n262 0.189894
R1860 commonsourceibias.n262 commonsourceibias.n261 0.189894
R1861 commonsourceibias.n261 commonsourceibias.n201 0.189894
R1862 commonsourceibias.n256 commonsourceibias.n201 0.189894
R1863 commonsourceibias.n256 commonsourceibias.n255 0.189894
R1864 commonsourceibias.n255 commonsourceibias.n254 0.189894
R1865 commonsourceibias.n254 commonsourceibias.n203 0.189894
R1866 commonsourceibias.n249 commonsourceibias.n203 0.189894
R1867 commonsourceibias.n249 commonsourceibias.n248 0.189894
R1868 commonsourceibias.n248 commonsourceibias.n247 0.189894
R1869 commonsourceibias.n247 commonsourceibias.n206 0.189894
R1870 commonsourceibias.n242 commonsourceibias.n206 0.189894
R1871 commonsourceibias.n242 commonsourceibias.n241 0.189894
R1872 commonsourceibias.n241 commonsourceibias.n208 0.189894
R1873 commonsourceibias.n237 commonsourceibias.n208 0.189894
R1874 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1875 commonsourceibias.n236 commonsourceibias.n210 0.189894
R1876 commonsourceibias.n232 commonsourceibias.n210 0.189894
R1877 commonsourceibias.n232 commonsourceibias.n231 0.189894
R1878 commonsourceibias.n231 commonsourceibias.n212 0.189894
R1879 commonsourceibias.n226 commonsourceibias.n212 0.189894
R1880 commonsourceibias.n226 commonsourceibias.n225 0.189894
R1881 commonsourceibias.n225 commonsourceibias.n224 0.189894
R1882 commonsourceibias.n224 commonsourceibias.n214 0.189894
R1883 commonsourceibias.n219 commonsourceibias.n214 0.189894
R1884 commonsourceibias.n219 commonsourceibias.n218 0.189894
R1885 commonsourceibias.n366 commonsourceibias.n365 0.189894
R1886 commonsourceibias.n366 commonsourceibias.n361 0.189894
R1887 commonsourceibias.n371 commonsourceibias.n361 0.189894
R1888 commonsourceibias.n372 commonsourceibias.n371 0.189894
R1889 commonsourceibias.n373 commonsourceibias.n372 0.189894
R1890 commonsourceibias.n373 commonsourceibias.n359 0.189894
R1891 commonsourceibias.n378 commonsourceibias.n359 0.189894
R1892 commonsourceibias.n379 commonsourceibias.n378 0.189894
R1893 commonsourceibias.n379 commonsourceibias.n357 0.189894
R1894 commonsourceibias.n383 commonsourceibias.n357 0.189894
R1895 commonsourceibias.n384 commonsourceibias.n383 0.189894
R1896 commonsourceibias.n384 commonsourceibias.n355 0.189894
R1897 commonsourceibias.n388 commonsourceibias.n355 0.189894
R1898 commonsourceibias.n389 commonsourceibias.n388 0.189894
R1899 commonsourceibias.n389 commonsourceibias.n353 0.189894
R1900 commonsourceibias.n394 commonsourceibias.n353 0.189894
R1901 commonsourceibias.n395 commonsourceibias.n394 0.189894
R1902 commonsourceibias.n396 commonsourceibias.n395 0.189894
R1903 commonsourceibias.n396 commonsourceibias.n351 0.189894
R1904 commonsourceibias.n402 commonsourceibias.n351 0.189894
R1905 commonsourceibias.n403 commonsourceibias.n402 0.189894
R1906 commonsourceibias.n404 commonsourceibias.n403 0.189894
R1907 commonsourceibias.n404 commonsourceibias.n349 0.189894
R1908 commonsourceibias.n409 commonsourceibias.n349 0.189894
R1909 commonsourceibias.n410 commonsourceibias.n409 0.189894
R1910 commonsourceibias.n411 commonsourceibias.n410 0.189894
R1911 commonsourceibias.n411 commonsourceibias.n347 0.189894
R1912 commonsourceibias.n417 commonsourceibias.n347 0.189894
R1913 commonsourceibias.n418 commonsourceibias.n417 0.189894
R1914 commonsourceibias.n419 commonsourceibias.n418 0.189894
R1915 commonsourceibias.n419 commonsourceibias.n345 0.189894
R1916 commonsourceibias.n424 commonsourceibias.n345 0.189894
R1917 commonsourceibias.n425 commonsourceibias.n424 0.189894
R1918 commonsourceibias.n426 commonsourceibias.n425 0.189894
R1919 commonsourceibias.n426 commonsourceibias.n343 0.189894
R1920 commonsourceibias.n307 commonsourceibias.n306 0.189894
R1921 commonsourceibias.n307 commonsourceibias.n302 0.189894
R1922 commonsourceibias.n312 commonsourceibias.n302 0.189894
R1923 commonsourceibias.n313 commonsourceibias.n312 0.189894
R1924 commonsourceibias.n314 commonsourceibias.n313 0.189894
R1925 commonsourceibias.n314 commonsourceibias.n300 0.189894
R1926 commonsourceibias.n319 commonsourceibias.n300 0.189894
R1927 commonsourceibias.n320 commonsourceibias.n319 0.189894
R1928 commonsourceibias.n320 commonsourceibias.n298 0.189894
R1929 commonsourceibias.n324 commonsourceibias.n298 0.189894
R1930 commonsourceibias.n325 commonsourceibias.n324 0.189894
R1931 commonsourceibias.n325 commonsourceibias.n296 0.189894
R1932 commonsourceibias.n329 commonsourceibias.n296 0.189894
R1933 commonsourceibias.n330 commonsourceibias.n329 0.189894
R1934 commonsourceibias.n330 commonsourceibias.n294 0.189894
R1935 commonsourceibias.n335 commonsourceibias.n294 0.189894
R1936 commonsourceibias.n442 commonsourceibias.n292 0.189894
R1937 commonsourceibias.n448 commonsourceibias.n292 0.189894
R1938 commonsourceibias.n449 commonsourceibias.n448 0.189894
R1939 commonsourceibias.n450 commonsourceibias.n449 0.189894
R1940 commonsourceibias.n450 commonsourceibias.n290 0.189894
R1941 commonsourceibias.n455 commonsourceibias.n290 0.189894
R1942 commonsourceibias.n456 commonsourceibias.n455 0.189894
R1943 commonsourceibias.n457 commonsourceibias.n456 0.189894
R1944 commonsourceibias.n457 commonsourceibias.n288 0.189894
R1945 commonsourceibias.n463 commonsourceibias.n288 0.189894
R1946 commonsourceibias.n464 commonsourceibias.n463 0.189894
R1947 commonsourceibias.n465 commonsourceibias.n464 0.189894
R1948 commonsourceibias.n465 commonsourceibias.n286 0.189894
R1949 commonsourceibias.n470 commonsourceibias.n286 0.189894
R1950 commonsourceibias.n471 commonsourceibias.n470 0.189894
R1951 commonsourceibias.n472 commonsourceibias.n471 0.189894
R1952 commonsourceibias.n472 commonsourceibias.n284 0.189894
R1953 commonsourceibias.n501 commonsourceibias.n500 0.189894
R1954 commonsourceibias.n501 commonsourceibias.n496 0.189894
R1955 commonsourceibias.n506 commonsourceibias.n496 0.189894
R1956 commonsourceibias.n507 commonsourceibias.n506 0.189894
R1957 commonsourceibias.n508 commonsourceibias.n507 0.189894
R1958 commonsourceibias.n508 commonsourceibias.n494 0.189894
R1959 commonsourceibias.n513 commonsourceibias.n494 0.189894
R1960 commonsourceibias.n514 commonsourceibias.n513 0.189894
R1961 commonsourceibias.n514 commonsourceibias.n492 0.189894
R1962 commonsourceibias.n518 commonsourceibias.n492 0.189894
R1963 commonsourceibias.n519 commonsourceibias.n518 0.189894
R1964 commonsourceibias.n519 commonsourceibias.n490 0.189894
R1965 commonsourceibias.n523 commonsourceibias.n490 0.189894
R1966 commonsourceibias.n524 commonsourceibias.n523 0.189894
R1967 commonsourceibias.n524 commonsourceibias.n488 0.189894
R1968 commonsourceibias.n529 commonsourceibias.n488 0.189894
R1969 commonsourceibias.n530 commonsourceibias.n529 0.189894
R1970 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1971 commonsourceibias.n531 commonsourceibias.n486 0.189894
R1972 commonsourceibias.n537 commonsourceibias.n486 0.189894
R1973 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1974 commonsourceibias.n539 commonsourceibias.n538 0.189894
R1975 commonsourceibias.n539 commonsourceibias.n484 0.189894
R1976 commonsourceibias.n544 commonsourceibias.n484 0.189894
R1977 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1978 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1979 commonsourceibias.n546 commonsourceibias.n482 0.189894
R1980 commonsourceibias.n552 commonsourceibias.n482 0.189894
R1981 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1982 commonsourceibias.n554 commonsourceibias.n553 0.189894
R1983 commonsourceibias.n554 commonsourceibias.n480 0.189894
R1984 commonsourceibias.n559 commonsourceibias.n480 0.189894
R1985 commonsourceibias.n560 commonsourceibias.n559 0.189894
R1986 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1987 commonsourceibias.n561 commonsourceibias.n478 0.189894
R1988 commonsourceibias.n159 commonsourceibias.n158 0.170955
R1989 commonsourceibias.n160 commonsourceibias.n159 0.170955
R1990 commonsourceibias.n441 commonsourceibias.n335 0.170955
R1991 commonsourceibias.n442 commonsourceibias.n441 0.170955
R1992 gnd.n6713 gnd.n446 1223.7
R1993 gnd.n6123 gnd.n6076 939.716
R1994 gnd.n7117 gnd.n103 795.207
R1995 gnd.n7281 gnd.n99 795.207
R1996 gnd.n2773 gnd.n2720 795.207
R1997 gnd.n5621 gnd.n2775 795.207
R1998 gnd.n5837 gnd.n2573 795.207
R1999 gnd.n4379 gnd.n2571 795.207
R2000 gnd.n3802 gnd.n2258 795.207
R2001 gnd.n3864 gnd.n3803 795.207
R2002 gnd.n7279 gnd.n105 775.989
R2003 gnd.n173 gnd.n101 775.989
R2004 gnd.n5624 gnd.n5623 775.989
R2005 gnd.n5696 gnd.n2724 775.989
R2006 gnd.n5839 gnd.n2568 775.989
R2007 gnd.n3632 gnd.n2570 775.989
R2008 gnd.n5998 gnd.n5997 775.989
R2009 gnd.n6074 gnd.n2262 775.989
R2010 gnd.n3511 gnd.n2578 771.183
R2011 gnd.n5708 gnd.n2681 771.183
R2012 gnd.n4424 gnd.n3431 771.183
R2013 gnd.n5408 gnd.n2684 771.183
R2014 gnd.n6138 gnd.n873 766.379
R2015 gnd.n2229 gnd.n870 766.379
R2016 gnd.n1745 gnd.n1648 766.379
R2017 gnd.n1741 gnd.n1646 766.379
R2018 gnd.n6122 gnd.n867 756.769
R2019 gnd.n6133 gnd.n6132 756.769
R2020 gnd.n1838 gnd.n1555 756.769
R2021 gnd.n1836 gnd.n1558 756.769
R2022 gnd.n6321 gnd.n678 723.135
R2023 gnd.n6712 gnd.n447 723.135
R2024 gnd.n6924 gnd.n6923 723.135
R2025 gnd.n3688 gnd.n3687 723.135
R2026 gnd.n6321 gnd.n6320 585
R2027 gnd.n6322 gnd.n6321 585
R2028 gnd.n6319 gnd.n680 585
R2029 gnd.n680 gnd.n679 585
R2030 gnd.n6318 gnd.n6317 585
R2031 gnd.n6317 gnd.n6316 585
R2032 gnd.n685 gnd.n684 585
R2033 gnd.n6315 gnd.n685 585
R2034 gnd.n6313 gnd.n6312 585
R2035 gnd.n6314 gnd.n6313 585
R2036 gnd.n6311 gnd.n687 585
R2037 gnd.n687 gnd.n686 585
R2038 gnd.n6310 gnd.n6309 585
R2039 gnd.n6309 gnd.n6308 585
R2040 gnd.n693 gnd.n692 585
R2041 gnd.n6307 gnd.n693 585
R2042 gnd.n6305 gnd.n6304 585
R2043 gnd.n6306 gnd.n6305 585
R2044 gnd.n6303 gnd.n695 585
R2045 gnd.n695 gnd.n694 585
R2046 gnd.n6302 gnd.n6301 585
R2047 gnd.n6301 gnd.n6300 585
R2048 gnd.n701 gnd.n700 585
R2049 gnd.n6299 gnd.n701 585
R2050 gnd.n6297 gnd.n6296 585
R2051 gnd.n6298 gnd.n6297 585
R2052 gnd.n6295 gnd.n703 585
R2053 gnd.n703 gnd.n702 585
R2054 gnd.n6294 gnd.n6293 585
R2055 gnd.n6293 gnd.n6292 585
R2056 gnd.n709 gnd.n708 585
R2057 gnd.n6291 gnd.n709 585
R2058 gnd.n6289 gnd.n6288 585
R2059 gnd.n6290 gnd.n6289 585
R2060 gnd.n6287 gnd.n711 585
R2061 gnd.n711 gnd.n710 585
R2062 gnd.n6286 gnd.n6285 585
R2063 gnd.n6285 gnd.n6284 585
R2064 gnd.n717 gnd.n716 585
R2065 gnd.n6283 gnd.n717 585
R2066 gnd.n6281 gnd.n6280 585
R2067 gnd.n6282 gnd.n6281 585
R2068 gnd.n6279 gnd.n719 585
R2069 gnd.n719 gnd.n718 585
R2070 gnd.n6278 gnd.n6277 585
R2071 gnd.n6277 gnd.n6276 585
R2072 gnd.n725 gnd.n724 585
R2073 gnd.n6275 gnd.n725 585
R2074 gnd.n6273 gnd.n6272 585
R2075 gnd.n6274 gnd.n6273 585
R2076 gnd.n6271 gnd.n727 585
R2077 gnd.n727 gnd.n726 585
R2078 gnd.n6270 gnd.n6269 585
R2079 gnd.n6269 gnd.n6268 585
R2080 gnd.n733 gnd.n732 585
R2081 gnd.n6267 gnd.n733 585
R2082 gnd.n6265 gnd.n6264 585
R2083 gnd.n6266 gnd.n6265 585
R2084 gnd.n6263 gnd.n735 585
R2085 gnd.n735 gnd.n734 585
R2086 gnd.n6262 gnd.n6261 585
R2087 gnd.n6261 gnd.n6260 585
R2088 gnd.n741 gnd.n740 585
R2089 gnd.n6259 gnd.n741 585
R2090 gnd.n6257 gnd.n6256 585
R2091 gnd.n6258 gnd.n6257 585
R2092 gnd.n6255 gnd.n743 585
R2093 gnd.n743 gnd.n742 585
R2094 gnd.n6254 gnd.n6253 585
R2095 gnd.n6253 gnd.n6252 585
R2096 gnd.n749 gnd.n748 585
R2097 gnd.n6251 gnd.n749 585
R2098 gnd.n6249 gnd.n6248 585
R2099 gnd.n6250 gnd.n6249 585
R2100 gnd.n6247 gnd.n751 585
R2101 gnd.n751 gnd.n750 585
R2102 gnd.n6246 gnd.n6245 585
R2103 gnd.n6245 gnd.n6244 585
R2104 gnd.n757 gnd.n756 585
R2105 gnd.n6243 gnd.n757 585
R2106 gnd.n6241 gnd.n6240 585
R2107 gnd.n6242 gnd.n6241 585
R2108 gnd.n6239 gnd.n759 585
R2109 gnd.n759 gnd.n758 585
R2110 gnd.n6238 gnd.n6237 585
R2111 gnd.n6237 gnd.n6236 585
R2112 gnd.n765 gnd.n764 585
R2113 gnd.n6235 gnd.n765 585
R2114 gnd.n6233 gnd.n6232 585
R2115 gnd.n6234 gnd.n6233 585
R2116 gnd.n6231 gnd.n767 585
R2117 gnd.n767 gnd.n766 585
R2118 gnd.n6230 gnd.n6229 585
R2119 gnd.n6229 gnd.n6228 585
R2120 gnd.n773 gnd.n772 585
R2121 gnd.n6227 gnd.n773 585
R2122 gnd.n6225 gnd.n6224 585
R2123 gnd.n6226 gnd.n6225 585
R2124 gnd.n6223 gnd.n775 585
R2125 gnd.n775 gnd.n774 585
R2126 gnd.n6222 gnd.n6221 585
R2127 gnd.n6221 gnd.n6220 585
R2128 gnd.n781 gnd.n780 585
R2129 gnd.n6219 gnd.n781 585
R2130 gnd.n6217 gnd.n6216 585
R2131 gnd.n6218 gnd.n6217 585
R2132 gnd.n6215 gnd.n783 585
R2133 gnd.n783 gnd.n782 585
R2134 gnd.n6214 gnd.n6213 585
R2135 gnd.n6213 gnd.n6212 585
R2136 gnd.n789 gnd.n788 585
R2137 gnd.n6211 gnd.n789 585
R2138 gnd.n6209 gnd.n6208 585
R2139 gnd.n6210 gnd.n6209 585
R2140 gnd.n6207 gnd.n791 585
R2141 gnd.n791 gnd.n790 585
R2142 gnd.n6206 gnd.n6205 585
R2143 gnd.n6205 gnd.n6204 585
R2144 gnd.n797 gnd.n796 585
R2145 gnd.n6203 gnd.n797 585
R2146 gnd.n6201 gnd.n6200 585
R2147 gnd.n6202 gnd.n6201 585
R2148 gnd.n6199 gnd.n799 585
R2149 gnd.n799 gnd.n798 585
R2150 gnd.n6198 gnd.n6197 585
R2151 gnd.n6197 gnd.n6196 585
R2152 gnd.n805 gnd.n804 585
R2153 gnd.n6195 gnd.n805 585
R2154 gnd.n6193 gnd.n6192 585
R2155 gnd.n6194 gnd.n6193 585
R2156 gnd.n6191 gnd.n807 585
R2157 gnd.n807 gnd.n806 585
R2158 gnd.n6190 gnd.n6189 585
R2159 gnd.n6189 gnd.n6188 585
R2160 gnd.n813 gnd.n812 585
R2161 gnd.n6187 gnd.n813 585
R2162 gnd.n6185 gnd.n6184 585
R2163 gnd.n6186 gnd.n6185 585
R2164 gnd.n6183 gnd.n815 585
R2165 gnd.n815 gnd.n814 585
R2166 gnd.n6182 gnd.n6181 585
R2167 gnd.n6181 gnd.n6180 585
R2168 gnd.n821 gnd.n820 585
R2169 gnd.n6179 gnd.n821 585
R2170 gnd.n6177 gnd.n6176 585
R2171 gnd.n6178 gnd.n6177 585
R2172 gnd.n6175 gnd.n823 585
R2173 gnd.n823 gnd.n822 585
R2174 gnd.n6174 gnd.n6173 585
R2175 gnd.n6173 gnd.n6172 585
R2176 gnd.n829 gnd.n828 585
R2177 gnd.n6171 gnd.n829 585
R2178 gnd.n6169 gnd.n6168 585
R2179 gnd.n6170 gnd.n6169 585
R2180 gnd.n6167 gnd.n831 585
R2181 gnd.n831 gnd.n830 585
R2182 gnd.n6166 gnd.n6165 585
R2183 gnd.n6165 gnd.n6164 585
R2184 gnd.n837 gnd.n836 585
R2185 gnd.n6163 gnd.n837 585
R2186 gnd.n6161 gnd.n6160 585
R2187 gnd.n6162 gnd.n6161 585
R2188 gnd.n6159 gnd.n839 585
R2189 gnd.n839 gnd.n838 585
R2190 gnd.n6158 gnd.n6157 585
R2191 gnd.n6157 gnd.n6156 585
R2192 gnd.n845 gnd.n844 585
R2193 gnd.n6155 gnd.n845 585
R2194 gnd.n678 gnd.n677 585
R2195 gnd.n6323 gnd.n678 585
R2196 gnd.n6326 gnd.n6325 585
R2197 gnd.n6325 gnd.n6324 585
R2198 gnd.n675 gnd.n674 585
R2199 gnd.n674 gnd.n673 585
R2200 gnd.n6331 gnd.n6330 585
R2201 gnd.n6332 gnd.n6331 585
R2202 gnd.n672 gnd.n671 585
R2203 gnd.n6333 gnd.n672 585
R2204 gnd.n6336 gnd.n6335 585
R2205 gnd.n6335 gnd.n6334 585
R2206 gnd.n669 gnd.n668 585
R2207 gnd.n668 gnd.n667 585
R2208 gnd.n6341 gnd.n6340 585
R2209 gnd.n6342 gnd.n6341 585
R2210 gnd.n666 gnd.n665 585
R2211 gnd.n6343 gnd.n666 585
R2212 gnd.n6346 gnd.n6345 585
R2213 gnd.n6345 gnd.n6344 585
R2214 gnd.n663 gnd.n662 585
R2215 gnd.n662 gnd.n661 585
R2216 gnd.n6351 gnd.n6350 585
R2217 gnd.n6352 gnd.n6351 585
R2218 gnd.n660 gnd.n659 585
R2219 gnd.n6353 gnd.n660 585
R2220 gnd.n6356 gnd.n6355 585
R2221 gnd.n6355 gnd.n6354 585
R2222 gnd.n657 gnd.n656 585
R2223 gnd.n656 gnd.n655 585
R2224 gnd.n6361 gnd.n6360 585
R2225 gnd.n6362 gnd.n6361 585
R2226 gnd.n654 gnd.n653 585
R2227 gnd.n6363 gnd.n654 585
R2228 gnd.n6366 gnd.n6365 585
R2229 gnd.n6365 gnd.n6364 585
R2230 gnd.n651 gnd.n650 585
R2231 gnd.n650 gnd.n649 585
R2232 gnd.n6371 gnd.n6370 585
R2233 gnd.n6372 gnd.n6371 585
R2234 gnd.n648 gnd.n647 585
R2235 gnd.n6373 gnd.n648 585
R2236 gnd.n6376 gnd.n6375 585
R2237 gnd.n6375 gnd.n6374 585
R2238 gnd.n645 gnd.n644 585
R2239 gnd.n644 gnd.n643 585
R2240 gnd.n6381 gnd.n6380 585
R2241 gnd.n6382 gnd.n6381 585
R2242 gnd.n642 gnd.n641 585
R2243 gnd.n6383 gnd.n642 585
R2244 gnd.n6386 gnd.n6385 585
R2245 gnd.n6385 gnd.n6384 585
R2246 gnd.n639 gnd.n638 585
R2247 gnd.n638 gnd.n637 585
R2248 gnd.n6391 gnd.n6390 585
R2249 gnd.n6392 gnd.n6391 585
R2250 gnd.n636 gnd.n635 585
R2251 gnd.n6393 gnd.n636 585
R2252 gnd.n6396 gnd.n6395 585
R2253 gnd.n6395 gnd.n6394 585
R2254 gnd.n633 gnd.n632 585
R2255 gnd.n632 gnd.n631 585
R2256 gnd.n6401 gnd.n6400 585
R2257 gnd.n6402 gnd.n6401 585
R2258 gnd.n630 gnd.n629 585
R2259 gnd.n6403 gnd.n630 585
R2260 gnd.n6406 gnd.n6405 585
R2261 gnd.n6405 gnd.n6404 585
R2262 gnd.n627 gnd.n626 585
R2263 gnd.n626 gnd.n625 585
R2264 gnd.n6411 gnd.n6410 585
R2265 gnd.n6412 gnd.n6411 585
R2266 gnd.n624 gnd.n623 585
R2267 gnd.n6413 gnd.n624 585
R2268 gnd.n6416 gnd.n6415 585
R2269 gnd.n6415 gnd.n6414 585
R2270 gnd.n621 gnd.n620 585
R2271 gnd.n620 gnd.n619 585
R2272 gnd.n6421 gnd.n6420 585
R2273 gnd.n6422 gnd.n6421 585
R2274 gnd.n618 gnd.n617 585
R2275 gnd.n6423 gnd.n618 585
R2276 gnd.n6426 gnd.n6425 585
R2277 gnd.n6425 gnd.n6424 585
R2278 gnd.n615 gnd.n614 585
R2279 gnd.n614 gnd.n613 585
R2280 gnd.n6431 gnd.n6430 585
R2281 gnd.n6432 gnd.n6431 585
R2282 gnd.n612 gnd.n611 585
R2283 gnd.n6433 gnd.n612 585
R2284 gnd.n6436 gnd.n6435 585
R2285 gnd.n6435 gnd.n6434 585
R2286 gnd.n609 gnd.n608 585
R2287 gnd.n608 gnd.n607 585
R2288 gnd.n6441 gnd.n6440 585
R2289 gnd.n6442 gnd.n6441 585
R2290 gnd.n606 gnd.n605 585
R2291 gnd.n6443 gnd.n606 585
R2292 gnd.n6446 gnd.n6445 585
R2293 gnd.n6445 gnd.n6444 585
R2294 gnd.n603 gnd.n602 585
R2295 gnd.n602 gnd.n601 585
R2296 gnd.n6451 gnd.n6450 585
R2297 gnd.n6452 gnd.n6451 585
R2298 gnd.n600 gnd.n599 585
R2299 gnd.n6453 gnd.n600 585
R2300 gnd.n6456 gnd.n6455 585
R2301 gnd.n6455 gnd.n6454 585
R2302 gnd.n597 gnd.n596 585
R2303 gnd.n596 gnd.n595 585
R2304 gnd.n6461 gnd.n6460 585
R2305 gnd.n6462 gnd.n6461 585
R2306 gnd.n594 gnd.n593 585
R2307 gnd.n6463 gnd.n594 585
R2308 gnd.n6466 gnd.n6465 585
R2309 gnd.n6465 gnd.n6464 585
R2310 gnd.n591 gnd.n590 585
R2311 gnd.n590 gnd.n589 585
R2312 gnd.n6471 gnd.n6470 585
R2313 gnd.n6472 gnd.n6471 585
R2314 gnd.n588 gnd.n587 585
R2315 gnd.n6473 gnd.n588 585
R2316 gnd.n6476 gnd.n6475 585
R2317 gnd.n6475 gnd.n6474 585
R2318 gnd.n585 gnd.n584 585
R2319 gnd.n584 gnd.n583 585
R2320 gnd.n6481 gnd.n6480 585
R2321 gnd.n6482 gnd.n6481 585
R2322 gnd.n582 gnd.n581 585
R2323 gnd.n6483 gnd.n582 585
R2324 gnd.n6486 gnd.n6485 585
R2325 gnd.n6485 gnd.n6484 585
R2326 gnd.n579 gnd.n578 585
R2327 gnd.n578 gnd.n577 585
R2328 gnd.n6491 gnd.n6490 585
R2329 gnd.n6492 gnd.n6491 585
R2330 gnd.n576 gnd.n575 585
R2331 gnd.n6493 gnd.n576 585
R2332 gnd.n6496 gnd.n6495 585
R2333 gnd.n6495 gnd.n6494 585
R2334 gnd.n573 gnd.n572 585
R2335 gnd.n572 gnd.n571 585
R2336 gnd.n6501 gnd.n6500 585
R2337 gnd.n6502 gnd.n6501 585
R2338 gnd.n570 gnd.n569 585
R2339 gnd.n6503 gnd.n570 585
R2340 gnd.n6506 gnd.n6505 585
R2341 gnd.n6505 gnd.n6504 585
R2342 gnd.n567 gnd.n566 585
R2343 gnd.n566 gnd.n565 585
R2344 gnd.n6511 gnd.n6510 585
R2345 gnd.n6512 gnd.n6511 585
R2346 gnd.n564 gnd.n563 585
R2347 gnd.n6513 gnd.n564 585
R2348 gnd.n6516 gnd.n6515 585
R2349 gnd.n6515 gnd.n6514 585
R2350 gnd.n561 gnd.n560 585
R2351 gnd.n560 gnd.n559 585
R2352 gnd.n6521 gnd.n6520 585
R2353 gnd.n6522 gnd.n6521 585
R2354 gnd.n558 gnd.n557 585
R2355 gnd.n6523 gnd.n558 585
R2356 gnd.n6526 gnd.n6525 585
R2357 gnd.n6525 gnd.n6524 585
R2358 gnd.n555 gnd.n554 585
R2359 gnd.n554 gnd.n553 585
R2360 gnd.n6531 gnd.n6530 585
R2361 gnd.n6532 gnd.n6531 585
R2362 gnd.n552 gnd.n551 585
R2363 gnd.n6533 gnd.n552 585
R2364 gnd.n6536 gnd.n6535 585
R2365 gnd.n6535 gnd.n6534 585
R2366 gnd.n549 gnd.n548 585
R2367 gnd.n548 gnd.n547 585
R2368 gnd.n6541 gnd.n6540 585
R2369 gnd.n6542 gnd.n6541 585
R2370 gnd.n546 gnd.n545 585
R2371 gnd.n6543 gnd.n546 585
R2372 gnd.n6546 gnd.n6545 585
R2373 gnd.n6545 gnd.n6544 585
R2374 gnd.n543 gnd.n542 585
R2375 gnd.n542 gnd.n541 585
R2376 gnd.n6551 gnd.n6550 585
R2377 gnd.n6552 gnd.n6551 585
R2378 gnd.n540 gnd.n539 585
R2379 gnd.n6553 gnd.n540 585
R2380 gnd.n6556 gnd.n6555 585
R2381 gnd.n6555 gnd.n6554 585
R2382 gnd.n537 gnd.n536 585
R2383 gnd.n536 gnd.n535 585
R2384 gnd.n6561 gnd.n6560 585
R2385 gnd.n6562 gnd.n6561 585
R2386 gnd.n534 gnd.n533 585
R2387 gnd.n6563 gnd.n534 585
R2388 gnd.n6566 gnd.n6565 585
R2389 gnd.n6565 gnd.n6564 585
R2390 gnd.n531 gnd.n530 585
R2391 gnd.n530 gnd.n529 585
R2392 gnd.n6571 gnd.n6570 585
R2393 gnd.n6572 gnd.n6571 585
R2394 gnd.n528 gnd.n527 585
R2395 gnd.n6573 gnd.n528 585
R2396 gnd.n6576 gnd.n6575 585
R2397 gnd.n6575 gnd.n6574 585
R2398 gnd.n525 gnd.n524 585
R2399 gnd.n524 gnd.n523 585
R2400 gnd.n6581 gnd.n6580 585
R2401 gnd.n6582 gnd.n6581 585
R2402 gnd.n522 gnd.n521 585
R2403 gnd.n6583 gnd.n522 585
R2404 gnd.n6586 gnd.n6585 585
R2405 gnd.n6585 gnd.n6584 585
R2406 gnd.n519 gnd.n518 585
R2407 gnd.n518 gnd.n517 585
R2408 gnd.n6591 gnd.n6590 585
R2409 gnd.n6592 gnd.n6591 585
R2410 gnd.n516 gnd.n515 585
R2411 gnd.n6593 gnd.n516 585
R2412 gnd.n6596 gnd.n6595 585
R2413 gnd.n6595 gnd.n6594 585
R2414 gnd.n513 gnd.n512 585
R2415 gnd.n512 gnd.n511 585
R2416 gnd.n6601 gnd.n6600 585
R2417 gnd.n6602 gnd.n6601 585
R2418 gnd.n510 gnd.n509 585
R2419 gnd.n6603 gnd.n510 585
R2420 gnd.n6606 gnd.n6605 585
R2421 gnd.n6605 gnd.n6604 585
R2422 gnd.n507 gnd.n506 585
R2423 gnd.n506 gnd.n505 585
R2424 gnd.n6611 gnd.n6610 585
R2425 gnd.n6612 gnd.n6611 585
R2426 gnd.n504 gnd.n503 585
R2427 gnd.n6613 gnd.n504 585
R2428 gnd.n6616 gnd.n6615 585
R2429 gnd.n6615 gnd.n6614 585
R2430 gnd.n501 gnd.n500 585
R2431 gnd.n500 gnd.n499 585
R2432 gnd.n6621 gnd.n6620 585
R2433 gnd.n6622 gnd.n6621 585
R2434 gnd.n498 gnd.n497 585
R2435 gnd.n6623 gnd.n498 585
R2436 gnd.n6626 gnd.n6625 585
R2437 gnd.n6625 gnd.n6624 585
R2438 gnd.n495 gnd.n494 585
R2439 gnd.n494 gnd.n493 585
R2440 gnd.n6631 gnd.n6630 585
R2441 gnd.n6632 gnd.n6631 585
R2442 gnd.n492 gnd.n491 585
R2443 gnd.n6633 gnd.n492 585
R2444 gnd.n6636 gnd.n6635 585
R2445 gnd.n6635 gnd.n6634 585
R2446 gnd.n489 gnd.n488 585
R2447 gnd.n488 gnd.n487 585
R2448 gnd.n6641 gnd.n6640 585
R2449 gnd.n6642 gnd.n6641 585
R2450 gnd.n486 gnd.n485 585
R2451 gnd.n6643 gnd.n486 585
R2452 gnd.n6646 gnd.n6645 585
R2453 gnd.n6645 gnd.n6644 585
R2454 gnd.n483 gnd.n482 585
R2455 gnd.n482 gnd.n481 585
R2456 gnd.n6651 gnd.n6650 585
R2457 gnd.n6652 gnd.n6651 585
R2458 gnd.n480 gnd.n479 585
R2459 gnd.n6653 gnd.n480 585
R2460 gnd.n6656 gnd.n6655 585
R2461 gnd.n6655 gnd.n6654 585
R2462 gnd.n477 gnd.n476 585
R2463 gnd.n476 gnd.n475 585
R2464 gnd.n6661 gnd.n6660 585
R2465 gnd.n6662 gnd.n6661 585
R2466 gnd.n474 gnd.n473 585
R2467 gnd.n6663 gnd.n474 585
R2468 gnd.n6666 gnd.n6665 585
R2469 gnd.n6665 gnd.n6664 585
R2470 gnd.n471 gnd.n470 585
R2471 gnd.n470 gnd.n469 585
R2472 gnd.n6671 gnd.n6670 585
R2473 gnd.n6672 gnd.n6671 585
R2474 gnd.n468 gnd.n467 585
R2475 gnd.n6673 gnd.n468 585
R2476 gnd.n6676 gnd.n6675 585
R2477 gnd.n6675 gnd.n6674 585
R2478 gnd.n465 gnd.n464 585
R2479 gnd.n464 gnd.n463 585
R2480 gnd.n6681 gnd.n6680 585
R2481 gnd.n6682 gnd.n6681 585
R2482 gnd.n462 gnd.n461 585
R2483 gnd.n6683 gnd.n462 585
R2484 gnd.n6686 gnd.n6685 585
R2485 gnd.n6685 gnd.n6684 585
R2486 gnd.n459 gnd.n458 585
R2487 gnd.n458 gnd.n457 585
R2488 gnd.n6691 gnd.n6690 585
R2489 gnd.n6692 gnd.n6691 585
R2490 gnd.n456 gnd.n455 585
R2491 gnd.n6693 gnd.n456 585
R2492 gnd.n6696 gnd.n6695 585
R2493 gnd.n6695 gnd.n6694 585
R2494 gnd.n453 gnd.n452 585
R2495 gnd.n452 gnd.n451 585
R2496 gnd.n6702 gnd.n6701 585
R2497 gnd.n6703 gnd.n6702 585
R2498 gnd.n450 gnd.n449 585
R2499 gnd.n6704 gnd.n450 585
R2500 gnd.n6707 gnd.n6706 585
R2501 gnd.n6706 gnd.n6705 585
R2502 gnd.n6708 gnd.n447 585
R2503 gnd.n447 gnd.n446 585
R2504 gnd.n322 gnd.n321 585
R2505 gnd.n6915 gnd.n321 585
R2506 gnd.n6918 gnd.n6917 585
R2507 gnd.n6917 gnd.n6916 585
R2508 gnd.n325 gnd.n324 585
R2509 gnd.n6914 gnd.n325 585
R2510 gnd.n6912 gnd.n6911 585
R2511 gnd.n6913 gnd.n6912 585
R2512 gnd.n328 gnd.n327 585
R2513 gnd.n327 gnd.n326 585
R2514 gnd.n6907 gnd.n6906 585
R2515 gnd.n6906 gnd.n6905 585
R2516 gnd.n331 gnd.n330 585
R2517 gnd.n6904 gnd.n331 585
R2518 gnd.n6902 gnd.n6901 585
R2519 gnd.n6903 gnd.n6902 585
R2520 gnd.n334 gnd.n333 585
R2521 gnd.n333 gnd.n332 585
R2522 gnd.n6897 gnd.n6896 585
R2523 gnd.n6896 gnd.n6895 585
R2524 gnd.n337 gnd.n336 585
R2525 gnd.n6894 gnd.n337 585
R2526 gnd.n6892 gnd.n6891 585
R2527 gnd.n6893 gnd.n6892 585
R2528 gnd.n340 gnd.n339 585
R2529 gnd.n339 gnd.n338 585
R2530 gnd.n6887 gnd.n6886 585
R2531 gnd.n6886 gnd.n6885 585
R2532 gnd.n343 gnd.n342 585
R2533 gnd.n6884 gnd.n343 585
R2534 gnd.n6882 gnd.n6881 585
R2535 gnd.n6883 gnd.n6882 585
R2536 gnd.n346 gnd.n345 585
R2537 gnd.n345 gnd.n344 585
R2538 gnd.n6877 gnd.n6876 585
R2539 gnd.n6876 gnd.n6875 585
R2540 gnd.n349 gnd.n348 585
R2541 gnd.n6874 gnd.n349 585
R2542 gnd.n6872 gnd.n6871 585
R2543 gnd.n6873 gnd.n6872 585
R2544 gnd.n352 gnd.n351 585
R2545 gnd.n351 gnd.n350 585
R2546 gnd.n6867 gnd.n6866 585
R2547 gnd.n6866 gnd.n6865 585
R2548 gnd.n355 gnd.n354 585
R2549 gnd.n6864 gnd.n355 585
R2550 gnd.n6862 gnd.n6861 585
R2551 gnd.n6863 gnd.n6862 585
R2552 gnd.n358 gnd.n357 585
R2553 gnd.n357 gnd.n356 585
R2554 gnd.n6857 gnd.n6856 585
R2555 gnd.n6856 gnd.n6855 585
R2556 gnd.n361 gnd.n360 585
R2557 gnd.n6854 gnd.n361 585
R2558 gnd.n6852 gnd.n6851 585
R2559 gnd.n6853 gnd.n6852 585
R2560 gnd.n364 gnd.n363 585
R2561 gnd.n363 gnd.n362 585
R2562 gnd.n6847 gnd.n6846 585
R2563 gnd.n6846 gnd.n6845 585
R2564 gnd.n367 gnd.n366 585
R2565 gnd.n6844 gnd.n367 585
R2566 gnd.n6842 gnd.n6841 585
R2567 gnd.n6843 gnd.n6842 585
R2568 gnd.n370 gnd.n369 585
R2569 gnd.n369 gnd.n368 585
R2570 gnd.n6837 gnd.n6836 585
R2571 gnd.n6836 gnd.n6835 585
R2572 gnd.n373 gnd.n372 585
R2573 gnd.n6834 gnd.n373 585
R2574 gnd.n6832 gnd.n6831 585
R2575 gnd.n6833 gnd.n6832 585
R2576 gnd.n376 gnd.n375 585
R2577 gnd.n375 gnd.n374 585
R2578 gnd.n6827 gnd.n6826 585
R2579 gnd.n6826 gnd.n6825 585
R2580 gnd.n379 gnd.n378 585
R2581 gnd.n6824 gnd.n379 585
R2582 gnd.n6822 gnd.n6821 585
R2583 gnd.n6823 gnd.n6822 585
R2584 gnd.n382 gnd.n381 585
R2585 gnd.n381 gnd.n380 585
R2586 gnd.n6817 gnd.n6816 585
R2587 gnd.n6816 gnd.n6815 585
R2588 gnd.n385 gnd.n384 585
R2589 gnd.n6814 gnd.n385 585
R2590 gnd.n6812 gnd.n6811 585
R2591 gnd.n6813 gnd.n6812 585
R2592 gnd.n388 gnd.n387 585
R2593 gnd.n387 gnd.n386 585
R2594 gnd.n6807 gnd.n6806 585
R2595 gnd.n6806 gnd.n6805 585
R2596 gnd.n391 gnd.n390 585
R2597 gnd.n6804 gnd.n391 585
R2598 gnd.n6802 gnd.n6801 585
R2599 gnd.n6803 gnd.n6802 585
R2600 gnd.n394 gnd.n393 585
R2601 gnd.n393 gnd.n392 585
R2602 gnd.n6797 gnd.n6796 585
R2603 gnd.n6796 gnd.n6795 585
R2604 gnd.n397 gnd.n396 585
R2605 gnd.n6794 gnd.n397 585
R2606 gnd.n6792 gnd.n6791 585
R2607 gnd.n6793 gnd.n6792 585
R2608 gnd.n400 gnd.n399 585
R2609 gnd.n399 gnd.n398 585
R2610 gnd.n6787 gnd.n6786 585
R2611 gnd.n6786 gnd.n6785 585
R2612 gnd.n403 gnd.n402 585
R2613 gnd.n6784 gnd.n403 585
R2614 gnd.n6782 gnd.n6781 585
R2615 gnd.n6783 gnd.n6782 585
R2616 gnd.n406 gnd.n405 585
R2617 gnd.n405 gnd.n404 585
R2618 gnd.n6777 gnd.n6776 585
R2619 gnd.n6776 gnd.n6775 585
R2620 gnd.n409 gnd.n408 585
R2621 gnd.n6774 gnd.n409 585
R2622 gnd.n6772 gnd.n6771 585
R2623 gnd.n6773 gnd.n6772 585
R2624 gnd.n412 gnd.n411 585
R2625 gnd.n411 gnd.n410 585
R2626 gnd.n6767 gnd.n6766 585
R2627 gnd.n6766 gnd.n6765 585
R2628 gnd.n415 gnd.n414 585
R2629 gnd.n6764 gnd.n415 585
R2630 gnd.n6762 gnd.n6761 585
R2631 gnd.n6763 gnd.n6762 585
R2632 gnd.n418 gnd.n417 585
R2633 gnd.n417 gnd.n416 585
R2634 gnd.n6757 gnd.n6756 585
R2635 gnd.n6756 gnd.n6755 585
R2636 gnd.n421 gnd.n420 585
R2637 gnd.n6754 gnd.n421 585
R2638 gnd.n6752 gnd.n6751 585
R2639 gnd.n6753 gnd.n6752 585
R2640 gnd.n424 gnd.n423 585
R2641 gnd.n423 gnd.n422 585
R2642 gnd.n6747 gnd.n6746 585
R2643 gnd.n6746 gnd.n6745 585
R2644 gnd.n427 gnd.n426 585
R2645 gnd.n6744 gnd.n427 585
R2646 gnd.n6742 gnd.n6741 585
R2647 gnd.n6743 gnd.n6742 585
R2648 gnd.n430 gnd.n429 585
R2649 gnd.n429 gnd.n428 585
R2650 gnd.n6737 gnd.n6736 585
R2651 gnd.n6736 gnd.n6735 585
R2652 gnd.n433 gnd.n432 585
R2653 gnd.n6734 gnd.n433 585
R2654 gnd.n6732 gnd.n6731 585
R2655 gnd.n6733 gnd.n6732 585
R2656 gnd.n436 gnd.n435 585
R2657 gnd.n435 gnd.n434 585
R2658 gnd.n6727 gnd.n6726 585
R2659 gnd.n6726 gnd.n6725 585
R2660 gnd.n439 gnd.n438 585
R2661 gnd.n6724 gnd.n439 585
R2662 gnd.n6722 gnd.n6721 585
R2663 gnd.n6723 gnd.n6722 585
R2664 gnd.n442 gnd.n441 585
R2665 gnd.n441 gnd.n440 585
R2666 gnd.n6717 gnd.n6716 585
R2667 gnd.n6716 gnd.n6715 585
R2668 gnd.n445 gnd.n444 585
R2669 gnd.n6714 gnd.n445 585
R2670 gnd.n6712 gnd.n6711 585
R2671 gnd.n6713 gnd.n6712 585
R2672 gnd.n5837 gnd.n5836 585
R2673 gnd.n5838 gnd.n5837 585
R2674 gnd.n2559 gnd.n2558 585
R2675 gnd.n4092 gnd.n2559 585
R2676 gnd.n5846 gnd.n5845 585
R2677 gnd.n5845 gnd.n5844 585
R2678 gnd.n5847 gnd.n2553 585
R2679 gnd.n4084 gnd.n2553 585
R2680 gnd.n5849 gnd.n5848 585
R2681 gnd.n5850 gnd.n5849 585
R2682 gnd.n2537 gnd.n2536 585
R2683 gnd.n4075 gnd.n2537 585
R2684 gnd.n5858 gnd.n5857 585
R2685 gnd.n5857 gnd.n5856 585
R2686 gnd.n5859 gnd.n2531 585
R2687 gnd.n4067 gnd.n2531 585
R2688 gnd.n5861 gnd.n5860 585
R2689 gnd.n5862 gnd.n5861 585
R2690 gnd.n2515 gnd.n2514 585
R2691 gnd.n4059 gnd.n2515 585
R2692 gnd.n5870 gnd.n5869 585
R2693 gnd.n5869 gnd.n5868 585
R2694 gnd.n5871 gnd.n2509 585
R2695 gnd.n4051 gnd.n2509 585
R2696 gnd.n5873 gnd.n5872 585
R2697 gnd.n5874 gnd.n5873 585
R2698 gnd.n2494 gnd.n2493 585
R2699 gnd.n4043 gnd.n2494 585
R2700 gnd.n5882 gnd.n5881 585
R2701 gnd.n5881 gnd.n5880 585
R2702 gnd.n5883 gnd.n2488 585
R2703 gnd.n4035 gnd.n2488 585
R2704 gnd.n5885 gnd.n5884 585
R2705 gnd.n5886 gnd.n5885 585
R2706 gnd.n2472 gnd.n2471 585
R2707 gnd.n4027 gnd.n2472 585
R2708 gnd.n5894 gnd.n5893 585
R2709 gnd.n5893 gnd.n5892 585
R2710 gnd.n5895 gnd.n2466 585
R2711 gnd.n4019 gnd.n2466 585
R2712 gnd.n5897 gnd.n5896 585
R2713 gnd.n5898 gnd.n5897 585
R2714 gnd.n2452 gnd.n2451 585
R2715 gnd.n4011 gnd.n2452 585
R2716 gnd.n5906 gnd.n5905 585
R2717 gnd.n5905 gnd.n5904 585
R2718 gnd.n5907 gnd.n2446 585
R2719 gnd.n4003 gnd.n2446 585
R2720 gnd.n5909 gnd.n5908 585
R2721 gnd.n5910 gnd.n5909 585
R2722 gnd.n2433 gnd.n2432 585
R2723 gnd.n3995 gnd.n2433 585
R2724 gnd.n5919 gnd.n5918 585
R2725 gnd.n5918 gnd.n5917 585
R2726 gnd.n5920 gnd.n2427 585
R2727 gnd.n3986 gnd.n2427 585
R2728 gnd.n5922 gnd.n5921 585
R2729 gnd.n5923 gnd.n5922 585
R2730 gnd.n2415 gnd.n2414 585
R2731 gnd.n3976 gnd.n2415 585
R2732 gnd.n5931 gnd.n5930 585
R2733 gnd.n5930 gnd.n5929 585
R2734 gnd.n5932 gnd.n2409 585
R2735 gnd.n3968 gnd.n2409 585
R2736 gnd.n5934 gnd.n5933 585
R2737 gnd.n5935 gnd.n5934 585
R2738 gnd.n2394 gnd.n2393 585
R2739 gnd.n2405 gnd.n2394 585
R2740 gnd.n5943 gnd.n5942 585
R2741 gnd.n5942 gnd.n5941 585
R2742 gnd.n5944 gnd.n2388 585
R2743 gnd.n2395 gnd.n2388 585
R2744 gnd.n5946 gnd.n5945 585
R2745 gnd.n5947 gnd.n5946 585
R2746 gnd.n2375 gnd.n2374 585
R2747 gnd.n2378 gnd.n2375 585
R2748 gnd.n5955 gnd.n5954 585
R2749 gnd.n5954 gnd.n5953 585
R2750 gnd.n5956 gnd.n2369 585
R2751 gnd.n2369 gnd.n2368 585
R2752 gnd.n5958 gnd.n5957 585
R2753 gnd.n5959 gnd.n5958 585
R2754 gnd.n2354 gnd.n2353 585
R2755 gnd.n2365 gnd.n2354 585
R2756 gnd.n5967 gnd.n5966 585
R2757 gnd.n5966 gnd.n5965 585
R2758 gnd.n5968 gnd.n2348 585
R2759 gnd.n2355 gnd.n2348 585
R2760 gnd.n5970 gnd.n5969 585
R2761 gnd.n5971 gnd.n5970 585
R2762 gnd.n2335 gnd.n2334 585
R2763 gnd.n2338 gnd.n2335 585
R2764 gnd.n5979 gnd.n5978 585
R2765 gnd.n5978 gnd.n5977 585
R2766 gnd.n5980 gnd.n2329 585
R2767 gnd.n2329 gnd.n2327 585
R2768 gnd.n5982 gnd.n5981 585
R2769 gnd.n5983 gnd.n5982 585
R2770 gnd.n2330 gnd.n2328 585
R2771 gnd.n2328 gnd.n2315 585
R2772 gnd.n3869 gnd.n2316 585
R2773 gnd.n5989 gnd.n2316 585
R2774 gnd.n3806 gnd.n3804 585
R2775 gnd.n3804 gnd.n2313 585
R2776 gnd.n3874 gnd.n3873 585
R2777 gnd.n3881 gnd.n3874 585
R2778 gnd.n3805 gnd.n3803 585
R2779 gnd.n3803 gnd.n2259 585
R2780 gnd.n3865 gnd.n3864 585
R2781 gnd.n3863 gnd.n3862 585
R2782 gnd.n3861 gnd.n3860 585
R2783 gnd.n3859 gnd.n3858 585
R2784 gnd.n3857 gnd.n3856 585
R2785 gnd.n3855 gnd.n3854 585
R2786 gnd.n3853 gnd.n3852 585
R2787 gnd.n3851 gnd.n3850 585
R2788 gnd.n3849 gnd.n3848 585
R2789 gnd.n3847 gnd.n3846 585
R2790 gnd.n3845 gnd.n3844 585
R2791 gnd.n3843 gnd.n3842 585
R2792 gnd.n3841 gnd.n3840 585
R2793 gnd.n3839 gnd.n3838 585
R2794 gnd.n3837 gnd.n3836 585
R2795 gnd.n3835 gnd.n3834 585
R2796 gnd.n3833 gnd.n3832 585
R2797 gnd.n3825 gnd.n3822 585
R2798 gnd.n3828 gnd.n2258 585
R2799 gnd.n6076 gnd.n2258 585
R2800 gnd.n4380 gnd.n4379 585
R2801 gnd.n4381 gnd.n3471 585
R2802 gnd.n3570 gnd.n3468 585
R2803 gnd.n3569 gnd.n3568 585
R2804 gnd.n3481 gnd.n3480 585
R2805 gnd.n3557 gnd.n3556 585
R2806 gnd.n3555 gnd.n3554 585
R2807 gnd.n3543 gnd.n3488 585
R2808 gnd.n3545 gnd.n3544 585
R2809 gnd.n3542 gnd.n3494 585
R2810 gnd.n3493 gnd.n3492 585
R2811 gnd.n3533 gnd.n3532 585
R2812 gnd.n3531 gnd.n3530 585
R2813 gnd.n3519 gnd.n3500 585
R2814 gnd.n3521 gnd.n3520 585
R2815 gnd.n3518 gnd.n3508 585
R2816 gnd.n3507 gnd.n3506 585
R2817 gnd.n3505 gnd.n3504 585
R2818 gnd.n2575 gnd.n2573 585
R2819 gnd.n4377 gnd.n2573 585
R2820 gnd.n3640 gnd.n2571 585
R2821 gnd.n5838 gnd.n2571 585
R2822 gnd.n4091 gnd.n4090 585
R2823 gnd.n4092 gnd.n4091 585
R2824 gnd.n3639 gnd.n2562 585
R2825 gnd.n5844 gnd.n2562 585
R2826 gnd.n4086 gnd.n4085 585
R2827 gnd.n4085 gnd.n4084 585
R2828 gnd.n3642 gnd.n2551 585
R2829 gnd.n5850 gnd.n2551 585
R2830 gnd.n4074 gnd.n4073 585
R2831 gnd.n4075 gnd.n4074 585
R2832 gnd.n3646 gnd.n2540 585
R2833 gnd.n5856 gnd.n2540 585
R2834 gnd.n4069 gnd.n4068 585
R2835 gnd.n4068 gnd.n4067 585
R2836 gnd.n3648 gnd.n2529 585
R2837 gnd.n5862 gnd.n2529 585
R2838 gnd.n4058 gnd.n4057 585
R2839 gnd.n4059 gnd.n4058 585
R2840 gnd.n3652 gnd.n2518 585
R2841 gnd.n5868 gnd.n2518 585
R2842 gnd.n4053 gnd.n4052 585
R2843 gnd.n4052 gnd.n4051 585
R2844 gnd.n3654 gnd.n2508 585
R2845 gnd.n5874 gnd.n2508 585
R2846 gnd.n4042 gnd.n4041 585
R2847 gnd.n4043 gnd.n4042 585
R2848 gnd.n3659 gnd.n2497 585
R2849 gnd.n5880 gnd.n2497 585
R2850 gnd.n4037 gnd.n4036 585
R2851 gnd.n4036 gnd.n4035 585
R2852 gnd.n3661 gnd.n2486 585
R2853 gnd.n5886 gnd.n2486 585
R2854 gnd.n4026 gnd.n4025 585
R2855 gnd.n4027 gnd.n4026 585
R2856 gnd.n3665 gnd.n2475 585
R2857 gnd.n5892 gnd.n2475 585
R2858 gnd.n4021 gnd.n4020 585
R2859 gnd.n4020 gnd.n4019 585
R2860 gnd.n3667 gnd.n2465 585
R2861 gnd.n5898 gnd.n2465 585
R2862 gnd.n4010 gnd.n4009 585
R2863 gnd.n4011 gnd.n4010 585
R2864 gnd.n3672 gnd.n2455 585
R2865 gnd.n5904 gnd.n2455 585
R2866 gnd.n4005 gnd.n4004 585
R2867 gnd.n4004 gnd.n4003 585
R2868 gnd.n3674 gnd.n2444 585
R2869 gnd.n5910 gnd.n2444 585
R2870 gnd.n3994 gnd.n3993 585
R2871 gnd.n3995 gnd.n3994 585
R2872 gnd.n3678 gnd.n2436 585
R2873 gnd.n5917 gnd.n2436 585
R2874 gnd.n3988 gnd.n3987 585
R2875 gnd.n3987 gnd.n3986 585
R2876 gnd.n3680 gnd.n2426 585
R2877 gnd.n5923 gnd.n2426 585
R2878 gnd.n3975 gnd.n3974 585
R2879 gnd.n3976 gnd.n3975 585
R2880 gnd.n3789 gnd.n2417 585
R2881 gnd.n5929 gnd.n2417 585
R2882 gnd.n3970 gnd.n3969 585
R2883 gnd.n3969 gnd.n3968 585
R2884 gnd.n3922 gnd.n2407 585
R2885 gnd.n5935 gnd.n2407 585
R2886 gnd.n3921 gnd.n3920 585
R2887 gnd.n3920 gnd.n2405 585
R2888 gnd.n3791 gnd.n2397 585
R2889 gnd.n5941 gnd.n2397 585
R2890 gnd.n3916 gnd.n3915 585
R2891 gnd.n3915 gnd.n2395 585
R2892 gnd.n3914 gnd.n2387 585
R2893 gnd.n5947 gnd.n2387 585
R2894 gnd.n3913 gnd.n3912 585
R2895 gnd.n3912 gnd.n2378 585
R2896 gnd.n3793 gnd.n2377 585
R2897 gnd.n5953 gnd.n2377 585
R2898 gnd.n3908 gnd.n3907 585
R2899 gnd.n3907 gnd.n2368 585
R2900 gnd.n3906 gnd.n2367 585
R2901 gnd.n5959 gnd.n2367 585
R2902 gnd.n3905 gnd.n3904 585
R2903 gnd.n3904 gnd.n2365 585
R2904 gnd.n3795 gnd.n2357 585
R2905 gnd.n5965 gnd.n2357 585
R2906 gnd.n3900 gnd.n3899 585
R2907 gnd.n3899 gnd.n2355 585
R2908 gnd.n3898 gnd.n2347 585
R2909 gnd.n5971 gnd.n2347 585
R2910 gnd.n3897 gnd.n3896 585
R2911 gnd.n3896 gnd.n2338 585
R2912 gnd.n3797 gnd.n2337 585
R2913 gnd.n5977 gnd.n2337 585
R2914 gnd.n3892 gnd.n3891 585
R2915 gnd.n3891 gnd.n2327 585
R2916 gnd.n3890 gnd.n2326 585
R2917 gnd.n5983 gnd.n2326 585
R2918 gnd.n3889 gnd.n3888 585
R2919 gnd.n3888 gnd.n2315 585
R2920 gnd.n3799 gnd.n2314 585
R2921 gnd.n5989 gnd.n2314 585
R2922 gnd.n3884 gnd.n3883 585
R2923 gnd.n3883 gnd.n2313 585
R2924 gnd.n3882 gnd.n3801 585
R2925 gnd.n3882 gnd.n3881 585
R2926 gnd.n3826 gnd.n3802 585
R2927 gnd.n3802 gnd.n2259 585
R2928 gnd.n7184 gnd.n103 585
R2929 gnd.n7280 gnd.n103 585
R2930 gnd.n7185 gnd.n7115 585
R2931 gnd.n7115 gnd.n100 585
R2932 gnd.n7186 gnd.n182 585
R2933 gnd.n7200 gnd.n182 585
R2934 gnd.n194 gnd.n192 585
R2935 gnd.n192 gnd.n181 585
R2936 gnd.n7191 gnd.n7190 585
R2937 gnd.n7192 gnd.n7191 585
R2938 gnd.n193 gnd.n191 585
R2939 gnd.n191 gnd.n188 585
R2940 gnd.n7111 gnd.n7110 585
R2941 gnd.n7110 gnd.n7109 585
R2942 gnd.n197 gnd.n196 585
R2943 gnd.n207 gnd.n197 585
R2944 gnd.n7100 gnd.n7099 585
R2945 gnd.n7101 gnd.n7100 585
R2946 gnd.n209 gnd.n208 585
R2947 gnd.n208 gnd.n204 585
R2948 gnd.n7095 gnd.n7094 585
R2949 gnd.n7094 gnd.n7093 585
R2950 gnd.n212 gnd.n211 585
R2951 gnd.n214 gnd.n212 585
R2952 gnd.n7084 gnd.n7083 585
R2953 gnd.n7085 gnd.n7084 585
R2954 gnd.n224 gnd.n223 585
R2955 gnd.n223 gnd.n221 585
R2956 gnd.n7079 gnd.n7078 585
R2957 gnd.n7078 gnd.n7077 585
R2958 gnd.n227 gnd.n226 585
R2959 gnd.n237 gnd.n227 585
R2960 gnd.n7068 gnd.n7067 585
R2961 gnd.n7069 gnd.n7068 585
R2962 gnd.n239 gnd.n238 585
R2963 gnd.n238 gnd.n234 585
R2964 gnd.n7063 gnd.n7062 585
R2965 gnd.n7062 gnd.n7061 585
R2966 gnd.n242 gnd.n241 585
R2967 gnd.n244 gnd.n242 585
R2968 gnd.n7052 gnd.n7051 585
R2969 gnd.n7053 gnd.n7052 585
R2970 gnd.n254 gnd.n253 585
R2971 gnd.n253 gnd.n251 585
R2972 gnd.n7047 gnd.n7046 585
R2973 gnd.n7046 gnd.n7045 585
R2974 gnd.n257 gnd.n256 585
R2975 gnd.n7011 gnd.n257 585
R2976 gnd.n7024 gnd.n7023 585
R2977 gnd.n7023 gnd.n7022 585
R2978 gnd.n7025 gnd.n288 585
R2979 gnd.n7017 gnd.n288 585
R2980 gnd.n6928 gnd.n285 585
R2981 gnd.n6929 gnd.n6928 585
R2982 gnd.n7030 gnd.n284 585
R2983 gnd.n6952 gnd.n284 585
R2984 gnd.n7031 gnd.n283 585
R2985 gnd.n6947 gnd.n283 585
R2986 gnd.n7032 gnd.n282 585
R2987 gnd.n308 gnd.n282 585
R2988 gnd.n279 gnd.n277 585
R2989 gnd.n6939 gnd.n277 585
R2990 gnd.n7037 gnd.n7036 585
R2991 gnd.n7038 gnd.n7037 585
R2992 gnd.n278 gnd.n276 585
R2993 gnd.n5548 gnd.n276 585
R2994 gnd.n5590 gnd.n5588 585
R2995 gnd.n5588 gnd.n5587 585
R2996 gnd.n5591 gnd.n2801 585
R2997 gnd.n2813 gnd.n2801 585
R2998 gnd.n5592 gnd.n2800 585
R2999 gnd.n5579 gnd.n2800 585
R3000 gnd.n5559 gnd.n2798 585
R3001 gnd.n5560 gnd.n5559 585
R3002 gnd.n5596 gnd.n2797 585
R3003 gnd.n2821 gnd.n2797 585
R3004 gnd.n5597 gnd.n2796 585
R3005 gnd.n5525 gnd.n2796 585
R3006 gnd.n5598 gnd.n2795 585
R3007 gnd.n2847 gnd.n2795 585
R3008 gnd.n5514 gnd.n2793 585
R3009 gnd.n5515 gnd.n5514 585
R3010 gnd.n5602 gnd.n2792 585
R3011 gnd.n5502 gnd.n2792 585
R3012 gnd.n5603 gnd.n2791 585
R3013 gnd.n2855 gnd.n2791 585
R3014 gnd.n5604 gnd.n2790 585
R3015 gnd.n5488 gnd.n2790 585
R3016 gnd.n2875 gnd.n2788 585
R3017 gnd.n2876 gnd.n2875 585
R3018 gnd.n5608 gnd.n2787 585
R3019 gnd.n5478 gnd.n2787 585
R3020 gnd.n5609 gnd.n2786 585
R3021 gnd.n5466 gnd.n2786 585
R3022 gnd.n5610 gnd.n2785 585
R3023 gnd.n2883 gnd.n2785 585
R3024 gnd.n2894 gnd.n2783 585
R3025 gnd.n5457 gnd.n2894 585
R3026 gnd.n5614 gnd.n2782 585
R3027 gnd.n2904 gnd.n2782 585
R3028 gnd.n5615 gnd.n2781 585
R3029 gnd.n5447 gnd.n2781 585
R3030 gnd.n5616 gnd.n2780 585
R3031 gnd.n5435 gnd.n2780 585
R3032 gnd.n2777 gnd.n2776 585
R3033 gnd.n2923 gnd.n2776 585
R3034 gnd.n5621 gnd.n5620 585
R3035 gnd.n5622 gnd.n5621 585
R3036 gnd.n3002 gnd.n2775 585
R3037 gnd.n3006 gnd.n3005 585
R3038 gnd.n3008 gnd.n3007 585
R3039 gnd.n2997 gnd.n2996 585
R3040 gnd.n3020 gnd.n2998 585
R3041 gnd.n3022 gnd.n3021 585
R3042 gnd.n3024 gnd.n3023 585
R3043 gnd.n2988 gnd.n2987 585
R3044 gnd.n3037 gnd.n2989 585
R3045 gnd.n3039 gnd.n3038 585
R3046 gnd.n3041 gnd.n3040 585
R3047 gnd.n2979 gnd.n2978 585
R3048 gnd.n3054 gnd.n2980 585
R3049 gnd.n3056 gnd.n3055 585
R3050 gnd.n3058 gnd.n3057 585
R3051 gnd.n2970 gnd.n2969 585
R3052 gnd.n3071 gnd.n2971 585
R3053 gnd.n3072 gnd.n2966 585
R3054 gnd.n3073 gnd.n2720 585
R3055 gnd.n5698 gnd.n2720 585
R3056 gnd.n7155 gnd.n99 585
R3057 gnd.n7156 gnd.n7153 585
R3058 gnd.n7157 gnd.n7149 585
R3059 gnd.n7147 gnd.n7145 585
R3060 gnd.n7161 gnd.n7144 585
R3061 gnd.n7162 gnd.n7142 585
R3062 gnd.n7163 gnd.n7141 585
R3063 gnd.n7139 gnd.n7137 585
R3064 gnd.n7167 gnd.n7136 585
R3065 gnd.n7168 gnd.n7134 585
R3066 gnd.n7169 gnd.n7133 585
R3067 gnd.n7131 gnd.n7129 585
R3068 gnd.n7173 gnd.n7128 585
R3069 gnd.n7174 gnd.n7126 585
R3070 gnd.n7175 gnd.n7125 585
R3071 gnd.n7123 gnd.n7121 585
R3072 gnd.n7179 gnd.n7120 585
R3073 gnd.n7180 gnd.n7118 585
R3074 gnd.n7181 gnd.n7117 585
R3075 gnd.n7117 gnd.n102 585
R3076 gnd.n7282 gnd.n7281 585
R3077 gnd.n7281 gnd.n7280 585
R3078 gnd.n7283 gnd.n97 585
R3079 gnd.n100 gnd.n97 585
R3080 gnd.n7284 gnd.n96 585
R3081 gnd.n7200 gnd.n96 585
R3082 gnd.n180 gnd.n94 585
R3083 gnd.n181 gnd.n180 585
R3084 gnd.n7288 gnd.n93 585
R3085 gnd.n7192 gnd.n93 585
R3086 gnd.n7289 gnd.n92 585
R3087 gnd.n188 gnd.n92 585
R3088 gnd.n7290 gnd.n91 585
R3089 gnd.n7109 gnd.n91 585
R3090 gnd.n206 gnd.n89 585
R3091 gnd.n207 gnd.n206 585
R3092 gnd.n7294 gnd.n88 585
R3093 gnd.n7101 gnd.n88 585
R3094 gnd.n7295 gnd.n87 585
R3095 gnd.n204 gnd.n87 585
R3096 gnd.n7296 gnd.n86 585
R3097 gnd.n7093 gnd.n86 585
R3098 gnd.n213 gnd.n84 585
R3099 gnd.n214 gnd.n213 585
R3100 gnd.n7300 gnd.n83 585
R3101 gnd.n7085 gnd.n83 585
R3102 gnd.n7301 gnd.n82 585
R3103 gnd.n221 gnd.n82 585
R3104 gnd.n7302 gnd.n81 585
R3105 gnd.n7077 gnd.n81 585
R3106 gnd.n236 gnd.n79 585
R3107 gnd.n237 gnd.n236 585
R3108 gnd.n7306 gnd.n78 585
R3109 gnd.n7069 gnd.n78 585
R3110 gnd.n7307 gnd.n77 585
R3111 gnd.n234 gnd.n77 585
R3112 gnd.n7308 gnd.n76 585
R3113 gnd.n7061 gnd.n76 585
R3114 gnd.n243 gnd.n74 585
R3115 gnd.n244 gnd.n243 585
R3116 gnd.n7312 gnd.n73 585
R3117 gnd.n7053 gnd.n73 585
R3118 gnd.n7313 gnd.n72 585
R3119 gnd.n251 gnd.n72 585
R3120 gnd.n7314 gnd.n71 585
R3121 gnd.n7045 gnd.n71 585
R3122 gnd.n7010 gnd.n69 585
R3123 gnd.n7011 gnd.n7010 585
R3124 gnd.n7318 gnd.n68 585
R3125 gnd.n7022 gnd.n68 585
R3126 gnd.n7319 gnd.n67 585
R3127 gnd.n7017 gnd.n67 585
R3128 gnd.n7320 gnd.n66 585
R3129 gnd.n6929 gnd.n66 585
R3130 gnd.n298 gnd.n65 585
R3131 gnd.n6952 gnd.n298 585
R3132 gnd.n6946 gnd.n6945 585
R3133 gnd.n6947 gnd.n6946 585
R3134 gnd.n304 gnd.n303 585
R3135 gnd.n308 gnd.n303 585
R3136 gnd.n6941 gnd.n6940 585
R3137 gnd.n6940 gnd.n6939 585
R3138 gnd.n306 gnd.n274 585
R3139 gnd.n7038 gnd.n274 585
R3140 gnd.n5551 gnd.n5549 585
R3141 gnd.n5549 gnd.n5548 585
R3142 gnd.n5552 gnd.n2803 585
R3143 gnd.n5587 gnd.n2803 585
R3144 gnd.n5553 gnd.n2828 585
R3145 gnd.n2828 gnd.n2813 585
R3146 gnd.n2825 gnd.n2812 585
R3147 gnd.n5579 gnd.n2812 585
R3148 gnd.n5558 gnd.n5557 585
R3149 gnd.n5560 gnd.n5558 585
R3150 gnd.n2824 gnd.n2823 585
R3151 gnd.n2823 gnd.n2821 585
R3152 gnd.n5495 gnd.n2836 585
R3153 gnd.n5525 gnd.n2836 585
R3154 gnd.n5496 gnd.n5494 585
R3155 gnd.n5494 gnd.n2847 585
R3156 gnd.n2859 gnd.n2846 585
R3157 gnd.n5515 gnd.n2846 585
R3158 gnd.n5501 gnd.n5500 585
R3159 gnd.n5502 gnd.n5501 585
R3160 gnd.n2858 gnd.n2857 585
R3161 gnd.n2857 gnd.n2855 585
R3162 gnd.n5490 gnd.n5489 585
R3163 gnd.n5489 gnd.n5488 585
R3164 gnd.n2862 gnd.n2861 585
R3165 gnd.n2876 gnd.n2862 585
R3166 gnd.n2887 gnd.n2874 585
R3167 gnd.n5478 gnd.n2874 585
R3168 gnd.n5465 gnd.n5464 585
R3169 gnd.n5466 gnd.n5465 585
R3170 gnd.n2886 gnd.n2885 585
R3171 gnd.n2885 gnd.n2883 585
R3172 gnd.n5459 gnd.n5458 585
R3173 gnd.n5458 gnd.n5457 585
R3174 gnd.n2890 gnd.n2889 585
R3175 gnd.n2904 gnd.n2890 585
R3176 gnd.n2957 gnd.n2903 585
R3177 gnd.n5447 gnd.n2903 585
R3178 gnd.n5434 gnd.n5433 585
R3179 gnd.n5435 gnd.n5434 585
R3180 gnd.n2956 gnd.n2955 585
R3181 gnd.n2955 gnd.n2923 585
R3182 gnd.n5428 gnd.n2773 585
R3183 gnd.n5622 gnd.n2773 585
R3184 gnd.n6138 gnd.n6137 585
R3185 gnd.n6139 gnd.n6138 585
R3186 gnd.n874 gnd.n872 585
R3187 gnd.n872 gnd.n868 585
R3188 gnd.n856 gnd.n855 585
R3189 gnd.n2221 gnd.n856 585
R3190 gnd.n6149 gnd.n6148 585
R3191 gnd.n6148 gnd.n6147 585
R3192 gnd.n6150 gnd.n850 585
R3193 gnd.n2175 gnd.n850 585
R3194 gnd.n6152 gnd.n6151 585
R3195 gnd.n6153 gnd.n6152 585
R3196 gnd.n851 gnd.n849 585
R3197 gnd.n2179 gnd.n849 585
R3198 gnd.n2203 gnd.n2202 585
R3199 gnd.n2202 gnd.n2201 585
R3200 gnd.n1242 gnd.n1241 585
R3201 gnd.n2185 gnd.n1242 585
R3202 gnd.n2159 gnd.n1261 585
R3203 gnd.n1261 gnd.n1260 585
R3204 gnd.n2161 gnd.n2160 585
R3205 gnd.n2162 gnd.n2161 585
R3206 gnd.n1262 gnd.n1259 585
R3207 gnd.n1270 gnd.n1259 585
R3208 gnd.n2135 gnd.n1282 585
R3209 gnd.n1282 gnd.n1269 585
R3210 gnd.n2137 gnd.n2136 585
R3211 gnd.n2138 gnd.n2137 585
R3212 gnd.n1283 gnd.n1281 585
R3213 gnd.n1281 gnd.n1277 585
R3214 gnd.n2123 gnd.n2122 585
R3215 gnd.n2122 gnd.n2121 585
R3216 gnd.n1288 gnd.n1287 585
R3217 gnd.n1298 gnd.n1288 585
R3218 gnd.n2112 gnd.n2111 585
R3219 gnd.n2111 gnd.n2110 585
R3220 gnd.n1295 gnd.n1294 585
R3221 gnd.n2098 gnd.n1295 585
R3222 gnd.n2072 gnd.n1316 585
R3223 gnd.n1316 gnd.n1305 585
R3224 gnd.n2074 gnd.n2073 585
R3225 gnd.n2075 gnd.n2074 585
R3226 gnd.n1317 gnd.n1315 585
R3227 gnd.n1325 gnd.n1315 585
R3228 gnd.n2050 gnd.n1337 585
R3229 gnd.n1337 gnd.n1324 585
R3230 gnd.n2052 gnd.n2051 585
R3231 gnd.n2053 gnd.n2052 585
R3232 gnd.n1338 gnd.n1336 585
R3233 gnd.n1336 gnd.n1332 585
R3234 gnd.n2038 gnd.n2037 585
R3235 gnd.n2037 gnd.n2036 585
R3236 gnd.n1343 gnd.n1342 585
R3237 gnd.n1352 gnd.n1343 585
R3238 gnd.n2027 gnd.n2026 585
R3239 gnd.n2026 gnd.n2025 585
R3240 gnd.n1350 gnd.n1349 585
R3241 gnd.n2013 gnd.n1350 585
R3242 gnd.n1451 gnd.n1450 585
R3243 gnd.n1451 gnd.n1359 585
R3244 gnd.n1970 gnd.n1969 585
R3245 gnd.n1969 gnd.n1968 585
R3246 gnd.n1971 gnd.n1445 585
R3247 gnd.n1456 gnd.n1445 585
R3248 gnd.n1973 gnd.n1972 585
R3249 gnd.n1974 gnd.n1973 585
R3250 gnd.n1446 gnd.n1444 585
R3251 gnd.n1469 gnd.n1444 585
R3252 gnd.n1429 gnd.n1428 585
R3253 gnd.n1432 gnd.n1429 585
R3254 gnd.n1984 gnd.n1983 585
R3255 gnd.n1983 gnd.n1982 585
R3256 gnd.n1985 gnd.n1423 585
R3257 gnd.n1944 gnd.n1423 585
R3258 gnd.n1987 gnd.n1986 585
R3259 gnd.n1988 gnd.n1987 585
R3260 gnd.n1424 gnd.n1422 585
R3261 gnd.n1483 gnd.n1422 585
R3262 gnd.n1936 gnd.n1935 585
R3263 gnd.n1935 gnd.n1934 585
R3264 gnd.n1480 gnd.n1479 585
R3265 gnd.n1918 gnd.n1480 585
R3266 gnd.n1905 gnd.n1499 585
R3267 gnd.n1499 gnd.n1498 585
R3268 gnd.n1907 gnd.n1906 585
R3269 gnd.n1908 gnd.n1907 585
R3270 gnd.n1500 gnd.n1497 585
R3271 gnd.n1506 gnd.n1497 585
R3272 gnd.n1886 gnd.n1885 585
R3273 gnd.n1887 gnd.n1886 585
R3274 gnd.n1517 gnd.n1516 585
R3275 gnd.n1516 gnd.n1512 585
R3276 gnd.n1876 gnd.n1875 585
R3277 gnd.n1877 gnd.n1876 585
R3278 gnd.n1527 gnd.n1526 585
R3279 gnd.n1532 gnd.n1526 585
R3280 gnd.n1854 gnd.n1545 585
R3281 gnd.n1545 gnd.n1531 585
R3282 gnd.n1856 gnd.n1855 585
R3283 gnd.n1857 gnd.n1856 585
R3284 gnd.n1546 gnd.n1544 585
R3285 gnd.n1544 gnd.n1540 585
R3286 gnd.n1845 gnd.n1844 585
R3287 gnd.n1846 gnd.n1845 585
R3288 gnd.n1553 gnd.n1552 585
R3289 gnd.n1557 gnd.n1552 585
R3290 gnd.n1822 gnd.n1574 585
R3291 gnd.n1574 gnd.n1556 585
R3292 gnd.n1824 gnd.n1823 585
R3293 gnd.n1825 gnd.n1824 585
R3294 gnd.n1575 gnd.n1573 585
R3295 gnd.n1573 gnd.n1564 585
R3296 gnd.n1817 gnd.n1816 585
R3297 gnd.n1816 gnd.n1815 585
R3298 gnd.n1622 gnd.n1621 585
R3299 gnd.n1623 gnd.n1622 585
R3300 gnd.n1776 gnd.n1775 585
R3301 gnd.n1777 gnd.n1776 585
R3302 gnd.n1632 gnd.n1631 585
R3303 gnd.n1631 gnd.n1630 585
R3304 gnd.n1771 gnd.n1770 585
R3305 gnd.n1770 gnd.n1769 585
R3306 gnd.n1635 gnd.n1634 585
R3307 gnd.n1636 gnd.n1635 585
R3308 gnd.n1760 gnd.n1759 585
R3309 gnd.n1761 gnd.n1760 585
R3310 gnd.n1643 gnd.n1642 585
R3311 gnd.n1752 gnd.n1642 585
R3312 gnd.n1755 gnd.n1754 585
R3313 gnd.n1754 gnd.n1753 585
R3314 gnd.n1646 gnd.n1645 585
R3315 gnd.n1647 gnd.n1646 585
R3316 gnd.n1741 gnd.n1740 585
R3317 gnd.n1739 gnd.n1665 585
R3318 gnd.n1738 gnd.n1664 585
R3319 gnd.n1743 gnd.n1664 585
R3320 gnd.n1737 gnd.n1736 585
R3321 gnd.n1735 gnd.n1734 585
R3322 gnd.n1733 gnd.n1732 585
R3323 gnd.n1731 gnd.n1730 585
R3324 gnd.n1729 gnd.n1728 585
R3325 gnd.n1727 gnd.n1726 585
R3326 gnd.n1725 gnd.n1724 585
R3327 gnd.n1723 gnd.n1722 585
R3328 gnd.n1721 gnd.n1720 585
R3329 gnd.n1719 gnd.n1718 585
R3330 gnd.n1717 gnd.n1716 585
R3331 gnd.n1715 gnd.n1714 585
R3332 gnd.n1713 gnd.n1712 585
R3333 gnd.n1711 gnd.n1710 585
R3334 gnd.n1709 gnd.n1708 585
R3335 gnd.n1707 gnd.n1706 585
R3336 gnd.n1705 gnd.n1704 585
R3337 gnd.n1703 gnd.n1702 585
R3338 gnd.n1701 gnd.n1700 585
R3339 gnd.n1699 gnd.n1698 585
R3340 gnd.n1697 gnd.n1696 585
R3341 gnd.n1695 gnd.n1694 585
R3342 gnd.n1652 gnd.n1651 585
R3343 gnd.n1746 gnd.n1745 585
R3344 gnd.n2229 gnd.n2228 585
R3345 gnd.n898 gnd.n897 585
R3346 gnd.n974 gnd.n973 585
R3347 gnd.n972 gnd.n971 585
R3348 gnd.n970 gnd.n969 585
R3349 gnd.n963 gnd.n903 585
R3350 gnd.n965 gnd.n964 585
R3351 gnd.n962 gnd.n961 585
R3352 gnd.n960 gnd.n959 585
R3353 gnd.n953 gnd.n905 585
R3354 gnd.n955 gnd.n954 585
R3355 gnd.n952 gnd.n951 585
R3356 gnd.n950 gnd.n949 585
R3357 gnd.n943 gnd.n907 585
R3358 gnd.n945 gnd.n944 585
R3359 gnd.n942 gnd.n941 585
R3360 gnd.n940 gnd.n939 585
R3361 gnd.n933 gnd.n909 585
R3362 gnd.n935 gnd.n934 585
R3363 gnd.n932 gnd.n931 585
R3364 gnd.n930 gnd.n929 585
R3365 gnd.n923 gnd.n911 585
R3366 gnd.n925 gnd.n924 585
R3367 gnd.n922 gnd.n921 585
R3368 gnd.n920 gnd.n919 585
R3369 gnd.n914 gnd.n913 585
R3370 gnd.n915 gnd.n873 585
R3371 gnd.n6123 gnd.n873 585
R3372 gnd.n2225 gnd.n870 585
R3373 gnd.n6139 gnd.n870 585
R3374 gnd.n2224 gnd.n2223 585
R3375 gnd.n2223 gnd.n868 585
R3376 gnd.n2222 gnd.n978 585
R3377 gnd.n2222 gnd.n2221 585
R3378 gnd.n2174 gnd.n858 585
R3379 gnd.n6147 gnd.n858 585
R3380 gnd.n2177 gnd.n2176 585
R3381 gnd.n2176 gnd.n2175 585
R3382 gnd.n2178 gnd.n847 585
R3383 gnd.n6153 gnd.n847 585
R3384 gnd.n2181 gnd.n2180 585
R3385 gnd.n2180 gnd.n2179 585
R3386 gnd.n2182 gnd.n1244 585
R3387 gnd.n2201 gnd.n1244 585
R3388 gnd.n2184 gnd.n2183 585
R3389 gnd.n2185 gnd.n2184 585
R3390 gnd.n1253 gnd.n1252 585
R3391 gnd.n1260 gnd.n1252 585
R3392 gnd.n2164 gnd.n2163 585
R3393 gnd.n2163 gnd.n2162 585
R3394 gnd.n1256 gnd.n1255 585
R3395 gnd.n1270 gnd.n1256 585
R3396 gnd.n2088 gnd.n2087 585
R3397 gnd.n2087 gnd.n1269 585
R3398 gnd.n2089 gnd.n1279 585
R3399 gnd.n2138 gnd.n1279 585
R3400 gnd.n2091 gnd.n2090 585
R3401 gnd.n2090 gnd.n1277 585
R3402 gnd.n2092 gnd.n1290 585
R3403 gnd.n2121 gnd.n1290 585
R3404 gnd.n2094 gnd.n2093 585
R3405 gnd.n2093 gnd.n1298 585
R3406 gnd.n2095 gnd.n1297 585
R3407 gnd.n2110 gnd.n1297 585
R3408 gnd.n2097 gnd.n2096 585
R3409 gnd.n2098 gnd.n2097 585
R3410 gnd.n1309 gnd.n1308 585
R3411 gnd.n1308 gnd.n1305 585
R3412 gnd.n2077 gnd.n2076 585
R3413 gnd.n2076 gnd.n2075 585
R3414 gnd.n1312 gnd.n1311 585
R3415 gnd.n1325 gnd.n1312 585
R3416 gnd.n2001 gnd.n2000 585
R3417 gnd.n2000 gnd.n1324 585
R3418 gnd.n2002 gnd.n1334 585
R3419 gnd.n2053 gnd.n1334 585
R3420 gnd.n2004 gnd.n2003 585
R3421 gnd.n2003 gnd.n1332 585
R3422 gnd.n2005 gnd.n1345 585
R3423 gnd.n2036 gnd.n1345 585
R3424 gnd.n2007 gnd.n2006 585
R3425 gnd.n2006 gnd.n1352 585
R3426 gnd.n2008 gnd.n1351 585
R3427 gnd.n2025 gnd.n1351 585
R3428 gnd.n2010 gnd.n2009 585
R3429 gnd.n2013 gnd.n2010 585
R3430 gnd.n1362 gnd.n1361 585
R3431 gnd.n1361 gnd.n1359 585
R3432 gnd.n1453 gnd.n1452 585
R3433 gnd.n1968 gnd.n1452 585
R3434 gnd.n1455 gnd.n1454 585
R3435 gnd.n1456 gnd.n1455 585
R3436 gnd.n1466 gnd.n1442 585
R3437 gnd.n1974 gnd.n1442 585
R3438 gnd.n1468 gnd.n1467 585
R3439 gnd.n1469 gnd.n1468 585
R3440 gnd.n1465 gnd.n1464 585
R3441 gnd.n1465 gnd.n1432 585
R3442 gnd.n1463 gnd.n1430 585
R3443 gnd.n1982 gnd.n1430 585
R3444 gnd.n1419 gnd.n1417 585
R3445 gnd.n1944 gnd.n1419 585
R3446 gnd.n1990 gnd.n1989 585
R3447 gnd.n1989 gnd.n1988 585
R3448 gnd.n1418 gnd.n1416 585
R3449 gnd.n1483 gnd.n1418 585
R3450 gnd.n1915 gnd.n1482 585
R3451 gnd.n1934 gnd.n1482 585
R3452 gnd.n1917 gnd.n1916 585
R3453 gnd.n1918 gnd.n1917 585
R3454 gnd.n1492 gnd.n1491 585
R3455 gnd.n1498 gnd.n1491 585
R3456 gnd.n1910 gnd.n1909 585
R3457 gnd.n1909 gnd.n1908 585
R3458 gnd.n1495 gnd.n1494 585
R3459 gnd.n1506 gnd.n1495 585
R3460 gnd.n1795 gnd.n1514 585
R3461 gnd.n1887 gnd.n1514 585
R3462 gnd.n1797 gnd.n1796 585
R3463 gnd.n1796 gnd.n1512 585
R3464 gnd.n1798 gnd.n1525 585
R3465 gnd.n1877 gnd.n1525 585
R3466 gnd.n1800 gnd.n1799 585
R3467 gnd.n1800 gnd.n1532 585
R3468 gnd.n1802 gnd.n1801 585
R3469 gnd.n1801 gnd.n1531 585
R3470 gnd.n1803 gnd.n1542 585
R3471 gnd.n1857 gnd.n1542 585
R3472 gnd.n1805 gnd.n1804 585
R3473 gnd.n1804 gnd.n1540 585
R3474 gnd.n1806 gnd.n1551 585
R3475 gnd.n1846 gnd.n1551 585
R3476 gnd.n1808 gnd.n1807 585
R3477 gnd.n1808 gnd.n1557 585
R3478 gnd.n1810 gnd.n1809 585
R3479 gnd.n1809 gnd.n1556 585
R3480 gnd.n1811 gnd.n1572 585
R3481 gnd.n1825 gnd.n1572 585
R3482 gnd.n1812 gnd.n1625 585
R3483 gnd.n1625 gnd.n1564 585
R3484 gnd.n1814 gnd.n1813 585
R3485 gnd.n1815 gnd.n1814 585
R3486 gnd.n1626 gnd.n1624 585
R3487 gnd.n1624 gnd.n1623 585
R3488 gnd.n1779 gnd.n1778 585
R3489 gnd.n1778 gnd.n1777 585
R3490 gnd.n1629 gnd.n1628 585
R3491 gnd.n1630 gnd.n1629 585
R3492 gnd.n1768 gnd.n1767 585
R3493 gnd.n1769 gnd.n1768 585
R3494 gnd.n1638 gnd.n1637 585
R3495 gnd.n1637 gnd.n1636 585
R3496 gnd.n1763 gnd.n1762 585
R3497 gnd.n1762 gnd.n1761 585
R3498 gnd.n1641 gnd.n1640 585
R3499 gnd.n1752 gnd.n1641 585
R3500 gnd.n1751 gnd.n1750 585
R3501 gnd.n1753 gnd.n1751 585
R3502 gnd.n1649 gnd.n1648 585
R3503 gnd.n1648 gnd.n1647 585
R3504 gnd.n867 gnd.n866 585
R3505 gnd.n871 gnd.n867 585
R3506 gnd.n6142 gnd.n6141 585
R3507 gnd.n6141 gnd.n6140 585
R3508 gnd.n6143 gnd.n861 585
R3509 gnd.n2220 gnd.n861 585
R3510 gnd.n6145 gnd.n6144 585
R3511 gnd.n6146 gnd.n6145 585
R3512 gnd.n862 gnd.n860 585
R3513 gnd.n860 gnd.n857 585
R3514 gnd.n2196 gnd.n2195 585
R3515 gnd.n2195 gnd.n848 585
R3516 gnd.n2197 gnd.n1246 585
R3517 gnd.n1246 gnd.n846 585
R3518 gnd.n2199 gnd.n2198 585
R3519 gnd.n2200 gnd.n2199 585
R3520 gnd.n1247 gnd.n1245 585
R3521 gnd.n1245 gnd.n1243 585
R3522 gnd.n2188 gnd.n2187 585
R3523 gnd.n2187 gnd.n2186 585
R3524 gnd.n1250 gnd.n1249 585
R3525 gnd.n1258 gnd.n1250 585
R3526 gnd.n2146 gnd.n1272 585
R3527 gnd.n1272 gnd.n1257 585
R3528 gnd.n2148 gnd.n2147 585
R3529 gnd.n2149 gnd.n2148 585
R3530 gnd.n1273 gnd.n1271 585
R3531 gnd.n1280 gnd.n1271 585
R3532 gnd.n2141 gnd.n2140 585
R3533 gnd.n2140 gnd.n2139 585
R3534 gnd.n1276 gnd.n1275 585
R3535 gnd.n2120 gnd.n1276 585
R3536 gnd.n2106 gnd.n1300 585
R3537 gnd.n1300 gnd.n1289 585
R3538 gnd.n2108 gnd.n2107 585
R3539 gnd.n2109 gnd.n2108 585
R3540 gnd.n1301 gnd.n1299 585
R3541 gnd.n1299 gnd.n1296 585
R3542 gnd.n2101 gnd.n2100 585
R3543 gnd.n2100 gnd.n2099 585
R3544 gnd.n1304 gnd.n1303 585
R3545 gnd.n1314 gnd.n1304 585
R3546 gnd.n2061 gnd.n1327 585
R3547 gnd.n1327 gnd.n1313 585
R3548 gnd.n2063 gnd.n2062 585
R3549 gnd.n2064 gnd.n2063 585
R3550 gnd.n1328 gnd.n1326 585
R3551 gnd.n1335 gnd.n1326 585
R3552 gnd.n2056 gnd.n2055 585
R3553 gnd.n2055 gnd.n2054 585
R3554 gnd.n1331 gnd.n1330 585
R3555 gnd.n2035 gnd.n1331 585
R3556 gnd.n2021 gnd.n1354 585
R3557 gnd.n1354 gnd.n1344 585
R3558 gnd.n2023 gnd.n2022 585
R3559 gnd.n2024 gnd.n2023 585
R3560 gnd.n1355 gnd.n1353 585
R3561 gnd.n2012 gnd.n1353 585
R3562 gnd.n2016 gnd.n2015 585
R3563 gnd.n2015 gnd.n2014 585
R3564 gnd.n1358 gnd.n1357 585
R3565 gnd.n1967 gnd.n1358 585
R3566 gnd.n1460 gnd.n1459 585
R3567 gnd.n1461 gnd.n1460 585
R3568 gnd.n1440 gnd.n1439 585
R3569 gnd.n1443 gnd.n1440 585
R3570 gnd.n1977 gnd.n1976 585
R3571 gnd.n1976 gnd.n1975 585
R3572 gnd.n1978 gnd.n1434 585
R3573 gnd.n1470 gnd.n1434 585
R3574 gnd.n1980 gnd.n1979 585
R3575 gnd.n1981 gnd.n1980 585
R3576 gnd.n1435 gnd.n1433 585
R3577 gnd.n1945 gnd.n1433 585
R3578 gnd.n1929 gnd.n1928 585
R3579 gnd.n1928 gnd.n1421 585
R3580 gnd.n1930 gnd.n1485 585
R3581 gnd.n1485 gnd.n1420 585
R3582 gnd.n1932 gnd.n1931 585
R3583 gnd.n1933 gnd.n1932 585
R3584 gnd.n1486 gnd.n1484 585
R3585 gnd.n1484 gnd.n1481 585
R3586 gnd.n1921 gnd.n1920 585
R3587 gnd.n1920 gnd.n1919 585
R3588 gnd.n1489 gnd.n1488 585
R3589 gnd.n1496 gnd.n1489 585
R3590 gnd.n1895 gnd.n1894 585
R3591 gnd.n1896 gnd.n1895 585
R3592 gnd.n1508 gnd.n1507 585
R3593 gnd.n1515 gnd.n1507 585
R3594 gnd.n1890 gnd.n1889 585
R3595 gnd.n1889 gnd.n1888 585
R3596 gnd.n1511 gnd.n1510 585
R3597 gnd.n1878 gnd.n1511 585
R3598 gnd.n1865 gnd.n1535 585
R3599 gnd.n1535 gnd.n1534 585
R3600 gnd.n1867 gnd.n1866 585
R3601 gnd.n1868 gnd.n1867 585
R3602 gnd.n1536 gnd.n1533 585
R3603 gnd.n1543 gnd.n1533 585
R3604 gnd.n1860 gnd.n1859 585
R3605 gnd.n1859 gnd.n1858 585
R3606 gnd.n1539 gnd.n1538 585
R3607 gnd.n1847 gnd.n1539 585
R3608 gnd.n1834 gnd.n1560 585
R3609 gnd.n1560 gnd.n1559 585
R3610 gnd.n1836 gnd.n1835 585
R3611 gnd.n1837 gnd.n1836 585
R3612 gnd.n1830 gnd.n1558 585
R3613 gnd.n1829 gnd.n1828 585
R3614 gnd.n1563 gnd.n1562 585
R3615 gnd.n1826 gnd.n1563 585
R3616 gnd.n1585 gnd.n1584 585
R3617 gnd.n1588 gnd.n1587 585
R3618 gnd.n1586 gnd.n1581 585
R3619 gnd.n1593 gnd.n1592 585
R3620 gnd.n1595 gnd.n1594 585
R3621 gnd.n1598 gnd.n1597 585
R3622 gnd.n1596 gnd.n1579 585
R3623 gnd.n1603 gnd.n1602 585
R3624 gnd.n1605 gnd.n1604 585
R3625 gnd.n1608 gnd.n1607 585
R3626 gnd.n1606 gnd.n1577 585
R3627 gnd.n1613 gnd.n1612 585
R3628 gnd.n1617 gnd.n1614 585
R3629 gnd.n1618 gnd.n1555 585
R3630 gnd.n6132 gnd.n6131 585
R3631 gnd.n6125 gnd.n881 585
R3632 gnd.n6127 gnd.n6126 585
R3633 gnd.n884 gnd.n883 585
R3634 gnd.n6097 gnd.n6096 585
R3635 gnd.n6099 gnd.n6098 585
R3636 gnd.n6101 gnd.n6100 585
R3637 gnd.n6103 gnd.n6102 585
R3638 gnd.n6105 gnd.n6104 585
R3639 gnd.n6107 gnd.n6106 585
R3640 gnd.n6109 gnd.n6108 585
R3641 gnd.n6111 gnd.n6110 585
R3642 gnd.n6113 gnd.n6112 585
R3643 gnd.n6116 gnd.n6115 585
R3644 gnd.n6114 gnd.n6086 585
R3645 gnd.n6120 gnd.n6083 585
R3646 gnd.n6122 gnd.n6121 585
R3647 gnd.n6123 gnd.n6122 585
R3648 gnd.n6134 gnd.n6133 585
R3649 gnd.n6133 gnd.n871 585
R3650 gnd.n877 gnd.n869 585
R3651 gnd.n6140 gnd.n869 585
R3652 gnd.n2219 gnd.n2218 585
R3653 gnd.n2220 gnd.n2219 585
R3654 gnd.n2213 gnd.n859 585
R3655 gnd.n6146 gnd.n859 585
R3656 gnd.n2212 gnd.n2211 585
R3657 gnd.n2211 gnd.n857 585
R3658 gnd.n2210 gnd.n1236 585
R3659 gnd.n2210 gnd.n848 585
R3660 gnd.n2209 gnd.n2208 585
R3661 gnd.n2209 gnd.n846 585
R3662 gnd.n1239 gnd.n1238 585
R3663 gnd.n2200 gnd.n1238 585
R3664 gnd.n2155 gnd.n2154 585
R3665 gnd.n2154 gnd.n1243 585
R3666 gnd.n2156 gnd.n1251 585
R3667 gnd.n2186 gnd.n1251 585
R3668 gnd.n2153 gnd.n2152 585
R3669 gnd.n2152 gnd.n1258 585
R3670 gnd.n2151 gnd.n1266 585
R3671 gnd.n2151 gnd.n1257 585
R3672 gnd.n2150 gnd.n1268 585
R3673 gnd.n2150 gnd.n2149 585
R3674 gnd.n2129 gnd.n1267 585
R3675 gnd.n1280 gnd.n1267 585
R3676 gnd.n2128 gnd.n1278 585
R3677 gnd.n2139 gnd.n1278 585
R3678 gnd.n2119 gnd.n1285 585
R3679 gnd.n2120 gnd.n2119 585
R3680 gnd.n2118 gnd.n2117 585
R3681 gnd.n2118 gnd.n1289 585
R3682 gnd.n2116 gnd.n1291 585
R3683 gnd.n2109 gnd.n1291 585
R3684 gnd.n1306 gnd.n1292 585
R3685 gnd.n1306 gnd.n1296 585
R3686 gnd.n2069 gnd.n1307 585
R3687 gnd.n2099 gnd.n1307 585
R3688 gnd.n2068 gnd.n2067 585
R3689 gnd.n2067 gnd.n1314 585
R3690 gnd.n2066 gnd.n1321 585
R3691 gnd.n2066 gnd.n1313 585
R3692 gnd.n2065 gnd.n1323 585
R3693 gnd.n2065 gnd.n2064 585
R3694 gnd.n2044 gnd.n1322 585
R3695 gnd.n1335 gnd.n1322 585
R3696 gnd.n2043 gnd.n1333 585
R3697 gnd.n2054 gnd.n1333 585
R3698 gnd.n2034 gnd.n1340 585
R3699 gnd.n2035 gnd.n2034 585
R3700 gnd.n2033 gnd.n2032 585
R3701 gnd.n2033 gnd.n1344 585
R3702 gnd.n2031 gnd.n1346 585
R3703 gnd.n2024 gnd.n1346 585
R3704 gnd.n2011 gnd.n1347 585
R3705 gnd.n2012 gnd.n2011 585
R3706 gnd.n1964 gnd.n1360 585
R3707 gnd.n2014 gnd.n1360 585
R3708 gnd.n1966 gnd.n1965 585
R3709 gnd.n1967 gnd.n1966 585
R3710 gnd.n1959 gnd.n1462 585
R3711 gnd.n1462 gnd.n1461 585
R3712 gnd.n1957 gnd.n1956 585
R3713 gnd.n1956 gnd.n1443 585
R3714 gnd.n1954 gnd.n1441 585
R3715 gnd.n1975 gnd.n1441 585
R3716 gnd.n1472 gnd.n1471 585
R3717 gnd.n1471 gnd.n1470 585
R3718 gnd.n1948 gnd.n1431 585
R3719 gnd.n1981 gnd.n1431 585
R3720 gnd.n1947 gnd.n1946 585
R3721 gnd.n1946 gnd.n1945 585
R3722 gnd.n1943 gnd.n1474 585
R3723 gnd.n1943 gnd.n1421 585
R3724 gnd.n1942 gnd.n1941 585
R3725 gnd.n1942 gnd.n1420 585
R3726 gnd.n1477 gnd.n1476 585
R3727 gnd.n1933 gnd.n1476 585
R3728 gnd.n1901 gnd.n1900 585
R3729 gnd.n1900 gnd.n1481 585
R3730 gnd.n1902 gnd.n1490 585
R3731 gnd.n1919 gnd.n1490 585
R3732 gnd.n1899 gnd.n1898 585
R3733 gnd.n1898 gnd.n1496 585
R3734 gnd.n1897 gnd.n1504 585
R3735 gnd.n1897 gnd.n1896 585
R3736 gnd.n1882 gnd.n1505 585
R3737 gnd.n1515 gnd.n1505 585
R3738 gnd.n1881 gnd.n1513 585
R3739 gnd.n1888 gnd.n1513 585
R3740 gnd.n1880 gnd.n1879 585
R3741 gnd.n1879 gnd.n1878 585
R3742 gnd.n1524 gnd.n1521 585
R3743 gnd.n1534 gnd.n1524 585
R3744 gnd.n1870 gnd.n1869 585
R3745 gnd.n1869 gnd.n1868 585
R3746 gnd.n1530 gnd.n1529 585
R3747 gnd.n1543 gnd.n1530 585
R3748 gnd.n1850 gnd.n1541 585
R3749 gnd.n1858 gnd.n1541 585
R3750 gnd.n1849 gnd.n1848 585
R3751 gnd.n1848 gnd.n1847 585
R3752 gnd.n1550 gnd.n1548 585
R3753 gnd.n1559 gnd.n1550 585
R3754 gnd.n1839 gnd.n1838 585
R3755 gnd.n1838 gnd.n1837 585
R3756 gnd.n5840 gnd.n5839 585
R3757 gnd.n5839 gnd.n5838 585
R3758 gnd.n5841 gnd.n2563 585
R3759 gnd.n4092 gnd.n2563 585
R3760 gnd.n5843 gnd.n5842 585
R3761 gnd.n5844 gnd.n5843 585
R3762 gnd.n2548 gnd.n2547 585
R3763 gnd.n4084 gnd.n2548 585
R3764 gnd.n5852 gnd.n5851 585
R3765 gnd.n5851 gnd.n5850 585
R3766 gnd.n5853 gnd.n2542 585
R3767 gnd.n4075 gnd.n2542 585
R3768 gnd.n5855 gnd.n5854 585
R3769 gnd.n5856 gnd.n5855 585
R3770 gnd.n2526 gnd.n2525 585
R3771 gnd.n4067 gnd.n2526 585
R3772 gnd.n5864 gnd.n5863 585
R3773 gnd.n5863 gnd.n5862 585
R3774 gnd.n5865 gnd.n2520 585
R3775 gnd.n4059 gnd.n2520 585
R3776 gnd.n5867 gnd.n5866 585
R3777 gnd.n5868 gnd.n5867 585
R3778 gnd.n2505 gnd.n2504 585
R3779 gnd.n4051 gnd.n2505 585
R3780 gnd.n5876 gnd.n5875 585
R3781 gnd.n5875 gnd.n5874 585
R3782 gnd.n5877 gnd.n2499 585
R3783 gnd.n4043 gnd.n2499 585
R3784 gnd.n5879 gnd.n5878 585
R3785 gnd.n5880 gnd.n5879 585
R3786 gnd.n2483 gnd.n2482 585
R3787 gnd.n4035 gnd.n2483 585
R3788 gnd.n5888 gnd.n5887 585
R3789 gnd.n5887 gnd.n5886 585
R3790 gnd.n5889 gnd.n2477 585
R3791 gnd.n4027 gnd.n2477 585
R3792 gnd.n5891 gnd.n5890 585
R3793 gnd.n5892 gnd.n5891 585
R3794 gnd.n2462 gnd.n2461 585
R3795 gnd.n4019 gnd.n2462 585
R3796 gnd.n5900 gnd.n5899 585
R3797 gnd.n5899 gnd.n5898 585
R3798 gnd.n5901 gnd.n2457 585
R3799 gnd.n4011 gnd.n2457 585
R3800 gnd.n5903 gnd.n5902 585
R3801 gnd.n5904 gnd.n5903 585
R3802 gnd.n2458 gnd.n2441 585
R3803 gnd.n4003 gnd.n2441 585
R3804 gnd.n5912 gnd.n5911 585
R3805 gnd.n5911 gnd.n5910 585
R3806 gnd.n5913 gnd.n2438 585
R3807 gnd.n3995 gnd.n2438 585
R3808 gnd.n5916 gnd.n5915 585
R3809 gnd.n5917 gnd.n5916 585
R3810 gnd.n2439 gnd.n2423 585
R3811 gnd.n3986 gnd.n2423 585
R3812 gnd.n5925 gnd.n5924 585
R3813 gnd.n5924 gnd.n5923 585
R3814 gnd.n5926 gnd.n2419 585
R3815 gnd.n3976 gnd.n2419 585
R3816 gnd.n5928 gnd.n5927 585
R3817 gnd.n5929 gnd.n5928 585
R3818 gnd.n2404 gnd.n2403 585
R3819 gnd.n3968 gnd.n2404 585
R3820 gnd.n5937 gnd.n5936 585
R3821 gnd.n5936 gnd.n5935 585
R3822 gnd.n5938 gnd.n2398 585
R3823 gnd.n2405 gnd.n2398 585
R3824 gnd.n5940 gnd.n5939 585
R3825 gnd.n5941 gnd.n5940 585
R3826 gnd.n2385 gnd.n2384 585
R3827 gnd.n2395 gnd.n2385 585
R3828 gnd.n5949 gnd.n5948 585
R3829 gnd.n5948 gnd.n5947 585
R3830 gnd.n5950 gnd.n2379 585
R3831 gnd.n2379 gnd.n2378 585
R3832 gnd.n5952 gnd.n5951 585
R3833 gnd.n5953 gnd.n5952 585
R3834 gnd.n2364 gnd.n2363 585
R3835 gnd.n2368 gnd.n2364 585
R3836 gnd.n5961 gnd.n5960 585
R3837 gnd.n5960 gnd.n5959 585
R3838 gnd.n5962 gnd.n2358 585
R3839 gnd.n2365 gnd.n2358 585
R3840 gnd.n5964 gnd.n5963 585
R3841 gnd.n5965 gnd.n5964 585
R3842 gnd.n2345 gnd.n2344 585
R3843 gnd.n2355 gnd.n2345 585
R3844 gnd.n5973 gnd.n5972 585
R3845 gnd.n5972 gnd.n5971 585
R3846 gnd.n5974 gnd.n2339 585
R3847 gnd.n2339 gnd.n2338 585
R3848 gnd.n5976 gnd.n5975 585
R3849 gnd.n5977 gnd.n5976 585
R3850 gnd.n2324 gnd.n2323 585
R3851 gnd.n2327 gnd.n2324 585
R3852 gnd.n5985 gnd.n5984 585
R3853 gnd.n5984 gnd.n5983 585
R3854 gnd.n5986 gnd.n2318 585
R3855 gnd.n2318 gnd.n2315 585
R3856 gnd.n5988 gnd.n5987 585
R3857 gnd.n5989 gnd.n5988 585
R3858 gnd.n2319 gnd.n2317 585
R3859 gnd.n2317 gnd.n2313 585
R3860 gnd.n3880 gnd.n3879 585
R3861 gnd.n3881 gnd.n3880 585
R3862 gnd.n3875 gnd.n2262 585
R3863 gnd.n2262 gnd.n2259 585
R3864 gnd.n6074 gnd.n6073 585
R3865 gnd.n6072 gnd.n2261 585
R3866 gnd.n6071 gnd.n2260 585
R3867 gnd.n6076 gnd.n2260 585
R3868 gnd.n6070 gnd.n6069 585
R3869 gnd.n6068 gnd.n6067 585
R3870 gnd.n6066 gnd.n6065 585
R3871 gnd.n6064 gnd.n6063 585
R3872 gnd.n6062 gnd.n6061 585
R3873 gnd.n6060 gnd.n6059 585
R3874 gnd.n6058 gnd.n6057 585
R3875 gnd.n6056 gnd.n6055 585
R3876 gnd.n6054 gnd.n6053 585
R3877 gnd.n6052 gnd.n6051 585
R3878 gnd.n6050 gnd.n6049 585
R3879 gnd.n6048 gnd.n6047 585
R3880 gnd.n6046 gnd.n6045 585
R3881 gnd.n6044 gnd.n6043 585
R3882 gnd.n6042 gnd.n6041 585
R3883 gnd.n6039 gnd.n6038 585
R3884 gnd.n6037 gnd.n6036 585
R3885 gnd.n6035 gnd.n6034 585
R3886 gnd.n6033 gnd.n6032 585
R3887 gnd.n6031 gnd.n6030 585
R3888 gnd.n6029 gnd.n6028 585
R3889 gnd.n6027 gnd.n6026 585
R3890 gnd.n6025 gnd.n6024 585
R3891 gnd.n6023 gnd.n6022 585
R3892 gnd.n6021 gnd.n6020 585
R3893 gnd.n6019 gnd.n6018 585
R3894 gnd.n6017 gnd.n6016 585
R3895 gnd.n6015 gnd.n6014 585
R3896 gnd.n6013 gnd.n6012 585
R3897 gnd.n6011 gnd.n6010 585
R3898 gnd.n6009 gnd.n6008 585
R3899 gnd.n6007 gnd.n6006 585
R3900 gnd.n6005 gnd.n6004 585
R3901 gnd.n6003 gnd.n2301 585
R3902 gnd.n2305 gnd.n2302 585
R3903 gnd.n5999 gnd.n5998 585
R3904 gnd.n3633 gnd.n3632 585
R3905 gnd.n4100 gnd.n4099 585
R3906 gnd.n4102 gnd.n4101 585
R3907 gnd.n4104 gnd.n4103 585
R3908 gnd.n4106 gnd.n4105 585
R3909 gnd.n4108 gnd.n4107 585
R3910 gnd.n4110 gnd.n4109 585
R3911 gnd.n4112 gnd.n4111 585
R3912 gnd.n4114 gnd.n4113 585
R3913 gnd.n4116 gnd.n4115 585
R3914 gnd.n4118 gnd.n4117 585
R3915 gnd.n4120 gnd.n4119 585
R3916 gnd.n4122 gnd.n4121 585
R3917 gnd.n4124 gnd.n4123 585
R3918 gnd.n4126 gnd.n4125 585
R3919 gnd.n4128 gnd.n4127 585
R3920 gnd.n4130 gnd.n4129 585
R3921 gnd.n4132 gnd.n4131 585
R3922 gnd.n4134 gnd.n4133 585
R3923 gnd.n4137 gnd.n4136 585
R3924 gnd.n4135 gnd.n3611 585
R3925 gnd.n4350 gnd.n4349 585
R3926 gnd.n4352 gnd.n4351 585
R3927 gnd.n4354 gnd.n4353 585
R3928 gnd.n4356 gnd.n4355 585
R3929 gnd.n4358 gnd.n4357 585
R3930 gnd.n4360 gnd.n4359 585
R3931 gnd.n4362 gnd.n4361 585
R3932 gnd.n4364 gnd.n4363 585
R3933 gnd.n4366 gnd.n4365 585
R3934 gnd.n4368 gnd.n4367 585
R3935 gnd.n4370 gnd.n4369 585
R3936 gnd.n4372 gnd.n4371 585
R3937 gnd.n4373 gnd.n3592 585
R3938 gnd.n4375 gnd.n4374 585
R3939 gnd.n3593 gnd.n3591 585
R3940 gnd.n3594 gnd.n2568 585
R3941 gnd.n4377 gnd.n2568 585
R3942 gnd.n4095 gnd.n2570 585
R3943 gnd.n5838 gnd.n2570 585
R3944 gnd.n4094 gnd.n4093 585
R3945 gnd.n4093 gnd.n4092 585
R3946 gnd.n3637 gnd.n2561 585
R3947 gnd.n5844 gnd.n2561 585
R3948 gnd.n4083 gnd.n4082 585
R3949 gnd.n4084 gnd.n4083 585
R3950 gnd.n3643 gnd.n2550 585
R3951 gnd.n5850 gnd.n2550 585
R3952 gnd.n4077 gnd.n4076 585
R3953 gnd.n4076 gnd.n4075 585
R3954 gnd.n3645 gnd.n2539 585
R3955 gnd.n5856 gnd.n2539 585
R3956 gnd.n4066 gnd.n4065 585
R3957 gnd.n4067 gnd.n4066 585
R3958 gnd.n3649 gnd.n2528 585
R3959 gnd.n5862 gnd.n2528 585
R3960 gnd.n4061 gnd.n4060 585
R3961 gnd.n4060 gnd.n4059 585
R3962 gnd.n3651 gnd.n2517 585
R3963 gnd.n5868 gnd.n2517 585
R3964 gnd.n4050 gnd.n4049 585
R3965 gnd.n4051 gnd.n4050 585
R3966 gnd.n3656 gnd.n2507 585
R3967 gnd.n5874 gnd.n2507 585
R3968 gnd.n4045 gnd.n4044 585
R3969 gnd.n4044 gnd.n4043 585
R3970 gnd.n3658 gnd.n2496 585
R3971 gnd.n5880 gnd.n2496 585
R3972 gnd.n4034 gnd.n4033 585
R3973 gnd.n4035 gnd.n4034 585
R3974 gnd.n3662 gnd.n2485 585
R3975 gnd.n5886 gnd.n2485 585
R3976 gnd.n4029 gnd.n4028 585
R3977 gnd.n4028 gnd.n4027 585
R3978 gnd.n3664 gnd.n2474 585
R3979 gnd.n5892 gnd.n2474 585
R3980 gnd.n4018 gnd.n4017 585
R3981 gnd.n4019 gnd.n4018 585
R3982 gnd.n3669 gnd.n2464 585
R3983 gnd.n5898 gnd.n2464 585
R3984 gnd.n4013 gnd.n4012 585
R3985 gnd.n4012 gnd.n4011 585
R3986 gnd.n3671 gnd.n2454 585
R3987 gnd.n5904 gnd.n2454 585
R3988 gnd.n4002 gnd.n4001 585
R3989 gnd.n4003 gnd.n4002 585
R3990 gnd.n3675 gnd.n2443 585
R3991 gnd.n5910 gnd.n2443 585
R3992 gnd.n3997 gnd.n3996 585
R3993 gnd.n3996 gnd.n3995 585
R3994 gnd.n3677 gnd.n2435 585
R3995 gnd.n5917 gnd.n2435 585
R3996 gnd.n3985 gnd.n3984 585
R3997 gnd.n3986 gnd.n3985 585
R3998 gnd.n3786 gnd.n2425 585
R3999 gnd.n5923 gnd.n2425 585
R4000 gnd.n3978 gnd.n3977 585
R4001 gnd.n3977 gnd.n3976 585
R4002 gnd.n3788 gnd.n2416 585
R4003 gnd.n5929 gnd.n2416 585
R4004 gnd.n3967 gnd.n3966 585
R4005 gnd.n3968 gnd.n3967 585
R4006 gnd.n3923 gnd.n2406 585
R4007 gnd.n5935 gnd.n2406 585
R4008 gnd.n3962 gnd.n3961 585
R4009 gnd.n3961 gnd.n2405 585
R4010 gnd.n3960 gnd.n2396 585
R4011 gnd.n5941 gnd.n2396 585
R4012 gnd.n3959 gnd.n3958 585
R4013 gnd.n3958 gnd.n2395 585
R4014 gnd.n3925 gnd.n2386 585
R4015 gnd.n5947 gnd.n2386 585
R4016 gnd.n3954 gnd.n3953 585
R4017 gnd.n3953 gnd.n2378 585
R4018 gnd.n3952 gnd.n2376 585
R4019 gnd.n5953 gnd.n2376 585
R4020 gnd.n3951 gnd.n3950 585
R4021 gnd.n3950 gnd.n2368 585
R4022 gnd.n3927 gnd.n2366 585
R4023 gnd.n5959 gnd.n2366 585
R4024 gnd.n3946 gnd.n3945 585
R4025 gnd.n3945 gnd.n2365 585
R4026 gnd.n3944 gnd.n2356 585
R4027 gnd.n5965 gnd.n2356 585
R4028 gnd.n3943 gnd.n3942 585
R4029 gnd.n3942 gnd.n2355 585
R4030 gnd.n3929 gnd.n2346 585
R4031 gnd.n5971 gnd.n2346 585
R4032 gnd.n3938 gnd.n3937 585
R4033 gnd.n3937 gnd.n2338 585
R4034 gnd.n3936 gnd.n2336 585
R4035 gnd.n5977 gnd.n2336 585
R4036 gnd.n3935 gnd.n3934 585
R4037 gnd.n3934 gnd.n2327 585
R4038 gnd.n3931 gnd.n2325 585
R4039 gnd.n5983 gnd.n2325 585
R4040 gnd.n2312 gnd.n2310 585
R4041 gnd.n2315 gnd.n2312 585
R4042 gnd.n5991 gnd.n5990 585
R4043 gnd.n5990 gnd.n5989 585
R4044 gnd.n2311 gnd.n2308 585
R4045 gnd.n2313 gnd.n2311 585
R4046 gnd.n5995 gnd.n2307 585
R4047 gnd.n3881 gnd.n2307 585
R4048 gnd.n5997 gnd.n5996 585
R4049 gnd.n5997 gnd.n2259 585
R4050 gnd.n7279 gnd.n7278 585
R4051 gnd.n7280 gnd.n7279 585
R4052 gnd.n106 gnd.n104 585
R4053 gnd.n104 gnd.n100 585
R4054 gnd.n7199 gnd.n7198 585
R4055 gnd.n7200 gnd.n7199 585
R4056 gnd.n184 gnd.n183 585
R4057 gnd.n183 gnd.n181 585
R4058 gnd.n7194 gnd.n7193 585
R4059 gnd.n7193 gnd.n7192 585
R4060 gnd.n187 gnd.n186 585
R4061 gnd.n188 gnd.n187 585
R4062 gnd.n7108 gnd.n7107 585
R4063 gnd.n7109 gnd.n7108 585
R4064 gnd.n200 gnd.n199 585
R4065 gnd.n207 gnd.n199 585
R4066 gnd.n7103 gnd.n7102 585
R4067 gnd.n7102 gnd.n7101 585
R4068 gnd.n203 gnd.n202 585
R4069 gnd.n204 gnd.n203 585
R4070 gnd.n7092 gnd.n7091 585
R4071 gnd.n7093 gnd.n7092 585
R4072 gnd.n217 gnd.n216 585
R4073 gnd.n216 gnd.n214 585
R4074 gnd.n7087 gnd.n7086 585
R4075 gnd.n7086 gnd.n7085 585
R4076 gnd.n220 gnd.n219 585
R4077 gnd.n221 gnd.n220 585
R4078 gnd.n7076 gnd.n7075 585
R4079 gnd.n7077 gnd.n7076 585
R4080 gnd.n230 gnd.n229 585
R4081 gnd.n237 gnd.n229 585
R4082 gnd.n7071 gnd.n7070 585
R4083 gnd.n7070 gnd.n7069 585
R4084 gnd.n233 gnd.n232 585
R4085 gnd.n234 gnd.n233 585
R4086 gnd.n7060 gnd.n7059 585
R4087 gnd.n7061 gnd.n7060 585
R4088 gnd.n247 gnd.n246 585
R4089 gnd.n246 gnd.n244 585
R4090 gnd.n7055 gnd.n7054 585
R4091 gnd.n7054 gnd.n7053 585
R4092 gnd.n250 gnd.n249 585
R4093 gnd.n251 gnd.n250 585
R4094 gnd.n7044 gnd.n7043 585
R4095 gnd.n7045 gnd.n7044 585
R4096 gnd.n261 gnd.n260 585
R4097 gnd.n7011 gnd.n260 585
R4098 gnd.n7021 gnd.n7020 585
R4099 gnd.n7022 gnd.n7021 585
R4100 gnd.n7019 gnd.n7018 585
R4101 gnd.n7018 gnd.n7017 585
R4102 gnd.n6949 gnd.n292 585
R4103 gnd.n6929 gnd.n292 585
R4104 gnd.n6951 gnd.n6950 585
R4105 gnd.n6952 gnd.n6951 585
R4106 gnd.n6948 gnd.n301 585
R4107 gnd.n6948 gnd.n6947 585
R4108 gnd.n300 gnd.n267 585
R4109 gnd.n308 gnd.n300 585
R4110 gnd.n271 gnd.n268 585
R4111 gnd.n6939 gnd.n271 585
R4112 gnd.n7040 gnd.n7039 585
R4113 gnd.n7039 gnd.n7038 585
R4114 gnd.n270 gnd.n269 585
R4115 gnd.n5548 gnd.n270 585
R4116 gnd.n5586 gnd.n5585 585
R4117 gnd.n5587 gnd.n5586 585
R4118 gnd.n2806 gnd.n2805 585
R4119 gnd.n2813 gnd.n2805 585
R4120 gnd.n5581 gnd.n5580 585
R4121 gnd.n5580 gnd.n5579 585
R4122 gnd.n2809 gnd.n2808 585
R4123 gnd.n5560 gnd.n2809 585
R4124 gnd.n5522 gnd.n2839 585
R4125 gnd.n2839 gnd.n2821 585
R4126 gnd.n5524 gnd.n5523 585
R4127 gnd.n5525 gnd.n5524 585
R4128 gnd.n2840 gnd.n2838 585
R4129 gnd.n2847 gnd.n2838 585
R4130 gnd.n5517 gnd.n5516 585
R4131 gnd.n5516 gnd.n5515 585
R4132 gnd.n2843 gnd.n2842 585
R4133 gnd.n5502 gnd.n2843 585
R4134 gnd.n5485 gnd.n2867 585
R4135 gnd.n2867 gnd.n2855 585
R4136 gnd.n5487 gnd.n5486 585
R4137 gnd.n5488 gnd.n5487 585
R4138 gnd.n2868 gnd.n2866 585
R4139 gnd.n2876 gnd.n2866 585
R4140 gnd.n5480 gnd.n5479 585
R4141 gnd.n5479 gnd.n5478 585
R4142 gnd.n2871 gnd.n2870 585
R4143 gnd.n5466 gnd.n2871 585
R4144 gnd.n5454 gnd.n2896 585
R4145 gnd.n2896 gnd.n2883 585
R4146 gnd.n5456 gnd.n5455 585
R4147 gnd.n5457 gnd.n5456 585
R4148 gnd.n2897 gnd.n2895 585
R4149 gnd.n2904 gnd.n2895 585
R4150 gnd.n5449 gnd.n5448 585
R4151 gnd.n5448 gnd.n5447 585
R4152 gnd.n2900 gnd.n2899 585
R4153 gnd.n5435 gnd.n2900 585
R4154 gnd.n2922 gnd.n2921 585
R4155 gnd.n2923 gnd.n2922 585
R4156 gnd.n2918 gnd.n2724 585
R4157 gnd.n5622 gnd.n2724 585
R4158 gnd.n5696 gnd.n5695 585
R4159 gnd.n5694 gnd.n2723 585
R4160 gnd.n5693 gnd.n2722 585
R4161 gnd.n5698 gnd.n2722 585
R4162 gnd.n5692 gnd.n5691 585
R4163 gnd.n5690 gnd.n5689 585
R4164 gnd.n5688 gnd.n5687 585
R4165 gnd.n5686 gnd.n5685 585
R4166 gnd.n5684 gnd.n5683 585
R4167 gnd.n5682 gnd.n5681 585
R4168 gnd.n5680 gnd.n5679 585
R4169 gnd.n5678 gnd.n5677 585
R4170 gnd.n5676 gnd.n5675 585
R4171 gnd.n5674 gnd.n5673 585
R4172 gnd.n5672 gnd.n5671 585
R4173 gnd.n5670 gnd.n5669 585
R4174 gnd.n5668 gnd.n5667 585
R4175 gnd.n5665 gnd.n5664 585
R4176 gnd.n5663 gnd.n5662 585
R4177 gnd.n5661 gnd.n5660 585
R4178 gnd.n5659 gnd.n5658 585
R4179 gnd.n5657 gnd.n5656 585
R4180 gnd.n5655 gnd.n5654 585
R4181 gnd.n5653 gnd.n5652 585
R4182 gnd.n5651 gnd.n5650 585
R4183 gnd.n5649 gnd.n5648 585
R4184 gnd.n5647 gnd.n5646 585
R4185 gnd.n5645 gnd.n5644 585
R4186 gnd.n5643 gnd.n5642 585
R4187 gnd.n5641 gnd.n5640 585
R4188 gnd.n5639 gnd.n5638 585
R4189 gnd.n5637 gnd.n5636 585
R4190 gnd.n5635 gnd.n5634 585
R4191 gnd.n5633 gnd.n5632 585
R4192 gnd.n5631 gnd.n5630 585
R4193 gnd.n5629 gnd.n2764 585
R4194 gnd.n2768 gnd.n2765 585
R4195 gnd.n5625 gnd.n5624 585
R4196 gnd.n174 gnd.n173 585
R4197 gnd.n7208 gnd.n169 585
R4198 gnd.n7210 gnd.n7209 585
R4199 gnd.n7212 gnd.n167 585
R4200 gnd.n7214 gnd.n7213 585
R4201 gnd.n7215 gnd.n162 585
R4202 gnd.n7217 gnd.n7216 585
R4203 gnd.n7219 gnd.n160 585
R4204 gnd.n7221 gnd.n7220 585
R4205 gnd.n7222 gnd.n155 585
R4206 gnd.n7224 gnd.n7223 585
R4207 gnd.n7226 gnd.n153 585
R4208 gnd.n7228 gnd.n7227 585
R4209 gnd.n7229 gnd.n148 585
R4210 gnd.n7231 gnd.n7230 585
R4211 gnd.n7233 gnd.n146 585
R4212 gnd.n7235 gnd.n7234 585
R4213 gnd.n7236 gnd.n141 585
R4214 gnd.n7238 gnd.n7237 585
R4215 gnd.n7240 gnd.n139 585
R4216 gnd.n7242 gnd.n7241 585
R4217 gnd.n7246 gnd.n134 585
R4218 gnd.n7248 gnd.n7247 585
R4219 gnd.n7250 gnd.n132 585
R4220 gnd.n7252 gnd.n7251 585
R4221 gnd.n7253 gnd.n127 585
R4222 gnd.n7255 gnd.n7254 585
R4223 gnd.n7257 gnd.n125 585
R4224 gnd.n7259 gnd.n7258 585
R4225 gnd.n7260 gnd.n120 585
R4226 gnd.n7262 gnd.n7261 585
R4227 gnd.n7264 gnd.n118 585
R4228 gnd.n7266 gnd.n7265 585
R4229 gnd.n7267 gnd.n113 585
R4230 gnd.n7269 gnd.n7268 585
R4231 gnd.n7271 gnd.n111 585
R4232 gnd.n7273 gnd.n7272 585
R4233 gnd.n7274 gnd.n109 585
R4234 gnd.n7275 gnd.n105 585
R4235 gnd.n105 gnd.n102 585
R4236 gnd.n7204 gnd.n101 585
R4237 gnd.n7280 gnd.n101 585
R4238 gnd.n7203 gnd.n7202 585
R4239 gnd.n7202 gnd.n100 585
R4240 gnd.n7201 gnd.n178 585
R4241 gnd.n7201 gnd.n7200 585
R4242 gnd.n6981 gnd.n179 585
R4243 gnd.n181 gnd.n179 585
R4244 gnd.n6982 gnd.n189 585
R4245 gnd.n7192 gnd.n189 585
R4246 gnd.n6984 gnd.n6983 585
R4247 gnd.n6983 gnd.n188 585
R4248 gnd.n6985 gnd.n198 585
R4249 gnd.n7109 gnd.n198 585
R4250 gnd.n6987 gnd.n6986 585
R4251 gnd.n6986 gnd.n207 585
R4252 gnd.n6988 gnd.n205 585
R4253 gnd.n7101 gnd.n205 585
R4254 gnd.n6990 gnd.n6989 585
R4255 gnd.n6989 gnd.n204 585
R4256 gnd.n6991 gnd.n215 585
R4257 gnd.n7093 gnd.n215 585
R4258 gnd.n6993 gnd.n6992 585
R4259 gnd.n6992 gnd.n214 585
R4260 gnd.n6994 gnd.n222 585
R4261 gnd.n7085 gnd.n222 585
R4262 gnd.n6996 gnd.n6995 585
R4263 gnd.n6995 gnd.n221 585
R4264 gnd.n6997 gnd.n228 585
R4265 gnd.n7077 gnd.n228 585
R4266 gnd.n6999 gnd.n6998 585
R4267 gnd.n6998 gnd.n237 585
R4268 gnd.n7000 gnd.n235 585
R4269 gnd.n7069 gnd.n235 585
R4270 gnd.n7002 gnd.n7001 585
R4271 gnd.n7001 gnd.n234 585
R4272 gnd.n7003 gnd.n245 585
R4273 gnd.n7061 gnd.n245 585
R4274 gnd.n7005 gnd.n7004 585
R4275 gnd.n7004 gnd.n244 585
R4276 gnd.n7006 gnd.n252 585
R4277 gnd.n7053 gnd.n252 585
R4278 gnd.n7008 gnd.n7007 585
R4279 gnd.n7007 gnd.n251 585
R4280 gnd.n7009 gnd.n258 585
R4281 gnd.n7045 gnd.n258 585
R4282 gnd.n7013 gnd.n7012 585
R4283 gnd.n7012 gnd.n7011 585
R4284 gnd.n7014 gnd.n290 585
R4285 gnd.n7022 gnd.n290 585
R4286 gnd.n7016 gnd.n7015 585
R4287 gnd.n7017 gnd.n7016 585
R4288 gnd.n6955 gnd.n293 585
R4289 gnd.n6929 gnd.n293 585
R4290 gnd.n6954 gnd.n6953 585
R4291 gnd.n6953 gnd.n6952 585
R4292 gnd.n296 gnd.n294 585
R4293 gnd.n6947 gnd.n296 585
R4294 gnd.n5543 gnd.n5542 585
R4295 gnd.n5542 gnd.n308 585
R4296 gnd.n5544 gnd.n307 585
R4297 gnd.n6939 gnd.n307 585
R4298 gnd.n5545 gnd.n273 585
R4299 gnd.n7038 gnd.n273 585
R4300 gnd.n5547 gnd.n5546 585
R4301 gnd.n5548 gnd.n5547 585
R4302 gnd.n2829 gnd.n2802 585
R4303 gnd.n5587 gnd.n2802 585
R4304 gnd.n5534 gnd.n5533 585
R4305 gnd.n5533 gnd.n2813 585
R4306 gnd.n5532 gnd.n2811 585
R4307 gnd.n5579 gnd.n2811 585
R4308 gnd.n5531 gnd.n2822 585
R4309 gnd.n5560 gnd.n2822 585
R4310 gnd.n2835 gnd.n2831 585
R4311 gnd.n2835 gnd.n2821 585
R4312 gnd.n5527 gnd.n5526 585
R4313 gnd.n5526 gnd.n5525 585
R4314 gnd.n2834 gnd.n2833 585
R4315 gnd.n2847 gnd.n2834 585
R4316 gnd.n2938 gnd.n2845 585
R4317 gnd.n5515 gnd.n2845 585
R4318 gnd.n2939 gnd.n2856 585
R4319 gnd.n5502 gnd.n2856 585
R4320 gnd.n2941 gnd.n2940 585
R4321 gnd.n2940 gnd.n2855 585
R4322 gnd.n2942 gnd.n2864 585
R4323 gnd.n5488 gnd.n2864 585
R4324 gnd.n2944 gnd.n2943 585
R4325 gnd.n2943 gnd.n2876 585
R4326 gnd.n2945 gnd.n2873 585
R4327 gnd.n5478 gnd.n2873 585
R4328 gnd.n2946 gnd.n2884 585
R4329 gnd.n5466 gnd.n2884 585
R4330 gnd.n2948 gnd.n2947 585
R4331 gnd.n2947 gnd.n2883 585
R4332 gnd.n2949 gnd.n2892 585
R4333 gnd.n5457 gnd.n2892 585
R4334 gnd.n2951 gnd.n2950 585
R4335 gnd.n2950 gnd.n2904 585
R4336 gnd.n2952 gnd.n2902 585
R4337 gnd.n5447 gnd.n2902 585
R4338 gnd.n2954 gnd.n2953 585
R4339 gnd.n5435 gnd.n2954 585
R4340 gnd.n2924 gnd.n2770 585
R4341 gnd.n2923 gnd.n2770 585
R4342 gnd.n5623 gnd.n2771 585
R4343 gnd.n5623 gnd.n5622 585
R4344 gnd.n5233 gnd.n5232 585
R4345 gnd.n5232 gnd.n5231 585
R4346 gnd.n5234 gnd.n5032 585
R4347 gnd.n5032 gnd.n3104 585
R4348 gnd.n5236 gnd.n5235 585
R4349 gnd.n5237 gnd.n5236 585
R4350 gnd.n5034 gnd.n5031 585
R4351 gnd.n5031 gnd.n3112 585
R4352 gnd.n5033 gnd.n5022 585
R4353 gnd.n5022 gnd.n3111 585
R4354 gnd.n5245 gnd.n5021 585
R4355 gnd.n5245 gnd.n5244 585
R4356 gnd.n5247 gnd.n5246 585
R4357 gnd.n5246 gnd.n3119 585
R4358 gnd.n5248 gnd.n5018 585
R4359 gnd.n5018 gnd.n3118 585
R4360 gnd.n5250 gnd.n5249 585
R4361 gnd.n5251 gnd.n5250 585
R4362 gnd.n5020 gnd.n5017 585
R4363 gnd.n5017 gnd.n3126 585
R4364 gnd.n5019 gnd.n5010 585
R4365 gnd.n5010 gnd.n3125 585
R4366 gnd.n5261 gnd.n5009 585
R4367 gnd.n5261 gnd.n5260 585
R4368 gnd.n5263 gnd.n5262 585
R4369 gnd.n5262 gnd.n3133 585
R4370 gnd.n5264 gnd.n5006 585
R4371 gnd.n5006 gnd.n3132 585
R4372 gnd.n5266 gnd.n5265 585
R4373 gnd.n5267 gnd.n5266 585
R4374 gnd.n5008 gnd.n5005 585
R4375 gnd.n5005 gnd.n3139 585
R4376 gnd.n5007 gnd.n4994 585
R4377 gnd.n5273 gnd.n4994 585
R4378 gnd.n5276 gnd.n4993 585
R4379 gnd.n5276 gnd.n5275 585
R4380 gnd.n5278 gnd.n5277 585
R4381 gnd.n5277 gnd.n3146 585
R4382 gnd.n5279 gnd.n4990 585
R4383 gnd.n4990 gnd.n3145 585
R4384 gnd.n5281 gnd.n5280 585
R4385 gnd.n5282 gnd.n5281 585
R4386 gnd.n4992 gnd.n4989 585
R4387 gnd.n4989 gnd.n3153 585
R4388 gnd.n4991 gnd.n4981 585
R4389 gnd.n4981 gnd.n3152 585
R4390 gnd.n5291 gnd.n4980 585
R4391 gnd.n5291 gnd.n5290 585
R4392 gnd.n5293 gnd.n5292 585
R4393 gnd.n5292 gnd.n3159 585
R4394 gnd.n5294 gnd.n3184 585
R4395 gnd.n3184 gnd.n3183 585
R4396 gnd.n5296 gnd.n5295 585
R4397 gnd.n5297 gnd.n5296 585
R4398 gnd.n4979 gnd.n3182 585
R4399 gnd.n3182 gnd.n3166 585
R4400 gnd.n4978 gnd.n4977 585
R4401 gnd.n4977 gnd.n3165 585
R4402 gnd.n4976 gnd.n4972 585
R4403 gnd.n4976 gnd.n4975 585
R4404 gnd.n4971 gnd.n3173 585
R4405 gnd.n5305 gnd.n3173 585
R4406 gnd.n4970 gnd.n4969 585
R4407 gnd.n4969 gnd.n3172 585
R4408 gnd.n4968 gnd.n3185 585
R4409 gnd.n4968 gnd.n4967 585
R4410 gnd.n4836 gnd.n3186 585
R4411 gnd.n4846 gnd.n3186 585
R4412 gnd.n4837 gnd.n4835 585
R4413 gnd.n4835 gnd.n3197 585
R4414 gnd.n4839 gnd.n4838 585
R4415 gnd.n4839 gnd.n3195 585
R4416 gnd.n4840 gnd.n4834 585
R4417 gnd.n4854 gnd.n4840 585
R4418 gnd.n4857 gnd.n4856 585
R4419 gnd.n4856 gnd.n4855 585
R4420 gnd.n4858 gnd.n4831 585
R4421 gnd.n4831 gnd.n3204 585
R4422 gnd.n4860 gnd.n4859 585
R4423 gnd.n4861 gnd.n4860 585
R4424 gnd.n4833 gnd.n4830 585
R4425 gnd.n4830 gnd.n3211 585
R4426 gnd.n4832 gnd.n4820 585
R4427 gnd.n4867 gnd.n4820 585
R4428 gnd.n4870 gnd.n4819 585
R4429 gnd.n4870 gnd.n4869 585
R4430 gnd.n4872 gnd.n4871 585
R4431 gnd.n4871 gnd.n3218 585
R4432 gnd.n4873 gnd.n4816 585
R4433 gnd.n4816 gnd.n3217 585
R4434 gnd.n4875 gnd.n4874 585
R4435 gnd.n4876 gnd.n4875 585
R4436 gnd.n4818 gnd.n4815 585
R4437 gnd.n4815 gnd.n3226 585
R4438 gnd.n4817 gnd.n4807 585
R4439 gnd.n4807 gnd.n3224 585
R4440 gnd.n4885 gnd.n4806 585
R4441 gnd.n4885 gnd.n4884 585
R4442 gnd.n4887 gnd.n4886 585
R4443 gnd.n4886 gnd.n3233 585
R4444 gnd.n4888 gnd.n3260 585
R4445 gnd.n3260 gnd.n3232 585
R4446 gnd.n4890 gnd.n4889 585
R4447 gnd.n4891 gnd.n4890 585
R4448 gnd.n4805 gnd.n3259 585
R4449 gnd.n3259 gnd.n3241 585
R4450 gnd.n4804 gnd.n4803 585
R4451 gnd.n4803 gnd.n3239 585
R4452 gnd.n4802 gnd.n4801 585
R4453 gnd.n4802 gnd.n3250 585
R4454 gnd.n4800 gnd.n3248 585
R4455 gnd.n4899 gnd.n3248 585
R4456 gnd.n4799 gnd.n4798 585
R4457 gnd.n4798 gnd.n3247 585
R4458 gnd.n4797 gnd.n3261 585
R4459 gnd.n4797 gnd.n4796 585
R4460 gnd.n4665 gnd.n3262 585
R4461 gnd.n4675 gnd.n3262 585
R4462 gnd.n4666 gnd.n4664 585
R4463 gnd.n4664 gnd.n3273 585
R4464 gnd.n4668 gnd.n4667 585
R4465 gnd.n4668 gnd.n3272 585
R4466 gnd.n4669 gnd.n4663 585
R4467 gnd.n4683 gnd.n4669 585
R4468 gnd.n4686 gnd.n4685 585
R4469 gnd.n4685 gnd.n4684 585
R4470 gnd.n4687 gnd.n4660 585
R4471 gnd.n4660 gnd.n3280 585
R4472 gnd.n4689 gnd.n4688 585
R4473 gnd.n4690 gnd.n4689 585
R4474 gnd.n4662 gnd.n4659 585
R4475 gnd.n4659 gnd.n4656 585
R4476 gnd.n4661 gnd.n4648 585
R4477 gnd.n4696 gnd.n4648 585
R4478 gnd.n4699 gnd.n4647 585
R4479 gnd.n4699 gnd.n4698 585
R4480 gnd.n4701 gnd.n4700 585
R4481 gnd.n4700 gnd.n3292 585
R4482 gnd.n4702 gnd.n4644 585
R4483 gnd.n4644 gnd.n3291 585
R4484 gnd.n4704 gnd.n4703 585
R4485 gnd.n4705 gnd.n4704 585
R4486 gnd.n4646 gnd.n4643 585
R4487 gnd.n4643 gnd.n3298 585
R4488 gnd.n4645 gnd.n4632 585
R4489 gnd.n4711 gnd.n4632 585
R4490 gnd.n4714 gnd.n4631 585
R4491 gnd.n4714 gnd.n4713 585
R4492 gnd.n4716 gnd.n4715 585
R4493 gnd.n4715 gnd.n3305 585
R4494 gnd.n4717 gnd.n3331 585
R4495 gnd.n3331 gnd.n3304 585
R4496 gnd.n4719 gnd.n4718 585
R4497 gnd.n4720 gnd.n4719 585
R4498 gnd.n4630 gnd.n3330 585
R4499 gnd.n3330 gnd.n3312 585
R4500 gnd.n4629 gnd.n4628 585
R4501 gnd.n4628 gnd.n3311 585
R4502 gnd.n4627 gnd.n4626 585
R4503 gnd.n4627 gnd.n3320 585
R4504 gnd.n4625 gnd.n3318 585
R4505 gnd.n4728 gnd.n3318 585
R4506 gnd.n4624 gnd.n4623 585
R4507 gnd.n4623 gnd.n4622 585
R4508 gnd.n3333 gnd.n3332 585
R4509 gnd.n3334 gnd.n3333 585
R4510 gnd.n4501 gnd.n4500 585
R4511 gnd.n4502 gnd.n4501 585
R4512 gnd.n4499 gnd.n4497 585
R4513 gnd.n4497 gnd.n3343 585
R4514 gnd.n4498 gnd.n4489 585
R4515 gnd.n4489 gnd.n3342 585
R4516 gnd.n4511 gnd.n4488 585
R4517 gnd.n4511 gnd.n4510 585
R4518 gnd.n4513 gnd.n4512 585
R4519 gnd.n4512 gnd.n3352 585
R4520 gnd.n4514 gnd.n4485 585
R4521 gnd.n4485 gnd.n3350 585
R4522 gnd.n4516 gnd.n4515 585
R4523 gnd.n4517 gnd.n4516 585
R4524 gnd.n4487 gnd.n4484 585
R4525 gnd.n4484 gnd.n3358 585
R4526 gnd.n4486 gnd.n4474 585
R4527 gnd.n4523 gnd.n4474 585
R4528 gnd.n4526 gnd.n4473 585
R4529 gnd.n4526 gnd.n4525 585
R4530 gnd.n4528 gnd.n4527 585
R4531 gnd.n4527 gnd.n3366 585
R4532 gnd.n4529 gnd.n4470 585
R4533 gnd.n4470 gnd.n3364 585
R4534 gnd.n4531 gnd.n4530 585
R4535 gnd.n4532 gnd.n4531 585
R4536 gnd.n4472 gnd.n4469 585
R4537 gnd.n4469 gnd.n3373 585
R4538 gnd.n4471 gnd.n4461 585
R4539 gnd.n4461 gnd.n3372 585
R4540 gnd.n4541 gnd.n4460 585
R4541 gnd.n4541 gnd.n4540 585
R4542 gnd.n4543 gnd.n4542 585
R4543 gnd.n4542 gnd.n3380 585
R4544 gnd.n4544 gnd.n3407 585
R4545 gnd.n3407 gnd.n3406 585
R4546 gnd.n4546 gnd.n4545 585
R4547 gnd.n4547 gnd.n4546 585
R4548 gnd.n4459 gnd.n3404 585
R4549 gnd.n3404 gnd.n3387 585
R4550 gnd.n4458 gnd.n4457 585
R4551 gnd.n4457 gnd.n3386 585
R4552 gnd.n4456 gnd.n4455 585
R4553 gnd.n4456 gnd.n3396 585
R4554 gnd.n4454 gnd.n3393 585
R4555 gnd.n4555 gnd.n3393 585
R4556 gnd.n4453 gnd.n4452 585
R4557 gnd.n4452 gnd.n4451 585
R4558 gnd.n3409 gnd.n3408 585
R4559 gnd.n3410 gnd.n3409 585
R4560 gnd.n4271 gnd.n4270 585
R4561 gnd.n4272 gnd.n4271 585
R4562 gnd.n4269 gnd.n4163 585
R4563 gnd.n4163 gnd.n3418 585
R4564 gnd.n4268 gnd.n4267 585
R4565 gnd.n4267 gnd.n3417 585
R4566 gnd.n4266 gnd.n4265 585
R4567 gnd.n4264 gnd.n4263 585
R4568 gnd.n4262 gnd.n4186 585
R4569 gnd.n4262 gnd.n3427 585
R4570 gnd.n4261 gnd.n4260 585
R4571 gnd.n4259 gnd.n4258 585
R4572 gnd.n4257 gnd.n4188 585
R4573 gnd.n4255 gnd.n4254 585
R4574 gnd.n4253 gnd.n4189 585
R4575 gnd.n4252 gnd.n4251 585
R4576 gnd.n4249 gnd.n4190 585
R4577 gnd.n4247 gnd.n4246 585
R4578 gnd.n4245 gnd.n4191 585
R4579 gnd.n4244 gnd.n4243 585
R4580 gnd.n4241 gnd.n4192 585
R4581 gnd.n4239 gnd.n4238 585
R4582 gnd.n4237 gnd.n4193 585
R4583 gnd.n4236 gnd.n4235 585
R4584 gnd.n4233 gnd.n4194 585
R4585 gnd.n4231 gnd.n4230 585
R4586 gnd.n4229 gnd.n4195 585
R4587 gnd.n4228 gnd.n4227 585
R4588 gnd.n4225 gnd.n4196 585
R4589 gnd.n4223 gnd.n4222 585
R4590 gnd.n4221 gnd.n4197 585
R4591 gnd.n4220 gnd.n4219 585
R4592 gnd.n4217 gnd.n4198 585
R4593 gnd.n4215 gnd.n4214 585
R4594 gnd.n4213 gnd.n4199 585
R4595 gnd.n4212 gnd.n4211 585
R4596 gnd.n4209 gnd.n4208 585
R4597 gnd.n4207 gnd.n4206 585
R4598 gnd.n4205 gnd.n4142 585
R4599 gnd.n4347 gnd.n4346 585
R4600 gnd.n4344 gnd.n4141 585
R4601 gnd.n4342 gnd.n4341 585
R4602 gnd.n4340 gnd.n4144 585
R4603 gnd.n4338 gnd.n4337 585
R4604 gnd.n4335 gnd.n4147 585
R4605 gnd.n4333 gnd.n4332 585
R4606 gnd.n4331 gnd.n4148 585
R4607 gnd.n4330 gnd.n4329 585
R4608 gnd.n4327 gnd.n4149 585
R4609 gnd.n4325 gnd.n4324 585
R4610 gnd.n4323 gnd.n4150 585
R4611 gnd.n4322 gnd.n4321 585
R4612 gnd.n4319 gnd.n4151 585
R4613 gnd.n4317 gnd.n4316 585
R4614 gnd.n4315 gnd.n4152 585
R4615 gnd.n4314 gnd.n4313 585
R4616 gnd.n4311 gnd.n4153 585
R4617 gnd.n4309 gnd.n4308 585
R4618 gnd.n4307 gnd.n4154 585
R4619 gnd.n4306 gnd.n4305 585
R4620 gnd.n4303 gnd.n4155 585
R4621 gnd.n4301 gnd.n4300 585
R4622 gnd.n4299 gnd.n4156 585
R4623 gnd.n4298 gnd.n4297 585
R4624 gnd.n4295 gnd.n4157 585
R4625 gnd.n4293 gnd.n4292 585
R4626 gnd.n4291 gnd.n4158 585
R4627 gnd.n4290 gnd.n4289 585
R4628 gnd.n4287 gnd.n4159 585
R4629 gnd.n4285 gnd.n4284 585
R4630 gnd.n4283 gnd.n4160 585
R4631 gnd.n4282 gnd.n4281 585
R4632 gnd.n5164 gnd.n5163 585
R4633 gnd.n5166 gnd.n5165 585
R4634 gnd.n5168 gnd.n5167 585
R4635 gnd.n5170 gnd.n5169 585
R4636 gnd.n5172 gnd.n5171 585
R4637 gnd.n5174 gnd.n5173 585
R4638 gnd.n5176 gnd.n5175 585
R4639 gnd.n5178 gnd.n5177 585
R4640 gnd.n5180 gnd.n5179 585
R4641 gnd.n5182 gnd.n5181 585
R4642 gnd.n5184 gnd.n5183 585
R4643 gnd.n5186 gnd.n5185 585
R4644 gnd.n5188 gnd.n5187 585
R4645 gnd.n5190 gnd.n5189 585
R4646 gnd.n5192 gnd.n5191 585
R4647 gnd.n5194 gnd.n5193 585
R4648 gnd.n5196 gnd.n5195 585
R4649 gnd.n5198 gnd.n5197 585
R4650 gnd.n5200 gnd.n5199 585
R4651 gnd.n5202 gnd.n5201 585
R4652 gnd.n5204 gnd.n5203 585
R4653 gnd.n5206 gnd.n5205 585
R4654 gnd.n5208 gnd.n5207 585
R4655 gnd.n5210 gnd.n5209 585
R4656 gnd.n5212 gnd.n5211 585
R4657 gnd.n5214 gnd.n5213 585
R4658 gnd.n5216 gnd.n5215 585
R4659 gnd.n5218 gnd.n5217 585
R4660 gnd.n5220 gnd.n5219 585
R4661 gnd.n5223 gnd.n5222 585
R4662 gnd.n5225 gnd.n5224 585
R4663 gnd.n5227 gnd.n5226 585
R4664 gnd.n5229 gnd.n5228 585
R4665 gnd.n5140 gnd.n2741 585
R4666 gnd.n5139 gnd.n5138 585
R4667 gnd.n5137 gnd.n5136 585
R4668 gnd.n5135 gnd.n5134 585
R4669 gnd.n5132 gnd.n5131 585
R4670 gnd.n5130 gnd.n5129 585
R4671 gnd.n5128 gnd.n5127 585
R4672 gnd.n5126 gnd.n5125 585
R4673 gnd.n5124 gnd.n5123 585
R4674 gnd.n5122 gnd.n5121 585
R4675 gnd.n5120 gnd.n5119 585
R4676 gnd.n5118 gnd.n5117 585
R4677 gnd.n5116 gnd.n5115 585
R4678 gnd.n5114 gnd.n5113 585
R4679 gnd.n5112 gnd.n5111 585
R4680 gnd.n5110 gnd.n5109 585
R4681 gnd.n5108 gnd.n5107 585
R4682 gnd.n5106 gnd.n5105 585
R4683 gnd.n5104 gnd.n5103 585
R4684 gnd.n5102 gnd.n5101 585
R4685 gnd.n5100 gnd.n5099 585
R4686 gnd.n5098 gnd.n5097 585
R4687 gnd.n5096 gnd.n5095 585
R4688 gnd.n5094 gnd.n5093 585
R4689 gnd.n5092 gnd.n5091 585
R4690 gnd.n5090 gnd.n5089 585
R4691 gnd.n5088 gnd.n5087 585
R4692 gnd.n5086 gnd.n5085 585
R4693 gnd.n5084 gnd.n5083 585
R4694 gnd.n5082 gnd.n5081 585
R4695 gnd.n5080 gnd.n5079 585
R4696 gnd.n5078 gnd.n5077 585
R4697 gnd.n5076 gnd.n5055 585
R4698 gnd.n5162 gnd.n5056 585
R4699 gnd.n5231 gnd.n5056 585
R4700 gnd.n5161 gnd.n5029 585
R4701 gnd.n5029 gnd.n3104 585
R4702 gnd.n5238 gnd.n5028 585
R4703 gnd.n5238 gnd.n5237 585
R4704 gnd.n5240 gnd.n5239 585
R4705 gnd.n5239 gnd.n3112 585
R4706 gnd.n5241 gnd.n5025 585
R4707 gnd.n5025 gnd.n3111 585
R4708 gnd.n5243 gnd.n5242 585
R4709 gnd.n5244 gnd.n5243 585
R4710 gnd.n5027 gnd.n5024 585
R4711 gnd.n5024 gnd.n3119 585
R4712 gnd.n5026 gnd.n5015 585
R4713 gnd.n5015 gnd.n3118 585
R4714 gnd.n5252 gnd.n5014 585
R4715 gnd.n5252 gnd.n5251 585
R4716 gnd.n5254 gnd.n5253 585
R4717 gnd.n5253 gnd.n3126 585
R4718 gnd.n5255 gnd.n5012 585
R4719 gnd.n5012 gnd.n3125 585
R4720 gnd.n5257 gnd.n5256 585
R4721 gnd.n5260 gnd.n5257 585
R4722 gnd.n5013 gnd.n5011 585
R4723 gnd.n5011 gnd.n3133 585
R4724 gnd.n5003 gnd.n5002 585
R4725 gnd.n5003 gnd.n3132 585
R4726 gnd.n5269 gnd.n5268 585
R4727 gnd.n5268 gnd.n5267 585
R4728 gnd.n5270 gnd.n4997 585
R4729 gnd.n4997 gnd.n3139 585
R4730 gnd.n5272 gnd.n5271 585
R4731 gnd.n5273 gnd.n5272 585
R4732 gnd.n5001 gnd.n4995 585
R4733 gnd.n5275 gnd.n4995 585
R4734 gnd.n5000 gnd.n4999 585
R4735 gnd.n4999 gnd.n3146 585
R4736 gnd.n4998 gnd.n4987 585
R4737 gnd.n4987 gnd.n3145 585
R4738 gnd.n5283 gnd.n4986 585
R4739 gnd.n5283 gnd.n5282 585
R4740 gnd.n5285 gnd.n5284 585
R4741 gnd.n5284 gnd.n3153 585
R4742 gnd.n5286 gnd.n4983 585
R4743 gnd.n4983 gnd.n3152 585
R4744 gnd.n5288 gnd.n5287 585
R4745 gnd.n5290 gnd.n5288 585
R4746 gnd.n4985 gnd.n4982 585
R4747 gnd.n4982 gnd.n3159 585
R4748 gnd.n4984 gnd.n3179 585
R4749 gnd.n3183 gnd.n3179 585
R4750 gnd.n5298 gnd.n3180 585
R4751 gnd.n5298 gnd.n5297 585
R4752 gnd.n5299 gnd.n3178 585
R4753 gnd.n5299 gnd.n3166 585
R4754 gnd.n5301 gnd.n5300 585
R4755 gnd.n5300 gnd.n3165 585
R4756 gnd.n5302 gnd.n3176 585
R4757 gnd.n4975 gnd.n3176 585
R4758 gnd.n5304 gnd.n5303 585
R4759 gnd.n5305 gnd.n5304 585
R4760 gnd.n3177 gnd.n3175 585
R4761 gnd.n3175 gnd.n3172 585
R4762 gnd.n4844 gnd.n3188 585
R4763 gnd.n4967 gnd.n3188 585
R4764 gnd.n4847 gnd.n4845 585
R4765 gnd.n4847 gnd.n4846 585
R4766 gnd.n4849 gnd.n4848 585
R4767 gnd.n4848 gnd.n3197 585
R4768 gnd.n4850 gnd.n4842 585
R4769 gnd.n4842 gnd.n3195 585
R4770 gnd.n4852 gnd.n4851 585
R4771 gnd.n4854 gnd.n4852 585
R4772 gnd.n4843 gnd.n4841 585
R4773 gnd.n4855 gnd.n4841 585
R4774 gnd.n4828 gnd.n4827 585
R4775 gnd.n4828 gnd.n3204 585
R4776 gnd.n4863 gnd.n4862 585
R4777 gnd.n4862 gnd.n4861 585
R4778 gnd.n4864 gnd.n4822 585
R4779 gnd.n4822 gnd.n3211 585
R4780 gnd.n4866 gnd.n4865 585
R4781 gnd.n4867 gnd.n4866 585
R4782 gnd.n4826 gnd.n4821 585
R4783 gnd.n4869 gnd.n4821 585
R4784 gnd.n4825 gnd.n4824 585
R4785 gnd.n4824 gnd.n3218 585
R4786 gnd.n4823 gnd.n4813 585
R4787 gnd.n4813 gnd.n3217 585
R4788 gnd.n4877 gnd.n4812 585
R4789 gnd.n4877 gnd.n4876 585
R4790 gnd.n4879 gnd.n4878 585
R4791 gnd.n4878 gnd.n3226 585
R4792 gnd.n4880 gnd.n4809 585
R4793 gnd.n4809 gnd.n3224 585
R4794 gnd.n4882 gnd.n4881 585
R4795 gnd.n4884 gnd.n4882 585
R4796 gnd.n4811 gnd.n4808 585
R4797 gnd.n4808 gnd.n3233 585
R4798 gnd.n4810 gnd.n3256 585
R4799 gnd.n3256 gnd.n3232 585
R4800 gnd.n4892 gnd.n3257 585
R4801 gnd.n4892 gnd.n4891 585
R4802 gnd.n4893 gnd.n3255 585
R4803 gnd.n4893 gnd.n3241 585
R4804 gnd.n4895 gnd.n4894 585
R4805 gnd.n4894 gnd.n3239 585
R4806 gnd.n4896 gnd.n3253 585
R4807 gnd.n3253 gnd.n3250 585
R4808 gnd.n4898 gnd.n4897 585
R4809 gnd.n4899 gnd.n4898 585
R4810 gnd.n3254 gnd.n3252 585
R4811 gnd.n3252 gnd.n3247 585
R4812 gnd.n4673 gnd.n3265 585
R4813 gnd.n4796 gnd.n3265 585
R4814 gnd.n4676 gnd.n4674 585
R4815 gnd.n4676 gnd.n4675 585
R4816 gnd.n4678 gnd.n4677 585
R4817 gnd.n4677 gnd.n3273 585
R4818 gnd.n4679 gnd.n4671 585
R4819 gnd.n4671 gnd.n3272 585
R4820 gnd.n4681 gnd.n4680 585
R4821 gnd.n4683 gnd.n4681 585
R4822 gnd.n4672 gnd.n4670 585
R4823 gnd.n4684 gnd.n4670 585
R4824 gnd.n4655 gnd.n4654 585
R4825 gnd.n4655 gnd.n3280 585
R4826 gnd.n4692 gnd.n4691 585
R4827 gnd.n4691 gnd.n4690 585
R4828 gnd.n4693 gnd.n4650 585
R4829 gnd.n4656 gnd.n4650 585
R4830 gnd.n4695 gnd.n4694 585
R4831 gnd.n4696 gnd.n4695 585
R4832 gnd.n4653 gnd.n4649 585
R4833 gnd.n4698 gnd.n4649 585
R4834 gnd.n4652 gnd.n4651 585
R4835 gnd.n4651 gnd.n3292 585
R4836 gnd.n4640 gnd.n4639 585
R4837 gnd.n4640 gnd.n3291 585
R4838 gnd.n4707 gnd.n4706 585
R4839 gnd.n4706 gnd.n4705 585
R4840 gnd.n4708 gnd.n4634 585
R4841 gnd.n4634 gnd.n3298 585
R4842 gnd.n4710 gnd.n4709 585
R4843 gnd.n4711 gnd.n4710 585
R4844 gnd.n4638 gnd.n4633 585
R4845 gnd.n4713 gnd.n4633 585
R4846 gnd.n4637 gnd.n4636 585
R4847 gnd.n4636 gnd.n3305 585
R4848 gnd.n4635 gnd.n3326 585
R4849 gnd.n3326 gnd.n3304 585
R4850 gnd.n4721 gnd.n3327 585
R4851 gnd.n4721 gnd.n4720 585
R4852 gnd.n4722 gnd.n3325 585
R4853 gnd.n4722 gnd.n3312 585
R4854 gnd.n4724 gnd.n4723 585
R4855 gnd.n4723 gnd.n3311 585
R4856 gnd.n4725 gnd.n3323 585
R4857 gnd.n3323 gnd.n3320 585
R4858 gnd.n4727 gnd.n4726 585
R4859 gnd.n4728 gnd.n4727 585
R4860 gnd.n3324 gnd.n3322 585
R4861 gnd.n4622 gnd.n3322 585
R4862 gnd.n4495 gnd.n4494 585
R4863 gnd.n4495 gnd.n3334 585
R4864 gnd.n4503 gnd.n4493 585
R4865 gnd.n4503 gnd.n4502 585
R4866 gnd.n4505 gnd.n4504 585
R4867 gnd.n4504 gnd.n3343 585
R4868 gnd.n4506 gnd.n4491 585
R4869 gnd.n4491 gnd.n3342 585
R4870 gnd.n4508 gnd.n4507 585
R4871 gnd.n4510 gnd.n4508 585
R4872 gnd.n4492 gnd.n4490 585
R4873 gnd.n4490 gnd.n3352 585
R4874 gnd.n4482 gnd.n4481 585
R4875 gnd.n4482 gnd.n3350 585
R4876 gnd.n4519 gnd.n4518 585
R4877 gnd.n4518 gnd.n4517 585
R4878 gnd.n4520 gnd.n4476 585
R4879 gnd.n4476 gnd.n3358 585
R4880 gnd.n4522 gnd.n4521 585
R4881 gnd.n4523 gnd.n4522 585
R4882 gnd.n4480 gnd.n4475 585
R4883 gnd.n4525 gnd.n4475 585
R4884 gnd.n4479 gnd.n4478 585
R4885 gnd.n4478 gnd.n3366 585
R4886 gnd.n4477 gnd.n4467 585
R4887 gnd.n4467 gnd.n3364 585
R4888 gnd.n4533 gnd.n4466 585
R4889 gnd.n4533 gnd.n4532 585
R4890 gnd.n4535 gnd.n4534 585
R4891 gnd.n4534 gnd.n3373 585
R4892 gnd.n4536 gnd.n4463 585
R4893 gnd.n4463 gnd.n3372 585
R4894 gnd.n4538 gnd.n4537 585
R4895 gnd.n4540 gnd.n4538 585
R4896 gnd.n4465 gnd.n4462 585
R4897 gnd.n4462 gnd.n3380 585
R4898 gnd.n4464 gnd.n3402 585
R4899 gnd.n3406 gnd.n3402 585
R4900 gnd.n4548 gnd.n3403 585
R4901 gnd.n4548 gnd.n4547 585
R4902 gnd.n4549 gnd.n3401 585
R4903 gnd.n4549 gnd.n3387 585
R4904 gnd.n4551 gnd.n4550 585
R4905 gnd.n4550 gnd.n3386 585
R4906 gnd.n4552 gnd.n3399 585
R4907 gnd.n3399 gnd.n3396 585
R4908 gnd.n4554 gnd.n4553 585
R4909 gnd.n4555 gnd.n4554 585
R4910 gnd.n3400 gnd.n3398 585
R4911 gnd.n4451 gnd.n3398 585
R4912 gnd.n4275 gnd.n4274 585
R4913 gnd.n4274 gnd.n3410 585
R4914 gnd.n4276 gnd.n4273 585
R4915 gnd.n4273 gnd.n4272 585
R4916 gnd.n4278 gnd.n4277 585
R4917 gnd.n4278 gnd.n3418 585
R4918 gnd.n4279 gnd.n4161 585
R4919 gnd.n4279 gnd.n3417 585
R4920 gnd.n3687 gnd.n3686 585
R4921 gnd.n3687 gnd.n2408 585
R4922 gnd.n6923 gnd.n6922 585
R4923 gnd.n6923 gnd.n259 585
R4924 gnd.n6925 gnd.n6924 585
R4925 gnd.n6924 gnd.n291 585
R4926 gnd.n6926 gnd.n317 585
R4927 gnd.n317 gnd.n289 585
R4928 gnd.n6931 gnd.n6927 585
R4929 gnd.n6931 gnd.n6930 585
R4930 gnd.n6932 gnd.n316 585
R4931 gnd.n6932 gnd.n299 585
R4932 gnd.n6934 gnd.n6933 585
R4933 gnd.n6933 gnd.n297 585
R4934 gnd.n6935 gnd.n310 585
R4935 gnd.n310 gnd.n302 585
R4936 gnd.n6937 gnd.n6936 585
R4937 gnd.n6938 gnd.n6937 585
R4938 gnd.n311 gnd.n309 585
R4939 gnd.n309 gnd.n275 585
R4940 gnd.n5572 gnd.n5571 585
R4941 gnd.n5572 gnd.n272 585
R4942 gnd.n5574 gnd.n5573 585
R4943 gnd.n5573 gnd.n2804 585
R4944 gnd.n5575 gnd.n2816 585
R4945 gnd.n2816 gnd.n2815 585
R4946 gnd.n5577 gnd.n5576 585
R4947 gnd.n5578 gnd.n5577 585
R4948 gnd.n2817 gnd.n2814 585
R4949 gnd.n2814 gnd.n2810 585
R4950 gnd.n5563 gnd.n5562 585
R4951 gnd.n5562 gnd.n5561 585
R4952 gnd.n2820 gnd.n2819 585
R4953 gnd.n2837 gnd.n2820 585
R4954 gnd.n5510 gnd.n2850 585
R4955 gnd.n2850 gnd.n2849 585
R4956 gnd.n5512 gnd.n5511 585
R4957 gnd.n5513 gnd.n5512 585
R4958 gnd.n2851 gnd.n2848 585
R4959 gnd.n2848 gnd.n2844 585
R4960 gnd.n5505 gnd.n5504 585
R4961 gnd.n5504 gnd.n5503 585
R4962 gnd.n2854 gnd.n2853 585
R4963 gnd.n2865 gnd.n2854 585
R4964 gnd.n5474 gnd.n2878 585
R4965 gnd.n2878 gnd.n2863 585
R4966 gnd.n5476 gnd.n5475 585
R4967 gnd.n5477 gnd.n5476 585
R4968 gnd.n2879 gnd.n2877 585
R4969 gnd.n2877 gnd.n2872 585
R4970 gnd.n5469 gnd.n5468 585
R4971 gnd.n5468 gnd.n5467 585
R4972 gnd.n2882 gnd.n2881 585
R4973 gnd.n2893 gnd.n2882 585
R4974 gnd.n5443 gnd.n2906 585
R4975 gnd.n2906 gnd.n2891 585
R4976 gnd.n5445 gnd.n5444 585
R4977 gnd.n5446 gnd.n5445 585
R4978 gnd.n2907 gnd.n2905 585
R4979 gnd.n2905 gnd.n2901 585
R4980 gnd.n5438 gnd.n5437 585
R4981 gnd.n5437 gnd.n5436 585
R4982 gnd.n2917 gnd.n2909 585
R4983 gnd.n2917 gnd.n2774 585
R4984 gnd.n2916 gnd.n2915 585
R4985 gnd.n2916 gnd.n2772 585
R4986 gnd.n2911 gnd.n2910 585
R4987 gnd.n2910 gnd.n2721 585
R4988 gnd.n2692 gnd.n2691 585
R4989 gnd.n5699 gnd.n2692 585
R4990 gnd.n5702 gnd.n5701 585
R4991 gnd.n5701 gnd.n5700 585
R4992 gnd.n5703 gnd.n2686 585
R4993 gnd.n2686 gnd.n2685 585
R4994 gnd.n5705 gnd.n5704 585
R4995 gnd.n5706 gnd.n5705 585
R4996 gnd.n2687 gnd.n2683 585
R4997 gnd.n5707 gnd.n2683 585
R4998 gnd.n5395 gnd.n3099 585
R4999 gnd.n3099 gnd.n2682 585
R5000 gnd.n5397 gnd.n5396 585
R5001 gnd.n5398 gnd.n5397 585
R5002 gnd.n3100 gnd.n3098 585
R5003 gnd.n5230 gnd.n3098 585
R5004 gnd.n5389 gnd.n5388 585
R5005 gnd.n5388 gnd.n5387 585
R5006 gnd.n3103 gnd.n3102 585
R5007 gnd.n5030 gnd.n3103 585
R5008 gnd.n5376 gnd.n5375 585
R5009 gnd.n5377 gnd.n5376 585
R5010 gnd.n3114 gnd.n3113 585
R5011 gnd.n5244 gnd.n3113 585
R5012 gnd.n5371 gnd.n5370 585
R5013 gnd.n5370 gnd.n5369 585
R5014 gnd.n3117 gnd.n3116 585
R5015 gnd.n5016 gnd.n3117 585
R5016 gnd.n5360 gnd.n5359 585
R5017 gnd.n5361 gnd.n5360 585
R5018 gnd.n3128 gnd.n3127 585
R5019 gnd.n5259 gnd.n3127 585
R5020 gnd.n5355 gnd.n5354 585
R5021 gnd.n5354 gnd.n5353 585
R5022 gnd.n3131 gnd.n3130 585
R5023 gnd.n5004 gnd.n3131 585
R5024 gnd.n5344 gnd.n5343 585
R5025 gnd.n5345 gnd.n5344 585
R5026 gnd.n3141 gnd.n3140 585
R5027 gnd.n5274 gnd.n3140 585
R5028 gnd.n5339 gnd.n5338 585
R5029 gnd.n5338 gnd.n5337 585
R5030 gnd.n3144 gnd.n3143 585
R5031 gnd.n4988 gnd.n3144 585
R5032 gnd.n5328 gnd.n5327 585
R5033 gnd.n5329 gnd.n5328 585
R5034 gnd.n3155 gnd.n3154 585
R5035 gnd.t298 gnd.n3154 585
R5036 gnd.n5323 gnd.n5322 585
R5037 gnd.n5322 gnd.n5321 585
R5038 gnd.n3158 gnd.n3157 585
R5039 gnd.n3181 gnd.n3158 585
R5040 gnd.n5312 gnd.n5311 585
R5041 gnd.n5313 gnd.n5312 585
R5042 gnd.n3168 gnd.n3167 585
R5043 gnd.n4974 gnd.n3167 585
R5044 gnd.n5307 gnd.n5306 585
R5045 gnd.n5306 gnd.n5305 585
R5046 gnd.n3171 gnd.n3170 585
R5047 gnd.n4966 gnd.n3171 585
R5048 gnd.n4954 gnd.n3199 585
R5049 gnd.n3199 gnd.n3187 585
R5050 gnd.n4956 gnd.n4955 585
R5051 gnd.n4957 gnd.n4956 585
R5052 gnd.n3200 gnd.n3198 585
R5053 gnd.n4853 gnd.n3198 585
R5054 gnd.n4949 gnd.n4948 585
R5055 gnd.n4948 gnd.n4947 585
R5056 gnd.n3203 gnd.n3202 585
R5057 gnd.n4829 gnd.n3203 585
R5058 gnd.n4938 gnd.n4937 585
R5059 gnd.n4939 gnd.n4938 585
R5060 gnd.n3213 gnd.n3212 585
R5061 gnd.n4868 gnd.n3212 585
R5062 gnd.n4933 gnd.n4932 585
R5063 gnd.n4932 gnd.n4931 585
R5064 gnd.n3216 gnd.n3215 585
R5065 gnd.n4814 gnd.n3216 585
R5066 gnd.n4922 gnd.n4921 585
R5067 gnd.n4923 gnd.n4922 585
R5068 gnd.n3228 gnd.n3227 585
R5069 gnd.n4883 gnd.n3227 585
R5070 gnd.n4917 gnd.n4916 585
R5071 gnd.n4916 gnd.n4915 585
R5072 gnd.n3231 gnd.n3230 585
R5073 gnd.n3258 gnd.n3231 585
R5074 gnd.n4906 gnd.n4905 585
R5075 gnd.n4907 gnd.n4906 585
R5076 gnd.n3243 gnd.n3242 585
R5077 gnd.n3249 gnd.n3242 585
R5078 gnd.n4901 gnd.n4900 585
R5079 gnd.n4900 gnd.n4899 585
R5080 gnd.n3246 gnd.n3245 585
R5081 gnd.n4795 gnd.n3246 585
R5082 gnd.n4783 gnd.n3275 585
R5083 gnd.n3275 gnd.n3264 585
R5084 gnd.n4785 gnd.n4784 585
R5085 gnd.n4786 gnd.n4785 585
R5086 gnd.n3276 gnd.n3274 585
R5087 gnd.n4682 gnd.n3274 585
R5088 gnd.n4778 gnd.n4777 585
R5089 gnd.n4777 gnd.n4776 585
R5090 gnd.n3279 gnd.n3278 585
R5091 gnd.n4658 gnd.n3279 585
R5092 gnd.n4767 gnd.n4766 585
R5093 gnd.n4768 gnd.n4767 585
R5094 gnd.n3287 gnd.n3286 585
R5095 gnd.n4697 gnd.n3286 585
R5096 gnd.n4762 gnd.n4761 585
R5097 gnd.n4761 gnd.n4760 585
R5098 gnd.n3290 gnd.n3289 585
R5099 gnd.n4642 gnd.n3290 585
R5100 gnd.n4751 gnd.n4750 585
R5101 gnd.n4752 gnd.n4751 585
R5102 gnd.n3300 gnd.n3299 585
R5103 gnd.n4712 gnd.n3299 585
R5104 gnd.n4746 gnd.n4745 585
R5105 gnd.n4745 gnd.n4744 585
R5106 gnd.n3303 gnd.n3302 585
R5107 gnd.n3329 gnd.n3303 585
R5108 gnd.n4735 gnd.n4734 585
R5109 gnd.n4736 gnd.n4735 585
R5110 gnd.n3314 gnd.n3313 585
R5111 gnd.n3319 gnd.n3313 585
R5112 gnd.n4730 gnd.n4729 585
R5113 gnd.n4729 gnd.n4728 585
R5114 gnd.n3317 gnd.n3316 585
R5115 gnd.n4621 gnd.n3317 585
R5116 gnd.n4609 gnd.n3345 585
R5117 gnd.n4496 gnd.n3345 585
R5118 gnd.n4611 gnd.n4610 585
R5119 gnd.n4612 gnd.n4611 585
R5120 gnd.n3346 gnd.n3344 585
R5121 gnd.n4509 gnd.n3344 585
R5122 gnd.n4604 gnd.n4603 585
R5123 gnd.n4603 gnd.t6 585
R5124 gnd.n3349 gnd.n3348 585
R5125 gnd.n4483 gnd.n3349 585
R5126 gnd.n4594 gnd.n4593 585
R5127 gnd.n4595 gnd.n4594 585
R5128 gnd.n3360 gnd.n3359 585
R5129 gnd.n4524 gnd.n3359 585
R5130 gnd.n4589 gnd.n4588 585
R5131 gnd.n4588 gnd.n4587 585
R5132 gnd.n3363 gnd.n3362 585
R5133 gnd.n4468 gnd.n3363 585
R5134 gnd.n4578 gnd.n4577 585
R5135 gnd.n4579 gnd.n4578 585
R5136 gnd.n3375 gnd.n3374 585
R5137 gnd.n4539 gnd.n3374 585
R5138 gnd.n4573 gnd.n4572 585
R5139 gnd.n4572 gnd.n4571 585
R5140 gnd.n3378 gnd.n3377 585
R5141 gnd.n3405 gnd.n3378 585
R5142 gnd.n4562 gnd.n4561 585
R5143 gnd.n4563 gnd.n4562 585
R5144 gnd.n3389 gnd.n3388 585
R5145 gnd.n3395 gnd.n3388 585
R5146 gnd.n4557 gnd.n4556 585
R5147 gnd.n4556 gnd.n4555 585
R5148 gnd.n3392 gnd.n3391 585
R5149 gnd.n4450 gnd.n3392 585
R5150 gnd.n4438 gnd.n3420 585
R5151 gnd.n4162 gnd.n3420 585
R5152 gnd.n4440 gnd.n4439 585
R5153 gnd.n4441 gnd.n4440 585
R5154 gnd.n3421 gnd.n3419 585
R5155 gnd.n3426 gnd.n3419 585
R5156 gnd.n4433 gnd.n4432 585
R5157 gnd.n4432 gnd.n4431 585
R5158 gnd.n3424 gnd.n3423 585
R5159 gnd.n3433 gnd.n3424 585
R5160 gnd.n4422 gnd.n4421 585
R5161 gnd.n4423 gnd.n4422 585
R5162 gnd.n3435 gnd.n3434 585
R5163 gnd.n3434 gnd.n3432 585
R5164 gnd.n4417 gnd.n4416 585
R5165 gnd.n4416 gnd.n4415 585
R5166 gnd.n3438 gnd.n3437 585
R5167 gnd.n3439 gnd.n3438 585
R5168 gnd.n3739 gnd.n3738 585
R5169 gnd.n3738 gnd.n3572 585
R5170 gnd.n3740 gnd.n3733 585
R5171 gnd.n3733 gnd.n3472 585
R5172 gnd.n3742 gnd.n3741 585
R5173 gnd.n3742 gnd.n2572 585
R5174 gnd.n3743 gnd.n3732 585
R5175 gnd.n3743 gnd.n2569 585
R5176 gnd.n3745 gnd.n3744 585
R5177 gnd.n3744 gnd.n3638 585
R5178 gnd.n3746 gnd.n3727 585
R5179 gnd.n3727 gnd.n2560 585
R5180 gnd.n3748 gnd.n3747 585
R5181 gnd.n3748 gnd.n2552 585
R5182 gnd.n3749 gnd.n3726 585
R5183 gnd.n3749 gnd.n2549 585
R5184 gnd.n3751 gnd.n3750 585
R5185 gnd.n3750 gnd.n2541 585
R5186 gnd.n3752 gnd.n3721 585
R5187 gnd.n3721 gnd.n2538 585
R5188 gnd.n3754 gnd.n3753 585
R5189 gnd.n3754 gnd.n2530 585
R5190 gnd.n3755 gnd.n3720 585
R5191 gnd.n3755 gnd.n2527 585
R5192 gnd.n3757 gnd.n3756 585
R5193 gnd.n3756 gnd.n2519 585
R5194 gnd.n3758 gnd.n3715 585
R5195 gnd.n3715 gnd.n2516 585
R5196 gnd.n3760 gnd.n3759 585
R5197 gnd.n3760 gnd.n3655 585
R5198 gnd.n3761 gnd.n3714 585
R5199 gnd.n3761 gnd.n2506 585
R5200 gnd.n3763 gnd.n3762 585
R5201 gnd.n3762 gnd.n2498 585
R5202 gnd.n3764 gnd.n3709 585
R5203 gnd.n3709 gnd.n2495 585
R5204 gnd.n3766 gnd.n3765 585
R5205 gnd.n3766 gnd.n2487 585
R5206 gnd.n3767 gnd.n3708 585
R5207 gnd.n3767 gnd.n2484 585
R5208 gnd.n3769 gnd.n3768 585
R5209 gnd.n3768 gnd.n2476 585
R5210 gnd.n3770 gnd.n3703 585
R5211 gnd.n3703 gnd.n2473 585
R5212 gnd.n3772 gnd.n3771 585
R5213 gnd.n3772 gnd.n3668 585
R5214 gnd.n3773 gnd.n3702 585
R5215 gnd.n3773 gnd.n2463 585
R5216 gnd.n3775 gnd.n3774 585
R5217 gnd.n3774 gnd.n2456 585
R5218 gnd.n3776 gnd.n3697 585
R5219 gnd.n3697 gnd.n2453 585
R5220 gnd.n3778 gnd.n3777 585
R5221 gnd.n3778 gnd.n2445 585
R5222 gnd.n3779 gnd.n3696 585
R5223 gnd.n3779 gnd.n2442 585
R5224 gnd.n3781 gnd.n3780 585
R5225 gnd.n3780 gnd.n2437 585
R5226 gnd.n3782 gnd.n3682 585
R5227 gnd.n3682 gnd.n2434 585
R5228 gnd.n3784 gnd.n3783 585
R5229 gnd.n3785 gnd.n3784 585
R5230 gnd.n3683 gnd.n3681 585
R5231 gnd.n3681 gnd.n2424 585
R5232 gnd.n3689 gnd.n3688 585
R5233 gnd.n3688 gnd.n2418 585
R5234 gnd.n5709 gnd.n5708 585
R5235 gnd.n5708 gnd.n5707 585
R5236 gnd.n5710 gnd.n2679 585
R5237 gnd.n2682 gnd.n2679 585
R5238 gnd.n5711 gnd.n2678 585
R5239 gnd.n5398 gnd.n2678 585
R5240 gnd.n5057 gnd.n2676 585
R5241 gnd.n5230 gnd.n5057 585
R5242 gnd.n5715 gnd.n2675 585
R5243 gnd.n5387 gnd.n2675 585
R5244 gnd.n5716 gnd.n2674 585
R5245 gnd.n5030 gnd.n2674 585
R5246 gnd.n5717 gnd.n2673 585
R5247 gnd.n5377 gnd.n2673 585
R5248 gnd.n5023 gnd.n2671 585
R5249 gnd.n5244 gnd.n5023 585
R5250 gnd.n5721 gnd.n2670 585
R5251 gnd.n5369 gnd.n2670 585
R5252 gnd.n5722 gnd.n2669 585
R5253 gnd.n5016 gnd.n2669 585
R5254 gnd.n5723 gnd.n2668 585
R5255 gnd.n5361 gnd.n2668 585
R5256 gnd.n5258 gnd.n2666 585
R5257 gnd.n5259 gnd.n5258 585
R5258 gnd.n5727 gnd.n2665 585
R5259 gnd.n5353 gnd.n2665 585
R5260 gnd.n5728 gnd.n2664 585
R5261 gnd.n5004 gnd.n2664 585
R5262 gnd.n5729 gnd.n2663 585
R5263 gnd.n5345 gnd.n2663 585
R5264 gnd.n4996 gnd.n2661 585
R5265 gnd.n5274 gnd.n4996 585
R5266 gnd.n5733 gnd.n2660 585
R5267 gnd.n5337 gnd.n2660 585
R5268 gnd.n5734 gnd.n2659 585
R5269 gnd.n4988 gnd.n2659 585
R5270 gnd.n5735 gnd.n2658 585
R5271 gnd.n5329 gnd.n2658 585
R5272 gnd.n5289 gnd.n2656 585
R5273 gnd.t298 gnd.n5289 585
R5274 gnd.n5739 gnd.n2655 585
R5275 gnd.n5321 gnd.n2655 585
R5276 gnd.n5740 gnd.n2654 585
R5277 gnd.n3181 gnd.n2654 585
R5278 gnd.n5741 gnd.n2653 585
R5279 gnd.n5313 gnd.n2653 585
R5280 gnd.n4973 gnd.n2651 585
R5281 gnd.n4974 gnd.n4973 585
R5282 gnd.n5745 gnd.n2650 585
R5283 gnd.n5305 gnd.n2650 585
R5284 gnd.n5746 gnd.n2649 585
R5285 gnd.n4966 gnd.n2649 585
R5286 gnd.n5747 gnd.n2648 585
R5287 gnd.n3187 gnd.n2648 585
R5288 gnd.n3196 gnd.n2646 585
R5289 gnd.n4957 gnd.n3196 585
R5290 gnd.n5751 gnd.n2645 585
R5291 gnd.n4853 gnd.n2645 585
R5292 gnd.n5752 gnd.n2644 585
R5293 gnd.n4947 gnd.n2644 585
R5294 gnd.n5753 gnd.n2643 585
R5295 gnd.n4829 gnd.n2643 585
R5296 gnd.n3210 gnd.n2641 585
R5297 gnd.n4939 gnd.n3210 585
R5298 gnd.n5757 gnd.n2640 585
R5299 gnd.n4868 gnd.n2640 585
R5300 gnd.n5758 gnd.n2639 585
R5301 gnd.n4931 gnd.n2639 585
R5302 gnd.n5759 gnd.n2638 585
R5303 gnd.n4814 gnd.n2638 585
R5304 gnd.n3225 gnd.n2636 585
R5305 gnd.n4923 gnd.n3225 585
R5306 gnd.n5763 gnd.n2635 585
R5307 gnd.n4883 gnd.n2635 585
R5308 gnd.n5764 gnd.n2634 585
R5309 gnd.n4915 gnd.n2634 585
R5310 gnd.n5765 gnd.n2633 585
R5311 gnd.n3258 gnd.n2633 585
R5312 gnd.n3240 gnd.n2631 585
R5313 gnd.n4907 gnd.n3240 585
R5314 gnd.n5769 gnd.n2630 585
R5315 gnd.n3249 gnd.n2630 585
R5316 gnd.n5770 gnd.n2629 585
R5317 gnd.n4899 gnd.n2629 585
R5318 gnd.n5771 gnd.n2628 585
R5319 gnd.n4795 gnd.n2628 585
R5320 gnd.n3263 gnd.n2626 585
R5321 gnd.n3264 gnd.n3263 585
R5322 gnd.n5775 gnd.n2625 585
R5323 gnd.n4786 gnd.n2625 585
R5324 gnd.n5776 gnd.n2624 585
R5325 gnd.n4682 gnd.n2624 585
R5326 gnd.n5777 gnd.n2623 585
R5327 gnd.n4776 gnd.n2623 585
R5328 gnd.n4657 gnd.n2621 585
R5329 gnd.n4658 gnd.n4657 585
R5330 gnd.n5781 gnd.n2620 585
R5331 gnd.n4768 gnd.n2620 585
R5332 gnd.n5782 gnd.n2619 585
R5333 gnd.n4697 gnd.n2619 585
R5334 gnd.n5783 gnd.n2618 585
R5335 gnd.n4760 gnd.n2618 585
R5336 gnd.n4641 gnd.n2616 585
R5337 gnd.n4642 gnd.n4641 585
R5338 gnd.n5787 gnd.n2615 585
R5339 gnd.n4752 gnd.n2615 585
R5340 gnd.n5788 gnd.n2614 585
R5341 gnd.n4712 gnd.n2614 585
R5342 gnd.n5789 gnd.n2613 585
R5343 gnd.n4744 gnd.n2613 585
R5344 gnd.n3328 gnd.n2611 585
R5345 gnd.n3329 gnd.n3328 585
R5346 gnd.n5793 gnd.n2610 585
R5347 gnd.n4736 gnd.n2610 585
R5348 gnd.n5794 gnd.n2609 585
R5349 gnd.n3319 gnd.n2609 585
R5350 gnd.n5795 gnd.n2608 585
R5351 gnd.n4728 gnd.n2608 585
R5352 gnd.n3335 gnd.n2606 585
R5353 gnd.n4621 gnd.n3335 585
R5354 gnd.n5799 gnd.n2605 585
R5355 gnd.n4496 gnd.n2605 585
R5356 gnd.n5800 gnd.n2604 585
R5357 gnd.n4612 gnd.n2604 585
R5358 gnd.n5801 gnd.n2603 585
R5359 gnd.n4509 gnd.n2603 585
R5360 gnd.n3351 gnd.n2601 585
R5361 gnd.t6 gnd.n3351 585
R5362 gnd.n5805 gnd.n2600 585
R5363 gnd.n4483 gnd.n2600 585
R5364 gnd.n5806 gnd.n2599 585
R5365 gnd.n4595 gnd.n2599 585
R5366 gnd.n5807 gnd.n2598 585
R5367 gnd.n4524 gnd.n2598 585
R5368 gnd.n3365 gnd.n2596 585
R5369 gnd.n4587 gnd.n3365 585
R5370 gnd.n5811 gnd.n2595 585
R5371 gnd.n4468 gnd.n2595 585
R5372 gnd.n5812 gnd.n2594 585
R5373 gnd.n4579 gnd.n2594 585
R5374 gnd.n5813 gnd.n2593 585
R5375 gnd.n4539 gnd.n2593 585
R5376 gnd.n3379 gnd.n2591 585
R5377 gnd.n4571 gnd.n3379 585
R5378 gnd.n5817 gnd.n2590 585
R5379 gnd.n3405 gnd.n2590 585
R5380 gnd.n5818 gnd.n2589 585
R5381 gnd.n4563 gnd.n2589 585
R5382 gnd.n5819 gnd.n2588 585
R5383 gnd.n3395 gnd.n2588 585
R5384 gnd.n3394 gnd.n2586 585
R5385 gnd.n4555 gnd.n3394 585
R5386 gnd.n5823 gnd.n2585 585
R5387 gnd.n4450 gnd.n2585 585
R5388 gnd.n5824 gnd.n2584 585
R5389 gnd.n4162 gnd.n2584 585
R5390 gnd.n5825 gnd.n2583 585
R5391 gnd.n4441 gnd.n2583 585
R5392 gnd.n3425 gnd.n2581 585
R5393 gnd.n3426 gnd.n3425 585
R5394 gnd.n5829 gnd.n2580 585
R5395 gnd.n4431 gnd.n2580 585
R5396 gnd.n5830 gnd.n2579 585
R5397 gnd.n3433 gnd.n2579 585
R5398 gnd.n5831 gnd.n2578 585
R5399 gnd.n4423 gnd.n2578 585
R5400 gnd.n3512 gnd.n3511 585
R5401 gnd.n3515 gnd.n3514 585
R5402 gnd.n3513 gnd.n3502 585
R5403 gnd.n3525 gnd.n3524 585
R5404 gnd.n3527 gnd.n3526 585
R5405 gnd.n3497 gnd.n3496 585
R5406 gnd.n3536 gnd.n3498 585
R5407 gnd.n3539 gnd.n3538 585
R5408 gnd.n3537 gnd.n3490 585
R5409 gnd.n3549 gnd.n3548 585
R5410 gnd.n3551 gnd.n3550 585
R5411 gnd.n3485 gnd.n3484 585
R5412 gnd.n3561 gnd.n3486 585
R5413 gnd.n3563 gnd.n3562 585
R5414 gnd.n3565 gnd.n3564 585
R5415 gnd.n3465 gnd.n3464 585
R5416 gnd.n4384 gnd.n3466 585
R5417 gnd.n4387 gnd.n4386 585
R5418 gnd.n4385 gnd.n3461 585
R5419 gnd.n4393 gnd.n4392 585
R5420 gnd.n4395 gnd.n4394 585
R5421 gnd.n4398 gnd.n4397 585
R5422 gnd.n4396 gnd.n3459 585
R5423 gnd.n4403 gnd.n4402 585
R5424 gnd.n4405 gnd.n4404 585
R5425 gnd.n4408 gnd.n4407 585
R5426 gnd.n3454 gnd.n3453 585
R5427 gnd.n4413 gnd.n4412 585
R5428 gnd.n3455 gnd.n3431 585
R5429 gnd.n4415 gnd.n3431 585
R5430 gnd.n5402 gnd.n2684 585
R5431 gnd.n5707 gnd.n2684 585
R5432 gnd.n5401 gnd.n5400 585
R5433 gnd.n5400 gnd.n2682 585
R5434 gnd.n5399 gnd.n3096 585
R5435 gnd.n5399 gnd.n5398 585
R5436 gnd.n3107 gnd.n3097 585
R5437 gnd.n5230 gnd.n3097 585
R5438 gnd.n5386 gnd.n5385 585
R5439 gnd.n5387 gnd.n5386 585
R5440 gnd.n3106 gnd.n3105 585
R5441 gnd.n5030 gnd.n3105 585
R5442 gnd.n5379 gnd.n5378 585
R5443 gnd.n5378 gnd.n5377 585
R5444 gnd.n3110 gnd.n3109 585
R5445 gnd.n5244 gnd.n3110 585
R5446 gnd.n5368 gnd.n5367 585
R5447 gnd.n5369 gnd.n5368 585
R5448 gnd.n3121 gnd.n3120 585
R5449 gnd.n5016 gnd.n3120 585
R5450 gnd.n5363 gnd.n5362 585
R5451 gnd.n5362 gnd.n5361 585
R5452 gnd.n3124 gnd.n3123 585
R5453 gnd.n5259 gnd.n3124 585
R5454 gnd.n5352 gnd.n5351 585
R5455 gnd.n5353 gnd.n5352 585
R5456 gnd.n3135 gnd.n3134 585
R5457 gnd.n5004 gnd.n3134 585
R5458 gnd.n5347 gnd.n5346 585
R5459 gnd.n5346 gnd.n5345 585
R5460 gnd.n3138 gnd.n3137 585
R5461 gnd.n5274 gnd.n3138 585
R5462 gnd.n5336 gnd.n5335 585
R5463 gnd.n5337 gnd.n5336 585
R5464 gnd.n3148 gnd.n3147 585
R5465 gnd.n4988 gnd.n3147 585
R5466 gnd.n5331 gnd.n5330 585
R5467 gnd.n5330 gnd.n5329 585
R5468 gnd.n3151 gnd.n3150 585
R5469 gnd.t298 gnd.n3151 585
R5470 gnd.n5320 gnd.n5319 585
R5471 gnd.n5321 gnd.n5320 585
R5472 gnd.n3161 gnd.n3160 585
R5473 gnd.n3181 gnd.n3160 585
R5474 gnd.n5315 gnd.n5314 585
R5475 gnd.n5314 gnd.n5313 585
R5476 gnd.n3164 gnd.n3163 585
R5477 gnd.n4974 gnd.n3164 585
R5478 gnd.n3191 gnd.n3174 585
R5479 gnd.n5305 gnd.n3174 585
R5480 gnd.n4965 gnd.n4964 585
R5481 gnd.n4966 gnd.n4965 585
R5482 gnd.n3190 gnd.n3189 585
R5483 gnd.n3189 gnd.n3187 585
R5484 gnd.n4959 gnd.n4958 585
R5485 gnd.n4958 gnd.n4957 585
R5486 gnd.n3194 gnd.n3193 585
R5487 gnd.n4853 gnd.n3194 585
R5488 gnd.n4946 gnd.n4945 585
R5489 gnd.n4947 gnd.n4946 585
R5490 gnd.n3206 gnd.n3205 585
R5491 gnd.n4829 gnd.n3205 585
R5492 gnd.n4941 gnd.n4940 585
R5493 gnd.n4940 gnd.n4939 585
R5494 gnd.n3209 gnd.n3208 585
R5495 gnd.n4868 gnd.n3209 585
R5496 gnd.n4930 gnd.n4929 585
R5497 gnd.n4931 gnd.n4930 585
R5498 gnd.n3220 gnd.n3219 585
R5499 gnd.n4814 gnd.n3219 585
R5500 gnd.n4925 gnd.n4924 585
R5501 gnd.n4924 gnd.n4923 585
R5502 gnd.n3223 gnd.n3222 585
R5503 gnd.n4883 gnd.n3223 585
R5504 gnd.n4914 gnd.n4913 585
R5505 gnd.n4915 gnd.n4914 585
R5506 gnd.n3235 gnd.n3234 585
R5507 gnd.n3258 gnd.n3234 585
R5508 gnd.n4909 gnd.n4908 585
R5509 gnd.n4908 gnd.n4907 585
R5510 gnd.n3238 gnd.n3237 585
R5511 gnd.n3249 gnd.n3238 585
R5512 gnd.n3268 gnd.n3251 585
R5513 gnd.n4899 gnd.n3251 585
R5514 gnd.n4794 gnd.n4793 585
R5515 gnd.n4795 gnd.n4794 585
R5516 gnd.n3267 gnd.n3266 585
R5517 gnd.n3266 gnd.n3264 585
R5518 gnd.n4788 gnd.n4787 585
R5519 gnd.n4787 gnd.n4786 585
R5520 gnd.n3271 gnd.n3270 585
R5521 gnd.n4682 gnd.n3271 585
R5522 gnd.n4775 gnd.n4774 585
R5523 gnd.n4776 gnd.n4775 585
R5524 gnd.n3282 gnd.n3281 585
R5525 gnd.n4658 gnd.n3281 585
R5526 gnd.n4770 gnd.n4769 585
R5527 gnd.n4769 gnd.n4768 585
R5528 gnd.n3285 gnd.n3284 585
R5529 gnd.n4697 gnd.n3285 585
R5530 gnd.n4759 gnd.n4758 585
R5531 gnd.n4760 gnd.n4759 585
R5532 gnd.n3294 gnd.n3293 585
R5533 gnd.n4642 gnd.n3293 585
R5534 gnd.n4754 gnd.n4753 585
R5535 gnd.n4753 gnd.n4752 585
R5536 gnd.n3297 gnd.n3296 585
R5537 gnd.n4712 gnd.n3297 585
R5538 gnd.n4743 gnd.n4742 585
R5539 gnd.n4744 gnd.n4743 585
R5540 gnd.n3307 gnd.n3306 585
R5541 gnd.n3329 gnd.n3306 585
R5542 gnd.n4738 gnd.n4737 585
R5543 gnd.n4737 gnd.n4736 585
R5544 gnd.n3310 gnd.n3309 585
R5545 gnd.n3319 gnd.n3310 585
R5546 gnd.n3338 gnd.n3321 585
R5547 gnd.n4728 gnd.n3321 585
R5548 gnd.n4620 gnd.n4619 585
R5549 gnd.n4621 gnd.n4620 585
R5550 gnd.n3337 gnd.n3336 585
R5551 gnd.n4496 gnd.n3336 585
R5552 gnd.n4614 gnd.n4613 585
R5553 gnd.n4613 gnd.n4612 585
R5554 gnd.n3341 gnd.n3340 585
R5555 gnd.n4509 gnd.n3341 585
R5556 gnd.n4602 gnd.n4601 585
R5557 gnd.t6 gnd.n4602 585
R5558 gnd.n3354 gnd.n3353 585
R5559 gnd.n4483 gnd.n3353 585
R5560 gnd.n4597 gnd.n4596 585
R5561 gnd.n4596 gnd.n4595 585
R5562 gnd.n3357 gnd.n3356 585
R5563 gnd.n4524 gnd.n3357 585
R5564 gnd.n4586 gnd.n4585 585
R5565 gnd.n4587 gnd.n4586 585
R5566 gnd.n3368 gnd.n3367 585
R5567 gnd.n4468 gnd.n3367 585
R5568 gnd.n4581 gnd.n4580 585
R5569 gnd.n4580 gnd.n4579 585
R5570 gnd.n3371 gnd.n3370 585
R5571 gnd.n4539 gnd.n3371 585
R5572 gnd.n4570 gnd.n4569 585
R5573 gnd.n4571 gnd.n4570 585
R5574 gnd.n3382 gnd.n3381 585
R5575 gnd.n3405 gnd.n3381 585
R5576 gnd.n4565 gnd.n4564 585
R5577 gnd.n4564 gnd.n4563 585
R5578 gnd.n3385 gnd.n3384 585
R5579 gnd.n3395 gnd.n3385 585
R5580 gnd.n3413 gnd.n3397 585
R5581 gnd.n4555 gnd.n3397 585
R5582 gnd.n4449 gnd.n4448 585
R5583 gnd.n4450 gnd.n4449 585
R5584 gnd.n3412 gnd.n3411 585
R5585 gnd.n4162 gnd.n3411 585
R5586 gnd.n4443 gnd.n4442 585
R5587 gnd.n4442 gnd.n4441 585
R5588 gnd.n3416 gnd.n3415 585
R5589 gnd.n3426 gnd.n3416 585
R5590 gnd.n4430 gnd.n4429 585
R5591 gnd.n4431 gnd.n4430 585
R5592 gnd.n3429 gnd.n3428 585
R5593 gnd.n3433 gnd.n3428 585
R5594 gnd.n4425 gnd.n4424 585
R5595 gnd.n4424 gnd.n4423 585
R5596 gnd.n5409 gnd.n5408 585
R5597 gnd.n5408 gnd.n2685 585
R5598 gnd.n5410 gnd.n5407 585
R5599 gnd.n5405 gnd.n3094 585
R5600 gnd.n5414 gnd.n3093 585
R5601 gnd.n5418 gnd.n3091 585
R5602 gnd.n5419 gnd.n3090 585
R5603 gnd.n3088 gnd.n3086 585
R5604 gnd.n5423 gnd.n3085 585
R5605 gnd.n5424 gnd.n3083 585
R5606 gnd.n5425 gnd.n3082 585
R5607 gnd.n3080 gnd.n2960 585
R5608 gnd.n3079 gnd.n2961 585
R5609 gnd.n3077 gnd.n3076 585
R5610 gnd.n2963 gnd.n2962 585
R5611 gnd.n3067 gnd.n3066 585
R5612 gnd.n3064 gnd.n2973 585
R5613 gnd.n3062 gnd.n3061 585
R5614 gnd.n2975 gnd.n2974 585
R5615 gnd.n3050 gnd.n3049 585
R5616 gnd.n3047 gnd.n2982 585
R5617 gnd.n3045 gnd.n3044 585
R5618 gnd.n2984 gnd.n2983 585
R5619 gnd.n3033 gnd.n3032 585
R5620 gnd.n3030 gnd.n2991 585
R5621 gnd.n3028 gnd.n3027 585
R5622 gnd.n2993 gnd.n2992 585
R5623 gnd.n3016 gnd.n3015 585
R5624 gnd.n3013 gnd.n3011 585
R5625 gnd.n3000 gnd.n2681 585
R5626 gnd.n5232 gnd.n5055 506.916
R5627 gnd.n5163 gnd.n5056 506.916
R5628 gnd.n4281 gnd.n4279 506.916
R5629 gnd.n4267 gnd.n4266 506.916
R5630 gnd.n6323 gnd.n6322 442.322
R5631 gnd.n4145 gnd.t115 389.64
R5632 gnd.n5159 gnd.t50 389.64
R5633 gnd.n4200 gnd.t57 389.64
R5634 gnd.n5074 gnd.t106 389.64
R5635 gnd.n3457 gnd.t95 371.625
R5636 gnd.n7150 gnd.t29 371.625
R5637 gnd.n2967 gnd.t64 371.625
R5638 gnd.n3469 gnd.t85 371.625
R5639 gnd.n2744 gnd.t61 371.625
R5640 gnd.n2766 gnd.t36 371.625
R5641 gnd.n175 gnd.t124 371.625
R5642 gnd.n7243 gnd.t40 371.625
R5643 gnd.n2281 gnd.t118 371.625
R5644 gnd.n2303 gnd.t112 371.625
R5645 gnd.n3634 gnd.t46 371.625
R5646 gnd.n3612 gnd.t82 371.625
R5647 gnd.n3823 gnd.t71 371.625
R5648 gnd.n5415 gnd.t78 371.625
R5649 gnd.n1615 gnd.t22 323.425
R5650 gnd.n879 gnd.t91 323.425
R5651 gnd.n1227 gnd.n1201 289.615
R5652 gnd.n1195 gnd.n1169 289.615
R5653 gnd.n1163 gnd.n1137 289.615
R5654 gnd.n1132 gnd.n1106 289.615
R5655 gnd.n1100 gnd.n1074 289.615
R5656 gnd.n1068 gnd.n1042 289.615
R5657 gnd.n1036 gnd.n1010 289.615
R5658 gnd.n1005 gnd.n979 289.615
R5659 gnd.n1689 gnd.t67 279.217
R5660 gnd.n900 gnd.t99 279.217
R5661 gnd.n4170 gnd.t105 260.649
R5662 gnd.n5046 gnd.t111 260.649
R5663 gnd.n4185 gnd.n3427 256.663
R5664 gnd.n4187 gnd.n3427 256.663
R5665 gnd.n4256 gnd.n3427 256.663
R5666 gnd.n4250 gnd.n3427 256.663
R5667 gnd.n4248 gnd.n3427 256.663
R5668 gnd.n4242 gnd.n3427 256.663
R5669 gnd.n4240 gnd.n3427 256.663
R5670 gnd.n4234 gnd.n3427 256.663
R5671 gnd.n4232 gnd.n3427 256.663
R5672 gnd.n4226 gnd.n3427 256.663
R5673 gnd.n4224 gnd.n3427 256.663
R5674 gnd.n4218 gnd.n3427 256.663
R5675 gnd.n4216 gnd.n3427 256.663
R5676 gnd.n4210 gnd.n3427 256.663
R5677 gnd.n4203 gnd.n3427 256.663
R5678 gnd.n4204 gnd.n3427 256.663
R5679 gnd.n4347 gnd.n4143 256.663
R5680 gnd.n4345 gnd.n3427 256.663
R5681 gnd.n4343 gnd.n3427 256.663
R5682 gnd.n4336 gnd.n3427 256.663
R5683 gnd.n4334 gnd.n3427 256.663
R5684 gnd.n4328 gnd.n3427 256.663
R5685 gnd.n4326 gnd.n3427 256.663
R5686 gnd.n4320 gnd.n3427 256.663
R5687 gnd.n4318 gnd.n3427 256.663
R5688 gnd.n4312 gnd.n3427 256.663
R5689 gnd.n4310 gnd.n3427 256.663
R5690 gnd.n4304 gnd.n3427 256.663
R5691 gnd.n4302 gnd.n3427 256.663
R5692 gnd.n4296 gnd.n3427 256.663
R5693 gnd.n4294 gnd.n3427 256.663
R5694 gnd.n4288 gnd.n3427 256.663
R5695 gnd.n4286 gnd.n3427 256.663
R5696 gnd.n4280 gnd.n3427 256.663
R5697 gnd.n5229 gnd.n5142 256.663
R5698 gnd.n5229 gnd.n5143 256.663
R5699 gnd.n5229 gnd.n5144 256.663
R5700 gnd.n5229 gnd.n5145 256.663
R5701 gnd.n5229 gnd.n5146 256.663
R5702 gnd.n5229 gnd.n5147 256.663
R5703 gnd.n5229 gnd.n5148 256.663
R5704 gnd.n5229 gnd.n5149 256.663
R5705 gnd.n5229 gnd.n5150 256.663
R5706 gnd.n5229 gnd.n5151 256.663
R5707 gnd.n5229 gnd.n5152 256.663
R5708 gnd.n5229 gnd.n5153 256.663
R5709 gnd.n5229 gnd.n5154 256.663
R5710 gnd.n5229 gnd.n5155 256.663
R5711 gnd.n5229 gnd.n5156 256.663
R5712 gnd.n5229 gnd.n5157 256.663
R5713 gnd.n5158 gnd.n2741 256.663
R5714 gnd.n5229 gnd.n5141 256.663
R5715 gnd.n5229 gnd.n5073 256.663
R5716 gnd.n5229 gnd.n5072 256.663
R5717 gnd.n5229 gnd.n5071 256.663
R5718 gnd.n5229 gnd.n5070 256.663
R5719 gnd.n5229 gnd.n5069 256.663
R5720 gnd.n5229 gnd.n5068 256.663
R5721 gnd.n5229 gnd.n5067 256.663
R5722 gnd.n5229 gnd.n5066 256.663
R5723 gnd.n5229 gnd.n5065 256.663
R5724 gnd.n5229 gnd.n5064 256.663
R5725 gnd.n5229 gnd.n5063 256.663
R5726 gnd.n5229 gnd.n5062 256.663
R5727 gnd.n5229 gnd.n5061 256.663
R5728 gnd.n5229 gnd.n5060 256.663
R5729 gnd.n5229 gnd.n5059 256.663
R5730 gnd.n5229 gnd.n5058 256.663
R5731 gnd.n6076 gnd.n2249 242.672
R5732 gnd.n6076 gnd.n2250 242.672
R5733 gnd.n6076 gnd.n2251 242.672
R5734 gnd.n6076 gnd.n2252 242.672
R5735 gnd.n6076 gnd.n2253 242.672
R5736 gnd.n6076 gnd.n2254 242.672
R5737 gnd.n6076 gnd.n2255 242.672
R5738 gnd.n6076 gnd.n2256 242.672
R5739 gnd.n6076 gnd.n2257 242.672
R5740 gnd.n4378 gnd.n4377 242.672
R5741 gnd.n4377 gnd.n3571 242.672
R5742 gnd.n4377 gnd.n3479 242.672
R5743 gnd.n4377 gnd.n3478 242.672
R5744 gnd.n4377 gnd.n3477 242.672
R5745 gnd.n4377 gnd.n3476 242.672
R5746 gnd.n4377 gnd.n3475 242.672
R5747 gnd.n4377 gnd.n3474 242.672
R5748 gnd.n4377 gnd.n3473 242.672
R5749 gnd.n5698 gnd.n2711 242.672
R5750 gnd.n5698 gnd.n2712 242.672
R5751 gnd.n5698 gnd.n2713 242.672
R5752 gnd.n5698 gnd.n2714 242.672
R5753 gnd.n5698 gnd.n2715 242.672
R5754 gnd.n5698 gnd.n2716 242.672
R5755 gnd.n5698 gnd.n2717 242.672
R5756 gnd.n5698 gnd.n2718 242.672
R5757 gnd.n5698 gnd.n2719 242.672
R5758 gnd.n7152 gnd.n102 242.672
R5759 gnd.n7148 gnd.n102 242.672
R5760 gnd.n7143 gnd.n102 242.672
R5761 gnd.n7140 gnd.n102 242.672
R5762 gnd.n7135 gnd.n102 242.672
R5763 gnd.n7132 gnd.n102 242.672
R5764 gnd.n7127 gnd.n102 242.672
R5765 gnd.n7124 gnd.n102 242.672
R5766 gnd.n7119 gnd.n102 242.672
R5767 gnd.n1743 gnd.n1742 242.672
R5768 gnd.n1743 gnd.n1653 242.672
R5769 gnd.n1743 gnd.n1654 242.672
R5770 gnd.n1743 gnd.n1655 242.672
R5771 gnd.n1743 gnd.n1656 242.672
R5772 gnd.n1743 gnd.n1657 242.672
R5773 gnd.n1743 gnd.n1658 242.672
R5774 gnd.n1743 gnd.n1659 242.672
R5775 gnd.n1743 gnd.n1660 242.672
R5776 gnd.n1743 gnd.n1661 242.672
R5777 gnd.n1743 gnd.n1662 242.672
R5778 gnd.n1743 gnd.n1663 242.672
R5779 gnd.n1744 gnd.n1743 242.672
R5780 gnd.n6123 gnd.n2230 242.672
R5781 gnd.n6123 gnd.n896 242.672
R5782 gnd.n6123 gnd.n895 242.672
R5783 gnd.n6123 gnd.n894 242.672
R5784 gnd.n6123 gnd.n893 242.672
R5785 gnd.n6123 gnd.n892 242.672
R5786 gnd.n6123 gnd.n891 242.672
R5787 gnd.n6123 gnd.n890 242.672
R5788 gnd.n6123 gnd.n889 242.672
R5789 gnd.n6123 gnd.n888 242.672
R5790 gnd.n6123 gnd.n887 242.672
R5791 gnd.n6123 gnd.n886 242.672
R5792 gnd.n6123 gnd.n885 242.672
R5793 gnd.n1827 gnd.n1826 242.672
R5794 gnd.n1826 gnd.n1565 242.672
R5795 gnd.n1826 gnd.n1566 242.672
R5796 gnd.n1826 gnd.n1567 242.672
R5797 gnd.n1826 gnd.n1568 242.672
R5798 gnd.n1826 gnd.n1569 242.672
R5799 gnd.n1826 gnd.n1570 242.672
R5800 gnd.n1826 gnd.n1571 242.672
R5801 gnd.n6123 gnd.n878 242.672
R5802 gnd.n6124 gnd.n6123 242.672
R5803 gnd.n6123 gnd.n6077 242.672
R5804 gnd.n6123 gnd.n6078 242.672
R5805 gnd.n6123 gnd.n6079 242.672
R5806 gnd.n6123 gnd.n6080 242.672
R5807 gnd.n6123 gnd.n6081 242.672
R5808 gnd.n6123 gnd.n6082 242.672
R5809 gnd.n6076 gnd.n6075 242.672
R5810 gnd.n6076 gnd.n2231 242.672
R5811 gnd.n6076 gnd.n2232 242.672
R5812 gnd.n6076 gnd.n2233 242.672
R5813 gnd.n6076 gnd.n2234 242.672
R5814 gnd.n6076 gnd.n2235 242.672
R5815 gnd.n6076 gnd.n2236 242.672
R5816 gnd.n6076 gnd.n2237 242.672
R5817 gnd.n6076 gnd.n2238 242.672
R5818 gnd.n6076 gnd.n2239 242.672
R5819 gnd.n6076 gnd.n2240 242.672
R5820 gnd.n6076 gnd.n2241 242.672
R5821 gnd.n6076 gnd.n2242 242.672
R5822 gnd.n6076 gnd.n2243 242.672
R5823 gnd.n6076 gnd.n2244 242.672
R5824 gnd.n6076 gnd.n2245 242.672
R5825 gnd.n6076 gnd.n2246 242.672
R5826 gnd.n6076 gnd.n2247 242.672
R5827 gnd.n6076 gnd.n2248 242.672
R5828 gnd.n4377 gnd.n3573 242.672
R5829 gnd.n4377 gnd.n3574 242.672
R5830 gnd.n4377 gnd.n3575 242.672
R5831 gnd.n4377 gnd.n3576 242.672
R5832 gnd.n4377 gnd.n3577 242.672
R5833 gnd.n4377 gnd.n3578 242.672
R5834 gnd.n4377 gnd.n3579 242.672
R5835 gnd.n4377 gnd.n3580 242.672
R5836 gnd.n4377 gnd.n3581 242.672
R5837 gnd.n4377 gnd.n3582 242.672
R5838 gnd.n4377 gnd.n3583 242.672
R5839 gnd.n4348 gnd.n3614 242.672
R5840 gnd.n4377 gnd.n3584 242.672
R5841 gnd.n4377 gnd.n3585 242.672
R5842 gnd.n4377 gnd.n3586 242.672
R5843 gnd.n4377 gnd.n3587 242.672
R5844 gnd.n4377 gnd.n3588 242.672
R5845 gnd.n4377 gnd.n3589 242.672
R5846 gnd.n4377 gnd.n3590 242.672
R5847 gnd.n4377 gnd.n4376 242.672
R5848 gnd.n5698 gnd.n5697 242.672
R5849 gnd.n5698 gnd.n2693 242.672
R5850 gnd.n5698 gnd.n2694 242.672
R5851 gnd.n5698 gnd.n2695 242.672
R5852 gnd.n5698 gnd.n2696 242.672
R5853 gnd.n5698 gnd.n2697 242.672
R5854 gnd.n5698 gnd.n2698 242.672
R5855 gnd.n5698 gnd.n2699 242.672
R5856 gnd.n5666 gnd.n2742 242.672
R5857 gnd.n5698 gnd.n2700 242.672
R5858 gnd.n5698 gnd.n2701 242.672
R5859 gnd.n5698 gnd.n2702 242.672
R5860 gnd.n5698 gnd.n2703 242.672
R5861 gnd.n5698 gnd.n2704 242.672
R5862 gnd.n5698 gnd.n2705 242.672
R5863 gnd.n5698 gnd.n2706 242.672
R5864 gnd.n5698 gnd.n2707 242.672
R5865 gnd.n5698 gnd.n2708 242.672
R5866 gnd.n5698 gnd.n2709 242.672
R5867 gnd.n5698 gnd.n2710 242.672
R5868 gnd.n172 gnd.n102 242.672
R5869 gnd.n7211 gnd.n102 242.672
R5870 gnd.n168 gnd.n102 242.672
R5871 gnd.n7218 gnd.n102 242.672
R5872 gnd.n161 gnd.n102 242.672
R5873 gnd.n7225 gnd.n102 242.672
R5874 gnd.n154 gnd.n102 242.672
R5875 gnd.n7232 gnd.n102 242.672
R5876 gnd.n147 gnd.n102 242.672
R5877 gnd.n7239 gnd.n102 242.672
R5878 gnd.n140 gnd.n102 242.672
R5879 gnd.n7249 gnd.n102 242.672
R5880 gnd.n133 gnd.n102 242.672
R5881 gnd.n7256 gnd.n102 242.672
R5882 gnd.n126 gnd.n102 242.672
R5883 gnd.n7263 gnd.n102 242.672
R5884 gnd.n119 gnd.n102 242.672
R5885 gnd.n7270 gnd.n102 242.672
R5886 gnd.n112 gnd.n102 242.672
R5887 gnd.n4415 gnd.n3440 242.672
R5888 gnd.n4415 gnd.n3441 242.672
R5889 gnd.n4415 gnd.n3442 242.672
R5890 gnd.n4415 gnd.n3443 242.672
R5891 gnd.n4415 gnd.n3444 242.672
R5892 gnd.n4415 gnd.n3445 242.672
R5893 gnd.n4415 gnd.n3446 242.672
R5894 gnd.n4415 gnd.n3447 242.672
R5895 gnd.n4415 gnd.n3448 242.672
R5896 gnd.n4415 gnd.n3449 242.672
R5897 gnd.n4415 gnd.n3450 242.672
R5898 gnd.n4415 gnd.n3451 242.672
R5899 gnd.n4415 gnd.n3452 242.672
R5900 gnd.n4415 gnd.n4414 242.672
R5901 gnd.n5406 gnd.n2685 242.672
R5902 gnd.n3092 gnd.n2685 242.672
R5903 gnd.n3089 gnd.n2685 242.672
R5904 gnd.n3084 gnd.n2685 242.672
R5905 gnd.n3081 gnd.n2685 242.672
R5906 gnd.n3078 gnd.n2685 242.672
R5907 gnd.n3065 gnd.n2685 242.672
R5908 gnd.n3063 gnd.n2685 242.672
R5909 gnd.n3048 gnd.n2685 242.672
R5910 gnd.n3046 gnd.n2685 242.672
R5911 gnd.n3031 gnd.n2685 242.672
R5912 gnd.n3029 gnd.n2685 242.672
R5913 gnd.n3014 gnd.n2685 242.672
R5914 gnd.n3012 gnd.n2685 242.672
R5915 gnd.n109 gnd.n105 240.244
R5916 gnd.n7272 gnd.n7271 240.244
R5917 gnd.n7269 gnd.n113 240.244
R5918 gnd.n7265 gnd.n7264 240.244
R5919 gnd.n7262 gnd.n120 240.244
R5920 gnd.n7258 gnd.n7257 240.244
R5921 gnd.n7255 gnd.n127 240.244
R5922 gnd.n7251 gnd.n7250 240.244
R5923 gnd.n7248 gnd.n134 240.244
R5924 gnd.n7241 gnd.n7240 240.244
R5925 gnd.n7238 gnd.n141 240.244
R5926 gnd.n7234 gnd.n7233 240.244
R5927 gnd.n7231 gnd.n148 240.244
R5928 gnd.n7227 gnd.n7226 240.244
R5929 gnd.n7224 gnd.n155 240.244
R5930 gnd.n7220 gnd.n7219 240.244
R5931 gnd.n7217 gnd.n162 240.244
R5932 gnd.n7213 gnd.n7212 240.244
R5933 gnd.n7210 gnd.n169 240.244
R5934 gnd.n5623 gnd.n2770 240.244
R5935 gnd.n2954 gnd.n2770 240.244
R5936 gnd.n2954 gnd.n2902 240.244
R5937 gnd.n2950 gnd.n2902 240.244
R5938 gnd.n2950 gnd.n2892 240.244
R5939 gnd.n2947 gnd.n2892 240.244
R5940 gnd.n2947 gnd.n2884 240.244
R5941 gnd.n2884 gnd.n2873 240.244
R5942 gnd.n2943 gnd.n2873 240.244
R5943 gnd.n2943 gnd.n2864 240.244
R5944 gnd.n2940 gnd.n2864 240.244
R5945 gnd.n2940 gnd.n2856 240.244
R5946 gnd.n2856 gnd.n2845 240.244
R5947 gnd.n2845 gnd.n2834 240.244
R5948 gnd.n5526 gnd.n2834 240.244
R5949 gnd.n5526 gnd.n2835 240.244
R5950 gnd.n2835 gnd.n2822 240.244
R5951 gnd.n2822 gnd.n2811 240.244
R5952 gnd.n5533 gnd.n2811 240.244
R5953 gnd.n5533 gnd.n2802 240.244
R5954 gnd.n5547 gnd.n2802 240.244
R5955 gnd.n5547 gnd.n273 240.244
R5956 gnd.n307 gnd.n273 240.244
R5957 gnd.n5542 gnd.n307 240.244
R5958 gnd.n5542 gnd.n296 240.244
R5959 gnd.n6953 gnd.n296 240.244
R5960 gnd.n6953 gnd.n293 240.244
R5961 gnd.n7016 gnd.n293 240.244
R5962 gnd.n7016 gnd.n290 240.244
R5963 gnd.n7012 gnd.n290 240.244
R5964 gnd.n7012 gnd.n258 240.244
R5965 gnd.n7007 gnd.n258 240.244
R5966 gnd.n7007 gnd.n252 240.244
R5967 gnd.n7004 gnd.n252 240.244
R5968 gnd.n7004 gnd.n245 240.244
R5969 gnd.n7001 gnd.n245 240.244
R5970 gnd.n7001 gnd.n235 240.244
R5971 gnd.n6998 gnd.n235 240.244
R5972 gnd.n6998 gnd.n228 240.244
R5973 gnd.n6995 gnd.n228 240.244
R5974 gnd.n6995 gnd.n222 240.244
R5975 gnd.n6992 gnd.n222 240.244
R5976 gnd.n6992 gnd.n215 240.244
R5977 gnd.n6989 gnd.n215 240.244
R5978 gnd.n6989 gnd.n205 240.244
R5979 gnd.n6986 gnd.n205 240.244
R5980 gnd.n6986 gnd.n198 240.244
R5981 gnd.n6983 gnd.n198 240.244
R5982 gnd.n6983 gnd.n189 240.244
R5983 gnd.n189 gnd.n179 240.244
R5984 gnd.n7201 gnd.n179 240.244
R5985 gnd.n7202 gnd.n7201 240.244
R5986 gnd.n7202 gnd.n101 240.244
R5987 gnd.n2723 gnd.n2722 240.244
R5988 gnd.n5691 gnd.n2722 240.244
R5989 gnd.n5689 gnd.n5688 240.244
R5990 gnd.n5685 gnd.n5684 240.244
R5991 gnd.n5681 gnd.n5680 240.244
R5992 gnd.n5677 gnd.n5676 240.244
R5993 gnd.n5673 gnd.n5672 240.244
R5994 gnd.n5669 gnd.n5668 240.244
R5995 gnd.n5664 gnd.n5663 240.244
R5996 gnd.n5660 gnd.n5659 240.244
R5997 gnd.n5656 gnd.n5655 240.244
R5998 gnd.n5652 gnd.n5651 240.244
R5999 gnd.n5648 gnd.n5647 240.244
R6000 gnd.n5644 gnd.n5643 240.244
R6001 gnd.n5640 gnd.n5639 240.244
R6002 gnd.n5636 gnd.n5635 240.244
R6003 gnd.n5632 gnd.n5631 240.244
R6004 gnd.n2765 gnd.n2764 240.244
R6005 gnd.n2922 gnd.n2724 240.244
R6006 gnd.n2922 gnd.n2900 240.244
R6007 gnd.n5448 gnd.n2900 240.244
R6008 gnd.n5448 gnd.n2895 240.244
R6009 gnd.n5456 gnd.n2895 240.244
R6010 gnd.n5456 gnd.n2896 240.244
R6011 gnd.n2896 gnd.n2871 240.244
R6012 gnd.n5479 gnd.n2871 240.244
R6013 gnd.n5479 gnd.n2866 240.244
R6014 gnd.n5487 gnd.n2866 240.244
R6015 gnd.n5487 gnd.n2867 240.244
R6016 gnd.n2867 gnd.n2843 240.244
R6017 gnd.n5516 gnd.n2843 240.244
R6018 gnd.n5516 gnd.n2838 240.244
R6019 gnd.n5524 gnd.n2838 240.244
R6020 gnd.n5524 gnd.n2839 240.244
R6021 gnd.n2839 gnd.n2809 240.244
R6022 gnd.n5580 gnd.n2809 240.244
R6023 gnd.n5580 gnd.n2805 240.244
R6024 gnd.n5586 gnd.n2805 240.244
R6025 gnd.n5586 gnd.n270 240.244
R6026 gnd.n7039 gnd.n270 240.244
R6027 gnd.n7039 gnd.n271 240.244
R6028 gnd.n300 gnd.n271 240.244
R6029 gnd.n6948 gnd.n300 240.244
R6030 gnd.n6951 gnd.n6948 240.244
R6031 gnd.n6951 gnd.n292 240.244
R6032 gnd.n7018 gnd.n292 240.244
R6033 gnd.n7021 gnd.n7018 240.244
R6034 gnd.n7021 gnd.n260 240.244
R6035 gnd.n7044 gnd.n260 240.244
R6036 gnd.n7044 gnd.n250 240.244
R6037 gnd.n7054 gnd.n250 240.244
R6038 gnd.n7054 gnd.n246 240.244
R6039 gnd.n7060 gnd.n246 240.244
R6040 gnd.n7060 gnd.n233 240.244
R6041 gnd.n7070 gnd.n233 240.244
R6042 gnd.n7070 gnd.n229 240.244
R6043 gnd.n7076 gnd.n229 240.244
R6044 gnd.n7076 gnd.n220 240.244
R6045 gnd.n7086 gnd.n220 240.244
R6046 gnd.n7086 gnd.n216 240.244
R6047 gnd.n7092 gnd.n216 240.244
R6048 gnd.n7092 gnd.n203 240.244
R6049 gnd.n7102 gnd.n203 240.244
R6050 gnd.n7102 gnd.n199 240.244
R6051 gnd.n7108 gnd.n199 240.244
R6052 gnd.n7108 gnd.n187 240.244
R6053 gnd.n7193 gnd.n187 240.244
R6054 gnd.n7193 gnd.n183 240.244
R6055 gnd.n7199 gnd.n183 240.244
R6056 gnd.n7199 gnd.n104 240.244
R6057 gnd.n7279 gnd.n104 240.244
R6058 gnd.n3591 gnd.n2568 240.244
R6059 gnd.n4375 gnd.n3592 240.244
R6060 gnd.n4371 gnd.n4370 240.244
R6061 gnd.n4367 gnd.n4366 240.244
R6062 gnd.n4363 gnd.n4362 240.244
R6063 gnd.n4359 gnd.n4358 240.244
R6064 gnd.n4355 gnd.n4354 240.244
R6065 gnd.n4351 gnd.n4350 240.244
R6066 gnd.n4136 gnd.n4135 240.244
R6067 gnd.n4133 gnd.n4132 240.244
R6068 gnd.n4129 gnd.n4128 240.244
R6069 gnd.n4125 gnd.n4124 240.244
R6070 gnd.n4121 gnd.n4120 240.244
R6071 gnd.n4117 gnd.n4116 240.244
R6072 gnd.n4113 gnd.n4112 240.244
R6073 gnd.n4109 gnd.n4108 240.244
R6074 gnd.n4105 gnd.n4104 240.244
R6075 gnd.n4101 gnd.n4100 240.244
R6076 gnd.n5997 gnd.n2307 240.244
R6077 gnd.n2311 gnd.n2307 240.244
R6078 gnd.n5990 gnd.n2311 240.244
R6079 gnd.n5990 gnd.n2312 240.244
R6080 gnd.n2325 gnd.n2312 240.244
R6081 gnd.n3934 gnd.n2325 240.244
R6082 gnd.n3934 gnd.n2336 240.244
R6083 gnd.n3937 gnd.n2336 240.244
R6084 gnd.n3937 gnd.n2346 240.244
R6085 gnd.n3942 gnd.n2346 240.244
R6086 gnd.n3942 gnd.n2356 240.244
R6087 gnd.n3945 gnd.n2356 240.244
R6088 gnd.n3945 gnd.n2366 240.244
R6089 gnd.n3950 gnd.n2366 240.244
R6090 gnd.n3950 gnd.n2376 240.244
R6091 gnd.n3953 gnd.n2376 240.244
R6092 gnd.n3953 gnd.n2386 240.244
R6093 gnd.n3958 gnd.n2386 240.244
R6094 gnd.n3958 gnd.n2396 240.244
R6095 gnd.n3961 gnd.n2396 240.244
R6096 gnd.n3961 gnd.n2406 240.244
R6097 gnd.n3967 gnd.n2406 240.244
R6098 gnd.n3967 gnd.n2416 240.244
R6099 gnd.n3977 gnd.n2416 240.244
R6100 gnd.n3977 gnd.n2425 240.244
R6101 gnd.n3985 gnd.n2425 240.244
R6102 gnd.n3985 gnd.n2435 240.244
R6103 gnd.n3996 gnd.n2435 240.244
R6104 gnd.n3996 gnd.n2443 240.244
R6105 gnd.n4002 gnd.n2443 240.244
R6106 gnd.n4002 gnd.n2454 240.244
R6107 gnd.n4012 gnd.n2454 240.244
R6108 gnd.n4012 gnd.n2464 240.244
R6109 gnd.n4018 gnd.n2464 240.244
R6110 gnd.n4018 gnd.n2474 240.244
R6111 gnd.n4028 gnd.n2474 240.244
R6112 gnd.n4028 gnd.n2485 240.244
R6113 gnd.n4034 gnd.n2485 240.244
R6114 gnd.n4034 gnd.n2496 240.244
R6115 gnd.n4044 gnd.n2496 240.244
R6116 gnd.n4044 gnd.n2507 240.244
R6117 gnd.n4050 gnd.n2507 240.244
R6118 gnd.n4050 gnd.n2517 240.244
R6119 gnd.n4060 gnd.n2517 240.244
R6120 gnd.n4060 gnd.n2528 240.244
R6121 gnd.n4066 gnd.n2528 240.244
R6122 gnd.n4066 gnd.n2539 240.244
R6123 gnd.n4076 gnd.n2539 240.244
R6124 gnd.n4076 gnd.n2550 240.244
R6125 gnd.n4083 gnd.n2550 240.244
R6126 gnd.n4083 gnd.n2561 240.244
R6127 gnd.n4093 gnd.n2561 240.244
R6128 gnd.n4093 gnd.n2570 240.244
R6129 gnd.n2261 gnd.n2260 240.244
R6130 gnd.n6069 gnd.n2260 240.244
R6131 gnd.n6067 gnd.n6066 240.244
R6132 gnd.n6063 gnd.n6062 240.244
R6133 gnd.n6059 gnd.n6058 240.244
R6134 gnd.n6055 gnd.n6054 240.244
R6135 gnd.n6051 gnd.n6050 240.244
R6136 gnd.n6047 gnd.n6046 240.244
R6137 gnd.n6043 gnd.n6042 240.244
R6138 gnd.n6038 gnd.n6037 240.244
R6139 gnd.n6034 gnd.n6033 240.244
R6140 gnd.n6030 gnd.n6029 240.244
R6141 gnd.n6026 gnd.n6025 240.244
R6142 gnd.n6022 gnd.n6021 240.244
R6143 gnd.n6018 gnd.n6017 240.244
R6144 gnd.n6014 gnd.n6013 240.244
R6145 gnd.n6010 gnd.n6009 240.244
R6146 gnd.n6006 gnd.n6005 240.244
R6147 gnd.n2302 gnd.n2301 240.244
R6148 gnd.n3880 gnd.n2262 240.244
R6149 gnd.n3880 gnd.n2317 240.244
R6150 gnd.n5988 gnd.n2317 240.244
R6151 gnd.n5988 gnd.n2318 240.244
R6152 gnd.n5984 gnd.n2318 240.244
R6153 gnd.n5984 gnd.n2324 240.244
R6154 gnd.n5976 gnd.n2324 240.244
R6155 gnd.n5976 gnd.n2339 240.244
R6156 gnd.n5972 gnd.n2339 240.244
R6157 gnd.n5972 gnd.n2345 240.244
R6158 gnd.n5964 gnd.n2345 240.244
R6159 gnd.n5964 gnd.n2358 240.244
R6160 gnd.n5960 gnd.n2358 240.244
R6161 gnd.n5960 gnd.n2364 240.244
R6162 gnd.n5952 gnd.n2364 240.244
R6163 gnd.n5952 gnd.n2379 240.244
R6164 gnd.n5948 gnd.n2379 240.244
R6165 gnd.n5948 gnd.n2385 240.244
R6166 gnd.n5940 gnd.n2385 240.244
R6167 gnd.n5940 gnd.n2398 240.244
R6168 gnd.n5936 gnd.n2398 240.244
R6169 gnd.n5936 gnd.n2404 240.244
R6170 gnd.n5928 gnd.n2404 240.244
R6171 gnd.n5928 gnd.n2419 240.244
R6172 gnd.n5924 gnd.n2419 240.244
R6173 gnd.n5924 gnd.n2423 240.244
R6174 gnd.n5916 gnd.n2423 240.244
R6175 gnd.n5916 gnd.n2438 240.244
R6176 gnd.n5911 gnd.n2438 240.244
R6177 gnd.n5911 gnd.n2441 240.244
R6178 gnd.n5903 gnd.n2441 240.244
R6179 gnd.n5903 gnd.n2457 240.244
R6180 gnd.n5899 gnd.n2457 240.244
R6181 gnd.n5899 gnd.n2462 240.244
R6182 gnd.n5891 gnd.n2462 240.244
R6183 gnd.n5891 gnd.n2477 240.244
R6184 gnd.n5887 gnd.n2477 240.244
R6185 gnd.n5887 gnd.n2483 240.244
R6186 gnd.n5879 gnd.n2483 240.244
R6187 gnd.n5879 gnd.n2499 240.244
R6188 gnd.n5875 gnd.n2499 240.244
R6189 gnd.n5875 gnd.n2505 240.244
R6190 gnd.n5867 gnd.n2505 240.244
R6191 gnd.n5867 gnd.n2520 240.244
R6192 gnd.n5863 gnd.n2520 240.244
R6193 gnd.n5863 gnd.n2526 240.244
R6194 gnd.n5855 gnd.n2526 240.244
R6195 gnd.n5855 gnd.n2542 240.244
R6196 gnd.n5851 gnd.n2542 240.244
R6197 gnd.n5851 gnd.n2548 240.244
R6198 gnd.n5843 gnd.n2548 240.244
R6199 gnd.n5843 gnd.n2563 240.244
R6200 gnd.n5839 gnd.n2563 240.244
R6201 gnd.n6122 gnd.n6083 240.244
R6202 gnd.n6115 gnd.n6114 240.244
R6203 gnd.n6112 gnd.n6111 240.244
R6204 gnd.n6108 gnd.n6107 240.244
R6205 gnd.n6104 gnd.n6103 240.244
R6206 gnd.n6100 gnd.n6099 240.244
R6207 gnd.n6096 gnd.n884 240.244
R6208 gnd.n6126 gnd.n6125 240.244
R6209 gnd.n1838 gnd.n1550 240.244
R6210 gnd.n1848 gnd.n1550 240.244
R6211 gnd.n1848 gnd.n1541 240.244
R6212 gnd.n1541 gnd.n1530 240.244
R6213 gnd.n1869 gnd.n1530 240.244
R6214 gnd.n1869 gnd.n1524 240.244
R6215 gnd.n1879 gnd.n1524 240.244
R6216 gnd.n1879 gnd.n1513 240.244
R6217 gnd.n1513 gnd.n1505 240.244
R6218 gnd.n1897 gnd.n1505 240.244
R6219 gnd.n1898 gnd.n1897 240.244
R6220 gnd.n1898 gnd.n1490 240.244
R6221 gnd.n1900 gnd.n1490 240.244
R6222 gnd.n1900 gnd.n1476 240.244
R6223 gnd.n1942 gnd.n1476 240.244
R6224 gnd.n1943 gnd.n1942 240.244
R6225 gnd.n1946 gnd.n1943 240.244
R6226 gnd.n1946 gnd.n1431 240.244
R6227 gnd.n1471 gnd.n1431 240.244
R6228 gnd.n1471 gnd.n1441 240.244
R6229 gnd.n1956 gnd.n1441 240.244
R6230 gnd.n1956 gnd.n1462 240.244
R6231 gnd.n1966 gnd.n1462 240.244
R6232 gnd.n1966 gnd.n1360 240.244
R6233 gnd.n2011 gnd.n1360 240.244
R6234 gnd.n2011 gnd.n1346 240.244
R6235 gnd.n2033 gnd.n1346 240.244
R6236 gnd.n2034 gnd.n2033 240.244
R6237 gnd.n2034 gnd.n1333 240.244
R6238 gnd.n1333 gnd.n1322 240.244
R6239 gnd.n2065 gnd.n1322 240.244
R6240 gnd.n2066 gnd.n2065 240.244
R6241 gnd.n2067 gnd.n2066 240.244
R6242 gnd.n2067 gnd.n1307 240.244
R6243 gnd.n1307 gnd.n1306 240.244
R6244 gnd.n1306 gnd.n1291 240.244
R6245 gnd.n2118 gnd.n1291 240.244
R6246 gnd.n2119 gnd.n2118 240.244
R6247 gnd.n2119 gnd.n1278 240.244
R6248 gnd.n1278 gnd.n1267 240.244
R6249 gnd.n2150 gnd.n1267 240.244
R6250 gnd.n2151 gnd.n2150 240.244
R6251 gnd.n2152 gnd.n2151 240.244
R6252 gnd.n2152 gnd.n1251 240.244
R6253 gnd.n2154 gnd.n1251 240.244
R6254 gnd.n2154 gnd.n1238 240.244
R6255 gnd.n2209 gnd.n1238 240.244
R6256 gnd.n2210 gnd.n2209 240.244
R6257 gnd.n2211 gnd.n2210 240.244
R6258 gnd.n2211 gnd.n859 240.244
R6259 gnd.n2219 gnd.n859 240.244
R6260 gnd.n2219 gnd.n869 240.244
R6261 gnd.n6133 gnd.n869 240.244
R6262 gnd.n1828 gnd.n1563 240.244
R6263 gnd.n1584 gnd.n1563 240.244
R6264 gnd.n1587 gnd.n1586 240.244
R6265 gnd.n1594 gnd.n1593 240.244
R6266 gnd.n1597 gnd.n1596 240.244
R6267 gnd.n1604 gnd.n1603 240.244
R6268 gnd.n1607 gnd.n1606 240.244
R6269 gnd.n1614 gnd.n1613 240.244
R6270 gnd.n1836 gnd.n1560 240.244
R6271 gnd.n1560 gnd.n1539 240.244
R6272 gnd.n1859 gnd.n1539 240.244
R6273 gnd.n1859 gnd.n1533 240.244
R6274 gnd.n1867 gnd.n1533 240.244
R6275 gnd.n1867 gnd.n1535 240.244
R6276 gnd.n1535 gnd.n1511 240.244
R6277 gnd.n1889 gnd.n1511 240.244
R6278 gnd.n1889 gnd.n1507 240.244
R6279 gnd.n1895 gnd.n1507 240.244
R6280 gnd.n1895 gnd.n1489 240.244
R6281 gnd.n1920 gnd.n1489 240.244
R6282 gnd.n1920 gnd.n1484 240.244
R6283 gnd.n1932 gnd.n1484 240.244
R6284 gnd.n1932 gnd.n1485 240.244
R6285 gnd.n1928 gnd.n1485 240.244
R6286 gnd.n1928 gnd.n1433 240.244
R6287 gnd.n1980 gnd.n1433 240.244
R6288 gnd.n1980 gnd.n1434 240.244
R6289 gnd.n1976 gnd.n1434 240.244
R6290 gnd.n1976 gnd.n1440 240.244
R6291 gnd.n1460 gnd.n1440 240.244
R6292 gnd.n1460 gnd.n1358 240.244
R6293 gnd.n2015 gnd.n1358 240.244
R6294 gnd.n2015 gnd.n1353 240.244
R6295 gnd.n2023 gnd.n1353 240.244
R6296 gnd.n2023 gnd.n1354 240.244
R6297 gnd.n1354 gnd.n1331 240.244
R6298 gnd.n2055 gnd.n1331 240.244
R6299 gnd.n2055 gnd.n1326 240.244
R6300 gnd.n2063 gnd.n1326 240.244
R6301 gnd.n2063 gnd.n1327 240.244
R6302 gnd.n1327 gnd.n1304 240.244
R6303 gnd.n2100 gnd.n1304 240.244
R6304 gnd.n2100 gnd.n1299 240.244
R6305 gnd.n2108 gnd.n1299 240.244
R6306 gnd.n2108 gnd.n1300 240.244
R6307 gnd.n1300 gnd.n1276 240.244
R6308 gnd.n2140 gnd.n1276 240.244
R6309 gnd.n2140 gnd.n1271 240.244
R6310 gnd.n2148 gnd.n1271 240.244
R6311 gnd.n2148 gnd.n1272 240.244
R6312 gnd.n1272 gnd.n1250 240.244
R6313 gnd.n2187 gnd.n1250 240.244
R6314 gnd.n2187 gnd.n1245 240.244
R6315 gnd.n2199 gnd.n1245 240.244
R6316 gnd.n2199 gnd.n1246 240.244
R6317 gnd.n2195 gnd.n1246 240.244
R6318 gnd.n2195 gnd.n860 240.244
R6319 gnd.n6145 gnd.n860 240.244
R6320 gnd.n6145 gnd.n861 240.244
R6321 gnd.n6141 gnd.n861 240.244
R6322 gnd.n6141 gnd.n867 240.244
R6323 gnd.n913 gnd.n873 240.244
R6324 gnd.n921 gnd.n920 240.244
R6325 gnd.n924 gnd.n923 240.244
R6326 gnd.n931 gnd.n930 240.244
R6327 gnd.n934 gnd.n933 240.244
R6328 gnd.n941 gnd.n940 240.244
R6329 gnd.n944 gnd.n943 240.244
R6330 gnd.n951 gnd.n950 240.244
R6331 gnd.n954 gnd.n953 240.244
R6332 gnd.n961 gnd.n960 240.244
R6333 gnd.n964 gnd.n963 240.244
R6334 gnd.n971 gnd.n970 240.244
R6335 gnd.n973 gnd.n897 240.244
R6336 gnd.n1751 gnd.n1648 240.244
R6337 gnd.n1751 gnd.n1641 240.244
R6338 gnd.n1762 gnd.n1641 240.244
R6339 gnd.n1762 gnd.n1637 240.244
R6340 gnd.n1768 gnd.n1637 240.244
R6341 gnd.n1768 gnd.n1629 240.244
R6342 gnd.n1778 gnd.n1629 240.244
R6343 gnd.n1778 gnd.n1624 240.244
R6344 gnd.n1814 gnd.n1624 240.244
R6345 gnd.n1814 gnd.n1625 240.244
R6346 gnd.n1625 gnd.n1572 240.244
R6347 gnd.n1809 gnd.n1572 240.244
R6348 gnd.n1809 gnd.n1808 240.244
R6349 gnd.n1808 gnd.n1551 240.244
R6350 gnd.n1804 gnd.n1551 240.244
R6351 gnd.n1804 gnd.n1542 240.244
R6352 gnd.n1801 gnd.n1542 240.244
R6353 gnd.n1801 gnd.n1800 240.244
R6354 gnd.n1800 gnd.n1525 240.244
R6355 gnd.n1796 gnd.n1525 240.244
R6356 gnd.n1796 gnd.n1514 240.244
R6357 gnd.n1514 gnd.n1495 240.244
R6358 gnd.n1909 gnd.n1495 240.244
R6359 gnd.n1909 gnd.n1491 240.244
R6360 gnd.n1917 gnd.n1491 240.244
R6361 gnd.n1917 gnd.n1482 240.244
R6362 gnd.n1482 gnd.n1418 240.244
R6363 gnd.n1989 gnd.n1418 240.244
R6364 gnd.n1989 gnd.n1419 240.244
R6365 gnd.n1430 gnd.n1419 240.244
R6366 gnd.n1465 gnd.n1430 240.244
R6367 gnd.n1468 gnd.n1465 240.244
R6368 gnd.n1468 gnd.n1442 240.244
R6369 gnd.n1455 gnd.n1442 240.244
R6370 gnd.n1455 gnd.n1452 240.244
R6371 gnd.n1452 gnd.n1361 240.244
R6372 gnd.n2010 gnd.n1361 240.244
R6373 gnd.n2010 gnd.n1351 240.244
R6374 gnd.n2006 gnd.n1351 240.244
R6375 gnd.n2006 gnd.n1345 240.244
R6376 gnd.n2003 gnd.n1345 240.244
R6377 gnd.n2003 gnd.n1334 240.244
R6378 gnd.n2000 gnd.n1334 240.244
R6379 gnd.n2000 gnd.n1312 240.244
R6380 gnd.n2076 gnd.n1312 240.244
R6381 gnd.n2076 gnd.n1308 240.244
R6382 gnd.n2097 gnd.n1308 240.244
R6383 gnd.n2097 gnd.n1297 240.244
R6384 gnd.n2093 gnd.n1297 240.244
R6385 gnd.n2093 gnd.n1290 240.244
R6386 gnd.n2090 gnd.n1290 240.244
R6387 gnd.n2090 gnd.n1279 240.244
R6388 gnd.n2087 gnd.n1279 240.244
R6389 gnd.n2087 gnd.n1256 240.244
R6390 gnd.n2163 gnd.n1256 240.244
R6391 gnd.n2163 gnd.n1252 240.244
R6392 gnd.n2184 gnd.n1252 240.244
R6393 gnd.n2184 gnd.n1244 240.244
R6394 gnd.n2180 gnd.n1244 240.244
R6395 gnd.n2180 gnd.n847 240.244
R6396 gnd.n2176 gnd.n847 240.244
R6397 gnd.n2176 gnd.n858 240.244
R6398 gnd.n2222 gnd.n858 240.244
R6399 gnd.n2223 gnd.n2222 240.244
R6400 gnd.n2223 gnd.n870 240.244
R6401 gnd.n1665 gnd.n1664 240.244
R6402 gnd.n1736 gnd.n1664 240.244
R6403 gnd.n1734 gnd.n1733 240.244
R6404 gnd.n1730 gnd.n1729 240.244
R6405 gnd.n1726 gnd.n1725 240.244
R6406 gnd.n1722 gnd.n1721 240.244
R6407 gnd.n1718 gnd.n1717 240.244
R6408 gnd.n1714 gnd.n1713 240.244
R6409 gnd.n1710 gnd.n1709 240.244
R6410 gnd.n1706 gnd.n1705 240.244
R6411 gnd.n1702 gnd.n1701 240.244
R6412 gnd.n1698 gnd.n1697 240.244
R6413 gnd.n1694 gnd.n1652 240.244
R6414 gnd.n1754 gnd.n1646 240.244
R6415 gnd.n1754 gnd.n1642 240.244
R6416 gnd.n1760 gnd.n1642 240.244
R6417 gnd.n1760 gnd.n1635 240.244
R6418 gnd.n1770 gnd.n1635 240.244
R6419 gnd.n1770 gnd.n1631 240.244
R6420 gnd.n1776 gnd.n1631 240.244
R6421 gnd.n1776 gnd.n1622 240.244
R6422 gnd.n1816 gnd.n1622 240.244
R6423 gnd.n1816 gnd.n1573 240.244
R6424 gnd.n1824 gnd.n1573 240.244
R6425 gnd.n1824 gnd.n1574 240.244
R6426 gnd.n1574 gnd.n1552 240.244
R6427 gnd.n1845 gnd.n1552 240.244
R6428 gnd.n1845 gnd.n1544 240.244
R6429 gnd.n1856 gnd.n1544 240.244
R6430 gnd.n1856 gnd.n1545 240.244
R6431 gnd.n1545 gnd.n1526 240.244
R6432 gnd.n1876 gnd.n1526 240.244
R6433 gnd.n1876 gnd.n1516 240.244
R6434 gnd.n1886 gnd.n1516 240.244
R6435 gnd.n1886 gnd.n1497 240.244
R6436 gnd.n1907 gnd.n1497 240.244
R6437 gnd.n1907 gnd.n1499 240.244
R6438 gnd.n1499 gnd.n1480 240.244
R6439 gnd.n1935 gnd.n1480 240.244
R6440 gnd.n1935 gnd.n1422 240.244
R6441 gnd.n1987 gnd.n1422 240.244
R6442 gnd.n1987 gnd.n1423 240.244
R6443 gnd.n1983 gnd.n1423 240.244
R6444 gnd.n1983 gnd.n1429 240.244
R6445 gnd.n1444 gnd.n1429 240.244
R6446 gnd.n1973 gnd.n1444 240.244
R6447 gnd.n1973 gnd.n1445 240.244
R6448 gnd.n1969 gnd.n1445 240.244
R6449 gnd.n1969 gnd.n1451 240.244
R6450 gnd.n1451 gnd.n1350 240.244
R6451 gnd.n2026 gnd.n1350 240.244
R6452 gnd.n2026 gnd.n1343 240.244
R6453 gnd.n2037 gnd.n1343 240.244
R6454 gnd.n2037 gnd.n1336 240.244
R6455 gnd.n2052 gnd.n1336 240.244
R6456 gnd.n2052 gnd.n1337 240.244
R6457 gnd.n1337 gnd.n1315 240.244
R6458 gnd.n2074 gnd.n1315 240.244
R6459 gnd.n2074 gnd.n1316 240.244
R6460 gnd.n1316 gnd.n1295 240.244
R6461 gnd.n2111 gnd.n1295 240.244
R6462 gnd.n2111 gnd.n1288 240.244
R6463 gnd.n2122 gnd.n1288 240.244
R6464 gnd.n2122 gnd.n1281 240.244
R6465 gnd.n2137 gnd.n1281 240.244
R6466 gnd.n2137 gnd.n1282 240.244
R6467 gnd.n1282 gnd.n1259 240.244
R6468 gnd.n2161 gnd.n1259 240.244
R6469 gnd.n2161 gnd.n1261 240.244
R6470 gnd.n1261 gnd.n1242 240.244
R6471 gnd.n2202 gnd.n1242 240.244
R6472 gnd.n2202 gnd.n849 240.244
R6473 gnd.n6152 gnd.n849 240.244
R6474 gnd.n6152 gnd.n850 240.244
R6475 gnd.n6148 gnd.n850 240.244
R6476 gnd.n6148 gnd.n856 240.244
R6477 gnd.n872 gnd.n856 240.244
R6478 gnd.n6138 gnd.n872 240.244
R6479 gnd.n7118 gnd.n7117 240.244
R6480 gnd.n7123 gnd.n7120 240.244
R6481 gnd.n7126 gnd.n7125 240.244
R6482 gnd.n7131 gnd.n7128 240.244
R6483 gnd.n7134 gnd.n7133 240.244
R6484 gnd.n7139 gnd.n7136 240.244
R6485 gnd.n7142 gnd.n7141 240.244
R6486 gnd.n7147 gnd.n7144 240.244
R6487 gnd.n7153 gnd.n7149 240.244
R6488 gnd.n2955 gnd.n2773 240.244
R6489 gnd.n5434 gnd.n2955 240.244
R6490 gnd.n5434 gnd.n2903 240.244
R6491 gnd.n2903 gnd.n2890 240.244
R6492 gnd.n5458 gnd.n2890 240.244
R6493 gnd.n5458 gnd.n2885 240.244
R6494 gnd.n5465 gnd.n2885 240.244
R6495 gnd.n5465 gnd.n2874 240.244
R6496 gnd.n2874 gnd.n2862 240.244
R6497 gnd.n5489 gnd.n2862 240.244
R6498 gnd.n5489 gnd.n2857 240.244
R6499 gnd.n5501 gnd.n2857 240.244
R6500 gnd.n5501 gnd.n2846 240.244
R6501 gnd.n5494 gnd.n2846 240.244
R6502 gnd.n5494 gnd.n2836 240.244
R6503 gnd.n2836 gnd.n2823 240.244
R6504 gnd.n5558 gnd.n2823 240.244
R6505 gnd.n5558 gnd.n2812 240.244
R6506 gnd.n2828 gnd.n2812 240.244
R6507 gnd.n2828 gnd.n2803 240.244
R6508 gnd.n5549 gnd.n2803 240.244
R6509 gnd.n5549 gnd.n274 240.244
R6510 gnd.n6940 gnd.n274 240.244
R6511 gnd.n6940 gnd.n303 240.244
R6512 gnd.n6946 gnd.n303 240.244
R6513 gnd.n6946 gnd.n298 240.244
R6514 gnd.n298 gnd.n66 240.244
R6515 gnd.n67 gnd.n66 240.244
R6516 gnd.n68 gnd.n67 240.244
R6517 gnd.n7010 gnd.n68 240.244
R6518 gnd.n7010 gnd.n71 240.244
R6519 gnd.n72 gnd.n71 240.244
R6520 gnd.n73 gnd.n72 240.244
R6521 gnd.n243 gnd.n73 240.244
R6522 gnd.n243 gnd.n76 240.244
R6523 gnd.n77 gnd.n76 240.244
R6524 gnd.n78 gnd.n77 240.244
R6525 gnd.n236 gnd.n78 240.244
R6526 gnd.n236 gnd.n81 240.244
R6527 gnd.n82 gnd.n81 240.244
R6528 gnd.n83 gnd.n82 240.244
R6529 gnd.n213 gnd.n83 240.244
R6530 gnd.n213 gnd.n86 240.244
R6531 gnd.n87 gnd.n86 240.244
R6532 gnd.n88 gnd.n87 240.244
R6533 gnd.n206 gnd.n88 240.244
R6534 gnd.n206 gnd.n91 240.244
R6535 gnd.n92 gnd.n91 240.244
R6536 gnd.n93 gnd.n92 240.244
R6537 gnd.n180 gnd.n93 240.244
R6538 gnd.n180 gnd.n96 240.244
R6539 gnd.n97 gnd.n96 240.244
R6540 gnd.n7281 gnd.n97 240.244
R6541 gnd.n3007 gnd.n3006 240.244
R6542 gnd.n2998 gnd.n2997 240.244
R6543 gnd.n3023 gnd.n3022 240.244
R6544 gnd.n2989 gnd.n2988 240.244
R6545 gnd.n3040 gnd.n3039 240.244
R6546 gnd.n2980 gnd.n2979 240.244
R6547 gnd.n3057 gnd.n3056 240.244
R6548 gnd.n2971 gnd.n2970 240.244
R6549 gnd.n2966 gnd.n2720 240.244
R6550 gnd.n5621 gnd.n2776 240.244
R6551 gnd.n2780 gnd.n2776 240.244
R6552 gnd.n2781 gnd.n2780 240.244
R6553 gnd.n2782 gnd.n2781 240.244
R6554 gnd.n2894 gnd.n2782 240.244
R6555 gnd.n2894 gnd.n2785 240.244
R6556 gnd.n2786 gnd.n2785 240.244
R6557 gnd.n2787 gnd.n2786 240.244
R6558 gnd.n2875 gnd.n2787 240.244
R6559 gnd.n2875 gnd.n2790 240.244
R6560 gnd.n2791 gnd.n2790 240.244
R6561 gnd.n2792 gnd.n2791 240.244
R6562 gnd.n5514 gnd.n2792 240.244
R6563 gnd.n5514 gnd.n2795 240.244
R6564 gnd.n2796 gnd.n2795 240.244
R6565 gnd.n2797 gnd.n2796 240.244
R6566 gnd.n5559 gnd.n2797 240.244
R6567 gnd.n5559 gnd.n2800 240.244
R6568 gnd.n2801 gnd.n2800 240.244
R6569 gnd.n5588 gnd.n2801 240.244
R6570 gnd.n5588 gnd.n276 240.244
R6571 gnd.n7037 gnd.n276 240.244
R6572 gnd.n7037 gnd.n277 240.244
R6573 gnd.n282 gnd.n277 240.244
R6574 gnd.n283 gnd.n282 240.244
R6575 gnd.n284 gnd.n283 240.244
R6576 gnd.n6928 gnd.n284 240.244
R6577 gnd.n6928 gnd.n288 240.244
R6578 gnd.n7023 gnd.n288 240.244
R6579 gnd.n7023 gnd.n257 240.244
R6580 gnd.n7046 gnd.n257 240.244
R6581 gnd.n7046 gnd.n253 240.244
R6582 gnd.n7052 gnd.n253 240.244
R6583 gnd.n7052 gnd.n242 240.244
R6584 gnd.n7062 gnd.n242 240.244
R6585 gnd.n7062 gnd.n238 240.244
R6586 gnd.n7068 gnd.n238 240.244
R6587 gnd.n7068 gnd.n227 240.244
R6588 gnd.n7078 gnd.n227 240.244
R6589 gnd.n7078 gnd.n223 240.244
R6590 gnd.n7084 gnd.n223 240.244
R6591 gnd.n7084 gnd.n212 240.244
R6592 gnd.n7094 gnd.n212 240.244
R6593 gnd.n7094 gnd.n208 240.244
R6594 gnd.n7100 gnd.n208 240.244
R6595 gnd.n7100 gnd.n197 240.244
R6596 gnd.n7110 gnd.n197 240.244
R6597 gnd.n7110 gnd.n191 240.244
R6598 gnd.n7191 gnd.n191 240.244
R6599 gnd.n7191 gnd.n192 240.244
R6600 gnd.n192 gnd.n182 240.244
R6601 gnd.n7115 gnd.n182 240.244
R6602 gnd.n7115 gnd.n103 240.244
R6603 gnd.n3504 gnd.n2573 240.244
R6604 gnd.n3508 gnd.n3507 240.244
R6605 gnd.n3520 gnd.n3519 240.244
R6606 gnd.n3532 gnd.n3531 240.244
R6607 gnd.n3494 gnd.n3493 240.244
R6608 gnd.n3544 gnd.n3543 240.244
R6609 gnd.n3556 gnd.n3555 240.244
R6610 gnd.n3569 gnd.n3480 240.244
R6611 gnd.n3570 gnd.n3471 240.244
R6612 gnd.n3882 gnd.n3802 240.244
R6613 gnd.n3883 gnd.n3882 240.244
R6614 gnd.n3883 gnd.n2314 240.244
R6615 gnd.n3888 gnd.n2314 240.244
R6616 gnd.n3888 gnd.n2326 240.244
R6617 gnd.n3891 gnd.n2326 240.244
R6618 gnd.n3891 gnd.n2337 240.244
R6619 gnd.n3896 gnd.n2337 240.244
R6620 gnd.n3896 gnd.n2347 240.244
R6621 gnd.n3899 gnd.n2347 240.244
R6622 gnd.n3899 gnd.n2357 240.244
R6623 gnd.n3904 gnd.n2357 240.244
R6624 gnd.n3904 gnd.n2367 240.244
R6625 gnd.n3907 gnd.n2367 240.244
R6626 gnd.n3907 gnd.n2377 240.244
R6627 gnd.n3912 gnd.n2377 240.244
R6628 gnd.n3912 gnd.n2387 240.244
R6629 gnd.n3915 gnd.n2387 240.244
R6630 gnd.n3915 gnd.n2397 240.244
R6631 gnd.n3920 gnd.n2397 240.244
R6632 gnd.n3920 gnd.n2407 240.244
R6633 gnd.n3969 gnd.n2407 240.244
R6634 gnd.n3969 gnd.n2417 240.244
R6635 gnd.n3975 gnd.n2417 240.244
R6636 gnd.n3975 gnd.n2426 240.244
R6637 gnd.n3987 gnd.n2426 240.244
R6638 gnd.n3987 gnd.n2436 240.244
R6639 gnd.n3994 gnd.n2436 240.244
R6640 gnd.n3994 gnd.n2444 240.244
R6641 gnd.n4004 gnd.n2444 240.244
R6642 gnd.n4004 gnd.n2455 240.244
R6643 gnd.n4010 gnd.n2455 240.244
R6644 gnd.n4010 gnd.n2465 240.244
R6645 gnd.n4020 gnd.n2465 240.244
R6646 gnd.n4020 gnd.n2475 240.244
R6647 gnd.n4026 gnd.n2475 240.244
R6648 gnd.n4026 gnd.n2486 240.244
R6649 gnd.n4036 gnd.n2486 240.244
R6650 gnd.n4036 gnd.n2497 240.244
R6651 gnd.n4042 gnd.n2497 240.244
R6652 gnd.n4042 gnd.n2508 240.244
R6653 gnd.n4052 gnd.n2508 240.244
R6654 gnd.n4052 gnd.n2518 240.244
R6655 gnd.n4058 gnd.n2518 240.244
R6656 gnd.n4058 gnd.n2529 240.244
R6657 gnd.n4068 gnd.n2529 240.244
R6658 gnd.n4068 gnd.n2540 240.244
R6659 gnd.n4074 gnd.n2540 240.244
R6660 gnd.n4074 gnd.n2551 240.244
R6661 gnd.n4085 gnd.n2551 240.244
R6662 gnd.n4085 gnd.n2562 240.244
R6663 gnd.n4091 gnd.n2562 240.244
R6664 gnd.n4091 gnd.n2571 240.244
R6665 gnd.n3862 gnd.n3861 240.244
R6666 gnd.n3858 gnd.n3857 240.244
R6667 gnd.n3854 gnd.n3853 240.244
R6668 gnd.n3850 gnd.n3849 240.244
R6669 gnd.n3846 gnd.n3845 240.244
R6670 gnd.n3842 gnd.n3841 240.244
R6671 gnd.n3838 gnd.n3837 240.244
R6672 gnd.n3834 gnd.n3833 240.244
R6673 gnd.n3822 gnd.n2258 240.244
R6674 gnd.n3874 gnd.n3803 240.244
R6675 gnd.n3874 gnd.n3804 240.244
R6676 gnd.n3804 gnd.n2316 240.244
R6677 gnd.n2328 gnd.n2316 240.244
R6678 gnd.n5982 gnd.n2328 240.244
R6679 gnd.n5982 gnd.n2329 240.244
R6680 gnd.n5978 gnd.n2329 240.244
R6681 gnd.n5978 gnd.n2335 240.244
R6682 gnd.n5970 gnd.n2335 240.244
R6683 gnd.n5970 gnd.n2348 240.244
R6684 gnd.n5966 gnd.n2348 240.244
R6685 gnd.n5966 gnd.n2354 240.244
R6686 gnd.n5958 gnd.n2354 240.244
R6687 gnd.n5958 gnd.n2369 240.244
R6688 gnd.n5954 gnd.n2369 240.244
R6689 gnd.n5954 gnd.n2375 240.244
R6690 gnd.n5946 gnd.n2375 240.244
R6691 gnd.n5946 gnd.n2388 240.244
R6692 gnd.n5942 gnd.n2388 240.244
R6693 gnd.n5942 gnd.n2394 240.244
R6694 gnd.n5934 gnd.n2394 240.244
R6695 gnd.n5934 gnd.n2409 240.244
R6696 gnd.n5930 gnd.n2409 240.244
R6697 gnd.n5930 gnd.n2415 240.244
R6698 gnd.n5922 gnd.n2415 240.244
R6699 gnd.n5922 gnd.n2427 240.244
R6700 gnd.n5918 gnd.n2427 240.244
R6701 gnd.n5918 gnd.n2433 240.244
R6702 gnd.n5909 gnd.n2433 240.244
R6703 gnd.n5909 gnd.n2446 240.244
R6704 gnd.n5905 gnd.n2446 240.244
R6705 gnd.n5905 gnd.n2452 240.244
R6706 gnd.n5897 gnd.n2452 240.244
R6707 gnd.n5897 gnd.n2466 240.244
R6708 gnd.n5893 gnd.n2466 240.244
R6709 gnd.n5893 gnd.n2472 240.244
R6710 gnd.n5885 gnd.n2472 240.244
R6711 gnd.n5885 gnd.n2488 240.244
R6712 gnd.n5881 gnd.n2488 240.244
R6713 gnd.n5881 gnd.n2494 240.244
R6714 gnd.n5873 gnd.n2494 240.244
R6715 gnd.n5873 gnd.n2509 240.244
R6716 gnd.n5869 gnd.n2509 240.244
R6717 gnd.n5869 gnd.n2515 240.244
R6718 gnd.n5861 gnd.n2515 240.244
R6719 gnd.n5861 gnd.n2531 240.244
R6720 gnd.n5857 gnd.n2531 240.244
R6721 gnd.n5857 gnd.n2537 240.244
R6722 gnd.n5849 gnd.n2537 240.244
R6723 gnd.n5849 gnd.n2553 240.244
R6724 gnd.n5845 gnd.n2553 240.244
R6725 gnd.n5845 gnd.n2559 240.244
R6726 gnd.n5837 gnd.n2559 240.244
R6727 gnd.n6325 gnd.n678 240.244
R6728 gnd.n6325 gnd.n674 240.244
R6729 gnd.n6331 gnd.n674 240.244
R6730 gnd.n6331 gnd.n672 240.244
R6731 gnd.n6335 gnd.n672 240.244
R6732 gnd.n6335 gnd.n668 240.244
R6733 gnd.n6341 gnd.n668 240.244
R6734 gnd.n6341 gnd.n666 240.244
R6735 gnd.n6345 gnd.n666 240.244
R6736 gnd.n6345 gnd.n662 240.244
R6737 gnd.n6351 gnd.n662 240.244
R6738 gnd.n6351 gnd.n660 240.244
R6739 gnd.n6355 gnd.n660 240.244
R6740 gnd.n6355 gnd.n656 240.244
R6741 gnd.n6361 gnd.n656 240.244
R6742 gnd.n6361 gnd.n654 240.244
R6743 gnd.n6365 gnd.n654 240.244
R6744 gnd.n6365 gnd.n650 240.244
R6745 gnd.n6371 gnd.n650 240.244
R6746 gnd.n6371 gnd.n648 240.244
R6747 gnd.n6375 gnd.n648 240.244
R6748 gnd.n6375 gnd.n644 240.244
R6749 gnd.n6381 gnd.n644 240.244
R6750 gnd.n6381 gnd.n642 240.244
R6751 gnd.n6385 gnd.n642 240.244
R6752 gnd.n6385 gnd.n638 240.244
R6753 gnd.n6391 gnd.n638 240.244
R6754 gnd.n6391 gnd.n636 240.244
R6755 gnd.n6395 gnd.n636 240.244
R6756 gnd.n6395 gnd.n632 240.244
R6757 gnd.n6401 gnd.n632 240.244
R6758 gnd.n6401 gnd.n630 240.244
R6759 gnd.n6405 gnd.n630 240.244
R6760 gnd.n6405 gnd.n626 240.244
R6761 gnd.n6411 gnd.n626 240.244
R6762 gnd.n6411 gnd.n624 240.244
R6763 gnd.n6415 gnd.n624 240.244
R6764 gnd.n6415 gnd.n620 240.244
R6765 gnd.n6421 gnd.n620 240.244
R6766 gnd.n6421 gnd.n618 240.244
R6767 gnd.n6425 gnd.n618 240.244
R6768 gnd.n6425 gnd.n614 240.244
R6769 gnd.n6431 gnd.n614 240.244
R6770 gnd.n6431 gnd.n612 240.244
R6771 gnd.n6435 gnd.n612 240.244
R6772 gnd.n6435 gnd.n608 240.244
R6773 gnd.n6441 gnd.n608 240.244
R6774 gnd.n6441 gnd.n606 240.244
R6775 gnd.n6445 gnd.n606 240.244
R6776 gnd.n6445 gnd.n602 240.244
R6777 gnd.n6451 gnd.n602 240.244
R6778 gnd.n6451 gnd.n600 240.244
R6779 gnd.n6455 gnd.n600 240.244
R6780 gnd.n6455 gnd.n596 240.244
R6781 gnd.n6461 gnd.n596 240.244
R6782 gnd.n6461 gnd.n594 240.244
R6783 gnd.n6465 gnd.n594 240.244
R6784 gnd.n6465 gnd.n590 240.244
R6785 gnd.n6471 gnd.n590 240.244
R6786 gnd.n6471 gnd.n588 240.244
R6787 gnd.n6475 gnd.n588 240.244
R6788 gnd.n6475 gnd.n584 240.244
R6789 gnd.n6481 gnd.n584 240.244
R6790 gnd.n6481 gnd.n582 240.244
R6791 gnd.n6485 gnd.n582 240.244
R6792 gnd.n6485 gnd.n578 240.244
R6793 gnd.n6491 gnd.n578 240.244
R6794 gnd.n6491 gnd.n576 240.244
R6795 gnd.n6495 gnd.n576 240.244
R6796 gnd.n6495 gnd.n572 240.244
R6797 gnd.n6501 gnd.n572 240.244
R6798 gnd.n6501 gnd.n570 240.244
R6799 gnd.n6505 gnd.n570 240.244
R6800 gnd.n6505 gnd.n566 240.244
R6801 gnd.n6511 gnd.n566 240.244
R6802 gnd.n6511 gnd.n564 240.244
R6803 gnd.n6515 gnd.n564 240.244
R6804 gnd.n6515 gnd.n560 240.244
R6805 gnd.n6521 gnd.n560 240.244
R6806 gnd.n6521 gnd.n558 240.244
R6807 gnd.n6525 gnd.n558 240.244
R6808 gnd.n6525 gnd.n554 240.244
R6809 gnd.n6531 gnd.n554 240.244
R6810 gnd.n6531 gnd.n552 240.244
R6811 gnd.n6535 gnd.n552 240.244
R6812 gnd.n6535 gnd.n548 240.244
R6813 gnd.n6541 gnd.n548 240.244
R6814 gnd.n6541 gnd.n546 240.244
R6815 gnd.n6545 gnd.n546 240.244
R6816 gnd.n6545 gnd.n542 240.244
R6817 gnd.n6551 gnd.n542 240.244
R6818 gnd.n6551 gnd.n540 240.244
R6819 gnd.n6555 gnd.n540 240.244
R6820 gnd.n6555 gnd.n536 240.244
R6821 gnd.n6561 gnd.n536 240.244
R6822 gnd.n6561 gnd.n534 240.244
R6823 gnd.n6565 gnd.n534 240.244
R6824 gnd.n6565 gnd.n530 240.244
R6825 gnd.n6571 gnd.n530 240.244
R6826 gnd.n6571 gnd.n528 240.244
R6827 gnd.n6575 gnd.n528 240.244
R6828 gnd.n6575 gnd.n524 240.244
R6829 gnd.n6581 gnd.n524 240.244
R6830 gnd.n6581 gnd.n522 240.244
R6831 gnd.n6585 gnd.n522 240.244
R6832 gnd.n6585 gnd.n518 240.244
R6833 gnd.n6591 gnd.n518 240.244
R6834 gnd.n6591 gnd.n516 240.244
R6835 gnd.n6595 gnd.n516 240.244
R6836 gnd.n6595 gnd.n512 240.244
R6837 gnd.n6601 gnd.n512 240.244
R6838 gnd.n6601 gnd.n510 240.244
R6839 gnd.n6605 gnd.n510 240.244
R6840 gnd.n6605 gnd.n506 240.244
R6841 gnd.n6611 gnd.n506 240.244
R6842 gnd.n6611 gnd.n504 240.244
R6843 gnd.n6615 gnd.n504 240.244
R6844 gnd.n6615 gnd.n500 240.244
R6845 gnd.n6621 gnd.n500 240.244
R6846 gnd.n6621 gnd.n498 240.244
R6847 gnd.n6625 gnd.n498 240.244
R6848 gnd.n6625 gnd.n494 240.244
R6849 gnd.n6631 gnd.n494 240.244
R6850 gnd.n6631 gnd.n492 240.244
R6851 gnd.n6635 gnd.n492 240.244
R6852 gnd.n6635 gnd.n488 240.244
R6853 gnd.n6641 gnd.n488 240.244
R6854 gnd.n6641 gnd.n486 240.244
R6855 gnd.n6645 gnd.n486 240.244
R6856 gnd.n6645 gnd.n482 240.244
R6857 gnd.n6651 gnd.n482 240.244
R6858 gnd.n6651 gnd.n480 240.244
R6859 gnd.n6655 gnd.n480 240.244
R6860 gnd.n6655 gnd.n476 240.244
R6861 gnd.n6661 gnd.n476 240.244
R6862 gnd.n6661 gnd.n474 240.244
R6863 gnd.n6665 gnd.n474 240.244
R6864 gnd.n6665 gnd.n470 240.244
R6865 gnd.n6671 gnd.n470 240.244
R6866 gnd.n6671 gnd.n468 240.244
R6867 gnd.n6675 gnd.n468 240.244
R6868 gnd.n6675 gnd.n464 240.244
R6869 gnd.n6681 gnd.n464 240.244
R6870 gnd.n6681 gnd.n462 240.244
R6871 gnd.n6685 gnd.n462 240.244
R6872 gnd.n6685 gnd.n458 240.244
R6873 gnd.n6691 gnd.n458 240.244
R6874 gnd.n6691 gnd.n456 240.244
R6875 gnd.n6695 gnd.n456 240.244
R6876 gnd.n6695 gnd.n452 240.244
R6877 gnd.n6702 gnd.n452 240.244
R6878 gnd.n6702 gnd.n450 240.244
R6879 gnd.n6706 gnd.n450 240.244
R6880 gnd.n6706 gnd.n447 240.244
R6881 gnd.n6712 gnd.n445 240.244
R6882 gnd.n6716 gnd.n445 240.244
R6883 gnd.n6716 gnd.n441 240.244
R6884 gnd.n6722 gnd.n441 240.244
R6885 gnd.n6722 gnd.n439 240.244
R6886 gnd.n6726 gnd.n439 240.244
R6887 gnd.n6726 gnd.n435 240.244
R6888 gnd.n6732 gnd.n435 240.244
R6889 gnd.n6732 gnd.n433 240.244
R6890 gnd.n6736 gnd.n433 240.244
R6891 gnd.n6736 gnd.n429 240.244
R6892 gnd.n6742 gnd.n429 240.244
R6893 gnd.n6742 gnd.n427 240.244
R6894 gnd.n6746 gnd.n427 240.244
R6895 gnd.n6746 gnd.n423 240.244
R6896 gnd.n6752 gnd.n423 240.244
R6897 gnd.n6752 gnd.n421 240.244
R6898 gnd.n6756 gnd.n421 240.244
R6899 gnd.n6756 gnd.n417 240.244
R6900 gnd.n6762 gnd.n417 240.244
R6901 gnd.n6762 gnd.n415 240.244
R6902 gnd.n6766 gnd.n415 240.244
R6903 gnd.n6766 gnd.n411 240.244
R6904 gnd.n6772 gnd.n411 240.244
R6905 gnd.n6772 gnd.n409 240.244
R6906 gnd.n6776 gnd.n409 240.244
R6907 gnd.n6776 gnd.n405 240.244
R6908 gnd.n6782 gnd.n405 240.244
R6909 gnd.n6782 gnd.n403 240.244
R6910 gnd.n6786 gnd.n403 240.244
R6911 gnd.n6786 gnd.n399 240.244
R6912 gnd.n6792 gnd.n399 240.244
R6913 gnd.n6792 gnd.n397 240.244
R6914 gnd.n6796 gnd.n397 240.244
R6915 gnd.n6796 gnd.n393 240.244
R6916 gnd.n6802 gnd.n393 240.244
R6917 gnd.n6802 gnd.n391 240.244
R6918 gnd.n6806 gnd.n391 240.244
R6919 gnd.n6806 gnd.n387 240.244
R6920 gnd.n6812 gnd.n387 240.244
R6921 gnd.n6812 gnd.n385 240.244
R6922 gnd.n6816 gnd.n385 240.244
R6923 gnd.n6816 gnd.n381 240.244
R6924 gnd.n6822 gnd.n381 240.244
R6925 gnd.n6822 gnd.n379 240.244
R6926 gnd.n6826 gnd.n379 240.244
R6927 gnd.n6826 gnd.n375 240.244
R6928 gnd.n6832 gnd.n375 240.244
R6929 gnd.n6832 gnd.n373 240.244
R6930 gnd.n6836 gnd.n373 240.244
R6931 gnd.n6836 gnd.n369 240.244
R6932 gnd.n6842 gnd.n369 240.244
R6933 gnd.n6842 gnd.n367 240.244
R6934 gnd.n6846 gnd.n367 240.244
R6935 gnd.n6846 gnd.n363 240.244
R6936 gnd.n6852 gnd.n363 240.244
R6937 gnd.n6852 gnd.n361 240.244
R6938 gnd.n6856 gnd.n361 240.244
R6939 gnd.n6856 gnd.n357 240.244
R6940 gnd.n6862 gnd.n357 240.244
R6941 gnd.n6862 gnd.n355 240.244
R6942 gnd.n6866 gnd.n355 240.244
R6943 gnd.n6866 gnd.n351 240.244
R6944 gnd.n6872 gnd.n351 240.244
R6945 gnd.n6872 gnd.n349 240.244
R6946 gnd.n6876 gnd.n349 240.244
R6947 gnd.n6876 gnd.n345 240.244
R6948 gnd.n6882 gnd.n345 240.244
R6949 gnd.n6882 gnd.n343 240.244
R6950 gnd.n6886 gnd.n343 240.244
R6951 gnd.n6886 gnd.n339 240.244
R6952 gnd.n6892 gnd.n339 240.244
R6953 gnd.n6892 gnd.n337 240.244
R6954 gnd.n6896 gnd.n337 240.244
R6955 gnd.n6896 gnd.n333 240.244
R6956 gnd.n6902 gnd.n333 240.244
R6957 gnd.n6902 gnd.n331 240.244
R6958 gnd.n6906 gnd.n331 240.244
R6959 gnd.n6906 gnd.n327 240.244
R6960 gnd.n6912 gnd.n327 240.244
R6961 gnd.n6912 gnd.n325 240.244
R6962 gnd.n6917 gnd.n325 240.244
R6963 gnd.n6917 gnd.n321 240.244
R6964 gnd.n6923 gnd.n321 240.244
R6965 gnd.n3688 gnd.n3681 240.244
R6966 gnd.n3784 gnd.n3681 240.244
R6967 gnd.n3784 gnd.n3682 240.244
R6968 gnd.n3780 gnd.n3682 240.244
R6969 gnd.n3780 gnd.n3779 240.244
R6970 gnd.n3779 gnd.n3778 240.244
R6971 gnd.n3778 gnd.n3697 240.244
R6972 gnd.n3774 gnd.n3697 240.244
R6973 gnd.n3774 gnd.n3773 240.244
R6974 gnd.n3773 gnd.n3772 240.244
R6975 gnd.n3772 gnd.n3703 240.244
R6976 gnd.n3768 gnd.n3703 240.244
R6977 gnd.n3768 gnd.n3767 240.244
R6978 gnd.n3767 gnd.n3766 240.244
R6979 gnd.n3766 gnd.n3709 240.244
R6980 gnd.n3762 gnd.n3709 240.244
R6981 gnd.n3762 gnd.n3761 240.244
R6982 gnd.n3761 gnd.n3760 240.244
R6983 gnd.n3760 gnd.n3715 240.244
R6984 gnd.n3756 gnd.n3715 240.244
R6985 gnd.n3756 gnd.n3755 240.244
R6986 gnd.n3755 gnd.n3754 240.244
R6987 gnd.n3754 gnd.n3721 240.244
R6988 gnd.n3750 gnd.n3721 240.244
R6989 gnd.n3750 gnd.n3749 240.244
R6990 gnd.n3749 gnd.n3748 240.244
R6991 gnd.n3748 gnd.n3727 240.244
R6992 gnd.n3744 gnd.n3727 240.244
R6993 gnd.n3744 gnd.n3743 240.244
R6994 gnd.n3743 gnd.n3742 240.244
R6995 gnd.n3742 gnd.n3733 240.244
R6996 gnd.n3738 gnd.n3733 240.244
R6997 gnd.n3738 gnd.n3438 240.244
R6998 gnd.n4416 gnd.n3438 240.244
R6999 gnd.n4416 gnd.n3434 240.244
R7000 gnd.n4422 gnd.n3434 240.244
R7001 gnd.n4422 gnd.n3424 240.244
R7002 gnd.n4432 gnd.n3424 240.244
R7003 gnd.n4432 gnd.n3419 240.244
R7004 gnd.n4440 gnd.n3419 240.244
R7005 gnd.n4440 gnd.n3420 240.244
R7006 gnd.n3420 gnd.n3392 240.244
R7007 gnd.n4556 gnd.n3392 240.244
R7008 gnd.n4556 gnd.n3388 240.244
R7009 gnd.n4562 gnd.n3388 240.244
R7010 gnd.n4562 gnd.n3378 240.244
R7011 gnd.n4572 gnd.n3378 240.244
R7012 gnd.n4572 gnd.n3374 240.244
R7013 gnd.n4578 gnd.n3374 240.244
R7014 gnd.n4578 gnd.n3363 240.244
R7015 gnd.n4588 gnd.n3363 240.244
R7016 gnd.n4588 gnd.n3359 240.244
R7017 gnd.n4594 gnd.n3359 240.244
R7018 gnd.n4594 gnd.n3349 240.244
R7019 gnd.n4603 gnd.n3349 240.244
R7020 gnd.n4603 gnd.n3344 240.244
R7021 gnd.n4611 gnd.n3344 240.244
R7022 gnd.n4611 gnd.n3345 240.244
R7023 gnd.n3345 gnd.n3317 240.244
R7024 gnd.n4729 gnd.n3317 240.244
R7025 gnd.n4729 gnd.n3313 240.244
R7026 gnd.n4735 gnd.n3313 240.244
R7027 gnd.n4735 gnd.n3303 240.244
R7028 gnd.n4745 gnd.n3303 240.244
R7029 gnd.n4745 gnd.n3299 240.244
R7030 gnd.n4751 gnd.n3299 240.244
R7031 gnd.n4751 gnd.n3290 240.244
R7032 gnd.n4761 gnd.n3290 240.244
R7033 gnd.n4761 gnd.n3286 240.244
R7034 gnd.n4767 gnd.n3286 240.244
R7035 gnd.n4767 gnd.n3279 240.244
R7036 gnd.n4777 gnd.n3279 240.244
R7037 gnd.n4777 gnd.n3274 240.244
R7038 gnd.n4785 gnd.n3274 240.244
R7039 gnd.n4785 gnd.n3275 240.244
R7040 gnd.n3275 gnd.n3246 240.244
R7041 gnd.n4900 gnd.n3246 240.244
R7042 gnd.n4900 gnd.n3242 240.244
R7043 gnd.n4906 gnd.n3242 240.244
R7044 gnd.n4906 gnd.n3231 240.244
R7045 gnd.n4916 gnd.n3231 240.244
R7046 gnd.n4916 gnd.n3227 240.244
R7047 gnd.n4922 gnd.n3227 240.244
R7048 gnd.n4922 gnd.n3216 240.244
R7049 gnd.n4932 gnd.n3216 240.244
R7050 gnd.n4932 gnd.n3212 240.244
R7051 gnd.n4938 gnd.n3212 240.244
R7052 gnd.n4938 gnd.n3203 240.244
R7053 gnd.n4948 gnd.n3203 240.244
R7054 gnd.n4948 gnd.n3198 240.244
R7055 gnd.n4956 gnd.n3198 240.244
R7056 gnd.n4956 gnd.n3199 240.244
R7057 gnd.n3199 gnd.n3171 240.244
R7058 gnd.n5306 gnd.n3171 240.244
R7059 gnd.n5306 gnd.n3167 240.244
R7060 gnd.n5312 gnd.n3167 240.244
R7061 gnd.n5312 gnd.n3158 240.244
R7062 gnd.n5322 gnd.n3158 240.244
R7063 gnd.n5322 gnd.n3154 240.244
R7064 gnd.n5328 gnd.n3154 240.244
R7065 gnd.n5328 gnd.n3144 240.244
R7066 gnd.n5338 gnd.n3144 240.244
R7067 gnd.n5338 gnd.n3140 240.244
R7068 gnd.n5344 gnd.n3140 240.244
R7069 gnd.n5344 gnd.n3131 240.244
R7070 gnd.n5354 gnd.n3131 240.244
R7071 gnd.n5354 gnd.n3127 240.244
R7072 gnd.n5360 gnd.n3127 240.244
R7073 gnd.n5360 gnd.n3117 240.244
R7074 gnd.n5370 gnd.n3117 240.244
R7075 gnd.n5370 gnd.n3113 240.244
R7076 gnd.n5376 gnd.n3113 240.244
R7077 gnd.n5376 gnd.n3103 240.244
R7078 gnd.n5388 gnd.n3103 240.244
R7079 gnd.n5388 gnd.n3098 240.244
R7080 gnd.n5397 gnd.n3098 240.244
R7081 gnd.n5397 gnd.n3099 240.244
R7082 gnd.n3099 gnd.n2683 240.244
R7083 gnd.n5705 gnd.n2683 240.244
R7084 gnd.n5705 gnd.n2686 240.244
R7085 gnd.n5701 gnd.n2686 240.244
R7086 gnd.n5701 gnd.n2692 240.244
R7087 gnd.n2910 gnd.n2692 240.244
R7088 gnd.n2916 gnd.n2910 240.244
R7089 gnd.n2917 gnd.n2916 240.244
R7090 gnd.n5437 gnd.n2917 240.244
R7091 gnd.n5437 gnd.n2905 240.244
R7092 gnd.n5445 gnd.n2905 240.244
R7093 gnd.n5445 gnd.n2906 240.244
R7094 gnd.n2906 gnd.n2882 240.244
R7095 gnd.n5468 gnd.n2882 240.244
R7096 gnd.n5468 gnd.n2877 240.244
R7097 gnd.n5476 gnd.n2877 240.244
R7098 gnd.n5476 gnd.n2878 240.244
R7099 gnd.n2878 gnd.n2854 240.244
R7100 gnd.n5504 gnd.n2854 240.244
R7101 gnd.n5504 gnd.n2848 240.244
R7102 gnd.n5512 gnd.n2848 240.244
R7103 gnd.n5512 gnd.n2850 240.244
R7104 gnd.n2850 gnd.n2820 240.244
R7105 gnd.n5562 gnd.n2820 240.244
R7106 gnd.n5562 gnd.n2814 240.244
R7107 gnd.n5577 gnd.n2814 240.244
R7108 gnd.n5577 gnd.n2816 240.244
R7109 gnd.n5573 gnd.n2816 240.244
R7110 gnd.n5573 gnd.n5572 240.244
R7111 gnd.n5572 gnd.n309 240.244
R7112 gnd.n6937 gnd.n309 240.244
R7113 gnd.n6937 gnd.n310 240.244
R7114 gnd.n6933 gnd.n310 240.244
R7115 gnd.n6933 gnd.n6932 240.244
R7116 gnd.n6932 gnd.n6931 240.244
R7117 gnd.n6931 gnd.n317 240.244
R7118 gnd.n6924 gnd.n317 240.244
R7119 gnd.n6321 gnd.n680 240.244
R7120 gnd.n6317 gnd.n680 240.244
R7121 gnd.n6317 gnd.n685 240.244
R7122 gnd.n6313 gnd.n685 240.244
R7123 gnd.n6313 gnd.n687 240.244
R7124 gnd.n6309 gnd.n687 240.244
R7125 gnd.n6309 gnd.n693 240.244
R7126 gnd.n6305 gnd.n693 240.244
R7127 gnd.n6305 gnd.n695 240.244
R7128 gnd.n6301 gnd.n695 240.244
R7129 gnd.n6301 gnd.n701 240.244
R7130 gnd.n6297 gnd.n701 240.244
R7131 gnd.n6297 gnd.n703 240.244
R7132 gnd.n6293 gnd.n703 240.244
R7133 gnd.n6293 gnd.n709 240.244
R7134 gnd.n6289 gnd.n709 240.244
R7135 gnd.n6289 gnd.n711 240.244
R7136 gnd.n6285 gnd.n711 240.244
R7137 gnd.n6285 gnd.n717 240.244
R7138 gnd.n6281 gnd.n717 240.244
R7139 gnd.n6281 gnd.n719 240.244
R7140 gnd.n6277 gnd.n719 240.244
R7141 gnd.n6277 gnd.n725 240.244
R7142 gnd.n6273 gnd.n725 240.244
R7143 gnd.n6273 gnd.n727 240.244
R7144 gnd.n6269 gnd.n727 240.244
R7145 gnd.n6269 gnd.n733 240.244
R7146 gnd.n6265 gnd.n733 240.244
R7147 gnd.n6265 gnd.n735 240.244
R7148 gnd.n6261 gnd.n735 240.244
R7149 gnd.n6261 gnd.n741 240.244
R7150 gnd.n6257 gnd.n741 240.244
R7151 gnd.n6257 gnd.n743 240.244
R7152 gnd.n6253 gnd.n743 240.244
R7153 gnd.n6253 gnd.n749 240.244
R7154 gnd.n6249 gnd.n749 240.244
R7155 gnd.n6249 gnd.n751 240.244
R7156 gnd.n6245 gnd.n751 240.244
R7157 gnd.n6245 gnd.n757 240.244
R7158 gnd.n6241 gnd.n757 240.244
R7159 gnd.n6241 gnd.n759 240.244
R7160 gnd.n6237 gnd.n759 240.244
R7161 gnd.n6237 gnd.n765 240.244
R7162 gnd.n6233 gnd.n765 240.244
R7163 gnd.n6233 gnd.n767 240.244
R7164 gnd.n6229 gnd.n767 240.244
R7165 gnd.n6229 gnd.n773 240.244
R7166 gnd.n6225 gnd.n773 240.244
R7167 gnd.n6225 gnd.n775 240.244
R7168 gnd.n6221 gnd.n775 240.244
R7169 gnd.n6221 gnd.n781 240.244
R7170 gnd.n6217 gnd.n781 240.244
R7171 gnd.n6217 gnd.n783 240.244
R7172 gnd.n6213 gnd.n783 240.244
R7173 gnd.n6213 gnd.n789 240.244
R7174 gnd.n6209 gnd.n789 240.244
R7175 gnd.n6209 gnd.n791 240.244
R7176 gnd.n6205 gnd.n791 240.244
R7177 gnd.n6205 gnd.n797 240.244
R7178 gnd.n6201 gnd.n797 240.244
R7179 gnd.n6201 gnd.n799 240.244
R7180 gnd.n6197 gnd.n799 240.244
R7181 gnd.n6197 gnd.n805 240.244
R7182 gnd.n6193 gnd.n805 240.244
R7183 gnd.n6193 gnd.n807 240.244
R7184 gnd.n6189 gnd.n807 240.244
R7185 gnd.n6189 gnd.n813 240.244
R7186 gnd.n6185 gnd.n813 240.244
R7187 gnd.n6185 gnd.n815 240.244
R7188 gnd.n6181 gnd.n815 240.244
R7189 gnd.n6181 gnd.n821 240.244
R7190 gnd.n6177 gnd.n821 240.244
R7191 gnd.n6177 gnd.n823 240.244
R7192 gnd.n6173 gnd.n823 240.244
R7193 gnd.n6173 gnd.n829 240.244
R7194 gnd.n6169 gnd.n829 240.244
R7195 gnd.n6169 gnd.n831 240.244
R7196 gnd.n6165 gnd.n831 240.244
R7197 gnd.n6165 gnd.n837 240.244
R7198 gnd.n6161 gnd.n837 240.244
R7199 gnd.n6161 gnd.n839 240.244
R7200 gnd.n6157 gnd.n839 240.244
R7201 gnd.n6157 gnd.n845 240.244
R7202 gnd.n3687 gnd.n845 240.244
R7203 gnd.n2579 gnd.n2578 240.244
R7204 gnd.n2580 gnd.n2579 240.244
R7205 gnd.n3425 gnd.n2580 240.244
R7206 gnd.n3425 gnd.n2583 240.244
R7207 gnd.n2584 gnd.n2583 240.244
R7208 gnd.n2585 gnd.n2584 240.244
R7209 gnd.n3394 gnd.n2585 240.244
R7210 gnd.n3394 gnd.n2588 240.244
R7211 gnd.n2589 gnd.n2588 240.244
R7212 gnd.n2590 gnd.n2589 240.244
R7213 gnd.n3379 gnd.n2590 240.244
R7214 gnd.n3379 gnd.n2593 240.244
R7215 gnd.n2594 gnd.n2593 240.244
R7216 gnd.n2595 gnd.n2594 240.244
R7217 gnd.n3365 gnd.n2595 240.244
R7218 gnd.n3365 gnd.n2598 240.244
R7219 gnd.n2599 gnd.n2598 240.244
R7220 gnd.n2600 gnd.n2599 240.244
R7221 gnd.n3351 gnd.n2600 240.244
R7222 gnd.n3351 gnd.n2603 240.244
R7223 gnd.n2604 gnd.n2603 240.244
R7224 gnd.n2605 gnd.n2604 240.244
R7225 gnd.n3335 gnd.n2605 240.244
R7226 gnd.n3335 gnd.n2608 240.244
R7227 gnd.n2609 gnd.n2608 240.244
R7228 gnd.n2610 gnd.n2609 240.244
R7229 gnd.n3328 gnd.n2610 240.244
R7230 gnd.n3328 gnd.n2613 240.244
R7231 gnd.n2614 gnd.n2613 240.244
R7232 gnd.n2615 gnd.n2614 240.244
R7233 gnd.n4641 gnd.n2615 240.244
R7234 gnd.n4641 gnd.n2618 240.244
R7235 gnd.n2619 gnd.n2618 240.244
R7236 gnd.n2620 gnd.n2619 240.244
R7237 gnd.n4657 gnd.n2620 240.244
R7238 gnd.n4657 gnd.n2623 240.244
R7239 gnd.n2624 gnd.n2623 240.244
R7240 gnd.n2625 gnd.n2624 240.244
R7241 gnd.n3263 gnd.n2625 240.244
R7242 gnd.n3263 gnd.n2628 240.244
R7243 gnd.n2629 gnd.n2628 240.244
R7244 gnd.n2630 gnd.n2629 240.244
R7245 gnd.n3240 gnd.n2630 240.244
R7246 gnd.n3240 gnd.n2633 240.244
R7247 gnd.n2634 gnd.n2633 240.244
R7248 gnd.n2635 gnd.n2634 240.244
R7249 gnd.n3225 gnd.n2635 240.244
R7250 gnd.n3225 gnd.n2638 240.244
R7251 gnd.n2639 gnd.n2638 240.244
R7252 gnd.n2640 gnd.n2639 240.244
R7253 gnd.n3210 gnd.n2640 240.244
R7254 gnd.n3210 gnd.n2643 240.244
R7255 gnd.n2644 gnd.n2643 240.244
R7256 gnd.n2645 gnd.n2644 240.244
R7257 gnd.n3196 gnd.n2645 240.244
R7258 gnd.n3196 gnd.n2648 240.244
R7259 gnd.n2649 gnd.n2648 240.244
R7260 gnd.n2650 gnd.n2649 240.244
R7261 gnd.n4973 gnd.n2650 240.244
R7262 gnd.n4973 gnd.n2653 240.244
R7263 gnd.n2654 gnd.n2653 240.244
R7264 gnd.n2655 gnd.n2654 240.244
R7265 gnd.n5289 gnd.n2655 240.244
R7266 gnd.n5289 gnd.n2658 240.244
R7267 gnd.n2659 gnd.n2658 240.244
R7268 gnd.n2660 gnd.n2659 240.244
R7269 gnd.n4996 gnd.n2660 240.244
R7270 gnd.n4996 gnd.n2663 240.244
R7271 gnd.n2664 gnd.n2663 240.244
R7272 gnd.n2665 gnd.n2664 240.244
R7273 gnd.n5258 gnd.n2665 240.244
R7274 gnd.n5258 gnd.n2668 240.244
R7275 gnd.n2669 gnd.n2668 240.244
R7276 gnd.n2670 gnd.n2669 240.244
R7277 gnd.n5023 gnd.n2670 240.244
R7278 gnd.n5023 gnd.n2673 240.244
R7279 gnd.n2674 gnd.n2673 240.244
R7280 gnd.n2675 gnd.n2674 240.244
R7281 gnd.n5057 gnd.n2675 240.244
R7282 gnd.n5057 gnd.n2678 240.244
R7283 gnd.n2679 gnd.n2678 240.244
R7284 gnd.n5708 gnd.n2679 240.244
R7285 gnd.n3514 gnd.n3513 240.244
R7286 gnd.n3526 gnd.n3525 240.244
R7287 gnd.n3498 gnd.n3497 240.244
R7288 gnd.n3538 gnd.n3537 240.244
R7289 gnd.n3550 gnd.n3549 240.244
R7290 gnd.n3486 gnd.n3485 240.244
R7291 gnd.n3564 gnd.n3563 240.244
R7292 gnd.n3466 gnd.n3465 240.244
R7293 gnd.n4386 gnd.n4385 240.244
R7294 gnd.n4394 gnd.n4393 240.244
R7295 gnd.n4397 gnd.n4396 240.244
R7296 gnd.n4404 gnd.n4403 240.244
R7297 gnd.n4407 gnd.n3453 240.244
R7298 gnd.n4413 gnd.n3431 240.244
R7299 gnd.n4424 gnd.n3428 240.244
R7300 gnd.n4430 gnd.n3428 240.244
R7301 gnd.n4430 gnd.n3416 240.244
R7302 gnd.n4442 gnd.n3416 240.244
R7303 gnd.n4442 gnd.n3411 240.244
R7304 gnd.n4449 gnd.n3411 240.244
R7305 gnd.n4449 gnd.n3397 240.244
R7306 gnd.n3397 gnd.n3385 240.244
R7307 gnd.n4564 gnd.n3385 240.244
R7308 gnd.n4564 gnd.n3381 240.244
R7309 gnd.n4570 gnd.n3381 240.244
R7310 gnd.n4570 gnd.n3371 240.244
R7311 gnd.n4580 gnd.n3371 240.244
R7312 gnd.n4580 gnd.n3367 240.244
R7313 gnd.n4586 gnd.n3367 240.244
R7314 gnd.n4586 gnd.n3357 240.244
R7315 gnd.n4596 gnd.n3357 240.244
R7316 gnd.n4596 gnd.n3353 240.244
R7317 gnd.n4602 gnd.n3353 240.244
R7318 gnd.n4602 gnd.n3341 240.244
R7319 gnd.n4613 gnd.n3341 240.244
R7320 gnd.n4613 gnd.n3336 240.244
R7321 gnd.n4620 gnd.n3336 240.244
R7322 gnd.n4620 gnd.n3321 240.244
R7323 gnd.n3321 gnd.n3310 240.244
R7324 gnd.n4737 gnd.n3310 240.244
R7325 gnd.n4737 gnd.n3306 240.244
R7326 gnd.n4743 gnd.n3306 240.244
R7327 gnd.n4743 gnd.n3297 240.244
R7328 gnd.n4753 gnd.n3297 240.244
R7329 gnd.n4753 gnd.n3293 240.244
R7330 gnd.n4759 gnd.n3293 240.244
R7331 gnd.n4759 gnd.n3285 240.244
R7332 gnd.n4769 gnd.n3285 240.244
R7333 gnd.n4769 gnd.n3281 240.244
R7334 gnd.n4775 gnd.n3281 240.244
R7335 gnd.n4775 gnd.n3271 240.244
R7336 gnd.n4787 gnd.n3271 240.244
R7337 gnd.n4787 gnd.n3266 240.244
R7338 gnd.n4794 gnd.n3266 240.244
R7339 gnd.n4794 gnd.n3251 240.244
R7340 gnd.n3251 gnd.n3238 240.244
R7341 gnd.n4908 gnd.n3238 240.244
R7342 gnd.n4908 gnd.n3234 240.244
R7343 gnd.n4914 gnd.n3234 240.244
R7344 gnd.n4914 gnd.n3223 240.244
R7345 gnd.n4924 gnd.n3223 240.244
R7346 gnd.n4924 gnd.n3219 240.244
R7347 gnd.n4930 gnd.n3219 240.244
R7348 gnd.n4930 gnd.n3209 240.244
R7349 gnd.n4940 gnd.n3209 240.244
R7350 gnd.n4940 gnd.n3205 240.244
R7351 gnd.n4946 gnd.n3205 240.244
R7352 gnd.n4946 gnd.n3194 240.244
R7353 gnd.n4958 gnd.n3194 240.244
R7354 gnd.n4958 gnd.n3189 240.244
R7355 gnd.n4965 gnd.n3189 240.244
R7356 gnd.n4965 gnd.n3174 240.244
R7357 gnd.n3174 gnd.n3164 240.244
R7358 gnd.n5314 gnd.n3164 240.244
R7359 gnd.n5314 gnd.n3160 240.244
R7360 gnd.n5320 gnd.n3160 240.244
R7361 gnd.n5320 gnd.n3151 240.244
R7362 gnd.n5330 gnd.n3151 240.244
R7363 gnd.n5330 gnd.n3147 240.244
R7364 gnd.n5336 gnd.n3147 240.244
R7365 gnd.n5336 gnd.n3138 240.244
R7366 gnd.n5346 gnd.n3138 240.244
R7367 gnd.n5346 gnd.n3134 240.244
R7368 gnd.n5352 gnd.n3134 240.244
R7369 gnd.n5352 gnd.n3124 240.244
R7370 gnd.n5362 gnd.n3124 240.244
R7371 gnd.n5362 gnd.n3120 240.244
R7372 gnd.n5368 gnd.n3120 240.244
R7373 gnd.n5368 gnd.n3110 240.244
R7374 gnd.n5378 gnd.n3110 240.244
R7375 gnd.n5378 gnd.n3105 240.244
R7376 gnd.n5386 gnd.n3105 240.244
R7377 gnd.n5386 gnd.n3097 240.244
R7378 gnd.n5399 gnd.n3097 240.244
R7379 gnd.n5400 gnd.n5399 240.244
R7380 gnd.n5400 gnd.n2684 240.244
R7381 gnd.n3015 gnd.n3013 240.244
R7382 gnd.n3028 gnd.n2992 240.244
R7383 gnd.n3032 gnd.n3030 240.244
R7384 gnd.n3045 gnd.n2983 240.244
R7385 gnd.n3049 gnd.n3047 240.244
R7386 gnd.n3062 gnd.n2974 240.244
R7387 gnd.n3066 gnd.n3064 240.244
R7388 gnd.n3077 gnd.n2962 240.244
R7389 gnd.n3080 gnd.n3079 240.244
R7390 gnd.n3083 gnd.n3082 240.244
R7391 gnd.n3088 gnd.n3085 240.244
R7392 gnd.n3091 gnd.n3090 240.244
R7393 gnd.n5405 gnd.n3093 240.244
R7394 gnd.n5408 gnd.n5407 240.244
R7395 gnd.n4170 gnd.n4169 240.132
R7396 gnd.n5046 gnd.n5045 240.132
R7397 gnd.n6324 gnd.n6323 225.874
R7398 gnd.n6324 gnd.n673 225.874
R7399 gnd.n6332 gnd.n673 225.874
R7400 gnd.n6333 gnd.n6332 225.874
R7401 gnd.n6334 gnd.n6333 225.874
R7402 gnd.n6334 gnd.n667 225.874
R7403 gnd.n6342 gnd.n667 225.874
R7404 gnd.n6343 gnd.n6342 225.874
R7405 gnd.n6344 gnd.n6343 225.874
R7406 gnd.n6344 gnd.n661 225.874
R7407 gnd.n6352 gnd.n661 225.874
R7408 gnd.n6353 gnd.n6352 225.874
R7409 gnd.n6354 gnd.n6353 225.874
R7410 gnd.n6354 gnd.n655 225.874
R7411 gnd.n6362 gnd.n655 225.874
R7412 gnd.n6363 gnd.n6362 225.874
R7413 gnd.n6364 gnd.n6363 225.874
R7414 gnd.n6364 gnd.n649 225.874
R7415 gnd.n6372 gnd.n649 225.874
R7416 gnd.n6373 gnd.n6372 225.874
R7417 gnd.n6374 gnd.n6373 225.874
R7418 gnd.n6374 gnd.n643 225.874
R7419 gnd.n6382 gnd.n643 225.874
R7420 gnd.n6383 gnd.n6382 225.874
R7421 gnd.n6384 gnd.n6383 225.874
R7422 gnd.n6384 gnd.n637 225.874
R7423 gnd.n6392 gnd.n637 225.874
R7424 gnd.n6393 gnd.n6392 225.874
R7425 gnd.n6394 gnd.n6393 225.874
R7426 gnd.n6394 gnd.n631 225.874
R7427 gnd.n6402 gnd.n631 225.874
R7428 gnd.n6403 gnd.n6402 225.874
R7429 gnd.n6404 gnd.n6403 225.874
R7430 gnd.n6404 gnd.n625 225.874
R7431 gnd.n6412 gnd.n625 225.874
R7432 gnd.n6413 gnd.n6412 225.874
R7433 gnd.n6414 gnd.n6413 225.874
R7434 gnd.n6414 gnd.n619 225.874
R7435 gnd.n6422 gnd.n619 225.874
R7436 gnd.n6423 gnd.n6422 225.874
R7437 gnd.n6424 gnd.n6423 225.874
R7438 gnd.n6424 gnd.n613 225.874
R7439 gnd.n6432 gnd.n613 225.874
R7440 gnd.n6433 gnd.n6432 225.874
R7441 gnd.n6434 gnd.n6433 225.874
R7442 gnd.n6434 gnd.n607 225.874
R7443 gnd.n6442 gnd.n607 225.874
R7444 gnd.n6443 gnd.n6442 225.874
R7445 gnd.n6444 gnd.n6443 225.874
R7446 gnd.n6444 gnd.n601 225.874
R7447 gnd.n6452 gnd.n601 225.874
R7448 gnd.n6453 gnd.n6452 225.874
R7449 gnd.n6454 gnd.n6453 225.874
R7450 gnd.n6454 gnd.n595 225.874
R7451 gnd.n6462 gnd.n595 225.874
R7452 gnd.n6463 gnd.n6462 225.874
R7453 gnd.n6464 gnd.n6463 225.874
R7454 gnd.n6464 gnd.n589 225.874
R7455 gnd.n6472 gnd.n589 225.874
R7456 gnd.n6473 gnd.n6472 225.874
R7457 gnd.n6474 gnd.n6473 225.874
R7458 gnd.n6474 gnd.n583 225.874
R7459 gnd.n6482 gnd.n583 225.874
R7460 gnd.n6483 gnd.n6482 225.874
R7461 gnd.n6484 gnd.n6483 225.874
R7462 gnd.n6484 gnd.n577 225.874
R7463 gnd.n6492 gnd.n577 225.874
R7464 gnd.n6493 gnd.n6492 225.874
R7465 gnd.n6494 gnd.n6493 225.874
R7466 gnd.n6494 gnd.n571 225.874
R7467 gnd.n6502 gnd.n571 225.874
R7468 gnd.n6503 gnd.n6502 225.874
R7469 gnd.n6504 gnd.n6503 225.874
R7470 gnd.n6504 gnd.n565 225.874
R7471 gnd.n6512 gnd.n565 225.874
R7472 gnd.n6513 gnd.n6512 225.874
R7473 gnd.n6514 gnd.n6513 225.874
R7474 gnd.n6514 gnd.n559 225.874
R7475 gnd.n6522 gnd.n559 225.874
R7476 gnd.n6523 gnd.n6522 225.874
R7477 gnd.n6524 gnd.n6523 225.874
R7478 gnd.n6524 gnd.n553 225.874
R7479 gnd.n6532 gnd.n553 225.874
R7480 gnd.n6533 gnd.n6532 225.874
R7481 gnd.n6534 gnd.n6533 225.874
R7482 gnd.n6534 gnd.n547 225.874
R7483 gnd.n6542 gnd.n547 225.874
R7484 gnd.n6543 gnd.n6542 225.874
R7485 gnd.n6544 gnd.n6543 225.874
R7486 gnd.n6544 gnd.n541 225.874
R7487 gnd.n6552 gnd.n541 225.874
R7488 gnd.n6553 gnd.n6552 225.874
R7489 gnd.n6554 gnd.n6553 225.874
R7490 gnd.n6554 gnd.n535 225.874
R7491 gnd.n6562 gnd.n535 225.874
R7492 gnd.n6563 gnd.n6562 225.874
R7493 gnd.n6564 gnd.n6563 225.874
R7494 gnd.n6564 gnd.n529 225.874
R7495 gnd.n6572 gnd.n529 225.874
R7496 gnd.n6573 gnd.n6572 225.874
R7497 gnd.n6574 gnd.n6573 225.874
R7498 gnd.n6574 gnd.n523 225.874
R7499 gnd.n6582 gnd.n523 225.874
R7500 gnd.n6583 gnd.n6582 225.874
R7501 gnd.n6584 gnd.n6583 225.874
R7502 gnd.n6584 gnd.n517 225.874
R7503 gnd.n6592 gnd.n517 225.874
R7504 gnd.n6593 gnd.n6592 225.874
R7505 gnd.n6594 gnd.n6593 225.874
R7506 gnd.n6594 gnd.n511 225.874
R7507 gnd.n6602 gnd.n511 225.874
R7508 gnd.n6603 gnd.n6602 225.874
R7509 gnd.n6604 gnd.n6603 225.874
R7510 gnd.n6604 gnd.n505 225.874
R7511 gnd.n6612 gnd.n505 225.874
R7512 gnd.n6613 gnd.n6612 225.874
R7513 gnd.n6614 gnd.n6613 225.874
R7514 gnd.n6614 gnd.n499 225.874
R7515 gnd.n6622 gnd.n499 225.874
R7516 gnd.n6623 gnd.n6622 225.874
R7517 gnd.n6624 gnd.n6623 225.874
R7518 gnd.n6624 gnd.n493 225.874
R7519 gnd.n6632 gnd.n493 225.874
R7520 gnd.n6633 gnd.n6632 225.874
R7521 gnd.n6634 gnd.n6633 225.874
R7522 gnd.n6634 gnd.n487 225.874
R7523 gnd.n6642 gnd.n487 225.874
R7524 gnd.n6643 gnd.n6642 225.874
R7525 gnd.n6644 gnd.n6643 225.874
R7526 gnd.n6644 gnd.n481 225.874
R7527 gnd.n6652 gnd.n481 225.874
R7528 gnd.n6653 gnd.n6652 225.874
R7529 gnd.n6654 gnd.n6653 225.874
R7530 gnd.n6654 gnd.n475 225.874
R7531 gnd.n6662 gnd.n475 225.874
R7532 gnd.n6663 gnd.n6662 225.874
R7533 gnd.n6664 gnd.n6663 225.874
R7534 gnd.n6664 gnd.n469 225.874
R7535 gnd.n6672 gnd.n469 225.874
R7536 gnd.n6673 gnd.n6672 225.874
R7537 gnd.n6674 gnd.n6673 225.874
R7538 gnd.n6674 gnd.n463 225.874
R7539 gnd.n6682 gnd.n463 225.874
R7540 gnd.n6683 gnd.n6682 225.874
R7541 gnd.n6684 gnd.n6683 225.874
R7542 gnd.n6684 gnd.n457 225.874
R7543 gnd.n6692 gnd.n457 225.874
R7544 gnd.n6693 gnd.n6692 225.874
R7545 gnd.n6694 gnd.n6693 225.874
R7546 gnd.n6694 gnd.n451 225.874
R7547 gnd.n6703 gnd.n451 225.874
R7548 gnd.n6704 gnd.n6703 225.874
R7549 gnd.n6705 gnd.n6704 225.874
R7550 gnd.n6705 gnd.n446 225.874
R7551 gnd.n1689 gnd.t70 224.174
R7552 gnd.n900 gnd.t101 224.174
R7553 gnd.n2742 gnd.n2699 199.319
R7554 gnd.n2742 gnd.n2700 199.319
R7555 gnd.n3614 gnd.n3584 199.319
R7556 gnd.n3614 gnd.n3583 199.319
R7557 gnd.n4171 gnd.n4168 186.49
R7558 gnd.n5047 gnd.n5044 186.49
R7559 gnd.n1228 gnd.n1227 185
R7560 gnd.n1226 gnd.n1225 185
R7561 gnd.n1205 gnd.n1204 185
R7562 gnd.n1220 gnd.n1219 185
R7563 gnd.n1218 gnd.n1217 185
R7564 gnd.n1209 gnd.n1208 185
R7565 gnd.n1212 gnd.n1211 185
R7566 gnd.n1196 gnd.n1195 185
R7567 gnd.n1194 gnd.n1193 185
R7568 gnd.n1173 gnd.n1172 185
R7569 gnd.n1188 gnd.n1187 185
R7570 gnd.n1186 gnd.n1185 185
R7571 gnd.n1177 gnd.n1176 185
R7572 gnd.n1180 gnd.n1179 185
R7573 gnd.n1164 gnd.n1163 185
R7574 gnd.n1162 gnd.n1161 185
R7575 gnd.n1141 gnd.n1140 185
R7576 gnd.n1156 gnd.n1155 185
R7577 gnd.n1154 gnd.n1153 185
R7578 gnd.n1145 gnd.n1144 185
R7579 gnd.n1148 gnd.n1147 185
R7580 gnd.n1133 gnd.n1132 185
R7581 gnd.n1131 gnd.n1130 185
R7582 gnd.n1110 gnd.n1109 185
R7583 gnd.n1125 gnd.n1124 185
R7584 gnd.n1123 gnd.n1122 185
R7585 gnd.n1114 gnd.n1113 185
R7586 gnd.n1117 gnd.n1116 185
R7587 gnd.n1101 gnd.n1100 185
R7588 gnd.n1099 gnd.n1098 185
R7589 gnd.n1078 gnd.n1077 185
R7590 gnd.n1093 gnd.n1092 185
R7591 gnd.n1091 gnd.n1090 185
R7592 gnd.n1082 gnd.n1081 185
R7593 gnd.n1085 gnd.n1084 185
R7594 gnd.n1069 gnd.n1068 185
R7595 gnd.n1067 gnd.n1066 185
R7596 gnd.n1046 gnd.n1045 185
R7597 gnd.n1061 gnd.n1060 185
R7598 gnd.n1059 gnd.n1058 185
R7599 gnd.n1050 gnd.n1049 185
R7600 gnd.n1053 gnd.n1052 185
R7601 gnd.n1037 gnd.n1036 185
R7602 gnd.n1035 gnd.n1034 185
R7603 gnd.n1014 gnd.n1013 185
R7604 gnd.n1029 gnd.n1028 185
R7605 gnd.n1027 gnd.n1026 185
R7606 gnd.n1018 gnd.n1017 185
R7607 gnd.n1021 gnd.n1020 185
R7608 gnd.n1006 gnd.n1005 185
R7609 gnd.n1004 gnd.n1003 185
R7610 gnd.n983 gnd.n982 185
R7611 gnd.n998 gnd.n997 185
R7612 gnd.n996 gnd.n995 185
R7613 gnd.n987 gnd.n986 185
R7614 gnd.n990 gnd.n989 185
R7615 gnd.n1690 gnd.t69 178.987
R7616 gnd.n901 gnd.t102 178.987
R7617 gnd.n1 gnd.t297 170.774
R7618 gnd.n7 gnd.t287 170.103
R7619 gnd.n6 gnd.t152 170.103
R7620 gnd.n5 gnd.t1 170.103
R7621 gnd.n4 gnd.t132 170.103
R7622 gnd.n3 gnd.t148 170.103
R7623 gnd.n2 gnd.t317 170.103
R7624 gnd.n1 gnd.t323 170.103
R7625 gnd.n5079 gnd.n5078 163.367
R7626 gnd.n5083 gnd.n5082 163.367
R7627 gnd.n5087 gnd.n5086 163.367
R7628 gnd.n5091 gnd.n5090 163.367
R7629 gnd.n5095 gnd.n5094 163.367
R7630 gnd.n5099 gnd.n5098 163.367
R7631 gnd.n5103 gnd.n5102 163.367
R7632 gnd.n5107 gnd.n5106 163.367
R7633 gnd.n5111 gnd.n5110 163.367
R7634 gnd.n5115 gnd.n5114 163.367
R7635 gnd.n5119 gnd.n5118 163.367
R7636 gnd.n5123 gnd.n5122 163.367
R7637 gnd.n5127 gnd.n5126 163.367
R7638 gnd.n5131 gnd.n5130 163.367
R7639 gnd.n5136 gnd.n5135 163.367
R7640 gnd.n5140 gnd.n5139 163.367
R7641 gnd.n5228 gnd.n5227 163.367
R7642 gnd.n5224 gnd.n5223 163.367
R7643 gnd.n5219 gnd.n5218 163.367
R7644 gnd.n5215 gnd.n5214 163.367
R7645 gnd.n5211 gnd.n5210 163.367
R7646 gnd.n5207 gnd.n5206 163.367
R7647 gnd.n5203 gnd.n5202 163.367
R7648 gnd.n5199 gnd.n5198 163.367
R7649 gnd.n5195 gnd.n5194 163.367
R7650 gnd.n5191 gnd.n5190 163.367
R7651 gnd.n5187 gnd.n5186 163.367
R7652 gnd.n5183 gnd.n5182 163.367
R7653 gnd.n5179 gnd.n5178 163.367
R7654 gnd.n5175 gnd.n5174 163.367
R7655 gnd.n5171 gnd.n5170 163.367
R7656 gnd.n5167 gnd.n5166 163.367
R7657 gnd.n4279 gnd.n4278 163.367
R7658 gnd.n4278 gnd.n4273 163.367
R7659 gnd.n4274 gnd.n4273 163.367
R7660 gnd.n4274 gnd.n3398 163.367
R7661 gnd.n4554 gnd.n3398 163.367
R7662 gnd.n4554 gnd.n3399 163.367
R7663 gnd.n4550 gnd.n3399 163.367
R7664 gnd.n4550 gnd.n4549 163.367
R7665 gnd.n4549 gnd.n4548 163.367
R7666 gnd.n4548 gnd.n3402 163.367
R7667 gnd.n4462 gnd.n3402 163.367
R7668 gnd.n4538 gnd.n4462 163.367
R7669 gnd.n4538 gnd.n4463 163.367
R7670 gnd.n4534 gnd.n4463 163.367
R7671 gnd.n4534 gnd.n4533 163.367
R7672 gnd.n4533 gnd.n4467 163.367
R7673 gnd.n4478 gnd.n4467 163.367
R7674 gnd.n4478 gnd.n4475 163.367
R7675 gnd.n4522 gnd.n4475 163.367
R7676 gnd.n4522 gnd.n4476 163.367
R7677 gnd.n4518 gnd.n4476 163.367
R7678 gnd.n4518 gnd.n4482 163.367
R7679 gnd.n4490 gnd.n4482 163.367
R7680 gnd.n4508 gnd.n4490 163.367
R7681 gnd.n4508 gnd.n4491 163.367
R7682 gnd.n4504 gnd.n4491 163.367
R7683 gnd.n4504 gnd.n4503 163.367
R7684 gnd.n4503 gnd.n4495 163.367
R7685 gnd.n4495 gnd.n3322 163.367
R7686 gnd.n4727 gnd.n3322 163.367
R7687 gnd.n4727 gnd.n3323 163.367
R7688 gnd.n4723 gnd.n3323 163.367
R7689 gnd.n4723 gnd.n4722 163.367
R7690 gnd.n4722 gnd.n4721 163.367
R7691 gnd.n4721 gnd.n3326 163.367
R7692 gnd.n4636 gnd.n3326 163.367
R7693 gnd.n4636 gnd.n4633 163.367
R7694 gnd.n4710 gnd.n4633 163.367
R7695 gnd.n4710 gnd.n4634 163.367
R7696 gnd.n4706 gnd.n4634 163.367
R7697 gnd.n4706 gnd.n4640 163.367
R7698 gnd.n4651 gnd.n4640 163.367
R7699 gnd.n4651 gnd.n4649 163.367
R7700 gnd.n4695 gnd.n4649 163.367
R7701 gnd.n4695 gnd.n4650 163.367
R7702 gnd.n4691 gnd.n4650 163.367
R7703 gnd.n4691 gnd.n4655 163.367
R7704 gnd.n4670 gnd.n4655 163.367
R7705 gnd.n4681 gnd.n4670 163.367
R7706 gnd.n4681 gnd.n4671 163.367
R7707 gnd.n4677 gnd.n4671 163.367
R7708 gnd.n4677 gnd.n4676 163.367
R7709 gnd.n4676 gnd.n3265 163.367
R7710 gnd.n3265 gnd.n3252 163.367
R7711 gnd.n4898 gnd.n3252 163.367
R7712 gnd.n4898 gnd.n3253 163.367
R7713 gnd.n4894 gnd.n3253 163.367
R7714 gnd.n4894 gnd.n4893 163.367
R7715 gnd.n4893 gnd.n4892 163.367
R7716 gnd.n4892 gnd.n3256 163.367
R7717 gnd.n4808 gnd.n3256 163.367
R7718 gnd.n4882 gnd.n4808 163.367
R7719 gnd.n4882 gnd.n4809 163.367
R7720 gnd.n4878 gnd.n4809 163.367
R7721 gnd.n4878 gnd.n4877 163.367
R7722 gnd.n4877 gnd.n4813 163.367
R7723 gnd.n4824 gnd.n4813 163.367
R7724 gnd.n4824 gnd.n4821 163.367
R7725 gnd.n4866 gnd.n4821 163.367
R7726 gnd.n4866 gnd.n4822 163.367
R7727 gnd.n4862 gnd.n4822 163.367
R7728 gnd.n4862 gnd.n4828 163.367
R7729 gnd.n4841 gnd.n4828 163.367
R7730 gnd.n4852 gnd.n4841 163.367
R7731 gnd.n4852 gnd.n4842 163.367
R7732 gnd.n4848 gnd.n4842 163.367
R7733 gnd.n4848 gnd.n4847 163.367
R7734 gnd.n4847 gnd.n3188 163.367
R7735 gnd.n3188 gnd.n3175 163.367
R7736 gnd.n5304 gnd.n3175 163.367
R7737 gnd.n5304 gnd.n3176 163.367
R7738 gnd.n5300 gnd.n3176 163.367
R7739 gnd.n5300 gnd.n5299 163.367
R7740 gnd.n5299 gnd.n5298 163.367
R7741 gnd.n5298 gnd.n3179 163.367
R7742 gnd.n4982 gnd.n3179 163.367
R7743 gnd.n5288 gnd.n4982 163.367
R7744 gnd.n5288 gnd.n4983 163.367
R7745 gnd.n5284 gnd.n4983 163.367
R7746 gnd.n5284 gnd.n5283 163.367
R7747 gnd.n5283 gnd.n4987 163.367
R7748 gnd.n4999 gnd.n4987 163.367
R7749 gnd.n4999 gnd.n4995 163.367
R7750 gnd.n5272 gnd.n4995 163.367
R7751 gnd.n5272 gnd.n4997 163.367
R7752 gnd.n5268 gnd.n4997 163.367
R7753 gnd.n5268 gnd.n5003 163.367
R7754 gnd.n5011 gnd.n5003 163.367
R7755 gnd.n5257 gnd.n5011 163.367
R7756 gnd.n5257 gnd.n5012 163.367
R7757 gnd.n5253 gnd.n5012 163.367
R7758 gnd.n5253 gnd.n5252 163.367
R7759 gnd.n5252 gnd.n5015 163.367
R7760 gnd.n5024 gnd.n5015 163.367
R7761 gnd.n5243 gnd.n5024 163.367
R7762 gnd.n5243 gnd.n5025 163.367
R7763 gnd.n5239 gnd.n5025 163.367
R7764 gnd.n5239 gnd.n5238 163.367
R7765 gnd.n5238 gnd.n5029 163.367
R7766 gnd.n5056 gnd.n5029 163.367
R7767 gnd.n4263 gnd.n4262 163.367
R7768 gnd.n4262 gnd.n4261 163.367
R7769 gnd.n4258 gnd.n4257 163.367
R7770 gnd.n4255 gnd.n4189 163.367
R7771 gnd.n4251 gnd.n4249 163.367
R7772 gnd.n4247 gnd.n4191 163.367
R7773 gnd.n4243 gnd.n4241 163.367
R7774 gnd.n4239 gnd.n4193 163.367
R7775 gnd.n4235 gnd.n4233 163.367
R7776 gnd.n4231 gnd.n4195 163.367
R7777 gnd.n4227 gnd.n4225 163.367
R7778 gnd.n4223 gnd.n4197 163.367
R7779 gnd.n4219 gnd.n4217 163.367
R7780 gnd.n4215 gnd.n4199 163.367
R7781 gnd.n4211 gnd.n4209 163.367
R7782 gnd.n4206 gnd.n4205 163.367
R7783 gnd.n4346 gnd.n4344 163.367
R7784 gnd.n4342 gnd.n4144 163.367
R7785 gnd.n4337 gnd.n4335 163.367
R7786 gnd.n4333 gnd.n4148 163.367
R7787 gnd.n4329 gnd.n4327 163.367
R7788 gnd.n4325 gnd.n4150 163.367
R7789 gnd.n4321 gnd.n4319 163.367
R7790 gnd.n4317 gnd.n4152 163.367
R7791 gnd.n4313 gnd.n4311 163.367
R7792 gnd.n4309 gnd.n4154 163.367
R7793 gnd.n4305 gnd.n4303 163.367
R7794 gnd.n4301 gnd.n4156 163.367
R7795 gnd.n4297 gnd.n4295 163.367
R7796 gnd.n4293 gnd.n4158 163.367
R7797 gnd.n4289 gnd.n4287 163.367
R7798 gnd.n4285 gnd.n4160 163.367
R7799 gnd.n4267 gnd.n4163 163.367
R7800 gnd.n4271 gnd.n4163 163.367
R7801 gnd.n4271 gnd.n3409 163.367
R7802 gnd.n4452 gnd.n3409 163.367
R7803 gnd.n4452 gnd.n3393 163.367
R7804 gnd.n4456 gnd.n3393 163.367
R7805 gnd.n4457 gnd.n4456 163.367
R7806 gnd.n4457 gnd.n3404 163.367
R7807 gnd.n4546 gnd.n3404 163.367
R7808 gnd.n4546 gnd.n3407 163.367
R7809 gnd.n4542 gnd.n3407 163.367
R7810 gnd.n4542 gnd.n4541 163.367
R7811 gnd.n4541 gnd.n4461 163.367
R7812 gnd.n4469 gnd.n4461 163.367
R7813 gnd.n4531 gnd.n4469 163.367
R7814 gnd.n4531 gnd.n4470 163.367
R7815 gnd.n4527 gnd.n4470 163.367
R7816 gnd.n4527 gnd.n4526 163.367
R7817 gnd.n4526 gnd.n4474 163.367
R7818 gnd.n4484 gnd.n4474 163.367
R7819 gnd.n4516 gnd.n4484 163.367
R7820 gnd.n4516 gnd.n4485 163.367
R7821 gnd.n4512 gnd.n4485 163.367
R7822 gnd.n4512 gnd.n4511 163.367
R7823 gnd.n4511 gnd.n4489 163.367
R7824 gnd.n4497 gnd.n4489 163.367
R7825 gnd.n4501 gnd.n4497 163.367
R7826 gnd.n4501 gnd.n3333 163.367
R7827 gnd.n4623 gnd.n3333 163.367
R7828 gnd.n4623 gnd.n3318 163.367
R7829 gnd.n4627 gnd.n3318 163.367
R7830 gnd.n4628 gnd.n4627 163.367
R7831 gnd.n4628 gnd.n3330 163.367
R7832 gnd.n4719 gnd.n3330 163.367
R7833 gnd.n4719 gnd.n3331 163.367
R7834 gnd.n4715 gnd.n3331 163.367
R7835 gnd.n4715 gnd.n4714 163.367
R7836 gnd.n4714 gnd.n4632 163.367
R7837 gnd.n4643 gnd.n4632 163.367
R7838 gnd.n4704 gnd.n4643 163.367
R7839 gnd.n4704 gnd.n4644 163.367
R7840 gnd.n4700 gnd.n4644 163.367
R7841 gnd.n4700 gnd.n4699 163.367
R7842 gnd.n4699 gnd.n4648 163.367
R7843 gnd.n4659 gnd.n4648 163.367
R7844 gnd.n4689 gnd.n4659 163.367
R7845 gnd.n4689 gnd.n4660 163.367
R7846 gnd.n4685 gnd.n4660 163.367
R7847 gnd.n4685 gnd.n4669 163.367
R7848 gnd.n4669 gnd.n4668 163.367
R7849 gnd.n4668 gnd.n4664 163.367
R7850 gnd.n4664 gnd.n3262 163.367
R7851 gnd.n4797 gnd.n3262 163.367
R7852 gnd.n4798 gnd.n4797 163.367
R7853 gnd.n4798 gnd.n3248 163.367
R7854 gnd.n4802 gnd.n3248 163.367
R7855 gnd.n4803 gnd.n4802 163.367
R7856 gnd.n4803 gnd.n3259 163.367
R7857 gnd.n4890 gnd.n3259 163.367
R7858 gnd.n4890 gnd.n3260 163.367
R7859 gnd.n4886 gnd.n3260 163.367
R7860 gnd.n4886 gnd.n4885 163.367
R7861 gnd.n4885 gnd.n4807 163.367
R7862 gnd.n4815 gnd.n4807 163.367
R7863 gnd.n4875 gnd.n4815 163.367
R7864 gnd.n4875 gnd.n4816 163.367
R7865 gnd.n4871 gnd.n4816 163.367
R7866 gnd.n4871 gnd.n4870 163.367
R7867 gnd.n4870 gnd.n4820 163.367
R7868 gnd.n4830 gnd.n4820 163.367
R7869 gnd.n4860 gnd.n4830 163.367
R7870 gnd.n4860 gnd.n4831 163.367
R7871 gnd.n4856 gnd.n4831 163.367
R7872 gnd.n4856 gnd.n4840 163.367
R7873 gnd.n4840 gnd.n4839 163.367
R7874 gnd.n4839 gnd.n4835 163.367
R7875 gnd.n4835 gnd.n3186 163.367
R7876 gnd.n4968 gnd.n3186 163.367
R7877 gnd.n4969 gnd.n4968 163.367
R7878 gnd.n4969 gnd.n3173 163.367
R7879 gnd.n4976 gnd.n3173 163.367
R7880 gnd.n4977 gnd.n4976 163.367
R7881 gnd.n4977 gnd.n3182 163.367
R7882 gnd.n5296 gnd.n3182 163.367
R7883 gnd.n5296 gnd.n3184 163.367
R7884 gnd.n5292 gnd.n3184 163.367
R7885 gnd.n5292 gnd.n5291 163.367
R7886 gnd.n5291 gnd.n4981 163.367
R7887 gnd.n4989 gnd.n4981 163.367
R7888 gnd.n5281 gnd.n4989 163.367
R7889 gnd.n5281 gnd.n4990 163.367
R7890 gnd.n5277 gnd.n4990 163.367
R7891 gnd.n5277 gnd.n5276 163.367
R7892 gnd.n5276 gnd.n4994 163.367
R7893 gnd.n5005 gnd.n4994 163.367
R7894 gnd.n5266 gnd.n5005 163.367
R7895 gnd.n5266 gnd.n5006 163.367
R7896 gnd.n5262 gnd.n5006 163.367
R7897 gnd.n5262 gnd.n5261 163.367
R7898 gnd.n5261 gnd.n5010 163.367
R7899 gnd.n5017 gnd.n5010 163.367
R7900 gnd.n5250 gnd.n5017 163.367
R7901 gnd.n5250 gnd.n5018 163.367
R7902 gnd.n5246 gnd.n5018 163.367
R7903 gnd.n5246 gnd.n5245 163.367
R7904 gnd.n5245 gnd.n5022 163.367
R7905 gnd.n5031 gnd.n5022 163.367
R7906 gnd.n5236 gnd.n5031 163.367
R7907 gnd.n5236 gnd.n5032 163.367
R7908 gnd.n5232 gnd.n5032 163.367
R7909 gnd.n5053 gnd.n5052 156.462
R7910 gnd.n1168 gnd.n1136 153.042
R7911 gnd.n1232 gnd.n1231 152.079
R7912 gnd.n1200 gnd.n1199 152.079
R7913 gnd.n1168 gnd.n1167 152.079
R7914 gnd.n4176 gnd.n4175 152
R7915 gnd.n4177 gnd.n4166 152
R7916 gnd.n4179 gnd.n4178 152
R7917 gnd.n4181 gnd.n4164 152
R7918 gnd.n4183 gnd.n4182 152
R7919 gnd.n5051 gnd.n5035 152
R7920 gnd.n5043 gnd.n5036 152
R7921 gnd.n5042 gnd.n5041 152
R7922 gnd.n5040 gnd.n5037 152
R7923 gnd.n5038 gnd.t109 150.546
R7924 gnd.t319 gnd.n1210 147.661
R7925 gnd.t150 gnd.n1178 147.661
R7926 gnd.t321 gnd.n1146 147.661
R7927 gnd.t144 gnd.n1115 147.661
R7928 gnd.t156 gnd.n1083 147.661
R7929 gnd.t293 gnd.n1051 147.661
R7930 gnd.t130 gnd.n1019 147.661
R7931 gnd.t138 gnd.n988 147.661
R7932 gnd.n5158 gnd.n5141 143.351
R7933 gnd.n4204 gnd.n4143 143.351
R7934 gnd.n4345 gnd.n4143 143.351
R7935 gnd.n4173 gnd.t33 130.484
R7936 gnd.n4182 gnd.t103 126.766
R7937 gnd.n4180 gnd.t26 126.766
R7938 gnd.n4166 gnd.t54 126.766
R7939 gnd.n4174 gnd.t121 126.766
R7940 gnd.n5039 gnd.t88 126.766
R7941 gnd.n5041 gnd.t19 126.766
R7942 gnd.n5050 gnd.t75 126.766
R7943 gnd.n5052 gnd.t43 126.766
R7944 gnd.n6714 gnd.n6713 114.019
R7945 gnd.n6715 gnd.n6714 114.019
R7946 gnd.n6715 gnd.n440 114.019
R7947 gnd.n6723 gnd.n440 114.019
R7948 gnd.n6724 gnd.n6723 114.019
R7949 gnd.n6725 gnd.n6724 114.019
R7950 gnd.n6725 gnd.n434 114.019
R7951 gnd.n6733 gnd.n434 114.019
R7952 gnd.n6734 gnd.n6733 114.019
R7953 gnd.n6735 gnd.n6734 114.019
R7954 gnd.n6735 gnd.n428 114.019
R7955 gnd.n6743 gnd.n428 114.019
R7956 gnd.n6744 gnd.n6743 114.019
R7957 gnd.n6745 gnd.n6744 114.019
R7958 gnd.n6745 gnd.n422 114.019
R7959 gnd.n6753 gnd.n422 114.019
R7960 gnd.n6754 gnd.n6753 114.019
R7961 gnd.n6755 gnd.n6754 114.019
R7962 gnd.n6755 gnd.n416 114.019
R7963 gnd.n6763 gnd.n416 114.019
R7964 gnd.n6764 gnd.n6763 114.019
R7965 gnd.n6765 gnd.n6764 114.019
R7966 gnd.n6765 gnd.n410 114.019
R7967 gnd.n6773 gnd.n410 114.019
R7968 gnd.n6774 gnd.n6773 114.019
R7969 gnd.n6775 gnd.n6774 114.019
R7970 gnd.n6775 gnd.n404 114.019
R7971 gnd.n6783 gnd.n404 114.019
R7972 gnd.n6784 gnd.n6783 114.019
R7973 gnd.n6785 gnd.n6784 114.019
R7974 gnd.n6785 gnd.n398 114.019
R7975 gnd.n6793 gnd.n398 114.019
R7976 gnd.n6794 gnd.n6793 114.019
R7977 gnd.n6795 gnd.n6794 114.019
R7978 gnd.n6795 gnd.n392 114.019
R7979 gnd.n6803 gnd.n392 114.019
R7980 gnd.n6804 gnd.n6803 114.019
R7981 gnd.n6805 gnd.n6804 114.019
R7982 gnd.n6805 gnd.n386 114.019
R7983 gnd.n6813 gnd.n386 114.019
R7984 gnd.n6814 gnd.n6813 114.019
R7985 gnd.n6815 gnd.n6814 114.019
R7986 gnd.n6815 gnd.n380 114.019
R7987 gnd.n6823 gnd.n380 114.019
R7988 gnd.n6824 gnd.n6823 114.019
R7989 gnd.n6825 gnd.n6824 114.019
R7990 gnd.n6825 gnd.n374 114.019
R7991 gnd.n6833 gnd.n374 114.019
R7992 gnd.n6834 gnd.n6833 114.019
R7993 gnd.n6835 gnd.n6834 114.019
R7994 gnd.n6835 gnd.n368 114.019
R7995 gnd.n6843 gnd.n368 114.019
R7996 gnd.n6844 gnd.n6843 114.019
R7997 gnd.n6845 gnd.n6844 114.019
R7998 gnd.n6845 gnd.n362 114.019
R7999 gnd.n6853 gnd.n362 114.019
R8000 gnd.n6854 gnd.n6853 114.019
R8001 gnd.n6855 gnd.n6854 114.019
R8002 gnd.n6855 gnd.n356 114.019
R8003 gnd.n6863 gnd.n356 114.019
R8004 gnd.n6864 gnd.n6863 114.019
R8005 gnd.n6865 gnd.n6864 114.019
R8006 gnd.n6865 gnd.n350 114.019
R8007 gnd.n6873 gnd.n350 114.019
R8008 gnd.n6874 gnd.n6873 114.019
R8009 gnd.n6875 gnd.n6874 114.019
R8010 gnd.n6875 gnd.n344 114.019
R8011 gnd.n6883 gnd.n344 114.019
R8012 gnd.n6884 gnd.n6883 114.019
R8013 gnd.n6885 gnd.n6884 114.019
R8014 gnd.n6885 gnd.n338 114.019
R8015 gnd.n6893 gnd.n338 114.019
R8016 gnd.n6894 gnd.n6893 114.019
R8017 gnd.n6895 gnd.n6894 114.019
R8018 gnd.n6895 gnd.n332 114.019
R8019 gnd.n6903 gnd.n332 114.019
R8020 gnd.n6904 gnd.n6903 114.019
R8021 gnd.n6905 gnd.n6904 114.019
R8022 gnd.n6905 gnd.n326 114.019
R8023 gnd.n6913 gnd.n326 114.019
R8024 gnd.n6914 gnd.n6913 114.019
R8025 gnd.n6916 gnd.n6914 114.019
R8026 gnd.n6916 gnd.n6915 114.019
R8027 gnd.n1227 gnd.n1226 104.615
R8028 gnd.n1226 gnd.n1204 104.615
R8029 gnd.n1219 gnd.n1204 104.615
R8030 gnd.n1219 gnd.n1218 104.615
R8031 gnd.n1218 gnd.n1208 104.615
R8032 gnd.n1211 gnd.n1208 104.615
R8033 gnd.n1195 gnd.n1194 104.615
R8034 gnd.n1194 gnd.n1172 104.615
R8035 gnd.n1187 gnd.n1172 104.615
R8036 gnd.n1187 gnd.n1186 104.615
R8037 gnd.n1186 gnd.n1176 104.615
R8038 gnd.n1179 gnd.n1176 104.615
R8039 gnd.n1163 gnd.n1162 104.615
R8040 gnd.n1162 gnd.n1140 104.615
R8041 gnd.n1155 gnd.n1140 104.615
R8042 gnd.n1155 gnd.n1154 104.615
R8043 gnd.n1154 gnd.n1144 104.615
R8044 gnd.n1147 gnd.n1144 104.615
R8045 gnd.n1132 gnd.n1131 104.615
R8046 gnd.n1131 gnd.n1109 104.615
R8047 gnd.n1124 gnd.n1109 104.615
R8048 gnd.n1124 gnd.n1123 104.615
R8049 gnd.n1123 gnd.n1113 104.615
R8050 gnd.n1116 gnd.n1113 104.615
R8051 gnd.n1100 gnd.n1099 104.615
R8052 gnd.n1099 gnd.n1077 104.615
R8053 gnd.n1092 gnd.n1077 104.615
R8054 gnd.n1092 gnd.n1091 104.615
R8055 gnd.n1091 gnd.n1081 104.615
R8056 gnd.n1084 gnd.n1081 104.615
R8057 gnd.n1068 gnd.n1067 104.615
R8058 gnd.n1067 gnd.n1045 104.615
R8059 gnd.n1060 gnd.n1045 104.615
R8060 gnd.n1060 gnd.n1059 104.615
R8061 gnd.n1059 gnd.n1049 104.615
R8062 gnd.n1052 gnd.n1049 104.615
R8063 gnd.n1036 gnd.n1035 104.615
R8064 gnd.n1035 gnd.n1013 104.615
R8065 gnd.n1028 gnd.n1013 104.615
R8066 gnd.n1028 gnd.n1027 104.615
R8067 gnd.n1027 gnd.n1017 104.615
R8068 gnd.n1020 gnd.n1017 104.615
R8069 gnd.n1005 gnd.n1004 104.615
R8070 gnd.n1004 gnd.n982 104.615
R8071 gnd.n997 gnd.n982 104.615
R8072 gnd.n997 gnd.n996 104.615
R8073 gnd.n996 gnd.n986 104.615
R8074 gnd.n989 gnd.n986 104.615
R8075 gnd.n1615 gnd.t25 100.632
R8076 gnd.n879 gnd.t93 100.632
R8077 gnd.n7272 gnd.n112 99.6594
R8078 gnd.n7270 gnd.n7269 99.6594
R8079 gnd.n7265 gnd.n119 99.6594
R8080 gnd.n7263 gnd.n7262 99.6594
R8081 gnd.n7258 gnd.n126 99.6594
R8082 gnd.n7256 gnd.n7255 99.6594
R8083 gnd.n7251 gnd.n133 99.6594
R8084 gnd.n7249 gnd.n7248 99.6594
R8085 gnd.n7241 gnd.n140 99.6594
R8086 gnd.n7239 gnd.n7238 99.6594
R8087 gnd.n7234 gnd.n147 99.6594
R8088 gnd.n7232 gnd.n7231 99.6594
R8089 gnd.n7227 gnd.n154 99.6594
R8090 gnd.n7225 gnd.n7224 99.6594
R8091 gnd.n7220 gnd.n161 99.6594
R8092 gnd.n7218 gnd.n7217 99.6594
R8093 gnd.n7213 gnd.n168 99.6594
R8094 gnd.n7211 gnd.n7210 99.6594
R8095 gnd.n173 gnd.n172 99.6594
R8096 gnd.n5697 gnd.n5696 99.6594
R8097 gnd.n5691 gnd.n2693 99.6594
R8098 gnd.n5688 gnd.n2694 99.6594
R8099 gnd.n5684 gnd.n2695 99.6594
R8100 gnd.n5680 gnd.n2696 99.6594
R8101 gnd.n5676 gnd.n2697 99.6594
R8102 gnd.n5672 gnd.n2698 99.6594
R8103 gnd.n5668 gnd.n2699 99.6594
R8104 gnd.n5663 gnd.n2701 99.6594
R8105 gnd.n5659 gnd.n2702 99.6594
R8106 gnd.n5655 gnd.n2703 99.6594
R8107 gnd.n5651 gnd.n2704 99.6594
R8108 gnd.n5647 gnd.n2705 99.6594
R8109 gnd.n5643 gnd.n2706 99.6594
R8110 gnd.n5639 gnd.n2707 99.6594
R8111 gnd.n5635 gnd.n2708 99.6594
R8112 gnd.n5631 gnd.n2709 99.6594
R8113 gnd.n2765 gnd.n2710 99.6594
R8114 gnd.n4376 gnd.n4375 99.6594
R8115 gnd.n4371 gnd.n3590 99.6594
R8116 gnd.n4367 gnd.n3589 99.6594
R8117 gnd.n4363 gnd.n3588 99.6594
R8118 gnd.n4359 gnd.n3587 99.6594
R8119 gnd.n4355 gnd.n3586 99.6594
R8120 gnd.n4351 gnd.n3585 99.6594
R8121 gnd.n4135 gnd.n3583 99.6594
R8122 gnd.n4133 gnd.n3582 99.6594
R8123 gnd.n4129 gnd.n3581 99.6594
R8124 gnd.n4125 gnd.n3580 99.6594
R8125 gnd.n4121 gnd.n3579 99.6594
R8126 gnd.n4117 gnd.n3578 99.6594
R8127 gnd.n4113 gnd.n3577 99.6594
R8128 gnd.n4109 gnd.n3576 99.6594
R8129 gnd.n4105 gnd.n3575 99.6594
R8130 gnd.n4101 gnd.n3574 99.6594
R8131 gnd.n3632 gnd.n3573 99.6594
R8132 gnd.n6075 gnd.n6074 99.6594
R8133 gnd.n6069 gnd.n2231 99.6594
R8134 gnd.n6066 gnd.n2232 99.6594
R8135 gnd.n6062 gnd.n2233 99.6594
R8136 gnd.n6058 gnd.n2234 99.6594
R8137 gnd.n6054 gnd.n2235 99.6594
R8138 gnd.n6050 gnd.n2236 99.6594
R8139 gnd.n6046 gnd.n2237 99.6594
R8140 gnd.n6042 gnd.n2238 99.6594
R8141 gnd.n6037 gnd.n2239 99.6594
R8142 gnd.n6033 gnd.n2240 99.6594
R8143 gnd.n6029 gnd.n2241 99.6594
R8144 gnd.n6025 gnd.n2242 99.6594
R8145 gnd.n6021 gnd.n2243 99.6594
R8146 gnd.n6017 gnd.n2244 99.6594
R8147 gnd.n6013 gnd.n2245 99.6594
R8148 gnd.n6009 gnd.n2246 99.6594
R8149 gnd.n6005 gnd.n2247 99.6594
R8150 gnd.n2302 gnd.n2248 99.6594
R8151 gnd.n6114 gnd.n6082 99.6594
R8152 gnd.n6112 gnd.n6081 99.6594
R8153 gnd.n6108 gnd.n6080 99.6594
R8154 gnd.n6104 gnd.n6079 99.6594
R8155 gnd.n6100 gnd.n6078 99.6594
R8156 gnd.n6096 gnd.n6077 99.6594
R8157 gnd.n6126 gnd.n6124 99.6594
R8158 gnd.n6132 gnd.n878 99.6594
R8159 gnd.n1827 gnd.n1558 99.6594
R8160 gnd.n1584 gnd.n1565 99.6594
R8161 gnd.n1586 gnd.n1566 99.6594
R8162 gnd.n1594 gnd.n1567 99.6594
R8163 gnd.n1596 gnd.n1568 99.6594
R8164 gnd.n1604 gnd.n1569 99.6594
R8165 gnd.n1606 gnd.n1570 99.6594
R8166 gnd.n1614 gnd.n1571 99.6594
R8167 gnd.n920 gnd.n885 99.6594
R8168 gnd.n924 gnd.n886 99.6594
R8169 gnd.n930 gnd.n887 99.6594
R8170 gnd.n934 gnd.n888 99.6594
R8171 gnd.n940 gnd.n889 99.6594
R8172 gnd.n944 gnd.n890 99.6594
R8173 gnd.n950 gnd.n891 99.6594
R8174 gnd.n954 gnd.n892 99.6594
R8175 gnd.n960 gnd.n893 99.6594
R8176 gnd.n964 gnd.n894 99.6594
R8177 gnd.n970 gnd.n895 99.6594
R8178 gnd.n973 gnd.n896 99.6594
R8179 gnd.n2230 gnd.n2229 99.6594
R8180 gnd.n1742 gnd.n1741 99.6594
R8181 gnd.n1736 gnd.n1653 99.6594
R8182 gnd.n1733 gnd.n1654 99.6594
R8183 gnd.n1729 gnd.n1655 99.6594
R8184 gnd.n1725 gnd.n1656 99.6594
R8185 gnd.n1721 gnd.n1657 99.6594
R8186 gnd.n1717 gnd.n1658 99.6594
R8187 gnd.n1713 gnd.n1659 99.6594
R8188 gnd.n1709 gnd.n1660 99.6594
R8189 gnd.n1705 gnd.n1661 99.6594
R8190 gnd.n1701 gnd.n1662 99.6594
R8191 gnd.n1697 gnd.n1663 99.6594
R8192 gnd.n1744 gnd.n1652 99.6594
R8193 gnd.n7120 gnd.n7119 99.6594
R8194 gnd.n7125 gnd.n7124 99.6594
R8195 gnd.n7128 gnd.n7127 99.6594
R8196 gnd.n7133 gnd.n7132 99.6594
R8197 gnd.n7136 gnd.n7135 99.6594
R8198 gnd.n7141 gnd.n7140 99.6594
R8199 gnd.n7144 gnd.n7143 99.6594
R8200 gnd.n7149 gnd.n7148 99.6594
R8201 gnd.n7152 gnd.n99 99.6594
R8202 gnd.n2775 gnd.n2711 99.6594
R8203 gnd.n3007 gnd.n2712 99.6594
R8204 gnd.n2998 gnd.n2713 99.6594
R8205 gnd.n3023 gnd.n2714 99.6594
R8206 gnd.n2989 gnd.n2715 99.6594
R8207 gnd.n3040 gnd.n2716 99.6594
R8208 gnd.n2980 gnd.n2717 99.6594
R8209 gnd.n3057 gnd.n2718 99.6594
R8210 gnd.n2971 gnd.n2719 99.6594
R8211 gnd.n3507 gnd.n3473 99.6594
R8212 gnd.n3520 gnd.n3474 99.6594
R8213 gnd.n3531 gnd.n3475 99.6594
R8214 gnd.n3493 gnd.n3476 99.6594
R8215 gnd.n3544 gnd.n3477 99.6594
R8216 gnd.n3555 gnd.n3478 99.6594
R8217 gnd.n3480 gnd.n3479 99.6594
R8218 gnd.n3571 gnd.n3570 99.6594
R8219 gnd.n4379 gnd.n4378 99.6594
R8220 gnd.n3864 gnd.n2249 99.6594
R8221 gnd.n3861 gnd.n2250 99.6594
R8222 gnd.n3857 gnd.n2251 99.6594
R8223 gnd.n3853 gnd.n2252 99.6594
R8224 gnd.n3849 gnd.n2253 99.6594
R8225 gnd.n3845 gnd.n2254 99.6594
R8226 gnd.n3841 gnd.n2255 99.6594
R8227 gnd.n3837 gnd.n2256 99.6594
R8228 gnd.n3833 gnd.n2257 99.6594
R8229 gnd.n3862 gnd.n2249 99.6594
R8230 gnd.n3858 gnd.n2250 99.6594
R8231 gnd.n3854 gnd.n2251 99.6594
R8232 gnd.n3850 gnd.n2252 99.6594
R8233 gnd.n3846 gnd.n2253 99.6594
R8234 gnd.n3842 gnd.n2254 99.6594
R8235 gnd.n3838 gnd.n2255 99.6594
R8236 gnd.n3834 gnd.n2256 99.6594
R8237 gnd.n3822 gnd.n2257 99.6594
R8238 gnd.n4378 gnd.n3471 99.6594
R8239 gnd.n3571 gnd.n3569 99.6594
R8240 gnd.n3556 gnd.n3479 99.6594
R8241 gnd.n3543 gnd.n3478 99.6594
R8242 gnd.n3494 gnd.n3477 99.6594
R8243 gnd.n3532 gnd.n3476 99.6594
R8244 gnd.n3519 gnd.n3475 99.6594
R8245 gnd.n3508 gnd.n3474 99.6594
R8246 gnd.n3504 gnd.n3473 99.6594
R8247 gnd.n3006 gnd.n2711 99.6594
R8248 gnd.n2997 gnd.n2712 99.6594
R8249 gnd.n3022 gnd.n2713 99.6594
R8250 gnd.n2988 gnd.n2714 99.6594
R8251 gnd.n3039 gnd.n2715 99.6594
R8252 gnd.n2979 gnd.n2716 99.6594
R8253 gnd.n3056 gnd.n2717 99.6594
R8254 gnd.n2970 gnd.n2718 99.6594
R8255 gnd.n2966 gnd.n2719 99.6594
R8256 gnd.n7153 gnd.n7152 99.6594
R8257 gnd.n7148 gnd.n7147 99.6594
R8258 gnd.n7143 gnd.n7142 99.6594
R8259 gnd.n7140 gnd.n7139 99.6594
R8260 gnd.n7135 gnd.n7134 99.6594
R8261 gnd.n7132 gnd.n7131 99.6594
R8262 gnd.n7127 gnd.n7126 99.6594
R8263 gnd.n7124 gnd.n7123 99.6594
R8264 gnd.n7119 gnd.n7118 99.6594
R8265 gnd.n1742 gnd.n1665 99.6594
R8266 gnd.n1734 gnd.n1653 99.6594
R8267 gnd.n1730 gnd.n1654 99.6594
R8268 gnd.n1726 gnd.n1655 99.6594
R8269 gnd.n1722 gnd.n1656 99.6594
R8270 gnd.n1718 gnd.n1657 99.6594
R8271 gnd.n1714 gnd.n1658 99.6594
R8272 gnd.n1710 gnd.n1659 99.6594
R8273 gnd.n1706 gnd.n1660 99.6594
R8274 gnd.n1702 gnd.n1661 99.6594
R8275 gnd.n1698 gnd.n1662 99.6594
R8276 gnd.n1694 gnd.n1663 99.6594
R8277 gnd.n1745 gnd.n1744 99.6594
R8278 gnd.n2230 gnd.n897 99.6594
R8279 gnd.n971 gnd.n896 99.6594
R8280 gnd.n963 gnd.n895 99.6594
R8281 gnd.n961 gnd.n894 99.6594
R8282 gnd.n953 gnd.n893 99.6594
R8283 gnd.n951 gnd.n892 99.6594
R8284 gnd.n943 gnd.n891 99.6594
R8285 gnd.n941 gnd.n890 99.6594
R8286 gnd.n933 gnd.n889 99.6594
R8287 gnd.n931 gnd.n888 99.6594
R8288 gnd.n923 gnd.n887 99.6594
R8289 gnd.n921 gnd.n886 99.6594
R8290 gnd.n913 gnd.n885 99.6594
R8291 gnd.n1828 gnd.n1827 99.6594
R8292 gnd.n1587 gnd.n1565 99.6594
R8293 gnd.n1593 gnd.n1566 99.6594
R8294 gnd.n1597 gnd.n1567 99.6594
R8295 gnd.n1603 gnd.n1568 99.6594
R8296 gnd.n1607 gnd.n1569 99.6594
R8297 gnd.n1613 gnd.n1570 99.6594
R8298 gnd.n1571 gnd.n1555 99.6594
R8299 gnd.n6125 gnd.n878 99.6594
R8300 gnd.n6124 gnd.n884 99.6594
R8301 gnd.n6099 gnd.n6077 99.6594
R8302 gnd.n6103 gnd.n6078 99.6594
R8303 gnd.n6107 gnd.n6079 99.6594
R8304 gnd.n6111 gnd.n6080 99.6594
R8305 gnd.n6115 gnd.n6081 99.6594
R8306 gnd.n6083 gnd.n6082 99.6594
R8307 gnd.n6075 gnd.n2261 99.6594
R8308 gnd.n6067 gnd.n2231 99.6594
R8309 gnd.n6063 gnd.n2232 99.6594
R8310 gnd.n6059 gnd.n2233 99.6594
R8311 gnd.n6055 gnd.n2234 99.6594
R8312 gnd.n6051 gnd.n2235 99.6594
R8313 gnd.n6047 gnd.n2236 99.6594
R8314 gnd.n6043 gnd.n2237 99.6594
R8315 gnd.n6038 gnd.n2238 99.6594
R8316 gnd.n6034 gnd.n2239 99.6594
R8317 gnd.n6030 gnd.n2240 99.6594
R8318 gnd.n6026 gnd.n2241 99.6594
R8319 gnd.n6022 gnd.n2242 99.6594
R8320 gnd.n6018 gnd.n2243 99.6594
R8321 gnd.n6014 gnd.n2244 99.6594
R8322 gnd.n6010 gnd.n2245 99.6594
R8323 gnd.n6006 gnd.n2246 99.6594
R8324 gnd.n2301 gnd.n2247 99.6594
R8325 gnd.n5998 gnd.n2248 99.6594
R8326 gnd.n4100 gnd.n3573 99.6594
R8327 gnd.n4104 gnd.n3574 99.6594
R8328 gnd.n4108 gnd.n3575 99.6594
R8329 gnd.n4112 gnd.n3576 99.6594
R8330 gnd.n4116 gnd.n3577 99.6594
R8331 gnd.n4120 gnd.n3578 99.6594
R8332 gnd.n4124 gnd.n3579 99.6594
R8333 gnd.n4128 gnd.n3580 99.6594
R8334 gnd.n4132 gnd.n3581 99.6594
R8335 gnd.n4136 gnd.n3582 99.6594
R8336 gnd.n4350 gnd.n3584 99.6594
R8337 gnd.n4354 gnd.n3585 99.6594
R8338 gnd.n4358 gnd.n3586 99.6594
R8339 gnd.n4362 gnd.n3587 99.6594
R8340 gnd.n4366 gnd.n3588 99.6594
R8341 gnd.n4370 gnd.n3589 99.6594
R8342 gnd.n3592 gnd.n3590 99.6594
R8343 gnd.n4376 gnd.n3591 99.6594
R8344 gnd.n5697 gnd.n2723 99.6594
R8345 gnd.n5689 gnd.n2693 99.6594
R8346 gnd.n5685 gnd.n2694 99.6594
R8347 gnd.n5681 gnd.n2695 99.6594
R8348 gnd.n5677 gnd.n2696 99.6594
R8349 gnd.n5673 gnd.n2697 99.6594
R8350 gnd.n5669 gnd.n2698 99.6594
R8351 gnd.n5664 gnd.n2700 99.6594
R8352 gnd.n5660 gnd.n2701 99.6594
R8353 gnd.n5656 gnd.n2702 99.6594
R8354 gnd.n5652 gnd.n2703 99.6594
R8355 gnd.n5648 gnd.n2704 99.6594
R8356 gnd.n5644 gnd.n2705 99.6594
R8357 gnd.n5640 gnd.n2706 99.6594
R8358 gnd.n5636 gnd.n2707 99.6594
R8359 gnd.n5632 gnd.n2708 99.6594
R8360 gnd.n2764 gnd.n2709 99.6594
R8361 gnd.n5624 gnd.n2710 99.6594
R8362 gnd.n172 gnd.n169 99.6594
R8363 gnd.n7212 gnd.n7211 99.6594
R8364 gnd.n168 gnd.n162 99.6594
R8365 gnd.n7219 gnd.n7218 99.6594
R8366 gnd.n161 gnd.n155 99.6594
R8367 gnd.n7226 gnd.n7225 99.6594
R8368 gnd.n154 gnd.n148 99.6594
R8369 gnd.n7233 gnd.n7232 99.6594
R8370 gnd.n147 gnd.n141 99.6594
R8371 gnd.n7240 gnd.n7239 99.6594
R8372 gnd.n140 gnd.n134 99.6594
R8373 gnd.n7250 gnd.n7249 99.6594
R8374 gnd.n133 gnd.n127 99.6594
R8375 gnd.n7257 gnd.n7256 99.6594
R8376 gnd.n126 gnd.n120 99.6594
R8377 gnd.n7264 gnd.n7263 99.6594
R8378 gnd.n119 gnd.n113 99.6594
R8379 gnd.n7271 gnd.n7270 99.6594
R8380 gnd.n112 gnd.n109 99.6594
R8381 gnd.n3511 gnd.n3440 99.6594
R8382 gnd.n3513 gnd.n3441 99.6594
R8383 gnd.n3526 gnd.n3442 99.6594
R8384 gnd.n3498 gnd.n3443 99.6594
R8385 gnd.n3537 gnd.n3444 99.6594
R8386 gnd.n3550 gnd.n3445 99.6594
R8387 gnd.n3486 gnd.n3446 99.6594
R8388 gnd.n3564 gnd.n3447 99.6594
R8389 gnd.n3466 gnd.n3448 99.6594
R8390 gnd.n4385 gnd.n3449 99.6594
R8391 gnd.n4394 gnd.n3450 99.6594
R8392 gnd.n4396 gnd.n3451 99.6594
R8393 gnd.n4404 gnd.n3452 99.6594
R8394 gnd.n4414 gnd.n3453 99.6594
R8395 gnd.n3514 gnd.n3440 99.6594
R8396 gnd.n3525 gnd.n3441 99.6594
R8397 gnd.n3497 gnd.n3442 99.6594
R8398 gnd.n3538 gnd.n3443 99.6594
R8399 gnd.n3549 gnd.n3444 99.6594
R8400 gnd.n3485 gnd.n3445 99.6594
R8401 gnd.n3563 gnd.n3446 99.6594
R8402 gnd.n3465 gnd.n3447 99.6594
R8403 gnd.n4386 gnd.n3448 99.6594
R8404 gnd.n4393 gnd.n3449 99.6594
R8405 gnd.n4397 gnd.n3450 99.6594
R8406 gnd.n4403 gnd.n3451 99.6594
R8407 gnd.n4407 gnd.n3452 99.6594
R8408 gnd.n4414 gnd.n4413 99.6594
R8409 gnd.n3012 gnd.n2681 99.6594
R8410 gnd.n3015 gnd.n3014 99.6594
R8411 gnd.n3029 gnd.n3028 99.6594
R8412 gnd.n3032 gnd.n3031 99.6594
R8413 gnd.n3046 gnd.n3045 99.6594
R8414 gnd.n3049 gnd.n3048 99.6594
R8415 gnd.n3063 gnd.n3062 99.6594
R8416 gnd.n3066 gnd.n3065 99.6594
R8417 gnd.n3078 gnd.n3077 99.6594
R8418 gnd.n3081 gnd.n3080 99.6594
R8419 gnd.n3084 gnd.n3083 99.6594
R8420 gnd.n3089 gnd.n3088 99.6594
R8421 gnd.n3092 gnd.n3091 99.6594
R8422 gnd.n5406 gnd.n5405 99.6594
R8423 gnd.n5407 gnd.n5406 99.6594
R8424 gnd.n3093 gnd.n3092 99.6594
R8425 gnd.n3090 gnd.n3089 99.6594
R8426 gnd.n3085 gnd.n3084 99.6594
R8427 gnd.n3082 gnd.n3081 99.6594
R8428 gnd.n3079 gnd.n3078 99.6594
R8429 gnd.n3065 gnd.n2962 99.6594
R8430 gnd.n3064 gnd.n3063 99.6594
R8431 gnd.n3048 gnd.n2974 99.6594
R8432 gnd.n3047 gnd.n3046 99.6594
R8433 gnd.n3031 gnd.n2983 99.6594
R8434 gnd.n3030 gnd.n3029 99.6594
R8435 gnd.n3014 gnd.n2992 99.6594
R8436 gnd.n3013 gnd.n3012 99.6594
R8437 gnd.n3457 gnd.t98 98.63
R8438 gnd.n7150 gnd.t31 98.63
R8439 gnd.n2967 gnd.t66 98.63
R8440 gnd.n3469 gnd.t86 98.63
R8441 gnd.n2744 gnd.t63 98.63
R8442 gnd.n2766 gnd.t39 98.63
R8443 gnd.n175 gnd.t125 98.63
R8444 gnd.n7243 gnd.t41 98.63
R8445 gnd.n2281 gnd.t120 98.63
R8446 gnd.n2303 gnd.t114 98.63
R8447 gnd.n3634 gnd.t48 98.63
R8448 gnd.n3612 gnd.t83 98.63
R8449 gnd.n3823 gnd.t74 98.63
R8450 gnd.n5415 gnd.t80 98.63
R8451 gnd.n4145 gnd.t117 96.6984
R8452 gnd.n5159 gnd.t52 96.6984
R8453 gnd.n4200 gnd.t60 96.6906
R8454 gnd.n5074 gnd.t107 96.6906
R8455 gnd.n4173 gnd.n4172 81.8399
R8456 gnd.n1616 gnd.t24 74.8376
R8457 gnd.n880 gnd.t94 74.8376
R8458 gnd.n4146 gnd.t116 72.8438
R8459 gnd.n5160 gnd.t53 72.8438
R8460 gnd.n4174 gnd.n4167 72.8411
R8461 gnd.n4180 gnd.n4165 72.8411
R8462 gnd.n5050 gnd.n5049 72.8411
R8463 gnd.n3458 gnd.t97 72.836
R8464 gnd.n4201 gnd.t59 72.836
R8465 gnd.n5075 gnd.t108 72.836
R8466 gnd.n7151 gnd.t32 72.836
R8467 gnd.n2968 gnd.t65 72.836
R8468 gnd.n3470 gnd.t87 72.836
R8469 gnd.n2745 gnd.t62 72.836
R8470 gnd.n2767 gnd.t38 72.836
R8471 gnd.n176 gnd.t126 72.836
R8472 gnd.n7244 gnd.t42 72.836
R8473 gnd.n2282 gnd.t119 72.836
R8474 gnd.n2304 gnd.t113 72.836
R8475 gnd.n3635 gnd.t49 72.836
R8476 gnd.n3613 gnd.t84 72.836
R8477 gnd.n3824 gnd.t73 72.836
R8478 gnd.n5416 gnd.t81 72.836
R8479 gnd.n5078 gnd.n5058 71.676
R8480 gnd.n5082 gnd.n5059 71.676
R8481 gnd.n5086 gnd.n5060 71.676
R8482 gnd.n5090 gnd.n5061 71.676
R8483 gnd.n5094 gnd.n5062 71.676
R8484 gnd.n5098 gnd.n5063 71.676
R8485 gnd.n5102 gnd.n5064 71.676
R8486 gnd.n5106 gnd.n5065 71.676
R8487 gnd.n5110 gnd.n5066 71.676
R8488 gnd.n5114 gnd.n5067 71.676
R8489 gnd.n5118 gnd.n5068 71.676
R8490 gnd.n5122 gnd.n5069 71.676
R8491 gnd.n5126 gnd.n5070 71.676
R8492 gnd.n5130 gnd.n5071 71.676
R8493 gnd.n5135 gnd.n5072 71.676
R8494 gnd.n5139 gnd.n5073 71.676
R8495 gnd.n5228 gnd.n5158 71.676
R8496 gnd.n5224 gnd.n5157 71.676
R8497 gnd.n5219 gnd.n5156 71.676
R8498 gnd.n5215 gnd.n5155 71.676
R8499 gnd.n5211 gnd.n5154 71.676
R8500 gnd.n5207 gnd.n5153 71.676
R8501 gnd.n5203 gnd.n5152 71.676
R8502 gnd.n5199 gnd.n5151 71.676
R8503 gnd.n5195 gnd.n5150 71.676
R8504 gnd.n5191 gnd.n5149 71.676
R8505 gnd.n5187 gnd.n5148 71.676
R8506 gnd.n5183 gnd.n5147 71.676
R8507 gnd.n5179 gnd.n5146 71.676
R8508 gnd.n5175 gnd.n5145 71.676
R8509 gnd.n5171 gnd.n5144 71.676
R8510 gnd.n5167 gnd.n5143 71.676
R8511 gnd.n5163 gnd.n5142 71.676
R8512 gnd.n4266 gnd.n4185 71.676
R8513 gnd.n4261 gnd.n4187 71.676
R8514 gnd.n4257 gnd.n4256 71.676
R8515 gnd.n4250 gnd.n4189 71.676
R8516 gnd.n4249 gnd.n4248 71.676
R8517 gnd.n4242 gnd.n4191 71.676
R8518 gnd.n4241 gnd.n4240 71.676
R8519 gnd.n4234 gnd.n4193 71.676
R8520 gnd.n4233 gnd.n4232 71.676
R8521 gnd.n4226 gnd.n4195 71.676
R8522 gnd.n4225 gnd.n4224 71.676
R8523 gnd.n4218 gnd.n4197 71.676
R8524 gnd.n4217 gnd.n4216 71.676
R8525 gnd.n4210 gnd.n4199 71.676
R8526 gnd.n4209 gnd.n4203 71.676
R8527 gnd.n4205 gnd.n4204 71.676
R8528 gnd.n4344 gnd.n4343 71.676
R8529 gnd.n4336 gnd.n4144 71.676
R8530 gnd.n4335 gnd.n4334 71.676
R8531 gnd.n4328 gnd.n4148 71.676
R8532 gnd.n4327 gnd.n4326 71.676
R8533 gnd.n4320 gnd.n4150 71.676
R8534 gnd.n4319 gnd.n4318 71.676
R8535 gnd.n4312 gnd.n4152 71.676
R8536 gnd.n4311 gnd.n4310 71.676
R8537 gnd.n4304 gnd.n4154 71.676
R8538 gnd.n4303 gnd.n4302 71.676
R8539 gnd.n4296 gnd.n4156 71.676
R8540 gnd.n4295 gnd.n4294 71.676
R8541 gnd.n4288 gnd.n4158 71.676
R8542 gnd.n4287 gnd.n4286 71.676
R8543 gnd.n4280 gnd.n4160 71.676
R8544 gnd.n4263 gnd.n4185 71.676
R8545 gnd.n4258 gnd.n4187 71.676
R8546 gnd.n4256 gnd.n4255 71.676
R8547 gnd.n4251 gnd.n4250 71.676
R8548 gnd.n4248 gnd.n4247 71.676
R8549 gnd.n4243 gnd.n4242 71.676
R8550 gnd.n4240 gnd.n4239 71.676
R8551 gnd.n4235 gnd.n4234 71.676
R8552 gnd.n4232 gnd.n4231 71.676
R8553 gnd.n4227 gnd.n4226 71.676
R8554 gnd.n4224 gnd.n4223 71.676
R8555 gnd.n4219 gnd.n4218 71.676
R8556 gnd.n4216 gnd.n4215 71.676
R8557 gnd.n4211 gnd.n4210 71.676
R8558 gnd.n4206 gnd.n4203 71.676
R8559 gnd.n4346 gnd.n4345 71.676
R8560 gnd.n4343 gnd.n4342 71.676
R8561 gnd.n4337 gnd.n4336 71.676
R8562 gnd.n4334 gnd.n4333 71.676
R8563 gnd.n4329 gnd.n4328 71.676
R8564 gnd.n4326 gnd.n4325 71.676
R8565 gnd.n4321 gnd.n4320 71.676
R8566 gnd.n4318 gnd.n4317 71.676
R8567 gnd.n4313 gnd.n4312 71.676
R8568 gnd.n4310 gnd.n4309 71.676
R8569 gnd.n4305 gnd.n4304 71.676
R8570 gnd.n4302 gnd.n4301 71.676
R8571 gnd.n4297 gnd.n4296 71.676
R8572 gnd.n4294 gnd.n4293 71.676
R8573 gnd.n4289 gnd.n4288 71.676
R8574 gnd.n4286 gnd.n4285 71.676
R8575 gnd.n4281 gnd.n4280 71.676
R8576 gnd.n5166 gnd.n5142 71.676
R8577 gnd.n5170 gnd.n5143 71.676
R8578 gnd.n5174 gnd.n5144 71.676
R8579 gnd.n5178 gnd.n5145 71.676
R8580 gnd.n5182 gnd.n5146 71.676
R8581 gnd.n5186 gnd.n5147 71.676
R8582 gnd.n5190 gnd.n5148 71.676
R8583 gnd.n5194 gnd.n5149 71.676
R8584 gnd.n5198 gnd.n5150 71.676
R8585 gnd.n5202 gnd.n5151 71.676
R8586 gnd.n5206 gnd.n5152 71.676
R8587 gnd.n5210 gnd.n5153 71.676
R8588 gnd.n5214 gnd.n5154 71.676
R8589 gnd.n5218 gnd.n5155 71.676
R8590 gnd.n5223 gnd.n5156 71.676
R8591 gnd.n5227 gnd.n5157 71.676
R8592 gnd.n5141 gnd.n5140 71.676
R8593 gnd.n5136 gnd.n5073 71.676
R8594 gnd.n5131 gnd.n5072 71.676
R8595 gnd.n5127 gnd.n5071 71.676
R8596 gnd.n5123 gnd.n5070 71.676
R8597 gnd.n5119 gnd.n5069 71.676
R8598 gnd.n5115 gnd.n5068 71.676
R8599 gnd.n5111 gnd.n5067 71.676
R8600 gnd.n5107 gnd.n5066 71.676
R8601 gnd.n5103 gnd.n5065 71.676
R8602 gnd.n5099 gnd.n5064 71.676
R8603 gnd.n5095 gnd.n5063 71.676
R8604 gnd.n5091 gnd.n5062 71.676
R8605 gnd.n5087 gnd.n5061 71.676
R8606 gnd.n5083 gnd.n5060 71.676
R8607 gnd.n5079 gnd.n5059 71.676
R8608 gnd.n5058 gnd.n5055 71.676
R8609 gnd.n8 gnd.t3 69.1507
R8610 gnd.n14 gnd.t146 68.4792
R8611 gnd.n13 gnd.t289 68.4792
R8612 gnd.n12 gnd.t295 68.4792
R8613 gnd.n11 gnd.t134 68.4792
R8614 gnd.n10 gnd.t154 68.4792
R8615 gnd.n9 gnd.t14 68.4792
R8616 gnd.n8 gnd.t9 68.4792
R8617 gnd.n6915 gnd.n190 68.412
R8618 gnd.n1743 gnd.n1647 64.369
R8619 gnd.n4339 gnd.n4146 59.5399
R8620 gnd.n5221 gnd.n5160 59.5399
R8621 gnd.n4202 gnd.n4201 59.5399
R8622 gnd.n5133 gnd.n5075 59.5399
R8623 gnd.n4184 gnd.n4183 59.1804
R8624 gnd.n6123 gnd.n871 57.3586
R8625 gnd.n6076 gnd.n2259 57.3586
R8626 gnd.n7280 gnd.n102 57.3586
R8627 gnd.n1398 gnd.t160 56.607
R8628 gnd.n48 gnd.t263 56.607
R8629 gnd.n1367 gnd.t224 56.407
R8630 gnd.n1382 gnd.t201 56.407
R8631 gnd.n17 gnd.t258 56.407
R8632 gnd.n32 gnd.t234 56.407
R8633 gnd.n1411 gnd.t227 55.8337
R8634 gnd.n1380 gnd.t232 55.8337
R8635 gnd.n1395 gnd.t211 55.8337
R8636 gnd.n61 gnd.t241 55.8337
R8637 gnd.n30 gnd.t265 55.8337
R8638 gnd.n45 gnd.t244 55.8337
R8639 gnd.n4171 gnd.n4170 54.358
R8640 gnd.n5047 gnd.n5046 54.358
R8641 gnd.n1398 gnd.n1397 53.0052
R8642 gnd.n1400 gnd.n1399 53.0052
R8643 gnd.n1402 gnd.n1401 53.0052
R8644 gnd.n1404 gnd.n1403 53.0052
R8645 gnd.n1406 gnd.n1405 53.0052
R8646 gnd.n1408 gnd.n1407 53.0052
R8647 gnd.n1410 gnd.n1409 53.0052
R8648 gnd.n1367 gnd.n1366 53.0052
R8649 gnd.n1369 gnd.n1368 53.0052
R8650 gnd.n1371 gnd.n1370 53.0052
R8651 gnd.n1373 gnd.n1372 53.0052
R8652 gnd.n1375 gnd.n1374 53.0052
R8653 gnd.n1377 gnd.n1376 53.0052
R8654 gnd.n1379 gnd.n1378 53.0052
R8655 gnd.n1382 gnd.n1381 53.0052
R8656 gnd.n1384 gnd.n1383 53.0052
R8657 gnd.n1386 gnd.n1385 53.0052
R8658 gnd.n1388 gnd.n1387 53.0052
R8659 gnd.n1390 gnd.n1389 53.0052
R8660 gnd.n1392 gnd.n1391 53.0052
R8661 gnd.n1394 gnd.n1393 53.0052
R8662 gnd.n60 gnd.n59 53.0052
R8663 gnd.n58 gnd.n57 53.0052
R8664 gnd.n56 gnd.n55 53.0052
R8665 gnd.n54 gnd.n53 53.0052
R8666 gnd.n52 gnd.n51 53.0052
R8667 gnd.n50 gnd.n49 53.0052
R8668 gnd.n48 gnd.n47 53.0052
R8669 gnd.n29 gnd.n28 53.0052
R8670 gnd.n27 gnd.n26 53.0052
R8671 gnd.n25 gnd.n24 53.0052
R8672 gnd.n23 gnd.n22 53.0052
R8673 gnd.n21 gnd.n20 53.0052
R8674 gnd.n19 gnd.n18 53.0052
R8675 gnd.n17 gnd.n16 53.0052
R8676 gnd.n44 gnd.n43 53.0052
R8677 gnd.n42 gnd.n41 53.0052
R8678 gnd.n40 gnd.n39 53.0052
R8679 gnd.n38 gnd.n37 53.0052
R8680 gnd.n36 gnd.n35 53.0052
R8681 gnd.n34 gnd.n33 53.0052
R8682 gnd.n32 gnd.n31 53.0052
R8683 gnd.n5038 gnd.n5037 52.4801
R8684 gnd.n1211 gnd.t319 52.3082
R8685 gnd.n1179 gnd.t150 52.3082
R8686 gnd.n1147 gnd.t321 52.3082
R8687 gnd.n1116 gnd.t144 52.3082
R8688 gnd.n1084 gnd.t156 52.3082
R8689 gnd.n1052 gnd.t293 52.3082
R8690 gnd.n1020 gnd.t130 52.3082
R8691 gnd.n989 gnd.t138 52.3082
R8692 gnd.n1041 gnd.n1009 51.4173
R8693 gnd.n1105 gnd.n1104 50.455
R8694 gnd.n1073 gnd.n1072 50.455
R8695 gnd.n1041 gnd.n1040 50.455
R8696 gnd.n5666 gnd.n2741 45.6325
R8697 gnd.n4348 gnd.n4347 45.6325
R8698 gnd.n1690 gnd.n1689 45.1884
R8699 gnd.n901 gnd.n900 45.1884
R8700 gnd.n5054 gnd.n5053 44.3322
R8701 gnd.n4174 gnd.n4173 44.3189
R8702 gnd.n4406 gnd.n3458 42.2793
R8703 gnd.n1691 gnd.n1690 42.2793
R8704 gnd.n902 gnd.n901 42.2793
R8705 gnd.n1617 gnd.n1616 42.2793
R8706 gnd.n881 gnd.n880 42.2793
R8707 gnd.n7156 gnd.n7151 42.2793
R8708 gnd.n3072 gnd.n2968 42.2793
R8709 gnd.n4381 gnd.n3470 42.2793
R8710 gnd.n2768 gnd.n2767 42.2793
R8711 gnd.n7208 gnd.n176 42.2793
R8712 gnd.n7245 gnd.n7244 42.2793
R8713 gnd.n6040 gnd.n2282 42.2793
R8714 gnd.n2305 gnd.n2304 42.2793
R8715 gnd.n4099 gnd.n3635 42.2793
R8716 gnd.n3825 gnd.n3824 42.2793
R8717 gnd.n5417 gnd.n5416 42.2793
R8718 gnd.n4172 gnd.n4171 41.6274
R8719 gnd.n5048 gnd.n5047 41.6274
R8720 gnd.n4181 gnd.n4180 40.8975
R8721 gnd.n5051 gnd.n5050 40.8975
R8722 gnd.n5666 gnd.n2745 36.9518
R8723 gnd.n4348 gnd.n3613 36.9518
R8724 gnd.n6322 gnd.n679 35.4101
R8725 gnd.n6316 gnd.n679 35.4101
R8726 gnd.n6316 gnd.n6315 35.4101
R8727 gnd.n6315 gnd.n6314 35.4101
R8728 gnd.n6314 gnd.n686 35.4101
R8729 gnd.n6308 gnd.n686 35.4101
R8730 gnd.n6308 gnd.n6307 35.4101
R8731 gnd.n6307 gnd.n6306 35.4101
R8732 gnd.n6306 gnd.n694 35.4101
R8733 gnd.n6300 gnd.n694 35.4101
R8734 gnd.n6300 gnd.n6299 35.4101
R8735 gnd.n6299 gnd.n6298 35.4101
R8736 gnd.n6298 gnd.n702 35.4101
R8737 gnd.n6292 gnd.n702 35.4101
R8738 gnd.n6292 gnd.n6291 35.4101
R8739 gnd.n6291 gnd.n6290 35.4101
R8740 gnd.n6290 gnd.n710 35.4101
R8741 gnd.n6284 gnd.n710 35.4101
R8742 gnd.n6284 gnd.n6283 35.4101
R8743 gnd.n6283 gnd.n6282 35.4101
R8744 gnd.n6282 gnd.n718 35.4101
R8745 gnd.n6276 gnd.n718 35.4101
R8746 gnd.n6276 gnd.n6275 35.4101
R8747 gnd.n6275 gnd.n6274 35.4101
R8748 gnd.n6274 gnd.n726 35.4101
R8749 gnd.n6268 gnd.n726 35.4101
R8750 gnd.n6268 gnd.n6267 35.4101
R8751 gnd.n6267 gnd.n6266 35.4101
R8752 gnd.n6266 gnd.n734 35.4101
R8753 gnd.n6260 gnd.n734 35.4101
R8754 gnd.n6260 gnd.n6259 35.4101
R8755 gnd.n6259 gnd.n6258 35.4101
R8756 gnd.n6258 gnd.n742 35.4101
R8757 gnd.n6252 gnd.n742 35.4101
R8758 gnd.n6252 gnd.n6251 35.4101
R8759 gnd.n6251 gnd.n6250 35.4101
R8760 gnd.n6250 gnd.n750 35.4101
R8761 gnd.n6244 gnd.n750 35.4101
R8762 gnd.n6244 gnd.n6243 35.4101
R8763 gnd.n6243 gnd.n6242 35.4101
R8764 gnd.n6242 gnd.n758 35.4101
R8765 gnd.n6236 gnd.n758 35.4101
R8766 gnd.n6236 gnd.n6235 35.4101
R8767 gnd.n6235 gnd.n6234 35.4101
R8768 gnd.n6234 gnd.n766 35.4101
R8769 gnd.n6228 gnd.n766 35.4101
R8770 gnd.n6228 gnd.n6227 35.4101
R8771 gnd.n6227 gnd.n6226 35.4101
R8772 gnd.n6226 gnd.n774 35.4101
R8773 gnd.n6220 gnd.n774 35.4101
R8774 gnd.n6220 gnd.n6219 35.4101
R8775 gnd.n6219 gnd.n6218 35.4101
R8776 gnd.n6218 gnd.n782 35.4101
R8777 gnd.n6212 gnd.n782 35.4101
R8778 gnd.n6212 gnd.n6211 35.4101
R8779 gnd.n6211 gnd.n6210 35.4101
R8780 gnd.n6210 gnd.n790 35.4101
R8781 gnd.n6204 gnd.n790 35.4101
R8782 gnd.n6204 gnd.n6203 35.4101
R8783 gnd.n6203 gnd.n6202 35.4101
R8784 gnd.n6202 gnd.n798 35.4101
R8785 gnd.n6196 gnd.n798 35.4101
R8786 gnd.n6196 gnd.n6195 35.4101
R8787 gnd.n6195 gnd.n6194 35.4101
R8788 gnd.n6194 gnd.n806 35.4101
R8789 gnd.n6188 gnd.n806 35.4101
R8790 gnd.n6188 gnd.n6187 35.4101
R8791 gnd.n6187 gnd.n6186 35.4101
R8792 gnd.n6186 gnd.n814 35.4101
R8793 gnd.n6180 gnd.n814 35.4101
R8794 gnd.n6180 gnd.n6179 35.4101
R8795 gnd.n6179 gnd.n6178 35.4101
R8796 gnd.n6178 gnd.n822 35.4101
R8797 gnd.n6172 gnd.n822 35.4101
R8798 gnd.n6172 gnd.n6171 35.4101
R8799 gnd.n6171 gnd.n6170 35.4101
R8800 gnd.n6170 gnd.n830 35.4101
R8801 gnd.n6164 gnd.n830 35.4101
R8802 gnd.n6164 gnd.n6163 35.4101
R8803 gnd.n6163 gnd.n6162 35.4101
R8804 gnd.n6162 gnd.n838 35.4101
R8805 gnd.n6156 gnd.n838 35.4101
R8806 gnd.n6156 gnd.n6155 35.4101
R8807 gnd.n4180 gnd.n4179 35.055
R8808 gnd.n4175 gnd.n4174 35.055
R8809 gnd.n5040 gnd.n5039 35.055
R8810 gnd.n5050 gnd.n5036 35.055
R8811 gnd.n5164 gnd.n5162 32.9371
R8812 gnd.n4282 gnd.n4161 32.9371
R8813 gnd.n1753 gnd.n1647 31.8661
R8814 gnd.n1753 gnd.n1752 31.8661
R8815 gnd.n1761 gnd.n1636 31.8661
R8816 gnd.n1769 gnd.n1636 31.8661
R8817 gnd.n1769 gnd.n1630 31.8661
R8818 gnd.n1777 gnd.n1630 31.8661
R8819 gnd.n1777 gnd.n1623 31.8661
R8820 gnd.n1815 gnd.n1623 31.8661
R8821 gnd.n1825 gnd.n1556 31.8661
R8822 gnd.n3881 gnd.n2259 31.8661
R8823 gnd.n5989 gnd.n2313 31.8661
R8824 gnd.n5989 gnd.n2315 31.8661
R8825 gnd.n5983 gnd.n2315 31.8661
R8826 gnd.n5983 gnd.n2327 31.8661
R8827 gnd.n5977 gnd.n2338 31.8661
R8828 gnd.n5971 gnd.n2338 31.8661
R8829 gnd.n5965 gnd.n2355 31.8661
R8830 gnd.n5959 gnd.n2365 31.8661
R8831 gnd.n5959 gnd.n2368 31.8661
R8832 gnd.n5953 gnd.n2378 31.8661
R8833 gnd.n5947 gnd.n2378 31.8661
R8834 gnd.n5941 gnd.n2395 31.8661
R8835 gnd.n5935 gnd.n2405 31.8661
R8836 gnd.n3472 gnd.n2572 31.8661
R8837 gnd.n3572 gnd.n3439 31.8661
R8838 gnd.n4415 gnd.n3439 31.8661
R8839 gnd.n4415 gnd.n3432 31.8661
R8840 gnd.n4423 gnd.n3432 31.8661
R8841 gnd.n4423 gnd.n3433 31.8661
R8842 gnd.n5707 gnd.n2682 31.8661
R8843 gnd.n5707 gnd.n5706 31.8661
R8844 gnd.n5706 gnd.n2685 31.8661
R8845 gnd.n5700 gnd.n2685 31.8661
R8846 gnd.n5700 gnd.n5699 31.8661
R8847 gnd.n2772 gnd.n2721 31.8661
R8848 gnd.n7053 gnd.n251 31.8661
R8849 gnd.n7061 gnd.n244 31.8661
R8850 gnd.n7069 gnd.n234 31.8661
R8851 gnd.n7069 gnd.n237 31.8661
R8852 gnd.n7077 gnd.n221 31.8661
R8853 gnd.n7085 gnd.n221 31.8661
R8854 gnd.n7093 gnd.n214 31.8661
R8855 gnd.n7101 gnd.n204 31.8661
R8856 gnd.n7101 gnd.n207 31.8661
R8857 gnd.n7109 gnd.n188 31.8661
R8858 gnd.n7192 gnd.n188 31.8661
R8859 gnd.n7200 gnd.n181 31.8661
R8860 gnd.n7280 gnd.n100 31.8661
R8861 gnd.n190 gnd.n181 30.5915
R8862 gnd.n5965 gnd.t167 27.7236
R8863 gnd.t204 gnd.n214 27.7236
R8864 gnd.n4377 gnd.n3572 27.4049
R8865 gnd.n5699 gnd.n5698 27.4049
R8866 gnd.n5941 gnd.t169 27.0862
R8867 gnd.n5935 gnd.n2408 27.0862
R8868 gnd.n259 gnd.n251 27.0862
R8869 gnd.t248 gnd.n244 27.0862
R8870 gnd.n2395 gnd.t198 25.8116
R8871 gnd.n7061 gnd.t255 25.8116
R8872 gnd.n3458 gnd.n3457 25.7944
R8873 gnd.n1616 gnd.n1615 25.7944
R8874 gnd.n880 gnd.n879 25.7944
R8875 gnd.n7151 gnd.n7150 25.7944
R8876 gnd.n2968 gnd.n2967 25.7944
R8877 gnd.n3470 gnd.n3469 25.7944
R8878 gnd.n2745 gnd.n2744 25.7944
R8879 gnd.n2767 gnd.n2766 25.7944
R8880 gnd.n176 gnd.n175 25.7944
R8881 gnd.n7244 gnd.n7243 25.7944
R8882 gnd.n2282 gnd.n2281 25.7944
R8883 gnd.n2304 gnd.n2303 25.7944
R8884 gnd.n3635 gnd.n3634 25.7944
R8885 gnd.n3613 gnd.n3612 25.7944
R8886 gnd.n3824 gnd.n3823 25.7944
R8887 gnd.n5416 gnd.n5415 25.7944
R8888 gnd.n2355 gnd.t229 25.1743
R8889 gnd.n7093 gnd.t190 25.1743
R8890 gnd.n1837 gnd.n1557 24.8557
R8891 gnd.n1847 gnd.n1540 24.8557
R8892 gnd.n1543 gnd.n1531 24.8557
R8893 gnd.n1868 gnd.n1532 24.8557
R8894 gnd.n1878 gnd.n1512 24.8557
R8895 gnd.n1888 gnd.n1887 24.8557
R8896 gnd.n1498 gnd.n1496 24.8557
R8897 gnd.n1919 gnd.n1918 24.8557
R8898 gnd.n1934 gnd.n1481 24.8557
R8899 gnd.n1988 gnd.n1420 24.8557
R8900 gnd.n1944 gnd.n1421 24.8557
R8901 gnd.n1981 gnd.n1432 24.8557
R8902 gnd.n1470 gnd.n1469 24.8557
R8903 gnd.n1975 gnd.n1974 24.8557
R8904 gnd.n1456 gnd.n1443 24.8557
R8905 gnd.n2014 gnd.n2013 24.8557
R8906 gnd.n2024 gnd.n1352 24.8557
R8907 gnd.n2036 gnd.n1344 24.8557
R8908 gnd.n2035 gnd.n1332 24.8557
R8909 gnd.n2054 gnd.n2053 24.8557
R8910 gnd.n2064 gnd.n1325 24.8557
R8911 gnd.n2075 gnd.n1313 24.8557
R8912 gnd.n2099 gnd.n2098 24.8557
R8913 gnd.n2110 gnd.n1296 24.8557
R8914 gnd.n2109 gnd.n1298 24.8557
R8915 gnd.n2121 gnd.n1289 24.8557
R8916 gnd.n2139 gnd.n2138 24.8557
R8917 gnd.n1280 gnd.n1269 24.8557
R8918 gnd.n2162 gnd.n1257 24.8557
R8919 gnd.n2186 gnd.n2185 24.8557
R8920 gnd.n2201 gnd.n1243 24.8557
R8921 gnd.n2175 gnd.n848 24.8557
R8922 gnd.n6147 gnd.n857 24.8557
R8923 gnd.n6140 gnd.n6139 24.8557
R8924 gnd.n4146 gnd.n4145 23.855
R8925 gnd.n5160 gnd.n5159 23.855
R8926 gnd.n4201 gnd.n4200 23.855
R8927 gnd.n5075 gnd.n5074 23.855
R8928 gnd.n1858 gnd.t137 23.2624
R8929 gnd.n3427 gnd.n3426 23.2624
R8930 gnd.n5230 gnd.n5229 23.2624
R8931 gnd.n1559 gnd.t23 22.6251
R8932 gnd.n3881 gnd.t72 22.6251
R8933 gnd.t30 gnd.n100 22.6251
R8934 gnd.n4555 gnd.n3396 21.6691
R8935 gnd.n4547 gnd.n3387 21.6691
R8936 gnd.n4532 gnd.n3373 21.6691
R8937 gnd.n4517 gnd.n3358 21.6691
R8938 gnd.n4510 gnd.n3352 21.6691
R8939 gnd.n4728 gnd.n3320 21.6691
R8940 gnd.n4713 gnd.n3305 21.6691
R8941 gnd.n4705 gnd.n3298 21.6691
R8942 gnd.n4698 gnd.n3292 21.6691
R8943 gnd.n4690 gnd.n4656 21.6691
R8944 gnd.n4684 gnd.n4683 21.6691
R8945 gnd.n4899 gnd.n3247 21.6691
R8946 gnd.n4899 gnd.n3250 21.6691
R8947 gnd.n4884 gnd.n3233 21.6691
R8948 gnd.n4876 gnd.n3226 21.6691
R8949 gnd.n4869 gnd.n3218 21.6691
R8950 gnd.n4861 gnd.n3211 21.6691
R8951 gnd.n4855 gnd.n4854 21.6691
R8952 gnd.n5305 gnd.n3172 21.6691
R8953 gnd.n5290 gnd.n3159 21.6691
R8954 gnd.n5282 gnd.n3153 21.6691
R8955 gnd.n5267 gnd.n3139 21.6691
R8956 gnd.n5251 gnd.n3126 21.6691
R8957 gnd.n5237 gnd.n3104 21.6691
R8958 gnd.t143 gnd.n1564 21.3504
R8959 gnd.n6155 gnd.n6154 21.2463
R8960 gnd.n5929 gnd.n2418 21.0318
R8961 gnd.n3976 gnd.n2424 21.0318
R8962 gnd.n3986 gnd.n2434 21.0318
R8963 gnd.n5917 gnd.n2437 21.0318
R8964 gnd.n3995 gnd.n2442 21.0318
R8965 gnd.n5910 gnd.n2445 21.0318
R8966 gnd.n5904 gnd.n2456 21.0318
R8967 gnd.n4011 gnd.n2463 21.0318
R8968 gnd.n4019 gnd.n2473 21.0318
R8969 gnd.n5892 gnd.n2476 21.0318
R8970 gnd.n4027 gnd.n2484 21.0318
R8971 gnd.n5886 gnd.n2487 21.0318
R8972 gnd.n5880 gnd.n2498 21.0318
R8973 gnd.n4043 gnd.n2506 21.0318
R8974 gnd.n4051 gnd.n2516 21.0318
R8975 gnd.n5868 gnd.n2519 21.0318
R8976 gnd.n4059 gnd.n2527 21.0318
R8977 gnd.n5862 gnd.n2530 21.0318
R8978 gnd.n5856 gnd.n2541 21.0318
R8979 gnd.n4075 gnd.n2549 21.0318
R8980 gnd.n5850 gnd.n2552 21.0318
R8981 gnd.n4084 gnd.n2560 21.0318
R8982 gnd.n4092 gnd.n2569 21.0318
R8983 gnd.n5838 gnd.n2572 21.0318
R8984 gnd.n5622 gnd.n2772 21.0318
R8985 gnd.n2923 gnd.n2774 21.0318
R8986 gnd.n5447 gnd.n2901 21.0318
R8987 gnd.n5446 gnd.n2904 21.0318
R8988 gnd.n5457 gnd.n2891 21.0318
R8989 gnd.n2893 gnd.n2883 21.0318
R8990 gnd.n5478 gnd.n2872 21.0318
R8991 gnd.n5477 gnd.n2876 21.0318
R8992 gnd.n5488 gnd.n2863 21.0318
R8993 gnd.n2865 gnd.n2855 21.0318
R8994 gnd.n5515 gnd.n2844 21.0318
R8995 gnd.n5513 gnd.n2847 21.0318
R8996 gnd.n2837 gnd.n2821 21.0318
R8997 gnd.n5561 gnd.n5560 21.0318
R8998 gnd.n5579 gnd.n2810 21.0318
R8999 gnd.n5578 gnd.n2813 21.0318
R9000 gnd.n5548 gnd.n2804 21.0318
R9001 gnd.n7038 gnd.n272 21.0318
R9002 gnd.n6938 gnd.n308 21.0318
R9003 gnd.n6947 gnd.n302 21.0318
R9004 gnd.n6952 gnd.n297 21.0318
R9005 gnd.n6929 gnd.n299 21.0318
R9006 gnd.n7022 gnd.n289 21.0318
R9007 gnd.n7011 gnd.n291 21.0318
R9008 gnd.n4268 gnd.n4184 20.7615
R9009 gnd.n5233 gnd.n5054 20.7615
R9010 gnd.t302 gnd.n1270 20.7131
R9011 gnd.t27 gnd.n3418 20.3945
R9012 gnd.n4162 gnd.n3410 20.3945
R9013 gnd.n4563 gnd.n3386 20.3945
R9014 gnd.n4496 gnd.n3334 20.3945
R9015 gnd.n4736 gnd.n3311 20.3945
R9016 gnd.n4796 gnd.n3264 20.3945
R9017 gnd.n4907 gnd.n3239 20.3945
R9018 gnd.n4967 gnd.n3187 20.3945
R9019 gnd.n5313 gnd.n3165 20.3945
R9020 gnd.t304 gnd.n1305 20.0758
R9021 gnd.t51 gnd.t145 20.0758
R9022 gnd.n4168 gnd.t123 19.8005
R9023 gnd.n4168 gnd.t35 19.8005
R9024 gnd.n4169 gnd.t28 19.8005
R9025 gnd.n4169 gnd.t56 19.8005
R9026 gnd.n5044 gnd.t77 19.8005
R9027 gnd.n5044 gnd.t45 19.8005
R9028 gnd.n5045 gnd.t90 19.8005
R9029 gnd.n5045 gnd.t21 19.8005
R9030 gnd.n4165 gnd.n4164 19.5087
R9031 gnd.n4178 gnd.n4165 19.5087
R9032 gnd.n4176 gnd.n4167 19.5087
R9033 gnd.n5049 gnd.n5043 19.5087
R9034 gnd.n2025 gnd.t310 19.4385
R9035 gnd.n4425 gnd.n3429 19.3944
R9036 gnd.n4429 gnd.n3429 19.3944
R9037 gnd.n4429 gnd.n3415 19.3944
R9038 gnd.n4443 gnd.n3415 19.3944
R9039 gnd.n4443 gnd.n3412 19.3944
R9040 gnd.n4448 gnd.n3412 19.3944
R9041 gnd.n4448 gnd.n3413 19.3944
R9042 gnd.n3413 gnd.n3384 19.3944
R9043 gnd.n4565 gnd.n3384 19.3944
R9044 gnd.n4565 gnd.n3382 19.3944
R9045 gnd.n4569 gnd.n3382 19.3944
R9046 gnd.n4569 gnd.n3370 19.3944
R9047 gnd.n4581 gnd.n3370 19.3944
R9048 gnd.n4581 gnd.n3368 19.3944
R9049 gnd.n4585 gnd.n3368 19.3944
R9050 gnd.n4585 gnd.n3356 19.3944
R9051 gnd.n4597 gnd.n3356 19.3944
R9052 gnd.n4597 gnd.n3354 19.3944
R9053 gnd.n4601 gnd.n3354 19.3944
R9054 gnd.n4601 gnd.n3340 19.3944
R9055 gnd.n4614 gnd.n3340 19.3944
R9056 gnd.n4614 gnd.n3337 19.3944
R9057 gnd.n4619 gnd.n3337 19.3944
R9058 gnd.n4619 gnd.n3338 19.3944
R9059 gnd.n3338 gnd.n3309 19.3944
R9060 gnd.n4738 gnd.n3309 19.3944
R9061 gnd.n4738 gnd.n3307 19.3944
R9062 gnd.n4742 gnd.n3307 19.3944
R9063 gnd.n4742 gnd.n3296 19.3944
R9064 gnd.n4754 gnd.n3296 19.3944
R9065 gnd.n4754 gnd.n3294 19.3944
R9066 gnd.n4758 gnd.n3294 19.3944
R9067 gnd.n4758 gnd.n3284 19.3944
R9068 gnd.n4770 gnd.n3284 19.3944
R9069 gnd.n4770 gnd.n3282 19.3944
R9070 gnd.n4774 gnd.n3282 19.3944
R9071 gnd.n4774 gnd.n3270 19.3944
R9072 gnd.n4788 gnd.n3270 19.3944
R9073 gnd.n4788 gnd.n3267 19.3944
R9074 gnd.n4793 gnd.n3267 19.3944
R9075 gnd.n4793 gnd.n3268 19.3944
R9076 gnd.n3268 gnd.n3237 19.3944
R9077 gnd.n4909 gnd.n3237 19.3944
R9078 gnd.n4909 gnd.n3235 19.3944
R9079 gnd.n4913 gnd.n3235 19.3944
R9080 gnd.n4913 gnd.n3222 19.3944
R9081 gnd.n4925 gnd.n3222 19.3944
R9082 gnd.n4925 gnd.n3220 19.3944
R9083 gnd.n4929 gnd.n3220 19.3944
R9084 gnd.n4929 gnd.n3208 19.3944
R9085 gnd.n4941 gnd.n3208 19.3944
R9086 gnd.n4941 gnd.n3206 19.3944
R9087 gnd.n4945 gnd.n3206 19.3944
R9088 gnd.n4945 gnd.n3193 19.3944
R9089 gnd.n4959 gnd.n3193 19.3944
R9090 gnd.n4959 gnd.n3190 19.3944
R9091 gnd.n4964 gnd.n3190 19.3944
R9092 gnd.n4964 gnd.n3191 19.3944
R9093 gnd.n3191 gnd.n3163 19.3944
R9094 gnd.n5315 gnd.n3163 19.3944
R9095 gnd.n5315 gnd.n3161 19.3944
R9096 gnd.n5319 gnd.n3161 19.3944
R9097 gnd.n5319 gnd.n3150 19.3944
R9098 gnd.n5331 gnd.n3150 19.3944
R9099 gnd.n5331 gnd.n3148 19.3944
R9100 gnd.n5335 gnd.n3148 19.3944
R9101 gnd.n5335 gnd.n3137 19.3944
R9102 gnd.n5347 gnd.n3137 19.3944
R9103 gnd.n5347 gnd.n3135 19.3944
R9104 gnd.n5351 gnd.n3135 19.3944
R9105 gnd.n5351 gnd.n3123 19.3944
R9106 gnd.n5363 gnd.n3123 19.3944
R9107 gnd.n5363 gnd.n3121 19.3944
R9108 gnd.n5367 gnd.n3121 19.3944
R9109 gnd.n5367 gnd.n3109 19.3944
R9110 gnd.n5379 gnd.n3109 19.3944
R9111 gnd.n5379 gnd.n3106 19.3944
R9112 gnd.n5385 gnd.n3106 19.3944
R9113 gnd.n5385 gnd.n3107 19.3944
R9114 gnd.n3107 gnd.n3096 19.3944
R9115 gnd.n5401 gnd.n3096 19.3944
R9116 gnd.n5402 gnd.n5401 19.3944
R9117 gnd.n4408 gnd.n3454 19.3944
R9118 gnd.n4412 gnd.n3454 19.3944
R9119 gnd.n4412 gnd.n3455 19.3944
R9120 gnd.n3515 gnd.n3512 19.3944
R9121 gnd.n3515 gnd.n3502 19.3944
R9122 gnd.n3524 gnd.n3502 19.3944
R9123 gnd.n3527 gnd.n3524 19.3944
R9124 gnd.n3527 gnd.n3496 19.3944
R9125 gnd.n3536 gnd.n3496 19.3944
R9126 gnd.n3539 gnd.n3536 19.3944
R9127 gnd.n3539 gnd.n3490 19.3944
R9128 gnd.n3548 gnd.n3490 19.3944
R9129 gnd.n3551 gnd.n3548 19.3944
R9130 gnd.n3551 gnd.n3484 19.3944
R9131 gnd.n3561 gnd.n3484 19.3944
R9132 gnd.n3562 gnd.n3561 19.3944
R9133 gnd.n3565 gnd.n3562 19.3944
R9134 gnd.n3565 gnd.n3464 19.3944
R9135 gnd.n4384 gnd.n3464 19.3944
R9136 gnd.n4387 gnd.n4384 19.3944
R9137 gnd.n4387 gnd.n3461 19.3944
R9138 gnd.n4392 gnd.n3461 19.3944
R9139 gnd.n4395 gnd.n4392 19.3944
R9140 gnd.n4398 gnd.n4395 19.3944
R9141 gnd.n4398 gnd.n3459 19.3944
R9142 gnd.n4402 gnd.n3459 19.3944
R9143 gnd.n4405 gnd.n4402 19.3944
R9144 gnd.n1740 gnd.n1739 19.3944
R9145 gnd.n1739 gnd.n1738 19.3944
R9146 gnd.n1738 gnd.n1737 19.3944
R9147 gnd.n1737 gnd.n1735 19.3944
R9148 gnd.n1735 gnd.n1732 19.3944
R9149 gnd.n1732 gnd.n1731 19.3944
R9150 gnd.n1731 gnd.n1728 19.3944
R9151 gnd.n1728 gnd.n1727 19.3944
R9152 gnd.n1727 gnd.n1724 19.3944
R9153 gnd.n1724 gnd.n1723 19.3944
R9154 gnd.n1723 gnd.n1720 19.3944
R9155 gnd.n1720 gnd.n1719 19.3944
R9156 gnd.n1719 gnd.n1716 19.3944
R9157 gnd.n1716 gnd.n1715 19.3944
R9158 gnd.n1715 gnd.n1712 19.3944
R9159 gnd.n1712 gnd.n1711 19.3944
R9160 gnd.n1711 gnd.n1708 19.3944
R9161 gnd.n1708 gnd.n1707 19.3944
R9162 gnd.n1707 gnd.n1704 19.3944
R9163 gnd.n1704 gnd.n1703 19.3944
R9164 gnd.n1703 gnd.n1700 19.3944
R9165 gnd.n1700 gnd.n1699 19.3944
R9166 gnd.n1696 gnd.n1695 19.3944
R9167 gnd.n1695 gnd.n1651 19.3944
R9168 gnd.n1746 gnd.n1651 19.3944
R9169 gnd.n974 gnd.n972 19.3944
R9170 gnd.n974 gnd.n898 19.3944
R9171 gnd.n2228 gnd.n898 19.3944
R9172 gnd.n915 gnd.n914 19.3944
R9173 gnd.n919 gnd.n914 19.3944
R9174 gnd.n922 gnd.n919 19.3944
R9175 gnd.n925 gnd.n922 19.3944
R9176 gnd.n925 gnd.n911 19.3944
R9177 gnd.n929 gnd.n911 19.3944
R9178 gnd.n932 gnd.n929 19.3944
R9179 gnd.n935 gnd.n932 19.3944
R9180 gnd.n935 gnd.n909 19.3944
R9181 gnd.n939 gnd.n909 19.3944
R9182 gnd.n942 gnd.n939 19.3944
R9183 gnd.n945 gnd.n942 19.3944
R9184 gnd.n945 gnd.n907 19.3944
R9185 gnd.n949 gnd.n907 19.3944
R9186 gnd.n952 gnd.n949 19.3944
R9187 gnd.n955 gnd.n952 19.3944
R9188 gnd.n955 gnd.n905 19.3944
R9189 gnd.n959 gnd.n905 19.3944
R9190 gnd.n962 gnd.n959 19.3944
R9191 gnd.n965 gnd.n962 19.3944
R9192 gnd.n965 gnd.n903 19.3944
R9193 gnd.n969 gnd.n903 19.3944
R9194 gnd.n1839 gnd.n1548 19.3944
R9195 gnd.n1849 gnd.n1548 19.3944
R9196 gnd.n1850 gnd.n1849 19.3944
R9197 gnd.n1850 gnd.n1529 19.3944
R9198 gnd.n1870 gnd.n1529 19.3944
R9199 gnd.n1870 gnd.n1521 19.3944
R9200 gnd.n1880 gnd.n1521 19.3944
R9201 gnd.n1881 gnd.n1880 19.3944
R9202 gnd.n1882 gnd.n1881 19.3944
R9203 gnd.n1882 gnd.n1504 19.3944
R9204 gnd.n1899 gnd.n1504 19.3944
R9205 gnd.n1902 gnd.n1899 19.3944
R9206 gnd.n1902 gnd.n1901 19.3944
R9207 gnd.n1901 gnd.n1477 19.3944
R9208 gnd.n1941 gnd.n1477 19.3944
R9209 gnd.n1941 gnd.n1474 19.3944
R9210 gnd.n1947 gnd.n1474 19.3944
R9211 gnd.n1948 gnd.n1947 19.3944
R9212 gnd.n1948 gnd.n1472 19.3944
R9213 gnd.n1954 gnd.n1472 19.3944
R9214 gnd.n1957 gnd.n1954 19.3944
R9215 gnd.n1959 gnd.n1957 19.3944
R9216 gnd.n1965 gnd.n1959 19.3944
R9217 gnd.n1965 gnd.n1964 19.3944
R9218 gnd.n1964 gnd.n1347 19.3944
R9219 gnd.n2031 gnd.n1347 19.3944
R9220 gnd.n2032 gnd.n2031 19.3944
R9221 gnd.n2032 gnd.n1340 19.3944
R9222 gnd.n2043 gnd.n1340 19.3944
R9223 gnd.n2044 gnd.n2043 19.3944
R9224 gnd.n2044 gnd.n1323 19.3944
R9225 gnd.n1323 gnd.n1321 19.3944
R9226 gnd.n2068 gnd.n1321 19.3944
R9227 gnd.n2069 gnd.n2068 19.3944
R9228 gnd.n2069 gnd.n1292 19.3944
R9229 gnd.n2116 gnd.n1292 19.3944
R9230 gnd.n2117 gnd.n2116 19.3944
R9231 gnd.n2117 gnd.n1285 19.3944
R9232 gnd.n2128 gnd.n1285 19.3944
R9233 gnd.n2129 gnd.n2128 19.3944
R9234 gnd.n2129 gnd.n1268 19.3944
R9235 gnd.n1268 gnd.n1266 19.3944
R9236 gnd.n2153 gnd.n1266 19.3944
R9237 gnd.n2156 gnd.n2153 19.3944
R9238 gnd.n2156 gnd.n2155 19.3944
R9239 gnd.n2155 gnd.n1239 19.3944
R9240 gnd.n2208 gnd.n1239 19.3944
R9241 gnd.n2208 gnd.n1236 19.3944
R9242 gnd.n2212 gnd.n1236 19.3944
R9243 gnd.n2213 gnd.n2212 19.3944
R9244 gnd.n2218 gnd.n2213 19.3944
R9245 gnd.n2218 gnd.n877 19.3944
R9246 gnd.n6134 gnd.n877 19.3944
R9247 gnd.n1830 gnd.n1829 19.3944
R9248 gnd.n1829 gnd.n1562 19.3944
R9249 gnd.n1585 gnd.n1562 19.3944
R9250 gnd.n1588 gnd.n1585 19.3944
R9251 gnd.n1588 gnd.n1581 19.3944
R9252 gnd.n1592 gnd.n1581 19.3944
R9253 gnd.n1595 gnd.n1592 19.3944
R9254 gnd.n1598 gnd.n1595 19.3944
R9255 gnd.n1598 gnd.n1579 19.3944
R9256 gnd.n1602 gnd.n1579 19.3944
R9257 gnd.n1605 gnd.n1602 19.3944
R9258 gnd.n1608 gnd.n1605 19.3944
R9259 gnd.n1608 gnd.n1577 19.3944
R9260 gnd.n1612 gnd.n1577 19.3944
R9261 gnd.n1835 gnd.n1834 19.3944
R9262 gnd.n1834 gnd.n1538 19.3944
R9263 gnd.n1860 gnd.n1538 19.3944
R9264 gnd.n1860 gnd.n1536 19.3944
R9265 gnd.n1866 gnd.n1536 19.3944
R9266 gnd.n1866 gnd.n1865 19.3944
R9267 gnd.n1865 gnd.n1510 19.3944
R9268 gnd.n1890 gnd.n1510 19.3944
R9269 gnd.n1890 gnd.n1508 19.3944
R9270 gnd.n1894 gnd.n1508 19.3944
R9271 gnd.n1894 gnd.n1488 19.3944
R9272 gnd.n1921 gnd.n1488 19.3944
R9273 gnd.n1921 gnd.n1486 19.3944
R9274 gnd.n1931 gnd.n1486 19.3944
R9275 gnd.n1931 gnd.n1930 19.3944
R9276 gnd.n1930 gnd.n1929 19.3944
R9277 gnd.n1929 gnd.n1435 19.3944
R9278 gnd.n1979 gnd.n1435 19.3944
R9279 gnd.n1979 gnd.n1978 19.3944
R9280 gnd.n1978 gnd.n1977 19.3944
R9281 gnd.n1977 gnd.n1439 19.3944
R9282 gnd.n1459 gnd.n1439 19.3944
R9283 gnd.n1459 gnd.n1357 19.3944
R9284 gnd.n2016 gnd.n1357 19.3944
R9285 gnd.n2016 gnd.n1355 19.3944
R9286 gnd.n2022 gnd.n1355 19.3944
R9287 gnd.n2022 gnd.n2021 19.3944
R9288 gnd.n2021 gnd.n1330 19.3944
R9289 gnd.n2056 gnd.n1330 19.3944
R9290 gnd.n2056 gnd.n1328 19.3944
R9291 gnd.n2062 gnd.n1328 19.3944
R9292 gnd.n2062 gnd.n2061 19.3944
R9293 gnd.n2061 gnd.n1303 19.3944
R9294 gnd.n2101 gnd.n1303 19.3944
R9295 gnd.n2101 gnd.n1301 19.3944
R9296 gnd.n2107 gnd.n1301 19.3944
R9297 gnd.n2107 gnd.n2106 19.3944
R9298 gnd.n2106 gnd.n1275 19.3944
R9299 gnd.n2141 gnd.n1275 19.3944
R9300 gnd.n2141 gnd.n1273 19.3944
R9301 gnd.n2147 gnd.n1273 19.3944
R9302 gnd.n2147 gnd.n2146 19.3944
R9303 gnd.n2146 gnd.n1249 19.3944
R9304 gnd.n2188 gnd.n1249 19.3944
R9305 gnd.n2188 gnd.n1247 19.3944
R9306 gnd.n2198 gnd.n1247 19.3944
R9307 gnd.n2198 gnd.n2197 19.3944
R9308 gnd.n2197 gnd.n2196 19.3944
R9309 gnd.n2196 gnd.n862 19.3944
R9310 gnd.n6144 gnd.n862 19.3944
R9311 gnd.n6144 gnd.n6143 19.3944
R9312 gnd.n6143 gnd.n6142 19.3944
R9313 gnd.n6142 gnd.n866 19.3944
R9314 gnd.n6121 gnd.n6120 19.3944
R9315 gnd.n6120 gnd.n6086 19.3944
R9316 gnd.n6116 gnd.n6086 19.3944
R9317 gnd.n6116 gnd.n6113 19.3944
R9318 gnd.n6113 gnd.n6110 19.3944
R9319 gnd.n6110 gnd.n6109 19.3944
R9320 gnd.n6109 gnd.n6106 19.3944
R9321 gnd.n6106 gnd.n6105 19.3944
R9322 gnd.n6105 gnd.n6102 19.3944
R9323 gnd.n6102 gnd.n6101 19.3944
R9324 gnd.n6101 gnd.n6098 19.3944
R9325 gnd.n6098 gnd.n6097 19.3944
R9326 gnd.n6097 gnd.n883 19.3944
R9327 gnd.n6127 gnd.n883 19.3944
R9328 gnd.n1750 gnd.n1649 19.3944
R9329 gnd.n1750 gnd.n1640 19.3944
R9330 gnd.n1763 gnd.n1640 19.3944
R9331 gnd.n1763 gnd.n1638 19.3944
R9332 gnd.n1767 gnd.n1638 19.3944
R9333 gnd.n1767 gnd.n1628 19.3944
R9334 gnd.n1779 gnd.n1628 19.3944
R9335 gnd.n1779 gnd.n1626 19.3944
R9336 gnd.n1813 gnd.n1626 19.3944
R9337 gnd.n1813 gnd.n1812 19.3944
R9338 gnd.n1812 gnd.n1811 19.3944
R9339 gnd.n1811 gnd.n1810 19.3944
R9340 gnd.n1810 gnd.n1807 19.3944
R9341 gnd.n1807 gnd.n1806 19.3944
R9342 gnd.n1806 gnd.n1805 19.3944
R9343 gnd.n1805 gnd.n1803 19.3944
R9344 gnd.n1803 gnd.n1802 19.3944
R9345 gnd.n1802 gnd.n1799 19.3944
R9346 gnd.n1799 gnd.n1798 19.3944
R9347 gnd.n1798 gnd.n1797 19.3944
R9348 gnd.n1797 gnd.n1795 19.3944
R9349 gnd.n1795 gnd.n1494 19.3944
R9350 gnd.n1910 gnd.n1494 19.3944
R9351 gnd.n1910 gnd.n1492 19.3944
R9352 gnd.n1916 gnd.n1492 19.3944
R9353 gnd.n1916 gnd.n1915 19.3944
R9354 gnd.n1915 gnd.n1416 19.3944
R9355 gnd.n1990 gnd.n1416 19.3944
R9356 gnd.n1990 gnd.n1417 19.3944
R9357 gnd.n1464 gnd.n1463 19.3944
R9358 gnd.n1467 gnd.n1466 19.3944
R9359 gnd.n1454 gnd.n1453 19.3944
R9360 gnd.n2009 gnd.n1362 19.3944
R9361 gnd.n2009 gnd.n2008 19.3944
R9362 gnd.n2008 gnd.n2007 19.3944
R9363 gnd.n2007 gnd.n2005 19.3944
R9364 gnd.n2005 gnd.n2004 19.3944
R9365 gnd.n2004 gnd.n2002 19.3944
R9366 gnd.n2002 gnd.n2001 19.3944
R9367 gnd.n2001 gnd.n1311 19.3944
R9368 gnd.n2077 gnd.n1311 19.3944
R9369 gnd.n2077 gnd.n1309 19.3944
R9370 gnd.n2096 gnd.n1309 19.3944
R9371 gnd.n2096 gnd.n2095 19.3944
R9372 gnd.n2095 gnd.n2094 19.3944
R9373 gnd.n2094 gnd.n2092 19.3944
R9374 gnd.n2092 gnd.n2091 19.3944
R9375 gnd.n2091 gnd.n2089 19.3944
R9376 gnd.n2089 gnd.n2088 19.3944
R9377 gnd.n2088 gnd.n1255 19.3944
R9378 gnd.n2164 gnd.n1255 19.3944
R9379 gnd.n2164 gnd.n1253 19.3944
R9380 gnd.n2183 gnd.n1253 19.3944
R9381 gnd.n2183 gnd.n2182 19.3944
R9382 gnd.n2182 gnd.n2181 19.3944
R9383 gnd.n2181 gnd.n2178 19.3944
R9384 gnd.n2178 gnd.n2177 19.3944
R9385 gnd.n2177 gnd.n2174 19.3944
R9386 gnd.n2174 gnd.n978 19.3944
R9387 gnd.n2224 gnd.n978 19.3944
R9388 gnd.n2225 gnd.n2224 19.3944
R9389 gnd.n1755 gnd.n1645 19.3944
R9390 gnd.n1755 gnd.n1643 19.3944
R9391 gnd.n1759 gnd.n1643 19.3944
R9392 gnd.n1759 gnd.n1634 19.3944
R9393 gnd.n1771 gnd.n1634 19.3944
R9394 gnd.n1771 gnd.n1632 19.3944
R9395 gnd.n1775 gnd.n1632 19.3944
R9396 gnd.n1775 gnd.n1621 19.3944
R9397 gnd.n1817 gnd.n1621 19.3944
R9398 gnd.n1817 gnd.n1575 19.3944
R9399 gnd.n1823 gnd.n1575 19.3944
R9400 gnd.n1823 gnd.n1822 19.3944
R9401 gnd.n1822 gnd.n1553 19.3944
R9402 gnd.n1844 gnd.n1553 19.3944
R9403 gnd.n1844 gnd.n1546 19.3944
R9404 gnd.n1855 gnd.n1546 19.3944
R9405 gnd.n1855 gnd.n1854 19.3944
R9406 gnd.n1854 gnd.n1527 19.3944
R9407 gnd.n1875 gnd.n1527 19.3944
R9408 gnd.n1875 gnd.n1517 19.3944
R9409 gnd.n1885 gnd.n1517 19.3944
R9410 gnd.n1885 gnd.n1500 19.3944
R9411 gnd.n1906 gnd.n1500 19.3944
R9412 gnd.n1906 gnd.n1905 19.3944
R9413 gnd.n1905 gnd.n1479 19.3944
R9414 gnd.n1936 gnd.n1479 19.3944
R9415 gnd.n1936 gnd.n1424 19.3944
R9416 gnd.n1986 gnd.n1424 19.3944
R9417 gnd.n1986 gnd.n1985 19.3944
R9418 gnd.n1985 gnd.n1984 19.3944
R9419 gnd.n1984 gnd.n1428 19.3944
R9420 gnd.n1446 gnd.n1428 19.3944
R9421 gnd.n1972 gnd.n1446 19.3944
R9422 gnd.n1972 gnd.n1971 19.3944
R9423 gnd.n1971 gnd.n1970 19.3944
R9424 gnd.n1970 gnd.n1450 19.3944
R9425 gnd.n1450 gnd.n1349 19.3944
R9426 gnd.n2027 gnd.n1349 19.3944
R9427 gnd.n2027 gnd.n1342 19.3944
R9428 gnd.n2038 gnd.n1342 19.3944
R9429 gnd.n2038 gnd.n1338 19.3944
R9430 gnd.n2051 gnd.n1338 19.3944
R9431 gnd.n2051 gnd.n2050 19.3944
R9432 gnd.n2050 gnd.n1317 19.3944
R9433 gnd.n2073 gnd.n1317 19.3944
R9434 gnd.n2073 gnd.n2072 19.3944
R9435 gnd.n2072 gnd.n1294 19.3944
R9436 gnd.n2112 gnd.n1294 19.3944
R9437 gnd.n2112 gnd.n1287 19.3944
R9438 gnd.n2123 gnd.n1287 19.3944
R9439 gnd.n2123 gnd.n1283 19.3944
R9440 gnd.n2136 gnd.n1283 19.3944
R9441 gnd.n2136 gnd.n2135 19.3944
R9442 gnd.n2135 gnd.n1262 19.3944
R9443 gnd.n2160 gnd.n1262 19.3944
R9444 gnd.n2160 gnd.n2159 19.3944
R9445 gnd.n2159 gnd.n1241 19.3944
R9446 gnd.n2203 gnd.n1241 19.3944
R9447 gnd.n2203 gnd.n851 19.3944
R9448 gnd.n6151 gnd.n851 19.3944
R9449 gnd.n6151 gnd.n6150 19.3944
R9450 gnd.n6150 gnd.n6149 19.3944
R9451 gnd.n6149 gnd.n855 19.3944
R9452 gnd.n874 gnd.n855 19.3944
R9453 gnd.n6137 gnd.n874 19.3944
R9454 gnd.n5428 gnd.n2956 19.3944
R9455 gnd.n5433 gnd.n2956 19.3944
R9456 gnd.n5433 gnd.n2957 19.3944
R9457 gnd.n2957 gnd.n2889 19.3944
R9458 gnd.n5459 gnd.n2889 19.3944
R9459 gnd.n5459 gnd.n2886 19.3944
R9460 gnd.n5464 gnd.n2886 19.3944
R9461 gnd.n5464 gnd.n2887 19.3944
R9462 gnd.n2887 gnd.n2861 19.3944
R9463 gnd.n5490 gnd.n2861 19.3944
R9464 gnd.n5490 gnd.n2858 19.3944
R9465 gnd.n5500 gnd.n2858 19.3944
R9466 gnd.n5500 gnd.n2859 19.3944
R9467 gnd.n5496 gnd.n2859 19.3944
R9468 gnd.n5496 gnd.n5495 19.3944
R9469 gnd.n5495 gnd.n2824 19.3944
R9470 gnd.n5557 gnd.n2824 19.3944
R9471 gnd.n5557 gnd.n2825 19.3944
R9472 gnd.n5553 gnd.n2825 19.3944
R9473 gnd.n5553 gnd.n5552 19.3944
R9474 gnd.n5552 gnd.n5551 19.3944
R9475 gnd.n5551 gnd.n306 19.3944
R9476 gnd.n6941 gnd.n306 19.3944
R9477 gnd.n6941 gnd.n304 19.3944
R9478 gnd.n6945 gnd.n304 19.3944
R9479 gnd.n6945 gnd.n65 19.3944
R9480 gnd.n7320 gnd.n65 19.3944
R9481 gnd.n7320 gnd.n7319 19.3944
R9482 gnd.n7319 gnd.n7318 19.3944
R9483 gnd.n7318 gnd.n69 19.3944
R9484 gnd.n7314 gnd.n69 19.3944
R9485 gnd.n7314 gnd.n7313 19.3944
R9486 gnd.n7313 gnd.n7312 19.3944
R9487 gnd.n7312 gnd.n74 19.3944
R9488 gnd.n7308 gnd.n74 19.3944
R9489 gnd.n7308 gnd.n7307 19.3944
R9490 gnd.n7307 gnd.n7306 19.3944
R9491 gnd.n7306 gnd.n79 19.3944
R9492 gnd.n7302 gnd.n79 19.3944
R9493 gnd.n7302 gnd.n7301 19.3944
R9494 gnd.n7301 gnd.n7300 19.3944
R9495 gnd.n7300 gnd.n84 19.3944
R9496 gnd.n7296 gnd.n84 19.3944
R9497 gnd.n7296 gnd.n7295 19.3944
R9498 gnd.n7295 gnd.n7294 19.3944
R9499 gnd.n7294 gnd.n89 19.3944
R9500 gnd.n7290 gnd.n89 19.3944
R9501 gnd.n7290 gnd.n7289 19.3944
R9502 gnd.n7289 gnd.n7288 19.3944
R9503 gnd.n7288 gnd.n94 19.3944
R9504 gnd.n7284 gnd.n94 19.3944
R9505 gnd.n7284 gnd.n7283 19.3944
R9506 gnd.n7283 gnd.n7282 19.3944
R9507 gnd.n7181 gnd.n7180 19.3944
R9508 gnd.n7180 gnd.n7179 19.3944
R9509 gnd.n7179 gnd.n7121 19.3944
R9510 gnd.n7175 gnd.n7121 19.3944
R9511 gnd.n7175 gnd.n7174 19.3944
R9512 gnd.n7174 gnd.n7173 19.3944
R9513 gnd.n7173 gnd.n7129 19.3944
R9514 gnd.n7169 gnd.n7129 19.3944
R9515 gnd.n7169 gnd.n7168 19.3944
R9516 gnd.n7168 gnd.n7167 19.3944
R9517 gnd.n7167 gnd.n7137 19.3944
R9518 gnd.n7163 gnd.n7137 19.3944
R9519 gnd.n7163 gnd.n7162 19.3944
R9520 gnd.n7162 gnd.n7161 19.3944
R9521 gnd.n7161 gnd.n7145 19.3944
R9522 gnd.n7157 gnd.n7145 19.3944
R9523 gnd.n3005 gnd.n3002 19.3944
R9524 gnd.n3008 gnd.n3005 19.3944
R9525 gnd.n3008 gnd.n2996 19.3944
R9526 gnd.n3020 gnd.n2996 19.3944
R9527 gnd.n3021 gnd.n3020 19.3944
R9528 gnd.n3024 gnd.n3021 19.3944
R9529 gnd.n3024 gnd.n2987 19.3944
R9530 gnd.n3037 gnd.n2987 19.3944
R9531 gnd.n3038 gnd.n3037 19.3944
R9532 gnd.n3041 gnd.n3038 19.3944
R9533 gnd.n3041 gnd.n2978 19.3944
R9534 gnd.n3054 gnd.n2978 19.3944
R9535 gnd.n3055 gnd.n3054 19.3944
R9536 gnd.n3058 gnd.n3055 19.3944
R9537 gnd.n3058 gnd.n2969 19.3944
R9538 gnd.n3071 gnd.n2969 19.3944
R9539 gnd.n5620 gnd.n2777 19.3944
R9540 gnd.n5616 gnd.n2777 19.3944
R9541 gnd.n5616 gnd.n5615 19.3944
R9542 gnd.n5615 gnd.n5614 19.3944
R9543 gnd.n5614 gnd.n2783 19.3944
R9544 gnd.n5610 gnd.n2783 19.3944
R9545 gnd.n5610 gnd.n5609 19.3944
R9546 gnd.n5609 gnd.n5608 19.3944
R9547 gnd.n5608 gnd.n2788 19.3944
R9548 gnd.n5604 gnd.n2788 19.3944
R9549 gnd.n5604 gnd.n5603 19.3944
R9550 gnd.n5603 gnd.n5602 19.3944
R9551 gnd.n5602 gnd.n2793 19.3944
R9552 gnd.n5598 gnd.n2793 19.3944
R9553 gnd.n5598 gnd.n5597 19.3944
R9554 gnd.n5597 gnd.n5596 19.3944
R9555 gnd.n5596 gnd.n2798 19.3944
R9556 gnd.n5592 gnd.n2798 19.3944
R9557 gnd.n5592 gnd.n5591 19.3944
R9558 gnd.n5591 gnd.n5590 19.3944
R9559 gnd.n5590 gnd.n278 19.3944
R9560 gnd.n7036 gnd.n278 19.3944
R9561 gnd.n7036 gnd.n279 19.3944
R9562 gnd.n7032 gnd.n279 19.3944
R9563 gnd.n7032 gnd.n7031 19.3944
R9564 gnd.n7031 gnd.n7030 19.3944
R9565 gnd.n7030 gnd.n285 19.3944
R9566 gnd.n7025 gnd.n285 19.3944
R9567 gnd.n7025 gnd.n7024 19.3944
R9568 gnd.n7024 gnd.n256 19.3944
R9569 gnd.n7047 gnd.n256 19.3944
R9570 gnd.n7047 gnd.n254 19.3944
R9571 gnd.n7051 gnd.n254 19.3944
R9572 gnd.n7051 gnd.n241 19.3944
R9573 gnd.n7063 gnd.n241 19.3944
R9574 gnd.n7063 gnd.n239 19.3944
R9575 gnd.n7067 gnd.n239 19.3944
R9576 gnd.n7067 gnd.n226 19.3944
R9577 gnd.n7079 gnd.n226 19.3944
R9578 gnd.n7079 gnd.n224 19.3944
R9579 gnd.n7083 gnd.n224 19.3944
R9580 gnd.n7083 gnd.n211 19.3944
R9581 gnd.n7095 gnd.n211 19.3944
R9582 gnd.n7095 gnd.n209 19.3944
R9583 gnd.n7099 gnd.n209 19.3944
R9584 gnd.n7099 gnd.n196 19.3944
R9585 gnd.n7111 gnd.n196 19.3944
R9586 gnd.n7111 gnd.n193 19.3944
R9587 gnd.n7190 gnd.n193 19.3944
R9588 gnd.n7190 gnd.n194 19.3944
R9589 gnd.n7186 gnd.n194 19.3944
R9590 gnd.n7186 gnd.n7185 19.3944
R9591 gnd.n7185 gnd.n7184 19.3944
R9592 gnd.n3505 gnd.n2575 19.3944
R9593 gnd.n3506 gnd.n3505 19.3944
R9594 gnd.n3518 gnd.n3506 19.3944
R9595 gnd.n3521 gnd.n3518 19.3944
R9596 gnd.n3521 gnd.n3500 19.3944
R9597 gnd.n3530 gnd.n3500 19.3944
R9598 gnd.n3533 gnd.n3530 19.3944
R9599 gnd.n3533 gnd.n3492 19.3944
R9600 gnd.n3542 gnd.n3492 19.3944
R9601 gnd.n3545 gnd.n3542 19.3944
R9602 gnd.n3545 gnd.n3488 19.3944
R9603 gnd.n3554 gnd.n3488 19.3944
R9604 gnd.n3557 gnd.n3554 19.3944
R9605 gnd.n3557 gnd.n3481 19.3944
R9606 gnd.n3568 gnd.n3481 19.3944
R9607 gnd.n3568 gnd.n3468 19.3944
R9608 gnd.n3689 gnd.n3683 19.3944
R9609 gnd.n3783 gnd.n3683 19.3944
R9610 gnd.n3783 gnd.n3782 19.3944
R9611 gnd.n3782 gnd.n3781 19.3944
R9612 gnd.n3781 gnd.n3696 19.3944
R9613 gnd.n3777 gnd.n3696 19.3944
R9614 gnd.n3777 gnd.n3776 19.3944
R9615 gnd.n3776 gnd.n3775 19.3944
R9616 gnd.n3775 gnd.n3702 19.3944
R9617 gnd.n3771 gnd.n3702 19.3944
R9618 gnd.n3771 gnd.n3770 19.3944
R9619 gnd.n3770 gnd.n3769 19.3944
R9620 gnd.n3769 gnd.n3708 19.3944
R9621 gnd.n3765 gnd.n3708 19.3944
R9622 gnd.n3765 gnd.n3764 19.3944
R9623 gnd.n3764 gnd.n3763 19.3944
R9624 gnd.n3763 gnd.n3714 19.3944
R9625 gnd.n3759 gnd.n3714 19.3944
R9626 gnd.n3759 gnd.n3758 19.3944
R9627 gnd.n3758 gnd.n3757 19.3944
R9628 gnd.n3757 gnd.n3720 19.3944
R9629 gnd.n3753 gnd.n3720 19.3944
R9630 gnd.n3753 gnd.n3752 19.3944
R9631 gnd.n3752 gnd.n3751 19.3944
R9632 gnd.n3751 gnd.n3726 19.3944
R9633 gnd.n3747 gnd.n3726 19.3944
R9634 gnd.n3747 gnd.n3746 19.3944
R9635 gnd.n3746 gnd.n3745 19.3944
R9636 gnd.n3745 gnd.n3732 19.3944
R9637 gnd.n3741 gnd.n3732 19.3944
R9638 gnd.n3741 gnd.n3740 19.3944
R9639 gnd.n3740 gnd.n3739 19.3944
R9640 gnd.n3739 gnd.n3437 19.3944
R9641 gnd.n4417 gnd.n3437 19.3944
R9642 gnd.n4417 gnd.n3435 19.3944
R9643 gnd.n4421 gnd.n3435 19.3944
R9644 gnd.n4421 gnd.n3423 19.3944
R9645 gnd.n4433 gnd.n3423 19.3944
R9646 gnd.n4433 gnd.n3421 19.3944
R9647 gnd.n4439 gnd.n3421 19.3944
R9648 gnd.n4439 gnd.n4438 19.3944
R9649 gnd.n4438 gnd.n3391 19.3944
R9650 gnd.n4557 gnd.n3391 19.3944
R9651 gnd.n4557 gnd.n3389 19.3944
R9652 gnd.n4561 gnd.n3389 19.3944
R9653 gnd.n4561 gnd.n3377 19.3944
R9654 gnd.n4573 gnd.n3377 19.3944
R9655 gnd.n4573 gnd.n3375 19.3944
R9656 gnd.n4577 gnd.n3375 19.3944
R9657 gnd.n4577 gnd.n3362 19.3944
R9658 gnd.n4589 gnd.n3362 19.3944
R9659 gnd.n4589 gnd.n3360 19.3944
R9660 gnd.n4593 gnd.n3360 19.3944
R9661 gnd.n4593 gnd.n3348 19.3944
R9662 gnd.n4604 gnd.n3348 19.3944
R9663 gnd.n4604 gnd.n3346 19.3944
R9664 gnd.n4610 gnd.n3346 19.3944
R9665 gnd.n4610 gnd.n4609 19.3944
R9666 gnd.n4609 gnd.n3316 19.3944
R9667 gnd.n4730 gnd.n3316 19.3944
R9668 gnd.n4730 gnd.n3314 19.3944
R9669 gnd.n4734 gnd.n3314 19.3944
R9670 gnd.n4734 gnd.n3302 19.3944
R9671 gnd.n4746 gnd.n3302 19.3944
R9672 gnd.n4746 gnd.n3300 19.3944
R9673 gnd.n4750 gnd.n3300 19.3944
R9674 gnd.n4750 gnd.n3289 19.3944
R9675 gnd.n4762 gnd.n3289 19.3944
R9676 gnd.n4762 gnd.n3287 19.3944
R9677 gnd.n4766 gnd.n3287 19.3944
R9678 gnd.n4766 gnd.n3278 19.3944
R9679 gnd.n4778 gnd.n3278 19.3944
R9680 gnd.n4778 gnd.n3276 19.3944
R9681 gnd.n4784 gnd.n3276 19.3944
R9682 gnd.n4784 gnd.n4783 19.3944
R9683 gnd.n4783 gnd.n3245 19.3944
R9684 gnd.n4901 gnd.n3245 19.3944
R9685 gnd.n4901 gnd.n3243 19.3944
R9686 gnd.n4905 gnd.n3243 19.3944
R9687 gnd.n4905 gnd.n3230 19.3944
R9688 gnd.n4917 gnd.n3230 19.3944
R9689 gnd.n4917 gnd.n3228 19.3944
R9690 gnd.n4921 gnd.n3228 19.3944
R9691 gnd.n4921 gnd.n3215 19.3944
R9692 gnd.n4933 gnd.n3215 19.3944
R9693 gnd.n4933 gnd.n3213 19.3944
R9694 gnd.n4937 gnd.n3213 19.3944
R9695 gnd.n4937 gnd.n3202 19.3944
R9696 gnd.n4949 gnd.n3202 19.3944
R9697 gnd.n4949 gnd.n3200 19.3944
R9698 gnd.n4955 gnd.n3200 19.3944
R9699 gnd.n4955 gnd.n4954 19.3944
R9700 gnd.n4954 gnd.n3170 19.3944
R9701 gnd.n5307 gnd.n3170 19.3944
R9702 gnd.n5307 gnd.n3168 19.3944
R9703 gnd.n5311 gnd.n3168 19.3944
R9704 gnd.n5311 gnd.n3157 19.3944
R9705 gnd.n5323 gnd.n3157 19.3944
R9706 gnd.n5323 gnd.n3155 19.3944
R9707 gnd.n5327 gnd.n3155 19.3944
R9708 gnd.n5327 gnd.n3143 19.3944
R9709 gnd.n5339 gnd.n3143 19.3944
R9710 gnd.n5339 gnd.n3141 19.3944
R9711 gnd.n5343 gnd.n3141 19.3944
R9712 gnd.n5343 gnd.n3130 19.3944
R9713 gnd.n5355 gnd.n3130 19.3944
R9714 gnd.n5355 gnd.n3128 19.3944
R9715 gnd.n5359 gnd.n3128 19.3944
R9716 gnd.n5359 gnd.n3116 19.3944
R9717 gnd.n5371 gnd.n3116 19.3944
R9718 gnd.n5371 gnd.n3114 19.3944
R9719 gnd.n5375 gnd.n3114 19.3944
R9720 gnd.n5375 gnd.n3102 19.3944
R9721 gnd.n5389 gnd.n3102 19.3944
R9722 gnd.n5389 gnd.n3100 19.3944
R9723 gnd.n5396 gnd.n3100 19.3944
R9724 gnd.n5396 gnd.n5395 19.3944
R9725 gnd.n5395 gnd.n2687 19.3944
R9726 gnd.n5704 gnd.n2687 19.3944
R9727 gnd.n5704 gnd.n5703 19.3944
R9728 gnd.n5703 gnd.n5702 19.3944
R9729 gnd.n5702 gnd.n2691 19.3944
R9730 gnd.n2911 gnd.n2691 19.3944
R9731 gnd.n2915 gnd.n2911 19.3944
R9732 gnd.n2915 gnd.n2909 19.3944
R9733 gnd.n5438 gnd.n2909 19.3944
R9734 gnd.n5438 gnd.n2907 19.3944
R9735 gnd.n5444 gnd.n2907 19.3944
R9736 gnd.n5444 gnd.n5443 19.3944
R9737 gnd.n5443 gnd.n2881 19.3944
R9738 gnd.n5469 gnd.n2881 19.3944
R9739 gnd.n5469 gnd.n2879 19.3944
R9740 gnd.n5475 gnd.n2879 19.3944
R9741 gnd.n5475 gnd.n5474 19.3944
R9742 gnd.n5474 gnd.n2853 19.3944
R9743 gnd.n5505 gnd.n2853 19.3944
R9744 gnd.n5505 gnd.n2851 19.3944
R9745 gnd.n5511 gnd.n2851 19.3944
R9746 gnd.n5511 gnd.n5510 19.3944
R9747 gnd.n5510 gnd.n2819 19.3944
R9748 gnd.n5563 gnd.n2819 19.3944
R9749 gnd.n5563 gnd.n2817 19.3944
R9750 gnd.n5576 gnd.n2817 19.3944
R9751 gnd.n5576 gnd.n5575 19.3944
R9752 gnd.n5575 gnd.n5574 19.3944
R9753 gnd.n5574 gnd.n5571 19.3944
R9754 gnd.n5571 gnd.n311 19.3944
R9755 gnd.n6936 gnd.n311 19.3944
R9756 gnd.n6936 gnd.n6935 19.3944
R9757 gnd.n6935 gnd.n6934 19.3944
R9758 gnd.n6934 gnd.n316 19.3944
R9759 gnd.n6927 gnd.n316 19.3944
R9760 gnd.n6927 gnd.n6926 19.3944
R9761 gnd.n6926 gnd.n6925 19.3944
R9762 gnd.n6711 gnd.n444 19.3944
R9763 gnd.n6717 gnd.n444 19.3944
R9764 gnd.n6717 gnd.n442 19.3944
R9765 gnd.n6721 gnd.n442 19.3944
R9766 gnd.n6721 gnd.n438 19.3944
R9767 gnd.n6727 gnd.n438 19.3944
R9768 gnd.n6727 gnd.n436 19.3944
R9769 gnd.n6731 gnd.n436 19.3944
R9770 gnd.n6731 gnd.n432 19.3944
R9771 gnd.n6737 gnd.n432 19.3944
R9772 gnd.n6737 gnd.n430 19.3944
R9773 gnd.n6741 gnd.n430 19.3944
R9774 gnd.n6741 gnd.n426 19.3944
R9775 gnd.n6747 gnd.n426 19.3944
R9776 gnd.n6747 gnd.n424 19.3944
R9777 gnd.n6751 gnd.n424 19.3944
R9778 gnd.n6751 gnd.n420 19.3944
R9779 gnd.n6757 gnd.n420 19.3944
R9780 gnd.n6757 gnd.n418 19.3944
R9781 gnd.n6761 gnd.n418 19.3944
R9782 gnd.n6761 gnd.n414 19.3944
R9783 gnd.n6767 gnd.n414 19.3944
R9784 gnd.n6767 gnd.n412 19.3944
R9785 gnd.n6771 gnd.n412 19.3944
R9786 gnd.n6771 gnd.n408 19.3944
R9787 gnd.n6777 gnd.n408 19.3944
R9788 gnd.n6777 gnd.n406 19.3944
R9789 gnd.n6781 gnd.n406 19.3944
R9790 gnd.n6781 gnd.n402 19.3944
R9791 gnd.n6787 gnd.n402 19.3944
R9792 gnd.n6787 gnd.n400 19.3944
R9793 gnd.n6791 gnd.n400 19.3944
R9794 gnd.n6791 gnd.n396 19.3944
R9795 gnd.n6797 gnd.n396 19.3944
R9796 gnd.n6797 gnd.n394 19.3944
R9797 gnd.n6801 gnd.n394 19.3944
R9798 gnd.n6801 gnd.n390 19.3944
R9799 gnd.n6807 gnd.n390 19.3944
R9800 gnd.n6807 gnd.n388 19.3944
R9801 gnd.n6811 gnd.n388 19.3944
R9802 gnd.n6811 gnd.n384 19.3944
R9803 gnd.n6817 gnd.n384 19.3944
R9804 gnd.n6817 gnd.n382 19.3944
R9805 gnd.n6821 gnd.n382 19.3944
R9806 gnd.n6821 gnd.n378 19.3944
R9807 gnd.n6827 gnd.n378 19.3944
R9808 gnd.n6827 gnd.n376 19.3944
R9809 gnd.n6831 gnd.n376 19.3944
R9810 gnd.n6831 gnd.n372 19.3944
R9811 gnd.n6837 gnd.n372 19.3944
R9812 gnd.n6837 gnd.n370 19.3944
R9813 gnd.n6841 gnd.n370 19.3944
R9814 gnd.n6841 gnd.n366 19.3944
R9815 gnd.n6847 gnd.n366 19.3944
R9816 gnd.n6847 gnd.n364 19.3944
R9817 gnd.n6851 gnd.n364 19.3944
R9818 gnd.n6851 gnd.n360 19.3944
R9819 gnd.n6857 gnd.n360 19.3944
R9820 gnd.n6857 gnd.n358 19.3944
R9821 gnd.n6861 gnd.n358 19.3944
R9822 gnd.n6861 gnd.n354 19.3944
R9823 gnd.n6867 gnd.n354 19.3944
R9824 gnd.n6867 gnd.n352 19.3944
R9825 gnd.n6871 gnd.n352 19.3944
R9826 gnd.n6871 gnd.n348 19.3944
R9827 gnd.n6877 gnd.n348 19.3944
R9828 gnd.n6877 gnd.n346 19.3944
R9829 gnd.n6881 gnd.n346 19.3944
R9830 gnd.n6881 gnd.n342 19.3944
R9831 gnd.n6887 gnd.n342 19.3944
R9832 gnd.n6887 gnd.n340 19.3944
R9833 gnd.n6891 gnd.n340 19.3944
R9834 gnd.n6891 gnd.n336 19.3944
R9835 gnd.n6897 gnd.n336 19.3944
R9836 gnd.n6897 gnd.n334 19.3944
R9837 gnd.n6901 gnd.n334 19.3944
R9838 gnd.n6901 gnd.n330 19.3944
R9839 gnd.n6907 gnd.n330 19.3944
R9840 gnd.n6907 gnd.n328 19.3944
R9841 gnd.n6911 gnd.n328 19.3944
R9842 gnd.n6911 gnd.n324 19.3944
R9843 gnd.n6918 gnd.n324 19.3944
R9844 gnd.n6918 gnd.n322 19.3944
R9845 gnd.n6922 gnd.n322 19.3944
R9846 gnd.n6326 gnd.n677 19.3944
R9847 gnd.n6326 gnd.n675 19.3944
R9848 gnd.n6330 gnd.n675 19.3944
R9849 gnd.n6330 gnd.n671 19.3944
R9850 gnd.n6336 gnd.n671 19.3944
R9851 gnd.n6336 gnd.n669 19.3944
R9852 gnd.n6340 gnd.n669 19.3944
R9853 gnd.n6340 gnd.n665 19.3944
R9854 gnd.n6346 gnd.n665 19.3944
R9855 gnd.n6346 gnd.n663 19.3944
R9856 gnd.n6350 gnd.n663 19.3944
R9857 gnd.n6350 gnd.n659 19.3944
R9858 gnd.n6356 gnd.n659 19.3944
R9859 gnd.n6356 gnd.n657 19.3944
R9860 gnd.n6360 gnd.n657 19.3944
R9861 gnd.n6360 gnd.n653 19.3944
R9862 gnd.n6366 gnd.n653 19.3944
R9863 gnd.n6366 gnd.n651 19.3944
R9864 gnd.n6370 gnd.n651 19.3944
R9865 gnd.n6370 gnd.n647 19.3944
R9866 gnd.n6376 gnd.n647 19.3944
R9867 gnd.n6376 gnd.n645 19.3944
R9868 gnd.n6380 gnd.n645 19.3944
R9869 gnd.n6380 gnd.n641 19.3944
R9870 gnd.n6386 gnd.n641 19.3944
R9871 gnd.n6386 gnd.n639 19.3944
R9872 gnd.n6390 gnd.n639 19.3944
R9873 gnd.n6390 gnd.n635 19.3944
R9874 gnd.n6396 gnd.n635 19.3944
R9875 gnd.n6396 gnd.n633 19.3944
R9876 gnd.n6400 gnd.n633 19.3944
R9877 gnd.n6400 gnd.n629 19.3944
R9878 gnd.n6406 gnd.n629 19.3944
R9879 gnd.n6406 gnd.n627 19.3944
R9880 gnd.n6410 gnd.n627 19.3944
R9881 gnd.n6410 gnd.n623 19.3944
R9882 gnd.n6416 gnd.n623 19.3944
R9883 gnd.n6416 gnd.n621 19.3944
R9884 gnd.n6420 gnd.n621 19.3944
R9885 gnd.n6420 gnd.n617 19.3944
R9886 gnd.n6426 gnd.n617 19.3944
R9887 gnd.n6426 gnd.n615 19.3944
R9888 gnd.n6430 gnd.n615 19.3944
R9889 gnd.n6430 gnd.n611 19.3944
R9890 gnd.n6436 gnd.n611 19.3944
R9891 gnd.n6436 gnd.n609 19.3944
R9892 gnd.n6440 gnd.n609 19.3944
R9893 gnd.n6440 gnd.n605 19.3944
R9894 gnd.n6446 gnd.n605 19.3944
R9895 gnd.n6446 gnd.n603 19.3944
R9896 gnd.n6450 gnd.n603 19.3944
R9897 gnd.n6450 gnd.n599 19.3944
R9898 gnd.n6456 gnd.n599 19.3944
R9899 gnd.n6456 gnd.n597 19.3944
R9900 gnd.n6460 gnd.n597 19.3944
R9901 gnd.n6460 gnd.n593 19.3944
R9902 gnd.n6466 gnd.n593 19.3944
R9903 gnd.n6466 gnd.n591 19.3944
R9904 gnd.n6470 gnd.n591 19.3944
R9905 gnd.n6470 gnd.n587 19.3944
R9906 gnd.n6476 gnd.n587 19.3944
R9907 gnd.n6476 gnd.n585 19.3944
R9908 gnd.n6480 gnd.n585 19.3944
R9909 gnd.n6480 gnd.n581 19.3944
R9910 gnd.n6486 gnd.n581 19.3944
R9911 gnd.n6486 gnd.n579 19.3944
R9912 gnd.n6490 gnd.n579 19.3944
R9913 gnd.n6490 gnd.n575 19.3944
R9914 gnd.n6496 gnd.n575 19.3944
R9915 gnd.n6496 gnd.n573 19.3944
R9916 gnd.n6500 gnd.n573 19.3944
R9917 gnd.n6500 gnd.n569 19.3944
R9918 gnd.n6506 gnd.n569 19.3944
R9919 gnd.n6506 gnd.n567 19.3944
R9920 gnd.n6510 gnd.n567 19.3944
R9921 gnd.n6510 gnd.n563 19.3944
R9922 gnd.n6516 gnd.n563 19.3944
R9923 gnd.n6516 gnd.n561 19.3944
R9924 gnd.n6520 gnd.n561 19.3944
R9925 gnd.n6520 gnd.n557 19.3944
R9926 gnd.n6526 gnd.n557 19.3944
R9927 gnd.n6526 gnd.n555 19.3944
R9928 gnd.n6530 gnd.n555 19.3944
R9929 gnd.n6530 gnd.n551 19.3944
R9930 gnd.n6536 gnd.n551 19.3944
R9931 gnd.n6536 gnd.n549 19.3944
R9932 gnd.n6540 gnd.n549 19.3944
R9933 gnd.n6540 gnd.n545 19.3944
R9934 gnd.n6546 gnd.n545 19.3944
R9935 gnd.n6546 gnd.n543 19.3944
R9936 gnd.n6550 gnd.n543 19.3944
R9937 gnd.n6550 gnd.n539 19.3944
R9938 gnd.n6556 gnd.n539 19.3944
R9939 gnd.n6556 gnd.n537 19.3944
R9940 gnd.n6560 gnd.n537 19.3944
R9941 gnd.n6560 gnd.n533 19.3944
R9942 gnd.n6566 gnd.n533 19.3944
R9943 gnd.n6566 gnd.n531 19.3944
R9944 gnd.n6570 gnd.n531 19.3944
R9945 gnd.n6570 gnd.n527 19.3944
R9946 gnd.n6576 gnd.n527 19.3944
R9947 gnd.n6576 gnd.n525 19.3944
R9948 gnd.n6580 gnd.n525 19.3944
R9949 gnd.n6580 gnd.n521 19.3944
R9950 gnd.n6586 gnd.n521 19.3944
R9951 gnd.n6586 gnd.n519 19.3944
R9952 gnd.n6590 gnd.n519 19.3944
R9953 gnd.n6590 gnd.n515 19.3944
R9954 gnd.n6596 gnd.n515 19.3944
R9955 gnd.n6596 gnd.n513 19.3944
R9956 gnd.n6600 gnd.n513 19.3944
R9957 gnd.n6600 gnd.n509 19.3944
R9958 gnd.n6606 gnd.n509 19.3944
R9959 gnd.n6606 gnd.n507 19.3944
R9960 gnd.n6610 gnd.n507 19.3944
R9961 gnd.n6610 gnd.n503 19.3944
R9962 gnd.n6616 gnd.n503 19.3944
R9963 gnd.n6616 gnd.n501 19.3944
R9964 gnd.n6620 gnd.n501 19.3944
R9965 gnd.n6620 gnd.n497 19.3944
R9966 gnd.n6626 gnd.n497 19.3944
R9967 gnd.n6626 gnd.n495 19.3944
R9968 gnd.n6630 gnd.n495 19.3944
R9969 gnd.n6630 gnd.n491 19.3944
R9970 gnd.n6636 gnd.n491 19.3944
R9971 gnd.n6636 gnd.n489 19.3944
R9972 gnd.n6640 gnd.n489 19.3944
R9973 gnd.n6640 gnd.n485 19.3944
R9974 gnd.n6646 gnd.n485 19.3944
R9975 gnd.n6646 gnd.n483 19.3944
R9976 gnd.n6650 gnd.n483 19.3944
R9977 gnd.n6650 gnd.n479 19.3944
R9978 gnd.n6656 gnd.n479 19.3944
R9979 gnd.n6656 gnd.n477 19.3944
R9980 gnd.n6660 gnd.n477 19.3944
R9981 gnd.n6660 gnd.n473 19.3944
R9982 gnd.n6666 gnd.n473 19.3944
R9983 gnd.n6666 gnd.n471 19.3944
R9984 gnd.n6670 gnd.n471 19.3944
R9985 gnd.n6670 gnd.n467 19.3944
R9986 gnd.n6676 gnd.n467 19.3944
R9987 gnd.n6676 gnd.n465 19.3944
R9988 gnd.n6680 gnd.n465 19.3944
R9989 gnd.n6680 gnd.n461 19.3944
R9990 gnd.n6686 gnd.n461 19.3944
R9991 gnd.n6686 gnd.n459 19.3944
R9992 gnd.n6690 gnd.n459 19.3944
R9993 gnd.n6690 gnd.n455 19.3944
R9994 gnd.n6696 gnd.n455 19.3944
R9995 gnd.n6696 gnd.n453 19.3944
R9996 gnd.n6701 gnd.n453 19.3944
R9997 gnd.n6701 gnd.n449 19.3944
R9998 gnd.n6707 gnd.n449 19.3944
R9999 gnd.n6708 gnd.n6707 19.3944
R10000 gnd.n5695 gnd.n5694 19.3944
R10001 gnd.n5694 gnd.n5693 19.3944
R10002 gnd.n5693 gnd.n5692 19.3944
R10003 gnd.n5692 gnd.n5690 19.3944
R10004 gnd.n5690 gnd.n5687 19.3944
R10005 gnd.n5687 gnd.n5686 19.3944
R10006 gnd.n5686 gnd.n5683 19.3944
R10007 gnd.n5683 gnd.n5682 19.3944
R10008 gnd.n5682 gnd.n5679 19.3944
R10009 gnd.n5679 gnd.n5678 19.3944
R10010 gnd.n5678 gnd.n5675 19.3944
R10011 gnd.n5675 gnd.n5674 19.3944
R10012 gnd.n5674 gnd.n5671 19.3944
R10013 gnd.n5671 gnd.n5670 19.3944
R10014 gnd.n5670 gnd.n5667 19.3944
R10015 gnd.n5665 gnd.n5662 19.3944
R10016 gnd.n5662 gnd.n5661 19.3944
R10017 gnd.n5661 gnd.n5658 19.3944
R10018 gnd.n5658 gnd.n5657 19.3944
R10019 gnd.n5657 gnd.n5654 19.3944
R10020 gnd.n5654 gnd.n5653 19.3944
R10021 gnd.n5653 gnd.n5650 19.3944
R10022 gnd.n5650 gnd.n5649 19.3944
R10023 gnd.n5649 gnd.n5646 19.3944
R10024 gnd.n5646 gnd.n5645 19.3944
R10025 gnd.n5645 gnd.n5642 19.3944
R10026 gnd.n5642 gnd.n5641 19.3944
R10027 gnd.n5641 gnd.n5638 19.3944
R10028 gnd.n5638 gnd.n5637 19.3944
R10029 gnd.n5637 gnd.n5634 19.3944
R10030 gnd.n5634 gnd.n5633 19.3944
R10031 gnd.n5633 gnd.n5630 19.3944
R10032 gnd.n5630 gnd.n5629 19.3944
R10033 gnd.n2924 gnd.n2771 19.3944
R10034 gnd.n2953 gnd.n2924 19.3944
R10035 gnd.n2953 gnd.n2952 19.3944
R10036 gnd.n2952 gnd.n2951 19.3944
R10037 gnd.n2951 gnd.n2949 19.3944
R10038 gnd.n2949 gnd.n2948 19.3944
R10039 gnd.n2948 gnd.n2946 19.3944
R10040 gnd.n2946 gnd.n2945 19.3944
R10041 gnd.n2945 gnd.n2944 19.3944
R10042 gnd.n2944 gnd.n2942 19.3944
R10043 gnd.n2942 gnd.n2941 19.3944
R10044 gnd.n2941 gnd.n2939 19.3944
R10045 gnd.n2939 gnd.n2938 19.3944
R10046 gnd.n2938 gnd.n2833 19.3944
R10047 gnd.n5527 gnd.n2833 19.3944
R10048 gnd.n5527 gnd.n2831 19.3944
R10049 gnd.n5531 gnd.n2831 19.3944
R10050 gnd.n5532 gnd.n5531 19.3944
R10051 gnd.n5534 gnd.n5532 19.3944
R10052 gnd.n5534 gnd.n2829 19.3944
R10053 gnd.n5546 gnd.n2829 19.3944
R10054 gnd.n5546 gnd.n5545 19.3944
R10055 gnd.n5545 gnd.n5544 19.3944
R10056 gnd.n5544 gnd.n5543 19.3944
R10057 gnd.n5543 gnd.n294 19.3944
R10058 gnd.n6954 gnd.n294 19.3944
R10059 gnd.n6955 gnd.n6954 19.3944
R10060 gnd.n7015 gnd.n6955 19.3944
R10061 gnd.n7015 gnd.n7014 19.3944
R10062 gnd.n7014 gnd.n7013 19.3944
R10063 gnd.n7013 gnd.n7009 19.3944
R10064 gnd.n7009 gnd.n7008 19.3944
R10065 gnd.n7008 gnd.n7006 19.3944
R10066 gnd.n7006 gnd.n7005 19.3944
R10067 gnd.n7005 gnd.n7003 19.3944
R10068 gnd.n7003 gnd.n7002 19.3944
R10069 gnd.n7002 gnd.n7000 19.3944
R10070 gnd.n7000 gnd.n6999 19.3944
R10071 gnd.n6999 gnd.n6997 19.3944
R10072 gnd.n6997 gnd.n6996 19.3944
R10073 gnd.n6996 gnd.n6994 19.3944
R10074 gnd.n6994 gnd.n6993 19.3944
R10075 gnd.n6993 gnd.n6991 19.3944
R10076 gnd.n6991 gnd.n6990 19.3944
R10077 gnd.n6990 gnd.n6988 19.3944
R10078 gnd.n6988 gnd.n6987 19.3944
R10079 gnd.n6987 gnd.n6985 19.3944
R10080 gnd.n6985 gnd.n6984 19.3944
R10081 gnd.n6984 gnd.n6982 19.3944
R10082 gnd.n6982 gnd.n6981 19.3944
R10083 gnd.n6981 gnd.n178 19.3944
R10084 gnd.n7203 gnd.n178 19.3944
R10085 gnd.n7204 gnd.n7203 19.3944
R10086 gnd.n7242 gnd.n139 19.3944
R10087 gnd.n7237 gnd.n139 19.3944
R10088 gnd.n7237 gnd.n7236 19.3944
R10089 gnd.n7236 gnd.n7235 19.3944
R10090 gnd.n7235 gnd.n146 19.3944
R10091 gnd.n7230 gnd.n146 19.3944
R10092 gnd.n7230 gnd.n7229 19.3944
R10093 gnd.n7229 gnd.n7228 19.3944
R10094 gnd.n7228 gnd.n153 19.3944
R10095 gnd.n7223 gnd.n153 19.3944
R10096 gnd.n7223 gnd.n7222 19.3944
R10097 gnd.n7222 gnd.n7221 19.3944
R10098 gnd.n7221 gnd.n160 19.3944
R10099 gnd.n7216 gnd.n160 19.3944
R10100 gnd.n7216 gnd.n7215 19.3944
R10101 gnd.n7215 gnd.n7214 19.3944
R10102 gnd.n7214 gnd.n167 19.3944
R10103 gnd.n7209 gnd.n167 19.3944
R10104 gnd.n7275 gnd.n7274 19.3944
R10105 gnd.n7274 gnd.n7273 19.3944
R10106 gnd.n7273 gnd.n111 19.3944
R10107 gnd.n7268 gnd.n111 19.3944
R10108 gnd.n7268 gnd.n7267 19.3944
R10109 gnd.n7267 gnd.n7266 19.3944
R10110 gnd.n7266 gnd.n118 19.3944
R10111 gnd.n7261 gnd.n118 19.3944
R10112 gnd.n7261 gnd.n7260 19.3944
R10113 gnd.n7260 gnd.n7259 19.3944
R10114 gnd.n7259 gnd.n125 19.3944
R10115 gnd.n7254 gnd.n125 19.3944
R10116 gnd.n7254 gnd.n7253 19.3944
R10117 gnd.n7253 gnd.n7252 19.3944
R10118 gnd.n7252 gnd.n132 19.3944
R10119 gnd.n7247 gnd.n132 19.3944
R10120 gnd.n7247 gnd.n7246 19.3944
R10121 gnd.n2921 gnd.n2918 19.3944
R10122 gnd.n2921 gnd.n2899 19.3944
R10123 gnd.n5449 gnd.n2899 19.3944
R10124 gnd.n5449 gnd.n2897 19.3944
R10125 gnd.n5455 gnd.n2897 19.3944
R10126 gnd.n5455 gnd.n5454 19.3944
R10127 gnd.n5454 gnd.n2870 19.3944
R10128 gnd.n5480 gnd.n2870 19.3944
R10129 gnd.n5480 gnd.n2868 19.3944
R10130 gnd.n5486 gnd.n2868 19.3944
R10131 gnd.n5486 gnd.n5485 19.3944
R10132 gnd.n5485 gnd.n2842 19.3944
R10133 gnd.n5517 gnd.n2842 19.3944
R10134 gnd.n5517 gnd.n2840 19.3944
R10135 gnd.n5523 gnd.n2840 19.3944
R10136 gnd.n5523 gnd.n5522 19.3944
R10137 gnd.n5522 gnd.n2808 19.3944
R10138 gnd.n5581 gnd.n2808 19.3944
R10139 gnd.n5581 gnd.n2806 19.3944
R10140 gnd.n5585 gnd.n2806 19.3944
R10141 gnd.n5585 gnd.n269 19.3944
R10142 gnd.n7040 gnd.n269 19.3944
R10143 gnd.n268 gnd.n267 19.3944
R10144 gnd.n301 gnd.n267 19.3944
R10145 gnd.n6950 gnd.n6949 19.3944
R10146 gnd.n7020 gnd.n7019 19.3944
R10147 gnd.n7043 gnd.n261 19.3944
R10148 gnd.n7043 gnd.n249 19.3944
R10149 gnd.n7055 gnd.n249 19.3944
R10150 gnd.n7055 gnd.n247 19.3944
R10151 gnd.n7059 gnd.n247 19.3944
R10152 gnd.n7059 gnd.n232 19.3944
R10153 gnd.n7071 gnd.n232 19.3944
R10154 gnd.n7071 gnd.n230 19.3944
R10155 gnd.n7075 gnd.n230 19.3944
R10156 gnd.n7075 gnd.n219 19.3944
R10157 gnd.n7087 gnd.n219 19.3944
R10158 gnd.n7087 gnd.n217 19.3944
R10159 gnd.n7091 gnd.n217 19.3944
R10160 gnd.n7091 gnd.n202 19.3944
R10161 gnd.n7103 gnd.n202 19.3944
R10162 gnd.n7103 gnd.n200 19.3944
R10163 gnd.n7107 gnd.n200 19.3944
R10164 gnd.n7107 gnd.n186 19.3944
R10165 gnd.n7194 gnd.n186 19.3944
R10166 gnd.n7194 gnd.n184 19.3944
R10167 gnd.n7198 gnd.n184 19.3944
R10168 gnd.n7198 gnd.n106 19.3944
R10169 gnd.n7278 gnd.n106 19.3944
R10170 gnd.n6073 gnd.n6072 19.3944
R10171 gnd.n6072 gnd.n6071 19.3944
R10172 gnd.n6071 gnd.n6070 19.3944
R10173 gnd.n6070 gnd.n6068 19.3944
R10174 gnd.n6068 gnd.n6065 19.3944
R10175 gnd.n6065 gnd.n6064 19.3944
R10176 gnd.n6064 gnd.n6061 19.3944
R10177 gnd.n6061 gnd.n6060 19.3944
R10178 gnd.n6060 gnd.n6057 19.3944
R10179 gnd.n6057 gnd.n6056 19.3944
R10180 gnd.n6056 gnd.n6053 19.3944
R10181 gnd.n6053 gnd.n6052 19.3944
R10182 gnd.n6052 gnd.n6049 19.3944
R10183 gnd.n6049 gnd.n6048 19.3944
R10184 gnd.n6048 gnd.n6045 19.3944
R10185 gnd.n6045 gnd.n6044 19.3944
R10186 gnd.n6044 gnd.n6041 19.3944
R10187 gnd.n6039 gnd.n6036 19.3944
R10188 gnd.n6036 gnd.n6035 19.3944
R10189 gnd.n6035 gnd.n6032 19.3944
R10190 gnd.n6032 gnd.n6031 19.3944
R10191 gnd.n6031 gnd.n6028 19.3944
R10192 gnd.n6028 gnd.n6027 19.3944
R10193 gnd.n6027 gnd.n6024 19.3944
R10194 gnd.n6024 gnd.n6023 19.3944
R10195 gnd.n6023 gnd.n6020 19.3944
R10196 gnd.n6020 gnd.n6019 19.3944
R10197 gnd.n6019 gnd.n6016 19.3944
R10198 gnd.n6016 gnd.n6015 19.3944
R10199 gnd.n6015 gnd.n6012 19.3944
R10200 gnd.n6012 gnd.n6011 19.3944
R10201 gnd.n6011 gnd.n6008 19.3944
R10202 gnd.n6008 gnd.n6007 19.3944
R10203 gnd.n6007 gnd.n6004 19.3944
R10204 gnd.n6004 gnd.n6003 19.3944
R10205 gnd.n5996 gnd.n5995 19.3944
R10206 gnd.n5995 gnd.n2308 19.3944
R10207 gnd.n5991 gnd.n2308 19.3944
R10208 gnd.n5991 gnd.n2310 19.3944
R10209 gnd.n3931 gnd.n2310 19.3944
R10210 gnd.n3935 gnd.n3931 19.3944
R10211 gnd.n3936 gnd.n3935 19.3944
R10212 gnd.n3938 gnd.n3936 19.3944
R10213 gnd.n3938 gnd.n3929 19.3944
R10214 gnd.n3943 gnd.n3929 19.3944
R10215 gnd.n3944 gnd.n3943 19.3944
R10216 gnd.n3946 gnd.n3944 19.3944
R10217 gnd.n3946 gnd.n3927 19.3944
R10218 gnd.n3951 gnd.n3927 19.3944
R10219 gnd.n3952 gnd.n3951 19.3944
R10220 gnd.n3954 gnd.n3952 19.3944
R10221 gnd.n3954 gnd.n3925 19.3944
R10222 gnd.n3959 gnd.n3925 19.3944
R10223 gnd.n3960 gnd.n3959 19.3944
R10224 gnd.n3962 gnd.n3960 19.3944
R10225 gnd.n3962 gnd.n3923 19.3944
R10226 gnd.n3966 gnd.n3923 19.3944
R10227 gnd.n3966 gnd.n3788 19.3944
R10228 gnd.n3978 gnd.n3788 19.3944
R10229 gnd.n3978 gnd.n3786 19.3944
R10230 gnd.n3984 gnd.n3786 19.3944
R10231 gnd.n3984 gnd.n3677 19.3944
R10232 gnd.n3997 gnd.n3677 19.3944
R10233 gnd.n3997 gnd.n3675 19.3944
R10234 gnd.n4001 gnd.n3675 19.3944
R10235 gnd.n4001 gnd.n3671 19.3944
R10236 gnd.n4013 gnd.n3671 19.3944
R10237 gnd.n4013 gnd.n3669 19.3944
R10238 gnd.n4017 gnd.n3669 19.3944
R10239 gnd.n4017 gnd.n3664 19.3944
R10240 gnd.n4029 gnd.n3664 19.3944
R10241 gnd.n4029 gnd.n3662 19.3944
R10242 gnd.n4033 gnd.n3662 19.3944
R10243 gnd.n4033 gnd.n3658 19.3944
R10244 gnd.n4045 gnd.n3658 19.3944
R10245 gnd.n4045 gnd.n3656 19.3944
R10246 gnd.n4049 gnd.n3656 19.3944
R10247 gnd.n4049 gnd.n3651 19.3944
R10248 gnd.n4061 gnd.n3651 19.3944
R10249 gnd.n4061 gnd.n3649 19.3944
R10250 gnd.n4065 gnd.n3649 19.3944
R10251 gnd.n4065 gnd.n3645 19.3944
R10252 gnd.n4077 gnd.n3645 19.3944
R10253 gnd.n4077 gnd.n3643 19.3944
R10254 gnd.n4082 gnd.n3643 19.3944
R10255 gnd.n4082 gnd.n3637 19.3944
R10256 gnd.n4094 gnd.n3637 19.3944
R10257 gnd.n4095 gnd.n4094 19.3944
R10258 gnd.n4137 gnd.n3611 19.3944
R10259 gnd.n4137 gnd.n4134 19.3944
R10260 gnd.n4134 gnd.n4131 19.3944
R10261 gnd.n4131 gnd.n4130 19.3944
R10262 gnd.n4130 gnd.n4127 19.3944
R10263 gnd.n4127 gnd.n4126 19.3944
R10264 gnd.n4126 gnd.n4123 19.3944
R10265 gnd.n4123 gnd.n4122 19.3944
R10266 gnd.n4122 gnd.n4119 19.3944
R10267 gnd.n4119 gnd.n4118 19.3944
R10268 gnd.n4118 gnd.n4115 19.3944
R10269 gnd.n4115 gnd.n4114 19.3944
R10270 gnd.n4114 gnd.n4111 19.3944
R10271 gnd.n4111 gnd.n4110 19.3944
R10272 gnd.n4110 gnd.n4107 19.3944
R10273 gnd.n4107 gnd.n4106 19.3944
R10274 gnd.n4106 gnd.n4103 19.3944
R10275 gnd.n4103 gnd.n4102 19.3944
R10276 gnd.n3594 gnd.n3593 19.3944
R10277 gnd.n4374 gnd.n3593 19.3944
R10278 gnd.n4374 gnd.n4373 19.3944
R10279 gnd.n4373 gnd.n4372 19.3944
R10280 gnd.n4372 gnd.n4369 19.3944
R10281 gnd.n4369 gnd.n4368 19.3944
R10282 gnd.n4368 gnd.n4365 19.3944
R10283 gnd.n4365 gnd.n4364 19.3944
R10284 gnd.n4364 gnd.n4361 19.3944
R10285 gnd.n4361 gnd.n4360 19.3944
R10286 gnd.n4360 gnd.n4357 19.3944
R10287 gnd.n4357 gnd.n4356 19.3944
R10288 gnd.n4356 gnd.n4353 19.3944
R10289 gnd.n4353 gnd.n4352 19.3944
R10290 gnd.n4352 gnd.n4349 19.3944
R10291 gnd.n3873 gnd.n3805 19.3944
R10292 gnd.n3873 gnd.n3806 19.3944
R10293 gnd.n3869 gnd.n3806 19.3944
R10294 gnd.n3869 gnd.n2330 19.3944
R10295 gnd.n5981 gnd.n2330 19.3944
R10296 gnd.n5981 gnd.n5980 19.3944
R10297 gnd.n5980 gnd.n5979 19.3944
R10298 gnd.n5979 gnd.n2334 19.3944
R10299 gnd.n5969 gnd.n2334 19.3944
R10300 gnd.n5969 gnd.n5968 19.3944
R10301 gnd.n5968 gnd.n5967 19.3944
R10302 gnd.n5967 gnd.n2353 19.3944
R10303 gnd.n5957 gnd.n2353 19.3944
R10304 gnd.n5957 gnd.n5956 19.3944
R10305 gnd.n5956 gnd.n5955 19.3944
R10306 gnd.n5955 gnd.n2374 19.3944
R10307 gnd.n5945 gnd.n2374 19.3944
R10308 gnd.n5945 gnd.n5944 19.3944
R10309 gnd.n5944 gnd.n5943 19.3944
R10310 gnd.n5943 gnd.n2393 19.3944
R10311 gnd.n5933 gnd.n2393 19.3944
R10312 gnd.n5933 gnd.n5932 19.3944
R10313 gnd.n5932 gnd.n5931 19.3944
R10314 gnd.n5931 gnd.n2414 19.3944
R10315 gnd.n5921 gnd.n2414 19.3944
R10316 gnd.n5921 gnd.n5920 19.3944
R10317 gnd.n5920 gnd.n5919 19.3944
R10318 gnd.n5919 gnd.n2432 19.3944
R10319 gnd.n5908 gnd.n2432 19.3944
R10320 gnd.n5908 gnd.n5907 19.3944
R10321 gnd.n5907 gnd.n5906 19.3944
R10322 gnd.n5906 gnd.n2451 19.3944
R10323 gnd.n5896 gnd.n2451 19.3944
R10324 gnd.n5896 gnd.n5895 19.3944
R10325 gnd.n5895 gnd.n5894 19.3944
R10326 gnd.n5894 gnd.n2471 19.3944
R10327 gnd.n5884 gnd.n2471 19.3944
R10328 gnd.n5884 gnd.n5883 19.3944
R10329 gnd.n5883 gnd.n5882 19.3944
R10330 gnd.n5882 gnd.n2493 19.3944
R10331 gnd.n5872 gnd.n2493 19.3944
R10332 gnd.n5872 gnd.n5871 19.3944
R10333 gnd.n5871 gnd.n5870 19.3944
R10334 gnd.n5870 gnd.n2514 19.3944
R10335 gnd.n5860 gnd.n2514 19.3944
R10336 gnd.n5860 gnd.n5859 19.3944
R10337 gnd.n5859 gnd.n5858 19.3944
R10338 gnd.n5858 gnd.n2536 19.3944
R10339 gnd.n5848 gnd.n2536 19.3944
R10340 gnd.n5848 gnd.n5847 19.3944
R10341 gnd.n5847 gnd.n5846 19.3944
R10342 gnd.n5846 gnd.n2558 19.3944
R10343 gnd.n5836 gnd.n2558 19.3944
R10344 gnd.n3865 gnd.n3863 19.3944
R10345 gnd.n3863 gnd.n3860 19.3944
R10346 gnd.n3860 gnd.n3859 19.3944
R10347 gnd.n3859 gnd.n3856 19.3944
R10348 gnd.n3856 gnd.n3855 19.3944
R10349 gnd.n3855 gnd.n3852 19.3944
R10350 gnd.n3852 gnd.n3851 19.3944
R10351 gnd.n3851 gnd.n3848 19.3944
R10352 gnd.n3848 gnd.n3847 19.3944
R10353 gnd.n3847 gnd.n3844 19.3944
R10354 gnd.n3844 gnd.n3843 19.3944
R10355 gnd.n3843 gnd.n3840 19.3944
R10356 gnd.n3840 gnd.n3839 19.3944
R10357 gnd.n3839 gnd.n3836 19.3944
R10358 gnd.n3836 gnd.n3835 19.3944
R10359 gnd.n3835 gnd.n3832 19.3944
R10360 gnd.n3826 gnd.n3801 19.3944
R10361 gnd.n3884 gnd.n3801 19.3944
R10362 gnd.n3884 gnd.n3799 19.3944
R10363 gnd.n3889 gnd.n3799 19.3944
R10364 gnd.n3890 gnd.n3889 19.3944
R10365 gnd.n3892 gnd.n3890 19.3944
R10366 gnd.n3892 gnd.n3797 19.3944
R10367 gnd.n3897 gnd.n3797 19.3944
R10368 gnd.n3898 gnd.n3897 19.3944
R10369 gnd.n3900 gnd.n3898 19.3944
R10370 gnd.n3900 gnd.n3795 19.3944
R10371 gnd.n3905 gnd.n3795 19.3944
R10372 gnd.n3906 gnd.n3905 19.3944
R10373 gnd.n3908 gnd.n3906 19.3944
R10374 gnd.n3908 gnd.n3793 19.3944
R10375 gnd.n3913 gnd.n3793 19.3944
R10376 gnd.n3914 gnd.n3913 19.3944
R10377 gnd.n3916 gnd.n3914 19.3944
R10378 gnd.n3916 gnd.n3791 19.3944
R10379 gnd.n3921 gnd.n3791 19.3944
R10380 gnd.n3922 gnd.n3921 19.3944
R10381 gnd.n3970 gnd.n3922 19.3944
R10382 gnd.n3970 gnd.n3789 19.3944
R10383 gnd.n3974 gnd.n3789 19.3944
R10384 gnd.n3974 gnd.n3680 19.3944
R10385 gnd.n3988 gnd.n3680 19.3944
R10386 gnd.n3988 gnd.n3678 19.3944
R10387 gnd.n3993 gnd.n3678 19.3944
R10388 gnd.n3993 gnd.n3674 19.3944
R10389 gnd.n4005 gnd.n3674 19.3944
R10390 gnd.n4005 gnd.n3672 19.3944
R10391 gnd.n4009 gnd.n3672 19.3944
R10392 gnd.n4009 gnd.n3667 19.3944
R10393 gnd.n4021 gnd.n3667 19.3944
R10394 gnd.n4021 gnd.n3665 19.3944
R10395 gnd.n4025 gnd.n3665 19.3944
R10396 gnd.n4025 gnd.n3661 19.3944
R10397 gnd.n4037 gnd.n3661 19.3944
R10398 gnd.n4037 gnd.n3659 19.3944
R10399 gnd.n4041 gnd.n3659 19.3944
R10400 gnd.n4041 gnd.n3654 19.3944
R10401 gnd.n4053 gnd.n3654 19.3944
R10402 gnd.n4053 gnd.n3652 19.3944
R10403 gnd.n4057 gnd.n3652 19.3944
R10404 gnd.n4057 gnd.n3648 19.3944
R10405 gnd.n4069 gnd.n3648 19.3944
R10406 gnd.n4069 gnd.n3646 19.3944
R10407 gnd.n4073 gnd.n3646 19.3944
R10408 gnd.n4073 gnd.n3642 19.3944
R10409 gnd.n4086 gnd.n3642 19.3944
R10410 gnd.n4086 gnd.n3639 19.3944
R10411 gnd.n4090 gnd.n3639 19.3944
R10412 gnd.n4090 gnd.n3640 19.3944
R10413 gnd.n3879 gnd.n3875 19.3944
R10414 gnd.n3879 gnd.n2319 19.3944
R10415 gnd.n5987 gnd.n2319 19.3944
R10416 gnd.n5987 gnd.n5986 19.3944
R10417 gnd.n5986 gnd.n5985 19.3944
R10418 gnd.n5985 gnd.n2323 19.3944
R10419 gnd.n5975 gnd.n2323 19.3944
R10420 gnd.n5975 gnd.n5974 19.3944
R10421 gnd.n5974 gnd.n5973 19.3944
R10422 gnd.n5973 gnd.n2344 19.3944
R10423 gnd.n5963 gnd.n2344 19.3944
R10424 gnd.n5963 gnd.n5962 19.3944
R10425 gnd.n5962 gnd.n5961 19.3944
R10426 gnd.n5961 gnd.n2363 19.3944
R10427 gnd.n5951 gnd.n2363 19.3944
R10428 gnd.n5951 gnd.n5950 19.3944
R10429 gnd.n5950 gnd.n5949 19.3944
R10430 gnd.n5949 gnd.n2384 19.3944
R10431 gnd.n5939 gnd.n2384 19.3944
R10432 gnd.n5939 gnd.n5938 19.3944
R10433 gnd.n5938 gnd.n5937 19.3944
R10434 gnd.n5937 gnd.n2403 19.3944
R10435 gnd.n5927 gnd.n5926 19.3944
R10436 gnd.n5926 gnd.n5925 19.3944
R10437 gnd.n5915 gnd.n2439 19.3944
R10438 gnd.n5913 gnd.n5912 19.3944
R10439 gnd.n5902 gnd.n2458 19.3944
R10440 gnd.n5902 gnd.n5901 19.3944
R10441 gnd.n5901 gnd.n5900 19.3944
R10442 gnd.n5900 gnd.n2461 19.3944
R10443 gnd.n5890 gnd.n2461 19.3944
R10444 gnd.n5890 gnd.n5889 19.3944
R10445 gnd.n5889 gnd.n5888 19.3944
R10446 gnd.n5888 gnd.n2482 19.3944
R10447 gnd.n5878 gnd.n2482 19.3944
R10448 gnd.n5878 gnd.n5877 19.3944
R10449 gnd.n5877 gnd.n5876 19.3944
R10450 gnd.n5876 gnd.n2504 19.3944
R10451 gnd.n5866 gnd.n2504 19.3944
R10452 gnd.n5866 gnd.n5865 19.3944
R10453 gnd.n5865 gnd.n5864 19.3944
R10454 gnd.n5864 gnd.n2525 19.3944
R10455 gnd.n5854 gnd.n2525 19.3944
R10456 gnd.n5854 gnd.n5853 19.3944
R10457 gnd.n5853 gnd.n5852 19.3944
R10458 gnd.n5852 gnd.n2547 19.3944
R10459 gnd.n5842 gnd.n2547 19.3944
R10460 gnd.n5842 gnd.n5841 19.3944
R10461 gnd.n5841 gnd.n5840 19.3944
R10462 gnd.n6320 gnd.n6319 19.3944
R10463 gnd.n6319 gnd.n6318 19.3944
R10464 gnd.n6318 gnd.n684 19.3944
R10465 gnd.n6312 gnd.n684 19.3944
R10466 gnd.n6312 gnd.n6311 19.3944
R10467 gnd.n6311 gnd.n6310 19.3944
R10468 gnd.n6310 gnd.n692 19.3944
R10469 gnd.n6304 gnd.n692 19.3944
R10470 gnd.n6304 gnd.n6303 19.3944
R10471 gnd.n6303 gnd.n6302 19.3944
R10472 gnd.n6302 gnd.n700 19.3944
R10473 gnd.n6296 gnd.n700 19.3944
R10474 gnd.n6296 gnd.n6295 19.3944
R10475 gnd.n6295 gnd.n6294 19.3944
R10476 gnd.n6294 gnd.n708 19.3944
R10477 gnd.n6288 gnd.n708 19.3944
R10478 gnd.n6288 gnd.n6287 19.3944
R10479 gnd.n6287 gnd.n6286 19.3944
R10480 gnd.n6286 gnd.n716 19.3944
R10481 gnd.n6280 gnd.n716 19.3944
R10482 gnd.n6280 gnd.n6279 19.3944
R10483 gnd.n6279 gnd.n6278 19.3944
R10484 gnd.n6278 gnd.n724 19.3944
R10485 gnd.n6272 gnd.n724 19.3944
R10486 gnd.n6272 gnd.n6271 19.3944
R10487 gnd.n6271 gnd.n6270 19.3944
R10488 gnd.n6270 gnd.n732 19.3944
R10489 gnd.n6264 gnd.n732 19.3944
R10490 gnd.n6264 gnd.n6263 19.3944
R10491 gnd.n6263 gnd.n6262 19.3944
R10492 gnd.n6262 gnd.n740 19.3944
R10493 gnd.n6256 gnd.n740 19.3944
R10494 gnd.n6256 gnd.n6255 19.3944
R10495 gnd.n6255 gnd.n6254 19.3944
R10496 gnd.n6254 gnd.n748 19.3944
R10497 gnd.n6248 gnd.n748 19.3944
R10498 gnd.n6248 gnd.n6247 19.3944
R10499 gnd.n6247 gnd.n6246 19.3944
R10500 gnd.n6246 gnd.n756 19.3944
R10501 gnd.n6240 gnd.n756 19.3944
R10502 gnd.n6240 gnd.n6239 19.3944
R10503 gnd.n6239 gnd.n6238 19.3944
R10504 gnd.n6238 gnd.n764 19.3944
R10505 gnd.n6232 gnd.n764 19.3944
R10506 gnd.n6232 gnd.n6231 19.3944
R10507 gnd.n6231 gnd.n6230 19.3944
R10508 gnd.n6230 gnd.n772 19.3944
R10509 gnd.n6224 gnd.n772 19.3944
R10510 gnd.n6224 gnd.n6223 19.3944
R10511 gnd.n6223 gnd.n6222 19.3944
R10512 gnd.n6222 gnd.n780 19.3944
R10513 gnd.n6216 gnd.n780 19.3944
R10514 gnd.n6216 gnd.n6215 19.3944
R10515 gnd.n6215 gnd.n6214 19.3944
R10516 gnd.n6214 gnd.n788 19.3944
R10517 gnd.n6208 gnd.n788 19.3944
R10518 gnd.n6208 gnd.n6207 19.3944
R10519 gnd.n6207 gnd.n6206 19.3944
R10520 gnd.n6206 gnd.n796 19.3944
R10521 gnd.n6200 gnd.n796 19.3944
R10522 gnd.n6200 gnd.n6199 19.3944
R10523 gnd.n6199 gnd.n6198 19.3944
R10524 gnd.n6198 gnd.n804 19.3944
R10525 gnd.n6192 gnd.n804 19.3944
R10526 gnd.n6192 gnd.n6191 19.3944
R10527 gnd.n6191 gnd.n6190 19.3944
R10528 gnd.n6190 gnd.n812 19.3944
R10529 gnd.n6184 gnd.n812 19.3944
R10530 gnd.n6184 gnd.n6183 19.3944
R10531 gnd.n6183 gnd.n6182 19.3944
R10532 gnd.n6182 gnd.n820 19.3944
R10533 gnd.n6176 gnd.n820 19.3944
R10534 gnd.n6176 gnd.n6175 19.3944
R10535 gnd.n6175 gnd.n6174 19.3944
R10536 gnd.n6174 gnd.n828 19.3944
R10537 gnd.n6168 gnd.n828 19.3944
R10538 gnd.n6168 gnd.n6167 19.3944
R10539 gnd.n6167 gnd.n6166 19.3944
R10540 gnd.n6166 gnd.n836 19.3944
R10541 gnd.n6160 gnd.n836 19.3944
R10542 gnd.n6160 gnd.n6159 19.3944
R10543 gnd.n6159 gnd.n6158 19.3944
R10544 gnd.n6158 gnd.n844 19.3944
R10545 gnd.n3686 gnd.n844 19.3944
R10546 gnd.n5831 gnd.n5830 19.3944
R10547 gnd.n5830 gnd.n5829 19.3944
R10548 gnd.n5829 gnd.n2581 19.3944
R10549 gnd.n5825 gnd.n2581 19.3944
R10550 gnd.n5825 gnd.n5824 19.3944
R10551 gnd.n5824 gnd.n5823 19.3944
R10552 gnd.n5823 gnd.n2586 19.3944
R10553 gnd.n5819 gnd.n2586 19.3944
R10554 gnd.n5819 gnd.n5818 19.3944
R10555 gnd.n5818 gnd.n5817 19.3944
R10556 gnd.n5817 gnd.n2591 19.3944
R10557 gnd.n5813 gnd.n2591 19.3944
R10558 gnd.n5813 gnd.n5812 19.3944
R10559 gnd.n5812 gnd.n5811 19.3944
R10560 gnd.n5811 gnd.n2596 19.3944
R10561 gnd.n5807 gnd.n2596 19.3944
R10562 gnd.n5807 gnd.n5806 19.3944
R10563 gnd.n5806 gnd.n5805 19.3944
R10564 gnd.n5805 gnd.n2601 19.3944
R10565 gnd.n5801 gnd.n2601 19.3944
R10566 gnd.n5801 gnd.n5800 19.3944
R10567 gnd.n5800 gnd.n5799 19.3944
R10568 gnd.n5799 gnd.n2606 19.3944
R10569 gnd.n5795 gnd.n2606 19.3944
R10570 gnd.n5795 gnd.n5794 19.3944
R10571 gnd.n5794 gnd.n5793 19.3944
R10572 gnd.n5793 gnd.n2611 19.3944
R10573 gnd.n5789 gnd.n2611 19.3944
R10574 gnd.n5789 gnd.n5788 19.3944
R10575 gnd.n5788 gnd.n5787 19.3944
R10576 gnd.n5787 gnd.n2616 19.3944
R10577 gnd.n5783 gnd.n2616 19.3944
R10578 gnd.n5783 gnd.n5782 19.3944
R10579 gnd.n5782 gnd.n5781 19.3944
R10580 gnd.n5781 gnd.n2621 19.3944
R10581 gnd.n5777 gnd.n2621 19.3944
R10582 gnd.n5777 gnd.n5776 19.3944
R10583 gnd.n5776 gnd.n5775 19.3944
R10584 gnd.n5775 gnd.n2626 19.3944
R10585 gnd.n5771 gnd.n2626 19.3944
R10586 gnd.n5771 gnd.n5770 19.3944
R10587 gnd.n5770 gnd.n5769 19.3944
R10588 gnd.n5769 gnd.n2631 19.3944
R10589 gnd.n5765 gnd.n2631 19.3944
R10590 gnd.n5765 gnd.n5764 19.3944
R10591 gnd.n5764 gnd.n5763 19.3944
R10592 gnd.n5763 gnd.n2636 19.3944
R10593 gnd.n5759 gnd.n2636 19.3944
R10594 gnd.n5759 gnd.n5758 19.3944
R10595 gnd.n5758 gnd.n5757 19.3944
R10596 gnd.n5757 gnd.n2641 19.3944
R10597 gnd.n5753 gnd.n2641 19.3944
R10598 gnd.n5753 gnd.n5752 19.3944
R10599 gnd.n5752 gnd.n5751 19.3944
R10600 gnd.n5751 gnd.n2646 19.3944
R10601 gnd.n5747 gnd.n2646 19.3944
R10602 gnd.n5747 gnd.n5746 19.3944
R10603 gnd.n5746 gnd.n5745 19.3944
R10604 gnd.n5745 gnd.n2651 19.3944
R10605 gnd.n5741 gnd.n2651 19.3944
R10606 gnd.n5741 gnd.n5740 19.3944
R10607 gnd.n5740 gnd.n5739 19.3944
R10608 gnd.n5739 gnd.n2656 19.3944
R10609 gnd.n5735 gnd.n2656 19.3944
R10610 gnd.n5735 gnd.n5734 19.3944
R10611 gnd.n5734 gnd.n5733 19.3944
R10612 gnd.n5733 gnd.n2661 19.3944
R10613 gnd.n5729 gnd.n2661 19.3944
R10614 gnd.n5729 gnd.n5728 19.3944
R10615 gnd.n5728 gnd.n5727 19.3944
R10616 gnd.n5727 gnd.n2666 19.3944
R10617 gnd.n5723 gnd.n2666 19.3944
R10618 gnd.n5723 gnd.n5722 19.3944
R10619 gnd.n5722 gnd.n5721 19.3944
R10620 gnd.n5721 gnd.n2671 19.3944
R10621 gnd.n5717 gnd.n2671 19.3944
R10622 gnd.n5717 gnd.n5716 19.3944
R10623 gnd.n5716 gnd.n5715 19.3944
R10624 gnd.n5715 gnd.n2676 19.3944
R10625 gnd.n5711 gnd.n2676 19.3944
R10626 gnd.n5711 gnd.n5710 19.3944
R10627 gnd.n5710 gnd.n5709 19.3944
R10628 gnd.n5414 gnd.n3094 19.3944
R10629 gnd.n5410 gnd.n3094 19.3944
R10630 gnd.n5410 gnd.n5409 19.3944
R10631 gnd.n3011 gnd.n3000 19.3944
R10632 gnd.n3016 gnd.n3011 19.3944
R10633 gnd.n3016 gnd.n2993 19.3944
R10634 gnd.n3027 gnd.n2993 19.3944
R10635 gnd.n3027 gnd.n2991 19.3944
R10636 gnd.n3033 gnd.n2991 19.3944
R10637 gnd.n3033 gnd.n2984 19.3944
R10638 gnd.n3044 gnd.n2984 19.3944
R10639 gnd.n3044 gnd.n2982 19.3944
R10640 gnd.n3050 gnd.n2982 19.3944
R10641 gnd.n3050 gnd.n2975 19.3944
R10642 gnd.n3061 gnd.n2975 19.3944
R10643 gnd.n3061 gnd.n2973 19.3944
R10644 gnd.n3067 gnd.n2973 19.3944
R10645 gnd.n3067 gnd.n2963 19.3944
R10646 gnd.n3076 gnd.n2963 19.3944
R10647 gnd.n3076 gnd.n2961 19.3944
R10648 gnd.n2961 gnd.n2960 19.3944
R10649 gnd.n5425 gnd.n2960 19.3944
R10650 gnd.n5425 gnd.n5424 19.3944
R10651 gnd.n5424 gnd.n5423 19.3944
R10652 gnd.n5423 gnd.n3086 19.3944
R10653 gnd.n5419 gnd.n3086 19.3944
R10654 gnd.n5419 gnd.n5418 19.3944
R10655 gnd.n4622 gnd.t5 19.1199
R10656 gnd.n4744 gnd.n3304 19.1199
R10657 gnd.n4682 gnd.n3272 19.1199
R10658 gnd.n4915 gnd.n3232 19.1199
R10659 gnd.n4853 gnd.n3195 19.1199
R10660 gnd.n4975 gnd.t4 19.1199
R10661 gnd.n5231 gnd.n5230 19.1199
R10662 gnd.n1982 gnd.t300 18.8012
R10663 gnd.n1967 gnd.t149 18.8012
R10664 gnd.n1826 gnd.n1825 18.4825
R10665 gnd.t89 gnd.n3119 18.4825
R10666 gnd.n5667 gnd.n5666 18.4247
R10667 gnd.n4349 gnd.n4348 18.4247
R10668 gnd.n7157 gnd.n7156 18.2308
R10669 gnd.n3072 gnd.n3071 18.2308
R10670 gnd.n4381 gnd.n3468 18.2308
R10671 gnd.n3832 gnd.n3825 18.2308
R10672 gnd.t301 gnd.n1506 18.1639
R10673 gnd.n3406 gnd.t2 18.1639
R10674 gnd.t286 gnd.n3125 18.1639
R10675 gnd.n6154 gnd.n6153 17.8452
R10676 gnd.n4579 gnd.n3372 17.8452
R10677 gnd.n4483 gnd.n3350 17.8452
R10678 gnd.n4658 gnd.n3280 17.8452
R10679 gnd.n4923 gnd.n3224 17.8452
R10680 gnd.n5329 gnd.n3152 17.8452
R10681 gnd.n5004 gnd.n3132 17.8452
R10682 gnd.n1534 gnd.t314 17.5266
R10683 gnd.t210 gnd.n2327 17.5266
R10684 gnd.n4752 gnd.t13 17.5266
R10685 gnd.n4829 gnd.t0 17.5266
R10686 gnd.n7109 gnd.t240 17.5266
R10687 gnd.t291 gnd.n3380 17.2079
R10688 gnd.n5260 gnd.t18 17.2079
R10689 gnd.n1933 gnd.t309 16.8893
R10690 gnd.t196 gnd.n2368 16.8893
R10691 gnd.n3655 gnd.t174 16.8893
R10692 gnd.n5503 gnd.t251 16.8893
R10693 gnd.n7077 gnd.t207 16.8893
R10694 gnd.n4587 gnd.n3364 16.5706
R10695 gnd.n4524 gnd.n4523 16.5706
R10696 gnd.n4760 gnd.n3291 16.5706
R10697 gnd.n4697 gnd.n4696 16.5706
R10698 gnd.n4931 gnd.n3217 16.5706
R10699 gnd.n4868 gnd.n4867 16.5706
R10700 gnd.n5337 gnd.n3145 16.5706
R10701 gnd.n5274 gnd.n5273 16.5706
R10702 gnd.n1761 gnd.t68 16.2519
R10703 gnd.n1461 gnd.t308 16.2519
R10704 gnd.n3968 gnd.t183 16.2519
R10705 gnd.n3668 gnd.t163 16.2519
R10706 gnd.n3433 gnd.t96 16.2519
R10707 gnd.t79 gnd.n2682 16.2519
R10708 gnd.n2815 gnd.t194 16.2519
R10709 gnd.n7045 gnd.t178 16.2519
R10710 gnd.n4502 gnd.t141 15.9333
R10711 gnd.t135 gnd.n3166 15.9333
R10712 gnd.n1212 gnd.n1210 15.6674
R10713 gnd.n1180 gnd.n1178 15.6674
R10714 gnd.n1148 gnd.n1146 15.6674
R10715 gnd.n1117 gnd.n1115 15.6674
R10716 gnd.n1085 gnd.n1083 15.6674
R10717 gnd.n1053 gnd.n1051 15.6674
R10718 gnd.n1021 gnd.n1019 15.6674
R10719 gnd.n990 gnd.n988 15.6674
R10720 gnd.n1752 gnd.t68 15.6146
R10721 gnd.n2221 gnd.t100 15.6146
R10722 gnd.t92 gnd.n868 15.6146
R10723 gnd.n5929 gnd.t183 15.6146
R10724 gnd.n3785 gnd.t161 15.6146
R10725 gnd.n4003 gnd.t171 15.6146
R10726 gnd.n4431 gnd.t96 15.6146
R10727 gnd.n5398 gnd.t79 15.6146
R10728 gnd.n6939 gnd.t181 15.6146
R10729 gnd.n6930 gnd.t242 15.6146
R10730 gnd.n7011 gnd.t178 15.6146
R10731 gnd.n5039 gnd.n5038 15.0827
R10732 gnd.n4172 gnd.n4167 15.0481
R10733 gnd.n5049 gnd.n5048 15.0481
R10734 gnd.n2120 gnd.t303 14.9773
R10735 gnd.n5953 gnd.t196 14.9773
R10736 gnd.n4035 gnd.t157 14.9773
R10737 gnd.n5525 gnd.t165 14.9773
R10738 gnd.n237 gnd.t207 14.9773
R10739 gnd.n4595 gnd.t16 14.6587
R10740 gnd.n4988 gnd.t128 14.6587
R10741 gnd.t155 gnd.n1258 14.34
R10742 gnd.n2200 gnd.t313 14.34
R10743 gnd.n5977 gnd.t210 14.34
R10744 gnd.n4067 gnd.t159 14.34
R10745 gnd.t233 gnd.n5466 14.34
R10746 gnd.n207 gnd.t240 14.34
R10747 gnd.n4539 gnd.n3372 14.0214
R10748 gnd.t6 gnd.n3350 14.0214
R10749 gnd.n4712 gnd.n4711 14.0214
R10750 gnd.n4776 gnd.n3280 14.0214
R10751 gnd.n4883 gnd.n3224 14.0214
R10752 gnd.n4947 gnd.n3204 14.0214
R10753 gnd.t298 gnd.n3152 14.0214
R10754 gnd.n5353 gnd.n3132 14.0214
R10755 gnd.n5030 gnd.t20 14.0214
R10756 gnd.n1908 gnd.t320 13.7027
R10757 gnd.t322 gnd.n3366 13.7027
R10758 gnd.n5275 gnd.t288 13.7027
R10759 gnd.n1618 gnd.n1617 13.5763
R10760 gnd.n6131 gnd.n881 13.5763
R10761 gnd.n5629 gnd.n2768 13.5763
R10762 gnd.n7209 gnd.n7208 13.5763
R10763 gnd.n6003 gnd.n2305 13.5763
R10764 gnd.n4102 gnd.n4099 13.5763
R10765 gnd.n1826 gnd.n1564 13.384
R10766 gnd.n4183 gnd.n4164 13.1884
R10767 gnd.n4178 gnd.n4177 13.1884
R10768 gnd.n4177 gnd.n4176 13.1884
R10769 gnd.n5042 gnd.n5037 13.1884
R10770 gnd.n5043 gnd.n5042 13.1884
R10771 gnd.n4179 gnd.n4166 13.146
R10772 gnd.n4175 gnd.n4166 13.146
R10773 gnd.n5041 gnd.n5040 13.146
R10774 gnd.n5041 gnd.n5036 13.146
R10775 gnd.n1213 gnd.n1209 12.8005
R10776 gnd.n1181 gnd.n1177 12.8005
R10777 gnd.n1149 gnd.n1145 12.8005
R10778 gnd.n1118 gnd.n1114 12.8005
R10779 gnd.n1086 gnd.n1082 12.8005
R10780 gnd.n1054 gnd.n1050 12.8005
R10781 gnd.n1022 gnd.n1018 12.8005
R10782 gnd.n991 gnd.n987 12.8005
R10783 gnd.n4441 gnd.n3417 12.7467
R10784 gnd.t55 gnd.t58 12.7467
R10785 gnd.n3406 gnd.n3405 12.7467
R10786 gnd.t12 gnd.n3364 12.7467
R10787 gnd.n4612 gnd.n3342 12.7467
R10788 gnd.n3329 gnd.n3304 12.7467
R10789 gnd.n4786 gnd.n3272 12.7467
R10790 gnd.t290 gnd.n3273 12.7467
R10791 gnd.n4891 gnd.t11 12.7467
R10792 gnd.n3258 gnd.n3232 12.7467
R10793 gnd.n4957 gnd.n3195 12.7467
R10794 gnd.n3183 gnd.n3181 12.7467
R10795 gnd.n5273 gnd.t15 12.7467
R10796 gnd.n5361 gnd.n3125 12.7467
R10797 gnd.t110 gnd.n3118 12.7467
R10798 gnd.t8 gnd.n3342 12.4281
R10799 gnd.n3183 gnd.t151 12.4281
R10800 gnd.n1617 gnd.n1612 12.4126
R10801 gnd.n6127 gnd.n881 12.4126
R10802 gnd.n5625 gnd.n2768 12.4126
R10803 gnd.n7208 gnd.n174 12.4126
R10804 gnd.n5999 gnd.n2305 12.4126
R10805 gnd.n4099 gnd.n3633 12.4126
R10806 gnd.n4265 gnd.n4184 12.1761
R10807 gnd.n5076 gnd.n5054 12.1761
R10808 gnd.n1217 gnd.n1216 12.0247
R10809 gnd.n1185 gnd.n1184 12.0247
R10810 gnd.n1153 gnd.n1152 12.0247
R10811 gnd.n1122 gnd.n1121 12.0247
R10812 gnd.n1090 gnd.n1089 12.0247
R10813 gnd.n1058 gnd.n1057 12.0247
R10814 gnd.n1026 gnd.n1025 12.0247
R10815 gnd.n995 gnd.n994 12.0247
R10816 gnd.n3638 gnd.t47 11.7908
R10817 gnd.n5436 gnd.t37 11.7908
R10818 gnd.n4450 gnd.n3410 11.4721
R10819 gnd.n4621 gnd.n3334 11.4721
R10820 gnd.n3319 gnd.n3311 11.4721
R10821 gnd.n4796 gnd.n4795 11.4721
R10822 gnd.n3249 gnd.n3239 11.4721
R10823 gnd.n4967 gnd.n4966 11.4721
R10824 gnd.n4974 gnd.n3165 11.4721
R10825 gnd.n5369 gnd.n3118 11.4721
R10826 gnd.n5377 gnd.n3112 11.4721
R10827 gnd.n1220 gnd.n1207 11.249
R10828 gnd.n1188 gnd.n1175 11.249
R10829 gnd.n1156 gnd.n1143 11.249
R10830 gnd.n1125 gnd.n1112 11.249
R10831 gnd.n1093 gnd.n1080 11.249
R10832 gnd.n1061 gnd.n1048 11.249
R10833 gnd.n1029 gnd.n1016 11.249
R10834 gnd.n998 gnd.n985 11.249
R10835 gnd.n1896 gnd.t320 11.1535
R10836 gnd.n3976 gnd.n2418 10.8348
R10837 gnd.n5923 gnd.n2424 10.8348
R10838 gnd.n3986 gnd.n3785 10.8348
R10839 gnd.n5917 gnd.n2434 10.8348
R10840 gnd.n5910 gnd.n2442 10.8348
R10841 gnd.n4003 gnd.n2445 10.8348
R10842 gnd.n5904 gnd.n2453 10.8348
R10843 gnd.n4011 gnd.n2456 10.8348
R10844 gnd.n5898 gnd.n2463 10.8348
R10845 gnd.n4019 gnd.n3668 10.8348
R10846 gnd.n5892 gnd.n2473 10.8348
R10847 gnd.n5886 gnd.n2484 10.8348
R10848 gnd.n4035 gnd.n2487 10.8348
R10849 gnd.n5880 gnd.n2495 10.8348
R10850 gnd.n4043 gnd.n2498 10.8348
R10851 gnd.n5874 gnd.n2506 10.8348
R10852 gnd.n4051 gnd.n3655 10.8348
R10853 gnd.n5868 gnd.n2516 10.8348
R10854 gnd.n5862 gnd.n2527 10.8348
R10855 gnd.n4067 gnd.n2530 10.8348
R10856 gnd.n5856 gnd.n2538 10.8348
R10857 gnd.n4075 gnd.n2541 10.8348
R10858 gnd.n5850 gnd.n2549 10.8348
R10859 gnd.n4084 gnd.n2552 10.8348
R10860 gnd.n5844 gnd.n2560 10.8348
R10861 gnd.n4092 gnd.n3638 10.8348
R10862 gnd.n5838 gnd.n2569 10.8348
R10863 gnd.t104 gnd.n3417 10.8348
R10864 gnd.t17 gnd.n3312 10.8348
R10865 gnd.n4720 gnd.t17 10.8348
R10866 gnd.t10 gnd.n3197 10.8348
R10867 gnd.n4846 gnd.t10 10.8348
R10868 gnd.n5622 gnd.n2774 10.8348
R10869 gnd.n5436 gnd.n2923 10.8348
R10870 gnd.n5435 gnd.n2901 10.8348
R10871 gnd.n5447 gnd.n5446 10.8348
R10872 gnd.n2904 gnd.n2891 10.8348
R10873 gnd.n5457 gnd.n2893 10.8348
R10874 gnd.n5467 gnd.n2883 10.8348
R10875 gnd.n5466 gnd.n2872 10.8348
R10876 gnd.n5478 gnd.n5477 10.8348
R10877 gnd.n5488 gnd.n2865 10.8348
R10878 gnd.n5503 gnd.n2855 10.8348
R10879 gnd.n5502 gnd.n2844 10.8348
R10880 gnd.n5515 gnd.n5513 10.8348
R10881 gnd.n2849 gnd.n2847 10.8348
R10882 gnd.n5525 gnd.n2837 10.8348
R10883 gnd.n5561 gnd.n2821 10.8348
R10884 gnd.n5579 gnd.n5578 10.8348
R10885 gnd.n2815 gnd.n2813 10.8348
R10886 gnd.n5587 gnd.n2804 10.8348
R10887 gnd.n5548 gnd.n272 10.8348
R10888 gnd.n7038 gnd.n275 10.8348
R10889 gnd.n6939 gnd.n6938 10.8348
R10890 gnd.n308 gnd.n302 10.8348
R10891 gnd.n6952 gnd.n299 10.8348
R10892 gnd.n6930 gnd.n6929 10.8348
R10893 gnd.n7017 gnd.n289 10.8348
R10894 gnd.n7022 gnd.n291 10.8348
R10895 gnd.n5226 gnd.n5225 10.6151
R10896 gnd.n5225 gnd.n5222 10.6151
R10897 gnd.n5220 gnd.n5217 10.6151
R10898 gnd.n5217 gnd.n5216 10.6151
R10899 gnd.n5216 gnd.n5213 10.6151
R10900 gnd.n5213 gnd.n5212 10.6151
R10901 gnd.n5212 gnd.n5209 10.6151
R10902 gnd.n5209 gnd.n5208 10.6151
R10903 gnd.n5208 gnd.n5205 10.6151
R10904 gnd.n5205 gnd.n5204 10.6151
R10905 gnd.n5204 gnd.n5201 10.6151
R10906 gnd.n5201 gnd.n5200 10.6151
R10907 gnd.n5200 gnd.n5197 10.6151
R10908 gnd.n5197 gnd.n5196 10.6151
R10909 gnd.n5196 gnd.n5193 10.6151
R10910 gnd.n5193 gnd.n5192 10.6151
R10911 gnd.n5192 gnd.n5189 10.6151
R10912 gnd.n5189 gnd.n5188 10.6151
R10913 gnd.n5188 gnd.n5185 10.6151
R10914 gnd.n5185 gnd.n5184 10.6151
R10915 gnd.n5184 gnd.n5181 10.6151
R10916 gnd.n5181 gnd.n5180 10.6151
R10917 gnd.n5180 gnd.n5177 10.6151
R10918 gnd.n5177 gnd.n5176 10.6151
R10919 gnd.n5176 gnd.n5173 10.6151
R10920 gnd.n5173 gnd.n5172 10.6151
R10921 gnd.n5172 gnd.n5169 10.6151
R10922 gnd.n5169 gnd.n5168 10.6151
R10923 gnd.n5168 gnd.n5165 10.6151
R10924 gnd.n5165 gnd.n5164 10.6151
R10925 gnd.n4277 gnd.n4161 10.6151
R10926 gnd.n4277 gnd.n4276 10.6151
R10927 gnd.n4276 gnd.n4275 10.6151
R10928 gnd.n4275 gnd.n3400 10.6151
R10929 gnd.n4553 gnd.n3400 10.6151
R10930 gnd.n4553 gnd.n4552 10.6151
R10931 gnd.n4552 gnd.n4551 10.6151
R10932 gnd.n4551 gnd.n3401 10.6151
R10933 gnd.n3403 gnd.n3401 10.6151
R10934 gnd.n4464 gnd.n3403 10.6151
R10935 gnd.n4465 gnd.n4464 10.6151
R10936 gnd.n4537 gnd.n4465 10.6151
R10937 gnd.n4537 gnd.n4536 10.6151
R10938 gnd.n4536 gnd.n4535 10.6151
R10939 gnd.n4535 gnd.n4466 10.6151
R10940 gnd.n4477 gnd.n4466 10.6151
R10941 gnd.n4479 gnd.n4477 10.6151
R10942 gnd.n4480 gnd.n4479 10.6151
R10943 gnd.n4521 gnd.n4480 10.6151
R10944 gnd.n4521 gnd.n4520 10.6151
R10945 gnd.n4520 gnd.n4519 10.6151
R10946 gnd.n4519 gnd.n4481 10.6151
R10947 gnd.n4492 gnd.n4481 10.6151
R10948 gnd.n4507 gnd.n4492 10.6151
R10949 gnd.n4507 gnd.n4506 10.6151
R10950 gnd.n4506 gnd.n4505 10.6151
R10951 gnd.n4505 gnd.n4493 10.6151
R10952 gnd.n4494 gnd.n4493 10.6151
R10953 gnd.n4494 gnd.n3324 10.6151
R10954 gnd.n4726 gnd.n3324 10.6151
R10955 gnd.n4726 gnd.n4725 10.6151
R10956 gnd.n4725 gnd.n4724 10.6151
R10957 gnd.n4724 gnd.n3325 10.6151
R10958 gnd.n3327 gnd.n3325 10.6151
R10959 gnd.n4635 gnd.n3327 10.6151
R10960 gnd.n4637 gnd.n4635 10.6151
R10961 gnd.n4638 gnd.n4637 10.6151
R10962 gnd.n4709 gnd.n4638 10.6151
R10963 gnd.n4709 gnd.n4708 10.6151
R10964 gnd.n4708 gnd.n4707 10.6151
R10965 gnd.n4707 gnd.n4639 10.6151
R10966 gnd.n4652 gnd.n4639 10.6151
R10967 gnd.n4653 gnd.n4652 10.6151
R10968 gnd.n4694 gnd.n4653 10.6151
R10969 gnd.n4694 gnd.n4693 10.6151
R10970 gnd.n4693 gnd.n4692 10.6151
R10971 gnd.n4692 gnd.n4654 10.6151
R10972 gnd.n4672 gnd.n4654 10.6151
R10973 gnd.n4680 gnd.n4672 10.6151
R10974 gnd.n4680 gnd.n4679 10.6151
R10975 gnd.n4679 gnd.n4678 10.6151
R10976 gnd.n4678 gnd.n4674 10.6151
R10977 gnd.n4674 gnd.n4673 10.6151
R10978 gnd.n4673 gnd.n3254 10.6151
R10979 gnd.n4897 gnd.n3254 10.6151
R10980 gnd.n4897 gnd.n4896 10.6151
R10981 gnd.n4896 gnd.n4895 10.6151
R10982 gnd.n4895 gnd.n3255 10.6151
R10983 gnd.n3257 gnd.n3255 10.6151
R10984 gnd.n4810 gnd.n3257 10.6151
R10985 gnd.n4811 gnd.n4810 10.6151
R10986 gnd.n4881 gnd.n4811 10.6151
R10987 gnd.n4881 gnd.n4880 10.6151
R10988 gnd.n4880 gnd.n4879 10.6151
R10989 gnd.n4879 gnd.n4812 10.6151
R10990 gnd.n4823 gnd.n4812 10.6151
R10991 gnd.n4825 gnd.n4823 10.6151
R10992 gnd.n4826 gnd.n4825 10.6151
R10993 gnd.n4865 gnd.n4826 10.6151
R10994 gnd.n4865 gnd.n4864 10.6151
R10995 gnd.n4864 gnd.n4863 10.6151
R10996 gnd.n4863 gnd.n4827 10.6151
R10997 gnd.n4843 gnd.n4827 10.6151
R10998 gnd.n4851 gnd.n4843 10.6151
R10999 gnd.n4851 gnd.n4850 10.6151
R11000 gnd.n4850 gnd.n4849 10.6151
R11001 gnd.n4849 gnd.n4845 10.6151
R11002 gnd.n4845 gnd.n4844 10.6151
R11003 gnd.n4844 gnd.n3177 10.6151
R11004 gnd.n5303 gnd.n3177 10.6151
R11005 gnd.n5303 gnd.n5302 10.6151
R11006 gnd.n5302 gnd.n5301 10.6151
R11007 gnd.n5301 gnd.n3178 10.6151
R11008 gnd.n3180 gnd.n3178 10.6151
R11009 gnd.n4984 gnd.n3180 10.6151
R11010 gnd.n4985 gnd.n4984 10.6151
R11011 gnd.n5287 gnd.n4985 10.6151
R11012 gnd.n5287 gnd.n5286 10.6151
R11013 gnd.n5286 gnd.n5285 10.6151
R11014 gnd.n5285 gnd.n4986 10.6151
R11015 gnd.n4998 gnd.n4986 10.6151
R11016 gnd.n5000 gnd.n4998 10.6151
R11017 gnd.n5001 gnd.n5000 10.6151
R11018 gnd.n5271 gnd.n5001 10.6151
R11019 gnd.n5271 gnd.n5270 10.6151
R11020 gnd.n5270 gnd.n5269 10.6151
R11021 gnd.n5269 gnd.n5002 10.6151
R11022 gnd.n5013 gnd.n5002 10.6151
R11023 gnd.n5256 gnd.n5013 10.6151
R11024 gnd.n5256 gnd.n5255 10.6151
R11025 gnd.n5255 gnd.n5254 10.6151
R11026 gnd.n5254 gnd.n5014 10.6151
R11027 gnd.n5026 gnd.n5014 10.6151
R11028 gnd.n5027 gnd.n5026 10.6151
R11029 gnd.n5242 gnd.n5027 10.6151
R11030 gnd.n5242 gnd.n5241 10.6151
R11031 gnd.n5241 gnd.n5240 10.6151
R11032 gnd.n5240 gnd.n5028 10.6151
R11033 gnd.n5161 gnd.n5028 10.6151
R11034 gnd.n5162 gnd.n5161 10.6151
R11035 gnd.n4341 gnd.n4141 10.6151
R11036 gnd.n4341 gnd.n4340 10.6151
R11037 gnd.n4338 gnd.n4147 10.6151
R11038 gnd.n4332 gnd.n4147 10.6151
R11039 gnd.n4332 gnd.n4331 10.6151
R11040 gnd.n4331 gnd.n4330 10.6151
R11041 gnd.n4330 gnd.n4149 10.6151
R11042 gnd.n4324 gnd.n4149 10.6151
R11043 gnd.n4324 gnd.n4323 10.6151
R11044 gnd.n4323 gnd.n4322 10.6151
R11045 gnd.n4322 gnd.n4151 10.6151
R11046 gnd.n4316 gnd.n4151 10.6151
R11047 gnd.n4316 gnd.n4315 10.6151
R11048 gnd.n4315 gnd.n4314 10.6151
R11049 gnd.n4314 gnd.n4153 10.6151
R11050 gnd.n4308 gnd.n4153 10.6151
R11051 gnd.n4308 gnd.n4307 10.6151
R11052 gnd.n4307 gnd.n4306 10.6151
R11053 gnd.n4306 gnd.n4155 10.6151
R11054 gnd.n4300 gnd.n4155 10.6151
R11055 gnd.n4300 gnd.n4299 10.6151
R11056 gnd.n4299 gnd.n4298 10.6151
R11057 gnd.n4298 gnd.n4157 10.6151
R11058 gnd.n4292 gnd.n4157 10.6151
R11059 gnd.n4292 gnd.n4291 10.6151
R11060 gnd.n4291 gnd.n4290 10.6151
R11061 gnd.n4290 gnd.n4159 10.6151
R11062 gnd.n4284 gnd.n4159 10.6151
R11063 gnd.n4284 gnd.n4283 10.6151
R11064 gnd.n4283 gnd.n4282 10.6151
R11065 gnd.n4265 gnd.n4264 10.6151
R11066 gnd.n4264 gnd.n4186 10.6151
R11067 gnd.n4260 gnd.n4186 10.6151
R11068 gnd.n4260 gnd.n4259 10.6151
R11069 gnd.n4259 gnd.n4188 10.6151
R11070 gnd.n4254 gnd.n4188 10.6151
R11071 gnd.n4254 gnd.n4253 10.6151
R11072 gnd.n4253 gnd.n4252 10.6151
R11073 gnd.n4252 gnd.n4190 10.6151
R11074 gnd.n4246 gnd.n4190 10.6151
R11075 gnd.n4246 gnd.n4245 10.6151
R11076 gnd.n4245 gnd.n4244 10.6151
R11077 gnd.n4244 gnd.n4192 10.6151
R11078 gnd.n4238 gnd.n4192 10.6151
R11079 gnd.n4238 gnd.n4237 10.6151
R11080 gnd.n4237 gnd.n4236 10.6151
R11081 gnd.n4236 gnd.n4194 10.6151
R11082 gnd.n4230 gnd.n4194 10.6151
R11083 gnd.n4230 gnd.n4229 10.6151
R11084 gnd.n4229 gnd.n4228 10.6151
R11085 gnd.n4228 gnd.n4196 10.6151
R11086 gnd.n4222 gnd.n4196 10.6151
R11087 gnd.n4222 gnd.n4221 10.6151
R11088 gnd.n4221 gnd.n4220 10.6151
R11089 gnd.n4220 gnd.n4198 10.6151
R11090 gnd.n4214 gnd.n4198 10.6151
R11091 gnd.n4214 gnd.n4213 10.6151
R11092 gnd.n4213 gnd.n4212 10.6151
R11093 gnd.n4208 gnd.n4207 10.6151
R11094 gnd.n4207 gnd.n4142 10.6151
R11095 gnd.n5077 gnd.n5076 10.6151
R11096 gnd.n5080 gnd.n5077 10.6151
R11097 gnd.n5081 gnd.n5080 10.6151
R11098 gnd.n5084 gnd.n5081 10.6151
R11099 gnd.n5085 gnd.n5084 10.6151
R11100 gnd.n5088 gnd.n5085 10.6151
R11101 gnd.n5089 gnd.n5088 10.6151
R11102 gnd.n5092 gnd.n5089 10.6151
R11103 gnd.n5093 gnd.n5092 10.6151
R11104 gnd.n5096 gnd.n5093 10.6151
R11105 gnd.n5097 gnd.n5096 10.6151
R11106 gnd.n5100 gnd.n5097 10.6151
R11107 gnd.n5101 gnd.n5100 10.6151
R11108 gnd.n5104 gnd.n5101 10.6151
R11109 gnd.n5105 gnd.n5104 10.6151
R11110 gnd.n5108 gnd.n5105 10.6151
R11111 gnd.n5109 gnd.n5108 10.6151
R11112 gnd.n5112 gnd.n5109 10.6151
R11113 gnd.n5113 gnd.n5112 10.6151
R11114 gnd.n5116 gnd.n5113 10.6151
R11115 gnd.n5117 gnd.n5116 10.6151
R11116 gnd.n5120 gnd.n5117 10.6151
R11117 gnd.n5121 gnd.n5120 10.6151
R11118 gnd.n5124 gnd.n5121 10.6151
R11119 gnd.n5125 gnd.n5124 10.6151
R11120 gnd.n5128 gnd.n5125 10.6151
R11121 gnd.n5129 gnd.n5128 10.6151
R11122 gnd.n5132 gnd.n5129 10.6151
R11123 gnd.n5137 gnd.n5134 10.6151
R11124 gnd.n5138 gnd.n5137 10.6151
R11125 gnd.n4269 gnd.n4268 10.6151
R11126 gnd.n4270 gnd.n4269 10.6151
R11127 gnd.n4270 gnd.n3408 10.6151
R11128 gnd.n4453 gnd.n3408 10.6151
R11129 gnd.n4454 gnd.n4453 10.6151
R11130 gnd.n4455 gnd.n4454 10.6151
R11131 gnd.n4458 gnd.n4455 10.6151
R11132 gnd.n4459 gnd.n4458 10.6151
R11133 gnd.n4545 gnd.n4459 10.6151
R11134 gnd.n4545 gnd.n4544 10.6151
R11135 gnd.n4544 gnd.n4543 10.6151
R11136 gnd.n4543 gnd.n4460 10.6151
R11137 gnd.n4471 gnd.n4460 10.6151
R11138 gnd.n4472 gnd.n4471 10.6151
R11139 gnd.n4530 gnd.n4472 10.6151
R11140 gnd.n4530 gnd.n4529 10.6151
R11141 gnd.n4529 gnd.n4528 10.6151
R11142 gnd.n4528 gnd.n4473 10.6151
R11143 gnd.n4486 gnd.n4473 10.6151
R11144 gnd.n4487 gnd.n4486 10.6151
R11145 gnd.n4515 gnd.n4487 10.6151
R11146 gnd.n4515 gnd.n4514 10.6151
R11147 gnd.n4514 gnd.n4513 10.6151
R11148 gnd.n4513 gnd.n4488 10.6151
R11149 gnd.n4498 gnd.n4488 10.6151
R11150 gnd.n4499 gnd.n4498 10.6151
R11151 gnd.n4500 gnd.n4499 10.6151
R11152 gnd.n4500 gnd.n3332 10.6151
R11153 gnd.n4624 gnd.n3332 10.6151
R11154 gnd.n4625 gnd.n4624 10.6151
R11155 gnd.n4626 gnd.n4625 10.6151
R11156 gnd.n4629 gnd.n4626 10.6151
R11157 gnd.n4630 gnd.n4629 10.6151
R11158 gnd.n4718 gnd.n4630 10.6151
R11159 gnd.n4718 gnd.n4717 10.6151
R11160 gnd.n4717 gnd.n4716 10.6151
R11161 gnd.n4716 gnd.n4631 10.6151
R11162 gnd.n4645 gnd.n4631 10.6151
R11163 gnd.n4646 gnd.n4645 10.6151
R11164 gnd.n4703 gnd.n4646 10.6151
R11165 gnd.n4703 gnd.n4702 10.6151
R11166 gnd.n4702 gnd.n4701 10.6151
R11167 gnd.n4701 gnd.n4647 10.6151
R11168 gnd.n4661 gnd.n4647 10.6151
R11169 gnd.n4662 gnd.n4661 10.6151
R11170 gnd.n4688 gnd.n4662 10.6151
R11171 gnd.n4688 gnd.n4687 10.6151
R11172 gnd.n4687 gnd.n4686 10.6151
R11173 gnd.n4686 gnd.n4663 10.6151
R11174 gnd.n4667 gnd.n4663 10.6151
R11175 gnd.n4667 gnd.n4666 10.6151
R11176 gnd.n4666 gnd.n4665 10.6151
R11177 gnd.n4665 gnd.n3261 10.6151
R11178 gnd.n4799 gnd.n3261 10.6151
R11179 gnd.n4800 gnd.n4799 10.6151
R11180 gnd.n4801 gnd.n4800 10.6151
R11181 gnd.n4804 gnd.n4801 10.6151
R11182 gnd.n4805 gnd.n4804 10.6151
R11183 gnd.n4889 gnd.n4805 10.6151
R11184 gnd.n4889 gnd.n4888 10.6151
R11185 gnd.n4888 gnd.n4887 10.6151
R11186 gnd.n4887 gnd.n4806 10.6151
R11187 gnd.n4817 gnd.n4806 10.6151
R11188 gnd.n4818 gnd.n4817 10.6151
R11189 gnd.n4874 gnd.n4818 10.6151
R11190 gnd.n4874 gnd.n4873 10.6151
R11191 gnd.n4873 gnd.n4872 10.6151
R11192 gnd.n4872 gnd.n4819 10.6151
R11193 gnd.n4832 gnd.n4819 10.6151
R11194 gnd.n4833 gnd.n4832 10.6151
R11195 gnd.n4859 gnd.n4833 10.6151
R11196 gnd.n4859 gnd.n4858 10.6151
R11197 gnd.n4858 gnd.n4857 10.6151
R11198 gnd.n4857 gnd.n4834 10.6151
R11199 gnd.n4838 gnd.n4834 10.6151
R11200 gnd.n4838 gnd.n4837 10.6151
R11201 gnd.n4837 gnd.n4836 10.6151
R11202 gnd.n4836 gnd.n3185 10.6151
R11203 gnd.n4970 gnd.n3185 10.6151
R11204 gnd.n4971 gnd.n4970 10.6151
R11205 gnd.n4972 gnd.n4971 10.6151
R11206 gnd.n4978 gnd.n4972 10.6151
R11207 gnd.n4979 gnd.n4978 10.6151
R11208 gnd.n5295 gnd.n4979 10.6151
R11209 gnd.n5295 gnd.n5294 10.6151
R11210 gnd.n5294 gnd.n5293 10.6151
R11211 gnd.n5293 gnd.n4980 10.6151
R11212 gnd.n4991 gnd.n4980 10.6151
R11213 gnd.n4992 gnd.n4991 10.6151
R11214 gnd.n5280 gnd.n4992 10.6151
R11215 gnd.n5280 gnd.n5279 10.6151
R11216 gnd.n5279 gnd.n5278 10.6151
R11217 gnd.n5278 gnd.n4993 10.6151
R11218 gnd.n5007 gnd.n4993 10.6151
R11219 gnd.n5008 gnd.n5007 10.6151
R11220 gnd.n5265 gnd.n5008 10.6151
R11221 gnd.n5265 gnd.n5264 10.6151
R11222 gnd.n5264 gnd.n5263 10.6151
R11223 gnd.n5263 gnd.n5009 10.6151
R11224 gnd.n5019 gnd.n5009 10.6151
R11225 gnd.n5020 gnd.n5019 10.6151
R11226 gnd.n5249 gnd.n5020 10.6151
R11227 gnd.n5249 gnd.n5248 10.6151
R11228 gnd.n5248 gnd.n5247 10.6151
R11229 gnd.n5247 gnd.n5021 10.6151
R11230 gnd.n5033 gnd.n5021 10.6151
R11231 gnd.n5034 gnd.n5033 10.6151
R11232 gnd.n5235 gnd.n5034 10.6151
R11233 gnd.n5235 gnd.n5234 10.6151
R11234 gnd.n5234 gnd.n5233 10.6151
R11235 gnd.n1815 gnd.t143 10.5161
R11236 gnd.n1260 gnd.t155 10.5161
R11237 gnd.n2179 gnd.t313 10.5161
R11238 gnd.n1221 gnd.n1205 10.4732
R11239 gnd.n1189 gnd.n1173 10.4732
R11240 gnd.n1157 gnd.n1141 10.4732
R11241 gnd.n1126 gnd.n1110 10.4732
R11242 gnd.n1094 gnd.n1078 10.4732
R11243 gnd.n1062 gnd.n1046 10.4732
R11244 gnd.n1030 gnd.n1014 10.4732
R11245 gnd.n999 gnd.n983 10.4732
R11246 gnd.n4451 gnd.n4450 10.1975
R11247 gnd.n3396 gnd.n3395 10.1975
R11248 gnd.n4622 gnd.n4621 10.1975
R11249 gnd.n4795 gnd.n3247 10.1975
R11250 gnd.n3250 gnd.n3249 10.1975
R11251 gnd.n4975 gnd.n4974 10.1975
R11252 gnd.n5369 gnd.n3119 10.1975
R11253 gnd.n5377 gnd.n3111 10.1975
R11254 gnd.t303 gnd.n1277 9.87883
R11255 gnd.n7323 gnd.n62 9.73455
R11256 gnd.n1225 gnd.n1224 9.69747
R11257 gnd.n1193 gnd.n1192 9.69747
R11258 gnd.n1161 gnd.n1160 9.69747
R11259 gnd.n1130 gnd.n1129 9.69747
R11260 gnd.n1098 gnd.n1097 9.69747
R11261 gnd.n1066 gnd.n1065 9.69747
R11262 gnd.n1034 gnd.n1033 9.69747
R11263 gnd.n1003 gnd.n1002 9.69747
R11264 gnd.n4642 gnd.t142 9.56018
R11265 gnd.n4939 gnd.t285 9.56018
R11266 gnd.n5834 gnd.n2575 9.45599
R11267 gnd.n3002 gnd.n2778 9.45599
R11268 gnd.n1231 gnd.n1230 9.45567
R11269 gnd.n1199 gnd.n1198 9.45567
R11270 gnd.n1167 gnd.n1166 9.45567
R11271 gnd.n1136 gnd.n1135 9.45567
R11272 gnd.n1104 gnd.n1103 9.45567
R11273 gnd.n1072 gnd.n1071 9.45567
R11274 gnd.n1040 gnd.n1039 9.45567
R11275 gnd.n1009 gnd.n1008 9.45567
R11276 gnd.n1413 gnd.n1412 9.39724
R11277 gnd.n1230 gnd.n1229 9.3005
R11278 gnd.n1203 gnd.n1202 9.3005
R11279 gnd.n1224 gnd.n1223 9.3005
R11280 gnd.n1222 gnd.n1221 9.3005
R11281 gnd.n1207 gnd.n1206 9.3005
R11282 gnd.n1216 gnd.n1215 9.3005
R11283 gnd.n1214 gnd.n1213 9.3005
R11284 gnd.n1198 gnd.n1197 9.3005
R11285 gnd.n1171 gnd.n1170 9.3005
R11286 gnd.n1192 gnd.n1191 9.3005
R11287 gnd.n1190 gnd.n1189 9.3005
R11288 gnd.n1175 gnd.n1174 9.3005
R11289 gnd.n1184 gnd.n1183 9.3005
R11290 gnd.n1182 gnd.n1181 9.3005
R11291 gnd.n1166 gnd.n1165 9.3005
R11292 gnd.n1139 gnd.n1138 9.3005
R11293 gnd.n1160 gnd.n1159 9.3005
R11294 gnd.n1158 gnd.n1157 9.3005
R11295 gnd.n1143 gnd.n1142 9.3005
R11296 gnd.n1152 gnd.n1151 9.3005
R11297 gnd.n1150 gnd.n1149 9.3005
R11298 gnd.n1135 gnd.n1134 9.3005
R11299 gnd.n1108 gnd.n1107 9.3005
R11300 gnd.n1129 gnd.n1128 9.3005
R11301 gnd.n1127 gnd.n1126 9.3005
R11302 gnd.n1112 gnd.n1111 9.3005
R11303 gnd.n1121 gnd.n1120 9.3005
R11304 gnd.n1119 gnd.n1118 9.3005
R11305 gnd.n1103 gnd.n1102 9.3005
R11306 gnd.n1076 gnd.n1075 9.3005
R11307 gnd.n1097 gnd.n1096 9.3005
R11308 gnd.n1095 gnd.n1094 9.3005
R11309 gnd.n1080 gnd.n1079 9.3005
R11310 gnd.n1089 gnd.n1088 9.3005
R11311 gnd.n1087 gnd.n1086 9.3005
R11312 gnd.n1071 gnd.n1070 9.3005
R11313 gnd.n1044 gnd.n1043 9.3005
R11314 gnd.n1065 gnd.n1064 9.3005
R11315 gnd.n1063 gnd.n1062 9.3005
R11316 gnd.n1048 gnd.n1047 9.3005
R11317 gnd.n1057 gnd.n1056 9.3005
R11318 gnd.n1055 gnd.n1054 9.3005
R11319 gnd.n1039 gnd.n1038 9.3005
R11320 gnd.n1012 gnd.n1011 9.3005
R11321 gnd.n1033 gnd.n1032 9.3005
R11322 gnd.n1031 gnd.n1030 9.3005
R11323 gnd.n1016 gnd.n1015 9.3005
R11324 gnd.n1025 gnd.n1024 9.3005
R11325 gnd.n1023 gnd.n1022 9.3005
R11326 gnd.n1008 gnd.n1007 9.3005
R11327 gnd.n981 gnd.n980 9.3005
R11328 gnd.n1002 gnd.n1001 9.3005
R11329 gnd.n1000 gnd.n999 9.3005
R11330 gnd.n985 gnd.n984 9.3005
R11331 gnd.n994 gnd.n993 9.3005
R11332 gnd.n992 gnd.n991 9.3005
R11333 gnd.n6120 gnd.n6119 9.3005
R11334 gnd.n6118 gnd.n6086 9.3005
R11335 gnd.n6117 gnd.n6116 9.3005
R11336 gnd.n6113 gnd.n6087 9.3005
R11337 gnd.n6110 gnd.n6088 9.3005
R11338 gnd.n6109 gnd.n6089 9.3005
R11339 gnd.n6106 gnd.n6090 9.3005
R11340 gnd.n6105 gnd.n6091 9.3005
R11341 gnd.n6102 gnd.n6092 9.3005
R11342 gnd.n6101 gnd.n6093 9.3005
R11343 gnd.n6098 gnd.n6094 9.3005
R11344 gnd.n6097 gnd.n6095 9.3005
R11345 gnd.n883 gnd.n882 9.3005
R11346 gnd.n6128 gnd.n6127 9.3005
R11347 gnd.n6129 gnd.n881 9.3005
R11348 gnd.n6131 gnd.n6130 9.3005
R11349 gnd.n6121 gnd.n6085 9.3005
R11350 gnd.n1834 gnd.n1833 9.3005
R11351 gnd.n1538 gnd.n1537 9.3005
R11352 gnd.n1861 gnd.n1860 9.3005
R11353 gnd.n1862 gnd.n1536 9.3005
R11354 gnd.n1866 gnd.n1863 9.3005
R11355 gnd.n1865 gnd.n1864 9.3005
R11356 gnd.n1510 gnd.n1509 9.3005
R11357 gnd.n1891 gnd.n1890 9.3005
R11358 gnd.n1892 gnd.n1508 9.3005
R11359 gnd.n1894 gnd.n1893 9.3005
R11360 gnd.n1488 gnd.n1487 9.3005
R11361 gnd.n1922 gnd.n1921 9.3005
R11362 gnd.n1923 gnd.n1486 9.3005
R11363 gnd.n1931 gnd.n1924 9.3005
R11364 gnd.n1930 gnd.n1925 9.3005
R11365 gnd.n1929 gnd.n1927 9.3005
R11366 gnd.n1926 gnd.n1435 9.3005
R11367 gnd.n1979 gnd.n1436 9.3005
R11368 gnd.n1978 gnd.n1437 9.3005
R11369 gnd.n1977 gnd.n1438 9.3005
R11370 gnd.n1457 gnd.n1439 9.3005
R11371 gnd.n1459 gnd.n1458 9.3005
R11372 gnd.n1357 gnd.n1356 9.3005
R11373 gnd.n2017 gnd.n2016 9.3005
R11374 gnd.n2018 gnd.n1355 9.3005
R11375 gnd.n2022 gnd.n2019 9.3005
R11376 gnd.n2021 gnd.n2020 9.3005
R11377 gnd.n1330 gnd.n1329 9.3005
R11378 gnd.n2057 gnd.n2056 9.3005
R11379 gnd.n2058 gnd.n1328 9.3005
R11380 gnd.n2062 gnd.n2059 9.3005
R11381 gnd.n2061 gnd.n2060 9.3005
R11382 gnd.n1303 gnd.n1302 9.3005
R11383 gnd.n2102 gnd.n2101 9.3005
R11384 gnd.n2103 gnd.n1301 9.3005
R11385 gnd.n2107 gnd.n2104 9.3005
R11386 gnd.n2106 gnd.n2105 9.3005
R11387 gnd.n1275 gnd.n1274 9.3005
R11388 gnd.n2142 gnd.n2141 9.3005
R11389 gnd.n2143 gnd.n1273 9.3005
R11390 gnd.n2147 gnd.n2144 9.3005
R11391 gnd.n2146 gnd.n2145 9.3005
R11392 gnd.n1249 gnd.n1248 9.3005
R11393 gnd.n2189 gnd.n2188 9.3005
R11394 gnd.n2190 gnd.n1247 9.3005
R11395 gnd.n2198 gnd.n2191 9.3005
R11396 gnd.n2197 gnd.n2192 9.3005
R11397 gnd.n2196 gnd.n2194 9.3005
R11398 gnd.n2193 gnd.n862 9.3005
R11399 gnd.n6144 gnd.n863 9.3005
R11400 gnd.n6143 gnd.n864 9.3005
R11401 gnd.n6142 gnd.n865 9.3005
R11402 gnd.n6084 gnd.n866 9.3005
R11403 gnd.n1835 gnd.n1832 9.3005
R11404 gnd.n1617 gnd.n1576 9.3005
R11405 gnd.n1612 gnd.n1611 9.3005
R11406 gnd.n1610 gnd.n1577 9.3005
R11407 gnd.n1609 gnd.n1608 9.3005
R11408 gnd.n1605 gnd.n1578 9.3005
R11409 gnd.n1602 gnd.n1601 9.3005
R11410 gnd.n1600 gnd.n1579 9.3005
R11411 gnd.n1599 gnd.n1598 9.3005
R11412 gnd.n1595 gnd.n1580 9.3005
R11413 gnd.n1592 gnd.n1591 9.3005
R11414 gnd.n1590 gnd.n1581 9.3005
R11415 gnd.n1589 gnd.n1588 9.3005
R11416 gnd.n1585 gnd.n1583 9.3005
R11417 gnd.n1582 gnd.n1562 9.3005
R11418 gnd.n1829 gnd.n1561 9.3005
R11419 gnd.n1831 gnd.n1830 9.3005
R11420 gnd.n1619 gnd.n1618 9.3005
R11421 gnd.n1842 gnd.n1548 9.3005
R11422 gnd.n1849 gnd.n1549 9.3005
R11423 gnd.n1851 gnd.n1850 9.3005
R11424 gnd.n1852 gnd.n1529 9.3005
R11425 gnd.n1871 gnd.n1870 9.3005
R11426 gnd.n1873 gnd.n1521 9.3005
R11427 gnd.n1880 gnd.n1523 9.3005
R11428 gnd.n1881 gnd.n1518 9.3005
R11429 gnd.n1883 gnd.n1882 9.3005
R11430 gnd.n1519 gnd.n1504 9.3005
R11431 gnd.n1899 gnd.n1502 9.3005
R11432 gnd.n1903 gnd.n1902 9.3005
R11433 gnd.n1901 gnd.n1478 9.3005
R11434 gnd.n1938 gnd.n1477 9.3005
R11435 gnd.n1941 gnd.n1940 9.3005
R11436 gnd.n1474 gnd.n1473 9.3005
R11437 gnd.n1947 gnd.n1475 9.3005
R11438 gnd.n1949 gnd.n1948 9.3005
R11439 gnd.n1951 gnd.n1472 9.3005
R11440 gnd.n1954 gnd.n1953 9.3005
R11441 gnd.n1957 gnd.n1955 9.3005
R11442 gnd.n1959 gnd.n1958 9.3005
R11443 gnd.n1965 gnd.n1960 9.3005
R11444 gnd.n1964 gnd.n1963 9.3005
R11445 gnd.n1348 gnd.n1347 9.3005
R11446 gnd.n2031 gnd.n2030 9.3005
R11447 gnd.n2032 gnd.n1341 9.3005
R11448 gnd.n2040 gnd.n1340 9.3005
R11449 gnd.n2043 gnd.n2042 9.3005
R11450 gnd.n2045 gnd.n2044 9.3005
R11451 gnd.n2048 gnd.n1323 9.3005
R11452 gnd.n2046 gnd.n1321 9.3005
R11453 gnd.n2068 gnd.n1319 9.3005
R11454 gnd.n2070 gnd.n2069 9.3005
R11455 gnd.n1293 gnd.n1292 9.3005
R11456 gnd.n2116 gnd.n2115 9.3005
R11457 gnd.n2117 gnd.n1286 9.3005
R11458 gnd.n2125 gnd.n1285 9.3005
R11459 gnd.n2128 gnd.n2127 9.3005
R11460 gnd.n2130 gnd.n2129 9.3005
R11461 gnd.n2133 gnd.n1268 9.3005
R11462 gnd.n2131 gnd.n1266 9.3005
R11463 gnd.n2153 gnd.n1264 9.3005
R11464 gnd.n2157 gnd.n2156 9.3005
R11465 gnd.n2155 gnd.n1240 9.3005
R11466 gnd.n2205 gnd.n1239 9.3005
R11467 gnd.n2208 gnd.n2207 9.3005
R11468 gnd.n1236 gnd.n1235 9.3005
R11469 gnd.n2212 gnd.n1237 9.3005
R11470 gnd.n2214 gnd.n2213 9.3005
R11471 gnd.n2218 gnd.n2217 9.3005
R11472 gnd.n877 gnd.n875 9.3005
R11473 gnd.n6135 gnd.n6134 9.3005
R11474 gnd.n1840 gnd.n1839 9.3005
R11475 gnd.n917 gnd.n914 9.3005
R11476 gnd.n919 gnd.n918 9.3005
R11477 gnd.n922 gnd.n912 9.3005
R11478 gnd.n926 gnd.n925 9.3005
R11479 gnd.n927 gnd.n911 9.3005
R11480 gnd.n929 gnd.n928 9.3005
R11481 gnd.n932 gnd.n910 9.3005
R11482 gnd.n936 gnd.n935 9.3005
R11483 gnd.n937 gnd.n909 9.3005
R11484 gnd.n939 gnd.n938 9.3005
R11485 gnd.n942 gnd.n908 9.3005
R11486 gnd.n946 gnd.n945 9.3005
R11487 gnd.n947 gnd.n907 9.3005
R11488 gnd.n949 gnd.n948 9.3005
R11489 gnd.n952 gnd.n906 9.3005
R11490 gnd.n956 gnd.n955 9.3005
R11491 gnd.n957 gnd.n905 9.3005
R11492 gnd.n959 gnd.n958 9.3005
R11493 gnd.n962 gnd.n904 9.3005
R11494 gnd.n966 gnd.n965 9.3005
R11495 gnd.n967 gnd.n903 9.3005
R11496 gnd.n969 gnd.n968 9.3005
R11497 gnd.n972 gnd.n899 9.3005
R11498 gnd.n975 gnd.n974 9.3005
R11499 gnd.n976 gnd.n898 9.3005
R11500 gnd.n2228 gnd.n2227 9.3005
R11501 gnd.n916 gnd.n915 9.3005
R11502 gnd.n2009 gnd.n1993 9.3005
R11503 gnd.n2008 gnd.n1994 9.3005
R11504 gnd.n2007 gnd.n1995 9.3005
R11505 gnd.n2005 gnd.n1996 9.3005
R11506 gnd.n2004 gnd.n1997 9.3005
R11507 gnd.n2002 gnd.n1998 9.3005
R11508 gnd.n2001 gnd.n1999 9.3005
R11509 gnd.n1311 gnd.n1310 9.3005
R11510 gnd.n2078 gnd.n2077 9.3005
R11511 gnd.n2079 gnd.n1309 9.3005
R11512 gnd.n2096 gnd.n2080 9.3005
R11513 gnd.n2095 gnd.n2081 9.3005
R11514 gnd.n2094 gnd.n2082 9.3005
R11515 gnd.n2092 gnd.n2083 9.3005
R11516 gnd.n2091 gnd.n2084 9.3005
R11517 gnd.n2089 gnd.n2085 9.3005
R11518 gnd.n2088 gnd.n2086 9.3005
R11519 gnd.n1255 gnd.n1254 9.3005
R11520 gnd.n2165 gnd.n2164 9.3005
R11521 gnd.n2166 gnd.n1253 9.3005
R11522 gnd.n2183 gnd.n2167 9.3005
R11523 gnd.n2182 gnd.n2168 9.3005
R11524 gnd.n2181 gnd.n2169 9.3005
R11525 gnd.n2178 gnd.n2170 9.3005
R11526 gnd.n2177 gnd.n2171 9.3005
R11527 gnd.n2174 gnd.n2173 9.3005
R11528 gnd.n2172 gnd.n978 9.3005
R11529 gnd.n2224 gnd.n977 9.3005
R11530 gnd.n2226 gnd.n2225 9.3005
R11531 gnd.n1750 gnd.n1749 9.3005
R11532 gnd.n1640 gnd.n1639 9.3005
R11533 gnd.n1764 gnd.n1763 9.3005
R11534 gnd.n1765 gnd.n1638 9.3005
R11535 gnd.n1767 gnd.n1766 9.3005
R11536 gnd.n1628 gnd.n1627 9.3005
R11537 gnd.n1780 gnd.n1779 9.3005
R11538 gnd.n1781 gnd.n1626 9.3005
R11539 gnd.n1813 gnd.n1782 9.3005
R11540 gnd.n1812 gnd.n1783 9.3005
R11541 gnd.n1811 gnd.n1784 9.3005
R11542 gnd.n1810 gnd.n1785 9.3005
R11543 gnd.n1807 gnd.n1786 9.3005
R11544 gnd.n1806 gnd.n1787 9.3005
R11545 gnd.n1805 gnd.n1788 9.3005
R11546 gnd.n1803 gnd.n1789 9.3005
R11547 gnd.n1802 gnd.n1790 9.3005
R11548 gnd.n1799 gnd.n1791 9.3005
R11549 gnd.n1798 gnd.n1792 9.3005
R11550 gnd.n1797 gnd.n1793 9.3005
R11551 gnd.n1795 gnd.n1794 9.3005
R11552 gnd.n1494 gnd.n1493 9.3005
R11553 gnd.n1911 gnd.n1910 9.3005
R11554 gnd.n1912 gnd.n1492 9.3005
R11555 gnd.n1916 gnd.n1913 9.3005
R11556 gnd.n1915 gnd.n1914 9.3005
R11557 gnd.n1416 gnd.n1415 9.3005
R11558 gnd.n1991 gnd.n1990 9.3005
R11559 gnd.n1748 gnd.n1649 9.3005
R11560 gnd.n1651 gnd.n1650 9.3005
R11561 gnd.n1695 gnd.n1693 9.3005
R11562 gnd.n1696 gnd.n1692 9.3005
R11563 gnd.n1699 gnd.n1688 9.3005
R11564 gnd.n1700 gnd.n1687 9.3005
R11565 gnd.n1703 gnd.n1686 9.3005
R11566 gnd.n1704 gnd.n1685 9.3005
R11567 gnd.n1707 gnd.n1684 9.3005
R11568 gnd.n1708 gnd.n1683 9.3005
R11569 gnd.n1711 gnd.n1682 9.3005
R11570 gnd.n1712 gnd.n1681 9.3005
R11571 gnd.n1715 gnd.n1680 9.3005
R11572 gnd.n1716 gnd.n1679 9.3005
R11573 gnd.n1719 gnd.n1678 9.3005
R11574 gnd.n1720 gnd.n1677 9.3005
R11575 gnd.n1723 gnd.n1676 9.3005
R11576 gnd.n1724 gnd.n1675 9.3005
R11577 gnd.n1727 gnd.n1674 9.3005
R11578 gnd.n1728 gnd.n1673 9.3005
R11579 gnd.n1731 gnd.n1672 9.3005
R11580 gnd.n1732 gnd.n1671 9.3005
R11581 gnd.n1735 gnd.n1670 9.3005
R11582 gnd.n1737 gnd.n1669 9.3005
R11583 gnd.n1738 gnd.n1668 9.3005
R11584 gnd.n1739 gnd.n1667 9.3005
R11585 gnd.n1740 gnd.n1666 9.3005
R11586 gnd.n1747 gnd.n1746 9.3005
R11587 gnd.n1756 gnd.n1755 9.3005
R11588 gnd.n1757 gnd.n1643 9.3005
R11589 gnd.n1759 gnd.n1758 9.3005
R11590 gnd.n1634 gnd.n1633 9.3005
R11591 gnd.n1772 gnd.n1771 9.3005
R11592 gnd.n1773 gnd.n1632 9.3005
R11593 gnd.n1775 gnd.n1774 9.3005
R11594 gnd.n1621 gnd.n1620 9.3005
R11595 gnd.n1818 gnd.n1817 9.3005
R11596 gnd.n1819 gnd.n1575 9.3005
R11597 gnd.n1823 gnd.n1821 9.3005
R11598 gnd.n1822 gnd.n1554 9.3005
R11599 gnd.n1841 gnd.n1553 9.3005
R11600 gnd.n1844 gnd.n1843 9.3005
R11601 gnd.n1547 gnd.n1546 9.3005
R11602 gnd.n1855 gnd.n1853 9.3005
R11603 gnd.n1854 gnd.n1528 9.3005
R11604 gnd.n1872 gnd.n1527 9.3005
R11605 gnd.n1875 gnd.n1874 9.3005
R11606 gnd.n1522 gnd.n1517 9.3005
R11607 gnd.n1885 gnd.n1884 9.3005
R11608 gnd.n1520 gnd.n1500 9.3005
R11609 gnd.n1906 gnd.n1501 9.3005
R11610 gnd.n1905 gnd.n1904 9.3005
R11611 gnd.n1503 gnd.n1479 9.3005
R11612 gnd.n1937 gnd.n1936 9.3005
R11613 gnd.n1939 gnd.n1424 9.3005
R11614 gnd.n1986 gnd.n1425 9.3005
R11615 gnd.n1985 gnd.n1426 9.3005
R11616 gnd.n1984 gnd.n1427 9.3005
R11617 gnd.n1950 gnd.n1428 9.3005
R11618 gnd.n1952 gnd.n1446 9.3005
R11619 gnd.n1972 gnd.n1447 9.3005
R11620 gnd.n1971 gnd.n1448 9.3005
R11621 gnd.n1970 gnd.n1449 9.3005
R11622 gnd.n1961 gnd.n1450 9.3005
R11623 gnd.n1962 gnd.n1349 9.3005
R11624 gnd.n2028 gnd.n2027 9.3005
R11625 gnd.n2029 gnd.n1342 9.3005
R11626 gnd.n2039 gnd.n2038 9.3005
R11627 gnd.n2041 gnd.n1338 9.3005
R11628 gnd.n2051 gnd.n1339 9.3005
R11629 gnd.n2050 gnd.n2049 9.3005
R11630 gnd.n2047 gnd.n1317 9.3005
R11631 gnd.n2073 gnd.n1318 9.3005
R11632 gnd.n2072 gnd.n2071 9.3005
R11633 gnd.n1320 gnd.n1294 9.3005
R11634 gnd.n2113 gnd.n2112 9.3005
R11635 gnd.n2114 gnd.n1287 9.3005
R11636 gnd.n2124 gnd.n2123 9.3005
R11637 gnd.n2126 gnd.n1283 9.3005
R11638 gnd.n2136 gnd.n1284 9.3005
R11639 gnd.n2135 gnd.n2134 9.3005
R11640 gnd.n2132 gnd.n1262 9.3005
R11641 gnd.n2160 gnd.n1263 9.3005
R11642 gnd.n2159 gnd.n2158 9.3005
R11643 gnd.n1265 gnd.n1241 9.3005
R11644 gnd.n2204 gnd.n2203 9.3005
R11645 gnd.n2206 gnd.n851 9.3005
R11646 gnd.n6151 gnd.n852 9.3005
R11647 gnd.n6150 gnd.n853 9.3005
R11648 gnd.n6149 gnd.n854 9.3005
R11649 gnd.n2215 gnd.n855 9.3005
R11650 gnd.n2216 gnd.n874 9.3005
R11651 gnd.n6137 gnd.n6136 9.3005
R11652 gnd.n1645 gnd.n1644 9.3005
R11653 gnd.n677 gnd.n676 9.3005
R11654 gnd.n6327 gnd.n6326 9.3005
R11655 gnd.n6328 gnd.n675 9.3005
R11656 gnd.n6330 gnd.n6329 9.3005
R11657 gnd.n671 gnd.n670 9.3005
R11658 gnd.n6337 gnd.n6336 9.3005
R11659 gnd.n6338 gnd.n669 9.3005
R11660 gnd.n6340 gnd.n6339 9.3005
R11661 gnd.n665 gnd.n664 9.3005
R11662 gnd.n6347 gnd.n6346 9.3005
R11663 gnd.n6348 gnd.n663 9.3005
R11664 gnd.n6350 gnd.n6349 9.3005
R11665 gnd.n659 gnd.n658 9.3005
R11666 gnd.n6357 gnd.n6356 9.3005
R11667 gnd.n6358 gnd.n657 9.3005
R11668 gnd.n6360 gnd.n6359 9.3005
R11669 gnd.n653 gnd.n652 9.3005
R11670 gnd.n6367 gnd.n6366 9.3005
R11671 gnd.n6368 gnd.n651 9.3005
R11672 gnd.n6370 gnd.n6369 9.3005
R11673 gnd.n647 gnd.n646 9.3005
R11674 gnd.n6377 gnd.n6376 9.3005
R11675 gnd.n6378 gnd.n645 9.3005
R11676 gnd.n6380 gnd.n6379 9.3005
R11677 gnd.n641 gnd.n640 9.3005
R11678 gnd.n6387 gnd.n6386 9.3005
R11679 gnd.n6388 gnd.n639 9.3005
R11680 gnd.n6390 gnd.n6389 9.3005
R11681 gnd.n635 gnd.n634 9.3005
R11682 gnd.n6397 gnd.n6396 9.3005
R11683 gnd.n6398 gnd.n633 9.3005
R11684 gnd.n6400 gnd.n6399 9.3005
R11685 gnd.n629 gnd.n628 9.3005
R11686 gnd.n6407 gnd.n6406 9.3005
R11687 gnd.n6408 gnd.n627 9.3005
R11688 gnd.n6410 gnd.n6409 9.3005
R11689 gnd.n623 gnd.n622 9.3005
R11690 gnd.n6417 gnd.n6416 9.3005
R11691 gnd.n6418 gnd.n621 9.3005
R11692 gnd.n6420 gnd.n6419 9.3005
R11693 gnd.n617 gnd.n616 9.3005
R11694 gnd.n6427 gnd.n6426 9.3005
R11695 gnd.n6428 gnd.n615 9.3005
R11696 gnd.n6430 gnd.n6429 9.3005
R11697 gnd.n611 gnd.n610 9.3005
R11698 gnd.n6437 gnd.n6436 9.3005
R11699 gnd.n6438 gnd.n609 9.3005
R11700 gnd.n6440 gnd.n6439 9.3005
R11701 gnd.n605 gnd.n604 9.3005
R11702 gnd.n6447 gnd.n6446 9.3005
R11703 gnd.n6448 gnd.n603 9.3005
R11704 gnd.n6450 gnd.n6449 9.3005
R11705 gnd.n599 gnd.n598 9.3005
R11706 gnd.n6457 gnd.n6456 9.3005
R11707 gnd.n6458 gnd.n597 9.3005
R11708 gnd.n6460 gnd.n6459 9.3005
R11709 gnd.n593 gnd.n592 9.3005
R11710 gnd.n6467 gnd.n6466 9.3005
R11711 gnd.n6468 gnd.n591 9.3005
R11712 gnd.n6470 gnd.n6469 9.3005
R11713 gnd.n587 gnd.n586 9.3005
R11714 gnd.n6477 gnd.n6476 9.3005
R11715 gnd.n6478 gnd.n585 9.3005
R11716 gnd.n6480 gnd.n6479 9.3005
R11717 gnd.n581 gnd.n580 9.3005
R11718 gnd.n6487 gnd.n6486 9.3005
R11719 gnd.n6488 gnd.n579 9.3005
R11720 gnd.n6490 gnd.n6489 9.3005
R11721 gnd.n575 gnd.n574 9.3005
R11722 gnd.n6497 gnd.n6496 9.3005
R11723 gnd.n6498 gnd.n573 9.3005
R11724 gnd.n6500 gnd.n6499 9.3005
R11725 gnd.n569 gnd.n568 9.3005
R11726 gnd.n6507 gnd.n6506 9.3005
R11727 gnd.n6508 gnd.n567 9.3005
R11728 gnd.n6510 gnd.n6509 9.3005
R11729 gnd.n563 gnd.n562 9.3005
R11730 gnd.n6517 gnd.n6516 9.3005
R11731 gnd.n6518 gnd.n561 9.3005
R11732 gnd.n6520 gnd.n6519 9.3005
R11733 gnd.n557 gnd.n556 9.3005
R11734 gnd.n6527 gnd.n6526 9.3005
R11735 gnd.n6528 gnd.n555 9.3005
R11736 gnd.n6530 gnd.n6529 9.3005
R11737 gnd.n551 gnd.n550 9.3005
R11738 gnd.n6537 gnd.n6536 9.3005
R11739 gnd.n6538 gnd.n549 9.3005
R11740 gnd.n6540 gnd.n6539 9.3005
R11741 gnd.n545 gnd.n544 9.3005
R11742 gnd.n6547 gnd.n6546 9.3005
R11743 gnd.n6548 gnd.n543 9.3005
R11744 gnd.n6550 gnd.n6549 9.3005
R11745 gnd.n539 gnd.n538 9.3005
R11746 gnd.n6557 gnd.n6556 9.3005
R11747 gnd.n6558 gnd.n537 9.3005
R11748 gnd.n6560 gnd.n6559 9.3005
R11749 gnd.n533 gnd.n532 9.3005
R11750 gnd.n6567 gnd.n6566 9.3005
R11751 gnd.n6568 gnd.n531 9.3005
R11752 gnd.n6570 gnd.n6569 9.3005
R11753 gnd.n527 gnd.n526 9.3005
R11754 gnd.n6577 gnd.n6576 9.3005
R11755 gnd.n6578 gnd.n525 9.3005
R11756 gnd.n6580 gnd.n6579 9.3005
R11757 gnd.n521 gnd.n520 9.3005
R11758 gnd.n6587 gnd.n6586 9.3005
R11759 gnd.n6588 gnd.n519 9.3005
R11760 gnd.n6590 gnd.n6589 9.3005
R11761 gnd.n515 gnd.n514 9.3005
R11762 gnd.n6597 gnd.n6596 9.3005
R11763 gnd.n6598 gnd.n513 9.3005
R11764 gnd.n6600 gnd.n6599 9.3005
R11765 gnd.n509 gnd.n508 9.3005
R11766 gnd.n6607 gnd.n6606 9.3005
R11767 gnd.n6608 gnd.n507 9.3005
R11768 gnd.n6610 gnd.n6609 9.3005
R11769 gnd.n503 gnd.n502 9.3005
R11770 gnd.n6617 gnd.n6616 9.3005
R11771 gnd.n6618 gnd.n501 9.3005
R11772 gnd.n6620 gnd.n6619 9.3005
R11773 gnd.n497 gnd.n496 9.3005
R11774 gnd.n6627 gnd.n6626 9.3005
R11775 gnd.n6628 gnd.n495 9.3005
R11776 gnd.n6630 gnd.n6629 9.3005
R11777 gnd.n491 gnd.n490 9.3005
R11778 gnd.n6637 gnd.n6636 9.3005
R11779 gnd.n6638 gnd.n489 9.3005
R11780 gnd.n6640 gnd.n6639 9.3005
R11781 gnd.n485 gnd.n484 9.3005
R11782 gnd.n6647 gnd.n6646 9.3005
R11783 gnd.n6648 gnd.n483 9.3005
R11784 gnd.n6650 gnd.n6649 9.3005
R11785 gnd.n479 gnd.n478 9.3005
R11786 gnd.n6657 gnd.n6656 9.3005
R11787 gnd.n6658 gnd.n477 9.3005
R11788 gnd.n6660 gnd.n6659 9.3005
R11789 gnd.n473 gnd.n472 9.3005
R11790 gnd.n6667 gnd.n6666 9.3005
R11791 gnd.n6668 gnd.n471 9.3005
R11792 gnd.n6670 gnd.n6669 9.3005
R11793 gnd.n467 gnd.n466 9.3005
R11794 gnd.n6677 gnd.n6676 9.3005
R11795 gnd.n6678 gnd.n465 9.3005
R11796 gnd.n6680 gnd.n6679 9.3005
R11797 gnd.n461 gnd.n460 9.3005
R11798 gnd.n6687 gnd.n6686 9.3005
R11799 gnd.n6688 gnd.n459 9.3005
R11800 gnd.n6690 gnd.n6689 9.3005
R11801 gnd.n455 gnd.n454 9.3005
R11802 gnd.n6697 gnd.n6696 9.3005
R11803 gnd.n6698 gnd.n453 9.3005
R11804 gnd.n6701 gnd.n6700 9.3005
R11805 gnd.n6699 gnd.n449 9.3005
R11806 gnd.n6707 gnd.n448 9.3005
R11807 gnd.n6709 gnd.n6708 9.3005
R11808 gnd.n444 gnd.n443 9.3005
R11809 gnd.n6718 gnd.n6717 9.3005
R11810 gnd.n6719 gnd.n442 9.3005
R11811 gnd.n6721 gnd.n6720 9.3005
R11812 gnd.n438 gnd.n437 9.3005
R11813 gnd.n6728 gnd.n6727 9.3005
R11814 gnd.n6729 gnd.n436 9.3005
R11815 gnd.n6731 gnd.n6730 9.3005
R11816 gnd.n432 gnd.n431 9.3005
R11817 gnd.n6738 gnd.n6737 9.3005
R11818 gnd.n6739 gnd.n430 9.3005
R11819 gnd.n6741 gnd.n6740 9.3005
R11820 gnd.n426 gnd.n425 9.3005
R11821 gnd.n6748 gnd.n6747 9.3005
R11822 gnd.n6749 gnd.n424 9.3005
R11823 gnd.n6751 gnd.n6750 9.3005
R11824 gnd.n420 gnd.n419 9.3005
R11825 gnd.n6758 gnd.n6757 9.3005
R11826 gnd.n6759 gnd.n418 9.3005
R11827 gnd.n6761 gnd.n6760 9.3005
R11828 gnd.n414 gnd.n413 9.3005
R11829 gnd.n6768 gnd.n6767 9.3005
R11830 gnd.n6769 gnd.n412 9.3005
R11831 gnd.n6771 gnd.n6770 9.3005
R11832 gnd.n408 gnd.n407 9.3005
R11833 gnd.n6778 gnd.n6777 9.3005
R11834 gnd.n6779 gnd.n406 9.3005
R11835 gnd.n6781 gnd.n6780 9.3005
R11836 gnd.n402 gnd.n401 9.3005
R11837 gnd.n6788 gnd.n6787 9.3005
R11838 gnd.n6789 gnd.n400 9.3005
R11839 gnd.n6791 gnd.n6790 9.3005
R11840 gnd.n396 gnd.n395 9.3005
R11841 gnd.n6798 gnd.n6797 9.3005
R11842 gnd.n6799 gnd.n394 9.3005
R11843 gnd.n6801 gnd.n6800 9.3005
R11844 gnd.n390 gnd.n389 9.3005
R11845 gnd.n6808 gnd.n6807 9.3005
R11846 gnd.n6809 gnd.n388 9.3005
R11847 gnd.n6811 gnd.n6810 9.3005
R11848 gnd.n384 gnd.n383 9.3005
R11849 gnd.n6818 gnd.n6817 9.3005
R11850 gnd.n6819 gnd.n382 9.3005
R11851 gnd.n6821 gnd.n6820 9.3005
R11852 gnd.n378 gnd.n377 9.3005
R11853 gnd.n6828 gnd.n6827 9.3005
R11854 gnd.n6829 gnd.n376 9.3005
R11855 gnd.n6831 gnd.n6830 9.3005
R11856 gnd.n372 gnd.n371 9.3005
R11857 gnd.n6838 gnd.n6837 9.3005
R11858 gnd.n6839 gnd.n370 9.3005
R11859 gnd.n6841 gnd.n6840 9.3005
R11860 gnd.n366 gnd.n365 9.3005
R11861 gnd.n6848 gnd.n6847 9.3005
R11862 gnd.n6849 gnd.n364 9.3005
R11863 gnd.n6851 gnd.n6850 9.3005
R11864 gnd.n360 gnd.n359 9.3005
R11865 gnd.n6858 gnd.n6857 9.3005
R11866 gnd.n6859 gnd.n358 9.3005
R11867 gnd.n6861 gnd.n6860 9.3005
R11868 gnd.n354 gnd.n353 9.3005
R11869 gnd.n6868 gnd.n6867 9.3005
R11870 gnd.n6869 gnd.n352 9.3005
R11871 gnd.n6871 gnd.n6870 9.3005
R11872 gnd.n348 gnd.n347 9.3005
R11873 gnd.n6878 gnd.n6877 9.3005
R11874 gnd.n6879 gnd.n346 9.3005
R11875 gnd.n6881 gnd.n6880 9.3005
R11876 gnd.n342 gnd.n341 9.3005
R11877 gnd.n6888 gnd.n6887 9.3005
R11878 gnd.n6889 gnd.n340 9.3005
R11879 gnd.n6891 gnd.n6890 9.3005
R11880 gnd.n336 gnd.n335 9.3005
R11881 gnd.n6898 gnd.n6897 9.3005
R11882 gnd.n6899 gnd.n334 9.3005
R11883 gnd.n6901 gnd.n6900 9.3005
R11884 gnd.n330 gnd.n329 9.3005
R11885 gnd.n6908 gnd.n6907 9.3005
R11886 gnd.n6909 gnd.n328 9.3005
R11887 gnd.n6911 gnd.n6910 9.3005
R11888 gnd.n324 gnd.n323 9.3005
R11889 gnd.n6919 gnd.n6918 9.3005
R11890 gnd.n6920 gnd.n322 9.3005
R11891 gnd.n6922 gnd.n6921 9.3005
R11892 gnd.n6711 gnd.n6710 9.3005
R11893 gnd.n7274 gnd.n108 9.3005
R11894 gnd.n7273 gnd.n110 9.3005
R11895 gnd.n114 gnd.n111 9.3005
R11896 gnd.n7268 gnd.n115 9.3005
R11897 gnd.n7267 gnd.n116 9.3005
R11898 gnd.n7266 gnd.n117 9.3005
R11899 gnd.n121 gnd.n118 9.3005
R11900 gnd.n7261 gnd.n122 9.3005
R11901 gnd.n7260 gnd.n123 9.3005
R11902 gnd.n7259 gnd.n124 9.3005
R11903 gnd.n128 gnd.n125 9.3005
R11904 gnd.n7254 gnd.n129 9.3005
R11905 gnd.n7253 gnd.n130 9.3005
R11906 gnd.n7252 gnd.n131 9.3005
R11907 gnd.n135 gnd.n132 9.3005
R11908 gnd.n7247 gnd.n136 9.3005
R11909 gnd.n7246 gnd.n137 9.3005
R11910 gnd.n7242 gnd.n138 9.3005
R11911 gnd.n142 gnd.n139 9.3005
R11912 gnd.n7237 gnd.n143 9.3005
R11913 gnd.n7236 gnd.n144 9.3005
R11914 gnd.n7235 gnd.n145 9.3005
R11915 gnd.n149 gnd.n146 9.3005
R11916 gnd.n7230 gnd.n150 9.3005
R11917 gnd.n7229 gnd.n151 9.3005
R11918 gnd.n7228 gnd.n152 9.3005
R11919 gnd.n156 gnd.n153 9.3005
R11920 gnd.n7223 gnd.n157 9.3005
R11921 gnd.n7222 gnd.n158 9.3005
R11922 gnd.n7221 gnd.n159 9.3005
R11923 gnd.n163 gnd.n160 9.3005
R11924 gnd.n7216 gnd.n164 9.3005
R11925 gnd.n7215 gnd.n165 9.3005
R11926 gnd.n7214 gnd.n166 9.3005
R11927 gnd.n170 gnd.n167 9.3005
R11928 gnd.n7209 gnd.n171 9.3005
R11929 gnd.n7208 gnd.n7207 9.3005
R11930 gnd.n7206 gnd.n174 9.3005
R11931 gnd.n7276 gnd.n7275 9.3005
R11932 gnd.n2925 gnd.n2924 9.3005
R11933 gnd.n2953 gnd.n2926 9.3005
R11934 gnd.n2952 gnd.n2927 9.3005
R11935 gnd.n2951 gnd.n2928 9.3005
R11936 gnd.n2949 gnd.n2929 9.3005
R11937 gnd.n2948 gnd.n2930 9.3005
R11938 gnd.n2946 gnd.n2931 9.3005
R11939 gnd.n2945 gnd.n2932 9.3005
R11940 gnd.n2944 gnd.n2933 9.3005
R11941 gnd.n2942 gnd.n2934 9.3005
R11942 gnd.n2941 gnd.n2935 9.3005
R11943 gnd.n2939 gnd.n2936 9.3005
R11944 gnd.n2938 gnd.n2937 9.3005
R11945 gnd.n2833 gnd.n2832 9.3005
R11946 gnd.n5528 gnd.n5527 9.3005
R11947 gnd.n5529 gnd.n2831 9.3005
R11948 gnd.n5531 gnd.n5530 9.3005
R11949 gnd.n5532 gnd.n2830 9.3005
R11950 gnd.n5535 gnd.n5534 9.3005
R11951 gnd.n5536 gnd.n2829 9.3005
R11952 gnd.n5546 gnd.n5537 9.3005
R11953 gnd.n5545 gnd.n5538 9.3005
R11954 gnd.n5544 gnd.n5539 9.3005
R11955 gnd.n5543 gnd.n5541 9.3005
R11956 gnd.n5540 gnd.n294 9.3005
R11957 gnd.n6954 gnd.n295 9.3005
R11958 gnd.n6956 gnd.n6955 9.3005
R11959 gnd.n7015 gnd.n6957 9.3005
R11960 gnd.n7014 gnd.n6958 9.3005
R11961 gnd.n7013 gnd.n6959 9.3005
R11962 gnd.n7009 gnd.n6960 9.3005
R11963 gnd.n7008 gnd.n6961 9.3005
R11964 gnd.n7006 gnd.n6962 9.3005
R11965 gnd.n7005 gnd.n6963 9.3005
R11966 gnd.n7003 gnd.n6964 9.3005
R11967 gnd.n7002 gnd.n6965 9.3005
R11968 gnd.n7000 gnd.n6966 9.3005
R11969 gnd.n6999 gnd.n6967 9.3005
R11970 gnd.n6997 gnd.n6968 9.3005
R11971 gnd.n6996 gnd.n6969 9.3005
R11972 gnd.n6994 gnd.n6970 9.3005
R11973 gnd.n6993 gnd.n6971 9.3005
R11974 gnd.n6991 gnd.n6972 9.3005
R11975 gnd.n6990 gnd.n6973 9.3005
R11976 gnd.n6988 gnd.n6974 9.3005
R11977 gnd.n6987 gnd.n6975 9.3005
R11978 gnd.n6985 gnd.n6976 9.3005
R11979 gnd.n6984 gnd.n6977 9.3005
R11980 gnd.n6982 gnd.n6978 9.3005
R11981 gnd.n6981 gnd.n6980 9.3005
R11982 gnd.n6979 gnd.n178 9.3005
R11983 gnd.n7203 gnd.n177 9.3005
R11984 gnd.n7205 gnd.n7204 9.3005
R11985 gnd.n2771 gnd.n2769 9.3005
R11986 gnd.n5629 gnd.n5628 9.3005
R11987 gnd.n5630 gnd.n2763 9.3005
R11988 gnd.n5633 gnd.n2762 9.3005
R11989 gnd.n5634 gnd.n2761 9.3005
R11990 gnd.n5637 gnd.n2760 9.3005
R11991 gnd.n5638 gnd.n2759 9.3005
R11992 gnd.n5641 gnd.n2758 9.3005
R11993 gnd.n5642 gnd.n2757 9.3005
R11994 gnd.n5645 gnd.n2756 9.3005
R11995 gnd.n5646 gnd.n2755 9.3005
R11996 gnd.n5649 gnd.n2754 9.3005
R11997 gnd.n5650 gnd.n2753 9.3005
R11998 gnd.n5653 gnd.n2752 9.3005
R11999 gnd.n5654 gnd.n2751 9.3005
R12000 gnd.n5657 gnd.n2750 9.3005
R12001 gnd.n5658 gnd.n2749 9.3005
R12002 gnd.n5661 gnd.n2748 9.3005
R12003 gnd.n5662 gnd.n2747 9.3005
R12004 gnd.n5665 gnd.n2746 9.3005
R12005 gnd.n5667 gnd.n2740 9.3005
R12006 gnd.n5670 gnd.n2739 9.3005
R12007 gnd.n5671 gnd.n2738 9.3005
R12008 gnd.n5674 gnd.n2737 9.3005
R12009 gnd.n5675 gnd.n2736 9.3005
R12010 gnd.n5678 gnd.n2735 9.3005
R12011 gnd.n5679 gnd.n2734 9.3005
R12012 gnd.n5682 gnd.n2733 9.3005
R12013 gnd.n5683 gnd.n2732 9.3005
R12014 gnd.n5686 gnd.n2731 9.3005
R12015 gnd.n5687 gnd.n2730 9.3005
R12016 gnd.n5690 gnd.n2729 9.3005
R12017 gnd.n5692 gnd.n2728 9.3005
R12018 gnd.n5693 gnd.n2727 9.3005
R12019 gnd.n5694 gnd.n2726 9.3005
R12020 gnd.n5695 gnd.n2725 9.3005
R12021 gnd.n5627 gnd.n2768 9.3005
R12022 gnd.n5626 gnd.n5625 9.3005
R12023 gnd.n2921 gnd.n2920 9.3005
R12024 gnd.n2899 gnd.n2898 9.3005
R12025 gnd.n5450 gnd.n5449 9.3005
R12026 gnd.n5451 gnd.n2897 9.3005
R12027 gnd.n5455 gnd.n5452 9.3005
R12028 gnd.n5454 gnd.n5453 9.3005
R12029 gnd.n2870 gnd.n2869 9.3005
R12030 gnd.n5481 gnd.n5480 9.3005
R12031 gnd.n5482 gnd.n2868 9.3005
R12032 gnd.n5486 gnd.n5483 9.3005
R12033 gnd.n5485 gnd.n5484 9.3005
R12034 gnd.n2842 gnd.n2841 9.3005
R12035 gnd.n5518 gnd.n5517 9.3005
R12036 gnd.n5519 gnd.n2840 9.3005
R12037 gnd.n5523 gnd.n5520 9.3005
R12038 gnd.n5522 gnd.n5521 9.3005
R12039 gnd.n2808 gnd.n2807 9.3005
R12040 gnd.n5582 gnd.n5581 9.3005
R12041 gnd.n5583 gnd.n2806 9.3005
R12042 gnd.n5585 gnd.n5584 9.3005
R12043 gnd.n269 gnd.n262 9.3005
R12044 gnd.n249 gnd.n248 9.3005
R12045 gnd.n7056 gnd.n7055 9.3005
R12046 gnd.n7057 gnd.n247 9.3005
R12047 gnd.n7059 gnd.n7058 9.3005
R12048 gnd.n232 gnd.n231 9.3005
R12049 gnd.n7072 gnd.n7071 9.3005
R12050 gnd.n7073 gnd.n230 9.3005
R12051 gnd.n7075 gnd.n7074 9.3005
R12052 gnd.n219 gnd.n218 9.3005
R12053 gnd.n7088 gnd.n7087 9.3005
R12054 gnd.n7089 gnd.n217 9.3005
R12055 gnd.n7091 gnd.n7090 9.3005
R12056 gnd.n202 gnd.n201 9.3005
R12057 gnd.n7104 gnd.n7103 9.3005
R12058 gnd.n7105 gnd.n200 9.3005
R12059 gnd.n7107 gnd.n7106 9.3005
R12060 gnd.n186 gnd.n185 9.3005
R12061 gnd.n7195 gnd.n7194 9.3005
R12062 gnd.n7196 gnd.n184 9.3005
R12063 gnd.n7198 gnd.n7197 9.3005
R12064 gnd.n107 gnd.n106 9.3005
R12065 gnd.n7278 gnd.n7277 9.3005
R12066 gnd.n2919 gnd.n2918 9.3005
R12067 gnd.n7042 gnd.n267 9.3005
R12068 gnd.n7043 gnd.n7042 9.3005
R12069 gnd.n5569 gnd.n311 9.3005
R12070 gnd.n6936 gnd.n312 9.3005
R12071 gnd.n6935 gnd.n313 9.3005
R12072 gnd.n6934 gnd.n314 9.3005
R12073 gnd.n316 gnd.n315 9.3005
R12074 gnd.n6927 gnd.n318 9.3005
R12075 gnd.n6926 gnd.n319 9.3005
R12076 gnd.n6925 gnd.n320 9.3005
R12077 gnd.n3775 gnd.n3701 9.3005
R12078 gnd.n3704 gnd.n3702 9.3005
R12079 gnd.n3771 gnd.n3705 9.3005
R12080 gnd.n3770 gnd.n3706 9.3005
R12081 gnd.n3769 gnd.n3707 9.3005
R12082 gnd.n3710 gnd.n3708 9.3005
R12083 gnd.n3765 gnd.n3711 9.3005
R12084 gnd.n3764 gnd.n3712 9.3005
R12085 gnd.n3763 gnd.n3713 9.3005
R12086 gnd.n3716 gnd.n3714 9.3005
R12087 gnd.n3759 gnd.n3717 9.3005
R12088 gnd.n3758 gnd.n3718 9.3005
R12089 gnd.n3757 gnd.n3719 9.3005
R12090 gnd.n3722 gnd.n3720 9.3005
R12091 gnd.n3753 gnd.n3723 9.3005
R12092 gnd.n3752 gnd.n3724 9.3005
R12093 gnd.n3751 gnd.n3725 9.3005
R12094 gnd.n3728 gnd.n3726 9.3005
R12095 gnd.n3747 gnd.n3729 9.3005
R12096 gnd.n3746 gnd.n3730 9.3005
R12097 gnd.n3745 gnd.n3731 9.3005
R12098 gnd.n3734 gnd.n3732 9.3005
R12099 gnd.n3741 gnd.n3735 9.3005
R12100 gnd.n3740 gnd.n3736 9.3005
R12101 gnd.n3739 gnd.n3737 9.3005
R12102 gnd.n3437 gnd.n3436 9.3005
R12103 gnd.n4418 gnd.n4417 9.3005
R12104 gnd.n4419 gnd.n3435 9.3005
R12105 gnd.n4421 gnd.n4420 9.3005
R12106 gnd.n3423 gnd.n3422 9.3005
R12107 gnd.n4434 gnd.n4433 9.3005
R12108 gnd.n4435 gnd.n3421 9.3005
R12109 gnd.n4439 gnd.n4436 9.3005
R12110 gnd.n4438 gnd.n4437 9.3005
R12111 gnd.n3391 gnd.n3390 9.3005
R12112 gnd.n4558 gnd.n4557 9.3005
R12113 gnd.n4559 gnd.n3389 9.3005
R12114 gnd.n4561 gnd.n4560 9.3005
R12115 gnd.n3377 gnd.n3376 9.3005
R12116 gnd.n4574 gnd.n4573 9.3005
R12117 gnd.n4575 gnd.n3375 9.3005
R12118 gnd.n4577 gnd.n4576 9.3005
R12119 gnd.n3362 gnd.n3361 9.3005
R12120 gnd.n4590 gnd.n4589 9.3005
R12121 gnd.n4591 gnd.n3360 9.3005
R12122 gnd.n4593 gnd.n4592 9.3005
R12123 gnd.n3348 gnd.n3347 9.3005
R12124 gnd.n4605 gnd.n4604 9.3005
R12125 gnd.n4606 gnd.n3346 9.3005
R12126 gnd.n4610 gnd.n4607 9.3005
R12127 gnd.n4609 gnd.n4608 9.3005
R12128 gnd.n3316 gnd.n3315 9.3005
R12129 gnd.n4731 gnd.n4730 9.3005
R12130 gnd.n4732 gnd.n3314 9.3005
R12131 gnd.n4734 gnd.n4733 9.3005
R12132 gnd.n3302 gnd.n3301 9.3005
R12133 gnd.n4747 gnd.n4746 9.3005
R12134 gnd.n4748 gnd.n3300 9.3005
R12135 gnd.n4750 gnd.n4749 9.3005
R12136 gnd.n3289 gnd.n3288 9.3005
R12137 gnd.n4763 gnd.n4762 9.3005
R12138 gnd.n4764 gnd.n3287 9.3005
R12139 gnd.n4766 gnd.n4765 9.3005
R12140 gnd.n3278 gnd.n3277 9.3005
R12141 gnd.n4779 gnd.n4778 9.3005
R12142 gnd.n4780 gnd.n3276 9.3005
R12143 gnd.n4784 gnd.n4781 9.3005
R12144 gnd.n4783 gnd.n4782 9.3005
R12145 gnd.n3245 gnd.n3244 9.3005
R12146 gnd.n4902 gnd.n4901 9.3005
R12147 gnd.n4903 gnd.n3243 9.3005
R12148 gnd.n4905 gnd.n4904 9.3005
R12149 gnd.n3230 gnd.n3229 9.3005
R12150 gnd.n4918 gnd.n4917 9.3005
R12151 gnd.n4919 gnd.n3228 9.3005
R12152 gnd.n4921 gnd.n4920 9.3005
R12153 gnd.n3215 gnd.n3214 9.3005
R12154 gnd.n4934 gnd.n4933 9.3005
R12155 gnd.n4935 gnd.n3213 9.3005
R12156 gnd.n4937 gnd.n4936 9.3005
R12157 gnd.n3202 gnd.n3201 9.3005
R12158 gnd.n4950 gnd.n4949 9.3005
R12159 gnd.n4951 gnd.n3200 9.3005
R12160 gnd.n4955 gnd.n4952 9.3005
R12161 gnd.n4954 gnd.n4953 9.3005
R12162 gnd.n3170 gnd.n3169 9.3005
R12163 gnd.n5308 gnd.n5307 9.3005
R12164 gnd.n5309 gnd.n3168 9.3005
R12165 gnd.n5311 gnd.n5310 9.3005
R12166 gnd.n3157 gnd.n3156 9.3005
R12167 gnd.n5324 gnd.n5323 9.3005
R12168 gnd.n5325 gnd.n3155 9.3005
R12169 gnd.n5327 gnd.n5326 9.3005
R12170 gnd.n3143 gnd.n3142 9.3005
R12171 gnd.n5340 gnd.n5339 9.3005
R12172 gnd.n5341 gnd.n3141 9.3005
R12173 gnd.n5343 gnd.n5342 9.3005
R12174 gnd.n3130 gnd.n3129 9.3005
R12175 gnd.n5356 gnd.n5355 9.3005
R12176 gnd.n5357 gnd.n3128 9.3005
R12177 gnd.n5359 gnd.n5358 9.3005
R12178 gnd.n3116 gnd.n3115 9.3005
R12179 gnd.n5372 gnd.n5371 9.3005
R12180 gnd.n5373 gnd.n3114 9.3005
R12181 gnd.n5375 gnd.n5374 9.3005
R12182 gnd.n3102 gnd.n3101 9.3005
R12183 gnd.n5390 gnd.n5389 9.3005
R12184 gnd.n5391 gnd.n3100 9.3005
R12185 gnd.n5396 gnd.n5392 9.3005
R12186 gnd.n5395 gnd.n5394 9.3005
R12187 gnd.n5393 gnd.n2687 9.3005
R12188 gnd.n5704 gnd.n2688 9.3005
R12189 gnd.n5703 gnd.n2689 9.3005
R12190 gnd.n5702 gnd.n2690 9.3005
R12191 gnd.n2912 gnd.n2691 9.3005
R12192 gnd.n2913 gnd.n2911 9.3005
R12193 gnd.n2915 gnd.n2914 9.3005
R12194 gnd.n2909 gnd.n2908 9.3005
R12195 gnd.n5439 gnd.n5438 9.3005
R12196 gnd.n5440 gnd.n2907 9.3005
R12197 gnd.n5444 gnd.n5441 9.3005
R12198 gnd.n5443 gnd.n5442 9.3005
R12199 gnd.n2881 gnd.n2880 9.3005
R12200 gnd.n5470 gnd.n5469 9.3005
R12201 gnd.n5471 gnd.n2879 9.3005
R12202 gnd.n5475 gnd.n5472 9.3005
R12203 gnd.n5474 gnd.n5473 9.3005
R12204 gnd.n2853 gnd.n2852 9.3005
R12205 gnd.n5506 gnd.n5505 9.3005
R12206 gnd.n5507 gnd.n2851 9.3005
R12207 gnd.n5511 gnd.n5508 9.3005
R12208 gnd.n5510 gnd.n5509 9.3005
R12209 gnd.n2819 gnd.n2818 9.3005
R12210 gnd.n5564 gnd.n5563 9.3005
R12211 gnd.n5565 gnd.n2817 9.3005
R12212 gnd.n5576 gnd.n5566 9.3005
R12213 gnd.n5575 gnd.n5567 9.3005
R12214 gnd.n5574 gnd.n5568 9.3005
R12215 gnd.n5571 gnd.n5570 9.3005
R12216 gnd.n4349 gnd.n3610 9.3005
R12217 gnd.n4352 gnd.n3609 9.3005
R12218 gnd.n4353 gnd.n3608 9.3005
R12219 gnd.n4356 gnd.n3607 9.3005
R12220 gnd.n4357 gnd.n3606 9.3005
R12221 gnd.n4360 gnd.n3605 9.3005
R12222 gnd.n4361 gnd.n3604 9.3005
R12223 gnd.n4364 gnd.n3603 9.3005
R12224 gnd.n4365 gnd.n3602 9.3005
R12225 gnd.n4368 gnd.n3601 9.3005
R12226 gnd.n4369 gnd.n3600 9.3005
R12227 gnd.n4372 gnd.n3599 9.3005
R12228 gnd.n4373 gnd.n3598 9.3005
R12229 gnd.n4374 gnd.n3597 9.3005
R12230 gnd.n3596 gnd.n3593 9.3005
R12231 gnd.n3595 gnd.n3594 9.3005
R12232 gnd.n4138 gnd.n4137 9.3005
R12233 gnd.n4134 gnd.n3615 9.3005
R12234 gnd.n4131 gnd.n3616 9.3005
R12235 gnd.n4130 gnd.n3617 9.3005
R12236 gnd.n4127 gnd.n3618 9.3005
R12237 gnd.n4126 gnd.n3619 9.3005
R12238 gnd.n4123 gnd.n3620 9.3005
R12239 gnd.n4122 gnd.n3621 9.3005
R12240 gnd.n4119 gnd.n3622 9.3005
R12241 gnd.n4118 gnd.n3623 9.3005
R12242 gnd.n4115 gnd.n3624 9.3005
R12243 gnd.n4114 gnd.n3625 9.3005
R12244 gnd.n4111 gnd.n3626 9.3005
R12245 gnd.n4110 gnd.n3627 9.3005
R12246 gnd.n4107 gnd.n3628 9.3005
R12247 gnd.n4106 gnd.n3629 9.3005
R12248 gnd.n4103 gnd.n3630 9.3005
R12249 gnd.n4102 gnd.n3631 9.3005
R12250 gnd.n4099 gnd.n4098 9.3005
R12251 gnd.n4097 gnd.n3633 9.3005
R12252 gnd.n4139 gnd.n3611 9.3005
R12253 gnd.n3801 gnd.n3800 9.3005
R12254 gnd.n3885 gnd.n3884 9.3005
R12255 gnd.n3886 gnd.n3799 9.3005
R12256 gnd.n3889 gnd.n3887 9.3005
R12257 gnd.n3890 gnd.n3798 9.3005
R12258 gnd.n3893 gnd.n3892 9.3005
R12259 gnd.n3894 gnd.n3797 9.3005
R12260 gnd.n3897 gnd.n3895 9.3005
R12261 gnd.n3898 gnd.n3796 9.3005
R12262 gnd.n3901 gnd.n3900 9.3005
R12263 gnd.n3902 gnd.n3795 9.3005
R12264 gnd.n3905 gnd.n3903 9.3005
R12265 gnd.n3906 gnd.n3794 9.3005
R12266 gnd.n3909 gnd.n3908 9.3005
R12267 gnd.n3910 gnd.n3793 9.3005
R12268 gnd.n3913 gnd.n3911 9.3005
R12269 gnd.n3914 gnd.n3792 9.3005
R12270 gnd.n3917 gnd.n3916 9.3005
R12271 gnd.n3918 gnd.n3791 9.3005
R12272 gnd.n3921 gnd.n3919 9.3005
R12273 gnd.n3922 gnd.n3790 9.3005
R12274 gnd.n3971 gnd.n3970 9.3005
R12275 gnd.n3972 gnd.n3789 9.3005
R12276 gnd.n3974 gnd.n3973 9.3005
R12277 gnd.n3680 gnd.n3679 9.3005
R12278 gnd.n3989 gnd.n3988 9.3005
R12279 gnd.n3827 gnd.n3826 9.3005
R12280 gnd.n3832 gnd.n3831 9.3005
R12281 gnd.n3835 gnd.n3821 9.3005
R12282 gnd.n3836 gnd.n3820 9.3005
R12283 gnd.n3839 gnd.n3819 9.3005
R12284 gnd.n3840 gnd.n3818 9.3005
R12285 gnd.n3843 gnd.n3817 9.3005
R12286 gnd.n3844 gnd.n3816 9.3005
R12287 gnd.n3847 gnd.n3815 9.3005
R12288 gnd.n3848 gnd.n3814 9.3005
R12289 gnd.n3851 gnd.n3813 9.3005
R12290 gnd.n3852 gnd.n3812 9.3005
R12291 gnd.n3855 gnd.n3811 9.3005
R12292 gnd.n3856 gnd.n3810 9.3005
R12293 gnd.n3859 gnd.n3809 9.3005
R12294 gnd.n3860 gnd.n3808 9.3005
R12295 gnd.n3863 gnd.n3807 9.3005
R12296 gnd.n3866 gnd.n3865 9.3005
R12297 gnd.n3830 gnd.n3825 9.3005
R12298 gnd.n3829 gnd.n3828 9.3005
R12299 gnd.n3873 gnd.n3872 9.3005
R12300 gnd.n3871 gnd.n3806 9.3005
R12301 gnd.n3870 gnd.n3869 9.3005
R12302 gnd.n3868 gnd.n2330 9.3005
R12303 gnd.n5981 gnd.n2331 9.3005
R12304 gnd.n5980 gnd.n2332 9.3005
R12305 gnd.n5979 gnd.n2333 9.3005
R12306 gnd.n2349 gnd.n2334 9.3005
R12307 gnd.n5969 gnd.n2350 9.3005
R12308 gnd.n5968 gnd.n2351 9.3005
R12309 gnd.n5967 gnd.n2352 9.3005
R12310 gnd.n2370 gnd.n2353 9.3005
R12311 gnd.n5957 gnd.n2371 9.3005
R12312 gnd.n5956 gnd.n2372 9.3005
R12313 gnd.n5955 gnd.n2373 9.3005
R12314 gnd.n2389 gnd.n2374 9.3005
R12315 gnd.n5945 gnd.n2390 9.3005
R12316 gnd.n5944 gnd.n2391 9.3005
R12317 gnd.n5943 gnd.n2392 9.3005
R12318 gnd.n2410 gnd.n2393 9.3005
R12319 gnd.n5933 gnd.n2411 9.3005
R12320 gnd.n5932 gnd.n2412 9.3005
R12321 gnd.n5931 gnd.n2413 9.3005
R12322 gnd.n2428 gnd.n2414 9.3005
R12323 gnd.n5921 gnd.n2429 9.3005
R12324 gnd.n5920 gnd.n2430 9.3005
R12325 gnd.n5919 gnd.n2431 9.3005
R12326 gnd.n2447 gnd.n2432 9.3005
R12327 gnd.n5908 gnd.n2448 9.3005
R12328 gnd.n5907 gnd.n2449 9.3005
R12329 gnd.n5906 gnd.n2450 9.3005
R12330 gnd.n2467 gnd.n2451 9.3005
R12331 gnd.n5896 gnd.n2468 9.3005
R12332 gnd.n5895 gnd.n2469 9.3005
R12333 gnd.n5894 gnd.n2470 9.3005
R12334 gnd.n2489 gnd.n2471 9.3005
R12335 gnd.n5884 gnd.n2490 9.3005
R12336 gnd.n5883 gnd.n2491 9.3005
R12337 gnd.n5882 gnd.n2492 9.3005
R12338 gnd.n2510 gnd.n2493 9.3005
R12339 gnd.n5872 gnd.n2511 9.3005
R12340 gnd.n5871 gnd.n2512 9.3005
R12341 gnd.n5870 gnd.n2513 9.3005
R12342 gnd.n2532 gnd.n2514 9.3005
R12343 gnd.n5860 gnd.n2533 9.3005
R12344 gnd.n5859 gnd.n2534 9.3005
R12345 gnd.n5858 gnd.n2535 9.3005
R12346 gnd.n2554 gnd.n2536 9.3005
R12347 gnd.n5848 gnd.n2555 9.3005
R12348 gnd.n5847 gnd.n2556 9.3005
R12349 gnd.n5846 gnd.n2557 9.3005
R12350 gnd.n2574 gnd.n2558 9.3005
R12351 gnd.n5836 gnd.n5835 9.3005
R12352 gnd.n3867 gnd.n3805 9.3005
R12353 gnd.n5995 gnd.n5994 9.3005
R12354 gnd.n5993 gnd.n2308 9.3005
R12355 gnd.n5992 gnd.n5991 9.3005
R12356 gnd.n2310 gnd.n2309 9.3005
R12357 gnd.n3932 gnd.n3931 9.3005
R12358 gnd.n3935 gnd.n3933 9.3005
R12359 gnd.n3936 gnd.n3930 9.3005
R12360 gnd.n3939 gnd.n3938 9.3005
R12361 gnd.n3940 gnd.n3929 9.3005
R12362 gnd.n3943 gnd.n3941 9.3005
R12363 gnd.n3944 gnd.n3928 9.3005
R12364 gnd.n3947 gnd.n3946 9.3005
R12365 gnd.n3948 gnd.n3927 9.3005
R12366 gnd.n3951 gnd.n3949 9.3005
R12367 gnd.n3952 gnd.n3926 9.3005
R12368 gnd.n3955 gnd.n3954 9.3005
R12369 gnd.n3956 gnd.n3925 9.3005
R12370 gnd.n3959 gnd.n3957 9.3005
R12371 gnd.n3960 gnd.n3924 9.3005
R12372 gnd.n3963 gnd.n3962 9.3005
R12373 gnd.n3964 gnd.n3923 9.3005
R12374 gnd.n3966 gnd.n3965 9.3005
R12375 gnd.n3788 gnd.n3787 9.3005
R12376 gnd.n3979 gnd.n3978 9.3005
R12377 gnd.n3980 gnd.n3786 9.3005
R12378 gnd.n3984 gnd.n3983 9.3005
R12379 gnd.n3677 gnd.n3676 9.3005
R12380 gnd.n3998 gnd.n3997 9.3005
R12381 gnd.n3999 gnd.n3675 9.3005
R12382 gnd.n4001 gnd.n4000 9.3005
R12383 gnd.n3671 gnd.n3670 9.3005
R12384 gnd.n4014 gnd.n4013 9.3005
R12385 gnd.n4015 gnd.n3669 9.3005
R12386 gnd.n4017 gnd.n4016 9.3005
R12387 gnd.n3664 gnd.n3663 9.3005
R12388 gnd.n4030 gnd.n4029 9.3005
R12389 gnd.n4031 gnd.n3662 9.3005
R12390 gnd.n4033 gnd.n4032 9.3005
R12391 gnd.n3658 gnd.n3657 9.3005
R12392 gnd.n4046 gnd.n4045 9.3005
R12393 gnd.n4047 gnd.n3656 9.3005
R12394 gnd.n4049 gnd.n4048 9.3005
R12395 gnd.n3651 gnd.n3650 9.3005
R12396 gnd.n4062 gnd.n4061 9.3005
R12397 gnd.n4063 gnd.n3649 9.3005
R12398 gnd.n4065 gnd.n4064 9.3005
R12399 gnd.n3645 gnd.n3644 9.3005
R12400 gnd.n4078 gnd.n4077 9.3005
R12401 gnd.n4079 gnd.n3643 9.3005
R12402 gnd.n4082 gnd.n4081 9.3005
R12403 gnd.n4080 gnd.n3637 9.3005
R12404 gnd.n4094 gnd.n3636 9.3005
R12405 gnd.n4096 gnd.n4095 9.3005
R12406 gnd.n5996 gnd.n2306 9.3005
R12407 gnd.n6003 gnd.n6002 9.3005
R12408 gnd.n6004 gnd.n2300 9.3005
R12409 gnd.n6007 gnd.n2299 9.3005
R12410 gnd.n6008 gnd.n2298 9.3005
R12411 gnd.n6011 gnd.n2297 9.3005
R12412 gnd.n6012 gnd.n2296 9.3005
R12413 gnd.n6015 gnd.n2295 9.3005
R12414 gnd.n6016 gnd.n2294 9.3005
R12415 gnd.n6019 gnd.n2293 9.3005
R12416 gnd.n6020 gnd.n2292 9.3005
R12417 gnd.n6023 gnd.n2291 9.3005
R12418 gnd.n6024 gnd.n2290 9.3005
R12419 gnd.n6027 gnd.n2289 9.3005
R12420 gnd.n6028 gnd.n2288 9.3005
R12421 gnd.n6031 gnd.n2287 9.3005
R12422 gnd.n6032 gnd.n2286 9.3005
R12423 gnd.n6035 gnd.n2285 9.3005
R12424 gnd.n6036 gnd.n2284 9.3005
R12425 gnd.n6039 gnd.n2283 9.3005
R12426 gnd.n6041 gnd.n2280 9.3005
R12427 gnd.n6044 gnd.n2279 9.3005
R12428 gnd.n6045 gnd.n2278 9.3005
R12429 gnd.n6048 gnd.n2277 9.3005
R12430 gnd.n6049 gnd.n2276 9.3005
R12431 gnd.n6052 gnd.n2275 9.3005
R12432 gnd.n6053 gnd.n2274 9.3005
R12433 gnd.n6056 gnd.n2273 9.3005
R12434 gnd.n6057 gnd.n2272 9.3005
R12435 gnd.n6060 gnd.n2271 9.3005
R12436 gnd.n6061 gnd.n2270 9.3005
R12437 gnd.n6064 gnd.n2269 9.3005
R12438 gnd.n6065 gnd.n2268 9.3005
R12439 gnd.n6068 gnd.n2267 9.3005
R12440 gnd.n6070 gnd.n2266 9.3005
R12441 gnd.n6071 gnd.n2265 9.3005
R12442 gnd.n6072 gnd.n2264 9.3005
R12443 gnd.n6073 gnd.n2263 9.3005
R12444 gnd.n6001 gnd.n2305 9.3005
R12445 gnd.n6000 gnd.n5999 9.3005
R12446 gnd.n3879 gnd.n3878 9.3005
R12447 gnd.n3877 gnd.n2319 9.3005
R12448 gnd.n5987 gnd.n2320 9.3005
R12449 gnd.n5986 gnd.n2321 9.3005
R12450 gnd.n5985 gnd.n2322 9.3005
R12451 gnd.n2340 gnd.n2323 9.3005
R12452 gnd.n5975 gnd.n2341 9.3005
R12453 gnd.n5974 gnd.n2342 9.3005
R12454 gnd.n5973 gnd.n2343 9.3005
R12455 gnd.n2359 gnd.n2344 9.3005
R12456 gnd.n5963 gnd.n2360 9.3005
R12457 gnd.n5962 gnd.n2361 9.3005
R12458 gnd.n5961 gnd.n2362 9.3005
R12459 gnd.n2380 gnd.n2363 9.3005
R12460 gnd.n5951 gnd.n2381 9.3005
R12461 gnd.n5950 gnd.n2382 9.3005
R12462 gnd.n5949 gnd.n2383 9.3005
R12463 gnd.n2399 gnd.n2384 9.3005
R12464 gnd.n5939 gnd.n2400 9.3005
R12465 gnd.n5938 gnd.n2401 9.3005
R12466 gnd.n5937 gnd.n2402 9.3005
R12467 gnd.n5901 gnd.n2459 9.3005
R12468 gnd.n5900 gnd.n2460 9.3005
R12469 gnd.n2478 gnd.n2461 9.3005
R12470 gnd.n5890 gnd.n2479 9.3005
R12471 gnd.n5889 gnd.n2480 9.3005
R12472 gnd.n5888 gnd.n2481 9.3005
R12473 gnd.n2500 gnd.n2482 9.3005
R12474 gnd.n5878 gnd.n2501 9.3005
R12475 gnd.n5877 gnd.n2502 9.3005
R12476 gnd.n5876 gnd.n2503 9.3005
R12477 gnd.n2521 gnd.n2504 9.3005
R12478 gnd.n5866 gnd.n2522 9.3005
R12479 gnd.n5865 gnd.n2523 9.3005
R12480 gnd.n5864 gnd.n2524 9.3005
R12481 gnd.n2543 gnd.n2525 9.3005
R12482 gnd.n5854 gnd.n2544 9.3005
R12483 gnd.n5853 gnd.n2545 9.3005
R12484 gnd.n5852 gnd.n2546 9.3005
R12485 gnd.n2564 gnd.n2547 9.3005
R12486 gnd.n5842 gnd.n2565 9.3005
R12487 gnd.n5841 gnd.n2566 9.3005
R12488 gnd.n5840 gnd.n2567 9.3005
R12489 gnd.n3876 gnd.n3875 9.3005
R12490 gnd.n5926 gnd.n2421 9.3005
R12491 gnd.n5902 gnd.n2421 9.3005
R12492 gnd.n3691 gnd.n3683 9.3005
R12493 gnd.n3783 gnd.n3692 9.3005
R12494 gnd.n3782 gnd.n3694 9.3005
R12495 gnd.n3781 gnd.n3695 9.3005
R12496 gnd.n3698 gnd.n3696 9.3005
R12497 gnd.n3777 gnd.n3699 9.3005
R12498 gnd.n3776 gnd.n3700 9.3005
R12499 gnd.n3690 gnd.n3689 9.3005
R12500 gnd.n3684 gnd.n844 9.3005
R12501 gnd.n6158 gnd.n843 9.3005
R12502 gnd.n6159 gnd.n842 9.3005
R12503 gnd.n6160 gnd.n841 9.3005
R12504 gnd.n840 gnd.n836 9.3005
R12505 gnd.n6166 gnd.n835 9.3005
R12506 gnd.n6167 gnd.n834 9.3005
R12507 gnd.n6168 gnd.n833 9.3005
R12508 gnd.n832 gnd.n828 9.3005
R12509 gnd.n6174 gnd.n827 9.3005
R12510 gnd.n6175 gnd.n826 9.3005
R12511 gnd.n6176 gnd.n825 9.3005
R12512 gnd.n824 gnd.n820 9.3005
R12513 gnd.n6182 gnd.n819 9.3005
R12514 gnd.n6183 gnd.n818 9.3005
R12515 gnd.n6184 gnd.n817 9.3005
R12516 gnd.n816 gnd.n812 9.3005
R12517 gnd.n6190 gnd.n811 9.3005
R12518 gnd.n6191 gnd.n810 9.3005
R12519 gnd.n6192 gnd.n809 9.3005
R12520 gnd.n808 gnd.n804 9.3005
R12521 gnd.n6198 gnd.n803 9.3005
R12522 gnd.n6199 gnd.n802 9.3005
R12523 gnd.n6200 gnd.n801 9.3005
R12524 gnd.n800 gnd.n796 9.3005
R12525 gnd.n6206 gnd.n795 9.3005
R12526 gnd.n6207 gnd.n794 9.3005
R12527 gnd.n6208 gnd.n793 9.3005
R12528 gnd.n792 gnd.n788 9.3005
R12529 gnd.n6214 gnd.n787 9.3005
R12530 gnd.n6215 gnd.n786 9.3005
R12531 gnd.n6216 gnd.n785 9.3005
R12532 gnd.n784 gnd.n780 9.3005
R12533 gnd.n6222 gnd.n779 9.3005
R12534 gnd.n6223 gnd.n778 9.3005
R12535 gnd.n6224 gnd.n777 9.3005
R12536 gnd.n776 gnd.n772 9.3005
R12537 gnd.n6230 gnd.n771 9.3005
R12538 gnd.n6231 gnd.n770 9.3005
R12539 gnd.n6232 gnd.n769 9.3005
R12540 gnd.n768 gnd.n764 9.3005
R12541 gnd.n6238 gnd.n763 9.3005
R12542 gnd.n6239 gnd.n762 9.3005
R12543 gnd.n6240 gnd.n761 9.3005
R12544 gnd.n760 gnd.n756 9.3005
R12545 gnd.n6246 gnd.n755 9.3005
R12546 gnd.n6247 gnd.n754 9.3005
R12547 gnd.n6248 gnd.n753 9.3005
R12548 gnd.n752 gnd.n748 9.3005
R12549 gnd.n6254 gnd.n747 9.3005
R12550 gnd.n6255 gnd.n746 9.3005
R12551 gnd.n6256 gnd.n745 9.3005
R12552 gnd.n744 gnd.n740 9.3005
R12553 gnd.n6262 gnd.n739 9.3005
R12554 gnd.n6263 gnd.n738 9.3005
R12555 gnd.n6264 gnd.n737 9.3005
R12556 gnd.n736 gnd.n732 9.3005
R12557 gnd.n6270 gnd.n731 9.3005
R12558 gnd.n6271 gnd.n730 9.3005
R12559 gnd.n6272 gnd.n729 9.3005
R12560 gnd.n728 gnd.n724 9.3005
R12561 gnd.n6278 gnd.n723 9.3005
R12562 gnd.n6279 gnd.n722 9.3005
R12563 gnd.n6280 gnd.n721 9.3005
R12564 gnd.n720 gnd.n716 9.3005
R12565 gnd.n6286 gnd.n715 9.3005
R12566 gnd.n6287 gnd.n714 9.3005
R12567 gnd.n6288 gnd.n713 9.3005
R12568 gnd.n712 gnd.n708 9.3005
R12569 gnd.n6294 gnd.n707 9.3005
R12570 gnd.n6295 gnd.n706 9.3005
R12571 gnd.n6296 gnd.n705 9.3005
R12572 gnd.n704 gnd.n700 9.3005
R12573 gnd.n6302 gnd.n699 9.3005
R12574 gnd.n6303 gnd.n698 9.3005
R12575 gnd.n6304 gnd.n697 9.3005
R12576 gnd.n696 gnd.n692 9.3005
R12577 gnd.n6310 gnd.n691 9.3005
R12578 gnd.n6311 gnd.n690 9.3005
R12579 gnd.n6312 gnd.n689 9.3005
R12580 gnd.n688 gnd.n684 9.3005
R12581 gnd.n6318 gnd.n683 9.3005
R12582 gnd.n6319 gnd.n682 9.3005
R12583 gnd.n6320 gnd.n681 9.3005
R12584 gnd.n3686 gnd.n3685 9.3005
R12585 gnd.n3011 gnd.n3010 9.3005
R12586 gnd.n3017 gnd.n3016 9.3005
R12587 gnd.n3018 gnd.n2993 9.3005
R12588 gnd.n3027 gnd.n3026 9.3005
R12589 gnd.n2995 gnd.n2991 9.3005
R12590 gnd.n3034 gnd.n3033 9.3005
R12591 gnd.n3035 gnd.n2984 9.3005
R12592 gnd.n3044 gnd.n3043 9.3005
R12593 gnd.n2986 gnd.n2982 9.3005
R12594 gnd.n3051 gnd.n3050 9.3005
R12595 gnd.n3052 gnd.n2975 9.3005
R12596 gnd.n3061 gnd.n3060 9.3005
R12597 gnd.n2977 gnd.n2973 9.3005
R12598 gnd.n3068 gnd.n3067 9.3005
R12599 gnd.n3069 gnd.n2963 9.3005
R12600 gnd.n3076 gnd.n3075 9.3005
R12601 gnd.n2965 gnd.n2961 9.3005
R12602 gnd.n2960 gnd.n2958 9.3005
R12603 gnd.n3001 gnd.n3000 9.3005
R12604 gnd.n3071 gnd.n3070 9.3005
R12605 gnd.n2972 gnd.n2969 9.3005
R12606 gnd.n3059 gnd.n3058 9.3005
R12607 gnd.n3055 gnd.n2976 9.3005
R12608 gnd.n3054 gnd.n3053 9.3005
R12609 gnd.n2981 gnd.n2978 9.3005
R12610 gnd.n3042 gnd.n3041 9.3005
R12611 gnd.n3038 gnd.n2985 9.3005
R12612 gnd.n3037 gnd.n3036 9.3005
R12613 gnd.n2990 gnd.n2987 9.3005
R12614 gnd.n3025 gnd.n3024 9.3005
R12615 gnd.n3021 gnd.n2994 9.3005
R12616 gnd.n3020 gnd.n3019 9.3005
R12617 gnd.n2999 gnd.n2996 9.3005
R12618 gnd.n3009 gnd.n3008 9.3005
R12619 gnd.n3005 gnd.n3004 9.3005
R12620 gnd.n3072 gnd.n2964 9.3005
R12621 gnd.n3074 gnd.n3073 9.3005
R12622 gnd.n5426 gnd.n5425 9.3005
R12623 gnd.n5424 gnd.n2959 9.3005
R12624 gnd.n5423 gnd.n5422 9.3005
R12625 gnd.n5421 gnd.n3086 9.3005
R12626 gnd.n5420 gnd.n5419 9.3005
R12627 gnd.n5418 gnd.n3087 9.3005
R12628 gnd.n5414 gnd.n5413 9.3005
R12629 gnd.n5412 gnd.n3094 9.3005
R12630 gnd.n5411 gnd.n5410 9.3005
R12631 gnd.n5409 gnd.n5404 9.3005
R12632 gnd.n4427 gnd.n3429 9.3005
R12633 gnd.n4429 gnd.n4428 9.3005
R12634 gnd.n3415 gnd.n3414 9.3005
R12635 gnd.n4444 gnd.n4443 9.3005
R12636 gnd.n4445 gnd.n3412 9.3005
R12637 gnd.n4448 gnd.n4447 9.3005
R12638 gnd.n4446 gnd.n3413 9.3005
R12639 gnd.n3384 gnd.n3383 9.3005
R12640 gnd.n4566 gnd.n4565 9.3005
R12641 gnd.n4567 gnd.n3382 9.3005
R12642 gnd.n4569 gnd.n4568 9.3005
R12643 gnd.n3370 gnd.n3369 9.3005
R12644 gnd.n4582 gnd.n4581 9.3005
R12645 gnd.n4583 gnd.n3368 9.3005
R12646 gnd.n4585 gnd.n4584 9.3005
R12647 gnd.n3356 gnd.n3355 9.3005
R12648 gnd.n4598 gnd.n4597 9.3005
R12649 gnd.n4599 gnd.n3354 9.3005
R12650 gnd.n4601 gnd.n4600 9.3005
R12651 gnd.n3340 gnd.n3339 9.3005
R12652 gnd.n4615 gnd.n4614 9.3005
R12653 gnd.n4616 gnd.n3337 9.3005
R12654 gnd.n4619 gnd.n4618 9.3005
R12655 gnd.n4617 gnd.n3338 9.3005
R12656 gnd.n3309 gnd.n3308 9.3005
R12657 gnd.n4739 gnd.n4738 9.3005
R12658 gnd.n4740 gnd.n3307 9.3005
R12659 gnd.n4742 gnd.n4741 9.3005
R12660 gnd.n3296 gnd.n3295 9.3005
R12661 gnd.n4755 gnd.n4754 9.3005
R12662 gnd.n4756 gnd.n3294 9.3005
R12663 gnd.n4758 gnd.n4757 9.3005
R12664 gnd.n3284 gnd.n3283 9.3005
R12665 gnd.n4771 gnd.n4770 9.3005
R12666 gnd.n4772 gnd.n3282 9.3005
R12667 gnd.n4774 gnd.n4773 9.3005
R12668 gnd.n3270 gnd.n3269 9.3005
R12669 gnd.n4789 gnd.n4788 9.3005
R12670 gnd.n4790 gnd.n3267 9.3005
R12671 gnd.n4793 gnd.n4792 9.3005
R12672 gnd.n4791 gnd.n3268 9.3005
R12673 gnd.n3237 gnd.n3236 9.3005
R12674 gnd.n4910 gnd.n4909 9.3005
R12675 gnd.n4911 gnd.n3235 9.3005
R12676 gnd.n4913 gnd.n4912 9.3005
R12677 gnd.n3222 gnd.n3221 9.3005
R12678 gnd.n4926 gnd.n4925 9.3005
R12679 gnd.n4927 gnd.n3220 9.3005
R12680 gnd.n4929 gnd.n4928 9.3005
R12681 gnd.n3208 gnd.n3207 9.3005
R12682 gnd.n4942 gnd.n4941 9.3005
R12683 gnd.n4943 gnd.n3206 9.3005
R12684 gnd.n4945 gnd.n4944 9.3005
R12685 gnd.n3193 gnd.n3192 9.3005
R12686 gnd.n4960 gnd.n4959 9.3005
R12687 gnd.n4961 gnd.n3190 9.3005
R12688 gnd.n4964 gnd.n4963 9.3005
R12689 gnd.n4962 gnd.n3191 9.3005
R12690 gnd.n3163 gnd.n3162 9.3005
R12691 gnd.n5316 gnd.n5315 9.3005
R12692 gnd.n5317 gnd.n3161 9.3005
R12693 gnd.n5319 gnd.n5318 9.3005
R12694 gnd.n3150 gnd.n3149 9.3005
R12695 gnd.n5332 gnd.n5331 9.3005
R12696 gnd.n5333 gnd.n3148 9.3005
R12697 gnd.n5335 gnd.n5334 9.3005
R12698 gnd.n3137 gnd.n3136 9.3005
R12699 gnd.n5348 gnd.n5347 9.3005
R12700 gnd.n5349 gnd.n3135 9.3005
R12701 gnd.n5351 gnd.n5350 9.3005
R12702 gnd.n3123 gnd.n3122 9.3005
R12703 gnd.n5364 gnd.n5363 9.3005
R12704 gnd.n5365 gnd.n3121 9.3005
R12705 gnd.n5367 gnd.n5366 9.3005
R12706 gnd.n3109 gnd.n3108 9.3005
R12707 gnd.n5380 gnd.n5379 9.3005
R12708 gnd.n5381 gnd.n3106 9.3005
R12709 gnd.n5385 gnd.n5384 9.3005
R12710 gnd.n5383 gnd.n3107 9.3005
R12711 gnd.n5382 gnd.n3096 9.3005
R12712 gnd.n5401 gnd.n3095 9.3005
R12713 gnd.n5403 gnd.n5402 9.3005
R12714 gnd.n4426 gnd.n4425 9.3005
R12715 gnd.n4412 gnd.n4411 9.3005
R12716 gnd.n4410 gnd.n3454 9.3005
R12717 gnd.n4409 gnd.n4408 9.3005
R12718 gnd.n4405 gnd.n3456 9.3005
R12719 gnd.n4402 gnd.n4401 9.3005
R12720 gnd.n4400 gnd.n3459 9.3005
R12721 gnd.n4399 gnd.n4398 9.3005
R12722 gnd.n4395 gnd.n3460 9.3005
R12723 gnd.n4392 gnd.n4391 9.3005
R12724 gnd.n3455 gnd.n3430 9.3005
R12725 gnd.n3991 gnd.n3678 9.3005
R12726 gnd.n3993 gnd.n3992 9.3005
R12727 gnd.n3674 gnd.n3673 9.3005
R12728 gnd.n4006 gnd.n4005 9.3005
R12729 gnd.n4007 gnd.n3672 9.3005
R12730 gnd.n4009 gnd.n4008 9.3005
R12731 gnd.n3667 gnd.n3666 9.3005
R12732 gnd.n4022 gnd.n4021 9.3005
R12733 gnd.n4023 gnd.n3665 9.3005
R12734 gnd.n4025 gnd.n4024 9.3005
R12735 gnd.n3661 gnd.n3660 9.3005
R12736 gnd.n4038 gnd.n4037 9.3005
R12737 gnd.n4039 gnd.n3659 9.3005
R12738 gnd.n4041 gnd.n4040 9.3005
R12739 gnd.n3654 gnd.n3653 9.3005
R12740 gnd.n4054 gnd.n4053 9.3005
R12741 gnd.n4055 gnd.n3652 9.3005
R12742 gnd.n4057 gnd.n4056 9.3005
R12743 gnd.n3648 gnd.n3647 9.3005
R12744 gnd.n4070 gnd.n4069 9.3005
R12745 gnd.n4071 gnd.n3646 9.3005
R12746 gnd.n4073 gnd.n4072 9.3005
R12747 gnd.n3642 gnd.n3641 9.3005
R12748 gnd.n4087 gnd.n4086 9.3005
R12749 gnd.n4088 gnd.n3639 9.3005
R12750 gnd.n4090 gnd.n4089 9.3005
R12751 gnd.n3640 gnd.n3462 9.3005
R12752 gnd.n4389 gnd.n3461 9.3005
R12753 gnd.n4388 gnd.n4387 9.3005
R12754 gnd.n4384 gnd.n4383 9.3005
R12755 gnd.n3467 gnd.n3464 9.3005
R12756 gnd.n3566 gnd.n3565 9.3005
R12757 gnd.n3562 gnd.n3482 9.3005
R12758 gnd.n3561 gnd.n3560 9.3005
R12759 gnd.n3487 gnd.n3484 9.3005
R12760 gnd.n3552 gnd.n3551 9.3005
R12761 gnd.n3548 gnd.n3547 9.3005
R12762 gnd.n3491 gnd.n3490 9.3005
R12763 gnd.n3540 gnd.n3539 9.3005
R12764 gnd.n3536 gnd.n3535 9.3005
R12765 gnd.n3499 gnd.n3496 9.3005
R12766 gnd.n3528 gnd.n3527 9.3005
R12767 gnd.n3524 gnd.n3523 9.3005
R12768 gnd.n3503 gnd.n3502 9.3005
R12769 gnd.n3516 gnd.n3515 9.3005
R12770 gnd.n3512 gnd.n3510 9.3005
R12771 gnd.n3505 gnd.n2576 9.3005
R12772 gnd.n3509 gnd.n3506 9.3005
R12773 gnd.n3518 gnd.n3517 9.3005
R12774 gnd.n3522 gnd.n3521 9.3005
R12775 gnd.n3501 gnd.n3500 9.3005
R12776 gnd.n3530 gnd.n3529 9.3005
R12777 gnd.n3534 gnd.n3533 9.3005
R12778 gnd.n3495 gnd.n3492 9.3005
R12779 gnd.n3542 gnd.n3541 9.3005
R12780 gnd.n3546 gnd.n3545 9.3005
R12781 gnd.n3489 gnd.n3488 9.3005
R12782 gnd.n3554 gnd.n3553 9.3005
R12783 gnd.n3558 gnd.n3557 9.3005
R12784 gnd.n3559 gnd.n3481 9.3005
R12785 gnd.n3568 gnd.n3567 9.3005
R12786 gnd.n3483 gnd.n3468 9.3005
R12787 gnd.n4382 gnd.n4381 9.3005
R12788 gnd.n4380 gnd.n3463 9.3005
R12789 gnd.n5830 gnd.n2577 9.3005
R12790 gnd.n5829 gnd.n5828 9.3005
R12791 gnd.n5827 gnd.n2581 9.3005
R12792 gnd.n5826 gnd.n5825 9.3005
R12793 gnd.n5824 gnd.n2582 9.3005
R12794 gnd.n5823 gnd.n5822 9.3005
R12795 gnd.n5821 gnd.n2586 9.3005
R12796 gnd.n5820 gnd.n5819 9.3005
R12797 gnd.n5818 gnd.n2587 9.3005
R12798 gnd.n5817 gnd.n5816 9.3005
R12799 gnd.n5815 gnd.n2591 9.3005
R12800 gnd.n5814 gnd.n5813 9.3005
R12801 gnd.n5812 gnd.n2592 9.3005
R12802 gnd.n5811 gnd.n5810 9.3005
R12803 gnd.n5809 gnd.n2596 9.3005
R12804 gnd.n5808 gnd.n5807 9.3005
R12805 gnd.n5806 gnd.n2597 9.3005
R12806 gnd.n5805 gnd.n5804 9.3005
R12807 gnd.n5803 gnd.n2601 9.3005
R12808 gnd.n5802 gnd.n5801 9.3005
R12809 gnd.n5800 gnd.n2602 9.3005
R12810 gnd.n5799 gnd.n5798 9.3005
R12811 gnd.n5797 gnd.n2606 9.3005
R12812 gnd.n5796 gnd.n5795 9.3005
R12813 gnd.n5794 gnd.n2607 9.3005
R12814 gnd.n5793 gnd.n5792 9.3005
R12815 gnd.n5791 gnd.n2611 9.3005
R12816 gnd.n5790 gnd.n5789 9.3005
R12817 gnd.n5788 gnd.n2612 9.3005
R12818 gnd.n5787 gnd.n5786 9.3005
R12819 gnd.n5785 gnd.n2616 9.3005
R12820 gnd.n5784 gnd.n5783 9.3005
R12821 gnd.n5782 gnd.n2617 9.3005
R12822 gnd.n5781 gnd.n5780 9.3005
R12823 gnd.n5779 gnd.n2621 9.3005
R12824 gnd.n5778 gnd.n5777 9.3005
R12825 gnd.n5776 gnd.n2622 9.3005
R12826 gnd.n5775 gnd.n5774 9.3005
R12827 gnd.n5773 gnd.n2626 9.3005
R12828 gnd.n5772 gnd.n5771 9.3005
R12829 gnd.n5770 gnd.n2627 9.3005
R12830 gnd.n5769 gnd.n5768 9.3005
R12831 gnd.n5767 gnd.n2631 9.3005
R12832 gnd.n5766 gnd.n5765 9.3005
R12833 gnd.n5764 gnd.n2632 9.3005
R12834 gnd.n5763 gnd.n5762 9.3005
R12835 gnd.n5761 gnd.n2636 9.3005
R12836 gnd.n5760 gnd.n5759 9.3005
R12837 gnd.n5758 gnd.n2637 9.3005
R12838 gnd.n5757 gnd.n5756 9.3005
R12839 gnd.n5755 gnd.n2641 9.3005
R12840 gnd.n5754 gnd.n5753 9.3005
R12841 gnd.n5752 gnd.n2642 9.3005
R12842 gnd.n5751 gnd.n5750 9.3005
R12843 gnd.n5749 gnd.n2646 9.3005
R12844 gnd.n5748 gnd.n5747 9.3005
R12845 gnd.n5746 gnd.n2647 9.3005
R12846 gnd.n5745 gnd.n5744 9.3005
R12847 gnd.n5743 gnd.n2651 9.3005
R12848 gnd.n5742 gnd.n5741 9.3005
R12849 gnd.n5740 gnd.n2652 9.3005
R12850 gnd.n5739 gnd.n5738 9.3005
R12851 gnd.n5737 gnd.n2656 9.3005
R12852 gnd.n5736 gnd.n5735 9.3005
R12853 gnd.n5734 gnd.n2657 9.3005
R12854 gnd.n5733 gnd.n5732 9.3005
R12855 gnd.n5731 gnd.n2661 9.3005
R12856 gnd.n5730 gnd.n5729 9.3005
R12857 gnd.n5728 gnd.n2662 9.3005
R12858 gnd.n5727 gnd.n5726 9.3005
R12859 gnd.n5725 gnd.n2666 9.3005
R12860 gnd.n5724 gnd.n5723 9.3005
R12861 gnd.n5722 gnd.n2667 9.3005
R12862 gnd.n5721 gnd.n5720 9.3005
R12863 gnd.n5719 gnd.n2671 9.3005
R12864 gnd.n5718 gnd.n5717 9.3005
R12865 gnd.n5716 gnd.n2672 9.3005
R12866 gnd.n5715 gnd.n5714 9.3005
R12867 gnd.n5713 gnd.n2676 9.3005
R12868 gnd.n5712 gnd.n5711 9.3005
R12869 gnd.n5710 gnd.n2677 9.3005
R12870 gnd.n5709 gnd.n2680 9.3005
R12871 gnd.n5832 gnd.n5831 9.3005
R12872 gnd.n5618 gnd.n2777 9.3005
R12873 gnd.n5617 gnd.n5616 9.3005
R12874 gnd.n5615 gnd.n2779 9.3005
R12875 gnd.n5614 gnd.n5613 9.3005
R12876 gnd.n5612 gnd.n2783 9.3005
R12877 gnd.n5611 gnd.n5610 9.3005
R12878 gnd.n5609 gnd.n2784 9.3005
R12879 gnd.n5608 gnd.n5607 9.3005
R12880 gnd.n5606 gnd.n2788 9.3005
R12881 gnd.n5605 gnd.n5604 9.3005
R12882 gnd.n5603 gnd.n2789 9.3005
R12883 gnd.n5602 gnd.n5601 9.3005
R12884 gnd.n5600 gnd.n2793 9.3005
R12885 gnd.n5599 gnd.n5598 9.3005
R12886 gnd.n5597 gnd.n2794 9.3005
R12887 gnd.n5596 gnd.n5595 9.3005
R12888 gnd.n5594 gnd.n2798 9.3005
R12889 gnd.n5593 gnd.n5592 9.3005
R12890 gnd.n5591 gnd.n2799 9.3005
R12891 gnd.n5590 gnd.n5589 9.3005
R12892 gnd.n280 gnd.n278 9.3005
R12893 gnd.n7036 gnd.n7035 9.3005
R12894 gnd.n7034 gnd.n279 9.3005
R12895 gnd.n7033 gnd.n7032 9.3005
R12896 gnd.n7031 gnd.n281 9.3005
R12897 gnd.n7030 gnd.n7029 9.3005
R12898 gnd.n7027 gnd.n285 9.3005
R12899 gnd.n7026 gnd.n7025 9.3005
R12900 gnd.n7024 gnd.n287 9.3005
R12901 gnd.n256 gnd.n255 9.3005
R12902 gnd.n7048 gnd.n7047 9.3005
R12903 gnd.n7049 gnd.n254 9.3005
R12904 gnd.n7051 gnd.n7050 9.3005
R12905 gnd.n241 gnd.n240 9.3005
R12906 gnd.n7064 gnd.n7063 9.3005
R12907 gnd.n7065 gnd.n239 9.3005
R12908 gnd.n7067 gnd.n7066 9.3005
R12909 gnd.n226 gnd.n225 9.3005
R12910 gnd.n7080 gnd.n7079 9.3005
R12911 gnd.n7081 gnd.n224 9.3005
R12912 gnd.n7083 gnd.n7082 9.3005
R12913 gnd.n211 gnd.n210 9.3005
R12914 gnd.n7096 gnd.n7095 9.3005
R12915 gnd.n7097 gnd.n209 9.3005
R12916 gnd.n7099 gnd.n7098 9.3005
R12917 gnd.n196 gnd.n195 9.3005
R12918 gnd.n7112 gnd.n7111 9.3005
R12919 gnd.n7113 gnd.n193 9.3005
R12920 gnd.n7190 gnd.n7189 9.3005
R12921 gnd.n7188 gnd.n194 9.3005
R12922 gnd.n7187 gnd.n7186 9.3005
R12923 gnd.n7185 gnd.n7114 9.3005
R12924 gnd.n7184 gnd.n7183 9.3005
R12925 gnd.n5620 gnd.n5619 9.3005
R12926 gnd.n7180 gnd.n7116 9.3005
R12927 gnd.n7179 gnd.n7178 9.3005
R12928 gnd.n7177 gnd.n7121 9.3005
R12929 gnd.n7176 gnd.n7175 9.3005
R12930 gnd.n7174 gnd.n7122 9.3005
R12931 gnd.n7173 gnd.n7172 9.3005
R12932 gnd.n7171 gnd.n7129 9.3005
R12933 gnd.n7170 gnd.n7169 9.3005
R12934 gnd.n7168 gnd.n7130 9.3005
R12935 gnd.n7167 gnd.n7166 9.3005
R12936 gnd.n7165 gnd.n7137 9.3005
R12937 gnd.n7164 gnd.n7163 9.3005
R12938 gnd.n7162 gnd.n7138 9.3005
R12939 gnd.n7161 gnd.n7160 9.3005
R12940 gnd.n7159 gnd.n7145 9.3005
R12941 gnd.n7158 gnd.n7157 9.3005
R12942 gnd.n7156 gnd.n7146 9.3005
R12943 gnd.n7155 gnd.n7154 9.3005
R12944 gnd.n7182 gnd.n7181 9.3005
R12945 gnd.n5430 gnd.n2956 9.3005
R12946 gnd.n5433 gnd.n5432 9.3005
R12947 gnd.n5431 gnd.n2957 9.3005
R12948 gnd.n2889 gnd.n2888 9.3005
R12949 gnd.n5460 gnd.n5459 9.3005
R12950 gnd.n5461 gnd.n2886 9.3005
R12951 gnd.n5464 gnd.n5463 9.3005
R12952 gnd.n5462 gnd.n2887 9.3005
R12953 gnd.n2861 gnd.n2860 9.3005
R12954 gnd.n5491 gnd.n5490 9.3005
R12955 gnd.n5492 gnd.n2858 9.3005
R12956 gnd.n5500 gnd.n5499 9.3005
R12957 gnd.n5498 gnd.n2859 9.3005
R12958 gnd.n5497 gnd.n5496 9.3005
R12959 gnd.n5495 gnd.n5493 9.3005
R12960 gnd.n2826 gnd.n2824 9.3005
R12961 gnd.n5557 gnd.n5556 9.3005
R12962 gnd.n5555 gnd.n2825 9.3005
R12963 gnd.n5554 gnd.n5553 9.3005
R12964 gnd.n5552 gnd.n2827 9.3005
R12965 gnd.n5551 gnd.n5550 9.3005
R12966 gnd.n306 gnd.n305 9.3005
R12967 gnd.n6942 gnd.n6941 9.3005
R12968 gnd.n6943 gnd.n304 9.3005
R12969 gnd.n6945 gnd.n6944 9.3005
R12970 gnd.n65 gnd.n63 9.3005
R12971 gnd.n7321 gnd.n7320 9.3005
R12972 gnd.n7319 gnd.n64 9.3005
R12973 gnd.n7318 gnd.n7317 9.3005
R12974 gnd.n7316 gnd.n69 9.3005
R12975 gnd.n7315 gnd.n7314 9.3005
R12976 gnd.n7313 gnd.n70 9.3005
R12977 gnd.n7312 gnd.n7311 9.3005
R12978 gnd.n7310 gnd.n74 9.3005
R12979 gnd.n7309 gnd.n7308 9.3005
R12980 gnd.n7307 gnd.n75 9.3005
R12981 gnd.n7306 gnd.n7305 9.3005
R12982 gnd.n7304 gnd.n79 9.3005
R12983 gnd.n7303 gnd.n7302 9.3005
R12984 gnd.n7301 gnd.n80 9.3005
R12985 gnd.n7300 gnd.n7299 9.3005
R12986 gnd.n7298 gnd.n84 9.3005
R12987 gnd.n7297 gnd.n7296 9.3005
R12988 gnd.n7295 gnd.n85 9.3005
R12989 gnd.n7294 gnd.n7293 9.3005
R12990 gnd.n7292 gnd.n89 9.3005
R12991 gnd.n7291 gnd.n7290 9.3005
R12992 gnd.n7289 gnd.n90 9.3005
R12993 gnd.n7288 gnd.n7287 9.3005
R12994 gnd.n7286 gnd.n94 9.3005
R12995 gnd.n7285 gnd.n7284 9.3005
R12996 gnd.n7283 gnd.n95 9.3005
R12997 gnd.n7282 gnd.n98 9.3005
R12998 gnd.n5429 gnd.n5428 9.3005
R12999 gnd.t306 gnd.n1324 9.24152
R13000 gnd.n6146 gnd.t100 9.24152
R13001 gnd.n2220 gnd.t92 9.24152
R13002 gnd.t72 gnd.n2313 9.24152
R13003 gnd.n5844 gnd.t47 9.24152
R13004 gnd.t37 gnd.n5435 9.24152
R13005 gnd.n7200 gnd.t30 9.24152
R13006 gnd.t292 gnd.t306 8.92286
R13007 gnd.n4441 gnd.n3418 8.92286
R13008 gnd.n4612 gnd.n3343 8.92286
R13009 gnd.n4720 gnd.n3329 8.92286
R13010 gnd.n4786 gnd.n3273 8.92286
R13011 gnd.n4891 gnd.n3258 8.92286
R13012 gnd.n4957 gnd.n3197 8.92286
R13013 gnd.n5297 gnd.n3181 8.92286
R13014 gnd.n5361 gnd.n3126 8.92286
R13015 gnd.n5387 gnd.n3104 8.92286
R13016 gnd.n1228 gnd.n1203 8.92171
R13017 gnd.n1196 gnd.n1171 8.92171
R13018 gnd.n1164 gnd.n1139 8.92171
R13019 gnd.n1133 gnd.n1108 8.92171
R13020 gnd.n1101 gnd.n1076 8.92171
R13021 gnd.n1069 gnd.n1044 8.92171
R13022 gnd.n1037 gnd.n1012 8.92171
R13023 gnd.n1006 gnd.n981 8.92171
R13024 gnd.n5053 gnd.n5035 8.72777
R13025 gnd.n1968 gnd.t308 8.60421
R13026 gnd.n4431 gnd.n3427 8.60421
R13027 gnd.n4675 gnd.t153 8.60421
R13028 gnd.t131 gnd.n3241 8.60421
R13029 gnd.n1396 gnd.n1380 8.43467
R13030 gnd.n46 gnd.n30 8.43467
R13031 gnd.n3990 gnd.n0 8.41456
R13032 gnd.n7323 gnd.n7322 8.41456
R13033 gnd.n3426 gnd.t104 8.28555
R13034 gnd.n1229 gnd.n1201 8.14595
R13035 gnd.n1197 gnd.n1169 8.14595
R13036 gnd.n1165 gnd.n1137 8.14595
R13037 gnd.n1134 gnd.n1106 8.14595
R13038 gnd.n1102 gnd.n1074 8.14595
R13039 gnd.n1070 gnd.n1042 8.14595
R13040 gnd.n1038 gnd.n1010 8.14595
R13041 gnd.n1007 gnd.n979 8.14595
R13042 gnd.n1234 gnd.n1233 7.97301
R13043 gnd.t309 gnd.n1483 7.9669
R13044 gnd.n4525 gnd.t322 7.9669
R13045 gnd.t288 gnd.n3146 7.9669
R13046 gnd.n7156 gnd.n7155 7.75808
R13047 gnd.n3073 gnd.n3072 7.75808
R13048 gnd.n4381 gnd.n4380 7.75808
R13049 gnd.n3828 gnd.n3825 7.75808
R13050 gnd.n3395 gnd.t122 7.64824
R13051 gnd.n4540 gnd.n4539 7.64824
R13052 gnd.t6 gnd.n3352 7.64824
R13053 gnd.n4696 gnd.t136 7.64824
R13054 gnd.n4768 gnd.t136 7.64824
R13055 gnd.n4814 gnd.t7 7.64824
R13056 gnd.t7 gnd.n3217 7.64824
R13057 gnd.n5290 gnd.t298 7.64824
R13058 gnd.n5353 gnd.n3133 7.64824
R13059 gnd.n5016 gnd.t110 7.64824
R13060 gnd.n1877 gnd.t314 7.32958
R13061 gnd.t296 gnd.t55 7.32958
R13062 gnd.n4182 gnd.n4181 7.30353
R13063 gnd.n5052 gnd.n5051 7.30353
R13064 gnd.n1837 gnd.n1556 7.01093
R13065 gnd.n1559 gnd.n1557 7.01093
R13066 gnd.n1847 gnd.n1846 7.01093
R13067 gnd.n1858 gnd.n1540 7.01093
R13068 gnd.n1857 gnd.n1543 7.01093
R13069 gnd.n1868 gnd.n1531 7.01093
R13070 gnd.n1534 gnd.n1532 7.01093
R13071 gnd.n1878 gnd.n1877 7.01093
R13072 gnd.n1888 gnd.n1512 7.01093
R13073 gnd.n1887 gnd.n1515 7.01093
R13074 gnd.n1896 gnd.n1506 7.01093
R13075 gnd.n1908 gnd.n1496 7.01093
R13076 gnd.n1918 gnd.n1481 7.01093
R13077 gnd.n1934 gnd.n1933 7.01093
R13078 gnd.n1483 gnd.n1420 7.01093
R13079 gnd.n1988 gnd.n1421 7.01093
R13080 gnd.n1982 gnd.n1981 7.01093
R13081 gnd.n1470 gnd.n1432 7.01093
R13082 gnd.n1974 gnd.n1443 7.01093
R13083 gnd.n1461 gnd.n1456 7.01093
R13084 gnd.n1968 gnd.n1967 7.01093
R13085 gnd.n2014 gnd.n1359 7.01093
R13086 gnd.n2013 gnd.n2012 7.01093
R13087 gnd.n2025 gnd.n2024 7.01093
R13088 gnd.n1352 gnd.n1344 7.01093
R13089 gnd.n2054 gnd.n1332 7.01093
R13090 gnd.n2053 gnd.n1335 7.01093
R13091 gnd.n2064 gnd.n1324 7.01093
R13092 gnd.n1325 gnd.n1313 7.01093
R13093 gnd.n2075 gnd.n1314 7.01093
R13094 gnd.n2099 gnd.n1305 7.01093
R13095 gnd.n2098 gnd.n1296 7.01093
R13096 gnd.n2121 gnd.n2120 7.01093
R13097 gnd.n2139 gnd.n1277 7.01093
R13098 gnd.n2138 gnd.n1280 7.01093
R13099 gnd.n2149 gnd.n1269 7.01093
R13100 gnd.n1270 gnd.n1257 7.01093
R13101 gnd.n2162 gnd.n1258 7.01093
R13102 gnd.n2185 gnd.n1243 7.01093
R13103 gnd.n2201 gnd.n2200 7.01093
R13104 gnd.n2179 gnd.n846 7.01093
R13105 gnd.n6154 gnd.n846 7.01093
R13106 gnd.n6153 gnd.n848 7.01093
R13107 gnd.n2175 gnd.n857 7.01093
R13108 gnd.n6147 gnd.n6146 7.01093
R13109 gnd.n2221 gnd.n2220 7.01093
R13110 gnd.n6140 gnd.n868 7.01093
R13111 gnd.n6139 gnd.n871 7.01093
R13112 gnd.n4776 gnd.t140 7.01093
R13113 gnd.t299 gnd.n4883 7.01093
R13114 gnd.n5387 gnd.t76 7.01093
R13115 gnd.n1515 gnd.t301 6.69227
R13116 gnd.n1335 gnd.t292 6.69227
R13117 gnd.n2186 gnd.t307 6.69227
R13118 gnd.n5971 gnd.t229 6.69227
R13119 gnd.n4059 gnd.t176 6.69227
R13120 gnd.t159 gnd.n2538 6.69227
R13121 gnd.n4509 gnd.t8 6.69227
R13122 gnd.n5321 gnd.t151 6.69227
R13123 gnd.n5467 gnd.t233 6.69227
R13124 gnd.n2876 gnd.t186 6.69227
R13125 gnd.t190 gnd.n204 6.69227
R13126 gnd.n5222 gnd.n5221 6.5566
R13127 gnd.n4340 gnd.n4339 6.5566
R13128 gnd.n4208 gnd.n4202 6.5566
R13129 gnd.n5134 gnd.n5133 6.5566
R13130 gnd.n4532 gnd.n4468 6.37362
R13131 gnd.n4595 gnd.n3358 6.37362
R13132 gnd.n4705 gnd.n4642 6.37362
R13133 gnd.n4939 gnd.n3211 6.37362
R13134 gnd.n5282 gnd.n4988 6.37362
R13135 gnd.n5345 gnd.n3139 6.37362
R13136 gnd.t20 gnd.n3112 6.37362
R13137 gnd.n4408 gnd.n4406 6.20656
R13138 gnd.n7245 gnd.n7242 6.20656
R13139 gnd.n6040 gnd.n6039 6.20656
R13140 gnd.n5417 gnd.n5414 6.20656
R13141 gnd.t129 gnd.n1944 6.05496
R13142 gnd.n1945 gnd.t300 6.05496
R13143 gnd.t149 gnd.n1359 6.05496
R13144 gnd.t311 gnd.n2109 6.05496
R13145 gnd.n5947 gnd.t198 6.05496
R13146 gnd.n4027 gnd.t188 6.05496
R13147 gnd.t157 gnd.n2495 6.05496
R13148 gnd.n2849 gnd.t165 6.05496
R13149 gnd.n5560 gnd.t217 6.05496
R13150 gnd.t255 gnd.n234 6.05496
R13151 gnd.n1231 gnd.n1201 5.81868
R13152 gnd.n1199 gnd.n1169 5.81868
R13153 gnd.n1167 gnd.n1137 5.81868
R13154 gnd.n1136 gnd.n1106 5.81868
R13155 gnd.n1104 gnd.n1074 5.81868
R13156 gnd.n1072 gnd.n1042 5.81868
R13157 gnd.n1040 gnd.n1010 5.81868
R13158 gnd.n1009 gnd.n979 5.81868
R13159 gnd.n4547 gnd.t34 5.73631
R13160 gnd.t141 gnd.n3343 5.73631
R13161 gnd.t142 gnd.n3291 5.73631
R13162 gnd.n4867 gnd.t285 5.73631
R13163 gnd.n5297 gnd.t135 5.73631
R13164 gnd.n5231 gnd.t76 5.73631
R13165 gnd.n5226 gnd.n2741 5.62001
R13166 gnd.n4347 gnd.n4141 5.62001
R13167 gnd.n4347 gnd.n4142 5.62001
R13168 gnd.n5138 gnd.n2741 5.62001
R13169 gnd.n1696 gnd.n1691 5.4308
R13170 gnd.n972 gnd.n902 5.4308
R13171 gnd.n2012 gnd.t310 5.41765
R13172 gnd.t312 gnd.n2035 5.41765
R13173 gnd.t318 gnd.n1289 5.41765
R13174 gnd.n5923 gnd.t161 5.41765
R13175 gnd.t202 gnd.n2437 5.41765
R13176 gnd.n3995 gnd.t202 5.41765
R13177 gnd.t171 gnd.n2453 5.41765
R13178 gnd.t316 gnd.n3319 5.41765
R13179 gnd.n4966 gnd.t294 5.41765
R13180 gnd.t181 gnd.n275 5.41765
R13181 gnd.n6947 gnd.t236 5.41765
R13182 gnd.t236 gnd.n297 5.41765
R13183 gnd.n7017 gnd.t242 5.41765
R13184 gnd.n4587 gnd.n3366 5.09899
R13185 gnd.n4525 gnd.n4524 5.09899
R13186 gnd.t127 gnd.n4712 5.09899
R13187 gnd.n4760 gnd.n3292 5.09899
R13188 gnd.n4698 gnd.n4697 5.09899
R13189 gnd.n4931 gnd.n3218 5.09899
R13190 gnd.n4869 gnd.n4868 5.09899
R13191 gnd.n4947 gnd.t139 5.09899
R13192 gnd.n5337 gnd.n3146 5.09899
R13193 gnd.n5275 gnd.n5274 5.09899
R13194 gnd.n1229 gnd.n1228 5.04292
R13195 gnd.n1197 gnd.n1196 5.04292
R13196 gnd.n1165 gnd.n1164 5.04292
R13197 gnd.n1134 gnd.n1133 5.04292
R13198 gnd.n1102 gnd.n1101 5.04292
R13199 gnd.n1070 gnd.n1069 5.04292
R13200 gnd.n1038 gnd.n1037 5.04292
R13201 gnd.n1007 gnd.n1006 5.04292
R13202 gnd.n1412 gnd.n1411 4.82753
R13203 gnd.n62 gnd.n61 4.82753
R13204 gnd.n1975 gnd.t315 4.78034
R13205 gnd.n1314 gnd.t304 4.78034
R13206 gnd.n2405 gnd.t169 4.78034
R13207 gnd.n3968 gnd.n2408 4.78034
R13208 gnd.n5898 gnd.t163 4.78034
R13209 gnd.t188 gnd.n2476 4.78034
R13210 gnd.n3320 gnd.t316 4.78034
R13211 gnd.t294 gnd.n3172 4.78034
R13212 gnd.n5229 gnd.t44 4.78034
R13213 gnd.t217 gnd.n2810 4.78034
R13214 gnd.n5587 gnd.t194 4.78034
R13215 gnd.n7045 gnd.n259 4.78034
R13216 gnd.n7053 gnd.t248 4.78034
R13217 gnd.n1417 gnd.n1414 4.74817
R13218 gnd.n1467 gnd.n1365 4.74817
R13219 gnd.n1454 gnd.n1364 4.74817
R13220 gnd.n1363 gnd.n1362 4.74817
R13221 gnd.n1463 gnd.n1414 4.74817
R13222 gnd.n1464 gnd.n1365 4.74817
R13223 gnd.n1466 gnd.n1364 4.74817
R13224 gnd.n1453 gnd.n1363 4.74817
R13225 gnd.n7041 gnd.n7040 4.74817
R13226 gnd.n6950 gnd.n266 4.74817
R13227 gnd.n7019 gnd.n265 4.74817
R13228 gnd.n264 gnd.n261 4.74817
R13229 gnd.n7041 gnd.n268 4.74817
R13230 gnd.n301 gnd.n266 4.74817
R13231 gnd.n6949 gnd.n265 4.74817
R13232 gnd.n7020 gnd.n264 4.74817
R13233 gnd.n2420 gnd.n2403 4.74817
R13234 gnd.n2439 gnd.n2422 4.74817
R13235 gnd.n5914 gnd.n5913 4.74817
R13236 gnd.n2458 gnd.n2440 4.74817
R13237 gnd.n5927 gnd.n2420 4.74817
R13238 gnd.n5925 gnd.n2422 4.74817
R13239 gnd.n5915 gnd.n5914 4.74817
R13240 gnd.n5912 gnd.n2440 4.74817
R13241 gnd.n1396 gnd.n1395 4.7074
R13242 gnd.n46 gnd.n45 4.7074
R13243 gnd.n1412 gnd.n1396 4.65959
R13244 gnd.n62 gnd.n46 4.65959
R13245 gnd.n5666 gnd.n2743 4.6132
R13246 gnd.n4348 gnd.n4140 4.6132
R13247 gnd.n4377 gnd.n3472 4.46168
R13248 gnd.n4540 gnd.t291 4.46168
R13249 gnd.t18 gnd.n3133 4.46168
R13250 gnd.n5698 gnd.n2721 4.46168
R13251 gnd.n5048 gnd.n5035 4.46111
R13252 gnd.n1214 gnd.n1210 4.38594
R13253 gnd.n1182 gnd.n1178 4.38594
R13254 gnd.n1150 gnd.n1146 4.38594
R13255 gnd.n1119 gnd.n1115 4.38594
R13256 gnd.n1087 gnd.n1083 4.38594
R13257 gnd.n1055 gnd.n1051 4.38594
R13258 gnd.n1023 gnd.n1019 4.38594
R13259 gnd.n992 gnd.n988 4.38594
R13260 gnd.n1225 gnd.n1203 4.26717
R13261 gnd.n1193 gnd.n1171 4.26717
R13262 gnd.n1161 gnd.n1139 4.26717
R13263 gnd.n1130 gnd.n1108 4.26717
R13264 gnd.n1098 gnd.n1076 4.26717
R13265 gnd.n1066 gnd.n1044 4.26717
R13266 gnd.n1034 gnd.n1012 4.26717
R13267 gnd.n1003 gnd.n981 4.26717
R13268 gnd.n1919 gnd.t305 4.14303
R13269 gnd.n2149 gnd.t302 4.14303
R13270 gnd.n2365 gnd.t167 4.14303
R13271 gnd.n5874 gnd.t174 4.14303
R13272 gnd.t176 gnd.n2519 4.14303
R13273 gnd.n4656 gnd.t147 4.14303
R13274 gnd.n4876 gnd.t133 4.14303
R13275 gnd.t186 gnd.n2863 4.14303
R13276 gnd.t251 gnd.n5502 4.14303
R13277 gnd.n7085 gnd.t204 4.14303
R13278 gnd.n1233 gnd.n1232 4.08274
R13279 gnd.n5221 gnd.n5220 4.05904
R13280 gnd.n4339 gnd.n4338 4.05904
R13281 gnd.n4212 gnd.n4202 4.05904
R13282 gnd.n5133 gnd.n5132 4.05904
R13283 gnd.n15 gnd.n7 3.99943
R13284 gnd.t122 gnd.n3386 3.82437
R13285 gnd.n4579 gnd.n3373 3.82437
R13286 gnd.n4517 gnd.n4483 3.82437
R13287 gnd.n4752 gnd.n3298 3.82437
R13288 gnd.n4690 gnd.n4658 3.82437
R13289 gnd.n4923 gnd.n3226 3.82437
R13290 gnd.n4861 gnd.n4829 3.82437
R13291 gnd.n5329 gnd.n3153 3.82437
R13292 gnd.n5267 gnd.n5004 3.82437
R13293 gnd.n5398 gnd.t44 3.82437
R13294 gnd.n1233 gnd.n1105 3.70378
R13295 gnd.n1992 gnd.n1413 3.65935
R13296 gnd.n15 gnd.n14 3.60163
R13297 gnd.n1224 gnd.n1205 3.49141
R13298 gnd.n1192 gnd.n1173 3.49141
R13299 gnd.n1160 gnd.n1141 3.49141
R13300 gnd.n1129 gnd.n1110 3.49141
R13301 gnd.n1097 gnd.n1078 3.49141
R13302 gnd.n1065 gnd.n1046 3.49141
R13303 gnd.n1033 gnd.n1014 3.49141
R13304 gnd.n1002 gnd.n983 3.49141
R13305 gnd.n3405 gnd.t34 3.18706
R13306 gnd.n5244 gnd.t89 3.18706
R13307 gnd.n1498 gnd.t305 2.8684
R13308 gnd.n1397 gnd.t269 2.82907
R13309 gnd.n1397 gnd.t222 2.82907
R13310 gnd.n1399 gnd.t257 2.82907
R13311 gnd.n1399 gnd.t158 2.82907
R13312 gnd.n1401 gnd.t180 2.82907
R13313 gnd.n1401 gnd.t164 2.82907
R13314 gnd.n1403 gnd.t162 2.82907
R13315 gnd.n1403 gnd.t278 2.82907
R13316 gnd.n1405 gnd.t170 2.82907
R13317 gnd.n1405 gnd.t214 2.82907
R13318 gnd.n1407 gnd.t246 2.82907
R13319 gnd.n1407 gnd.t199 2.82907
R13320 gnd.n1409 gnd.t230 2.82907
R13321 gnd.n1409 gnd.t168 2.82907
R13322 gnd.n1366 gnd.t175 2.82907
R13323 gnd.n1366 gnd.t200 2.82907
R13324 gnd.n1368 gnd.t213 2.82907
R13325 gnd.n1368 gnd.t271 2.82907
R13326 gnd.n1370 gnd.t193 2.82907
R13327 gnd.n1370 gnd.t185 2.82907
R13328 gnd.n1372 gnd.t235 2.82907
R13329 gnd.n1372 gnd.t223 2.82907
R13330 gnd.n1374 gnd.t275 2.82907
R13331 gnd.n1374 gnd.t206 2.82907
R13332 gnd.n1376 gnd.t219 2.82907
R13333 gnd.n1376 gnd.t247 2.82907
R13334 gnd.n1378 gnd.t260 2.82907
R13335 gnd.n1378 gnd.t192 2.82907
R13336 gnd.n1381 gnd.t277 2.82907
R13337 gnd.n1381 gnd.t177 2.82907
R13338 gnd.n1383 gnd.t189 2.82907
R13339 gnd.n1383 gnd.t250 2.82907
R13340 gnd.n1385 gnd.t172 2.82907
R13341 gnd.n1385 gnd.t283 2.82907
R13342 gnd.n1387 gnd.t212 2.82907
R13343 gnd.n1387 gnd.t203 2.82907
R13344 gnd.n1389 gnd.t261 2.82907
R13345 gnd.n1389 gnd.t184 2.82907
R13346 gnd.n1391 gnd.t197 2.82907
R13347 gnd.n1391 gnd.t221 2.82907
R13348 gnd.n1393 gnd.t238 2.82907
R13349 gnd.n1393 gnd.t173 2.82907
R13350 gnd.n59 gnd.t226 2.82907
R13351 gnd.n59 gnd.t191 2.82907
R13352 gnd.n57 gnd.t284 2.82907
R13353 gnd.n57 gnd.t208 2.82907
R13354 gnd.n55 gnd.t179 2.82907
R13355 gnd.n55 gnd.t276 2.82907
R13356 gnd.n53 gnd.t253 2.82907
R13357 gnd.n53 gnd.t264 2.82907
R13358 gnd.n51 gnd.t266 2.82907
R13359 gnd.n51 gnd.t281 2.82907
R13360 gnd.n49 gnd.t262 2.82907
R13361 gnd.n49 gnd.t218 2.82907
R13362 gnd.n47 gnd.t187 2.82907
R13363 gnd.n47 gnd.t252 2.82907
R13364 gnd.n28 gnd.t225 2.82907
R13365 gnd.n28 gnd.t279 2.82907
R13366 gnd.n26 gnd.t273 2.82907
R13367 gnd.n26 gnd.t254 2.82907
R13368 gnd.n24 gnd.t239 2.82907
R13369 gnd.n24 gnd.t270 2.82907
R13370 gnd.n22 gnd.t259 2.82907
R13371 gnd.n22 gnd.t267 2.82907
R13372 gnd.n20 gnd.t216 2.82907
R13373 gnd.n20 gnd.t182 2.82907
R13374 gnd.n18 gnd.t166 2.82907
R13375 gnd.n18 gnd.t245 2.82907
R13376 gnd.n16 gnd.t231 2.82907
R13377 gnd.n16 gnd.t282 2.82907
R13378 gnd.n43 gnd.t205 2.82907
R13379 gnd.n43 gnd.t268 2.82907
R13380 gnd.n41 gnd.t256 2.82907
R13381 gnd.n41 gnd.t228 2.82907
R13382 gnd.n39 gnd.t215 2.82907
R13383 gnd.n39 gnd.t249 2.82907
R13384 gnd.n37 gnd.t237 2.82907
R13385 gnd.n37 gnd.t243 2.82907
R13386 gnd.n35 gnd.t195 2.82907
R13387 gnd.n35 gnd.t280 2.82907
R13388 gnd.n33 gnd.t274 2.82907
R13389 gnd.n33 gnd.t220 2.82907
R13390 gnd.n31 gnd.t209 2.82907
R13391 gnd.n31 gnd.t272 2.82907
R13392 gnd.n1221 gnd.n1220 2.71565
R13393 gnd.n1189 gnd.n1188 2.71565
R13394 gnd.n1157 gnd.n1156 2.71565
R13395 gnd.n1126 gnd.n1125 2.71565
R13396 gnd.n1094 gnd.n1093 2.71565
R13397 gnd.n1062 gnd.n1061 2.71565
R13398 gnd.n1030 gnd.n1029 2.71565
R13399 gnd.n999 gnd.n998 2.71565
R13400 gnd.n4571 gnd.n3380 2.54975
R13401 gnd.n4468 gnd.t12 2.54975
R13402 gnd.n4510 gnd.n4509 2.54975
R13403 gnd.n4728 gnd.t5 2.54975
R13404 gnd.n4744 gnd.n3305 2.54975
R13405 gnd.n4713 gnd.t127 2.54975
R13406 gnd.n4683 gnd.n4682 2.54975
R13407 gnd.n4915 gnd.n3233 2.54975
R13408 gnd.n4855 gnd.t139 2.54975
R13409 gnd.n4854 gnd.n4853 2.54975
R13410 gnd.n5305 gnd.t4 2.54975
R13411 gnd.n5321 gnd.n3159 2.54975
R13412 gnd.n5345 gnd.t15 2.54975
R13413 gnd.n5260 gnd.n5259 2.54975
R13414 gnd.n1992 gnd.n1414 2.27742
R13415 gnd.n1992 gnd.n1365 2.27742
R13416 gnd.n1992 gnd.n1364 2.27742
R13417 gnd.n1992 gnd.n1363 2.27742
R13418 gnd.n7042 gnd.n7041 2.27742
R13419 gnd.n7042 gnd.n266 2.27742
R13420 gnd.n7042 gnd.n265 2.27742
R13421 gnd.n7042 gnd.n264 2.27742
R13422 gnd.n2421 gnd.n2420 2.27742
R13423 gnd.n2422 gnd.n2421 2.27742
R13424 gnd.n5914 gnd.n2421 2.27742
R13425 gnd.n2440 gnd.n2421 2.27742
R13426 gnd.n1846 gnd.t23 2.23109
R13427 gnd.n1469 gnd.t315 2.23109
R13428 gnd.n4768 gnd.t147 2.23109
R13429 gnd.t133 gnd.n4814 2.23109
R13430 gnd.n1217 gnd.n1207 1.93989
R13431 gnd.n1185 gnd.n1175 1.93989
R13432 gnd.n1153 gnd.n1143 1.93989
R13433 gnd.n1122 gnd.n1112 1.93989
R13434 gnd.n1090 gnd.n1080 1.93989
R13435 gnd.n1058 gnd.n1048 1.93989
R13436 gnd.n1026 gnd.n1016 1.93989
R13437 gnd.n995 gnd.n985 1.93989
R13438 gnd.t137 gnd.n1857 1.59378
R13439 gnd.n2036 gnd.t312 1.59378
R13440 gnd.n1298 gnd.t318 1.59378
R13441 gnd.n4272 gnd.t27 1.27512
R13442 gnd.n4272 gnd.n4162 1.27512
R13443 gnd.n4563 gnd.n3387 1.27512
R13444 gnd.n4502 gnd.n4496 1.27512
R13445 gnd.n4736 gnd.n3312 1.27512
R13446 gnd.n4675 gnd.n3264 1.27512
R13447 gnd.n4907 gnd.n3241 1.27512
R13448 gnd.n4846 gnd.n3187 1.27512
R13449 gnd.n5313 gnd.n3166 1.27512
R13450 gnd.n5251 gnd.n5016 1.27512
R13451 gnd.n5237 gnd.n5030 1.27512
R13452 gnd.n7192 gnd.n190 1.27512
R13453 gnd.n1699 gnd.n1691 1.16414
R13454 gnd.n969 gnd.n902 1.16414
R13455 gnd.n1216 gnd.n1209 1.16414
R13456 gnd.n1184 gnd.n1177 1.16414
R13457 gnd.n1152 gnd.n1145 1.16414
R13458 gnd.n1121 gnd.n1114 1.16414
R13459 gnd.n1089 gnd.n1082 1.16414
R13460 gnd.n1057 gnd.n1050 1.16414
R13461 gnd.n1025 gnd.n1018 1.16414
R13462 gnd.n994 gnd.n987 1.16414
R13463 gnd.n5666 gnd.n5665 0.970197
R13464 gnd.n4348 gnd.n3611 0.970197
R13465 gnd.n1200 gnd.n1168 0.962709
R13466 gnd.n1232 gnd.n1200 0.962709
R13467 gnd.n1073 gnd.n1041 0.962709
R13468 gnd.n1105 gnd.n1073 0.962709
R13469 gnd.n1945 gnd.t129 0.956468
R13470 gnd.n2110 gnd.t311 0.956468
R13471 gnd.n4451 gnd.t296 0.956468
R13472 gnd.n4571 gnd.t2 0.956468
R13473 gnd.n5259 gnd.t286 0.956468
R13474 gnd.t145 gnd.n3111 0.956468
R13475 gnd.n1406 gnd.n1404 0.773756
R13476 gnd.n56 gnd.n54 0.773756
R13477 gnd.n1411 gnd.n1410 0.773756
R13478 gnd.n1410 gnd.n1408 0.773756
R13479 gnd.n1408 gnd.n1406 0.773756
R13480 gnd.n1404 gnd.n1402 0.773756
R13481 gnd.n1402 gnd.n1400 0.773756
R13482 gnd.n1400 gnd.n1398 0.773756
R13483 gnd.n50 gnd.n48 0.773756
R13484 gnd.n52 gnd.n50 0.773756
R13485 gnd.n54 gnd.n52 0.773756
R13486 gnd.n58 gnd.n56 0.773756
R13487 gnd.n60 gnd.n58 0.773756
R13488 gnd.n61 gnd.n60 0.773756
R13489 gnd.n2 gnd.n1 0.672012
R13490 gnd.n3 gnd.n2 0.672012
R13491 gnd.n4 gnd.n3 0.672012
R13492 gnd.n5 gnd.n4 0.672012
R13493 gnd.n6 gnd.n5 0.672012
R13494 gnd.n7 gnd.n6 0.672012
R13495 gnd.n9 gnd.n8 0.672012
R13496 gnd.n10 gnd.n9 0.672012
R13497 gnd.n11 gnd.n10 0.672012
R13498 gnd.n12 gnd.n11 0.672012
R13499 gnd.n13 gnd.n12 0.672012
R13500 gnd.n14 gnd.n13 0.672012
R13501 gnd.n4555 gnd.t58 0.637812
R13502 gnd.n4523 gnd.t16 0.637812
R13503 gnd.n4684 gnd.t140 0.637812
R13504 gnd.n4884 gnd.t299 0.637812
R13505 gnd.t128 gnd.n3145 0.637812
R13506 gnd.n5244 gnd.t51 0.637812
R13507 gnd gnd.n0 0.59317
R13508 gnd.n1380 gnd.n1379 0.573776
R13509 gnd.n1379 gnd.n1377 0.573776
R13510 gnd.n1377 gnd.n1375 0.573776
R13511 gnd.n1375 gnd.n1373 0.573776
R13512 gnd.n1373 gnd.n1371 0.573776
R13513 gnd.n1371 gnd.n1369 0.573776
R13514 gnd.n1369 gnd.n1367 0.573776
R13515 gnd.n1395 gnd.n1394 0.573776
R13516 gnd.n1394 gnd.n1392 0.573776
R13517 gnd.n1392 gnd.n1390 0.573776
R13518 gnd.n1390 gnd.n1388 0.573776
R13519 gnd.n1388 gnd.n1386 0.573776
R13520 gnd.n1386 gnd.n1384 0.573776
R13521 gnd.n1384 gnd.n1382 0.573776
R13522 gnd.n19 gnd.n17 0.573776
R13523 gnd.n21 gnd.n19 0.573776
R13524 gnd.n23 gnd.n21 0.573776
R13525 gnd.n25 gnd.n23 0.573776
R13526 gnd.n27 gnd.n25 0.573776
R13527 gnd.n29 gnd.n27 0.573776
R13528 gnd.n30 gnd.n29 0.573776
R13529 gnd.n34 gnd.n32 0.573776
R13530 gnd.n36 gnd.n34 0.573776
R13531 gnd.n38 gnd.n36 0.573776
R13532 gnd.n40 gnd.n38 0.573776
R13533 gnd.n42 gnd.n40 0.573776
R13534 gnd.n44 gnd.n42 0.573776
R13535 gnd.n45 gnd.n44 0.573776
R13536 gnd.n7324 gnd.n7323 0.553533
R13537 gnd.n7042 gnd.n263 0.5435
R13538 gnd.n3693 gnd.n2421 0.5435
R13539 gnd.n5833 gnd.n5832 0.523366
R13540 gnd.n3003 gnd.n2680 0.523366
R13541 gnd.n3829 gnd.n3827 0.505073
R13542 gnd.n3867 gnd.n3866 0.505073
R13543 gnd.n7183 gnd.n7182 0.505073
R13544 gnd.n7154 gnd.n98 0.505073
R13545 gnd.n7277 gnd.n7276 0.492878
R13546 gnd.n7206 gnd.n7205 0.492878
R13547 gnd.n5626 gnd.n2769 0.492878
R13548 gnd.n2919 gnd.n2725 0.492878
R13549 gnd.n3595 gnd.n2567 0.492878
R13550 gnd.n4097 gnd.n4096 0.492878
R13551 gnd.n6000 gnd.n2306 0.492878
R13552 gnd.n3876 gnd.n2263 0.492878
R13553 gnd.n5404 gnd.n5403 0.489829
R13554 gnd.n4426 gnd.n3430 0.489829
R13555 gnd.n2227 gnd.n2226 0.486781
R13556 gnd.n1748 gnd.n1747 0.48678
R13557 gnd.n6085 gnd.n6084 0.480683
R13558 gnd.n1832 gnd.n1831 0.480683
R13559 gnd.n681 gnd.n676 0.459342
R13560 gnd.n6710 gnd.n6709 0.459342
R13561 gnd.n6921 gnd.n320 0.459342
R13562 gnd.n3690 gnd.n3685 0.459342
R13563 gnd.n5835 gnd.n5834 0.404992
R13564 gnd.n5619 gnd.n2778 0.404992
R13565 gnd.n4406 gnd.n4405 0.388379
R13566 gnd.n1213 gnd.n1212 0.388379
R13567 gnd.n1181 gnd.n1180 0.388379
R13568 gnd.n1149 gnd.n1148 0.388379
R13569 gnd.n1118 gnd.n1117 0.388379
R13570 gnd.n1086 gnd.n1085 0.388379
R13571 gnd.n1054 gnd.n1053 0.388379
R13572 gnd.n1022 gnd.n1021 0.388379
R13573 gnd.n991 gnd.n990 0.388379
R13574 gnd.n7246 gnd.n7245 0.388379
R13575 gnd.n6041 gnd.n6040 0.388379
R13576 gnd.n5418 gnd.n5417 0.388379
R13577 gnd.n7324 gnd.n15 0.374463
R13578 gnd.n1260 gnd.t307 0.319156
R13579 gnd.n4711 gnd.t13 0.319156
R13580 gnd.t153 gnd.t290 0.319156
R13581 gnd.t11 gnd.t131 0.319156
R13582 gnd.t0 gnd.n3204 0.319156
R13583 gnd.n1666 gnd.n1644 0.311721
R13584 gnd gnd.n7324 0.295112
R13585 gnd.n4390 gnd.n3462 0.27489
R13586 gnd.n5429 gnd.n5427 0.27489
R13587 gnd.n6130 gnd.n876 0.268793
R13588 gnd.n916 gnd.n876 0.241354
R13589 gnd.n2743 gnd.n2740 0.229039
R13590 gnd.n2746 gnd.n2743 0.229039
R13591 gnd.n4140 gnd.n3610 0.229039
R13592 gnd.n4140 gnd.n4139 0.229039
R13593 gnd.n1820 gnd.n1619 0.206293
R13594 gnd.n1413 gnd.n0 0.169152
R13595 gnd.n1230 gnd.n1202 0.155672
R13596 gnd.n1223 gnd.n1202 0.155672
R13597 gnd.n1223 gnd.n1222 0.155672
R13598 gnd.n1222 gnd.n1206 0.155672
R13599 gnd.n1215 gnd.n1206 0.155672
R13600 gnd.n1215 gnd.n1214 0.155672
R13601 gnd.n1198 gnd.n1170 0.155672
R13602 gnd.n1191 gnd.n1170 0.155672
R13603 gnd.n1191 gnd.n1190 0.155672
R13604 gnd.n1190 gnd.n1174 0.155672
R13605 gnd.n1183 gnd.n1174 0.155672
R13606 gnd.n1183 gnd.n1182 0.155672
R13607 gnd.n1166 gnd.n1138 0.155672
R13608 gnd.n1159 gnd.n1138 0.155672
R13609 gnd.n1159 gnd.n1158 0.155672
R13610 gnd.n1158 gnd.n1142 0.155672
R13611 gnd.n1151 gnd.n1142 0.155672
R13612 gnd.n1151 gnd.n1150 0.155672
R13613 gnd.n1135 gnd.n1107 0.155672
R13614 gnd.n1128 gnd.n1107 0.155672
R13615 gnd.n1128 gnd.n1127 0.155672
R13616 gnd.n1127 gnd.n1111 0.155672
R13617 gnd.n1120 gnd.n1111 0.155672
R13618 gnd.n1120 gnd.n1119 0.155672
R13619 gnd.n1103 gnd.n1075 0.155672
R13620 gnd.n1096 gnd.n1075 0.155672
R13621 gnd.n1096 gnd.n1095 0.155672
R13622 gnd.n1095 gnd.n1079 0.155672
R13623 gnd.n1088 gnd.n1079 0.155672
R13624 gnd.n1088 gnd.n1087 0.155672
R13625 gnd.n1071 gnd.n1043 0.155672
R13626 gnd.n1064 gnd.n1043 0.155672
R13627 gnd.n1064 gnd.n1063 0.155672
R13628 gnd.n1063 gnd.n1047 0.155672
R13629 gnd.n1056 gnd.n1047 0.155672
R13630 gnd.n1056 gnd.n1055 0.155672
R13631 gnd.n1039 gnd.n1011 0.155672
R13632 gnd.n1032 gnd.n1011 0.155672
R13633 gnd.n1032 gnd.n1031 0.155672
R13634 gnd.n1031 gnd.n1015 0.155672
R13635 gnd.n1024 gnd.n1015 0.155672
R13636 gnd.n1024 gnd.n1023 0.155672
R13637 gnd.n1008 gnd.n980 0.155672
R13638 gnd.n1001 gnd.n980 0.155672
R13639 gnd.n1001 gnd.n1000 0.155672
R13640 gnd.n1000 gnd.n984 0.155672
R13641 gnd.n993 gnd.n984 0.155672
R13642 gnd.n993 gnd.n992 0.155672
R13643 gnd.n6119 gnd.n6085 0.152939
R13644 gnd.n6119 gnd.n6118 0.152939
R13645 gnd.n6118 gnd.n6117 0.152939
R13646 gnd.n6117 gnd.n6087 0.152939
R13647 gnd.n6088 gnd.n6087 0.152939
R13648 gnd.n6089 gnd.n6088 0.152939
R13649 gnd.n6090 gnd.n6089 0.152939
R13650 gnd.n6091 gnd.n6090 0.152939
R13651 gnd.n6092 gnd.n6091 0.152939
R13652 gnd.n6093 gnd.n6092 0.152939
R13653 gnd.n6094 gnd.n6093 0.152939
R13654 gnd.n6095 gnd.n6094 0.152939
R13655 gnd.n6095 gnd.n882 0.152939
R13656 gnd.n6128 gnd.n882 0.152939
R13657 gnd.n6129 gnd.n6128 0.152939
R13658 gnd.n6130 gnd.n6129 0.152939
R13659 gnd.n1833 gnd.n1832 0.152939
R13660 gnd.n1833 gnd.n1537 0.152939
R13661 gnd.n1861 gnd.n1537 0.152939
R13662 gnd.n1862 gnd.n1861 0.152939
R13663 gnd.n1863 gnd.n1862 0.152939
R13664 gnd.n1864 gnd.n1863 0.152939
R13665 gnd.n1864 gnd.n1509 0.152939
R13666 gnd.n1891 gnd.n1509 0.152939
R13667 gnd.n1892 gnd.n1891 0.152939
R13668 gnd.n1893 gnd.n1892 0.152939
R13669 gnd.n1893 gnd.n1487 0.152939
R13670 gnd.n1922 gnd.n1487 0.152939
R13671 gnd.n1923 gnd.n1922 0.152939
R13672 gnd.n1924 gnd.n1923 0.152939
R13673 gnd.n1925 gnd.n1924 0.152939
R13674 gnd.n1927 gnd.n1925 0.152939
R13675 gnd.n1927 gnd.n1926 0.152939
R13676 gnd.n1926 gnd.n1436 0.152939
R13677 gnd.n1437 gnd.n1436 0.152939
R13678 gnd.n1438 gnd.n1437 0.152939
R13679 gnd.n1457 gnd.n1438 0.152939
R13680 gnd.n1458 gnd.n1457 0.152939
R13681 gnd.n1458 gnd.n1356 0.152939
R13682 gnd.n2017 gnd.n1356 0.152939
R13683 gnd.n2018 gnd.n2017 0.152939
R13684 gnd.n2019 gnd.n2018 0.152939
R13685 gnd.n2020 gnd.n2019 0.152939
R13686 gnd.n2020 gnd.n1329 0.152939
R13687 gnd.n2057 gnd.n1329 0.152939
R13688 gnd.n2058 gnd.n2057 0.152939
R13689 gnd.n2059 gnd.n2058 0.152939
R13690 gnd.n2060 gnd.n2059 0.152939
R13691 gnd.n2060 gnd.n1302 0.152939
R13692 gnd.n2102 gnd.n1302 0.152939
R13693 gnd.n2103 gnd.n2102 0.152939
R13694 gnd.n2104 gnd.n2103 0.152939
R13695 gnd.n2105 gnd.n2104 0.152939
R13696 gnd.n2105 gnd.n1274 0.152939
R13697 gnd.n2142 gnd.n1274 0.152939
R13698 gnd.n2143 gnd.n2142 0.152939
R13699 gnd.n2144 gnd.n2143 0.152939
R13700 gnd.n2145 gnd.n2144 0.152939
R13701 gnd.n2145 gnd.n1248 0.152939
R13702 gnd.n2189 gnd.n1248 0.152939
R13703 gnd.n2190 gnd.n2189 0.152939
R13704 gnd.n2191 gnd.n2190 0.152939
R13705 gnd.n2192 gnd.n2191 0.152939
R13706 gnd.n2194 gnd.n2192 0.152939
R13707 gnd.n2194 gnd.n2193 0.152939
R13708 gnd.n2193 gnd.n863 0.152939
R13709 gnd.n864 gnd.n863 0.152939
R13710 gnd.n865 gnd.n864 0.152939
R13711 gnd.n6084 gnd.n865 0.152939
R13712 gnd.n1831 gnd.n1561 0.152939
R13713 gnd.n1582 gnd.n1561 0.152939
R13714 gnd.n1583 gnd.n1582 0.152939
R13715 gnd.n1589 gnd.n1583 0.152939
R13716 gnd.n1590 gnd.n1589 0.152939
R13717 gnd.n1591 gnd.n1590 0.152939
R13718 gnd.n1591 gnd.n1580 0.152939
R13719 gnd.n1599 gnd.n1580 0.152939
R13720 gnd.n1600 gnd.n1599 0.152939
R13721 gnd.n1601 gnd.n1600 0.152939
R13722 gnd.n1601 gnd.n1578 0.152939
R13723 gnd.n1609 gnd.n1578 0.152939
R13724 gnd.n1610 gnd.n1609 0.152939
R13725 gnd.n1611 gnd.n1610 0.152939
R13726 gnd.n1611 gnd.n1576 0.152939
R13727 gnd.n1619 gnd.n1576 0.152939
R13728 gnd.n917 gnd.n916 0.152939
R13729 gnd.n918 gnd.n917 0.152939
R13730 gnd.n918 gnd.n912 0.152939
R13731 gnd.n926 gnd.n912 0.152939
R13732 gnd.n927 gnd.n926 0.152939
R13733 gnd.n928 gnd.n927 0.152939
R13734 gnd.n928 gnd.n910 0.152939
R13735 gnd.n936 gnd.n910 0.152939
R13736 gnd.n937 gnd.n936 0.152939
R13737 gnd.n938 gnd.n937 0.152939
R13738 gnd.n938 gnd.n908 0.152939
R13739 gnd.n946 gnd.n908 0.152939
R13740 gnd.n947 gnd.n946 0.152939
R13741 gnd.n948 gnd.n947 0.152939
R13742 gnd.n948 gnd.n906 0.152939
R13743 gnd.n956 gnd.n906 0.152939
R13744 gnd.n957 gnd.n956 0.152939
R13745 gnd.n958 gnd.n957 0.152939
R13746 gnd.n958 gnd.n904 0.152939
R13747 gnd.n966 gnd.n904 0.152939
R13748 gnd.n967 gnd.n966 0.152939
R13749 gnd.n968 gnd.n967 0.152939
R13750 gnd.n968 gnd.n899 0.152939
R13751 gnd.n975 gnd.n899 0.152939
R13752 gnd.n976 gnd.n975 0.152939
R13753 gnd.n2227 gnd.n976 0.152939
R13754 gnd.n1994 gnd.n1993 0.152939
R13755 gnd.n1995 gnd.n1994 0.152939
R13756 gnd.n1996 gnd.n1995 0.152939
R13757 gnd.n1997 gnd.n1996 0.152939
R13758 gnd.n1998 gnd.n1997 0.152939
R13759 gnd.n1999 gnd.n1998 0.152939
R13760 gnd.n1999 gnd.n1310 0.152939
R13761 gnd.n2078 gnd.n1310 0.152939
R13762 gnd.n2079 gnd.n2078 0.152939
R13763 gnd.n2080 gnd.n2079 0.152939
R13764 gnd.n2081 gnd.n2080 0.152939
R13765 gnd.n2082 gnd.n2081 0.152939
R13766 gnd.n2083 gnd.n2082 0.152939
R13767 gnd.n2084 gnd.n2083 0.152939
R13768 gnd.n2085 gnd.n2084 0.152939
R13769 gnd.n2086 gnd.n2085 0.152939
R13770 gnd.n2086 gnd.n1254 0.152939
R13771 gnd.n2165 gnd.n1254 0.152939
R13772 gnd.n2166 gnd.n2165 0.152939
R13773 gnd.n2167 gnd.n2166 0.152939
R13774 gnd.n2168 gnd.n2167 0.152939
R13775 gnd.n2169 gnd.n2168 0.152939
R13776 gnd.n2170 gnd.n2169 0.152939
R13777 gnd.n2171 gnd.n2170 0.152939
R13778 gnd.n2173 gnd.n2171 0.152939
R13779 gnd.n2173 gnd.n2172 0.152939
R13780 gnd.n2172 gnd.n977 0.152939
R13781 gnd.n2226 gnd.n977 0.152939
R13782 gnd.n1749 gnd.n1748 0.152939
R13783 gnd.n1749 gnd.n1639 0.152939
R13784 gnd.n1764 gnd.n1639 0.152939
R13785 gnd.n1765 gnd.n1764 0.152939
R13786 gnd.n1766 gnd.n1765 0.152939
R13787 gnd.n1766 gnd.n1627 0.152939
R13788 gnd.n1780 gnd.n1627 0.152939
R13789 gnd.n1781 gnd.n1780 0.152939
R13790 gnd.n1782 gnd.n1781 0.152939
R13791 gnd.n1783 gnd.n1782 0.152939
R13792 gnd.n1784 gnd.n1783 0.152939
R13793 gnd.n1785 gnd.n1784 0.152939
R13794 gnd.n1786 gnd.n1785 0.152939
R13795 gnd.n1787 gnd.n1786 0.152939
R13796 gnd.n1788 gnd.n1787 0.152939
R13797 gnd.n1789 gnd.n1788 0.152939
R13798 gnd.n1790 gnd.n1789 0.152939
R13799 gnd.n1791 gnd.n1790 0.152939
R13800 gnd.n1792 gnd.n1791 0.152939
R13801 gnd.n1793 gnd.n1792 0.152939
R13802 gnd.n1794 gnd.n1793 0.152939
R13803 gnd.n1794 gnd.n1493 0.152939
R13804 gnd.n1911 gnd.n1493 0.152939
R13805 gnd.n1912 gnd.n1911 0.152939
R13806 gnd.n1913 gnd.n1912 0.152939
R13807 gnd.n1914 gnd.n1913 0.152939
R13808 gnd.n1914 gnd.n1415 0.152939
R13809 gnd.n1991 gnd.n1415 0.152939
R13810 gnd.n1667 gnd.n1666 0.152939
R13811 gnd.n1668 gnd.n1667 0.152939
R13812 gnd.n1669 gnd.n1668 0.152939
R13813 gnd.n1670 gnd.n1669 0.152939
R13814 gnd.n1671 gnd.n1670 0.152939
R13815 gnd.n1672 gnd.n1671 0.152939
R13816 gnd.n1673 gnd.n1672 0.152939
R13817 gnd.n1674 gnd.n1673 0.152939
R13818 gnd.n1675 gnd.n1674 0.152939
R13819 gnd.n1676 gnd.n1675 0.152939
R13820 gnd.n1677 gnd.n1676 0.152939
R13821 gnd.n1678 gnd.n1677 0.152939
R13822 gnd.n1679 gnd.n1678 0.152939
R13823 gnd.n1680 gnd.n1679 0.152939
R13824 gnd.n1681 gnd.n1680 0.152939
R13825 gnd.n1682 gnd.n1681 0.152939
R13826 gnd.n1683 gnd.n1682 0.152939
R13827 gnd.n1684 gnd.n1683 0.152939
R13828 gnd.n1685 gnd.n1684 0.152939
R13829 gnd.n1686 gnd.n1685 0.152939
R13830 gnd.n1687 gnd.n1686 0.152939
R13831 gnd.n1688 gnd.n1687 0.152939
R13832 gnd.n1692 gnd.n1688 0.152939
R13833 gnd.n1693 gnd.n1692 0.152939
R13834 gnd.n1693 gnd.n1650 0.152939
R13835 gnd.n1747 gnd.n1650 0.152939
R13836 gnd.n6327 gnd.n676 0.152939
R13837 gnd.n6328 gnd.n6327 0.152939
R13838 gnd.n6329 gnd.n6328 0.152939
R13839 gnd.n6329 gnd.n670 0.152939
R13840 gnd.n6337 gnd.n670 0.152939
R13841 gnd.n6338 gnd.n6337 0.152939
R13842 gnd.n6339 gnd.n6338 0.152939
R13843 gnd.n6339 gnd.n664 0.152939
R13844 gnd.n6347 gnd.n664 0.152939
R13845 gnd.n6348 gnd.n6347 0.152939
R13846 gnd.n6349 gnd.n6348 0.152939
R13847 gnd.n6349 gnd.n658 0.152939
R13848 gnd.n6357 gnd.n658 0.152939
R13849 gnd.n6358 gnd.n6357 0.152939
R13850 gnd.n6359 gnd.n6358 0.152939
R13851 gnd.n6359 gnd.n652 0.152939
R13852 gnd.n6367 gnd.n652 0.152939
R13853 gnd.n6368 gnd.n6367 0.152939
R13854 gnd.n6369 gnd.n6368 0.152939
R13855 gnd.n6369 gnd.n646 0.152939
R13856 gnd.n6377 gnd.n646 0.152939
R13857 gnd.n6378 gnd.n6377 0.152939
R13858 gnd.n6379 gnd.n6378 0.152939
R13859 gnd.n6379 gnd.n640 0.152939
R13860 gnd.n6387 gnd.n640 0.152939
R13861 gnd.n6388 gnd.n6387 0.152939
R13862 gnd.n6389 gnd.n6388 0.152939
R13863 gnd.n6389 gnd.n634 0.152939
R13864 gnd.n6397 gnd.n634 0.152939
R13865 gnd.n6398 gnd.n6397 0.152939
R13866 gnd.n6399 gnd.n6398 0.152939
R13867 gnd.n6399 gnd.n628 0.152939
R13868 gnd.n6407 gnd.n628 0.152939
R13869 gnd.n6408 gnd.n6407 0.152939
R13870 gnd.n6409 gnd.n6408 0.152939
R13871 gnd.n6409 gnd.n622 0.152939
R13872 gnd.n6417 gnd.n622 0.152939
R13873 gnd.n6418 gnd.n6417 0.152939
R13874 gnd.n6419 gnd.n6418 0.152939
R13875 gnd.n6419 gnd.n616 0.152939
R13876 gnd.n6427 gnd.n616 0.152939
R13877 gnd.n6428 gnd.n6427 0.152939
R13878 gnd.n6429 gnd.n6428 0.152939
R13879 gnd.n6429 gnd.n610 0.152939
R13880 gnd.n6437 gnd.n610 0.152939
R13881 gnd.n6438 gnd.n6437 0.152939
R13882 gnd.n6439 gnd.n6438 0.152939
R13883 gnd.n6439 gnd.n604 0.152939
R13884 gnd.n6447 gnd.n604 0.152939
R13885 gnd.n6448 gnd.n6447 0.152939
R13886 gnd.n6449 gnd.n6448 0.152939
R13887 gnd.n6449 gnd.n598 0.152939
R13888 gnd.n6457 gnd.n598 0.152939
R13889 gnd.n6458 gnd.n6457 0.152939
R13890 gnd.n6459 gnd.n6458 0.152939
R13891 gnd.n6459 gnd.n592 0.152939
R13892 gnd.n6467 gnd.n592 0.152939
R13893 gnd.n6468 gnd.n6467 0.152939
R13894 gnd.n6469 gnd.n6468 0.152939
R13895 gnd.n6469 gnd.n586 0.152939
R13896 gnd.n6477 gnd.n586 0.152939
R13897 gnd.n6478 gnd.n6477 0.152939
R13898 gnd.n6479 gnd.n6478 0.152939
R13899 gnd.n6479 gnd.n580 0.152939
R13900 gnd.n6487 gnd.n580 0.152939
R13901 gnd.n6488 gnd.n6487 0.152939
R13902 gnd.n6489 gnd.n6488 0.152939
R13903 gnd.n6489 gnd.n574 0.152939
R13904 gnd.n6497 gnd.n574 0.152939
R13905 gnd.n6498 gnd.n6497 0.152939
R13906 gnd.n6499 gnd.n6498 0.152939
R13907 gnd.n6499 gnd.n568 0.152939
R13908 gnd.n6507 gnd.n568 0.152939
R13909 gnd.n6508 gnd.n6507 0.152939
R13910 gnd.n6509 gnd.n6508 0.152939
R13911 gnd.n6509 gnd.n562 0.152939
R13912 gnd.n6517 gnd.n562 0.152939
R13913 gnd.n6518 gnd.n6517 0.152939
R13914 gnd.n6519 gnd.n6518 0.152939
R13915 gnd.n6519 gnd.n556 0.152939
R13916 gnd.n6527 gnd.n556 0.152939
R13917 gnd.n6528 gnd.n6527 0.152939
R13918 gnd.n6529 gnd.n6528 0.152939
R13919 gnd.n6529 gnd.n550 0.152939
R13920 gnd.n6537 gnd.n550 0.152939
R13921 gnd.n6538 gnd.n6537 0.152939
R13922 gnd.n6539 gnd.n6538 0.152939
R13923 gnd.n6539 gnd.n544 0.152939
R13924 gnd.n6547 gnd.n544 0.152939
R13925 gnd.n6548 gnd.n6547 0.152939
R13926 gnd.n6549 gnd.n6548 0.152939
R13927 gnd.n6549 gnd.n538 0.152939
R13928 gnd.n6557 gnd.n538 0.152939
R13929 gnd.n6558 gnd.n6557 0.152939
R13930 gnd.n6559 gnd.n6558 0.152939
R13931 gnd.n6559 gnd.n532 0.152939
R13932 gnd.n6567 gnd.n532 0.152939
R13933 gnd.n6568 gnd.n6567 0.152939
R13934 gnd.n6569 gnd.n6568 0.152939
R13935 gnd.n6569 gnd.n526 0.152939
R13936 gnd.n6577 gnd.n526 0.152939
R13937 gnd.n6578 gnd.n6577 0.152939
R13938 gnd.n6579 gnd.n6578 0.152939
R13939 gnd.n6579 gnd.n520 0.152939
R13940 gnd.n6587 gnd.n520 0.152939
R13941 gnd.n6588 gnd.n6587 0.152939
R13942 gnd.n6589 gnd.n6588 0.152939
R13943 gnd.n6589 gnd.n514 0.152939
R13944 gnd.n6597 gnd.n514 0.152939
R13945 gnd.n6598 gnd.n6597 0.152939
R13946 gnd.n6599 gnd.n6598 0.152939
R13947 gnd.n6599 gnd.n508 0.152939
R13948 gnd.n6607 gnd.n508 0.152939
R13949 gnd.n6608 gnd.n6607 0.152939
R13950 gnd.n6609 gnd.n6608 0.152939
R13951 gnd.n6609 gnd.n502 0.152939
R13952 gnd.n6617 gnd.n502 0.152939
R13953 gnd.n6618 gnd.n6617 0.152939
R13954 gnd.n6619 gnd.n6618 0.152939
R13955 gnd.n6619 gnd.n496 0.152939
R13956 gnd.n6627 gnd.n496 0.152939
R13957 gnd.n6628 gnd.n6627 0.152939
R13958 gnd.n6629 gnd.n6628 0.152939
R13959 gnd.n6629 gnd.n490 0.152939
R13960 gnd.n6637 gnd.n490 0.152939
R13961 gnd.n6638 gnd.n6637 0.152939
R13962 gnd.n6639 gnd.n6638 0.152939
R13963 gnd.n6639 gnd.n484 0.152939
R13964 gnd.n6647 gnd.n484 0.152939
R13965 gnd.n6648 gnd.n6647 0.152939
R13966 gnd.n6649 gnd.n6648 0.152939
R13967 gnd.n6649 gnd.n478 0.152939
R13968 gnd.n6657 gnd.n478 0.152939
R13969 gnd.n6658 gnd.n6657 0.152939
R13970 gnd.n6659 gnd.n6658 0.152939
R13971 gnd.n6659 gnd.n472 0.152939
R13972 gnd.n6667 gnd.n472 0.152939
R13973 gnd.n6668 gnd.n6667 0.152939
R13974 gnd.n6669 gnd.n6668 0.152939
R13975 gnd.n6669 gnd.n466 0.152939
R13976 gnd.n6677 gnd.n466 0.152939
R13977 gnd.n6678 gnd.n6677 0.152939
R13978 gnd.n6679 gnd.n6678 0.152939
R13979 gnd.n6679 gnd.n460 0.152939
R13980 gnd.n6687 gnd.n460 0.152939
R13981 gnd.n6688 gnd.n6687 0.152939
R13982 gnd.n6689 gnd.n6688 0.152939
R13983 gnd.n6689 gnd.n454 0.152939
R13984 gnd.n6697 gnd.n454 0.152939
R13985 gnd.n6698 gnd.n6697 0.152939
R13986 gnd.n6700 gnd.n6698 0.152939
R13987 gnd.n6700 gnd.n6699 0.152939
R13988 gnd.n6699 gnd.n448 0.152939
R13989 gnd.n6709 gnd.n448 0.152939
R13990 gnd.n6710 gnd.n443 0.152939
R13991 gnd.n6718 gnd.n443 0.152939
R13992 gnd.n6719 gnd.n6718 0.152939
R13993 gnd.n6720 gnd.n6719 0.152939
R13994 gnd.n6720 gnd.n437 0.152939
R13995 gnd.n6728 gnd.n437 0.152939
R13996 gnd.n6729 gnd.n6728 0.152939
R13997 gnd.n6730 gnd.n6729 0.152939
R13998 gnd.n6730 gnd.n431 0.152939
R13999 gnd.n6738 gnd.n431 0.152939
R14000 gnd.n6739 gnd.n6738 0.152939
R14001 gnd.n6740 gnd.n6739 0.152939
R14002 gnd.n6740 gnd.n425 0.152939
R14003 gnd.n6748 gnd.n425 0.152939
R14004 gnd.n6749 gnd.n6748 0.152939
R14005 gnd.n6750 gnd.n6749 0.152939
R14006 gnd.n6750 gnd.n419 0.152939
R14007 gnd.n6758 gnd.n419 0.152939
R14008 gnd.n6759 gnd.n6758 0.152939
R14009 gnd.n6760 gnd.n6759 0.152939
R14010 gnd.n6760 gnd.n413 0.152939
R14011 gnd.n6768 gnd.n413 0.152939
R14012 gnd.n6769 gnd.n6768 0.152939
R14013 gnd.n6770 gnd.n6769 0.152939
R14014 gnd.n6770 gnd.n407 0.152939
R14015 gnd.n6778 gnd.n407 0.152939
R14016 gnd.n6779 gnd.n6778 0.152939
R14017 gnd.n6780 gnd.n6779 0.152939
R14018 gnd.n6780 gnd.n401 0.152939
R14019 gnd.n6788 gnd.n401 0.152939
R14020 gnd.n6789 gnd.n6788 0.152939
R14021 gnd.n6790 gnd.n6789 0.152939
R14022 gnd.n6790 gnd.n395 0.152939
R14023 gnd.n6798 gnd.n395 0.152939
R14024 gnd.n6799 gnd.n6798 0.152939
R14025 gnd.n6800 gnd.n6799 0.152939
R14026 gnd.n6800 gnd.n389 0.152939
R14027 gnd.n6808 gnd.n389 0.152939
R14028 gnd.n6809 gnd.n6808 0.152939
R14029 gnd.n6810 gnd.n6809 0.152939
R14030 gnd.n6810 gnd.n383 0.152939
R14031 gnd.n6818 gnd.n383 0.152939
R14032 gnd.n6819 gnd.n6818 0.152939
R14033 gnd.n6820 gnd.n6819 0.152939
R14034 gnd.n6820 gnd.n377 0.152939
R14035 gnd.n6828 gnd.n377 0.152939
R14036 gnd.n6829 gnd.n6828 0.152939
R14037 gnd.n6830 gnd.n6829 0.152939
R14038 gnd.n6830 gnd.n371 0.152939
R14039 gnd.n6838 gnd.n371 0.152939
R14040 gnd.n6839 gnd.n6838 0.152939
R14041 gnd.n6840 gnd.n6839 0.152939
R14042 gnd.n6840 gnd.n365 0.152939
R14043 gnd.n6848 gnd.n365 0.152939
R14044 gnd.n6849 gnd.n6848 0.152939
R14045 gnd.n6850 gnd.n6849 0.152939
R14046 gnd.n6850 gnd.n359 0.152939
R14047 gnd.n6858 gnd.n359 0.152939
R14048 gnd.n6859 gnd.n6858 0.152939
R14049 gnd.n6860 gnd.n6859 0.152939
R14050 gnd.n6860 gnd.n353 0.152939
R14051 gnd.n6868 gnd.n353 0.152939
R14052 gnd.n6869 gnd.n6868 0.152939
R14053 gnd.n6870 gnd.n6869 0.152939
R14054 gnd.n6870 gnd.n347 0.152939
R14055 gnd.n6878 gnd.n347 0.152939
R14056 gnd.n6879 gnd.n6878 0.152939
R14057 gnd.n6880 gnd.n6879 0.152939
R14058 gnd.n6880 gnd.n341 0.152939
R14059 gnd.n6888 gnd.n341 0.152939
R14060 gnd.n6889 gnd.n6888 0.152939
R14061 gnd.n6890 gnd.n6889 0.152939
R14062 gnd.n6890 gnd.n335 0.152939
R14063 gnd.n6898 gnd.n335 0.152939
R14064 gnd.n6899 gnd.n6898 0.152939
R14065 gnd.n6900 gnd.n6899 0.152939
R14066 gnd.n6900 gnd.n329 0.152939
R14067 gnd.n6908 gnd.n329 0.152939
R14068 gnd.n6909 gnd.n6908 0.152939
R14069 gnd.n6910 gnd.n6909 0.152939
R14070 gnd.n6910 gnd.n323 0.152939
R14071 gnd.n6919 gnd.n323 0.152939
R14072 gnd.n6920 gnd.n6919 0.152939
R14073 gnd.n6921 gnd.n6920 0.152939
R14074 gnd.n7056 gnd.n248 0.152939
R14075 gnd.n7057 gnd.n7056 0.152939
R14076 gnd.n7058 gnd.n7057 0.152939
R14077 gnd.n7058 gnd.n231 0.152939
R14078 gnd.n7072 gnd.n231 0.152939
R14079 gnd.n7073 gnd.n7072 0.152939
R14080 gnd.n7074 gnd.n7073 0.152939
R14081 gnd.n7074 gnd.n218 0.152939
R14082 gnd.n7088 gnd.n218 0.152939
R14083 gnd.n7089 gnd.n7088 0.152939
R14084 gnd.n7090 gnd.n7089 0.152939
R14085 gnd.n7090 gnd.n201 0.152939
R14086 gnd.n7104 gnd.n201 0.152939
R14087 gnd.n7105 gnd.n7104 0.152939
R14088 gnd.n7106 gnd.n7105 0.152939
R14089 gnd.n7106 gnd.n185 0.152939
R14090 gnd.n7195 gnd.n185 0.152939
R14091 gnd.n7196 gnd.n7195 0.152939
R14092 gnd.n7197 gnd.n7196 0.152939
R14093 gnd.n7197 gnd.n107 0.152939
R14094 gnd.n7277 gnd.n107 0.152939
R14095 gnd.n7276 gnd.n108 0.152939
R14096 gnd.n110 gnd.n108 0.152939
R14097 gnd.n114 gnd.n110 0.152939
R14098 gnd.n115 gnd.n114 0.152939
R14099 gnd.n116 gnd.n115 0.152939
R14100 gnd.n117 gnd.n116 0.152939
R14101 gnd.n121 gnd.n117 0.152939
R14102 gnd.n122 gnd.n121 0.152939
R14103 gnd.n123 gnd.n122 0.152939
R14104 gnd.n124 gnd.n123 0.152939
R14105 gnd.n128 gnd.n124 0.152939
R14106 gnd.n129 gnd.n128 0.152939
R14107 gnd.n130 gnd.n129 0.152939
R14108 gnd.n131 gnd.n130 0.152939
R14109 gnd.n135 gnd.n131 0.152939
R14110 gnd.n136 gnd.n135 0.152939
R14111 gnd.n137 gnd.n136 0.152939
R14112 gnd.n138 gnd.n137 0.152939
R14113 gnd.n142 gnd.n138 0.152939
R14114 gnd.n143 gnd.n142 0.152939
R14115 gnd.n144 gnd.n143 0.152939
R14116 gnd.n145 gnd.n144 0.152939
R14117 gnd.n149 gnd.n145 0.152939
R14118 gnd.n150 gnd.n149 0.152939
R14119 gnd.n151 gnd.n150 0.152939
R14120 gnd.n152 gnd.n151 0.152939
R14121 gnd.n156 gnd.n152 0.152939
R14122 gnd.n157 gnd.n156 0.152939
R14123 gnd.n158 gnd.n157 0.152939
R14124 gnd.n159 gnd.n158 0.152939
R14125 gnd.n163 gnd.n159 0.152939
R14126 gnd.n164 gnd.n163 0.152939
R14127 gnd.n165 gnd.n164 0.152939
R14128 gnd.n166 gnd.n165 0.152939
R14129 gnd.n170 gnd.n166 0.152939
R14130 gnd.n171 gnd.n170 0.152939
R14131 gnd.n7207 gnd.n171 0.152939
R14132 gnd.n7207 gnd.n7206 0.152939
R14133 gnd.n2925 gnd.n2769 0.152939
R14134 gnd.n2926 gnd.n2925 0.152939
R14135 gnd.n2927 gnd.n2926 0.152939
R14136 gnd.n2928 gnd.n2927 0.152939
R14137 gnd.n2929 gnd.n2928 0.152939
R14138 gnd.n2930 gnd.n2929 0.152939
R14139 gnd.n2931 gnd.n2930 0.152939
R14140 gnd.n2932 gnd.n2931 0.152939
R14141 gnd.n2933 gnd.n2932 0.152939
R14142 gnd.n2934 gnd.n2933 0.152939
R14143 gnd.n2935 gnd.n2934 0.152939
R14144 gnd.n2936 gnd.n2935 0.152939
R14145 gnd.n2937 gnd.n2936 0.152939
R14146 gnd.n2937 gnd.n2832 0.152939
R14147 gnd.n5528 gnd.n2832 0.152939
R14148 gnd.n5529 gnd.n5528 0.152939
R14149 gnd.n5530 gnd.n5529 0.152939
R14150 gnd.n5530 gnd.n2830 0.152939
R14151 gnd.n5535 gnd.n2830 0.152939
R14152 gnd.n5536 gnd.n5535 0.152939
R14153 gnd.n5537 gnd.n5536 0.152939
R14154 gnd.n5538 gnd.n5537 0.152939
R14155 gnd.n5539 gnd.n5538 0.152939
R14156 gnd.n5541 gnd.n5539 0.152939
R14157 gnd.n5541 gnd.n5540 0.152939
R14158 gnd.n5540 gnd.n295 0.152939
R14159 gnd.n6957 gnd.n6956 0.152939
R14160 gnd.n6958 gnd.n6957 0.152939
R14161 gnd.n6959 gnd.n6958 0.152939
R14162 gnd.n6960 gnd.n6959 0.152939
R14163 gnd.n6961 gnd.n6960 0.152939
R14164 gnd.n6962 gnd.n6961 0.152939
R14165 gnd.n6963 gnd.n6962 0.152939
R14166 gnd.n6964 gnd.n6963 0.152939
R14167 gnd.n6965 gnd.n6964 0.152939
R14168 gnd.n6966 gnd.n6965 0.152939
R14169 gnd.n6967 gnd.n6966 0.152939
R14170 gnd.n6968 gnd.n6967 0.152939
R14171 gnd.n6969 gnd.n6968 0.152939
R14172 gnd.n6970 gnd.n6969 0.152939
R14173 gnd.n6971 gnd.n6970 0.152939
R14174 gnd.n6972 gnd.n6971 0.152939
R14175 gnd.n6973 gnd.n6972 0.152939
R14176 gnd.n6974 gnd.n6973 0.152939
R14177 gnd.n6975 gnd.n6974 0.152939
R14178 gnd.n6976 gnd.n6975 0.152939
R14179 gnd.n6977 gnd.n6976 0.152939
R14180 gnd.n6978 gnd.n6977 0.152939
R14181 gnd.n6980 gnd.n6978 0.152939
R14182 gnd.n6980 gnd.n6979 0.152939
R14183 gnd.n6979 gnd.n177 0.152939
R14184 gnd.n7205 gnd.n177 0.152939
R14185 gnd.n2726 gnd.n2725 0.152939
R14186 gnd.n2727 gnd.n2726 0.152939
R14187 gnd.n2728 gnd.n2727 0.152939
R14188 gnd.n2729 gnd.n2728 0.152939
R14189 gnd.n2730 gnd.n2729 0.152939
R14190 gnd.n2731 gnd.n2730 0.152939
R14191 gnd.n2732 gnd.n2731 0.152939
R14192 gnd.n2733 gnd.n2732 0.152939
R14193 gnd.n2734 gnd.n2733 0.152939
R14194 gnd.n2735 gnd.n2734 0.152939
R14195 gnd.n2736 gnd.n2735 0.152939
R14196 gnd.n2737 gnd.n2736 0.152939
R14197 gnd.n2738 gnd.n2737 0.152939
R14198 gnd.n2739 gnd.n2738 0.152939
R14199 gnd.n2740 gnd.n2739 0.152939
R14200 gnd.n2747 gnd.n2746 0.152939
R14201 gnd.n2748 gnd.n2747 0.152939
R14202 gnd.n2749 gnd.n2748 0.152939
R14203 gnd.n2750 gnd.n2749 0.152939
R14204 gnd.n2751 gnd.n2750 0.152939
R14205 gnd.n2752 gnd.n2751 0.152939
R14206 gnd.n2753 gnd.n2752 0.152939
R14207 gnd.n2754 gnd.n2753 0.152939
R14208 gnd.n2755 gnd.n2754 0.152939
R14209 gnd.n2756 gnd.n2755 0.152939
R14210 gnd.n2757 gnd.n2756 0.152939
R14211 gnd.n2758 gnd.n2757 0.152939
R14212 gnd.n2759 gnd.n2758 0.152939
R14213 gnd.n2760 gnd.n2759 0.152939
R14214 gnd.n2761 gnd.n2760 0.152939
R14215 gnd.n2762 gnd.n2761 0.152939
R14216 gnd.n2763 gnd.n2762 0.152939
R14217 gnd.n5628 gnd.n2763 0.152939
R14218 gnd.n5628 gnd.n5627 0.152939
R14219 gnd.n5627 gnd.n5626 0.152939
R14220 gnd.n2920 gnd.n2919 0.152939
R14221 gnd.n2920 gnd.n2898 0.152939
R14222 gnd.n5450 gnd.n2898 0.152939
R14223 gnd.n5451 gnd.n5450 0.152939
R14224 gnd.n5452 gnd.n5451 0.152939
R14225 gnd.n5453 gnd.n5452 0.152939
R14226 gnd.n5453 gnd.n2869 0.152939
R14227 gnd.n5481 gnd.n2869 0.152939
R14228 gnd.n5482 gnd.n5481 0.152939
R14229 gnd.n5483 gnd.n5482 0.152939
R14230 gnd.n5484 gnd.n5483 0.152939
R14231 gnd.n5484 gnd.n2841 0.152939
R14232 gnd.n5518 gnd.n2841 0.152939
R14233 gnd.n5519 gnd.n5518 0.152939
R14234 gnd.n5520 gnd.n5519 0.152939
R14235 gnd.n5521 gnd.n5520 0.152939
R14236 gnd.n5521 gnd.n2807 0.152939
R14237 gnd.n5582 gnd.n2807 0.152939
R14238 gnd.n5583 gnd.n5582 0.152939
R14239 gnd.n5584 gnd.n5583 0.152939
R14240 gnd.n5584 gnd.n262 0.152939
R14241 gnd.n5570 gnd.n5569 0.152939
R14242 gnd.n5569 gnd.n312 0.152939
R14243 gnd.n313 gnd.n312 0.152939
R14244 gnd.n314 gnd.n313 0.152939
R14245 gnd.n315 gnd.n314 0.152939
R14246 gnd.n319 gnd.n318 0.152939
R14247 gnd.n320 gnd.n319 0.152939
R14248 gnd.n3701 gnd.n3700 0.152939
R14249 gnd.n3704 gnd.n3701 0.152939
R14250 gnd.n3705 gnd.n3704 0.152939
R14251 gnd.n3706 gnd.n3705 0.152939
R14252 gnd.n3707 gnd.n3706 0.152939
R14253 gnd.n3710 gnd.n3707 0.152939
R14254 gnd.n3711 gnd.n3710 0.152939
R14255 gnd.n3712 gnd.n3711 0.152939
R14256 gnd.n3713 gnd.n3712 0.152939
R14257 gnd.n3716 gnd.n3713 0.152939
R14258 gnd.n3717 gnd.n3716 0.152939
R14259 gnd.n3718 gnd.n3717 0.152939
R14260 gnd.n3719 gnd.n3718 0.152939
R14261 gnd.n3722 gnd.n3719 0.152939
R14262 gnd.n3723 gnd.n3722 0.152939
R14263 gnd.n3724 gnd.n3723 0.152939
R14264 gnd.n3725 gnd.n3724 0.152939
R14265 gnd.n3728 gnd.n3725 0.152939
R14266 gnd.n3729 gnd.n3728 0.152939
R14267 gnd.n3730 gnd.n3729 0.152939
R14268 gnd.n3731 gnd.n3730 0.152939
R14269 gnd.n3734 gnd.n3731 0.152939
R14270 gnd.n3735 gnd.n3734 0.152939
R14271 gnd.n3736 gnd.n3735 0.152939
R14272 gnd.n3737 gnd.n3736 0.152939
R14273 gnd.n3737 gnd.n3436 0.152939
R14274 gnd.n4418 gnd.n3436 0.152939
R14275 gnd.n4419 gnd.n4418 0.152939
R14276 gnd.n4420 gnd.n4419 0.152939
R14277 gnd.n4420 gnd.n3422 0.152939
R14278 gnd.n4434 gnd.n3422 0.152939
R14279 gnd.n4435 gnd.n4434 0.152939
R14280 gnd.n4436 gnd.n4435 0.152939
R14281 gnd.n4437 gnd.n4436 0.152939
R14282 gnd.n4437 gnd.n3390 0.152939
R14283 gnd.n4558 gnd.n3390 0.152939
R14284 gnd.n4559 gnd.n4558 0.152939
R14285 gnd.n4560 gnd.n4559 0.152939
R14286 gnd.n4560 gnd.n3376 0.152939
R14287 gnd.n4574 gnd.n3376 0.152939
R14288 gnd.n4575 gnd.n4574 0.152939
R14289 gnd.n4576 gnd.n4575 0.152939
R14290 gnd.n4576 gnd.n3361 0.152939
R14291 gnd.n4590 gnd.n3361 0.152939
R14292 gnd.n4591 gnd.n4590 0.152939
R14293 gnd.n4592 gnd.n4591 0.152939
R14294 gnd.n4592 gnd.n3347 0.152939
R14295 gnd.n4605 gnd.n3347 0.152939
R14296 gnd.n4606 gnd.n4605 0.152939
R14297 gnd.n4607 gnd.n4606 0.152939
R14298 gnd.n4608 gnd.n4607 0.152939
R14299 gnd.n4608 gnd.n3315 0.152939
R14300 gnd.n4731 gnd.n3315 0.152939
R14301 gnd.n4732 gnd.n4731 0.152939
R14302 gnd.n4733 gnd.n4732 0.152939
R14303 gnd.n4733 gnd.n3301 0.152939
R14304 gnd.n4747 gnd.n3301 0.152939
R14305 gnd.n4748 gnd.n4747 0.152939
R14306 gnd.n4749 gnd.n4748 0.152939
R14307 gnd.n4749 gnd.n3288 0.152939
R14308 gnd.n4763 gnd.n3288 0.152939
R14309 gnd.n4764 gnd.n4763 0.152939
R14310 gnd.n4765 gnd.n4764 0.152939
R14311 gnd.n4765 gnd.n3277 0.152939
R14312 gnd.n4779 gnd.n3277 0.152939
R14313 gnd.n4780 gnd.n4779 0.152939
R14314 gnd.n4781 gnd.n4780 0.152939
R14315 gnd.n4782 gnd.n4781 0.152939
R14316 gnd.n4782 gnd.n3244 0.152939
R14317 gnd.n4902 gnd.n3244 0.152939
R14318 gnd.n4903 gnd.n4902 0.152939
R14319 gnd.n4904 gnd.n4903 0.152939
R14320 gnd.n4904 gnd.n3229 0.152939
R14321 gnd.n4918 gnd.n3229 0.152939
R14322 gnd.n4919 gnd.n4918 0.152939
R14323 gnd.n4920 gnd.n4919 0.152939
R14324 gnd.n4920 gnd.n3214 0.152939
R14325 gnd.n4934 gnd.n3214 0.152939
R14326 gnd.n4935 gnd.n4934 0.152939
R14327 gnd.n4936 gnd.n4935 0.152939
R14328 gnd.n4936 gnd.n3201 0.152939
R14329 gnd.n4950 gnd.n3201 0.152939
R14330 gnd.n4951 gnd.n4950 0.152939
R14331 gnd.n4952 gnd.n4951 0.152939
R14332 gnd.n4953 gnd.n4952 0.152939
R14333 gnd.n4953 gnd.n3169 0.152939
R14334 gnd.n5308 gnd.n3169 0.152939
R14335 gnd.n5309 gnd.n5308 0.152939
R14336 gnd.n5310 gnd.n5309 0.152939
R14337 gnd.n5310 gnd.n3156 0.152939
R14338 gnd.n5324 gnd.n3156 0.152939
R14339 gnd.n5325 gnd.n5324 0.152939
R14340 gnd.n5326 gnd.n5325 0.152939
R14341 gnd.n5326 gnd.n3142 0.152939
R14342 gnd.n5340 gnd.n3142 0.152939
R14343 gnd.n5341 gnd.n5340 0.152939
R14344 gnd.n5342 gnd.n5341 0.152939
R14345 gnd.n5342 gnd.n3129 0.152939
R14346 gnd.n5356 gnd.n3129 0.152939
R14347 gnd.n5357 gnd.n5356 0.152939
R14348 gnd.n5358 gnd.n5357 0.152939
R14349 gnd.n5358 gnd.n3115 0.152939
R14350 gnd.n5372 gnd.n3115 0.152939
R14351 gnd.n5373 gnd.n5372 0.152939
R14352 gnd.n5374 gnd.n5373 0.152939
R14353 gnd.n5374 gnd.n3101 0.152939
R14354 gnd.n5390 gnd.n3101 0.152939
R14355 gnd.n5391 gnd.n5390 0.152939
R14356 gnd.n5392 gnd.n5391 0.152939
R14357 gnd.n5394 gnd.n5392 0.152939
R14358 gnd.n5394 gnd.n5393 0.152939
R14359 gnd.n5393 gnd.n2688 0.152939
R14360 gnd.n2689 gnd.n2688 0.152939
R14361 gnd.n2690 gnd.n2689 0.152939
R14362 gnd.n2912 gnd.n2690 0.152939
R14363 gnd.n2913 gnd.n2912 0.152939
R14364 gnd.n2914 gnd.n2913 0.152939
R14365 gnd.n2914 gnd.n2908 0.152939
R14366 gnd.n5439 gnd.n2908 0.152939
R14367 gnd.n5440 gnd.n5439 0.152939
R14368 gnd.n5441 gnd.n5440 0.152939
R14369 gnd.n5442 gnd.n5441 0.152939
R14370 gnd.n5442 gnd.n2880 0.152939
R14371 gnd.n5470 gnd.n2880 0.152939
R14372 gnd.n5471 gnd.n5470 0.152939
R14373 gnd.n5472 gnd.n5471 0.152939
R14374 gnd.n5473 gnd.n5472 0.152939
R14375 gnd.n5473 gnd.n2852 0.152939
R14376 gnd.n5506 gnd.n2852 0.152939
R14377 gnd.n5507 gnd.n5506 0.152939
R14378 gnd.n5508 gnd.n5507 0.152939
R14379 gnd.n5509 gnd.n5508 0.152939
R14380 gnd.n5509 gnd.n2818 0.152939
R14381 gnd.n5564 gnd.n2818 0.152939
R14382 gnd.n5565 gnd.n5564 0.152939
R14383 gnd.n5566 gnd.n5565 0.152939
R14384 gnd.n5567 gnd.n5566 0.152939
R14385 gnd.n5568 gnd.n5567 0.152939
R14386 gnd.n5570 gnd.n5568 0.152939
R14387 gnd.n2460 gnd.n2459 0.152939
R14388 gnd.n2478 gnd.n2460 0.152939
R14389 gnd.n2479 gnd.n2478 0.152939
R14390 gnd.n2480 gnd.n2479 0.152939
R14391 gnd.n2481 gnd.n2480 0.152939
R14392 gnd.n2500 gnd.n2481 0.152939
R14393 gnd.n2501 gnd.n2500 0.152939
R14394 gnd.n2502 gnd.n2501 0.152939
R14395 gnd.n2503 gnd.n2502 0.152939
R14396 gnd.n2521 gnd.n2503 0.152939
R14397 gnd.n2522 gnd.n2521 0.152939
R14398 gnd.n2523 gnd.n2522 0.152939
R14399 gnd.n2524 gnd.n2523 0.152939
R14400 gnd.n2543 gnd.n2524 0.152939
R14401 gnd.n2544 gnd.n2543 0.152939
R14402 gnd.n2545 gnd.n2544 0.152939
R14403 gnd.n2546 gnd.n2545 0.152939
R14404 gnd.n2564 gnd.n2546 0.152939
R14405 gnd.n2565 gnd.n2564 0.152939
R14406 gnd.n2566 gnd.n2565 0.152939
R14407 gnd.n2567 gnd.n2566 0.152939
R14408 gnd.n3596 gnd.n3595 0.152939
R14409 gnd.n3597 gnd.n3596 0.152939
R14410 gnd.n3598 gnd.n3597 0.152939
R14411 gnd.n3599 gnd.n3598 0.152939
R14412 gnd.n3600 gnd.n3599 0.152939
R14413 gnd.n3601 gnd.n3600 0.152939
R14414 gnd.n3602 gnd.n3601 0.152939
R14415 gnd.n3603 gnd.n3602 0.152939
R14416 gnd.n3604 gnd.n3603 0.152939
R14417 gnd.n3605 gnd.n3604 0.152939
R14418 gnd.n3606 gnd.n3605 0.152939
R14419 gnd.n3607 gnd.n3606 0.152939
R14420 gnd.n3608 gnd.n3607 0.152939
R14421 gnd.n3609 gnd.n3608 0.152939
R14422 gnd.n3610 gnd.n3609 0.152939
R14423 gnd.n4139 gnd.n4138 0.152939
R14424 gnd.n4138 gnd.n3615 0.152939
R14425 gnd.n3616 gnd.n3615 0.152939
R14426 gnd.n3617 gnd.n3616 0.152939
R14427 gnd.n3618 gnd.n3617 0.152939
R14428 gnd.n3619 gnd.n3618 0.152939
R14429 gnd.n3620 gnd.n3619 0.152939
R14430 gnd.n3621 gnd.n3620 0.152939
R14431 gnd.n3622 gnd.n3621 0.152939
R14432 gnd.n3623 gnd.n3622 0.152939
R14433 gnd.n3624 gnd.n3623 0.152939
R14434 gnd.n3625 gnd.n3624 0.152939
R14435 gnd.n3626 gnd.n3625 0.152939
R14436 gnd.n3627 gnd.n3626 0.152939
R14437 gnd.n3628 gnd.n3627 0.152939
R14438 gnd.n3629 gnd.n3628 0.152939
R14439 gnd.n3630 gnd.n3629 0.152939
R14440 gnd.n3631 gnd.n3630 0.152939
R14441 gnd.n4098 gnd.n3631 0.152939
R14442 gnd.n4098 gnd.n4097 0.152939
R14443 gnd.n3827 gnd.n3800 0.152939
R14444 gnd.n3885 gnd.n3800 0.152939
R14445 gnd.n3886 gnd.n3885 0.152939
R14446 gnd.n3887 gnd.n3886 0.152939
R14447 gnd.n3887 gnd.n3798 0.152939
R14448 gnd.n3893 gnd.n3798 0.152939
R14449 gnd.n3894 gnd.n3893 0.152939
R14450 gnd.n3895 gnd.n3894 0.152939
R14451 gnd.n3895 gnd.n3796 0.152939
R14452 gnd.n3901 gnd.n3796 0.152939
R14453 gnd.n3902 gnd.n3901 0.152939
R14454 gnd.n3903 gnd.n3902 0.152939
R14455 gnd.n3903 gnd.n3794 0.152939
R14456 gnd.n3909 gnd.n3794 0.152939
R14457 gnd.n3910 gnd.n3909 0.152939
R14458 gnd.n3911 gnd.n3910 0.152939
R14459 gnd.n3911 gnd.n3792 0.152939
R14460 gnd.n3917 gnd.n3792 0.152939
R14461 gnd.n3918 gnd.n3917 0.152939
R14462 gnd.n3919 gnd.n3918 0.152939
R14463 gnd.n3919 gnd.n3790 0.152939
R14464 gnd.n3971 gnd.n3790 0.152939
R14465 gnd.n3972 gnd.n3971 0.152939
R14466 gnd.n3973 gnd.n3972 0.152939
R14467 gnd.n3973 gnd.n3679 0.152939
R14468 gnd.n3989 gnd.n3679 0.152939
R14469 gnd.n3866 gnd.n3807 0.152939
R14470 gnd.n3808 gnd.n3807 0.152939
R14471 gnd.n3809 gnd.n3808 0.152939
R14472 gnd.n3810 gnd.n3809 0.152939
R14473 gnd.n3811 gnd.n3810 0.152939
R14474 gnd.n3812 gnd.n3811 0.152939
R14475 gnd.n3813 gnd.n3812 0.152939
R14476 gnd.n3814 gnd.n3813 0.152939
R14477 gnd.n3815 gnd.n3814 0.152939
R14478 gnd.n3816 gnd.n3815 0.152939
R14479 gnd.n3817 gnd.n3816 0.152939
R14480 gnd.n3818 gnd.n3817 0.152939
R14481 gnd.n3819 gnd.n3818 0.152939
R14482 gnd.n3820 gnd.n3819 0.152939
R14483 gnd.n3821 gnd.n3820 0.152939
R14484 gnd.n3831 gnd.n3821 0.152939
R14485 gnd.n3831 gnd.n3830 0.152939
R14486 gnd.n3830 gnd.n3829 0.152939
R14487 gnd.n3872 gnd.n3867 0.152939
R14488 gnd.n3872 gnd.n3871 0.152939
R14489 gnd.n3871 gnd.n3870 0.152939
R14490 gnd.n3870 gnd.n3868 0.152939
R14491 gnd.n3868 gnd.n2331 0.152939
R14492 gnd.n2332 gnd.n2331 0.152939
R14493 gnd.n2333 gnd.n2332 0.152939
R14494 gnd.n2349 gnd.n2333 0.152939
R14495 gnd.n2350 gnd.n2349 0.152939
R14496 gnd.n2351 gnd.n2350 0.152939
R14497 gnd.n2352 gnd.n2351 0.152939
R14498 gnd.n2370 gnd.n2352 0.152939
R14499 gnd.n2371 gnd.n2370 0.152939
R14500 gnd.n2372 gnd.n2371 0.152939
R14501 gnd.n2373 gnd.n2372 0.152939
R14502 gnd.n2389 gnd.n2373 0.152939
R14503 gnd.n2390 gnd.n2389 0.152939
R14504 gnd.n2391 gnd.n2390 0.152939
R14505 gnd.n2392 gnd.n2391 0.152939
R14506 gnd.n2410 gnd.n2392 0.152939
R14507 gnd.n2411 gnd.n2410 0.152939
R14508 gnd.n2412 gnd.n2411 0.152939
R14509 gnd.n2413 gnd.n2412 0.152939
R14510 gnd.n2428 gnd.n2413 0.152939
R14511 gnd.n2429 gnd.n2428 0.152939
R14512 gnd.n2430 gnd.n2429 0.152939
R14513 gnd.n2447 gnd.n2431 0.152939
R14514 gnd.n2448 gnd.n2447 0.152939
R14515 gnd.n2449 gnd.n2448 0.152939
R14516 gnd.n2450 gnd.n2449 0.152939
R14517 gnd.n2467 gnd.n2450 0.152939
R14518 gnd.n2468 gnd.n2467 0.152939
R14519 gnd.n2469 gnd.n2468 0.152939
R14520 gnd.n2470 gnd.n2469 0.152939
R14521 gnd.n2489 gnd.n2470 0.152939
R14522 gnd.n2490 gnd.n2489 0.152939
R14523 gnd.n2491 gnd.n2490 0.152939
R14524 gnd.n2492 gnd.n2491 0.152939
R14525 gnd.n2510 gnd.n2492 0.152939
R14526 gnd.n2511 gnd.n2510 0.152939
R14527 gnd.n2512 gnd.n2511 0.152939
R14528 gnd.n2513 gnd.n2512 0.152939
R14529 gnd.n2532 gnd.n2513 0.152939
R14530 gnd.n2533 gnd.n2532 0.152939
R14531 gnd.n2534 gnd.n2533 0.152939
R14532 gnd.n2535 gnd.n2534 0.152939
R14533 gnd.n2554 gnd.n2535 0.152939
R14534 gnd.n2555 gnd.n2554 0.152939
R14535 gnd.n2556 gnd.n2555 0.152939
R14536 gnd.n2557 gnd.n2556 0.152939
R14537 gnd.n2574 gnd.n2557 0.152939
R14538 gnd.n5835 gnd.n2574 0.152939
R14539 gnd.n5994 gnd.n2306 0.152939
R14540 gnd.n5994 gnd.n5993 0.152939
R14541 gnd.n5993 gnd.n5992 0.152939
R14542 gnd.n5992 gnd.n2309 0.152939
R14543 gnd.n3932 gnd.n2309 0.152939
R14544 gnd.n3933 gnd.n3932 0.152939
R14545 gnd.n3933 gnd.n3930 0.152939
R14546 gnd.n3939 gnd.n3930 0.152939
R14547 gnd.n3940 gnd.n3939 0.152939
R14548 gnd.n3941 gnd.n3940 0.152939
R14549 gnd.n3941 gnd.n3928 0.152939
R14550 gnd.n3947 gnd.n3928 0.152939
R14551 gnd.n3948 gnd.n3947 0.152939
R14552 gnd.n3949 gnd.n3948 0.152939
R14553 gnd.n3949 gnd.n3926 0.152939
R14554 gnd.n3955 gnd.n3926 0.152939
R14555 gnd.n3956 gnd.n3955 0.152939
R14556 gnd.n3957 gnd.n3956 0.152939
R14557 gnd.n3957 gnd.n3924 0.152939
R14558 gnd.n3963 gnd.n3924 0.152939
R14559 gnd.n3964 gnd.n3963 0.152939
R14560 gnd.n3965 gnd.n3964 0.152939
R14561 gnd.n3965 gnd.n3787 0.152939
R14562 gnd.n3979 gnd.n3787 0.152939
R14563 gnd.n3980 gnd.n3979 0.152939
R14564 gnd.n3983 gnd.n3980 0.152939
R14565 gnd.n3998 gnd.n3676 0.152939
R14566 gnd.n3999 gnd.n3998 0.152939
R14567 gnd.n4000 gnd.n3999 0.152939
R14568 gnd.n4000 gnd.n3670 0.152939
R14569 gnd.n4014 gnd.n3670 0.152939
R14570 gnd.n4015 gnd.n4014 0.152939
R14571 gnd.n4016 gnd.n4015 0.152939
R14572 gnd.n4016 gnd.n3663 0.152939
R14573 gnd.n4030 gnd.n3663 0.152939
R14574 gnd.n4031 gnd.n4030 0.152939
R14575 gnd.n4032 gnd.n4031 0.152939
R14576 gnd.n4032 gnd.n3657 0.152939
R14577 gnd.n4046 gnd.n3657 0.152939
R14578 gnd.n4047 gnd.n4046 0.152939
R14579 gnd.n4048 gnd.n4047 0.152939
R14580 gnd.n4048 gnd.n3650 0.152939
R14581 gnd.n4062 gnd.n3650 0.152939
R14582 gnd.n4063 gnd.n4062 0.152939
R14583 gnd.n4064 gnd.n4063 0.152939
R14584 gnd.n4064 gnd.n3644 0.152939
R14585 gnd.n4078 gnd.n3644 0.152939
R14586 gnd.n4079 gnd.n4078 0.152939
R14587 gnd.n4081 gnd.n4079 0.152939
R14588 gnd.n4081 gnd.n4080 0.152939
R14589 gnd.n4080 gnd.n3636 0.152939
R14590 gnd.n4096 gnd.n3636 0.152939
R14591 gnd.n2264 gnd.n2263 0.152939
R14592 gnd.n2265 gnd.n2264 0.152939
R14593 gnd.n2266 gnd.n2265 0.152939
R14594 gnd.n2267 gnd.n2266 0.152939
R14595 gnd.n2268 gnd.n2267 0.152939
R14596 gnd.n2269 gnd.n2268 0.152939
R14597 gnd.n2270 gnd.n2269 0.152939
R14598 gnd.n2271 gnd.n2270 0.152939
R14599 gnd.n2272 gnd.n2271 0.152939
R14600 gnd.n2273 gnd.n2272 0.152939
R14601 gnd.n2274 gnd.n2273 0.152939
R14602 gnd.n2275 gnd.n2274 0.152939
R14603 gnd.n2276 gnd.n2275 0.152939
R14604 gnd.n2277 gnd.n2276 0.152939
R14605 gnd.n2278 gnd.n2277 0.152939
R14606 gnd.n2279 gnd.n2278 0.152939
R14607 gnd.n2280 gnd.n2279 0.152939
R14608 gnd.n2283 gnd.n2280 0.152939
R14609 gnd.n2284 gnd.n2283 0.152939
R14610 gnd.n2285 gnd.n2284 0.152939
R14611 gnd.n2286 gnd.n2285 0.152939
R14612 gnd.n2287 gnd.n2286 0.152939
R14613 gnd.n2288 gnd.n2287 0.152939
R14614 gnd.n2289 gnd.n2288 0.152939
R14615 gnd.n2290 gnd.n2289 0.152939
R14616 gnd.n2291 gnd.n2290 0.152939
R14617 gnd.n2292 gnd.n2291 0.152939
R14618 gnd.n2293 gnd.n2292 0.152939
R14619 gnd.n2294 gnd.n2293 0.152939
R14620 gnd.n2295 gnd.n2294 0.152939
R14621 gnd.n2296 gnd.n2295 0.152939
R14622 gnd.n2297 gnd.n2296 0.152939
R14623 gnd.n2298 gnd.n2297 0.152939
R14624 gnd.n2299 gnd.n2298 0.152939
R14625 gnd.n2300 gnd.n2299 0.152939
R14626 gnd.n6002 gnd.n2300 0.152939
R14627 gnd.n6002 gnd.n6001 0.152939
R14628 gnd.n6001 gnd.n6000 0.152939
R14629 gnd.n3878 gnd.n3876 0.152939
R14630 gnd.n3878 gnd.n3877 0.152939
R14631 gnd.n3877 gnd.n2320 0.152939
R14632 gnd.n2321 gnd.n2320 0.152939
R14633 gnd.n2322 gnd.n2321 0.152939
R14634 gnd.n2340 gnd.n2322 0.152939
R14635 gnd.n2341 gnd.n2340 0.152939
R14636 gnd.n2342 gnd.n2341 0.152939
R14637 gnd.n2343 gnd.n2342 0.152939
R14638 gnd.n2359 gnd.n2343 0.152939
R14639 gnd.n2360 gnd.n2359 0.152939
R14640 gnd.n2361 gnd.n2360 0.152939
R14641 gnd.n2362 gnd.n2361 0.152939
R14642 gnd.n2380 gnd.n2362 0.152939
R14643 gnd.n2381 gnd.n2380 0.152939
R14644 gnd.n2382 gnd.n2381 0.152939
R14645 gnd.n2383 gnd.n2382 0.152939
R14646 gnd.n2399 gnd.n2383 0.152939
R14647 gnd.n2400 gnd.n2399 0.152939
R14648 gnd.n2401 gnd.n2400 0.152939
R14649 gnd.n2402 gnd.n2401 0.152939
R14650 gnd.n3691 gnd.n3690 0.152939
R14651 gnd.n3692 gnd.n3691 0.152939
R14652 gnd.n3695 gnd.n3694 0.152939
R14653 gnd.n3698 gnd.n3695 0.152939
R14654 gnd.n3699 gnd.n3698 0.152939
R14655 gnd.n3700 gnd.n3699 0.152939
R14656 gnd.n682 gnd.n681 0.152939
R14657 gnd.n683 gnd.n682 0.152939
R14658 gnd.n688 gnd.n683 0.152939
R14659 gnd.n689 gnd.n688 0.152939
R14660 gnd.n690 gnd.n689 0.152939
R14661 gnd.n691 gnd.n690 0.152939
R14662 gnd.n696 gnd.n691 0.152939
R14663 gnd.n697 gnd.n696 0.152939
R14664 gnd.n698 gnd.n697 0.152939
R14665 gnd.n699 gnd.n698 0.152939
R14666 gnd.n704 gnd.n699 0.152939
R14667 gnd.n705 gnd.n704 0.152939
R14668 gnd.n706 gnd.n705 0.152939
R14669 gnd.n707 gnd.n706 0.152939
R14670 gnd.n712 gnd.n707 0.152939
R14671 gnd.n713 gnd.n712 0.152939
R14672 gnd.n714 gnd.n713 0.152939
R14673 gnd.n715 gnd.n714 0.152939
R14674 gnd.n720 gnd.n715 0.152939
R14675 gnd.n721 gnd.n720 0.152939
R14676 gnd.n722 gnd.n721 0.152939
R14677 gnd.n723 gnd.n722 0.152939
R14678 gnd.n728 gnd.n723 0.152939
R14679 gnd.n729 gnd.n728 0.152939
R14680 gnd.n730 gnd.n729 0.152939
R14681 gnd.n731 gnd.n730 0.152939
R14682 gnd.n736 gnd.n731 0.152939
R14683 gnd.n737 gnd.n736 0.152939
R14684 gnd.n738 gnd.n737 0.152939
R14685 gnd.n739 gnd.n738 0.152939
R14686 gnd.n744 gnd.n739 0.152939
R14687 gnd.n745 gnd.n744 0.152939
R14688 gnd.n746 gnd.n745 0.152939
R14689 gnd.n747 gnd.n746 0.152939
R14690 gnd.n752 gnd.n747 0.152939
R14691 gnd.n753 gnd.n752 0.152939
R14692 gnd.n754 gnd.n753 0.152939
R14693 gnd.n755 gnd.n754 0.152939
R14694 gnd.n760 gnd.n755 0.152939
R14695 gnd.n761 gnd.n760 0.152939
R14696 gnd.n762 gnd.n761 0.152939
R14697 gnd.n763 gnd.n762 0.152939
R14698 gnd.n768 gnd.n763 0.152939
R14699 gnd.n769 gnd.n768 0.152939
R14700 gnd.n770 gnd.n769 0.152939
R14701 gnd.n771 gnd.n770 0.152939
R14702 gnd.n776 gnd.n771 0.152939
R14703 gnd.n777 gnd.n776 0.152939
R14704 gnd.n778 gnd.n777 0.152939
R14705 gnd.n779 gnd.n778 0.152939
R14706 gnd.n784 gnd.n779 0.152939
R14707 gnd.n785 gnd.n784 0.152939
R14708 gnd.n786 gnd.n785 0.152939
R14709 gnd.n787 gnd.n786 0.152939
R14710 gnd.n792 gnd.n787 0.152939
R14711 gnd.n793 gnd.n792 0.152939
R14712 gnd.n794 gnd.n793 0.152939
R14713 gnd.n795 gnd.n794 0.152939
R14714 gnd.n800 gnd.n795 0.152939
R14715 gnd.n801 gnd.n800 0.152939
R14716 gnd.n802 gnd.n801 0.152939
R14717 gnd.n803 gnd.n802 0.152939
R14718 gnd.n808 gnd.n803 0.152939
R14719 gnd.n809 gnd.n808 0.152939
R14720 gnd.n810 gnd.n809 0.152939
R14721 gnd.n811 gnd.n810 0.152939
R14722 gnd.n816 gnd.n811 0.152939
R14723 gnd.n817 gnd.n816 0.152939
R14724 gnd.n818 gnd.n817 0.152939
R14725 gnd.n819 gnd.n818 0.152939
R14726 gnd.n824 gnd.n819 0.152939
R14727 gnd.n825 gnd.n824 0.152939
R14728 gnd.n826 gnd.n825 0.152939
R14729 gnd.n827 gnd.n826 0.152939
R14730 gnd.n832 gnd.n827 0.152939
R14731 gnd.n833 gnd.n832 0.152939
R14732 gnd.n834 gnd.n833 0.152939
R14733 gnd.n835 gnd.n834 0.152939
R14734 gnd.n840 gnd.n835 0.152939
R14735 gnd.n841 gnd.n840 0.152939
R14736 gnd.n842 gnd.n841 0.152939
R14737 gnd.n843 gnd.n842 0.152939
R14738 gnd.n3684 gnd.n843 0.152939
R14739 gnd.n3685 gnd.n3684 0.152939
R14740 gnd.n5426 gnd.n2959 0.152939
R14741 gnd.n5422 gnd.n2959 0.152939
R14742 gnd.n5422 gnd.n5421 0.152939
R14743 gnd.n5421 gnd.n5420 0.152939
R14744 gnd.n5420 gnd.n3087 0.152939
R14745 gnd.n5413 gnd.n3087 0.152939
R14746 gnd.n5413 gnd.n5412 0.152939
R14747 gnd.n5412 gnd.n5411 0.152939
R14748 gnd.n5411 gnd.n5404 0.152939
R14749 gnd.n4427 gnd.n4426 0.152939
R14750 gnd.n4428 gnd.n4427 0.152939
R14751 gnd.n4428 gnd.n3414 0.152939
R14752 gnd.n4444 gnd.n3414 0.152939
R14753 gnd.n4445 gnd.n4444 0.152939
R14754 gnd.n4447 gnd.n4445 0.152939
R14755 gnd.n4447 gnd.n4446 0.152939
R14756 gnd.n4446 gnd.n3383 0.152939
R14757 gnd.n4566 gnd.n3383 0.152939
R14758 gnd.n4567 gnd.n4566 0.152939
R14759 gnd.n4568 gnd.n4567 0.152939
R14760 gnd.n4568 gnd.n3369 0.152939
R14761 gnd.n4582 gnd.n3369 0.152939
R14762 gnd.n4583 gnd.n4582 0.152939
R14763 gnd.n4584 gnd.n4583 0.152939
R14764 gnd.n4584 gnd.n3355 0.152939
R14765 gnd.n4598 gnd.n3355 0.152939
R14766 gnd.n4599 gnd.n4598 0.152939
R14767 gnd.n4600 gnd.n4599 0.152939
R14768 gnd.n4600 gnd.n3339 0.152939
R14769 gnd.n4615 gnd.n3339 0.152939
R14770 gnd.n4616 gnd.n4615 0.152939
R14771 gnd.n4618 gnd.n4616 0.152939
R14772 gnd.n4618 gnd.n4617 0.152939
R14773 gnd.n4617 gnd.n3308 0.152939
R14774 gnd.n4739 gnd.n3308 0.152939
R14775 gnd.n4740 gnd.n4739 0.152939
R14776 gnd.n4741 gnd.n4740 0.152939
R14777 gnd.n4741 gnd.n3295 0.152939
R14778 gnd.n4755 gnd.n3295 0.152939
R14779 gnd.n4756 gnd.n4755 0.152939
R14780 gnd.n4757 gnd.n4756 0.152939
R14781 gnd.n4757 gnd.n3283 0.152939
R14782 gnd.n4771 gnd.n3283 0.152939
R14783 gnd.n4772 gnd.n4771 0.152939
R14784 gnd.n4773 gnd.n4772 0.152939
R14785 gnd.n4773 gnd.n3269 0.152939
R14786 gnd.n4789 gnd.n3269 0.152939
R14787 gnd.n4790 gnd.n4789 0.152939
R14788 gnd.n4792 gnd.n4790 0.152939
R14789 gnd.n4792 gnd.n4791 0.152939
R14790 gnd.n4791 gnd.n3236 0.152939
R14791 gnd.n4910 gnd.n3236 0.152939
R14792 gnd.n4911 gnd.n4910 0.152939
R14793 gnd.n4912 gnd.n4911 0.152939
R14794 gnd.n4912 gnd.n3221 0.152939
R14795 gnd.n4926 gnd.n3221 0.152939
R14796 gnd.n4927 gnd.n4926 0.152939
R14797 gnd.n4928 gnd.n4927 0.152939
R14798 gnd.n4928 gnd.n3207 0.152939
R14799 gnd.n4942 gnd.n3207 0.152939
R14800 gnd.n4943 gnd.n4942 0.152939
R14801 gnd.n4944 gnd.n4943 0.152939
R14802 gnd.n4944 gnd.n3192 0.152939
R14803 gnd.n4960 gnd.n3192 0.152939
R14804 gnd.n4961 gnd.n4960 0.152939
R14805 gnd.n4963 gnd.n4961 0.152939
R14806 gnd.n4963 gnd.n4962 0.152939
R14807 gnd.n4962 gnd.n3162 0.152939
R14808 gnd.n5316 gnd.n3162 0.152939
R14809 gnd.n5317 gnd.n5316 0.152939
R14810 gnd.n5318 gnd.n5317 0.152939
R14811 gnd.n5318 gnd.n3149 0.152939
R14812 gnd.n5332 gnd.n3149 0.152939
R14813 gnd.n5333 gnd.n5332 0.152939
R14814 gnd.n5334 gnd.n5333 0.152939
R14815 gnd.n5334 gnd.n3136 0.152939
R14816 gnd.n5348 gnd.n3136 0.152939
R14817 gnd.n5349 gnd.n5348 0.152939
R14818 gnd.n5350 gnd.n5349 0.152939
R14819 gnd.n5350 gnd.n3122 0.152939
R14820 gnd.n5364 gnd.n3122 0.152939
R14821 gnd.n5365 gnd.n5364 0.152939
R14822 gnd.n5366 gnd.n5365 0.152939
R14823 gnd.n5366 gnd.n3108 0.152939
R14824 gnd.n5380 gnd.n3108 0.152939
R14825 gnd.n5381 gnd.n5380 0.152939
R14826 gnd.n5384 gnd.n5381 0.152939
R14827 gnd.n5384 gnd.n5383 0.152939
R14828 gnd.n5383 gnd.n5382 0.152939
R14829 gnd.n5382 gnd.n3095 0.152939
R14830 gnd.n5403 gnd.n3095 0.152939
R14831 gnd.n4391 gnd.n3460 0.152939
R14832 gnd.n4399 gnd.n3460 0.152939
R14833 gnd.n4400 gnd.n4399 0.152939
R14834 gnd.n4401 gnd.n4400 0.152939
R14835 gnd.n4401 gnd.n3456 0.152939
R14836 gnd.n4409 gnd.n3456 0.152939
R14837 gnd.n4410 gnd.n4409 0.152939
R14838 gnd.n4411 gnd.n4410 0.152939
R14839 gnd.n4411 gnd.n3430 0.152939
R14840 gnd.n3992 gnd.n3991 0.152939
R14841 gnd.n3992 gnd.n3673 0.152939
R14842 gnd.n4006 gnd.n3673 0.152939
R14843 gnd.n4007 gnd.n4006 0.152939
R14844 gnd.n4008 gnd.n4007 0.152939
R14845 gnd.n4008 gnd.n3666 0.152939
R14846 gnd.n4022 gnd.n3666 0.152939
R14847 gnd.n4023 gnd.n4022 0.152939
R14848 gnd.n4024 gnd.n4023 0.152939
R14849 gnd.n4024 gnd.n3660 0.152939
R14850 gnd.n4038 gnd.n3660 0.152939
R14851 gnd.n4039 gnd.n4038 0.152939
R14852 gnd.n4040 gnd.n4039 0.152939
R14853 gnd.n4040 gnd.n3653 0.152939
R14854 gnd.n4054 gnd.n3653 0.152939
R14855 gnd.n4055 gnd.n4054 0.152939
R14856 gnd.n4056 gnd.n4055 0.152939
R14857 gnd.n4056 gnd.n3647 0.152939
R14858 gnd.n4070 gnd.n3647 0.152939
R14859 gnd.n4071 gnd.n4070 0.152939
R14860 gnd.n4072 gnd.n4071 0.152939
R14861 gnd.n4072 gnd.n3641 0.152939
R14862 gnd.n4087 gnd.n3641 0.152939
R14863 gnd.n4088 gnd.n4087 0.152939
R14864 gnd.n4089 gnd.n4088 0.152939
R14865 gnd.n4089 gnd.n3462 0.152939
R14866 gnd.n5832 gnd.n2577 0.152939
R14867 gnd.n5828 gnd.n2577 0.152939
R14868 gnd.n5828 gnd.n5827 0.152939
R14869 gnd.n5827 gnd.n5826 0.152939
R14870 gnd.n5826 gnd.n2582 0.152939
R14871 gnd.n5822 gnd.n2582 0.152939
R14872 gnd.n5822 gnd.n5821 0.152939
R14873 gnd.n5821 gnd.n5820 0.152939
R14874 gnd.n5820 gnd.n2587 0.152939
R14875 gnd.n5816 gnd.n2587 0.152939
R14876 gnd.n5816 gnd.n5815 0.152939
R14877 gnd.n5815 gnd.n5814 0.152939
R14878 gnd.n5814 gnd.n2592 0.152939
R14879 gnd.n5810 gnd.n2592 0.152939
R14880 gnd.n5810 gnd.n5809 0.152939
R14881 gnd.n5809 gnd.n5808 0.152939
R14882 gnd.n5808 gnd.n2597 0.152939
R14883 gnd.n5804 gnd.n2597 0.152939
R14884 gnd.n5804 gnd.n5803 0.152939
R14885 gnd.n5803 gnd.n5802 0.152939
R14886 gnd.n5802 gnd.n2602 0.152939
R14887 gnd.n5798 gnd.n2602 0.152939
R14888 gnd.n5798 gnd.n5797 0.152939
R14889 gnd.n5797 gnd.n5796 0.152939
R14890 gnd.n5796 gnd.n2607 0.152939
R14891 gnd.n5792 gnd.n2607 0.152939
R14892 gnd.n5792 gnd.n5791 0.152939
R14893 gnd.n5791 gnd.n5790 0.152939
R14894 gnd.n5790 gnd.n2612 0.152939
R14895 gnd.n5786 gnd.n2612 0.152939
R14896 gnd.n5786 gnd.n5785 0.152939
R14897 gnd.n5785 gnd.n5784 0.152939
R14898 gnd.n5784 gnd.n2617 0.152939
R14899 gnd.n5780 gnd.n2617 0.152939
R14900 gnd.n5780 gnd.n5779 0.152939
R14901 gnd.n5779 gnd.n5778 0.152939
R14902 gnd.n5778 gnd.n2622 0.152939
R14903 gnd.n5774 gnd.n2622 0.152939
R14904 gnd.n5774 gnd.n5773 0.152939
R14905 gnd.n5773 gnd.n5772 0.152939
R14906 gnd.n5772 gnd.n2627 0.152939
R14907 gnd.n5768 gnd.n2627 0.152939
R14908 gnd.n5768 gnd.n5767 0.152939
R14909 gnd.n5767 gnd.n5766 0.152939
R14910 gnd.n5766 gnd.n2632 0.152939
R14911 gnd.n5762 gnd.n2632 0.152939
R14912 gnd.n5762 gnd.n5761 0.152939
R14913 gnd.n5761 gnd.n5760 0.152939
R14914 gnd.n5760 gnd.n2637 0.152939
R14915 gnd.n5756 gnd.n2637 0.152939
R14916 gnd.n5756 gnd.n5755 0.152939
R14917 gnd.n5755 gnd.n5754 0.152939
R14918 gnd.n5754 gnd.n2642 0.152939
R14919 gnd.n5750 gnd.n2642 0.152939
R14920 gnd.n5750 gnd.n5749 0.152939
R14921 gnd.n5749 gnd.n5748 0.152939
R14922 gnd.n5748 gnd.n2647 0.152939
R14923 gnd.n5744 gnd.n2647 0.152939
R14924 gnd.n5744 gnd.n5743 0.152939
R14925 gnd.n5743 gnd.n5742 0.152939
R14926 gnd.n5742 gnd.n2652 0.152939
R14927 gnd.n5738 gnd.n2652 0.152939
R14928 gnd.n5738 gnd.n5737 0.152939
R14929 gnd.n5737 gnd.n5736 0.152939
R14930 gnd.n5736 gnd.n2657 0.152939
R14931 gnd.n5732 gnd.n2657 0.152939
R14932 gnd.n5732 gnd.n5731 0.152939
R14933 gnd.n5731 gnd.n5730 0.152939
R14934 gnd.n5730 gnd.n2662 0.152939
R14935 gnd.n5726 gnd.n2662 0.152939
R14936 gnd.n5726 gnd.n5725 0.152939
R14937 gnd.n5725 gnd.n5724 0.152939
R14938 gnd.n5724 gnd.n2667 0.152939
R14939 gnd.n5720 gnd.n2667 0.152939
R14940 gnd.n5720 gnd.n5719 0.152939
R14941 gnd.n5719 gnd.n5718 0.152939
R14942 gnd.n5718 gnd.n2672 0.152939
R14943 gnd.n5714 gnd.n2672 0.152939
R14944 gnd.n5714 gnd.n5713 0.152939
R14945 gnd.n5713 gnd.n5712 0.152939
R14946 gnd.n5712 gnd.n2677 0.152939
R14947 gnd.n2680 gnd.n2677 0.152939
R14948 gnd.n5619 gnd.n5618 0.152939
R14949 gnd.n5618 gnd.n5617 0.152939
R14950 gnd.n5617 gnd.n2779 0.152939
R14951 gnd.n5613 gnd.n2779 0.152939
R14952 gnd.n5613 gnd.n5612 0.152939
R14953 gnd.n5612 gnd.n5611 0.152939
R14954 gnd.n5611 gnd.n2784 0.152939
R14955 gnd.n5607 gnd.n2784 0.152939
R14956 gnd.n5607 gnd.n5606 0.152939
R14957 gnd.n5606 gnd.n5605 0.152939
R14958 gnd.n5605 gnd.n2789 0.152939
R14959 gnd.n5601 gnd.n2789 0.152939
R14960 gnd.n5601 gnd.n5600 0.152939
R14961 gnd.n5600 gnd.n5599 0.152939
R14962 gnd.n5599 gnd.n2794 0.152939
R14963 gnd.n5595 gnd.n2794 0.152939
R14964 gnd.n5595 gnd.n5594 0.152939
R14965 gnd.n5594 gnd.n5593 0.152939
R14966 gnd.n5593 gnd.n2799 0.152939
R14967 gnd.n5589 gnd.n2799 0.152939
R14968 gnd.n5589 gnd.n280 0.152939
R14969 gnd.n7035 gnd.n280 0.152939
R14970 gnd.n7035 gnd.n7034 0.152939
R14971 gnd.n7034 gnd.n7033 0.152939
R14972 gnd.n7033 gnd.n281 0.152939
R14973 gnd.n7029 gnd.n281 0.152939
R14974 gnd.n7027 gnd.n7026 0.152939
R14975 gnd.n7026 gnd.n287 0.152939
R14976 gnd.n287 gnd.n255 0.152939
R14977 gnd.n7048 gnd.n255 0.152939
R14978 gnd.n7049 gnd.n7048 0.152939
R14979 gnd.n7050 gnd.n7049 0.152939
R14980 gnd.n7050 gnd.n240 0.152939
R14981 gnd.n7064 gnd.n240 0.152939
R14982 gnd.n7065 gnd.n7064 0.152939
R14983 gnd.n7066 gnd.n7065 0.152939
R14984 gnd.n7066 gnd.n225 0.152939
R14985 gnd.n7080 gnd.n225 0.152939
R14986 gnd.n7081 gnd.n7080 0.152939
R14987 gnd.n7082 gnd.n7081 0.152939
R14988 gnd.n7082 gnd.n210 0.152939
R14989 gnd.n7096 gnd.n210 0.152939
R14990 gnd.n7097 gnd.n7096 0.152939
R14991 gnd.n7098 gnd.n7097 0.152939
R14992 gnd.n7098 gnd.n195 0.152939
R14993 gnd.n7112 gnd.n195 0.152939
R14994 gnd.n7113 gnd.n7112 0.152939
R14995 gnd.n7189 gnd.n7113 0.152939
R14996 gnd.n7189 gnd.n7188 0.152939
R14997 gnd.n7188 gnd.n7187 0.152939
R14998 gnd.n7187 gnd.n7114 0.152939
R14999 gnd.n7183 gnd.n7114 0.152939
R15000 gnd.n7182 gnd.n7116 0.152939
R15001 gnd.n7178 gnd.n7116 0.152939
R15002 gnd.n7178 gnd.n7177 0.152939
R15003 gnd.n7177 gnd.n7176 0.152939
R15004 gnd.n7176 gnd.n7122 0.152939
R15005 gnd.n7172 gnd.n7122 0.152939
R15006 gnd.n7172 gnd.n7171 0.152939
R15007 gnd.n7171 gnd.n7170 0.152939
R15008 gnd.n7170 gnd.n7130 0.152939
R15009 gnd.n7166 gnd.n7130 0.152939
R15010 gnd.n7166 gnd.n7165 0.152939
R15011 gnd.n7165 gnd.n7164 0.152939
R15012 gnd.n7164 gnd.n7138 0.152939
R15013 gnd.n7160 gnd.n7138 0.152939
R15014 gnd.n7160 gnd.n7159 0.152939
R15015 gnd.n7159 gnd.n7158 0.152939
R15016 gnd.n7158 gnd.n7146 0.152939
R15017 gnd.n7154 gnd.n7146 0.152939
R15018 gnd.n5430 gnd.n5429 0.152939
R15019 gnd.n5432 gnd.n5430 0.152939
R15020 gnd.n5432 gnd.n5431 0.152939
R15021 gnd.n5431 gnd.n2888 0.152939
R15022 gnd.n5460 gnd.n2888 0.152939
R15023 gnd.n5461 gnd.n5460 0.152939
R15024 gnd.n5463 gnd.n5461 0.152939
R15025 gnd.n5463 gnd.n5462 0.152939
R15026 gnd.n5462 gnd.n2860 0.152939
R15027 gnd.n5491 gnd.n2860 0.152939
R15028 gnd.n5492 gnd.n5491 0.152939
R15029 gnd.n5499 gnd.n5492 0.152939
R15030 gnd.n5499 gnd.n5498 0.152939
R15031 gnd.n5498 gnd.n5497 0.152939
R15032 gnd.n5497 gnd.n5493 0.152939
R15033 gnd.n5493 gnd.n2826 0.152939
R15034 gnd.n5556 gnd.n2826 0.152939
R15035 gnd.n5556 gnd.n5555 0.152939
R15036 gnd.n5555 gnd.n5554 0.152939
R15037 gnd.n5554 gnd.n2827 0.152939
R15038 gnd.n5550 gnd.n2827 0.152939
R15039 gnd.n5550 gnd.n305 0.152939
R15040 gnd.n6942 gnd.n305 0.152939
R15041 gnd.n6943 gnd.n6942 0.152939
R15042 gnd.n6944 gnd.n6943 0.152939
R15043 gnd.n6944 gnd.n63 0.152939
R15044 gnd.n7321 gnd.n64 0.152939
R15045 gnd.n7317 gnd.n64 0.152939
R15046 gnd.n7317 gnd.n7316 0.152939
R15047 gnd.n7316 gnd.n7315 0.152939
R15048 gnd.n7315 gnd.n70 0.152939
R15049 gnd.n7311 gnd.n70 0.152939
R15050 gnd.n7311 gnd.n7310 0.152939
R15051 gnd.n7310 gnd.n7309 0.152939
R15052 gnd.n7309 gnd.n75 0.152939
R15053 gnd.n7305 gnd.n75 0.152939
R15054 gnd.n7305 gnd.n7304 0.152939
R15055 gnd.n7304 gnd.n7303 0.152939
R15056 gnd.n7303 gnd.n80 0.152939
R15057 gnd.n7299 gnd.n80 0.152939
R15058 gnd.n7299 gnd.n7298 0.152939
R15059 gnd.n7298 gnd.n7297 0.152939
R15060 gnd.n7297 gnd.n85 0.152939
R15061 gnd.n7293 gnd.n85 0.152939
R15062 gnd.n7293 gnd.n7292 0.152939
R15063 gnd.n7292 gnd.n7291 0.152939
R15064 gnd.n7291 gnd.n90 0.152939
R15065 gnd.n7287 gnd.n90 0.152939
R15066 gnd.n7287 gnd.n7286 0.152939
R15067 gnd.n7286 gnd.n7285 0.152939
R15068 gnd.n7285 gnd.n95 0.152939
R15069 gnd.n98 gnd.n95 0.152939
R15070 gnd.n5427 gnd.n5426 0.151415
R15071 gnd.n4391 gnd.n4390 0.151415
R15072 gnd.n318 gnd.n263 0.128549
R15073 gnd.n3693 gnd.n3692 0.128549
R15074 gnd.n1993 gnd.n1992 0.0767195
R15075 gnd.n1992 gnd.n1991 0.0767195
R15076 gnd.n7042 gnd.n248 0.0767195
R15077 gnd.n295 gnd.n286 0.0767195
R15078 gnd.n6956 gnd.n286 0.0767195
R15079 gnd.n7042 gnd.n262 0.0767195
R15080 gnd.n2459 gnd.n2421 0.0767195
R15081 gnd.n3981 gnd.n2430 0.0767195
R15082 gnd.n3981 gnd.n2431 0.0767195
R15083 gnd.n3983 gnd.n3982 0.0767195
R15084 gnd.n3982 gnd.n3676 0.0767195
R15085 gnd.n2421 gnd.n2402 0.0767195
R15086 gnd.n7029 gnd.n7028 0.0767195
R15087 gnd.n7028 gnd.n7027 0.0767195
R15088 gnd.n7322 gnd.n63 0.0767195
R15089 gnd.n7322 gnd.n7321 0.0767195
R15090 gnd.n3990 gnd.n3989 0.0695946
R15091 gnd.n3991 gnd.n3990 0.0695946
R15092 gnd.n5834 gnd.n5833 0.063
R15093 gnd.n3003 gnd.n2778 0.063
R15094 gnd.n6135 gnd.n876 0.0477147
R15095 gnd.n1756 gnd.n1644 0.0442063
R15096 gnd.n1757 gnd.n1756 0.0442063
R15097 gnd.n1758 gnd.n1757 0.0442063
R15098 gnd.n1758 gnd.n1633 0.0442063
R15099 gnd.n1772 gnd.n1633 0.0442063
R15100 gnd.n1773 gnd.n1772 0.0442063
R15101 gnd.n1774 gnd.n1773 0.0442063
R15102 gnd.n1774 gnd.n1620 0.0442063
R15103 gnd.n1818 gnd.n1620 0.0442063
R15104 gnd.n1819 gnd.n1818 0.0442063
R15105 gnd.n1821 gnd.n1554 0.0344674
R15106 gnd.n2965 gnd.n2958 0.0344674
R15107 gnd.n4389 gnd.n4388 0.0344674
R15108 gnd.n1841 gnd.n1840 0.0269946
R15109 gnd.n1843 gnd.n1842 0.0269946
R15110 gnd.n1549 gnd.n1547 0.0269946
R15111 gnd.n1853 gnd.n1851 0.0269946
R15112 gnd.n1852 gnd.n1528 0.0269946
R15113 gnd.n1872 gnd.n1871 0.0269946
R15114 gnd.n1874 gnd.n1873 0.0269946
R15115 gnd.n1523 gnd.n1522 0.0269946
R15116 gnd.n1884 gnd.n1518 0.0269946
R15117 gnd.n1883 gnd.n1520 0.0269946
R15118 gnd.n1519 gnd.n1501 0.0269946
R15119 gnd.n1904 gnd.n1502 0.0269946
R15120 gnd.n1903 gnd.n1503 0.0269946
R15121 gnd.n1937 gnd.n1478 0.0269946
R15122 gnd.n1939 gnd.n1938 0.0269946
R15123 gnd.n1940 gnd.n1425 0.0269946
R15124 gnd.n1473 gnd.n1426 0.0269946
R15125 gnd.n1475 gnd.n1427 0.0269946
R15126 gnd.n1950 gnd.n1949 0.0269946
R15127 gnd.n1952 gnd.n1951 0.0269946
R15128 gnd.n1953 gnd.n1447 0.0269946
R15129 gnd.n1955 gnd.n1448 0.0269946
R15130 gnd.n1958 gnd.n1449 0.0269946
R15131 gnd.n1961 gnd.n1960 0.0269946
R15132 gnd.n1963 gnd.n1962 0.0269946
R15133 gnd.n2028 gnd.n1348 0.0269946
R15134 gnd.n2030 gnd.n2029 0.0269946
R15135 gnd.n2039 gnd.n1341 0.0269946
R15136 gnd.n2041 gnd.n2040 0.0269946
R15137 gnd.n2042 gnd.n1339 0.0269946
R15138 gnd.n2049 gnd.n2045 0.0269946
R15139 gnd.n2048 gnd.n2047 0.0269946
R15140 gnd.n2046 gnd.n1318 0.0269946
R15141 gnd.n2071 gnd.n1319 0.0269946
R15142 gnd.n2070 gnd.n1320 0.0269946
R15143 gnd.n2113 gnd.n1293 0.0269946
R15144 gnd.n2115 gnd.n2114 0.0269946
R15145 gnd.n2124 gnd.n1286 0.0269946
R15146 gnd.n2126 gnd.n2125 0.0269946
R15147 gnd.n2127 gnd.n1284 0.0269946
R15148 gnd.n2134 gnd.n2130 0.0269946
R15149 gnd.n2133 gnd.n2132 0.0269946
R15150 gnd.n2131 gnd.n1263 0.0269946
R15151 gnd.n2158 gnd.n1264 0.0269946
R15152 gnd.n2157 gnd.n1265 0.0269946
R15153 gnd.n2204 gnd.n1240 0.0269946
R15154 gnd.n2206 gnd.n2205 0.0269946
R15155 gnd.n2207 gnd.n852 0.0269946
R15156 gnd.n1237 gnd.n854 0.0269946
R15157 gnd.n2215 gnd.n2214 0.0269946
R15158 gnd.n2217 gnd.n2216 0.0269946
R15159 gnd.n6136 gnd.n875 0.0269946
R15160 gnd.n315 gnd.n263 0.0248902
R15161 gnd.n3694 gnd.n3693 0.0248902
R15162 gnd.n3004 gnd.n3003 0.0246168
R15163 gnd.n5833 gnd.n2576 0.0246168
R15164 gnd.n1821 gnd.n1820 0.0202011
R15165 gnd.n3004 gnd.n3001 0.0174837
R15166 gnd.n3009 gnd.n3001 0.0174837
R15167 gnd.n3010 gnd.n3009 0.0174837
R15168 gnd.n3010 gnd.n2999 0.0174837
R15169 gnd.n3017 gnd.n2999 0.0174837
R15170 gnd.n3019 gnd.n3017 0.0174837
R15171 gnd.n3019 gnd.n3018 0.0174837
R15172 gnd.n3018 gnd.n2994 0.0174837
R15173 gnd.n3026 gnd.n2994 0.0174837
R15174 gnd.n3026 gnd.n3025 0.0174837
R15175 gnd.n3025 gnd.n2995 0.0174837
R15176 gnd.n2995 gnd.n2990 0.0174837
R15177 gnd.n3034 gnd.n2990 0.0174837
R15178 gnd.n3036 gnd.n3034 0.0174837
R15179 gnd.n3036 gnd.n3035 0.0174837
R15180 gnd.n3035 gnd.n2985 0.0174837
R15181 gnd.n3043 gnd.n2985 0.0174837
R15182 gnd.n3043 gnd.n3042 0.0174837
R15183 gnd.n3042 gnd.n2986 0.0174837
R15184 gnd.n2986 gnd.n2981 0.0174837
R15185 gnd.n3051 gnd.n2981 0.0174837
R15186 gnd.n3053 gnd.n3051 0.0174837
R15187 gnd.n3053 gnd.n3052 0.0174837
R15188 gnd.n3052 gnd.n2976 0.0174837
R15189 gnd.n3060 gnd.n2976 0.0174837
R15190 gnd.n3060 gnd.n3059 0.0174837
R15191 gnd.n3059 gnd.n2977 0.0174837
R15192 gnd.n2977 gnd.n2972 0.0174837
R15193 gnd.n3068 gnd.n2972 0.0174837
R15194 gnd.n3070 gnd.n3068 0.0174837
R15195 gnd.n3070 gnd.n3069 0.0174837
R15196 gnd.n3069 gnd.n2964 0.0174837
R15197 gnd.n3075 gnd.n2964 0.0174837
R15198 gnd.n3075 gnd.n3074 0.0174837
R15199 gnd.n3074 gnd.n2965 0.0174837
R15200 gnd.n3510 gnd.n2576 0.0174837
R15201 gnd.n3510 gnd.n3509 0.0174837
R15202 gnd.n3516 gnd.n3509 0.0174837
R15203 gnd.n3517 gnd.n3516 0.0174837
R15204 gnd.n3517 gnd.n3503 0.0174837
R15205 gnd.n3522 gnd.n3503 0.0174837
R15206 gnd.n3523 gnd.n3522 0.0174837
R15207 gnd.n3523 gnd.n3501 0.0174837
R15208 gnd.n3528 gnd.n3501 0.0174837
R15209 gnd.n3529 gnd.n3528 0.0174837
R15210 gnd.n3529 gnd.n3499 0.0174837
R15211 gnd.n3534 gnd.n3499 0.0174837
R15212 gnd.n3535 gnd.n3534 0.0174837
R15213 gnd.n3535 gnd.n3495 0.0174837
R15214 gnd.n3540 gnd.n3495 0.0174837
R15215 gnd.n3541 gnd.n3540 0.0174837
R15216 gnd.n3541 gnd.n3491 0.0174837
R15217 gnd.n3546 gnd.n3491 0.0174837
R15218 gnd.n3547 gnd.n3546 0.0174837
R15219 gnd.n3547 gnd.n3489 0.0174837
R15220 gnd.n3552 gnd.n3489 0.0174837
R15221 gnd.n3553 gnd.n3552 0.0174837
R15222 gnd.n3553 gnd.n3487 0.0174837
R15223 gnd.n3558 gnd.n3487 0.0174837
R15224 gnd.n3560 gnd.n3558 0.0174837
R15225 gnd.n3560 gnd.n3559 0.0174837
R15226 gnd.n3559 gnd.n3482 0.0174837
R15227 gnd.n3567 gnd.n3482 0.0174837
R15228 gnd.n3567 gnd.n3566 0.0174837
R15229 gnd.n3566 gnd.n3483 0.0174837
R15230 gnd.n3483 gnd.n3467 0.0174837
R15231 gnd.n4382 gnd.n3467 0.0174837
R15232 gnd.n4383 gnd.n4382 0.0174837
R15233 gnd.n4383 gnd.n3463 0.0174837
R15234 gnd.n4388 gnd.n3463 0.0174837
R15235 gnd.n1820 gnd.n1819 0.0148637
R15236 gnd.n1235 gnd.n1234 0.0144266
R15237 gnd.n1234 gnd.n853 0.0130679
R15238 gnd.n1840 gnd.n1554 0.00797283
R15239 gnd.n1842 gnd.n1841 0.00797283
R15240 gnd.n1843 gnd.n1549 0.00797283
R15241 gnd.n1851 gnd.n1547 0.00797283
R15242 gnd.n1853 gnd.n1852 0.00797283
R15243 gnd.n1871 gnd.n1528 0.00797283
R15244 gnd.n1873 gnd.n1872 0.00797283
R15245 gnd.n1874 gnd.n1523 0.00797283
R15246 gnd.n1522 gnd.n1518 0.00797283
R15247 gnd.n1884 gnd.n1883 0.00797283
R15248 gnd.n1520 gnd.n1519 0.00797283
R15249 gnd.n1502 gnd.n1501 0.00797283
R15250 gnd.n1904 gnd.n1903 0.00797283
R15251 gnd.n1503 gnd.n1478 0.00797283
R15252 gnd.n1938 gnd.n1937 0.00797283
R15253 gnd.n1940 gnd.n1939 0.00797283
R15254 gnd.n1473 gnd.n1425 0.00797283
R15255 gnd.n1475 gnd.n1426 0.00797283
R15256 gnd.n1949 gnd.n1427 0.00797283
R15257 gnd.n1951 gnd.n1950 0.00797283
R15258 gnd.n1953 gnd.n1952 0.00797283
R15259 gnd.n1955 gnd.n1447 0.00797283
R15260 gnd.n1958 gnd.n1448 0.00797283
R15261 gnd.n1960 gnd.n1449 0.00797283
R15262 gnd.n1963 gnd.n1961 0.00797283
R15263 gnd.n1962 gnd.n1348 0.00797283
R15264 gnd.n2030 gnd.n2028 0.00797283
R15265 gnd.n2029 gnd.n1341 0.00797283
R15266 gnd.n2040 gnd.n2039 0.00797283
R15267 gnd.n2042 gnd.n2041 0.00797283
R15268 gnd.n2045 gnd.n1339 0.00797283
R15269 gnd.n2049 gnd.n2048 0.00797283
R15270 gnd.n2047 gnd.n2046 0.00797283
R15271 gnd.n1319 gnd.n1318 0.00797283
R15272 gnd.n2071 gnd.n2070 0.00797283
R15273 gnd.n1320 gnd.n1293 0.00797283
R15274 gnd.n2115 gnd.n2113 0.00797283
R15275 gnd.n2114 gnd.n1286 0.00797283
R15276 gnd.n2125 gnd.n2124 0.00797283
R15277 gnd.n2127 gnd.n2126 0.00797283
R15278 gnd.n2130 gnd.n1284 0.00797283
R15279 gnd.n2134 gnd.n2133 0.00797283
R15280 gnd.n2132 gnd.n2131 0.00797283
R15281 gnd.n1264 gnd.n1263 0.00797283
R15282 gnd.n2158 gnd.n2157 0.00797283
R15283 gnd.n1265 gnd.n1240 0.00797283
R15284 gnd.n2205 gnd.n2204 0.00797283
R15285 gnd.n2207 gnd.n2206 0.00797283
R15286 gnd.n1235 gnd.n852 0.00797283
R15287 gnd.n1237 gnd.n853 0.00797283
R15288 gnd.n2214 gnd.n854 0.00797283
R15289 gnd.n2217 gnd.n2215 0.00797283
R15290 gnd.n2216 gnd.n875 0.00797283
R15291 gnd.n6136 gnd.n6135 0.00797283
R15292 gnd.n7028 gnd.n286 0.00507153
R15293 gnd.n3982 gnd.n3981 0.00507153
R15294 gnd.n5427 gnd.n2958 0.000839674
R15295 gnd.n4390 gnd.n4389 0.000839674
R15296 a_n6972_8799.n185 a_n6972_8799.t57 485.149
R15297 a_n6972_8799.n201 a_n6972_8799.t71 485.149
R15298 a_n6972_8799.n218 a_n6972_8799.t120 485.149
R15299 a_n6972_8799.n134 a_n6972_8799.t115 485.149
R15300 a_n6972_8799.n150 a_n6972_8799.t125 485.149
R15301 a_n6972_8799.n167 a_n6972_8799.t118 485.149
R15302 a_n6972_8799.n195 a_n6972_8799.t80 464.166
R15303 a_n6972_8799.n194 a_n6972_8799.t79 464.166
R15304 a_n6972_8799.n180 a_n6972_8799.t58 464.166
R15305 a_n6972_8799.n193 a_n6972_8799.t116 464.166
R15306 a_n6972_8799.n192 a_n6972_8799.t81 464.166
R15307 a_n6972_8799.n181 a_n6972_8799.t63 464.166
R15308 a_n6972_8799.n191 a_n6972_8799.t119 464.166
R15309 a_n6972_8799.n190 a_n6972_8799.t95 464.166
R15310 a_n6972_8799.n182 a_n6972_8799.t93 464.166
R15311 a_n6972_8799.n189 a_n6972_8799.t40 464.166
R15312 a_n6972_8799.n188 a_n6972_8799.t99 464.166
R15313 a_n6972_8799.n183 a_n6972_8799.t98 464.166
R15314 a_n6972_8799.n187 a_n6972_8799.t42 464.166
R15315 a_n6972_8799.n186 a_n6972_8799.t41 464.166
R15316 a_n6972_8799.n184 a_n6972_8799.t112 464.166
R15317 a_n6972_8799.n211 a_n6972_8799.t87 464.166
R15318 a_n6972_8799.n210 a_n6972_8799.t86 464.166
R15319 a_n6972_8799.n196 a_n6972_8799.t70 464.166
R15320 a_n6972_8799.n209 a_n6972_8799.t128 464.166
R15321 a_n6972_8799.n208 a_n6972_8799.t92 464.166
R15322 a_n6972_8799.n197 a_n6972_8799.t72 464.166
R15323 a_n6972_8799.n207 a_n6972_8799.t36 464.166
R15324 a_n6972_8799.n206 a_n6972_8799.t105 464.166
R15325 a_n6972_8799.n198 a_n6972_8799.t104 464.166
R15326 a_n6972_8799.n205 a_n6972_8799.t49 464.166
R15327 a_n6972_8799.n204 a_n6972_8799.t108 464.166
R15328 a_n6972_8799.n199 a_n6972_8799.t107 464.166
R15329 a_n6972_8799.n203 a_n6972_8799.t53 464.166
R15330 a_n6972_8799.n202 a_n6972_8799.t52 464.166
R15331 a_n6972_8799.n200 a_n6972_8799.t123 464.166
R15332 a_n6972_8799.n228 a_n6972_8799.t130 464.166
R15333 a_n6972_8799.n227 a_n6972_8799.t51 464.166
R15334 a_n6972_8799.n213 a_n6972_8799.t90 464.166
R15335 a_n6972_8799.n226 a_n6972_8799.t38 464.166
R15336 a_n6972_8799.n225 a_n6972_8799.t110 464.166
R15337 a_n6972_8799.n214 a_n6972_8799.t62 464.166
R15338 a_n6972_8799.n224 a_n6972_8799.t96 464.166
R15339 a_n6972_8799.n223 a_n6972_8799.t43 464.166
R15340 a_n6972_8799.n215 a_n6972_8799.t66 464.166
R15341 a_n6972_8799.n222 a_n6972_8799.t126 464.166
R15342 a_n6972_8799.n221 a_n6972_8799.t102 464.166
R15343 a_n6972_8799.n216 a_n6972_8799.t122 464.166
R15344 a_n6972_8799.n220 a_n6972_8799.t89 464.166
R15345 a_n6972_8799.n219 a_n6972_8799.t106 464.166
R15346 a_n6972_8799.n217 a_n6972_8799.t56 464.166
R15347 a_n6972_8799.n133 a_n6972_8799.t78 464.166
R15348 a_n6972_8799.n136 a_n6972_8799.t77 464.166
R15349 a_n6972_8799.n132 a_n6972_8799.t101 464.166
R15350 a_n6972_8799.n137 a_n6972_8799.t68 464.166
R15351 a_n6972_8799.n138 a_n6972_8799.t69 464.166
R15352 a_n6972_8799.n139 a_n6972_8799.t100 464.166
R15353 a_n6972_8799.n140 a_n6972_8799.t37 464.166
R15354 a_n6972_8799.n131 a_n6972_8799.t65 464.166
R15355 a_n6972_8799.n141 a_n6972_8799.t83 464.166
R15356 a_n6972_8799.n142 a_n6972_8799.t117 464.166
R15357 a_n6972_8799.n143 a_n6972_8799.t47 464.166
R15358 a_n6972_8799.n144 a_n6972_8799.t64 464.166
R15359 a_n6972_8799.n130 a_n6972_8799.t114 464.166
R15360 a_n6972_8799.n145 a_n6972_8799.t46 464.166
R15361 a_n6972_8799.n149 a_n6972_8799.t84 464.166
R15362 a_n6972_8799.n152 a_n6972_8799.t85 464.166
R15363 a_n6972_8799.n148 a_n6972_8799.t113 464.166
R15364 a_n6972_8799.n153 a_n6972_8799.t75 464.166
R15365 a_n6972_8799.n154 a_n6972_8799.t76 464.166
R15366 a_n6972_8799.n155 a_n6972_8799.t109 464.166
R15367 a_n6972_8799.n156 a_n6972_8799.t48 464.166
R15368 a_n6972_8799.n147 a_n6972_8799.t74 464.166
R15369 a_n6972_8799.n157 a_n6972_8799.t94 464.166
R15370 a_n6972_8799.n158 a_n6972_8799.t129 464.166
R15371 a_n6972_8799.n159 a_n6972_8799.t61 464.166
R15372 a_n6972_8799.n160 a_n6972_8799.t73 464.166
R15373 a_n6972_8799.n146 a_n6972_8799.t124 464.166
R15374 a_n6972_8799.n161 a_n6972_8799.t55 464.166
R15375 a_n6972_8799.n166 a_n6972_8799.t54 464.166
R15376 a_n6972_8799.n169 a_n6972_8799.t39 464.166
R15377 a_n6972_8799.n165 a_n6972_8799.t88 464.166
R15378 a_n6972_8799.n170 a_n6972_8799.t121 464.166
R15379 a_n6972_8799.n171 a_n6972_8799.t103 464.166
R15380 a_n6972_8799.n172 a_n6972_8799.t127 464.166
R15381 a_n6972_8799.n173 a_n6972_8799.t82 464.166
R15382 a_n6972_8799.n164 a_n6972_8799.t44 464.166
R15383 a_n6972_8799.n174 a_n6972_8799.t97 464.166
R15384 a_n6972_8799.n175 a_n6972_8799.t60 464.166
R15385 a_n6972_8799.n176 a_n6972_8799.t111 464.166
R15386 a_n6972_8799.n177 a_n6972_8799.t67 464.166
R15387 a_n6972_8799.n163 a_n6972_8799.t91 464.166
R15388 a_n6972_8799.n178 a_n6972_8799.t50 464.166
R15389 a_n6972_8799.n52 a_n6972_8799.n30 74.4178
R15390 a_n6972_8799.n186 a_n6972_8799.n52 12.4674
R15391 a_n6972_8799.n51 a_n6972_8799.n30 80.107
R15392 a_n6972_8799.n51 a_n6972_8799.n187 1.08907
R15393 a_n6972_8799.n31 a_n6972_8799.n50 75.3623
R15394 a_n6972_8799.n49 a_n6972_8799.n31 70.3058
R15395 a_n6972_8799.n33 a_n6972_8799.n48 70.1674
R15396 a_n6972_8799.n48 a_n6972_8799.n182 20.9683
R15397 a_n6972_8799.n47 a_n6972_8799.n33 75.0448
R15398 a_n6972_8799.n190 a_n6972_8799.n47 11.2134
R15399 a_n6972_8799.n46 a_n6972_8799.n32 80.4688
R15400 a_n6972_8799.n32 a_n6972_8799.n45 74.73
R15401 a_n6972_8799.n44 a_n6972_8799.n34 70.1674
R15402 a_n6972_8799.n193 a_n6972_8799.n44 20.9683
R15403 a_n6972_8799.n34 a_n6972_8799.n43 70.5844
R15404 a_n6972_8799.n43 a_n6972_8799.n180 20.1342
R15405 a_n6972_8799.n42 a_n6972_8799.n35 75.6825
R15406 a_n6972_8799.n194 a_n6972_8799.n42 9.93802
R15407 a_n6972_8799.n35 a_n6972_8799.n195 161.3
R15408 a_n6972_8799.n63 a_n6972_8799.n24 74.4178
R15409 a_n6972_8799.n202 a_n6972_8799.n63 12.4674
R15410 a_n6972_8799.n62 a_n6972_8799.n24 80.107
R15411 a_n6972_8799.n62 a_n6972_8799.n203 1.08907
R15412 a_n6972_8799.n25 a_n6972_8799.n61 75.3623
R15413 a_n6972_8799.n60 a_n6972_8799.n25 70.3058
R15414 a_n6972_8799.n27 a_n6972_8799.n59 70.1674
R15415 a_n6972_8799.n59 a_n6972_8799.n198 20.9683
R15416 a_n6972_8799.n58 a_n6972_8799.n27 75.0448
R15417 a_n6972_8799.n206 a_n6972_8799.n58 11.2134
R15418 a_n6972_8799.n57 a_n6972_8799.n26 80.4688
R15419 a_n6972_8799.n26 a_n6972_8799.n56 74.73
R15420 a_n6972_8799.n55 a_n6972_8799.n28 70.1674
R15421 a_n6972_8799.n209 a_n6972_8799.n55 20.9683
R15422 a_n6972_8799.n28 a_n6972_8799.n54 70.5844
R15423 a_n6972_8799.n54 a_n6972_8799.n196 20.1342
R15424 a_n6972_8799.n53 a_n6972_8799.n29 75.6825
R15425 a_n6972_8799.n210 a_n6972_8799.n53 9.93802
R15426 a_n6972_8799.n29 a_n6972_8799.n211 161.3
R15427 a_n6972_8799.n74 a_n6972_8799.n18 74.4178
R15428 a_n6972_8799.n219 a_n6972_8799.n74 12.4674
R15429 a_n6972_8799.n73 a_n6972_8799.n18 80.107
R15430 a_n6972_8799.n73 a_n6972_8799.n220 1.08907
R15431 a_n6972_8799.n19 a_n6972_8799.n72 75.3623
R15432 a_n6972_8799.n71 a_n6972_8799.n19 70.3058
R15433 a_n6972_8799.n21 a_n6972_8799.n70 70.1674
R15434 a_n6972_8799.n70 a_n6972_8799.n215 20.9683
R15435 a_n6972_8799.n69 a_n6972_8799.n21 75.0448
R15436 a_n6972_8799.n223 a_n6972_8799.n69 11.2134
R15437 a_n6972_8799.n68 a_n6972_8799.n20 80.4688
R15438 a_n6972_8799.n20 a_n6972_8799.n67 74.73
R15439 a_n6972_8799.n66 a_n6972_8799.n22 70.1674
R15440 a_n6972_8799.n226 a_n6972_8799.n66 20.9683
R15441 a_n6972_8799.n22 a_n6972_8799.n65 70.5844
R15442 a_n6972_8799.n65 a_n6972_8799.n213 20.1342
R15443 a_n6972_8799.n64 a_n6972_8799.n23 75.6825
R15444 a_n6972_8799.n227 a_n6972_8799.n64 9.93802
R15445 a_n6972_8799.n23 a_n6972_8799.n228 161.3
R15446 a_n6972_8799.n13 a_n6972_8799.n85 70.1674
R15447 a_n6972_8799.n145 a_n6972_8799.n85 20.9683
R15448 a_n6972_8799.n84 a_n6972_8799.n13 74.4178
R15449 a_n6972_8799.n84 a_n6972_8799.n130 12.4674
R15450 a_n6972_8799.n12 a_n6972_8799.n83 80.107
R15451 a_n6972_8799.n144 a_n6972_8799.n83 1.08907
R15452 a_n6972_8799.n82 a_n6972_8799.n12 75.3623
R15453 a_n6972_8799.n14 a_n6972_8799.n81 70.3058
R15454 a_n6972_8799.n80 a_n6972_8799.n14 70.1674
R15455 a_n6972_8799.n80 a_n6972_8799.n131 20.9683
R15456 a_n6972_8799.n15 a_n6972_8799.n79 75.0448
R15457 a_n6972_8799.n140 a_n6972_8799.n79 11.2134
R15458 a_n6972_8799.n78 a_n6972_8799.n15 80.4688
R15459 a_n6972_8799.n16 a_n6972_8799.n77 74.73
R15460 a_n6972_8799.n76 a_n6972_8799.n16 70.1674
R15461 a_n6972_8799.n76 a_n6972_8799.n132 20.9683
R15462 a_n6972_8799.n17 a_n6972_8799.n75 70.5844
R15463 a_n6972_8799.n136 a_n6972_8799.n75 20.1342
R15464 a_n6972_8799.n135 a_n6972_8799.n17 161.3
R15465 a_n6972_8799.n7 a_n6972_8799.n96 70.1674
R15466 a_n6972_8799.n161 a_n6972_8799.n96 20.9683
R15467 a_n6972_8799.n95 a_n6972_8799.n7 74.4178
R15468 a_n6972_8799.n95 a_n6972_8799.n146 12.4674
R15469 a_n6972_8799.n6 a_n6972_8799.n94 80.107
R15470 a_n6972_8799.n160 a_n6972_8799.n94 1.08907
R15471 a_n6972_8799.n93 a_n6972_8799.n6 75.3623
R15472 a_n6972_8799.n8 a_n6972_8799.n92 70.3058
R15473 a_n6972_8799.n91 a_n6972_8799.n8 70.1674
R15474 a_n6972_8799.n91 a_n6972_8799.n147 20.9683
R15475 a_n6972_8799.n9 a_n6972_8799.n90 75.0448
R15476 a_n6972_8799.n156 a_n6972_8799.n90 11.2134
R15477 a_n6972_8799.n89 a_n6972_8799.n9 80.4688
R15478 a_n6972_8799.n10 a_n6972_8799.n88 74.73
R15479 a_n6972_8799.n87 a_n6972_8799.n10 70.1674
R15480 a_n6972_8799.n87 a_n6972_8799.n148 20.9683
R15481 a_n6972_8799.n11 a_n6972_8799.n86 70.5844
R15482 a_n6972_8799.n152 a_n6972_8799.n86 20.1342
R15483 a_n6972_8799.n151 a_n6972_8799.n11 161.3
R15484 a_n6972_8799.n1 a_n6972_8799.n107 70.1674
R15485 a_n6972_8799.n178 a_n6972_8799.n107 20.9683
R15486 a_n6972_8799.n106 a_n6972_8799.n1 74.4178
R15487 a_n6972_8799.n106 a_n6972_8799.n163 12.4674
R15488 a_n6972_8799.n0 a_n6972_8799.n105 80.107
R15489 a_n6972_8799.n177 a_n6972_8799.n105 1.08907
R15490 a_n6972_8799.n104 a_n6972_8799.n0 75.3623
R15491 a_n6972_8799.n2 a_n6972_8799.n103 70.3058
R15492 a_n6972_8799.n102 a_n6972_8799.n2 70.1674
R15493 a_n6972_8799.n102 a_n6972_8799.n164 20.9683
R15494 a_n6972_8799.n3 a_n6972_8799.n101 75.0448
R15495 a_n6972_8799.n173 a_n6972_8799.n101 11.2134
R15496 a_n6972_8799.n100 a_n6972_8799.n3 80.4688
R15497 a_n6972_8799.n4 a_n6972_8799.n99 74.73
R15498 a_n6972_8799.n98 a_n6972_8799.n4 70.1674
R15499 a_n6972_8799.n98 a_n6972_8799.n165 20.9683
R15500 a_n6972_8799.n5 a_n6972_8799.n97 70.5844
R15501 a_n6972_8799.n169 a_n6972_8799.n97 20.1342
R15502 a_n6972_8799.n168 a_n6972_8799.n5 161.3
R15503 a_n6972_8799.n37 a_n6972_8799.n108 98.9633
R15504 a_n6972_8799.n36 a_n6972_8799.n110 98.9631
R15505 a_n6972_8799.n37 a_n6972_8799.n109 98.6055
R15506 a_n6972_8799.n36 a_n6972_8799.n111 98.6055
R15507 a_n6972_8799.n36 a_n6972_8799.n112 98.6055
R15508 a_n6972_8799.n233 a_n6972_8799.n37 98.6054
R15509 a_n6972_8799.n115 a_n6972_8799.n113 81.4626
R15510 a_n6972_8799.n123 a_n6972_8799.n121 81.4626
R15511 a_n6972_8799.n119 a_n6972_8799.n117 81.4626
R15512 a_n6972_8799.n126 a_n6972_8799.n125 80.9324
R15513 a_n6972_8799.n128 a_n6972_8799.n127 80.9324
R15514 a_n6972_8799.n41 a_n6972_8799.n129 80.9324
R15515 a_n6972_8799.n40 a_n6972_8799.n116 80.9324
R15516 a_n6972_8799.n115 a_n6972_8799.n114 80.9324
R15517 a_n6972_8799.n123 a_n6972_8799.n122 80.9324
R15518 a_n6972_8799.n39 a_n6972_8799.n124 80.9324
R15519 a_n6972_8799.n38 a_n6972_8799.n120 80.9324
R15520 a_n6972_8799.n119 a_n6972_8799.n118 80.9324
R15521 a_n6972_8799.n30 a_n6972_8799.n185 70.4033
R15522 a_n6972_8799.n24 a_n6972_8799.n201 70.4033
R15523 a_n6972_8799.n18 a_n6972_8799.n218 70.4033
R15524 a_n6972_8799.n17 a_n6972_8799.n134 70.4033
R15525 a_n6972_8799.n11 a_n6972_8799.n150 70.4033
R15526 a_n6972_8799.n5 a_n6972_8799.n167 70.4033
R15527 a_n6972_8799.n195 a_n6972_8799.n194 48.2005
R15528 a_n6972_8799.n44 a_n6972_8799.n192 20.9683
R15529 a_n6972_8799.n191 a_n6972_8799.n190 48.2005
R15530 a_n6972_8799.n189 a_n6972_8799.n48 20.9683
R15531 a_n6972_8799.n187 a_n6972_8799.n183 48.2005
R15532 a_n6972_8799.n211 a_n6972_8799.n210 48.2005
R15533 a_n6972_8799.n55 a_n6972_8799.n208 20.9683
R15534 a_n6972_8799.n207 a_n6972_8799.n206 48.2005
R15535 a_n6972_8799.n205 a_n6972_8799.n59 20.9683
R15536 a_n6972_8799.n203 a_n6972_8799.n199 48.2005
R15537 a_n6972_8799.n228 a_n6972_8799.n227 48.2005
R15538 a_n6972_8799.n66 a_n6972_8799.n225 20.9683
R15539 a_n6972_8799.n224 a_n6972_8799.n223 48.2005
R15540 a_n6972_8799.n222 a_n6972_8799.n70 20.9683
R15541 a_n6972_8799.n220 a_n6972_8799.n216 48.2005
R15542 a_n6972_8799.n137 a_n6972_8799.n76 20.9683
R15543 a_n6972_8799.n140 a_n6972_8799.n139 48.2005
R15544 a_n6972_8799.n141 a_n6972_8799.n80 20.9683
R15545 a_n6972_8799.n144 a_n6972_8799.n143 48.2005
R15546 a_n6972_8799.t45 a_n6972_8799.n85 485.135
R15547 a_n6972_8799.n153 a_n6972_8799.n87 20.9683
R15548 a_n6972_8799.n156 a_n6972_8799.n155 48.2005
R15549 a_n6972_8799.n157 a_n6972_8799.n91 20.9683
R15550 a_n6972_8799.n160 a_n6972_8799.n159 48.2005
R15551 a_n6972_8799.t59 a_n6972_8799.n96 485.135
R15552 a_n6972_8799.n170 a_n6972_8799.n98 20.9683
R15553 a_n6972_8799.n173 a_n6972_8799.n172 48.2005
R15554 a_n6972_8799.n174 a_n6972_8799.n102 20.9683
R15555 a_n6972_8799.n177 a_n6972_8799.n176 48.2005
R15556 a_n6972_8799.t131 a_n6972_8799.n107 485.135
R15557 a_n6972_8799.n46 a_n6972_8799.n181 47.835
R15558 a_n6972_8799.n49 a_n6972_8799.n188 20.6913
R15559 a_n6972_8799.n57 a_n6972_8799.n197 47.835
R15560 a_n6972_8799.n60 a_n6972_8799.n204 20.6913
R15561 a_n6972_8799.n68 a_n6972_8799.n214 47.835
R15562 a_n6972_8799.n71 a_n6972_8799.n221 20.6913
R15563 a_n6972_8799.n138 a_n6972_8799.n78 47.835
R15564 a_n6972_8799.n142 a_n6972_8799.n81 20.6913
R15565 a_n6972_8799.n154 a_n6972_8799.n89 47.835
R15566 a_n6972_8799.n158 a_n6972_8799.n92 20.6913
R15567 a_n6972_8799.n171 a_n6972_8799.n100 47.835
R15568 a_n6972_8799.n175 a_n6972_8799.n103 20.6913
R15569 a_n6972_8799.n193 a_n6972_8799.n43 22.3251
R15570 a_n6972_8799.n209 a_n6972_8799.n54 22.3251
R15571 a_n6972_8799.n226 a_n6972_8799.n65 22.3251
R15572 a_n6972_8799.n132 a_n6972_8799.n75 22.3251
R15573 a_n6972_8799.n148 a_n6972_8799.n86 22.3251
R15574 a_n6972_8799.n165 a_n6972_8799.n97 22.3251
R15575 a_n6972_8799.n126 a_n6972_8799.n39 34.3237
R15576 a_n6972_8799.n52 a_n6972_8799.n184 33.6462
R15577 a_n6972_8799.n63 a_n6972_8799.n200 33.6462
R15578 a_n6972_8799.n74 a_n6972_8799.n217 33.6462
R15579 a_n6972_8799.n136 a_n6972_8799.n135 27.0217
R15580 a_n6972_8799.n145 a_n6972_8799.n84 33.6462
R15581 a_n6972_8799.n152 a_n6972_8799.n151 27.0217
R15582 a_n6972_8799.n161 a_n6972_8799.n95 33.6462
R15583 a_n6972_8799.n169 a_n6972_8799.n168 27.0217
R15584 a_n6972_8799.n178 a_n6972_8799.n106 33.6462
R15585 a_n6972_8799.n45 a_n6972_8799.n181 11.843
R15586 a_n6972_8799.n188 a_n6972_8799.n50 36.139
R15587 a_n6972_8799.n56 a_n6972_8799.n197 11.843
R15588 a_n6972_8799.n204 a_n6972_8799.n61 36.139
R15589 a_n6972_8799.n67 a_n6972_8799.n214 11.843
R15590 a_n6972_8799.n221 a_n6972_8799.n72 36.139
R15591 a_n6972_8799.n138 a_n6972_8799.n77 11.843
R15592 a_n6972_8799.n142 a_n6972_8799.n82 36.139
R15593 a_n6972_8799.n154 a_n6972_8799.n88 11.843
R15594 a_n6972_8799.n158 a_n6972_8799.n93 36.139
R15595 a_n6972_8799.n171 a_n6972_8799.n99 11.843
R15596 a_n6972_8799.n175 a_n6972_8799.n104 36.139
R15597 a_n6972_8799.n47 a_n6972_8799.n182 35.3134
R15598 a_n6972_8799.n58 a_n6972_8799.n198 35.3134
R15599 a_n6972_8799.n69 a_n6972_8799.n215 35.3134
R15600 a_n6972_8799.n131 a_n6972_8799.n79 35.3134
R15601 a_n6972_8799.n147 a_n6972_8799.n90 35.3134
R15602 a_n6972_8799.n164 a_n6972_8799.n101 35.3134
R15603 a_n6972_8799.n192 a_n6972_8799.n45 34.4824
R15604 a_n6972_8799.n50 a_n6972_8799.n183 10.5784
R15605 a_n6972_8799.n208 a_n6972_8799.n56 34.4824
R15606 a_n6972_8799.n61 a_n6972_8799.n199 10.5784
R15607 a_n6972_8799.n225 a_n6972_8799.n67 34.4824
R15608 a_n6972_8799.n72 a_n6972_8799.n216 10.5784
R15609 a_n6972_8799.n77 a_n6972_8799.n137 34.4824
R15610 a_n6972_8799.n143 a_n6972_8799.n82 10.5784
R15611 a_n6972_8799.n88 a_n6972_8799.n153 34.4824
R15612 a_n6972_8799.n159 a_n6972_8799.n93 10.5784
R15613 a_n6972_8799.n99 a_n6972_8799.n170 34.4824
R15614 a_n6972_8799.n176 a_n6972_8799.n104 10.5784
R15615 a_n6972_8799.n42 a_n6972_8799.n180 36.9592
R15616 a_n6972_8799.n53 a_n6972_8799.n196 36.9592
R15617 a_n6972_8799.n64 a_n6972_8799.n213 36.9592
R15618 a_n6972_8799.n135 a_n6972_8799.n133 21.1793
R15619 a_n6972_8799.n151 a_n6972_8799.n149 21.1793
R15620 a_n6972_8799.n168 a_n6972_8799.n166 21.1793
R15621 a_n6972_8799.n185 a_n6972_8799.n184 20.9576
R15622 a_n6972_8799.n201 a_n6972_8799.n200 20.9576
R15623 a_n6972_8799.n218 a_n6972_8799.n217 20.9576
R15624 a_n6972_8799.n134 a_n6972_8799.n133 20.9576
R15625 a_n6972_8799.n150 a_n6972_8799.n149 20.9576
R15626 a_n6972_8799.n167 a_n6972_8799.n166 20.9576
R15627 a_n6972_8799.n231 a_n6972_8799.n41 12.3339
R15628 a_n6972_8799.n232 a_n6972_8799.n231 11.4887
R15629 a_n6972_8799.n212 a_n6972_8799.n35 9.07815
R15630 a_n6972_8799.n162 a_n6972_8799.n13 9.07815
R15631 a_n6972_8799.n230 a_n6972_8799.n179 6.93972
R15632 a_n6972_8799.n230 a_n6972_8799.n229 6.44309
R15633 a_n6972_8799.n212 a_n6972_8799.n29 4.9702
R15634 a_n6972_8799.n229 a_n6972_8799.n23 4.9702
R15635 a_n6972_8799.n162 a_n6972_8799.n7 4.9702
R15636 a_n6972_8799.n179 a_n6972_8799.n1 4.9702
R15637 a_n6972_8799.n229 a_n6972_8799.n212 4.10845
R15638 a_n6972_8799.n179 a_n6972_8799.n162 4.10845
R15639 a_n6972_8799.n109 a_n6972_8799.t10 3.61217
R15640 a_n6972_8799.n109 a_n6972_8799.t5 3.61217
R15641 a_n6972_8799.n108 a_n6972_8799.t33 3.61217
R15642 a_n6972_8799.n108 a_n6972_8799.t34 3.61217
R15643 a_n6972_8799.n110 a_n6972_8799.t7 3.61217
R15644 a_n6972_8799.n110 a_n6972_8799.t9 3.61217
R15645 a_n6972_8799.n111 a_n6972_8799.t8 3.61217
R15646 a_n6972_8799.n111 a_n6972_8799.t2 3.61217
R15647 a_n6972_8799.n112 a_n6972_8799.t11 3.61217
R15648 a_n6972_8799.n112 a_n6972_8799.t12 3.61217
R15649 a_n6972_8799.t0 a_n6972_8799.n233 3.61217
R15650 a_n6972_8799.n233 a_n6972_8799.t4 3.61217
R15651 a_n6972_8799.n231 a_n6972_8799.n230 3.4105
R15652 a_n6972_8799.n125 a_n6972_8799.t35 2.82907
R15653 a_n6972_8799.n125 a_n6972_8799.t25 2.82907
R15654 a_n6972_8799.n127 a_n6972_8799.t19 2.82907
R15655 a_n6972_8799.n127 a_n6972_8799.t28 2.82907
R15656 a_n6972_8799.n129 a_n6972_8799.t30 2.82907
R15657 a_n6972_8799.n129 a_n6972_8799.t29 2.82907
R15658 a_n6972_8799.n116 a_n6972_8799.t20 2.82907
R15659 a_n6972_8799.n116 a_n6972_8799.t18 2.82907
R15660 a_n6972_8799.n114 a_n6972_8799.t1 2.82907
R15661 a_n6972_8799.n114 a_n6972_8799.t13 2.82907
R15662 a_n6972_8799.n113 a_n6972_8799.t22 2.82907
R15663 a_n6972_8799.n113 a_n6972_8799.t27 2.82907
R15664 a_n6972_8799.n121 a_n6972_8799.t16 2.82907
R15665 a_n6972_8799.n121 a_n6972_8799.t14 2.82907
R15666 a_n6972_8799.n122 a_n6972_8799.t32 2.82907
R15667 a_n6972_8799.n122 a_n6972_8799.t24 2.82907
R15668 a_n6972_8799.n124 a_n6972_8799.t31 2.82907
R15669 a_n6972_8799.n124 a_n6972_8799.t23 2.82907
R15670 a_n6972_8799.n120 a_n6972_8799.t17 2.82907
R15671 a_n6972_8799.n120 a_n6972_8799.t26 2.82907
R15672 a_n6972_8799.n118 a_n6972_8799.t6 2.82907
R15673 a_n6972_8799.n118 a_n6972_8799.t21 2.82907
R15674 a_n6972_8799.n117 a_n6972_8799.t15 2.82907
R15675 a_n6972_8799.n117 a_n6972_8799.t3 2.82907
R15676 a_n6972_8799.n51 a_n6972_8799.n186 47.0982
R15677 a_n6972_8799.n62 a_n6972_8799.n202 47.0982
R15678 a_n6972_8799.n73 a_n6972_8799.n219 47.0982
R15679 a_n6972_8799.n130 a_n6972_8799.n83 47.0982
R15680 a_n6972_8799.n146 a_n6972_8799.n94 47.0982
R15681 a_n6972_8799.n163 a_n6972_8799.n105 47.0982
R15682 a_n6972_8799.n232 a_n6972_8799.n36 31.5519
R15683 a_n6972_8799.n46 a_n6972_8799.n191 0.365327
R15684 a_n6972_8799.n189 a_n6972_8799.n49 21.4216
R15685 a_n6972_8799.n57 a_n6972_8799.n207 0.365327
R15686 a_n6972_8799.n205 a_n6972_8799.n60 21.4216
R15687 a_n6972_8799.n68 a_n6972_8799.n224 0.365327
R15688 a_n6972_8799.n222 a_n6972_8799.n71 21.4216
R15689 a_n6972_8799.n139 a_n6972_8799.n78 0.365327
R15690 a_n6972_8799.n81 a_n6972_8799.n141 21.4216
R15691 a_n6972_8799.n155 a_n6972_8799.n89 0.365327
R15692 a_n6972_8799.n92 a_n6972_8799.n157 21.4216
R15693 a_n6972_8799.n172 a_n6972_8799.n100 0.365327
R15694 a_n6972_8799.n103 a_n6972_8799.n174 21.4216
R15695 a_n6972_8799.n37 a_n6972_8799.n232 17.6132
R15696 a_n6972_8799.n31 a_n6972_8799.n30 1.13686
R15697 a_n6972_8799.n25 a_n6972_8799.n24 1.13686
R15698 a_n6972_8799.n19 a_n6972_8799.n18 1.13686
R15699 a_n6972_8799.n13 a_n6972_8799.n12 1.13686
R15700 a_n6972_8799.n7 a_n6972_8799.n6 1.13686
R15701 a_n6972_8799.n1 a_n6972_8799.n0 1.13686
R15702 a_n6972_8799.n35 a_n6972_8799.n34 0.758076
R15703 a_n6972_8799.n32 a_n6972_8799.n34 0.758076
R15704 a_n6972_8799.n33 a_n6972_8799.n32 0.758076
R15705 a_n6972_8799.n33 a_n6972_8799.n31 0.758076
R15706 a_n6972_8799.n29 a_n6972_8799.n28 0.758076
R15707 a_n6972_8799.n26 a_n6972_8799.n28 0.758076
R15708 a_n6972_8799.n27 a_n6972_8799.n26 0.758076
R15709 a_n6972_8799.n27 a_n6972_8799.n25 0.758076
R15710 a_n6972_8799.n23 a_n6972_8799.n22 0.758076
R15711 a_n6972_8799.n20 a_n6972_8799.n22 0.758076
R15712 a_n6972_8799.n21 a_n6972_8799.n20 0.758076
R15713 a_n6972_8799.n21 a_n6972_8799.n19 0.758076
R15714 a_n6972_8799.n16 a_n6972_8799.n17 0.758076
R15715 a_n6972_8799.n15 a_n6972_8799.n16 0.758076
R15716 a_n6972_8799.n14 a_n6972_8799.n15 0.758076
R15717 a_n6972_8799.n12 a_n6972_8799.n14 0.758076
R15718 a_n6972_8799.n10 a_n6972_8799.n11 0.758076
R15719 a_n6972_8799.n9 a_n6972_8799.n10 0.758076
R15720 a_n6972_8799.n8 a_n6972_8799.n9 0.758076
R15721 a_n6972_8799.n6 a_n6972_8799.n8 0.758076
R15722 a_n6972_8799.n4 a_n6972_8799.n5 0.758076
R15723 a_n6972_8799.n3 a_n6972_8799.n4 0.758076
R15724 a_n6972_8799.n2 a_n6972_8799.n3 0.758076
R15725 a_n6972_8799.n0 a_n6972_8799.n2 0.758076
R15726 a_n6972_8799.n38 a_n6972_8799.n119 0.530672
R15727 a_n6972_8799.n39 a_n6972_8799.n123 0.530672
R15728 a_n6972_8799.n40 a_n6972_8799.n115 0.530672
R15729 a_n6972_8799.n41 a_n6972_8799.n128 0.530672
R15730 a_n6972_8799.n128 a_n6972_8799.n126 0.530672
R15731 a_n6972_8799.n41 a_n6972_8799.n40 0.530672
R15732 a_n6972_8799.n39 a_n6972_8799.n38 0.530672
R15733 vdd.n315 vdd.n279 756.745
R15734 vdd.n260 vdd.n224 756.745
R15735 vdd.n217 vdd.n181 756.745
R15736 vdd.n162 vdd.n126 756.745
R15737 vdd.n120 vdd.n84 756.745
R15738 vdd.n65 vdd.n29 756.745
R15739 vdd.n1684 vdd.n1648 756.745
R15740 vdd.n1739 vdd.n1703 756.745
R15741 vdd.n1586 vdd.n1550 756.745
R15742 vdd.n1641 vdd.n1605 756.745
R15743 vdd.n1489 vdd.n1453 756.745
R15744 vdd.n1544 vdd.n1508 756.745
R15745 vdd.n2094 vdd.t214 640.208
R15746 vdd.n936 vdd.t199 640.208
R15747 vdd.n2068 vdd.t237 640.208
R15748 vdd.n928 vdd.t225 640.208
R15749 vdd.n2839 vdd.t186 640.208
R15750 vdd.n2559 vdd.t222 640.208
R15751 vdd.n804 vdd.t203 640.208
R15752 vdd.n2556 vdd.t207 640.208
R15753 vdd.n768 vdd.t211 640.208
R15754 vdd.n998 vdd.t218 640.208
R15755 vdd.n1148 vdd.t168 592.009
R15756 vdd.n1304 vdd.t183 592.009
R15757 vdd.n1340 vdd.t190 592.009
R15758 vdd.n2250 vdd.t179 592.009
R15759 vdd.n1887 vdd.t193 592.009
R15760 vdd.n1847 vdd.t196 592.009
R15761 vdd.n405 vdd.t172 592.009
R15762 vdd.n419 vdd.t228 592.009
R15763 vdd.n431 vdd.t234 592.009
R15764 vdd.n723 vdd.t164 592.009
R15765 vdd.n686 vdd.t176 592.009
R15766 vdd.n3013 vdd.t231 592.009
R15767 vdd.n316 vdd.n315 585
R15768 vdd.n314 vdd.n281 585
R15769 vdd.n313 vdd.n312 585
R15770 vdd.n284 vdd.n282 585
R15771 vdd.n307 vdd.n306 585
R15772 vdd.n305 vdd.n304 585
R15773 vdd.n288 vdd.n287 585
R15774 vdd.n299 vdd.n298 585
R15775 vdd.n297 vdd.n296 585
R15776 vdd.n292 vdd.n291 585
R15777 vdd.n261 vdd.n260 585
R15778 vdd.n259 vdd.n226 585
R15779 vdd.n258 vdd.n257 585
R15780 vdd.n229 vdd.n227 585
R15781 vdd.n252 vdd.n251 585
R15782 vdd.n250 vdd.n249 585
R15783 vdd.n233 vdd.n232 585
R15784 vdd.n244 vdd.n243 585
R15785 vdd.n242 vdd.n241 585
R15786 vdd.n237 vdd.n236 585
R15787 vdd.n218 vdd.n217 585
R15788 vdd.n216 vdd.n183 585
R15789 vdd.n215 vdd.n214 585
R15790 vdd.n186 vdd.n184 585
R15791 vdd.n209 vdd.n208 585
R15792 vdd.n207 vdd.n206 585
R15793 vdd.n190 vdd.n189 585
R15794 vdd.n201 vdd.n200 585
R15795 vdd.n199 vdd.n198 585
R15796 vdd.n194 vdd.n193 585
R15797 vdd.n163 vdd.n162 585
R15798 vdd.n161 vdd.n128 585
R15799 vdd.n160 vdd.n159 585
R15800 vdd.n131 vdd.n129 585
R15801 vdd.n154 vdd.n153 585
R15802 vdd.n152 vdd.n151 585
R15803 vdd.n135 vdd.n134 585
R15804 vdd.n146 vdd.n145 585
R15805 vdd.n144 vdd.n143 585
R15806 vdd.n139 vdd.n138 585
R15807 vdd.n121 vdd.n120 585
R15808 vdd.n119 vdd.n86 585
R15809 vdd.n118 vdd.n117 585
R15810 vdd.n89 vdd.n87 585
R15811 vdd.n112 vdd.n111 585
R15812 vdd.n110 vdd.n109 585
R15813 vdd.n93 vdd.n92 585
R15814 vdd.n104 vdd.n103 585
R15815 vdd.n102 vdd.n101 585
R15816 vdd.n97 vdd.n96 585
R15817 vdd.n66 vdd.n65 585
R15818 vdd.n64 vdd.n31 585
R15819 vdd.n63 vdd.n62 585
R15820 vdd.n34 vdd.n32 585
R15821 vdd.n57 vdd.n56 585
R15822 vdd.n55 vdd.n54 585
R15823 vdd.n38 vdd.n37 585
R15824 vdd.n49 vdd.n48 585
R15825 vdd.n47 vdd.n46 585
R15826 vdd.n42 vdd.n41 585
R15827 vdd.n1685 vdd.n1684 585
R15828 vdd.n1683 vdd.n1650 585
R15829 vdd.n1682 vdd.n1681 585
R15830 vdd.n1653 vdd.n1651 585
R15831 vdd.n1676 vdd.n1675 585
R15832 vdd.n1674 vdd.n1673 585
R15833 vdd.n1657 vdd.n1656 585
R15834 vdd.n1668 vdd.n1667 585
R15835 vdd.n1666 vdd.n1665 585
R15836 vdd.n1661 vdd.n1660 585
R15837 vdd.n1740 vdd.n1739 585
R15838 vdd.n1738 vdd.n1705 585
R15839 vdd.n1737 vdd.n1736 585
R15840 vdd.n1708 vdd.n1706 585
R15841 vdd.n1731 vdd.n1730 585
R15842 vdd.n1729 vdd.n1728 585
R15843 vdd.n1712 vdd.n1711 585
R15844 vdd.n1723 vdd.n1722 585
R15845 vdd.n1721 vdd.n1720 585
R15846 vdd.n1716 vdd.n1715 585
R15847 vdd.n1587 vdd.n1586 585
R15848 vdd.n1585 vdd.n1552 585
R15849 vdd.n1584 vdd.n1583 585
R15850 vdd.n1555 vdd.n1553 585
R15851 vdd.n1578 vdd.n1577 585
R15852 vdd.n1576 vdd.n1575 585
R15853 vdd.n1559 vdd.n1558 585
R15854 vdd.n1570 vdd.n1569 585
R15855 vdd.n1568 vdd.n1567 585
R15856 vdd.n1563 vdd.n1562 585
R15857 vdd.n1642 vdd.n1641 585
R15858 vdd.n1640 vdd.n1607 585
R15859 vdd.n1639 vdd.n1638 585
R15860 vdd.n1610 vdd.n1608 585
R15861 vdd.n1633 vdd.n1632 585
R15862 vdd.n1631 vdd.n1630 585
R15863 vdd.n1614 vdd.n1613 585
R15864 vdd.n1625 vdd.n1624 585
R15865 vdd.n1623 vdd.n1622 585
R15866 vdd.n1618 vdd.n1617 585
R15867 vdd.n1490 vdd.n1489 585
R15868 vdd.n1488 vdd.n1455 585
R15869 vdd.n1487 vdd.n1486 585
R15870 vdd.n1458 vdd.n1456 585
R15871 vdd.n1481 vdd.n1480 585
R15872 vdd.n1479 vdd.n1478 585
R15873 vdd.n1462 vdd.n1461 585
R15874 vdd.n1473 vdd.n1472 585
R15875 vdd.n1471 vdd.n1470 585
R15876 vdd.n1466 vdd.n1465 585
R15877 vdd.n1545 vdd.n1544 585
R15878 vdd.n1543 vdd.n1510 585
R15879 vdd.n1542 vdd.n1541 585
R15880 vdd.n1513 vdd.n1511 585
R15881 vdd.n1536 vdd.n1535 585
R15882 vdd.n1534 vdd.n1533 585
R15883 vdd.n1517 vdd.n1516 585
R15884 vdd.n1528 vdd.n1527 585
R15885 vdd.n1526 vdd.n1525 585
R15886 vdd.n1521 vdd.n1520 585
R15887 vdd.n445 vdd.n370 462.44
R15888 vdd.n3251 vdd.n372 462.44
R15889 vdd.n3146 vdd.n657 462.44
R15890 vdd.n3144 vdd.n660 462.44
R15891 vdd.n2245 vdd.n1047 462.44
R15892 vdd.n2248 vdd.n2247 462.44
R15893 vdd.n1375 vdd.n1145 462.44
R15894 vdd.n1372 vdd.n1143 462.44
R15895 vdd.n293 vdd.t124 329.043
R15896 vdd.n238 vdd.t98 329.043
R15897 vdd.n195 vdd.t110 329.043
R15898 vdd.n140 vdd.t87 329.043
R15899 vdd.n98 vdd.t42 329.043
R15900 vdd.n43 vdd.t22 329.043
R15901 vdd.n1662 vdd.t137 329.043
R15902 vdd.n1717 vdd.t48 329.043
R15903 vdd.n1564 vdd.t122 329.043
R15904 vdd.n1619 vdd.t32 329.043
R15905 vdd.n1467 vdd.t20 329.043
R15906 vdd.n1522 vdd.t45 329.043
R15907 vdd.n1148 vdd.t171 319.788
R15908 vdd.n1304 vdd.t185 319.788
R15909 vdd.n1340 vdd.t192 319.788
R15910 vdd.n2250 vdd.t181 319.788
R15911 vdd.n1887 vdd.t194 319.788
R15912 vdd.n1847 vdd.t197 319.788
R15913 vdd.n405 vdd.t174 319.788
R15914 vdd.n419 vdd.t229 319.788
R15915 vdd.n431 vdd.t235 319.788
R15916 vdd.n723 vdd.t167 319.788
R15917 vdd.n686 vdd.t178 319.788
R15918 vdd.n3013 vdd.t233 319.788
R15919 vdd.n1149 vdd.t170 303.69
R15920 vdd.n1305 vdd.t184 303.69
R15921 vdd.n1341 vdd.t191 303.69
R15922 vdd.n2251 vdd.t182 303.69
R15923 vdd.n1888 vdd.t195 303.69
R15924 vdd.n1848 vdd.t198 303.69
R15925 vdd.n406 vdd.t175 303.69
R15926 vdd.n420 vdd.t230 303.69
R15927 vdd.n432 vdd.t236 303.69
R15928 vdd.n724 vdd.t166 303.69
R15929 vdd.n687 vdd.t177 303.69
R15930 vdd.n3014 vdd.t232 303.69
R15931 vdd.n2782 vdd.n884 297.074
R15932 vdd.n2975 vdd.n778 297.074
R15933 vdd.n2912 vdd.n775 297.074
R15934 vdd.n2705 vdd.n885 297.074
R15935 vdd.n2520 vdd.n925 297.074
R15936 vdd.n2451 vdd.n2450 297.074
R15937 vdd.n2197 vdd.n1021 297.074
R15938 vdd.n2293 vdd.n1019 297.074
R15939 vdd.n2891 vdd.n776 297.074
R15940 vdd.n2978 vdd.n2977 297.074
R15941 vdd.n2554 vdd.n886 297.074
R15942 vdd.n2780 vdd.n887 297.074
R15943 vdd.n2448 vdd.n934 297.074
R15944 vdd.n932 vdd.n907 297.074
R15945 vdd.n2134 vdd.n1022 297.074
R15946 vdd.n2291 vdd.n1023 297.074
R15947 vdd.n2893 vdd.n776 185
R15948 vdd.n2976 vdd.n776 185
R15949 vdd.n2895 vdd.n2894 185
R15950 vdd.n2894 vdd.n774 185
R15951 vdd.n2896 vdd.n810 185
R15952 vdd.n2906 vdd.n810 185
R15953 vdd.n2897 vdd.n819 185
R15954 vdd.n819 vdd.n817 185
R15955 vdd.n2899 vdd.n2898 185
R15956 vdd.n2900 vdd.n2899 185
R15957 vdd.n2852 vdd.n818 185
R15958 vdd.n818 vdd.n814 185
R15959 vdd.n2851 vdd.n2850 185
R15960 vdd.n2850 vdd.n2849 185
R15961 vdd.n821 vdd.n820 185
R15962 vdd.n822 vdd.n821 185
R15963 vdd.n2842 vdd.n2841 185
R15964 vdd.n2843 vdd.n2842 185
R15965 vdd.n2838 vdd.n831 185
R15966 vdd.n831 vdd.n828 185
R15967 vdd.n2837 vdd.n2836 185
R15968 vdd.n2836 vdd.n2835 185
R15969 vdd.n833 vdd.n832 185
R15970 vdd.n841 vdd.n833 185
R15971 vdd.n2828 vdd.n2827 185
R15972 vdd.n2829 vdd.n2828 185
R15973 vdd.n2826 vdd.n842 185
R15974 vdd.n2677 vdd.n842 185
R15975 vdd.n2825 vdd.n2824 185
R15976 vdd.n2824 vdd.n2823 185
R15977 vdd.n844 vdd.n843 185
R15978 vdd.n845 vdd.n844 185
R15979 vdd.n2816 vdd.n2815 185
R15980 vdd.n2817 vdd.n2816 185
R15981 vdd.n2814 vdd.n854 185
R15982 vdd.n854 vdd.n851 185
R15983 vdd.n2813 vdd.n2812 185
R15984 vdd.n2812 vdd.n2811 185
R15985 vdd.n856 vdd.n855 185
R15986 vdd.n864 vdd.n856 185
R15987 vdd.n2804 vdd.n2803 185
R15988 vdd.n2805 vdd.n2804 185
R15989 vdd.n2802 vdd.n865 185
R15990 vdd.n871 vdd.n865 185
R15991 vdd.n2801 vdd.n2800 185
R15992 vdd.n2800 vdd.n2799 185
R15993 vdd.n867 vdd.n866 185
R15994 vdd.n868 vdd.n867 185
R15995 vdd.n2792 vdd.n2791 185
R15996 vdd.n2793 vdd.n2792 185
R15997 vdd.n2790 vdd.n877 185
R15998 vdd.n2698 vdd.n877 185
R15999 vdd.n2789 vdd.n2788 185
R16000 vdd.n2788 vdd.n2787 185
R16001 vdd.n879 vdd.n878 185
R16002 vdd.t157 vdd.n879 185
R16003 vdd.n2780 vdd.n2779 185
R16004 vdd.n2781 vdd.n2780 185
R16005 vdd.n2778 vdd.n887 185
R16006 vdd.n2777 vdd.n2776 185
R16007 vdd.n889 vdd.n888 185
R16008 vdd.n2563 vdd.n2562 185
R16009 vdd.n2565 vdd.n2564 185
R16010 vdd.n2567 vdd.n2566 185
R16011 vdd.n2569 vdd.n2568 185
R16012 vdd.n2571 vdd.n2570 185
R16013 vdd.n2573 vdd.n2572 185
R16014 vdd.n2575 vdd.n2574 185
R16015 vdd.n2577 vdd.n2576 185
R16016 vdd.n2579 vdd.n2578 185
R16017 vdd.n2581 vdd.n2580 185
R16018 vdd.n2583 vdd.n2582 185
R16019 vdd.n2585 vdd.n2584 185
R16020 vdd.n2587 vdd.n2586 185
R16021 vdd.n2589 vdd.n2588 185
R16022 vdd.n2591 vdd.n2590 185
R16023 vdd.n2593 vdd.n2592 185
R16024 vdd.n2595 vdd.n2594 185
R16025 vdd.n2597 vdd.n2596 185
R16026 vdd.n2599 vdd.n2598 185
R16027 vdd.n2601 vdd.n2600 185
R16028 vdd.n2603 vdd.n2602 185
R16029 vdd.n2605 vdd.n2604 185
R16030 vdd.n2607 vdd.n2606 185
R16031 vdd.n2609 vdd.n2608 185
R16032 vdd.n2611 vdd.n2610 185
R16033 vdd.n2613 vdd.n2612 185
R16034 vdd.n2615 vdd.n2614 185
R16035 vdd.n2617 vdd.n2616 185
R16036 vdd.n2619 vdd.n2618 185
R16037 vdd.n2621 vdd.n2620 185
R16038 vdd.n2623 vdd.n2622 185
R16039 vdd.n2624 vdd.n2554 185
R16040 vdd.n2774 vdd.n2554 185
R16041 vdd.n2979 vdd.n2978 185
R16042 vdd.n2980 vdd.n767 185
R16043 vdd.n2982 vdd.n2981 185
R16044 vdd.n2984 vdd.n765 185
R16045 vdd.n2986 vdd.n2985 185
R16046 vdd.n2987 vdd.n764 185
R16047 vdd.n2989 vdd.n2988 185
R16048 vdd.n2991 vdd.n762 185
R16049 vdd.n2993 vdd.n2992 185
R16050 vdd.n2994 vdd.n761 185
R16051 vdd.n2996 vdd.n2995 185
R16052 vdd.n2998 vdd.n759 185
R16053 vdd.n3000 vdd.n2999 185
R16054 vdd.n3001 vdd.n758 185
R16055 vdd.n3003 vdd.n3002 185
R16056 vdd.n3005 vdd.n757 185
R16057 vdd.n3006 vdd.n754 185
R16058 vdd.n3009 vdd.n3008 185
R16059 vdd.n755 vdd.n753 185
R16060 vdd.n2865 vdd.n2864 185
R16061 vdd.n2867 vdd.n2866 185
R16062 vdd.n2869 vdd.n2861 185
R16063 vdd.n2871 vdd.n2870 185
R16064 vdd.n2872 vdd.n2860 185
R16065 vdd.n2874 vdd.n2873 185
R16066 vdd.n2876 vdd.n2858 185
R16067 vdd.n2878 vdd.n2877 185
R16068 vdd.n2879 vdd.n2857 185
R16069 vdd.n2881 vdd.n2880 185
R16070 vdd.n2883 vdd.n2855 185
R16071 vdd.n2885 vdd.n2884 185
R16072 vdd.n2886 vdd.n2854 185
R16073 vdd.n2888 vdd.n2887 185
R16074 vdd.n2890 vdd.n2853 185
R16075 vdd.n2892 vdd.n2891 185
R16076 vdd.n2891 vdd.n756 185
R16077 vdd.n2977 vdd.n771 185
R16078 vdd.n2977 vdd.n2976 185
R16079 vdd.n2629 vdd.n773 185
R16080 vdd.n774 vdd.n773 185
R16081 vdd.n2630 vdd.n809 185
R16082 vdd.n2906 vdd.n809 185
R16083 vdd.n2632 vdd.n2631 185
R16084 vdd.n2631 vdd.n817 185
R16085 vdd.n2633 vdd.n816 185
R16086 vdd.n2900 vdd.n816 185
R16087 vdd.n2635 vdd.n2634 185
R16088 vdd.n2634 vdd.n814 185
R16089 vdd.n2636 vdd.n824 185
R16090 vdd.n2849 vdd.n824 185
R16091 vdd.n2638 vdd.n2637 185
R16092 vdd.n2637 vdd.n822 185
R16093 vdd.n2639 vdd.n830 185
R16094 vdd.n2843 vdd.n830 185
R16095 vdd.n2641 vdd.n2640 185
R16096 vdd.n2640 vdd.n828 185
R16097 vdd.n2642 vdd.n835 185
R16098 vdd.n2835 vdd.n835 185
R16099 vdd.n2644 vdd.n2643 185
R16100 vdd.n2643 vdd.n841 185
R16101 vdd.n2645 vdd.n840 185
R16102 vdd.n2829 vdd.n840 185
R16103 vdd.n2679 vdd.n2678 185
R16104 vdd.n2678 vdd.n2677 185
R16105 vdd.n2680 vdd.n847 185
R16106 vdd.n2823 vdd.n847 185
R16107 vdd.n2682 vdd.n2681 185
R16108 vdd.n2681 vdd.n845 185
R16109 vdd.n2683 vdd.n853 185
R16110 vdd.n2817 vdd.n853 185
R16111 vdd.n2685 vdd.n2684 185
R16112 vdd.n2684 vdd.n851 185
R16113 vdd.n2686 vdd.n858 185
R16114 vdd.n2811 vdd.n858 185
R16115 vdd.n2688 vdd.n2687 185
R16116 vdd.n2687 vdd.n864 185
R16117 vdd.n2689 vdd.n863 185
R16118 vdd.n2805 vdd.n863 185
R16119 vdd.n2691 vdd.n2690 185
R16120 vdd.n2690 vdd.n871 185
R16121 vdd.n2692 vdd.n870 185
R16122 vdd.n2799 vdd.n870 185
R16123 vdd.n2694 vdd.n2693 185
R16124 vdd.n2693 vdd.n868 185
R16125 vdd.n2695 vdd.n876 185
R16126 vdd.n2793 vdd.n876 185
R16127 vdd.n2697 vdd.n2696 185
R16128 vdd.n2698 vdd.n2697 185
R16129 vdd.n2628 vdd.n881 185
R16130 vdd.n2787 vdd.n881 185
R16131 vdd.n2627 vdd.n2626 185
R16132 vdd.n2626 vdd.t157 185
R16133 vdd.n2625 vdd.n886 185
R16134 vdd.n2781 vdd.n886 185
R16135 vdd.n2245 vdd.n2244 185
R16136 vdd.n2246 vdd.n2245 185
R16137 vdd.n1048 vdd.n1046 185
R16138 vdd.n1046 vdd.n1044 185
R16139 vdd.n1814 vdd.n1813 185
R16140 vdd.n1813 vdd.n1812 185
R16141 vdd.n1051 vdd.n1050 185
R16142 vdd.n1052 vdd.n1051 185
R16143 vdd.n1801 vdd.n1800 185
R16144 vdd.n1802 vdd.n1801 185
R16145 vdd.n1060 vdd.n1059 185
R16146 vdd.n1793 vdd.n1059 185
R16147 vdd.n1796 vdd.n1795 185
R16148 vdd.n1795 vdd.n1794 185
R16149 vdd.n1063 vdd.n1062 185
R16150 vdd.n1069 vdd.n1063 185
R16151 vdd.n1784 vdd.n1783 185
R16152 vdd.n1785 vdd.n1784 185
R16153 vdd.n1071 vdd.n1070 185
R16154 vdd.n1776 vdd.n1070 185
R16155 vdd.n1779 vdd.n1778 185
R16156 vdd.n1778 vdd.n1777 185
R16157 vdd.n1074 vdd.n1073 185
R16158 vdd.n1075 vdd.n1074 185
R16159 vdd.n1767 vdd.n1766 185
R16160 vdd.n1768 vdd.n1767 185
R16161 vdd.n1083 vdd.n1082 185
R16162 vdd.n1082 vdd.n1081 185
R16163 vdd.n1762 vdd.n1761 185
R16164 vdd.n1761 vdd.n1760 185
R16165 vdd.n1086 vdd.n1085 185
R16166 vdd.n1092 vdd.n1086 185
R16167 vdd.n1751 vdd.n1750 185
R16168 vdd.n1752 vdd.n1751 185
R16169 vdd.n1094 vdd.n1093 185
R16170 vdd.n1448 vdd.n1093 185
R16171 vdd.n1451 vdd.n1450 185
R16172 vdd.n1450 vdd.n1449 185
R16173 vdd.n1097 vdd.n1096 185
R16174 vdd.n1104 vdd.n1097 185
R16175 vdd.n1439 vdd.n1438 185
R16176 vdd.n1440 vdd.n1439 185
R16177 vdd.n1106 vdd.n1105 185
R16178 vdd.n1105 vdd.n1103 185
R16179 vdd.n1434 vdd.n1433 185
R16180 vdd.n1433 vdd.n1432 185
R16181 vdd.n1109 vdd.n1108 185
R16182 vdd.n1110 vdd.n1109 185
R16183 vdd.n1423 vdd.n1422 185
R16184 vdd.n1424 vdd.n1423 185
R16185 vdd.n1117 vdd.n1116 185
R16186 vdd.n1415 vdd.n1116 185
R16187 vdd.n1418 vdd.n1417 185
R16188 vdd.n1417 vdd.n1416 185
R16189 vdd.n1120 vdd.n1119 185
R16190 vdd.n1126 vdd.n1120 185
R16191 vdd.n1406 vdd.n1405 185
R16192 vdd.n1407 vdd.n1406 185
R16193 vdd.n1128 vdd.n1127 185
R16194 vdd.n1398 vdd.n1127 185
R16195 vdd.n1401 vdd.n1400 185
R16196 vdd.n1400 vdd.n1399 185
R16197 vdd.n1131 vdd.n1130 185
R16198 vdd.n1132 vdd.n1131 185
R16199 vdd.n1389 vdd.n1388 185
R16200 vdd.n1390 vdd.n1389 185
R16201 vdd.n1140 vdd.n1139 185
R16202 vdd.n1139 vdd.n1138 185
R16203 vdd.n1384 vdd.n1383 185
R16204 vdd.n1383 vdd.n1382 185
R16205 vdd.n1143 vdd.n1142 185
R16206 vdd.n1144 vdd.n1143 185
R16207 vdd.n1372 vdd.n1371 185
R16208 vdd.n1370 vdd.n1183 185
R16209 vdd.n1185 vdd.n1182 185
R16210 vdd.n1374 vdd.n1182 185
R16211 vdd.n1366 vdd.n1187 185
R16212 vdd.n1365 vdd.n1188 185
R16213 vdd.n1364 vdd.n1189 185
R16214 vdd.n1192 vdd.n1190 185
R16215 vdd.n1360 vdd.n1193 185
R16216 vdd.n1359 vdd.n1194 185
R16217 vdd.n1358 vdd.n1195 185
R16218 vdd.n1198 vdd.n1196 185
R16219 vdd.n1354 vdd.n1199 185
R16220 vdd.n1353 vdd.n1200 185
R16221 vdd.n1352 vdd.n1201 185
R16222 vdd.n1204 vdd.n1202 185
R16223 vdd.n1348 vdd.n1205 185
R16224 vdd.n1347 vdd.n1206 185
R16225 vdd.n1346 vdd.n1207 185
R16226 vdd.n1338 vdd.n1208 185
R16227 vdd.n1342 vdd.n1339 185
R16228 vdd.n1337 vdd.n1210 185
R16229 vdd.n1336 vdd.n1211 185
R16230 vdd.n1214 vdd.n1212 185
R16231 vdd.n1332 vdd.n1215 185
R16232 vdd.n1331 vdd.n1216 185
R16233 vdd.n1330 vdd.n1217 185
R16234 vdd.n1220 vdd.n1218 185
R16235 vdd.n1326 vdd.n1221 185
R16236 vdd.n1325 vdd.n1222 185
R16237 vdd.n1324 vdd.n1223 185
R16238 vdd.n1226 vdd.n1224 185
R16239 vdd.n1320 vdd.n1227 185
R16240 vdd.n1319 vdd.n1228 185
R16241 vdd.n1318 vdd.n1229 185
R16242 vdd.n1232 vdd.n1230 185
R16243 vdd.n1314 vdd.n1233 185
R16244 vdd.n1313 vdd.n1234 185
R16245 vdd.n1312 vdd.n1235 185
R16246 vdd.n1238 vdd.n1236 185
R16247 vdd.n1308 vdd.n1239 185
R16248 vdd.n1307 vdd.n1240 185
R16249 vdd.n1306 vdd.n1303 185
R16250 vdd.n1243 vdd.n1241 185
R16251 vdd.n1299 vdd.n1244 185
R16252 vdd.n1298 vdd.n1245 185
R16253 vdd.n1297 vdd.n1246 185
R16254 vdd.n1249 vdd.n1247 185
R16255 vdd.n1293 vdd.n1250 185
R16256 vdd.n1292 vdd.n1251 185
R16257 vdd.n1291 vdd.n1252 185
R16258 vdd.n1255 vdd.n1253 185
R16259 vdd.n1287 vdd.n1256 185
R16260 vdd.n1286 vdd.n1257 185
R16261 vdd.n1285 vdd.n1258 185
R16262 vdd.n1261 vdd.n1259 185
R16263 vdd.n1281 vdd.n1262 185
R16264 vdd.n1280 vdd.n1263 185
R16265 vdd.n1279 vdd.n1264 185
R16266 vdd.n1267 vdd.n1265 185
R16267 vdd.n1275 vdd.n1268 185
R16268 vdd.n1274 vdd.n1269 185
R16269 vdd.n1273 vdd.n1270 185
R16270 vdd.n1271 vdd.n1151 185
R16271 vdd.n1376 vdd.n1375 185
R16272 vdd.n1375 vdd.n1374 185
R16273 vdd.n2249 vdd.n2248 185
R16274 vdd.n2253 vdd.n1040 185
R16275 vdd.n1916 vdd.n1039 185
R16276 vdd.n1919 vdd.n1918 185
R16277 vdd.n1921 vdd.n1920 185
R16278 vdd.n1924 vdd.n1923 185
R16279 vdd.n1926 vdd.n1925 185
R16280 vdd.n1928 vdd.n1914 185
R16281 vdd.n1930 vdd.n1929 185
R16282 vdd.n1931 vdd.n1908 185
R16283 vdd.n1933 vdd.n1932 185
R16284 vdd.n1935 vdd.n1906 185
R16285 vdd.n1937 vdd.n1936 185
R16286 vdd.n1938 vdd.n1901 185
R16287 vdd.n1940 vdd.n1939 185
R16288 vdd.n1942 vdd.n1899 185
R16289 vdd.n1944 vdd.n1943 185
R16290 vdd.n1945 vdd.n1895 185
R16291 vdd.n1947 vdd.n1946 185
R16292 vdd.n1949 vdd.n1892 185
R16293 vdd.n1951 vdd.n1950 185
R16294 vdd.n1893 vdd.n1886 185
R16295 vdd.n1955 vdd.n1890 185
R16296 vdd.n1956 vdd.n1882 185
R16297 vdd.n1958 vdd.n1957 185
R16298 vdd.n1960 vdd.n1880 185
R16299 vdd.n1962 vdd.n1961 185
R16300 vdd.n1963 vdd.n1875 185
R16301 vdd.n1965 vdd.n1964 185
R16302 vdd.n1967 vdd.n1873 185
R16303 vdd.n1969 vdd.n1968 185
R16304 vdd.n1970 vdd.n1868 185
R16305 vdd.n1972 vdd.n1971 185
R16306 vdd.n1974 vdd.n1866 185
R16307 vdd.n1976 vdd.n1975 185
R16308 vdd.n1977 vdd.n1861 185
R16309 vdd.n1979 vdd.n1978 185
R16310 vdd.n1981 vdd.n1859 185
R16311 vdd.n1983 vdd.n1982 185
R16312 vdd.n1984 vdd.n1855 185
R16313 vdd.n1986 vdd.n1985 185
R16314 vdd.n1988 vdd.n1852 185
R16315 vdd.n1990 vdd.n1989 185
R16316 vdd.n1853 vdd.n1846 185
R16317 vdd.n1994 vdd.n1850 185
R16318 vdd.n1995 vdd.n1842 185
R16319 vdd.n1997 vdd.n1996 185
R16320 vdd.n1999 vdd.n1840 185
R16321 vdd.n2001 vdd.n2000 185
R16322 vdd.n2002 vdd.n1835 185
R16323 vdd.n2004 vdd.n2003 185
R16324 vdd.n2006 vdd.n1833 185
R16325 vdd.n2008 vdd.n2007 185
R16326 vdd.n2009 vdd.n1828 185
R16327 vdd.n2011 vdd.n2010 185
R16328 vdd.n2013 vdd.n1827 185
R16329 vdd.n2014 vdd.n1824 185
R16330 vdd.n2017 vdd.n2016 185
R16331 vdd.n1826 vdd.n1822 185
R16332 vdd.n2234 vdd.n1820 185
R16333 vdd.n2236 vdd.n2235 185
R16334 vdd.n2238 vdd.n1818 185
R16335 vdd.n2240 vdd.n2239 185
R16336 vdd.n2241 vdd.n1047 185
R16337 vdd.n2247 vdd.n1043 185
R16338 vdd.n2247 vdd.n2246 185
R16339 vdd.n1055 vdd.n1042 185
R16340 vdd.n1044 vdd.n1042 185
R16341 vdd.n1811 vdd.n1810 185
R16342 vdd.n1812 vdd.n1811 185
R16343 vdd.n1054 vdd.n1053 185
R16344 vdd.n1053 vdd.n1052 185
R16345 vdd.n1804 vdd.n1803 185
R16346 vdd.n1803 vdd.n1802 185
R16347 vdd.n1058 vdd.n1057 185
R16348 vdd.n1793 vdd.n1058 185
R16349 vdd.n1792 vdd.n1791 185
R16350 vdd.n1794 vdd.n1792 185
R16351 vdd.n1065 vdd.n1064 185
R16352 vdd.n1069 vdd.n1064 185
R16353 vdd.n1787 vdd.n1786 185
R16354 vdd.n1786 vdd.n1785 185
R16355 vdd.n1068 vdd.n1067 185
R16356 vdd.n1776 vdd.n1068 185
R16357 vdd.n1775 vdd.n1774 185
R16358 vdd.n1777 vdd.n1775 185
R16359 vdd.n1077 vdd.n1076 185
R16360 vdd.n1076 vdd.n1075 185
R16361 vdd.n1770 vdd.n1769 185
R16362 vdd.n1769 vdd.n1768 185
R16363 vdd.n1080 vdd.n1079 185
R16364 vdd.n1081 vdd.n1080 185
R16365 vdd.n1759 vdd.n1758 185
R16366 vdd.n1760 vdd.n1759 185
R16367 vdd.n1088 vdd.n1087 185
R16368 vdd.n1092 vdd.n1087 185
R16369 vdd.n1754 vdd.n1753 185
R16370 vdd.n1753 vdd.n1752 185
R16371 vdd.n1091 vdd.n1090 185
R16372 vdd.n1448 vdd.n1091 185
R16373 vdd.n1447 vdd.n1446 185
R16374 vdd.n1449 vdd.n1447 185
R16375 vdd.n1099 vdd.n1098 185
R16376 vdd.n1104 vdd.n1098 185
R16377 vdd.n1442 vdd.n1441 185
R16378 vdd.n1441 vdd.n1440 185
R16379 vdd.n1102 vdd.n1101 185
R16380 vdd.n1103 vdd.n1102 185
R16381 vdd.n1431 vdd.n1430 185
R16382 vdd.n1432 vdd.n1431 185
R16383 vdd.n1112 vdd.n1111 185
R16384 vdd.n1111 vdd.n1110 185
R16385 vdd.n1426 vdd.n1425 185
R16386 vdd.n1425 vdd.n1424 185
R16387 vdd.n1115 vdd.n1114 185
R16388 vdd.n1415 vdd.n1115 185
R16389 vdd.n1414 vdd.n1413 185
R16390 vdd.n1416 vdd.n1414 185
R16391 vdd.n1122 vdd.n1121 185
R16392 vdd.n1126 vdd.n1121 185
R16393 vdd.n1409 vdd.n1408 185
R16394 vdd.n1408 vdd.n1407 185
R16395 vdd.n1125 vdd.n1124 185
R16396 vdd.n1398 vdd.n1125 185
R16397 vdd.n1397 vdd.n1396 185
R16398 vdd.n1399 vdd.n1397 185
R16399 vdd.n1134 vdd.n1133 185
R16400 vdd.n1133 vdd.n1132 185
R16401 vdd.n1392 vdd.n1391 185
R16402 vdd.n1391 vdd.n1390 185
R16403 vdd.n1137 vdd.n1136 185
R16404 vdd.n1138 vdd.n1137 185
R16405 vdd.n1381 vdd.n1380 185
R16406 vdd.n1382 vdd.n1381 185
R16407 vdd.n1146 vdd.n1145 185
R16408 vdd.n1145 vdd.n1144 185
R16409 vdd.n927 vdd.n925 185
R16410 vdd.n2449 vdd.n925 185
R16411 vdd.n2371 vdd.n944 185
R16412 vdd.n944 vdd.t15 185
R16413 vdd.n2373 vdd.n2372 185
R16414 vdd.n2374 vdd.n2373 185
R16415 vdd.n2370 vdd.n943 185
R16416 vdd.n2073 vdd.n943 185
R16417 vdd.n2369 vdd.n2368 185
R16418 vdd.n2368 vdd.n2367 185
R16419 vdd.n946 vdd.n945 185
R16420 vdd.n947 vdd.n946 185
R16421 vdd.n2358 vdd.n2357 185
R16422 vdd.n2359 vdd.n2358 185
R16423 vdd.n2356 vdd.n957 185
R16424 vdd.n957 vdd.n954 185
R16425 vdd.n2355 vdd.n2354 185
R16426 vdd.n2354 vdd.n2353 185
R16427 vdd.n959 vdd.n958 185
R16428 vdd.n960 vdd.n959 185
R16429 vdd.n2346 vdd.n2345 185
R16430 vdd.n2347 vdd.n2346 185
R16431 vdd.n2344 vdd.n968 185
R16432 vdd.n973 vdd.n968 185
R16433 vdd.n2343 vdd.n2342 185
R16434 vdd.n2342 vdd.n2341 185
R16435 vdd.n970 vdd.n969 185
R16436 vdd.n979 vdd.n970 185
R16437 vdd.n2334 vdd.n2333 185
R16438 vdd.n2335 vdd.n2334 185
R16439 vdd.n2332 vdd.n980 185
R16440 vdd.n2174 vdd.n980 185
R16441 vdd.n2331 vdd.n2330 185
R16442 vdd.n2330 vdd.n2329 185
R16443 vdd.n982 vdd.n981 185
R16444 vdd.n983 vdd.n982 185
R16445 vdd.n2322 vdd.n2321 185
R16446 vdd.n2323 vdd.n2322 185
R16447 vdd.n2320 vdd.n992 185
R16448 vdd.n992 vdd.n989 185
R16449 vdd.n2319 vdd.n2318 185
R16450 vdd.n2318 vdd.n2317 185
R16451 vdd.n994 vdd.n993 185
R16452 vdd.n1004 vdd.n994 185
R16453 vdd.n2309 vdd.n2308 185
R16454 vdd.n2310 vdd.n2309 185
R16455 vdd.n2307 vdd.n1005 185
R16456 vdd.n1005 vdd.n1001 185
R16457 vdd.n2306 vdd.n2305 185
R16458 vdd.n2305 vdd.n2304 185
R16459 vdd.n1007 vdd.n1006 185
R16460 vdd.n1008 vdd.n1007 185
R16461 vdd.n2297 vdd.n2296 185
R16462 vdd.n2298 vdd.n2297 185
R16463 vdd.n2295 vdd.n1017 185
R16464 vdd.n1017 vdd.n1014 185
R16465 vdd.n2294 vdd.n2293 185
R16466 vdd.n2293 vdd.n2292 185
R16467 vdd.n1019 vdd.n1018 185
R16468 vdd.n2029 vdd.n2028 185
R16469 vdd.n2030 vdd.n2026 185
R16470 vdd.n2026 vdd.n1020 185
R16471 vdd.n2032 vdd.n2031 185
R16472 vdd.n2034 vdd.n2025 185
R16473 vdd.n2037 vdd.n2036 185
R16474 vdd.n2038 vdd.n2024 185
R16475 vdd.n2040 vdd.n2039 185
R16476 vdd.n2042 vdd.n2023 185
R16477 vdd.n2045 vdd.n2044 185
R16478 vdd.n2046 vdd.n2022 185
R16479 vdd.n2048 vdd.n2047 185
R16480 vdd.n2050 vdd.n2021 185
R16481 vdd.n2053 vdd.n2052 185
R16482 vdd.n2054 vdd.n2020 185
R16483 vdd.n2056 vdd.n2055 185
R16484 vdd.n2058 vdd.n2019 185
R16485 vdd.n2231 vdd.n2059 185
R16486 vdd.n2230 vdd.n2229 185
R16487 vdd.n2227 vdd.n2060 185
R16488 vdd.n2225 vdd.n2224 185
R16489 vdd.n2223 vdd.n2061 185
R16490 vdd.n2222 vdd.n2221 185
R16491 vdd.n2219 vdd.n2062 185
R16492 vdd.n2217 vdd.n2216 185
R16493 vdd.n2215 vdd.n2063 185
R16494 vdd.n2214 vdd.n2213 185
R16495 vdd.n2211 vdd.n2064 185
R16496 vdd.n2209 vdd.n2208 185
R16497 vdd.n2207 vdd.n2065 185
R16498 vdd.n2206 vdd.n2205 185
R16499 vdd.n2203 vdd.n2066 185
R16500 vdd.n2201 vdd.n2200 185
R16501 vdd.n2199 vdd.n2067 185
R16502 vdd.n2198 vdd.n2197 185
R16503 vdd.n2452 vdd.n2451 185
R16504 vdd.n2454 vdd.n2453 185
R16505 vdd.n2456 vdd.n2455 185
R16506 vdd.n2459 vdd.n2458 185
R16507 vdd.n2461 vdd.n2460 185
R16508 vdd.n2463 vdd.n2462 185
R16509 vdd.n2465 vdd.n2464 185
R16510 vdd.n2467 vdd.n2466 185
R16511 vdd.n2469 vdd.n2468 185
R16512 vdd.n2471 vdd.n2470 185
R16513 vdd.n2473 vdd.n2472 185
R16514 vdd.n2475 vdd.n2474 185
R16515 vdd.n2477 vdd.n2476 185
R16516 vdd.n2479 vdd.n2478 185
R16517 vdd.n2481 vdd.n2480 185
R16518 vdd.n2483 vdd.n2482 185
R16519 vdd.n2485 vdd.n2484 185
R16520 vdd.n2487 vdd.n2486 185
R16521 vdd.n2489 vdd.n2488 185
R16522 vdd.n2491 vdd.n2490 185
R16523 vdd.n2493 vdd.n2492 185
R16524 vdd.n2495 vdd.n2494 185
R16525 vdd.n2497 vdd.n2496 185
R16526 vdd.n2499 vdd.n2498 185
R16527 vdd.n2501 vdd.n2500 185
R16528 vdd.n2503 vdd.n2502 185
R16529 vdd.n2505 vdd.n2504 185
R16530 vdd.n2507 vdd.n2506 185
R16531 vdd.n2509 vdd.n2508 185
R16532 vdd.n2511 vdd.n2510 185
R16533 vdd.n2513 vdd.n2512 185
R16534 vdd.n2515 vdd.n2514 185
R16535 vdd.n2517 vdd.n2516 185
R16536 vdd.n2518 vdd.n926 185
R16537 vdd.n2520 vdd.n2519 185
R16538 vdd.n2521 vdd.n2520 185
R16539 vdd.n2450 vdd.n930 185
R16540 vdd.n2450 vdd.n2449 185
R16541 vdd.n2071 vdd.n931 185
R16542 vdd.t15 vdd.n931 185
R16543 vdd.n2072 vdd.n941 185
R16544 vdd.n2374 vdd.n941 185
R16545 vdd.n2075 vdd.n2074 185
R16546 vdd.n2074 vdd.n2073 185
R16547 vdd.n2076 vdd.n948 185
R16548 vdd.n2367 vdd.n948 185
R16549 vdd.n2078 vdd.n2077 185
R16550 vdd.n2077 vdd.n947 185
R16551 vdd.n2079 vdd.n955 185
R16552 vdd.n2359 vdd.n955 185
R16553 vdd.n2081 vdd.n2080 185
R16554 vdd.n2080 vdd.n954 185
R16555 vdd.n2082 vdd.n961 185
R16556 vdd.n2353 vdd.n961 185
R16557 vdd.n2084 vdd.n2083 185
R16558 vdd.n2083 vdd.n960 185
R16559 vdd.n2085 vdd.n966 185
R16560 vdd.n2347 vdd.n966 185
R16561 vdd.n2087 vdd.n2086 185
R16562 vdd.n2086 vdd.n973 185
R16563 vdd.n2088 vdd.n971 185
R16564 vdd.n2341 vdd.n971 185
R16565 vdd.n2090 vdd.n2089 185
R16566 vdd.n2089 vdd.n979 185
R16567 vdd.n2091 vdd.n977 185
R16568 vdd.n2335 vdd.n977 185
R16569 vdd.n2176 vdd.n2175 185
R16570 vdd.n2175 vdd.n2174 185
R16571 vdd.n2177 vdd.n984 185
R16572 vdd.n2329 vdd.n984 185
R16573 vdd.n2179 vdd.n2178 185
R16574 vdd.n2178 vdd.n983 185
R16575 vdd.n2180 vdd.n990 185
R16576 vdd.n2323 vdd.n990 185
R16577 vdd.n2182 vdd.n2181 185
R16578 vdd.n2181 vdd.n989 185
R16579 vdd.n2183 vdd.n995 185
R16580 vdd.n2317 vdd.n995 185
R16581 vdd.n2185 vdd.n2184 185
R16582 vdd.n2184 vdd.n1004 185
R16583 vdd.n2186 vdd.n1002 185
R16584 vdd.n2310 vdd.n1002 185
R16585 vdd.n2188 vdd.n2187 185
R16586 vdd.n2187 vdd.n1001 185
R16587 vdd.n2189 vdd.n1009 185
R16588 vdd.n2304 vdd.n1009 185
R16589 vdd.n2191 vdd.n2190 185
R16590 vdd.n2190 vdd.n1008 185
R16591 vdd.n2192 vdd.n1015 185
R16592 vdd.n2298 vdd.n1015 185
R16593 vdd.n2194 vdd.n2193 185
R16594 vdd.n2193 vdd.n1014 185
R16595 vdd.n2195 vdd.n1021 185
R16596 vdd.n2292 vdd.n1021 185
R16597 vdd.n370 vdd.n369 185
R16598 vdd.n3254 vdd.n370 185
R16599 vdd.n3257 vdd.n3256 185
R16600 vdd.n3256 vdd.n3255 185
R16601 vdd.n3258 vdd.n364 185
R16602 vdd.n364 vdd.n363 185
R16603 vdd.n3260 vdd.n3259 185
R16604 vdd.n3261 vdd.n3260 185
R16605 vdd.n359 vdd.n358 185
R16606 vdd.n3262 vdd.n359 185
R16607 vdd.n3265 vdd.n3264 185
R16608 vdd.n3264 vdd.n3263 185
R16609 vdd.n3266 vdd.n353 185
R16610 vdd.n3236 vdd.n353 185
R16611 vdd.n3268 vdd.n3267 185
R16612 vdd.n3269 vdd.n3268 185
R16613 vdd.n348 vdd.n347 185
R16614 vdd.n3270 vdd.n348 185
R16615 vdd.n3273 vdd.n3272 185
R16616 vdd.n3272 vdd.n3271 185
R16617 vdd.n3274 vdd.n342 185
R16618 vdd.n349 vdd.n342 185
R16619 vdd.n3276 vdd.n3275 185
R16620 vdd.n3277 vdd.n3276 185
R16621 vdd.n338 vdd.n337 185
R16622 vdd.n3278 vdd.n338 185
R16623 vdd.n3281 vdd.n3280 185
R16624 vdd.n3280 vdd.n3279 185
R16625 vdd.n3282 vdd.n333 185
R16626 vdd.n333 vdd.n332 185
R16627 vdd.n3284 vdd.n3283 185
R16628 vdd.n3285 vdd.n3284 185
R16629 vdd.n327 vdd.n325 185
R16630 vdd.n3286 vdd.n327 185
R16631 vdd.n3289 vdd.n3288 185
R16632 vdd.n3288 vdd.n3287 185
R16633 vdd.n326 vdd.n324 185
R16634 vdd.n328 vdd.n326 185
R16635 vdd.n3212 vdd.n3211 185
R16636 vdd.n3213 vdd.n3212 185
R16637 vdd.n615 vdd.n614 185
R16638 vdd.n614 vdd.n613 185
R16639 vdd.n3207 vdd.n3206 185
R16640 vdd.n3206 vdd.n3205 185
R16641 vdd.n618 vdd.n617 185
R16642 vdd.n624 vdd.n618 185
R16643 vdd.n3193 vdd.n3192 185
R16644 vdd.n3194 vdd.n3193 185
R16645 vdd.n626 vdd.n625 185
R16646 vdd.n3185 vdd.n625 185
R16647 vdd.n3188 vdd.n3187 185
R16648 vdd.n3187 vdd.n3186 185
R16649 vdd.n629 vdd.n628 185
R16650 vdd.n636 vdd.n629 185
R16651 vdd.n3176 vdd.n3175 185
R16652 vdd.n3177 vdd.n3176 185
R16653 vdd.n638 vdd.n637 185
R16654 vdd.n637 vdd.n635 185
R16655 vdd.n3171 vdd.n3170 185
R16656 vdd.n3170 vdd.n3169 185
R16657 vdd.n641 vdd.n640 185
R16658 vdd.n642 vdd.n641 185
R16659 vdd.n3160 vdd.n3159 185
R16660 vdd.n3161 vdd.n3160 185
R16661 vdd.n650 vdd.n649 185
R16662 vdd.n649 vdd.n648 185
R16663 vdd.n3155 vdd.n3154 185
R16664 vdd.n3154 vdd.n3153 185
R16665 vdd.n653 vdd.n652 185
R16666 vdd.n659 vdd.n653 185
R16667 vdd.n3144 vdd.n3143 185
R16668 vdd.n3145 vdd.n3144 185
R16669 vdd.n3140 vdd.n660 185
R16670 vdd.n3139 vdd.n3138 185
R16671 vdd.n3136 vdd.n662 185
R16672 vdd.n3136 vdd.n658 185
R16673 vdd.n3135 vdd.n3134 185
R16674 vdd.n3133 vdd.n3132 185
R16675 vdd.n3131 vdd.n3130 185
R16676 vdd.n3129 vdd.n3128 185
R16677 vdd.n3127 vdd.n668 185
R16678 vdd.n3125 vdd.n3124 185
R16679 vdd.n3123 vdd.n669 185
R16680 vdd.n3122 vdd.n3121 185
R16681 vdd.n3119 vdd.n674 185
R16682 vdd.n3117 vdd.n3116 185
R16683 vdd.n3115 vdd.n675 185
R16684 vdd.n3114 vdd.n3113 185
R16685 vdd.n3111 vdd.n680 185
R16686 vdd.n3109 vdd.n3108 185
R16687 vdd.n3107 vdd.n681 185
R16688 vdd.n3106 vdd.n3105 185
R16689 vdd.n3103 vdd.n688 185
R16690 vdd.n3101 vdd.n3100 185
R16691 vdd.n3099 vdd.n689 185
R16692 vdd.n3098 vdd.n3097 185
R16693 vdd.n3095 vdd.n694 185
R16694 vdd.n3093 vdd.n3092 185
R16695 vdd.n3091 vdd.n695 185
R16696 vdd.n3090 vdd.n3089 185
R16697 vdd.n3087 vdd.n700 185
R16698 vdd.n3085 vdd.n3084 185
R16699 vdd.n3083 vdd.n701 185
R16700 vdd.n3082 vdd.n3081 185
R16701 vdd.n3079 vdd.n706 185
R16702 vdd.n3077 vdd.n3076 185
R16703 vdd.n3075 vdd.n707 185
R16704 vdd.n3074 vdd.n3073 185
R16705 vdd.n3071 vdd.n712 185
R16706 vdd.n3069 vdd.n3068 185
R16707 vdd.n3067 vdd.n713 185
R16708 vdd.n3066 vdd.n3065 185
R16709 vdd.n3063 vdd.n718 185
R16710 vdd.n3061 vdd.n3060 185
R16711 vdd.n3059 vdd.n719 185
R16712 vdd.n728 vdd.n722 185
R16713 vdd.n3055 vdd.n3054 185
R16714 vdd.n3052 vdd.n726 185
R16715 vdd.n3051 vdd.n3050 185
R16716 vdd.n3049 vdd.n3048 185
R16717 vdd.n3047 vdd.n732 185
R16718 vdd.n3045 vdd.n3044 185
R16719 vdd.n3043 vdd.n733 185
R16720 vdd.n3042 vdd.n3041 185
R16721 vdd.n3039 vdd.n738 185
R16722 vdd.n3037 vdd.n3036 185
R16723 vdd.n3035 vdd.n739 185
R16724 vdd.n3034 vdd.n3033 185
R16725 vdd.n3031 vdd.n744 185
R16726 vdd.n3029 vdd.n3028 185
R16727 vdd.n3027 vdd.n745 185
R16728 vdd.n3026 vdd.n3025 185
R16729 vdd.n3023 vdd.n3022 185
R16730 vdd.n3021 vdd.n3020 185
R16731 vdd.n3019 vdd.n3018 185
R16732 vdd.n3017 vdd.n3016 185
R16733 vdd.n3012 vdd.n657 185
R16734 vdd.n658 vdd.n657 185
R16735 vdd.n3251 vdd.n3250 185
R16736 vdd.n599 vdd.n404 185
R16737 vdd.n598 vdd.n597 185
R16738 vdd.n596 vdd.n595 185
R16739 vdd.n594 vdd.n409 185
R16740 vdd.n590 vdd.n589 185
R16741 vdd.n588 vdd.n587 185
R16742 vdd.n586 vdd.n585 185
R16743 vdd.n584 vdd.n411 185
R16744 vdd.n580 vdd.n579 185
R16745 vdd.n578 vdd.n577 185
R16746 vdd.n576 vdd.n575 185
R16747 vdd.n574 vdd.n413 185
R16748 vdd.n570 vdd.n569 185
R16749 vdd.n568 vdd.n567 185
R16750 vdd.n566 vdd.n565 185
R16751 vdd.n564 vdd.n415 185
R16752 vdd.n560 vdd.n559 185
R16753 vdd.n558 vdd.n557 185
R16754 vdd.n556 vdd.n555 185
R16755 vdd.n554 vdd.n417 185
R16756 vdd.n550 vdd.n549 185
R16757 vdd.n548 vdd.n547 185
R16758 vdd.n546 vdd.n545 185
R16759 vdd.n544 vdd.n421 185
R16760 vdd.n540 vdd.n539 185
R16761 vdd.n538 vdd.n537 185
R16762 vdd.n536 vdd.n535 185
R16763 vdd.n534 vdd.n423 185
R16764 vdd.n530 vdd.n529 185
R16765 vdd.n528 vdd.n527 185
R16766 vdd.n526 vdd.n525 185
R16767 vdd.n524 vdd.n425 185
R16768 vdd.n520 vdd.n519 185
R16769 vdd.n518 vdd.n517 185
R16770 vdd.n516 vdd.n515 185
R16771 vdd.n514 vdd.n427 185
R16772 vdd.n510 vdd.n509 185
R16773 vdd.n508 vdd.n507 185
R16774 vdd.n506 vdd.n505 185
R16775 vdd.n504 vdd.n429 185
R16776 vdd.n500 vdd.n499 185
R16777 vdd.n498 vdd.n497 185
R16778 vdd.n496 vdd.n495 185
R16779 vdd.n494 vdd.n433 185
R16780 vdd.n490 vdd.n489 185
R16781 vdd.n488 vdd.n487 185
R16782 vdd.n486 vdd.n485 185
R16783 vdd.n484 vdd.n435 185
R16784 vdd.n480 vdd.n479 185
R16785 vdd.n478 vdd.n477 185
R16786 vdd.n476 vdd.n475 185
R16787 vdd.n474 vdd.n437 185
R16788 vdd.n470 vdd.n469 185
R16789 vdd.n468 vdd.n467 185
R16790 vdd.n466 vdd.n465 185
R16791 vdd.n464 vdd.n439 185
R16792 vdd.n460 vdd.n459 185
R16793 vdd.n458 vdd.n457 185
R16794 vdd.n456 vdd.n455 185
R16795 vdd.n454 vdd.n441 185
R16796 vdd.n450 vdd.n449 185
R16797 vdd.n448 vdd.n447 185
R16798 vdd.n446 vdd.n445 185
R16799 vdd.n3247 vdd.n372 185
R16800 vdd.n3254 vdd.n372 185
R16801 vdd.n3246 vdd.n371 185
R16802 vdd.n3255 vdd.n371 185
R16803 vdd.n3245 vdd.n3244 185
R16804 vdd.n3244 vdd.n363 185
R16805 vdd.n602 vdd.n362 185
R16806 vdd.n3261 vdd.n362 185
R16807 vdd.n3240 vdd.n361 185
R16808 vdd.n3262 vdd.n361 185
R16809 vdd.n3239 vdd.n360 185
R16810 vdd.n3263 vdd.n360 185
R16811 vdd.n3238 vdd.n3237 185
R16812 vdd.n3237 vdd.n3236 185
R16813 vdd.n604 vdd.n352 185
R16814 vdd.n3269 vdd.n352 185
R16815 vdd.n3232 vdd.n351 185
R16816 vdd.n3270 vdd.n351 185
R16817 vdd.n3231 vdd.n350 185
R16818 vdd.n3271 vdd.n350 185
R16819 vdd.n3230 vdd.n3229 185
R16820 vdd.n3229 vdd.n349 185
R16821 vdd.n606 vdd.n341 185
R16822 vdd.n3277 vdd.n341 185
R16823 vdd.n3225 vdd.n340 185
R16824 vdd.n3278 vdd.n340 185
R16825 vdd.n3224 vdd.n339 185
R16826 vdd.n3279 vdd.n339 185
R16827 vdd.n3223 vdd.n3222 185
R16828 vdd.n3222 vdd.n332 185
R16829 vdd.n608 vdd.n331 185
R16830 vdd.n3285 vdd.n331 185
R16831 vdd.n3218 vdd.n330 185
R16832 vdd.n3286 vdd.n330 185
R16833 vdd.n3217 vdd.n329 185
R16834 vdd.n3287 vdd.n329 185
R16835 vdd.n3216 vdd.n3215 185
R16836 vdd.n3215 vdd.n328 185
R16837 vdd.n3214 vdd.n610 185
R16838 vdd.n3214 vdd.n3213 185
R16839 vdd.n3202 vdd.n612 185
R16840 vdd.n613 vdd.n612 185
R16841 vdd.n3204 vdd.n3203 185
R16842 vdd.n3205 vdd.n3204 185
R16843 vdd.n620 vdd.n619 185
R16844 vdd.n624 vdd.n619 185
R16845 vdd.n3196 vdd.n3195 185
R16846 vdd.n3195 vdd.n3194 185
R16847 vdd.n623 vdd.n622 185
R16848 vdd.n3185 vdd.n623 185
R16849 vdd.n3184 vdd.n3183 185
R16850 vdd.n3186 vdd.n3184 185
R16851 vdd.n631 vdd.n630 185
R16852 vdd.n636 vdd.n630 185
R16853 vdd.n3179 vdd.n3178 185
R16854 vdd.n3178 vdd.n3177 185
R16855 vdd.n634 vdd.n633 185
R16856 vdd.n635 vdd.n634 185
R16857 vdd.n3168 vdd.n3167 185
R16858 vdd.n3169 vdd.n3168 185
R16859 vdd.n644 vdd.n643 185
R16860 vdd.n643 vdd.n642 185
R16861 vdd.n3163 vdd.n3162 185
R16862 vdd.n3162 vdd.n3161 185
R16863 vdd.n647 vdd.n646 185
R16864 vdd.n648 vdd.n647 185
R16865 vdd.n3152 vdd.n3151 185
R16866 vdd.n3153 vdd.n3152 185
R16867 vdd.n655 vdd.n654 185
R16868 vdd.n659 vdd.n654 185
R16869 vdd.n3147 vdd.n3146 185
R16870 vdd.n3146 vdd.n3145 185
R16871 vdd.n884 vdd.n883 185
R16872 vdd.n2772 vdd.n2771 185
R16873 vdd.n2770 vdd.n2555 185
R16874 vdd.n2774 vdd.n2555 185
R16875 vdd.n2769 vdd.n2768 185
R16876 vdd.n2767 vdd.n2766 185
R16877 vdd.n2765 vdd.n2764 185
R16878 vdd.n2763 vdd.n2762 185
R16879 vdd.n2761 vdd.n2760 185
R16880 vdd.n2759 vdd.n2758 185
R16881 vdd.n2757 vdd.n2756 185
R16882 vdd.n2755 vdd.n2754 185
R16883 vdd.n2753 vdd.n2752 185
R16884 vdd.n2751 vdd.n2750 185
R16885 vdd.n2749 vdd.n2748 185
R16886 vdd.n2747 vdd.n2746 185
R16887 vdd.n2745 vdd.n2744 185
R16888 vdd.n2743 vdd.n2742 185
R16889 vdd.n2741 vdd.n2740 185
R16890 vdd.n2739 vdd.n2738 185
R16891 vdd.n2737 vdd.n2736 185
R16892 vdd.n2735 vdd.n2734 185
R16893 vdd.n2733 vdd.n2732 185
R16894 vdd.n2731 vdd.n2730 185
R16895 vdd.n2729 vdd.n2728 185
R16896 vdd.n2727 vdd.n2726 185
R16897 vdd.n2725 vdd.n2724 185
R16898 vdd.n2723 vdd.n2722 185
R16899 vdd.n2721 vdd.n2720 185
R16900 vdd.n2719 vdd.n2718 185
R16901 vdd.n2717 vdd.n2716 185
R16902 vdd.n2715 vdd.n2714 185
R16903 vdd.n2713 vdd.n2712 185
R16904 vdd.n2710 vdd.n2709 185
R16905 vdd.n2708 vdd.n2707 185
R16906 vdd.n2706 vdd.n2705 185
R16907 vdd.n2913 vdd.n2912 185
R16908 vdd.n2914 vdd.n803 185
R16909 vdd.n2916 vdd.n2915 185
R16910 vdd.n2918 vdd.n801 185
R16911 vdd.n2920 vdd.n2919 185
R16912 vdd.n2921 vdd.n800 185
R16913 vdd.n2923 vdd.n2922 185
R16914 vdd.n2925 vdd.n798 185
R16915 vdd.n2927 vdd.n2926 185
R16916 vdd.n2928 vdd.n797 185
R16917 vdd.n2930 vdd.n2929 185
R16918 vdd.n2932 vdd.n795 185
R16919 vdd.n2934 vdd.n2933 185
R16920 vdd.n2935 vdd.n794 185
R16921 vdd.n2937 vdd.n2936 185
R16922 vdd.n2939 vdd.n792 185
R16923 vdd.n2941 vdd.n2940 185
R16924 vdd.n2943 vdd.n791 185
R16925 vdd.n2945 vdd.n2944 185
R16926 vdd.n2947 vdd.n789 185
R16927 vdd.n2949 vdd.n2948 185
R16928 vdd.n2950 vdd.n788 185
R16929 vdd.n2952 vdd.n2951 185
R16930 vdd.n2954 vdd.n786 185
R16931 vdd.n2956 vdd.n2955 185
R16932 vdd.n2957 vdd.n785 185
R16933 vdd.n2959 vdd.n2958 185
R16934 vdd.n2961 vdd.n783 185
R16935 vdd.n2963 vdd.n2962 185
R16936 vdd.n2964 vdd.n782 185
R16937 vdd.n2966 vdd.n2965 185
R16938 vdd.n2968 vdd.n781 185
R16939 vdd.n2969 vdd.n780 185
R16940 vdd.n2972 vdd.n2971 185
R16941 vdd.n2973 vdd.n778 185
R16942 vdd.n778 vdd.n756 185
R16943 vdd.n2910 vdd.n775 185
R16944 vdd.n2976 vdd.n775 185
R16945 vdd.n2909 vdd.n2908 185
R16946 vdd.n2908 vdd.n774 185
R16947 vdd.n2907 vdd.n807 185
R16948 vdd.n2907 vdd.n2906 185
R16949 vdd.n2661 vdd.n808 185
R16950 vdd.n817 vdd.n808 185
R16951 vdd.n2662 vdd.n815 185
R16952 vdd.n2900 vdd.n815 185
R16953 vdd.n2664 vdd.n2663 185
R16954 vdd.n2663 vdd.n814 185
R16955 vdd.n2665 vdd.n823 185
R16956 vdd.n2849 vdd.n823 185
R16957 vdd.n2667 vdd.n2666 185
R16958 vdd.n2666 vdd.n822 185
R16959 vdd.n2668 vdd.n829 185
R16960 vdd.n2843 vdd.n829 185
R16961 vdd.n2670 vdd.n2669 185
R16962 vdd.n2669 vdd.n828 185
R16963 vdd.n2671 vdd.n834 185
R16964 vdd.n2835 vdd.n834 185
R16965 vdd.n2673 vdd.n2672 185
R16966 vdd.n2672 vdd.n841 185
R16967 vdd.n2674 vdd.n839 185
R16968 vdd.n2829 vdd.n839 185
R16969 vdd.n2676 vdd.n2675 185
R16970 vdd.n2677 vdd.n2676 185
R16971 vdd.n2660 vdd.n846 185
R16972 vdd.n2823 vdd.n846 185
R16973 vdd.n2659 vdd.n2658 185
R16974 vdd.n2658 vdd.n845 185
R16975 vdd.n2657 vdd.n852 185
R16976 vdd.n2817 vdd.n852 185
R16977 vdd.n2656 vdd.n2655 185
R16978 vdd.n2655 vdd.n851 185
R16979 vdd.n2654 vdd.n857 185
R16980 vdd.n2811 vdd.n857 185
R16981 vdd.n2653 vdd.n2652 185
R16982 vdd.n2652 vdd.n864 185
R16983 vdd.n2651 vdd.n862 185
R16984 vdd.n2805 vdd.n862 185
R16985 vdd.n2650 vdd.n2649 185
R16986 vdd.n2649 vdd.n871 185
R16987 vdd.n2648 vdd.n869 185
R16988 vdd.n2799 vdd.n869 185
R16989 vdd.n2647 vdd.n2646 185
R16990 vdd.n2646 vdd.n868 185
R16991 vdd.n2558 vdd.n875 185
R16992 vdd.n2793 vdd.n875 185
R16993 vdd.n2700 vdd.n2699 185
R16994 vdd.n2699 vdd.n2698 185
R16995 vdd.n2701 vdd.n880 185
R16996 vdd.n2787 vdd.n880 185
R16997 vdd.n2703 vdd.n2702 185
R16998 vdd.n2702 vdd.t157 185
R16999 vdd.n2704 vdd.n885 185
R17000 vdd.n2781 vdd.n885 185
R17001 vdd.n2783 vdd.n2782 185
R17002 vdd.n2782 vdd.n2781 185
R17003 vdd.n2784 vdd.n882 185
R17004 vdd.n882 vdd.t157 185
R17005 vdd.n2786 vdd.n2785 185
R17006 vdd.n2787 vdd.n2786 185
R17007 vdd.n874 vdd.n873 185
R17008 vdd.n2698 vdd.n874 185
R17009 vdd.n2795 vdd.n2794 185
R17010 vdd.n2794 vdd.n2793 185
R17011 vdd.n2796 vdd.n872 185
R17012 vdd.n872 vdd.n868 185
R17013 vdd.n2798 vdd.n2797 185
R17014 vdd.n2799 vdd.n2798 185
R17015 vdd.n861 vdd.n860 185
R17016 vdd.n871 vdd.n861 185
R17017 vdd.n2807 vdd.n2806 185
R17018 vdd.n2806 vdd.n2805 185
R17019 vdd.n2808 vdd.n859 185
R17020 vdd.n864 vdd.n859 185
R17021 vdd.n2810 vdd.n2809 185
R17022 vdd.n2811 vdd.n2810 185
R17023 vdd.n850 vdd.n849 185
R17024 vdd.n851 vdd.n850 185
R17025 vdd.n2819 vdd.n2818 185
R17026 vdd.n2818 vdd.n2817 185
R17027 vdd.n2820 vdd.n848 185
R17028 vdd.n848 vdd.n845 185
R17029 vdd.n2822 vdd.n2821 185
R17030 vdd.n2823 vdd.n2822 185
R17031 vdd.n838 vdd.n837 185
R17032 vdd.n2677 vdd.n838 185
R17033 vdd.n2831 vdd.n2830 185
R17034 vdd.n2830 vdd.n2829 185
R17035 vdd.n2832 vdd.n836 185
R17036 vdd.n841 vdd.n836 185
R17037 vdd.n2834 vdd.n2833 185
R17038 vdd.n2835 vdd.n2834 185
R17039 vdd.n827 vdd.n826 185
R17040 vdd.n828 vdd.n827 185
R17041 vdd.n2845 vdd.n2844 185
R17042 vdd.n2844 vdd.n2843 185
R17043 vdd.n2846 vdd.n825 185
R17044 vdd.n825 vdd.n822 185
R17045 vdd.n2848 vdd.n2847 185
R17046 vdd.n2849 vdd.n2848 185
R17047 vdd.n813 vdd.n812 185
R17048 vdd.n814 vdd.n813 185
R17049 vdd.n2902 vdd.n2901 185
R17050 vdd.n2901 vdd.n2900 185
R17051 vdd.n2903 vdd.n811 185
R17052 vdd.n817 vdd.n811 185
R17053 vdd.n2905 vdd.n2904 185
R17054 vdd.n2906 vdd.n2905 185
R17055 vdd.n779 vdd.n777 185
R17056 vdd.n777 vdd.n774 185
R17057 vdd.n2975 vdd.n2974 185
R17058 vdd.n2976 vdd.n2975 185
R17059 vdd.n2448 vdd.n2447 185
R17060 vdd.n2449 vdd.n2448 185
R17061 vdd.n935 vdd.n933 185
R17062 vdd.n933 vdd.t15 185
R17063 vdd.n2363 vdd.n942 185
R17064 vdd.n2374 vdd.n942 185
R17065 vdd.n2364 vdd.n951 185
R17066 vdd.n2073 vdd.n951 185
R17067 vdd.n2366 vdd.n2365 185
R17068 vdd.n2367 vdd.n2366 185
R17069 vdd.n2362 vdd.n950 185
R17070 vdd.n950 vdd.n947 185
R17071 vdd.n2361 vdd.n2360 185
R17072 vdd.n2360 vdd.n2359 185
R17073 vdd.n953 vdd.n952 185
R17074 vdd.n954 vdd.n953 185
R17075 vdd.n2352 vdd.n2351 185
R17076 vdd.n2353 vdd.n2352 185
R17077 vdd.n2350 vdd.n963 185
R17078 vdd.n963 vdd.n960 185
R17079 vdd.n2349 vdd.n2348 185
R17080 vdd.n2348 vdd.n2347 185
R17081 vdd.n965 vdd.n964 185
R17082 vdd.n973 vdd.n965 185
R17083 vdd.n2340 vdd.n2339 185
R17084 vdd.n2341 vdd.n2340 185
R17085 vdd.n2338 vdd.n974 185
R17086 vdd.n979 vdd.n974 185
R17087 vdd.n2337 vdd.n2336 185
R17088 vdd.n2336 vdd.n2335 185
R17089 vdd.n976 vdd.n975 185
R17090 vdd.n2174 vdd.n976 185
R17091 vdd.n2328 vdd.n2327 185
R17092 vdd.n2329 vdd.n2328 185
R17093 vdd.n2326 vdd.n986 185
R17094 vdd.n986 vdd.n983 185
R17095 vdd.n2325 vdd.n2324 185
R17096 vdd.n2324 vdd.n2323 185
R17097 vdd.n988 vdd.n987 185
R17098 vdd.n989 vdd.n988 185
R17099 vdd.n2316 vdd.n2315 185
R17100 vdd.n2317 vdd.n2316 185
R17101 vdd.n2313 vdd.n997 185
R17102 vdd.n1004 vdd.n997 185
R17103 vdd.n2312 vdd.n2311 185
R17104 vdd.n2311 vdd.n2310 185
R17105 vdd.n1000 vdd.n999 185
R17106 vdd.n1001 vdd.n1000 185
R17107 vdd.n2303 vdd.n2302 185
R17108 vdd.n2304 vdd.n2303 185
R17109 vdd.n2301 vdd.n1011 185
R17110 vdd.n1011 vdd.n1008 185
R17111 vdd.n2300 vdd.n2299 185
R17112 vdd.n2299 vdd.n2298 185
R17113 vdd.n1013 vdd.n1012 185
R17114 vdd.n1014 vdd.n1013 185
R17115 vdd.n2291 vdd.n2290 185
R17116 vdd.n2292 vdd.n2291 185
R17117 vdd.n2379 vdd.n907 185
R17118 vdd.n2521 vdd.n907 185
R17119 vdd.n2381 vdd.n2380 185
R17120 vdd.n2383 vdd.n2382 185
R17121 vdd.n2385 vdd.n2384 185
R17122 vdd.n2387 vdd.n2386 185
R17123 vdd.n2389 vdd.n2388 185
R17124 vdd.n2391 vdd.n2390 185
R17125 vdd.n2393 vdd.n2392 185
R17126 vdd.n2395 vdd.n2394 185
R17127 vdd.n2397 vdd.n2396 185
R17128 vdd.n2399 vdd.n2398 185
R17129 vdd.n2401 vdd.n2400 185
R17130 vdd.n2403 vdd.n2402 185
R17131 vdd.n2405 vdd.n2404 185
R17132 vdd.n2407 vdd.n2406 185
R17133 vdd.n2409 vdd.n2408 185
R17134 vdd.n2411 vdd.n2410 185
R17135 vdd.n2413 vdd.n2412 185
R17136 vdd.n2415 vdd.n2414 185
R17137 vdd.n2417 vdd.n2416 185
R17138 vdd.n2419 vdd.n2418 185
R17139 vdd.n2421 vdd.n2420 185
R17140 vdd.n2423 vdd.n2422 185
R17141 vdd.n2425 vdd.n2424 185
R17142 vdd.n2427 vdd.n2426 185
R17143 vdd.n2429 vdd.n2428 185
R17144 vdd.n2431 vdd.n2430 185
R17145 vdd.n2433 vdd.n2432 185
R17146 vdd.n2435 vdd.n2434 185
R17147 vdd.n2437 vdd.n2436 185
R17148 vdd.n2439 vdd.n2438 185
R17149 vdd.n2441 vdd.n2440 185
R17150 vdd.n2443 vdd.n2442 185
R17151 vdd.n2445 vdd.n2444 185
R17152 vdd.n2446 vdd.n934 185
R17153 vdd.n2378 vdd.n932 185
R17154 vdd.n2449 vdd.n932 185
R17155 vdd.n2377 vdd.n2376 185
R17156 vdd.n2376 vdd.t15 185
R17157 vdd.n2375 vdd.n939 185
R17158 vdd.n2375 vdd.n2374 185
R17159 vdd.n2155 vdd.n940 185
R17160 vdd.n2073 vdd.n940 185
R17161 vdd.n2156 vdd.n949 185
R17162 vdd.n2367 vdd.n949 185
R17163 vdd.n2158 vdd.n2157 185
R17164 vdd.n2157 vdd.n947 185
R17165 vdd.n2159 vdd.n956 185
R17166 vdd.n2359 vdd.n956 185
R17167 vdd.n2161 vdd.n2160 185
R17168 vdd.n2160 vdd.n954 185
R17169 vdd.n2162 vdd.n962 185
R17170 vdd.n2353 vdd.n962 185
R17171 vdd.n2164 vdd.n2163 185
R17172 vdd.n2163 vdd.n960 185
R17173 vdd.n2165 vdd.n967 185
R17174 vdd.n2347 vdd.n967 185
R17175 vdd.n2167 vdd.n2166 185
R17176 vdd.n2166 vdd.n973 185
R17177 vdd.n2168 vdd.n972 185
R17178 vdd.n2341 vdd.n972 185
R17179 vdd.n2170 vdd.n2169 185
R17180 vdd.n2169 vdd.n979 185
R17181 vdd.n2171 vdd.n978 185
R17182 vdd.n2335 vdd.n978 185
R17183 vdd.n2173 vdd.n2172 185
R17184 vdd.n2174 vdd.n2173 185
R17185 vdd.n2154 vdd.n985 185
R17186 vdd.n2329 vdd.n985 185
R17187 vdd.n2153 vdd.n2152 185
R17188 vdd.n2152 vdd.n983 185
R17189 vdd.n2151 vdd.n991 185
R17190 vdd.n2323 vdd.n991 185
R17191 vdd.n2150 vdd.n2149 185
R17192 vdd.n2149 vdd.n989 185
R17193 vdd.n2148 vdd.n996 185
R17194 vdd.n2317 vdd.n996 185
R17195 vdd.n2147 vdd.n2146 185
R17196 vdd.n2146 vdd.n1004 185
R17197 vdd.n2145 vdd.n1003 185
R17198 vdd.n2310 vdd.n1003 185
R17199 vdd.n2144 vdd.n2143 185
R17200 vdd.n2143 vdd.n1001 185
R17201 vdd.n2142 vdd.n1010 185
R17202 vdd.n2304 vdd.n1010 185
R17203 vdd.n2141 vdd.n2140 185
R17204 vdd.n2140 vdd.n1008 185
R17205 vdd.n2139 vdd.n1016 185
R17206 vdd.n2298 vdd.n1016 185
R17207 vdd.n2138 vdd.n2137 185
R17208 vdd.n2137 vdd.n1014 185
R17209 vdd.n2136 vdd.n1022 185
R17210 vdd.n2292 vdd.n1022 185
R17211 vdd.n2289 vdd.n1023 185
R17212 vdd.n2288 vdd.n2287 185
R17213 vdd.n2285 vdd.n1024 185
R17214 vdd.n2283 vdd.n2282 185
R17215 vdd.n2281 vdd.n1025 185
R17216 vdd.n2280 vdd.n2279 185
R17217 vdd.n2277 vdd.n1026 185
R17218 vdd.n2275 vdd.n2274 185
R17219 vdd.n2273 vdd.n1027 185
R17220 vdd.n2272 vdd.n2271 185
R17221 vdd.n2269 vdd.n1028 185
R17222 vdd.n2267 vdd.n2266 185
R17223 vdd.n2265 vdd.n1029 185
R17224 vdd.n2264 vdd.n2263 185
R17225 vdd.n2261 vdd.n1030 185
R17226 vdd.n2259 vdd.n2258 185
R17227 vdd.n2257 vdd.n1031 185
R17228 vdd.n2256 vdd.n1033 185
R17229 vdd.n2101 vdd.n1034 185
R17230 vdd.n2104 vdd.n2103 185
R17231 vdd.n2106 vdd.n2105 185
R17232 vdd.n2108 vdd.n2100 185
R17233 vdd.n2111 vdd.n2110 185
R17234 vdd.n2112 vdd.n2099 185
R17235 vdd.n2114 vdd.n2113 185
R17236 vdd.n2116 vdd.n2098 185
R17237 vdd.n2119 vdd.n2118 185
R17238 vdd.n2120 vdd.n2097 185
R17239 vdd.n2122 vdd.n2121 185
R17240 vdd.n2124 vdd.n2096 185
R17241 vdd.n2127 vdd.n2126 185
R17242 vdd.n2128 vdd.n2093 185
R17243 vdd.n2131 vdd.n2130 185
R17244 vdd.n2133 vdd.n2092 185
R17245 vdd.n2135 vdd.n2134 185
R17246 vdd.n2134 vdd.n1020 185
R17247 vdd.n315 vdd.n314 171.744
R17248 vdd.n314 vdd.n313 171.744
R17249 vdd.n313 vdd.n282 171.744
R17250 vdd.n306 vdd.n282 171.744
R17251 vdd.n306 vdd.n305 171.744
R17252 vdd.n305 vdd.n287 171.744
R17253 vdd.n298 vdd.n287 171.744
R17254 vdd.n298 vdd.n297 171.744
R17255 vdd.n297 vdd.n291 171.744
R17256 vdd.n260 vdd.n259 171.744
R17257 vdd.n259 vdd.n258 171.744
R17258 vdd.n258 vdd.n227 171.744
R17259 vdd.n251 vdd.n227 171.744
R17260 vdd.n251 vdd.n250 171.744
R17261 vdd.n250 vdd.n232 171.744
R17262 vdd.n243 vdd.n232 171.744
R17263 vdd.n243 vdd.n242 171.744
R17264 vdd.n242 vdd.n236 171.744
R17265 vdd.n217 vdd.n216 171.744
R17266 vdd.n216 vdd.n215 171.744
R17267 vdd.n215 vdd.n184 171.744
R17268 vdd.n208 vdd.n184 171.744
R17269 vdd.n208 vdd.n207 171.744
R17270 vdd.n207 vdd.n189 171.744
R17271 vdd.n200 vdd.n189 171.744
R17272 vdd.n200 vdd.n199 171.744
R17273 vdd.n199 vdd.n193 171.744
R17274 vdd.n162 vdd.n161 171.744
R17275 vdd.n161 vdd.n160 171.744
R17276 vdd.n160 vdd.n129 171.744
R17277 vdd.n153 vdd.n129 171.744
R17278 vdd.n153 vdd.n152 171.744
R17279 vdd.n152 vdd.n134 171.744
R17280 vdd.n145 vdd.n134 171.744
R17281 vdd.n145 vdd.n144 171.744
R17282 vdd.n144 vdd.n138 171.744
R17283 vdd.n120 vdd.n119 171.744
R17284 vdd.n119 vdd.n118 171.744
R17285 vdd.n118 vdd.n87 171.744
R17286 vdd.n111 vdd.n87 171.744
R17287 vdd.n111 vdd.n110 171.744
R17288 vdd.n110 vdd.n92 171.744
R17289 vdd.n103 vdd.n92 171.744
R17290 vdd.n103 vdd.n102 171.744
R17291 vdd.n102 vdd.n96 171.744
R17292 vdd.n65 vdd.n64 171.744
R17293 vdd.n64 vdd.n63 171.744
R17294 vdd.n63 vdd.n32 171.744
R17295 vdd.n56 vdd.n32 171.744
R17296 vdd.n56 vdd.n55 171.744
R17297 vdd.n55 vdd.n37 171.744
R17298 vdd.n48 vdd.n37 171.744
R17299 vdd.n48 vdd.n47 171.744
R17300 vdd.n47 vdd.n41 171.744
R17301 vdd.n1684 vdd.n1683 171.744
R17302 vdd.n1683 vdd.n1682 171.744
R17303 vdd.n1682 vdd.n1651 171.744
R17304 vdd.n1675 vdd.n1651 171.744
R17305 vdd.n1675 vdd.n1674 171.744
R17306 vdd.n1674 vdd.n1656 171.744
R17307 vdd.n1667 vdd.n1656 171.744
R17308 vdd.n1667 vdd.n1666 171.744
R17309 vdd.n1666 vdd.n1660 171.744
R17310 vdd.n1739 vdd.n1738 171.744
R17311 vdd.n1738 vdd.n1737 171.744
R17312 vdd.n1737 vdd.n1706 171.744
R17313 vdd.n1730 vdd.n1706 171.744
R17314 vdd.n1730 vdd.n1729 171.744
R17315 vdd.n1729 vdd.n1711 171.744
R17316 vdd.n1722 vdd.n1711 171.744
R17317 vdd.n1722 vdd.n1721 171.744
R17318 vdd.n1721 vdd.n1715 171.744
R17319 vdd.n1586 vdd.n1585 171.744
R17320 vdd.n1585 vdd.n1584 171.744
R17321 vdd.n1584 vdd.n1553 171.744
R17322 vdd.n1577 vdd.n1553 171.744
R17323 vdd.n1577 vdd.n1576 171.744
R17324 vdd.n1576 vdd.n1558 171.744
R17325 vdd.n1569 vdd.n1558 171.744
R17326 vdd.n1569 vdd.n1568 171.744
R17327 vdd.n1568 vdd.n1562 171.744
R17328 vdd.n1641 vdd.n1640 171.744
R17329 vdd.n1640 vdd.n1639 171.744
R17330 vdd.n1639 vdd.n1608 171.744
R17331 vdd.n1632 vdd.n1608 171.744
R17332 vdd.n1632 vdd.n1631 171.744
R17333 vdd.n1631 vdd.n1613 171.744
R17334 vdd.n1624 vdd.n1613 171.744
R17335 vdd.n1624 vdd.n1623 171.744
R17336 vdd.n1623 vdd.n1617 171.744
R17337 vdd.n1489 vdd.n1488 171.744
R17338 vdd.n1488 vdd.n1487 171.744
R17339 vdd.n1487 vdd.n1456 171.744
R17340 vdd.n1480 vdd.n1456 171.744
R17341 vdd.n1480 vdd.n1479 171.744
R17342 vdd.n1479 vdd.n1461 171.744
R17343 vdd.n1472 vdd.n1461 171.744
R17344 vdd.n1472 vdd.n1471 171.744
R17345 vdd.n1471 vdd.n1465 171.744
R17346 vdd.n1544 vdd.n1543 171.744
R17347 vdd.n1543 vdd.n1542 171.744
R17348 vdd.n1542 vdd.n1511 171.744
R17349 vdd.n1535 vdd.n1511 171.744
R17350 vdd.n1535 vdd.n1534 171.744
R17351 vdd.n1534 vdd.n1516 171.744
R17352 vdd.n1527 vdd.n1516 171.744
R17353 vdd.n1527 vdd.n1526 171.744
R17354 vdd.n1526 vdd.n1520 171.744
R17355 vdd.n449 vdd.n448 146.341
R17356 vdd.n455 vdd.n454 146.341
R17357 vdd.n459 vdd.n458 146.341
R17358 vdd.n465 vdd.n464 146.341
R17359 vdd.n469 vdd.n468 146.341
R17360 vdd.n475 vdd.n474 146.341
R17361 vdd.n479 vdd.n478 146.341
R17362 vdd.n485 vdd.n484 146.341
R17363 vdd.n489 vdd.n488 146.341
R17364 vdd.n495 vdd.n494 146.341
R17365 vdd.n499 vdd.n498 146.341
R17366 vdd.n505 vdd.n504 146.341
R17367 vdd.n509 vdd.n508 146.341
R17368 vdd.n515 vdd.n514 146.341
R17369 vdd.n519 vdd.n518 146.341
R17370 vdd.n525 vdd.n524 146.341
R17371 vdd.n529 vdd.n528 146.341
R17372 vdd.n535 vdd.n534 146.341
R17373 vdd.n539 vdd.n538 146.341
R17374 vdd.n545 vdd.n544 146.341
R17375 vdd.n549 vdd.n548 146.341
R17376 vdd.n555 vdd.n554 146.341
R17377 vdd.n559 vdd.n558 146.341
R17378 vdd.n565 vdd.n564 146.341
R17379 vdd.n569 vdd.n568 146.341
R17380 vdd.n575 vdd.n574 146.341
R17381 vdd.n579 vdd.n578 146.341
R17382 vdd.n585 vdd.n584 146.341
R17383 vdd.n589 vdd.n588 146.341
R17384 vdd.n595 vdd.n594 146.341
R17385 vdd.n597 vdd.n404 146.341
R17386 vdd.n3146 vdd.n654 146.341
R17387 vdd.n3152 vdd.n654 146.341
R17388 vdd.n3152 vdd.n647 146.341
R17389 vdd.n3162 vdd.n647 146.341
R17390 vdd.n3162 vdd.n643 146.341
R17391 vdd.n3168 vdd.n643 146.341
R17392 vdd.n3168 vdd.n634 146.341
R17393 vdd.n3178 vdd.n634 146.341
R17394 vdd.n3178 vdd.n630 146.341
R17395 vdd.n3184 vdd.n630 146.341
R17396 vdd.n3184 vdd.n623 146.341
R17397 vdd.n3195 vdd.n623 146.341
R17398 vdd.n3195 vdd.n619 146.341
R17399 vdd.n3204 vdd.n619 146.341
R17400 vdd.n3204 vdd.n612 146.341
R17401 vdd.n3214 vdd.n612 146.341
R17402 vdd.n3215 vdd.n3214 146.341
R17403 vdd.n3215 vdd.n329 146.341
R17404 vdd.n330 vdd.n329 146.341
R17405 vdd.n331 vdd.n330 146.341
R17406 vdd.n3222 vdd.n331 146.341
R17407 vdd.n3222 vdd.n339 146.341
R17408 vdd.n340 vdd.n339 146.341
R17409 vdd.n341 vdd.n340 146.341
R17410 vdd.n3229 vdd.n341 146.341
R17411 vdd.n3229 vdd.n350 146.341
R17412 vdd.n351 vdd.n350 146.341
R17413 vdd.n352 vdd.n351 146.341
R17414 vdd.n3237 vdd.n352 146.341
R17415 vdd.n3237 vdd.n360 146.341
R17416 vdd.n361 vdd.n360 146.341
R17417 vdd.n362 vdd.n361 146.341
R17418 vdd.n3244 vdd.n362 146.341
R17419 vdd.n3244 vdd.n371 146.341
R17420 vdd.n372 vdd.n371 146.341
R17421 vdd.n3138 vdd.n3136 146.341
R17422 vdd.n3136 vdd.n3135 146.341
R17423 vdd.n3132 vdd.n3131 146.341
R17424 vdd.n3128 vdd.n3127 146.341
R17425 vdd.n3125 vdd.n669 146.341
R17426 vdd.n3121 vdd.n3119 146.341
R17427 vdd.n3117 vdd.n675 146.341
R17428 vdd.n3113 vdd.n3111 146.341
R17429 vdd.n3109 vdd.n681 146.341
R17430 vdd.n3105 vdd.n3103 146.341
R17431 vdd.n3101 vdd.n689 146.341
R17432 vdd.n3097 vdd.n3095 146.341
R17433 vdd.n3093 vdd.n695 146.341
R17434 vdd.n3089 vdd.n3087 146.341
R17435 vdd.n3085 vdd.n701 146.341
R17436 vdd.n3081 vdd.n3079 146.341
R17437 vdd.n3077 vdd.n707 146.341
R17438 vdd.n3073 vdd.n3071 146.341
R17439 vdd.n3069 vdd.n713 146.341
R17440 vdd.n3065 vdd.n3063 146.341
R17441 vdd.n3061 vdd.n719 146.341
R17442 vdd.n3054 vdd.n728 146.341
R17443 vdd.n3052 vdd.n3051 146.341
R17444 vdd.n3048 vdd.n3047 146.341
R17445 vdd.n3045 vdd.n733 146.341
R17446 vdd.n3041 vdd.n3039 146.341
R17447 vdd.n3037 vdd.n739 146.341
R17448 vdd.n3033 vdd.n3031 146.341
R17449 vdd.n3029 vdd.n745 146.341
R17450 vdd.n3025 vdd.n3023 146.341
R17451 vdd.n3020 vdd.n3019 146.341
R17452 vdd.n3016 vdd.n657 146.341
R17453 vdd.n3144 vdd.n653 146.341
R17454 vdd.n3154 vdd.n653 146.341
R17455 vdd.n3154 vdd.n649 146.341
R17456 vdd.n3160 vdd.n649 146.341
R17457 vdd.n3160 vdd.n641 146.341
R17458 vdd.n3170 vdd.n641 146.341
R17459 vdd.n3170 vdd.n637 146.341
R17460 vdd.n3176 vdd.n637 146.341
R17461 vdd.n3176 vdd.n629 146.341
R17462 vdd.n3187 vdd.n629 146.341
R17463 vdd.n3187 vdd.n625 146.341
R17464 vdd.n3193 vdd.n625 146.341
R17465 vdd.n3193 vdd.n618 146.341
R17466 vdd.n3206 vdd.n618 146.341
R17467 vdd.n3206 vdd.n614 146.341
R17468 vdd.n3212 vdd.n614 146.341
R17469 vdd.n3212 vdd.n326 146.341
R17470 vdd.n3288 vdd.n326 146.341
R17471 vdd.n3288 vdd.n327 146.341
R17472 vdd.n3284 vdd.n327 146.341
R17473 vdd.n3284 vdd.n333 146.341
R17474 vdd.n3280 vdd.n333 146.341
R17475 vdd.n3280 vdd.n338 146.341
R17476 vdd.n3276 vdd.n338 146.341
R17477 vdd.n3276 vdd.n342 146.341
R17478 vdd.n3272 vdd.n342 146.341
R17479 vdd.n3272 vdd.n348 146.341
R17480 vdd.n3268 vdd.n348 146.341
R17481 vdd.n3268 vdd.n353 146.341
R17482 vdd.n3264 vdd.n353 146.341
R17483 vdd.n3264 vdd.n359 146.341
R17484 vdd.n3260 vdd.n359 146.341
R17485 vdd.n3260 vdd.n364 146.341
R17486 vdd.n3256 vdd.n364 146.341
R17487 vdd.n3256 vdd.n370 146.341
R17488 vdd.n2239 vdd.n2238 146.341
R17489 vdd.n2236 vdd.n1820 146.341
R17490 vdd.n2016 vdd.n1826 146.341
R17491 vdd.n2014 vdd.n2013 146.341
R17492 vdd.n2011 vdd.n1828 146.341
R17493 vdd.n2007 vdd.n2006 146.341
R17494 vdd.n2004 vdd.n1835 146.341
R17495 vdd.n2000 vdd.n1999 146.341
R17496 vdd.n1997 vdd.n1842 146.341
R17497 vdd.n1853 vdd.n1850 146.341
R17498 vdd.n1989 vdd.n1988 146.341
R17499 vdd.n1986 vdd.n1855 146.341
R17500 vdd.n1982 vdd.n1981 146.341
R17501 vdd.n1979 vdd.n1861 146.341
R17502 vdd.n1975 vdd.n1974 146.341
R17503 vdd.n1972 vdd.n1868 146.341
R17504 vdd.n1968 vdd.n1967 146.341
R17505 vdd.n1965 vdd.n1875 146.341
R17506 vdd.n1961 vdd.n1960 146.341
R17507 vdd.n1958 vdd.n1882 146.341
R17508 vdd.n1893 vdd.n1890 146.341
R17509 vdd.n1950 vdd.n1949 146.341
R17510 vdd.n1947 vdd.n1895 146.341
R17511 vdd.n1943 vdd.n1942 146.341
R17512 vdd.n1940 vdd.n1901 146.341
R17513 vdd.n1936 vdd.n1935 146.341
R17514 vdd.n1933 vdd.n1908 146.341
R17515 vdd.n1929 vdd.n1928 146.341
R17516 vdd.n1926 vdd.n1923 146.341
R17517 vdd.n1921 vdd.n1918 146.341
R17518 vdd.n1916 vdd.n1040 146.341
R17519 vdd.n1381 vdd.n1145 146.341
R17520 vdd.n1381 vdd.n1137 146.341
R17521 vdd.n1391 vdd.n1137 146.341
R17522 vdd.n1391 vdd.n1133 146.341
R17523 vdd.n1397 vdd.n1133 146.341
R17524 vdd.n1397 vdd.n1125 146.341
R17525 vdd.n1408 vdd.n1125 146.341
R17526 vdd.n1408 vdd.n1121 146.341
R17527 vdd.n1414 vdd.n1121 146.341
R17528 vdd.n1414 vdd.n1115 146.341
R17529 vdd.n1425 vdd.n1115 146.341
R17530 vdd.n1425 vdd.n1111 146.341
R17531 vdd.n1431 vdd.n1111 146.341
R17532 vdd.n1431 vdd.n1102 146.341
R17533 vdd.n1441 vdd.n1102 146.341
R17534 vdd.n1441 vdd.n1098 146.341
R17535 vdd.n1447 vdd.n1098 146.341
R17536 vdd.n1447 vdd.n1091 146.341
R17537 vdd.n1753 vdd.n1091 146.341
R17538 vdd.n1753 vdd.n1087 146.341
R17539 vdd.n1759 vdd.n1087 146.341
R17540 vdd.n1759 vdd.n1080 146.341
R17541 vdd.n1769 vdd.n1080 146.341
R17542 vdd.n1769 vdd.n1076 146.341
R17543 vdd.n1775 vdd.n1076 146.341
R17544 vdd.n1775 vdd.n1068 146.341
R17545 vdd.n1786 vdd.n1068 146.341
R17546 vdd.n1786 vdd.n1064 146.341
R17547 vdd.n1792 vdd.n1064 146.341
R17548 vdd.n1792 vdd.n1058 146.341
R17549 vdd.n1803 vdd.n1058 146.341
R17550 vdd.n1803 vdd.n1053 146.341
R17551 vdd.n1811 vdd.n1053 146.341
R17552 vdd.n1811 vdd.n1042 146.341
R17553 vdd.n2247 vdd.n1042 146.341
R17554 vdd.n1183 vdd.n1182 146.341
R17555 vdd.n1187 vdd.n1182 146.341
R17556 vdd.n1189 vdd.n1188 146.341
R17557 vdd.n1193 vdd.n1192 146.341
R17558 vdd.n1195 vdd.n1194 146.341
R17559 vdd.n1199 vdd.n1198 146.341
R17560 vdd.n1201 vdd.n1200 146.341
R17561 vdd.n1205 vdd.n1204 146.341
R17562 vdd.n1207 vdd.n1206 146.341
R17563 vdd.n1339 vdd.n1338 146.341
R17564 vdd.n1211 vdd.n1210 146.341
R17565 vdd.n1215 vdd.n1214 146.341
R17566 vdd.n1217 vdd.n1216 146.341
R17567 vdd.n1221 vdd.n1220 146.341
R17568 vdd.n1223 vdd.n1222 146.341
R17569 vdd.n1227 vdd.n1226 146.341
R17570 vdd.n1229 vdd.n1228 146.341
R17571 vdd.n1233 vdd.n1232 146.341
R17572 vdd.n1235 vdd.n1234 146.341
R17573 vdd.n1239 vdd.n1238 146.341
R17574 vdd.n1303 vdd.n1240 146.341
R17575 vdd.n1244 vdd.n1243 146.341
R17576 vdd.n1246 vdd.n1245 146.341
R17577 vdd.n1250 vdd.n1249 146.341
R17578 vdd.n1252 vdd.n1251 146.341
R17579 vdd.n1256 vdd.n1255 146.341
R17580 vdd.n1258 vdd.n1257 146.341
R17581 vdd.n1262 vdd.n1261 146.341
R17582 vdd.n1264 vdd.n1263 146.341
R17583 vdd.n1268 vdd.n1267 146.341
R17584 vdd.n1270 vdd.n1269 146.341
R17585 vdd.n1375 vdd.n1151 146.341
R17586 vdd.n1383 vdd.n1143 146.341
R17587 vdd.n1383 vdd.n1139 146.341
R17588 vdd.n1389 vdd.n1139 146.341
R17589 vdd.n1389 vdd.n1131 146.341
R17590 vdd.n1400 vdd.n1131 146.341
R17591 vdd.n1400 vdd.n1127 146.341
R17592 vdd.n1406 vdd.n1127 146.341
R17593 vdd.n1406 vdd.n1120 146.341
R17594 vdd.n1417 vdd.n1120 146.341
R17595 vdd.n1417 vdd.n1116 146.341
R17596 vdd.n1423 vdd.n1116 146.341
R17597 vdd.n1423 vdd.n1109 146.341
R17598 vdd.n1433 vdd.n1109 146.341
R17599 vdd.n1433 vdd.n1105 146.341
R17600 vdd.n1439 vdd.n1105 146.341
R17601 vdd.n1439 vdd.n1097 146.341
R17602 vdd.n1450 vdd.n1097 146.341
R17603 vdd.n1450 vdd.n1093 146.341
R17604 vdd.n1751 vdd.n1093 146.341
R17605 vdd.n1751 vdd.n1086 146.341
R17606 vdd.n1761 vdd.n1086 146.341
R17607 vdd.n1761 vdd.n1082 146.341
R17608 vdd.n1767 vdd.n1082 146.341
R17609 vdd.n1767 vdd.n1074 146.341
R17610 vdd.n1778 vdd.n1074 146.341
R17611 vdd.n1778 vdd.n1070 146.341
R17612 vdd.n1784 vdd.n1070 146.341
R17613 vdd.n1784 vdd.n1063 146.341
R17614 vdd.n1795 vdd.n1063 146.341
R17615 vdd.n1795 vdd.n1059 146.341
R17616 vdd.n1801 vdd.n1059 146.341
R17617 vdd.n1801 vdd.n1051 146.341
R17618 vdd.n1813 vdd.n1051 146.341
R17619 vdd.n1813 vdd.n1046 146.341
R17620 vdd.n2245 vdd.n1046 146.341
R17621 vdd.n1045 vdd.n1020 141.707
R17622 vdd.n756 vdd.n658 141.707
R17623 vdd.n2094 vdd.t217 127.284
R17624 vdd.n936 vdd.t201 127.284
R17625 vdd.n2068 vdd.t239 127.284
R17626 vdd.n928 vdd.t226 127.284
R17627 vdd.n2839 vdd.t188 127.284
R17628 vdd.n2839 vdd.t189 127.284
R17629 vdd.n2559 vdd.t224 127.284
R17630 vdd.n804 vdd.t205 127.284
R17631 vdd.n2556 vdd.t210 127.284
R17632 vdd.n768 vdd.t212 127.284
R17633 vdd.n998 vdd.t220 127.284
R17634 vdd.n998 vdd.t221 127.284
R17635 vdd.n22 vdd.n20 117.314
R17636 vdd.n17 vdd.n15 117.314
R17637 vdd.n27 vdd.n26 116.927
R17638 vdd.n24 vdd.n23 116.927
R17639 vdd.n22 vdd.n21 116.927
R17640 vdd.n17 vdd.n16 116.927
R17641 vdd.n19 vdd.n18 116.927
R17642 vdd.n27 vdd.n25 116.927
R17643 vdd.n2095 vdd.t216 111.188
R17644 vdd.n937 vdd.t202 111.188
R17645 vdd.n2069 vdd.t238 111.188
R17646 vdd.n929 vdd.t227 111.188
R17647 vdd.n2560 vdd.t223 111.188
R17648 vdd.n805 vdd.t206 111.188
R17649 vdd.n2557 vdd.t209 111.188
R17650 vdd.n769 vdd.t213 111.188
R17651 vdd.n2782 vdd.n882 99.5127
R17652 vdd.n2786 vdd.n882 99.5127
R17653 vdd.n2786 vdd.n874 99.5127
R17654 vdd.n2794 vdd.n874 99.5127
R17655 vdd.n2794 vdd.n872 99.5127
R17656 vdd.n2798 vdd.n872 99.5127
R17657 vdd.n2798 vdd.n861 99.5127
R17658 vdd.n2806 vdd.n861 99.5127
R17659 vdd.n2806 vdd.n859 99.5127
R17660 vdd.n2810 vdd.n859 99.5127
R17661 vdd.n2810 vdd.n850 99.5127
R17662 vdd.n2818 vdd.n850 99.5127
R17663 vdd.n2818 vdd.n848 99.5127
R17664 vdd.n2822 vdd.n848 99.5127
R17665 vdd.n2822 vdd.n838 99.5127
R17666 vdd.n2830 vdd.n838 99.5127
R17667 vdd.n2830 vdd.n836 99.5127
R17668 vdd.n2834 vdd.n836 99.5127
R17669 vdd.n2834 vdd.n827 99.5127
R17670 vdd.n2844 vdd.n827 99.5127
R17671 vdd.n2844 vdd.n825 99.5127
R17672 vdd.n2848 vdd.n825 99.5127
R17673 vdd.n2848 vdd.n813 99.5127
R17674 vdd.n2901 vdd.n813 99.5127
R17675 vdd.n2901 vdd.n811 99.5127
R17676 vdd.n2905 vdd.n811 99.5127
R17677 vdd.n2905 vdd.n777 99.5127
R17678 vdd.n2975 vdd.n777 99.5127
R17679 vdd.n2971 vdd.n778 99.5127
R17680 vdd.n2969 vdd.n2968 99.5127
R17681 vdd.n2966 vdd.n782 99.5127
R17682 vdd.n2962 vdd.n2961 99.5127
R17683 vdd.n2959 vdd.n785 99.5127
R17684 vdd.n2955 vdd.n2954 99.5127
R17685 vdd.n2952 vdd.n788 99.5127
R17686 vdd.n2948 vdd.n2947 99.5127
R17687 vdd.n2945 vdd.n791 99.5127
R17688 vdd.n2940 vdd.n2939 99.5127
R17689 vdd.n2937 vdd.n794 99.5127
R17690 vdd.n2933 vdd.n2932 99.5127
R17691 vdd.n2930 vdd.n797 99.5127
R17692 vdd.n2926 vdd.n2925 99.5127
R17693 vdd.n2923 vdd.n800 99.5127
R17694 vdd.n2919 vdd.n2918 99.5127
R17695 vdd.n2916 vdd.n803 99.5127
R17696 vdd.n2702 vdd.n885 99.5127
R17697 vdd.n2702 vdd.n880 99.5127
R17698 vdd.n2699 vdd.n880 99.5127
R17699 vdd.n2699 vdd.n875 99.5127
R17700 vdd.n2646 vdd.n875 99.5127
R17701 vdd.n2646 vdd.n869 99.5127
R17702 vdd.n2649 vdd.n869 99.5127
R17703 vdd.n2649 vdd.n862 99.5127
R17704 vdd.n2652 vdd.n862 99.5127
R17705 vdd.n2652 vdd.n857 99.5127
R17706 vdd.n2655 vdd.n857 99.5127
R17707 vdd.n2655 vdd.n852 99.5127
R17708 vdd.n2658 vdd.n852 99.5127
R17709 vdd.n2658 vdd.n846 99.5127
R17710 vdd.n2676 vdd.n846 99.5127
R17711 vdd.n2676 vdd.n839 99.5127
R17712 vdd.n2672 vdd.n839 99.5127
R17713 vdd.n2672 vdd.n834 99.5127
R17714 vdd.n2669 vdd.n834 99.5127
R17715 vdd.n2669 vdd.n829 99.5127
R17716 vdd.n2666 vdd.n829 99.5127
R17717 vdd.n2666 vdd.n823 99.5127
R17718 vdd.n2663 vdd.n823 99.5127
R17719 vdd.n2663 vdd.n815 99.5127
R17720 vdd.n815 vdd.n808 99.5127
R17721 vdd.n2907 vdd.n808 99.5127
R17722 vdd.n2908 vdd.n2907 99.5127
R17723 vdd.n2908 vdd.n775 99.5127
R17724 vdd.n2772 vdd.n2555 99.5127
R17725 vdd.n2768 vdd.n2555 99.5127
R17726 vdd.n2766 vdd.n2765 99.5127
R17727 vdd.n2762 vdd.n2761 99.5127
R17728 vdd.n2758 vdd.n2757 99.5127
R17729 vdd.n2754 vdd.n2753 99.5127
R17730 vdd.n2750 vdd.n2749 99.5127
R17731 vdd.n2746 vdd.n2745 99.5127
R17732 vdd.n2742 vdd.n2741 99.5127
R17733 vdd.n2738 vdd.n2737 99.5127
R17734 vdd.n2734 vdd.n2733 99.5127
R17735 vdd.n2730 vdd.n2729 99.5127
R17736 vdd.n2726 vdd.n2725 99.5127
R17737 vdd.n2722 vdd.n2721 99.5127
R17738 vdd.n2718 vdd.n2717 99.5127
R17739 vdd.n2714 vdd.n2713 99.5127
R17740 vdd.n2709 vdd.n2708 99.5127
R17741 vdd.n2520 vdd.n926 99.5127
R17742 vdd.n2516 vdd.n2515 99.5127
R17743 vdd.n2512 vdd.n2511 99.5127
R17744 vdd.n2508 vdd.n2507 99.5127
R17745 vdd.n2504 vdd.n2503 99.5127
R17746 vdd.n2500 vdd.n2499 99.5127
R17747 vdd.n2496 vdd.n2495 99.5127
R17748 vdd.n2492 vdd.n2491 99.5127
R17749 vdd.n2488 vdd.n2487 99.5127
R17750 vdd.n2484 vdd.n2483 99.5127
R17751 vdd.n2480 vdd.n2479 99.5127
R17752 vdd.n2476 vdd.n2475 99.5127
R17753 vdd.n2472 vdd.n2471 99.5127
R17754 vdd.n2468 vdd.n2467 99.5127
R17755 vdd.n2464 vdd.n2463 99.5127
R17756 vdd.n2460 vdd.n2459 99.5127
R17757 vdd.n2455 vdd.n2454 99.5127
R17758 vdd.n2193 vdd.n1021 99.5127
R17759 vdd.n2193 vdd.n1015 99.5127
R17760 vdd.n2190 vdd.n1015 99.5127
R17761 vdd.n2190 vdd.n1009 99.5127
R17762 vdd.n2187 vdd.n1009 99.5127
R17763 vdd.n2187 vdd.n1002 99.5127
R17764 vdd.n2184 vdd.n1002 99.5127
R17765 vdd.n2184 vdd.n995 99.5127
R17766 vdd.n2181 vdd.n995 99.5127
R17767 vdd.n2181 vdd.n990 99.5127
R17768 vdd.n2178 vdd.n990 99.5127
R17769 vdd.n2178 vdd.n984 99.5127
R17770 vdd.n2175 vdd.n984 99.5127
R17771 vdd.n2175 vdd.n977 99.5127
R17772 vdd.n2089 vdd.n977 99.5127
R17773 vdd.n2089 vdd.n971 99.5127
R17774 vdd.n2086 vdd.n971 99.5127
R17775 vdd.n2086 vdd.n966 99.5127
R17776 vdd.n2083 vdd.n966 99.5127
R17777 vdd.n2083 vdd.n961 99.5127
R17778 vdd.n2080 vdd.n961 99.5127
R17779 vdd.n2080 vdd.n955 99.5127
R17780 vdd.n2077 vdd.n955 99.5127
R17781 vdd.n2077 vdd.n948 99.5127
R17782 vdd.n2074 vdd.n948 99.5127
R17783 vdd.n2074 vdd.n941 99.5127
R17784 vdd.n941 vdd.n931 99.5127
R17785 vdd.n2450 vdd.n931 99.5127
R17786 vdd.n2028 vdd.n2026 99.5127
R17787 vdd.n2032 vdd.n2026 99.5127
R17788 vdd.n2036 vdd.n2034 99.5127
R17789 vdd.n2040 vdd.n2024 99.5127
R17790 vdd.n2044 vdd.n2042 99.5127
R17791 vdd.n2048 vdd.n2022 99.5127
R17792 vdd.n2052 vdd.n2050 99.5127
R17793 vdd.n2056 vdd.n2020 99.5127
R17794 vdd.n2059 vdd.n2058 99.5127
R17795 vdd.n2229 vdd.n2227 99.5127
R17796 vdd.n2225 vdd.n2061 99.5127
R17797 vdd.n2221 vdd.n2219 99.5127
R17798 vdd.n2217 vdd.n2063 99.5127
R17799 vdd.n2213 vdd.n2211 99.5127
R17800 vdd.n2209 vdd.n2065 99.5127
R17801 vdd.n2205 vdd.n2203 99.5127
R17802 vdd.n2201 vdd.n2067 99.5127
R17803 vdd.n2293 vdd.n1017 99.5127
R17804 vdd.n2297 vdd.n1017 99.5127
R17805 vdd.n2297 vdd.n1007 99.5127
R17806 vdd.n2305 vdd.n1007 99.5127
R17807 vdd.n2305 vdd.n1005 99.5127
R17808 vdd.n2309 vdd.n1005 99.5127
R17809 vdd.n2309 vdd.n994 99.5127
R17810 vdd.n2318 vdd.n994 99.5127
R17811 vdd.n2318 vdd.n992 99.5127
R17812 vdd.n2322 vdd.n992 99.5127
R17813 vdd.n2322 vdd.n982 99.5127
R17814 vdd.n2330 vdd.n982 99.5127
R17815 vdd.n2330 vdd.n980 99.5127
R17816 vdd.n2334 vdd.n980 99.5127
R17817 vdd.n2334 vdd.n970 99.5127
R17818 vdd.n2342 vdd.n970 99.5127
R17819 vdd.n2342 vdd.n968 99.5127
R17820 vdd.n2346 vdd.n968 99.5127
R17821 vdd.n2346 vdd.n959 99.5127
R17822 vdd.n2354 vdd.n959 99.5127
R17823 vdd.n2354 vdd.n957 99.5127
R17824 vdd.n2358 vdd.n957 99.5127
R17825 vdd.n2358 vdd.n946 99.5127
R17826 vdd.n2368 vdd.n946 99.5127
R17827 vdd.n2368 vdd.n943 99.5127
R17828 vdd.n2373 vdd.n943 99.5127
R17829 vdd.n2373 vdd.n944 99.5127
R17830 vdd.n944 vdd.n925 99.5127
R17831 vdd.n2891 vdd.n2890 99.5127
R17832 vdd.n2888 vdd.n2854 99.5127
R17833 vdd.n2884 vdd.n2883 99.5127
R17834 vdd.n2881 vdd.n2857 99.5127
R17835 vdd.n2877 vdd.n2876 99.5127
R17836 vdd.n2874 vdd.n2860 99.5127
R17837 vdd.n2870 vdd.n2869 99.5127
R17838 vdd.n2867 vdd.n2864 99.5127
R17839 vdd.n3008 vdd.n755 99.5127
R17840 vdd.n3006 vdd.n3005 99.5127
R17841 vdd.n3003 vdd.n758 99.5127
R17842 vdd.n2999 vdd.n2998 99.5127
R17843 vdd.n2996 vdd.n761 99.5127
R17844 vdd.n2992 vdd.n2991 99.5127
R17845 vdd.n2989 vdd.n764 99.5127
R17846 vdd.n2985 vdd.n2984 99.5127
R17847 vdd.n2982 vdd.n767 99.5127
R17848 vdd.n2626 vdd.n886 99.5127
R17849 vdd.n2626 vdd.n881 99.5127
R17850 vdd.n2697 vdd.n881 99.5127
R17851 vdd.n2697 vdd.n876 99.5127
R17852 vdd.n2693 vdd.n876 99.5127
R17853 vdd.n2693 vdd.n870 99.5127
R17854 vdd.n2690 vdd.n870 99.5127
R17855 vdd.n2690 vdd.n863 99.5127
R17856 vdd.n2687 vdd.n863 99.5127
R17857 vdd.n2687 vdd.n858 99.5127
R17858 vdd.n2684 vdd.n858 99.5127
R17859 vdd.n2684 vdd.n853 99.5127
R17860 vdd.n2681 vdd.n853 99.5127
R17861 vdd.n2681 vdd.n847 99.5127
R17862 vdd.n2678 vdd.n847 99.5127
R17863 vdd.n2678 vdd.n840 99.5127
R17864 vdd.n2643 vdd.n840 99.5127
R17865 vdd.n2643 vdd.n835 99.5127
R17866 vdd.n2640 vdd.n835 99.5127
R17867 vdd.n2640 vdd.n830 99.5127
R17868 vdd.n2637 vdd.n830 99.5127
R17869 vdd.n2637 vdd.n824 99.5127
R17870 vdd.n2634 vdd.n824 99.5127
R17871 vdd.n2634 vdd.n816 99.5127
R17872 vdd.n2631 vdd.n816 99.5127
R17873 vdd.n2631 vdd.n809 99.5127
R17874 vdd.n809 vdd.n773 99.5127
R17875 vdd.n2977 vdd.n773 99.5127
R17876 vdd.n2776 vdd.n889 99.5127
R17877 vdd.n2564 vdd.n2563 99.5127
R17878 vdd.n2568 vdd.n2567 99.5127
R17879 vdd.n2572 vdd.n2571 99.5127
R17880 vdd.n2576 vdd.n2575 99.5127
R17881 vdd.n2580 vdd.n2579 99.5127
R17882 vdd.n2584 vdd.n2583 99.5127
R17883 vdd.n2588 vdd.n2587 99.5127
R17884 vdd.n2592 vdd.n2591 99.5127
R17885 vdd.n2596 vdd.n2595 99.5127
R17886 vdd.n2600 vdd.n2599 99.5127
R17887 vdd.n2604 vdd.n2603 99.5127
R17888 vdd.n2608 vdd.n2607 99.5127
R17889 vdd.n2612 vdd.n2611 99.5127
R17890 vdd.n2616 vdd.n2615 99.5127
R17891 vdd.n2620 vdd.n2619 99.5127
R17892 vdd.n2622 vdd.n2554 99.5127
R17893 vdd.n2780 vdd.n879 99.5127
R17894 vdd.n2788 vdd.n879 99.5127
R17895 vdd.n2788 vdd.n877 99.5127
R17896 vdd.n2792 vdd.n877 99.5127
R17897 vdd.n2792 vdd.n867 99.5127
R17898 vdd.n2800 vdd.n867 99.5127
R17899 vdd.n2800 vdd.n865 99.5127
R17900 vdd.n2804 vdd.n865 99.5127
R17901 vdd.n2804 vdd.n856 99.5127
R17902 vdd.n2812 vdd.n856 99.5127
R17903 vdd.n2812 vdd.n854 99.5127
R17904 vdd.n2816 vdd.n854 99.5127
R17905 vdd.n2816 vdd.n844 99.5127
R17906 vdd.n2824 vdd.n844 99.5127
R17907 vdd.n2824 vdd.n842 99.5127
R17908 vdd.n2828 vdd.n842 99.5127
R17909 vdd.n2828 vdd.n833 99.5127
R17910 vdd.n2836 vdd.n833 99.5127
R17911 vdd.n2836 vdd.n831 99.5127
R17912 vdd.n2842 vdd.n831 99.5127
R17913 vdd.n2842 vdd.n821 99.5127
R17914 vdd.n2850 vdd.n821 99.5127
R17915 vdd.n2850 vdd.n818 99.5127
R17916 vdd.n2899 vdd.n818 99.5127
R17917 vdd.n2899 vdd.n819 99.5127
R17918 vdd.n819 vdd.n810 99.5127
R17919 vdd.n2894 vdd.n810 99.5127
R17920 vdd.n2894 vdd.n776 99.5127
R17921 vdd.n2444 vdd.n2443 99.5127
R17922 vdd.n2440 vdd.n2439 99.5127
R17923 vdd.n2436 vdd.n2435 99.5127
R17924 vdd.n2432 vdd.n2431 99.5127
R17925 vdd.n2428 vdd.n2427 99.5127
R17926 vdd.n2424 vdd.n2423 99.5127
R17927 vdd.n2420 vdd.n2419 99.5127
R17928 vdd.n2416 vdd.n2415 99.5127
R17929 vdd.n2412 vdd.n2411 99.5127
R17930 vdd.n2408 vdd.n2407 99.5127
R17931 vdd.n2404 vdd.n2403 99.5127
R17932 vdd.n2400 vdd.n2399 99.5127
R17933 vdd.n2396 vdd.n2395 99.5127
R17934 vdd.n2392 vdd.n2391 99.5127
R17935 vdd.n2388 vdd.n2387 99.5127
R17936 vdd.n2384 vdd.n2383 99.5127
R17937 vdd.n2380 vdd.n907 99.5127
R17938 vdd.n2137 vdd.n1022 99.5127
R17939 vdd.n2137 vdd.n1016 99.5127
R17940 vdd.n2140 vdd.n1016 99.5127
R17941 vdd.n2140 vdd.n1010 99.5127
R17942 vdd.n2143 vdd.n1010 99.5127
R17943 vdd.n2143 vdd.n1003 99.5127
R17944 vdd.n2146 vdd.n1003 99.5127
R17945 vdd.n2146 vdd.n996 99.5127
R17946 vdd.n2149 vdd.n996 99.5127
R17947 vdd.n2149 vdd.n991 99.5127
R17948 vdd.n2152 vdd.n991 99.5127
R17949 vdd.n2152 vdd.n985 99.5127
R17950 vdd.n2173 vdd.n985 99.5127
R17951 vdd.n2173 vdd.n978 99.5127
R17952 vdd.n2169 vdd.n978 99.5127
R17953 vdd.n2169 vdd.n972 99.5127
R17954 vdd.n2166 vdd.n972 99.5127
R17955 vdd.n2166 vdd.n967 99.5127
R17956 vdd.n2163 vdd.n967 99.5127
R17957 vdd.n2163 vdd.n962 99.5127
R17958 vdd.n2160 vdd.n962 99.5127
R17959 vdd.n2160 vdd.n956 99.5127
R17960 vdd.n2157 vdd.n956 99.5127
R17961 vdd.n2157 vdd.n949 99.5127
R17962 vdd.n949 vdd.n940 99.5127
R17963 vdd.n2375 vdd.n940 99.5127
R17964 vdd.n2376 vdd.n2375 99.5127
R17965 vdd.n2376 vdd.n932 99.5127
R17966 vdd.n2287 vdd.n2285 99.5127
R17967 vdd.n2283 vdd.n1025 99.5127
R17968 vdd.n2279 vdd.n2277 99.5127
R17969 vdd.n2275 vdd.n1027 99.5127
R17970 vdd.n2271 vdd.n2269 99.5127
R17971 vdd.n2267 vdd.n1029 99.5127
R17972 vdd.n2263 vdd.n2261 99.5127
R17973 vdd.n2259 vdd.n1031 99.5127
R17974 vdd.n2101 vdd.n1033 99.5127
R17975 vdd.n2106 vdd.n2103 99.5127
R17976 vdd.n2110 vdd.n2108 99.5127
R17977 vdd.n2114 vdd.n2099 99.5127
R17978 vdd.n2118 vdd.n2116 99.5127
R17979 vdd.n2122 vdd.n2097 99.5127
R17980 vdd.n2126 vdd.n2124 99.5127
R17981 vdd.n2131 vdd.n2093 99.5127
R17982 vdd.n2134 vdd.n2133 99.5127
R17983 vdd.n2291 vdd.n1013 99.5127
R17984 vdd.n2299 vdd.n1013 99.5127
R17985 vdd.n2299 vdd.n1011 99.5127
R17986 vdd.n2303 vdd.n1011 99.5127
R17987 vdd.n2303 vdd.n1000 99.5127
R17988 vdd.n2311 vdd.n1000 99.5127
R17989 vdd.n2311 vdd.n997 99.5127
R17990 vdd.n2316 vdd.n997 99.5127
R17991 vdd.n2316 vdd.n988 99.5127
R17992 vdd.n2324 vdd.n988 99.5127
R17993 vdd.n2324 vdd.n986 99.5127
R17994 vdd.n2328 vdd.n986 99.5127
R17995 vdd.n2328 vdd.n976 99.5127
R17996 vdd.n2336 vdd.n976 99.5127
R17997 vdd.n2336 vdd.n974 99.5127
R17998 vdd.n2340 vdd.n974 99.5127
R17999 vdd.n2340 vdd.n965 99.5127
R18000 vdd.n2348 vdd.n965 99.5127
R18001 vdd.n2348 vdd.n963 99.5127
R18002 vdd.n2352 vdd.n963 99.5127
R18003 vdd.n2352 vdd.n953 99.5127
R18004 vdd.n2360 vdd.n953 99.5127
R18005 vdd.n2360 vdd.n950 99.5127
R18006 vdd.n2366 vdd.n950 99.5127
R18007 vdd.n2366 vdd.n951 99.5127
R18008 vdd.n951 vdd.n942 99.5127
R18009 vdd.n942 vdd.n933 99.5127
R18010 vdd.n2448 vdd.n933 99.5127
R18011 vdd.n9 vdd.n7 98.9633
R18012 vdd.n2 vdd.n0 98.9633
R18013 vdd.n9 vdd.n8 98.6055
R18014 vdd.n11 vdd.n10 98.6055
R18015 vdd.n13 vdd.n12 98.6055
R18016 vdd.n6 vdd.n5 98.6055
R18017 vdd.n4 vdd.n3 98.6055
R18018 vdd.n2 vdd.n1 98.6055
R18019 vdd.t124 vdd.n291 85.8723
R18020 vdd.t98 vdd.n236 85.8723
R18021 vdd.t110 vdd.n193 85.8723
R18022 vdd.t87 vdd.n138 85.8723
R18023 vdd.t42 vdd.n96 85.8723
R18024 vdd.t22 vdd.n41 85.8723
R18025 vdd.t137 vdd.n1660 85.8723
R18026 vdd.t48 vdd.n1715 85.8723
R18027 vdd.t122 vdd.n1562 85.8723
R18028 vdd.t32 vdd.n1617 85.8723
R18029 vdd.t20 vdd.n1465 85.8723
R18030 vdd.t45 vdd.n1520 85.8723
R18031 vdd.n2840 vdd.n2839 78.546
R18032 vdd.n2314 vdd.n998 78.546
R18033 vdd.n278 vdd.n277 75.1835
R18034 vdd.n276 vdd.n275 75.1835
R18035 vdd.n274 vdd.n273 75.1835
R18036 vdd.n272 vdd.n271 75.1835
R18037 vdd.n270 vdd.n269 75.1835
R18038 vdd.n268 vdd.n267 75.1835
R18039 vdd.n266 vdd.n265 75.1835
R18040 vdd.n180 vdd.n179 75.1835
R18041 vdd.n178 vdd.n177 75.1835
R18042 vdd.n176 vdd.n175 75.1835
R18043 vdd.n174 vdd.n173 75.1835
R18044 vdd.n172 vdd.n171 75.1835
R18045 vdd.n170 vdd.n169 75.1835
R18046 vdd.n168 vdd.n167 75.1835
R18047 vdd.n83 vdd.n82 75.1835
R18048 vdd.n81 vdd.n80 75.1835
R18049 vdd.n79 vdd.n78 75.1835
R18050 vdd.n77 vdd.n76 75.1835
R18051 vdd.n75 vdd.n74 75.1835
R18052 vdd.n73 vdd.n72 75.1835
R18053 vdd.n71 vdd.n70 75.1835
R18054 vdd.n1690 vdd.n1689 75.1835
R18055 vdd.n1692 vdd.n1691 75.1835
R18056 vdd.n1694 vdd.n1693 75.1835
R18057 vdd.n1696 vdd.n1695 75.1835
R18058 vdd.n1698 vdd.n1697 75.1835
R18059 vdd.n1700 vdd.n1699 75.1835
R18060 vdd.n1702 vdd.n1701 75.1835
R18061 vdd.n1592 vdd.n1591 75.1835
R18062 vdd.n1594 vdd.n1593 75.1835
R18063 vdd.n1596 vdd.n1595 75.1835
R18064 vdd.n1598 vdd.n1597 75.1835
R18065 vdd.n1600 vdd.n1599 75.1835
R18066 vdd.n1602 vdd.n1601 75.1835
R18067 vdd.n1604 vdd.n1603 75.1835
R18068 vdd.n1495 vdd.n1494 75.1835
R18069 vdd.n1497 vdd.n1496 75.1835
R18070 vdd.n1499 vdd.n1498 75.1835
R18071 vdd.n1501 vdd.n1500 75.1835
R18072 vdd.n1503 vdd.n1502 75.1835
R18073 vdd.n1505 vdd.n1504 75.1835
R18074 vdd.n1507 vdd.n1506 75.1835
R18075 vdd.n2775 vdd.n2774 72.8958
R18076 vdd.n2774 vdd.n2538 72.8958
R18077 vdd.n2774 vdd.n2539 72.8958
R18078 vdd.n2774 vdd.n2540 72.8958
R18079 vdd.n2774 vdd.n2541 72.8958
R18080 vdd.n2774 vdd.n2542 72.8958
R18081 vdd.n2774 vdd.n2543 72.8958
R18082 vdd.n2774 vdd.n2544 72.8958
R18083 vdd.n2774 vdd.n2545 72.8958
R18084 vdd.n2774 vdd.n2546 72.8958
R18085 vdd.n2774 vdd.n2547 72.8958
R18086 vdd.n2774 vdd.n2548 72.8958
R18087 vdd.n2774 vdd.n2549 72.8958
R18088 vdd.n2774 vdd.n2550 72.8958
R18089 vdd.n2774 vdd.n2551 72.8958
R18090 vdd.n2774 vdd.n2552 72.8958
R18091 vdd.n2774 vdd.n2553 72.8958
R18092 vdd.n772 vdd.n756 72.8958
R18093 vdd.n2983 vdd.n756 72.8958
R18094 vdd.n766 vdd.n756 72.8958
R18095 vdd.n2990 vdd.n756 72.8958
R18096 vdd.n763 vdd.n756 72.8958
R18097 vdd.n2997 vdd.n756 72.8958
R18098 vdd.n760 vdd.n756 72.8958
R18099 vdd.n3004 vdd.n756 72.8958
R18100 vdd.n3007 vdd.n756 72.8958
R18101 vdd.n2863 vdd.n756 72.8958
R18102 vdd.n2868 vdd.n756 72.8958
R18103 vdd.n2862 vdd.n756 72.8958
R18104 vdd.n2875 vdd.n756 72.8958
R18105 vdd.n2859 vdd.n756 72.8958
R18106 vdd.n2882 vdd.n756 72.8958
R18107 vdd.n2856 vdd.n756 72.8958
R18108 vdd.n2889 vdd.n756 72.8958
R18109 vdd.n2027 vdd.n1020 72.8958
R18110 vdd.n2033 vdd.n1020 72.8958
R18111 vdd.n2035 vdd.n1020 72.8958
R18112 vdd.n2041 vdd.n1020 72.8958
R18113 vdd.n2043 vdd.n1020 72.8958
R18114 vdd.n2049 vdd.n1020 72.8958
R18115 vdd.n2051 vdd.n1020 72.8958
R18116 vdd.n2057 vdd.n1020 72.8958
R18117 vdd.n2228 vdd.n1020 72.8958
R18118 vdd.n2226 vdd.n1020 72.8958
R18119 vdd.n2220 vdd.n1020 72.8958
R18120 vdd.n2218 vdd.n1020 72.8958
R18121 vdd.n2212 vdd.n1020 72.8958
R18122 vdd.n2210 vdd.n1020 72.8958
R18123 vdd.n2204 vdd.n1020 72.8958
R18124 vdd.n2202 vdd.n1020 72.8958
R18125 vdd.n2196 vdd.n1020 72.8958
R18126 vdd.n2521 vdd.n908 72.8958
R18127 vdd.n2521 vdd.n909 72.8958
R18128 vdd.n2521 vdd.n910 72.8958
R18129 vdd.n2521 vdd.n911 72.8958
R18130 vdd.n2521 vdd.n912 72.8958
R18131 vdd.n2521 vdd.n913 72.8958
R18132 vdd.n2521 vdd.n914 72.8958
R18133 vdd.n2521 vdd.n915 72.8958
R18134 vdd.n2521 vdd.n916 72.8958
R18135 vdd.n2521 vdd.n917 72.8958
R18136 vdd.n2521 vdd.n918 72.8958
R18137 vdd.n2521 vdd.n919 72.8958
R18138 vdd.n2521 vdd.n920 72.8958
R18139 vdd.n2521 vdd.n921 72.8958
R18140 vdd.n2521 vdd.n922 72.8958
R18141 vdd.n2521 vdd.n923 72.8958
R18142 vdd.n2521 vdd.n924 72.8958
R18143 vdd.n2774 vdd.n2773 72.8958
R18144 vdd.n2774 vdd.n2522 72.8958
R18145 vdd.n2774 vdd.n2523 72.8958
R18146 vdd.n2774 vdd.n2524 72.8958
R18147 vdd.n2774 vdd.n2525 72.8958
R18148 vdd.n2774 vdd.n2526 72.8958
R18149 vdd.n2774 vdd.n2527 72.8958
R18150 vdd.n2774 vdd.n2528 72.8958
R18151 vdd.n2774 vdd.n2529 72.8958
R18152 vdd.n2774 vdd.n2530 72.8958
R18153 vdd.n2774 vdd.n2531 72.8958
R18154 vdd.n2774 vdd.n2532 72.8958
R18155 vdd.n2774 vdd.n2533 72.8958
R18156 vdd.n2774 vdd.n2534 72.8958
R18157 vdd.n2774 vdd.n2535 72.8958
R18158 vdd.n2774 vdd.n2536 72.8958
R18159 vdd.n2774 vdd.n2537 72.8958
R18160 vdd.n2911 vdd.n756 72.8958
R18161 vdd.n2917 vdd.n756 72.8958
R18162 vdd.n802 vdd.n756 72.8958
R18163 vdd.n2924 vdd.n756 72.8958
R18164 vdd.n799 vdd.n756 72.8958
R18165 vdd.n2931 vdd.n756 72.8958
R18166 vdd.n796 vdd.n756 72.8958
R18167 vdd.n2938 vdd.n756 72.8958
R18168 vdd.n793 vdd.n756 72.8958
R18169 vdd.n2946 vdd.n756 72.8958
R18170 vdd.n790 vdd.n756 72.8958
R18171 vdd.n2953 vdd.n756 72.8958
R18172 vdd.n787 vdd.n756 72.8958
R18173 vdd.n2960 vdd.n756 72.8958
R18174 vdd.n784 vdd.n756 72.8958
R18175 vdd.n2967 vdd.n756 72.8958
R18176 vdd.n2970 vdd.n756 72.8958
R18177 vdd.n2521 vdd.n906 72.8958
R18178 vdd.n2521 vdd.n905 72.8958
R18179 vdd.n2521 vdd.n904 72.8958
R18180 vdd.n2521 vdd.n903 72.8958
R18181 vdd.n2521 vdd.n902 72.8958
R18182 vdd.n2521 vdd.n901 72.8958
R18183 vdd.n2521 vdd.n900 72.8958
R18184 vdd.n2521 vdd.n899 72.8958
R18185 vdd.n2521 vdd.n898 72.8958
R18186 vdd.n2521 vdd.n897 72.8958
R18187 vdd.n2521 vdd.n896 72.8958
R18188 vdd.n2521 vdd.n895 72.8958
R18189 vdd.n2521 vdd.n894 72.8958
R18190 vdd.n2521 vdd.n893 72.8958
R18191 vdd.n2521 vdd.n892 72.8958
R18192 vdd.n2521 vdd.n891 72.8958
R18193 vdd.n2521 vdd.n890 72.8958
R18194 vdd.n2286 vdd.n1020 72.8958
R18195 vdd.n2284 vdd.n1020 72.8958
R18196 vdd.n2278 vdd.n1020 72.8958
R18197 vdd.n2276 vdd.n1020 72.8958
R18198 vdd.n2270 vdd.n1020 72.8958
R18199 vdd.n2268 vdd.n1020 72.8958
R18200 vdd.n2262 vdd.n1020 72.8958
R18201 vdd.n2260 vdd.n1020 72.8958
R18202 vdd.n1032 vdd.n1020 72.8958
R18203 vdd.n2102 vdd.n1020 72.8958
R18204 vdd.n2107 vdd.n1020 72.8958
R18205 vdd.n2109 vdd.n1020 72.8958
R18206 vdd.n2115 vdd.n1020 72.8958
R18207 vdd.n2117 vdd.n1020 72.8958
R18208 vdd.n2123 vdd.n1020 72.8958
R18209 vdd.n2125 vdd.n1020 72.8958
R18210 vdd.n2132 vdd.n1020 72.8958
R18211 vdd.n1374 vdd.n1373 66.2847
R18212 vdd.n1374 vdd.n1152 66.2847
R18213 vdd.n1374 vdd.n1153 66.2847
R18214 vdd.n1374 vdd.n1154 66.2847
R18215 vdd.n1374 vdd.n1155 66.2847
R18216 vdd.n1374 vdd.n1156 66.2847
R18217 vdd.n1374 vdd.n1157 66.2847
R18218 vdd.n1374 vdd.n1158 66.2847
R18219 vdd.n1374 vdd.n1159 66.2847
R18220 vdd.n1374 vdd.n1160 66.2847
R18221 vdd.n1374 vdd.n1161 66.2847
R18222 vdd.n1374 vdd.n1162 66.2847
R18223 vdd.n1374 vdd.n1163 66.2847
R18224 vdd.n1374 vdd.n1164 66.2847
R18225 vdd.n1374 vdd.n1165 66.2847
R18226 vdd.n1374 vdd.n1166 66.2847
R18227 vdd.n1374 vdd.n1167 66.2847
R18228 vdd.n1374 vdd.n1168 66.2847
R18229 vdd.n1374 vdd.n1169 66.2847
R18230 vdd.n1374 vdd.n1170 66.2847
R18231 vdd.n1374 vdd.n1171 66.2847
R18232 vdd.n1374 vdd.n1172 66.2847
R18233 vdd.n1374 vdd.n1173 66.2847
R18234 vdd.n1374 vdd.n1174 66.2847
R18235 vdd.n1374 vdd.n1175 66.2847
R18236 vdd.n1374 vdd.n1176 66.2847
R18237 vdd.n1374 vdd.n1177 66.2847
R18238 vdd.n1374 vdd.n1178 66.2847
R18239 vdd.n1374 vdd.n1179 66.2847
R18240 vdd.n1374 vdd.n1180 66.2847
R18241 vdd.n1374 vdd.n1181 66.2847
R18242 vdd.n1045 vdd.n1041 66.2847
R18243 vdd.n1917 vdd.n1045 66.2847
R18244 vdd.n1922 vdd.n1045 66.2847
R18245 vdd.n1927 vdd.n1045 66.2847
R18246 vdd.n1915 vdd.n1045 66.2847
R18247 vdd.n1934 vdd.n1045 66.2847
R18248 vdd.n1907 vdd.n1045 66.2847
R18249 vdd.n1941 vdd.n1045 66.2847
R18250 vdd.n1900 vdd.n1045 66.2847
R18251 vdd.n1948 vdd.n1045 66.2847
R18252 vdd.n1894 vdd.n1045 66.2847
R18253 vdd.n1889 vdd.n1045 66.2847
R18254 vdd.n1959 vdd.n1045 66.2847
R18255 vdd.n1881 vdd.n1045 66.2847
R18256 vdd.n1966 vdd.n1045 66.2847
R18257 vdd.n1874 vdd.n1045 66.2847
R18258 vdd.n1973 vdd.n1045 66.2847
R18259 vdd.n1867 vdd.n1045 66.2847
R18260 vdd.n1980 vdd.n1045 66.2847
R18261 vdd.n1860 vdd.n1045 66.2847
R18262 vdd.n1987 vdd.n1045 66.2847
R18263 vdd.n1854 vdd.n1045 66.2847
R18264 vdd.n1849 vdd.n1045 66.2847
R18265 vdd.n1998 vdd.n1045 66.2847
R18266 vdd.n1841 vdd.n1045 66.2847
R18267 vdd.n2005 vdd.n1045 66.2847
R18268 vdd.n1834 vdd.n1045 66.2847
R18269 vdd.n2012 vdd.n1045 66.2847
R18270 vdd.n2015 vdd.n1045 66.2847
R18271 vdd.n1825 vdd.n1045 66.2847
R18272 vdd.n2237 vdd.n1045 66.2847
R18273 vdd.n1819 vdd.n1045 66.2847
R18274 vdd.n3137 vdd.n658 66.2847
R18275 vdd.n663 vdd.n658 66.2847
R18276 vdd.n666 vdd.n658 66.2847
R18277 vdd.n3126 vdd.n658 66.2847
R18278 vdd.n3120 vdd.n658 66.2847
R18279 vdd.n3118 vdd.n658 66.2847
R18280 vdd.n3112 vdd.n658 66.2847
R18281 vdd.n3110 vdd.n658 66.2847
R18282 vdd.n3104 vdd.n658 66.2847
R18283 vdd.n3102 vdd.n658 66.2847
R18284 vdd.n3096 vdd.n658 66.2847
R18285 vdd.n3094 vdd.n658 66.2847
R18286 vdd.n3088 vdd.n658 66.2847
R18287 vdd.n3086 vdd.n658 66.2847
R18288 vdd.n3080 vdd.n658 66.2847
R18289 vdd.n3078 vdd.n658 66.2847
R18290 vdd.n3072 vdd.n658 66.2847
R18291 vdd.n3070 vdd.n658 66.2847
R18292 vdd.n3064 vdd.n658 66.2847
R18293 vdd.n3062 vdd.n658 66.2847
R18294 vdd.n727 vdd.n658 66.2847
R18295 vdd.n3053 vdd.n658 66.2847
R18296 vdd.n729 vdd.n658 66.2847
R18297 vdd.n3046 vdd.n658 66.2847
R18298 vdd.n3040 vdd.n658 66.2847
R18299 vdd.n3038 vdd.n658 66.2847
R18300 vdd.n3032 vdd.n658 66.2847
R18301 vdd.n3030 vdd.n658 66.2847
R18302 vdd.n3024 vdd.n658 66.2847
R18303 vdd.n750 vdd.n658 66.2847
R18304 vdd.n752 vdd.n658 66.2847
R18305 vdd.n3253 vdd.n3252 66.2847
R18306 vdd.n3253 vdd.n403 66.2847
R18307 vdd.n3253 vdd.n402 66.2847
R18308 vdd.n3253 vdd.n401 66.2847
R18309 vdd.n3253 vdd.n400 66.2847
R18310 vdd.n3253 vdd.n399 66.2847
R18311 vdd.n3253 vdd.n398 66.2847
R18312 vdd.n3253 vdd.n397 66.2847
R18313 vdd.n3253 vdd.n396 66.2847
R18314 vdd.n3253 vdd.n395 66.2847
R18315 vdd.n3253 vdd.n394 66.2847
R18316 vdd.n3253 vdd.n393 66.2847
R18317 vdd.n3253 vdd.n392 66.2847
R18318 vdd.n3253 vdd.n391 66.2847
R18319 vdd.n3253 vdd.n390 66.2847
R18320 vdd.n3253 vdd.n389 66.2847
R18321 vdd.n3253 vdd.n388 66.2847
R18322 vdd.n3253 vdd.n387 66.2847
R18323 vdd.n3253 vdd.n386 66.2847
R18324 vdd.n3253 vdd.n385 66.2847
R18325 vdd.n3253 vdd.n384 66.2847
R18326 vdd.n3253 vdd.n383 66.2847
R18327 vdd.n3253 vdd.n382 66.2847
R18328 vdd.n3253 vdd.n381 66.2847
R18329 vdd.n3253 vdd.n380 66.2847
R18330 vdd.n3253 vdd.n379 66.2847
R18331 vdd.n3253 vdd.n378 66.2847
R18332 vdd.n3253 vdd.n377 66.2847
R18333 vdd.n3253 vdd.n376 66.2847
R18334 vdd.n3253 vdd.n375 66.2847
R18335 vdd.n3253 vdd.n374 66.2847
R18336 vdd.n3253 vdd.n373 66.2847
R18337 vdd.n448 vdd.n373 52.4337
R18338 vdd.n454 vdd.n374 52.4337
R18339 vdd.n458 vdd.n375 52.4337
R18340 vdd.n464 vdd.n376 52.4337
R18341 vdd.n468 vdd.n377 52.4337
R18342 vdd.n474 vdd.n378 52.4337
R18343 vdd.n478 vdd.n379 52.4337
R18344 vdd.n484 vdd.n380 52.4337
R18345 vdd.n488 vdd.n381 52.4337
R18346 vdd.n494 vdd.n382 52.4337
R18347 vdd.n498 vdd.n383 52.4337
R18348 vdd.n504 vdd.n384 52.4337
R18349 vdd.n508 vdd.n385 52.4337
R18350 vdd.n514 vdd.n386 52.4337
R18351 vdd.n518 vdd.n387 52.4337
R18352 vdd.n524 vdd.n388 52.4337
R18353 vdd.n528 vdd.n389 52.4337
R18354 vdd.n534 vdd.n390 52.4337
R18355 vdd.n538 vdd.n391 52.4337
R18356 vdd.n544 vdd.n392 52.4337
R18357 vdd.n548 vdd.n393 52.4337
R18358 vdd.n554 vdd.n394 52.4337
R18359 vdd.n558 vdd.n395 52.4337
R18360 vdd.n564 vdd.n396 52.4337
R18361 vdd.n568 vdd.n397 52.4337
R18362 vdd.n574 vdd.n398 52.4337
R18363 vdd.n578 vdd.n399 52.4337
R18364 vdd.n584 vdd.n400 52.4337
R18365 vdd.n588 vdd.n401 52.4337
R18366 vdd.n594 vdd.n402 52.4337
R18367 vdd.n597 vdd.n403 52.4337
R18368 vdd.n3252 vdd.n3251 52.4337
R18369 vdd.n3137 vdd.n660 52.4337
R18370 vdd.n3135 vdd.n663 52.4337
R18371 vdd.n3131 vdd.n666 52.4337
R18372 vdd.n3127 vdd.n3126 52.4337
R18373 vdd.n3120 vdd.n669 52.4337
R18374 vdd.n3119 vdd.n3118 52.4337
R18375 vdd.n3112 vdd.n675 52.4337
R18376 vdd.n3111 vdd.n3110 52.4337
R18377 vdd.n3104 vdd.n681 52.4337
R18378 vdd.n3103 vdd.n3102 52.4337
R18379 vdd.n3096 vdd.n689 52.4337
R18380 vdd.n3095 vdd.n3094 52.4337
R18381 vdd.n3088 vdd.n695 52.4337
R18382 vdd.n3087 vdd.n3086 52.4337
R18383 vdd.n3080 vdd.n701 52.4337
R18384 vdd.n3079 vdd.n3078 52.4337
R18385 vdd.n3072 vdd.n707 52.4337
R18386 vdd.n3071 vdd.n3070 52.4337
R18387 vdd.n3064 vdd.n713 52.4337
R18388 vdd.n3063 vdd.n3062 52.4337
R18389 vdd.n727 vdd.n719 52.4337
R18390 vdd.n3054 vdd.n3053 52.4337
R18391 vdd.n3051 vdd.n729 52.4337
R18392 vdd.n3047 vdd.n3046 52.4337
R18393 vdd.n3040 vdd.n733 52.4337
R18394 vdd.n3039 vdd.n3038 52.4337
R18395 vdd.n3032 vdd.n739 52.4337
R18396 vdd.n3031 vdd.n3030 52.4337
R18397 vdd.n3024 vdd.n745 52.4337
R18398 vdd.n3023 vdd.n750 52.4337
R18399 vdd.n3019 vdd.n752 52.4337
R18400 vdd.n2239 vdd.n1819 52.4337
R18401 vdd.n2237 vdd.n2236 52.4337
R18402 vdd.n1826 vdd.n1825 52.4337
R18403 vdd.n2015 vdd.n2014 52.4337
R18404 vdd.n2012 vdd.n2011 52.4337
R18405 vdd.n2007 vdd.n1834 52.4337
R18406 vdd.n2005 vdd.n2004 52.4337
R18407 vdd.n2000 vdd.n1841 52.4337
R18408 vdd.n1998 vdd.n1997 52.4337
R18409 vdd.n1850 vdd.n1849 52.4337
R18410 vdd.n1989 vdd.n1854 52.4337
R18411 vdd.n1987 vdd.n1986 52.4337
R18412 vdd.n1982 vdd.n1860 52.4337
R18413 vdd.n1980 vdd.n1979 52.4337
R18414 vdd.n1975 vdd.n1867 52.4337
R18415 vdd.n1973 vdd.n1972 52.4337
R18416 vdd.n1968 vdd.n1874 52.4337
R18417 vdd.n1966 vdd.n1965 52.4337
R18418 vdd.n1961 vdd.n1881 52.4337
R18419 vdd.n1959 vdd.n1958 52.4337
R18420 vdd.n1890 vdd.n1889 52.4337
R18421 vdd.n1950 vdd.n1894 52.4337
R18422 vdd.n1948 vdd.n1947 52.4337
R18423 vdd.n1943 vdd.n1900 52.4337
R18424 vdd.n1941 vdd.n1940 52.4337
R18425 vdd.n1936 vdd.n1907 52.4337
R18426 vdd.n1934 vdd.n1933 52.4337
R18427 vdd.n1929 vdd.n1915 52.4337
R18428 vdd.n1927 vdd.n1926 52.4337
R18429 vdd.n1922 vdd.n1921 52.4337
R18430 vdd.n1917 vdd.n1916 52.4337
R18431 vdd.n2248 vdd.n1041 52.4337
R18432 vdd.n1373 vdd.n1372 52.4337
R18433 vdd.n1187 vdd.n1152 52.4337
R18434 vdd.n1189 vdd.n1153 52.4337
R18435 vdd.n1193 vdd.n1154 52.4337
R18436 vdd.n1195 vdd.n1155 52.4337
R18437 vdd.n1199 vdd.n1156 52.4337
R18438 vdd.n1201 vdd.n1157 52.4337
R18439 vdd.n1205 vdd.n1158 52.4337
R18440 vdd.n1207 vdd.n1159 52.4337
R18441 vdd.n1339 vdd.n1160 52.4337
R18442 vdd.n1211 vdd.n1161 52.4337
R18443 vdd.n1215 vdd.n1162 52.4337
R18444 vdd.n1217 vdd.n1163 52.4337
R18445 vdd.n1221 vdd.n1164 52.4337
R18446 vdd.n1223 vdd.n1165 52.4337
R18447 vdd.n1227 vdd.n1166 52.4337
R18448 vdd.n1229 vdd.n1167 52.4337
R18449 vdd.n1233 vdd.n1168 52.4337
R18450 vdd.n1235 vdd.n1169 52.4337
R18451 vdd.n1239 vdd.n1170 52.4337
R18452 vdd.n1303 vdd.n1171 52.4337
R18453 vdd.n1244 vdd.n1172 52.4337
R18454 vdd.n1246 vdd.n1173 52.4337
R18455 vdd.n1250 vdd.n1174 52.4337
R18456 vdd.n1252 vdd.n1175 52.4337
R18457 vdd.n1256 vdd.n1176 52.4337
R18458 vdd.n1258 vdd.n1177 52.4337
R18459 vdd.n1262 vdd.n1178 52.4337
R18460 vdd.n1264 vdd.n1179 52.4337
R18461 vdd.n1268 vdd.n1180 52.4337
R18462 vdd.n1270 vdd.n1181 52.4337
R18463 vdd.n1373 vdd.n1183 52.4337
R18464 vdd.n1188 vdd.n1152 52.4337
R18465 vdd.n1192 vdd.n1153 52.4337
R18466 vdd.n1194 vdd.n1154 52.4337
R18467 vdd.n1198 vdd.n1155 52.4337
R18468 vdd.n1200 vdd.n1156 52.4337
R18469 vdd.n1204 vdd.n1157 52.4337
R18470 vdd.n1206 vdd.n1158 52.4337
R18471 vdd.n1338 vdd.n1159 52.4337
R18472 vdd.n1210 vdd.n1160 52.4337
R18473 vdd.n1214 vdd.n1161 52.4337
R18474 vdd.n1216 vdd.n1162 52.4337
R18475 vdd.n1220 vdd.n1163 52.4337
R18476 vdd.n1222 vdd.n1164 52.4337
R18477 vdd.n1226 vdd.n1165 52.4337
R18478 vdd.n1228 vdd.n1166 52.4337
R18479 vdd.n1232 vdd.n1167 52.4337
R18480 vdd.n1234 vdd.n1168 52.4337
R18481 vdd.n1238 vdd.n1169 52.4337
R18482 vdd.n1240 vdd.n1170 52.4337
R18483 vdd.n1243 vdd.n1171 52.4337
R18484 vdd.n1245 vdd.n1172 52.4337
R18485 vdd.n1249 vdd.n1173 52.4337
R18486 vdd.n1251 vdd.n1174 52.4337
R18487 vdd.n1255 vdd.n1175 52.4337
R18488 vdd.n1257 vdd.n1176 52.4337
R18489 vdd.n1261 vdd.n1177 52.4337
R18490 vdd.n1263 vdd.n1178 52.4337
R18491 vdd.n1267 vdd.n1179 52.4337
R18492 vdd.n1269 vdd.n1180 52.4337
R18493 vdd.n1181 vdd.n1151 52.4337
R18494 vdd.n1041 vdd.n1040 52.4337
R18495 vdd.n1918 vdd.n1917 52.4337
R18496 vdd.n1923 vdd.n1922 52.4337
R18497 vdd.n1928 vdd.n1927 52.4337
R18498 vdd.n1915 vdd.n1908 52.4337
R18499 vdd.n1935 vdd.n1934 52.4337
R18500 vdd.n1907 vdd.n1901 52.4337
R18501 vdd.n1942 vdd.n1941 52.4337
R18502 vdd.n1900 vdd.n1895 52.4337
R18503 vdd.n1949 vdd.n1948 52.4337
R18504 vdd.n1894 vdd.n1893 52.4337
R18505 vdd.n1889 vdd.n1882 52.4337
R18506 vdd.n1960 vdd.n1959 52.4337
R18507 vdd.n1881 vdd.n1875 52.4337
R18508 vdd.n1967 vdd.n1966 52.4337
R18509 vdd.n1874 vdd.n1868 52.4337
R18510 vdd.n1974 vdd.n1973 52.4337
R18511 vdd.n1867 vdd.n1861 52.4337
R18512 vdd.n1981 vdd.n1980 52.4337
R18513 vdd.n1860 vdd.n1855 52.4337
R18514 vdd.n1988 vdd.n1987 52.4337
R18515 vdd.n1854 vdd.n1853 52.4337
R18516 vdd.n1849 vdd.n1842 52.4337
R18517 vdd.n1999 vdd.n1998 52.4337
R18518 vdd.n1841 vdd.n1835 52.4337
R18519 vdd.n2006 vdd.n2005 52.4337
R18520 vdd.n1834 vdd.n1828 52.4337
R18521 vdd.n2013 vdd.n2012 52.4337
R18522 vdd.n2016 vdd.n2015 52.4337
R18523 vdd.n1825 vdd.n1820 52.4337
R18524 vdd.n2238 vdd.n2237 52.4337
R18525 vdd.n1819 vdd.n1047 52.4337
R18526 vdd.n3138 vdd.n3137 52.4337
R18527 vdd.n3132 vdd.n663 52.4337
R18528 vdd.n3128 vdd.n666 52.4337
R18529 vdd.n3126 vdd.n3125 52.4337
R18530 vdd.n3121 vdd.n3120 52.4337
R18531 vdd.n3118 vdd.n3117 52.4337
R18532 vdd.n3113 vdd.n3112 52.4337
R18533 vdd.n3110 vdd.n3109 52.4337
R18534 vdd.n3105 vdd.n3104 52.4337
R18535 vdd.n3102 vdd.n3101 52.4337
R18536 vdd.n3097 vdd.n3096 52.4337
R18537 vdd.n3094 vdd.n3093 52.4337
R18538 vdd.n3089 vdd.n3088 52.4337
R18539 vdd.n3086 vdd.n3085 52.4337
R18540 vdd.n3081 vdd.n3080 52.4337
R18541 vdd.n3078 vdd.n3077 52.4337
R18542 vdd.n3073 vdd.n3072 52.4337
R18543 vdd.n3070 vdd.n3069 52.4337
R18544 vdd.n3065 vdd.n3064 52.4337
R18545 vdd.n3062 vdd.n3061 52.4337
R18546 vdd.n728 vdd.n727 52.4337
R18547 vdd.n3053 vdd.n3052 52.4337
R18548 vdd.n3048 vdd.n729 52.4337
R18549 vdd.n3046 vdd.n3045 52.4337
R18550 vdd.n3041 vdd.n3040 52.4337
R18551 vdd.n3038 vdd.n3037 52.4337
R18552 vdd.n3033 vdd.n3032 52.4337
R18553 vdd.n3030 vdd.n3029 52.4337
R18554 vdd.n3025 vdd.n3024 52.4337
R18555 vdd.n3020 vdd.n750 52.4337
R18556 vdd.n3016 vdd.n752 52.4337
R18557 vdd.n3252 vdd.n404 52.4337
R18558 vdd.n595 vdd.n403 52.4337
R18559 vdd.n589 vdd.n402 52.4337
R18560 vdd.n585 vdd.n401 52.4337
R18561 vdd.n579 vdd.n400 52.4337
R18562 vdd.n575 vdd.n399 52.4337
R18563 vdd.n569 vdd.n398 52.4337
R18564 vdd.n565 vdd.n397 52.4337
R18565 vdd.n559 vdd.n396 52.4337
R18566 vdd.n555 vdd.n395 52.4337
R18567 vdd.n549 vdd.n394 52.4337
R18568 vdd.n545 vdd.n393 52.4337
R18569 vdd.n539 vdd.n392 52.4337
R18570 vdd.n535 vdd.n391 52.4337
R18571 vdd.n529 vdd.n390 52.4337
R18572 vdd.n525 vdd.n389 52.4337
R18573 vdd.n519 vdd.n388 52.4337
R18574 vdd.n515 vdd.n387 52.4337
R18575 vdd.n509 vdd.n386 52.4337
R18576 vdd.n505 vdd.n385 52.4337
R18577 vdd.n499 vdd.n384 52.4337
R18578 vdd.n495 vdd.n383 52.4337
R18579 vdd.n489 vdd.n382 52.4337
R18580 vdd.n485 vdd.n381 52.4337
R18581 vdd.n479 vdd.n380 52.4337
R18582 vdd.n475 vdd.n379 52.4337
R18583 vdd.n469 vdd.n378 52.4337
R18584 vdd.n465 vdd.n377 52.4337
R18585 vdd.n459 vdd.n376 52.4337
R18586 vdd.n455 vdd.n375 52.4337
R18587 vdd.n449 vdd.n374 52.4337
R18588 vdd.n445 vdd.n373 52.4337
R18589 vdd.t12 vdd.t151 51.4683
R18590 vdd.n266 vdd.n264 42.0461
R18591 vdd.n168 vdd.n166 42.0461
R18592 vdd.n71 vdd.n69 42.0461
R18593 vdd.n1690 vdd.n1688 42.0461
R18594 vdd.n1592 vdd.n1590 42.0461
R18595 vdd.n1495 vdd.n1493 42.0461
R18596 vdd.n320 vdd.n319 41.6884
R18597 vdd.n222 vdd.n221 41.6884
R18598 vdd.n125 vdd.n124 41.6884
R18599 vdd.n1744 vdd.n1743 41.6884
R18600 vdd.n1646 vdd.n1645 41.6884
R18601 vdd.n1549 vdd.n1548 41.6884
R18602 vdd.n1150 vdd.n1149 41.1157
R18603 vdd.n1306 vdd.n1305 41.1157
R18604 vdd.n1342 vdd.n1341 41.1157
R18605 vdd.n407 vdd.n406 41.1157
R18606 vdd.n547 vdd.n420 41.1157
R18607 vdd.n433 vdd.n432 41.1157
R18608 vdd.n2970 vdd.n2969 39.2114
R18609 vdd.n2967 vdd.n2966 39.2114
R18610 vdd.n2962 vdd.n784 39.2114
R18611 vdd.n2960 vdd.n2959 39.2114
R18612 vdd.n2955 vdd.n787 39.2114
R18613 vdd.n2953 vdd.n2952 39.2114
R18614 vdd.n2948 vdd.n790 39.2114
R18615 vdd.n2946 vdd.n2945 39.2114
R18616 vdd.n2940 vdd.n793 39.2114
R18617 vdd.n2938 vdd.n2937 39.2114
R18618 vdd.n2933 vdd.n796 39.2114
R18619 vdd.n2931 vdd.n2930 39.2114
R18620 vdd.n2926 vdd.n799 39.2114
R18621 vdd.n2924 vdd.n2923 39.2114
R18622 vdd.n2919 vdd.n802 39.2114
R18623 vdd.n2917 vdd.n2916 39.2114
R18624 vdd.n2912 vdd.n2911 39.2114
R18625 vdd.n2773 vdd.n884 39.2114
R18626 vdd.n2768 vdd.n2522 39.2114
R18627 vdd.n2765 vdd.n2523 39.2114
R18628 vdd.n2761 vdd.n2524 39.2114
R18629 vdd.n2757 vdd.n2525 39.2114
R18630 vdd.n2753 vdd.n2526 39.2114
R18631 vdd.n2749 vdd.n2527 39.2114
R18632 vdd.n2745 vdd.n2528 39.2114
R18633 vdd.n2741 vdd.n2529 39.2114
R18634 vdd.n2737 vdd.n2530 39.2114
R18635 vdd.n2733 vdd.n2531 39.2114
R18636 vdd.n2729 vdd.n2532 39.2114
R18637 vdd.n2725 vdd.n2533 39.2114
R18638 vdd.n2721 vdd.n2534 39.2114
R18639 vdd.n2717 vdd.n2535 39.2114
R18640 vdd.n2713 vdd.n2536 39.2114
R18641 vdd.n2708 vdd.n2537 39.2114
R18642 vdd.n2516 vdd.n924 39.2114
R18643 vdd.n2512 vdd.n923 39.2114
R18644 vdd.n2508 vdd.n922 39.2114
R18645 vdd.n2504 vdd.n921 39.2114
R18646 vdd.n2500 vdd.n920 39.2114
R18647 vdd.n2496 vdd.n919 39.2114
R18648 vdd.n2492 vdd.n918 39.2114
R18649 vdd.n2488 vdd.n917 39.2114
R18650 vdd.n2484 vdd.n916 39.2114
R18651 vdd.n2480 vdd.n915 39.2114
R18652 vdd.n2476 vdd.n914 39.2114
R18653 vdd.n2472 vdd.n913 39.2114
R18654 vdd.n2468 vdd.n912 39.2114
R18655 vdd.n2464 vdd.n911 39.2114
R18656 vdd.n2460 vdd.n910 39.2114
R18657 vdd.n2455 vdd.n909 39.2114
R18658 vdd.n2451 vdd.n908 39.2114
R18659 vdd.n2027 vdd.n1019 39.2114
R18660 vdd.n2033 vdd.n2032 39.2114
R18661 vdd.n2036 vdd.n2035 39.2114
R18662 vdd.n2041 vdd.n2040 39.2114
R18663 vdd.n2044 vdd.n2043 39.2114
R18664 vdd.n2049 vdd.n2048 39.2114
R18665 vdd.n2052 vdd.n2051 39.2114
R18666 vdd.n2057 vdd.n2056 39.2114
R18667 vdd.n2228 vdd.n2059 39.2114
R18668 vdd.n2227 vdd.n2226 39.2114
R18669 vdd.n2220 vdd.n2061 39.2114
R18670 vdd.n2219 vdd.n2218 39.2114
R18671 vdd.n2212 vdd.n2063 39.2114
R18672 vdd.n2211 vdd.n2210 39.2114
R18673 vdd.n2204 vdd.n2065 39.2114
R18674 vdd.n2203 vdd.n2202 39.2114
R18675 vdd.n2196 vdd.n2067 39.2114
R18676 vdd.n2889 vdd.n2888 39.2114
R18677 vdd.n2884 vdd.n2856 39.2114
R18678 vdd.n2882 vdd.n2881 39.2114
R18679 vdd.n2877 vdd.n2859 39.2114
R18680 vdd.n2875 vdd.n2874 39.2114
R18681 vdd.n2870 vdd.n2862 39.2114
R18682 vdd.n2868 vdd.n2867 39.2114
R18683 vdd.n2863 vdd.n755 39.2114
R18684 vdd.n3007 vdd.n3006 39.2114
R18685 vdd.n3004 vdd.n3003 39.2114
R18686 vdd.n2999 vdd.n760 39.2114
R18687 vdd.n2997 vdd.n2996 39.2114
R18688 vdd.n2992 vdd.n763 39.2114
R18689 vdd.n2990 vdd.n2989 39.2114
R18690 vdd.n2985 vdd.n766 39.2114
R18691 vdd.n2983 vdd.n2982 39.2114
R18692 vdd.n2978 vdd.n772 39.2114
R18693 vdd.n2775 vdd.n887 39.2114
R18694 vdd.n2538 vdd.n889 39.2114
R18695 vdd.n2564 vdd.n2539 39.2114
R18696 vdd.n2568 vdd.n2540 39.2114
R18697 vdd.n2572 vdd.n2541 39.2114
R18698 vdd.n2576 vdd.n2542 39.2114
R18699 vdd.n2580 vdd.n2543 39.2114
R18700 vdd.n2584 vdd.n2544 39.2114
R18701 vdd.n2588 vdd.n2545 39.2114
R18702 vdd.n2592 vdd.n2546 39.2114
R18703 vdd.n2596 vdd.n2547 39.2114
R18704 vdd.n2600 vdd.n2548 39.2114
R18705 vdd.n2604 vdd.n2549 39.2114
R18706 vdd.n2608 vdd.n2550 39.2114
R18707 vdd.n2612 vdd.n2551 39.2114
R18708 vdd.n2616 vdd.n2552 39.2114
R18709 vdd.n2620 vdd.n2553 39.2114
R18710 vdd.n2776 vdd.n2775 39.2114
R18711 vdd.n2563 vdd.n2538 39.2114
R18712 vdd.n2567 vdd.n2539 39.2114
R18713 vdd.n2571 vdd.n2540 39.2114
R18714 vdd.n2575 vdd.n2541 39.2114
R18715 vdd.n2579 vdd.n2542 39.2114
R18716 vdd.n2583 vdd.n2543 39.2114
R18717 vdd.n2587 vdd.n2544 39.2114
R18718 vdd.n2591 vdd.n2545 39.2114
R18719 vdd.n2595 vdd.n2546 39.2114
R18720 vdd.n2599 vdd.n2547 39.2114
R18721 vdd.n2603 vdd.n2548 39.2114
R18722 vdd.n2607 vdd.n2549 39.2114
R18723 vdd.n2611 vdd.n2550 39.2114
R18724 vdd.n2615 vdd.n2551 39.2114
R18725 vdd.n2619 vdd.n2552 39.2114
R18726 vdd.n2622 vdd.n2553 39.2114
R18727 vdd.n772 vdd.n767 39.2114
R18728 vdd.n2984 vdd.n2983 39.2114
R18729 vdd.n766 vdd.n764 39.2114
R18730 vdd.n2991 vdd.n2990 39.2114
R18731 vdd.n763 vdd.n761 39.2114
R18732 vdd.n2998 vdd.n2997 39.2114
R18733 vdd.n760 vdd.n758 39.2114
R18734 vdd.n3005 vdd.n3004 39.2114
R18735 vdd.n3008 vdd.n3007 39.2114
R18736 vdd.n2864 vdd.n2863 39.2114
R18737 vdd.n2869 vdd.n2868 39.2114
R18738 vdd.n2862 vdd.n2860 39.2114
R18739 vdd.n2876 vdd.n2875 39.2114
R18740 vdd.n2859 vdd.n2857 39.2114
R18741 vdd.n2883 vdd.n2882 39.2114
R18742 vdd.n2856 vdd.n2854 39.2114
R18743 vdd.n2890 vdd.n2889 39.2114
R18744 vdd.n2028 vdd.n2027 39.2114
R18745 vdd.n2034 vdd.n2033 39.2114
R18746 vdd.n2035 vdd.n2024 39.2114
R18747 vdd.n2042 vdd.n2041 39.2114
R18748 vdd.n2043 vdd.n2022 39.2114
R18749 vdd.n2050 vdd.n2049 39.2114
R18750 vdd.n2051 vdd.n2020 39.2114
R18751 vdd.n2058 vdd.n2057 39.2114
R18752 vdd.n2229 vdd.n2228 39.2114
R18753 vdd.n2226 vdd.n2225 39.2114
R18754 vdd.n2221 vdd.n2220 39.2114
R18755 vdd.n2218 vdd.n2217 39.2114
R18756 vdd.n2213 vdd.n2212 39.2114
R18757 vdd.n2210 vdd.n2209 39.2114
R18758 vdd.n2205 vdd.n2204 39.2114
R18759 vdd.n2202 vdd.n2201 39.2114
R18760 vdd.n2197 vdd.n2196 39.2114
R18761 vdd.n2454 vdd.n908 39.2114
R18762 vdd.n2459 vdd.n909 39.2114
R18763 vdd.n2463 vdd.n910 39.2114
R18764 vdd.n2467 vdd.n911 39.2114
R18765 vdd.n2471 vdd.n912 39.2114
R18766 vdd.n2475 vdd.n913 39.2114
R18767 vdd.n2479 vdd.n914 39.2114
R18768 vdd.n2483 vdd.n915 39.2114
R18769 vdd.n2487 vdd.n916 39.2114
R18770 vdd.n2491 vdd.n917 39.2114
R18771 vdd.n2495 vdd.n918 39.2114
R18772 vdd.n2499 vdd.n919 39.2114
R18773 vdd.n2503 vdd.n920 39.2114
R18774 vdd.n2507 vdd.n921 39.2114
R18775 vdd.n2511 vdd.n922 39.2114
R18776 vdd.n2515 vdd.n923 39.2114
R18777 vdd.n926 vdd.n924 39.2114
R18778 vdd.n2773 vdd.n2772 39.2114
R18779 vdd.n2766 vdd.n2522 39.2114
R18780 vdd.n2762 vdd.n2523 39.2114
R18781 vdd.n2758 vdd.n2524 39.2114
R18782 vdd.n2754 vdd.n2525 39.2114
R18783 vdd.n2750 vdd.n2526 39.2114
R18784 vdd.n2746 vdd.n2527 39.2114
R18785 vdd.n2742 vdd.n2528 39.2114
R18786 vdd.n2738 vdd.n2529 39.2114
R18787 vdd.n2734 vdd.n2530 39.2114
R18788 vdd.n2730 vdd.n2531 39.2114
R18789 vdd.n2726 vdd.n2532 39.2114
R18790 vdd.n2722 vdd.n2533 39.2114
R18791 vdd.n2718 vdd.n2534 39.2114
R18792 vdd.n2714 vdd.n2535 39.2114
R18793 vdd.n2709 vdd.n2536 39.2114
R18794 vdd.n2705 vdd.n2537 39.2114
R18795 vdd.n2911 vdd.n803 39.2114
R18796 vdd.n2918 vdd.n2917 39.2114
R18797 vdd.n802 vdd.n800 39.2114
R18798 vdd.n2925 vdd.n2924 39.2114
R18799 vdd.n799 vdd.n797 39.2114
R18800 vdd.n2932 vdd.n2931 39.2114
R18801 vdd.n796 vdd.n794 39.2114
R18802 vdd.n2939 vdd.n2938 39.2114
R18803 vdd.n793 vdd.n791 39.2114
R18804 vdd.n2947 vdd.n2946 39.2114
R18805 vdd.n790 vdd.n788 39.2114
R18806 vdd.n2954 vdd.n2953 39.2114
R18807 vdd.n787 vdd.n785 39.2114
R18808 vdd.n2961 vdd.n2960 39.2114
R18809 vdd.n784 vdd.n782 39.2114
R18810 vdd.n2968 vdd.n2967 39.2114
R18811 vdd.n2971 vdd.n2970 39.2114
R18812 vdd.n934 vdd.n890 39.2114
R18813 vdd.n2443 vdd.n891 39.2114
R18814 vdd.n2439 vdd.n892 39.2114
R18815 vdd.n2435 vdd.n893 39.2114
R18816 vdd.n2431 vdd.n894 39.2114
R18817 vdd.n2427 vdd.n895 39.2114
R18818 vdd.n2423 vdd.n896 39.2114
R18819 vdd.n2419 vdd.n897 39.2114
R18820 vdd.n2415 vdd.n898 39.2114
R18821 vdd.n2411 vdd.n899 39.2114
R18822 vdd.n2407 vdd.n900 39.2114
R18823 vdd.n2403 vdd.n901 39.2114
R18824 vdd.n2399 vdd.n902 39.2114
R18825 vdd.n2395 vdd.n903 39.2114
R18826 vdd.n2391 vdd.n904 39.2114
R18827 vdd.n2387 vdd.n905 39.2114
R18828 vdd.n2383 vdd.n906 39.2114
R18829 vdd.n2286 vdd.n1023 39.2114
R18830 vdd.n2285 vdd.n2284 39.2114
R18831 vdd.n2278 vdd.n1025 39.2114
R18832 vdd.n2277 vdd.n2276 39.2114
R18833 vdd.n2270 vdd.n1027 39.2114
R18834 vdd.n2269 vdd.n2268 39.2114
R18835 vdd.n2262 vdd.n1029 39.2114
R18836 vdd.n2261 vdd.n2260 39.2114
R18837 vdd.n1032 vdd.n1031 39.2114
R18838 vdd.n2102 vdd.n2101 39.2114
R18839 vdd.n2107 vdd.n2106 39.2114
R18840 vdd.n2110 vdd.n2109 39.2114
R18841 vdd.n2115 vdd.n2114 39.2114
R18842 vdd.n2118 vdd.n2117 39.2114
R18843 vdd.n2123 vdd.n2122 39.2114
R18844 vdd.n2126 vdd.n2125 39.2114
R18845 vdd.n2132 vdd.n2131 39.2114
R18846 vdd.n2380 vdd.n906 39.2114
R18847 vdd.n2384 vdd.n905 39.2114
R18848 vdd.n2388 vdd.n904 39.2114
R18849 vdd.n2392 vdd.n903 39.2114
R18850 vdd.n2396 vdd.n902 39.2114
R18851 vdd.n2400 vdd.n901 39.2114
R18852 vdd.n2404 vdd.n900 39.2114
R18853 vdd.n2408 vdd.n899 39.2114
R18854 vdd.n2412 vdd.n898 39.2114
R18855 vdd.n2416 vdd.n897 39.2114
R18856 vdd.n2420 vdd.n896 39.2114
R18857 vdd.n2424 vdd.n895 39.2114
R18858 vdd.n2428 vdd.n894 39.2114
R18859 vdd.n2432 vdd.n893 39.2114
R18860 vdd.n2436 vdd.n892 39.2114
R18861 vdd.n2440 vdd.n891 39.2114
R18862 vdd.n2444 vdd.n890 39.2114
R18863 vdd.n2287 vdd.n2286 39.2114
R18864 vdd.n2284 vdd.n2283 39.2114
R18865 vdd.n2279 vdd.n2278 39.2114
R18866 vdd.n2276 vdd.n2275 39.2114
R18867 vdd.n2271 vdd.n2270 39.2114
R18868 vdd.n2268 vdd.n2267 39.2114
R18869 vdd.n2263 vdd.n2262 39.2114
R18870 vdd.n2260 vdd.n2259 39.2114
R18871 vdd.n1033 vdd.n1032 39.2114
R18872 vdd.n2103 vdd.n2102 39.2114
R18873 vdd.n2108 vdd.n2107 39.2114
R18874 vdd.n2109 vdd.n2099 39.2114
R18875 vdd.n2116 vdd.n2115 39.2114
R18876 vdd.n2117 vdd.n2097 39.2114
R18877 vdd.n2124 vdd.n2123 39.2114
R18878 vdd.n2125 vdd.n2093 39.2114
R18879 vdd.n2133 vdd.n2132 39.2114
R18880 vdd.n2252 vdd.n2251 37.2369
R18881 vdd.n1955 vdd.n1888 37.2369
R18882 vdd.n1994 vdd.n1848 37.2369
R18883 vdd.n3059 vdd.n724 37.2369
R18884 vdd.n688 vdd.n687 37.2369
R18885 vdd.n3015 vdd.n3014 37.2369
R18886 vdd.n2294 vdd.n1018 31.6883
R18887 vdd.n2519 vdd.n927 31.6883
R18888 vdd.n2452 vdd.n930 31.6883
R18889 vdd.n2198 vdd.n2195 31.6883
R18890 vdd.n2706 vdd.n2704 31.6883
R18891 vdd.n2913 vdd.n2910 31.6883
R18892 vdd.n2783 vdd.n883 31.6883
R18893 vdd.n2974 vdd.n2973 31.6883
R18894 vdd.n2893 vdd.n2892 31.6883
R18895 vdd.n2979 vdd.n771 31.6883
R18896 vdd.n2625 vdd.n2624 31.6883
R18897 vdd.n2779 vdd.n2778 31.6883
R18898 vdd.n2290 vdd.n2289 31.6883
R18899 vdd.n2447 vdd.n2446 31.6883
R18900 vdd.n2379 vdd.n2378 31.6883
R18901 vdd.n2136 vdd.n2135 31.6883
R18902 vdd.n2129 vdd.n2095 30.449
R18903 vdd.n938 vdd.n937 30.449
R18904 vdd.n2070 vdd.n2069 30.449
R18905 vdd.n2457 vdd.n929 30.449
R18906 vdd.n2561 vdd.n2560 30.449
R18907 vdd.n806 vdd.n805 30.449
R18908 vdd.n2711 vdd.n2557 30.449
R18909 vdd.n770 vdd.n769 30.449
R18910 vdd.n1380 vdd.n1146 19.3944
R18911 vdd.n1380 vdd.n1136 19.3944
R18912 vdd.n1392 vdd.n1136 19.3944
R18913 vdd.n1392 vdd.n1134 19.3944
R18914 vdd.n1396 vdd.n1134 19.3944
R18915 vdd.n1396 vdd.n1124 19.3944
R18916 vdd.n1409 vdd.n1124 19.3944
R18917 vdd.n1409 vdd.n1122 19.3944
R18918 vdd.n1413 vdd.n1122 19.3944
R18919 vdd.n1413 vdd.n1114 19.3944
R18920 vdd.n1426 vdd.n1114 19.3944
R18921 vdd.n1426 vdd.n1112 19.3944
R18922 vdd.n1430 vdd.n1112 19.3944
R18923 vdd.n1430 vdd.n1101 19.3944
R18924 vdd.n1442 vdd.n1101 19.3944
R18925 vdd.n1442 vdd.n1099 19.3944
R18926 vdd.n1446 vdd.n1099 19.3944
R18927 vdd.n1446 vdd.n1090 19.3944
R18928 vdd.n1754 vdd.n1090 19.3944
R18929 vdd.n1754 vdd.n1088 19.3944
R18930 vdd.n1758 vdd.n1088 19.3944
R18931 vdd.n1758 vdd.n1079 19.3944
R18932 vdd.n1770 vdd.n1079 19.3944
R18933 vdd.n1770 vdd.n1077 19.3944
R18934 vdd.n1774 vdd.n1077 19.3944
R18935 vdd.n1774 vdd.n1067 19.3944
R18936 vdd.n1787 vdd.n1067 19.3944
R18937 vdd.n1787 vdd.n1065 19.3944
R18938 vdd.n1791 vdd.n1065 19.3944
R18939 vdd.n1791 vdd.n1057 19.3944
R18940 vdd.n1804 vdd.n1057 19.3944
R18941 vdd.n1804 vdd.n1054 19.3944
R18942 vdd.n1810 vdd.n1054 19.3944
R18943 vdd.n1810 vdd.n1055 19.3944
R18944 vdd.n1055 vdd.n1043 19.3944
R18945 vdd.n1299 vdd.n1241 19.3944
R18946 vdd.n1299 vdd.n1298 19.3944
R18947 vdd.n1298 vdd.n1297 19.3944
R18948 vdd.n1297 vdd.n1247 19.3944
R18949 vdd.n1293 vdd.n1247 19.3944
R18950 vdd.n1293 vdd.n1292 19.3944
R18951 vdd.n1292 vdd.n1291 19.3944
R18952 vdd.n1291 vdd.n1253 19.3944
R18953 vdd.n1287 vdd.n1253 19.3944
R18954 vdd.n1287 vdd.n1286 19.3944
R18955 vdd.n1286 vdd.n1285 19.3944
R18956 vdd.n1285 vdd.n1259 19.3944
R18957 vdd.n1281 vdd.n1259 19.3944
R18958 vdd.n1281 vdd.n1280 19.3944
R18959 vdd.n1280 vdd.n1279 19.3944
R18960 vdd.n1279 vdd.n1265 19.3944
R18961 vdd.n1275 vdd.n1265 19.3944
R18962 vdd.n1275 vdd.n1274 19.3944
R18963 vdd.n1274 vdd.n1273 19.3944
R18964 vdd.n1273 vdd.n1271 19.3944
R18965 vdd.n1337 vdd.n1336 19.3944
R18966 vdd.n1336 vdd.n1212 19.3944
R18967 vdd.n1332 vdd.n1212 19.3944
R18968 vdd.n1332 vdd.n1331 19.3944
R18969 vdd.n1331 vdd.n1330 19.3944
R18970 vdd.n1330 vdd.n1218 19.3944
R18971 vdd.n1326 vdd.n1218 19.3944
R18972 vdd.n1326 vdd.n1325 19.3944
R18973 vdd.n1325 vdd.n1324 19.3944
R18974 vdd.n1324 vdd.n1224 19.3944
R18975 vdd.n1320 vdd.n1224 19.3944
R18976 vdd.n1320 vdd.n1319 19.3944
R18977 vdd.n1319 vdd.n1318 19.3944
R18978 vdd.n1318 vdd.n1230 19.3944
R18979 vdd.n1314 vdd.n1230 19.3944
R18980 vdd.n1314 vdd.n1313 19.3944
R18981 vdd.n1313 vdd.n1312 19.3944
R18982 vdd.n1312 vdd.n1236 19.3944
R18983 vdd.n1308 vdd.n1236 19.3944
R18984 vdd.n1308 vdd.n1307 19.3944
R18985 vdd.n1371 vdd.n1370 19.3944
R18986 vdd.n1370 vdd.n1185 19.3944
R18987 vdd.n1366 vdd.n1185 19.3944
R18988 vdd.n1366 vdd.n1365 19.3944
R18989 vdd.n1365 vdd.n1364 19.3944
R18990 vdd.n1364 vdd.n1190 19.3944
R18991 vdd.n1360 vdd.n1190 19.3944
R18992 vdd.n1360 vdd.n1359 19.3944
R18993 vdd.n1359 vdd.n1358 19.3944
R18994 vdd.n1358 vdd.n1196 19.3944
R18995 vdd.n1354 vdd.n1196 19.3944
R18996 vdd.n1354 vdd.n1353 19.3944
R18997 vdd.n1353 vdd.n1352 19.3944
R18998 vdd.n1352 vdd.n1202 19.3944
R18999 vdd.n1348 vdd.n1202 19.3944
R19000 vdd.n1348 vdd.n1347 19.3944
R19001 vdd.n1347 vdd.n1346 19.3944
R19002 vdd.n1346 vdd.n1208 19.3944
R19003 vdd.n1951 vdd.n1886 19.3944
R19004 vdd.n1951 vdd.n1892 19.3944
R19005 vdd.n1946 vdd.n1892 19.3944
R19006 vdd.n1946 vdd.n1945 19.3944
R19007 vdd.n1945 vdd.n1944 19.3944
R19008 vdd.n1944 vdd.n1899 19.3944
R19009 vdd.n1939 vdd.n1899 19.3944
R19010 vdd.n1939 vdd.n1938 19.3944
R19011 vdd.n1938 vdd.n1937 19.3944
R19012 vdd.n1937 vdd.n1906 19.3944
R19013 vdd.n1932 vdd.n1906 19.3944
R19014 vdd.n1932 vdd.n1931 19.3944
R19015 vdd.n1931 vdd.n1930 19.3944
R19016 vdd.n1930 vdd.n1914 19.3944
R19017 vdd.n1925 vdd.n1914 19.3944
R19018 vdd.n1925 vdd.n1924 19.3944
R19019 vdd.n1920 vdd.n1919 19.3944
R19020 vdd.n2253 vdd.n1039 19.3944
R19021 vdd.n1990 vdd.n1846 19.3944
R19022 vdd.n1990 vdd.n1852 19.3944
R19023 vdd.n1985 vdd.n1852 19.3944
R19024 vdd.n1985 vdd.n1984 19.3944
R19025 vdd.n1984 vdd.n1983 19.3944
R19026 vdd.n1983 vdd.n1859 19.3944
R19027 vdd.n1978 vdd.n1859 19.3944
R19028 vdd.n1978 vdd.n1977 19.3944
R19029 vdd.n1977 vdd.n1976 19.3944
R19030 vdd.n1976 vdd.n1866 19.3944
R19031 vdd.n1971 vdd.n1866 19.3944
R19032 vdd.n1971 vdd.n1970 19.3944
R19033 vdd.n1970 vdd.n1969 19.3944
R19034 vdd.n1969 vdd.n1873 19.3944
R19035 vdd.n1964 vdd.n1873 19.3944
R19036 vdd.n1964 vdd.n1963 19.3944
R19037 vdd.n1963 vdd.n1962 19.3944
R19038 vdd.n1962 vdd.n1880 19.3944
R19039 vdd.n1957 vdd.n1880 19.3944
R19040 vdd.n1957 vdd.n1956 19.3944
R19041 vdd.n2241 vdd.n2240 19.3944
R19042 vdd.n2240 vdd.n1818 19.3944
R19043 vdd.n2235 vdd.n2234 19.3944
R19044 vdd.n2017 vdd.n1822 19.3944
R19045 vdd.n2017 vdd.n1824 19.3944
R19046 vdd.n1827 vdd.n1824 19.3944
R19047 vdd.n2010 vdd.n1827 19.3944
R19048 vdd.n2010 vdd.n2009 19.3944
R19049 vdd.n2009 vdd.n2008 19.3944
R19050 vdd.n2008 vdd.n1833 19.3944
R19051 vdd.n2003 vdd.n1833 19.3944
R19052 vdd.n2003 vdd.n2002 19.3944
R19053 vdd.n2002 vdd.n2001 19.3944
R19054 vdd.n2001 vdd.n1840 19.3944
R19055 vdd.n1996 vdd.n1840 19.3944
R19056 vdd.n1996 vdd.n1995 19.3944
R19057 vdd.n1384 vdd.n1142 19.3944
R19058 vdd.n1384 vdd.n1140 19.3944
R19059 vdd.n1388 vdd.n1140 19.3944
R19060 vdd.n1388 vdd.n1130 19.3944
R19061 vdd.n1401 vdd.n1130 19.3944
R19062 vdd.n1401 vdd.n1128 19.3944
R19063 vdd.n1405 vdd.n1128 19.3944
R19064 vdd.n1405 vdd.n1119 19.3944
R19065 vdd.n1418 vdd.n1119 19.3944
R19066 vdd.n1418 vdd.n1117 19.3944
R19067 vdd.n1422 vdd.n1117 19.3944
R19068 vdd.n1422 vdd.n1108 19.3944
R19069 vdd.n1434 vdd.n1108 19.3944
R19070 vdd.n1434 vdd.n1106 19.3944
R19071 vdd.n1438 vdd.n1106 19.3944
R19072 vdd.n1438 vdd.n1096 19.3944
R19073 vdd.n1451 vdd.n1096 19.3944
R19074 vdd.n1451 vdd.n1094 19.3944
R19075 vdd.n1750 vdd.n1094 19.3944
R19076 vdd.n1750 vdd.n1085 19.3944
R19077 vdd.n1762 vdd.n1085 19.3944
R19078 vdd.n1762 vdd.n1083 19.3944
R19079 vdd.n1766 vdd.n1083 19.3944
R19080 vdd.n1766 vdd.n1073 19.3944
R19081 vdd.n1779 vdd.n1073 19.3944
R19082 vdd.n1779 vdd.n1071 19.3944
R19083 vdd.n1783 vdd.n1071 19.3944
R19084 vdd.n1783 vdd.n1062 19.3944
R19085 vdd.n1796 vdd.n1062 19.3944
R19086 vdd.n1796 vdd.n1060 19.3944
R19087 vdd.n1800 vdd.n1060 19.3944
R19088 vdd.n1800 vdd.n1050 19.3944
R19089 vdd.n1814 vdd.n1050 19.3944
R19090 vdd.n1814 vdd.n1048 19.3944
R19091 vdd.n2244 vdd.n1048 19.3944
R19092 vdd.n3147 vdd.n655 19.3944
R19093 vdd.n3151 vdd.n655 19.3944
R19094 vdd.n3151 vdd.n646 19.3944
R19095 vdd.n3163 vdd.n646 19.3944
R19096 vdd.n3163 vdd.n644 19.3944
R19097 vdd.n3167 vdd.n644 19.3944
R19098 vdd.n3167 vdd.n633 19.3944
R19099 vdd.n3179 vdd.n633 19.3944
R19100 vdd.n3179 vdd.n631 19.3944
R19101 vdd.n3183 vdd.n631 19.3944
R19102 vdd.n3183 vdd.n622 19.3944
R19103 vdd.n3196 vdd.n622 19.3944
R19104 vdd.n3196 vdd.n620 19.3944
R19105 vdd.n3203 vdd.n620 19.3944
R19106 vdd.n3203 vdd.n3202 19.3944
R19107 vdd.n3202 vdd.n610 19.3944
R19108 vdd.n3216 vdd.n610 19.3944
R19109 vdd.n3217 vdd.n3216 19.3944
R19110 vdd.n3218 vdd.n3217 19.3944
R19111 vdd.n3218 vdd.n608 19.3944
R19112 vdd.n3223 vdd.n608 19.3944
R19113 vdd.n3224 vdd.n3223 19.3944
R19114 vdd.n3225 vdd.n3224 19.3944
R19115 vdd.n3225 vdd.n606 19.3944
R19116 vdd.n3230 vdd.n606 19.3944
R19117 vdd.n3231 vdd.n3230 19.3944
R19118 vdd.n3232 vdd.n3231 19.3944
R19119 vdd.n3232 vdd.n604 19.3944
R19120 vdd.n3238 vdd.n604 19.3944
R19121 vdd.n3239 vdd.n3238 19.3944
R19122 vdd.n3240 vdd.n3239 19.3944
R19123 vdd.n3240 vdd.n602 19.3944
R19124 vdd.n3245 vdd.n602 19.3944
R19125 vdd.n3246 vdd.n3245 19.3944
R19126 vdd.n3247 vdd.n3246 19.3944
R19127 vdd.n550 vdd.n417 19.3944
R19128 vdd.n556 vdd.n417 19.3944
R19129 vdd.n557 vdd.n556 19.3944
R19130 vdd.n560 vdd.n557 19.3944
R19131 vdd.n560 vdd.n415 19.3944
R19132 vdd.n566 vdd.n415 19.3944
R19133 vdd.n567 vdd.n566 19.3944
R19134 vdd.n570 vdd.n567 19.3944
R19135 vdd.n570 vdd.n413 19.3944
R19136 vdd.n576 vdd.n413 19.3944
R19137 vdd.n577 vdd.n576 19.3944
R19138 vdd.n580 vdd.n577 19.3944
R19139 vdd.n580 vdd.n411 19.3944
R19140 vdd.n586 vdd.n411 19.3944
R19141 vdd.n587 vdd.n586 19.3944
R19142 vdd.n590 vdd.n587 19.3944
R19143 vdd.n590 vdd.n409 19.3944
R19144 vdd.n596 vdd.n409 19.3944
R19145 vdd.n598 vdd.n596 19.3944
R19146 vdd.n599 vdd.n598 19.3944
R19147 vdd.n497 vdd.n496 19.3944
R19148 vdd.n500 vdd.n497 19.3944
R19149 vdd.n500 vdd.n429 19.3944
R19150 vdd.n506 vdd.n429 19.3944
R19151 vdd.n507 vdd.n506 19.3944
R19152 vdd.n510 vdd.n507 19.3944
R19153 vdd.n510 vdd.n427 19.3944
R19154 vdd.n516 vdd.n427 19.3944
R19155 vdd.n517 vdd.n516 19.3944
R19156 vdd.n520 vdd.n517 19.3944
R19157 vdd.n520 vdd.n425 19.3944
R19158 vdd.n526 vdd.n425 19.3944
R19159 vdd.n527 vdd.n526 19.3944
R19160 vdd.n530 vdd.n527 19.3944
R19161 vdd.n530 vdd.n423 19.3944
R19162 vdd.n536 vdd.n423 19.3944
R19163 vdd.n537 vdd.n536 19.3944
R19164 vdd.n540 vdd.n537 19.3944
R19165 vdd.n540 vdd.n421 19.3944
R19166 vdd.n546 vdd.n421 19.3944
R19167 vdd.n447 vdd.n446 19.3944
R19168 vdd.n450 vdd.n447 19.3944
R19169 vdd.n450 vdd.n441 19.3944
R19170 vdd.n456 vdd.n441 19.3944
R19171 vdd.n457 vdd.n456 19.3944
R19172 vdd.n460 vdd.n457 19.3944
R19173 vdd.n460 vdd.n439 19.3944
R19174 vdd.n466 vdd.n439 19.3944
R19175 vdd.n467 vdd.n466 19.3944
R19176 vdd.n470 vdd.n467 19.3944
R19177 vdd.n470 vdd.n437 19.3944
R19178 vdd.n476 vdd.n437 19.3944
R19179 vdd.n477 vdd.n476 19.3944
R19180 vdd.n480 vdd.n477 19.3944
R19181 vdd.n480 vdd.n435 19.3944
R19182 vdd.n486 vdd.n435 19.3944
R19183 vdd.n487 vdd.n486 19.3944
R19184 vdd.n490 vdd.n487 19.3944
R19185 vdd.n3143 vdd.n652 19.3944
R19186 vdd.n3155 vdd.n652 19.3944
R19187 vdd.n3155 vdd.n650 19.3944
R19188 vdd.n3159 vdd.n650 19.3944
R19189 vdd.n3159 vdd.n640 19.3944
R19190 vdd.n3171 vdd.n640 19.3944
R19191 vdd.n3171 vdd.n638 19.3944
R19192 vdd.n3175 vdd.n638 19.3944
R19193 vdd.n3175 vdd.n628 19.3944
R19194 vdd.n3188 vdd.n628 19.3944
R19195 vdd.n3188 vdd.n626 19.3944
R19196 vdd.n3192 vdd.n626 19.3944
R19197 vdd.n3192 vdd.n617 19.3944
R19198 vdd.n3207 vdd.n617 19.3944
R19199 vdd.n3207 vdd.n615 19.3944
R19200 vdd.n3211 vdd.n615 19.3944
R19201 vdd.n3211 vdd.n324 19.3944
R19202 vdd.n3289 vdd.n324 19.3944
R19203 vdd.n3289 vdd.n325 19.3944
R19204 vdd.n3283 vdd.n325 19.3944
R19205 vdd.n3283 vdd.n3282 19.3944
R19206 vdd.n3282 vdd.n3281 19.3944
R19207 vdd.n3281 vdd.n337 19.3944
R19208 vdd.n3275 vdd.n337 19.3944
R19209 vdd.n3275 vdd.n3274 19.3944
R19210 vdd.n3274 vdd.n3273 19.3944
R19211 vdd.n3273 vdd.n347 19.3944
R19212 vdd.n3267 vdd.n347 19.3944
R19213 vdd.n3267 vdd.n3266 19.3944
R19214 vdd.n3266 vdd.n3265 19.3944
R19215 vdd.n3265 vdd.n358 19.3944
R19216 vdd.n3259 vdd.n358 19.3944
R19217 vdd.n3259 vdd.n3258 19.3944
R19218 vdd.n3258 vdd.n3257 19.3944
R19219 vdd.n3257 vdd.n369 19.3944
R19220 vdd.n3100 vdd.n3099 19.3944
R19221 vdd.n3099 vdd.n3098 19.3944
R19222 vdd.n3098 vdd.n694 19.3944
R19223 vdd.n3092 vdd.n694 19.3944
R19224 vdd.n3092 vdd.n3091 19.3944
R19225 vdd.n3091 vdd.n3090 19.3944
R19226 vdd.n3090 vdd.n700 19.3944
R19227 vdd.n3084 vdd.n700 19.3944
R19228 vdd.n3084 vdd.n3083 19.3944
R19229 vdd.n3083 vdd.n3082 19.3944
R19230 vdd.n3082 vdd.n706 19.3944
R19231 vdd.n3076 vdd.n706 19.3944
R19232 vdd.n3076 vdd.n3075 19.3944
R19233 vdd.n3075 vdd.n3074 19.3944
R19234 vdd.n3074 vdd.n712 19.3944
R19235 vdd.n3068 vdd.n712 19.3944
R19236 vdd.n3068 vdd.n3067 19.3944
R19237 vdd.n3067 vdd.n3066 19.3944
R19238 vdd.n3066 vdd.n718 19.3944
R19239 vdd.n3060 vdd.n718 19.3944
R19240 vdd.n3140 vdd.n3139 19.3944
R19241 vdd.n3139 vdd.n662 19.3944
R19242 vdd.n3134 vdd.n3133 19.3944
R19243 vdd.n3130 vdd.n3129 19.3944
R19244 vdd.n3129 vdd.n668 19.3944
R19245 vdd.n3124 vdd.n668 19.3944
R19246 vdd.n3124 vdd.n3123 19.3944
R19247 vdd.n3123 vdd.n3122 19.3944
R19248 vdd.n3122 vdd.n674 19.3944
R19249 vdd.n3116 vdd.n674 19.3944
R19250 vdd.n3116 vdd.n3115 19.3944
R19251 vdd.n3115 vdd.n3114 19.3944
R19252 vdd.n3114 vdd.n680 19.3944
R19253 vdd.n3108 vdd.n680 19.3944
R19254 vdd.n3108 vdd.n3107 19.3944
R19255 vdd.n3107 vdd.n3106 19.3944
R19256 vdd.n3055 vdd.n722 19.3944
R19257 vdd.n3055 vdd.n726 19.3944
R19258 vdd.n3050 vdd.n726 19.3944
R19259 vdd.n3050 vdd.n3049 19.3944
R19260 vdd.n3049 vdd.n732 19.3944
R19261 vdd.n3044 vdd.n732 19.3944
R19262 vdd.n3044 vdd.n3043 19.3944
R19263 vdd.n3043 vdd.n3042 19.3944
R19264 vdd.n3042 vdd.n738 19.3944
R19265 vdd.n3036 vdd.n738 19.3944
R19266 vdd.n3036 vdd.n3035 19.3944
R19267 vdd.n3035 vdd.n3034 19.3944
R19268 vdd.n3034 vdd.n744 19.3944
R19269 vdd.n3028 vdd.n744 19.3944
R19270 vdd.n3028 vdd.n3027 19.3944
R19271 vdd.n3027 vdd.n3026 19.3944
R19272 vdd.n3022 vdd.n3021 19.3944
R19273 vdd.n3018 vdd.n3017 19.3944
R19274 vdd.n1306 vdd.n1241 19.0066
R19275 vdd.n1955 vdd.n1886 19.0066
R19276 vdd.n550 vdd.n547 19.0066
R19277 vdd.n3059 vdd.n722 19.0066
R19278 vdd.n1374 vdd.n1144 18.5924
R19279 vdd.n2246 vdd.n1045 18.5924
R19280 vdd.n3145 vdd.n658 18.5924
R19281 vdd.n3254 vdd.n3253 18.5924
R19282 vdd.n2095 vdd.n2094 16.0975
R19283 vdd.n937 vdd.n936 16.0975
R19284 vdd.n1149 vdd.n1148 16.0975
R19285 vdd.n1305 vdd.n1304 16.0975
R19286 vdd.n1341 vdd.n1340 16.0975
R19287 vdd.n2251 vdd.n2250 16.0975
R19288 vdd.n1888 vdd.n1887 16.0975
R19289 vdd.n1848 vdd.n1847 16.0975
R19290 vdd.n2069 vdd.n2068 16.0975
R19291 vdd.n929 vdd.n928 16.0975
R19292 vdd.n2560 vdd.n2559 16.0975
R19293 vdd.n406 vdd.n405 16.0975
R19294 vdd.n420 vdd.n419 16.0975
R19295 vdd.n432 vdd.n431 16.0975
R19296 vdd.n724 vdd.n723 16.0975
R19297 vdd.n687 vdd.n686 16.0975
R19298 vdd.n805 vdd.n804 16.0975
R19299 vdd.n2557 vdd.n2556 16.0975
R19300 vdd.n3014 vdd.n3013 16.0975
R19301 vdd.n769 vdd.n768 16.0975
R19302 vdd.t151 vdd.n2521 15.4182
R19303 vdd.n2774 vdd.t12 15.4182
R19304 vdd.n28 vdd.n27 14.6905
R19305 vdd.n2292 vdd.n1020 14.5112
R19306 vdd.n2976 vdd.n756 14.5112
R19307 vdd.n316 vdd.n281 13.1884
R19308 vdd.n261 vdd.n226 13.1884
R19309 vdd.n218 vdd.n183 13.1884
R19310 vdd.n163 vdd.n128 13.1884
R19311 vdd.n121 vdd.n86 13.1884
R19312 vdd.n66 vdd.n31 13.1884
R19313 vdd.n1685 vdd.n1650 13.1884
R19314 vdd.n1740 vdd.n1705 13.1884
R19315 vdd.n1587 vdd.n1552 13.1884
R19316 vdd.n1642 vdd.n1607 13.1884
R19317 vdd.n1490 vdd.n1455 13.1884
R19318 vdd.n1545 vdd.n1510 13.1884
R19319 vdd.n1342 vdd.n1337 12.9944
R19320 vdd.n1342 vdd.n1208 12.9944
R19321 vdd.n1994 vdd.n1846 12.9944
R19322 vdd.n1995 vdd.n1994 12.9944
R19323 vdd.n496 vdd.n433 12.9944
R19324 vdd.n490 vdd.n433 12.9944
R19325 vdd.n3100 vdd.n688 12.9944
R19326 vdd.n3106 vdd.n688 12.9944
R19327 vdd.n317 vdd.n279 12.8005
R19328 vdd.n312 vdd.n283 12.8005
R19329 vdd.n262 vdd.n224 12.8005
R19330 vdd.n257 vdd.n228 12.8005
R19331 vdd.n219 vdd.n181 12.8005
R19332 vdd.n214 vdd.n185 12.8005
R19333 vdd.n164 vdd.n126 12.8005
R19334 vdd.n159 vdd.n130 12.8005
R19335 vdd.n122 vdd.n84 12.8005
R19336 vdd.n117 vdd.n88 12.8005
R19337 vdd.n67 vdd.n29 12.8005
R19338 vdd.n62 vdd.n33 12.8005
R19339 vdd.n1686 vdd.n1648 12.8005
R19340 vdd.n1681 vdd.n1652 12.8005
R19341 vdd.n1741 vdd.n1703 12.8005
R19342 vdd.n1736 vdd.n1707 12.8005
R19343 vdd.n1588 vdd.n1550 12.8005
R19344 vdd.n1583 vdd.n1554 12.8005
R19345 vdd.n1643 vdd.n1605 12.8005
R19346 vdd.n1638 vdd.n1609 12.8005
R19347 vdd.n1491 vdd.n1453 12.8005
R19348 vdd.n1486 vdd.n1457 12.8005
R19349 vdd.n1546 vdd.n1508 12.8005
R19350 vdd.n1541 vdd.n1512 12.8005
R19351 vdd.n311 vdd.n284 12.0247
R19352 vdd.n256 vdd.n229 12.0247
R19353 vdd.n213 vdd.n186 12.0247
R19354 vdd.n158 vdd.n131 12.0247
R19355 vdd.n116 vdd.n89 12.0247
R19356 vdd.n61 vdd.n34 12.0247
R19357 vdd.n1680 vdd.n1653 12.0247
R19358 vdd.n1735 vdd.n1708 12.0247
R19359 vdd.n1582 vdd.n1555 12.0247
R19360 vdd.n1637 vdd.n1610 12.0247
R19361 vdd.n1485 vdd.n1458 12.0247
R19362 vdd.n1540 vdd.n1513 12.0247
R19363 vdd.n1382 vdd.n1144 11.337
R19364 vdd.n1390 vdd.n1138 11.337
R19365 vdd.n1390 vdd.n1132 11.337
R19366 vdd.n1399 vdd.n1132 11.337
R19367 vdd.n1407 vdd.n1126 11.337
R19368 vdd.n1416 vdd.n1415 11.337
R19369 vdd.n1432 vdd.n1110 11.337
R19370 vdd.n1440 vdd.n1103 11.337
R19371 vdd.n1449 vdd.n1448 11.337
R19372 vdd.n1752 vdd.n1092 11.337
R19373 vdd.n1768 vdd.n1081 11.337
R19374 vdd.n1777 vdd.n1075 11.337
R19375 vdd.n1785 vdd.n1069 11.337
R19376 vdd.n1794 vdd.n1793 11.337
R19377 vdd.n1802 vdd.n1052 11.337
R19378 vdd.n1812 vdd.n1052 11.337
R19379 vdd.n2246 vdd.n1044 11.337
R19380 vdd.n3145 vdd.n659 11.337
R19381 vdd.n3153 vdd.n648 11.337
R19382 vdd.n3161 vdd.n648 11.337
R19383 vdd.n3169 vdd.n642 11.337
R19384 vdd.n3177 vdd.n635 11.337
R19385 vdd.n3186 vdd.n3185 11.337
R19386 vdd.n3194 vdd.n624 11.337
R19387 vdd.n3213 vdd.n613 11.337
R19388 vdd.n3287 vdd.n328 11.337
R19389 vdd.n3285 vdd.n332 11.337
R19390 vdd.n3279 vdd.n3278 11.337
R19391 vdd.n3271 vdd.n349 11.337
R19392 vdd.n3270 vdd.n3269 11.337
R19393 vdd.n3263 vdd.n3262 11.337
R19394 vdd.n3262 vdd.n3261 11.337
R19395 vdd.n3261 vdd.n363 11.337
R19396 vdd.n3255 vdd.n3254 11.337
R19397 vdd.n308 vdd.n307 11.249
R19398 vdd.n253 vdd.n252 11.249
R19399 vdd.n210 vdd.n209 11.249
R19400 vdd.n155 vdd.n154 11.249
R19401 vdd.n113 vdd.n112 11.249
R19402 vdd.n58 vdd.n57 11.249
R19403 vdd.n1677 vdd.n1676 11.249
R19404 vdd.n1732 vdd.n1731 11.249
R19405 vdd.n1579 vdd.n1578 11.249
R19406 vdd.n1634 vdd.n1633 11.249
R19407 vdd.n1482 vdd.n1481 11.249
R19408 vdd.n1537 vdd.n1536 11.249
R19409 vdd.n2449 vdd.t6 11.1103
R19410 vdd.n2781 vdd.t159 11.1103
R19411 vdd.n1802 vdd.t19 10.7702
R19412 vdd.n3161 vdd.t21 10.7702
R19413 vdd.n293 vdd.n292 10.7238
R19414 vdd.n238 vdd.n237 10.7238
R19415 vdd.n195 vdd.n194 10.7238
R19416 vdd.n140 vdd.n139 10.7238
R19417 vdd.n98 vdd.n97 10.7238
R19418 vdd.n43 vdd.n42 10.7238
R19419 vdd.n1662 vdd.n1661 10.7238
R19420 vdd.n1717 vdd.n1716 10.7238
R19421 vdd.n1564 vdd.n1563 10.7238
R19422 vdd.n1619 vdd.n1618 10.7238
R19423 vdd.n1467 vdd.n1466 10.7238
R19424 vdd.n1522 vdd.n1521 10.7238
R19425 vdd.n2295 vdd.n2294 10.6151
R19426 vdd.n2296 vdd.n2295 10.6151
R19427 vdd.n2296 vdd.n1006 10.6151
R19428 vdd.n2306 vdd.n1006 10.6151
R19429 vdd.n2307 vdd.n2306 10.6151
R19430 vdd.n2308 vdd.n2307 10.6151
R19431 vdd.n2308 vdd.n993 10.6151
R19432 vdd.n2319 vdd.n993 10.6151
R19433 vdd.n2320 vdd.n2319 10.6151
R19434 vdd.n2321 vdd.n2320 10.6151
R19435 vdd.n2321 vdd.n981 10.6151
R19436 vdd.n2331 vdd.n981 10.6151
R19437 vdd.n2332 vdd.n2331 10.6151
R19438 vdd.n2333 vdd.n2332 10.6151
R19439 vdd.n2333 vdd.n969 10.6151
R19440 vdd.n2343 vdd.n969 10.6151
R19441 vdd.n2344 vdd.n2343 10.6151
R19442 vdd.n2345 vdd.n2344 10.6151
R19443 vdd.n2345 vdd.n958 10.6151
R19444 vdd.n2355 vdd.n958 10.6151
R19445 vdd.n2356 vdd.n2355 10.6151
R19446 vdd.n2357 vdd.n2356 10.6151
R19447 vdd.n2357 vdd.n945 10.6151
R19448 vdd.n2369 vdd.n945 10.6151
R19449 vdd.n2370 vdd.n2369 10.6151
R19450 vdd.n2372 vdd.n2370 10.6151
R19451 vdd.n2372 vdd.n2371 10.6151
R19452 vdd.n2371 vdd.n927 10.6151
R19453 vdd.n2519 vdd.n2518 10.6151
R19454 vdd.n2518 vdd.n2517 10.6151
R19455 vdd.n2517 vdd.n2514 10.6151
R19456 vdd.n2514 vdd.n2513 10.6151
R19457 vdd.n2513 vdd.n2510 10.6151
R19458 vdd.n2510 vdd.n2509 10.6151
R19459 vdd.n2509 vdd.n2506 10.6151
R19460 vdd.n2506 vdd.n2505 10.6151
R19461 vdd.n2505 vdd.n2502 10.6151
R19462 vdd.n2502 vdd.n2501 10.6151
R19463 vdd.n2501 vdd.n2498 10.6151
R19464 vdd.n2498 vdd.n2497 10.6151
R19465 vdd.n2497 vdd.n2494 10.6151
R19466 vdd.n2494 vdd.n2493 10.6151
R19467 vdd.n2493 vdd.n2490 10.6151
R19468 vdd.n2490 vdd.n2489 10.6151
R19469 vdd.n2489 vdd.n2486 10.6151
R19470 vdd.n2486 vdd.n2485 10.6151
R19471 vdd.n2485 vdd.n2482 10.6151
R19472 vdd.n2482 vdd.n2481 10.6151
R19473 vdd.n2481 vdd.n2478 10.6151
R19474 vdd.n2478 vdd.n2477 10.6151
R19475 vdd.n2477 vdd.n2474 10.6151
R19476 vdd.n2474 vdd.n2473 10.6151
R19477 vdd.n2473 vdd.n2470 10.6151
R19478 vdd.n2470 vdd.n2469 10.6151
R19479 vdd.n2469 vdd.n2466 10.6151
R19480 vdd.n2466 vdd.n2465 10.6151
R19481 vdd.n2465 vdd.n2462 10.6151
R19482 vdd.n2462 vdd.n2461 10.6151
R19483 vdd.n2461 vdd.n2458 10.6151
R19484 vdd.n2456 vdd.n2453 10.6151
R19485 vdd.n2453 vdd.n2452 10.6151
R19486 vdd.n2195 vdd.n2194 10.6151
R19487 vdd.n2194 vdd.n2192 10.6151
R19488 vdd.n2192 vdd.n2191 10.6151
R19489 vdd.n2191 vdd.n2189 10.6151
R19490 vdd.n2189 vdd.n2188 10.6151
R19491 vdd.n2188 vdd.n2186 10.6151
R19492 vdd.n2186 vdd.n2185 10.6151
R19493 vdd.n2185 vdd.n2183 10.6151
R19494 vdd.n2183 vdd.n2182 10.6151
R19495 vdd.n2182 vdd.n2180 10.6151
R19496 vdd.n2180 vdd.n2179 10.6151
R19497 vdd.n2179 vdd.n2177 10.6151
R19498 vdd.n2177 vdd.n2176 10.6151
R19499 vdd.n2176 vdd.n2091 10.6151
R19500 vdd.n2091 vdd.n2090 10.6151
R19501 vdd.n2090 vdd.n2088 10.6151
R19502 vdd.n2088 vdd.n2087 10.6151
R19503 vdd.n2087 vdd.n2085 10.6151
R19504 vdd.n2085 vdd.n2084 10.6151
R19505 vdd.n2084 vdd.n2082 10.6151
R19506 vdd.n2082 vdd.n2081 10.6151
R19507 vdd.n2081 vdd.n2079 10.6151
R19508 vdd.n2079 vdd.n2078 10.6151
R19509 vdd.n2078 vdd.n2076 10.6151
R19510 vdd.n2076 vdd.n2075 10.6151
R19511 vdd.n2075 vdd.n2072 10.6151
R19512 vdd.n2072 vdd.n2071 10.6151
R19513 vdd.n2071 vdd.n930 10.6151
R19514 vdd.n2029 vdd.n1018 10.6151
R19515 vdd.n2030 vdd.n2029 10.6151
R19516 vdd.n2031 vdd.n2030 10.6151
R19517 vdd.n2031 vdd.n2025 10.6151
R19518 vdd.n2037 vdd.n2025 10.6151
R19519 vdd.n2038 vdd.n2037 10.6151
R19520 vdd.n2039 vdd.n2038 10.6151
R19521 vdd.n2039 vdd.n2023 10.6151
R19522 vdd.n2045 vdd.n2023 10.6151
R19523 vdd.n2046 vdd.n2045 10.6151
R19524 vdd.n2047 vdd.n2046 10.6151
R19525 vdd.n2047 vdd.n2021 10.6151
R19526 vdd.n2053 vdd.n2021 10.6151
R19527 vdd.n2054 vdd.n2053 10.6151
R19528 vdd.n2055 vdd.n2054 10.6151
R19529 vdd.n2055 vdd.n2019 10.6151
R19530 vdd.n2231 vdd.n2019 10.6151
R19531 vdd.n2231 vdd.n2230 10.6151
R19532 vdd.n2230 vdd.n2060 10.6151
R19533 vdd.n2224 vdd.n2060 10.6151
R19534 vdd.n2224 vdd.n2223 10.6151
R19535 vdd.n2223 vdd.n2222 10.6151
R19536 vdd.n2222 vdd.n2062 10.6151
R19537 vdd.n2216 vdd.n2062 10.6151
R19538 vdd.n2216 vdd.n2215 10.6151
R19539 vdd.n2215 vdd.n2214 10.6151
R19540 vdd.n2214 vdd.n2064 10.6151
R19541 vdd.n2208 vdd.n2064 10.6151
R19542 vdd.n2208 vdd.n2207 10.6151
R19543 vdd.n2207 vdd.n2206 10.6151
R19544 vdd.n2206 vdd.n2066 10.6151
R19545 vdd.n2200 vdd.n2199 10.6151
R19546 vdd.n2199 vdd.n2198 10.6151
R19547 vdd.n2704 vdd.n2703 10.6151
R19548 vdd.n2703 vdd.n2701 10.6151
R19549 vdd.n2701 vdd.n2700 10.6151
R19550 vdd.n2700 vdd.n2558 10.6151
R19551 vdd.n2647 vdd.n2558 10.6151
R19552 vdd.n2648 vdd.n2647 10.6151
R19553 vdd.n2650 vdd.n2648 10.6151
R19554 vdd.n2651 vdd.n2650 10.6151
R19555 vdd.n2653 vdd.n2651 10.6151
R19556 vdd.n2654 vdd.n2653 10.6151
R19557 vdd.n2656 vdd.n2654 10.6151
R19558 vdd.n2657 vdd.n2656 10.6151
R19559 vdd.n2659 vdd.n2657 10.6151
R19560 vdd.n2660 vdd.n2659 10.6151
R19561 vdd.n2675 vdd.n2660 10.6151
R19562 vdd.n2675 vdd.n2674 10.6151
R19563 vdd.n2674 vdd.n2673 10.6151
R19564 vdd.n2673 vdd.n2671 10.6151
R19565 vdd.n2671 vdd.n2670 10.6151
R19566 vdd.n2670 vdd.n2668 10.6151
R19567 vdd.n2668 vdd.n2667 10.6151
R19568 vdd.n2667 vdd.n2665 10.6151
R19569 vdd.n2665 vdd.n2664 10.6151
R19570 vdd.n2664 vdd.n2662 10.6151
R19571 vdd.n2662 vdd.n2661 10.6151
R19572 vdd.n2661 vdd.n807 10.6151
R19573 vdd.n2909 vdd.n807 10.6151
R19574 vdd.n2910 vdd.n2909 10.6151
R19575 vdd.n2771 vdd.n883 10.6151
R19576 vdd.n2771 vdd.n2770 10.6151
R19577 vdd.n2770 vdd.n2769 10.6151
R19578 vdd.n2769 vdd.n2767 10.6151
R19579 vdd.n2767 vdd.n2764 10.6151
R19580 vdd.n2764 vdd.n2763 10.6151
R19581 vdd.n2763 vdd.n2760 10.6151
R19582 vdd.n2760 vdd.n2759 10.6151
R19583 vdd.n2759 vdd.n2756 10.6151
R19584 vdd.n2756 vdd.n2755 10.6151
R19585 vdd.n2755 vdd.n2752 10.6151
R19586 vdd.n2752 vdd.n2751 10.6151
R19587 vdd.n2751 vdd.n2748 10.6151
R19588 vdd.n2748 vdd.n2747 10.6151
R19589 vdd.n2747 vdd.n2744 10.6151
R19590 vdd.n2744 vdd.n2743 10.6151
R19591 vdd.n2743 vdd.n2740 10.6151
R19592 vdd.n2740 vdd.n2739 10.6151
R19593 vdd.n2739 vdd.n2736 10.6151
R19594 vdd.n2736 vdd.n2735 10.6151
R19595 vdd.n2735 vdd.n2732 10.6151
R19596 vdd.n2732 vdd.n2731 10.6151
R19597 vdd.n2731 vdd.n2728 10.6151
R19598 vdd.n2728 vdd.n2727 10.6151
R19599 vdd.n2727 vdd.n2724 10.6151
R19600 vdd.n2724 vdd.n2723 10.6151
R19601 vdd.n2723 vdd.n2720 10.6151
R19602 vdd.n2720 vdd.n2719 10.6151
R19603 vdd.n2719 vdd.n2716 10.6151
R19604 vdd.n2716 vdd.n2715 10.6151
R19605 vdd.n2715 vdd.n2712 10.6151
R19606 vdd.n2710 vdd.n2707 10.6151
R19607 vdd.n2707 vdd.n2706 10.6151
R19608 vdd.n2784 vdd.n2783 10.6151
R19609 vdd.n2785 vdd.n2784 10.6151
R19610 vdd.n2785 vdd.n873 10.6151
R19611 vdd.n2795 vdd.n873 10.6151
R19612 vdd.n2796 vdd.n2795 10.6151
R19613 vdd.n2797 vdd.n2796 10.6151
R19614 vdd.n2797 vdd.n860 10.6151
R19615 vdd.n2807 vdd.n860 10.6151
R19616 vdd.n2808 vdd.n2807 10.6151
R19617 vdd.n2809 vdd.n2808 10.6151
R19618 vdd.n2809 vdd.n849 10.6151
R19619 vdd.n2819 vdd.n849 10.6151
R19620 vdd.n2820 vdd.n2819 10.6151
R19621 vdd.n2821 vdd.n2820 10.6151
R19622 vdd.n2821 vdd.n837 10.6151
R19623 vdd.n2831 vdd.n837 10.6151
R19624 vdd.n2832 vdd.n2831 10.6151
R19625 vdd.n2833 vdd.n2832 10.6151
R19626 vdd.n2833 vdd.n826 10.6151
R19627 vdd.n2845 vdd.n826 10.6151
R19628 vdd.n2846 vdd.n2845 10.6151
R19629 vdd.n2847 vdd.n2846 10.6151
R19630 vdd.n2847 vdd.n812 10.6151
R19631 vdd.n2902 vdd.n812 10.6151
R19632 vdd.n2903 vdd.n2902 10.6151
R19633 vdd.n2904 vdd.n2903 10.6151
R19634 vdd.n2904 vdd.n779 10.6151
R19635 vdd.n2974 vdd.n779 10.6151
R19636 vdd.n2973 vdd.n2972 10.6151
R19637 vdd.n2972 vdd.n780 10.6151
R19638 vdd.n781 vdd.n780 10.6151
R19639 vdd.n2965 vdd.n781 10.6151
R19640 vdd.n2965 vdd.n2964 10.6151
R19641 vdd.n2964 vdd.n2963 10.6151
R19642 vdd.n2963 vdd.n783 10.6151
R19643 vdd.n2958 vdd.n783 10.6151
R19644 vdd.n2958 vdd.n2957 10.6151
R19645 vdd.n2957 vdd.n2956 10.6151
R19646 vdd.n2956 vdd.n786 10.6151
R19647 vdd.n2951 vdd.n786 10.6151
R19648 vdd.n2951 vdd.n2950 10.6151
R19649 vdd.n2950 vdd.n2949 10.6151
R19650 vdd.n2949 vdd.n789 10.6151
R19651 vdd.n2944 vdd.n789 10.6151
R19652 vdd.n2944 vdd.n2943 10.6151
R19653 vdd.n2943 vdd.n2941 10.6151
R19654 vdd.n2941 vdd.n792 10.6151
R19655 vdd.n2936 vdd.n792 10.6151
R19656 vdd.n2936 vdd.n2935 10.6151
R19657 vdd.n2935 vdd.n2934 10.6151
R19658 vdd.n2934 vdd.n795 10.6151
R19659 vdd.n2929 vdd.n795 10.6151
R19660 vdd.n2929 vdd.n2928 10.6151
R19661 vdd.n2928 vdd.n2927 10.6151
R19662 vdd.n2927 vdd.n798 10.6151
R19663 vdd.n2922 vdd.n798 10.6151
R19664 vdd.n2922 vdd.n2921 10.6151
R19665 vdd.n2921 vdd.n2920 10.6151
R19666 vdd.n2920 vdd.n801 10.6151
R19667 vdd.n2915 vdd.n2914 10.6151
R19668 vdd.n2914 vdd.n2913 10.6151
R19669 vdd.n2892 vdd.n2853 10.6151
R19670 vdd.n2887 vdd.n2853 10.6151
R19671 vdd.n2887 vdd.n2886 10.6151
R19672 vdd.n2886 vdd.n2885 10.6151
R19673 vdd.n2885 vdd.n2855 10.6151
R19674 vdd.n2880 vdd.n2855 10.6151
R19675 vdd.n2880 vdd.n2879 10.6151
R19676 vdd.n2879 vdd.n2878 10.6151
R19677 vdd.n2878 vdd.n2858 10.6151
R19678 vdd.n2873 vdd.n2858 10.6151
R19679 vdd.n2873 vdd.n2872 10.6151
R19680 vdd.n2872 vdd.n2871 10.6151
R19681 vdd.n2871 vdd.n2861 10.6151
R19682 vdd.n2866 vdd.n2861 10.6151
R19683 vdd.n2866 vdd.n2865 10.6151
R19684 vdd.n2865 vdd.n753 10.6151
R19685 vdd.n3009 vdd.n753 10.6151
R19686 vdd.n3009 vdd.n754 10.6151
R19687 vdd.n757 vdd.n754 10.6151
R19688 vdd.n3002 vdd.n757 10.6151
R19689 vdd.n3002 vdd.n3001 10.6151
R19690 vdd.n3001 vdd.n3000 10.6151
R19691 vdd.n3000 vdd.n759 10.6151
R19692 vdd.n2995 vdd.n759 10.6151
R19693 vdd.n2995 vdd.n2994 10.6151
R19694 vdd.n2994 vdd.n2993 10.6151
R19695 vdd.n2993 vdd.n762 10.6151
R19696 vdd.n2988 vdd.n762 10.6151
R19697 vdd.n2988 vdd.n2987 10.6151
R19698 vdd.n2987 vdd.n2986 10.6151
R19699 vdd.n2986 vdd.n765 10.6151
R19700 vdd.n2981 vdd.n2980 10.6151
R19701 vdd.n2980 vdd.n2979 10.6151
R19702 vdd.n2627 vdd.n2625 10.6151
R19703 vdd.n2628 vdd.n2627 10.6151
R19704 vdd.n2696 vdd.n2628 10.6151
R19705 vdd.n2696 vdd.n2695 10.6151
R19706 vdd.n2695 vdd.n2694 10.6151
R19707 vdd.n2694 vdd.n2692 10.6151
R19708 vdd.n2692 vdd.n2691 10.6151
R19709 vdd.n2691 vdd.n2689 10.6151
R19710 vdd.n2689 vdd.n2688 10.6151
R19711 vdd.n2688 vdd.n2686 10.6151
R19712 vdd.n2686 vdd.n2685 10.6151
R19713 vdd.n2685 vdd.n2683 10.6151
R19714 vdd.n2683 vdd.n2682 10.6151
R19715 vdd.n2682 vdd.n2680 10.6151
R19716 vdd.n2680 vdd.n2679 10.6151
R19717 vdd.n2679 vdd.n2645 10.6151
R19718 vdd.n2645 vdd.n2644 10.6151
R19719 vdd.n2644 vdd.n2642 10.6151
R19720 vdd.n2642 vdd.n2641 10.6151
R19721 vdd.n2641 vdd.n2639 10.6151
R19722 vdd.n2639 vdd.n2638 10.6151
R19723 vdd.n2638 vdd.n2636 10.6151
R19724 vdd.n2636 vdd.n2635 10.6151
R19725 vdd.n2635 vdd.n2633 10.6151
R19726 vdd.n2633 vdd.n2632 10.6151
R19727 vdd.n2632 vdd.n2630 10.6151
R19728 vdd.n2630 vdd.n2629 10.6151
R19729 vdd.n2629 vdd.n771 10.6151
R19730 vdd.n2778 vdd.n2777 10.6151
R19731 vdd.n2777 vdd.n888 10.6151
R19732 vdd.n2562 vdd.n888 10.6151
R19733 vdd.n2565 vdd.n2562 10.6151
R19734 vdd.n2566 vdd.n2565 10.6151
R19735 vdd.n2569 vdd.n2566 10.6151
R19736 vdd.n2570 vdd.n2569 10.6151
R19737 vdd.n2573 vdd.n2570 10.6151
R19738 vdd.n2574 vdd.n2573 10.6151
R19739 vdd.n2577 vdd.n2574 10.6151
R19740 vdd.n2578 vdd.n2577 10.6151
R19741 vdd.n2581 vdd.n2578 10.6151
R19742 vdd.n2582 vdd.n2581 10.6151
R19743 vdd.n2585 vdd.n2582 10.6151
R19744 vdd.n2586 vdd.n2585 10.6151
R19745 vdd.n2589 vdd.n2586 10.6151
R19746 vdd.n2590 vdd.n2589 10.6151
R19747 vdd.n2593 vdd.n2590 10.6151
R19748 vdd.n2594 vdd.n2593 10.6151
R19749 vdd.n2597 vdd.n2594 10.6151
R19750 vdd.n2598 vdd.n2597 10.6151
R19751 vdd.n2601 vdd.n2598 10.6151
R19752 vdd.n2602 vdd.n2601 10.6151
R19753 vdd.n2605 vdd.n2602 10.6151
R19754 vdd.n2606 vdd.n2605 10.6151
R19755 vdd.n2609 vdd.n2606 10.6151
R19756 vdd.n2610 vdd.n2609 10.6151
R19757 vdd.n2613 vdd.n2610 10.6151
R19758 vdd.n2614 vdd.n2613 10.6151
R19759 vdd.n2617 vdd.n2614 10.6151
R19760 vdd.n2618 vdd.n2617 10.6151
R19761 vdd.n2623 vdd.n2621 10.6151
R19762 vdd.n2624 vdd.n2623 10.6151
R19763 vdd.n2779 vdd.n878 10.6151
R19764 vdd.n2789 vdd.n878 10.6151
R19765 vdd.n2790 vdd.n2789 10.6151
R19766 vdd.n2791 vdd.n2790 10.6151
R19767 vdd.n2791 vdd.n866 10.6151
R19768 vdd.n2801 vdd.n866 10.6151
R19769 vdd.n2802 vdd.n2801 10.6151
R19770 vdd.n2803 vdd.n2802 10.6151
R19771 vdd.n2803 vdd.n855 10.6151
R19772 vdd.n2813 vdd.n855 10.6151
R19773 vdd.n2814 vdd.n2813 10.6151
R19774 vdd.n2815 vdd.n2814 10.6151
R19775 vdd.n2815 vdd.n843 10.6151
R19776 vdd.n2825 vdd.n843 10.6151
R19777 vdd.n2826 vdd.n2825 10.6151
R19778 vdd.n2827 vdd.n2826 10.6151
R19779 vdd.n2827 vdd.n832 10.6151
R19780 vdd.n2837 vdd.n832 10.6151
R19781 vdd.n2838 vdd.n2837 10.6151
R19782 vdd.n2841 vdd.n2838 10.6151
R19783 vdd.n2851 vdd.n820 10.6151
R19784 vdd.n2852 vdd.n2851 10.6151
R19785 vdd.n2898 vdd.n2852 10.6151
R19786 vdd.n2898 vdd.n2897 10.6151
R19787 vdd.n2897 vdd.n2896 10.6151
R19788 vdd.n2896 vdd.n2895 10.6151
R19789 vdd.n2895 vdd.n2893 10.6151
R19790 vdd.n2290 vdd.n1012 10.6151
R19791 vdd.n2300 vdd.n1012 10.6151
R19792 vdd.n2301 vdd.n2300 10.6151
R19793 vdd.n2302 vdd.n2301 10.6151
R19794 vdd.n2302 vdd.n999 10.6151
R19795 vdd.n2312 vdd.n999 10.6151
R19796 vdd.n2313 vdd.n2312 10.6151
R19797 vdd.n2315 vdd.n987 10.6151
R19798 vdd.n2325 vdd.n987 10.6151
R19799 vdd.n2326 vdd.n2325 10.6151
R19800 vdd.n2327 vdd.n2326 10.6151
R19801 vdd.n2327 vdd.n975 10.6151
R19802 vdd.n2337 vdd.n975 10.6151
R19803 vdd.n2338 vdd.n2337 10.6151
R19804 vdd.n2339 vdd.n2338 10.6151
R19805 vdd.n2339 vdd.n964 10.6151
R19806 vdd.n2349 vdd.n964 10.6151
R19807 vdd.n2350 vdd.n2349 10.6151
R19808 vdd.n2351 vdd.n2350 10.6151
R19809 vdd.n2351 vdd.n952 10.6151
R19810 vdd.n2361 vdd.n952 10.6151
R19811 vdd.n2362 vdd.n2361 10.6151
R19812 vdd.n2365 vdd.n2362 10.6151
R19813 vdd.n2365 vdd.n2364 10.6151
R19814 vdd.n2364 vdd.n2363 10.6151
R19815 vdd.n2363 vdd.n935 10.6151
R19816 vdd.n2447 vdd.n935 10.6151
R19817 vdd.n2446 vdd.n2445 10.6151
R19818 vdd.n2445 vdd.n2442 10.6151
R19819 vdd.n2442 vdd.n2441 10.6151
R19820 vdd.n2441 vdd.n2438 10.6151
R19821 vdd.n2438 vdd.n2437 10.6151
R19822 vdd.n2437 vdd.n2434 10.6151
R19823 vdd.n2434 vdd.n2433 10.6151
R19824 vdd.n2433 vdd.n2430 10.6151
R19825 vdd.n2430 vdd.n2429 10.6151
R19826 vdd.n2429 vdd.n2426 10.6151
R19827 vdd.n2426 vdd.n2425 10.6151
R19828 vdd.n2425 vdd.n2422 10.6151
R19829 vdd.n2422 vdd.n2421 10.6151
R19830 vdd.n2421 vdd.n2418 10.6151
R19831 vdd.n2418 vdd.n2417 10.6151
R19832 vdd.n2417 vdd.n2414 10.6151
R19833 vdd.n2414 vdd.n2413 10.6151
R19834 vdd.n2413 vdd.n2410 10.6151
R19835 vdd.n2410 vdd.n2409 10.6151
R19836 vdd.n2409 vdd.n2406 10.6151
R19837 vdd.n2406 vdd.n2405 10.6151
R19838 vdd.n2405 vdd.n2402 10.6151
R19839 vdd.n2402 vdd.n2401 10.6151
R19840 vdd.n2401 vdd.n2398 10.6151
R19841 vdd.n2398 vdd.n2397 10.6151
R19842 vdd.n2397 vdd.n2394 10.6151
R19843 vdd.n2394 vdd.n2393 10.6151
R19844 vdd.n2393 vdd.n2390 10.6151
R19845 vdd.n2390 vdd.n2389 10.6151
R19846 vdd.n2389 vdd.n2386 10.6151
R19847 vdd.n2386 vdd.n2385 10.6151
R19848 vdd.n2382 vdd.n2381 10.6151
R19849 vdd.n2381 vdd.n2379 10.6151
R19850 vdd.n2138 vdd.n2136 10.6151
R19851 vdd.n2139 vdd.n2138 10.6151
R19852 vdd.n2141 vdd.n2139 10.6151
R19853 vdd.n2142 vdd.n2141 10.6151
R19854 vdd.n2144 vdd.n2142 10.6151
R19855 vdd.n2145 vdd.n2144 10.6151
R19856 vdd.n2147 vdd.n2145 10.6151
R19857 vdd.n2148 vdd.n2147 10.6151
R19858 vdd.n2150 vdd.n2148 10.6151
R19859 vdd.n2151 vdd.n2150 10.6151
R19860 vdd.n2153 vdd.n2151 10.6151
R19861 vdd.n2154 vdd.n2153 10.6151
R19862 vdd.n2172 vdd.n2154 10.6151
R19863 vdd.n2172 vdd.n2171 10.6151
R19864 vdd.n2171 vdd.n2170 10.6151
R19865 vdd.n2170 vdd.n2168 10.6151
R19866 vdd.n2168 vdd.n2167 10.6151
R19867 vdd.n2167 vdd.n2165 10.6151
R19868 vdd.n2165 vdd.n2164 10.6151
R19869 vdd.n2164 vdd.n2162 10.6151
R19870 vdd.n2162 vdd.n2161 10.6151
R19871 vdd.n2161 vdd.n2159 10.6151
R19872 vdd.n2159 vdd.n2158 10.6151
R19873 vdd.n2158 vdd.n2156 10.6151
R19874 vdd.n2156 vdd.n2155 10.6151
R19875 vdd.n2155 vdd.n939 10.6151
R19876 vdd.n2377 vdd.n939 10.6151
R19877 vdd.n2378 vdd.n2377 10.6151
R19878 vdd.n2289 vdd.n2288 10.6151
R19879 vdd.n2288 vdd.n1024 10.6151
R19880 vdd.n2282 vdd.n1024 10.6151
R19881 vdd.n2282 vdd.n2281 10.6151
R19882 vdd.n2281 vdd.n2280 10.6151
R19883 vdd.n2280 vdd.n1026 10.6151
R19884 vdd.n2274 vdd.n1026 10.6151
R19885 vdd.n2274 vdd.n2273 10.6151
R19886 vdd.n2273 vdd.n2272 10.6151
R19887 vdd.n2272 vdd.n1028 10.6151
R19888 vdd.n2266 vdd.n1028 10.6151
R19889 vdd.n2266 vdd.n2265 10.6151
R19890 vdd.n2265 vdd.n2264 10.6151
R19891 vdd.n2264 vdd.n1030 10.6151
R19892 vdd.n2258 vdd.n1030 10.6151
R19893 vdd.n2258 vdd.n2257 10.6151
R19894 vdd.n2257 vdd.n2256 10.6151
R19895 vdd.n2256 vdd.n1034 10.6151
R19896 vdd.n2104 vdd.n1034 10.6151
R19897 vdd.n2105 vdd.n2104 10.6151
R19898 vdd.n2105 vdd.n2100 10.6151
R19899 vdd.n2111 vdd.n2100 10.6151
R19900 vdd.n2112 vdd.n2111 10.6151
R19901 vdd.n2113 vdd.n2112 10.6151
R19902 vdd.n2113 vdd.n2098 10.6151
R19903 vdd.n2119 vdd.n2098 10.6151
R19904 vdd.n2120 vdd.n2119 10.6151
R19905 vdd.n2121 vdd.n2120 10.6151
R19906 vdd.n2121 vdd.n2096 10.6151
R19907 vdd.n2127 vdd.n2096 10.6151
R19908 vdd.n2128 vdd.n2127 10.6151
R19909 vdd.n2130 vdd.n2092 10.6151
R19910 vdd.n2135 vdd.n2092 10.6151
R19911 vdd.t106 vdd.n1776 10.5435
R19912 vdd.n636 vdd.t25 10.5435
R19913 vdd.n304 vdd.n286 10.4732
R19914 vdd.n249 vdd.n231 10.4732
R19915 vdd.n206 vdd.n188 10.4732
R19916 vdd.n151 vdd.n133 10.4732
R19917 vdd.n109 vdd.n91 10.4732
R19918 vdd.n54 vdd.n36 10.4732
R19919 vdd.n1673 vdd.n1655 10.4732
R19920 vdd.n1728 vdd.n1710 10.4732
R19921 vdd.n1575 vdd.n1557 10.4732
R19922 vdd.n1630 vdd.n1612 10.4732
R19923 vdd.n1478 vdd.n1460 10.4732
R19924 vdd.n1533 vdd.n1515 10.4732
R19925 vdd.n1760 vdd.t74 10.3167
R19926 vdd.n3205 vdd.t43 10.3167
R19927 vdd.t27 vdd.n1104 10.09
R19928 vdd.n1812 vdd.t180 10.09
R19929 vdd.n3153 vdd.t165 10.09
R19930 vdd.n3286 vdd.t29 10.09
R19931 vdd.n1424 vdd.t50 9.86327
R19932 vdd.n3277 vdd.t84 9.86327
R19933 vdd.n303 vdd.n288 9.69747
R19934 vdd.n248 vdd.n233 9.69747
R19935 vdd.n205 vdd.n190 9.69747
R19936 vdd.n150 vdd.n135 9.69747
R19937 vdd.n108 vdd.n93 9.69747
R19938 vdd.n53 vdd.n38 9.69747
R19939 vdd.n1672 vdd.n1657 9.69747
R19940 vdd.n1727 vdd.n1712 9.69747
R19941 vdd.n1574 vdd.n1559 9.69747
R19942 vdd.n1629 vdd.n1614 9.69747
R19943 vdd.n1477 vdd.n1462 9.69747
R19944 vdd.n1532 vdd.n1517 9.69747
R19945 vdd.n2232 vdd.n2231 9.67831
R19946 vdd.n2943 vdd.n2942 9.67831
R19947 vdd.n3010 vdd.n3009 9.67831
R19948 vdd.n2256 vdd.n2255 9.67831
R19949 vdd.t31 vdd.n1398 9.63654
R19950 vdd.n3236 vdd.t41 9.63654
R19951 vdd.n319 vdd.n318 9.45567
R19952 vdd.n264 vdd.n263 9.45567
R19953 vdd.n221 vdd.n220 9.45567
R19954 vdd.n166 vdd.n165 9.45567
R19955 vdd.n124 vdd.n123 9.45567
R19956 vdd.n69 vdd.n68 9.45567
R19957 vdd.n1688 vdd.n1687 9.45567
R19958 vdd.n1743 vdd.n1742 9.45567
R19959 vdd.n1590 vdd.n1589 9.45567
R19960 vdd.n1645 vdd.n1644 9.45567
R19961 vdd.n1493 vdd.n1492 9.45567
R19962 vdd.n1548 vdd.n1547 9.45567
R19963 vdd.n1992 vdd.n1846 9.3005
R19964 vdd.n1991 vdd.n1990 9.3005
R19965 vdd.n1852 vdd.n1851 9.3005
R19966 vdd.n1985 vdd.n1856 9.3005
R19967 vdd.n1984 vdd.n1857 9.3005
R19968 vdd.n1983 vdd.n1858 9.3005
R19969 vdd.n1862 vdd.n1859 9.3005
R19970 vdd.n1978 vdd.n1863 9.3005
R19971 vdd.n1977 vdd.n1864 9.3005
R19972 vdd.n1976 vdd.n1865 9.3005
R19973 vdd.n1869 vdd.n1866 9.3005
R19974 vdd.n1971 vdd.n1870 9.3005
R19975 vdd.n1970 vdd.n1871 9.3005
R19976 vdd.n1969 vdd.n1872 9.3005
R19977 vdd.n1876 vdd.n1873 9.3005
R19978 vdd.n1964 vdd.n1877 9.3005
R19979 vdd.n1963 vdd.n1878 9.3005
R19980 vdd.n1962 vdd.n1879 9.3005
R19981 vdd.n1883 vdd.n1880 9.3005
R19982 vdd.n1957 vdd.n1884 9.3005
R19983 vdd.n1956 vdd.n1885 9.3005
R19984 vdd.n1955 vdd.n1954 9.3005
R19985 vdd.n1953 vdd.n1886 9.3005
R19986 vdd.n1952 vdd.n1951 9.3005
R19987 vdd.n1892 vdd.n1891 9.3005
R19988 vdd.n1946 vdd.n1896 9.3005
R19989 vdd.n1945 vdd.n1897 9.3005
R19990 vdd.n1944 vdd.n1898 9.3005
R19991 vdd.n1902 vdd.n1899 9.3005
R19992 vdd.n1939 vdd.n1903 9.3005
R19993 vdd.n1938 vdd.n1904 9.3005
R19994 vdd.n1937 vdd.n1905 9.3005
R19995 vdd.n1909 vdd.n1906 9.3005
R19996 vdd.n1932 vdd.n1910 9.3005
R19997 vdd.n1931 vdd.n1911 9.3005
R19998 vdd.n1930 vdd.n1912 9.3005
R19999 vdd.n1914 vdd.n1913 9.3005
R20000 vdd.n1925 vdd.n1035 9.3005
R20001 vdd.n1994 vdd.n1993 9.3005
R20002 vdd.n2018 vdd.n2017 9.3005
R20003 vdd.n1824 vdd.n1823 9.3005
R20004 vdd.n1829 vdd.n1827 9.3005
R20005 vdd.n2010 vdd.n1830 9.3005
R20006 vdd.n2009 vdd.n1831 9.3005
R20007 vdd.n2008 vdd.n1832 9.3005
R20008 vdd.n1836 vdd.n1833 9.3005
R20009 vdd.n2003 vdd.n1837 9.3005
R20010 vdd.n2002 vdd.n1838 9.3005
R20011 vdd.n2001 vdd.n1839 9.3005
R20012 vdd.n1843 vdd.n1840 9.3005
R20013 vdd.n1996 vdd.n1844 9.3005
R20014 vdd.n1995 vdd.n1845 9.3005
R20015 vdd.n2240 vdd.n1817 9.3005
R20016 vdd.n2242 vdd.n2241 9.3005
R20017 vdd.n1748 vdd.n1094 9.3005
R20018 vdd.n1750 vdd.n1749 9.3005
R20019 vdd.n1085 vdd.n1084 9.3005
R20020 vdd.n1763 vdd.n1762 9.3005
R20021 vdd.n1764 vdd.n1083 9.3005
R20022 vdd.n1766 vdd.n1765 9.3005
R20023 vdd.n1073 vdd.n1072 9.3005
R20024 vdd.n1780 vdd.n1779 9.3005
R20025 vdd.n1781 vdd.n1071 9.3005
R20026 vdd.n1783 vdd.n1782 9.3005
R20027 vdd.n1062 vdd.n1061 9.3005
R20028 vdd.n1797 vdd.n1796 9.3005
R20029 vdd.n1798 vdd.n1060 9.3005
R20030 vdd.n1800 vdd.n1799 9.3005
R20031 vdd.n1050 vdd.n1049 9.3005
R20032 vdd.n1815 vdd.n1814 9.3005
R20033 vdd.n1816 vdd.n1048 9.3005
R20034 vdd.n2244 vdd.n2243 9.3005
R20035 vdd.n295 vdd.n294 9.3005
R20036 vdd.n290 vdd.n289 9.3005
R20037 vdd.n301 vdd.n300 9.3005
R20038 vdd.n303 vdd.n302 9.3005
R20039 vdd.n286 vdd.n285 9.3005
R20040 vdd.n309 vdd.n308 9.3005
R20041 vdd.n311 vdd.n310 9.3005
R20042 vdd.n283 vdd.n280 9.3005
R20043 vdd.n318 vdd.n317 9.3005
R20044 vdd.n240 vdd.n239 9.3005
R20045 vdd.n235 vdd.n234 9.3005
R20046 vdd.n246 vdd.n245 9.3005
R20047 vdd.n248 vdd.n247 9.3005
R20048 vdd.n231 vdd.n230 9.3005
R20049 vdd.n254 vdd.n253 9.3005
R20050 vdd.n256 vdd.n255 9.3005
R20051 vdd.n228 vdd.n225 9.3005
R20052 vdd.n263 vdd.n262 9.3005
R20053 vdd.n197 vdd.n196 9.3005
R20054 vdd.n192 vdd.n191 9.3005
R20055 vdd.n203 vdd.n202 9.3005
R20056 vdd.n205 vdd.n204 9.3005
R20057 vdd.n188 vdd.n187 9.3005
R20058 vdd.n211 vdd.n210 9.3005
R20059 vdd.n213 vdd.n212 9.3005
R20060 vdd.n185 vdd.n182 9.3005
R20061 vdd.n220 vdd.n219 9.3005
R20062 vdd.n142 vdd.n141 9.3005
R20063 vdd.n137 vdd.n136 9.3005
R20064 vdd.n148 vdd.n147 9.3005
R20065 vdd.n150 vdd.n149 9.3005
R20066 vdd.n133 vdd.n132 9.3005
R20067 vdd.n156 vdd.n155 9.3005
R20068 vdd.n158 vdd.n157 9.3005
R20069 vdd.n130 vdd.n127 9.3005
R20070 vdd.n165 vdd.n164 9.3005
R20071 vdd.n100 vdd.n99 9.3005
R20072 vdd.n95 vdd.n94 9.3005
R20073 vdd.n106 vdd.n105 9.3005
R20074 vdd.n108 vdd.n107 9.3005
R20075 vdd.n91 vdd.n90 9.3005
R20076 vdd.n114 vdd.n113 9.3005
R20077 vdd.n116 vdd.n115 9.3005
R20078 vdd.n88 vdd.n85 9.3005
R20079 vdd.n123 vdd.n122 9.3005
R20080 vdd.n45 vdd.n44 9.3005
R20081 vdd.n40 vdd.n39 9.3005
R20082 vdd.n51 vdd.n50 9.3005
R20083 vdd.n53 vdd.n52 9.3005
R20084 vdd.n36 vdd.n35 9.3005
R20085 vdd.n59 vdd.n58 9.3005
R20086 vdd.n61 vdd.n60 9.3005
R20087 vdd.n33 vdd.n30 9.3005
R20088 vdd.n68 vdd.n67 9.3005
R20089 vdd.n3059 vdd.n3058 9.3005
R20090 vdd.n3060 vdd.n721 9.3005
R20091 vdd.n720 vdd.n718 9.3005
R20092 vdd.n3066 vdd.n717 9.3005
R20093 vdd.n3067 vdd.n716 9.3005
R20094 vdd.n3068 vdd.n715 9.3005
R20095 vdd.n714 vdd.n712 9.3005
R20096 vdd.n3074 vdd.n711 9.3005
R20097 vdd.n3075 vdd.n710 9.3005
R20098 vdd.n3076 vdd.n709 9.3005
R20099 vdd.n708 vdd.n706 9.3005
R20100 vdd.n3082 vdd.n705 9.3005
R20101 vdd.n3083 vdd.n704 9.3005
R20102 vdd.n3084 vdd.n703 9.3005
R20103 vdd.n702 vdd.n700 9.3005
R20104 vdd.n3090 vdd.n699 9.3005
R20105 vdd.n3091 vdd.n698 9.3005
R20106 vdd.n3092 vdd.n697 9.3005
R20107 vdd.n696 vdd.n694 9.3005
R20108 vdd.n3098 vdd.n693 9.3005
R20109 vdd.n3099 vdd.n692 9.3005
R20110 vdd.n3100 vdd.n691 9.3005
R20111 vdd.n690 vdd.n688 9.3005
R20112 vdd.n3106 vdd.n685 9.3005
R20113 vdd.n3107 vdd.n684 9.3005
R20114 vdd.n3108 vdd.n683 9.3005
R20115 vdd.n682 vdd.n680 9.3005
R20116 vdd.n3114 vdd.n679 9.3005
R20117 vdd.n3115 vdd.n678 9.3005
R20118 vdd.n3116 vdd.n677 9.3005
R20119 vdd.n676 vdd.n674 9.3005
R20120 vdd.n3122 vdd.n673 9.3005
R20121 vdd.n3123 vdd.n672 9.3005
R20122 vdd.n3124 vdd.n671 9.3005
R20123 vdd.n670 vdd.n668 9.3005
R20124 vdd.n3129 vdd.n667 9.3005
R20125 vdd.n3139 vdd.n661 9.3005
R20126 vdd.n3141 vdd.n3140 9.3005
R20127 vdd.n652 vdd.n651 9.3005
R20128 vdd.n3156 vdd.n3155 9.3005
R20129 vdd.n3157 vdd.n650 9.3005
R20130 vdd.n3159 vdd.n3158 9.3005
R20131 vdd.n640 vdd.n639 9.3005
R20132 vdd.n3172 vdd.n3171 9.3005
R20133 vdd.n3173 vdd.n638 9.3005
R20134 vdd.n3175 vdd.n3174 9.3005
R20135 vdd.n628 vdd.n627 9.3005
R20136 vdd.n3189 vdd.n3188 9.3005
R20137 vdd.n3190 vdd.n626 9.3005
R20138 vdd.n3192 vdd.n3191 9.3005
R20139 vdd.n617 vdd.n616 9.3005
R20140 vdd.n3208 vdd.n3207 9.3005
R20141 vdd.n3209 vdd.n615 9.3005
R20142 vdd.n3211 vdd.n3210 9.3005
R20143 vdd.n324 vdd.n322 9.3005
R20144 vdd.n3143 vdd.n3142 9.3005
R20145 vdd.n3290 vdd.n3289 9.3005
R20146 vdd.n325 vdd.n323 9.3005
R20147 vdd.n3283 vdd.n334 9.3005
R20148 vdd.n3282 vdd.n335 9.3005
R20149 vdd.n3281 vdd.n336 9.3005
R20150 vdd.n343 vdd.n337 9.3005
R20151 vdd.n3275 vdd.n344 9.3005
R20152 vdd.n3274 vdd.n345 9.3005
R20153 vdd.n3273 vdd.n346 9.3005
R20154 vdd.n354 vdd.n347 9.3005
R20155 vdd.n3267 vdd.n355 9.3005
R20156 vdd.n3266 vdd.n356 9.3005
R20157 vdd.n3265 vdd.n357 9.3005
R20158 vdd.n365 vdd.n358 9.3005
R20159 vdd.n3259 vdd.n366 9.3005
R20160 vdd.n3258 vdd.n367 9.3005
R20161 vdd.n3257 vdd.n368 9.3005
R20162 vdd.n443 vdd.n369 9.3005
R20163 vdd.n447 vdd.n442 9.3005
R20164 vdd.n451 vdd.n450 9.3005
R20165 vdd.n452 vdd.n441 9.3005
R20166 vdd.n456 vdd.n453 9.3005
R20167 vdd.n457 vdd.n440 9.3005
R20168 vdd.n461 vdd.n460 9.3005
R20169 vdd.n462 vdd.n439 9.3005
R20170 vdd.n466 vdd.n463 9.3005
R20171 vdd.n467 vdd.n438 9.3005
R20172 vdd.n471 vdd.n470 9.3005
R20173 vdd.n472 vdd.n437 9.3005
R20174 vdd.n476 vdd.n473 9.3005
R20175 vdd.n477 vdd.n436 9.3005
R20176 vdd.n481 vdd.n480 9.3005
R20177 vdd.n482 vdd.n435 9.3005
R20178 vdd.n486 vdd.n483 9.3005
R20179 vdd.n487 vdd.n434 9.3005
R20180 vdd.n491 vdd.n490 9.3005
R20181 vdd.n492 vdd.n433 9.3005
R20182 vdd.n496 vdd.n493 9.3005
R20183 vdd.n497 vdd.n430 9.3005
R20184 vdd.n501 vdd.n500 9.3005
R20185 vdd.n502 vdd.n429 9.3005
R20186 vdd.n506 vdd.n503 9.3005
R20187 vdd.n507 vdd.n428 9.3005
R20188 vdd.n511 vdd.n510 9.3005
R20189 vdd.n512 vdd.n427 9.3005
R20190 vdd.n516 vdd.n513 9.3005
R20191 vdd.n517 vdd.n426 9.3005
R20192 vdd.n521 vdd.n520 9.3005
R20193 vdd.n522 vdd.n425 9.3005
R20194 vdd.n526 vdd.n523 9.3005
R20195 vdd.n527 vdd.n424 9.3005
R20196 vdd.n531 vdd.n530 9.3005
R20197 vdd.n532 vdd.n423 9.3005
R20198 vdd.n536 vdd.n533 9.3005
R20199 vdd.n537 vdd.n422 9.3005
R20200 vdd.n541 vdd.n540 9.3005
R20201 vdd.n542 vdd.n421 9.3005
R20202 vdd.n546 vdd.n543 9.3005
R20203 vdd.n547 vdd.n418 9.3005
R20204 vdd.n551 vdd.n550 9.3005
R20205 vdd.n552 vdd.n417 9.3005
R20206 vdd.n556 vdd.n553 9.3005
R20207 vdd.n557 vdd.n416 9.3005
R20208 vdd.n561 vdd.n560 9.3005
R20209 vdd.n562 vdd.n415 9.3005
R20210 vdd.n566 vdd.n563 9.3005
R20211 vdd.n567 vdd.n414 9.3005
R20212 vdd.n571 vdd.n570 9.3005
R20213 vdd.n572 vdd.n413 9.3005
R20214 vdd.n576 vdd.n573 9.3005
R20215 vdd.n577 vdd.n412 9.3005
R20216 vdd.n581 vdd.n580 9.3005
R20217 vdd.n582 vdd.n411 9.3005
R20218 vdd.n586 vdd.n583 9.3005
R20219 vdd.n587 vdd.n410 9.3005
R20220 vdd.n591 vdd.n590 9.3005
R20221 vdd.n592 vdd.n409 9.3005
R20222 vdd.n596 vdd.n593 9.3005
R20223 vdd.n598 vdd.n408 9.3005
R20224 vdd.n600 vdd.n599 9.3005
R20225 vdd.n3250 vdd.n3249 9.3005
R20226 vdd.n446 vdd.n444 9.3005
R20227 vdd.n3149 vdd.n655 9.3005
R20228 vdd.n3151 vdd.n3150 9.3005
R20229 vdd.n646 vdd.n645 9.3005
R20230 vdd.n3164 vdd.n3163 9.3005
R20231 vdd.n3165 vdd.n644 9.3005
R20232 vdd.n3167 vdd.n3166 9.3005
R20233 vdd.n633 vdd.n632 9.3005
R20234 vdd.n3180 vdd.n3179 9.3005
R20235 vdd.n3181 vdd.n631 9.3005
R20236 vdd.n3183 vdd.n3182 9.3005
R20237 vdd.n622 vdd.n621 9.3005
R20238 vdd.n3197 vdd.n3196 9.3005
R20239 vdd.n3198 vdd.n620 9.3005
R20240 vdd.n3203 vdd.n3199 9.3005
R20241 vdd.n3202 vdd.n3201 9.3005
R20242 vdd.n3200 vdd.n610 9.3005
R20243 vdd.n3216 vdd.n611 9.3005
R20244 vdd.n3217 vdd.n609 9.3005
R20245 vdd.n3219 vdd.n3218 9.3005
R20246 vdd.n3220 vdd.n608 9.3005
R20247 vdd.n3223 vdd.n3221 9.3005
R20248 vdd.n3224 vdd.n607 9.3005
R20249 vdd.n3226 vdd.n3225 9.3005
R20250 vdd.n3227 vdd.n606 9.3005
R20251 vdd.n3230 vdd.n3228 9.3005
R20252 vdd.n3231 vdd.n605 9.3005
R20253 vdd.n3233 vdd.n3232 9.3005
R20254 vdd.n3234 vdd.n604 9.3005
R20255 vdd.n3238 vdd.n3235 9.3005
R20256 vdd.n3239 vdd.n603 9.3005
R20257 vdd.n3241 vdd.n3240 9.3005
R20258 vdd.n3242 vdd.n602 9.3005
R20259 vdd.n3245 vdd.n3243 9.3005
R20260 vdd.n3246 vdd.n601 9.3005
R20261 vdd.n3248 vdd.n3247 9.3005
R20262 vdd.n3148 vdd.n3147 9.3005
R20263 vdd.n3012 vdd.n656 9.3005
R20264 vdd.n3017 vdd.n3011 9.3005
R20265 vdd.n3027 vdd.n748 9.3005
R20266 vdd.n3028 vdd.n747 9.3005
R20267 vdd.n746 vdd.n744 9.3005
R20268 vdd.n3034 vdd.n743 9.3005
R20269 vdd.n3035 vdd.n742 9.3005
R20270 vdd.n3036 vdd.n741 9.3005
R20271 vdd.n740 vdd.n738 9.3005
R20272 vdd.n3042 vdd.n737 9.3005
R20273 vdd.n3043 vdd.n736 9.3005
R20274 vdd.n3044 vdd.n735 9.3005
R20275 vdd.n734 vdd.n732 9.3005
R20276 vdd.n3049 vdd.n731 9.3005
R20277 vdd.n3050 vdd.n730 9.3005
R20278 vdd.n726 vdd.n725 9.3005
R20279 vdd.n3056 vdd.n3055 9.3005
R20280 vdd.n3057 vdd.n722 9.3005
R20281 vdd.n2254 vdd.n2253 9.3005
R20282 vdd.n2249 vdd.n1038 9.3005
R20283 vdd.n1380 vdd.n1379 9.3005
R20284 vdd.n1136 vdd.n1135 9.3005
R20285 vdd.n1393 vdd.n1392 9.3005
R20286 vdd.n1394 vdd.n1134 9.3005
R20287 vdd.n1396 vdd.n1395 9.3005
R20288 vdd.n1124 vdd.n1123 9.3005
R20289 vdd.n1410 vdd.n1409 9.3005
R20290 vdd.n1411 vdd.n1122 9.3005
R20291 vdd.n1413 vdd.n1412 9.3005
R20292 vdd.n1114 vdd.n1113 9.3005
R20293 vdd.n1427 vdd.n1426 9.3005
R20294 vdd.n1428 vdd.n1112 9.3005
R20295 vdd.n1430 vdd.n1429 9.3005
R20296 vdd.n1101 vdd.n1100 9.3005
R20297 vdd.n1443 vdd.n1442 9.3005
R20298 vdd.n1444 vdd.n1099 9.3005
R20299 vdd.n1446 vdd.n1445 9.3005
R20300 vdd.n1090 vdd.n1089 9.3005
R20301 vdd.n1755 vdd.n1754 9.3005
R20302 vdd.n1756 vdd.n1088 9.3005
R20303 vdd.n1758 vdd.n1757 9.3005
R20304 vdd.n1079 vdd.n1078 9.3005
R20305 vdd.n1771 vdd.n1770 9.3005
R20306 vdd.n1772 vdd.n1077 9.3005
R20307 vdd.n1774 vdd.n1773 9.3005
R20308 vdd.n1067 vdd.n1066 9.3005
R20309 vdd.n1788 vdd.n1787 9.3005
R20310 vdd.n1789 vdd.n1065 9.3005
R20311 vdd.n1791 vdd.n1790 9.3005
R20312 vdd.n1057 vdd.n1056 9.3005
R20313 vdd.n1805 vdd.n1804 9.3005
R20314 vdd.n1806 vdd.n1054 9.3005
R20315 vdd.n1810 vdd.n1809 9.3005
R20316 vdd.n1808 vdd.n1055 9.3005
R20317 vdd.n1807 vdd.n1043 9.3005
R20318 vdd.n1378 vdd.n1146 9.3005
R20319 vdd.n1271 vdd.n1147 9.3005
R20320 vdd.n1273 vdd.n1272 9.3005
R20321 vdd.n1274 vdd.n1266 9.3005
R20322 vdd.n1276 vdd.n1275 9.3005
R20323 vdd.n1277 vdd.n1265 9.3005
R20324 vdd.n1279 vdd.n1278 9.3005
R20325 vdd.n1280 vdd.n1260 9.3005
R20326 vdd.n1282 vdd.n1281 9.3005
R20327 vdd.n1283 vdd.n1259 9.3005
R20328 vdd.n1285 vdd.n1284 9.3005
R20329 vdd.n1286 vdd.n1254 9.3005
R20330 vdd.n1288 vdd.n1287 9.3005
R20331 vdd.n1289 vdd.n1253 9.3005
R20332 vdd.n1291 vdd.n1290 9.3005
R20333 vdd.n1292 vdd.n1248 9.3005
R20334 vdd.n1294 vdd.n1293 9.3005
R20335 vdd.n1295 vdd.n1247 9.3005
R20336 vdd.n1297 vdd.n1296 9.3005
R20337 vdd.n1298 vdd.n1242 9.3005
R20338 vdd.n1300 vdd.n1299 9.3005
R20339 vdd.n1301 vdd.n1241 9.3005
R20340 vdd.n1306 vdd.n1302 9.3005
R20341 vdd.n1307 vdd.n1237 9.3005
R20342 vdd.n1309 vdd.n1308 9.3005
R20343 vdd.n1310 vdd.n1236 9.3005
R20344 vdd.n1312 vdd.n1311 9.3005
R20345 vdd.n1313 vdd.n1231 9.3005
R20346 vdd.n1315 vdd.n1314 9.3005
R20347 vdd.n1316 vdd.n1230 9.3005
R20348 vdd.n1318 vdd.n1317 9.3005
R20349 vdd.n1319 vdd.n1225 9.3005
R20350 vdd.n1321 vdd.n1320 9.3005
R20351 vdd.n1322 vdd.n1224 9.3005
R20352 vdd.n1324 vdd.n1323 9.3005
R20353 vdd.n1325 vdd.n1219 9.3005
R20354 vdd.n1327 vdd.n1326 9.3005
R20355 vdd.n1328 vdd.n1218 9.3005
R20356 vdd.n1330 vdd.n1329 9.3005
R20357 vdd.n1331 vdd.n1213 9.3005
R20358 vdd.n1333 vdd.n1332 9.3005
R20359 vdd.n1334 vdd.n1212 9.3005
R20360 vdd.n1336 vdd.n1335 9.3005
R20361 vdd.n1337 vdd.n1209 9.3005
R20362 vdd.n1343 vdd.n1342 9.3005
R20363 vdd.n1344 vdd.n1208 9.3005
R20364 vdd.n1346 vdd.n1345 9.3005
R20365 vdd.n1347 vdd.n1203 9.3005
R20366 vdd.n1349 vdd.n1348 9.3005
R20367 vdd.n1350 vdd.n1202 9.3005
R20368 vdd.n1352 vdd.n1351 9.3005
R20369 vdd.n1353 vdd.n1197 9.3005
R20370 vdd.n1355 vdd.n1354 9.3005
R20371 vdd.n1356 vdd.n1196 9.3005
R20372 vdd.n1358 vdd.n1357 9.3005
R20373 vdd.n1359 vdd.n1191 9.3005
R20374 vdd.n1361 vdd.n1360 9.3005
R20375 vdd.n1362 vdd.n1190 9.3005
R20376 vdd.n1364 vdd.n1363 9.3005
R20377 vdd.n1365 vdd.n1186 9.3005
R20378 vdd.n1367 vdd.n1366 9.3005
R20379 vdd.n1368 vdd.n1185 9.3005
R20380 vdd.n1370 vdd.n1369 9.3005
R20381 vdd.n1371 vdd.n1184 9.3005
R20382 vdd.n1377 vdd.n1376 9.3005
R20383 vdd.n1385 vdd.n1384 9.3005
R20384 vdd.n1386 vdd.n1140 9.3005
R20385 vdd.n1388 vdd.n1387 9.3005
R20386 vdd.n1130 vdd.n1129 9.3005
R20387 vdd.n1402 vdd.n1401 9.3005
R20388 vdd.n1403 vdd.n1128 9.3005
R20389 vdd.n1405 vdd.n1404 9.3005
R20390 vdd.n1119 vdd.n1118 9.3005
R20391 vdd.n1419 vdd.n1418 9.3005
R20392 vdd.n1420 vdd.n1117 9.3005
R20393 vdd.n1422 vdd.n1421 9.3005
R20394 vdd.n1108 vdd.n1107 9.3005
R20395 vdd.n1435 vdd.n1434 9.3005
R20396 vdd.n1436 vdd.n1106 9.3005
R20397 vdd.n1438 vdd.n1437 9.3005
R20398 vdd.n1096 vdd.n1095 9.3005
R20399 vdd.n1452 vdd.n1451 9.3005
R20400 vdd.n1142 vdd.n1141 9.3005
R20401 vdd.n1664 vdd.n1663 9.3005
R20402 vdd.n1659 vdd.n1658 9.3005
R20403 vdd.n1670 vdd.n1669 9.3005
R20404 vdd.n1672 vdd.n1671 9.3005
R20405 vdd.n1655 vdd.n1654 9.3005
R20406 vdd.n1678 vdd.n1677 9.3005
R20407 vdd.n1680 vdd.n1679 9.3005
R20408 vdd.n1652 vdd.n1649 9.3005
R20409 vdd.n1687 vdd.n1686 9.3005
R20410 vdd.n1719 vdd.n1718 9.3005
R20411 vdd.n1714 vdd.n1713 9.3005
R20412 vdd.n1725 vdd.n1724 9.3005
R20413 vdd.n1727 vdd.n1726 9.3005
R20414 vdd.n1710 vdd.n1709 9.3005
R20415 vdd.n1733 vdd.n1732 9.3005
R20416 vdd.n1735 vdd.n1734 9.3005
R20417 vdd.n1707 vdd.n1704 9.3005
R20418 vdd.n1742 vdd.n1741 9.3005
R20419 vdd.n1566 vdd.n1565 9.3005
R20420 vdd.n1561 vdd.n1560 9.3005
R20421 vdd.n1572 vdd.n1571 9.3005
R20422 vdd.n1574 vdd.n1573 9.3005
R20423 vdd.n1557 vdd.n1556 9.3005
R20424 vdd.n1580 vdd.n1579 9.3005
R20425 vdd.n1582 vdd.n1581 9.3005
R20426 vdd.n1554 vdd.n1551 9.3005
R20427 vdd.n1589 vdd.n1588 9.3005
R20428 vdd.n1621 vdd.n1620 9.3005
R20429 vdd.n1616 vdd.n1615 9.3005
R20430 vdd.n1627 vdd.n1626 9.3005
R20431 vdd.n1629 vdd.n1628 9.3005
R20432 vdd.n1612 vdd.n1611 9.3005
R20433 vdd.n1635 vdd.n1634 9.3005
R20434 vdd.n1637 vdd.n1636 9.3005
R20435 vdd.n1609 vdd.n1606 9.3005
R20436 vdd.n1644 vdd.n1643 9.3005
R20437 vdd.n1469 vdd.n1468 9.3005
R20438 vdd.n1464 vdd.n1463 9.3005
R20439 vdd.n1475 vdd.n1474 9.3005
R20440 vdd.n1477 vdd.n1476 9.3005
R20441 vdd.n1460 vdd.n1459 9.3005
R20442 vdd.n1483 vdd.n1482 9.3005
R20443 vdd.n1485 vdd.n1484 9.3005
R20444 vdd.n1457 vdd.n1454 9.3005
R20445 vdd.n1492 vdd.n1491 9.3005
R20446 vdd.n1524 vdd.n1523 9.3005
R20447 vdd.n1519 vdd.n1518 9.3005
R20448 vdd.n1530 vdd.n1529 9.3005
R20449 vdd.n1532 vdd.n1531 9.3005
R20450 vdd.n1515 vdd.n1514 9.3005
R20451 vdd.n1538 vdd.n1537 9.3005
R20452 vdd.n1540 vdd.n1539 9.3005
R20453 vdd.n1512 vdd.n1509 9.3005
R20454 vdd.n1547 vdd.n1546 9.3005
R20455 vdd.n1398 vdd.t92 9.18308
R20456 vdd.n3236 vdd.t35 9.18308
R20457 vdd.n1424 vdd.t39 8.95635
R20458 vdd.t37 vdd.n3277 8.95635
R20459 vdd.n300 vdd.n299 8.92171
R20460 vdd.n245 vdd.n244 8.92171
R20461 vdd.n202 vdd.n201 8.92171
R20462 vdd.n147 vdd.n146 8.92171
R20463 vdd.n105 vdd.n104 8.92171
R20464 vdd.n50 vdd.n49 8.92171
R20465 vdd.n1669 vdd.n1668 8.92171
R20466 vdd.n1724 vdd.n1723 8.92171
R20467 vdd.n1571 vdd.n1570 8.92171
R20468 vdd.n1626 vdd.n1625 8.92171
R20469 vdd.n1474 vdd.n1473 8.92171
R20470 vdd.n1529 vdd.n1528 8.92171
R20471 vdd.n223 vdd.n125 8.81535
R20472 vdd.n1647 vdd.n1549 8.81535
R20473 vdd.n1104 vdd.t95 8.72962
R20474 vdd.t65 vdd.n3286 8.72962
R20475 vdd.n1760 vdd.t23 8.50289
R20476 vdd.n3205 vdd.t108 8.50289
R20477 vdd.n28 vdd.n14 8.42249
R20478 vdd.n1776 vdd.t33 8.27616
R20479 vdd.t82 vdd.n636 8.27616
R20480 vdd.n3292 vdd.n3291 8.16225
R20481 vdd.n1747 vdd.n1746 8.16225
R20482 vdd.n296 vdd.n290 8.14595
R20483 vdd.n241 vdd.n235 8.14595
R20484 vdd.n198 vdd.n192 8.14595
R20485 vdd.n143 vdd.n137 8.14595
R20486 vdd.n101 vdd.n95 8.14595
R20487 vdd.n46 vdd.n40 8.14595
R20488 vdd.n1665 vdd.n1659 8.14595
R20489 vdd.n1720 vdd.n1714 8.14595
R20490 vdd.n1567 vdd.n1561 8.14595
R20491 vdd.n1622 vdd.n1616 8.14595
R20492 vdd.n1470 vdd.n1464 8.14595
R20493 vdd.n1525 vdd.n1519 8.14595
R20494 vdd.n2840 vdd.n820 8.11757
R20495 vdd.n2314 vdd.n2313 8.11757
R20496 vdd.t169 vdd.n1138 7.8227
R20497 vdd.t173 vdd.n363 7.8227
R20498 vdd.n2292 vdd.n1014 7.70933
R20499 vdd.n2298 vdd.n1014 7.70933
R20500 vdd.n2304 vdd.n1008 7.70933
R20501 vdd.n2304 vdd.n1001 7.70933
R20502 vdd.n2310 vdd.n1001 7.70933
R20503 vdd.n2310 vdd.n1004 7.70933
R20504 vdd.n2317 vdd.n989 7.70933
R20505 vdd.n2323 vdd.n989 7.70933
R20506 vdd.n2329 vdd.n983 7.70933
R20507 vdd.n2335 vdd.n979 7.70933
R20508 vdd.n2341 vdd.n973 7.70933
R20509 vdd.n2353 vdd.n960 7.70933
R20510 vdd.n2359 vdd.n954 7.70933
R20511 vdd.n2359 vdd.n947 7.70933
R20512 vdd.n2367 vdd.n947 7.70933
R20513 vdd.n2374 vdd.t15 7.70933
R20514 vdd.n2449 vdd.t15 7.70933
R20515 vdd.n2781 vdd.t157 7.70933
R20516 vdd.n2787 vdd.t157 7.70933
R20517 vdd.n2793 vdd.n868 7.70933
R20518 vdd.n2799 vdd.n868 7.70933
R20519 vdd.n2799 vdd.n871 7.70933
R20520 vdd.n2805 vdd.n864 7.70933
R20521 vdd.n2817 vdd.n851 7.70933
R20522 vdd.n2823 vdd.n845 7.70933
R20523 vdd.n2829 vdd.n841 7.70933
R20524 vdd.n2835 vdd.n828 7.70933
R20525 vdd.n2843 vdd.n828 7.70933
R20526 vdd.n2849 vdd.n822 7.70933
R20527 vdd.n2849 vdd.n814 7.70933
R20528 vdd.n2900 vdd.n814 7.70933
R20529 vdd.n2900 vdd.n817 7.70933
R20530 vdd.n2906 vdd.n774 7.70933
R20531 vdd.n2976 vdd.n774 7.70933
R20532 vdd.n295 vdd.n292 7.3702
R20533 vdd.n240 vdd.n237 7.3702
R20534 vdd.n197 vdd.n194 7.3702
R20535 vdd.n142 vdd.n139 7.3702
R20536 vdd.n100 vdd.n97 7.3702
R20537 vdd.n45 vdd.n42 7.3702
R20538 vdd.n1664 vdd.n1661 7.3702
R20539 vdd.n1719 vdd.n1716 7.3702
R20540 vdd.n1566 vdd.n1563 7.3702
R20541 vdd.n1621 vdd.n1618 7.3702
R20542 vdd.n1469 vdd.n1466 7.3702
R20543 vdd.n1524 vdd.n1521 7.3702
R20544 vdd.n1307 vdd.n1306 6.98232
R20545 vdd.n1956 vdd.n1955 6.98232
R20546 vdd.n547 vdd.n546 6.98232
R20547 vdd.n3060 vdd.n3059 6.98232
R20548 vdd.n1794 vdd.t126 6.91577
R20549 vdd.n3169 vdd.t88 6.91577
R20550 vdd.t53 vdd.n1075 6.68904
R20551 vdd.n3185 vdd.t55 6.68904
R20552 vdd.n1752 vdd.t104 6.46231
R20553 vdd.n3213 vdd.t63 6.46231
R20554 vdd.n3292 vdd.n321 6.32949
R20555 vdd.n1746 vdd.n1745 6.32949
R20556 vdd.t67 vdd.n1103 6.23558
R20557 vdd.t58 vdd.n332 6.23558
R20558 vdd.n1416 vdd.t90 6.00885
R20559 vdd.n2329 vdd.t18 6.00885
R20560 vdd.n2829 vdd.t11 6.00885
R20561 vdd.n3271 vdd.t61 6.00885
R20562 vdd.n1004 vdd.t219 5.89549
R20563 vdd.t187 vdd.n822 5.89549
R20564 vdd.n296 vdd.n295 5.81868
R20565 vdd.n241 vdd.n240 5.81868
R20566 vdd.n198 vdd.n197 5.81868
R20567 vdd.n143 vdd.n142 5.81868
R20568 vdd.n101 vdd.n100 5.81868
R20569 vdd.n46 vdd.n45 5.81868
R20570 vdd.n1665 vdd.n1664 5.81868
R20571 vdd.n1720 vdd.n1719 5.81868
R20572 vdd.n1567 vdd.n1566 5.81868
R20573 vdd.n1622 vdd.n1621 5.81868
R20574 vdd.n1470 vdd.n1469 5.81868
R20575 vdd.n1525 vdd.n1524 5.81868
R20576 vdd.t215 vdd.n1008 5.78212
R20577 vdd.n2073 vdd.t200 5.78212
R20578 vdd.n2698 vdd.t208 5.78212
R20579 vdd.n817 vdd.t204 5.78212
R20580 vdd.n2457 vdd.n2456 5.77611
R20581 vdd.n2200 vdd.n2070 5.77611
R20582 vdd.n2711 vdd.n2710 5.77611
R20583 vdd.n2915 vdd.n806 5.77611
R20584 vdd.n2981 vdd.n770 5.77611
R20585 vdd.n2621 vdd.n2561 5.77611
R20586 vdd.n2382 vdd.n938 5.77611
R20587 vdd.n2130 vdd.n2129 5.77611
R20588 vdd.n1376 vdd.n1150 5.62474
R20589 vdd.n2252 vdd.n2249 5.62474
R20590 vdd.n3250 vdd.n407 5.62474
R20591 vdd.n3015 vdd.n3012 5.62474
R20592 vdd.t153 vdd.n960 5.44203
R20593 vdd.n864 vdd.t8 5.44203
R20594 vdd.n1126 vdd.t90 5.32866
R20595 vdd.t61 vdd.n3270 5.32866
R20596 vdd.n1432 vdd.t67 5.10193
R20597 vdd.t162 vdd.n983 5.10193
R20598 vdd.n973 vdd.t149 5.10193
R20599 vdd.t17 vdd.n851 5.10193
R20600 vdd.n841 vdd.t2 5.10193
R20601 vdd.n3279 vdd.t58 5.10193
R20602 vdd.n299 vdd.n290 5.04292
R20603 vdd.n244 vdd.n235 5.04292
R20604 vdd.n201 vdd.n192 5.04292
R20605 vdd.n146 vdd.n137 5.04292
R20606 vdd.n104 vdd.n95 5.04292
R20607 vdd.n49 vdd.n40 5.04292
R20608 vdd.n1668 vdd.n1659 5.04292
R20609 vdd.n1723 vdd.n1714 5.04292
R20610 vdd.n1570 vdd.n1561 5.04292
R20611 vdd.n1625 vdd.n1616 5.04292
R20612 vdd.n1473 vdd.n1464 5.04292
R20613 vdd.n1528 vdd.n1519 5.04292
R20614 vdd.n1448 vdd.t104 4.8752
R20615 vdd.t3 vdd.t0 4.8752
R20616 vdd.t150 vdd.t262 4.8752
R20617 vdd.t147 vdd.t161 4.8752
R20618 vdd.t155 vdd.t10 4.8752
R20619 vdd.t63 vdd.n328 4.8752
R20620 vdd.n2458 vdd.n2457 4.83952
R20621 vdd.n2070 vdd.n2066 4.83952
R20622 vdd.n2712 vdd.n2711 4.83952
R20623 vdd.n806 vdd.n801 4.83952
R20624 vdd.n770 vdd.n765 4.83952
R20625 vdd.n2618 vdd.n2561 4.83952
R20626 vdd.n2385 vdd.n938 4.83952
R20627 vdd.n2129 vdd.n2128 4.83952
R20628 vdd.n1924 vdd.n1036 4.74817
R20629 vdd.n1919 vdd.n1037 4.74817
R20630 vdd.n1821 vdd.n1818 4.74817
R20631 vdd.n2233 vdd.n1822 4.74817
R20632 vdd.n2235 vdd.n1821 4.74817
R20633 vdd.n2234 vdd.n2233 4.74817
R20634 vdd.n664 vdd.n662 4.74817
R20635 vdd.n3130 vdd.n665 4.74817
R20636 vdd.n3133 vdd.n665 4.74817
R20637 vdd.n3134 vdd.n664 4.74817
R20638 vdd.n3022 vdd.n749 4.74817
R20639 vdd.n3018 vdd.n751 4.74817
R20640 vdd.n3021 vdd.n751 4.74817
R20641 vdd.n3026 vdd.n749 4.74817
R20642 vdd.n1920 vdd.n1036 4.74817
R20643 vdd.n1039 vdd.n1037 4.74817
R20644 vdd.n321 vdd.n320 4.7074
R20645 vdd.n223 vdd.n222 4.7074
R20646 vdd.n1745 vdd.n1744 4.7074
R20647 vdd.n1647 vdd.n1646 4.7074
R20648 vdd.n1768 vdd.t53 4.64847
R20649 vdd.n3194 vdd.t55 4.64847
R20650 vdd.n2335 vdd.t4 4.53511
R20651 vdd.n2823 vdd.t260 4.53511
R20652 vdd.n1069 vdd.t126 4.42174
R20653 vdd.t88 vdd.n635 4.42174
R20654 vdd.n2367 vdd.t258 4.30838
R20655 vdd.n2793 vdd.t256 4.30838
R20656 vdd.n300 vdd.n288 4.26717
R20657 vdd.n245 vdd.n233 4.26717
R20658 vdd.n202 vdd.n190 4.26717
R20659 vdd.n147 vdd.n135 4.26717
R20660 vdd.n105 vdd.n93 4.26717
R20661 vdd.n50 vdd.n38 4.26717
R20662 vdd.n1669 vdd.n1657 4.26717
R20663 vdd.n1724 vdd.n1712 4.26717
R20664 vdd.n1571 vdd.n1559 4.26717
R20665 vdd.n1626 vdd.n1614 4.26717
R20666 vdd.n1474 vdd.n1462 4.26717
R20667 vdd.n1529 vdd.n1517 4.26717
R20668 vdd.n321 vdd.n223 4.10845
R20669 vdd.n1745 vdd.n1647 4.10845
R20670 vdd.n277 vdd.t141 4.06363
R20671 vdd.n277 vdd.t52 4.06363
R20672 vdd.n275 vdd.t73 4.06363
R20673 vdd.n275 vdd.t140 4.06363
R20674 vdd.n273 vdd.t142 4.06363
R20675 vdd.n273 vdd.t72 4.06363
R20676 vdd.n271 vdd.t77 4.06363
R20677 vdd.n271 vdd.t79 4.06363
R20678 vdd.n269 vdd.t118 4.06363
R20679 vdd.n269 vdd.t44 4.06363
R20680 vdd.n267 vdd.t47 4.06363
R20681 vdd.n267 vdd.t97 4.06363
R20682 vdd.n265 vdd.t99 4.06363
R20683 vdd.n265 vdd.t123 4.06363
R20684 vdd.n179 vdd.t130 4.06363
R20685 vdd.n179 vdd.t36 4.06363
R20686 vdd.n177 vdd.t60 4.06363
R20687 vdd.n177 vdd.t129 4.06363
R20688 vdd.n175 vdd.t133 4.06363
R20689 vdd.n175 vdd.t59 4.06363
R20690 vdd.n173 vdd.t64 4.06363
R20691 vdd.n173 vdd.t66 4.06363
R20692 vdd.n171 vdd.t109 4.06363
R20693 vdd.n171 vdd.t146 4.06363
R20694 vdd.n169 vdd.t26 4.06363
R20695 vdd.n169 vdd.t80 4.06363
R20696 vdd.n167 vdd.t89 4.06363
R20697 vdd.n167 vdd.t111 4.06363
R20698 vdd.n82 vdd.t62 4.06363
R20699 vdd.n82 vdd.t125 4.06363
R20700 vdd.n80 vdd.t38 4.06363
R20701 vdd.n80 vdd.t85 4.06363
R20702 vdd.n78 vdd.t30 4.06363
R20703 vdd.n78 vdd.t69 4.06363
R20704 vdd.n76 vdd.t139 4.06363
R20705 vdd.n76 vdd.t115 4.06363
R20706 vdd.n74 vdd.t119 4.06363
R20707 vdd.n74 vdd.t76 4.06363
R20708 vdd.n72 vdd.t144 4.06363
R20709 vdd.n72 vdd.t56 4.06363
R20710 vdd.n70 vdd.t131 4.06363
R20711 vdd.n70 vdd.t83 4.06363
R20712 vdd.n1689 vdd.t49 4.06363
R20713 vdd.n1689 vdd.t136 4.06363
R20714 vdd.n1691 vdd.t135 4.06363
R20715 vdd.n1691 vdd.t117 4.06363
R20716 vdd.n1693 vdd.t94 4.06363
R20717 vdd.n1693 vdd.t46 4.06363
R20718 vdd.n1695 vdd.t145 4.06363
R20719 vdd.n1695 vdd.t116 4.06363
R20720 vdd.n1697 vdd.t112 4.06363
R20721 vdd.n1697 vdd.t71 4.06363
R20722 vdd.n1699 vdd.t70 4.06363
R20723 vdd.n1699 vdd.t113 4.06363
R20724 vdd.n1701 vdd.t100 4.06363
R20725 vdd.n1701 vdd.t101 4.06363
R20726 vdd.n1591 vdd.t34 4.06363
R20727 vdd.n1591 vdd.t127 4.06363
R20728 vdd.n1593 vdd.t120 4.06363
R20729 vdd.n1593 vdd.t107 4.06363
R20730 vdd.n1595 vdd.t78 4.06363
R20731 vdd.n1595 vdd.t24 4.06363
R20732 vdd.n1597 vdd.t134 4.06363
R20733 vdd.n1597 vdd.t105 4.06363
R20734 vdd.n1599 vdd.t102 4.06363
R20735 vdd.n1599 vdd.t57 4.06363
R20736 vdd.n1601 vdd.t51 4.06363
R20737 vdd.n1601 vdd.t103 4.06363
R20738 vdd.n1603 vdd.t93 4.06363
R20739 vdd.n1603 vdd.t91 4.06363
R20740 vdd.n1494 vdd.t81 4.06363
R20741 vdd.n1494 vdd.t132 4.06363
R20742 vdd.n1496 vdd.t54 4.06363
R20743 vdd.n1496 vdd.t114 4.06363
R20744 vdd.n1498 vdd.t75 4.06363
R20745 vdd.n1498 vdd.t121 4.06363
R20746 vdd.n1500 vdd.t96 4.06363
R20747 vdd.n1500 vdd.t138 4.06363
R20748 vdd.n1502 vdd.t68 4.06363
R20749 vdd.n1502 vdd.t28 4.06363
R20750 vdd.n1504 vdd.t86 4.06363
R20751 vdd.n1504 vdd.t40 4.06363
R20752 vdd.n1506 vdd.t128 4.06363
R20753 vdd.n1506 vdd.t143 4.06363
R20754 vdd.n26 vdd.t249 3.9605
R20755 vdd.n26 vdd.t247 3.9605
R20756 vdd.n23 vdd.t248 3.9605
R20757 vdd.n23 vdd.t253 3.9605
R20758 vdd.n21 vdd.t246 3.9605
R20759 vdd.n21 vdd.t244 3.9605
R20760 vdd.n20 vdd.t252 3.9605
R20761 vdd.n20 vdd.t242 3.9605
R20762 vdd.n15 vdd.t251 3.9605
R20763 vdd.n15 vdd.t255 3.9605
R20764 vdd.n16 vdd.t254 3.9605
R20765 vdd.n16 vdd.t240 3.9605
R20766 vdd.n18 vdd.t245 3.9605
R20767 vdd.n18 vdd.t250 3.9605
R20768 vdd.n25 vdd.t241 3.9605
R20769 vdd.n25 vdd.t243 3.9605
R20770 vdd.n7 vdd.t156 3.61217
R20771 vdd.n7 vdd.t261 3.61217
R20772 vdd.n8 vdd.t148 3.61217
R20773 vdd.n8 vdd.t9 3.61217
R20774 vdd.n10 vdd.t158 3.61217
R20775 vdd.n10 vdd.t257 3.61217
R20776 vdd.n12 vdd.t13 3.61217
R20777 vdd.n12 vdd.t160 3.61217
R20778 vdd.n5 vdd.t7 3.61217
R20779 vdd.n5 vdd.t152 3.61217
R20780 vdd.n3 vdd.t259 3.61217
R20781 vdd.n3 vdd.t16 3.61217
R20782 vdd.n1 vdd.t154 3.61217
R20783 vdd.n1 vdd.t263 3.61217
R20784 vdd.n0 vdd.t5 3.61217
R20785 vdd.n0 vdd.t1 3.61217
R20786 vdd.n1382 vdd.t169 3.51482
R20787 vdd.n3255 vdd.t173 3.51482
R20788 vdd.n304 vdd.n303 3.49141
R20789 vdd.n249 vdd.n248 3.49141
R20790 vdd.n206 vdd.n205 3.49141
R20791 vdd.n151 vdd.n150 3.49141
R20792 vdd.n109 vdd.n108 3.49141
R20793 vdd.n54 vdd.n53 3.49141
R20794 vdd.n1673 vdd.n1672 3.49141
R20795 vdd.n1728 vdd.n1727 3.49141
R20796 vdd.n1575 vdd.n1574 3.49141
R20797 vdd.n1630 vdd.n1629 3.49141
R20798 vdd.n1478 vdd.n1477 3.49141
R20799 vdd.n1533 vdd.n1532 3.49141
R20800 vdd.n2073 vdd.t258 3.40145
R20801 vdd.n2521 vdd.t6 3.40145
R20802 vdd.n2774 vdd.t159 3.40145
R20803 vdd.n2698 vdd.t256 3.40145
R20804 vdd.n2174 vdd.t4 3.17472
R20805 vdd.n2677 vdd.t260 3.17472
R20806 vdd.n1785 vdd.t33 3.06136
R20807 vdd.n3177 vdd.t82 3.06136
R20808 vdd.t23 vdd.n1081 2.83463
R20809 vdd.n624 vdd.t108 2.83463
R20810 vdd.n307 vdd.n286 2.71565
R20811 vdd.n252 vdd.n231 2.71565
R20812 vdd.n209 vdd.n188 2.71565
R20813 vdd.n154 vdd.n133 2.71565
R20814 vdd.n112 vdd.n91 2.71565
R20815 vdd.n57 vdd.n36 2.71565
R20816 vdd.n1676 vdd.n1655 2.71565
R20817 vdd.n1731 vdd.n1710 2.71565
R20818 vdd.n1578 vdd.n1557 2.71565
R20819 vdd.n1633 vdd.n1612 2.71565
R20820 vdd.n1481 vdd.n1460 2.71565
R20821 vdd.n1536 vdd.n1515 2.71565
R20822 vdd.n1449 vdd.t95 2.6079
R20823 vdd.n2323 vdd.t162 2.6079
R20824 vdd.n2347 vdd.t149 2.6079
R20825 vdd.n2811 vdd.t17 2.6079
R20826 vdd.n2835 vdd.t2 2.6079
R20827 vdd.n3287 vdd.t65 2.6079
R20828 vdd.n2841 vdd.n2840 2.49806
R20829 vdd.n2315 vdd.n2314 2.49806
R20830 vdd.n294 vdd.n293 2.4129
R20831 vdd.n239 vdd.n238 2.4129
R20832 vdd.n196 vdd.n195 2.4129
R20833 vdd.n141 vdd.n140 2.4129
R20834 vdd.n99 vdd.n98 2.4129
R20835 vdd.n44 vdd.n43 2.4129
R20836 vdd.n1663 vdd.n1662 2.4129
R20837 vdd.n1718 vdd.n1717 2.4129
R20838 vdd.n1565 vdd.n1564 2.4129
R20839 vdd.n1620 vdd.n1619 2.4129
R20840 vdd.n1468 vdd.n1467 2.4129
R20841 vdd.n1523 vdd.n1522 2.4129
R20842 vdd.t39 vdd.n1110 2.38117
R20843 vdd.n3278 vdd.t37 2.38117
R20844 vdd.n2232 vdd.n1821 2.27742
R20845 vdd.n2233 vdd.n2232 2.27742
R20846 vdd.n2942 vdd.n665 2.27742
R20847 vdd.n2942 vdd.n664 2.27742
R20848 vdd.n3010 vdd.n751 2.27742
R20849 vdd.n3010 vdd.n749 2.27742
R20850 vdd.n2255 vdd.n1036 2.27742
R20851 vdd.n2255 vdd.n1037 2.27742
R20852 vdd.n2347 vdd.t153 2.2678
R20853 vdd.n2811 vdd.t8 2.2678
R20854 vdd.n1407 vdd.t92 2.15444
R20855 vdd.n3269 vdd.t35 2.15444
R20856 vdd.t262 vdd.n954 2.04107
R20857 vdd.n871 vdd.t147 2.04107
R20858 vdd.n308 vdd.n284 1.93989
R20859 vdd.n253 vdd.n229 1.93989
R20860 vdd.n210 vdd.n186 1.93989
R20861 vdd.n155 vdd.n131 1.93989
R20862 vdd.n113 vdd.n89 1.93989
R20863 vdd.n58 vdd.n34 1.93989
R20864 vdd.n1677 vdd.n1653 1.93989
R20865 vdd.n1732 vdd.n1708 1.93989
R20866 vdd.n1579 vdd.n1555 1.93989
R20867 vdd.n1634 vdd.n1610 1.93989
R20868 vdd.n1482 vdd.n1458 1.93989
R20869 vdd.n1537 vdd.n1513 1.93989
R20870 vdd.n2298 vdd.t215 1.92771
R20871 vdd.n2374 vdd.t200 1.92771
R20872 vdd.n2787 vdd.t208 1.92771
R20873 vdd.n2906 vdd.t204 1.92771
R20874 vdd.n1399 vdd.t31 1.70098
R20875 vdd.n2174 vdd.t18 1.70098
R20876 vdd.n979 vdd.t3 1.70098
R20877 vdd.t10 vdd.n845 1.70098
R20878 vdd.n2677 vdd.t11 1.70098
R20879 vdd.n3263 vdd.t41 1.70098
R20880 vdd.n1415 vdd.t50 1.47425
R20881 vdd.n349 vdd.t84 1.47425
R20882 vdd.n1440 vdd.t27 1.24752
R20883 vdd.t180 vdd.n1044 1.24752
R20884 vdd.n659 vdd.t165 1.24752
R20885 vdd.t29 vdd.n3285 1.24752
R20886 vdd.n319 vdd.n279 1.16414
R20887 vdd.n312 vdd.n311 1.16414
R20888 vdd.n264 vdd.n224 1.16414
R20889 vdd.n257 vdd.n256 1.16414
R20890 vdd.n221 vdd.n181 1.16414
R20891 vdd.n214 vdd.n213 1.16414
R20892 vdd.n166 vdd.n126 1.16414
R20893 vdd.n159 vdd.n158 1.16414
R20894 vdd.n124 vdd.n84 1.16414
R20895 vdd.n117 vdd.n116 1.16414
R20896 vdd.n69 vdd.n29 1.16414
R20897 vdd.n62 vdd.n61 1.16414
R20898 vdd.n1688 vdd.n1648 1.16414
R20899 vdd.n1681 vdd.n1680 1.16414
R20900 vdd.n1743 vdd.n1703 1.16414
R20901 vdd.n1736 vdd.n1735 1.16414
R20902 vdd.n1590 vdd.n1550 1.16414
R20903 vdd.n1583 vdd.n1582 1.16414
R20904 vdd.n1645 vdd.n1605 1.16414
R20905 vdd.n1638 vdd.n1637 1.16414
R20906 vdd.n1493 vdd.n1453 1.16414
R20907 vdd.n1486 vdd.n1485 1.16414
R20908 vdd.n1548 vdd.n1508 1.16414
R20909 vdd.n1541 vdd.n1540 1.16414
R20910 vdd.n2341 vdd.t0 1.13415
R20911 vdd.n2817 vdd.t155 1.13415
R20912 vdd.n1092 vdd.t74 1.02079
R20913 vdd.t219 vdd.t163 1.02079
R20914 vdd.t14 vdd.t187 1.02079
R20915 vdd.t43 vdd.n613 1.02079
R20916 vdd.n1271 vdd.n1150 0.970197
R20917 vdd.n2253 vdd.n2252 0.970197
R20918 vdd.n599 vdd.n407 0.970197
R20919 vdd.n3017 vdd.n3015 0.970197
R20920 vdd.n1746 vdd.n28 0.852297
R20921 vdd vdd.n3292 0.844463
R20922 vdd.n1777 vdd.t106 0.794056
R20923 vdd.n2317 vdd.t163 0.794056
R20924 vdd.n2353 vdd.t150 0.794056
R20925 vdd.n2805 vdd.t161 0.794056
R20926 vdd.n2843 vdd.t14 0.794056
R20927 vdd.n3186 vdd.t25 0.794056
R20928 vdd.n1793 vdd.t19 0.567326
R20929 vdd.t21 vdd.n642 0.567326
R20930 vdd.n2243 vdd.n2242 0.482207
R20931 vdd.n3142 vdd.n3141 0.482207
R20932 vdd.n444 vdd.n443 0.482207
R20933 vdd.n3249 vdd.n3248 0.482207
R20934 vdd.n3148 vdd.n656 0.482207
R20935 vdd.n1807 vdd.n1038 0.482207
R20936 vdd.n1378 vdd.n1377 0.482207
R20937 vdd.n1184 vdd.n1141 0.482207
R20938 vdd.n4 vdd.n2 0.459552
R20939 vdd.n11 vdd.n9 0.459552
R20940 vdd.n317 vdd.n316 0.388379
R20941 vdd.n283 vdd.n281 0.388379
R20942 vdd.n262 vdd.n261 0.388379
R20943 vdd.n228 vdd.n226 0.388379
R20944 vdd.n219 vdd.n218 0.388379
R20945 vdd.n185 vdd.n183 0.388379
R20946 vdd.n164 vdd.n163 0.388379
R20947 vdd.n130 vdd.n128 0.388379
R20948 vdd.n122 vdd.n121 0.388379
R20949 vdd.n88 vdd.n86 0.388379
R20950 vdd.n67 vdd.n66 0.388379
R20951 vdd.n33 vdd.n31 0.388379
R20952 vdd.n1686 vdd.n1685 0.388379
R20953 vdd.n1652 vdd.n1650 0.388379
R20954 vdd.n1741 vdd.n1740 0.388379
R20955 vdd.n1707 vdd.n1705 0.388379
R20956 vdd.n1588 vdd.n1587 0.388379
R20957 vdd.n1554 vdd.n1552 0.388379
R20958 vdd.n1643 vdd.n1642 0.388379
R20959 vdd.n1609 vdd.n1607 0.388379
R20960 vdd.n1491 vdd.n1490 0.388379
R20961 vdd.n1457 vdd.n1455 0.388379
R20962 vdd.n1546 vdd.n1545 0.388379
R20963 vdd.n1512 vdd.n1510 0.388379
R20964 vdd.n19 vdd.n17 0.387128
R20965 vdd.n24 vdd.n22 0.387128
R20966 vdd.n6 vdd.n4 0.358259
R20967 vdd.n13 vdd.n11 0.358259
R20968 vdd.n268 vdd.n266 0.358259
R20969 vdd.n270 vdd.n268 0.358259
R20970 vdd.n272 vdd.n270 0.358259
R20971 vdd.n274 vdd.n272 0.358259
R20972 vdd.n276 vdd.n274 0.358259
R20973 vdd.n278 vdd.n276 0.358259
R20974 vdd.n320 vdd.n278 0.358259
R20975 vdd.n170 vdd.n168 0.358259
R20976 vdd.n172 vdd.n170 0.358259
R20977 vdd.n174 vdd.n172 0.358259
R20978 vdd.n176 vdd.n174 0.358259
R20979 vdd.n178 vdd.n176 0.358259
R20980 vdd.n180 vdd.n178 0.358259
R20981 vdd.n222 vdd.n180 0.358259
R20982 vdd.n73 vdd.n71 0.358259
R20983 vdd.n75 vdd.n73 0.358259
R20984 vdd.n77 vdd.n75 0.358259
R20985 vdd.n79 vdd.n77 0.358259
R20986 vdd.n81 vdd.n79 0.358259
R20987 vdd.n83 vdd.n81 0.358259
R20988 vdd.n125 vdd.n83 0.358259
R20989 vdd.n1744 vdd.n1702 0.358259
R20990 vdd.n1702 vdd.n1700 0.358259
R20991 vdd.n1700 vdd.n1698 0.358259
R20992 vdd.n1698 vdd.n1696 0.358259
R20993 vdd.n1696 vdd.n1694 0.358259
R20994 vdd.n1694 vdd.n1692 0.358259
R20995 vdd.n1692 vdd.n1690 0.358259
R20996 vdd.n1646 vdd.n1604 0.358259
R20997 vdd.n1604 vdd.n1602 0.358259
R20998 vdd.n1602 vdd.n1600 0.358259
R20999 vdd.n1600 vdd.n1598 0.358259
R21000 vdd.n1598 vdd.n1596 0.358259
R21001 vdd.n1596 vdd.n1594 0.358259
R21002 vdd.n1594 vdd.n1592 0.358259
R21003 vdd.n1549 vdd.n1507 0.358259
R21004 vdd.n1507 vdd.n1505 0.358259
R21005 vdd.n1505 vdd.n1503 0.358259
R21006 vdd.n1503 vdd.n1501 0.358259
R21007 vdd.n1501 vdd.n1499 0.358259
R21008 vdd.n1499 vdd.n1497 0.358259
R21009 vdd.n1497 vdd.n1495 0.358259
R21010 vdd.n14 vdd.n6 0.334552
R21011 vdd.n14 vdd.n13 0.334552
R21012 vdd.n27 vdd.n19 0.21707
R21013 vdd.n27 vdd.n24 0.21707
R21014 vdd.n318 vdd.n280 0.155672
R21015 vdd.n310 vdd.n280 0.155672
R21016 vdd.n310 vdd.n309 0.155672
R21017 vdd.n309 vdd.n285 0.155672
R21018 vdd.n302 vdd.n285 0.155672
R21019 vdd.n302 vdd.n301 0.155672
R21020 vdd.n301 vdd.n289 0.155672
R21021 vdd.n294 vdd.n289 0.155672
R21022 vdd.n263 vdd.n225 0.155672
R21023 vdd.n255 vdd.n225 0.155672
R21024 vdd.n255 vdd.n254 0.155672
R21025 vdd.n254 vdd.n230 0.155672
R21026 vdd.n247 vdd.n230 0.155672
R21027 vdd.n247 vdd.n246 0.155672
R21028 vdd.n246 vdd.n234 0.155672
R21029 vdd.n239 vdd.n234 0.155672
R21030 vdd.n220 vdd.n182 0.155672
R21031 vdd.n212 vdd.n182 0.155672
R21032 vdd.n212 vdd.n211 0.155672
R21033 vdd.n211 vdd.n187 0.155672
R21034 vdd.n204 vdd.n187 0.155672
R21035 vdd.n204 vdd.n203 0.155672
R21036 vdd.n203 vdd.n191 0.155672
R21037 vdd.n196 vdd.n191 0.155672
R21038 vdd.n165 vdd.n127 0.155672
R21039 vdd.n157 vdd.n127 0.155672
R21040 vdd.n157 vdd.n156 0.155672
R21041 vdd.n156 vdd.n132 0.155672
R21042 vdd.n149 vdd.n132 0.155672
R21043 vdd.n149 vdd.n148 0.155672
R21044 vdd.n148 vdd.n136 0.155672
R21045 vdd.n141 vdd.n136 0.155672
R21046 vdd.n123 vdd.n85 0.155672
R21047 vdd.n115 vdd.n85 0.155672
R21048 vdd.n115 vdd.n114 0.155672
R21049 vdd.n114 vdd.n90 0.155672
R21050 vdd.n107 vdd.n90 0.155672
R21051 vdd.n107 vdd.n106 0.155672
R21052 vdd.n106 vdd.n94 0.155672
R21053 vdd.n99 vdd.n94 0.155672
R21054 vdd.n68 vdd.n30 0.155672
R21055 vdd.n60 vdd.n30 0.155672
R21056 vdd.n60 vdd.n59 0.155672
R21057 vdd.n59 vdd.n35 0.155672
R21058 vdd.n52 vdd.n35 0.155672
R21059 vdd.n52 vdd.n51 0.155672
R21060 vdd.n51 vdd.n39 0.155672
R21061 vdd.n44 vdd.n39 0.155672
R21062 vdd.n1687 vdd.n1649 0.155672
R21063 vdd.n1679 vdd.n1649 0.155672
R21064 vdd.n1679 vdd.n1678 0.155672
R21065 vdd.n1678 vdd.n1654 0.155672
R21066 vdd.n1671 vdd.n1654 0.155672
R21067 vdd.n1671 vdd.n1670 0.155672
R21068 vdd.n1670 vdd.n1658 0.155672
R21069 vdd.n1663 vdd.n1658 0.155672
R21070 vdd.n1742 vdd.n1704 0.155672
R21071 vdd.n1734 vdd.n1704 0.155672
R21072 vdd.n1734 vdd.n1733 0.155672
R21073 vdd.n1733 vdd.n1709 0.155672
R21074 vdd.n1726 vdd.n1709 0.155672
R21075 vdd.n1726 vdd.n1725 0.155672
R21076 vdd.n1725 vdd.n1713 0.155672
R21077 vdd.n1718 vdd.n1713 0.155672
R21078 vdd.n1589 vdd.n1551 0.155672
R21079 vdd.n1581 vdd.n1551 0.155672
R21080 vdd.n1581 vdd.n1580 0.155672
R21081 vdd.n1580 vdd.n1556 0.155672
R21082 vdd.n1573 vdd.n1556 0.155672
R21083 vdd.n1573 vdd.n1572 0.155672
R21084 vdd.n1572 vdd.n1560 0.155672
R21085 vdd.n1565 vdd.n1560 0.155672
R21086 vdd.n1644 vdd.n1606 0.155672
R21087 vdd.n1636 vdd.n1606 0.155672
R21088 vdd.n1636 vdd.n1635 0.155672
R21089 vdd.n1635 vdd.n1611 0.155672
R21090 vdd.n1628 vdd.n1611 0.155672
R21091 vdd.n1628 vdd.n1627 0.155672
R21092 vdd.n1627 vdd.n1615 0.155672
R21093 vdd.n1620 vdd.n1615 0.155672
R21094 vdd.n1492 vdd.n1454 0.155672
R21095 vdd.n1484 vdd.n1454 0.155672
R21096 vdd.n1484 vdd.n1483 0.155672
R21097 vdd.n1483 vdd.n1459 0.155672
R21098 vdd.n1476 vdd.n1459 0.155672
R21099 vdd.n1476 vdd.n1475 0.155672
R21100 vdd.n1475 vdd.n1463 0.155672
R21101 vdd.n1468 vdd.n1463 0.155672
R21102 vdd.n1547 vdd.n1509 0.155672
R21103 vdd.n1539 vdd.n1509 0.155672
R21104 vdd.n1539 vdd.n1538 0.155672
R21105 vdd.n1538 vdd.n1514 0.155672
R21106 vdd.n1531 vdd.n1514 0.155672
R21107 vdd.n1531 vdd.n1530 0.155672
R21108 vdd.n1530 vdd.n1518 0.155672
R21109 vdd.n1523 vdd.n1518 0.155672
R21110 vdd.n2018 vdd.n1823 0.152939
R21111 vdd.n1829 vdd.n1823 0.152939
R21112 vdd.n1830 vdd.n1829 0.152939
R21113 vdd.n1831 vdd.n1830 0.152939
R21114 vdd.n1832 vdd.n1831 0.152939
R21115 vdd.n1836 vdd.n1832 0.152939
R21116 vdd.n1837 vdd.n1836 0.152939
R21117 vdd.n1838 vdd.n1837 0.152939
R21118 vdd.n1839 vdd.n1838 0.152939
R21119 vdd.n1843 vdd.n1839 0.152939
R21120 vdd.n1844 vdd.n1843 0.152939
R21121 vdd.n1845 vdd.n1844 0.152939
R21122 vdd.n1993 vdd.n1845 0.152939
R21123 vdd.n1993 vdd.n1992 0.152939
R21124 vdd.n1992 vdd.n1991 0.152939
R21125 vdd.n1991 vdd.n1851 0.152939
R21126 vdd.n1856 vdd.n1851 0.152939
R21127 vdd.n1857 vdd.n1856 0.152939
R21128 vdd.n1858 vdd.n1857 0.152939
R21129 vdd.n1862 vdd.n1858 0.152939
R21130 vdd.n1863 vdd.n1862 0.152939
R21131 vdd.n1864 vdd.n1863 0.152939
R21132 vdd.n1865 vdd.n1864 0.152939
R21133 vdd.n1869 vdd.n1865 0.152939
R21134 vdd.n1870 vdd.n1869 0.152939
R21135 vdd.n1871 vdd.n1870 0.152939
R21136 vdd.n1872 vdd.n1871 0.152939
R21137 vdd.n1876 vdd.n1872 0.152939
R21138 vdd.n1877 vdd.n1876 0.152939
R21139 vdd.n1878 vdd.n1877 0.152939
R21140 vdd.n1879 vdd.n1878 0.152939
R21141 vdd.n1883 vdd.n1879 0.152939
R21142 vdd.n1884 vdd.n1883 0.152939
R21143 vdd.n1885 vdd.n1884 0.152939
R21144 vdd.n1954 vdd.n1885 0.152939
R21145 vdd.n1954 vdd.n1953 0.152939
R21146 vdd.n1953 vdd.n1952 0.152939
R21147 vdd.n1952 vdd.n1891 0.152939
R21148 vdd.n1896 vdd.n1891 0.152939
R21149 vdd.n1897 vdd.n1896 0.152939
R21150 vdd.n1898 vdd.n1897 0.152939
R21151 vdd.n1902 vdd.n1898 0.152939
R21152 vdd.n1903 vdd.n1902 0.152939
R21153 vdd.n1904 vdd.n1903 0.152939
R21154 vdd.n1905 vdd.n1904 0.152939
R21155 vdd.n1909 vdd.n1905 0.152939
R21156 vdd.n1910 vdd.n1909 0.152939
R21157 vdd.n1911 vdd.n1910 0.152939
R21158 vdd.n1912 vdd.n1911 0.152939
R21159 vdd.n1913 vdd.n1912 0.152939
R21160 vdd.n1913 vdd.n1035 0.152939
R21161 vdd.n2242 vdd.n1817 0.152939
R21162 vdd.n1749 vdd.n1748 0.152939
R21163 vdd.n1749 vdd.n1084 0.152939
R21164 vdd.n1763 vdd.n1084 0.152939
R21165 vdd.n1764 vdd.n1763 0.152939
R21166 vdd.n1765 vdd.n1764 0.152939
R21167 vdd.n1765 vdd.n1072 0.152939
R21168 vdd.n1780 vdd.n1072 0.152939
R21169 vdd.n1781 vdd.n1780 0.152939
R21170 vdd.n1782 vdd.n1781 0.152939
R21171 vdd.n1782 vdd.n1061 0.152939
R21172 vdd.n1797 vdd.n1061 0.152939
R21173 vdd.n1798 vdd.n1797 0.152939
R21174 vdd.n1799 vdd.n1798 0.152939
R21175 vdd.n1799 vdd.n1049 0.152939
R21176 vdd.n1815 vdd.n1049 0.152939
R21177 vdd.n1816 vdd.n1815 0.152939
R21178 vdd.n2243 vdd.n1816 0.152939
R21179 vdd.n670 vdd.n667 0.152939
R21180 vdd.n671 vdd.n670 0.152939
R21181 vdd.n672 vdd.n671 0.152939
R21182 vdd.n673 vdd.n672 0.152939
R21183 vdd.n676 vdd.n673 0.152939
R21184 vdd.n677 vdd.n676 0.152939
R21185 vdd.n678 vdd.n677 0.152939
R21186 vdd.n679 vdd.n678 0.152939
R21187 vdd.n682 vdd.n679 0.152939
R21188 vdd.n683 vdd.n682 0.152939
R21189 vdd.n684 vdd.n683 0.152939
R21190 vdd.n685 vdd.n684 0.152939
R21191 vdd.n690 vdd.n685 0.152939
R21192 vdd.n691 vdd.n690 0.152939
R21193 vdd.n692 vdd.n691 0.152939
R21194 vdd.n693 vdd.n692 0.152939
R21195 vdd.n696 vdd.n693 0.152939
R21196 vdd.n697 vdd.n696 0.152939
R21197 vdd.n698 vdd.n697 0.152939
R21198 vdd.n699 vdd.n698 0.152939
R21199 vdd.n702 vdd.n699 0.152939
R21200 vdd.n703 vdd.n702 0.152939
R21201 vdd.n704 vdd.n703 0.152939
R21202 vdd.n705 vdd.n704 0.152939
R21203 vdd.n708 vdd.n705 0.152939
R21204 vdd.n709 vdd.n708 0.152939
R21205 vdd.n710 vdd.n709 0.152939
R21206 vdd.n711 vdd.n710 0.152939
R21207 vdd.n714 vdd.n711 0.152939
R21208 vdd.n715 vdd.n714 0.152939
R21209 vdd.n716 vdd.n715 0.152939
R21210 vdd.n717 vdd.n716 0.152939
R21211 vdd.n720 vdd.n717 0.152939
R21212 vdd.n721 vdd.n720 0.152939
R21213 vdd.n3058 vdd.n721 0.152939
R21214 vdd.n3058 vdd.n3057 0.152939
R21215 vdd.n3057 vdd.n3056 0.152939
R21216 vdd.n3056 vdd.n725 0.152939
R21217 vdd.n730 vdd.n725 0.152939
R21218 vdd.n731 vdd.n730 0.152939
R21219 vdd.n734 vdd.n731 0.152939
R21220 vdd.n735 vdd.n734 0.152939
R21221 vdd.n736 vdd.n735 0.152939
R21222 vdd.n737 vdd.n736 0.152939
R21223 vdd.n740 vdd.n737 0.152939
R21224 vdd.n741 vdd.n740 0.152939
R21225 vdd.n742 vdd.n741 0.152939
R21226 vdd.n743 vdd.n742 0.152939
R21227 vdd.n746 vdd.n743 0.152939
R21228 vdd.n747 vdd.n746 0.152939
R21229 vdd.n748 vdd.n747 0.152939
R21230 vdd.n3141 vdd.n661 0.152939
R21231 vdd.n3142 vdd.n651 0.152939
R21232 vdd.n3156 vdd.n651 0.152939
R21233 vdd.n3157 vdd.n3156 0.152939
R21234 vdd.n3158 vdd.n3157 0.152939
R21235 vdd.n3158 vdd.n639 0.152939
R21236 vdd.n3172 vdd.n639 0.152939
R21237 vdd.n3173 vdd.n3172 0.152939
R21238 vdd.n3174 vdd.n3173 0.152939
R21239 vdd.n3174 vdd.n627 0.152939
R21240 vdd.n3189 vdd.n627 0.152939
R21241 vdd.n3190 vdd.n3189 0.152939
R21242 vdd.n3191 vdd.n3190 0.152939
R21243 vdd.n3191 vdd.n616 0.152939
R21244 vdd.n3208 vdd.n616 0.152939
R21245 vdd.n3209 vdd.n3208 0.152939
R21246 vdd.n3210 vdd.n3209 0.152939
R21247 vdd.n3210 vdd.n322 0.152939
R21248 vdd.n3290 vdd.n323 0.152939
R21249 vdd.n334 vdd.n323 0.152939
R21250 vdd.n335 vdd.n334 0.152939
R21251 vdd.n336 vdd.n335 0.152939
R21252 vdd.n343 vdd.n336 0.152939
R21253 vdd.n344 vdd.n343 0.152939
R21254 vdd.n345 vdd.n344 0.152939
R21255 vdd.n346 vdd.n345 0.152939
R21256 vdd.n354 vdd.n346 0.152939
R21257 vdd.n355 vdd.n354 0.152939
R21258 vdd.n356 vdd.n355 0.152939
R21259 vdd.n357 vdd.n356 0.152939
R21260 vdd.n365 vdd.n357 0.152939
R21261 vdd.n366 vdd.n365 0.152939
R21262 vdd.n367 vdd.n366 0.152939
R21263 vdd.n368 vdd.n367 0.152939
R21264 vdd.n443 vdd.n368 0.152939
R21265 vdd.n444 vdd.n442 0.152939
R21266 vdd.n451 vdd.n442 0.152939
R21267 vdd.n452 vdd.n451 0.152939
R21268 vdd.n453 vdd.n452 0.152939
R21269 vdd.n453 vdd.n440 0.152939
R21270 vdd.n461 vdd.n440 0.152939
R21271 vdd.n462 vdd.n461 0.152939
R21272 vdd.n463 vdd.n462 0.152939
R21273 vdd.n463 vdd.n438 0.152939
R21274 vdd.n471 vdd.n438 0.152939
R21275 vdd.n472 vdd.n471 0.152939
R21276 vdd.n473 vdd.n472 0.152939
R21277 vdd.n473 vdd.n436 0.152939
R21278 vdd.n481 vdd.n436 0.152939
R21279 vdd.n482 vdd.n481 0.152939
R21280 vdd.n483 vdd.n482 0.152939
R21281 vdd.n483 vdd.n434 0.152939
R21282 vdd.n491 vdd.n434 0.152939
R21283 vdd.n492 vdd.n491 0.152939
R21284 vdd.n493 vdd.n492 0.152939
R21285 vdd.n493 vdd.n430 0.152939
R21286 vdd.n501 vdd.n430 0.152939
R21287 vdd.n502 vdd.n501 0.152939
R21288 vdd.n503 vdd.n502 0.152939
R21289 vdd.n503 vdd.n428 0.152939
R21290 vdd.n511 vdd.n428 0.152939
R21291 vdd.n512 vdd.n511 0.152939
R21292 vdd.n513 vdd.n512 0.152939
R21293 vdd.n513 vdd.n426 0.152939
R21294 vdd.n521 vdd.n426 0.152939
R21295 vdd.n522 vdd.n521 0.152939
R21296 vdd.n523 vdd.n522 0.152939
R21297 vdd.n523 vdd.n424 0.152939
R21298 vdd.n531 vdd.n424 0.152939
R21299 vdd.n532 vdd.n531 0.152939
R21300 vdd.n533 vdd.n532 0.152939
R21301 vdd.n533 vdd.n422 0.152939
R21302 vdd.n541 vdd.n422 0.152939
R21303 vdd.n542 vdd.n541 0.152939
R21304 vdd.n543 vdd.n542 0.152939
R21305 vdd.n543 vdd.n418 0.152939
R21306 vdd.n551 vdd.n418 0.152939
R21307 vdd.n552 vdd.n551 0.152939
R21308 vdd.n553 vdd.n552 0.152939
R21309 vdd.n553 vdd.n416 0.152939
R21310 vdd.n561 vdd.n416 0.152939
R21311 vdd.n562 vdd.n561 0.152939
R21312 vdd.n563 vdd.n562 0.152939
R21313 vdd.n563 vdd.n414 0.152939
R21314 vdd.n571 vdd.n414 0.152939
R21315 vdd.n572 vdd.n571 0.152939
R21316 vdd.n573 vdd.n572 0.152939
R21317 vdd.n573 vdd.n412 0.152939
R21318 vdd.n581 vdd.n412 0.152939
R21319 vdd.n582 vdd.n581 0.152939
R21320 vdd.n583 vdd.n582 0.152939
R21321 vdd.n583 vdd.n410 0.152939
R21322 vdd.n591 vdd.n410 0.152939
R21323 vdd.n592 vdd.n591 0.152939
R21324 vdd.n593 vdd.n592 0.152939
R21325 vdd.n593 vdd.n408 0.152939
R21326 vdd.n600 vdd.n408 0.152939
R21327 vdd.n3249 vdd.n600 0.152939
R21328 vdd.n3149 vdd.n3148 0.152939
R21329 vdd.n3150 vdd.n3149 0.152939
R21330 vdd.n3150 vdd.n645 0.152939
R21331 vdd.n3164 vdd.n645 0.152939
R21332 vdd.n3165 vdd.n3164 0.152939
R21333 vdd.n3166 vdd.n3165 0.152939
R21334 vdd.n3166 vdd.n632 0.152939
R21335 vdd.n3180 vdd.n632 0.152939
R21336 vdd.n3181 vdd.n3180 0.152939
R21337 vdd.n3182 vdd.n3181 0.152939
R21338 vdd.n3182 vdd.n621 0.152939
R21339 vdd.n3197 vdd.n621 0.152939
R21340 vdd.n3198 vdd.n3197 0.152939
R21341 vdd.n3199 vdd.n3198 0.152939
R21342 vdd.n3201 vdd.n3199 0.152939
R21343 vdd.n3201 vdd.n3200 0.152939
R21344 vdd.n3200 vdd.n611 0.152939
R21345 vdd.n611 vdd.n609 0.152939
R21346 vdd.n3219 vdd.n609 0.152939
R21347 vdd.n3220 vdd.n3219 0.152939
R21348 vdd.n3221 vdd.n3220 0.152939
R21349 vdd.n3221 vdd.n607 0.152939
R21350 vdd.n3226 vdd.n607 0.152939
R21351 vdd.n3227 vdd.n3226 0.152939
R21352 vdd.n3228 vdd.n3227 0.152939
R21353 vdd.n3228 vdd.n605 0.152939
R21354 vdd.n3233 vdd.n605 0.152939
R21355 vdd.n3234 vdd.n3233 0.152939
R21356 vdd.n3235 vdd.n3234 0.152939
R21357 vdd.n3235 vdd.n603 0.152939
R21358 vdd.n3241 vdd.n603 0.152939
R21359 vdd.n3242 vdd.n3241 0.152939
R21360 vdd.n3243 vdd.n3242 0.152939
R21361 vdd.n3243 vdd.n601 0.152939
R21362 vdd.n3248 vdd.n601 0.152939
R21363 vdd.n3011 vdd.n656 0.152939
R21364 vdd.n2254 vdd.n1038 0.152939
R21365 vdd.n1379 vdd.n1378 0.152939
R21366 vdd.n1379 vdd.n1135 0.152939
R21367 vdd.n1393 vdd.n1135 0.152939
R21368 vdd.n1394 vdd.n1393 0.152939
R21369 vdd.n1395 vdd.n1394 0.152939
R21370 vdd.n1395 vdd.n1123 0.152939
R21371 vdd.n1410 vdd.n1123 0.152939
R21372 vdd.n1411 vdd.n1410 0.152939
R21373 vdd.n1412 vdd.n1411 0.152939
R21374 vdd.n1412 vdd.n1113 0.152939
R21375 vdd.n1427 vdd.n1113 0.152939
R21376 vdd.n1428 vdd.n1427 0.152939
R21377 vdd.n1429 vdd.n1428 0.152939
R21378 vdd.n1429 vdd.n1100 0.152939
R21379 vdd.n1443 vdd.n1100 0.152939
R21380 vdd.n1444 vdd.n1443 0.152939
R21381 vdd.n1445 vdd.n1444 0.152939
R21382 vdd.n1445 vdd.n1089 0.152939
R21383 vdd.n1755 vdd.n1089 0.152939
R21384 vdd.n1756 vdd.n1755 0.152939
R21385 vdd.n1757 vdd.n1756 0.152939
R21386 vdd.n1757 vdd.n1078 0.152939
R21387 vdd.n1771 vdd.n1078 0.152939
R21388 vdd.n1772 vdd.n1771 0.152939
R21389 vdd.n1773 vdd.n1772 0.152939
R21390 vdd.n1773 vdd.n1066 0.152939
R21391 vdd.n1788 vdd.n1066 0.152939
R21392 vdd.n1789 vdd.n1788 0.152939
R21393 vdd.n1790 vdd.n1789 0.152939
R21394 vdd.n1790 vdd.n1056 0.152939
R21395 vdd.n1805 vdd.n1056 0.152939
R21396 vdd.n1806 vdd.n1805 0.152939
R21397 vdd.n1809 vdd.n1806 0.152939
R21398 vdd.n1809 vdd.n1808 0.152939
R21399 vdd.n1808 vdd.n1807 0.152939
R21400 vdd.n1369 vdd.n1184 0.152939
R21401 vdd.n1369 vdd.n1368 0.152939
R21402 vdd.n1368 vdd.n1367 0.152939
R21403 vdd.n1367 vdd.n1186 0.152939
R21404 vdd.n1363 vdd.n1186 0.152939
R21405 vdd.n1363 vdd.n1362 0.152939
R21406 vdd.n1362 vdd.n1361 0.152939
R21407 vdd.n1361 vdd.n1191 0.152939
R21408 vdd.n1357 vdd.n1191 0.152939
R21409 vdd.n1357 vdd.n1356 0.152939
R21410 vdd.n1356 vdd.n1355 0.152939
R21411 vdd.n1355 vdd.n1197 0.152939
R21412 vdd.n1351 vdd.n1197 0.152939
R21413 vdd.n1351 vdd.n1350 0.152939
R21414 vdd.n1350 vdd.n1349 0.152939
R21415 vdd.n1349 vdd.n1203 0.152939
R21416 vdd.n1345 vdd.n1203 0.152939
R21417 vdd.n1345 vdd.n1344 0.152939
R21418 vdd.n1344 vdd.n1343 0.152939
R21419 vdd.n1343 vdd.n1209 0.152939
R21420 vdd.n1335 vdd.n1209 0.152939
R21421 vdd.n1335 vdd.n1334 0.152939
R21422 vdd.n1334 vdd.n1333 0.152939
R21423 vdd.n1333 vdd.n1213 0.152939
R21424 vdd.n1329 vdd.n1213 0.152939
R21425 vdd.n1329 vdd.n1328 0.152939
R21426 vdd.n1328 vdd.n1327 0.152939
R21427 vdd.n1327 vdd.n1219 0.152939
R21428 vdd.n1323 vdd.n1219 0.152939
R21429 vdd.n1323 vdd.n1322 0.152939
R21430 vdd.n1322 vdd.n1321 0.152939
R21431 vdd.n1321 vdd.n1225 0.152939
R21432 vdd.n1317 vdd.n1225 0.152939
R21433 vdd.n1317 vdd.n1316 0.152939
R21434 vdd.n1316 vdd.n1315 0.152939
R21435 vdd.n1315 vdd.n1231 0.152939
R21436 vdd.n1311 vdd.n1231 0.152939
R21437 vdd.n1311 vdd.n1310 0.152939
R21438 vdd.n1310 vdd.n1309 0.152939
R21439 vdd.n1309 vdd.n1237 0.152939
R21440 vdd.n1302 vdd.n1237 0.152939
R21441 vdd.n1302 vdd.n1301 0.152939
R21442 vdd.n1301 vdd.n1300 0.152939
R21443 vdd.n1300 vdd.n1242 0.152939
R21444 vdd.n1296 vdd.n1242 0.152939
R21445 vdd.n1296 vdd.n1295 0.152939
R21446 vdd.n1295 vdd.n1294 0.152939
R21447 vdd.n1294 vdd.n1248 0.152939
R21448 vdd.n1290 vdd.n1248 0.152939
R21449 vdd.n1290 vdd.n1289 0.152939
R21450 vdd.n1289 vdd.n1288 0.152939
R21451 vdd.n1288 vdd.n1254 0.152939
R21452 vdd.n1284 vdd.n1254 0.152939
R21453 vdd.n1284 vdd.n1283 0.152939
R21454 vdd.n1283 vdd.n1282 0.152939
R21455 vdd.n1282 vdd.n1260 0.152939
R21456 vdd.n1278 vdd.n1260 0.152939
R21457 vdd.n1278 vdd.n1277 0.152939
R21458 vdd.n1277 vdd.n1276 0.152939
R21459 vdd.n1276 vdd.n1266 0.152939
R21460 vdd.n1272 vdd.n1266 0.152939
R21461 vdd.n1272 vdd.n1147 0.152939
R21462 vdd.n1377 vdd.n1147 0.152939
R21463 vdd.n1385 vdd.n1141 0.152939
R21464 vdd.n1386 vdd.n1385 0.152939
R21465 vdd.n1387 vdd.n1386 0.152939
R21466 vdd.n1387 vdd.n1129 0.152939
R21467 vdd.n1402 vdd.n1129 0.152939
R21468 vdd.n1403 vdd.n1402 0.152939
R21469 vdd.n1404 vdd.n1403 0.152939
R21470 vdd.n1404 vdd.n1118 0.152939
R21471 vdd.n1419 vdd.n1118 0.152939
R21472 vdd.n1420 vdd.n1419 0.152939
R21473 vdd.n1421 vdd.n1420 0.152939
R21474 vdd.n1421 vdd.n1107 0.152939
R21475 vdd.n1435 vdd.n1107 0.152939
R21476 vdd.n1436 vdd.n1435 0.152939
R21477 vdd.n1437 vdd.n1436 0.152939
R21478 vdd.n1437 vdd.n1095 0.152939
R21479 vdd.n1452 vdd.n1095 0.152939
R21480 vdd.n2232 vdd.n1817 0.110256
R21481 vdd.n2942 vdd.n661 0.110256
R21482 vdd.n3011 vdd.n3010 0.110256
R21483 vdd.n2255 vdd.n2254 0.110256
R21484 vdd.n1748 vdd.n1747 0.0695946
R21485 vdd.n3291 vdd.n322 0.0695946
R21486 vdd.n3291 vdd.n3290 0.0695946
R21487 vdd.n1747 vdd.n1452 0.0695946
R21488 vdd.n2232 vdd.n2018 0.0431829
R21489 vdd.n2255 vdd.n1035 0.0431829
R21490 vdd.n2942 vdd.n667 0.0431829
R21491 vdd.n3010 vdd.n748 0.0431829
R21492 vdd vdd.n28 0.00833333
R21493 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R21494 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R21495 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R21496 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R21497 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R21498 a_n2848_n452.n1 a_n2848_n452.t23 533.058
R21499 a_n2848_n452.n101 a_n2848_n452.t25 512.366
R21500 a_n2848_n452.n100 a_n2848_n452.t19 512.366
R21501 a_n2848_n452.n69 a_n2848_n452.t37 512.366
R21502 a_n2848_n452.n98 a_n2848_n452.t33 512.366
R21503 a_n2848_n452.n19 a_n2848_n452.t29 539.01
R21504 a_n2848_n452.n78 a_n2848_n452.t27 512.366
R21505 a_n2848_n452.n79 a_n2848_n452.t35 512.366
R21506 a_n2848_n452.n73 a_n2848_n452.t17 512.366
R21507 a_n2848_n452.n80 a_n2848_n452.t21 512.366
R21508 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R21509 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R21510 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R21511 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R21512 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R21513 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R21514 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R21515 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R21516 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R21517 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R21518 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R21519 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R21520 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R21521 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R21522 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R21523 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R21524 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R21525 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R21526 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R21527 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R21528 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R21529 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R21530 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R21531 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R21532 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R21533 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R21534 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R21535 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R21536 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R21537 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R21538 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R21539 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R21540 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R21541 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R21542 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R21543 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R21544 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R21545 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R21546 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R21547 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R21548 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R21549 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R21550 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R21551 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R21552 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R21553 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R21554 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R21555 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R21556 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R21557 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R21558 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R21559 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R21560 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R21561 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R21562 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R21563 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R21564 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R21565 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R21566 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R21567 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R21568 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R21569 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R21570 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R21571 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R21572 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R21573 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R21574 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R21575 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R21576 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R21577 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R21578 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R21579 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R21580 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R21581 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R21582 a_n2848_n452.n24 a_n2848_n452.t30 74.6477
R21583 a_n2848_n452.t16 a_n2848_n452.n27 74.6477
R21584 a_n2848_n452.n26 a_n2848_n452.t24 74.2899
R21585 a_n2848_n452.n25 a_n2848_n452.t32 74.2897
R21586 a_n2848_n452.n27 a_n2848_n452.n104 70.6783
R21587 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R21588 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R21589 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R21590 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R21591 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R21592 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R21593 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R21594 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R21595 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R21596 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R21597 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R21598 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R21599 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R21600 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R21601 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R21602 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R21603 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R21604 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R21605 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R21606 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R21607 a_n2848_n452.n47 a_n2848_n452.t15 533.058
R21608 a_n2848_n452.t31 a_n2848_n452.n37 533.058
R21609 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R21610 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R21611 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R21612 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R21613 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R21614 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R21615 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R21616 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R21617 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R21618 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R21619 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R21620 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R21621 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R21622 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R21623 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R21624 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R21625 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R21626 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R21627 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R21628 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R21629 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R21630 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R21631 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R21632 a_n2848_n452.n104 a_n2848_n452.t38 3.61217
R21633 a_n2848_n452.n104 a_n2848_n452.t34 3.61217
R21634 a_n2848_n452.n103 a_n2848_n452.t26 3.61217
R21635 a_n2848_n452.n103 a_n2848_n452.t20 3.61217
R21636 a_n2848_n452.n72 a_n2848_n452.t18 3.61217
R21637 a_n2848_n452.n72 a_n2848_n452.t22 3.61217
R21638 a_n2848_n452.n71 a_n2848_n452.t28 3.61217
R21639 a_n2848_n452.n71 a_n2848_n452.t36 3.61217
R21640 a_n2848_n452.n65 a_n2848_n452.t39 2.82907
R21641 a_n2848_n452.n65 a_n2848_n452.t42 2.82907
R21642 a_n2848_n452.n66 a_n2848_n452.t41 2.82907
R21643 a_n2848_n452.n66 a_n2848_n452.t13 2.82907
R21644 a_n2848_n452.n68 a_n2848_n452.t7 2.82907
R21645 a_n2848_n452.n68 a_n2848_n452.t10 2.82907
R21646 a_n2848_n452.n64 a_n2848_n452.t40 2.82907
R21647 a_n2848_n452.n64 a_n2848_n452.t1 2.82907
R21648 a_n2848_n452.n62 a_n2848_n452.t6 2.82907
R21649 a_n2848_n452.n62 a_n2848_n452.t2 2.82907
R21650 a_n2848_n452.n60 a_n2848_n452.t43 2.82907
R21651 a_n2848_n452.n60 a_n2848_n452.t45 2.82907
R21652 a_n2848_n452.n56 a_n2848_n452.t5 2.82907
R21653 a_n2848_n452.n56 a_n2848_n452.t8 2.82907
R21654 a_n2848_n452.n57 a_n2848_n452.t46 2.82907
R21655 a_n2848_n452.n57 a_n2848_n452.t11 2.82907
R21656 a_n2848_n452.n59 a_n2848_n452.t0 2.82907
R21657 a_n2848_n452.n59 a_n2848_n452.t12 2.82907
R21658 a_n2848_n452.n55 a_n2848_n452.t14 2.82907
R21659 a_n2848_n452.n55 a_n2848_n452.t3 2.82907
R21660 a_n2848_n452.n53 a_n2848_n452.t9 2.82907
R21661 a_n2848_n452.n53 a_n2848_n452.t47 2.82907
R21662 a_n2848_n452.n52 a_n2848_n452.t4 2.82907
R21663 a_n2848_n452.n52 a_n2848_n452.t44 2.82907
R21664 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R21665 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R21666 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R21667 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R21668 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R21669 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R21670 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R21671 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R21672 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R21673 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R21674 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R21675 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R21676 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R21677 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R21678 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R21679 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R21680 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R21681 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R21682 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R21683 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R21684 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R21685 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R21686 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R21687 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R21688 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R21689 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R21690 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R21691 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R21692 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R21693 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R21694 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R21695 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R21696 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R21697 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R21698 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R21699 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R21700 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R21701 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R21702 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R21703 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R21704 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R21705 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R21706 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R21707 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R21708 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R21709 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R21710 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R21711 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R21712 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R21713 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R21714 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R21715 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R21716 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R21717 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R21718 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R21719 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R21720 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R21721 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R21722 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R21723 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R21724 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R21725 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R21726 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R21727 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R21728 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R21729 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R21730 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R21731 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R21732 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R21733 plus.n76 plus.t11 250.337
R21734 plus.n15 plus.t14 250.337
R21735 plus.n124 plus.t1 243.97
R21736 plus.n120 plus.t24 231.093
R21737 plus.n59 plus.t20 231.093
R21738 plus.n124 plus.n123 223.454
R21739 plus.n126 plus.n125 223.454
R21740 plus.n77 plus.t5 187.445
R21741 plus.n74 plus.t22 187.445
R21742 plus.n72 plus.t21 187.445
R21743 plus.n89 plus.t16 187.445
R21744 plus.n95 plus.t17 187.445
R21745 plus.n68 plus.t13 187.445
R21746 plus.n66 plus.t15 187.445
R21747 plus.n107 plus.t10 187.445
R21748 plus.n113 plus.t26 187.445
R21749 plus.n62 plus.t28 187.445
R21750 plus.n1 plus.t23 187.445
R21751 plus.n52 plus.t6 187.445
R21752 plus.n46 plus.t12 187.445
R21753 plus.n5 plus.t8 187.445
R21754 plus.n7 plus.t7 187.445
R21755 plus.n34 plus.t19 187.445
R21756 plus.n28 plus.t18 187.445
R21757 plus.n11 plus.t27 187.445
R21758 plus.n13 plus.t25 187.445
R21759 plus.n16 plus.t9 187.445
R21760 plus.n121 plus.n120 161.3
R21761 plus.n119 plus.n61 161.3
R21762 plus.n118 plus.n117 161.3
R21763 plus.n116 plus.n115 161.3
R21764 plus.n114 plus.n63 161.3
R21765 plus.n112 plus.n111 161.3
R21766 plus.n110 plus.n64 161.3
R21767 plus.n109 plus.n108 161.3
R21768 plus.n106 plus.n65 161.3
R21769 plus.n105 plus.n104 161.3
R21770 plus.n103 plus.n102 161.3
R21771 plus.n101 plus.n67 161.3
R21772 plus.n100 plus.n99 161.3
R21773 plus.n98 plus.n97 161.3
R21774 plus.n96 plus.n69 161.3
R21775 plus.n94 plus.n93 161.3
R21776 plus.n92 plus.n70 161.3
R21777 plus.n91 plus.n90 161.3
R21778 plus.n88 plus.n71 161.3
R21779 plus.n87 plus.n86 161.3
R21780 plus.n85 plus.n84 161.3
R21781 plus.n83 plus.n73 161.3
R21782 plus.n82 plus.n81 161.3
R21783 plus.n80 plus.n79 161.3
R21784 plus.n78 plus.n75 161.3
R21785 plus.n17 plus.n14 161.3
R21786 plus.n19 plus.n18 161.3
R21787 plus.n21 plus.n20 161.3
R21788 plus.n22 plus.n12 161.3
R21789 plus.n24 plus.n23 161.3
R21790 plus.n26 plus.n25 161.3
R21791 plus.n27 plus.n10 161.3
R21792 plus.n30 plus.n29 161.3
R21793 plus.n31 plus.n9 161.3
R21794 plus.n33 plus.n32 161.3
R21795 plus.n35 plus.n8 161.3
R21796 plus.n37 plus.n36 161.3
R21797 plus.n39 plus.n38 161.3
R21798 plus.n40 plus.n6 161.3
R21799 plus.n42 plus.n41 161.3
R21800 plus.n44 plus.n43 161.3
R21801 plus.n45 plus.n4 161.3
R21802 plus.n48 plus.n47 161.3
R21803 plus.n49 plus.n3 161.3
R21804 plus.n51 plus.n50 161.3
R21805 plus.n53 plus.n2 161.3
R21806 plus.n55 plus.n54 161.3
R21807 plus.n57 plus.n56 161.3
R21808 plus.n58 plus.n0 161.3
R21809 plus.n60 plus.n59 161.3
R21810 plus.n88 plus.n87 56.5617
R21811 plus.n97 plus.n96 56.5617
R21812 plus.n106 plus.n105 56.5617
R21813 plus.n45 plus.n44 56.5617
R21814 plus.n36 plus.n35 56.5617
R21815 plus.n27 plus.n26 56.5617
R21816 plus.n79 plus.n78 56.5617
R21817 plus.n115 plus.n114 56.5617
R21818 plus.n54 plus.n53 56.5617
R21819 plus.n18 plus.n17 56.5617
R21820 plus.n119 plus.n118 50.2647
R21821 plus.n58 plus.n57 50.2647
R21822 plus.n84 plus.n83 46.3896
R21823 plus.n108 plus.n64 46.3896
R21824 plus.n47 plus.n3 46.3896
R21825 plus.n23 plus.n22 46.3896
R21826 plus.n76 plus.n75 43.1929
R21827 plus.n15 plus.n14 43.1929
R21828 plus.n94 plus.n70 42.5146
R21829 plus.n101 plus.n100 42.5146
R21830 plus.n40 plus.n39 42.5146
R21831 plus.n33 plus.n9 42.5146
R21832 plus.n77 plus.n76 40.6041
R21833 plus.n16 plus.n15 40.6041
R21834 plus.n90 plus.n70 38.6395
R21835 plus.n102 plus.n101 38.6395
R21836 plus.n41 plus.n40 38.6395
R21837 plus.n29 plus.n9 38.6395
R21838 plus.n122 plus.n121 35.2031
R21839 plus.n83 plus.n82 34.7644
R21840 plus.n112 plus.n64 34.7644
R21841 plus.n51 plus.n3 34.7644
R21842 plus.n22 plus.n21 34.7644
R21843 plus.n79 plus.n74 21.8872
R21844 plus.n114 plus.n113 21.8872
R21845 plus.n53 plus.n52 21.8872
R21846 plus.n18 plus.n13 21.8872
R21847 plus.n89 plus.n88 19.9199
R21848 plus.n105 plus.n66 19.9199
R21849 plus.n44 plus.n5 19.9199
R21850 plus.n28 plus.n27 19.9199
R21851 plus.n123 plus.t2 19.8005
R21852 plus.n123 plus.t4 19.8005
R21853 plus.n125 plus.t3 19.8005
R21854 plus.n125 plus.t0 19.8005
R21855 plus.n96 plus.n95 17.9525
R21856 plus.n97 plus.n68 17.9525
R21857 plus.n36 plus.n7 17.9525
R21858 plus.n35 plus.n34 17.9525
R21859 plus.n87 plus.n72 15.9852
R21860 plus.n107 plus.n106 15.9852
R21861 plus.n46 plus.n45 15.9852
R21862 plus.n26 plus.n11 15.9852
R21863 plus plus.n127 14.7359
R21864 plus.n78 plus.n77 14.0178
R21865 plus.n115 plus.n62 14.0178
R21866 plus.n54 plus.n1 14.0178
R21867 plus.n17 plus.n16 14.0178
R21868 plus.n122 plus.n60 11.9342
R21869 plus.n118 plus.n62 10.575
R21870 plus.n57 plus.n1 10.575
R21871 plus.n120 plus.n119 9.49444
R21872 plus.n59 plus.n58 9.49444
R21873 plus.n84 plus.n72 8.60764
R21874 plus.n108 plus.n107 8.60764
R21875 plus.n47 plus.n46 8.60764
R21876 plus.n23 plus.n11 8.60764
R21877 plus.n95 plus.n94 6.6403
R21878 plus.n100 plus.n68 6.6403
R21879 plus.n39 plus.n7 6.6403
R21880 plus.n34 plus.n33 6.6403
R21881 plus.n127 plus.n126 5.40567
R21882 plus.n90 plus.n89 4.67295
R21883 plus.n102 plus.n66 4.67295
R21884 plus.n41 plus.n5 4.67295
R21885 plus.n29 plus.n28 4.67295
R21886 plus.n82 plus.n74 2.7056
R21887 plus.n113 plus.n112 2.7056
R21888 plus.n52 plus.n51 2.7056
R21889 plus.n21 plus.n13 2.7056
R21890 plus.n127 plus.n122 1.188
R21891 plus.n126 plus.n124 0.716017
R21892 plus.n80 plus.n75 0.189894
R21893 plus.n81 plus.n80 0.189894
R21894 plus.n81 plus.n73 0.189894
R21895 plus.n85 plus.n73 0.189894
R21896 plus.n86 plus.n85 0.189894
R21897 plus.n86 plus.n71 0.189894
R21898 plus.n91 plus.n71 0.189894
R21899 plus.n92 plus.n91 0.189894
R21900 plus.n93 plus.n92 0.189894
R21901 plus.n93 plus.n69 0.189894
R21902 plus.n98 plus.n69 0.189894
R21903 plus.n99 plus.n98 0.189894
R21904 plus.n99 plus.n67 0.189894
R21905 plus.n103 plus.n67 0.189894
R21906 plus.n104 plus.n103 0.189894
R21907 plus.n104 plus.n65 0.189894
R21908 plus.n109 plus.n65 0.189894
R21909 plus.n110 plus.n109 0.189894
R21910 plus.n111 plus.n110 0.189894
R21911 plus.n111 plus.n63 0.189894
R21912 plus.n116 plus.n63 0.189894
R21913 plus.n117 plus.n116 0.189894
R21914 plus.n117 plus.n61 0.189894
R21915 plus.n121 plus.n61 0.189894
R21916 plus.n60 plus.n0 0.189894
R21917 plus.n56 plus.n0 0.189894
R21918 plus.n56 plus.n55 0.189894
R21919 plus.n55 plus.n2 0.189894
R21920 plus.n50 plus.n2 0.189894
R21921 plus.n50 plus.n49 0.189894
R21922 plus.n49 plus.n48 0.189894
R21923 plus.n48 plus.n4 0.189894
R21924 plus.n43 plus.n4 0.189894
R21925 plus.n43 plus.n42 0.189894
R21926 plus.n42 plus.n6 0.189894
R21927 plus.n38 plus.n6 0.189894
R21928 plus.n38 plus.n37 0.189894
R21929 plus.n37 plus.n8 0.189894
R21930 plus.n32 plus.n8 0.189894
R21931 plus.n32 plus.n31 0.189894
R21932 plus.n31 plus.n30 0.189894
R21933 plus.n30 plus.n10 0.189894
R21934 plus.n25 plus.n10 0.189894
R21935 plus.n25 plus.n24 0.189894
R21936 plus.n24 plus.n12 0.189894
R21937 plus.n20 plus.n12 0.189894
R21938 plus.n20 plus.n19 0.189894
R21939 plus.n19 plus.n14 0.189894
R21940 a_n3106_n452.n1 a_n3106_n452.t22 214.321
R21941 a_n3106_n452.n14 a_n3106_n452.t21 214.321
R21942 a_n3106_n452.n15 a_n3106_n452.t0 214.321
R21943 a_n3106_n452.n16 a_n3106_n452.t13 214.321
R21944 a_n3106_n452.n17 a_n3106_n452.t20 214.321
R21945 a_n3106_n452.n18 a_n3106_n452.t54 214.321
R21946 a_n3106_n452.n19 a_n3106_n452.t55 214.321
R21947 a_n3106_n452.n20 a_n3106_n452.t25 214.321
R21948 a_n3106_n452.n0 a_n3106_n452.t46 55.8337
R21949 a_n3106_n452.n2 a_n3106_n452.t23 55.8337
R21950 a_n3106_n452.n13 a_n3106_n452.t24 55.8337
R21951 a_n3106_n452.n47 a_n3106_n452.t33 55.8335
R21952 a_n3106_n452.n45 a_n3106_n452.t9 55.8335
R21953 a_n3106_n452.n34 a_n3106_n452.t5 55.8335
R21954 a_n3106_n452.n33 a_n3106_n452.t43 55.8335
R21955 a_n3106_n452.n22 a_n3106_n452.t37 55.8335
R21956 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R21957 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R21958 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R21959 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R21960 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R21961 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R21962 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R21963 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R21964 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R21965 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R21966 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R21967 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R21968 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R21969 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R21970 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R21971 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R21972 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R21973 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R21974 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R21975 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R21976 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R21977 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R21978 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R21979 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R21980 a_n3106_n452.n48 a_n3106_n452.t31 2.82907
R21981 a_n3106_n452.n48 a_n3106_n452.t29 2.82907
R21982 a_n3106_n452.n50 a_n3106_n452.t42 2.82907
R21983 a_n3106_n452.n50 a_n3106_n452.t47 2.82907
R21984 a_n3106_n452.n52 a_n3106_n452.t40 2.82907
R21985 a_n3106_n452.n52 a_n3106_n452.t44 2.82907
R21986 a_n3106_n452.n54 a_n3106_n452.t36 2.82907
R21987 a_n3106_n452.n54 a_n3106_n452.t41 2.82907
R21988 a_n3106_n452.n3 a_n3106_n452.t15 2.82907
R21989 a_n3106_n452.n3 a_n3106_n452.t17 2.82907
R21990 a_n3106_n452.n5 a_n3106_n452.t11 2.82907
R21991 a_n3106_n452.n5 a_n3106_n452.t19 2.82907
R21992 a_n3106_n452.n7 a_n3106_n452.t2 2.82907
R21993 a_n3106_n452.n7 a_n3106_n452.t8 2.82907
R21994 a_n3106_n452.n9 a_n3106_n452.t3 2.82907
R21995 a_n3106_n452.n9 a_n3106_n452.t18 2.82907
R21996 a_n3106_n452.n11 a_n3106_n452.t27 2.82907
R21997 a_n3106_n452.n11 a_n3106_n452.t7 2.82907
R21998 a_n3106_n452.n43 a_n3106_n452.t12 2.82907
R21999 a_n3106_n452.n43 a_n3106_n452.t6 2.82907
R22000 a_n3106_n452.n41 a_n3106_n452.t14 2.82907
R22001 a_n3106_n452.n41 a_n3106_n452.t28 2.82907
R22002 a_n3106_n452.n39 a_n3106_n452.t4 2.82907
R22003 a_n3106_n452.n39 a_n3106_n452.t1 2.82907
R22004 a_n3106_n452.n37 a_n3106_n452.t53 2.82907
R22005 a_n3106_n452.n37 a_n3106_n452.t16 2.82907
R22006 a_n3106_n452.n35 a_n3106_n452.t26 2.82907
R22007 a_n3106_n452.n35 a_n3106_n452.t10 2.82907
R22008 a_n3106_n452.n31 a_n3106_n452.t32 2.82907
R22009 a_n3106_n452.n31 a_n3106_n452.t48 2.82907
R22010 a_n3106_n452.n29 a_n3106_n452.t39 2.82907
R22011 a_n3106_n452.n29 a_n3106_n452.t30 2.82907
R22012 a_n3106_n452.n27 a_n3106_n452.t50 2.82907
R22013 a_n3106_n452.n27 a_n3106_n452.t38 2.82907
R22014 a_n3106_n452.n25 a_n3106_n452.t45 2.82907
R22015 a_n3106_n452.n25 a_n3106_n452.t49 2.82907
R22016 a_n3106_n452.n23 a_n3106_n452.t34 2.82907
R22017 a_n3106_n452.n23 a_n3106_n452.t51 2.82907
R22018 a_n3106_n452.t52 a_n3106_n452.n57 2.82907
R22019 a_n3106_n452.n57 a_n3106_n452.t35 2.82907
R22020 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R22021 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R22022 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R22023 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R22024 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R22025 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R22026 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R22027 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R22028 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R22029 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R22030 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R22031 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R22032 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R22033 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R22034 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R22035 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R22036 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R22037 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R22038 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R22039 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R22040 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R22041 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R22042 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R22043 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R22044 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R22045 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R22046 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R22047 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R22048 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R22049 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R22050 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R22051 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R22052 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R22053 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R22054 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R22055 output.n41 output.n15 289.615
R22056 output.n72 output.n46 289.615
R22057 output.n104 output.n78 289.615
R22058 output.n136 output.n110 289.615
R22059 output.n77 output.n45 197.26
R22060 output.n77 output.n76 196.298
R22061 output.n109 output.n108 196.298
R22062 output.n141 output.n140 196.298
R22063 output.n42 output.n41 185
R22064 output.n40 output.n39 185
R22065 output.n19 output.n18 185
R22066 output.n34 output.n33 185
R22067 output.n32 output.n31 185
R22068 output.n23 output.n22 185
R22069 output.n26 output.n25 185
R22070 output.n73 output.n72 185
R22071 output.n71 output.n70 185
R22072 output.n50 output.n49 185
R22073 output.n65 output.n64 185
R22074 output.n63 output.n62 185
R22075 output.n54 output.n53 185
R22076 output.n57 output.n56 185
R22077 output.n105 output.n104 185
R22078 output.n103 output.n102 185
R22079 output.n82 output.n81 185
R22080 output.n97 output.n96 185
R22081 output.n95 output.n94 185
R22082 output.n86 output.n85 185
R22083 output.n89 output.n88 185
R22084 output.n137 output.n136 185
R22085 output.n135 output.n134 185
R22086 output.n114 output.n113 185
R22087 output.n129 output.n128 185
R22088 output.n127 output.n126 185
R22089 output.n118 output.n117 185
R22090 output.n121 output.n120 185
R22091 output.t18 output.n24 147.661
R22092 output.t1 output.n55 147.661
R22093 output.t19 output.n87 147.661
R22094 output.t0 output.n119 147.661
R22095 output.n41 output.n40 104.615
R22096 output.n40 output.n18 104.615
R22097 output.n33 output.n18 104.615
R22098 output.n33 output.n32 104.615
R22099 output.n32 output.n22 104.615
R22100 output.n25 output.n22 104.615
R22101 output.n72 output.n71 104.615
R22102 output.n71 output.n49 104.615
R22103 output.n64 output.n49 104.615
R22104 output.n64 output.n63 104.615
R22105 output.n63 output.n53 104.615
R22106 output.n56 output.n53 104.615
R22107 output.n104 output.n103 104.615
R22108 output.n103 output.n81 104.615
R22109 output.n96 output.n81 104.615
R22110 output.n96 output.n95 104.615
R22111 output.n95 output.n85 104.615
R22112 output.n88 output.n85 104.615
R22113 output.n136 output.n135 104.615
R22114 output.n135 output.n113 104.615
R22115 output.n128 output.n113 104.615
R22116 output.n128 output.n127 104.615
R22117 output.n127 output.n117 104.615
R22118 output.n120 output.n117 104.615
R22119 output.n1 output.t15 77.056
R22120 output.n14 output.t16 76.6694
R22121 output.n1 output.n0 72.7095
R22122 output.n3 output.n2 72.7095
R22123 output.n5 output.n4 72.7095
R22124 output.n7 output.n6 72.7095
R22125 output.n9 output.n8 72.7095
R22126 output.n11 output.n10 72.7095
R22127 output.n13 output.n12 72.7095
R22128 output.n25 output.t18 52.3082
R22129 output.n56 output.t1 52.3082
R22130 output.n88 output.t19 52.3082
R22131 output.n120 output.t0 52.3082
R22132 output.n26 output.n24 15.6674
R22133 output.n57 output.n55 15.6674
R22134 output.n89 output.n87 15.6674
R22135 output.n121 output.n119 15.6674
R22136 output.n27 output.n23 12.8005
R22137 output.n58 output.n54 12.8005
R22138 output.n90 output.n86 12.8005
R22139 output.n122 output.n118 12.8005
R22140 output.n31 output.n30 12.0247
R22141 output.n62 output.n61 12.0247
R22142 output.n94 output.n93 12.0247
R22143 output.n126 output.n125 12.0247
R22144 output.n34 output.n21 11.249
R22145 output.n65 output.n52 11.249
R22146 output.n97 output.n84 11.249
R22147 output.n129 output.n116 11.249
R22148 output.n35 output.n19 10.4732
R22149 output.n66 output.n50 10.4732
R22150 output.n98 output.n82 10.4732
R22151 output.n130 output.n114 10.4732
R22152 output.n39 output.n38 9.69747
R22153 output.n70 output.n69 9.69747
R22154 output.n102 output.n101 9.69747
R22155 output.n134 output.n133 9.69747
R22156 output.n45 output.n44 9.45567
R22157 output.n76 output.n75 9.45567
R22158 output.n108 output.n107 9.45567
R22159 output.n140 output.n139 9.45567
R22160 output.n44 output.n43 9.3005
R22161 output.n17 output.n16 9.3005
R22162 output.n38 output.n37 9.3005
R22163 output.n36 output.n35 9.3005
R22164 output.n21 output.n20 9.3005
R22165 output.n30 output.n29 9.3005
R22166 output.n28 output.n27 9.3005
R22167 output.n75 output.n74 9.3005
R22168 output.n48 output.n47 9.3005
R22169 output.n69 output.n68 9.3005
R22170 output.n67 output.n66 9.3005
R22171 output.n52 output.n51 9.3005
R22172 output.n61 output.n60 9.3005
R22173 output.n59 output.n58 9.3005
R22174 output.n107 output.n106 9.3005
R22175 output.n80 output.n79 9.3005
R22176 output.n101 output.n100 9.3005
R22177 output.n99 output.n98 9.3005
R22178 output.n84 output.n83 9.3005
R22179 output.n93 output.n92 9.3005
R22180 output.n91 output.n90 9.3005
R22181 output.n139 output.n138 9.3005
R22182 output.n112 output.n111 9.3005
R22183 output.n133 output.n132 9.3005
R22184 output.n131 output.n130 9.3005
R22185 output.n116 output.n115 9.3005
R22186 output.n125 output.n124 9.3005
R22187 output.n123 output.n122 9.3005
R22188 output.n42 output.n17 8.92171
R22189 output.n73 output.n48 8.92171
R22190 output.n105 output.n80 8.92171
R22191 output.n137 output.n112 8.92171
R22192 output output.n141 8.15037
R22193 output.n43 output.n15 8.14595
R22194 output.n74 output.n46 8.14595
R22195 output.n106 output.n78 8.14595
R22196 output.n138 output.n110 8.14595
R22197 output.n45 output.n15 5.81868
R22198 output.n76 output.n46 5.81868
R22199 output.n108 output.n78 5.81868
R22200 output.n140 output.n110 5.81868
R22201 output.n43 output.n42 5.04292
R22202 output.n74 output.n73 5.04292
R22203 output.n106 output.n105 5.04292
R22204 output.n138 output.n137 5.04292
R22205 output.n28 output.n24 4.38594
R22206 output.n59 output.n55 4.38594
R22207 output.n91 output.n87 4.38594
R22208 output.n123 output.n119 4.38594
R22209 output.n39 output.n17 4.26717
R22210 output.n70 output.n48 4.26717
R22211 output.n102 output.n80 4.26717
R22212 output.n134 output.n112 4.26717
R22213 output.n0 output.t4 3.9605
R22214 output.n0 output.t9 3.9605
R22215 output.n2 output.t13 3.9605
R22216 output.n2 output.t5 3.9605
R22217 output.n4 output.t8 3.9605
R22218 output.n4 output.t6 3.9605
R22219 output.n6 output.t12 3.9605
R22220 output.n6 output.t14 3.9605
R22221 output.n8 output.t17 3.9605
R22222 output.n8 output.t10 3.9605
R22223 output.n10 output.t11 3.9605
R22224 output.n10 output.t2 3.9605
R22225 output.n12 output.t3 3.9605
R22226 output.n12 output.t7 3.9605
R22227 output.n38 output.n19 3.49141
R22228 output.n69 output.n50 3.49141
R22229 output.n101 output.n82 3.49141
R22230 output.n133 output.n114 3.49141
R22231 output.n35 output.n34 2.71565
R22232 output.n66 output.n65 2.71565
R22233 output.n98 output.n97 2.71565
R22234 output.n130 output.n129 2.71565
R22235 output.n31 output.n21 1.93989
R22236 output.n62 output.n52 1.93989
R22237 output.n94 output.n84 1.93989
R22238 output.n126 output.n116 1.93989
R22239 output.n30 output.n23 1.16414
R22240 output.n61 output.n54 1.16414
R22241 output.n93 output.n86 1.16414
R22242 output.n125 output.n118 1.16414
R22243 output.n141 output.n109 0.962709
R22244 output.n109 output.n77 0.962709
R22245 output.n27 output.n26 0.388379
R22246 output.n58 output.n57 0.388379
R22247 output.n90 output.n89 0.388379
R22248 output.n122 output.n121 0.388379
R22249 output.n14 output.n13 0.387128
R22250 output.n13 output.n11 0.387128
R22251 output.n11 output.n9 0.387128
R22252 output.n9 output.n7 0.387128
R22253 output.n7 output.n5 0.387128
R22254 output.n5 output.n3 0.387128
R22255 output.n3 output.n1 0.387128
R22256 output.n44 output.n16 0.155672
R22257 output.n37 output.n16 0.155672
R22258 output.n37 output.n36 0.155672
R22259 output.n36 output.n20 0.155672
R22260 output.n29 output.n20 0.155672
R22261 output.n29 output.n28 0.155672
R22262 output.n75 output.n47 0.155672
R22263 output.n68 output.n47 0.155672
R22264 output.n68 output.n67 0.155672
R22265 output.n67 output.n51 0.155672
R22266 output.n60 output.n51 0.155672
R22267 output.n60 output.n59 0.155672
R22268 output.n107 output.n79 0.155672
R22269 output.n100 output.n79 0.155672
R22270 output.n100 output.n99 0.155672
R22271 output.n99 output.n83 0.155672
R22272 output.n92 output.n83 0.155672
R22273 output.n92 output.n91 0.155672
R22274 output.n139 output.n111 0.155672
R22275 output.n132 output.n111 0.155672
R22276 output.n132 output.n131 0.155672
R22277 output.n131 output.n115 0.155672
R22278 output.n124 output.n115 0.155672
R22279 output.n124 output.n123 0.155672
R22280 output output.n14 0.126227
R22281 minus.n76 minus.t28 250.337
R22282 minus.n15 minus.t20 250.337
R22283 minus.n126 minus.t1 243.255
R22284 minus.n120 minus.t8 231.093
R22285 minus.n59 minus.t10 231.093
R22286 minus.n125 minus.n123 224.169
R22287 minus.n125 minus.n124 223.454
R22288 minus.n62 minus.t12 187.445
R22289 minus.n113 minus.t18 187.445
R22290 minus.n107 minus.t25 187.445
R22291 minus.n66 minus.t22 187.445
R22292 minus.n68 minus.t19 187.445
R22293 minus.n95 minus.t7 187.445
R22294 minus.n89 minus.t6 187.445
R22295 minus.n72 minus.t16 187.445
R22296 minus.n74 minus.t15 187.445
R22297 minus.n77 minus.t23 187.445
R22298 minus.n16 minus.t14 187.445
R22299 minus.n13 minus.t9 187.445
R22300 minus.n11 minus.t5 187.445
R22301 minus.n28 minus.t26 187.445
R22302 minus.n34 minus.t27 187.445
R22303 minus.n7 minus.t21 187.445
R22304 minus.n5 minus.t24 187.445
R22305 minus.n46 minus.t17 187.445
R22306 minus.n52 minus.t11 187.445
R22307 minus.n1 minus.t13 187.445
R22308 minus.n78 minus.n75 161.3
R22309 minus.n80 minus.n79 161.3
R22310 minus.n82 minus.n81 161.3
R22311 minus.n83 minus.n73 161.3
R22312 minus.n85 minus.n84 161.3
R22313 minus.n87 minus.n86 161.3
R22314 minus.n88 minus.n71 161.3
R22315 minus.n91 minus.n90 161.3
R22316 minus.n92 minus.n70 161.3
R22317 minus.n94 minus.n93 161.3
R22318 minus.n96 minus.n69 161.3
R22319 minus.n98 minus.n97 161.3
R22320 minus.n100 minus.n99 161.3
R22321 minus.n101 minus.n67 161.3
R22322 minus.n103 minus.n102 161.3
R22323 minus.n105 minus.n104 161.3
R22324 minus.n106 minus.n65 161.3
R22325 minus.n109 minus.n108 161.3
R22326 minus.n110 minus.n64 161.3
R22327 minus.n112 minus.n111 161.3
R22328 minus.n114 minus.n63 161.3
R22329 minus.n116 minus.n115 161.3
R22330 minus.n118 minus.n117 161.3
R22331 minus.n119 minus.n61 161.3
R22332 minus.n121 minus.n120 161.3
R22333 minus.n60 minus.n59 161.3
R22334 minus.n58 minus.n0 161.3
R22335 minus.n57 minus.n56 161.3
R22336 minus.n55 minus.n54 161.3
R22337 minus.n53 minus.n2 161.3
R22338 minus.n51 minus.n50 161.3
R22339 minus.n49 minus.n3 161.3
R22340 minus.n48 minus.n47 161.3
R22341 minus.n45 minus.n4 161.3
R22342 minus.n44 minus.n43 161.3
R22343 minus.n42 minus.n41 161.3
R22344 minus.n40 minus.n6 161.3
R22345 minus.n39 minus.n38 161.3
R22346 minus.n37 minus.n36 161.3
R22347 minus.n35 minus.n8 161.3
R22348 minus.n33 minus.n32 161.3
R22349 minus.n31 minus.n9 161.3
R22350 minus.n30 minus.n29 161.3
R22351 minus.n27 minus.n10 161.3
R22352 minus.n26 minus.n25 161.3
R22353 minus.n24 minus.n23 161.3
R22354 minus.n22 minus.n12 161.3
R22355 minus.n21 minus.n20 161.3
R22356 minus.n19 minus.n18 161.3
R22357 minus.n17 minus.n14 161.3
R22358 minus.n106 minus.n105 56.5617
R22359 minus.n97 minus.n96 56.5617
R22360 minus.n88 minus.n87 56.5617
R22361 minus.n27 minus.n26 56.5617
R22362 minus.n36 minus.n35 56.5617
R22363 minus.n45 minus.n44 56.5617
R22364 minus.n115 minus.n114 56.5617
R22365 minus.n79 minus.n78 56.5617
R22366 minus.n18 minus.n17 56.5617
R22367 minus.n54 minus.n53 56.5617
R22368 minus.n119 minus.n118 50.2647
R22369 minus.n58 minus.n57 50.2647
R22370 minus.n108 minus.n64 46.3896
R22371 minus.n84 minus.n83 46.3896
R22372 minus.n23 minus.n22 46.3896
R22373 minus.n47 minus.n3 46.3896
R22374 minus.n76 minus.n75 43.1929
R22375 minus.n15 minus.n14 43.1929
R22376 minus.n101 minus.n100 42.5146
R22377 minus.n94 minus.n70 42.5146
R22378 minus.n33 minus.n9 42.5146
R22379 minus.n40 minus.n39 42.5146
R22380 minus.n77 minus.n76 40.6041
R22381 minus.n16 minus.n15 40.6041
R22382 minus.n102 minus.n101 38.6395
R22383 minus.n90 minus.n70 38.6395
R22384 minus.n29 minus.n9 38.6395
R22385 minus.n41 minus.n40 38.6395
R22386 minus.n122 minus.n121 35.4191
R22387 minus.n112 minus.n64 34.7644
R22388 minus.n83 minus.n82 34.7644
R22389 minus.n22 minus.n21 34.7644
R22390 minus.n51 minus.n3 34.7644
R22391 minus.n114 minus.n113 21.8872
R22392 minus.n79 minus.n74 21.8872
R22393 minus.n18 minus.n13 21.8872
R22394 minus.n53 minus.n52 21.8872
R22395 minus.n105 minus.n66 19.9199
R22396 minus.n89 minus.n88 19.9199
R22397 minus.n28 minus.n27 19.9199
R22398 minus.n44 minus.n5 19.9199
R22399 minus.n124 minus.t0 19.8005
R22400 minus.n124 minus.t2 19.8005
R22401 minus.n123 minus.t4 19.8005
R22402 minus.n123 minus.t3 19.8005
R22403 minus.n97 minus.n68 17.9525
R22404 minus.n96 minus.n95 17.9525
R22405 minus.n35 minus.n34 17.9525
R22406 minus.n36 minus.n7 17.9525
R22407 minus.n107 minus.n106 15.9852
R22408 minus.n87 minus.n72 15.9852
R22409 minus.n26 minus.n11 15.9852
R22410 minus.n46 minus.n45 15.9852
R22411 minus.n115 minus.n62 14.0178
R22412 minus.n78 minus.n77 14.0178
R22413 minus.n17 minus.n16 14.0178
R22414 minus.n54 minus.n1 14.0178
R22415 minus.n122 minus.n60 12.1501
R22416 minus minus.n127 11.2487
R22417 minus.n118 minus.n62 10.575
R22418 minus.n57 minus.n1 10.575
R22419 minus.n120 minus.n119 9.49444
R22420 minus.n59 minus.n58 9.49444
R22421 minus.n108 minus.n107 8.60764
R22422 minus.n84 minus.n72 8.60764
R22423 minus.n23 minus.n11 8.60764
R22424 minus.n47 minus.n46 8.60764
R22425 minus.n100 minus.n68 6.6403
R22426 minus.n95 minus.n94 6.6403
R22427 minus.n34 minus.n33 6.6403
R22428 minus.n39 minus.n7 6.6403
R22429 minus.n127 minus.n126 4.80222
R22430 minus.n102 minus.n66 4.67295
R22431 minus.n90 minus.n89 4.67295
R22432 minus.n29 minus.n28 4.67295
R22433 minus.n41 minus.n5 4.67295
R22434 minus.n113 minus.n112 2.7056
R22435 minus.n82 minus.n74 2.7056
R22436 minus.n21 minus.n13 2.7056
R22437 minus.n52 minus.n51 2.7056
R22438 minus.n127 minus.n122 0.972091
R22439 minus.n126 minus.n125 0.716017
R22440 minus.n121 minus.n61 0.189894
R22441 minus.n117 minus.n61 0.189894
R22442 minus.n117 minus.n116 0.189894
R22443 minus.n116 minus.n63 0.189894
R22444 minus.n111 minus.n63 0.189894
R22445 minus.n111 minus.n110 0.189894
R22446 minus.n110 minus.n109 0.189894
R22447 minus.n109 minus.n65 0.189894
R22448 minus.n104 minus.n65 0.189894
R22449 minus.n104 minus.n103 0.189894
R22450 minus.n103 minus.n67 0.189894
R22451 minus.n99 minus.n67 0.189894
R22452 minus.n99 minus.n98 0.189894
R22453 minus.n98 minus.n69 0.189894
R22454 minus.n93 minus.n69 0.189894
R22455 minus.n93 minus.n92 0.189894
R22456 minus.n92 minus.n91 0.189894
R22457 minus.n91 minus.n71 0.189894
R22458 minus.n86 minus.n71 0.189894
R22459 minus.n86 minus.n85 0.189894
R22460 minus.n85 minus.n73 0.189894
R22461 minus.n81 minus.n73 0.189894
R22462 minus.n81 minus.n80 0.189894
R22463 minus.n80 minus.n75 0.189894
R22464 minus.n19 minus.n14 0.189894
R22465 minus.n20 minus.n19 0.189894
R22466 minus.n20 minus.n12 0.189894
R22467 minus.n24 minus.n12 0.189894
R22468 minus.n25 minus.n24 0.189894
R22469 minus.n25 minus.n10 0.189894
R22470 minus.n30 minus.n10 0.189894
R22471 minus.n31 minus.n30 0.189894
R22472 minus.n32 minus.n31 0.189894
R22473 minus.n32 minus.n8 0.189894
R22474 minus.n37 minus.n8 0.189894
R22475 minus.n38 minus.n37 0.189894
R22476 minus.n38 minus.n6 0.189894
R22477 minus.n42 minus.n6 0.189894
R22478 minus.n43 minus.n42 0.189894
R22479 minus.n43 minus.n4 0.189894
R22480 minus.n48 minus.n4 0.189894
R22481 minus.n49 minus.n48 0.189894
R22482 minus.n50 minus.n49 0.189894
R22483 minus.n50 minus.n2 0.189894
R22484 minus.n55 minus.n2 0.189894
R22485 minus.n56 minus.n55 0.189894
R22486 minus.n56 minus.n0 0.189894
R22487 minus.n60 minus.n0 0.189894
R22488 outputibias.n27 outputibias.n1 289.615
R22489 outputibias.n58 outputibias.n32 289.615
R22490 outputibias.n90 outputibias.n64 289.615
R22491 outputibias.n122 outputibias.n96 289.615
R22492 outputibias.n28 outputibias.n27 185
R22493 outputibias.n26 outputibias.n25 185
R22494 outputibias.n5 outputibias.n4 185
R22495 outputibias.n20 outputibias.n19 185
R22496 outputibias.n18 outputibias.n17 185
R22497 outputibias.n9 outputibias.n8 185
R22498 outputibias.n12 outputibias.n11 185
R22499 outputibias.n59 outputibias.n58 185
R22500 outputibias.n57 outputibias.n56 185
R22501 outputibias.n36 outputibias.n35 185
R22502 outputibias.n51 outputibias.n50 185
R22503 outputibias.n49 outputibias.n48 185
R22504 outputibias.n40 outputibias.n39 185
R22505 outputibias.n43 outputibias.n42 185
R22506 outputibias.n91 outputibias.n90 185
R22507 outputibias.n89 outputibias.n88 185
R22508 outputibias.n68 outputibias.n67 185
R22509 outputibias.n83 outputibias.n82 185
R22510 outputibias.n81 outputibias.n80 185
R22511 outputibias.n72 outputibias.n71 185
R22512 outputibias.n75 outputibias.n74 185
R22513 outputibias.n123 outputibias.n122 185
R22514 outputibias.n121 outputibias.n120 185
R22515 outputibias.n100 outputibias.n99 185
R22516 outputibias.n115 outputibias.n114 185
R22517 outputibias.n113 outputibias.n112 185
R22518 outputibias.n104 outputibias.n103 185
R22519 outputibias.n107 outputibias.n106 185
R22520 outputibias.n0 outputibias.t8 178.945
R22521 outputibias.n133 outputibias.t9 177.018
R22522 outputibias.n132 outputibias.t10 177.018
R22523 outputibias.n0 outputibias.t11 177.018
R22524 outputibias.t7 outputibias.n10 147.661
R22525 outputibias.t5 outputibias.n41 147.661
R22526 outputibias.t1 outputibias.n73 147.661
R22527 outputibias.t3 outputibias.n105 147.661
R22528 outputibias.n128 outputibias.t6 132.363
R22529 outputibias.n128 outputibias.t4 130.436
R22530 outputibias.n129 outputibias.t0 130.436
R22531 outputibias.n130 outputibias.t2 130.436
R22532 outputibias.n27 outputibias.n26 104.615
R22533 outputibias.n26 outputibias.n4 104.615
R22534 outputibias.n19 outputibias.n4 104.615
R22535 outputibias.n19 outputibias.n18 104.615
R22536 outputibias.n18 outputibias.n8 104.615
R22537 outputibias.n11 outputibias.n8 104.615
R22538 outputibias.n58 outputibias.n57 104.615
R22539 outputibias.n57 outputibias.n35 104.615
R22540 outputibias.n50 outputibias.n35 104.615
R22541 outputibias.n50 outputibias.n49 104.615
R22542 outputibias.n49 outputibias.n39 104.615
R22543 outputibias.n42 outputibias.n39 104.615
R22544 outputibias.n90 outputibias.n89 104.615
R22545 outputibias.n89 outputibias.n67 104.615
R22546 outputibias.n82 outputibias.n67 104.615
R22547 outputibias.n82 outputibias.n81 104.615
R22548 outputibias.n81 outputibias.n71 104.615
R22549 outputibias.n74 outputibias.n71 104.615
R22550 outputibias.n122 outputibias.n121 104.615
R22551 outputibias.n121 outputibias.n99 104.615
R22552 outputibias.n114 outputibias.n99 104.615
R22553 outputibias.n114 outputibias.n113 104.615
R22554 outputibias.n113 outputibias.n103 104.615
R22555 outputibias.n106 outputibias.n103 104.615
R22556 outputibias.n63 outputibias.n31 95.6354
R22557 outputibias.n63 outputibias.n62 94.6732
R22558 outputibias.n95 outputibias.n94 94.6732
R22559 outputibias.n127 outputibias.n126 94.6732
R22560 outputibias.n11 outputibias.t7 52.3082
R22561 outputibias.n42 outputibias.t5 52.3082
R22562 outputibias.n74 outputibias.t1 52.3082
R22563 outputibias.n106 outputibias.t3 52.3082
R22564 outputibias.n12 outputibias.n10 15.6674
R22565 outputibias.n43 outputibias.n41 15.6674
R22566 outputibias.n75 outputibias.n73 15.6674
R22567 outputibias.n107 outputibias.n105 15.6674
R22568 outputibias.n13 outputibias.n9 12.8005
R22569 outputibias.n44 outputibias.n40 12.8005
R22570 outputibias.n76 outputibias.n72 12.8005
R22571 outputibias.n108 outputibias.n104 12.8005
R22572 outputibias.n17 outputibias.n16 12.0247
R22573 outputibias.n48 outputibias.n47 12.0247
R22574 outputibias.n80 outputibias.n79 12.0247
R22575 outputibias.n112 outputibias.n111 12.0247
R22576 outputibias.n20 outputibias.n7 11.249
R22577 outputibias.n51 outputibias.n38 11.249
R22578 outputibias.n83 outputibias.n70 11.249
R22579 outputibias.n115 outputibias.n102 11.249
R22580 outputibias.n21 outputibias.n5 10.4732
R22581 outputibias.n52 outputibias.n36 10.4732
R22582 outputibias.n84 outputibias.n68 10.4732
R22583 outputibias.n116 outputibias.n100 10.4732
R22584 outputibias.n25 outputibias.n24 9.69747
R22585 outputibias.n56 outputibias.n55 9.69747
R22586 outputibias.n88 outputibias.n87 9.69747
R22587 outputibias.n120 outputibias.n119 9.69747
R22588 outputibias.n31 outputibias.n30 9.45567
R22589 outputibias.n62 outputibias.n61 9.45567
R22590 outputibias.n94 outputibias.n93 9.45567
R22591 outputibias.n126 outputibias.n125 9.45567
R22592 outputibias.n30 outputibias.n29 9.3005
R22593 outputibias.n3 outputibias.n2 9.3005
R22594 outputibias.n24 outputibias.n23 9.3005
R22595 outputibias.n22 outputibias.n21 9.3005
R22596 outputibias.n7 outputibias.n6 9.3005
R22597 outputibias.n16 outputibias.n15 9.3005
R22598 outputibias.n14 outputibias.n13 9.3005
R22599 outputibias.n61 outputibias.n60 9.3005
R22600 outputibias.n34 outputibias.n33 9.3005
R22601 outputibias.n55 outputibias.n54 9.3005
R22602 outputibias.n53 outputibias.n52 9.3005
R22603 outputibias.n38 outputibias.n37 9.3005
R22604 outputibias.n47 outputibias.n46 9.3005
R22605 outputibias.n45 outputibias.n44 9.3005
R22606 outputibias.n93 outputibias.n92 9.3005
R22607 outputibias.n66 outputibias.n65 9.3005
R22608 outputibias.n87 outputibias.n86 9.3005
R22609 outputibias.n85 outputibias.n84 9.3005
R22610 outputibias.n70 outputibias.n69 9.3005
R22611 outputibias.n79 outputibias.n78 9.3005
R22612 outputibias.n77 outputibias.n76 9.3005
R22613 outputibias.n125 outputibias.n124 9.3005
R22614 outputibias.n98 outputibias.n97 9.3005
R22615 outputibias.n119 outputibias.n118 9.3005
R22616 outputibias.n117 outputibias.n116 9.3005
R22617 outputibias.n102 outputibias.n101 9.3005
R22618 outputibias.n111 outputibias.n110 9.3005
R22619 outputibias.n109 outputibias.n108 9.3005
R22620 outputibias.n28 outputibias.n3 8.92171
R22621 outputibias.n59 outputibias.n34 8.92171
R22622 outputibias.n91 outputibias.n66 8.92171
R22623 outputibias.n123 outputibias.n98 8.92171
R22624 outputibias.n29 outputibias.n1 8.14595
R22625 outputibias.n60 outputibias.n32 8.14595
R22626 outputibias.n92 outputibias.n64 8.14595
R22627 outputibias.n124 outputibias.n96 8.14595
R22628 outputibias.n31 outputibias.n1 5.81868
R22629 outputibias.n62 outputibias.n32 5.81868
R22630 outputibias.n94 outputibias.n64 5.81868
R22631 outputibias.n126 outputibias.n96 5.81868
R22632 outputibias.n131 outputibias.n130 5.20947
R22633 outputibias.n29 outputibias.n28 5.04292
R22634 outputibias.n60 outputibias.n59 5.04292
R22635 outputibias.n92 outputibias.n91 5.04292
R22636 outputibias.n124 outputibias.n123 5.04292
R22637 outputibias.n131 outputibias.n127 4.42209
R22638 outputibias.n14 outputibias.n10 4.38594
R22639 outputibias.n45 outputibias.n41 4.38594
R22640 outputibias.n77 outputibias.n73 4.38594
R22641 outputibias.n109 outputibias.n105 4.38594
R22642 outputibias.n132 outputibias.n131 4.28454
R22643 outputibias.n25 outputibias.n3 4.26717
R22644 outputibias.n56 outputibias.n34 4.26717
R22645 outputibias.n88 outputibias.n66 4.26717
R22646 outputibias.n120 outputibias.n98 4.26717
R22647 outputibias.n24 outputibias.n5 3.49141
R22648 outputibias.n55 outputibias.n36 3.49141
R22649 outputibias.n87 outputibias.n68 3.49141
R22650 outputibias.n119 outputibias.n100 3.49141
R22651 outputibias.n21 outputibias.n20 2.71565
R22652 outputibias.n52 outputibias.n51 2.71565
R22653 outputibias.n84 outputibias.n83 2.71565
R22654 outputibias.n116 outputibias.n115 2.71565
R22655 outputibias.n17 outputibias.n7 1.93989
R22656 outputibias.n48 outputibias.n38 1.93989
R22657 outputibias.n80 outputibias.n70 1.93989
R22658 outputibias.n112 outputibias.n102 1.93989
R22659 outputibias.n130 outputibias.n129 1.9266
R22660 outputibias.n129 outputibias.n128 1.9266
R22661 outputibias.n133 outputibias.n132 1.92658
R22662 outputibias.n134 outputibias.n133 1.29913
R22663 outputibias.n16 outputibias.n9 1.16414
R22664 outputibias.n47 outputibias.n40 1.16414
R22665 outputibias.n79 outputibias.n72 1.16414
R22666 outputibias.n111 outputibias.n104 1.16414
R22667 outputibias.n127 outputibias.n95 0.962709
R22668 outputibias.n95 outputibias.n63 0.962709
R22669 outputibias.n13 outputibias.n12 0.388379
R22670 outputibias.n44 outputibias.n43 0.388379
R22671 outputibias.n76 outputibias.n75 0.388379
R22672 outputibias.n108 outputibias.n107 0.388379
R22673 outputibias.n134 outputibias.n0 0.337251
R22674 outputibias outputibias.n134 0.302375
R22675 outputibias.n30 outputibias.n2 0.155672
R22676 outputibias.n23 outputibias.n2 0.155672
R22677 outputibias.n23 outputibias.n22 0.155672
R22678 outputibias.n22 outputibias.n6 0.155672
R22679 outputibias.n15 outputibias.n6 0.155672
R22680 outputibias.n15 outputibias.n14 0.155672
R22681 outputibias.n61 outputibias.n33 0.155672
R22682 outputibias.n54 outputibias.n33 0.155672
R22683 outputibias.n54 outputibias.n53 0.155672
R22684 outputibias.n53 outputibias.n37 0.155672
R22685 outputibias.n46 outputibias.n37 0.155672
R22686 outputibias.n46 outputibias.n45 0.155672
R22687 outputibias.n93 outputibias.n65 0.155672
R22688 outputibias.n86 outputibias.n65 0.155672
R22689 outputibias.n86 outputibias.n85 0.155672
R22690 outputibias.n85 outputibias.n69 0.155672
R22691 outputibias.n78 outputibias.n69 0.155672
R22692 outputibias.n78 outputibias.n77 0.155672
R22693 outputibias.n125 outputibias.n97 0.155672
R22694 outputibias.n118 outputibias.n97 0.155672
R22695 outputibias.n118 outputibias.n117 0.155672
R22696 outputibias.n117 outputibias.n101 0.155672
R22697 outputibias.n110 outputibias.n101 0.155672
R22698 outputibias.n110 outputibias.n109 0.155672
R22699 diffpairibias.n0 diffpairibias.t18 436.822
R22700 diffpairibias.n21 diffpairibias.t19 435.479
R22701 diffpairibias.n20 diffpairibias.t16 435.479
R22702 diffpairibias.n19 diffpairibias.t17 435.479
R22703 diffpairibias.n18 diffpairibias.t21 435.479
R22704 diffpairibias.n0 diffpairibias.t22 435.479
R22705 diffpairibias.n1 diffpairibias.t20 435.479
R22706 diffpairibias.n2 diffpairibias.t23 435.479
R22707 diffpairibias.n10 diffpairibias.t0 377.536
R22708 diffpairibias.n10 diffpairibias.t8 376.193
R22709 diffpairibias.n11 diffpairibias.t10 376.193
R22710 diffpairibias.n12 diffpairibias.t6 376.193
R22711 diffpairibias.n13 diffpairibias.t2 376.193
R22712 diffpairibias.n14 diffpairibias.t12 376.193
R22713 diffpairibias.n15 diffpairibias.t4 376.193
R22714 diffpairibias.n16 diffpairibias.t14 376.193
R22715 diffpairibias.n3 diffpairibias.t1 113.368
R22716 diffpairibias.n3 diffpairibias.t9 112.698
R22717 diffpairibias.n4 diffpairibias.t11 112.698
R22718 diffpairibias.n5 diffpairibias.t7 112.698
R22719 diffpairibias.n6 diffpairibias.t3 112.698
R22720 diffpairibias.n7 diffpairibias.t13 112.698
R22721 diffpairibias.n8 diffpairibias.t5 112.698
R22722 diffpairibias.n9 diffpairibias.t15 112.698
R22723 diffpairibias.n17 diffpairibias.n16 4.77242
R22724 diffpairibias.n17 diffpairibias.n9 4.30807
R22725 diffpairibias.n18 diffpairibias.n17 4.13945
R22726 diffpairibias.n16 diffpairibias.n15 1.34352
R22727 diffpairibias.n15 diffpairibias.n14 1.34352
R22728 diffpairibias.n14 diffpairibias.n13 1.34352
R22729 diffpairibias.n13 diffpairibias.n12 1.34352
R22730 diffpairibias.n12 diffpairibias.n11 1.34352
R22731 diffpairibias.n11 diffpairibias.n10 1.34352
R22732 diffpairibias.n2 diffpairibias.n1 1.34352
R22733 diffpairibias.n1 diffpairibias.n0 1.34352
R22734 diffpairibias.n19 diffpairibias.n18 1.34352
R22735 diffpairibias.n20 diffpairibias.n19 1.34352
R22736 diffpairibias.n21 diffpairibias.n20 1.34352
R22737 diffpairibias.n22 diffpairibias.n21 0.862419
R22738 diffpairibias diffpairibias.n22 0.684875
R22739 diffpairibias.n9 diffpairibias.n8 0.672012
R22740 diffpairibias.n8 diffpairibias.n7 0.672012
R22741 diffpairibias.n7 diffpairibias.n6 0.672012
R22742 diffpairibias.n6 diffpairibias.n5 0.672012
R22743 diffpairibias.n5 diffpairibias.n4 0.672012
R22744 diffpairibias.n4 diffpairibias.n3 0.672012
R22745 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.116309p
C2 minus diffpairibias 5.39e-19
C3 commonsourceibias output 0.006808f
C4 vdd plus 0.088406f
C5 CSoutput minus 2.52746f
C6 plus diffpairibias 4.4e-19
C7 commonsourceibias outputibias 0.003832f
C8 vdd commonsourceibias 0.004218f
C9 CSoutput plus 0.894824f
C10 commonsourceibias diffpairibias 0.052851f
C11 CSoutput commonsourceibias 36.982002f
C12 minus plus 10.0542f
C13 minus commonsourceibias 0.515369f
C14 plus commonsourceibias 0.498793f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13571f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.149395p
C22 plus gnd 38.458603f
C23 minus gnd 30.00252f
C24 CSoutput gnd 0.101442p
C25 vdd gnd 0.408415p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 outputibias.t11 gnd 0.11477f
C74 outputibias.t8 gnd 0.115567f
C75 outputibias.n0 gnd 0.130108f
C76 outputibias.n1 gnd 0.001372f
C77 outputibias.n2 gnd 9.76e-19
C78 outputibias.n3 gnd 5.24e-19
C79 outputibias.n4 gnd 0.001239f
C80 outputibias.n5 gnd 5.55e-19
C81 outputibias.n6 gnd 9.76e-19
C82 outputibias.n7 gnd 5.24e-19
C83 outputibias.n8 gnd 0.001239f
C84 outputibias.n9 gnd 5.55e-19
C85 outputibias.n10 gnd 0.004176f
C86 outputibias.t7 gnd 0.00202f
C87 outputibias.n11 gnd 9.3e-19
C88 outputibias.n12 gnd 7.32e-19
C89 outputibias.n13 gnd 5.24e-19
C90 outputibias.n14 gnd 0.02322f
C91 outputibias.n15 gnd 9.76e-19
C92 outputibias.n16 gnd 5.24e-19
C93 outputibias.n17 gnd 5.55e-19
C94 outputibias.n18 gnd 0.001239f
C95 outputibias.n19 gnd 0.001239f
C96 outputibias.n20 gnd 5.55e-19
C97 outputibias.n21 gnd 5.24e-19
C98 outputibias.n22 gnd 9.76e-19
C99 outputibias.n23 gnd 9.76e-19
C100 outputibias.n24 gnd 5.24e-19
C101 outputibias.n25 gnd 5.55e-19
C102 outputibias.n26 gnd 0.001239f
C103 outputibias.n27 gnd 0.002683f
C104 outputibias.n28 gnd 5.55e-19
C105 outputibias.n29 gnd 5.24e-19
C106 outputibias.n30 gnd 0.002256f
C107 outputibias.n31 gnd 0.005781f
C108 outputibias.n32 gnd 0.001372f
C109 outputibias.n33 gnd 9.76e-19
C110 outputibias.n34 gnd 5.24e-19
C111 outputibias.n35 gnd 0.001239f
C112 outputibias.n36 gnd 5.55e-19
C113 outputibias.n37 gnd 9.76e-19
C114 outputibias.n38 gnd 5.24e-19
C115 outputibias.n39 gnd 0.001239f
C116 outputibias.n40 gnd 5.55e-19
C117 outputibias.n41 gnd 0.004176f
C118 outputibias.t5 gnd 0.00202f
C119 outputibias.n42 gnd 9.3e-19
C120 outputibias.n43 gnd 7.32e-19
C121 outputibias.n44 gnd 5.24e-19
C122 outputibias.n45 gnd 0.02322f
C123 outputibias.n46 gnd 9.76e-19
C124 outputibias.n47 gnd 5.24e-19
C125 outputibias.n48 gnd 5.55e-19
C126 outputibias.n49 gnd 0.001239f
C127 outputibias.n50 gnd 0.001239f
C128 outputibias.n51 gnd 5.55e-19
C129 outputibias.n52 gnd 5.24e-19
C130 outputibias.n53 gnd 9.76e-19
C131 outputibias.n54 gnd 9.76e-19
C132 outputibias.n55 gnd 5.24e-19
C133 outputibias.n56 gnd 5.55e-19
C134 outputibias.n57 gnd 0.001239f
C135 outputibias.n58 gnd 0.002683f
C136 outputibias.n59 gnd 5.55e-19
C137 outputibias.n60 gnd 5.24e-19
C138 outputibias.n61 gnd 0.002256f
C139 outputibias.n62 gnd 0.005197f
C140 outputibias.n63 gnd 0.121892f
C141 outputibias.n64 gnd 0.001372f
C142 outputibias.n65 gnd 9.76e-19
C143 outputibias.n66 gnd 5.24e-19
C144 outputibias.n67 gnd 0.001239f
C145 outputibias.n68 gnd 5.55e-19
C146 outputibias.n69 gnd 9.76e-19
C147 outputibias.n70 gnd 5.24e-19
C148 outputibias.n71 gnd 0.001239f
C149 outputibias.n72 gnd 5.55e-19
C150 outputibias.n73 gnd 0.004176f
C151 outputibias.t1 gnd 0.00202f
C152 outputibias.n74 gnd 9.3e-19
C153 outputibias.n75 gnd 7.32e-19
C154 outputibias.n76 gnd 5.24e-19
C155 outputibias.n77 gnd 0.02322f
C156 outputibias.n78 gnd 9.76e-19
C157 outputibias.n79 gnd 5.24e-19
C158 outputibias.n80 gnd 5.55e-19
C159 outputibias.n81 gnd 0.001239f
C160 outputibias.n82 gnd 0.001239f
C161 outputibias.n83 gnd 5.55e-19
C162 outputibias.n84 gnd 5.24e-19
C163 outputibias.n85 gnd 9.76e-19
C164 outputibias.n86 gnd 9.76e-19
C165 outputibias.n87 gnd 5.24e-19
C166 outputibias.n88 gnd 5.55e-19
C167 outputibias.n89 gnd 0.001239f
C168 outputibias.n90 gnd 0.002683f
C169 outputibias.n91 gnd 5.55e-19
C170 outputibias.n92 gnd 5.24e-19
C171 outputibias.n93 gnd 0.002256f
C172 outputibias.n94 gnd 0.005197f
C173 outputibias.n95 gnd 0.064513f
C174 outputibias.n96 gnd 0.001372f
C175 outputibias.n97 gnd 9.76e-19
C176 outputibias.n98 gnd 5.24e-19
C177 outputibias.n99 gnd 0.001239f
C178 outputibias.n100 gnd 5.55e-19
C179 outputibias.n101 gnd 9.76e-19
C180 outputibias.n102 gnd 5.24e-19
C181 outputibias.n103 gnd 0.001239f
C182 outputibias.n104 gnd 5.55e-19
C183 outputibias.n105 gnd 0.004176f
C184 outputibias.t3 gnd 0.00202f
C185 outputibias.n106 gnd 9.3e-19
C186 outputibias.n107 gnd 7.32e-19
C187 outputibias.n108 gnd 5.24e-19
C188 outputibias.n109 gnd 0.02322f
C189 outputibias.n110 gnd 9.76e-19
C190 outputibias.n111 gnd 5.24e-19
C191 outputibias.n112 gnd 5.55e-19
C192 outputibias.n113 gnd 0.001239f
C193 outputibias.n114 gnd 0.001239f
C194 outputibias.n115 gnd 5.55e-19
C195 outputibias.n116 gnd 5.24e-19
C196 outputibias.n117 gnd 9.76e-19
C197 outputibias.n118 gnd 9.76e-19
C198 outputibias.n119 gnd 5.24e-19
C199 outputibias.n120 gnd 5.55e-19
C200 outputibias.n121 gnd 0.001239f
C201 outputibias.n122 gnd 0.002683f
C202 outputibias.n123 gnd 5.55e-19
C203 outputibias.n124 gnd 5.24e-19
C204 outputibias.n125 gnd 0.002256f
C205 outputibias.n126 gnd 0.005197f
C206 outputibias.n127 gnd 0.084814f
C207 outputibias.t2 gnd 0.108319f
C208 outputibias.t0 gnd 0.108319f
C209 outputibias.t4 gnd 0.108319f
C210 outputibias.t6 gnd 0.109238f
C211 outputibias.n128 gnd 0.134674f
C212 outputibias.n129 gnd 0.07244f
C213 outputibias.n130 gnd 0.079818f
C214 outputibias.n131 gnd 0.164901f
C215 outputibias.t10 gnd 0.11477f
C216 outputibias.n132 gnd 0.067481f
C217 outputibias.t9 gnd 0.11477f
C218 outputibias.n133 gnd 0.065115f
C219 outputibias.n134 gnd 0.029159f
C220 minus.n0 gnd 0.031226f
C221 minus.t13 gnd 0.525058f
C222 minus.n1 gnd 0.212357f
C223 minus.n2 gnd 0.031226f
C224 minus.t11 gnd 0.525058f
C225 minus.n3 gnd 0.026683f
C226 minus.n4 gnd 0.031226f
C227 minus.t17 gnd 0.525058f
C228 minus.t24 gnd 0.525058f
C229 minus.n5 gnd 0.212357f
C230 minus.n6 gnd 0.031226f
C231 minus.t21 gnd 0.525058f
C232 minus.n7 gnd 0.212357f
C233 minus.n8 gnd 0.031226f
C234 minus.t27 gnd 0.525058f
C235 minus.n9 gnd 0.02538f
C236 minus.n10 gnd 0.031226f
C237 minus.t26 gnd 0.525058f
C238 minus.t5 gnd 0.525058f
C239 minus.n11 gnd 0.212357f
C240 minus.n12 gnd 0.031226f
C241 minus.t9 gnd 0.525058f
C242 minus.n13 gnd 0.212357f
C243 minus.n14 gnd 0.132519f
C244 minus.t14 gnd 0.525058f
C245 minus.t20 gnd 0.587372f
C246 minus.n15 gnd 0.248266f
C247 minus.n16 gnd 0.243188f
C248 minus.n17 gnd 0.040011f
C249 minus.n18 gnd 0.035336f
C250 minus.n19 gnd 0.031226f
C251 minus.n20 gnd 0.031226f
C252 minus.n21 gnd 0.037315f
C253 minus.n22 gnd 0.026683f
C254 minus.n23 gnd 0.040668f
C255 minus.n24 gnd 0.031226f
C256 minus.n25 gnd 0.031226f
C257 minus.n26 gnd 0.038842f
C258 minus.n27 gnd 0.036505f
C259 minus.n28 gnd 0.212357f
C260 minus.n29 gnd 0.039115f
C261 minus.n30 gnd 0.031226f
C262 minus.n31 gnd 0.031226f
C263 minus.n32 gnd 0.031226f
C264 minus.n33 gnd 0.040171f
C265 minus.n34 gnd 0.212357f
C266 minus.n35 gnd 0.037673f
C267 minus.n36 gnd 0.037673f
C268 minus.n37 gnd 0.031226f
C269 minus.n38 gnd 0.031226f
C270 minus.n39 gnd 0.040171f
C271 minus.n40 gnd 0.02538f
C272 minus.n41 gnd 0.039115f
C273 minus.n42 gnd 0.031226f
C274 minus.n43 gnd 0.031226f
C275 minus.n44 gnd 0.036505f
C276 minus.n45 gnd 0.038842f
C277 minus.n46 gnd 0.212357f
C278 minus.n47 gnd 0.040668f
C279 minus.n48 gnd 0.031226f
C280 minus.n49 gnd 0.031226f
C281 minus.n50 gnd 0.031226f
C282 minus.n51 gnd 0.037315f
C283 minus.n52 gnd 0.212357f
C284 minus.n53 gnd 0.035336f
C285 minus.n54 gnd 0.040011f
C286 minus.n55 gnd 0.031226f
C287 minus.n56 gnd 0.031226f
C288 minus.n57 gnd 0.040735f
C289 minus.n58 gnd 0.011348f
C290 minus.t10 gnd 0.56785f
C291 minus.n59 gnd 0.245873f
C292 minus.n60 gnd 0.365799f
C293 minus.n61 gnd 0.031226f
C294 minus.t8 gnd 0.56785f
C295 minus.t12 gnd 0.525058f
C296 minus.n62 gnd 0.212357f
C297 minus.n63 gnd 0.031226f
C298 minus.t18 gnd 0.525058f
C299 minus.n64 gnd 0.026683f
C300 minus.n65 gnd 0.031226f
C301 minus.t25 gnd 0.525058f
C302 minus.t22 gnd 0.525058f
C303 minus.n66 gnd 0.212357f
C304 minus.n67 gnd 0.031226f
C305 minus.t19 gnd 0.525058f
C306 minus.n68 gnd 0.212357f
C307 minus.n69 gnd 0.031226f
C308 minus.t7 gnd 0.525058f
C309 minus.n70 gnd 0.02538f
C310 minus.n71 gnd 0.031226f
C311 minus.t6 gnd 0.525058f
C312 minus.t16 gnd 0.525058f
C313 minus.n72 gnd 0.212357f
C314 minus.n73 gnd 0.031226f
C315 minus.t15 gnd 0.525058f
C316 minus.n74 gnd 0.212357f
C317 minus.n75 gnd 0.132519f
C318 minus.t23 gnd 0.525058f
C319 minus.t28 gnd 0.587372f
C320 minus.n76 gnd 0.248266f
C321 minus.n77 gnd 0.243188f
C322 minus.n78 gnd 0.040011f
C323 minus.n79 gnd 0.035336f
C324 minus.n80 gnd 0.031226f
C325 minus.n81 gnd 0.031226f
C326 minus.n82 gnd 0.037315f
C327 minus.n83 gnd 0.026683f
C328 minus.n84 gnd 0.040668f
C329 minus.n85 gnd 0.031226f
C330 minus.n86 gnd 0.031226f
C331 minus.n87 gnd 0.038842f
C332 minus.n88 gnd 0.036505f
C333 minus.n89 gnd 0.212357f
C334 minus.n90 gnd 0.039115f
C335 minus.n91 gnd 0.031226f
C336 minus.n92 gnd 0.031226f
C337 minus.n93 gnd 0.031226f
C338 minus.n94 gnd 0.040171f
C339 minus.n95 gnd 0.212357f
C340 minus.n96 gnd 0.037673f
C341 minus.n97 gnd 0.037673f
C342 minus.n98 gnd 0.031226f
C343 minus.n99 gnd 0.031226f
C344 minus.n100 gnd 0.040171f
C345 minus.n101 gnd 0.02538f
C346 minus.n102 gnd 0.039115f
C347 minus.n103 gnd 0.031226f
C348 minus.n104 gnd 0.031226f
C349 minus.n105 gnd 0.036505f
C350 minus.n106 gnd 0.038842f
C351 minus.n107 gnd 0.212357f
C352 minus.n108 gnd 0.040668f
C353 minus.n109 gnd 0.031226f
C354 minus.n110 gnd 0.031226f
C355 minus.n111 gnd 0.031226f
C356 minus.n112 gnd 0.037315f
C357 minus.n113 gnd 0.212357f
C358 minus.n114 gnd 0.035336f
C359 minus.n115 gnd 0.040011f
C360 minus.n116 gnd 0.031226f
C361 minus.n117 gnd 0.031226f
C362 minus.n118 gnd 0.040735f
C363 minus.n119 gnd 0.011348f
C364 minus.n120 gnd 0.245873f
C365 minus.n121 gnd 1.1391f
C366 minus.n122 gnd 1.67326f
C367 minus.t4 gnd 0.009626f
C368 minus.t3 gnd 0.009626f
C369 minus.n123 gnd 0.031653f
C370 minus.t0 gnd 0.009626f
C371 minus.t2 gnd 0.009626f
C372 minus.n124 gnd 0.031219f
C373 minus.n125 gnd 0.266439f
C374 minus.t1 gnd 0.053577f
C375 minus.n126 gnd 0.145393f
C376 minus.n127 gnd 1.77594f
C377 output.t15 gnd 0.464308f
C378 output.t4 gnd 0.044422f
C379 output.t9 gnd 0.044422f
C380 output.n0 gnd 0.364624f
C381 output.n1 gnd 0.614102f
C382 output.t13 gnd 0.044422f
C383 output.t5 gnd 0.044422f
C384 output.n2 gnd 0.364624f
C385 output.n3 gnd 0.350265f
C386 output.t8 gnd 0.044422f
C387 output.t6 gnd 0.044422f
C388 output.n4 gnd 0.364624f
C389 output.n5 gnd 0.350265f
C390 output.t12 gnd 0.044422f
C391 output.t14 gnd 0.044422f
C392 output.n6 gnd 0.364624f
C393 output.n7 gnd 0.350265f
C394 output.t17 gnd 0.044422f
C395 output.t10 gnd 0.044422f
C396 output.n8 gnd 0.364624f
C397 output.n9 gnd 0.350265f
C398 output.t11 gnd 0.044422f
C399 output.t2 gnd 0.044422f
C400 output.n10 gnd 0.364624f
C401 output.n11 gnd 0.350265f
C402 output.t3 gnd 0.044422f
C403 output.t7 gnd 0.044422f
C404 output.n12 gnd 0.364624f
C405 output.n13 gnd 0.350265f
C406 output.t16 gnd 0.462979f
C407 output.n14 gnd 0.28994f
C408 output.n15 gnd 0.015803f
C409 output.n16 gnd 0.011243f
C410 output.n17 gnd 0.006041f
C411 output.n18 gnd 0.01428f
C412 output.n19 gnd 0.006397f
C413 output.n20 gnd 0.011243f
C414 output.n21 gnd 0.006041f
C415 output.n22 gnd 0.01428f
C416 output.n23 gnd 0.006397f
C417 output.n24 gnd 0.048111f
C418 output.t18 gnd 0.023274f
C419 output.n25 gnd 0.01071f
C420 output.n26 gnd 0.008435f
C421 output.n27 gnd 0.006041f
C422 output.n28 gnd 0.267512f
C423 output.n29 gnd 0.011243f
C424 output.n30 gnd 0.006041f
C425 output.n31 gnd 0.006397f
C426 output.n32 gnd 0.01428f
C427 output.n33 gnd 0.01428f
C428 output.n34 gnd 0.006397f
C429 output.n35 gnd 0.006041f
C430 output.n36 gnd 0.011243f
C431 output.n37 gnd 0.011243f
C432 output.n38 gnd 0.006041f
C433 output.n39 gnd 0.006397f
C434 output.n40 gnd 0.01428f
C435 output.n41 gnd 0.030913f
C436 output.n42 gnd 0.006397f
C437 output.n43 gnd 0.006041f
C438 output.n44 gnd 0.025987f
C439 output.n45 gnd 0.097665f
C440 output.n46 gnd 0.015803f
C441 output.n47 gnd 0.011243f
C442 output.n48 gnd 0.006041f
C443 output.n49 gnd 0.01428f
C444 output.n50 gnd 0.006397f
C445 output.n51 gnd 0.011243f
C446 output.n52 gnd 0.006041f
C447 output.n53 gnd 0.01428f
C448 output.n54 gnd 0.006397f
C449 output.n55 gnd 0.048111f
C450 output.t1 gnd 0.023274f
C451 output.n56 gnd 0.01071f
C452 output.n57 gnd 0.008435f
C453 output.n58 gnd 0.006041f
C454 output.n59 gnd 0.267512f
C455 output.n60 gnd 0.011243f
C456 output.n61 gnd 0.006041f
C457 output.n62 gnd 0.006397f
C458 output.n63 gnd 0.01428f
C459 output.n64 gnd 0.01428f
C460 output.n65 gnd 0.006397f
C461 output.n66 gnd 0.006041f
C462 output.n67 gnd 0.011243f
C463 output.n68 gnd 0.011243f
C464 output.n69 gnd 0.006041f
C465 output.n70 gnd 0.006397f
C466 output.n71 gnd 0.01428f
C467 output.n72 gnd 0.030913f
C468 output.n73 gnd 0.006397f
C469 output.n74 gnd 0.006041f
C470 output.n75 gnd 0.025987f
C471 output.n76 gnd 0.09306f
C472 output.n77 gnd 1.65264f
C473 output.n78 gnd 0.015803f
C474 output.n79 gnd 0.011243f
C475 output.n80 gnd 0.006041f
C476 output.n81 gnd 0.01428f
C477 output.n82 gnd 0.006397f
C478 output.n83 gnd 0.011243f
C479 output.n84 gnd 0.006041f
C480 output.n85 gnd 0.01428f
C481 output.n86 gnd 0.006397f
C482 output.n87 gnd 0.048111f
C483 output.t19 gnd 0.023274f
C484 output.n88 gnd 0.01071f
C485 output.n89 gnd 0.008435f
C486 output.n90 gnd 0.006041f
C487 output.n91 gnd 0.267512f
C488 output.n92 gnd 0.011243f
C489 output.n93 gnd 0.006041f
C490 output.n94 gnd 0.006397f
C491 output.n95 gnd 0.01428f
C492 output.n96 gnd 0.01428f
C493 output.n97 gnd 0.006397f
C494 output.n98 gnd 0.006041f
C495 output.n99 gnd 0.011243f
C496 output.n100 gnd 0.011243f
C497 output.n101 gnd 0.006041f
C498 output.n102 gnd 0.006397f
C499 output.n103 gnd 0.01428f
C500 output.n104 gnd 0.030913f
C501 output.n105 gnd 0.006397f
C502 output.n106 gnd 0.006041f
C503 output.n107 gnd 0.025987f
C504 output.n108 gnd 0.09306f
C505 output.n109 gnd 0.713089f
C506 output.n110 gnd 0.015803f
C507 output.n111 gnd 0.011243f
C508 output.n112 gnd 0.006041f
C509 output.n113 gnd 0.01428f
C510 output.n114 gnd 0.006397f
C511 output.n115 gnd 0.011243f
C512 output.n116 gnd 0.006041f
C513 output.n117 gnd 0.01428f
C514 output.n118 gnd 0.006397f
C515 output.n119 gnd 0.048111f
C516 output.t0 gnd 0.023274f
C517 output.n120 gnd 0.01071f
C518 output.n121 gnd 0.008435f
C519 output.n122 gnd 0.006041f
C520 output.n123 gnd 0.267512f
C521 output.n124 gnd 0.011243f
C522 output.n125 gnd 0.006041f
C523 output.n126 gnd 0.006397f
C524 output.n127 gnd 0.01428f
C525 output.n128 gnd 0.01428f
C526 output.n129 gnd 0.006397f
C527 output.n130 gnd 0.006041f
C528 output.n131 gnd 0.011243f
C529 output.n132 gnd 0.011243f
C530 output.n133 gnd 0.006041f
C531 output.n134 gnd 0.006397f
C532 output.n135 gnd 0.01428f
C533 output.n136 gnd 0.030913f
C534 output.n137 gnd 0.006397f
C535 output.n138 gnd 0.006041f
C536 output.n139 gnd 0.025987f
C537 output.n140 gnd 0.09306f
C538 output.n141 gnd 1.67353f
C539 a_n3106_n452.t35 gnd 0.10001f
C540 a_n3106_n452.t46 gnd 1.03942f
C541 a_n3106_n452.n0 gnd 0.392946f
C542 a_n3106_n452.t22 gnd 1.29145f
C543 a_n3106_n452.n1 gnd 1.22854f
C544 a_n3106_n452.t23 gnd 1.03942f
C545 a_n3106_n452.n2 gnd 0.392946f
C546 a_n3106_n452.t15 gnd 0.10001f
C547 a_n3106_n452.t17 gnd 0.10001f
C548 a_n3106_n452.n3 gnd 0.816794f
C549 a_n3106_n452.n4 gnd 0.411618f
C550 a_n3106_n452.t11 gnd 0.10001f
C551 a_n3106_n452.t19 gnd 0.10001f
C552 a_n3106_n452.n5 gnd 0.816794f
C553 a_n3106_n452.n6 gnd 0.411618f
C554 a_n3106_n452.t2 gnd 0.10001f
C555 a_n3106_n452.t8 gnd 0.10001f
C556 a_n3106_n452.n7 gnd 0.816794f
C557 a_n3106_n452.n8 gnd 0.411618f
C558 a_n3106_n452.t3 gnd 0.10001f
C559 a_n3106_n452.t18 gnd 0.10001f
C560 a_n3106_n452.n9 gnd 0.816794f
C561 a_n3106_n452.n10 gnd 0.411618f
C562 a_n3106_n452.t27 gnd 0.10001f
C563 a_n3106_n452.t7 gnd 0.10001f
C564 a_n3106_n452.n11 gnd 0.816794f
C565 a_n3106_n452.n12 gnd 0.411618f
C566 a_n3106_n452.t24 gnd 1.03942f
C567 a_n3106_n452.n13 gnd 0.972974f
C568 a_n3106_n452.t21 gnd 1.29145f
C569 a_n3106_n452.n14 gnd 0.909591f
C570 a_n3106_n452.t0 gnd 1.29145f
C571 a_n3106_n452.n15 gnd 0.909591f
C572 a_n3106_n452.t13 gnd 1.29145f
C573 a_n3106_n452.n16 gnd 0.909591f
C574 a_n3106_n452.t20 gnd 1.29145f
C575 a_n3106_n452.n17 gnd 0.909591f
C576 a_n3106_n452.t54 gnd 1.29145f
C577 a_n3106_n452.n18 gnd 0.909591f
C578 a_n3106_n452.t55 gnd 1.29145f
C579 a_n3106_n452.n19 gnd 0.909591f
C580 a_n3106_n452.t25 gnd 1.29145f
C581 a_n3106_n452.n20 gnd 0.789472f
C582 a_n3106_n452.n21 gnd 0.948419f
C583 a_n3106_n452.t37 gnd 1.03941f
C584 a_n3106_n452.n22 gnd 0.645631f
C585 a_n3106_n452.t34 gnd 0.10001f
C586 a_n3106_n452.t51 gnd 0.10001f
C587 a_n3106_n452.n23 gnd 0.816793f
C588 a_n3106_n452.n24 gnd 0.41162f
C589 a_n3106_n452.t45 gnd 0.10001f
C590 a_n3106_n452.t49 gnd 0.10001f
C591 a_n3106_n452.n25 gnd 0.816793f
C592 a_n3106_n452.n26 gnd 0.41162f
C593 a_n3106_n452.t50 gnd 0.10001f
C594 a_n3106_n452.t38 gnd 0.10001f
C595 a_n3106_n452.n27 gnd 0.816793f
C596 a_n3106_n452.n28 gnd 0.41162f
C597 a_n3106_n452.t39 gnd 0.10001f
C598 a_n3106_n452.t30 gnd 0.10001f
C599 a_n3106_n452.n29 gnd 0.816793f
C600 a_n3106_n452.n30 gnd 0.41162f
C601 a_n3106_n452.t32 gnd 0.10001f
C602 a_n3106_n452.t48 gnd 0.10001f
C603 a_n3106_n452.n31 gnd 0.816793f
C604 a_n3106_n452.n32 gnd 0.41162f
C605 a_n3106_n452.t43 gnd 1.03941f
C606 a_n3106_n452.n33 gnd 0.39295f
C607 a_n3106_n452.t5 gnd 1.03941f
C608 a_n3106_n452.n34 gnd 0.39295f
C609 a_n3106_n452.t26 gnd 0.10001f
C610 a_n3106_n452.t10 gnd 0.10001f
C611 a_n3106_n452.n35 gnd 0.816793f
C612 a_n3106_n452.n36 gnd 0.41162f
C613 a_n3106_n452.t53 gnd 0.10001f
C614 a_n3106_n452.t16 gnd 0.10001f
C615 a_n3106_n452.n37 gnd 0.816793f
C616 a_n3106_n452.n38 gnd 0.41162f
C617 a_n3106_n452.t4 gnd 0.10001f
C618 a_n3106_n452.t1 gnd 0.10001f
C619 a_n3106_n452.n39 gnd 0.816793f
C620 a_n3106_n452.n40 gnd 0.41162f
C621 a_n3106_n452.t14 gnd 0.10001f
C622 a_n3106_n452.t28 gnd 0.10001f
C623 a_n3106_n452.n41 gnd 0.816793f
C624 a_n3106_n452.n42 gnd 0.41162f
C625 a_n3106_n452.t12 gnd 0.10001f
C626 a_n3106_n452.t6 gnd 0.10001f
C627 a_n3106_n452.n43 gnd 0.816793f
C628 a_n3106_n452.n44 gnd 0.41162f
C629 a_n3106_n452.t9 gnd 1.03941f
C630 a_n3106_n452.n45 gnd 0.645631f
C631 a_n3106_n452.n46 gnd 1.05146f
C632 a_n3106_n452.t33 gnd 1.03941f
C633 a_n3106_n452.n47 gnd 0.972978f
C634 a_n3106_n452.t31 gnd 0.10001f
C635 a_n3106_n452.t29 gnd 0.10001f
C636 a_n3106_n452.n48 gnd 0.816794f
C637 a_n3106_n452.n49 gnd 0.411618f
C638 a_n3106_n452.t42 gnd 0.10001f
C639 a_n3106_n452.t47 gnd 0.10001f
C640 a_n3106_n452.n50 gnd 0.816794f
C641 a_n3106_n452.n51 gnd 0.411618f
C642 a_n3106_n452.t40 gnd 0.10001f
C643 a_n3106_n452.t44 gnd 0.10001f
C644 a_n3106_n452.n52 gnd 0.816794f
C645 a_n3106_n452.n53 gnd 0.411618f
C646 a_n3106_n452.t36 gnd 0.10001f
C647 a_n3106_n452.t41 gnd 0.10001f
C648 a_n3106_n452.n54 gnd 0.816794f
C649 a_n3106_n452.n55 gnd 0.411618f
C650 a_n3106_n452.n56 gnd 0.411617f
C651 a_n3106_n452.n57 gnd 0.816796f
C652 a_n3106_n452.t52 gnd 0.10001f
C653 plus.n0 gnd 0.023269f
C654 plus.t20 gnd 0.423154f
C655 plus.t23 gnd 0.391266f
C656 plus.n1 gnd 0.158245f
C657 plus.n2 gnd 0.023269f
C658 plus.t6 gnd 0.391266f
C659 plus.n3 gnd 0.019884f
C660 plus.n4 gnd 0.023269f
C661 plus.t12 gnd 0.391266f
C662 plus.t8 gnd 0.391266f
C663 plus.n5 gnd 0.158245f
C664 plus.n6 gnd 0.023269f
C665 plus.t7 gnd 0.391266f
C666 plus.n7 gnd 0.158245f
C667 plus.n8 gnd 0.023269f
C668 plus.t19 gnd 0.391266f
C669 plus.n9 gnd 0.018913f
C670 plus.n10 gnd 0.023269f
C671 plus.t18 gnd 0.391266f
C672 plus.t27 gnd 0.391266f
C673 plus.n11 gnd 0.158245f
C674 plus.n12 gnd 0.023269f
C675 plus.t25 gnd 0.391266f
C676 plus.n13 gnd 0.158245f
C677 plus.n14 gnd 0.098752f
C678 plus.t9 gnd 0.391266f
C679 plus.t14 gnd 0.437702f
C680 plus.n15 gnd 0.185005f
C681 plus.n16 gnd 0.181221f
C682 plus.n17 gnd 0.029816f
C683 plus.n18 gnd 0.026332f
C684 plus.n19 gnd 0.023269f
C685 plus.n20 gnd 0.023269f
C686 plus.n21 gnd 0.027807f
C687 plus.n22 gnd 0.019884f
C688 plus.n23 gnd 0.030305f
C689 plus.n24 gnd 0.023269f
C690 plus.n25 gnd 0.023269f
C691 plus.n26 gnd 0.028945f
C692 plus.n27 gnd 0.027203f
C693 plus.n28 gnd 0.158245f
C694 plus.n29 gnd 0.029148f
C695 plus.n30 gnd 0.023269f
C696 plus.n31 gnd 0.023269f
C697 plus.n32 gnd 0.023269f
C698 plus.n33 gnd 0.029935f
C699 plus.n34 gnd 0.158245f
C700 plus.n35 gnd 0.028074f
C701 plus.n36 gnd 0.028074f
C702 plus.n37 gnd 0.023269f
C703 plus.n38 gnd 0.023269f
C704 plus.n39 gnd 0.029935f
C705 plus.n40 gnd 0.018913f
C706 plus.n41 gnd 0.029148f
C707 plus.n42 gnd 0.023269f
C708 plus.n43 gnd 0.023269f
C709 plus.n44 gnd 0.027203f
C710 plus.n45 gnd 0.028945f
C711 plus.n46 gnd 0.158245f
C712 plus.n47 gnd 0.030305f
C713 plus.n48 gnd 0.023269f
C714 plus.n49 gnd 0.023269f
C715 plus.n50 gnd 0.023269f
C716 plus.n51 gnd 0.027807f
C717 plus.n52 gnd 0.158245f
C718 plus.n53 gnd 0.026332f
C719 plus.n54 gnd 0.029816f
C720 plus.n55 gnd 0.023269f
C721 plus.n56 gnd 0.023269f
C722 plus.n57 gnd 0.030355f
C723 plus.n58 gnd 0.008457f
C724 plus.n59 gnd 0.183222f
C725 plus.n60 gnd 0.266602f
C726 plus.n61 gnd 0.023269f
C727 plus.t28 gnd 0.391266f
C728 plus.n62 gnd 0.158245f
C729 plus.n63 gnd 0.023269f
C730 plus.t26 gnd 0.391266f
C731 plus.n64 gnd 0.019884f
C732 plus.n65 gnd 0.023269f
C733 plus.t10 gnd 0.391266f
C734 plus.t15 gnd 0.391266f
C735 plus.n66 gnd 0.158245f
C736 plus.n67 gnd 0.023269f
C737 plus.t13 gnd 0.391266f
C738 plus.n68 gnd 0.158245f
C739 plus.n69 gnd 0.023269f
C740 plus.t17 gnd 0.391266f
C741 plus.n70 gnd 0.018913f
C742 plus.n71 gnd 0.023269f
C743 plus.t16 gnd 0.391266f
C744 plus.t21 gnd 0.391266f
C745 plus.n72 gnd 0.158245f
C746 plus.n73 gnd 0.023269f
C747 plus.t22 gnd 0.391266f
C748 plus.n74 gnd 0.158245f
C749 plus.n75 gnd 0.098752f
C750 plus.t5 gnd 0.391266f
C751 plus.t11 gnd 0.437702f
C752 plus.n76 gnd 0.185005f
C753 plus.n77 gnd 0.181221f
C754 plus.n78 gnd 0.029816f
C755 plus.n79 gnd 0.026332f
C756 plus.n80 gnd 0.023269f
C757 plus.n81 gnd 0.023269f
C758 plus.n82 gnd 0.027807f
C759 plus.n83 gnd 0.019884f
C760 plus.n84 gnd 0.030305f
C761 plus.n85 gnd 0.023269f
C762 plus.n86 gnd 0.023269f
C763 plus.n87 gnd 0.028945f
C764 plus.n88 gnd 0.027203f
C765 plus.n89 gnd 0.158245f
C766 plus.n90 gnd 0.029148f
C767 plus.n91 gnd 0.023269f
C768 plus.n92 gnd 0.023269f
C769 plus.n93 gnd 0.023269f
C770 plus.n94 gnd 0.029935f
C771 plus.n95 gnd 0.158245f
C772 plus.n96 gnd 0.028074f
C773 plus.n97 gnd 0.028074f
C774 plus.n98 gnd 0.023269f
C775 plus.n99 gnd 0.023269f
C776 plus.n100 gnd 0.029935f
C777 plus.n101 gnd 0.018913f
C778 plus.n102 gnd 0.029148f
C779 plus.n103 gnd 0.023269f
C780 plus.n104 gnd 0.023269f
C781 plus.n105 gnd 0.027203f
C782 plus.n106 gnd 0.028945f
C783 plus.n107 gnd 0.158245f
C784 plus.n108 gnd 0.030305f
C785 plus.n109 gnd 0.023269f
C786 plus.n110 gnd 0.023269f
C787 plus.n111 gnd 0.023269f
C788 plus.n112 gnd 0.027807f
C789 plus.n113 gnd 0.158245f
C790 plus.n114 gnd 0.026332f
C791 plus.n115 gnd 0.029816f
C792 plus.n116 gnd 0.023269f
C793 plus.n117 gnd 0.023269f
C794 plus.n118 gnd 0.030355f
C795 plus.n119 gnd 0.008457f
C796 plus.t24 gnd 0.423154f
C797 plus.n120 gnd 0.183222f
C798 plus.n121 gnd 0.83954f
C799 plus.n122 gnd 1.23765f
C800 plus.t1 gnd 0.040169f
C801 plus.t2 gnd 0.007173f
C802 plus.t4 gnd 0.007173f
C803 plus.n123 gnd 0.023264f
C804 plus.n124 gnd 0.1806f
C805 plus.t3 gnd 0.007173f
C806 plus.t0 gnd 0.007173f
C807 plus.n125 gnd 0.023264f
C808 plus.n126 gnd 0.135562f
C809 plus.n127 gnd 2.83926f
C810 a_n1808_13878.t4 gnd 0.185195f
C811 a_n1808_13878.t0 gnd 0.185195f
C812 a_n1808_13878.t2 gnd 0.185195f
C813 a_n1808_13878.n0 gnd 1.4598f
C814 a_n1808_13878.t6 gnd 0.185195f
C815 a_n1808_13878.t1 gnd 0.185195f
C816 a_n1808_13878.n1 gnd 1.45825f
C817 a_n1808_13878.n2 gnd 2.03762f
C818 a_n1808_13878.t5 gnd 0.185195f
C819 a_n1808_13878.t9 gnd 0.185195f
C820 a_n1808_13878.n3 gnd 1.46067f
C821 a_n1808_13878.t10 gnd 0.185195f
C822 a_n1808_13878.t3 gnd 0.185195f
C823 a_n1808_13878.n4 gnd 1.45825f
C824 a_n1808_13878.n5 gnd 1.31079f
C825 a_n1808_13878.t7 gnd 0.185195f
C826 a_n1808_13878.t8 gnd 0.185195f
C827 a_n1808_13878.n6 gnd 1.45825f
C828 a_n1808_13878.n7 gnd 1.80025f
C829 a_n1808_13878.t13 gnd 1.73408f
C830 a_n1808_13878.t16 gnd 0.185195f
C831 a_n1808_13878.t17 gnd 0.185195f
C832 a_n1808_13878.n8 gnd 1.30452f
C833 a_n1808_13878.n9 gnd 1.4576f
C834 a_n1808_13878.t12 gnd 1.73062f
C835 a_n1808_13878.n10 gnd 0.733487f
C836 a_n1808_13878.t15 gnd 1.73062f
C837 a_n1808_13878.n11 gnd 0.733487f
C838 a_n1808_13878.t18 gnd 0.185195f
C839 a_n1808_13878.t19 gnd 0.185195f
C840 a_n1808_13878.n12 gnd 1.30452f
C841 a_n1808_13878.n13 gnd 0.74059f
C842 a_n1808_13878.t14 gnd 1.73062f
C843 a_n1808_13878.n14 gnd 1.7272f
C844 a_n1808_13878.n15 gnd 2.51438f
C845 a_n1808_13878.n16 gnd 3.69301f
C846 a_n1808_13878.n17 gnd 1.45826f
C847 a_n1808_13878.t11 gnd 0.185195f
C848 a_n2848_n452.n0 gnd 3.415f
C849 a_n2848_n452.n1 gnd 0.285666f
C850 a_n2848_n452.n2 gnd 0.492471f
C851 a_n2848_n452.n3 gnd 0.664435f
C852 a_n2848_n452.n4 gnd 0.215942f
C853 a_n2848_n452.n5 gnd 0.282512f
C854 a_n2848_n452.n6 gnd 0.546457f
C855 a_n2848_n452.n7 gnd 0.526038f
C856 a_n2848_n452.n8 gnd 0.204894f
C857 a_n2848_n452.n9 gnd 0.150908f
C858 a_n2848_n452.n10 gnd 0.23718f
C859 a_n2848_n452.n11 gnd 0.183194f
C860 a_n2848_n452.n12 gnd 0.204894f
C861 a_n2848_n452.n13 gnd 1.0063f
C862 a_n2848_n452.n14 gnd 0.150908f
C863 a_n2848_n452.n15 gnd 0.580023f
C864 a_n2848_n452.n16 gnd 0.432289f
C865 a_n2848_n452.n17 gnd 0.215942f
C866 a_n2848_n452.n18 gnd 0.492471f
C867 a_n2848_n452.n19 gnd 0.282512f
C868 a_n2848_n452.n20 gnd 0.438486f
C869 a_n2848_n452.n21 gnd 0.215942f
C870 a_n2848_n452.n22 gnd 0.731535f
C871 a_n2848_n452.n23 gnd 0.282512f
C872 a_n2848_n452.n24 gnd 1.17886f
C873 a_n2848_n452.n25 gnd 1.91568f
C874 a_n2848_n452.n26 gnd 1.14458f
C875 a_n2848_n452.n27 gnd 1.77783f
C876 a_n2848_n452.n28 gnd 0.377489f
C877 a_n2848_n452.n29 gnd 3.11576f
C878 a_n2848_n452.n30 gnd 0.377488f
C879 a_n2848_n452.n31 gnd 3.20158f
C880 a_n2848_n452.n32 gnd 0.008361f
C881 a_n2848_n452.n34 gnd 0.285666f
C882 a_n2848_n452.n35 gnd 0.008361f
C883 a_n2848_n452.n37 gnd 0.285666f
C884 a_n2848_n452.n38 gnd 0.008361f
C885 a_n2848_n452.n39 gnd 0.28526f
C886 a_n2848_n452.n40 gnd 0.008361f
C887 a_n2848_n452.n41 gnd 0.28526f
C888 a_n2848_n452.n42 gnd 0.008361f
C889 a_n2848_n452.n43 gnd 0.28526f
C890 a_n2848_n452.n44 gnd 0.008361f
C891 a_n2848_n452.n45 gnd 0.28526f
C892 a_n2848_n452.n47 gnd 0.285666f
C893 a_n2848_n452.n48 gnd 0.008361f
C894 a_n2848_n452.n50 gnd 0.285666f
C895 a_n2848_n452.t23 gnd 0.708223f
C896 a_n2848_n452.t25 gnd 0.696704f
C897 a_n2848_n452.t19 gnd 0.696704f
C898 a_n2848_n452.t4 gnd 0.116496f
C899 a_n2848_n452.t44 gnd 0.116496f
C900 a_n2848_n452.n52 gnd 1.03243f
C901 a_n2848_n452.t9 gnd 0.116496f
C902 a_n2848_n452.t47 gnd 0.116496f
C903 a_n2848_n452.n53 gnd 1.0294f
C904 a_n2848_n452.n54 gnd 0.912817f
C905 a_n2848_n452.t14 gnd 0.116496f
C906 a_n2848_n452.t3 gnd 0.116496f
C907 a_n2848_n452.n55 gnd 1.0294f
C908 a_n2848_n452.t5 gnd 0.116496f
C909 a_n2848_n452.t8 gnd 0.116496f
C910 a_n2848_n452.n56 gnd 1.03243f
C911 a_n2848_n452.t46 gnd 0.116496f
C912 a_n2848_n452.t11 gnd 0.116496f
C913 a_n2848_n452.n57 gnd 1.0294f
C914 a_n2848_n452.n58 gnd 0.912817f
C915 a_n2848_n452.t0 gnd 0.116496f
C916 a_n2848_n452.t12 gnd 0.116496f
C917 a_n2848_n452.n59 gnd 1.0294f
C918 a_n2848_n452.t43 gnd 0.116496f
C919 a_n2848_n452.t45 gnd 0.116496f
C920 a_n2848_n452.n60 gnd 1.0294f
C921 a_n2848_n452.n61 gnd 3.15028f
C922 a_n2848_n452.t6 gnd 0.116496f
C923 a_n2848_n452.t2 gnd 0.116496f
C924 a_n2848_n452.n62 gnd 1.0294f
C925 a_n2848_n452.n63 gnd 0.449443f
C926 a_n2848_n452.t40 gnd 0.116496f
C927 a_n2848_n452.t1 gnd 0.116496f
C928 a_n2848_n452.n64 gnd 1.0294f
C929 a_n2848_n452.t39 gnd 0.116496f
C930 a_n2848_n452.t42 gnd 0.116496f
C931 a_n2848_n452.n65 gnd 1.03243f
C932 a_n2848_n452.t41 gnd 0.116496f
C933 a_n2848_n452.t13 gnd 0.116496f
C934 a_n2848_n452.n66 gnd 1.0294f
C935 a_n2848_n452.n67 gnd 0.912814f
C936 a_n2848_n452.t7 gnd 0.116496f
C937 a_n2848_n452.t10 gnd 0.116496f
C938 a_n2848_n452.n68 gnd 1.0294f
C939 a_n2848_n452.t37 gnd 0.696704f
C940 a_n2848_n452.n69 gnd 0.302425f
C941 a_n2848_n452.t33 gnd 0.696704f
C942 a_n2848_n452.t15 gnd 0.708223f
C943 a_n2848_n452.t75 gnd 0.711378f
C944 a_n2848_n452.t58 gnd 0.696704f
C945 a_n2848_n452.t62 gnd 0.696704f
C946 a_n2848_n452.t52 gnd 0.696704f
C947 a_n2848_n452.n70 gnd 0.306315f
C948 a_n2848_n452.t67 gnd 0.696704f
C949 a_n2848_n452.t73 gnd 0.708223f
C950 a_n2848_n452.t30 gnd 1.40246f
C951 a_n2848_n452.t28 gnd 0.14978f
C952 a_n2848_n452.t36 gnd 0.14978f
C953 a_n2848_n452.n71 gnd 1.05505f
C954 a_n2848_n452.t18 gnd 0.14978f
C955 a_n2848_n452.t22 gnd 0.14978f
C956 a_n2848_n452.n72 gnd 1.05505f
C957 a_n2848_n452.t32 gnd 1.39967f
C958 a_n2848_n452.t17 gnd 0.696704f
C959 a_n2848_n452.n73 gnd 0.306315f
C960 a_n2848_n452.t21 gnd 0.696704f
C961 a_n2848_n452.t27 gnd 0.696704f
C962 a_n2848_n452.t56 gnd 0.696704f
C963 a_n2848_n452.n74 gnd 0.306315f
C964 a_n2848_n452.t65 gnd 0.696704f
C965 a_n2848_n452.t71 gnd 0.696704f
C966 a_n2848_n452.t70 gnd 0.711378f
C967 a_n2848_n452.n75 gnd 0.308932f
C968 a_n2848_n452.t50 gnd 0.696704f
C969 a_n2848_n452.n76 gnd 0.302425f
C970 a_n2848_n452.n77 gnd 0.308933f
C971 a_n2848_n452.t51 gnd 0.708223f
C972 a_n2848_n452.t29 gnd 0.711378f
C973 a_n2848_n452.n78 gnd 0.308932f
C974 a_n2848_n452.t35 gnd 0.696704f
C975 a_n2848_n452.n79 gnd 0.302425f
C976 a_n2848_n452.n80 gnd 0.308933f
C977 a_n2848_n452.t31 gnd 0.708223f
C978 a_n2848_n452.n81 gnd 1.13204f
C979 a_n2848_n452.t55 gnd 0.696704f
C980 a_n2848_n452.n82 gnd 0.302425f
C981 a_n2848_n452.t61 gnd 0.696704f
C982 a_n2848_n452.n83 gnd 0.302425f
C983 a_n2848_n452.t53 gnd 0.696704f
C984 a_n2848_n452.n84 gnd 0.302425f
C985 a_n2848_n452.t66 gnd 0.696704f
C986 a_n2848_n452.n85 gnd 0.302425f
C987 a_n2848_n452.t57 gnd 0.696704f
C988 a_n2848_n452.n86 gnd 0.296933f
C989 a_n2848_n452.t48 gnd 0.696704f
C990 a_n2848_n452.n87 gnd 0.306315f
C991 a_n2848_n452.t59 gnd 0.708378f
C992 a_n2848_n452.t68 gnd 0.696704f
C993 a_n2848_n452.n88 gnd 0.296933f
C994 a_n2848_n452.t54 gnd 0.696704f
C995 a_n2848_n452.n89 gnd 0.306315f
C996 a_n2848_n452.t63 gnd 0.708378f
C997 a_n2848_n452.t72 gnd 0.696704f
C998 a_n2848_n452.n90 gnd 0.296933f
C999 a_n2848_n452.t60 gnd 0.696704f
C1000 a_n2848_n452.n91 gnd 0.306315f
C1001 a_n2848_n452.t74 gnd 0.708378f
C1002 a_n2848_n452.t64 gnd 0.696704f
C1003 a_n2848_n452.n92 gnd 0.296933f
C1004 a_n2848_n452.t49 gnd 0.696704f
C1005 a_n2848_n452.n93 gnd 0.306315f
C1006 a_n2848_n452.t69 gnd 0.708378f
C1007 a_n2848_n452.n94 gnd 1.33845f
C1008 a_n2848_n452.n95 gnd 0.308933f
C1009 a_n2848_n452.n96 gnd 0.302425f
C1010 a_n2848_n452.n97 gnd 0.308932f
C1011 a_n2848_n452.n98 gnd 0.308933f
C1012 a_n2848_n452.n99 gnd 0.01225f
C1013 a_n2848_n452.n100 gnd 0.302425f
C1014 a_n2848_n452.n101 gnd 0.308933f
C1015 a_n2848_n452.n102 gnd 0.786935f
C1016 a_n2848_n452.t24 gnd 1.39967f
C1017 a_n2848_n452.t26 gnd 0.14978f
C1018 a_n2848_n452.t20 gnd 0.14978f
C1019 a_n2848_n452.n103 gnd 1.05505f
C1020 a_n2848_n452.t38 gnd 0.14978f
C1021 a_n2848_n452.t34 gnd 0.14978f
C1022 a_n2848_n452.n104 gnd 1.05505f
C1023 a_n2848_n452.t16 gnd 1.40246f
C1024 vdd.t5 gnd 0.038352f
C1025 vdd.t1 gnd 0.038352f
C1026 vdd.n0 gnd 0.302486f
C1027 vdd.t154 gnd 0.038352f
C1028 vdd.t263 gnd 0.038352f
C1029 vdd.n1 gnd 0.301987f
C1030 vdd.n2 gnd 0.278489f
C1031 vdd.t259 gnd 0.038352f
C1032 vdd.t16 gnd 0.038352f
C1033 vdd.n3 gnd 0.301987f
C1034 vdd.n4 gnd 0.140842f
C1035 vdd.t7 gnd 0.038352f
C1036 vdd.t152 gnd 0.038352f
C1037 vdd.n5 gnd 0.301987f
C1038 vdd.n6 gnd 0.132155f
C1039 vdd.t156 gnd 0.038352f
C1040 vdd.t261 gnd 0.038352f
C1041 vdd.n7 gnd 0.302486f
C1042 vdd.t148 gnd 0.038352f
C1043 vdd.t9 gnd 0.038352f
C1044 vdd.n8 gnd 0.301987f
C1045 vdd.n9 gnd 0.278489f
C1046 vdd.t158 gnd 0.038352f
C1047 vdd.t257 gnd 0.038352f
C1048 vdd.n10 gnd 0.301987f
C1049 vdd.n11 gnd 0.140842f
C1050 vdd.t13 gnd 0.038352f
C1051 vdd.t160 gnd 0.038352f
C1052 vdd.n12 gnd 0.301987f
C1053 vdd.n13 gnd 0.132155f
C1054 vdd.n14 gnd 0.093431f
C1055 vdd.t251 gnd 0.021306f
C1056 vdd.t255 gnd 0.021306f
C1057 vdd.n15 gnd 0.196117f
C1058 vdd.t254 gnd 0.021306f
C1059 vdd.t240 gnd 0.021306f
C1060 vdd.n16 gnd 0.195543f
C1061 vdd.n17 gnd 0.340307f
C1062 vdd.t245 gnd 0.021306f
C1063 vdd.t250 gnd 0.021306f
C1064 vdd.n18 gnd 0.195543f
C1065 vdd.n19 gnd 0.140789f
C1066 vdd.t252 gnd 0.021306f
C1067 vdd.t242 gnd 0.021306f
C1068 vdd.n20 gnd 0.196117f
C1069 vdd.t246 gnd 0.021306f
C1070 vdd.t244 gnd 0.021306f
C1071 vdd.n21 gnd 0.195543f
C1072 vdd.n22 gnd 0.340307f
C1073 vdd.t248 gnd 0.021306f
C1074 vdd.t253 gnd 0.021306f
C1075 vdd.n23 gnd 0.195543f
C1076 vdd.n24 gnd 0.140789f
C1077 vdd.t241 gnd 0.021306f
C1078 vdd.t243 gnd 0.021306f
C1079 vdd.n25 gnd 0.195543f
C1080 vdd.t249 gnd 0.021306f
C1081 vdd.t247 gnd 0.021306f
C1082 vdd.n26 gnd 0.195543f
C1083 vdd.n27 gnd 22.528301f
C1084 vdd.n28 gnd 8.31901f
C1085 vdd.n29 gnd 0.005811f
C1086 vdd.n30 gnd 0.005392f
C1087 vdd.n31 gnd 0.002983f
C1088 vdd.n32 gnd 0.006849f
C1089 vdd.n33 gnd 0.002898f
C1090 vdd.n34 gnd 0.003068f
C1091 vdd.n35 gnd 0.005392f
C1092 vdd.n36 gnd 0.002898f
C1093 vdd.n37 gnd 0.006849f
C1094 vdd.n38 gnd 0.003068f
C1095 vdd.n39 gnd 0.005392f
C1096 vdd.n40 gnd 0.002898f
C1097 vdd.n41 gnd 0.005137f
C1098 vdd.n42 gnd 0.005152f
C1099 vdd.t22 gnd 0.014715f
C1100 vdd.n43 gnd 0.03274f
C1101 vdd.n44 gnd 0.170386f
C1102 vdd.n45 gnd 0.002898f
C1103 vdd.n46 gnd 0.003068f
C1104 vdd.n47 gnd 0.006849f
C1105 vdd.n48 gnd 0.006849f
C1106 vdd.n49 gnd 0.003068f
C1107 vdd.n50 gnd 0.002898f
C1108 vdd.n51 gnd 0.005392f
C1109 vdd.n52 gnd 0.005392f
C1110 vdd.n53 gnd 0.002898f
C1111 vdd.n54 gnd 0.003068f
C1112 vdd.n55 gnd 0.006849f
C1113 vdd.n56 gnd 0.006849f
C1114 vdd.n57 gnd 0.003068f
C1115 vdd.n58 gnd 0.002898f
C1116 vdd.n59 gnd 0.005392f
C1117 vdd.n60 gnd 0.005392f
C1118 vdd.n61 gnd 0.002898f
C1119 vdd.n62 gnd 0.003068f
C1120 vdd.n63 gnd 0.006849f
C1121 vdd.n64 gnd 0.006849f
C1122 vdd.n65 gnd 0.016193f
C1123 vdd.n66 gnd 0.002983f
C1124 vdd.n67 gnd 0.002898f
C1125 vdd.n68 gnd 0.013938f
C1126 vdd.n69 gnd 0.009731f
C1127 vdd.t131 gnd 0.03409f
C1128 vdd.t83 gnd 0.03409f
C1129 vdd.n70 gnd 0.234293f
C1130 vdd.n71 gnd 0.184235f
C1131 vdd.t144 gnd 0.03409f
C1132 vdd.t56 gnd 0.03409f
C1133 vdd.n72 gnd 0.234293f
C1134 vdd.n73 gnd 0.148677f
C1135 vdd.t119 gnd 0.03409f
C1136 vdd.t76 gnd 0.03409f
C1137 vdd.n74 gnd 0.234293f
C1138 vdd.n75 gnd 0.148677f
C1139 vdd.t139 gnd 0.03409f
C1140 vdd.t115 gnd 0.03409f
C1141 vdd.n76 gnd 0.234293f
C1142 vdd.n77 gnd 0.148677f
C1143 vdd.t30 gnd 0.03409f
C1144 vdd.t69 gnd 0.03409f
C1145 vdd.n78 gnd 0.234293f
C1146 vdd.n79 gnd 0.148677f
C1147 vdd.t38 gnd 0.03409f
C1148 vdd.t85 gnd 0.03409f
C1149 vdd.n80 gnd 0.234293f
C1150 vdd.n81 gnd 0.148677f
C1151 vdd.t62 gnd 0.03409f
C1152 vdd.t125 gnd 0.03409f
C1153 vdd.n82 gnd 0.234293f
C1154 vdd.n83 gnd 0.148677f
C1155 vdd.n84 gnd 0.005811f
C1156 vdd.n85 gnd 0.005392f
C1157 vdd.n86 gnd 0.002983f
C1158 vdd.n87 gnd 0.006849f
C1159 vdd.n88 gnd 0.002898f
C1160 vdd.n89 gnd 0.003068f
C1161 vdd.n90 gnd 0.005392f
C1162 vdd.n91 gnd 0.002898f
C1163 vdd.n92 gnd 0.006849f
C1164 vdd.n93 gnd 0.003068f
C1165 vdd.n94 gnd 0.005392f
C1166 vdd.n95 gnd 0.002898f
C1167 vdd.n96 gnd 0.005137f
C1168 vdd.n97 gnd 0.005152f
C1169 vdd.t42 gnd 0.014715f
C1170 vdd.n98 gnd 0.03274f
C1171 vdd.n99 gnd 0.170386f
C1172 vdd.n100 gnd 0.002898f
C1173 vdd.n101 gnd 0.003068f
C1174 vdd.n102 gnd 0.006849f
C1175 vdd.n103 gnd 0.006849f
C1176 vdd.n104 gnd 0.003068f
C1177 vdd.n105 gnd 0.002898f
C1178 vdd.n106 gnd 0.005392f
C1179 vdd.n107 gnd 0.005392f
C1180 vdd.n108 gnd 0.002898f
C1181 vdd.n109 gnd 0.003068f
C1182 vdd.n110 gnd 0.006849f
C1183 vdd.n111 gnd 0.006849f
C1184 vdd.n112 gnd 0.003068f
C1185 vdd.n113 gnd 0.002898f
C1186 vdd.n114 gnd 0.005392f
C1187 vdd.n115 gnd 0.005392f
C1188 vdd.n116 gnd 0.002898f
C1189 vdd.n117 gnd 0.003068f
C1190 vdd.n118 gnd 0.006849f
C1191 vdd.n119 gnd 0.006849f
C1192 vdd.n120 gnd 0.016193f
C1193 vdd.n121 gnd 0.002983f
C1194 vdd.n122 gnd 0.002898f
C1195 vdd.n123 gnd 0.013938f
C1196 vdd.n124 gnd 0.009425f
C1197 vdd.n125 gnd 0.110616f
C1198 vdd.n126 gnd 0.005811f
C1199 vdd.n127 gnd 0.005392f
C1200 vdd.n128 gnd 0.002983f
C1201 vdd.n129 gnd 0.006849f
C1202 vdd.n130 gnd 0.002898f
C1203 vdd.n131 gnd 0.003068f
C1204 vdd.n132 gnd 0.005392f
C1205 vdd.n133 gnd 0.002898f
C1206 vdd.n134 gnd 0.006849f
C1207 vdd.n135 gnd 0.003068f
C1208 vdd.n136 gnd 0.005392f
C1209 vdd.n137 gnd 0.002898f
C1210 vdd.n138 gnd 0.005137f
C1211 vdd.n139 gnd 0.005152f
C1212 vdd.t87 gnd 0.014715f
C1213 vdd.n140 gnd 0.03274f
C1214 vdd.n141 gnd 0.170386f
C1215 vdd.n142 gnd 0.002898f
C1216 vdd.n143 gnd 0.003068f
C1217 vdd.n144 gnd 0.006849f
C1218 vdd.n145 gnd 0.006849f
C1219 vdd.n146 gnd 0.003068f
C1220 vdd.n147 gnd 0.002898f
C1221 vdd.n148 gnd 0.005392f
C1222 vdd.n149 gnd 0.005392f
C1223 vdd.n150 gnd 0.002898f
C1224 vdd.n151 gnd 0.003068f
C1225 vdd.n152 gnd 0.006849f
C1226 vdd.n153 gnd 0.006849f
C1227 vdd.n154 gnd 0.003068f
C1228 vdd.n155 gnd 0.002898f
C1229 vdd.n156 gnd 0.005392f
C1230 vdd.n157 gnd 0.005392f
C1231 vdd.n158 gnd 0.002898f
C1232 vdd.n159 gnd 0.003068f
C1233 vdd.n160 gnd 0.006849f
C1234 vdd.n161 gnd 0.006849f
C1235 vdd.n162 gnd 0.016193f
C1236 vdd.n163 gnd 0.002983f
C1237 vdd.n164 gnd 0.002898f
C1238 vdd.n165 gnd 0.013938f
C1239 vdd.n166 gnd 0.009731f
C1240 vdd.t89 gnd 0.03409f
C1241 vdd.t111 gnd 0.03409f
C1242 vdd.n167 gnd 0.234293f
C1243 vdd.n168 gnd 0.184235f
C1244 vdd.t26 gnd 0.03409f
C1245 vdd.t80 gnd 0.03409f
C1246 vdd.n169 gnd 0.234293f
C1247 vdd.n170 gnd 0.148677f
C1248 vdd.t109 gnd 0.03409f
C1249 vdd.t146 gnd 0.03409f
C1250 vdd.n171 gnd 0.234293f
C1251 vdd.n172 gnd 0.148677f
C1252 vdd.t64 gnd 0.03409f
C1253 vdd.t66 gnd 0.03409f
C1254 vdd.n173 gnd 0.234293f
C1255 vdd.n174 gnd 0.148677f
C1256 vdd.t133 gnd 0.03409f
C1257 vdd.t59 gnd 0.03409f
C1258 vdd.n175 gnd 0.234293f
C1259 vdd.n176 gnd 0.148677f
C1260 vdd.t60 gnd 0.03409f
C1261 vdd.t129 gnd 0.03409f
C1262 vdd.n177 gnd 0.234293f
C1263 vdd.n178 gnd 0.148677f
C1264 vdd.t130 gnd 0.03409f
C1265 vdd.t36 gnd 0.03409f
C1266 vdd.n179 gnd 0.234293f
C1267 vdd.n180 gnd 0.148677f
C1268 vdd.n181 gnd 0.005811f
C1269 vdd.n182 gnd 0.005392f
C1270 vdd.n183 gnd 0.002983f
C1271 vdd.n184 gnd 0.006849f
C1272 vdd.n185 gnd 0.002898f
C1273 vdd.n186 gnd 0.003068f
C1274 vdd.n187 gnd 0.005392f
C1275 vdd.n188 gnd 0.002898f
C1276 vdd.n189 gnd 0.006849f
C1277 vdd.n190 gnd 0.003068f
C1278 vdd.n191 gnd 0.005392f
C1279 vdd.n192 gnd 0.002898f
C1280 vdd.n193 gnd 0.005137f
C1281 vdd.n194 gnd 0.005152f
C1282 vdd.t110 gnd 0.014715f
C1283 vdd.n195 gnd 0.03274f
C1284 vdd.n196 gnd 0.170386f
C1285 vdd.n197 gnd 0.002898f
C1286 vdd.n198 gnd 0.003068f
C1287 vdd.n199 gnd 0.006849f
C1288 vdd.n200 gnd 0.006849f
C1289 vdd.n201 gnd 0.003068f
C1290 vdd.n202 gnd 0.002898f
C1291 vdd.n203 gnd 0.005392f
C1292 vdd.n204 gnd 0.005392f
C1293 vdd.n205 gnd 0.002898f
C1294 vdd.n206 gnd 0.003068f
C1295 vdd.n207 gnd 0.006849f
C1296 vdd.n208 gnd 0.006849f
C1297 vdd.n209 gnd 0.003068f
C1298 vdd.n210 gnd 0.002898f
C1299 vdd.n211 gnd 0.005392f
C1300 vdd.n212 gnd 0.005392f
C1301 vdd.n213 gnd 0.002898f
C1302 vdd.n214 gnd 0.003068f
C1303 vdd.n215 gnd 0.006849f
C1304 vdd.n216 gnd 0.006849f
C1305 vdd.n217 gnd 0.016193f
C1306 vdd.n218 gnd 0.002983f
C1307 vdd.n219 gnd 0.002898f
C1308 vdd.n220 gnd 0.013938f
C1309 vdd.n221 gnd 0.009425f
C1310 vdd.n222 gnd 0.065805f
C1311 vdd.n223 gnd 0.237115f
C1312 vdd.n224 gnd 0.005811f
C1313 vdd.n225 gnd 0.005392f
C1314 vdd.n226 gnd 0.002983f
C1315 vdd.n227 gnd 0.006849f
C1316 vdd.n228 gnd 0.002898f
C1317 vdd.n229 gnd 0.003068f
C1318 vdd.n230 gnd 0.005392f
C1319 vdd.n231 gnd 0.002898f
C1320 vdd.n232 gnd 0.006849f
C1321 vdd.n233 gnd 0.003068f
C1322 vdd.n234 gnd 0.005392f
C1323 vdd.n235 gnd 0.002898f
C1324 vdd.n236 gnd 0.005137f
C1325 vdd.n237 gnd 0.005152f
C1326 vdd.t98 gnd 0.014715f
C1327 vdd.n238 gnd 0.03274f
C1328 vdd.n239 gnd 0.170386f
C1329 vdd.n240 gnd 0.002898f
C1330 vdd.n241 gnd 0.003068f
C1331 vdd.n242 gnd 0.006849f
C1332 vdd.n243 gnd 0.006849f
C1333 vdd.n244 gnd 0.003068f
C1334 vdd.n245 gnd 0.002898f
C1335 vdd.n246 gnd 0.005392f
C1336 vdd.n247 gnd 0.005392f
C1337 vdd.n248 gnd 0.002898f
C1338 vdd.n249 gnd 0.003068f
C1339 vdd.n250 gnd 0.006849f
C1340 vdd.n251 gnd 0.006849f
C1341 vdd.n252 gnd 0.003068f
C1342 vdd.n253 gnd 0.002898f
C1343 vdd.n254 gnd 0.005392f
C1344 vdd.n255 gnd 0.005392f
C1345 vdd.n256 gnd 0.002898f
C1346 vdd.n257 gnd 0.003068f
C1347 vdd.n258 gnd 0.006849f
C1348 vdd.n259 gnd 0.006849f
C1349 vdd.n260 gnd 0.016193f
C1350 vdd.n261 gnd 0.002983f
C1351 vdd.n262 gnd 0.002898f
C1352 vdd.n263 gnd 0.013938f
C1353 vdd.n264 gnd 0.009731f
C1354 vdd.t99 gnd 0.03409f
C1355 vdd.t123 gnd 0.03409f
C1356 vdd.n265 gnd 0.234293f
C1357 vdd.n266 gnd 0.184235f
C1358 vdd.t47 gnd 0.03409f
C1359 vdd.t97 gnd 0.03409f
C1360 vdd.n267 gnd 0.234293f
C1361 vdd.n268 gnd 0.148677f
C1362 vdd.t118 gnd 0.03409f
C1363 vdd.t44 gnd 0.03409f
C1364 vdd.n269 gnd 0.234293f
C1365 vdd.n270 gnd 0.148677f
C1366 vdd.t77 gnd 0.03409f
C1367 vdd.t79 gnd 0.03409f
C1368 vdd.n271 gnd 0.234293f
C1369 vdd.n272 gnd 0.148677f
C1370 vdd.t142 gnd 0.03409f
C1371 vdd.t72 gnd 0.03409f
C1372 vdd.n273 gnd 0.234293f
C1373 vdd.n274 gnd 0.148677f
C1374 vdd.t73 gnd 0.03409f
C1375 vdd.t140 gnd 0.03409f
C1376 vdd.n275 gnd 0.234293f
C1377 vdd.n276 gnd 0.148677f
C1378 vdd.t141 gnd 0.03409f
C1379 vdd.t52 gnd 0.03409f
C1380 vdd.n277 gnd 0.234293f
C1381 vdd.n278 gnd 0.148677f
C1382 vdd.n279 gnd 0.005811f
C1383 vdd.n280 gnd 0.005392f
C1384 vdd.n281 gnd 0.002983f
C1385 vdd.n282 gnd 0.006849f
C1386 vdd.n283 gnd 0.002898f
C1387 vdd.n284 gnd 0.003068f
C1388 vdd.n285 gnd 0.005392f
C1389 vdd.n286 gnd 0.002898f
C1390 vdd.n287 gnd 0.006849f
C1391 vdd.n288 gnd 0.003068f
C1392 vdd.n289 gnd 0.005392f
C1393 vdd.n290 gnd 0.002898f
C1394 vdd.n291 gnd 0.005137f
C1395 vdd.n292 gnd 0.005152f
C1396 vdd.t124 gnd 0.014715f
C1397 vdd.n293 gnd 0.03274f
C1398 vdd.n294 gnd 0.170386f
C1399 vdd.n295 gnd 0.002898f
C1400 vdd.n296 gnd 0.003068f
C1401 vdd.n297 gnd 0.006849f
C1402 vdd.n298 gnd 0.006849f
C1403 vdd.n299 gnd 0.003068f
C1404 vdd.n300 gnd 0.002898f
C1405 vdd.n301 gnd 0.005392f
C1406 vdd.n302 gnd 0.005392f
C1407 vdd.n303 gnd 0.002898f
C1408 vdd.n304 gnd 0.003068f
C1409 vdd.n305 gnd 0.006849f
C1410 vdd.n306 gnd 0.006849f
C1411 vdd.n307 gnd 0.003068f
C1412 vdd.n308 gnd 0.002898f
C1413 vdd.n309 gnd 0.005392f
C1414 vdd.n310 gnd 0.005392f
C1415 vdd.n311 gnd 0.002898f
C1416 vdd.n312 gnd 0.003068f
C1417 vdd.n313 gnd 0.006849f
C1418 vdd.n314 gnd 0.006849f
C1419 vdd.n315 gnd 0.016193f
C1420 vdd.n316 gnd 0.002983f
C1421 vdd.n317 gnd 0.002898f
C1422 vdd.n318 gnd 0.013938f
C1423 vdd.n319 gnd 0.009425f
C1424 vdd.n320 gnd 0.065805f
C1425 vdd.n321 gnd 0.265537f
C1426 vdd.n322 gnd 0.008138f
C1427 vdd.n323 gnd 0.010589f
C1428 vdd.n324 gnd 0.008523f
C1429 vdd.n325 gnd 0.008523f
C1430 vdd.n326 gnd 0.010589f
C1431 vdd.n327 gnd 0.010589f
C1432 vdd.n328 gnd 0.77371f
C1433 vdd.n329 gnd 0.010589f
C1434 vdd.n330 gnd 0.010589f
C1435 vdd.n331 gnd 0.010589f
C1436 vdd.n332 gnd 0.838637f
C1437 vdd.n333 gnd 0.010589f
C1438 vdd.n334 gnd 0.010589f
C1439 vdd.n335 gnd 0.010589f
C1440 vdd.n336 gnd 0.010589f
C1441 vdd.n337 gnd 0.008523f
C1442 vdd.n338 gnd 0.010589f
C1443 vdd.t58 gnd 0.541056f
C1444 vdd.n339 gnd 0.010589f
C1445 vdd.n340 gnd 0.010589f
C1446 vdd.n341 gnd 0.010589f
C1447 vdd.t84 gnd 0.541056f
C1448 vdd.n342 gnd 0.010589f
C1449 vdd.n343 gnd 0.010589f
C1450 vdd.n344 gnd 0.010589f
C1451 vdd.n345 gnd 0.010589f
C1452 vdd.n346 gnd 0.010589f
C1453 vdd.n347 gnd 0.008523f
C1454 vdd.n348 gnd 0.010589f
C1455 vdd.n349 gnd 0.611393f
C1456 vdd.n350 gnd 0.010589f
C1457 vdd.n351 gnd 0.010589f
C1458 vdd.n352 gnd 0.010589f
C1459 vdd.t35 gnd 0.541056f
C1460 vdd.n353 gnd 0.010589f
C1461 vdd.n354 gnd 0.010589f
C1462 vdd.n355 gnd 0.010589f
C1463 vdd.n356 gnd 0.010589f
C1464 vdd.n357 gnd 0.010589f
C1465 vdd.n358 gnd 0.008523f
C1466 vdd.n359 gnd 0.010589f
C1467 vdd.t41 gnd 0.541056f
C1468 vdd.n360 gnd 0.010589f
C1469 vdd.n361 gnd 0.010589f
C1470 vdd.n362 gnd 0.010589f
C1471 vdd.n363 gnd 0.914385f
C1472 vdd.n364 gnd 0.010589f
C1473 vdd.n365 gnd 0.010589f
C1474 vdd.n366 gnd 0.010589f
C1475 vdd.n367 gnd 0.010589f
C1476 vdd.n368 gnd 0.010589f
C1477 vdd.n369 gnd 0.007074f
C1478 vdd.n370 gnd 0.024113f
C1479 vdd.t173 gnd 0.541056f
C1480 vdd.n371 gnd 0.010589f
C1481 vdd.n372 gnd 0.024113f
C1482 vdd.n404 gnd 0.010589f
C1483 vdd.t175 gnd 0.130268f
C1484 vdd.t174 gnd 0.139221f
C1485 vdd.t172 gnd 0.170129f
C1486 vdd.n405 gnd 0.218081f
C1487 vdd.n406 gnd 0.18408f
C1488 vdd.n407 gnd 0.013977f
C1489 vdd.n408 gnd 0.010589f
C1490 vdd.n409 gnd 0.008523f
C1491 vdd.n410 gnd 0.010589f
C1492 vdd.n411 gnd 0.008523f
C1493 vdd.n412 gnd 0.010589f
C1494 vdd.n413 gnd 0.008523f
C1495 vdd.n414 gnd 0.010589f
C1496 vdd.n415 gnd 0.008523f
C1497 vdd.n416 gnd 0.010589f
C1498 vdd.n417 gnd 0.008523f
C1499 vdd.n418 gnd 0.010589f
C1500 vdd.t230 gnd 0.130268f
C1501 vdd.t229 gnd 0.139221f
C1502 vdd.t228 gnd 0.170129f
C1503 vdd.n419 gnd 0.218081f
C1504 vdd.n420 gnd 0.18408f
C1505 vdd.n421 gnd 0.008523f
C1506 vdd.n422 gnd 0.010589f
C1507 vdd.n423 gnd 0.008523f
C1508 vdd.n424 gnd 0.010589f
C1509 vdd.n425 gnd 0.008523f
C1510 vdd.n426 gnd 0.010589f
C1511 vdd.n427 gnd 0.008523f
C1512 vdd.n428 gnd 0.010589f
C1513 vdd.n429 gnd 0.008523f
C1514 vdd.n430 gnd 0.010589f
C1515 vdd.t236 gnd 0.130268f
C1516 vdd.t235 gnd 0.139221f
C1517 vdd.t234 gnd 0.170129f
C1518 vdd.n431 gnd 0.218081f
C1519 vdd.n432 gnd 0.18408f
C1520 vdd.n433 gnd 0.018238f
C1521 vdd.n434 gnd 0.010589f
C1522 vdd.n435 gnd 0.008523f
C1523 vdd.n436 gnd 0.010589f
C1524 vdd.n437 gnd 0.008523f
C1525 vdd.n438 gnd 0.010589f
C1526 vdd.n439 gnd 0.008523f
C1527 vdd.n440 gnd 0.010589f
C1528 vdd.n441 gnd 0.008523f
C1529 vdd.n442 gnd 0.010589f
C1530 vdd.n443 gnd 0.024113f
C1531 vdd.n444 gnd 0.024278f
C1532 vdd.n445 gnd 0.024278f
C1533 vdd.n446 gnd 0.007074f
C1534 vdd.n447 gnd 0.008523f
C1535 vdd.n448 gnd 0.010589f
C1536 vdd.n449 gnd 0.010589f
C1537 vdd.n450 gnd 0.008523f
C1538 vdd.n451 gnd 0.010589f
C1539 vdd.n452 gnd 0.010589f
C1540 vdd.n453 gnd 0.010589f
C1541 vdd.n454 gnd 0.010589f
C1542 vdd.n455 gnd 0.010589f
C1543 vdd.n456 gnd 0.008523f
C1544 vdd.n457 gnd 0.008523f
C1545 vdd.n458 gnd 0.010589f
C1546 vdd.n459 gnd 0.010589f
C1547 vdd.n460 gnd 0.008523f
C1548 vdd.n461 gnd 0.010589f
C1549 vdd.n462 gnd 0.010589f
C1550 vdd.n463 gnd 0.010589f
C1551 vdd.n464 gnd 0.010589f
C1552 vdd.n465 gnd 0.010589f
C1553 vdd.n466 gnd 0.008523f
C1554 vdd.n467 gnd 0.008523f
C1555 vdd.n468 gnd 0.010589f
C1556 vdd.n469 gnd 0.010589f
C1557 vdd.n470 gnd 0.008523f
C1558 vdd.n471 gnd 0.010589f
C1559 vdd.n472 gnd 0.010589f
C1560 vdd.n473 gnd 0.010589f
C1561 vdd.n474 gnd 0.010589f
C1562 vdd.n475 gnd 0.010589f
C1563 vdd.n476 gnd 0.008523f
C1564 vdd.n477 gnd 0.008523f
C1565 vdd.n478 gnd 0.010589f
C1566 vdd.n479 gnd 0.010589f
C1567 vdd.n480 gnd 0.008523f
C1568 vdd.n481 gnd 0.010589f
C1569 vdd.n482 gnd 0.010589f
C1570 vdd.n483 gnd 0.010589f
C1571 vdd.n484 gnd 0.010589f
C1572 vdd.n485 gnd 0.010589f
C1573 vdd.n486 gnd 0.008523f
C1574 vdd.n487 gnd 0.008523f
C1575 vdd.n488 gnd 0.010589f
C1576 vdd.n489 gnd 0.010589f
C1577 vdd.n490 gnd 0.007116f
C1578 vdd.n491 gnd 0.010589f
C1579 vdd.n492 gnd 0.010589f
C1580 vdd.n493 gnd 0.010589f
C1581 vdd.n494 gnd 0.010589f
C1582 vdd.n495 gnd 0.010589f
C1583 vdd.n496 gnd 0.007116f
C1584 vdd.n497 gnd 0.008523f
C1585 vdd.n498 gnd 0.010589f
C1586 vdd.n499 gnd 0.010589f
C1587 vdd.n500 gnd 0.008523f
C1588 vdd.n501 gnd 0.010589f
C1589 vdd.n502 gnd 0.010589f
C1590 vdd.n503 gnd 0.010589f
C1591 vdd.n504 gnd 0.010589f
C1592 vdd.n505 gnd 0.010589f
C1593 vdd.n506 gnd 0.008523f
C1594 vdd.n507 gnd 0.008523f
C1595 vdd.n508 gnd 0.010589f
C1596 vdd.n509 gnd 0.010589f
C1597 vdd.n510 gnd 0.008523f
C1598 vdd.n511 gnd 0.010589f
C1599 vdd.n512 gnd 0.010589f
C1600 vdd.n513 gnd 0.010589f
C1601 vdd.n514 gnd 0.010589f
C1602 vdd.n515 gnd 0.010589f
C1603 vdd.n516 gnd 0.008523f
C1604 vdd.n517 gnd 0.008523f
C1605 vdd.n518 gnd 0.010589f
C1606 vdd.n519 gnd 0.010589f
C1607 vdd.n520 gnd 0.008523f
C1608 vdd.n521 gnd 0.010589f
C1609 vdd.n522 gnd 0.010589f
C1610 vdd.n523 gnd 0.010589f
C1611 vdd.n524 gnd 0.010589f
C1612 vdd.n525 gnd 0.010589f
C1613 vdd.n526 gnd 0.008523f
C1614 vdd.n527 gnd 0.008523f
C1615 vdd.n528 gnd 0.010589f
C1616 vdd.n529 gnd 0.010589f
C1617 vdd.n530 gnd 0.008523f
C1618 vdd.n531 gnd 0.010589f
C1619 vdd.n532 gnd 0.010589f
C1620 vdd.n533 gnd 0.010589f
C1621 vdd.n534 gnd 0.010589f
C1622 vdd.n535 gnd 0.010589f
C1623 vdd.n536 gnd 0.008523f
C1624 vdd.n537 gnd 0.008523f
C1625 vdd.n538 gnd 0.010589f
C1626 vdd.n539 gnd 0.010589f
C1627 vdd.n540 gnd 0.008523f
C1628 vdd.n541 gnd 0.010589f
C1629 vdd.n542 gnd 0.010589f
C1630 vdd.n543 gnd 0.010589f
C1631 vdd.n544 gnd 0.010589f
C1632 vdd.n545 gnd 0.010589f
C1633 vdd.n546 gnd 0.005795f
C1634 vdd.n547 gnd 0.018238f
C1635 vdd.n548 gnd 0.010589f
C1636 vdd.n549 gnd 0.010589f
C1637 vdd.n550 gnd 0.008437f
C1638 vdd.n551 gnd 0.010589f
C1639 vdd.n552 gnd 0.010589f
C1640 vdd.n553 gnd 0.010589f
C1641 vdd.n554 gnd 0.010589f
C1642 vdd.n555 gnd 0.010589f
C1643 vdd.n556 gnd 0.008523f
C1644 vdd.n557 gnd 0.008523f
C1645 vdd.n558 gnd 0.010589f
C1646 vdd.n559 gnd 0.010589f
C1647 vdd.n560 gnd 0.008523f
C1648 vdd.n561 gnd 0.010589f
C1649 vdd.n562 gnd 0.010589f
C1650 vdd.n563 gnd 0.010589f
C1651 vdd.n564 gnd 0.010589f
C1652 vdd.n565 gnd 0.010589f
C1653 vdd.n566 gnd 0.008523f
C1654 vdd.n567 gnd 0.008523f
C1655 vdd.n568 gnd 0.010589f
C1656 vdd.n569 gnd 0.010589f
C1657 vdd.n570 gnd 0.008523f
C1658 vdd.n571 gnd 0.010589f
C1659 vdd.n572 gnd 0.010589f
C1660 vdd.n573 gnd 0.010589f
C1661 vdd.n574 gnd 0.010589f
C1662 vdd.n575 gnd 0.010589f
C1663 vdd.n576 gnd 0.008523f
C1664 vdd.n577 gnd 0.008523f
C1665 vdd.n578 gnd 0.010589f
C1666 vdd.n579 gnd 0.010589f
C1667 vdd.n580 gnd 0.008523f
C1668 vdd.n581 gnd 0.010589f
C1669 vdd.n582 gnd 0.010589f
C1670 vdd.n583 gnd 0.010589f
C1671 vdd.n584 gnd 0.010589f
C1672 vdd.n585 gnd 0.010589f
C1673 vdd.n586 gnd 0.008523f
C1674 vdd.n587 gnd 0.008523f
C1675 vdd.n588 gnd 0.010589f
C1676 vdd.n589 gnd 0.010589f
C1677 vdd.n590 gnd 0.008523f
C1678 vdd.n591 gnd 0.010589f
C1679 vdd.n592 gnd 0.010589f
C1680 vdd.n593 gnd 0.010589f
C1681 vdd.n594 gnd 0.010589f
C1682 vdd.n595 gnd 0.010589f
C1683 vdd.n596 gnd 0.008523f
C1684 vdd.n597 gnd 0.010589f
C1685 vdd.n598 gnd 0.008523f
C1686 vdd.n599 gnd 0.004474f
C1687 vdd.n600 gnd 0.010589f
C1688 vdd.n601 gnd 0.010589f
C1689 vdd.n602 gnd 0.008523f
C1690 vdd.n603 gnd 0.010589f
C1691 vdd.n604 gnd 0.008523f
C1692 vdd.n605 gnd 0.010589f
C1693 vdd.n606 gnd 0.008523f
C1694 vdd.n607 gnd 0.010589f
C1695 vdd.n608 gnd 0.008523f
C1696 vdd.n609 gnd 0.010589f
C1697 vdd.n610 gnd 0.008523f
C1698 vdd.n611 gnd 0.010589f
C1699 vdd.n612 gnd 0.010589f
C1700 vdd.n613 gnd 0.589751f
C1701 vdd.t63 gnd 0.541056f
C1702 vdd.n614 gnd 0.010589f
C1703 vdd.n615 gnd 0.008523f
C1704 vdd.n616 gnd 0.010589f
C1705 vdd.n617 gnd 0.008523f
C1706 vdd.n618 gnd 0.010589f
C1707 vdd.t108 gnd 0.541056f
C1708 vdd.n619 gnd 0.010589f
C1709 vdd.n620 gnd 0.008523f
C1710 vdd.n621 gnd 0.010589f
C1711 vdd.n622 gnd 0.008523f
C1712 vdd.n623 gnd 0.010589f
C1713 vdd.t55 gnd 0.541056f
C1714 vdd.n624 gnd 0.67632f
C1715 vdd.n625 gnd 0.010589f
C1716 vdd.n626 gnd 0.008523f
C1717 vdd.n627 gnd 0.010589f
C1718 vdd.n628 gnd 0.008523f
C1719 vdd.n629 gnd 0.010589f
C1720 vdd.t25 gnd 0.541056f
C1721 vdd.n630 gnd 0.010589f
C1722 vdd.n631 gnd 0.008523f
C1723 vdd.n632 gnd 0.010589f
C1724 vdd.n633 gnd 0.008523f
C1725 vdd.n634 gnd 0.010589f
C1726 vdd.n635 gnd 0.752068f
C1727 vdd.n636 gnd 0.898153f
C1728 vdd.t82 gnd 0.541056f
C1729 vdd.n637 gnd 0.010589f
C1730 vdd.n638 gnd 0.008523f
C1731 vdd.n639 gnd 0.010589f
C1732 vdd.n640 gnd 0.008523f
C1733 vdd.n641 gnd 0.010589f
C1734 vdd.n642 gnd 0.568109f
C1735 vdd.n643 gnd 0.010589f
C1736 vdd.n644 gnd 0.008523f
C1737 vdd.n645 gnd 0.010589f
C1738 vdd.n646 gnd 0.008523f
C1739 vdd.n647 gnd 0.010589f
C1740 vdd.n648 gnd 1.08211f
C1741 vdd.t21 gnd 0.541056f
C1742 vdd.n649 gnd 0.010589f
C1743 vdd.n650 gnd 0.008523f
C1744 vdd.n651 gnd 0.010589f
C1745 vdd.n652 gnd 0.008523f
C1746 vdd.n653 gnd 0.010589f
C1747 vdd.t165 gnd 0.541056f
C1748 vdd.n654 gnd 0.010589f
C1749 vdd.n655 gnd 0.008523f
C1750 vdd.n656 gnd 0.024278f
C1751 vdd.n657 gnd 0.024278f
C1752 vdd.n658 gnd 7.650529f
C1753 vdd.n659 gnd 0.600572f
C1754 vdd.n660 gnd 0.024278f
C1755 vdd.n661 gnd 0.009106f
C1756 vdd.n662 gnd 0.008523f
C1757 vdd.n667 gnd 0.006777f
C1758 vdd.n668 gnd 0.008523f
C1759 vdd.n669 gnd 0.010589f
C1760 vdd.n670 gnd 0.010589f
C1761 vdd.n671 gnd 0.010589f
C1762 vdd.n672 gnd 0.010589f
C1763 vdd.n673 gnd 0.010589f
C1764 vdd.n674 gnd 0.008523f
C1765 vdd.n675 gnd 0.010589f
C1766 vdd.n676 gnd 0.010589f
C1767 vdd.n677 gnd 0.010589f
C1768 vdd.n678 gnd 0.010589f
C1769 vdd.n679 gnd 0.010589f
C1770 vdd.n680 gnd 0.008523f
C1771 vdd.n681 gnd 0.010589f
C1772 vdd.n682 gnd 0.010589f
C1773 vdd.n683 gnd 0.010589f
C1774 vdd.n684 gnd 0.010589f
C1775 vdd.n685 gnd 0.010589f
C1776 vdd.t177 gnd 0.130268f
C1777 vdd.t178 gnd 0.139221f
C1778 vdd.t176 gnd 0.170129f
C1779 vdd.n686 gnd 0.218081f
C1780 vdd.n687 gnd 0.183228f
C1781 vdd.n688 gnd 0.017386f
C1782 vdd.n689 gnd 0.010589f
C1783 vdd.n690 gnd 0.010589f
C1784 vdd.n691 gnd 0.010589f
C1785 vdd.n692 gnd 0.010589f
C1786 vdd.n693 gnd 0.010589f
C1787 vdd.n694 gnd 0.008523f
C1788 vdd.n695 gnd 0.010589f
C1789 vdd.n696 gnd 0.010589f
C1790 vdd.n697 gnd 0.010589f
C1791 vdd.n698 gnd 0.010589f
C1792 vdd.n699 gnd 0.010589f
C1793 vdd.n700 gnd 0.008523f
C1794 vdd.n701 gnd 0.010589f
C1795 vdd.n702 gnd 0.010589f
C1796 vdd.n703 gnd 0.010589f
C1797 vdd.n704 gnd 0.010589f
C1798 vdd.n705 gnd 0.010589f
C1799 vdd.n706 gnd 0.008523f
C1800 vdd.n707 gnd 0.010589f
C1801 vdd.n708 gnd 0.010589f
C1802 vdd.n709 gnd 0.010589f
C1803 vdd.n710 gnd 0.010589f
C1804 vdd.n711 gnd 0.010589f
C1805 vdd.n712 gnd 0.008523f
C1806 vdd.n713 gnd 0.010589f
C1807 vdd.n714 gnd 0.010589f
C1808 vdd.n715 gnd 0.010589f
C1809 vdd.n716 gnd 0.010589f
C1810 vdd.n717 gnd 0.010589f
C1811 vdd.n718 gnd 0.008523f
C1812 vdd.n719 gnd 0.010589f
C1813 vdd.n720 gnd 0.010589f
C1814 vdd.n721 gnd 0.010589f
C1815 vdd.n722 gnd 0.008437f
C1816 vdd.t166 gnd 0.130268f
C1817 vdd.t167 gnd 0.139221f
C1818 vdd.t164 gnd 0.170129f
C1819 vdd.n723 gnd 0.218081f
C1820 vdd.n724 gnd 0.183228f
C1821 vdd.n725 gnd 0.010589f
C1822 vdd.n726 gnd 0.008523f
C1823 vdd.n728 gnd 0.010589f
C1824 vdd.n730 gnd 0.010589f
C1825 vdd.n731 gnd 0.010589f
C1826 vdd.n732 gnd 0.008523f
C1827 vdd.n733 gnd 0.010589f
C1828 vdd.n734 gnd 0.010589f
C1829 vdd.n735 gnd 0.010589f
C1830 vdd.n736 gnd 0.010589f
C1831 vdd.n737 gnd 0.010589f
C1832 vdd.n738 gnd 0.008523f
C1833 vdd.n739 gnd 0.010589f
C1834 vdd.n740 gnd 0.010589f
C1835 vdd.n741 gnd 0.010589f
C1836 vdd.n742 gnd 0.010589f
C1837 vdd.n743 gnd 0.010589f
C1838 vdd.n744 gnd 0.008523f
C1839 vdd.n745 gnd 0.010589f
C1840 vdd.n746 gnd 0.010589f
C1841 vdd.n747 gnd 0.010589f
C1842 vdd.n748 gnd 0.006777f
C1843 vdd.n753 gnd 0.0072f
C1844 vdd.n754 gnd 0.0072f
C1845 vdd.n755 gnd 0.0072f
C1846 vdd.n756 gnd 7.45575f
C1847 vdd.n757 gnd 0.0072f
C1848 vdd.n758 gnd 0.0072f
C1849 vdd.n759 gnd 0.0072f
C1850 vdd.n761 gnd 0.0072f
C1851 vdd.n762 gnd 0.0072f
C1852 vdd.n764 gnd 0.0072f
C1853 vdd.n765 gnd 0.005241f
C1854 vdd.n767 gnd 0.0072f
C1855 vdd.t213 gnd 0.290963f
C1856 vdd.t212 gnd 0.297837f
C1857 vdd.t211 gnd 0.189952f
C1858 vdd.n768 gnd 0.102658f
C1859 vdd.n769 gnd 0.058231f
C1860 vdd.n770 gnd 0.01029f
C1861 vdd.n771 gnd 0.016828f
C1862 vdd.n773 gnd 0.0072f
C1863 vdd.n774 gnd 0.735836f
C1864 vdd.n775 gnd 0.015952f
C1865 vdd.n776 gnd 0.015952f
C1866 vdd.n777 gnd 0.0072f
C1867 vdd.n778 gnd 0.017085f
C1868 vdd.n779 gnd 0.0072f
C1869 vdd.n780 gnd 0.0072f
C1870 vdd.n781 gnd 0.0072f
C1871 vdd.n782 gnd 0.0072f
C1872 vdd.n783 gnd 0.0072f
C1873 vdd.n785 gnd 0.0072f
C1874 vdd.n786 gnd 0.0072f
C1875 vdd.n788 gnd 0.0072f
C1876 vdd.n789 gnd 0.0072f
C1877 vdd.n791 gnd 0.0072f
C1878 vdd.n792 gnd 0.0072f
C1879 vdd.n794 gnd 0.0072f
C1880 vdd.n795 gnd 0.0072f
C1881 vdd.n797 gnd 0.0072f
C1882 vdd.n798 gnd 0.0072f
C1883 vdd.n800 gnd 0.0072f
C1884 vdd.n801 gnd 0.005241f
C1885 vdd.n803 gnd 0.0072f
C1886 vdd.t206 gnd 0.290963f
C1887 vdd.t205 gnd 0.297837f
C1888 vdd.t203 gnd 0.189952f
C1889 vdd.n804 gnd 0.102658f
C1890 vdd.n805 gnd 0.058231f
C1891 vdd.n806 gnd 0.01029f
C1892 vdd.n807 gnd 0.0072f
C1893 vdd.n808 gnd 0.0072f
C1894 vdd.t204 gnd 0.367918f
C1895 vdd.n809 gnd 0.0072f
C1896 vdd.n810 gnd 0.0072f
C1897 vdd.n811 gnd 0.0072f
C1898 vdd.n812 gnd 0.0072f
C1899 vdd.n813 gnd 0.0072f
C1900 vdd.n814 gnd 0.735836f
C1901 vdd.n815 gnd 0.0072f
C1902 vdd.n816 gnd 0.0072f
C1903 vdd.n817 gnd 0.643857f
C1904 vdd.n818 gnd 0.0072f
C1905 vdd.n819 gnd 0.0072f
C1906 vdd.n820 gnd 0.006353f
C1907 vdd.n821 gnd 0.0072f
C1908 vdd.n822 gnd 0.649267f
C1909 vdd.n823 gnd 0.0072f
C1910 vdd.n824 gnd 0.0072f
C1911 vdd.n825 gnd 0.0072f
C1912 vdd.n826 gnd 0.0072f
C1913 vdd.n827 gnd 0.0072f
C1914 vdd.n828 gnd 0.735836f
C1915 vdd.n829 gnd 0.0072f
C1916 vdd.n830 gnd 0.0072f
C1917 vdd.t187 gnd 0.330044f
C1918 vdd.t14 gnd 0.086569f
C1919 vdd.n831 gnd 0.0072f
C1920 vdd.n832 gnd 0.0072f
C1921 vdd.n833 gnd 0.0072f
C1922 vdd.t2 gnd 0.367918f
C1923 vdd.n834 gnd 0.0072f
C1924 vdd.n835 gnd 0.0072f
C1925 vdd.n836 gnd 0.0072f
C1926 vdd.n837 gnd 0.0072f
C1927 vdd.n838 gnd 0.0072f
C1928 vdd.t11 gnd 0.367918f
C1929 vdd.n839 gnd 0.0072f
C1930 vdd.n840 gnd 0.0072f
C1931 vdd.n841 gnd 0.611393f
C1932 vdd.n842 gnd 0.0072f
C1933 vdd.n843 gnd 0.0072f
C1934 vdd.n844 gnd 0.0072f
C1935 vdd.n845 gnd 0.449076f
C1936 vdd.n846 gnd 0.0072f
C1937 vdd.n847 gnd 0.0072f
C1938 vdd.t260 gnd 0.367918f
C1939 vdd.n848 gnd 0.0072f
C1940 vdd.n849 gnd 0.0072f
C1941 vdd.n850 gnd 0.0072f
C1942 vdd.n851 gnd 0.611393f
C1943 vdd.n852 gnd 0.0072f
C1944 vdd.n853 gnd 0.0072f
C1945 vdd.t10 gnd 0.313812f
C1946 vdd.t155 gnd 0.28676f
C1947 vdd.n854 gnd 0.0072f
C1948 vdd.n855 gnd 0.0072f
C1949 vdd.n856 gnd 0.0072f
C1950 vdd.t8 gnd 0.367918f
C1951 vdd.n857 gnd 0.0072f
C1952 vdd.n858 gnd 0.0072f
C1953 vdd.t17 gnd 0.367918f
C1954 vdd.n859 gnd 0.0072f
C1955 vdd.n860 gnd 0.0072f
C1956 vdd.n861 gnd 0.0072f
C1957 vdd.t161 gnd 0.270528f
C1958 vdd.n862 gnd 0.0072f
C1959 vdd.n863 gnd 0.0072f
C1960 vdd.n864 gnd 0.627625f
C1961 vdd.n865 gnd 0.0072f
C1962 vdd.n866 gnd 0.0072f
C1963 vdd.n867 gnd 0.0072f
C1964 vdd.n868 gnd 0.735836f
C1965 vdd.n869 gnd 0.0072f
C1966 vdd.n870 gnd 0.0072f
C1967 vdd.t147 gnd 0.330044f
C1968 vdd.n871 gnd 0.465308f
C1969 vdd.n872 gnd 0.0072f
C1970 vdd.n873 gnd 0.0072f
C1971 vdd.n874 gnd 0.0072f
C1972 vdd.t256 gnd 0.367918f
C1973 vdd.n875 gnd 0.0072f
C1974 vdd.n876 gnd 0.0072f
C1975 vdd.n877 gnd 0.0072f
C1976 vdd.n878 gnd 0.0072f
C1977 vdd.n879 gnd 0.0072f
C1978 vdd.t157 gnd 0.735836f
C1979 vdd.n880 gnd 0.0072f
C1980 vdd.n881 gnd 0.0072f
C1981 vdd.t208 gnd 0.367918f
C1982 vdd.n882 gnd 0.0072f
C1983 vdd.n883 gnd 0.017085f
C1984 vdd.n884 gnd 0.017085f
C1985 vdd.t159 gnd 0.692552f
C1986 vdd.n885 gnd 0.015952f
C1987 vdd.n886 gnd 0.015952f
C1988 vdd.n887 gnd 0.017085f
C1989 vdd.n888 gnd 0.0072f
C1990 vdd.n889 gnd 0.0072f
C1991 vdd.t6 gnd 0.692552f
C1992 vdd.n907 gnd 0.017085f
C1993 vdd.n925 gnd 0.015952f
C1994 vdd.n926 gnd 0.0072f
C1995 vdd.n927 gnd 0.015952f
C1996 vdd.t227 gnd 0.290963f
C1997 vdd.t226 gnd 0.297837f
C1998 vdd.t225 gnd 0.189952f
C1999 vdd.n928 gnd 0.102658f
C2000 vdd.n929 gnd 0.058231f
C2001 vdd.n930 gnd 0.016828f
C2002 vdd.n931 gnd 0.0072f
C2003 vdd.t15 gnd 0.735836f
C2004 vdd.n932 gnd 0.015952f
C2005 vdd.n933 gnd 0.0072f
C2006 vdd.n934 gnd 0.017085f
C2007 vdd.n935 gnd 0.0072f
C2008 vdd.t202 gnd 0.290963f
C2009 vdd.t201 gnd 0.297837f
C2010 vdd.t199 gnd 0.189952f
C2011 vdd.n936 gnd 0.102658f
C2012 vdd.n937 gnd 0.058231f
C2013 vdd.n938 gnd 0.01029f
C2014 vdd.n939 gnd 0.0072f
C2015 vdd.n940 gnd 0.0072f
C2016 vdd.t200 gnd 0.367918f
C2017 vdd.n941 gnd 0.0072f
C2018 vdd.n942 gnd 0.0072f
C2019 vdd.n943 gnd 0.0072f
C2020 vdd.n944 gnd 0.0072f
C2021 vdd.n945 gnd 0.0072f
C2022 vdd.n946 gnd 0.0072f
C2023 vdd.n947 gnd 0.735836f
C2024 vdd.n948 gnd 0.0072f
C2025 vdd.n949 gnd 0.0072f
C2026 vdd.t258 gnd 0.367918f
C2027 vdd.n950 gnd 0.0072f
C2028 vdd.n951 gnd 0.0072f
C2029 vdd.n952 gnd 0.0072f
C2030 vdd.n953 gnd 0.0072f
C2031 vdd.n954 gnd 0.465308f
C2032 vdd.n955 gnd 0.0072f
C2033 vdd.n956 gnd 0.0072f
C2034 vdd.n957 gnd 0.0072f
C2035 vdd.n958 gnd 0.0072f
C2036 vdd.n959 gnd 0.0072f
C2037 vdd.n960 gnd 0.627625f
C2038 vdd.n961 gnd 0.0072f
C2039 vdd.n962 gnd 0.0072f
C2040 vdd.t262 gnd 0.330044f
C2041 vdd.t150 gnd 0.270528f
C2042 vdd.n963 gnd 0.0072f
C2043 vdd.n964 gnd 0.0072f
C2044 vdd.n965 gnd 0.0072f
C2045 vdd.t149 gnd 0.367918f
C2046 vdd.n966 gnd 0.0072f
C2047 vdd.n967 gnd 0.0072f
C2048 vdd.t153 gnd 0.367918f
C2049 vdd.n968 gnd 0.0072f
C2050 vdd.n969 gnd 0.0072f
C2051 vdd.n970 gnd 0.0072f
C2052 vdd.t0 gnd 0.28676f
C2053 vdd.n971 gnd 0.0072f
C2054 vdd.n972 gnd 0.0072f
C2055 vdd.n973 gnd 0.611393f
C2056 vdd.n974 gnd 0.0072f
C2057 vdd.n975 gnd 0.0072f
C2058 vdd.n976 gnd 0.0072f
C2059 vdd.t4 gnd 0.367918f
C2060 vdd.n977 gnd 0.0072f
C2061 vdd.n978 gnd 0.0072f
C2062 vdd.t3 gnd 0.313812f
C2063 vdd.n979 gnd 0.449076f
C2064 vdd.n980 gnd 0.0072f
C2065 vdd.n981 gnd 0.0072f
C2066 vdd.n982 gnd 0.0072f
C2067 vdd.n983 gnd 0.611393f
C2068 vdd.n984 gnd 0.0072f
C2069 vdd.n985 gnd 0.0072f
C2070 vdd.t18 gnd 0.367918f
C2071 vdd.n986 gnd 0.0072f
C2072 vdd.n987 gnd 0.0072f
C2073 vdd.n988 gnd 0.0072f
C2074 vdd.n989 gnd 0.735836f
C2075 vdd.n990 gnd 0.0072f
C2076 vdd.n991 gnd 0.0072f
C2077 vdd.t162 gnd 0.367918f
C2078 vdd.n992 gnd 0.0072f
C2079 vdd.n993 gnd 0.0072f
C2080 vdd.n994 gnd 0.0072f
C2081 vdd.t163 gnd 0.086569f
C2082 vdd.n995 gnd 0.0072f
C2083 vdd.n996 gnd 0.0072f
C2084 vdd.n997 gnd 0.0072f
C2085 vdd.t220 gnd 0.297837f
C2086 vdd.t218 gnd 0.189952f
C2087 vdd.t221 gnd 0.297837f
C2088 vdd.n998 gnd 0.167396f
C2089 vdd.n999 gnd 0.0072f
C2090 vdd.n1000 gnd 0.0072f
C2091 vdd.n1001 gnd 0.735836f
C2092 vdd.n1002 gnd 0.0072f
C2093 vdd.n1003 gnd 0.0072f
C2094 vdd.t219 gnd 0.330044f
C2095 vdd.n1004 gnd 0.649267f
C2096 vdd.n1005 gnd 0.0072f
C2097 vdd.n1006 gnd 0.0072f
C2098 vdd.n1007 gnd 0.0072f
C2099 vdd.n1008 gnd 0.643857f
C2100 vdd.n1009 gnd 0.0072f
C2101 vdd.n1010 gnd 0.0072f
C2102 vdd.n1011 gnd 0.0072f
C2103 vdd.n1012 gnd 0.0072f
C2104 vdd.n1013 gnd 0.0072f
C2105 vdd.n1014 gnd 0.735836f
C2106 vdd.n1015 gnd 0.0072f
C2107 vdd.n1016 gnd 0.0072f
C2108 vdd.t215 gnd 0.367918f
C2109 vdd.n1017 gnd 0.0072f
C2110 vdd.n1018 gnd 0.017085f
C2111 vdd.n1019 gnd 0.017085f
C2112 vdd.n1020 gnd 7.45575f
C2113 vdd.n1021 gnd 0.015952f
C2114 vdd.n1022 gnd 0.015952f
C2115 vdd.n1023 gnd 0.017085f
C2116 vdd.n1024 gnd 0.0072f
C2117 vdd.n1025 gnd 0.0072f
C2118 vdd.n1026 gnd 0.0072f
C2119 vdd.n1027 gnd 0.0072f
C2120 vdd.n1028 gnd 0.0072f
C2121 vdd.n1029 gnd 0.0072f
C2122 vdd.n1030 gnd 0.0072f
C2123 vdd.n1031 gnd 0.0072f
C2124 vdd.n1033 gnd 0.0072f
C2125 vdd.n1034 gnd 0.0072f
C2126 vdd.n1035 gnd 0.006777f
C2127 vdd.n1038 gnd 0.024278f
C2128 vdd.n1039 gnd 0.008523f
C2129 vdd.n1040 gnd 0.010589f
C2130 vdd.n1042 gnd 0.010589f
C2131 vdd.n1043 gnd 0.007074f
C2132 vdd.n1044 gnd 0.600572f
C2133 vdd.n1045 gnd 7.650529f
C2134 vdd.n1046 gnd 0.010589f
C2135 vdd.n1047 gnd 0.024278f
C2136 vdd.n1048 gnd 0.008523f
C2137 vdd.n1049 gnd 0.010589f
C2138 vdd.n1050 gnd 0.008523f
C2139 vdd.n1051 gnd 0.010589f
C2140 vdd.n1052 gnd 1.08211f
C2141 vdd.n1053 gnd 0.010589f
C2142 vdd.n1054 gnd 0.008523f
C2143 vdd.n1055 gnd 0.008523f
C2144 vdd.n1056 gnd 0.010589f
C2145 vdd.n1057 gnd 0.008523f
C2146 vdd.n1058 gnd 0.010589f
C2147 vdd.t19 gnd 0.541056f
C2148 vdd.n1059 gnd 0.010589f
C2149 vdd.n1060 gnd 0.008523f
C2150 vdd.n1061 gnd 0.010589f
C2151 vdd.n1062 gnd 0.008523f
C2152 vdd.n1063 gnd 0.010589f
C2153 vdd.t126 gnd 0.541056f
C2154 vdd.n1064 gnd 0.010589f
C2155 vdd.n1065 gnd 0.008523f
C2156 vdd.n1066 gnd 0.010589f
C2157 vdd.n1067 gnd 0.008523f
C2158 vdd.n1068 gnd 0.010589f
C2159 vdd.t33 gnd 0.541056f
C2160 vdd.n1069 gnd 0.752068f
C2161 vdd.n1070 gnd 0.010589f
C2162 vdd.n1071 gnd 0.008523f
C2163 vdd.n1072 gnd 0.010589f
C2164 vdd.n1073 gnd 0.008523f
C2165 vdd.n1074 gnd 0.010589f
C2166 vdd.n1075 gnd 0.860279f
C2167 vdd.n1076 gnd 0.010589f
C2168 vdd.n1077 gnd 0.008523f
C2169 vdd.n1078 gnd 0.010589f
C2170 vdd.n1079 gnd 0.008523f
C2171 vdd.n1080 gnd 0.010589f
C2172 vdd.n1081 gnd 0.67632f
C2173 vdd.t53 gnd 0.541056f
C2174 vdd.n1082 gnd 0.010589f
C2175 vdd.n1083 gnd 0.008523f
C2176 vdd.n1084 gnd 0.010589f
C2177 vdd.n1085 gnd 0.008523f
C2178 vdd.n1086 gnd 0.010589f
C2179 vdd.t74 gnd 0.541056f
C2180 vdd.n1087 gnd 0.010589f
C2181 vdd.n1088 gnd 0.008523f
C2182 vdd.n1089 gnd 0.010589f
C2183 vdd.n1090 gnd 0.008523f
C2184 vdd.n1091 gnd 0.010589f
C2185 vdd.t104 gnd 0.541056f
C2186 vdd.n1092 gnd 0.589751f
C2187 vdd.n1093 gnd 0.010589f
C2188 vdd.n1094 gnd 0.008523f
C2189 vdd.n1095 gnd 0.010589f
C2190 vdd.n1096 gnd 0.008523f
C2191 vdd.n1097 gnd 0.010589f
C2192 vdd.t95 gnd 0.541056f
C2193 vdd.n1098 gnd 0.010589f
C2194 vdd.n1099 gnd 0.008523f
C2195 vdd.n1100 gnd 0.010589f
C2196 vdd.n1101 gnd 0.008523f
C2197 vdd.n1102 gnd 0.010589f
C2198 vdd.n1103 gnd 0.838637f
C2199 vdd.n1104 gnd 0.898153f
C2200 vdd.t27 gnd 0.541056f
C2201 vdd.n1105 gnd 0.010589f
C2202 vdd.n1106 gnd 0.008523f
C2203 vdd.n1107 gnd 0.010589f
C2204 vdd.n1108 gnd 0.008523f
C2205 vdd.n1109 gnd 0.010589f
C2206 vdd.n1110 gnd 0.654678f
C2207 vdd.n1111 gnd 0.010589f
C2208 vdd.n1112 gnd 0.008523f
C2209 vdd.n1113 gnd 0.010589f
C2210 vdd.n1114 gnd 0.008523f
C2211 vdd.n1115 gnd 0.010589f
C2212 vdd.t50 gnd 0.541056f
C2213 vdd.t39 gnd 0.541056f
C2214 vdd.n1116 gnd 0.010589f
C2215 vdd.n1117 gnd 0.008523f
C2216 vdd.n1118 gnd 0.010589f
C2217 vdd.n1119 gnd 0.008523f
C2218 vdd.n1120 gnd 0.010589f
C2219 vdd.t90 gnd 0.541056f
C2220 vdd.n1121 gnd 0.010589f
C2221 vdd.n1122 gnd 0.008523f
C2222 vdd.n1123 gnd 0.010589f
C2223 vdd.n1124 gnd 0.008523f
C2224 vdd.n1125 gnd 0.010589f
C2225 vdd.t92 gnd 0.541056f
C2226 vdd.n1126 gnd 0.795352f
C2227 vdd.n1127 gnd 0.010589f
C2228 vdd.n1128 gnd 0.008523f
C2229 vdd.n1129 gnd 0.010589f
C2230 vdd.n1130 gnd 0.008523f
C2231 vdd.n1131 gnd 0.010589f
C2232 vdd.n1132 gnd 1.08211f
C2233 vdd.n1133 gnd 0.010589f
C2234 vdd.n1134 gnd 0.008523f
C2235 vdd.n1135 gnd 0.010589f
C2236 vdd.n1136 gnd 0.008523f
C2237 vdd.n1137 gnd 0.010589f
C2238 vdd.n1138 gnd 0.914385f
C2239 vdd.n1139 gnd 0.010589f
C2240 vdd.n1140 gnd 0.008523f
C2241 vdd.n1141 gnd 0.024113f
C2242 vdd.n1142 gnd 0.007074f
C2243 vdd.n1143 gnd 0.024113f
C2244 vdd.n1144 gnd 1.42839f
C2245 vdd.n1145 gnd 0.024113f
C2246 vdd.n1146 gnd 0.007074f
C2247 vdd.n1147 gnd 0.010589f
C2248 vdd.t170 gnd 0.130268f
C2249 vdd.t171 gnd 0.139221f
C2250 vdd.t168 gnd 0.170129f
C2251 vdd.n1148 gnd 0.218081f
C2252 vdd.n1149 gnd 0.18408f
C2253 vdd.n1150 gnd 0.013977f
C2254 vdd.n1151 gnd 0.010589f
C2255 vdd.n1182 gnd 0.010589f
C2256 vdd.n1183 gnd 0.010589f
C2257 vdd.n1184 gnd 0.024278f
C2258 vdd.n1185 gnd 0.008523f
C2259 vdd.n1186 gnd 0.010589f
C2260 vdd.n1187 gnd 0.010589f
C2261 vdd.n1188 gnd 0.010589f
C2262 vdd.n1189 gnd 0.010589f
C2263 vdd.n1190 gnd 0.008523f
C2264 vdd.n1191 gnd 0.010589f
C2265 vdd.n1192 gnd 0.010589f
C2266 vdd.n1193 gnd 0.010589f
C2267 vdd.n1194 gnd 0.010589f
C2268 vdd.n1195 gnd 0.010589f
C2269 vdd.n1196 gnd 0.008523f
C2270 vdd.n1197 gnd 0.010589f
C2271 vdd.n1198 gnd 0.010589f
C2272 vdd.n1199 gnd 0.010589f
C2273 vdd.n1200 gnd 0.010589f
C2274 vdd.n1201 gnd 0.010589f
C2275 vdd.n1202 gnd 0.008523f
C2276 vdd.n1203 gnd 0.010589f
C2277 vdd.n1204 gnd 0.010589f
C2278 vdd.n1205 gnd 0.010589f
C2279 vdd.n1206 gnd 0.010589f
C2280 vdd.n1207 gnd 0.010589f
C2281 vdd.n1208 gnd 0.007116f
C2282 vdd.n1209 gnd 0.010589f
C2283 vdd.n1210 gnd 0.010589f
C2284 vdd.n1211 gnd 0.010589f
C2285 vdd.n1212 gnd 0.008523f
C2286 vdd.n1213 gnd 0.010589f
C2287 vdd.n1214 gnd 0.010589f
C2288 vdd.n1215 gnd 0.010589f
C2289 vdd.n1216 gnd 0.010589f
C2290 vdd.n1217 gnd 0.010589f
C2291 vdd.n1218 gnd 0.008523f
C2292 vdd.n1219 gnd 0.010589f
C2293 vdd.n1220 gnd 0.010589f
C2294 vdd.n1221 gnd 0.010589f
C2295 vdd.n1222 gnd 0.010589f
C2296 vdd.n1223 gnd 0.010589f
C2297 vdd.n1224 gnd 0.008523f
C2298 vdd.n1225 gnd 0.010589f
C2299 vdd.n1226 gnd 0.010589f
C2300 vdd.n1227 gnd 0.010589f
C2301 vdd.n1228 gnd 0.010589f
C2302 vdd.n1229 gnd 0.010589f
C2303 vdd.n1230 gnd 0.008523f
C2304 vdd.n1231 gnd 0.010589f
C2305 vdd.n1232 gnd 0.010589f
C2306 vdd.n1233 gnd 0.010589f
C2307 vdd.n1234 gnd 0.010589f
C2308 vdd.n1235 gnd 0.010589f
C2309 vdd.n1236 gnd 0.008523f
C2310 vdd.n1237 gnd 0.010589f
C2311 vdd.n1238 gnd 0.010589f
C2312 vdd.n1239 gnd 0.010589f
C2313 vdd.n1240 gnd 0.010589f
C2314 vdd.n1241 gnd 0.008437f
C2315 vdd.n1242 gnd 0.010589f
C2316 vdd.n1243 gnd 0.010589f
C2317 vdd.n1244 gnd 0.010589f
C2318 vdd.n1245 gnd 0.010589f
C2319 vdd.n1246 gnd 0.010589f
C2320 vdd.n1247 gnd 0.008523f
C2321 vdd.n1248 gnd 0.010589f
C2322 vdd.n1249 gnd 0.010589f
C2323 vdd.n1250 gnd 0.010589f
C2324 vdd.n1251 gnd 0.010589f
C2325 vdd.n1252 gnd 0.010589f
C2326 vdd.n1253 gnd 0.008523f
C2327 vdd.n1254 gnd 0.010589f
C2328 vdd.n1255 gnd 0.010589f
C2329 vdd.n1256 gnd 0.010589f
C2330 vdd.n1257 gnd 0.010589f
C2331 vdd.n1258 gnd 0.010589f
C2332 vdd.n1259 gnd 0.008523f
C2333 vdd.n1260 gnd 0.010589f
C2334 vdd.n1261 gnd 0.010589f
C2335 vdd.n1262 gnd 0.010589f
C2336 vdd.n1263 gnd 0.010589f
C2337 vdd.n1264 gnd 0.010589f
C2338 vdd.n1265 gnd 0.008523f
C2339 vdd.n1266 gnd 0.010589f
C2340 vdd.n1267 gnd 0.010589f
C2341 vdd.n1268 gnd 0.010589f
C2342 vdd.n1269 gnd 0.010589f
C2343 vdd.n1270 gnd 0.010589f
C2344 vdd.n1271 gnd 0.004474f
C2345 vdd.n1272 gnd 0.010589f
C2346 vdd.n1273 gnd 0.008523f
C2347 vdd.n1274 gnd 0.008523f
C2348 vdd.n1275 gnd 0.008523f
C2349 vdd.n1276 gnd 0.010589f
C2350 vdd.n1277 gnd 0.010589f
C2351 vdd.n1278 gnd 0.010589f
C2352 vdd.n1279 gnd 0.008523f
C2353 vdd.n1280 gnd 0.008523f
C2354 vdd.n1281 gnd 0.008523f
C2355 vdd.n1282 gnd 0.010589f
C2356 vdd.n1283 gnd 0.010589f
C2357 vdd.n1284 gnd 0.010589f
C2358 vdd.n1285 gnd 0.008523f
C2359 vdd.n1286 gnd 0.008523f
C2360 vdd.n1287 gnd 0.008523f
C2361 vdd.n1288 gnd 0.010589f
C2362 vdd.n1289 gnd 0.010589f
C2363 vdd.n1290 gnd 0.010589f
C2364 vdd.n1291 gnd 0.008523f
C2365 vdd.n1292 gnd 0.008523f
C2366 vdd.n1293 gnd 0.008523f
C2367 vdd.n1294 gnd 0.010589f
C2368 vdd.n1295 gnd 0.010589f
C2369 vdd.n1296 gnd 0.010589f
C2370 vdd.n1297 gnd 0.008523f
C2371 vdd.n1298 gnd 0.008523f
C2372 vdd.n1299 gnd 0.008523f
C2373 vdd.n1300 gnd 0.010589f
C2374 vdd.n1301 gnd 0.010589f
C2375 vdd.n1302 gnd 0.010589f
C2376 vdd.n1303 gnd 0.010589f
C2377 vdd.t184 gnd 0.130268f
C2378 vdd.t185 gnd 0.139221f
C2379 vdd.t183 gnd 0.170129f
C2380 vdd.n1304 gnd 0.218081f
C2381 vdd.n1305 gnd 0.18408f
C2382 vdd.n1306 gnd 0.018238f
C2383 vdd.n1307 gnd 0.005795f
C2384 vdd.n1308 gnd 0.008523f
C2385 vdd.n1309 gnd 0.010589f
C2386 vdd.n1310 gnd 0.010589f
C2387 vdd.n1311 gnd 0.010589f
C2388 vdd.n1312 gnd 0.008523f
C2389 vdd.n1313 gnd 0.008523f
C2390 vdd.n1314 gnd 0.008523f
C2391 vdd.n1315 gnd 0.010589f
C2392 vdd.n1316 gnd 0.010589f
C2393 vdd.n1317 gnd 0.010589f
C2394 vdd.n1318 gnd 0.008523f
C2395 vdd.n1319 gnd 0.008523f
C2396 vdd.n1320 gnd 0.008523f
C2397 vdd.n1321 gnd 0.010589f
C2398 vdd.n1322 gnd 0.010589f
C2399 vdd.n1323 gnd 0.010589f
C2400 vdd.n1324 gnd 0.008523f
C2401 vdd.n1325 gnd 0.008523f
C2402 vdd.n1326 gnd 0.008523f
C2403 vdd.n1327 gnd 0.010589f
C2404 vdd.n1328 gnd 0.010589f
C2405 vdd.n1329 gnd 0.010589f
C2406 vdd.n1330 gnd 0.008523f
C2407 vdd.n1331 gnd 0.008523f
C2408 vdd.n1332 gnd 0.008523f
C2409 vdd.n1333 gnd 0.010589f
C2410 vdd.n1334 gnd 0.010589f
C2411 vdd.n1335 gnd 0.010589f
C2412 vdd.n1336 gnd 0.008523f
C2413 vdd.n1337 gnd 0.007116f
C2414 vdd.n1338 gnd 0.010589f
C2415 vdd.n1339 gnd 0.010589f
C2416 vdd.t191 gnd 0.130268f
C2417 vdd.t192 gnd 0.139221f
C2418 vdd.t190 gnd 0.170129f
C2419 vdd.n1340 gnd 0.218081f
C2420 vdd.n1341 gnd 0.18408f
C2421 vdd.n1342 gnd 0.018238f
C2422 vdd.n1343 gnd 0.010589f
C2423 vdd.n1344 gnd 0.010589f
C2424 vdd.n1345 gnd 0.010589f
C2425 vdd.n1346 gnd 0.008523f
C2426 vdd.n1347 gnd 0.008523f
C2427 vdd.n1348 gnd 0.008523f
C2428 vdd.n1349 gnd 0.010589f
C2429 vdd.n1350 gnd 0.010589f
C2430 vdd.n1351 gnd 0.010589f
C2431 vdd.n1352 gnd 0.008523f
C2432 vdd.n1353 gnd 0.008523f
C2433 vdd.n1354 gnd 0.008523f
C2434 vdd.n1355 gnd 0.010589f
C2435 vdd.n1356 gnd 0.010589f
C2436 vdd.n1357 gnd 0.010589f
C2437 vdd.n1358 gnd 0.008523f
C2438 vdd.n1359 gnd 0.008523f
C2439 vdd.n1360 gnd 0.008523f
C2440 vdd.n1361 gnd 0.010589f
C2441 vdd.n1362 gnd 0.010589f
C2442 vdd.n1363 gnd 0.010589f
C2443 vdd.n1364 gnd 0.008523f
C2444 vdd.n1365 gnd 0.008523f
C2445 vdd.n1366 gnd 0.008523f
C2446 vdd.n1367 gnd 0.010589f
C2447 vdd.n1368 gnd 0.010589f
C2448 vdd.n1369 gnd 0.010589f
C2449 vdd.n1370 gnd 0.008523f
C2450 vdd.n1371 gnd 0.007074f
C2451 vdd.n1372 gnd 0.024278f
C2452 vdd.n1374 gnd 2.39147f
C2453 vdd.n1375 gnd 0.024278f
C2454 vdd.n1376 gnd 0.004048f
C2455 vdd.n1377 gnd 0.024278f
C2456 vdd.n1378 gnd 0.024113f
C2457 vdd.n1379 gnd 0.010589f
C2458 vdd.n1380 gnd 0.008523f
C2459 vdd.n1381 gnd 0.010589f
C2460 vdd.t169 gnd 0.541056f
C2461 vdd.n1382 gnd 0.708783f
C2462 vdd.n1383 gnd 0.010589f
C2463 vdd.n1384 gnd 0.008523f
C2464 vdd.n1385 gnd 0.010589f
C2465 vdd.n1386 gnd 0.010589f
C2466 vdd.n1387 gnd 0.010589f
C2467 vdd.n1388 gnd 0.008523f
C2468 vdd.n1389 gnd 0.010589f
C2469 vdd.n1390 gnd 1.08211f
C2470 vdd.n1391 gnd 0.010589f
C2471 vdd.n1392 gnd 0.008523f
C2472 vdd.n1393 gnd 0.010589f
C2473 vdd.n1394 gnd 0.010589f
C2474 vdd.n1395 gnd 0.010589f
C2475 vdd.n1396 gnd 0.008523f
C2476 vdd.n1397 gnd 0.010589f
C2477 vdd.n1398 gnd 0.898153f
C2478 vdd.t31 gnd 0.541056f
C2479 vdd.n1399 gnd 0.622214f
C2480 vdd.n1400 gnd 0.010589f
C2481 vdd.n1401 gnd 0.008523f
C2482 vdd.n1402 gnd 0.010589f
C2483 vdd.n1403 gnd 0.010589f
C2484 vdd.n1404 gnd 0.010589f
C2485 vdd.n1405 gnd 0.008523f
C2486 vdd.n1406 gnd 0.010589f
C2487 vdd.n1407 gnd 0.643857f
C2488 vdd.n1408 gnd 0.010589f
C2489 vdd.n1409 gnd 0.008523f
C2490 vdd.n1410 gnd 0.010589f
C2491 vdd.n1411 gnd 0.010589f
C2492 vdd.n1412 gnd 0.010589f
C2493 vdd.n1413 gnd 0.008523f
C2494 vdd.n1414 gnd 0.010589f
C2495 vdd.n1415 gnd 0.611393f
C2496 vdd.n1416 gnd 0.827816f
C2497 vdd.n1417 gnd 0.010589f
C2498 vdd.n1418 gnd 0.008523f
C2499 vdd.n1419 gnd 0.010589f
C2500 vdd.n1420 gnd 0.010589f
C2501 vdd.n1421 gnd 0.010589f
C2502 vdd.n1422 gnd 0.008523f
C2503 vdd.n1423 gnd 0.010589f
C2504 vdd.n1424 gnd 0.898153f
C2505 vdd.n1425 gnd 0.010589f
C2506 vdd.n1426 gnd 0.008523f
C2507 vdd.n1427 gnd 0.010589f
C2508 vdd.n1428 gnd 0.010589f
C2509 vdd.n1429 gnd 0.010589f
C2510 vdd.n1430 gnd 0.008523f
C2511 vdd.n1431 gnd 0.010589f
C2512 vdd.t67 gnd 0.541056f
C2513 vdd.n1432 gnd 0.784531f
C2514 vdd.n1433 gnd 0.010589f
C2515 vdd.n1434 gnd 0.008523f
C2516 vdd.n1435 gnd 0.010589f
C2517 vdd.n1436 gnd 0.010589f
C2518 vdd.n1437 gnd 0.010589f
C2519 vdd.n1438 gnd 0.008523f
C2520 vdd.n1439 gnd 0.010589f
C2521 vdd.n1440 gnd 0.600572f
C2522 vdd.n1441 gnd 0.010589f
C2523 vdd.n1442 gnd 0.008523f
C2524 vdd.n1443 gnd 0.010589f
C2525 vdd.n1444 gnd 0.010589f
C2526 vdd.n1445 gnd 0.010589f
C2527 vdd.n1446 gnd 0.008523f
C2528 vdd.n1447 gnd 0.010589f
C2529 vdd.n1448 gnd 0.77371f
C2530 vdd.n1449 gnd 0.665499f
C2531 vdd.n1450 gnd 0.010589f
C2532 vdd.n1451 gnd 0.008523f
C2533 vdd.n1452 gnd 0.008138f
C2534 vdd.n1453 gnd 0.005811f
C2535 vdd.n1454 gnd 0.005392f
C2536 vdd.n1455 gnd 0.002983f
C2537 vdd.n1456 gnd 0.006849f
C2538 vdd.n1457 gnd 0.002898f
C2539 vdd.n1458 gnd 0.003068f
C2540 vdd.n1459 gnd 0.005392f
C2541 vdd.n1460 gnd 0.002898f
C2542 vdd.n1461 gnd 0.006849f
C2543 vdd.n1462 gnd 0.003068f
C2544 vdd.n1463 gnd 0.005392f
C2545 vdd.n1464 gnd 0.002898f
C2546 vdd.n1465 gnd 0.005137f
C2547 vdd.n1466 gnd 0.005152f
C2548 vdd.t20 gnd 0.014715f
C2549 vdd.n1467 gnd 0.03274f
C2550 vdd.n1468 gnd 0.170386f
C2551 vdd.n1469 gnd 0.002898f
C2552 vdd.n1470 gnd 0.003068f
C2553 vdd.n1471 gnd 0.006849f
C2554 vdd.n1472 gnd 0.006849f
C2555 vdd.n1473 gnd 0.003068f
C2556 vdd.n1474 gnd 0.002898f
C2557 vdd.n1475 gnd 0.005392f
C2558 vdd.n1476 gnd 0.005392f
C2559 vdd.n1477 gnd 0.002898f
C2560 vdd.n1478 gnd 0.003068f
C2561 vdd.n1479 gnd 0.006849f
C2562 vdd.n1480 gnd 0.006849f
C2563 vdd.n1481 gnd 0.003068f
C2564 vdd.n1482 gnd 0.002898f
C2565 vdd.n1483 gnd 0.005392f
C2566 vdd.n1484 gnd 0.005392f
C2567 vdd.n1485 gnd 0.002898f
C2568 vdd.n1486 gnd 0.003068f
C2569 vdd.n1487 gnd 0.006849f
C2570 vdd.n1488 gnd 0.006849f
C2571 vdd.n1489 gnd 0.016193f
C2572 vdd.n1490 gnd 0.002983f
C2573 vdd.n1491 gnd 0.002898f
C2574 vdd.n1492 gnd 0.013938f
C2575 vdd.n1493 gnd 0.009731f
C2576 vdd.t81 gnd 0.03409f
C2577 vdd.t132 gnd 0.03409f
C2578 vdd.n1494 gnd 0.234293f
C2579 vdd.n1495 gnd 0.184235f
C2580 vdd.t54 gnd 0.03409f
C2581 vdd.t114 gnd 0.03409f
C2582 vdd.n1496 gnd 0.234293f
C2583 vdd.n1497 gnd 0.148677f
C2584 vdd.t75 gnd 0.03409f
C2585 vdd.t121 gnd 0.03409f
C2586 vdd.n1498 gnd 0.234293f
C2587 vdd.n1499 gnd 0.148677f
C2588 vdd.t96 gnd 0.03409f
C2589 vdd.t138 gnd 0.03409f
C2590 vdd.n1500 gnd 0.234293f
C2591 vdd.n1501 gnd 0.148677f
C2592 vdd.t68 gnd 0.03409f
C2593 vdd.t28 gnd 0.03409f
C2594 vdd.n1502 gnd 0.234293f
C2595 vdd.n1503 gnd 0.148677f
C2596 vdd.t86 gnd 0.03409f
C2597 vdd.t40 gnd 0.03409f
C2598 vdd.n1504 gnd 0.234293f
C2599 vdd.n1505 gnd 0.148677f
C2600 vdd.t128 gnd 0.03409f
C2601 vdd.t143 gnd 0.03409f
C2602 vdd.n1506 gnd 0.234293f
C2603 vdd.n1507 gnd 0.148677f
C2604 vdd.n1508 gnd 0.005811f
C2605 vdd.n1509 gnd 0.005392f
C2606 vdd.n1510 gnd 0.002983f
C2607 vdd.n1511 gnd 0.006849f
C2608 vdd.n1512 gnd 0.002898f
C2609 vdd.n1513 gnd 0.003068f
C2610 vdd.n1514 gnd 0.005392f
C2611 vdd.n1515 gnd 0.002898f
C2612 vdd.n1516 gnd 0.006849f
C2613 vdd.n1517 gnd 0.003068f
C2614 vdd.n1518 gnd 0.005392f
C2615 vdd.n1519 gnd 0.002898f
C2616 vdd.n1520 gnd 0.005137f
C2617 vdd.n1521 gnd 0.005152f
C2618 vdd.t45 gnd 0.014715f
C2619 vdd.n1522 gnd 0.03274f
C2620 vdd.n1523 gnd 0.170386f
C2621 vdd.n1524 gnd 0.002898f
C2622 vdd.n1525 gnd 0.003068f
C2623 vdd.n1526 gnd 0.006849f
C2624 vdd.n1527 gnd 0.006849f
C2625 vdd.n1528 gnd 0.003068f
C2626 vdd.n1529 gnd 0.002898f
C2627 vdd.n1530 gnd 0.005392f
C2628 vdd.n1531 gnd 0.005392f
C2629 vdd.n1532 gnd 0.002898f
C2630 vdd.n1533 gnd 0.003068f
C2631 vdd.n1534 gnd 0.006849f
C2632 vdd.n1535 gnd 0.006849f
C2633 vdd.n1536 gnd 0.003068f
C2634 vdd.n1537 gnd 0.002898f
C2635 vdd.n1538 gnd 0.005392f
C2636 vdd.n1539 gnd 0.005392f
C2637 vdd.n1540 gnd 0.002898f
C2638 vdd.n1541 gnd 0.003068f
C2639 vdd.n1542 gnd 0.006849f
C2640 vdd.n1543 gnd 0.006849f
C2641 vdd.n1544 gnd 0.016193f
C2642 vdd.n1545 gnd 0.002983f
C2643 vdd.n1546 gnd 0.002898f
C2644 vdd.n1547 gnd 0.013938f
C2645 vdd.n1548 gnd 0.009425f
C2646 vdd.n1549 gnd 0.110616f
C2647 vdd.n1550 gnd 0.005811f
C2648 vdd.n1551 gnd 0.005392f
C2649 vdd.n1552 gnd 0.002983f
C2650 vdd.n1553 gnd 0.006849f
C2651 vdd.n1554 gnd 0.002898f
C2652 vdd.n1555 gnd 0.003068f
C2653 vdd.n1556 gnd 0.005392f
C2654 vdd.n1557 gnd 0.002898f
C2655 vdd.n1558 gnd 0.006849f
C2656 vdd.n1559 gnd 0.003068f
C2657 vdd.n1560 gnd 0.005392f
C2658 vdd.n1561 gnd 0.002898f
C2659 vdd.n1562 gnd 0.005137f
C2660 vdd.n1563 gnd 0.005152f
C2661 vdd.t122 gnd 0.014715f
C2662 vdd.n1564 gnd 0.03274f
C2663 vdd.n1565 gnd 0.170386f
C2664 vdd.n1566 gnd 0.002898f
C2665 vdd.n1567 gnd 0.003068f
C2666 vdd.n1568 gnd 0.006849f
C2667 vdd.n1569 gnd 0.006849f
C2668 vdd.n1570 gnd 0.003068f
C2669 vdd.n1571 gnd 0.002898f
C2670 vdd.n1572 gnd 0.005392f
C2671 vdd.n1573 gnd 0.005392f
C2672 vdd.n1574 gnd 0.002898f
C2673 vdd.n1575 gnd 0.003068f
C2674 vdd.n1576 gnd 0.006849f
C2675 vdd.n1577 gnd 0.006849f
C2676 vdd.n1578 gnd 0.003068f
C2677 vdd.n1579 gnd 0.002898f
C2678 vdd.n1580 gnd 0.005392f
C2679 vdd.n1581 gnd 0.005392f
C2680 vdd.n1582 gnd 0.002898f
C2681 vdd.n1583 gnd 0.003068f
C2682 vdd.n1584 gnd 0.006849f
C2683 vdd.n1585 gnd 0.006849f
C2684 vdd.n1586 gnd 0.016193f
C2685 vdd.n1587 gnd 0.002983f
C2686 vdd.n1588 gnd 0.002898f
C2687 vdd.n1589 gnd 0.013938f
C2688 vdd.n1590 gnd 0.009731f
C2689 vdd.t34 gnd 0.03409f
C2690 vdd.t127 gnd 0.03409f
C2691 vdd.n1591 gnd 0.234293f
C2692 vdd.n1592 gnd 0.184235f
C2693 vdd.t120 gnd 0.03409f
C2694 vdd.t107 gnd 0.03409f
C2695 vdd.n1593 gnd 0.234293f
C2696 vdd.n1594 gnd 0.148677f
C2697 vdd.t78 gnd 0.03409f
C2698 vdd.t24 gnd 0.03409f
C2699 vdd.n1595 gnd 0.234293f
C2700 vdd.n1596 gnd 0.148677f
C2701 vdd.t134 gnd 0.03409f
C2702 vdd.t105 gnd 0.03409f
C2703 vdd.n1597 gnd 0.234293f
C2704 vdd.n1598 gnd 0.148677f
C2705 vdd.t102 gnd 0.03409f
C2706 vdd.t57 gnd 0.03409f
C2707 vdd.n1599 gnd 0.234293f
C2708 vdd.n1600 gnd 0.148677f
C2709 vdd.t51 gnd 0.03409f
C2710 vdd.t103 gnd 0.03409f
C2711 vdd.n1601 gnd 0.234293f
C2712 vdd.n1602 gnd 0.148677f
C2713 vdd.t93 gnd 0.03409f
C2714 vdd.t91 gnd 0.03409f
C2715 vdd.n1603 gnd 0.234293f
C2716 vdd.n1604 gnd 0.148677f
C2717 vdd.n1605 gnd 0.005811f
C2718 vdd.n1606 gnd 0.005392f
C2719 vdd.n1607 gnd 0.002983f
C2720 vdd.n1608 gnd 0.006849f
C2721 vdd.n1609 gnd 0.002898f
C2722 vdd.n1610 gnd 0.003068f
C2723 vdd.n1611 gnd 0.005392f
C2724 vdd.n1612 gnd 0.002898f
C2725 vdd.n1613 gnd 0.006849f
C2726 vdd.n1614 gnd 0.003068f
C2727 vdd.n1615 gnd 0.005392f
C2728 vdd.n1616 gnd 0.002898f
C2729 vdd.n1617 gnd 0.005137f
C2730 vdd.n1618 gnd 0.005152f
C2731 vdd.t32 gnd 0.014715f
C2732 vdd.n1619 gnd 0.03274f
C2733 vdd.n1620 gnd 0.170386f
C2734 vdd.n1621 gnd 0.002898f
C2735 vdd.n1622 gnd 0.003068f
C2736 vdd.n1623 gnd 0.006849f
C2737 vdd.n1624 gnd 0.006849f
C2738 vdd.n1625 gnd 0.003068f
C2739 vdd.n1626 gnd 0.002898f
C2740 vdd.n1627 gnd 0.005392f
C2741 vdd.n1628 gnd 0.005392f
C2742 vdd.n1629 gnd 0.002898f
C2743 vdd.n1630 gnd 0.003068f
C2744 vdd.n1631 gnd 0.006849f
C2745 vdd.n1632 gnd 0.006849f
C2746 vdd.n1633 gnd 0.003068f
C2747 vdd.n1634 gnd 0.002898f
C2748 vdd.n1635 gnd 0.005392f
C2749 vdd.n1636 gnd 0.005392f
C2750 vdd.n1637 gnd 0.002898f
C2751 vdd.n1638 gnd 0.003068f
C2752 vdd.n1639 gnd 0.006849f
C2753 vdd.n1640 gnd 0.006849f
C2754 vdd.n1641 gnd 0.016193f
C2755 vdd.n1642 gnd 0.002983f
C2756 vdd.n1643 gnd 0.002898f
C2757 vdd.n1644 gnd 0.013938f
C2758 vdd.n1645 gnd 0.009425f
C2759 vdd.n1646 gnd 0.065805f
C2760 vdd.n1647 gnd 0.237115f
C2761 vdd.n1648 gnd 0.005811f
C2762 vdd.n1649 gnd 0.005392f
C2763 vdd.n1650 gnd 0.002983f
C2764 vdd.n1651 gnd 0.006849f
C2765 vdd.n1652 gnd 0.002898f
C2766 vdd.n1653 gnd 0.003068f
C2767 vdd.n1654 gnd 0.005392f
C2768 vdd.n1655 gnd 0.002898f
C2769 vdd.n1656 gnd 0.006849f
C2770 vdd.n1657 gnd 0.003068f
C2771 vdd.n1658 gnd 0.005392f
C2772 vdd.n1659 gnd 0.002898f
C2773 vdd.n1660 gnd 0.005137f
C2774 vdd.n1661 gnd 0.005152f
C2775 vdd.t137 gnd 0.014715f
C2776 vdd.n1662 gnd 0.03274f
C2777 vdd.n1663 gnd 0.170386f
C2778 vdd.n1664 gnd 0.002898f
C2779 vdd.n1665 gnd 0.003068f
C2780 vdd.n1666 gnd 0.006849f
C2781 vdd.n1667 gnd 0.006849f
C2782 vdd.n1668 gnd 0.003068f
C2783 vdd.n1669 gnd 0.002898f
C2784 vdd.n1670 gnd 0.005392f
C2785 vdd.n1671 gnd 0.005392f
C2786 vdd.n1672 gnd 0.002898f
C2787 vdd.n1673 gnd 0.003068f
C2788 vdd.n1674 gnd 0.006849f
C2789 vdd.n1675 gnd 0.006849f
C2790 vdd.n1676 gnd 0.003068f
C2791 vdd.n1677 gnd 0.002898f
C2792 vdd.n1678 gnd 0.005392f
C2793 vdd.n1679 gnd 0.005392f
C2794 vdd.n1680 gnd 0.002898f
C2795 vdd.n1681 gnd 0.003068f
C2796 vdd.n1682 gnd 0.006849f
C2797 vdd.n1683 gnd 0.006849f
C2798 vdd.n1684 gnd 0.016193f
C2799 vdd.n1685 gnd 0.002983f
C2800 vdd.n1686 gnd 0.002898f
C2801 vdd.n1687 gnd 0.013938f
C2802 vdd.n1688 gnd 0.009731f
C2803 vdd.t49 gnd 0.03409f
C2804 vdd.t136 gnd 0.03409f
C2805 vdd.n1689 gnd 0.234293f
C2806 vdd.n1690 gnd 0.184235f
C2807 vdd.t135 gnd 0.03409f
C2808 vdd.t117 gnd 0.03409f
C2809 vdd.n1691 gnd 0.234293f
C2810 vdd.n1692 gnd 0.148677f
C2811 vdd.t94 gnd 0.03409f
C2812 vdd.t46 gnd 0.03409f
C2813 vdd.n1693 gnd 0.234293f
C2814 vdd.n1694 gnd 0.148677f
C2815 vdd.t145 gnd 0.03409f
C2816 vdd.t116 gnd 0.03409f
C2817 vdd.n1695 gnd 0.234293f
C2818 vdd.n1696 gnd 0.148677f
C2819 vdd.t112 gnd 0.03409f
C2820 vdd.t71 gnd 0.03409f
C2821 vdd.n1697 gnd 0.234293f
C2822 vdd.n1698 gnd 0.148677f
C2823 vdd.t70 gnd 0.03409f
C2824 vdd.t113 gnd 0.03409f
C2825 vdd.n1699 gnd 0.234293f
C2826 vdd.n1700 gnd 0.148677f
C2827 vdd.t100 gnd 0.03409f
C2828 vdd.t101 gnd 0.03409f
C2829 vdd.n1701 gnd 0.234293f
C2830 vdd.n1702 gnd 0.148677f
C2831 vdd.n1703 gnd 0.005811f
C2832 vdd.n1704 gnd 0.005392f
C2833 vdd.n1705 gnd 0.002983f
C2834 vdd.n1706 gnd 0.006849f
C2835 vdd.n1707 gnd 0.002898f
C2836 vdd.n1708 gnd 0.003068f
C2837 vdd.n1709 gnd 0.005392f
C2838 vdd.n1710 gnd 0.002898f
C2839 vdd.n1711 gnd 0.006849f
C2840 vdd.n1712 gnd 0.003068f
C2841 vdd.n1713 gnd 0.005392f
C2842 vdd.n1714 gnd 0.002898f
C2843 vdd.n1715 gnd 0.005137f
C2844 vdd.n1716 gnd 0.005152f
C2845 vdd.t48 gnd 0.014715f
C2846 vdd.n1717 gnd 0.03274f
C2847 vdd.n1718 gnd 0.170386f
C2848 vdd.n1719 gnd 0.002898f
C2849 vdd.n1720 gnd 0.003068f
C2850 vdd.n1721 gnd 0.006849f
C2851 vdd.n1722 gnd 0.006849f
C2852 vdd.n1723 gnd 0.003068f
C2853 vdd.n1724 gnd 0.002898f
C2854 vdd.n1725 gnd 0.005392f
C2855 vdd.n1726 gnd 0.005392f
C2856 vdd.n1727 gnd 0.002898f
C2857 vdd.n1728 gnd 0.003068f
C2858 vdd.n1729 gnd 0.006849f
C2859 vdd.n1730 gnd 0.006849f
C2860 vdd.n1731 gnd 0.003068f
C2861 vdd.n1732 gnd 0.002898f
C2862 vdd.n1733 gnd 0.005392f
C2863 vdd.n1734 gnd 0.005392f
C2864 vdd.n1735 gnd 0.002898f
C2865 vdd.n1736 gnd 0.003068f
C2866 vdd.n1737 gnd 0.006849f
C2867 vdd.n1738 gnd 0.006849f
C2868 vdd.n1739 gnd 0.016193f
C2869 vdd.n1740 gnd 0.002983f
C2870 vdd.n1741 gnd 0.002898f
C2871 vdd.n1742 gnd 0.013938f
C2872 vdd.n1743 gnd 0.009425f
C2873 vdd.n1744 gnd 0.065805f
C2874 vdd.n1745 gnd 0.265537f
C2875 vdd.n1746 gnd 2.53296f
C2876 vdd.n1747 gnd 0.62456f
C2877 vdd.n1748 gnd 0.008138f
C2878 vdd.n1749 gnd 0.010589f
C2879 vdd.n1750 gnd 0.008523f
C2880 vdd.n1751 gnd 0.010589f
C2881 vdd.n1752 gnd 0.849458f
C2882 vdd.n1753 gnd 0.010589f
C2883 vdd.n1754 gnd 0.008523f
C2884 vdd.n1755 gnd 0.010589f
C2885 vdd.n1756 gnd 0.010589f
C2886 vdd.n1757 gnd 0.010589f
C2887 vdd.n1758 gnd 0.008523f
C2888 vdd.n1759 gnd 0.010589f
C2889 vdd.t23 gnd 0.541056f
C2890 vdd.n1760 gnd 0.898153f
C2891 vdd.n1761 gnd 0.010589f
C2892 vdd.n1762 gnd 0.008523f
C2893 vdd.n1763 gnd 0.010589f
C2894 vdd.n1764 gnd 0.010589f
C2895 vdd.n1765 gnd 0.010589f
C2896 vdd.n1766 gnd 0.008523f
C2897 vdd.n1767 gnd 0.010589f
C2898 vdd.n1768 gnd 0.762889f
C2899 vdd.n1769 gnd 0.010589f
C2900 vdd.n1770 gnd 0.008523f
C2901 vdd.n1771 gnd 0.010589f
C2902 vdd.n1772 gnd 0.010589f
C2903 vdd.n1773 gnd 0.010589f
C2904 vdd.n1774 gnd 0.008523f
C2905 vdd.n1775 gnd 0.010589f
C2906 vdd.n1776 gnd 0.898153f
C2907 vdd.t106 gnd 0.541056f
C2908 vdd.n1777 gnd 0.57893f
C2909 vdd.n1778 gnd 0.010589f
C2910 vdd.n1779 gnd 0.008523f
C2911 vdd.n1780 gnd 0.010589f
C2912 vdd.n1781 gnd 0.010589f
C2913 vdd.n1782 gnd 0.010589f
C2914 vdd.n1783 gnd 0.008523f
C2915 vdd.n1784 gnd 0.010589f
C2916 vdd.n1785 gnd 0.687141f
C2917 vdd.n1786 gnd 0.010589f
C2918 vdd.n1787 gnd 0.008523f
C2919 vdd.n1788 gnd 0.010589f
C2920 vdd.n1789 gnd 0.010589f
C2921 vdd.n1790 gnd 0.010589f
C2922 vdd.n1791 gnd 0.008523f
C2923 vdd.n1792 gnd 0.010589f
C2924 vdd.n1793 gnd 0.568109f
C2925 vdd.n1794 gnd 0.8711f
C2926 vdd.n1795 gnd 0.010589f
C2927 vdd.n1796 gnd 0.008523f
C2928 vdd.n1797 gnd 0.010589f
C2929 vdd.n1798 gnd 0.010589f
C2930 vdd.n1799 gnd 0.010589f
C2931 vdd.n1800 gnd 0.008523f
C2932 vdd.n1801 gnd 0.010589f
C2933 vdd.n1802 gnd 1.05506f
C2934 vdd.n1803 gnd 0.010589f
C2935 vdd.n1804 gnd 0.008523f
C2936 vdd.n1805 gnd 0.010589f
C2937 vdd.n1806 gnd 0.010589f
C2938 vdd.n1807 gnd 0.024113f
C2939 vdd.n1808 gnd 0.010589f
C2940 vdd.n1809 gnd 0.010589f
C2941 vdd.n1810 gnd 0.008523f
C2942 vdd.n1811 gnd 0.010589f
C2943 vdd.t180 gnd 0.541056f
C2944 vdd.n1812 gnd 1.0226f
C2945 vdd.n1813 gnd 0.010589f
C2946 vdd.n1814 gnd 0.008523f
C2947 vdd.n1815 gnd 0.010589f
C2948 vdd.n1816 gnd 0.010589f
C2949 vdd.n1817 gnd 0.009106f
C2950 vdd.n1818 gnd 0.008523f
C2951 vdd.n1820 gnd 0.010589f
C2952 vdd.n1822 gnd 0.008523f
C2953 vdd.n1823 gnd 0.010589f
C2954 vdd.n1824 gnd 0.008523f
C2955 vdd.n1826 gnd 0.010589f
C2956 vdd.n1827 gnd 0.008523f
C2957 vdd.n1828 gnd 0.010589f
C2958 vdd.n1829 gnd 0.010589f
C2959 vdd.n1830 gnd 0.010589f
C2960 vdd.n1831 gnd 0.010589f
C2961 vdd.n1832 gnd 0.010589f
C2962 vdd.n1833 gnd 0.008523f
C2963 vdd.n1835 gnd 0.010589f
C2964 vdd.n1836 gnd 0.010589f
C2965 vdd.n1837 gnd 0.010589f
C2966 vdd.n1838 gnd 0.010589f
C2967 vdd.n1839 gnd 0.010589f
C2968 vdd.n1840 gnd 0.008523f
C2969 vdd.n1842 gnd 0.010589f
C2970 vdd.n1843 gnd 0.010589f
C2971 vdd.n1844 gnd 0.010589f
C2972 vdd.n1845 gnd 0.010589f
C2973 vdd.n1846 gnd 0.007116f
C2974 vdd.t198 gnd 0.130268f
C2975 vdd.t197 gnd 0.139221f
C2976 vdd.t196 gnd 0.170129f
C2977 vdd.n1847 gnd 0.218081f
C2978 vdd.n1848 gnd 0.183228f
C2979 vdd.n1850 gnd 0.010589f
C2980 vdd.n1851 gnd 0.010589f
C2981 vdd.n1852 gnd 0.008523f
C2982 vdd.n1853 gnd 0.010589f
C2983 vdd.n1855 gnd 0.010589f
C2984 vdd.n1856 gnd 0.010589f
C2985 vdd.n1857 gnd 0.010589f
C2986 vdd.n1858 gnd 0.010589f
C2987 vdd.n1859 gnd 0.008523f
C2988 vdd.n1861 gnd 0.010589f
C2989 vdd.n1862 gnd 0.010589f
C2990 vdd.n1863 gnd 0.010589f
C2991 vdd.n1864 gnd 0.010589f
C2992 vdd.n1865 gnd 0.010589f
C2993 vdd.n1866 gnd 0.008523f
C2994 vdd.n1868 gnd 0.010589f
C2995 vdd.n1869 gnd 0.010589f
C2996 vdd.n1870 gnd 0.010589f
C2997 vdd.n1871 gnd 0.010589f
C2998 vdd.n1872 gnd 0.010589f
C2999 vdd.n1873 gnd 0.008523f
C3000 vdd.n1875 gnd 0.010589f
C3001 vdd.n1876 gnd 0.010589f
C3002 vdd.n1877 gnd 0.010589f
C3003 vdd.n1878 gnd 0.010589f
C3004 vdd.n1879 gnd 0.010589f
C3005 vdd.n1880 gnd 0.008523f
C3006 vdd.n1882 gnd 0.010589f
C3007 vdd.n1883 gnd 0.010589f
C3008 vdd.n1884 gnd 0.010589f
C3009 vdd.n1885 gnd 0.010589f
C3010 vdd.n1886 gnd 0.008437f
C3011 vdd.t195 gnd 0.130268f
C3012 vdd.t194 gnd 0.139221f
C3013 vdd.t193 gnd 0.170129f
C3014 vdd.n1887 gnd 0.218081f
C3015 vdd.n1888 gnd 0.183228f
C3016 vdd.n1890 gnd 0.010589f
C3017 vdd.n1891 gnd 0.010589f
C3018 vdd.n1892 gnd 0.008523f
C3019 vdd.n1893 gnd 0.010589f
C3020 vdd.n1895 gnd 0.010589f
C3021 vdd.n1896 gnd 0.010589f
C3022 vdd.n1897 gnd 0.010589f
C3023 vdd.n1898 gnd 0.010589f
C3024 vdd.n1899 gnd 0.008523f
C3025 vdd.n1901 gnd 0.010589f
C3026 vdd.n1902 gnd 0.010589f
C3027 vdd.n1903 gnd 0.010589f
C3028 vdd.n1904 gnd 0.010589f
C3029 vdd.n1905 gnd 0.010589f
C3030 vdd.n1906 gnd 0.008523f
C3031 vdd.n1908 gnd 0.010589f
C3032 vdd.n1909 gnd 0.010589f
C3033 vdd.n1910 gnd 0.010589f
C3034 vdd.n1911 gnd 0.010589f
C3035 vdd.n1912 gnd 0.010589f
C3036 vdd.n1913 gnd 0.010589f
C3037 vdd.n1914 gnd 0.008523f
C3038 vdd.n1916 gnd 0.010589f
C3039 vdd.n1918 gnd 0.010589f
C3040 vdd.n1919 gnd 0.008523f
C3041 vdd.n1920 gnd 0.008523f
C3042 vdd.n1921 gnd 0.010589f
C3043 vdd.n1923 gnd 0.010589f
C3044 vdd.n1924 gnd 0.008523f
C3045 vdd.n1925 gnd 0.008523f
C3046 vdd.n1926 gnd 0.010589f
C3047 vdd.n1928 gnd 0.010589f
C3048 vdd.n1929 gnd 0.010589f
C3049 vdd.n1930 gnd 0.008523f
C3050 vdd.n1931 gnd 0.008523f
C3051 vdd.n1932 gnd 0.008523f
C3052 vdd.n1933 gnd 0.010589f
C3053 vdd.n1935 gnd 0.010589f
C3054 vdd.n1936 gnd 0.010589f
C3055 vdd.n1937 gnd 0.008523f
C3056 vdd.n1938 gnd 0.008523f
C3057 vdd.n1939 gnd 0.008523f
C3058 vdd.n1940 gnd 0.010589f
C3059 vdd.n1942 gnd 0.010589f
C3060 vdd.n1943 gnd 0.010589f
C3061 vdd.n1944 gnd 0.008523f
C3062 vdd.n1945 gnd 0.008523f
C3063 vdd.n1946 gnd 0.008523f
C3064 vdd.n1947 gnd 0.010589f
C3065 vdd.n1949 gnd 0.010589f
C3066 vdd.n1950 gnd 0.010589f
C3067 vdd.n1951 gnd 0.008523f
C3068 vdd.n1952 gnd 0.010589f
C3069 vdd.n1953 gnd 0.010589f
C3070 vdd.n1954 gnd 0.010589f
C3071 vdd.n1955 gnd 0.017386f
C3072 vdd.n1956 gnd 0.005795f
C3073 vdd.n1957 gnd 0.008523f
C3074 vdd.n1958 gnd 0.010589f
C3075 vdd.n1960 gnd 0.010589f
C3076 vdd.n1961 gnd 0.010589f
C3077 vdd.n1962 gnd 0.008523f
C3078 vdd.n1963 gnd 0.008523f
C3079 vdd.n1964 gnd 0.008523f
C3080 vdd.n1965 gnd 0.010589f
C3081 vdd.n1967 gnd 0.010589f
C3082 vdd.n1968 gnd 0.010589f
C3083 vdd.n1969 gnd 0.008523f
C3084 vdd.n1970 gnd 0.008523f
C3085 vdd.n1971 gnd 0.008523f
C3086 vdd.n1972 gnd 0.010589f
C3087 vdd.n1974 gnd 0.010589f
C3088 vdd.n1975 gnd 0.010589f
C3089 vdd.n1976 gnd 0.008523f
C3090 vdd.n1977 gnd 0.008523f
C3091 vdd.n1978 gnd 0.008523f
C3092 vdd.n1979 gnd 0.010589f
C3093 vdd.n1981 gnd 0.010589f
C3094 vdd.n1982 gnd 0.010589f
C3095 vdd.n1983 gnd 0.008523f
C3096 vdd.n1984 gnd 0.008523f
C3097 vdd.n1985 gnd 0.008523f
C3098 vdd.n1986 gnd 0.010589f
C3099 vdd.n1988 gnd 0.010589f
C3100 vdd.n1989 gnd 0.010589f
C3101 vdd.n1990 gnd 0.008523f
C3102 vdd.n1991 gnd 0.010589f
C3103 vdd.n1992 gnd 0.010589f
C3104 vdd.n1993 gnd 0.010589f
C3105 vdd.n1994 gnd 0.017386f
C3106 vdd.n1995 gnd 0.007116f
C3107 vdd.n1996 gnd 0.008523f
C3108 vdd.n1997 gnd 0.010589f
C3109 vdd.n1999 gnd 0.010589f
C3110 vdd.n2000 gnd 0.010589f
C3111 vdd.n2001 gnd 0.008523f
C3112 vdd.n2002 gnd 0.008523f
C3113 vdd.n2003 gnd 0.008523f
C3114 vdd.n2004 gnd 0.010589f
C3115 vdd.n2006 gnd 0.010589f
C3116 vdd.n2007 gnd 0.010589f
C3117 vdd.n2008 gnd 0.008523f
C3118 vdd.n2009 gnd 0.008523f
C3119 vdd.n2010 gnd 0.008523f
C3120 vdd.n2011 gnd 0.010589f
C3121 vdd.n2013 gnd 0.010589f
C3122 vdd.n2014 gnd 0.010589f
C3123 vdd.n2016 gnd 0.010589f
C3124 vdd.n2017 gnd 0.008523f
C3125 vdd.n2018 gnd 0.006777f
C3126 vdd.n2019 gnd 0.0072f
C3127 vdd.n2020 gnd 0.0072f
C3128 vdd.n2021 gnd 0.0072f
C3129 vdd.n2022 gnd 0.0072f
C3130 vdd.n2023 gnd 0.0072f
C3131 vdd.n2024 gnd 0.0072f
C3132 vdd.n2025 gnd 0.0072f
C3133 vdd.n2026 gnd 0.0072f
C3134 vdd.n2028 gnd 0.0072f
C3135 vdd.n2029 gnd 0.0072f
C3136 vdd.n2030 gnd 0.0072f
C3137 vdd.n2031 gnd 0.0072f
C3138 vdd.n2032 gnd 0.0072f
C3139 vdd.n2034 gnd 0.0072f
C3140 vdd.n2036 gnd 0.0072f
C3141 vdd.n2037 gnd 0.0072f
C3142 vdd.n2038 gnd 0.0072f
C3143 vdd.n2039 gnd 0.0072f
C3144 vdd.n2040 gnd 0.0072f
C3145 vdd.n2042 gnd 0.0072f
C3146 vdd.n2044 gnd 0.0072f
C3147 vdd.n2045 gnd 0.0072f
C3148 vdd.n2046 gnd 0.0072f
C3149 vdd.n2047 gnd 0.0072f
C3150 vdd.n2048 gnd 0.0072f
C3151 vdd.n2050 gnd 0.0072f
C3152 vdd.n2052 gnd 0.0072f
C3153 vdd.n2053 gnd 0.0072f
C3154 vdd.n2054 gnd 0.0072f
C3155 vdd.n2055 gnd 0.0072f
C3156 vdd.n2056 gnd 0.0072f
C3157 vdd.n2058 gnd 0.0072f
C3158 vdd.n2059 gnd 0.0072f
C3159 vdd.n2060 gnd 0.0072f
C3160 vdd.n2061 gnd 0.0072f
C3161 vdd.n2062 gnd 0.0072f
C3162 vdd.n2063 gnd 0.0072f
C3163 vdd.n2064 gnd 0.0072f
C3164 vdd.n2065 gnd 0.0072f
C3165 vdd.n2066 gnd 0.005241f
C3166 vdd.n2067 gnd 0.0072f
C3167 vdd.t238 gnd 0.290963f
C3168 vdd.t239 gnd 0.297837f
C3169 vdd.t237 gnd 0.189952f
C3170 vdd.n2068 gnd 0.102658f
C3171 vdd.n2069 gnd 0.058231f
C3172 vdd.n2070 gnd 0.01029f
C3173 vdd.n2071 gnd 0.0072f
C3174 vdd.n2072 gnd 0.0072f
C3175 vdd.n2073 gnd 0.438255f
C3176 vdd.n2074 gnd 0.0072f
C3177 vdd.n2075 gnd 0.0072f
C3178 vdd.n2076 gnd 0.0072f
C3179 vdd.n2077 gnd 0.0072f
C3180 vdd.n2078 gnd 0.0072f
C3181 vdd.n2079 gnd 0.0072f
C3182 vdd.n2080 gnd 0.0072f
C3183 vdd.n2081 gnd 0.0072f
C3184 vdd.n2082 gnd 0.0072f
C3185 vdd.n2083 gnd 0.0072f
C3186 vdd.n2084 gnd 0.0072f
C3187 vdd.n2085 gnd 0.0072f
C3188 vdd.n2086 gnd 0.0072f
C3189 vdd.n2087 gnd 0.0072f
C3190 vdd.n2088 gnd 0.0072f
C3191 vdd.n2089 gnd 0.0072f
C3192 vdd.n2090 gnd 0.0072f
C3193 vdd.n2091 gnd 0.0072f
C3194 vdd.n2092 gnd 0.0072f
C3195 vdd.n2093 gnd 0.0072f
C3196 vdd.t216 gnd 0.290963f
C3197 vdd.t217 gnd 0.297837f
C3198 vdd.t214 gnd 0.189952f
C3199 vdd.n2094 gnd 0.102658f
C3200 vdd.n2095 gnd 0.058231f
C3201 vdd.n2096 gnd 0.0072f
C3202 vdd.n2097 gnd 0.0072f
C3203 vdd.n2098 gnd 0.0072f
C3204 vdd.n2099 gnd 0.0072f
C3205 vdd.n2100 gnd 0.0072f
C3206 vdd.n2101 gnd 0.0072f
C3207 vdd.n2103 gnd 0.0072f
C3208 vdd.n2104 gnd 0.0072f
C3209 vdd.n2105 gnd 0.0072f
C3210 vdd.n2106 gnd 0.0072f
C3211 vdd.n2108 gnd 0.0072f
C3212 vdd.n2110 gnd 0.0072f
C3213 vdd.n2111 gnd 0.0072f
C3214 vdd.n2112 gnd 0.0072f
C3215 vdd.n2113 gnd 0.0072f
C3216 vdd.n2114 gnd 0.0072f
C3217 vdd.n2116 gnd 0.0072f
C3218 vdd.n2118 gnd 0.0072f
C3219 vdd.n2119 gnd 0.0072f
C3220 vdd.n2120 gnd 0.0072f
C3221 vdd.n2121 gnd 0.0072f
C3222 vdd.n2122 gnd 0.0072f
C3223 vdd.n2124 gnd 0.0072f
C3224 vdd.n2126 gnd 0.0072f
C3225 vdd.n2127 gnd 0.0072f
C3226 vdd.n2128 gnd 0.005241f
C3227 vdd.n2129 gnd 0.01029f
C3228 vdd.n2130 gnd 0.005559f
C3229 vdd.n2131 gnd 0.0072f
C3230 vdd.n2133 gnd 0.0072f
C3231 vdd.n2134 gnd 0.017085f
C3232 vdd.n2135 gnd 0.017085f
C3233 vdd.n2136 gnd 0.015952f
C3234 vdd.n2137 gnd 0.0072f
C3235 vdd.n2138 gnd 0.0072f
C3236 vdd.n2139 gnd 0.0072f
C3237 vdd.n2140 gnd 0.0072f
C3238 vdd.n2141 gnd 0.0072f
C3239 vdd.n2142 gnd 0.0072f
C3240 vdd.n2143 gnd 0.0072f
C3241 vdd.n2144 gnd 0.0072f
C3242 vdd.n2145 gnd 0.0072f
C3243 vdd.n2146 gnd 0.0072f
C3244 vdd.n2147 gnd 0.0072f
C3245 vdd.n2148 gnd 0.0072f
C3246 vdd.n2149 gnd 0.0072f
C3247 vdd.n2150 gnd 0.0072f
C3248 vdd.n2151 gnd 0.0072f
C3249 vdd.n2152 gnd 0.0072f
C3250 vdd.n2153 gnd 0.0072f
C3251 vdd.n2154 gnd 0.0072f
C3252 vdd.n2155 gnd 0.0072f
C3253 vdd.n2156 gnd 0.0072f
C3254 vdd.n2157 gnd 0.0072f
C3255 vdd.n2158 gnd 0.0072f
C3256 vdd.n2159 gnd 0.0072f
C3257 vdd.n2160 gnd 0.0072f
C3258 vdd.n2161 gnd 0.0072f
C3259 vdd.n2162 gnd 0.0072f
C3260 vdd.n2163 gnd 0.0072f
C3261 vdd.n2164 gnd 0.0072f
C3262 vdd.n2165 gnd 0.0072f
C3263 vdd.n2166 gnd 0.0072f
C3264 vdd.n2167 gnd 0.0072f
C3265 vdd.n2168 gnd 0.0072f
C3266 vdd.n2169 gnd 0.0072f
C3267 vdd.n2170 gnd 0.0072f
C3268 vdd.n2171 gnd 0.0072f
C3269 vdd.n2172 gnd 0.0072f
C3270 vdd.n2173 gnd 0.0072f
C3271 vdd.n2174 gnd 0.232654f
C3272 vdd.n2175 gnd 0.0072f
C3273 vdd.n2176 gnd 0.0072f
C3274 vdd.n2177 gnd 0.0072f
C3275 vdd.n2178 gnd 0.0072f
C3276 vdd.n2179 gnd 0.0072f
C3277 vdd.n2180 gnd 0.0072f
C3278 vdd.n2181 gnd 0.0072f
C3279 vdd.n2182 gnd 0.0072f
C3280 vdd.n2183 gnd 0.0072f
C3281 vdd.n2184 gnd 0.0072f
C3282 vdd.n2185 gnd 0.0072f
C3283 vdd.n2186 gnd 0.0072f
C3284 vdd.n2187 gnd 0.0072f
C3285 vdd.n2188 gnd 0.0072f
C3286 vdd.n2189 gnd 0.0072f
C3287 vdd.n2190 gnd 0.0072f
C3288 vdd.n2191 gnd 0.0072f
C3289 vdd.n2192 gnd 0.0072f
C3290 vdd.n2193 gnd 0.0072f
C3291 vdd.n2194 gnd 0.0072f
C3292 vdd.n2195 gnd 0.015952f
C3293 vdd.n2197 gnd 0.017085f
C3294 vdd.n2198 gnd 0.017085f
C3295 vdd.n2199 gnd 0.0072f
C3296 vdd.n2200 gnd 0.005559f
C3297 vdd.n2201 gnd 0.0072f
C3298 vdd.n2203 gnd 0.0072f
C3299 vdd.n2205 gnd 0.0072f
C3300 vdd.n2206 gnd 0.0072f
C3301 vdd.n2207 gnd 0.0072f
C3302 vdd.n2208 gnd 0.0072f
C3303 vdd.n2209 gnd 0.0072f
C3304 vdd.n2211 gnd 0.0072f
C3305 vdd.n2213 gnd 0.0072f
C3306 vdd.n2214 gnd 0.0072f
C3307 vdd.n2215 gnd 0.0072f
C3308 vdd.n2216 gnd 0.0072f
C3309 vdd.n2217 gnd 0.0072f
C3310 vdd.n2219 gnd 0.0072f
C3311 vdd.n2221 gnd 0.0072f
C3312 vdd.n2222 gnd 0.0072f
C3313 vdd.n2223 gnd 0.0072f
C3314 vdd.n2224 gnd 0.0072f
C3315 vdd.n2225 gnd 0.0072f
C3316 vdd.n2227 gnd 0.0072f
C3317 vdd.n2229 gnd 0.0072f
C3318 vdd.n2230 gnd 0.0072f
C3319 vdd.n2231 gnd 0.021477f
C3320 vdd.n2232 gnd 0.636669f
C3321 vdd.n2234 gnd 0.008523f
C3322 vdd.n2235 gnd 0.008523f
C3323 vdd.n2236 gnd 0.010589f
C3324 vdd.n2238 gnd 0.010589f
C3325 vdd.n2239 gnd 0.010589f
C3326 vdd.n2240 gnd 0.008523f
C3327 vdd.n2241 gnd 0.007074f
C3328 vdd.n2242 gnd 0.024278f
C3329 vdd.n2243 gnd 0.024113f
C3330 vdd.n2244 gnd 0.007074f
C3331 vdd.n2245 gnd 0.024113f
C3332 vdd.n2246 gnd 1.42839f
C3333 vdd.n2247 gnd 0.024113f
C3334 vdd.n2248 gnd 0.024278f
C3335 vdd.n2249 gnd 0.004048f
C3336 vdd.t182 gnd 0.130268f
C3337 vdd.t181 gnd 0.139221f
C3338 vdd.t179 gnd 0.170129f
C3339 vdd.n2250 gnd 0.218081f
C3340 vdd.n2251 gnd 0.183228f
C3341 vdd.n2252 gnd 0.013125f
C3342 vdd.n2253 gnd 0.004474f
C3343 vdd.n2254 gnd 0.009106f
C3344 vdd.n2255 gnd 0.636669f
C3345 vdd.n2256 gnd 0.021477f
C3346 vdd.n2257 gnd 0.0072f
C3347 vdd.n2258 gnd 0.0072f
C3348 vdd.n2259 gnd 0.0072f
C3349 vdd.n2261 gnd 0.0072f
C3350 vdd.n2263 gnd 0.0072f
C3351 vdd.n2264 gnd 0.0072f
C3352 vdd.n2265 gnd 0.0072f
C3353 vdd.n2266 gnd 0.0072f
C3354 vdd.n2267 gnd 0.0072f
C3355 vdd.n2269 gnd 0.0072f
C3356 vdd.n2271 gnd 0.0072f
C3357 vdd.n2272 gnd 0.0072f
C3358 vdd.n2273 gnd 0.0072f
C3359 vdd.n2274 gnd 0.0072f
C3360 vdd.n2275 gnd 0.0072f
C3361 vdd.n2277 gnd 0.0072f
C3362 vdd.n2279 gnd 0.0072f
C3363 vdd.n2280 gnd 0.0072f
C3364 vdd.n2281 gnd 0.0072f
C3365 vdd.n2282 gnd 0.0072f
C3366 vdd.n2283 gnd 0.0072f
C3367 vdd.n2285 gnd 0.0072f
C3368 vdd.n2287 gnd 0.0072f
C3369 vdd.n2288 gnd 0.0072f
C3370 vdd.n2289 gnd 0.017085f
C3371 vdd.n2290 gnd 0.015952f
C3372 vdd.n2291 gnd 0.015952f
C3373 vdd.n2292 gnd 1.06047f
C3374 vdd.n2293 gnd 0.015952f
C3375 vdd.n2294 gnd 0.015952f
C3376 vdd.n2295 gnd 0.0072f
C3377 vdd.n2296 gnd 0.0072f
C3378 vdd.n2297 gnd 0.0072f
C3379 vdd.n2298 gnd 0.459898f
C3380 vdd.n2299 gnd 0.0072f
C3381 vdd.n2300 gnd 0.0072f
C3382 vdd.n2301 gnd 0.0072f
C3383 vdd.n2302 gnd 0.0072f
C3384 vdd.n2303 gnd 0.0072f
C3385 vdd.n2304 gnd 0.735836f
C3386 vdd.n2305 gnd 0.0072f
C3387 vdd.n2306 gnd 0.0072f
C3388 vdd.n2307 gnd 0.0072f
C3389 vdd.n2308 gnd 0.0072f
C3390 vdd.n2309 gnd 0.0072f
C3391 vdd.n2310 gnd 0.735836f
C3392 vdd.n2311 gnd 0.0072f
C3393 vdd.n2312 gnd 0.0072f
C3394 vdd.n2313 gnd 0.006353f
C3395 vdd.n2314 gnd 0.020858f
C3396 vdd.n2315 gnd 0.004447f
C3397 vdd.n2316 gnd 0.0072f
C3398 vdd.n2317 gnd 0.405792f
C3399 vdd.n2318 gnd 0.0072f
C3400 vdd.n2319 gnd 0.0072f
C3401 vdd.n2320 gnd 0.0072f
C3402 vdd.n2321 gnd 0.0072f
C3403 vdd.n2322 gnd 0.0072f
C3404 vdd.n2323 gnd 0.492361f
C3405 vdd.n2324 gnd 0.0072f
C3406 vdd.n2325 gnd 0.0072f
C3407 vdd.n2326 gnd 0.0072f
C3408 vdd.n2327 gnd 0.0072f
C3409 vdd.n2328 gnd 0.0072f
C3410 vdd.n2329 gnd 0.654678f
C3411 vdd.n2330 gnd 0.0072f
C3412 vdd.n2331 gnd 0.0072f
C3413 vdd.n2332 gnd 0.0072f
C3414 vdd.n2333 gnd 0.0072f
C3415 vdd.n2334 gnd 0.0072f
C3416 vdd.n2335 gnd 0.58434f
C3417 vdd.n2336 gnd 0.0072f
C3418 vdd.n2337 gnd 0.0072f
C3419 vdd.n2338 gnd 0.0072f
C3420 vdd.n2339 gnd 0.0072f
C3421 vdd.n2340 gnd 0.0072f
C3422 vdd.n2341 gnd 0.422024f
C3423 vdd.n2342 gnd 0.0072f
C3424 vdd.n2343 gnd 0.0072f
C3425 vdd.n2344 gnd 0.0072f
C3426 vdd.n2345 gnd 0.0072f
C3427 vdd.n2346 gnd 0.0072f
C3428 vdd.n2347 gnd 0.232654f
C3429 vdd.n2348 gnd 0.0072f
C3430 vdd.n2349 gnd 0.0072f
C3431 vdd.n2350 gnd 0.0072f
C3432 vdd.n2351 gnd 0.0072f
C3433 vdd.n2352 gnd 0.0072f
C3434 vdd.n2353 gnd 0.405792f
C3435 vdd.n2354 gnd 0.0072f
C3436 vdd.n2355 gnd 0.0072f
C3437 vdd.n2356 gnd 0.0072f
C3438 vdd.n2357 gnd 0.0072f
C3439 vdd.n2358 gnd 0.0072f
C3440 vdd.n2359 gnd 0.735836f
C3441 vdd.n2360 gnd 0.0072f
C3442 vdd.n2361 gnd 0.0072f
C3443 vdd.n2362 gnd 0.0072f
C3444 vdd.n2363 gnd 0.0072f
C3445 vdd.n2364 gnd 0.0072f
C3446 vdd.n2365 gnd 0.0072f
C3447 vdd.n2366 gnd 0.0072f
C3448 vdd.n2367 gnd 0.573519f
C3449 vdd.n2368 gnd 0.0072f
C3450 vdd.n2369 gnd 0.0072f
C3451 vdd.n2370 gnd 0.0072f
C3452 vdd.n2371 gnd 0.0072f
C3453 vdd.n2372 gnd 0.0072f
C3454 vdd.n2373 gnd 0.0072f
C3455 vdd.n2374 gnd 0.459898f
C3456 vdd.n2375 gnd 0.0072f
C3457 vdd.n2376 gnd 0.0072f
C3458 vdd.n2377 gnd 0.0072f
C3459 vdd.n2378 gnd 0.016828f
C3460 vdd.n2379 gnd 0.016208f
C3461 vdd.n2380 gnd 0.0072f
C3462 vdd.n2381 gnd 0.0072f
C3463 vdd.n2382 gnd 0.005559f
C3464 vdd.n2383 gnd 0.0072f
C3465 vdd.n2384 gnd 0.0072f
C3466 vdd.n2385 gnd 0.005241f
C3467 vdd.n2386 gnd 0.0072f
C3468 vdd.n2387 gnd 0.0072f
C3469 vdd.n2388 gnd 0.0072f
C3470 vdd.n2389 gnd 0.0072f
C3471 vdd.n2390 gnd 0.0072f
C3472 vdd.n2391 gnd 0.0072f
C3473 vdd.n2392 gnd 0.0072f
C3474 vdd.n2393 gnd 0.0072f
C3475 vdd.n2394 gnd 0.0072f
C3476 vdd.n2395 gnd 0.0072f
C3477 vdd.n2396 gnd 0.0072f
C3478 vdd.n2397 gnd 0.0072f
C3479 vdd.n2398 gnd 0.0072f
C3480 vdd.n2399 gnd 0.0072f
C3481 vdd.n2400 gnd 0.0072f
C3482 vdd.n2401 gnd 0.0072f
C3483 vdd.n2402 gnd 0.0072f
C3484 vdd.n2403 gnd 0.0072f
C3485 vdd.n2404 gnd 0.0072f
C3486 vdd.n2405 gnd 0.0072f
C3487 vdd.n2406 gnd 0.0072f
C3488 vdd.n2407 gnd 0.0072f
C3489 vdd.n2408 gnd 0.0072f
C3490 vdd.n2409 gnd 0.0072f
C3491 vdd.n2410 gnd 0.0072f
C3492 vdd.n2411 gnd 0.0072f
C3493 vdd.n2412 gnd 0.0072f
C3494 vdd.n2413 gnd 0.0072f
C3495 vdd.n2414 gnd 0.0072f
C3496 vdd.n2415 gnd 0.0072f
C3497 vdd.n2416 gnd 0.0072f
C3498 vdd.n2417 gnd 0.0072f
C3499 vdd.n2418 gnd 0.0072f
C3500 vdd.n2419 gnd 0.0072f
C3501 vdd.n2420 gnd 0.0072f
C3502 vdd.n2421 gnd 0.0072f
C3503 vdd.n2422 gnd 0.0072f
C3504 vdd.n2423 gnd 0.0072f
C3505 vdd.n2424 gnd 0.0072f
C3506 vdd.n2425 gnd 0.0072f
C3507 vdd.n2426 gnd 0.0072f
C3508 vdd.n2427 gnd 0.0072f
C3509 vdd.n2428 gnd 0.0072f
C3510 vdd.n2429 gnd 0.0072f
C3511 vdd.n2430 gnd 0.0072f
C3512 vdd.n2431 gnd 0.0072f
C3513 vdd.n2432 gnd 0.0072f
C3514 vdd.n2433 gnd 0.0072f
C3515 vdd.n2434 gnd 0.0072f
C3516 vdd.n2435 gnd 0.0072f
C3517 vdd.n2436 gnd 0.0072f
C3518 vdd.n2437 gnd 0.0072f
C3519 vdd.n2438 gnd 0.0072f
C3520 vdd.n2439 gnd 0.0072f
C3521 vdd.n2440 gnd 0.0072f
C3522 vdd.n2441 gnd 0.0072f
C3523 vdd.n2442 gnd 0.0072f
C3524 vdd.n2443 gnd 0.0072f
C3525 vdd.n2444 gnd 0.0072f
C3526 vdd.n2445 gnd 0.0072f
C3527 vdd.n2446 gnd 0.017085f
C3528 vdd.n2447 gnd 0.015952f
C3529 vdd.n2448 gnd 0.015952f
C3530 vdd.n2449 gnd 0.898153f
C3531 vdd.n2450 gnd 0.015952f
C3532 vdd.n2451 gnd 0.017085f
C3533 vdd.n2452 gnd 0.016208f
C3534 vdd.n2453 gnd 0.0072f
C3535 vdd.n2454 gnd 0.0072f
C3536 vdd.n2455 gnd 0.0072f
C3537 vdd.n2456 gnd 0.005559f
C3538 vdd.n2457 gnd 0.01029f
C3539 vdd.n2458 gnd 0.005241f
C3540 vdd.n2459 gnd 0.0072f
C3541 vdd.n2460 gnd 0.0072f
C3542 vdd.n2461 gnd 0.0072f
C3543 vdd.n2462 gnd 0.0072f
C3544 vdd.n2463 gnd 0.0072f
C3545 vdd.n2464 gnd 0.0072f
C3546 vdd.n2465 gnd 0.0072f
C3547 vdd.n2466 gnd 0.0072f
C3548 vdd.n2467 gnd 0.0072f
C3549 vdd.n2468 gnd 0.0072f
C3550 vdd.n2469 gnd 0.0072f
C3551 vdd.n2470 gnd 0.0072f
C3552 vdd.n2471 gnd 0.0072f
C3553 vdd.n2472 gnd 0.0072f
C3554 vdd.n2473 gnd 0.0072f
C3555 vdd.n2474 gnd 0.0072f
C3556 vdd.n2475 gnd 0.0072f
C3557 vdd.n2476 gnd 0.0072f
C3558 vdd.n2477 gnd 0.0072f
C3559 vdd.n2478 gnd 0.0072f
C3560 vdd.n2479 gnd 0.0072f
C3561 vdd.n2480 gnd 0.0072f
C3562 vdd.n2481 gnd 0.0072f
C3563 vdd.n2482 gnd 0.0072f
C3564 vdd.n2483 gnd 0.0072f
C3565 vdd.n2484 gnd 0.0072f
C3566 vdd.n2485 gnd 0.0072f
C3567 vdd.n2486 gnd 0.0072f
C3568 vdd.n2487 gnd 0.0072f
C3569 vdd.n2488 gnd 0.0072f
C3570 vdd.n2489 gnd 0.0072f
C3571 vdd.n2490 gnd 0.0072f
C3572 vdd.n2491 gnd 0.0072f
C3573 vdd.n2492 gnd 0.0072f
C3574 vdd.n2493 gnd 0.0072f
C3575 vdd.n2494 gnd 0.0072f
C3576 vdd.n2495 gnd 0.0072f
C3577 vdd.n2496 gnd 0.0072f
C3578 vdd.n2497 gnd 0.0072f
C3579 vdd.n2498 gnd 0.0072f
C3580 vdd.n2499 gnd 0.0072f
C3581 vdd.n2500 gnd 0.0072f
C3582 vdd.n2501 gnd 0.0072f
C3583 vdd.n2502 gnd 0.0072f
C3584 vdd.n2503 gnd 0.0072f
C3585 vdd.n2504 gnd 0.0072f
C3586 vdd.n2505 gnd 0.0072f
C3587 vdd.n2506 gnd 0.0072f
C3588 vdd.n2507 gnd 0.0072f
C3589 vdd.n2508 gnd 0.0072f
C3590 vdd.n2509 gnd 0.0072f
C3591 vdd.n2510 gnd 0.0072f
C3592 vdd.n2511 gnd 0.0072f
C3593 vdd.n2512 gnd 0.0072f
C3594 vdd.n2513 gnd 0.0072f
C3595 vdd.n2514 gnd 0.0072f
C3596 vdd.n2515 gnd 0.0072f
C3597 vdd.n2516 gnd 0.0072f
C3598 vdd.n2517 gnd 0.0072f
C3599 vdd.n2518 gnd 0.0072f
C3600 vdd.n2519 gnd 0.017085f
C3601 vdd.n2520 gnd 0.017085f
C3602 vdd.n2521 gnd 0.898153f
C3603 vdd.t151 gnd 3.19223f
C3604 vdd.t12 gnd 3.19223f
C3605 vdd.n2554 gnd 0.017085f
C3606 vdd.n2555 gnd 0.0072f
C3607 vdd.t209 gnd 0.290963f
C3608 vdd.t210 gnd 0.297837f
C3609 vdd.t207 gnd 0.189952f
C3610 vdd.n2556 gnd 0.102658f
C3611 vdd.n2557 gnd 0.058231f
C3612 vdd.n2558 gnd 0.0072f
C3613 vdd.t223 gnd 0.290963f
C3614 vdd.t224 gnd 0.297837f
C3615 vdd.t222 gnd 0.189952f
C3616 vdd.n2559 gnd 0.102658f
C3617 vdd.n2560 gnd 0.058231f
C3618 vdd.n2561 gnd 0.01029f
C3619 vdd.n2562 gnd 0.0072f
C3620 vdd.n2563 gnd 0.0072f
C3621 vdd.n2564 gnd 0.0072f
C3622 vdd.n2565 gnd 0.0072f
C3623 vdd.n2566 gnd 0.0072f
C3624 vdd.n2567 gnd 0.0072f
C3625 vdd.n2568 gnd 0.0072f
C3626 vdd.n2569 gnd 0.0072f
C3627 vdd.n2570 gnd 0.0072f
C3628 vdd.n2571 gnd 0.0072f
C3629 vdd.n2572 gnd 0.0072f
C3630 vdd.n2573 gnd 0.0072f
C3631 vdd.n2574 gnd 0.0072f
C3632 vdd.n2575 gnd 0.0072f
C3633 vdd.n2576 gnd 0.0072f
C3634 vdd.n2577 gnd 0.0072f
C3635 vdd.n2578 gnd 0.0072f
C3636 vdd.n2579 gnd 0.0072f
C3637 vdd.n2580 gnd 0.0072f
C3638 vdd.n2581 gnd 0.0072f
C3639 vdd.n2582 gnd 0.0072f
C3640 vdd.n2583 gnd 0.0072f
C3641 vdd.n2584 gnd 0.0072f
C3642 vdd.n2585 gnd 0.0072f
C3643 vdd.n2586 gnd 0.0072f
C3644 vdd.n2587 gnd 0.0072f
C3645 vdd.n2588 gnd 0.0072f
C3646 vdd.n2589 gnd 0.0072f
C3647 vdd.n2590 gnd 0.0072f
C3648 vdd.n2591 gnd 0.0072f
C3649 vdd.n2592 gnd 0.0072f
C3650 vdd.n2593 gnd 0.0072f
C3651 vdd.n2594 gnd 0.0072f
C3652 vdd.n2595 gnd 0.0072f
C3653 vdd.n2596 gnd 0.0072f
C3654 vdd.n2597 gnd 0.0072f
C3655 vdd.n2598 gnd 0.0072f
C3656 vdd.n2599 gnd 0.0072f
C3657 vdd.n2600 gnd 0.0072f
C3658 vdd.n2601 gnd 0.0072f
C3659 vdd.n2602 gnd 0.0072f
C3660 vdd.n2603 gnd 0.0072f
C3661 vdd.n2604 gnd 0.0072f
C3662 vdd.n2605 gnd 0.0072f
C3663 vdd.n2606 gnd 0.0072f
C3664 vdd.n2607 gnd 0.0072f
C3665 vdd.n2608 gnd 0.0072f
C3666 vdd.n2609 gnd 0.0072f
C3667 vdd.n2610 gnd 0.0072f
C3668 vdd.n2611 gnd 0.0072f
C3669 vdd.n2612 gnd 0.0072f
C3670 vdd.n2613 gnd 0.0072f
C3671 vdd.n2614 gnd 0.0072f
C3672 vdd.n2615 gnd 0.0072f
C3673 vdd.n2616 gnd 0.0072f
C3674 vdd.n2617 gnd 0.0072f
C3675 vdd.n2618 gnd 0.005241f
C3676 vdd.n2619 gnd 0.0072f
C3677 vdd.n2620 gnd 0.0072f
C3678 vdd.n2621 gnd 0.005559f
C3679 vdd.n2622 gnd 0.0072f
C3680 vdd.n2623 gnd 0.0072f
C3681 vdd.n2624 gnd 0.017085f
C3682 vdd.n2625 gnd 0.015952f
C3683 vdd.n2626 gnd 0.0072f
C3684 vdd.n2627 gnd 0.0072f
C3685 vdd.n2628 gnd 0.0072f
C3686 vdd.n2629 gnd 0.0072f
C3687 vdd.n2630 gnd 0.0072f
C3688 vdd.n2631 gnd 0.0072f
C3689 vdd.n2632 gnd 0.0072f
C3690 vdd.n2633 gnd 0.0072f
C3691 vdd.n2634 gnd 0.0072f
C3692 vdd.n2635 gnd 0.0072f
C3693 vdd.n2636 gnd 0.0072f
C3694 vdd.n2637 gnd 0.0072f
C3695 vdd.n2638 gnd 0.0072f
C3696 vdd.n2639 gnd 0.0072f
C3697 vdd.n2640 gnd 0.0072f
C3698 vdd.n2641 gnd 0.0072f
C3699 vdd.n2642 gnd 0.0072f
C3700 vdd.n2643 gnd 0.0072f
C3701 vdd.n2644 gnd 0.0072f
C3702 vdd.n2645 gnd 0.0072f
C3703 vdd.n2646 gnd 0.0072f
C3704 vdd.n2647 gnd 0.0072f
C3705 vdd.n2648 gnd 0.0072f
C3706 vdd.n2649 gnd 0.0072f
C3707 vdd.n2650 gnd 0.0072f
C3708 vdd.n2651 gnd 0.0072f
C3709 vdd.n2652 gnd 0.0072f
C3710 vdd.n2653 gnd 0.0072f
C3711 vdd.n2654 gnd 0.0072f
C3712 vdd.n2655 gnd 0.0072f
C3713 vdd.n2656 gnd 0.0072f
C3714 vdd.n2657 gnd 0.0072f
C3715 vdd.n2658 gnd 0.0072f
C3716 vdd.n2659 gnd 0.0072f
C3717 vdd.n2660 gnd 0.0072f
C3718 vdd.n2661 gnd 0.0072f
C3719 vdd.n2662 gnd 0.0072f
C3720 vdd.n2663 gnd 0.0072f
C3721 vdd.n2664 gnd 0.0072f
C3722 vdd.n2665 gnd 0.0072f
C3723 vdd.n2666 gnd 0.0072f
C3724 vdd.n2667 gnd 0.0072f
C3725 vdd.n2668 gnd 0.0072f
C3726 vdd.n2669 gnd 0.0072f
C3727 vdd.n2670 gnd 0.0072f
C3728 vdd.n2671 gnd 0.0072f
C3729 vdd.n2672 gnd 0.0072f
C3730 vdd.n2673 gnd 0.0072f
C3731 vdd.n2674 gnd 0.0072f
C3732 vdd.n2675 gnd 0.0072f
C3733 vdd.n2676 gnd 0.0072f
C3734 vdd.n2677 gnd 0.232654f
C3735 vdd.n2678 gnd 0.0072f
C3736 vdd.n2679 gnd 0.0072f
C3737 vdd.n2680 gnd 0.0072f
C3738 vdd.n2681 gnd 0.0072f
C3739 vdd.n2682 gnd 0.0072f
C3740 vdd.n2683 gnd 0.0072f
C3741 vdd.n2684 gnd 0.0072f
C3742 vdd.n2685 gnd 0.0072f
C3743 vdd.n2686 gnd 0.0072f
C3744 vdd.n2687 gnd 0.0072f
C3745 vdd.n2688 gnd 0.0072f
C3746 vdd.n2689 gnd 0.0072f
C3747 vdd.n2690 gnd 0.0072f
C3748 vdd.n2691 gnd 0.0072f
C3749 vdd.n2692 gnd 0.0072f
C3750 vdd.n2693 gnd 0.0072f
C3751 vdd.n2694 gnd 0.0072f
C3752 vdd.n2695 gnd 0.0072f
C3753 vdd.n2696 gnd 0.0072f
C3754 vdd.n2697 gnd 0.0072f
C3755 vdd.n2698 gnd 0.438255f
C3756 vdd.n2699 gnd 0.0072f
C3757 vdd.n2700 gnd 0.0072f
C3758 vdd.n2701 gnd 0.0072f
C3759 vdd.n2702 gnd 0.0072f
C3760 vdd.n2703 gnd 0.0072f
C3761 vdd.n2704 gnd 0.015952f
C3762 vdd.n2705 gnd 0.017085f
C3763 vdd.n2706 gnd 0.017085f
C3764 vdd.n2707 gnd 0.0072f
C3765 vdd.n2708 gnd 0.0072f
C3766 vdd.n2709 gnd 0.0072f
C3767 vdd.n2710 gnd 0.005559f
C3768 vdd.n2711 gnd 0.01029f
C3769 vdd.n2712 gnd 0.005241f
C3770 vdd.n2713 gnd 0.0072f
C3771 vdd.n2714 gnd 0.0072f
C3772 vdd.n2715 gnd 0.0072f
C3773 vdd.n2716 gnd 0.0072f
C3774 vdd.n2717 gnd 0.0072f
C3775 vdd.n2718 gnd 0.0072f
C3776 vdd.n2719 gnd 0.0072f
C3777 vdd.n2720 gnd 0.0072f
C3778 vdd.n2721 gnd 0.0072f
C3779 vdd.n2722 gnd 0.0072f
C3780 vdd.n2723 gnd 0.0072f
C3781 vdd.n2724 gnd 0.0072f
C3782 vdd.n2725 gnd 0.0072f
C3783 vdd.n2726 gnd 0.0072f
C3784 vdd.n2727 gnd 0.0072f
C3785 vdd.n2728 gnd 0.0072f
C3786 vdd.n2729 gnd 0.0072f
C3787 vdd.n2730 gnd 0.0072f
C3788 vdd.n2731 gnd 0.0072f
C3789 vdd.n2732 gnd 0.0072f
C3790 vdd.n2733 gnd 0.0072f
C3791 vdd.n2734 gnd 0.0072f
C3792 vdd.n2735 gnd 0.0072f
C3793 vdd.n2736 gnd 0.0072f
C3794 vdd.n2737 gnd 0.0072f
C3795 vdd.n2738 gnd 0.0072f
C3796 vdd.n2739 gnd 0.0072f
C3797 vdd.n2740 gnd 0.0072f
C3798 vdd.n2741 gnd 0.0072f
C3799 vdd.n2742 gnd 0.0072f
C3800 vdd.n2743 gnd 0.0072f
C3801 vdd.n2744 gnd 0.0072f
C3802 vdd.n2745 gnd 0.0072f
C3803 vdd.n2746 gnd 0.0072f
C3804 vdd.n2747 gnd 0.0072f
C3805 vdd.n2748 gnd 0.0072f
C3806 vdd.n2749 gnd 0.0072f
C3807 vdd.n2750 gnd 0.0072f
C3808 vdd.n2751 gnd 0.0072f
C3809 vdd.n2752 gnd 0.0072f
C3810 vdd.n2753 gnd 0.0072f
C3811 vdd.n2754 gnd 0.0072f
C3812 vdd.n2755 gnd 0.0072f
C3813 vdd.n2756 gnd 0.0072f
C3814 vdd.n2757 gnd 0.0072f
C3815 vdd.n2758 gnd 0.0072f
C3816 vdd.n2759 gnd 0.0072f
C3817 vdd.n2760 gnd 0.0072f
C3818 vdd.n2761 gnd 0.0072f
C3819 vdd.n2762 gnd 0.0072f
C3820 vdd.n2763 gnd 0.0072f
C3821 vdd.n2764 gnd 0.0072f
C3822 vdd.n2765 gnd 0.0072f
C3823 vdd.n2766 gnd 0.0072f
C3824 vdd.n2767 gnd 0.0072f
C3825 vdd.n2768 gnd 0.0072f
C3826 vdd.n2769 gnd 0.0072f
C3827 vdd.n2770 gnd 0.0072f
C3828 vdd.n2771 gnd 0.0072f
C3829 vdd.n2772 gnd 0.0072f
C3830 vdd.n2774 gnd 0.898153f
C3831 vdd.n2776 gnd 0.0072f
C3832 vdd.n2777 gnd 0.0072f
C3833 vdd.n2778 gnd 0.017085f
C3834 vdd.n2779 gnd 0.015952f
C3835 vdd.n2780 gnd 0.015952f
C3836 vdd.n2781 gnd 0.898153f
C3837 vdd.n2782 gnd 0.015952f
C3838 vdd.n2783 gnd 0.015952f
C3839 vdd.n2784 gnd 0.0072f
C3840 vdd.n2785 gnd 0.0072f
C3841 vdd.n2786 gnd 0.0072f
C3842 vdd.n2787 gnd 0.459898f
C3843 vdd.n2788 gnd 0.0072f
C3844 vdd.n2789 gnd 0.0072f
C3845 vdd.n2790 gnd 0.0072f
C3846 vdd.n2791 gnd 0.0072f
C3847 vdd.n2792 gnd 0.0072f
C3848 vdd.n2793 gnd 0.573519f
C3849 vdd.n2794 gnd 0.0072f
C3850 vdd.n2795 gnd 0.0072f
C3851 vdd.n2796 gnd 0.0072f
C3852 vdd.n2797 gnd 0.0072f
C3853 vdd.n2798 gnd 0.0072f
C3854 vdd.n2799 gnd 0.735836f
C3855 vdd.n2800 gnd 0.0072f
C3856 vdd.n2801 gnd 0.0072f
C3857 vdd.n2802 gnd 0.0072f
C3858 vdd.n2803 gnd 0.0072f
C3859 vdd.n2804 gnd 0.0072f
C3860 vdd.n2805 gnd 0.405792f
C3861 vdd.n2806 gnd 0.0072f
C3862 vdd.n2807 gnd 0.0072f
C3863 vdd.n2808 gnd 0.0072f
C3864 vdd.n2809 gnd 0.0072f
C3865 vdd.n2810 gnd 0.0072f
C3866 vdd.n2811 gnd 0.232654f
C3867 vdd.n2812 gnd 0.0072f
C3868 vdd.n2813 gnd 0.0072f
C3869 vdd.n2814 gnd 0.0072f
C3870 vdd.n2815 gnd 0.0072f
C3871 vdd.n2816 gnd 0.0072f
C3872 vdd.n2817 gnd 0.422024f
C3873 vdd.n2818 gnd 0.0072f
C3874 vdd.n2819 gnd 0.0072f
C3875 vdd.n2820 gnd 0.0072f
C3876 vdd.n2821 gnd 0.0072f
C3877 vdd.n2822 gnd 0.0072f
C3878 vdd.n2823 gnd 0.58434f
C3879 vdd.n2824 gnd 0.0072f
C3880 vdd.n2825 gnd 0.0072f
C3881 vdd.n2826 gnd 0.0072f
C3882 vdd.n2827 gnd 0.0072f
C3883 vdd.n2828 gnd 0.0072f
C3884 vdd.n2829 gnd 0.654678f
C3885 vdd.n2830 gnd 0.0072f
C3886 vdd.n2831 gnd 0.0072f
C3887 vdd.n2832 gnd 0.0072f
C3888 vdd.n2833 gnd 0.0072f
C3889 vdd.n2834 gnd 0.0072f
C3890 vdd.n2835 gnd 0.492361f
C3891 vdd.n2836 gnd 0.0072f
C3892 vdd.n2837 gnd 0.0072f
C3893 vdd.n2838 gnd 0.0072f
C3894 vdd.t188 gnd 0.297837f
C3895 vdd.t186 gnd 0.189952f
C3896 vdd.t189 gnd 0.297837f
C3897 vdd.n2839 gnd 0.167396f
C3898 vdd.n2840 gnd 0.020858f
C3899 vdd.n2841 gnd 0.004447f
C3900 vdd.n2842 gnd 0.0072f
C3901 vdd.n2843 gnd 0.405792f
C3902 vdd.n2844 gnd 0.0072f
C3903 vdd.n2845 gnd 0.0072f
C3904 vdd.n2846 gnd 0.0072f
C3905 vdd.n2847 gnd 0.0072f
C3906 vdd.n2848 gnd 0.0072f
C3907 vdd.n2849 gnd 0.735836f
C3908 vdd.n2850 gnd 0.0072f
C3909 vdd.n2851 gnd 0.0072f
C3910 vdd.n2852 gnd 0.0072f
C3911 vdd.n2853 gnd 0.0072f
C3912 vdd.n2854 gnd 0.0072f
C3913 vdd.n2855 gnd 0.0072f
C3914 vdd.n2857 gnd 0.0072f
C3915 vdd.n2858 gnd 0.0072f
C3916 vdd.n2860 gnd 0.0072f
C3917 vdd.n2861 gnd 0.0072f
C3918 vdd.n2864 gnd 0.0072f
C3919 vdd.n2865 gnd 0.0072f
C3920 vdd.n2866 gnd 0.0072f
C3921 vdd.n2867 gnd 0.0072f
C3922 vdd.n2869 gnd 0.0072f
C3923 vdd.n2870 gnd 0.0072f
C3924 vdd.n2871 gnd 0.0072f
C3925 vdd.n2872 gnd 0.0072f
C3926 vdd.n2873 gnd 0.0072f
C3927 vdd.n2874 gnd 0.0072f
C3928 vdd.n2876 gnd 0.0072f
C3929 vdd.n2877 gnd 0.0072f
C3930 vdd.n2878 gnd 0.0072f
C3931 vdd.n2879 gnd 0.0072f
C3932 vdd.n2880 gnd 0.0072f
C3933 vdd.n2881 gnd 0.0072f
C3934 vdd.n2883 gnd 0.0072f
C3935 vdd.n2884 gnd 0.0072f
C3936 vdd.n2885 gnd 0.0072f
C3937 vdd.n2886 gnd 0.0072f
C3938 vdd.n2887 gnd 0.0072f
C3939 vdd.n2888 gnd 0.0072f
C3940 vdd.n2890 gnd 0.0072f
C3941 vdd.n2891 gnd 0.017085f
C3942 vdd.n2892 gnd 0.017085f
C3943 vdd.n2893 gnd 0.015952f
C3944 vdd.n2894 gnd 0.0072f
C3945 vdd.n2895 gnd 0.0072f
C3946 vdd.n2896 gnd 0.0072f
C3947 vdd.n2897 gnd 0.0072f
C3948 vdd.n2898 gnd 0.0072f
C3949 vdd.n2899 gnd 0.0072f
C3950 vdd.n2900 gnd 0.735836f
C3951 vdd.n2901 gnd 0.0072f
C3952 vdd.n2902 gnd 0.0072f
C3953 vdd.n2903 gnd 0.0072f
C3954 vdd.n2904 gnd 0.0072f
C3955 vdd.n2905 gnd 0.0072f
C3956 vdd.n2906 gnd 0.459898f
C3957 vdd.n2907 gnd 0.0072f
C3958 vdd.n2908 gnd 0.0072f
C3959 vdd.n2909 gnd 0.0072f
C3960 vdd.n2910 gnd 0.016828f
C3961 vdd.n2912 gnd 0.017085f
C3962 vdd.n2913 gnd 0.016208f
C3963 vdd.n2914 gnd 0.0072f
C3964 vdd.n2915 gnd 0.005559f
C3965 vdd.n2916 gnd 0.0072f
C3966 vdd.n2918 gnd 0.0072f
C3967 vdd.n2919 gnd 0.0072f
C3968 vdd.n2920 gnd 0.0072f
C3969 vdd.n2921 gnd 0.0072f
C3970 vdd.n2922 gnd 0.0072f
C3971 vdd.n2923 gnd 0.0072f
C3972 vdd.n2925 gnd 0.0072f
C3973 vdd.n2926 gnd 0.0072f
C3974 vdd.n2927 gnd 0.0072f
C3975 vdd.n2928 gnd 0.0072f
C3976 vdd.n2929 gnd 0.0072f
C3977 vdd.n2930 gnd 0.0072f
C3978 vdd.n2932 gnd 0.0072f
C3979 vdd.n2933 gnd 0.0072f
C3980 vdd.n2934 gnd 0.0072f
C3981 vdd.n2935 gnd 0.0072f
C3982 vdd.n2936 gnd 0.0072f
C3983 vdd.n2937 gnd 0.0072f
C3984 vdd.n2939 gnd 0.0072f
C3985 vdd.n2940 gnd 0.0072f
C3986 vdd.n2941 gnd 0.0072f
C3987 vdd.n2942 gnd 0.640844f
C3988 vdd.n2943 gnd 0.017303f
C3989 vdd.n2944 gnd 0.0072f
C3990 vdd.n2945 gnd 0.0072f
C3991 vdd.n2947 gnd 0.0072f
C3992 vdd.n2948 gnd 0.0072f
C3993 vdd.n2949 gnd 0.0072f
C3994 vdd.n2950 gnd 0.0072f
C3995 vdd.n2951 gnd 0.0072f
C3996 vdd.n2952 gnd 0.0072f
C3997 vdd.n2954 gnd 0.0072f
C3998 vdd.n2955 gnd 0.0072f
C3999 vdd.n2956 gnd 0.0072f
C4000 vdd.n2957 gnd 0.0072f
C4001 vdd.n2958 gnd 0.0072f
C4002 vdd.n2959 gnd 0.0072f
C4003 vdd.n2961 gnd 0.0072f
C4004 vdd.n2962 gnd 0.0072f
C4005 vdd.n2963 gnd 0.0072f
C4006 vdd.n2964 gnd 0.0072f
C4007 vdd.n2965 gnd 0.0072f
C4008 vdd.n2966 gnd 0.0072f
C4009 vdd.n2968 gnd 0.0072f
C4010 vdd.n2969 gnd 0.0072f
C4011 vdd.n2971 gnd 0.0072f
C4012 vdd.n2972 gnd 0.0072f
C4013 vdd.n2973 gnd 0.017085f
C4014 vdd.n2974 gnd 0.015952f
C4015 vdd.n2975 gnd 0.015952f
C4016 vdd.n2976 gnd 1.06047f
C4017 vdd.n2977 gnd 0.015952f
C4018 vdd.n2978 gnd 0.017085f
C4019 vdd.n2979 gnd 0.016208f
C4020 vdd.n2980 gnd 0.0072f
C4021 vdd.n2981 gnd 0.005559f
C4022 vdd.n2982 gnd 0.0072f
C4023 vdd.n2984 gnd 0.0072f
C4024 vdd.n2985 gnd 0.0072f
C4025 vdd.n2986 gnd 0.0072f
C4026 vdd.n2987 gnd 0.0072f
C4027 vdd.n2988 gnd 0.0072f
C4028 vdd.n2989 gnd 0.0072f
C4029 vdd.n2991 gnd 0.0072f
C4030 vdd.n2992 gnd 0.0072f
C4031 vdd.n2993 gnd 0.0072f
C4032 vdd.n2994 gnd 0.0072f
C4033 vdd.n2995 gnd 0.0072f
C4034 vdd.n2996 gnd 0.0072f
C4035 vdd.n2998 gnd 0.0072f
C4036 vdd.n2999 gnd 0.0072f
C4037 vdd.n3000 gnd 0.0072f
C4038 vdd.n3001 gnd 0.0072f
C4039 vdd.n3002 gnd 0.0072f
C4040 vdd.n3003 gnd 0.0072f
C4041 vdd.n3005 gnd 0.0072f
C4042 vdd.n3006 gnd 0.0072f
C4043 vdd.n3008 gnd 0.0072f
C4044 vdd.n3009 gnd 0.017303f
C4045 vdd.n3010 gnd 0.640844f
C4046 vdd.n3011 gnd 0.009106f
C4047 vdd.n3012 gnd 0.004048f
C4048 vdd.t232 gnd 0.130268f
C4049 vdd.t233 gnd 0.139221f
C4050 vdd.t231 gnd 0.170129f
C4051 vdd.n3013 gnd 0.218081f
C4052 vdd.n3014 gnd 0.183228f
C4053 vdd.n3015 gnd 0.013125f
C4054 vdd.n3016 gnd 0.010589f
C4055 vdd.n3017 gnd 0.004474f
C4056 vdd.n3018 gnd 0.008523f
C4057 vdd.n3019 gnd 0.010589f
C4058 vdd.n3020 gnd 0.010589f
C4059 vdd.n3021 gnd 0.008523f
C4060 vdd.n3022 gnd 0.008523f
C4061 vdd.n3023 gnd 0.010589f
C4062 vdd.n3025 gnd 0.010589f
C4063 vdd.n3026 gnd 0.008523f
C4064 vdd.n3027 gnd 0.008523f
C4065 vdd.n3028 gnd 0.008523f
C4066 vdd.n3029 gnd 0.010589f
C4067 vdd.n3031 gnd 0.010589f
C4068 vdd.n3033 gnd 0.010589f
C4069 vdd.n3034 gnd 0.008523f
C4070 vdd.n3035 gnd 0.008523f
C4071 vdd.n3036 gnd 0.008523f
C4072 vdd.n3037 gnd 0.010589f
C4073 vdd.n3039 gnd 0.010589f
C4074 vdd.n3041 gnd 0.010589f
C4075 vdd.n3042 gnd 0.008523f
C4076 vdd.n3043 gnd 0.008523f
C4077 vdd.n3044 gnd 0.008523f
C4078 vdd.n3045 gnd 0.010589f
C4079 vdd.n3047 gnd 0.010589f
C4080 vdd.n3048 gnd 0.010589f
C4081 vdd.n3049 gnd 0.008523f
C4082 vdd.n3050 gnd 0.008523f
C4083 vdd.n3051 gnd 0.010589f
C4084 vdd.n3052 gnd 0.010589f
C4085 vdd.n3054 gnd 0.010589f
C4086 vdd.n3055 gnd 0.008523f
C4087 vdd.n3056 gnd 0.010589f
C4088 vdd.n3057 gnd 0.010589f
C4089 vdd.n3058 gnd 0.010589f
C4090 vdd.n3059 gnd 0.017386f
C4091 vdd.n3060 gnd 0.005795f
C4092 vdd.n3061 gnd 0.010589f
C4093 vdd.n3063 gnd 0.010589f
C4094 vdd.n3065 gnd 0.010589f
C4095 vdd.n3066 gnd 0.008523f
C4096 vdd.n3067 gnd 0.008523f
C4097 vdd.n3068 gnd 0.008523f
C4098 vdd.n3069 gnd 0.010589f
C4099 vdd.n3071 gnd 0.010589f
C4100 vdd.n3073 gnd 0.010589f
C4101 vdd.n3074 gnd 0.008523f
C4102 vdd.n3075 gnd 0.008523f
C4103 vdd.n3076 gnd 0.008523f
C4104 vdd.n3077 gnd 0.010589f
C4105 vdd.n3079 gnd 0.010589f
C4106 vdd.n3081 gnd 0.010589f
C4107 vdd.n3082 gnd 0.008523f
C4108 vdd.n3083 gnd 0.008523f
C4109 vdd.n3084 gnd 0.008523f
C4110 vdd.n3085 gnd 0.010589f
C4111 vdd.n3087 gnd 0.010589f
C4112 vdd.n3089 gnd 0.010589f
C4113 vdd.n3090 gnd 0.008523f
C4114 vdd.n3091 gnd 0.008523f
C4115 vdd.n3092 gnd 0.008523f
C4116 vdd.n3093 gnd 0.010589f
C4117 vdd.n3095 gnd 0.010589f
C4118 vdd.n3097 gnd 0.010589f
C4119 vdd.n3098 gnd 0.008523f
C4120 vdd.n3099 gnd 0.008523f
C4121 vdd.n3100 gnd 0.007116f
C4122 vdd.n3101 gnd 0.010589f
C4123 vdd.n3103 gnd 0.010589f
C4124 vdd.n3105 gnd 0.010589f
C4125 vdd.n3106 gnd 0.007116f
C4126 vdd.n3107 gnd 0.008523f
C4127 vdd.n3108 gnd 0.008523f
C4128 vdd.n3109 gnd 0.010589f
C4129 vdd.n3111 gnd 0.010589f
C4130 vdd.n3113 gnd 0.010589f
C4131 vdd.n3114 gnd 0.008523f
C4132 vdd.n3115 gnd 0.008523f
C4133 vdd.n3116 gnd 0.008523f
C4134 vdd.n3117 gnd 0.010589f
C4135 vdd.n3119 gnd 0.010589f
C4136 vdd.n3121 gnd 0.010589f
C4137 vdd.n3122 gnd 0.008523f
C4138 vdd.n3123 gnd 0.008523f
C4139 vdd.n3124 gnd 0.008523f
C4140 vdd.n3125 gnd 0.010589f
C4141 vdd.n3127 gnd 0.010589f
C4142 vdd.n3128 gnd 0.010589f
C4143 vdd.n3129 gnd 0.008523f
C4144 vdd.n3130 gnd 0.008523f
C4145 vdd.n3131 gnd 0.010589f
C4146 vdd.n3132 gnd 0.010589f
C4147 vdd.n3133 gnd 0.008523f
C4148 vdd.n3134 gnd 0.008523f
C4149 vdd.n3135 gnd 0.010589f
C4150 vdd.n3136 gnd 0.010589f
C4151 vdd.n3138 gnd 0.010589f
C4152 vdd.n3139 gnd 0.008523f
C4153 vdd.n3140 gnd 0.007074f
C4154 vdd.n3141 gnd 0.024278f
C4155 vdd.n3142 gnd 0.024113f
C4156 vdd.n3143 gnd 0.007074f
C4157 vdd.n3144 gnd 0.024113f
C4158 vdd.n3145 gnd 1.42839f
C4159 vdd.n3146 gnd 0.024113f
C4160 vdd.n3147 gnd 0.007074f
C4161 vdd.n3148 gnd 0.024113f
C4162 vdd.n3149 gnd 0.010589f
C4163 vdd.n3150 gnd 0.010589f
C4164 vdd.n3151 gnd 0.008523f
C4165 vdd.n3152 gnd 0.010589f
C4166 vdd.n3153 gnd 1.0226f
C4167 vdd.n3154 gnd 0.010589f
C4168 vdd.n3155 gnd 0.008523f
C4169 vdd.n3156 gnd 0.010589f
C4170 vdd.n3157 gnd 0.010589f
C4171 vdd.n3158 gnd 0.010589f
C4172 vdd.n3159 gnd 0.008523f
C4173 vdd.n3160 gnd 0.010589f
C4174 vdd.n3161 gnd 1.05506f
C4175 vdd.n3162 gnd 0.010589f
C4176 vdd.n3163 gnd 0.008523f
C4177 vdd.n3164 gnd 0.010589f
C4178 vdd.n3165 gnd 0.010589f
C4179 vdd.n3166 gnd 0.010589f
C4180 vdd.n3167 gnd 0.008523f
C4181 vdd.n3168 gnd 0.010589f
C4182 vdd.t88 gnd 0.541056f
C4183 vdd.n3169 gnd 0.8711f
C4184 vdd.n3170 gnd 0.010589f
C4185 vdd.n3171 gnd 0.008523f
C4186 vdd.n3172 gnd 0.010589f
C4187 vdd.n3173 gnd 0.010589f
C4188 vdd.n3174 gnd 0.010589f
C4189 vdd.n3175 gnd 0.008523f
C4190 vdd.n3176 gnd 0.010589f
C4191 vdd.n3177 gnd 0.687141f
C4192 vdd.n3178 gnd 0.010589f
C4193 vdd.n3179 gnd 0.008523f
C4194 vdd.n3180 gnd 0.010589f
C4195 vdd.n3181 gnd 0.010589f
C4196 vdd.n3182 gnd 0.010589f
C4197 vdd.n3183 gnd 0.008523f
C4198 vdd.n3184 gnd 0.010589f
C4199 vdd.n3185 gnd 0.860279f
C4200 vdd.n3186 gnd 0.57893f
C4201 vdd.n3187 gnd 0.010589f
C4202 vdd.n3188 gnd 0.008523f
C4203 vdd.n3189 gnd 0.010589f
C4204 vdd.n3190 gnd 0.010589f
C4205 vdd.n3191 gnd 0.010589f
C4206 vdd.n3192 gnd 0.008523f
C4207 vdd.n3193 gnd 0.010589f
C4208 vdd.n3194 gnd 0.762889f
C4209 vdd.n3195 gnd 0.010589f
C4210 vdd.n3196 gnd 0.008523f
C4211 vdd.n3197 gnd 0.010589f
C4212 vdd.n3198 gnd 0.010589f
C4213 vdd.n3199 gnd 0.010589f
C4214 vdd.n3200 gnd 0.010589f
C4215 vdd.n3201 gnd 0.010589f
C4216 vdd.n3202 gnd 0.008523f
C4217 vdd.n3203 gnd 0.008523f
C4218 vdd.n3204 gnd 0.010589f
C4219 vdd.t43 gnd 0.541056f
C4220 vdd.n3205 gnd 0.898153f
C4221 vdd.n3206 gnd 0.010589f
C4222 vdd.n3207 gnd 0.008523f
C4223 vdd.n3208 gnd 0.010589f
C4224 vdd.n3209 gnd 0.010589f
C4225 vdd.n3210 gnd 0.010589f
C4226 vdd.n3211 gnd 0.008523f
C4227 vdd.n3212 gnd 0.010589f
C4228 vdd.n3213 gnd 0.849458f
C4229 vdd.n3214 gnd 0.010589f
C4230 vdd.n3215 gnd 0.010589f
C4231 vdd.n3216 gnd 0.008523f
C4232 vdd.n3217 gnd 0.008523f
C4233 vdd.n3218 gnd 0.008523f
C4234 vdd.n3219 gnd 0.010589f
C4235 vdd.n3220 gnd 0.010589f
C4236 vdd.n3221 gnd 0.010589f
C4237 vdd.n3222 gnd 0.010589f
C4238 vdd.n3223 gnd 0.008523f
C4239 vdd.n3224 gnd 0.008523f
C4240 vdd.n3225 gnd 0.008523f
C4241 vdd.n3226 gnd 0.010589f
C4242 vdd.n3227 gnd 0.010589f
C4243 vdd.n3228 gnd 0.010589f
C4244 vdd.n3229 gnd 0.010589f
C4245 vdd.n3230 gnd 0.008523f
C4246 vdd.n3231 gnd 0.008523f
C4247 vdd.n3232 gnd 0.008523f
C4248 vdd.n3233 gnd 0.010589f
C4249 vdd.n3234 gnd 0.010589f
C4250 vdd.n3235 gnd 0.010589f
C4251 vdd.n3236 gnd 0.898153f
C4252 vdd.n3237 gnd 0.010589f
C4253 vdd.n3238 gnd 0.008523f
C4254 vdd.n3239 gnd 0.008523f
C4255 vdd.n3240 gnd 0.008523f
C4256 vdd.n3241 gnd 0.010589f
C4257 vdd.n3242 gnd 0.010589f
C4258 vdd.n3243 gnd 0.010589f
C4259 vdd.n3244 gnd 0.010589f
C4260 vdd.n3245 gnd 0.008523f
C4261 vdd.n3246 gnd 0.008523f
C4262 vdd.n3247 gnd 0.007074f
C4263 vdd.n3248 gnd 0.024113f
C4264 vdd.n3249 gnd 0.024278f
C4265 vdd.n3250 gnd 0.004048f
C4266 vdd.n3251 gnd 0.024278f
C4267 vdd.n3253 gnd 2.39147f
C4268 vdd.n3254 gnd 1.42839f
C4269 vdd.n3255 gnd 0.708783f
C4270 vdd.n3256 gnd 0.010589f
C4271 vdd.n3257 gnd 0.008523f
C4272 vdd.n3258 gnd 0.008523f
C4273 vdd.n3259 gnd 0.008523f
C4274 vdd.n3260 gnd 0.010589f
C4275 vdd.n3261 gnd 1.08211f
C4276 vdd.n3262 gnd 1.08211f
C4277 vdd.n3263 gnd 0.622214f
C4278 vdd.n3264 gnd 0.010589f
C4279 vdd.n3265 gnd 0.008523f
C4280 vdd.n3266 gnd 0.008523f
C4281 vdd.n3267 gnd 0.008523f
C4282 vdd.n3268 gnd 0.010589f
C4283 vdd.n3269 gnd 0.643857f
C4284 vdd.n3270 gnd 0.795352f
C4285 vdd.t61 gnd 0.541056f
C4286 vdd.n3271 gnd 0.827816f
C4287 vdd.n3272 gnd 0.010589f
C4288 vdd.n3273 gnd 0.008523f
C4289 vdd.n3274 gnd 0.008523f
C4290 vdd.n3275 gnd 0.008523f
C4291 vdd.n3276 gnd 0.010589f
C4292 vdd.n3277 gnd 0.898153f
C4293 vdd.t37 gnd 0.541056f
C4294 vdd.n3278 gnd 0.654678f
C4295 vdd.n3279 gnd 0.784531f
C4296 vdd.n3280 gnd 0.010589f
C4297 vdd.n3281 gnd 0.008523f
C4298 vdd.n3282 gnd 0.008523f
C4299 vdd.n3283 gnd 0.008523f
C4300 vdd.n3284 gnd 0.010589f
C4301 vdd.n3285 gnd 0.600572f
C4302 vdd.t29 gnd 0.541056f
C4303 vdd.n3286 gnd 0.898153f
C4304 vdd.t65 gnd 0.541056f
C4305 vdd.n3287 gnd 0.665499f
C4306 vdd.n3288 gnd 0.010589f
C4307 vdd.n3289 gnd 0.008523f
C4308 vdd.n3290 gnd 0.008138f
C4309 vdd.n3291 gnd 0.62456f
C4310 vdd.n3292 gnd 2.52091f
C4311 a_n6972_8799.n0 gnd 0.207737f
C4312 a_n6972_8799.n1 gnd 0.290352f
C4313 a_n6972_8799.n2 gnd 0.207737f
C4314 a_n6972_8799.n3 gnd 0.207737f
C4315 a_n6972_8799.n4 gnd 0.207737f
C4316 a_n6972_8799.n5 gnd 0.273684f
C4317 a_n6972_8799.n6 gnd 0.207737f
C4318 a_n6972_8799.n7 gnd 0.290352f
C4319 a_n6972_8799.n8 gnd 0.207737f
C4320 a_n6972_8799.n9 gnd 0.207737f
C4321 a_n6972_8799.n10 gnd 0.207737f
C4322 a_n6972_8799.n11 gnd 0.273684f
C4323 a_n6972_8799.n12 gnd 0.207737f
C4324 a_n6972_8799.n13 gnd 0.455038f
C4325 a_n6972_8799.n14 gnd 0.207737f
C4326 a_n6972_8799.n15 gnd 0.207737f
C4327 a_n6972_8799.n16 gnd 0.207737f
C4328 a_n6972_8799.n17 gnd 0.273684f
C4329 a_n6972_8799.n18 gnd 0.325619f
C4330 a_n6972_8799.n19 gnd 0.207737f
C4331 a_n6972_8799.n20 gnd 0.207737f
C4332 a_n6972_8799.n21 gnd 0.207737f
C4333 a_n6972_8799.n22 gnd 0.207737f
C4334 a_n6972_8799.n23 gnd 0.238418f
C4335 a_n6972_8799.n24 gnd 0.325619f
C4336 a_n6972_8799.n25 gnd 0.207737f
C4337 a_n6972_8799.n26 gnd 0.207737f
C4338 a_n6972_8799.n27 gnd 0.207737f
C4339 a_n6972_8799.n28 gnd 0.207737f
C4340 a_n6972_8799.n29 gnd 0.238418f
C4341 a_n6972_8799.n30 gnd 0.325619f
C4342 a_n6972_8799.n31 gnd 0.207737f
C4343 a_n6972_8799.n32 gnd 0.207737f
C4344 a_n6972_8799.n33 gnd 0.207737f
C4345 a_n6972_8799.n34 gnd 0.207737f
C4346 a_n6972_8799.n35 gnd 0.403104f
C4347 a_n6972_8799.n36 gnd 4.02811f
C4348 a_n6972_8799.n37 gnd 2.79029f
C4349 a_n6972_8799.n38 gnd 0.363145f
C4350 a_n6972_8799.n39 gnd 3.04349f
C4351 a_n6972_8799.n40 gnd 0.363144f
C4352 a_n6972_8799.n41 gnd 0.8559f
C4353 a_n6972_8799.n42 gnd 0.008616f
C4354 a_n6972_8799.n43 gnd 0.001157f
C4355 a_n6972_8799.n45 gnd 0.007738f
C4356 a_n6972_8799.n46 gnd 0.011695f
C4357 a_n6972_8799.n47 gnd 0.008043f
C4358 a_n6972_8799.n49 gnd 4.02e-19
C4359 a_n6972_8799.n50 gnd 0.008335f
C4360 a_n6972_8799.n51 gnd 0.011513f
C4361 a_n6972_8799.n52 gnd 0.007418f
C4362 a_n6972_8799.n53 gnd 0.008616f
C4363 a_n6972_8799.n54 gnd 0.001157f
C4364 a_n6972_8799.n56 gnd 0.007738f
C4365 a_n6972_8799.n57 gnd 0.011695f
C4366 a_n6972_8799.n58 gnd 0.008043f
C4367 a_n6972_8799.n60 gnd 4.02e-19
C4368 a_n6972_8799.n61 gnd 0.008335f
C4369 a_n6972_8799.n62 gnd 0.011513f
C4370 a_n6972_8799.n63 gnd 0.007418f
C4371 a_n6972_8799.n64 gnd 0.008616f
C4372 a_n6972_8799.n65 gnd 0.001157f
C4373 a_n6972_8799.n67 gnd 0.007738f
C4374 a_n6972_8799.n68 gnd 0.011695f
C4375 a_n6972_8799.n69 gnd 0.008043f
C4376 a_n6972_8799.n71 gnd 4.02e-19
C4377 a_n6972_8799.n72 gnd 0.008335f
C4378 a_n6972_8799.n73 gnd 0.011513f
C4379 a_n6972_8799.n74 gnd 0.007418f
C4380 a_n6972_8799.n75 gnd 0.001157f
C4381 a_n6972_8799.n77 gnd 0.007738f
C4382 a_n6972_8799.n78 gnd 0.011695f
C4383 a_n6972_8799.n79 gnd 0.008043f
C4384 a_n6972_8799.n81 gnd 4.02e-19
C4385 a_n6972_8799.n82 gnd 0.008335f
C4386 a_n6972_8799.n83 gnd 0.011513f
C4387 a_n6972_8799.n84 gnd 0.007418f
C4388 a_n6972_8799.n85 gnd 0.250096f
C4389 a_n6972_8799.n86 gnd 0.001157f
C4390 a_n6972_8799.n88 gnd 0.007738f
C4391 a_n6972_8799.n89 gnd 0.011695f
C4392 a_n6972_8799.n90 gnd 0.008043f
C4393 a_n6972_8799.n92 gnd 4.02e-19
C4394 a_n6972_8799.n93 gnd 0.008335f
C4395 a_n6972_8799.n94 gnd 0.011513f
C4396 a_n6972_8799.n95 gnd 0.007418f
C4397 a_n6972_8799.n96 gnd 0.250096f
C4398 a_n6972_8799.n97 gnd 0.001157f
C4399 a_n6972_8799.n99 gnd 0.007738f
C4400 a_n6972_8799.n100 gnd 0.011695f
C4401 a_n6972_8799.n101 gnd 0.008043f
C4402 a_n6972_8799.n103 gnd 4.02e-19
C4403 a_n6972_8799.n104 gnd 0.008335f
C4404 a_n6972_8799.n105 gnd 0.011513f
C4405 a_n6972_8799.n106 gnd 0.007418f
C4406 a_n6972_8799.n107 gnd 0.250096f
C4407 a_n6972_8799.t4 gnd 0.144089f
C4408 a_n6972_8799.t33 gnd 0.144089f
C4409 a_n6972_8799.t34 gnd 0.144089f
C4410 a_n6972_8799.n108 gnd 1.13645f
C4411 a_n6972_8799.t10 gnd 0.144089f
C4412 a_n6972_8799.t5 gnd 0.144089f
C4413 a_n6972_8799.n109 gnd 1.13457f
C4414 a_n6972_8799.t7 gnd 0.144089f
C4415 a_n6972_8799.t9 gnd 0.144089f
C4416 a_n6972_8799.n110 gnd 1.13645f
C4417 a_n6972_8799.t8 gnd 0.144089f
C4418 a_n6972_8799.t2 gnd 0.144089f
C4419 a_n6972_8799.n111 gnd 1.13457f
C4420 a_n6972_8799.t11 gnd 0.144089f
C4421 a_n6972_8799.t12 gnd 0.144089f
C4422 a_n6972_8799.n112 gnd 1.13457f
C4423 a_n6972_8799.t22 gnd 0.112069f
C4424 a_n6972_8799.t27 gnd 0.112069f
C4425 a_n6972_8799.n113 gnd 0.993201f
C4426 a_n6972_8799.t1 gnd 0.112069f
C4427 a_n6972_8799.t13 gnd 0.112069f
C4428 a_n6972_8799.n114 gnd 0.990281f
C4429 a_n6972_8799.n115 gnd 0.878129f
C4430 a_n6972_8799.t20 gnd 0.112069f
C4431 a_n6972_8799.t18 gnd 0.112069f
C4432 a_n6972_8799.n116 gnd 0.990281f
C4433 a_n6972_8799.t15 gnd 0.112069f
C4434 a_n6972_8799.t3 gnd 0.112069f
C4435 a_n6972_8799.n117 gnd 0.9932f
C4436 a_n6972_8799.t6 gnd 0.112069f
C4437 a_n6972_8799.t21 gnd 0.112069f
C4438 a_n6972_8799.n118 gnd 0.99028f
C4439 a_n6972_8799.n119 gnd 0.878131f
C4440 a_n6972_8799.t17 gnd 0.112069f
C4441 a_n6972_8799.t26 gnd 0.112069f
C4442 a_n6972_8799.n120 gnd 0.99028f
C4443 a_n6972_8799.t16 gnd 0.112069f
C4444 a_n6972_8799.t14 gnd 0.112069f
C4445 a_n6972_8799.n121 gnd 0.9932f
C4446 a_n6972_8799.t32 gnd 0.112069f
C4447 a_n6972_8799.t24 gnd 0.112069f
C4448 a_n6972_8799.n122 gnd 0.99028f
C4449 a_n6972_8799.n123 gnd 0.878131f
C4450 a_n6972_8799.t31 gnd 0.112069f
C4451 a_n6972_8799.t23 gnd 0.112069f
C4452 a_n6972_8799.n124 gnd 0.99028f
C4453 a_n6972_8799.t35 gnd 0.112069f
C4454 a_n6972_8799.t25 gnd 0.112069f
C4455 a_n6972_8799.n125 gnd 0.990281f
C4456 a_n6972_8799.n126 gnd 3.08917f
C4457 a_n6972_8799.t19 gnd 0.112069f
C4458 a_n6972_8799.t28 gnd 0.112069f
C4459 a_n6972_8799.n127 gnd 0.990281f
C4460 a_n6972_8799.n128 gnd 0.432365f
C4461 a_n6972_8799.t30 gnd 0.112069f
C4462 a_n6972_8799.t29 gnd 0.112069f
C4463 a_n6972_8799.n129 gnd 0.990281f
C4464 a_n6972_8799.t114 gnd 0.597459f
C4465 a_n6972_8799.n130 gnd 0.267109f
C4466 a_n6972_8799.t47 gnd 0.597459f
C4467 a_n6972_8799.t65 gnd 0.597459f
C4468 a_n6972_8799.n131 gnd 0.270418f
C4469 a_n6972_8799.t83 gnd 0.597459f
C4470 a_n6972_8799.t100 gnd 0.597459f
C4471 a_n6972_8799.t101 gnd 0.597459f
C4472 a_n6972_8799.n132 gnd 0.272502f
C4473 a_n6972_8799.t68 gnd 0.597459f
C4474 a_n6972_8799.t78 gnd 0.597459f
C4475 a_n6972_8799.n133 gnd 0.266036f
C4476 a_n6972_8799.t115 gnd 0.608767f
C4477 a_n6972_8799.n134 gnd 0.250481f
C4478 a_n6972_8799.n135 gnd 0.011785f
C4479 a_n6972_8799.t77 gnd 0.597459f
C4480 a_n6972_8799.n136 gnd 0.266837f
C4481 a_n6972_8799.n137 gnd 0.270404f
C4482 a_n6972_8799.t69 gnd 0.597459f
C4483 a_n6972_8799.n138 gnd 0.266926f
C4484 a_n6972_8799.n139 gnd 0.261553f
C4485 a_n6972_8799.t37 gnd 0.597459f
C4486 a_n6972_8799.n140 gnd 0.266676f
C4487 a_n6972_8799.n141 gnd 0.272936f
C4488 a_n6972_8799.t117 gnd 0.597459f
C4489 a_n6972_8799.n142 gnd 0.270286f
C4490 a_n6972_8799.n143 gnd 0.266356f
C4491 a_n6972_8799.t64 gnd 0.597459f
C4492 a_n6972_8799.n144 gnd 0.261873f
C4493 a_n6972_8799.t46 gnd 0.597459f
C4494 a_n6972_8799.n145 gnd 0.270403f
C4495 a_n6972_8799.t45 gnd 0.608756f
C4496 a_n6972_8799.t124 gnd 0.597459f
C4497 a_n6972_8799.n146 gnd 0.267109f
C4498 a_n6972_8799.t61 gnd 0.597459f
C4499 a_n6972_8799.t74 gnd 0.597459f
C4500 a_n6972_8799.n147 gnd 0.270418f
C4501 a_n6972_8799.t94 gnd 0.597459f
C4502 a_n6972_8799.t109 gnd 0.597459f
C4503 a_n6972_8799.t113 gnd 0.597459f
C4504 a_n6972_8799.n148 gnd 0.272502f
C4505 a_n6972_8799.t75 gnd 0.597459f
C4506 a_n6972_8799.t84 gnd 0.597459f
C4507 a_n6972_8799.n149 gnd 0.266036f
C4508 a_n6972_8799.t125 gnd 0.608767f
C4509 a_n6972_8799.n150 gnd 0.250481f
C4510 a_n6972_8799.n151 gnd 0.011785f
C4511 a_n6972_8799.t85 gnd 0.597459f
C4512 a_n6972_8799.n152 gnd 0.266837f
C4513 a_n6972_8799.n153 gnd 0.270404f
C4514 a_n6972_8799.t76 gnd 0.597459f
C4515 a_n6972_8799.n154 gnd 0.266926f
C4516 a_n6972_8799.n155 gnd 0.261553f
C4517 a_n6972_8799.t48 gnd 0.597459f
C4518 a_n6972_8799.n156 gnd 0.266676f
C4519 a_n6972_8799.n157 gnd 0.272936f
C4520 a_n6972_8799.t129 gnd 0.597459f
C4521 a_n6972_8799.n158 gnd 0.270286f
C4522 a_n6972_8799.n159 gnd 0.266356f
C4523 a_n6972_8799.t73 gnd 0.597459f
C4524 a_n6972_8799.n160 gnd 0.261873f
C4525 a_n6972_8799.t55 gnd 0.597459f
C4526 a_n6972_8799.n161 gnd 0.270403f
C4527 a_n6972_8799.t59 gnd 0.608756f
C4528 a_n6972_8799.n162 gnd 0.899839f
C4529 a_n6972_8799.t91 gnd 0.597459f
C4530 a_n6972_8799.n163 gnd 0.267109f
C4531 a_n6972_8799.t111 gnd 0.597459f
C4532 a_n6972_8799.t44 gnd 0.597459f
C4533 a_n6972_8799.n164 gnd 0.270418f
C4534 a_n6972_8799.t97 gnd 0.597459f
C4535 a_n6972_8799.t127 gnd 0.597459f
C4536 a_n6972_8799.t88 gnd 0.597459f
C4537 a_n6972_8799.n165 gnd 0.272502f
C4538 a_n6972_8799.t121 gnd 0.597459f
C4539 a_n6972_8799.t54 gnd 0.597459f
C4540 a_n6972_8799.n166 gnd 0.266036f
C4541 a_n6972_8799.t118 gnd 0.608767f
C4542 a_n6972_8799.n167 gnd 0.250481f
C4543 a_n6972_8799.n168 gnd 0.011785f
C4544 a_n6972_8799.t39 gnd 0.597459f
C4545 a_n6972_8799.n169 gnd 0.266837f
C4546 a_n6972_8799.n170 gnd 0.270404f
C4547 a_n6972_8799.t103 gnd 0.597459f
C4548 a_n6972_8799.n171 gnd 0.266926f
C4549 a_n6972_8799.n172 gnd 0.261553f
C4550 a_n6972_8799.t82 gnd 0.597459f
C4551 a_n6972_8799.n173 gnd 0.266676f
C4552 a_n6972_8799.n174 gnd 0.272936f
C4553 a_n6972_8799.t60 gnd 0.597459f
C4554 a_n6972_8799.n175 gnd 0.270286f
C4555 a_n6972_8799.n176 gnd 0.266356f
C4556 a_n6972_8799.t67 gnd 0.597459f
C4557 a_n6972_8799.n177 gnd 0.261873f
C4558 a_n6972_8799.t50 gnd 0.597459f
C4559 a_n6972_8799.n178 gnd 0.270403f
C4560 a_n6972_8799.t131 gnd 0.608756f
C4561 a_n6972_8799.n179 gnd 1.53901f
C4562 a_n6972_8799.t80 gnd 0.597459f
C4563 a_n6972_8799.t79 gnd 0.597459f
C4564 a_n6972_8799.t58 gnd 0.597459f
C4565 a_n6972_8799.n180 gnd 0.270005f
C4566 a_n6972_8799.t116 gnd 0.597459f
C4567 a_n6972_8799.t81 gnd 0.597459f
C4568 a_n6972_8799.t63 gnd 0.597459f
C4569 a_n6972_8799.n181 gnd 0.266926f
C4570 a_n6972_8799.t119 gnd 0.597459f
C4571 a_n6972_8799.t95 gnd 0.597459f
C4572 a_n6972_8799.t93 gnd 0.597459f
C4573 a_n6972_8799.n182 gnd 0.270418f
C4574 a_n6972_8799.t40 gnd 0.597459f
C4575 a_n6972_8799.t99 gnd 0.597459f
C4576 a_n6972_8799.t98 gnd 0.597459f
C4577 a_n6972_8799.n183 gnd 0.266356f
C4578 a_n6972_8799.t42 gnd 0.597459f
C4579 a_n6972_8799.t41 gnd 0.597459f
C4580 a_n6972_8799.t112 gnd 0.597459f
C4581 a_n6972_8799.n184 gnd 0.270403f
C4582 a_n6972_8799.t57 gnd 0.608767f
C4583 a_n6972_8799.n185 gnd 0.250481f
C4584 a_n6972_8799.n186 gnd 0.267109f
C4585 a_n6972_8799.n187 gnd 0.261873f
C4586 a_n6972_8799.n188 gnd 0.270286f
C4587 a_n6972_8799.n189 gnd 0.272936f
C4588 a_n6972_8799.n190 gnd 0.266676f
C4589 a_n6972_8799.n191 gnd 0.261553f
C4590 a_n6972_8799.n192 gnd 0.270404f
C4591 a_n6972_8799.n193 gnd 0.272502f
C4592 a_n6972_8799.n194 gnd 0.266036f
C4593 a_n6972_8799.n195 gnd 0.261393f
C4594 a_n6972_8799.t87 gnd 0.597459f
C4595 a_n6972_8799.t86 gnd 0.597459f
C4596 a_n6972_8799.t70 gnd 0.597459f
C4597 a_n6972_8799.n196 gnd 0.270005f
C4598 a_n6972_8799.t128 gnd 0.597459f
C4599 a_n6972_8799.t92 gnd 0.597459f
C4600 a_n6972_8799.t72 gnd 0.597459f
C4601 a_n6972_8799.n197 gnd 0.266926f
C4602 a_n6972_8799.t36 gnd 0.597459f
C4603 a_n6972_8799.t105 gnd 0.597459f
C4604 a_n6972_8799.t104 gnd 0.597459f
C4605 a_n6972_8799.n198 gnd 0.270418f
C4606 a_n6972_8799.t49 gnd 0.597459f
C4607 a_n6972_8799.t108 gnd 0.597459f
C4608 a_n6972_8799.t107 gnd 0.597459f
C4609 a_n6972_8799.n199 gnd 0.266356f
C4610 a_n6972_8799.t53 gnd 0.597459f
C4611 a_n6972_8799.t52 gnd 0.597459f
C4612 a_n6972_8799.t123 gnd 0.597459f
C4613 a_n6972_8799.n200 gnd 0.270403f
C4614 a_n6972_8799.t71 gnd 0.608767f
C4615 a_n6972_8799.n201 gnd 0.250481f
C4616 a_n6972_8799.n202 gnd 0.267109f
C4617 a_n6972_8799.n203 gnd 0.261873f
C4618 a_n6972_8799.n204 gnd 0.270286f
C4619 a_n6972_8799.n205 gnd 0.272936f
C4620 a_n6972_8799.n206 gnd 0.266676f
C4621 a_n6972_8799.n207 gnd 0.261553f
C4622 a_n6972_8799.n208 gnd 0.270404f
C4623 a_n6972_8799.n209 gnd 0.272502f
C4624 a_n6972_8799.n210 gnd 0.266036f
C4625 a_n6972_8799.n211 gnd 0.261393f
C4626 a_n6972_8799.n212 gnd 0.899839f
C4627 a_n6972_8799.t130 gnd 0.597459f
C4628 a_n6972_8799.t51 gnd 0.597459f
C4629 a_n6972_8799.t90 gnd 0.597459f
C4630 a_n6972_8799.n213 gnd 0.270005f
C4631 a_n6972_8799.t38 gnd 0.597459f
C4632 a_n6972_8799.t110 gnd 0.597459f
C4633 a_n6972_8799.t62 gnd 0.597459f
C4634 a_n6972_8799.n214 gnd 0.266926f
C4635 a_n6972_8799.t96 gnd 0.597459f
C4636 a_n6972_8799.t43 gnd 0.597459f
C4637 a_n6972_8799.t66 gnd 0.597459f
C4638 a_n6972_8799.n215 gnd 0.270418f
C4639 a_n6972_8799.t126 gnd 0.597459f
C4640 a_n6972_8799.t102 gnd 0.597459f
C4641 a_n6972_8799.t122 gnd 0.597459f
C4642 a_n6972_8799.n216 gnd 0.266356f
C4643 a_n6972_8799.t89 gnd 0.597459f
C4644 a_n6972_8799.t106 gnd 0.597459f
C4645 a_n6972_8799.t56 gnd 0.597459f
C4646 a_n6972_8799.n217 gnd 0.270403f
C4647 a_n6972_8799.t120 gnd 0.608767f
C4648 a_n6972_8799.n218 gnd 0.250481f
C4649 a_n6972_8799.n219 gnd 0.267109f
C4650 a_n6972_8799.n220 gnd 0.261873f
C4651 a_n6972_8799.n221 gnd 0.270286f
C4652 a_n6972_8799.n222 gnd 0.272936f
C4653 a_n6972_8799.n223 gnd 0.266676f
C4654 a_n6972_8799.n224 gnd 0.261553f
C4655 a_n6972_8799.n225 gnd 0.270404f
C4656 a_n6972_8799.n226 gnd 0.272502f
C4657 a_n6972_8799.n227 gnd 0.266036f
C4658 a_n6972_8799.n228 gnd 0.261393f
C4659 a_n6972_8799.n229 gnd 1.08613f
C4660 a_n6972_8799.n230 gnd 12.2028f
C4661 a_n6972_8799.n231 gnd 4.37253f
C4662 a_n6972_8799.n232 gnd 5.6731f
C4663 a_n6972_8799.n233 gnd 1.13458f
C4664 a_n6972_8799.t0 gnd 0.144089f
C4665 commonsourceibias.n0 gnd 0.010545f
C4666 commonsourceibias.t94 gnd 0.159685f
C4667 commonsourceibias.t109 gnd 0.147652f
C4668 commonsourceibias.n1 gnd 0.006423f
C4669 commonsourceibias.n2 gnd 0.007903f
C4670 commonsourceibias.t72 gnd 0.147652f
C4671 commonsourceibias.n3 gnd 0.008017f
C4672 commonsourceibias.n4 gnd 0.007903f
C4673 commonsourceibias.t70 gnd 0.147652f
C4674 commonsourceibias.n5 gnd 0.058913f
C4675 commonsourceibias.t102 gnd 0.147652f
C4676 commonsourceibias.n6 gnd 0.006393f
C4677 commonsourceibias.n7 gnd 0.007903f
C4678 commonsourceibias.t116 gnd 0.147652f
C4679 commonsourceibias.n8 gnd 0.00763f
C4680 commonsourceibias.n9 gnd 0.007903f
C4681 commonsourceibias.t66 gnd 0.147652f
C4682 commonsourceibias.n10 gnd 0.058913f
C4683 commonsourceibias.t92 gnd 0.147652f
C4684 commonsourceibias.n11 gnd 0.006383f
C4685 commonsourceibias.n12 gnd 0.010545f
C4686 commonsourceibias.t48 gnd 0.159685f
C4687 commonsourceibias.t18 gnd 0.147652f
C4688 commonsourceibias.n13 gnd 0.006423f
C4689 commonsourceibias.n14 gnd 0.007903f
C4690 commonsourceibias.t12 gnd 0.147652f
C4691 commonsourceibias.n15 gnd 0.008017f
C4692 commonsourceibias.n16 gnd 0.007903f
C4693 commonsourceibias.t46 gnd 0.147652f
C4694 commonsourceibias.n17 gnd 0.058913f
C4695 commonsourceibias.t24 gnd 0.147652f
C4696 commonsourceibias.n18 gnd 0.006393f
C4697 commonsourceibias.n19 gnd 0.007903f
C4698 commonsourceibias.t52 gnd 0.147652f
C4699 commonsourceibias.n20 gnd 0.00763f
C4700 commonsourceibias.n21 gnd 0.007903f
C4701 commonsourceibias.t60 gnd 0.147652f
C4702 commonsourceibias.n22 gnd 0.058913f
C4703 commonsourceibias.t14 gnd 0.147652f
C4704 commonsourceibias.n23 gnd 0.006383f
C4705 commonsourceibias.n24 gnd 0.007903f
C4706 commonsourceibias.t50 gnd 0.147652f
C4707 commonsourceibias.t42 gnd 0.147652f
C4708 commonsourceibias.n25 gnd 0.058913f
C4709 commonsourceibias.n26 gnd 0.007903f
C4710 commonsourceibias.t56 gnd 0.147652f
C4711 commonsourceibias.n27 gnd 0.058913f
C4712 commonsourceibias.n28 gnd 0.007903f
C4713 commonsourceibias.t62 gnd 0.147652f
C4714 commonsourceibias.n29 gnd 0.058913f
C4715 commonsourceibias.n30 gnd 0.007903f
C4716 commonsourceibias.t10 gnd 0.147652f
C4717 commonsourceibias.n31 gnd 0.008983f
C4718 commonsourceibias.n32 gnd 0.007903f
C4719 commonsourceibias.t28 gnd 0.147652f
C4720 commonsourceibias.n33 gnd 0.010623f
C4721 commonsourceibias.t34 gnd 0.164481f
C4722 commonsourceibias.t20 gnd 0.147652f
C4723 commonsourceibias.n34 gnd 0.065644f
C4724 commonsourceibias.n35 gnd 0.070328f
C4725 commonsourceibias.n36 gnd 0.033639f
C4726 commonsourceibias.n37 gnd 0.007903f
C4727 commonsourceibias.n38 gnd 0.006423f
C4728 commonsourceibias.n39 gnd 0.01089f
C4729 commonsourceibias.n40 gnd 0.058913f
C4730 commonsourceibias.n41 gnd 0.010937f
C4731 commonsourceibias.n42 gnd 0.007903f
C4732 commonsourceibias.n43 gnd 0.007903f
C4733 commonsourceibias.n44 gnd 0.007903f
C4734 commonsourceibias.n45 gnd 0.008017f
C4735 commonsourceibias.n46 gnd 0.058913f
C4736 commonsourceibias.n47 gnd 0.009741f
C4737 commonsourceibias.n48 gnd 0.010776f
C4738 commonsourceibias.n49 gnd 0.007903f
C4739 commonsourceibias.n50 gnd 0.007903f
C4740 commonsourceibias.n51 gnd 0.010705f
C4741 commonsourceibias.n52 gnd 0.006393f
C4742 commonsourceibias.n53 gnd 0.010838f
C4743 commonsourceibias.n54 gnd 0.007903f
C4744 commonsourceibias.n55 gnd 0.007903f
C4745 commonsourceibias.n56 gnd 0.010904f
C4746 commonsourceibias.n57 gnd 0.009403f
C4747 commonsourceibias.n58 gnd 0.00763f
C4748 commonsourceibias.n59 gnd 0.007903f
C4749 commonsourceibias.n60 gnd 0.007903f
C4750 commonsourceibias.n61 gnd 0.009667f
C4751 commonsourceibias.n62 gnd 0.01085f
C4752 commonsourceibias.n63 gnd 0.058913f
C4753 commonsourceibias.n64 gnd 0.010777f
C4754 commonsourceibias.n65 gnd 0.007903f
C4755 commonsourceibias.n66 gnd 0.007903f
C4756 commonsourceibias.n67 gnd 0.007903f
C4757 commonsourceibias.n68 gnd 0.010777f
C4758 commonsourceibias.n69 gnd 0.058913f
C4759 commonsourceibias.n70 gnd 0.01085f
C4760 commonsourceibias.n71 gnd 0.009667f
C4761 commonsourceibias.n72 gnd 0.007903f
C4762 commonsourceibias.n73 gnd 0.007903f
C4763 commonsourceibias.n74 gnd 0.007903f
C4764 commonsourceibias.n75 gnd 0.009403f
C4765 commonsourceibias.n76 gnd 0.010904f
C4766 commonsourceibias.n77 gnd 0.058913f
C4767 commonsourceibias.n78 gnd 0.010838f
C4768 commonsourceibias.n79 gnd 0.007903f
C4769 commonsourceibias.n80 gnd 0.007903f
C4770 commonsourceibias.n81 gnd 0.007903f
C4771 commonsourceibias.n82 gnd 0.010705f
C4772 commonsourceibias.n83 gnd 0.058913f
C4773 commonsourceibias.n84 gnd 0.010776f
C4774 commonsourceibias.n85 gnd 0.009741f
C4775 commonsourceibias.n86 gnd 0.007903f
C4776 commonsourceibias.n87 gnd 0.007903f
C4777 commonsourceibias.n88 gnd 0.007903f
C4778 commonsourceibias.n89 gnd 0.008983f
C4779 commonsourceibias.n90 gnd 0.010937f
C4780 commonsourceibias.n91 gnd 0.058913f
C4781 commonsourceibias.n92 gnd 0.01089f
C4782 commonsourceibias.n93 gnd 0.007903f
C4783 commonsourceibias.n94 gnd 0.007903f
C4784 commonsourceibias.n95 gnd 0.007903f
C4785 commonsourceibias.n96 gnd 0.010623f
C4786 commonsourceibias.n97 gnd 0.058913f
C4787 commonsourceibias.n98 gnd 0.010649f
C4788 commonsourceibias.n99 gnd 0.071041f
C4789 commonsourceibias.n100 gnd 0.079434f
C4790 commonsourceibias.t49 gnd 0.017054f
C4791 commonsourceibias.t19 gnd 0.017054f
C4792 commonsourceibias.n101 gnd 0.150693f
C4793 commonsourceibias.n102 gnd 0.130533f
C4794 commonsourceibias.t13 gnd 0.017054f
C4795 commonsourceibias.t47 gnd 0.017054f
C4796 commonsourceibias.n103 gnd 0.150693f
C4797 commonsourceibias.n104 gnd 0.069219f
C4798 commonsourceibias.t25 gnd 0.017054f
C4799 commonsourceibias.t53 gnd 0.017054f
C4800 commonsourceibias.n105 gnd 0.150693f
C4801 commonsourceibias.n106 gnd 0.069219f
C4802 commonsourceibias.t61 gnd 0.017054f
C4803 commonsourceibias.t15 gnd 0.017054f
C4804 commonsourceibias.n107 gnd 0.150693f
C4805 commonsourceibias.n108 gnd 0.057829f
C4806 commonsourceibias.t21 gnd 0.017054f
C4807 commonsourceibias.t35 gnd 0.017054f
C4808 commonsourceibias.n109 gnd 0.151197f
C4809 commonsourceibias.t11 gnd 0.017054f
C4810 commonsourceibias.t29 gnd 0.017054f
C4811 commonsourceibias.n110 gnd 0.150693f
C4812 commonsourceibias.n111 gnd 0.140418f
C4813 commonsourceibias.t57 gnd 0.017054f
C4814 commonsourceibias.t63 gnd 0.017054f
C4815 commonsourceibias.n112 gnd 0.150693f
C4816 commonsourceibias.n113 gnd 0.069219f
C4817 commonsourceibias.t51 gnd 0.017054f
C4818 commonsourceibias.t43 gnd 0.017054f
C4819 commonsourceibias.n114 gnd 0.150693f
C4820 commonsourceibias.n115 gnd 0.057829f
C4821 commonsourceibias.n116 gnd 0.070025f
C4822 commonsourceibias.n117 gnd 0.007903f
C4823 commonsourceibias.t89 gnd 0.147652f
C4824 commonsourceibias.t105 gnd 0.147652f
C4825 commonsourceibias.n118 gnd 0.058913f
C4826 commonsourceibias.n119 gnd 0.007903f
C4827 commonsourceibias.t85 gnd 0.147652f
C4828 commonsourceibias.n120 gnd 0.058913f
C4829 commonsourceibias.n121 gnd 0.007903f
C4830 commonsourceibias.t82 gnd 0.147652f
C4831 commonsourceibias.n122 gnd 0.058913f
C4832 commonsourceibias.n123 gnd 0.007903f
C4833 commonsourceibias.t97 gnd 0.147652f
C4834 commonsourceibias.n124 gnd 0.008983f
C4835 commonsourceibias.n125 gnd 0.007903f
C4836 commonsourceibias.t111 gnd 0.147652f
C4837 commonsourceibias.n126 gnd 0.010623f
C4838 commonsourceibias.t88 gnd 0.164481f
C4839 commonsourceibias.t75 gnd 0.147652f
C4840 commonsourceibias.n127 gnd 0.065644f
C4841 commonsourceibias.n128 gnd 0.070328f
C4842 commonsourceibias.n129 gnd 0.033639f
C4843 commonsourceibias.n130 gnd 0.007903f
C4844 commonsourceibias.n131 gnd 0.006423f
C4845 commonsourceibias.n132 gnd 0.01089f
C4846 commonsourceibias.n133 gnd 0.058913f
C4847 commonsourceibias.n134 gnd 0.010937f
C4848 commonsourceibias.n135 gnd 0.007903f
C4849 commonsourceibias.n136 gnd 0.007903f
C4850 commonsourceibias.n137 gnd 0.007903f
C4851 commonsourceibias.n138 gnd 0.008017f
C4852 commonsourceibias.n139 gnd 0.058913f
C4853 commonsourceibias.n140 gnd 0.009741f
C4854 commonsourceibias.n141 gnd 0.010776f
C4855 commonsourceibias.n142 gnd 0.007903f
C4856 commonsourceibias.n143 gnd 0.007903f
C4857 commonsourceibias.n144 gnd 0.010705f
C4858 commonsourceibias.n145 gnd 0.006393f
C4859 commonsourceibias.n146 gnd 0.010838f
C4860 commonsourceibias.n147 gnd 0.007903f
C4861 commonsourceibias.n148 gnd 0.007903f
C4862 commonsourceibias.n149 gnd 0.010904f
C4863 commonsourceibias.n150 gnd 0.009403f
C4864 commonsourceibias.n151 gnd 0.00763f
C4865 commonsourceibias.n152 gnd 0.007903f
C4866 commonsourceibias.n153 gnd 0.007903f
C4867 commonsourceibias.n154 gnd 0.009667f
C4868 commonsourceibias.n155 gnd 0.01085f
C4869 commonsourceibias.n156 gnd 0.058913f
C4870 commonsourceibias.n157 gnd 0.010777f
C4871 commonsourceibias.n158 gnd 0.007865f
C4872 commonsourceibias.n159 gnd 0.057129f
C4873 commonsourceibias.n160 gnd 0.007865f
C4874 commonsourceibias.n161 gnd 0.010777f
C4875 commonsourceibias.n162 gnd 0.058913f
C4876 commonsourceibias.n163 gnd 0.01085f
C4877 commonsourceibias.n164 gnd 0.009667f
C4878 commonsourceibias.n165 gnd 0.007903f
C4879 commonsourceibias.n166 gnd 0.007903f
C4880 commonsourceibias.n167 gnd 0.007903f
C4881 commonsourceibias.n168 gnd 0.009403f
C4882 commonsourceibias.n169 gnd 0.010904f
C4883 commonsourceibias.n170 gnd 0.058913f
C4884 commonsourceibias.n171 gnd 0.010838f
C4885 commonsourceibias.n172 gnd 0.007903f
C4886 commonsourceibias.n173 gnd 0.007903f
C4887 commonsourceibias.n174 gnd 0.007903f
C4888 commonsourceibias.n175 gnd 0.010705f
C4889 commonsourceibias.n176 gnd 0.058913f
C4890 commonsourceibias.n177 gnd 0.010776f
C4891 commonsourceibias.n178 gnd 0.009741f
C4892 commonsourceibias.n179 gnd 0.007903f
C4893 commonsourceibias.n180 gnd 0.007903f
C4894 commonsourceibias.n181 gnd 0.007903f
C4895 commonsourceibias.n182 gnd 0.008983f
C4896 commonsourceibias.n183 gnd 0.010937f
C4897 commonsourceibias.n184 gnd 0.058913f
C4898 commonsourceibias.n185 gnd 0.01089f
C4899 commonsourceibias.n186 gnd 0.007903f
C4900 commonsourceibias.n187 gnd 0.007903f
C4901 commonsourceibias.n188 gnd 0.007903f
C4902 commonsourceibias.n189 gnd 0.010623f
C4903 commonsourceibias.n190 gnd 0.058913f
C4904 commonsourceibias.n191 gnd 0.010649f
C4905 commonsourceibias.n192 gnd 0.071041f
C4906 commonsourceibias.n193 gnd 0.046914f
C4907 commonsourceibias.n194 gnd 0.010545f
C4908 commonsourceibias.t96 gnd 0.147652f
C4909 commonsourceibias.n195 gnd 0.006423f
C4910 commonsourceibias.n196 gnd 0.007903f
C4911 commonsourceibias.t65 gnd 0.147652f
C4912 commonsourceibias.n197 gnd 0.008017f
C4913 commonsourceibias.n198 gnd 0.007903f
C4914 commonsourceibias.t127 gnd 0.147652f
C4915 commonsourceibias.n199 gnd 0.058913f
C4916 commonsourceibias.t87 gnd 0.147652f
C4917 commonsourceibias.n200 gnd 0.006393f
C4918 commonsourceibias.n201 gnd 0.007903f
C4919 commonsourceibias.t104 gnd 0.147652f
C4920 commonsourceibias.n202 gnd 0.00763f
C4921 commonsourceibias.n203 gnd 0.007903f
C4922 commonsourceibias.t122 gnd 0.147652f
C4923 commonsourceibias.n204 gnd 0.058913f
C4924 commonsourceibias.t80 gnd 0.147652f
C4925 commonsourceibias.n205 gnd 0.006383f
C4926 commonsourceibias.n206 gnd 0.007903f
C4927 commonsourceibias.t76 gnd 0.147652f
C4928 commonsourceibias.t90 gnd 0.147652f
C4929 commonsourceibias.n207 gnd 0.058913f
C4930 commonsourceibias.n208 gnd 0.007903f
C4931 commonsourceibias.t74 gnd 0.147652f
C4932 commonsourceibias.n209 gnd 0.058913f
C4933 commonsourceibias.n210 gnd 0.007903f
C4934 commonsourceibias.t71 gnd 0.147652f
C4935 commonsourceibias.n211 gnd 0.058913f
C4936 commonsourceibias.n212 gnd 0.007903f
C4937 commonsourceibias.t83 gnd 0.147652f
C4938 commonsourceibias.n213 gnd 0.008983f
C4939 commonsourceibias.n214 gnd 0.007903f
C4940 commonsourceibias.t98 gnd 0.147652f
C4941 commonsourceibias.n215 gnd 0.010623f
C4942 commonsourceibias.t77 gnd 0.164481f
C4943 commonsourceibias.t67 gnd 0.147652f
C4944 commonsourceibias.n216 gnd 0.065644f
C4945 commonsourceibias.n217 gnd 0.070328f
C4946 commonsourceibias.n218 gnd 0.033639f
C4947 commonsourceibias.n219 gnd 0.007903f
C4948 commonsourceibias.n220 gnd 0.006423f
C4949 commonsourceibias.n221 gnd 0.01089f
C4950 commonsourceibias.n222 gnd 0.058913f
C4951 commonsourceibias.n223 gnd 0.010937f
C4952 commonsourceibias.n224 gnd 0.007903f
C4953 commonsourceibias.n225 gnd 0.007903f
C4954 commonsourceibias.n226 gnd 0.007903f
C4955 commonsourceibias.n227 gnd 0.008017f
C4956 commonsourceibias.n228 gnd 0.058913f
C4957 commonsourceibias.n229 gnd 0.009741f
C4958 commonsourceibias.n230 gnd 0.010776f
C4959 commonsourceibias.n231 gnd 0.007903f
C4960 commonsourceibias.n232 gnd 0.007903f
C4961 commonsourceibias.n233 gnd 0.010705f
C4962 commonsourceibias.n234 gnd 0.006393f
C4963 commonsourceibias.n235 gnd 0.010838f
C4964 commonsourceibias.n236 gnd 0.007903f
C4965 commonsourceibias.n237 gnd 0.007903f
C4966 commonsourceibias.n238 gnd 0.010904f
C4967 commonsourceibias.n239 gnd 0.009403f
C4968 commonsourceibias.n240 gnd 0.00763f
C4969 commonsourceibias.n241 gnd 0.007903f
C4970 commonsourceibias.n242 gnd 0.007903f
C4971 commonsourceibias.n243 gnd 0.009667f
C4972 commonsourceibias.n244 gnd 0.01085f
C4973 commonsourceibias.n245 gnd 0.058913f
C4974 commonsourceibias.n246 gnd 0.010777f
C4975 commonsourceibias.n247 gnd 0.007903f
C4976 commonsourceibias.n248 gnd 0.007903f
C4977 commonsourceibias.n249 gnd 0.007903f
C4978 commonsourceibias.n250 gnd 0.010777f
C4979 commonsourceibias.n251 gnd 0.058913f
C4980 commonsourceibias.n252 gnd 0.01085f
C4981 commonsourceibias.n253 gnd 0.009667f
C4982 commonsourceibias.n254 gnd 0.007903f
C4983 commonsourceibias.n255 gnd 0.007903f
C4984 commonsourceibias.n256 gnd 0.007903f
C4985 commonsourceibias.n257 gnd 0.009403f
C4986 commonsourceibias.n258 gnd 0.010904f
C4987 commonsourceibias.n259 gnd 0.058913f
C4988 commonsourceibias.n260 gnd 0.010838f
C4989 commonsourceibias.n261 gnd 0.007903f
C4990 commonsourceibias.n262 gnd 0.007903f
C4991 commonsourceibias.n263 gnd 0.007903f
C4992 commonsourceibias.n264 gnd 0.010705f
C4993 commonsourceibias.n265 gnd 0.058913f
C4994 commonsourceibias.n266 gnd 0.010776f
C4995 commonsourceibias.n267 gnd 0.009741f
C4996 commonsourceibias.n268 gnd 0.007903f
C4997 commonsourceibias.n269 gnd 0.007903f
C4998 commonsourceibias.n270 gnd 0.007903f
C4999 commonsourceibias.n271 gnd 0.008983f
C5000 commonsourceibias.n272 gnd 0.010937f
C5001 commonsourceibias.n273 gnd 0.058913f
C5002 commonsourceibias.n274 gnd 0.01089f
C5003 commonsourceibias.n275 gnd 0.007903f
C5004 commonsourceibias.n276 gnd 0.007903f
C5005 commonsourceibias.n277 gnd 0.007903f
C5006 commonsourceibias.n278 gnd 0.010623f
C5007 commonsourceibias.n279 gnd 0.058913f
C5008 commonsourceibias.n280 gnd 0.010649f
C5009 commonsourceibias.t81 gnd 0.159685f
C5010 commonsourceibias.n281 gnd 0.071041f
C5011 commonsourceibias.n282 gnd 0.02535f
C5012 commonsourceibias.n283 gnd 0.398385f
C5013 commonsourceibias.n284 gnd 0.010545f
C5014 commonsourceibias.t113 gnd 0.159685f
C5015 commonsourceibias.t123 gnd 0.147652f
C5016 commonsourceibias.n285 gnd 0.006423f
C5017 commonsourceibias.n286 gnd 0.007903f
C5018 commonsourceibias.t68 gnd 0.147652f
C5019 commonsourceibias.n287 gnd 0.008017f
C5020 commonsourceibias.n288 gnd 0.007903f
C5021 commonsourceibias.t119 gnd 0.147652f
C5022 commonsourceibias.n289 gnd 0.006393f
C5023 commonsourceibias.n290 gnd 0.007903f
C5024 commonsourceibias.t64 gnd 0.147652f
C5025 commonsourceibias.n291 gnd 0.00763f
C5026 commonsourceibias.n292 gnd 0.007903f
C5027 commonsourceibias.t112 gnd 0.147652f
C5028 commonsourceibias.n293 gnd 0.006383f
C5029 commonsourceibias.n294 gnd 0.007903f
C5030 commonsourceibias.t107 gnd 0.147652f
C5031 commonsourceibias.t121 gnd 0.147652f
C5032 commonsourceibias.n295 gnd 0.058913f
C5033 commonsourceibias.n296 gnd 0.007903f
C5034 commonsourceibias.t78 gnd 0.147652f
C5035 commonsourceibias.n297 gnd 0.058913f
C5036 commonsourceibias.n298 gnd 0.007903f
C5037 commonsourceibias.t101 gnd 0.147652f
C5038 commonsourceibias.n299 gnd 0.058913f
C5039 commonsourceibias.n300 gnd 0.007903f
C5040 commonsourceibias.t115 gnd 0.147652f
C5041 commonsourceibias.n301 gnd 0.008983f
C5042 commonsourceibias.n302 gnd 0.007903f
C5043 commonsourceibias.t125 gnd 0.147652f
C5044 commonsourceibias.n303 gnd 0.010623f
C5045 commonsourceibias.t108 gnd 0.164481f
C5046 commonsourceibias.t91 gnd 0.147652f
C5047 commonsourceibias.n304 gnd 0.065644f
C5048 commonsourceibias.n305 gnd 0.070328f
C5049 commonsourceibias.n306 gnd 0.033639f
C5050 commonsourceibias.n307 gnd 0.007903f
C5051 commonsourceibias.n308 gnd 0.006423f
C5052 commonsourceibias.n309 gnd 0.01089f
C5053 commonsourceibias.n310 gnd 0.058913f
C5054 commonsourceibias.n311 gnd 0.010937f
C5055 commonsourceibias.n312 gnd 0.007903f
C5056 commonsourceibias.n313 gnd 0.007903f
C5057 commonsourceibias.n314 gnd 0.007903f
C5058 commonsourceibias.n315 gnd 0.008017f
C5059 commonsourceibias.n316 gnd 0.058913f
C5060 commonsourceibias.n317 gnd 0.009741f
C5061 commonsourceibias.n318 gnd 0.010776f
C5062 commonsourceibias.n319 gnd 0.007903f
C5063 commonsourceibias.n320 gnd 0.007903f
C5064 commonsourceibias.n321 gnd 0.010705f
C5065 commonsourceibias.n322 gnd 0.006393f
C5066 commonsourceibias.n323 gnd 0.010838f
C5067 commonsourceibias.n324 gnd 0.007903f
C5068 commonsourceibias.n325 gnd 0.007903f
C5069 commonsourceibias.n326 gnd 0.010904f
C5070 commonsourceibias.n327 gnd 0.009403f
C5071 commonsourceibias.n328 gnd 0.00763f
C5072 commonsourceibias.n329 gnd 0.007903f
C5073 commonsourceibias.n330 gnd 0.007903f
C5074 commonsourceibias.n331 gnd 0.009667f
C5075 commonsourceibias.n332 gnd 0.01085f
C5076 commonsourceibias.n333 gnd 0.058913f
C5077 commonsourceibias.n334 gnd 0.010777f
C5078 commonsourceibias.n335 gnd 0.007865f
C5079 commonsourceibias.t31 gnd 0.017054f
C5080 commonsourceibias.t33 gnd 0.017054f
C5081 commonsourceibias.n336 gnd 0.151197f
C5082 commonsourceibias.t39 gnd 0.017054f
C5083 commonsourceibias.t37 gnd 0.017054f
C5084 commonsourceibias.n337 gnd 0.150693f
C5085 commonsourceibias.n338 gnd 0.140418f
C5086 commonsourceibias.t9 gnd 0.017054f
C5087 commonsourceibias.t41 gnd 0.017054f
C5088 commonsourceibias.n339 gnd 0.150693f
C5089 commonsourceibias.n340 gnd 0.069219f
C5090 commonsourceibias.t23 gnd 0.017054f
C5091 commonsourceibias.t5 gnd 0.017054f
C5092 commonsourceibias.n341 gnd 0.150693f
C5093 commonsourceibias.n342 gnd 0.057829f
C5094 commonsourceibias.n343 gnd 0.010545f
C5095 commonsourceibias.t26 gnd 0.147652f
C5096 commonsourceibias.n344 gnd 0.006423f
C5097 commonsourceibias.n345 gnd 0.007903f
C5098 commonsourceibias.t54 gnd 0.147652f
C5099 commonsourceibias.n346 gnd 0.008017f
C5100 commonsourceibias.n347 gnd 0.007903f
C5101 commonsourceibias.t16 gnd 0.147652f
C5102 commonsourceibias.n348 gnd 0.006393f
C5103 commonsourceibias.n349 gnd 0.007903f
C5104 commonsourceibias.t6 gnd 0.147652f
C5105 commonsourceibias.n350 gnd 0.00763f
C5106 commonsourceibias.n351 gnd 0.007903f
C5107 commonsourceibias.t58 gnd 0.147652f
C5108 commonsourceibias.n352 gnd 0.006383f
C5109 commonsourceibias.n353 gnd 0.007903f
C5110 commonsourceibias.t4 gnd 0.147652f
C5111 commonsourceibias.t22 gnd 0.147652f
C5112 commonsourceibias.n354 gnd 0.058913f
C5113 commonsourceibias.n355 gnd 0.007903f
C5114 commonsourceibias.t40 gnd 0.147652f
C5115 commonsourceibias.n356 gnd 0.058913f
C5116 commonsourceibias.n357 gnd 0.007903f
C5117 commonsourceibias.t8 gnd 0.147652f
C5118 commonsourceibias.n358 gnd 0.058913f
C5119 commonsourceibias.n359 gnd 0.007903f
C5120 commonsourceibias.t36 gnd 0.147652f
C5121 commonsourceibias.n360 gnd 0.008983f
C5122 commonsourceibias.n361 gnd 0.007903f
C5123 commonsourceibias.t38 gnd 0.147652f
C5124 commonsourceibias.n362 gnd 0.010623f
C5125 commonsourceibias.t30 gnd 0.164481f
C5126 commonsourceibias.t32 gnd 0.147652f
C5127 commonsourceibias.n363 gnd 0.065644f
C5128 commonsourceibias.n364 gnd 0.070328f
C5129 commonsourceibias.n365 gnd 0.033639f
C5130 commonsourceibias.n366 gnd 0.007903f
C5131 commonsourceibias.n367 gnd 0.006423f
C5132 commonsourceibias.n368 gnd 0.01089f
C5133 commonsourceibias.n369 gnd 0.058913f
C5134 commonsourceibias.n370 gnd 0.010937f
C5135 commonsourceibias.n371 gnd 0.007903f
C5136 commonsourceibias.n372 gnd 0.007903f
C5137 commonsourceibias.n373 gnd 0.007903f
C5138 commonsourceibias.n374 gnd 0.008017f
C5139 commonsourceibias.n375 gnd 0.058913f
C5140 commonsourceibias.n376 gnd 0.009741f
C5141 commonsourceibias.n377 gnd 0.010776f
C5142 commonsourceibias.n378 gnd 0.007903f
C5143 commonsourceibias.n379 gnd 0.007903f
C5144 commonsourceibias.n380 gnd 0.010705f
C5145 commonsourceibias.n381 gnd 0.006393f
C5146 commonsourceibias.n382 gnd 0.010838f
C5147 commonsourceibias.n383 gnd 0.007903f
C5148 commonsourceibias.n384 gnd 0.007903f
C5149 commonsourceibias.n385 gnd 0.010904f
C5150 commonsourceibias.n386 gnd 0.009403f
C5151 commonsourceibias.n387 gnd 0.00763f
C5152 commonsourceibias.n388 gnd 0.007903f
C5153 commonsourceibias.n389 gnd 0.007903f
C5154 commonsourceibias.n390 gnd 0.009667f
C5155 commonsourceibias.n391 gnd 0.01085f
C5156 commonsourceibias.n392 gnd 0.058913f
C5157 commonsourceibias.n393 gnd 0.010777f
C5158 commonsourceibias.n394 gnd 0.007903f
C5159 commonsourceibias.n395 gnd 0.007903f
C5160 commonsourceibias.n396 gnd 0.007903f
C5161 commonsourceibias.n397 gnd 0.010777f
C5162 commonsourceibias.n398 gnd 0.058913f
C5163 commonsourceibias.n399 gnd 0.01085f
C5164 commonsourceibias.t44 gnd 0.147652f
C5165 commonsourceibias.n400 gnd 0.058913f
C5166 commonsourceibias.n401 gnd 0.009667f
C5167 commonsourceibias.n402 gnd 0.007903f
C5168 commonsourceibias.n403 gnd 0.007903f
C5169 commonsourceibias.n404 gnd 0.007903f
C5170 commonsourceibias.n405 gnd 0.009403f
C5171 commonsourceibias.n406 gnd 0.010904f
C5172 commonsourceibias.n407 gnd 0.058913f
C5173 commonsourceibias.n408 gnd 0.010838f
C5174 commonsourceibias.n409 gnd 0.007903f
C5175 commonsourceibias.n410 gnd 0.007903f
C5176 commonsourceibias.n411 gnd 0.007903f
C5177 commonsourceibias.n412 gnd 0.010705f
C5178 commonsourceibias.n413 gnd 0.058913f
C5179 commonsourceibias.n414 gnd 0.010776f
C5180 commonsourceibias.t0 gnd 0.147652f
C5181 commonsourceibias.n415 gnd 0.058913f
C5182 commonsourceibias.n416 gnd 0.009741f
C5183 commonsourceibias.n417 gnd 0.007903f
C5184 commonsourceibias.n418 gnd 0.007903f
C5185 commonsourceibias.n419 gnd 0.007903f
C5186 commonsourceibias.n420 gnd 0.008983f
C5187 commonsourceibias.n421 gnd 0.010937f
C5188 commonsourceibias.n422 gnd 0.058913f
C5189 commonsourceibias.n423 gnd 0.01089f
C5190 commonsourceibias.n424 gnd 0.007903f
C5191 commonsourceibias.n425 gnd 0.007903f
C5192 commonsourceibias.n426 gnd 0.007903f
C5193 commonsourceibias.n427 gnd 0.010623f
C5194 commonsourceibias.n428 gnd 0.058913f
C5195 commonsourceibias.n429 gnd 0.010649f
C5196 commonsourceibias.t2 gnd 0.159685f
C5197 commonsourceibias.n430 gnd 0.071041f
C5198 commonsourceibias.n431 gnd 0.079434f
C5199 commonsourceibias.t27 gnd 0.017054f
C5200 commonsourceibias.t3 gnd 0.017054f
C5201 commonsourceibias.n432 gnd 0.150693f
C5202 commonsourceibias.n433 gnd 0.130533f
C5203 commonsourceibias.t1 gnd 0.017054f
C5204 commonsourceibias.t55 gnd 0.017054f
C5205 commonsourceibias.n434 gnd 0.150693f
C5206 commonsourceibias.n435 gnd 0.069219f
C5207 commonsourceibias.t7 gnd 0.017054f
C5208 commonsourceibias.t17 gnd 0.017054f
C5209 commonsourceibias.n436 gnd 0.150693f
C5210 commonsourceibias.n437 gnd 0.069219f
C5211 commonsourceibias.t59 gnd 0.017054f
C5212 commonsourceibias.t45 gnd 0.017054f
C5213 commonsourceibias.n438 gnd 0.150693f
C5214 commonsourceibias.n439 gnd 0.057829f
C5215 commonsourceibias.n440 gnd 0.070025f
C5216 commonsourceibias.n441 gnd 0.057129f
C5217 commonsourceibias.n442 gnd 0.007865f
C5218 commonsourceibias.n443 gnd 0.010777f
C5219 commonsourceibias.n444 gnd 0.058913f
C5220 commonsourceibias.n445 gnd 0.01085f
C5221 commonsourceibias.t126 gnd 0.147652f
C5222 commonsourceibias.n446 gnd 0.058913f
C5223 commonsourceibias.n447 gnd 0.009667f
C5224 commonsourceibias.n448 gnd 0.007903f
C5225 commonsourceibias.n449 gnd 0.007903f
C5226 commonsourceibias.n450 gnd 0.007903f
C5227 commonsourceibias.n451 gnd 0.009403f
C5228 commonsourceibias.n452 gnd 0.010904f
C5229 commonsourceibias.n453 gnd 0.058913f
C5230 commonsourceibias.n454 gnd 0.010838f
C5231 commonsourceibias.n455 gnd 0.007903f
C5232 commonsourceibias.n456 gnd 0.007903f
C5233 commonsourceibias.n457 gnd 0.007903f
C5234 commonsourceibias.n458 gnd 0.010705f
C5235 commonsourceibias.n459 gnd 0.058913f
C5236 commonsourceibias.n460 gnd 0.010776f
C5237 commonsourceibias.t84 gnd 0.147652f
C5238 commonsourceibias.n461 gnd 0.058913f
C5239 commonsourceibias.n462 gnd 0.009741f
C5240 commonsourceibias.n463 gnd 0.007903f
C5241 commonsourceibias.n464 gnd 0.007903f
C5242 commonsourceibias.n465 gnd 0.007903f
C5243 commonsourceibias.n466 gnd 0.008983f
C5244 commonsourceibias.n467 gnd 0.010937f
C5245 commonsourceibias.n468 gnd 0.058913f
C5246 commonsourceibias.n469 gnd 0.01089f
C5247 commonsourceibias.n470 gnd 0.007903f
C5248 commonsourceibias.n471 gnd 0.007903f
C5249 commonsourceibias.n472 gnd 0.007903f
C5250 commonsourceibias.n473 gnd 0.010623f
C5251 commonsourceibias.n474 gnd 0.058913f
C5252 commonsourceibias.n475 gnd 0.010649f
C5253 commonsourceibias.n476 gnd 0.071041f
C5254 commonsourceibias.n477 gnd 0.046914f
C5255 commonsourceibias.n478 gnd 0.010545f
C5256 commonsourceibias.t114 gnd 0.147652f
C5257 commonsourceibias.n479 gnd 0.006423f
C5258 commonsourceibias.n480 gnd 0.007903f
C5259 commonsourceibias.t124 gnd 0.147652f
C5260 commonsourceibias.n481 gnd 0.008017f
C5261 commonsourceibias.n482 gnd 0.007903f
C5262 commonsourceibias.t106 gnd 0.147652f
C5263 commonsourceibias.n483 gnd 0.006393f
C5264 commonsourceibias.n484 gnd 0.007903f
C5265 commonsourceibias.t120 gnd 0.147652f
C5266 commonsourceibias.n485 gnd 0.00763f
C5267 commonsourceibias.n486 gnd 0.007903f
C5268 commonsourceibias.t100 gnd 0.147652f
C5269 commonsourceibias.n487 gnd 0.006383f
C5270 commonsourceibias.n488 gnd 0.007903f
C5271 commonsourceibias.t93 gnd 0.147652f
C5272 commonsourceibias.t110 gnd 0.147652f
C5273 commonsourceibias.n489 gnd 0.058913f
C5274 commonsourceibias.n490 gnd 0.007903f
C5275 commonsourceibias.t69 gnd 0.147652f
C5276 commonsourceibias.n491 gnd 0.058913f
C5277 commonsourceibias.n492 gnd 0.007903f
C5278 commonsourceibias.t86 gnd 0.147652f
C5279 commonsourceibias.n493 gnd 0.058913f
C5280 commonsourceibias.n494 gnd 0.007903f
C5281 commonsourceibias.t103 gnd 0.147652f
C5282 commonsourceibias.n495 gnd 0.008983f
C5283 commonsourceibias.n496 gnd 0.007903f
C5284 commonsourceibias.t118 gnd 0.147652f
C5285 commonsourceibias.n497 gnd 0.010623f
C5286 commonsourceibias.t95 gnd 0.164481f
C5287 commonsourceibias.t79 gnd 0.147652f
C5288 commonsourceibias.n498 gnd 0.065644f
C5289 commonsourceibias.n499 gnd 0.070328f
C5290 commonsourceibias.n500 gnd 0.033639f
C5291 commonsourceibias.n501 gnd 0.007903f
C5292 commonsourceibias.n502 gnd 0.006423f
C5293 commonsourceibias.n503 gnd 0.01089f
C5294 commonsourceibias.n504 gnd 0.058913f
C5295 commonsourceibias.n505 gnd 0.010937f
C5296 commonsourceibias.n506 gnd 0.007903f
C5297 commonsourceibias.n507 gnd 0.007903f
C5298 commonsourceibias.n508 gnd 0.007903f
C5299 commonsourceibias.n509 gnd 0.008017f
C5300 commonsourceibias.n510 gnd 0.058913f
C5301 commonsourceibias.n511 gnd 0.009741f
C5302 commonsourceibias.n512 gnd 0.010776f
C5303 commonsourceibias.n513 gnd 0.007903f
C5304 commonsourceibias.n514 gnd 0.007903f
C5305 commonsourceibias.n515 gnd 0.010705f
C5306 commonsourceibias.n516 gnd 0.006393f
C5307 commonsourceibias.n517 gnd 0.010838f
C5308 commonsourceibias.n518 gnd 0.007903f
C5309 commonsourceibias.n519 gnd 0.007903f
C5310 commonsourceibias.n520 gnd 0.010904f
C5311 commonsourceibias.n521 gnd 0.009403f
C5312 commonsourceibias.n522 gnd 0.00763f
C5313 commonsourceibias.n523 gnd 0.007903f
C5314 commonsourceibias.n524 gnd 0.007903f
C5315 commonsourceibias.n525 gnd 0.009667f
C5316 commonsourceibias.n526 gnd 0.01085f
C5317 commonsourceibias.n527 gnd 0.058913f
C5318 commonsourceibias.n528 gnd 0.010777f
C5319 commonsourceibias.n529 gnd 0.007903f
C5320 commonsourceibias.n530 gnd 0.007903f
C5321 commonsourceibias.n531 gnd 0.007903f
C5322 commonsourceibias.n532 gnd 0.010777f
C5323 commonsourceibias.n533 gnd 0.058913f
C5324 commonsourceibias.n534 gnd 0.01085f
C5325 commonsourceibias.t117 gnd 0.147652f
C5326 commonsourceibias.n535 gnd 0.058913f
C5327 commonsourceibias.n536 gnd 0.009667f
C5328 commonsourceibias.n537 gnd 0.007903f
C5329 commonsourceibias.n538 gnd 0.007903f
C5330 commonsourceibias.n539 gnd 0.007903f
C5331 commonsourceibias.n540 gnd 0.009403f
C5332 commonsourceibias.n541 gnd 0.010904f
C5333 commonsourceibias.n542 gnd 0.058913f
C5334 commonsourceibias.n543 gnd 0.010838f
C5335 commonsourceibias.n544 gnd 0.007903f
C5336 commonsourceibias.n545 gnd 0.007903f
C5337 commonsourceibias.n546 gnd 0.007903f
C5338 commonsourceibias.n547 gnd 0.010705f
C5339 commonsourceibias.n548 gnd 0.058913f
C5340 commonsourceibias.n549 gnd 0.010776f
C5341 commonsourceibias.t73 gnd 0.147652f
C5342 commonsourceibias.n550 gnd 0.058913f
C5343 commonsourceibias.n551 gnd 0.009741f
C5344 commonsourceibias.n552 gnd 0.007903f
C5345 commonsourceibias.n553 gnd 0.007903f
C5346 commonsourceibias.n554 gnd 0.007903f
C5347 commonsourceibias.n555 gnd 0.008983f
C5348 commonsourceibias.n556 gnd 0.010937f
C5349 commonsourceibias.n557 gnd 0.058913f
C5350 commonsourceibias.n558 gnd 0.01089f
C5351 commonsourceibias.n559 gnd 0.007903f
C5352 commonsourceibias.n560 gnd 0.007903f
C5353 commonsourceibias.n561 gnd 0.007903f
C5354 commonsourceibias.n562 gnd 0.010623f
C5355 commonsourceibias.n563 gnd 0.058913f
C5356 commonsourceibias.n564 gnd 0.010649f
C5357 commonsourceibias.t99 gnd 0.159685f
C5358 commonsourceibias.n565 gnd 0.071041f
C5359 commonsourceibias.n566 gnd 0.02535f
C5360 commonsourceibias.n567 gnd 0.218509f
C5361 commonsourceibias.n568 gnd 4.2686f
C5362 a_n1986_8322.n0 gnd 1.11016f
C5363 a_n1986_8322.n1 gnd 1.11016f
C5364 a_n1986_8322.n2 gnd 1.477f
C5365 a_n1986_8322.n3 gnd 1.24631f
C5366 a_n1986_8322.t16 gnd 0.124841p
C5367 a_n1986_8322.t13 gnd 0.093529f
C5368 a_n1986_8322.t10 gnd 0.875759f
C5369 a_n1986_8322.t2 gnd 0.093529f
C5370 a_n1986_8322.t8 gnd 0.093529f
C5371 a_n1986_8322.n4 gnd 0.65882f
C5372 a_n1986_8322.t15 gnd 0.093529f
C5373 a_n1986_8322.t9 gnd 0.093529f
C5374 a_n1986_8322.n5 gnd 0.65882f
C5375 a_n1986_8322.t14 gnd 0.874017f
C5376 a_n1986_8322.n6 gnd 0.766493f
C5377 a_n1986_8322.n7 gnd 3.48702f
C5378 a_n1986_8322.t5 gnd 0.875761f
C5379 a_n1986_8322.t6 gnd 0.093529f
C5380 a_n1986_8322.t1 gnd 0.093529f
C5381 a_n1986_8322.n8 gnd 0.65882f
C5382 a_n1986_8322.t19 gnd 0.093529f
C5383 a_n1986_8322.t11 gnd 0.093529f
C5384 a_n1986_8322.n9 gnd 0.65882f
C5385 a_n1986_8322.t17 gnd 0.874017f
C5386 a_n1986_8322.n10 gnd 1.39891f
C5387 a_n1986_8322.n11 gnd 1.59065f
C5388 a_n1986_8322.t3 gnd 0.874017f
C5389 a_n1986_8322.t12 gnd 0.875761f
C5390 a_n1986_8322.t7 gnd 0.093529f
C5391 a_n1986_8322.t4 gnd 0.093529f
C5392 a_n1986_8322.n12 gnd 0.65882f
C5393 a_n1986_8322.t18 gnd 0.874017f
C5394 a_n1986_8322.t20 gnd 0.874017f
C5395 a_n1986_8322.n13 gnd 0.658822f
C5396 a_n1986_8322.t0 gnd 0.093529f
C5397 CSoutput.n0 gnd 0.044735f
C5398 CSoutput.t173 gnd 0.295914f
C5399 CSoutput.n1 gnd 0.13362f
C5400 CSoutput.n2 gnd 0.044735f
C5401 CSoutput.t178 gnd 0.295914f
C5402 CSoutput.n3 gnd 0.035456f
C5403 CSoutput.n4 gnd 0.044735f
C5404 CSoutput.t166 gnd 0.295914f
C5405 CSoutput.n5 gnd 0.030574f
C5406 CSoutput.n6 gnd 0.044735f
C5407 CSoutput.t176 gnd 0.295914f
C5408 CSoutput.t174 gnd 0.295914f
C5409 CSoutput.n7 gnd 0.132163f
C5410 CSoutput.n8 gnd 0.044735f
C5411 CSoutput.t165 gnd 0.295914f
C5412 CSoutput.n9 gnd 0.029151f
C5413 CSoutput.n10 gnd 0.044735f
C5414 CSoutput.t170 gnd 0.295914f
C5415 CSoutput.t172 gnd 0.295914f
C5416 CSoutput.n11 gnd 0.132163f
C5417 CSoutput.n12 gnd 0.044735f
C5418 CSoutput.t161 gnd 0.295914f
C5419 CSoutput.n13 gnd 0.030574f
C5420 CSoutput.n14 gnd 0.044735f
C5421 CSoutput.t181 gnd 0.295914f
C5422 CSoutput.t171 gnd 0.295914f
C5423 CSoutput.n15 gnd 0.132163f
C5424 CSoutput.n16 gnd 0.044735f
C5425 CSoutput.t175 gnd 0.295914f
C5426 CSoutput.n17 gnd 0.032655f
C5427 CSoutput.t162 gnd 0.353624f
C5428 CSoutput.t179 gnd 0.295914f
C5429 CSoutput.n18 gnd 0.168721f
C5430 CSoutput.n19 gnd 0.163718f
C5431 CSoutput.n20 gnd 0.189933f
C5432 CSoutput.n21 gnd 0.044735f
C5433 CSoutput.n22 gnd 0.037336f
C5434 CSoutput.n23 gnd 0.132163f
C5435 CSoutput.n24 gnd 0.035991f
C5436 CSoutput.n25 gnd 0.035456f
C5437 CSoutput.n26 gnd 0.044735f
C5438 CSoutput.n27 gnd 0.044735f
C5439 CSoutput.n28 gnd 0.037049f
C5440 CSoutput.n29 gnd 0.031456f
C5441 CSoutput.n30 gnd 0.135106f
C5442 CSoutput.n31 gnd 0.031889f
C5443 CSoutput.n32 gnd 0.044735f
C5444 CSoutput.n33 gnd 0.044735f
C5445 CSoutput.n34 gnd 0.044735f
C5446 CSoutput.n35 gnd 0.036655f
C5447 CSoutput.n36 gnd 0.132163f
C5448 CSoutput.n37 gnd 0.035055f
C5449 CSoutput.n38 gnd 0.036393f
C5450 CSoutput.n39 gnd 0.044735f
C5451 CSoutput.n40 gnd 0.044735f
C5452 CSoutput.n41 gnd 0.037329f
C5453 CSoutput.n42 gnd 0.034119f
C5454 CSoutput.n43 gnd 0.132163f
C5455 CSoutput.n44 gnd 0.034984f
C5456 CSoutput.n45 gnd 0.044735f
C5457 CSoutput.n46 gnd 0.044735f
C5458 CSoutput.n47 gnd 0.044735f
C5459 CSoutput.n48 gnd 0.034984f
C5460 CSoutput.n49 gnd 0.132163f
C5461 CSoutput.n50 gnd 0.034119f
C5462 CSoutput.n51 gnd 0.037329f
C5463 CSoutput.n52 gnd 0.044735f
C5464 CSoutput.n53 gnd 0.044735f
C5465 CSoutput.n54 gnd 0.036393f
C5466 CSoutput.n55 gnd 0.035055f
C5467 CSoutput.n56 gnd 0.132163f
C5468 CSoutput.n57 gnd 0.036655f
C5469 CSoutput.n58 gnd 0.044735f
C5470 CSoutput.n59 gnd 0.044735f
C5471 CSoutput.n60 gnd 0.044735f
C5472 CSoutput.n61 gnd 0.031889f
C5473 CSoutput.n62 gnd 0.135106f
C5474 CSoutput.n63 gnd 0.031456f
C5475 CSoutput.t177 gnd 0.295914f
C5476 CSoutput.n64 gnd 0.132163f
C5477 CSoutput.n65 gnd 0.037049f
C5478 CSoutput.n66 gnd 0.044735f
C5479 CSoutput.n67 gnd 0.044735f
C5480 CSoutput.n68 gnd 0.044735f
C5481 CSoutput.n69 gnd 0.035991f
C5482 CSoutput.n70 gnd 0.132163f
C5483 CSoutput.n71 gnd 0.037336f
C5484 CSoutput.n72 gnd 0.032655f
C5485 CSoutput.n73 gnd 0.044735f
C5486 CSoutput.n74 gnd 0.044735f
C5487 CSoutput.n75 gnd 0.033865f
C5488 CSoutput.n76 gnd 0.020113f
C5489 CSoutput.t164 gnd 0.33248f
C5490 CSoutput.n77 gnd 0.165163f
C5491 CSoutput.n78 gnd 0.706716f
C5492 CSoutput.t146 gnd 0.055801f
C5493 CSoutput.t55 gnd 0.055801f
C5494 CSoutput.n79 gnd 0.432029f
C5495 CSoutput.t105 gnd 0.055801f
C5496 CSoutput.t30 gnd 0.055801f
C5497 CSoutput.n80 gnd 0.431258f
C5498 CSoutput.n81 gnd 0.437727f
C5499 CSoutput.t44 gnd 0.055801f
C5500 CSoutput.t95 gnd 0.055801f
C5501 CSoutput.n82 gnd 0.431258f
C5502 CSoutput.n83 gnd 0.215693f
C5503 CSoutput.t14 gnd 0.055801f
C5504 CSoutput.t56 gnd 0.055801f
C5505 CSoutput.n84 gnd 0.431258f
C5506 CSoutput.n85 gnd 0.215693f
C5507 CSoutput.t68 gnd 0.055801f
C5508 CSoutput.t127 gnd 0.055801f
C5509 CSoutput.n86 gnd 0.431258f
C5510 CSoutput.n87 gnd 0.215693f
C5511 CSoutput.t7 gnd 0.055801f
C5512 CSoutput.t70 gnd 0.055801f
C5513 CSoutput.n88 gnd 0.431258f
C5514 CSoutput.n89 gnd 0.215693f
C5515 CSoutput.t143 gnd 0.055801f
C5516 CSoutput.t73 gnd 0.055801f
C5517 CSoutput.n90 gnd 0.431258f
C5518 CSoutput.n91 gnd 0.215693f
C5519 CSoutput.t135 gnd 0.055801f
C5520 CSoutput.t41 gnd 0.055801f
C5521 CSoutput.n92 gnd 0.431258f
C5522 CSoutput.n93 gnd 0.395531f
C5523 CSoutput.t155 gnd 0.055801f
C5524 CSoutput.t153 gnd 0.055801f
C5525 CSoutput.n94 gnd 0.432029f
C5526 CSoutput.t157 gnd 0.055801f
C5527 CSoutput.t152 gnd 0.055801f
C5528 CSoutput.n95 gnd 0.431258f
C5529 CSoutput.n96 gnd 0.437727f
C5530 CSoutput.t93 gnd 0.055801f
C5531 CSoutput.t61 gnd 0.055801f
C5532 CSoutput.n97 gnd 0.431258f
C5533 CSoutput.n98 gnd 0.215693f
C5534 CSoutput.t19 gnd 0.055801f
C5535 CSoutput.t53 gnd 0.055801f
C5536 CSoutput.n99 gnd 0.431258f
C5537 CSoutput.n100 gnd 0.215693f
C5538 CSoutput.t72 gnd 0.055801f
C5539 CSoutput.t43 gnd 0.055801f
C5540 CSoutput.n101 gnd 0.431258f
C5541 CSoutput.n102 gnd 0.215693f
C5542 CSoutput.t34 gnd 0.055801f
C5543 CSoutput.t66 gnd 0.055801f
C5544 CSoutput.n103 gnd 0.431258f
C5545 CSoutput.n104 gnd 0.215693f
C5546 CSoutput.t98 gnd 0.055801f
C5547 CSoutput.t52 gnd 0.055801f
C5548 CSoutput.n105 gnd 0.431258f
C5549 CSoutput.n106 gnd 0.215693f
C5550 CSoutput.t132 gnd 0.055801f
C5551 CSoutput.t130 gnd 0.055801f
C5552 CSoutput.n107 gnd 0.431258f
C5553 CSoutput.n108 gnd 0.321653f
C5554 CSoutput.n109 gnd 0.405602f
C5555 CSoutput.t65 gnd 0.055801f
C5556 CSoutput.t118 gnd 0.055801f
C5557 CSoutput.n110 gnd 0.432029f
C5558 CSoutput.t137 gnd 0.055801f
C5559 CSoutput.t104 gnd 0.055801f
C5560 CSoutput.n111 gnd 0.431258f
C5561 CSoutput.n112 gnd 0.437727f
C5562 CSoutput.t71 gnd 0.055801f
C5563 CSoutput.t99 gnd 0.055801f
C5564 CSoutput.n113 gnd 0.431258f
C5565 CSoutput.n114 gnd 0.215693f
C5566 CSoutput.t94 gnd 0.055801f
C5567 CSoutput.t116 gnd 0.055801f
C5568 CSoutput.n115 gnd 0.431258f
C5569 CSoutput.n116 gnd 0.215693f
C5570 CSoutput.t13 gnd 0.055801f
C5571 CSoutput.t147 gnd 0.055801f
C5572 CSoutput.n117 gnd 0.431258f
C5573 CSoutput.n118 gnd 0.215693f
C5574 CSoutput.t107 gnd 0.055801f
C5575 CSoutput.t82 gnd 0.055801f
C5576 CSoutput.n119 gnd 0.431258f
C5577 CSoutput.n120 gnd 0.215693f
C5578 CSoutput.t83 gnd 0.055801f
C5579 CSoutput.t85 gnd 0.055801f
C5580 CSoutput.n121 gnd 0.431258f
C5581 CSoutput.n122 gnd 0.215693f
C5582 CSoutput.t103 gnd 0.055801f
C5583 CSoutput.t158 gnd 0.055801f
C5584 CSoutput.n123 gnd 0.431258f
C5585 CSoutput.n124 gnd 0.321653f
C5586 CSoutput.n125 gnd 0.453359f
C5587 CSoutput.n126 gnd 8.323791f
C5588 CSoutput.n128 gnd 0.791357f
C5589 CSoutput.n129 gnd 0.593518f
C5590 CSoutput.n130 gnd 0.791357f
C5591 CSoutput.n131 gnd 0.791357f
C5592 CSoutput.n132 gnd 2.13058f
C5593 CSoutput.n133 gnd 0.791357f
C5594 CSoutput.n134 gnd 0.791357f
C5595 CSoutput.t168 gnd 0.989197f
C5596 CSoutput.n135 gnd 0.791357f
C5597 CSoutput.n136 gnd 0.791357f
C5598 CSoutput.n140 gnd 0.791357f
C5599 CSoutput.n144 gnd 0.791357f
C5600 CSoutput.n145 gnd 0.791357f
C5601 CSoutput.n147 gnd 0.791357f
C5602 CSoutput.n152 gnd 0.791357f
C5603 CSoutput.n154 gnd 0.791357f
C5604 CSoutput.n155 gnd 0.791357f
C5605 CSoutput.n157 gnd 0.791357f
C5606 CSoutput.n158 gnd 0.791357f
C5607 CSoutput.n160 gnd 0.791357f
C5608 CSoutput.t163 gnd 13.223499f
C5609 CSoutput.n162 gnd 0.791357f
C5610 CSoutput.n163 gnd 0.593518f
C5611 CSoutput.n164 gnd 0.791357f
C5612 CSoutput.n165 gnd 0.791357f
C5613 CSoutput.n166 gnd 2.13058f
C5614 CSoutput.n167 gnd 0.791357f
C5615 CSoutput.n168 gnd 0.791357f
C5616 CSoutput.t180 gnd 0.989197f
C5617 CSoutput.n169 gnd 0.791357f
C5618 CSoutput.n170 gnd 0.791357f
C5619 CSoutput.n174 gnd 0.791357f
C5620 CSoutput.n178 gnd 0.791357f
C5621 CSoutput.n179 gnd 0.791357f
C5622 CSoutput.n181 gnd 0.791357f
C5623 CSoutput.n186 gnd 0.791357f
C5624 CSoutput.n188 gnd 0.791357f
C5625 CSoutput.n189 gnd 0.791357f
C5626 CSoutput.n191 gnd 0.791357f
C5627 CSoutput.n192 gnd 0.791357f
C5628 CSoutput.n194 gnd 0.791357f
C5629 CSoutput.n195 gnd 0.593518f
C5630 CSoutput.n197 gnd 0.791357f
C5631 CSoutput.n198 gnd 0.593518f
C5632 CSoutput.n199 gnd 0.791357f
C5633 CSoutput.n200 gnd 0.791357f
C5634 CSoutput.n201 gnd 2.13058f
C5635 CSoutput.n202 gnd 0.791357f
C5636 CSoutput.n203 gnd 0.791357f
C5637 CSoutput.t160 gnd 0.989197f
C5638 CSoutput.n204 gnd 0.791357f
C5639 CSoutput.n205 gnd 2.13058f
C5640 CSoutput.n207 gnd 0.791357f
C5641 CSoutput.n208 gnd 0.791357f
C5642 CSoutput.n210 gnd 0.791357f
C5643 CSoutput.n211 gnd 0.791357f
C5644 CSoutput.t169 gnd 13.008f
C5645 CSoutput.t167 gnd 13.223499f
C5646 CSoutput.n217 gnd 2.4826f
C5647 CSoutput.n218 gnd 10.1132f
C5648 CSoutput.n219 gnd 10.536401f
C5649 CSoutput.n224 gnd 2.68933f
C5650 CSoutput.n230 gnd 0.791357f
C5651 CSoutput.n232 gnd 0.791357f
C5652 CSoutput.n234 gnd 0.791357f
C5653 CSoutput.n236 gnd 0.791357f
C5654 CSoutput.n238 gnd 0.791357f
C5655 CSoutput.n244 gnd 0.791357f
C5656 CSoutput.n251 gnd 1.45184f
C5657 CSoutput.n252 gnd 1.45184f
C5658 CSoutput.n253 gnd 0.791357f
C5659 CSoutput.n254 gnd 0.791357f
C5660 CSoutput.n256 gnd 0.593518f
C5661 CSoutput.n257 gnd 0.508295f
C5662 CSoutput.n259 gnd 0.593518f
C5663 CSoutput.n260 gnd 0.508295f
C5664 CSoutput.n261 gnd 0.593518f
C5665 CSoutput.n263 gnd 0.791357f
C5666 CSoutput.n265 gnd 2.13058f
C5667 CSoutput.n266 gnd 2.4826f
C5668 CSoutput.n267 gnd 9.30157f
C5669 CSoutput.n269 gnd 0.593518f
C5670 CSoutput.n270 gnd 1.52716f
C5671 CSoutput.n271 gnd 0.593518f
C5672 CSoutput.n273 gnd 0.791357f
C5673 CSoutput.n275 gnd 2.13058f
C5674 CSoutput.n276 gnd 4.64074f
C5675 CSoutput.t90 gnd 0.055801f
C5676 CSoutput.t125 gnd 0.055801f
C5677 CSoutput.n277 gnd 0.432029f
C5678 CSoutput.t2 gnd 0.055801f
C5679 CSoutput.t109 gnd 0.055801f
C5680 CSoutput.n278 gnd 0.431258f
C5681 CSoutput.n279 gnd 0.437727f
C5682 CSoutput.t108 gnd 0.055801f
C5683 CSoutput.t17 gnd 0.055801f
C5684 CSoutput.n280 gnd 0.431258f
C5685 CSoutput.n281 gnd 0.215693f
C5686 CSoutput.t29 gnd 0.055801f
C5687 CSoutput.t149 gnd 0.055801f
C5688 CSoutput.n282 gnd 0.431258f
C5689 CSoutput.n283 gnd 0.215693f
C5690 CSoutput.t60 gnd 0.055801f
C5691 CSoutput.t154 gnd 0.055801f
C5692 CSoutput.n284 gnd 0.431258f
C5693 CSoutput.n285 gnd 0.215693f
C5694 CSoutput.t100 gnd 0.055801f
C5695 CSoutput.t42 gnd 0.055801f
C5696 CSoutput.n286 gnd 0.431258f
C5697 CSoutput.n287 gnd 0.215693f
C5698 CSoutput.t4 gnd 0.055801f
C5699 CSoutput.t106 gnd 0.055801f
C5700 CSoutput.n288 gnd 0.431258f
C5701 CSoutput.n289 gnd 0.215693f
C5702 CSoutput.t10 gnd 0.055801f
C5703 CSoutput.t1 gnd 0.055801f
C5704 CSoutput.n290 gnd 0.431258f
C5705 CSoutput.n291 gnd 0.395531f
C5706 CSoutput.t126 gnd 0.055801f
C5707 CSoutput.t140 gnd 0.055801f
C5708 CSoutput.n292 gnd 0.432029f
C5709 CSoutput.t111 gnd 0.055801f
C5710 CSoutput.t139 gnd 0.055801f
C5711 CSoutput.n293 gnd 0.431258f
C5712 CSoutput.n294 gnd 0.437727f
C5713 CSoutput.t51 gnd 0.055801f
C5714 CSoutput.t63 gnd 0.055801f
C5715 CSoutput.n295 gnd 0.431258f
C5716 CSoutput.n296 gnd 0.215693f
C5717 CSoutput.t69 gnd 0.055801f
C5718 CSoutput.t86 gnd 0.055801f
C5719 CSoutput.n297 gnd 0.431258f
C5720 CSoutput.n298 gnd 0.215693f
C5721 CSoutput.t35 gnd 0.055801f
C5722 CSoutput.t36 gnd 0.055801f
C5723 CSoutput.n299 gnd 0.431258f
C5724 CSoutput.n300 gnd 0.215693f
C5725 CSoutput.t156 gnd 0.055801f
C5726 CSoutput.t67 gnd 0.055801f
C5727 CSoutput.n301 gnd 0.431258f
C5728 CSoutput.n302 gnd 0.215693f
C5729 CSoutput.t131 gnd 0.055801f
C5730 CSoutput.t87 gnd 0.055801f
C5731 CSoutput.n303 gnd 0.431258f
C5732 CSoutput.n304 gnd 0.215693f
C5733 CSoutput.t15 gnd 0.055801f
C5734 CSoutput.t18 gnd 0.055801f
C5735 CSoutput.n305 gnd 0.431258f
C5736 CSoutput.n306 gnd 0.321653f
C5737 CSoutput.n307 gnd 0.405602f
C5738 CSoutput.t5 gnd 0.055801f
C5739 CSoutput.t141 gnd 0.055801f
C5740 CSoutput.n308 gnd 0.432029f
C5741 CSoutput.t159 gnd 0.055801f
C5742 CSoutput.t124 gnd 0.055801f
C5743 CSoutput.n309 gnd 0.431258f
C5744 CSoutput.n310 gnd 0.437727f
C5745 CSoutput.t101 gnd 0.055801f
C5746 CSoutput.t57 gnd 0.055801f
C5747 CSoutput.n311 gnd 0.431258f
C5748 CSoutput.n312 gnd 0.215693f
C5749 CSoutput.t77 gnd 0.055801f
C5750 CSoutput.t12 gnd 0.055801f
C5751 CSoutput.n313 gnd 0.431258f
C5752 CSoutput.n314 gnd 0.215693f
C5753 CSoutput.t97 gnd 0.055801f
C5754 CSoutput.t62 gnd 0.055801f
C5755 CSoutput.n315 gnd 0.431258f
C5756 CSoutput.n316 gnd 0.215693f
C5757 CSoutput.t28 gnd 0.055801f
C5758 CSoutput.t88 gnd 0.055801f
C5759 CSoutput.n317 gnd 0.431258f
C5760 CSoutput.n318 gnd 0.215693f
C5761 CSoutput.t151 gnd 0.055801f
C5762 CSoutput.t150 gnd 0.055801f
C5763 CSoutput.n319 gnd 0.431258f
C5764 CSoutput.n320 gnd 0.215693f
C5765 CSoutput.t145 gnd 0.055801f
C5766 CSoutput.t16 gnd 0.055801f
C5767 CSoutput.n321 gnd 0.431257f
C5768 CSoutput.n322 gnd 0.321654f
C5769 CSoutput.n323 gnd 0.453359f
C5770 CSoutput.n324 gnd 11.9024f
C5771 CSoutput.t9 gnd 0.048826f
C5772 CSoutput.t31 gnd 0.048826f
C5773 CSoutput.n325 gnd 0.432885f
C5774 CSoutput.t115 gnd 0.048826f
C5775 CSoutput.t120 gnd 0.048826f
C5776 CSoutput.n326 gnd 0.431441f
C5777 CSoutput.n327 gnd 0.402023f
C5778 CSoutput.t114 gnd 0.048826f
C5779 CSoutput.t142 gnd 0.048826f
C5780 CSoutput.n328 gnd 0.431441f
C5781 CSoutput.n329 gnd 0.198178f
C5782 CSoutput.t48 gnd 0.048826f
C5783 CSoutput.t96 gnd 0.048826f
C5784 CSoutput.n330 gnd 0.431441f
C5785 CSoutput.n331 gnd 0.198178f
C5786 CSoutput.t136 gnd 0.048826f
C5787 CSoutput.t138 gnd 0.048826f
C5788 CSoutput.n332 gnd 0.431441f
C5789 CSoutput.n333 gnd 0.198178f
C5790 CSoutput.t134 gnd 0.048826f
C5791 CSoutput.t112 gnd 0.048826f
C5792 CSoutput.n334 gnd 0.431441f
C5793 CSoutput.n335 gnd 0.198178f
C5794 CSoutput.t64 gnd 0.048826f
C5795 CSoutput.t123 gnd 0.048826f
C5796 CSoutput.n336 gnd 0.431441f
C5797 CSoutput.n337 gnd 0.198178f
C5798 CSoutput.t6 gnd 0.048826f
C5799 CSoutput.t148 gnd 0.048826f
C5800 CSoutput.n338 gnd 0.431441f
C5801 CSoutput.n339 gnd 0.365481f
C5802 CSoutput.t22 gnd 0.048826f
C5803 CSoutput.t33 gnd 0.048826f
C5804 CSoutput.n340 gnd 0.432885f
C5805 CSoutput.t49 gnd 0.048826f
C5806 CSoutput.t133 gnd 0.048826f
C5807 CSoutput.n341 gnd 0.431441f
C5808 CSoutput.n342 gnd 0.402023f
C5809 CSoutput.t59 gnd 0.048826f
C5810 CSoutput.t32 gnd 0.048826f
C5811 CSoutput.n343 gnd 0.431441f
C5812 CSoutput.n344 gnd 0.198178f
C5813 CSoutput.t80 gnd 0.048826f
C5814 CSoutput.t119 gnd 0.048826f
C5815 CSoutput.n345 gnd 0.431441f
C5816 CSoutput.n346 gnd 0.198178f
C5817 CSoutput.t40 gnd 0.048826f
C5818 CSoutput.t78 gnd 0.048826f
C5819 CSoutput.n347 gnd 0.431441f
C5820 CSoutput.n348 gnd 0.198178f
C5821 CSoutput.t0 gnd 0.048826f
C5822 CSoutput.t76 gnd 0.048826f
C5823 CSoutput.n349 gnd 0.431441f
C5824 CSoutput.n350 gnd 0.198178f
C5825 CSoutput.t122 gnd 0.048826f
C5826 CSoutput.t26 gnd 0.048826f
C5827 CSoutput.n351 gnd 0.431441f
C5828 CSoutput.n352 gnd 0.198178f
C5829 CSoutput.t46 gnd 0.048826f
C5830 CSoutput.t74 gnd 0.048826f
C5831 CSoutput.n353 gnd 0.431441f
C5832 CSoutput.n354 gnd 0.300877f
C5833 CSoutput.n355 gnd 0.559052f
C5834 CSoutput.n356 gnd 12.459901f
C5835 CSoutput.t91 gnd 0.048826f
C5836 CSoutput.t92 gnd 0.048826f
C5837 CSoutput.n357 gnd 0.432885f
C5838 CSoutput.t27 gnd 0.048826f
C5839 CSoutput.t117 gnd 0.048826f
C5840 CSoutput.n358 gnd 0.431441f
C5841 CSoutput.n359 gnd 0.402023f
C5842 CSoutput.t89 gnd 0.048826f
C5843 CSoutput.t24 gnd 0.048826f
C5844 CSoutput.n360 gnd 0.431441f
C5845 CSoutput.n361 gnd 0.198178f
C5846 CSoutput.t102 gnd 0.048826f
C5847 CSoutput.t128 gnd 0.048826f
C5848 CSoutput.n362 gnd 0.431441f
C5849 CSoutput.n363 gnd 0.198178f
C5850 CSoutput.t75 gnd 0.048826f
C5851 CSoutput.t25 gnd 0.048826f
C5852 CSoutput.n364 gnd 0.431441f
C5853 CSoutput.n365 gnd 0.198178f
C5854 CSoutput.t20 gnd 0.048826f
C5855 CSoutput.t8 gnd 0.048826f
C5856 CSoutput.n366 gnd 0.431441f
C5857 CSoutput.n367 gnd 0.198178f
C5858 CSoutput.t129 gnd 0.048826f
C5859 CSoutput.t47 gnd 0.048826f
C5860 CSoutput.n368 gnd 0.431441f
C5861 CSoutput.n369 gnd 0.198178f
C5862 CSoutput.t38 gnd 0.048826f
C5863 CSoutput.t121 gnd 0.048826f
C5864 CSoutput.n370 gnd 0.431441f
C5865 CSoutput.n371 gnd 0.365481f
C5866 CSoutput.t84 gnd 0.048826f
C5867 CSoutput.t45 gnd 0.048826f
C5868 CSoutput.n372 gnd 0.432885f
C5869 CSoutput.t54 gnd 0.048826f
C5870 CSoutput.t50 gnd 0.048826f
C5871 CSoutput.n373 gnd 0.431441f
C5872 CSoutput.n374 gnd 0.402023f
C5873 CSoutput.t23 gnd 0.048826f
C5874 CSoutput.t11 gnd 0.048826f
C5875 CSoutput.n375 gnd 0.431441f
C5876 CSoutput.n376 gnd 0.198178f
C5877 CSoutput.t21 gnd 0.048826f
C5878 CSoutput.t113 gnd 0.048826f
C5879 CSoutput.n377 gnd 0.431441f
C5880 CSoutput.n378 gnd 0.198178f
C5881 CSoutput.t110 gnd 0.048826f
C5882 CSoutput.t3 gnd 0.048826f
C5883 CSoutput.n379 gnd 0.431441f
C5884 CSoutput.n380 gnd 0.198178f
C5885 CSoutput.t58 gnd 0.048826f
C5886 CSoutput.t144 gnd 0.048826f
C5887 CSoutput.n381 gnd 0.431441f
C5888 CSoutput.n382 gnd 0.198178f
C5889 CSoutput.t81 gnd 0.048826f
C5890 CSoutput.t37 gnd 0.048826f
C5891 CSoutput.n383 gnd 0.431441f
C5892 CSoutput.n384 gnd 0.198178f
C5893 CSoutput.t39 gnd 0.048826f
C5894 CSoutput.t79 gnd 0.048826f
C5895 CSoutput.n385 gnd 0.431441f
C5896 CSoutput.n386 gnd 0.300877f
C5897 CSoutput.n387 gnd 0.559052f
C5898 CSoutput.n388 gnd 7.18565f
C5899 CSoutput.n389 gnd 14.439799f
.ends

