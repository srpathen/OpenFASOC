* NGSPICE file created from opamp307.ext - technology: sky130A

.subckt opamp307 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n8300_8799.t37 plus.t5 a_n3827_n3924.t48 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t124 a_n8300_8799.t40 vdd.t176 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t15 a_n2408_n452.t19 a_n2408_n452.t20 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2140_13878.t23 a_n2408_n452.t56 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 gnd.t167 gnd.t165 gnd.t166 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 vdd.t175 a_n8300_8799.t41 CSoutput.t123 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 gnd.t164 gnd.t162 minus.t4 gnd.t163 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X7 CSoutput.t122 a_n8300_8799.t42 vdd.t174 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X8 gnd.t286 commonsourceibias.t64 CSoutput.t175 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 a_n3827_n3924.t1 diffpairibias.t20 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 CSoutput.t121 a_n8300_8799.t43 vdd.t173 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 a_n3827_n3924.t42 plus.t6 a_n8300_8799.t36 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X12 commonsourceibias.t63 commonsourceibias.t62 gnd.t280 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t161 gnd.t159 gnd.t160 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X14 a_n3827_n3924.t4 minus.t5 a_n2408_n452.t3 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X15 vdd.t177 CSoutput.t184 output.t18 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X16 a_n2318_8322.t15 a_n2408_n452.t57 a_n8300_8799.t2 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t158 gnd.t156 gnd.t157 gnd.t76 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X18 CSoutput.t130 commonsourceibias.t65 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t120 a_n8300_8799.t44 vdd.t172 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t195 commonsourceibias.t60 commonsourceibias.t61 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t128 commonsourceibias.t66 gnd.t41 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t171 a_n8300_8799.t45 CSoutput.t119 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 gnd.t155 gnd.t153 gnd.t154 gnd.t76 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X24 a_n2408_n452.t48 minus.t6 a_n3827_n3924.t22 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X25 commonsourceibias.t59 commonsourceibias.t58 gnd.t251 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n8300_8799.t3 a_n2408_n452.t58 a_n2318_8322.t14 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X27 CSoutput.t174 commonsourceibias.t67 gnd.t285 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 vdd.t170 a_n8300_8799.t46 CSoutput.t118 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 vdd.t169 a_n8300_8799.t47 CSoutput.t117 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 a_n2408_n452.t44 minus.t7 a_n3827_n3924.t15 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X31 CSoutput.t116 a_n8300_8799.t48 vdd.t168 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 vdd.t167 a_n8300_8799.t49 CSoutput.t115 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n8300_8799.t4 a_n2408_n452.t59 a_n2318_8322.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 commonsourceibias.t57 commonsourceibias.t56 gnd.t241 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 a_n3827_n3924.t56 minus.t8 a_n2408_n452.t55 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X36 vdd.t292 vdd.t290 vdd.t291 vdd.t218 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X37 gnd.t152 gnd.t150 gnd.t151 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 CSoutput.t185 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X39 CSoutput.t114 a_n8300_8799.t50 vdd.t166 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 CSoutput.t172 commonsourceibias.t68 gnd.t279 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n3827_n3924.t51 diffpairibias.t21 gnd.t304 gnd.t303 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 CSoutput.t113 a_n8300_8799.t51 vdd.t165 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X43 CSoutput.t112 a_n8300_8799.t52 vdd.t164 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 gnd.t149 gnd.t146 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X45 gnd.t221 commonsourceibias.t69 CSoutput.t152 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 vdd.t163 a_n8300_8799.t53 CSoutput.t111 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 gnd.t281 commonsourceibias.t54 commonsourceibias.t55 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X48 output.t17 CSoutput.t186 vdd.t178 gnd.t36 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X49 CSoutput.t110 a_n8300_8799.t54 vdd.t162 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 commonsourceibias.t53 commonsourceibias.t52 gnd.t307 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 a_n3827_n3924.t27 plus.t7 a_n8300_8799.t35 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X52 gnd.t278 commonsourceibias.t70 CSoutput.t171 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 a_n2140_13878.t14 a_n2408_n452.t9 a_n2408_n452.t10 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 a_n8300_8799.t34 plus.t8 a_n3827_n3924.t43 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X55 a_n2408_n452.t40 a_n2408_n452.t39 a_n2140_13878.t13 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X56 CSoutput.t187 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X57 gnd.t186 commonsourceibias.t71 CSoutput.t140 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 a_n8300_8799.t33 plus.t9 a_n3827_n3924.t45 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X59 CSoutput.t109 a_n8300_8799.t55 vdd.t161 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 output.t16 CSoutput.t188 vdd.t7 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X61 vdd.t289 vdd.t287 vdd.t288 vdd.t264 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 vdd.t160 a_n8300_8799.t56 CSoutput.t108 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 gnd.t242 commonsourceibias.t50 commonsourceibias.t51 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 diffpairibias.t19 diffpairibias.t18 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X65 a_n3827_n3924.t47 plus.t10 a_n8300_8799.t32 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X66 commonsourceibias.t49 commonsourceibias.t48 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 a_n2408_n452.t51 minus.t9 a_n3827_n3924.t52 gnd.t292 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X68 a_n8300_8799.t10 a_n2408_n452.t60 a_n2318_8322.t12 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X69 CSoutput.t107 a_n8300_8799.t57 vdd.t159 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 commonsourceibias.t47 commonsourceibias.t46 gnd.t245 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 gnd.t145 gnd.t143 plus.t0 gnd.t144 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X72 vdd.t158 a_n8300_8799.t58 CSoutput.t106 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 vdd.t157 a_n8300_8799.t59 CSoutput.t105 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 gnd.t142 gnd.t140 gnd.t141 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X75 diffpairibias.t17 diffpairibias.t16 gnd.t306 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 gnd.t308 commonsourceibias.t44 commonsourceibias.t45 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 CSoutput.t104 a_n8300_8799.t60 vdd.t156 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 CSoutput.t143 commonsourceibias.t72 gnd.t194 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 output.t1 outputibias.t8 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X80 vdd.t155 a_n8300_8799.t61 CSoutput.t103 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t102 a_n8300_8799.t62 vdd.t154 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 vdd.t286 vdd.t284 vdd.t285 vdd.t254 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X83 CSoutput.t101 a_n8300_8799.t63 vdd.t153 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X84 CSoutput.t100 a_n8300_8799.t64 vdd.t152 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 CSoutput.t99 a_n8300_8799.t65 vdd.t151 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t8 CSoutput.t189 output.t15 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X87 vdd.t9 CSoutput.t190 output.t14 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X88 gnd.t323 commonsourceibias.t42 commonsourceibias.t43 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t183 commonsourceibias.t73 gnd.t322 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t151 commonsourceibias.t74 gnd.t220 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t139 gnd.t137 gnd.t138 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X92 gnd.t136 gnd.t134 plus.t2 gnd.t135 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X93 a_n3827_n3924.t28 plus.t11 a_n8300_8799.t31 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X94 CSoutput.t133 commonsourceibias.t75 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 outputibias.t7 outputibias.t6 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X96 CSoutput.t155 commonsourceibias.t76 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 a_n3827_n3924.t5 diffpairibias.t22 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 vdd.t150 a_n8300_8799.t66 CSoutput.t98 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 vdd.t149 a_n8300_8799.t67 CSoutput.t97 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 a_n2408_n452.t34 a_n2408_n452.t33 a_n2140_13878.t12 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 vdd.t147 a_n8300_8799.t68 CSoutput.t96 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 vdd.t148 a_n8300_8799.t69 CSoutput.t95 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 a_n8300_8799.t11 a_n2408_n452.t61 a_n2318_8322.t11 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X104 vdd.t146 a_n8300_8799.t70 CSoutput.t94 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 a_n2408_n452.t12 a_n2408_n452.t11 a_n2140_13878.t11 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X106 gnd.t310 commonsourceibias.t40 commonsourceibias.t41 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 gnd.t327 commonsourceibias.t38 commonsourceibias.t39 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 vdd.t145 a_n8300_8799.t71 CSoutput.t93 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 CSoutput.t92 a_n8300_8799.t72 vdd.t144 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 diffpairibias.t15 diffpairibias.t14 gnd.t284 gnd.t283 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X111 a_n2408_n452.t4 minus.t10 a_n3827_n3924.t6 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X112 vdd.t283 vdd.t281 vdd.t282 vdd.t268 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 vdd.t280 vdd.t278 vdd.t279 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X114 CSoutput.t91 a_n8300_8799.t73 vdd.t143 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 gnd.t237 commonsourceibias.t77 CSoutput.t156 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 vdd.t277 vdd.t274 vdd.t276 vdd.t275 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 gnd.t297 commonsourceibias.t78 CSoutput.t177 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X118 gnd.t210 commonsourceibias.t79 CSoutput.t150 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t277 commonsourceibias.t80 CSoutput.t170 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 a_n3827_n3924.t23 minus.t11 a_n2408_n452.t49 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X121 CSoutput.t90 a_n8300_8799.t74 vdd.t142 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 output.t13 CSoutput.t191 vdd.t183 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X123 vdd.t141 a_n8300_8799.t75 CSoutput.t89 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 vdd.t184 CSoutput.t192 output.t12 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t207 a_n2408_n452.t62 a_n2318_8322.t23 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 a_n2408_n452.t14 a_n2408_n452.t13 a_n2140_13878.t10 vdd.t295 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X127 gnd.t316 commonsourceibias.t81 CSoutput.t181 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X128 vdd.t273 vdd.t271 vdd.t272 vdd.t254 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X129 gnd.t133 gnd.t131 gnd.t132 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X130 a_n2318_8322.t22 a_n2408_n452.t63 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 a_n3827_n3924.t57 diffpairibias.t23 gnd.t326 gnd.t325 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X132 CSoutput.t88 a_n8300_8799.t76 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 CSoutput.t87 a_n8300_8799.t77 vdd.t138 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 a_n3827_n3924.t12 minus.t12 a_n2408_n452.t41 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X135 a_n3827_n3924.t0 minus.t13 a_n2408_n452.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X136 vdd.t202 a_n2408_n452.t64 a_n2140_13878.t22 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 a_n2408_n452.t45 minus.t14 a_n3827_n3924.t16 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X138 a_n3827_n3924.t25 plus.t12 a_n8300_8799.t30 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X139 a_n3827_n3924.t31 plus.t13 a_n8300_8799.t29 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X140 gnd.t30 commonsourceibias.t82 CSoutput.t4 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t270 vdd.t267 vdd.t269 vdd.t268 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 a_n2408_n452.t6 minus.t15 a_n3827_n3924.t9 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X143 vdd.t137 a_n8300_8799.t78 CSoutput.t86 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 vdd.t135 a_n8300_8799.t79 CSoutput.t85 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 vdd.t134 a_n8300_8799.t80 CSoutput.t84 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 gnd.t130 gnd.t128 plus.t1 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X147 a_n8300_8799.t28 plus.t14 a_n3827_n3924.t34 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X148 a_n8300_8799.t27 plus.t15 a_n3827_n3924.t29 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X149 vdd.t266 vdd.t263 vdd.t265 vdd.t264 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 a_n2318_8322.t21 a_n2408_n452.t65 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X151 a_n8300_8799.t5 a_n2408_n452.t66 a_n2318_8322.t10 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 CSoutput.t83 a_n8300_8799.t81 vdd.t132 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X153 diffpairibias.t13 diffpairibias.t12 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X154 vdd.t131 a_n8300_8799.t82 CSoutput.t82 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 a_n2408_n452.t5 minus.t16 a_n3827_n3924.t8 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X156 a_n2408_n452.t32 a_n2408_n452.t31 a_n2140_13878.t9 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 vdd.t110 a_n8300_8799.t83 CSoutput.t81 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 a_n8300_8799.t6 a_n2408_n452.t67 a_n2318_8322.t9 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X159 CSoutput.t80 a_n8300_8799.t84 vdd.t129 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput.t161 commonsourceibias.t83 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n2140_13878.t8 a_n2408_n452.t35 a_n2408_n452.t36 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 commonsourceibias.t37 commonsourceibias.t36 gnd.t309 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 CSoutput.t142 commonsourceibias.t84 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 vdd.t262 vdd.t260 vdd.t261 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X165 a_n3827_n3924.t14 minus.t17 a_n2408_n452.t43 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X166 CSoutput.t169 commonsourceibias.t85 gnd.t276 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X167 vdd.t185 CSoutput.t193 output.t11 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X168 CSoutput.t149 commonsourceibias.t86 gnd.t209 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 gnd.t184 commonsourceibias.t87 CSoutput.t139 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 CSoutput.t79 a_n8300_8799.t85 vdd.t128 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 gnd.t324 commonsourceibias.t34 commonsourceibias.t35 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X173 vdd.t16 a_n2408_n452.t68 a_n2318_8322.t20 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X174 a_n2140_13878.t7 a_n2408_n452.t25 a_n2408_n452.t26 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X175 vdd.t127 a_n8300_8799.t86 CSoutput.t78 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X176 a_n2408_n452.t24 a_n2408_n452.t23 a_n2140_13878.t6 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 commonsourceibias.t33 commonsourceibias.t32 gnd.t311 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 gnd.t328 commonsourceibias.t30 commonsourceibias.t31 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 minus.t3 gnd.t121 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X180 a_n3827_n3924.t33 plus.t16 a_n8300_8799.t26 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X181 vdd.t126 a_n8300_8799.t87 CSoutput.t77 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 gnd.t329 commonsourceibias.t28 commonsourceibias.t29 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n3827_n3924.t21 diffpairibias.t24 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 commonsourceibias.t27 commonsourceibias.t26 gnd.t330 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n3827_n3924.t49 diffpairibias.t25 gnd.t300 gnd.t299 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 outputibias.t5 outputibias.t4 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X187 gnd.t182 commonsourceibias.t88 CSoutput.t138 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 vdd.t125 a_n8300_8799.t88 CSoutput.t76 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t124 a_n8300_8799.t89 CSoutput.t75 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X190 a_n8300_8799.t25 plus.t17 a_n3827_n3924.t26 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X191 gnd.t28 commonsourceibias.t89 CSoutput.t3 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t34 commonsourceibias.t90 CSoutput.t126 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 gnd.t8 commonsourceibias.t91 CSoutput.t0 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t43 commonsourceibias.t92 CSoutput.t129 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X195 CSoutput.t74 a_n8300_8799.t90 vdd.t123 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 commonsourceibias.t25 commonsourceibias.t24 gnd.t331 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 CSoutput.t73 a_n8300_8799.t91 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 outputibias.t3 outputibias.t2 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X199 CSoutput.t72 a_n8300_8799.t92 vdd.t120 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 gnd.t315 commonsourceibias.t93 CSoutput.t180 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 CSoutput.t2 commonsourceibias.t94 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 diffpairibias.t11 diffpairibias.t10 gnd.t240 gnd.t239 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 a_n2140_13878.t21 a_n2408_n452.t69 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 gnd.t256 commonsourceibias.t95 CSoutput.t160 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 vdd.t197 a_n2408_n452.t70 a_n2140_13878.t20 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 gnd.t232 commonsourceibias.t22 commonsourceibias.t23 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 CSoutput.t71 a_n8300_8799.t93 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 vdd.t117 a_n8300_8799.t94 CSoutput.t70 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 commonsourceibias.t21 commonsourceibias.t20 gnd.t223 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 vdd.t112 a_n8300_8799.t95 CSoutput.t69 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput.t141 commonsourceibias.t96 gnd.t191 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t68 a_n8300_8799.t96 vdd.t115 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 plus.t3 gnd.t118 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X214 a_n2140_13878.t5 a_n2408_n452.t29 a_n2408_n452.t30 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X215 diffpairibias.t9 diffpairibias.t8 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X216 a_n3827_n3924.t3 minus.t18 a_n2408_n452.t2 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X217 vdd.t114 a_n8300_8799.t97 CSoutput.t67 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 gnd.t226 commonsourceibias.t18 commonsourceibias.t19 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 CSoutput.t127 commonsourceibias.t97 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X220 a_n2408_n452.t8 minus.t19 a_n3827_n3924.t11 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X221 a_n2318_8322.t8 a_n2408_n452.t71 a_n8300_8799.t9 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 CSoutput.t66 a_n8300_8799.t98 vdd.t113 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 diffpairibias.t7 diffpairibias.t6 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 vdd.t109 a_n8300_8799.t99 CSoutput.t65 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 a_n2408_n452.t47 minus.t20 a_n3827_n3924.t20 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X226 a_n2408_n452.t42 minus.t21 a_n3827_n3924.t13 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X227 vdd.t259 vdd.t257 vdd.t258 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X228 vdd.t210 a_n2408_n452.t72 a_n2318_8322.t19 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X229 vdd.t107 a_n8300_8799.t100 CSoutput.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X230 vdd.t106 a_n8300_8799.t101 CSoutput.t63 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 a_n3827_n3924.t19 minus.t22 a_n2408_n452.t46 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X232 vdd.t186 CSoutput.t194 output.t10 gnd.t55 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X233 CSoutput.t195 a_n2318_8322.t27 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X234 CSoutput.t178 commonsourceibias.t98 gnd.t298 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n8300_8799.t24 plus.t18 a_n3827_n3924.t46 gnd.t292 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 CSoutput.t132 commonsourceibias.t99 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 gnd.t261 commonsourceibias.t100 CSoutput.t163 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 a_n3827_n3924.t24 minus.t23 a_n2408_n452.t50 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X239 CSoutput.t62 a_n8300_8799.t102 vdd.t104 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 gnd.t117 gnd.t114 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X241 a_n2140_13878.t19 a_n2408_n452.t73 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X242 outputibias.t1 outputibias.t0 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X243 vdd.t256 vdd.t253 vdd.t255 vdd.t254 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 CSoutput.t162 commonsourceibias.t101 gnd.t260 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 vdd.t252 vdd.t250 vdd.t251 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X246 commonsourceibias.t17 commonsourceibias.t16 gnd.t259 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X247 vdd.t103 a_n8300_8799.t103 CSoutput.t61 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t196 a_n2318_8322.t26 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X249 CSoutput.t60 a_n8300_8799.t104 vdd.t102 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t59 a_n8300_8799.t105 vdd.t101 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t58 a_n8300_8799.t106 vdd.t100 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 gnd.t113 gnd.t111 minus.t2 gnd.t112 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X253 gnd.t103 gnd.t101 gnd.t102 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 gnd.t110 gnd.t107 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X255 vdd.t99 a_n8300_8799.t107 CSoutput.t57 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X256 a_n3827_n3924.t50 diffpairibias.t26 gnd.t302 gnd.t301 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X257 vdd.t214 a_n2408_n452.t74 a_n2318_8322.t18 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X258 a_n2318_8322.t7 a_n2408_n452.t75 a_n8300_8799.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 CSoutput.t56 a_n8300_8799.t108 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 gnd.t282 commonsourceibias.t102 CSoutput.t173 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 vdd.t96 a_n8300_8799.t109 CSoutput.t55 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 CSoutput.t54 a_n8300_8799.t110 vdd.t95 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 vdd.t94 a_n8300_8799.t111 CSoutput.t53 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 vdd.t93 a_n8300_8799.t112 CSoutput.t52 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 a_n8300_8799.t23 plus.t19 a_n3827_n3924.t37 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X266 output.t2 outputibias.t9 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X267 gnd.t57 commonsourceibias.t103 CSoutput.t131 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 CSoutput.t179 commonsourceibias.t104 gnd.t314 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 vdd.t249 vdd.t247 vdd.t248 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X270 vdd.t246 vdd.t243 vdd.t245 vdd.t244 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X271 a_n3827_n3924.t40 plus.t20 a_n8300_8799.t22 gnd.t291 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X272 vdd.t92 a_n8300_8799.t113 CSoutput.t51 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t50 a_n8300_8799.t114 vdd.t91 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 gnd.t318 commonsourceibias.t105 CSoutput.t182 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2140_13878.t4 a_n2408_n452.t37 a_n2408_n452.t38 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 CSoutput.t49 a_n8300_8799.t115 vdd.t89 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t159 commonsourceibias.t106 gnd.t255 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 a_n2318_8322.t6 a_n2408_n452.t76 a_n8300_8799.t1 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X279 vdd.t242 vdd.t239 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X280 diffpairibias.t5 diffpairibias.t4 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X281 commonsourceibias.t15 commonsourceibias.t14 gnd.t319 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 gnd.t208 commonsourceibias.t107 CSoutput.t148 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 gnd.t106 gnd.t104 gnd.t105 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 CSoutput.t147 commonsourceibias.t108 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 gnd.t317 commonsourceibias.t12 commonsourceibias.t13 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t48 a_n8300_8799.t116 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 CSoutput.t47 a_n8300_8799.t117 vdd.t86 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t46 a_n8300_8799.t118 vdd.t84 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 a_n3827_n3924.t17 diffpairibias.t27 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X290 vdd.t83 a_n8300_8799.t119 CSoutput.t45 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 CSoutput.t137 commonsourceibias.t109 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 vdd.t82 a_n8300_8799.t120 CSoutput.t44 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 a_n2318_8322.t17 a_n2408_n452.t77 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 CSoutput.t43 a_n8300_8799.t121 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t42 a_n8300_8799.t122 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t157 commonsourceibias.t110 gnd.t238 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X297 vdd.t76 a_n8300_8799.t123 CSoutput.t41 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t238 vdd.t236 vdd.t237 vdd.t222 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X299 CSoutput.t40 a_n8300_8799.t124 vdd.t75 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X300 vdd.t190 a_n2408_n452.t78 a_n2140_13878.t18 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X301 gnd.t287 commonsourceibias.t10 commonsourceibias.t11 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 plus.t4 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X303 vdd.t74 a_n8300_8799.t125 CSoutput.t39 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t38 a_n8300_8799.t126 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 output.t9 CSoutput.t197 vdd.t192 gnd.t211 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X306 CSoutput.t158 commonsourceibias.t111 gnd.t250 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 CSoutput.t37 a_n8300_8799.t127 vdd.t70 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 gnd.t275 commonsourceibias.t112 CSoutput.t168 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 a_n3827_n3924.t36 plus.t21 a_n8300_8799.t21 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X310 vdd.t69 a_n8300_8799.t128 CSoutput.t36 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 vdd.t67 a_n8300_8799.t129 CSoutput.t35 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 CSoutput.t167 commonsourceibias.t113 gnd.t274 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 vdd.t235 vdd.t233 vdd.t234 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X314 commonsourceibias.t9 commonsourceibias.t8 gnd.t288 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X315 a_n3827_n3924.t53 minus.t24 a_n2408_n452.t52 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X316 a_n2318_8322.t5 a_n2408_n452.t79 a_n8300_8799.t7 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X317 CSoutput.t34 a_n8300_8799.t130 vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X318 CSoutput.t146 commonsourceibias.t114 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 a_n8300_8799.t8 a_n2408_n452.t80 a_n2318_8322.t4 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 output.t8 CSoutput.t198 vdd.t193 gnd.t212 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X321 gnd.t290 commonsourceibias.t6 commonsourceibias.t7 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 a_n8300_8799.t20 plus.t22 a_n3827_n3924.t38 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X323 vdd.t64 a_n8300_8799.t131 CSoutput.t33 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X324 a_n2140_13878.t17 a_n2408_n452.t81 vdd.t294 vdd.t293 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X325 gnd.t178 commonsourceibias.t115 CSoutput.t136 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 vdd.t62 a_n8300_8799.t132 CSoutput.t32 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 a_n2408_n452.t53 minus.t25 a_n3827_n3924.t54 gnd.t293 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X328 CSoutput.t31 a_n8300_8799.t133 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X330 commonsourceibias.t5 commonsourceibias.t4 gnd.t224 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 a_n8300_8799.t19 plus.t23 a_n3827_n3924.t44 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X332 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X333 gnd.t89 gnd.t87 minus.t1 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X334 a_n2318_8322.t3 a_n2408_n452.t82 a_n8300_8799.t12 vdd.t295 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 CSoutput.t199 a_n2318_8322.t25 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X336 a_n3827_n3924.t10 minus.t26 a_n2408_n452.t7 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X337 vdd.t59 a_n8300_8799.t134 CSoutput.t30 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 CSoutput.t29 a_n8300_8799.t135 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t28 a_n8300_8799.t136 vdd.t55 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 gnd.t227 commonsourceibias.t2 commonsourceibias.t3 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 CSoutput.t27 a_n8300_8799.t137 vdd.t54 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 a_n2140_13878.t3 a_n2408_n452.t21 a_n2408_n452.t22 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X343 a_n3827_n3924.t32 plus.t24 a_n8300_8799.t18 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X344 vdd.t53 a_n8300_8799.t138 CSoutput.t26 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 gnd.t176 commonsourceibias.t116 CSoutput.t135 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 CSoutput.t1 commonsourceibias.t117 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 vdd.t232 vdd.t229 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X348 vdd.t228 vdd.t225 vdd.t227 vdd.t226 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X349 output.t7 CSoutput.t200 vdd.t181 gnd.t44 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X350 gnd.t229 commonsourceibias.t118 CSoutput.t153 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 a_n3827_n3924.t18 diffpairibias.t28 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X352 vdd.t49 a_n8300_8799.t139 CSoutput.t25 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 vdd.t52 a_n8300_8799.t140 CSoutput.t24 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 gnd.t86 gnd.t83 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X355 CSoutput.t23 a_n8300_8799.t141 vdd.t51 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 gnd.t82 gnd.t79 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X357 a_n2408_n452.t28 a_n2408_n452.t27 a_n2140_13878.t2 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X358 gnd.t78 gnd.t75 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X359 a_n8300_8799.t13 a_n2408_n452.t83 a_n2318_8322.t2 vdd.t215 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X360 output.t19 outputibias.t10 gnd.t269 gnd.t268 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X361 vdd.t50 a_n8300_8799.t142 CSoutput.t22 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 gnd.t231 commonsourceibias.t119 CSoutput.t154 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 CSoutput.t21 a_n8300_8799.t143 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 a_n8300_8799.t17 plus.t25 a_n3827_n3924.t39 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X365 vdd.t182 CSoutput.t201 output.t6 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X366 vdd.t46 a_n8300_8799.t144 CSoutput.t20 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 gnd.t74 gnd.t71 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X368 CSoutput.t125 commonsourceibias.t120 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 CSoutput.t176 commonsourceibias.t121 gnd.t296 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 diffpairibias.t3 diffpairibias.t2 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X371 vdd.t45 a_n8300_8799.t145 CSoutput.t19 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 CSoutput.t18 a_n8300_8799.t146 vdd.t43 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 output.t0 outputibias.t11 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X374 CSoutput.t17 a_n8300_8799.t147 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 a_n2318_8322.t1 a_n2408_n452.t84 a_n8300_8799.t38 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X376 a_n3827_n3924.t30 plus.t26 a_n8300_8799.t16 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X377 vdd.t40 a_n8300_8799.t148 CSoutput.t16 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 CSoutput.t15 a_n8300_8799.t149 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X379 diffpairibias.t1 diffpairibias.t0 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X380 a_n3827_n3924.t41 plus.t27 a_n8300_8799.t15 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X381 CSoutput.t145 commonsourceibias.t122 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 CSoutput.t202 a_n2318_8322.t24 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X383 vdd.t224 vdd.t221 vdd.t223 vdd.t222 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X384 vdd.t299 a_n2408_n452.t85 a_n2140_13878.t16 vdd.t298 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X385 gnd.t273 commonsourceibias.t123 CSoutput.t166 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 a_n8300_8799.t14 plus.t28 a_n3827_n3924.t35 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X387 CSoutput.t14 a_n8300_8799.t150 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X389 vdd.t220 vdd.t217 vdd.t219 vdd.t218 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X390 gnd.t70 gnd.t67 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X391 a_n3827_n3924.t55 minus.t27 a_n2408_n452.t54 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X392 vdd.t4 CSoutput.t203 output.t5 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X393 vdd.t34 a_n8300_8799.t151 CSoutput.t13 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 vdd.t32 a_n8300_8799.t152 CSoutput.t12 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 CSoutput.t144 commonsourceibias.t124 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 CSoutput.t11 a_n8300_8799.t153 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 output.t4 CSoutput.t204 vdd.t5 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X398 gnd.t175 commonsourceibias.t125 CSoutput.t134 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 a_n2408_n452.t1 minus.t28 a_n3827_n3924.t2 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X400 gnd.t271 commonsourceibias.t126 CSoutput.t165 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 a_n2318_8322.t0 a_n2408_n452.t86 a_n8300_8799.t39 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X402 vdd.t28 a_n8300_8799.t154 CSoutput.t10 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 vdd.t26 a_n8300_8799.t155 CSoutput.t9 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X404 vdd.t20 a_n8300_8799.t156 CSoutput.t8 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 CSoutput.t7 a_n8300_8799.t157 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 output.t3 CSoutput.t205 vdd.t6 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X407 gnd.t270 commonsourceibias.t127 CSoutput.t164 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 a_n2318_8322.t16 a_n2408_n452.t87 vdd.t297 vdd.t296 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X409 a_n2140_13878.t1 a_n2408_n452.t17 a_n2408_n452.t18 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X410 vdd.t22 a_n8300_8799.t158 CSoutput.t6 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X411 minus.t0 gnd.t60 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X412 commonsourceibias.t1 commonsourceibias.t0 gnd.t230 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 a_n3827_n3924.t7 diffpairibias.t29 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X414 CSoutput.t5 a_n8300_8799.t159 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 a_n2408_n452.t16 a_n2408_n452.t15 a_n2140_13878.t0 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t1 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t2 19.8005
R93 plus.n85 plus.t3 19.8005
R94 plus.n87 plus.t0 19.8005
R95 plus.n87 plus.t4 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 14.8628
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n3827_n3924.n9 a_n3827_n3924.t1 214.994
R160 a_n3827_n3924.n6 a_n3827_n3924.t17 214.786
R161 a_n3827_n3924.n6 a_n3827_n3924.t57 214.321
R162 a_n3827_n3924.n6 a_n3827_n3924.t18 214.321
R163 a_n3827_n3924.n6 a_n3827_n3924.t49 214.321
R164 a_n3827_n3924.n8 a_n3827_n3924.t7 214.321
R165 a_n3827_n3924.n8 a_n3827_n3924.t21 214.321
R166 a_n3827_n3924.n7 a_n3827_n3924.t51 214.321
R167 a_n3827_n3924.n9 a_n3827_n3924.t5 214.321
R168 a_n3827_n3924.n9 a_n3827_n3924.t50 214.321
R169 a_n3827_n3924.n1 a_n3827_n3924.t40 55.8337
R170 a_n3827_n3924.n1 a_n3827_n3924.t2 55.8337
R171 a_n3827_n3924.t0 a_n3827_n3924.n12 55.8337
R172 a_n3827_n3924.n0 a_n3827_n3924.t43 55.8335
R173 a_n3827_n3924.n10 a_n3827_n3924.t11 55.8335
R174 a_n3827_n3924.n4 a_n3827_n3924.t56 55.8335
R175 a_n3827_n3924.n4 a_n3827_n3924.t29 55.8335
R176 a_n3827_n3924.n3 a_n3827_n3924.t36 55.8335
R177 a_n3827_n3924.n0 a_n3827_n3924.n24 53.0052
R178 a_n3827_n3924.n0 a_n3827_n3924.n25 53.0052
R179 a_n3827_n3924.n0 a_n3827_n3924.n26 53.0052
R180 a_n3827_n3924.n1 a_n3827_n3924.n27 53.0052
R181 a_n3827_n3924.n1 a_n3827_n3924.n28 53.0052
R182 a_n3827_n3924.n1 a_n3827_n3924.n29 53.0052
R183 a_n3827_n3924.n1 a_n3827_n3924.n30 53.0052
R184 a_n3827_n3924.n11 a_n3827_n3924.n31 53.0052
R185 a_n3827_n3924.n11 a_n3827_n3924.n32 53.0052
R186 a_n3827_n3924.n12 a_n3827_n3924.n33 53.0052
R187 a_n3827_n3924.n10 a_n3827_n3924.n22 53.0051
R188 a_n3827_n3924.n2 a_n3827_n3924.n21 53.0051
R189 a_n3827_n3924.n2 a_n3827_n3924.n20 53.0051
R190 a_n3827_n3924.n2 a_n3827_n3924.n19 53.0051
R191 a_n3827_n3924.n2 a_n3827_n3924.n18 53.0051
R192 a_n3827_n3924.n4 a_n3827_n3924.n17 53.0051
R193 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0051
R194 a_n3827_n3924.n4 a_n3827_n3924.n15 53.0051
R195 a_n3827_n3924.n3 a_n3827_n3924.n14 53.0051
R196 a_n3827_n3924.n3 a_n3827_n3924.n13 53.0051
R197 a_n3827_n3924.n12 a_n3827_n3924.n5 12.1986
R198 a_n3827_n3924.n0 a_n3827_n3924.n23 12.1986
R199 a_n3827_n3924.n3 a_n3827_n3924.n5 5.11903
R200 a_n3827_n3924.n23 a_n3827_n3924.n10 5.11903
R201 a_n3827_n3924.n24 a_n3827_n3924.t35 2.82907
R202 a_n3827_n3924.n24 a_n3827_n3924.t47 2.82907
R203 a_n3827_n3924.n25 a_n3827_n3924.t34 2.82907
R204 a_n3827_n3924.n25 a_n3827_n3924.t25 2.82907
R205 a_n3827_n3924.n26 a_n3827_n3924.t45 2.82907
R206 a_n3827_n3924.n26 a_n3827_n3924.t27 2.82907
R207 a_n3827_n3924.n27 a_n3827_n3924.t39 2.82907
R208 a_n3827_n3924.n27 a_n3827_n3924.t41 2.82907
R209 a_n3827_n3924.n28 a_n3827_n3924.t37 2.82907
R210 a_n3827_n3924.n28 a_n3827_n3924.t30 2.82907
R211 a_n3827_n3924.n29 a_n3827_n3924.t52 2.82907
R212 a_n3827_n3924.n29 a_n3827_n3924.t55 2.82907
R213 a_n3827_n3924.n30 a_n3827_n3924.t8 2.82907
R214 a_n3827_n3924.n30 a_n3827_n3924.t14 2.82907
R215 a_n3827_n3924.n31 a_n3827_n3924.t13 2.82907
R216 a_n3827_n3924.n31 a_n3827_n3924.t24 2.82907
R217 a_n3827_n3924.n32 a_n3827_n3924.t22 2.82907
R218 a_n3827_n3924.n32 a_n3827_n3924.t10 2.82907
R219 a_n3827_n3924.n33 a_n3827_n3924.t9 2.82907
R220 a_n3827_n3924.n33 a_n3827_n3924.t4 2.82907
R221 a_n3827_n3924.n22 a_n3827_n3924.t16 2.82907
R222 a_n3827_n3924.n22 a_n3827_n3924.t19 2.82907
R223 a_n3827_n3924.n21 a_n3827_n3924.t54 2.82907
R224 a_n3827_n3924.n21 a_n3827_n3924.t53 2.82907
R225 a_n3827_n3924.n20 a_n3827_n3924.t20 2.82907
R226 a_n3827_n3924.n20 a_n3827_n3924.t3 2.82907
R227 a_n3827_n3924.n19 a_n3827_n3924.t6 2.82907
R228 a_n3827_n3924.n19 a_n3827_n3924.t12 2.82907
R229 a_n3827_n3924.n18 a_n3827_n3924.t15 2.82907
R230 a_n3827_n3924.n18 a_n3827_n3924.t23 2.82907
R231 a_n3827_n3924.n17 a_n3827_n3924.t46 2.82907
R232 a_n3827_n3924.n17 a_n3827_n3924.t31 2.82907
R233 a_n3827_n3924.n16 a_n3827_n3924.t44 2.82907
R234 a_n3827_n3924.n16 a_n3827_n3924.t32 2.82907
R235 a_n3827_n3924.n15 a_n3827_n3924.t48 2.82907
R236 a_n3827_n3924.n15 a_n3827_n3924.t42 2.82907
R237 a_n3827_n3924.n14 a_n3827_n3924.t26 2.82907
R238 a_n3827_n3924.n14 a_n3827_n3924.t28 2.82907
R239 a_n3827_n3924.n13 a_n3827_n3924.t38 2.82907
R240 a_n3827_n3924.n13 a_n3827_n3924.t33 2.82907
R241 a_n3827_n3924.n1 a_n3827_n3924.n0 2.66429
R242 a_n3827_n3924.n6 a_n3827_n3924.n8 2.22216
R243 a_n3827_n3924.n2 a_n3827_n3924.n4 2.01128
R244 a_n3827_n3924.n23 a_n3827_n3924.n6 1.95694
R245 a_n3827_n3924.n9 a_n3827_n3924.n5 1.95694
R246 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R247 a_n3827_n3924.n10 a_n3827_n3924.n2 1.77636
R248 a_n3827_n3924.n11 a_n3827_n3924.n1 1.56731
R249 a_n3827_n3924.n8 a_n3827_n3924.n7 1.34352
R250 a_n3827_n3924.n7 a_n3827_n3924.n9 1.34352
R251 a_n3827_n3924.n12 a_n3827_n3924.n11 1.3324
R252 a_n8300_8799.n223 a_n8300_8799.t149 485.149
R253 a_n8300_8799.n285 a_n8300_8799.t42 485.149
R254 a_n8300_8799.n348 a_n8300_8799.t124 485.149
R255 a_n8300_8799.n33 a_n8300_8799.t107 485.149
R256 a_n8300_8799.n95 a_n8300_8799.t123 485.149
R257 a_n8300_8799.n158 a_n8300_8799.t125 485.149
R258 a_n8300_8799.n266 a_n8300_8799.t89 464.166
R259 a_n8300_8799.n265 a_n8300_8799.t65 464.166
R260 a_n8300_8799.n207 a_n8300_8799.t144 464.166
R261 a_n8300_8799.n259 a_n8300_8799.t106 464.166
R262 a_n8300_8799.n258 a_n8300_8799.t103 464.166
R263 a_n8300_8799.n210 a_n8300_8799.t43 464.166
R264 a_n8300_8799.n252 a_n8300_8799.t111 464.166
R265 a_n8300_8799.n251 a_n8300_8799.t110 464.166
R266 a_n8300_8799.n213 a_n8300_8799.t45 464.166
R267 a_n8300_8799.n245 a_n8300_8799.t44 464.166
R268 a_n8300_8799.n244 a_n8300_8799.t132 464.166
R269 a_n8300_8799.n216 a_n8300_8799.t60 464.166
R270 a_n8300_8799.n238 a_n8300_8799.t49 464.166
R271 a_n8300_8799.n237 a_n8300_8799.t136 464.166
R272 a_n8300_8799.n219 a_n8300_8799.t88 464.166
R273 a_n8300_8799.n231 a_n8300_8799.t64 464.166
R274 a_n8300_8799.n230 a_n8300_8799.t156 464.166
R275 a_n8300_8799.n222 a_n8300_8799.t105 464.166
R276 a_n8300_8799.n224 a_n8300_8799.t67 464.166
R277 a_n8300_8799.n328 a_n8300_8799.t100 464.166
R278 a_n8300_8799.n327 a_n8300_8799.t76 464.166
R279 a_n8300_8799.n269 a_n8300_8799.t158 464.166
R280 a_n8300_8799.n321 a_n8300_8799.t121 464.166
R281 a_n8300_8799.n320 a_n8300_8799.t120 464.166
R282 a_n8300_8799.n272 a_n8300_8799.t54 464.166
R283 a_n8300_8799.n314 a_n8300_8799.t128 464.166
R284 a_n8300_8799.n313 a_n8300_8799.t127 464.166
R285 a_n8300_8799.n275 a_n8300_8799.t56 464.166
R286 a_n8300_8799.n307 a_n8300_8799.t55 464.166
R287 a_n8300_8799.n306 a_n8300_8799.t148 464.166
R288 a_n8300_8799.n278 a_n8300_8799.t73 464.166
R289 a_n8300_8799.n300 a_n8300_8799.t59 464.166
R290 a_n8300_8799.n299 a_n8300_8799.t150 464.166
R291 a_n8300_8799.n281 a_n8300_8799.t101 464.166
R292 a_n8300_8799.n293 a_n8300_8799.t77 464.166
R293 a_n8300_8799.n292 a_n8300_8799.t47 464.166
R294 a_n8300_8799.n284 a_n8300_8799.t122 464.166
R295 a_n8300_8799.n286 a_n8300_8799.t78 464.166
R296 a_n8300_8799.n391 a_n8300_8799.t131 464.166
R297 a_n8300_8799.n390 a_n8300_8799.t62 464.166
R298 a_n8300_8799.n332 a_n8300_8799.t109 464.166
R299 a_n8300_8799.n384 a_n8300_8799.t48 464.166
R300 a_n8300_8799.n383 a_n8300_8799.t68 464.166
R301 a_n8300_8799.n335 a_n8300_8799.t153 464.166
R302 a_n8300_8799.n377 a_n8300_8799.t119 464.166
R303 a_n8300_8799.n376 a_n8300_8799.t147 464.166
R304 a_n8300_8799.n338 a_n8300_8799.t99 464.166
R305 a_n8300_8799.n370 a_n8300_8799.t126 464.166
R306 a_n8300_8799.n369 a_n8300_8799.t58 464.166
R307 a_n8300_8799.n341 a_n8300_8799.t143 464.166
R308 a_n8300_8799.n363 a_n8300_8799.t82 464.166
R309 a_n8300_8799.n362 a_n8300_8799.t137 464.166
R310 a_n8300_8799.n344 a_n8300_8799.t66 464.166
R311 a_n8300_8799.n356 a_n8300_8799.t114 464.166
R312 a_n8300_8799.n355 a_n8300_8799.t53 464.166
R313 a_n8300_8799.n347 a_n8300_8799.t96 464.166
R314 a_n8300_8799.n349 a_n8300_8799.t75 464.166
R315 a_n8300_8799.n34 a_n8300_8799.t146 464.166
R316 a_n8300_8799.n36 a_n8300_8799.t69 464.166
R317 a_n8300_8799.n40 a_n8300_8799.t102 464.166
R318 a_n8300_8799.n41 a_n8300_8799.t139 464.166
R319 a_n8300_8799.n29 a_n8300_8799.t141 464.166
R320 a_n8300_8799.n47 a_n8300_8799.t87 464.166
R321 a_n8300_8799.n48 a_n8300_8799.t118 464.166
R322 a_n8300_8799.n52 a_n8300_8799.t138 464.166
R323 a_n8300_8799.n54 a_n8300_8799.t85 464.166
R324 a_n8300_8799.n25 a_n8300_8799.t86 464.166
R325 a_n8300_8799.n59 a_n8300_8799.t115 464.166
R326 a_n8300_8799.n23 a_n8300_8799.t71 464.166
R327 a_n8300_8799.n64 a_n8300_8799.t72 464.166
R328 a_n8300_8799.n66 a_n8300_8799.t112 464.166
R329 a_n8300_8799.n70 a_n8300_8799.t40 464.166
R330 a_n8300_8799.n71 a_n8300_8799.t70 464.166
R331 a_n8300_8799.n19 a_n8300_8799.t92 464.166
R332 a_n8300_8799.n77 a_n8300_8799.t140 464.166
R333 a_n8300_8799.n78 a_n8300_8799.t51 464.166
R334 a_n8300_8799.n96 a_n8300_8799.t159 464.166
R335 a_n8300_8799.n98 a_n8300_8799.t79 464.166
R336 a_n8300_8799.n102 a_n8300_8799.t116 464.166
R337 a_n8300_8799.n103 a_n8300_8799.t154 464.166
R338 a_n8300_8799.n91 a_n8300_8799.t157 464.166
R339 a_n8300_8799.n109 a_n8300_8799.t97 464.166
R340 a_n8300_8799.n110 a_n8300_8799.t135 464.166
R341 a_n8300_8799.n114 a_n8300_8799.t152 464.166
R342 a_n8300_8799.n116 a_n8300_8799.t93 464.166
R343 a_n8300_8799.n87 a_n8300_8799.t94 464.166
R344 a_n8300_8799.n121 a_n8300_8799.t133 464.166
R345 a_n8300_8799.n85 a_n8300_8799.t83 464.166
R346 a_n8300_8799.n126 a_n8300_8799.t84 464.166
R347 a_n8300_8799.n128 a_n8300_8799.t129 464.166
R348 a_n8300_8799.n132 a_n8300_8799.t50 464.166
R349 a_n8300_8799.n133 a_n8300_8799.t80 464.166
R350 a_n8300_8799.n81 a_n8300_8799.t104 464.166
R351 a_n8300_8799.n139 a_n8300_8799.t155 464.166
R352 a_n8300_8799.n140 a_n8300_8799.t63 464.166
R353 a_n8300_8799.n159 a_n8300_8799.t74 464.166
R354 a_n8300_8799.n161 a_n8300_8799.t95 464.166
R355 a_n8300_8799.n165 a_n8300_8799.t52 464.166
R356 a_n8300_8799.n166 a_n8300_8799.t113 464.166
R357 a_n8300_8799.n154 a_n8300_8799.t90 464.166
R358 a_n8300_8799.n172 a_n8300_8799.t134 464.166
R359 a_n8300_8799.n173 a_n8300_8799.t81 464.166
R360 a_n8300_8799.n177 a_n8300_8799.t142 464.166
R361 a_n8300_8799.n179 a_n8300_8799.t57 464.166
R362 a_n8300_8799.n150 a_n8300_8799.t41 464.166
R363 a_n8300_8799.n184 a_n8300_8799.t98 464.166
R364 a_n8300_8799.n148 a_n8300_8799.t145 464.166
R365 a_n8300_8799.n189 a_n8300_8799.t117 464.166
R366 a_n8300_8799.n191 a_n8300_8799.t151 464.166
R367 a_n8300_8799.n195 a_n8300_8799.t91 464.166
R368 a_n8300_8799.n196 a_n8300_8799.t46 464.166
R369 a_n8300_8799.n144 a_n8300_8799.t108 464.166
R370 a_n8300_8799.n202 a_n8300_8799.t61 464.166
R371 a_n8300_8799.n203 a_n8300_8799.t130 464.166
R372 a_n8300_8799.n226 a_n8300_8799.n225 161.3
R373 a_n8300_8799.n227 a_n8300_8799.n222 161.3
R374 a_n8300_8799.n229 a_n8300_8799.n228 161.3
R375 a_n8300_8799.n230 a_n8300_8799.n221 161.3
R376 a_n8300_8799.n231 a_n8300_8799.n220 161.3
R377 a_n8300_8799.n233 a_n8300_8799.n232 161.3
R378 a_n8300_8799.n234 a_n8300_8799.n219 161.3
R379 a_n8300_8799.n236 a_n8300_8799.n235 161.3
R380 a_n8300_8799.n237 a_n8300_8799.n218 161.3
R381 a_n8300_8799.n238 a_n8300_8799.n217 161.3
R382 a_n8300_8799.n240 a_n8300_8799.n239 161.3
R383 a_n8300_8799.n241 a_n8300_8799.n216 161.3
R384 a_n8300_8799.n243 a_n8300_8799.n242 161.3
R385 a_n8300_8799.n244 a_n8300_8799.n215 161.3
R386 a_n8300_8799.n245 a_n8300_8799.n214 161.3
R387 a_n8300_8799.n247 a_n8300_8799.n246 161.3
R388 a_n8300_8799.n248 a_n8300_8799.n213 161.3
R389 a_n8300_8799.n250 a_n8300_8799.n249 161.3
R390 a_n8300_8799.n251 a_n8300_8799.n212 161.3
R391 a_n8300_8799.n252 a_n8300_8799.n211 161.3
R392 a_n8300_8799.n254 a_n8300_8799.n253 161.3
R393 a_n8300_8799.n255 a_n8300_8799.n210 161.3
R394 a_n8300_8799.n257 a_n8300_8799.n256 161.3
R395 a_n8300_8799.n258 a_n8300_8799.n209 161.3
R396 a_n8300_8799.n259 a_n8300_8799.n208 161.3
R397 a_n8300_8799.n261 a_n8300_8799.n260 161.3
R398 a_n8300_8799.n262 a_n8300_8799.n207 161.3
R399 a_n8300_8799.n264 a_n8300_8799.n263 161.3
R400 a_n8300_8799.n265 a_n8300_8799.n206 161.3
R401 a_n8300_8799.n267 a_n8300_8799.n266 161.3
R402 a_n8300_8799.n288 a_n8300_8799.n287 161.3
R403 a_n8300_8799.n289 a_n8300_8799.n284 161.3
R404 a_n8300_8799.n291 a_n8300_8799.n290 161.3
R405 a_n8300_8799.n292 a_n8300_8799.n283 161.3
R406 a_n8300_8799.n293 a_n8300_8799.n282 161.3
R407 a_n8300_8799.n295 a_n8300_8799.n294 161.3
R408 a_n8300_8799.n296 a_n8300_8799.n281 161.3
R409 a_n8300_8799.n298 a_n8300_8799.n297 161.3
R410 a_n8300_8799.n299 a_n8300_8799.n280 161.3
R411 a_n8300_8799.n300 a_n8300_8799.n279 161.3
R412 a_n8300_8799.n302 a_n8300_8799.n301 161.3
R413 a_n8300_8799.n303 a_n8300_8799.n278 161.3
R414 a_n8300_8799.n305 a_n8300_8799.n304 161.3
R415 a_n8300_8799.n306 a_n8300_8799.n277 161.3
R416 a_n8300_8799.n307 a_n8300_8799.n276 161.3
R417 a_n8300_8799.n309 a_n8300_8799.n308 161.3
R418 a_n8300_8799.n310 a_n8300_8799.n275 161.3
R419 a_n8300_8799.n312 a_n8300_8799.n311 161.3
R420 a_n8300_8799.n313 a_n8300_8799.n274 161.3
R421 a_n8300_8799.n314 a_n8300_8799.n273 161.3
R422 a_n8300_8799.n316 a_n8300_8799.n315 161.3
R423 a_n8300_8799.n317 a_n8300_8799.n272 161.3
R424 a_n8300_8799.n319 a_n8300_8799.n318 161.3
R425 a_n8300_8799.n320 a_n8300_8799.n271 161.3
R426 a_n8300_8799.n321 a_n8300_8799.n270 161.3
R427 a_n8300_8799.n323 a_n8300_8799.n322 161.3
R428 a_n8300_8799.n324 a_n8300_8799.n269 161.3
R429 a_n8300_8799.n326 a_n8300_8799.n325 161.3
R430 a_n8300_8799.n327 a_n8300_8799.n268 161.3
R431 a_n8300_8799.n329 a_n8300_8799.n328 161.3
R432 a_n8300_8799.n351 a_n8300_8799.n350 161.3
R433 a_n8300_8799.n352 a_n8300_8799.n347 161.3
R434 a_n8300_8799.n354 a_n8300_8799.n353 161.3
R435 a_n8300_8799.n355 a_n8300_8799.n346 161.3
R436 a_n8300_8799.n356 a_n8300_8799.n345 161.3
R437 a_n8300_8799.n358 a_n8300_8799.n357 161.3
R438 a_n8300_8799.n359 a_n8300_8799.n344 161.3
R439 a_n8300_8799.n361 a_n8300_8799.n360 161.3
R440 a_n8300_8799.n362 a_n8300_8799.n343 161.3
R441 a_n8300_8799.n363 a_n8300_8799.n342 161.3
R442 a_n8300_8799.n365 a_n8300_8799.n364 161.3
R443 a_n8300_8799.n366 a_n8300_8799.n341 161.3
R444 a_n8300_8799.n368 a_n8300_8799.n367 161.3
R445 a_n8300_8799.n369 a_n8300_8799.n340 161.3
R446 a_n8300_8799.n370 a_n8300_8799.n339 161.3
R447 a_n8300_8799.n372 a_n8300_8799.n371 161.3
R448 a_n8300_8799.n373 a_n8300_8799.n338 161.3
R449 a_n8300_8799.n375 a_n8300_8799.n374 161.3
R450 a_n8300_8799.n376 a_n8300_8799.n337 161.3
R451 a_n8300_8799.n377 a_n8300_8799.n336 161.3
R452 a_n8300_8799.n379 a_n8300_8799.n378 161.3
R453 a_n8300_8799.n380 a_n8300_8799.n335 161.3
R454 a_n8300_8799.n382 a_n8300_8799.n381 161.3
R455 a_n8300_8799.n383 a_n8300_8799.n334 161.3
R456 a_n8300_8799.n384 a_n8300_8799.n333 161.3
R457 a_n8300_8799.n386 a_n8300_8799.n385 161.3
R458 a_n8300_8799.n387 a_n8300_8799.n332 161.3
R459 a_n8300_8799.n389 a_n8300_8799.n388 161.3
R460 a_n8300_8799.n390 a_n8300_8799.n331 161.3
R461 a_n8300_8799.n392 a_n8300_8799.n391 161.3
R462 a_n8300_8799.n79 a_n8300_8799.n78 161.3
R463 a_n8300_8799.n77 a_n8300_8799.n18 161.3
R464 a_n8300_8799.n76 a_n8300_8799.n75 161.3
R465 a_n8300_8799.n74 a_n8300_8799.n19 161.3
R466 a_n8300_8799.n73 a_n8300_8799.n72 161.3
R467 a_n8300_8799.n71 a_n8300_8799.n20 161.3
R468 a_n8300_8799.n70 a_n8300_8799.n69 161.3
R469 a_n8300_8799.n68 a_n8300_8799.n21 161.3
R470 a_n8300_8799.n67 a_n8300_8799.n66 161.3
R471 a_n8300_8799.n65 a_n8300_8799.n22 161.3
R472 a_n8300_8799.n64 a_n8300_8799.n63 161.3
R473 a_n8300_8799.n62 a_n8300_8799.n23 161.3
R474 a_n8300_8799.n61 a_n8300_8799.n60 161.3
R475 a_n8300_8799.n59 a_n8300_8799.n24 161.3
R476 a_n8300_8799.n58 a_n8300_8799.n57 161.3
R477 a_n8300_8799.n56 a_n8300_8799.n25 161.3
R478 a_n8300_8799.n55 a_n8300_8799.n54 161.3
R479 a_n8300_8799.n53 a_n8300_8799.n26 161.3
R480 a_n8300_8799.n52 a_n8300_8799.n51 161.3
R481 a_n8300_8799.n50 a_n8300_8799.n27 161.3
R482 a_n8300_8799.n49 a_n8300_8799.n48 161.3
R483 a_n8300_8799.n47 a_n8300_8799.n28 161.3
R484 a_n8300_8799.n46 a_n8300_8799.n45 161.3
R485 a_n8300_8799.n44 a_n8300_8799.n29 161.3
R486 a_n8300_8799.n43 a_n8300_8799.n42 161.3
R487 a_n8300_8799.n41 a_n8300_8799.n30 161.3
R488 a_n8300_8799.n40 a_n8300_8799.n39 161.3
R489 a_n8300_8799.n38 a_n8300_8799.n31 161.3
R490 a_n8300_8799.n37 a_n8300_8799.n36 161.3
R491 a_n8300_8799.n35 a_n8300_8799.n32 161.3
R492 a_n8300_8799.n141 a_n8300_8799.n140 161.3
R493 a_n8300_8799.n139 a_n8300_8799.n80 161.3
R494 a_n8300_8799.n138 a_n8300_8799.n137 161.3
R495 a_n8300_8799.n136 a_n8300_8799.n81 161.3
R496 a_n8300_8799.n135 a_n8300_8799.n134 161.3
R497 a_n8300_8799.n133 a_n8300_8799.n82 161.3
R498 a_n8300_8799.n132 a_n8300_8799.n131 161.3
R499 a_n8300_8799.n130 a_n8300_8799.n83 161.3
R500 a_n8300_8799.n129 a_n8300_8799.n128 161.3
R501 a_n8300_8799.n127 a_n8300_8799.n84 161.3
R502 a_n8300_8799.n126 a_n8300_8799.n125 161.3
R503 a_n8300_8799.n124 a_n8300_8799.n85 161.3
R504 a_n8300_8799.n123 a_n8300_8799.n122 161.3
R505 a_n8300_8799.n121 a_n8300_8799.n86 161.3
R506 a_n8300_8799.n120 a_n8300_8799.n119 161.3
R507 a_n8300_8799.n118 a_n8300_8799.n87 161.3
R508 a_n8300_8799.n117 a_n8300_8799.n116 161.3
R509 a_n8300_8799.n115 a_n8300_8799.n88 161.3
R510 a_n8300_8799.n114 a_n8300_8799.n113 161.3
R511 a_n8300_8799.n112 a_n8300_8799.n89 161.3
R512 a_n8300_8799.n111 a_n8300_8799.n110 161.3
R513 a_n8300_8799.n109 a_n8300_8799.n90 161.3
R514 a_n8300_8799.n108 a_n8300_8799.n107 161.3
R515 a_n8300_8799.n106 a_n8300_8799.n91 161.3
R516 a_n8300_8799.n105 a_n8300_8799.n104 161.3
R517 a_n8300_8799.n103 a_n8300_8799.n92 161.3
R518 a_n8300_8799.n102 a_n8300_8799.n101 161.3
R519 a_n8300_8799.n100 a_n8300_8799.n93 161.3
R520 a_n8300_8799.n99 a_n8300_8799.n98 161.3
R521 a_n8300_8799.n97 a_n8300_8799.n94 161.3
R522 a_n8300_8799.n204 a_n8300_8799.n203 161.3
R523 a_n8300_8799.n202 a_n8300_8799.n143 161.3
R524 a_n8300_8799.n201 a_n8300_8799.n200 161.3
R525 a_n8300_8799.n199 a_n8300_8799.n144 161.3
R526 a_n8300_8799.n198 a_n8300_8799.n197 161.3
R527 a_n8300_8799.n196 a_n8300_8799.n145 161.3
R528 a_n8300_8799.n195 a_n8300_8799.n194 161.3
R529 a_n8300_8799.n193 a_n8300_8799.n146 161.3
R530 a_n8300_8799.n192 a_n8300_8799.n191 161.3
R531 a_n8300_8799.n190 a_n8300_8799.n147 161.3
R532 a_n8300_8799.n189 a_n8300_8799.n188 161.3
R533 a_n8300_8799.n187 a_n8300_8799.n148 161.3
R534 a_n8300_8799.n186 a_n8300_8799.n185 161.3
R535 a_n8300_8799.n184 a_n8300_8799.n149 161.3
R536 a_n8300_8799.n183 a_n8300_8799.n182 161.3
R537 a_n8300_8799.n181 a_n8300_8799.n150 161.3
R538 a_n8300_8799.n180 a_n8300_8799.n179 161.3
R539 a_n8300_8799.n178 a_n8300_8799.n151 161.3
R540 a_n8300_8799.n177 a_n8300_8799.n176 161.3
R541 a_n8300_8799.n175 a_n8300_8799.n152 161.3
R542 a_n8300_8799.n174 a_n8300_8799.n173 161.3
R543 a_n8300_8799.n172 a_n8300_8799.n153 161.3
R544 a_n8300_8799.n171 a_n8300_8799.n170 161.3
R545 a_n8300_8799.n169 a_n8300_8799.n154 161.3
R546 a_n8300_8799.n168 a_n8300_8799.n167 161.3
R547 a_n8300_8799.n166 a_n8300_8799.n155 161.3
R548 a_n8300_8799.n165 a_n8300_8799.n164 161.3
R549 a_n8300_8799.n163 a_n8300_8799.n156 161.3
R550 a_n8300_8799.n162 a_n8300_8799.n161 161.3
R551 a_n8300_8799.n160 a_n8300_8799.n157 161.3
R552 a_n8300_8799.n12 a_n8300_8799.n10 98.9633
R553 a_n8300_8799.n5 a_n8300_8799.n3 98.9631
R554 a_n8300_8799.n16 a_n8300_8799.n15 98.6055
R555 a_n8300_8799.n14 a_n8300_8799.n13 98.6055
R556 a_n8300_8799.n12 a_n8300_8799.n11 98.6055
R557 a_n8300_8799.n5 a_n8300_8799.n4 98.6055
R558 a_n8300_8799.n7 a_n8300_8799.n6 98.6055
R559 a_n8300_8799.n9 a_n8300_8799.n8 98.6055
R560 a_n8300_8799.n398 a_n8300_8799.n396 81.3764
R561 a_n8300_8799.n410 a_n8300_8799.n408 81.3764
R562 a_n8300_8799.n2 a_n8300_8799.n0 81.3764
R563 a_n8300_8799.n415 a_n8300_8799.n414 80.9326
R564 a_n8300_8799.n407 a_n8300_8799.n406 80.9324
R565 a_n8300_8799.n405 a_n8300_8799.n404 80.9324
R566 a_n8300_8799.n403 a_n8300_8799.n402 80.9324
R567 a_n8300_8799.n400 a_n8300_8799.n399 80.9324
R568 a_n8300_8799.n398 a_n8300_8799.n397 80.9324
R569 a_n8300_8799.n410 a_n8300_8799.n409 80.9324
R570 a_n8300_8799.n412 a_n8300_8799.n411 80.9324
R571 a_n8300_8799.n2 a_n8300_8799.n1 80.9324
R572 a_n8300_8799.n226 a_n8300_8799.n223 70.4033
R573 a_n8300_8799.n288 a_n8300_8799.n285 70.4033
R574 a_n8300_8799.n351 a_n8300_8799.n348 70.4033
R575 a_n8300_8799.n33 a_n8300_8799.n32 70.4033
R576 a_n8300_8799.n95 a_n8300_8799.n94 70.4033
R577 a_n8300_8799.n158 a_n8300_8799.n157 70.4033
R578 a_n8300_8799.n266 a_n8300_8799.n265 48.2005
R579 a_n8300_8799.n259 a_n8300_8799.n258 48.2005
R580 a_n8300_8799.n252 a_n8300_8799.n251 48.2005
R581 a_n8300_8799.n245 a_n8300_8799.n244 48.2005
R582 a_n8300_8799.n238 a_n8300_8799.n237 48.2005
R583 a_n8300_8799.n231 a_n8300_8799.n230 48.2005
R584 a_n8300_8799.n328 a_n8300_8799.n327 48.2005
R585 a_n8300_8799.n321 a_n8300_8799.n320 48.2005
R586 a_n8300_8799.n314 a_n8300_8799.n313 48.2005
R587 a_n8300_8799.n307 a_n8300_8799.n306 48.2005
R588 a_n8300_8799.n300 a_n8300_8799.n299 48.2005
R589 a_n8300_8799.n293 a_n8300_8799.n292 48.2005
R590 a_n8300_8799.n391 a_n8300_8799.n390 48.2005
R591 a_n8300_8799.n384 a_n8300_8799.n383 48.2005
R592 a_n8300_8799.n377 a_n8300_8799.n376 48.2005
R593 a_n8300_8799.n370 a_n8300_8799.n369 48.2005
R594 a_n8300_8799.n363 a_n8300_8799.n362 48.2005
R595 a_n8300_8799.n356 a_n8300_8799.n355 48.2005
R596 a_n8300_8799.n41 a_n8300_8799.n40 48.2005
R597 a_n8300_8799.n48 a_n8300_8799.n47 48.2005
R598 a_n8300_8799.n54 a_n8300_8799.n25 48.2005
R599 a_n8300_8799.n64 a_n8300_8799.n23 48.2005
R600 a_n8300_8799.n71 a_n8300_8799.n70 48.2005
R601 a_n8300_8799.n78 a_n8300_8799.n77 48.2005
R602 a_n8300_8799.n103 a_n8300_8799.n102 48.2005
R603 a_n8300_8799.n110 a_n8300_8799.n109 48.2005
R604 a_n8300_8799.n116 a_n8300_8799.n87 48.2005
R605 a_n8300_8799.n126 a_n8300_8799.n85 48.2005
R606 a_n8300_8799.n133 a_n8300_8799.n132 48.2005
R607 a_n8300_8799.n140 a_n8300_8799.n139 48.2005
R608 a_n8300_8799.n166 a_n8300_8799.n165 48.2005
R609 a_n8300_8799.n173 a_n8300_8799.n172 48.2005
R610 a_n8300_8799.n179 a_n8300_8799.n150 48.2005
R611 a_n8300_8799.n189 a_n8300_8799.n148 48.2005
R612 a_n8300_8799.n196 a_n8300_8799.n195 48.2005
R613 a_n8300_8799.n203 a_n8300_8799.n202 48.2005
R614 a_n8300_8799.n264 a_n8300_8799.n207 40.1672
R615 a_n8300_8799.n225 a_n8300_8799.n222 40.1672
R616 a_n8300_8799.n326 a_n8300_8799.n269 40.1672
R617 a_n8300_8799.n287 a_n8300_8799.n284 40.1672
R618 a_n8300_8799.n389 a_n8300_8799.n332 40.1672
R619 a_n8300_8799.n350 a_n8300_8799.n347 40.1672
R620 a_n8300_8799.n36 a_n8300_8799.n35 40.1672
R621 a_n8300_8799.n76 a_n8300_8799.n19 40.1672
R622 a_n8300_8799.n98 a_n8300_8799.n97 40.1672
R623 a_n8300_8799.n138 a_n8300_8799.n81 40.1672
R624 a_n8300_8799.n161 a_n8300_8799.n160 40.1672
R625 a_n8300_8799.n201 a_n8300_8799.n144 40.1672
R626 a_n8300_8799.n257 a_n8300_8799.n210 38.7066
R627 a_n8300_8799.n232 a_n8300_8799.n219 38.7066
R628 a_n8300_8799.n319 a_n8300_8799.n272 38.7066
R629 a_n8300_8799.n294 a_n8300_8799.n281 38.7066
R630 a_n8300_8799.n382 a_n8300_8799.n335 38.7066
R631 a_n8300_8799.n357 a_n8300_8799.n344 38.7066
R632 a_n8300_8799.n42 a_n8300_8799.n29 38.7066
R633 a_n8300_8799.n66 a_n8300_8799.n21 38.7066
R634 a_n8300_8799.n104 a_n8300_8799.n91 38.7066
R635 a_n8300_8799.n128 a_n8300_8799.n83 38.7066
R636 a_n8300_8799.n167 a_n8300_8799.n154 38.7066
R637 a_n8300_8799.n191 a_n8300_8799.n146 38.7066
R638 a_n8300_8799.n250 a_n8300_8799.n213 37.246
R639 a_n8300_8799.n239 a_n8300_8799.n216 37.246
R640 a_n8300_8799.n312 a_n8300_8799.n275 37.246
R641 a_n8300_8799.n301 a_n8300_8799.n278 37.246
R642 a_n8300_8799.n375 a_n8300_8799.n338 37.246
R643 a_n8300_8799.n364 a_n8300_8799.n341 37.246
R644 a_n8300_8799.n52 a_n8300_8799.n27 37.246
R645 a_n8300_8799.n60 a_n8300_8799.n59 37.246
R646 a_n8300_8799.n114 a_n8300_8799.n89 37.246
R647 a_n8300_8799.n122 a_n8300_8799.n121 37.246
R648 a_n8300_8799.n177 a_n8300_8799.n152 37.246
R649 a_n8300_8799.n185 a_n8300_8799.n184 37.246
R650 a_n8300_8799.n246 a_n8300_8799.n213 35.7853
R651 a_n8300_8799.n243 a_n8300_8799.n216 35.7853
R652 a_n8300_8799.n308 a_n8300_8799.n275 35.7853
R653 a_n8300_8799.n305 a_n8300_8799.n278 35.7853
R654 a_n8300_8799.n371 a_n8300_8799.n338 35.7853
R655 a_n8300_8799.n368 a_n8300_8799.n341 35.7853
R656 a_n8300_8799.n53 a_n8300_8799.n52 35.7853
R657 a_n8300_8799.n59 a_n8300_8799.n58 35.7853
R658 a_n8300_8799.n115 a_n8300_8799.n114 35.7853
R659 a_n8300_8799.n121 a_n8300_8799.n120 35.7853
R660 a_n8300_8799.n178 a_n8300_8799.n177 35.7853
R661 a_n8300_8799.n184 a_n8300_8799.n183 35.7853
R662 a_n8300_8799.n253 a_n8300_8799.n210 34.3247
R663 a_n8300_8799.n236 a_n8300_8799.n219 34.3247
R664 a_n8300_8799.n315 a_n8300_8799.n272 34.3247
R665 a_n8300_8799.n298 a_n8300_8799.n281 34.3247
R666 a_n8300_8799.n378 a_n8300_8799.n335 34.3247
R667 a_n8300_8799.n361 a_n8300_8799.n344 34.3247
R668 a_n8300_8799.n46 a_n8300_8799.n29 34.3247
R669 a_n8300_8799.n66 a_n8300_8799.n65 34.3247
R670 a_n8300_8799.n108 a_n8300_8799.n91 34.3247
R671 a_n8300_8799.n128 a_n8300_8799.n127 34.3247
R672 a_n8300_8799.n171 a_n8300_8799.n154 34.3247
R673 a_n8300_8799.n191 a_n8300_8799.n190 34.3247
R674 a_n8300_8799.n413 a_n8300_8799.n407 33.4185
R675 a_n8300_8799.n260 a_n8300_8799.n207 32.8641
R676 a_n8300_8799.n229 a_n8300_8799.n222 32.8641
R677 a_n8300_8799.n322 a_n8300_8799.n269 32.8641
R678 a_n8300_8799.n291 a_n8300_8799.n284 32.8641
R679 a_n8300_8799.n385 a_n8300_8799.n332 32.8641
R680 a_n8300_8799.n354 a_n8300_8799.n347 32.8641
R681 a_n8300_8799.n36 a_n8300_8799.n31 32.8641
R682 a_n8300_8799.n72 a_n8300_8799.n19 32.8641
R683 a_n8300_8799.n98 a_n8300_8799.n93 32.8641
R684 a_n8300_8799.n134 a_n8300_8799.n81 32.8641
R685 a_n8300_8799.n161 a_n8300_8799.n156 32.8641
R686 a_n8300_8799.n197 a_n8300_8799.n144 32.8641
R687 a_n8300_8799.n17 a_n8300_8799.n9 32.0088
R688 a_n8300_8799.n224 a_n8300_8799.n223 20.9576
R689 a_n8300_8799.n286 a_n8300_8799.n285 20.9576
R690 a_n8300_8799.n349 a_n8300_8799.n348 20.9576
R691 a_n8300_8799.n34 a_n8300_8799.n33 20.9576
R692 a_n8300_8799.n96 a_n8300_8799.n95 20.9576
R693 a_n8300_8799.n159 a_n8300_8799.n158 20.9576
R694 a_n8300_8799.n17 a_n8300_8799.n16 18.5874
R695 a_n8300_8799.n260 a_n8300_8799.n259 15.3369
R696 a_n8300_8799.n230 a_n8300_8799.n229 15.3369
R697 a_n8300_8799.n322 a_n8300_8799.n321 15.3369
R698 a_n8300_8799.n292 a_n8300_8799.n291 15.3369
R699 a_n8300_8799.n385 a_n8300_8799.n384 15.3369
R700 a_n8300_8799.n355 a_n8300_8799.n354 15.3369
R701 a_n8300_8799.n40 a_n8300_8799.n31 15.3369
R702 a_n8300_8799.n72 a_n8300_8799.n71 15.3369
R703 a_n8300_8799.n102 a_n8300_8799.n93 15.3369
R704 a_n8300_8799.n134 a_n8300_8799.n133 15.3369
R705 a_n8300_8799.n165 a_n8300_8799.n156 15.3369
R706 a_n8300_8799.n197 a_n8300_8799.n196 15.3369
R707 a_n8300_8799.n253 a_n8300_8799.n252 13.8763
R708 a_n8300_8799.n237 a_n8300_8799.n236 13.8763
R709 a_n8300_8799.n315 a_n8300_8799.n314 13.8763
R710 a_n8300_8799.n299 a_n8300_8799.n298 13.8763
R711 a_n8300_8799.n378 a_n8300_8799.n377 13.8763
R712 a_n8300_8799.n362 a_n8300_8799.n361 13.8763
R713 a_n8300_8799.n47 a_n8300_8799.n46 13.8763
R714 a_n8300_8799.n65 a_n8300_8799.n64 13.8763
R715 a_n8300_8799.n109 a_n8300_8799.n108 13.8763
R716 a_n8300_8799.n127 a_n8300_8799.n126 13.8763
R717 a_n8300_8799.n172 a_n8300_8799.n171 13.8763
R718 a_n8300_8799.n190 a_n8300_8799.n189 13.8763
R719 a_n8300_8799.n246 a_n8300_8799.n245 12.4157
R720 a_n8300_8799.n244 a_n8300_8799.n243 12.4157
R721 a_n8300_8799.n308 a_n8300_8799.n307 12.4157
R722 a_n8300_8799.n306 a_n8300_8799.n305 12.4157
R723 a_n8300_8799.n371 a_n8300_8799.n370 12.4157
R724 a_n8300_8799.n369 a_n8300_8799.n368 12.4157
R725 a_n8300_8799.n54 a_n8300_8799.n53 12.4157
R726 a_n8300_8799.n58 a_n8300_8799.n25 12.4157
R727 a_n8300_8799.n116 a_n8300_8799.n115 12.4157
R728 a_n8300_8799.n120 a_n8300_8799.n87 12.4157
R729 a_n8300_8799.n179 a_n8300_8799.n178 12.4157
R730 a_n8300_8799.n183 a_n8300_8799.n150 12.4157
R731 a_n8300_8799.n401 a_n8300_8799.n395 12.3339
R732 a_n8300_8799.n395 a_n8300_8799.n17 11.4887
R733 a_n8300_8799.n251 a_n8300_8799.n250 10.955
R734 a_n8300_8799.n239 a_n8300_8799.n238 10.955
R735 a_n8300_8799.n313 a_n8300_8799.n312 10.955
R736 a_n8300_8799.n301 a_n8300_8799.n300 10.955
R737 a_n8300_8799.n376 a_n8300_8799.n375 10.955
R738 a_n8300_8799.n364 a_n8300_8799.n363 10.955
R739 a_n8300_8799.n48 a_n8300_8799.n27 10.955
R740 a_n8300_8799.n60 a_n8300_8799.n23 10.955
R741 a_n8300_8799.n110 a_n8300_8799.n89 10.955
R742 a_n8300_8799.n122 a_n8300_8799.n85 10.955
R743 a_n8300_8799.n173 a_n8300_8799.n152 10.955
R744 a_n8300_8799.n185 a_n8300_8799.n148 10.955
R745 a_n8300_8799.n258 a_n8300_8799.n257 9.49444
R746 a_n8300_8799.n232 a_n8300_8799.n231 9.49444
R747 a_n8300_8799.n320 a_n8300_8799.n319 9.49444
R748 a_n8300_8799.n294 a_n8300_8799.n293 9.49444
R749 a_n8300_8799.n383 a_n8300_8799.n382 9.49444
R750 a_n8300_8799.n357 a_n8300_8799.n356 9.49444
R751 a_n8300_8799.n42 a_n8300_8799.n41 9.49444
R752 a_n8300_8799.n70 a_n8300_8799.n21 9.49444
R753 a_n8300_8799.n104 a_n8300_8799.n103 9.49444
R754 a_n8300_8799.n132 a_n8300_8799.n83 9.49444
R755 a_n8300_8799.n167 a_n8300_8799.n166 9.49444
R756 a_n8300_8799.n195 a_n8300_8799.n146 9.49444
R757 a_n8300_8799.n330 a_n8300_8799.n267 9.04406
R758 a_n8300_8799.n142 a_n8300_8799.n79 9.04406
R759 a_n8300_8799.n265 a_n8300_8799.n264 8.03383
R760 a_n8300_8799.n225 a_n8300_8799.n224 8.03383
R761 a_n8300_8799.n327 a_n8300_8799.n326 8.03383
R762 a_n8300_8799.n287 a_n8300_8799.n286 8.03383
R763 a_n8300_8799.n390 a_n8300_8799.n389 8.03383
R764 a_n8300_8799.n350 a_n8300_8799.n349 8.03383
R765 a_n8300_8799.n35 a_n8300_8799.n34 8.03383
R766 a_n8300_8799.n77 a_n8300_8799.n76 8.03383
R767 a_n8300_8799.n97 a_n8300_8799.n96 8.03383
R768 a_n8300_8799.n139 a_n8300_8799.n138 8.03383
R769 a_n8300_8799.n160 a_n8300_8799.n159 8.03383
R770 a_n8300_8799.n202 a_n8300_8799.n201 8.03383
R771 a_n8300_8799.n394 a_n8300_8799.n205 7.00615
R772 a_n8300_8799.n394 a_n8300_8799.n393 6.58471
R773 a_n8300_8799.n330 a_n8300_8799.n329 4.93611
R774 a_n8300_8799.n393 a_n8300_8799.n392 4.93611
R775 a_n8300_8799.n142 a_n8300_8799.n141 4.93611
R776 a_n8300_8799.n205 a_n8300_8799.n204 4.93611
R777 a_n8300_8799.n393 a_n8300_8799.n330 4.10845
R778 a_n8300_8799.n205 a_n8300_8799.n142 4.10845
R779 a_n8300_8799.n15 a_n8300_8799.t38 3.61217
R780 a_n8300_8799.n15 a_n8300_8799.t3 3.61217
R781 a_n8300_8799.n13 a_n8300_8799.t1 3.61217
R782 a_n8300_8799.n13 a_n8300_8799.t13 3.61217
R783 a_n8300_8799.n11 a_n8300_8799.t9 3.61217
R784 a_n8300_8799.n11 a_n8300_8799.t11 3.61217
R785 a_n8300_8799.n10 a_n8300_8799.t39 3.61217
R786 a_n8300_8799.n10 a_n8300_8799.t6 3.61217
R787 a_n8300_8799.n3 a_n8300_8799.t0 3.61217
R788 a_n8300_8799.n3 a_n8300_8799.t4 3.61217
R789 a_n8300_8799.n4 a_n8300_8799.t2 3.61217
R790 a_n8300_8799.n4 a_n8300_8799.t5 3.61217
R791 a_n8300_8799.n6 a_n8300_8799.t7 3.61217
R792 a_n8300_8799.n6 a_n8300_8799.t8 3.61217
R793 a_n8300_8799.n8 a_n8300_8799.t12 3.61217
R794 a_n8300_8799.n8 a_n8300_8799.t10 3.61217
R795 a_n8300_8799.n395 a_n8300_8799.n394 3.4105
R796 a_n8300_8799.n408 a_n8300_8799.t29 2.82907
R797 a_n8300_8799.n408 a_n8300_8799.t27 2.82907
R798 a_n8300_8799.n409 a_n8300_8799.t18 2.82907
R799 a_n8300_8799.n409 a_n8300_8799.t24 2.82907
R800 a_n8300_8799.n411 a_n8300_8799.t36 2.82907
R801 a_n8300_8799.n411 a_n8300_8799.t19 2.82907
R802 a_n8300_8799.n1 a_n8300_8799.t26 2.82907
R803 a_n8300_8799.n1 a_n8300_8799.t25 2.82907
R804 a_n8300_8799.n0 a_n8300_8799.t21 2.82907
R805 a_n8300_8799.n0 a_n8300_8799.t20 2.82907
R806 a_n8300_8799.n406 a_n8300_8799.t32 2.82907
R807 a_n8300_8799.n406 a_n8300_8799.t34 2.82907
R808 a_n8300_8799.n404 a_n8300_8799.t30 2.82907
R809 a_n8300_8799.n404 a_n8300_8799.t14 2.82907
R810 a_n8300_8799.n402 a_n8300_8799.t35 2.82907
R811 a_n8300_8799.n402 a_n8300_8799.t28 2.82907
R812 a_n8300_8799.n399 a_n8300_8799.t15 2.82907
R813 a_n8300_8799.n399 a_n8300_8799.t33 2.82907
R814 a_n8300_8799.n397 a_n8300_8799.t16 2.82907
R815 a_n8300_8799.n397 a_n8300_8799.t17 2.82907
R816 a_n8300_8799.n396 a_n8300_8799.t22 2.82907
R817 a_n8300_8799.n396 a_n8300_8799.t23 2.82907
R818 a_n8300_8799.n415 a_n8300_8799.t31 2.82907
R819 a_n8300_8799.t37 a_n8300_8799.n415 2.82907
R820 a_n8300_8799.n400 a_n8300_8799.n398 0.444466
R821 a_n8300_8799.n405 a_n8300_8799.n403 0.444466
R822 a_n8300_8799.n407 a_n8300_8799.n405 0.444466
R823 a_n8300_8799.n414 a_n8300_8799.n2 0.444466
R824 a_n8300_8799.n412 a_n8300_8799.n410 0.444466
R825 a_n8300_8799.n14 a_n8300_8799.n12 0.358259
R826 a_n8300_8799.n16 a_n8300_8799.n14 0.358259
R827 a_n8300_8799.n9 a_n8300_8799.n7 0.358259
R828 a_n8300_8799.n7 a_n8300_8799.n5 0.358259
R829 a_n8300_8799.n401 a_n8300_8799.n400 0.222483
R830 a_n8300_8799.n403 a_n8300_8799.n401 0.222483
R831 a_n8300_8799.n414 a_n8300_8799.n413 0.222483
R832 a_n8300_8799.n413 a_n8300_8799.n412 0.222483
R833 a_n8300_8799.n267 a_n8300_8799.n206 0.189894
R834 a_n8300_8799.n263 a_n8300_8799.n206 0.189894
R835 a_n8300_8799.n263 a_n8300_8799.n262 0.189894
R836 a_n8300_8799.n262 a_n8300_8799.n261 0.189894
R837 a_n8300_8799.n261 a_n8300_8799.n208 0.189894
R838 a_n8300_8799.n209 a_n8300_8799.n208 0.189894
R839 a_n8300_8799.n256 a_n8300_8799.n209 0.189894
R840 a_n8300_8799.n256 a_n8300_8799.n255 0.189894
R841 a_n8300_8799.n255 a_n8300_8799.n254 0.189894
R842 a_n8300_8799.n254 a_n8300_8799.n211 0.189894
R843 a_n8300_8799.n212 a_n8300_8799.n211 0.189894
R844 a_n8300_8799.n249 a_n8300_8799.n212 0.189894
R845 a_n8300_8799.n249 a_n8300_8799.n248 0.189894
R846 a_n8300_8799.n248 a_n8300_8799.n247 0.189894
R847 a_n8300_8799.n247 a_n8300_8799.n214 0.189894
R848 a_n8300_8799.n215 a_n8300_8799.n214 0.189894
R849 a_n8300_8799.n242 a_n8300_8799.n215 0.189894
R850 a_n8300_8799.n242 a_n8300_8799.n241 0.189894
R851 a_n8300_8799.n241 a_n8300_8799.n240 0.189894
R852 a_n8300_8799.n240 a_n8300_8799.n217 0.189894
R853 a_n8300_8799.n218 a_n8300_8799.n217 0.189894
R854 a_n8300_8799.n235 a_n8300_8799.n218 0.189894
R855 a_n8300_8799.n235 a_n8300_8799.n234 0.189894
R856 a_n8300_8799.n234 a_n8300_8799.n233 0.189894
R857 a_n8300_8799.n233 a_n8300_8799.n220 0.189894
R858 a_n8300_8799.n221 a_n8300_8799.n220 0.189894
R859 a_n8300_8799.n228 a_n8300_8799.n221 0.189894
R860 a_n8300_8799.n228 a_n8300_8799.n227 0.189894
R861 a_n8300_8799.n227 a_n8300_8799.n226 0.189894
R862 a_n8300_8799.n329 a_n8300_8799.n268 0.189894
R863 a_n8300_8799.n325 a_n8300_8799.n268 0.189894
R864 a_n8300_8799.n325 a_n8300_8799.n324 0.189894
R865 a_n8300_8799.n324 a_n8300_8799.n323 0.189894
R866 a_n8300_8799.n323 a_n8300_8799.n270 0.189894
R867 a_n8300_8799.n271 a_n8300_8799.n270 0.189894
R868 a_n8300_8799.n318 a_n8300_8799.n271 0.189894
R869 a_n8300_8799.n318 a_n8300_8799.n317 0.189894
R870 a_n8300_8799.n317 a_n8300_8799.n316 0.189894
R871 a_n8300_8799.n316 a_n8300_8799.n273 0.189894
R872 a_n8300_8799.n274 a_n8300_8799.n273 0.189894
R873 a_n8300_8799.n311 a_n8300_8799.n274 0.189894
R874 a_n8300_8799.n311 a_n8300_8799.n310 0.189894
R875 a_n8300_8799.n310 a_n8300_8799.n309 0.189894
R876 a_n8300_8799.n309 a_n8300_8799.n276 0.189894
R877 a_n8300_8799.n277 a_n8300_8799.n276 0.189894
R878 a_n8300_8799.n304 a_n8300_8799.n277 0.189894
R879 a_n8300_8799.n304 a_n8300_8799.n303 0.189894
R880 a_n8300_8799.n303 a_n8300_8799.n302 0.189894
R881 a_n8300_8799.n302 a_n8300_8799.n279 0.189894
R882 a_n8300_8799.n280 a_n8300_8799.n279 0.189894
R883 a_n8300_8799.n297 a_n8300_8799.n280 0.189894
R884 a_n8300_8799.n297 a_n8300_8799.n296 0.189894
R885 a_n8300_8799.n296 a_n8300_8799.n295 0.189894
R886 a_n8300_8799.n295 a_n8300_8799.n282 0.189894
R887 a_n8300_8799.n283 a_n8300_8799.n282 0.189894
R888 a_n8300_8799.n290 a_n8300_8799.n283 0.189894
R889 a_n8300_8799.n290 a_n8300_8799.n289 0.189894
R890 a_n8300_8799.n289 a_n8300_8799.n288 0.189894
R891 a_n8300_8799.n392 a_n8300_8799.n331 0.189894
R892 a_n8300_8799.n388 a_n8300_8799.n331 0.189894
R893 a_n8300_8799.n388 a_n8300_8799.n387 0.189894
R894 a_n8300_8799.n387 a_n8300_8799.n386 0.189894
R895 a_n8300_8799.n386 a_n8300_8799.n333 0.189894
R896 a_n8300_8799.n334 a_n8300_8799.n333 0.189894
R897 a_n8300_8799.n381 a_n8300_8799.n334 0.189894
R898 a_n8300_8799.n381 a_n8300_8799.n380 0.189894
R899 a_n8300_8799.n380 a_n8300_8799.n379 0.189894
R900 a_n8300_8799.n379 a_n8300_8799.n336 0.189894
R901 a_n8300_8799.n337 a_n8300_8799.n336 0.189894
R902 a_n8300_8799.n374 a_n8300_8799.n337 0.189894
R903 a_n8300_8799.n374 a_n8300_8799.n373 0.189894
R904 a_n8300_8799.n373 a_n8300_8799.n372 0.189894
R905 a_n8300_8799.n372 a_n8300_8799.n339 0.189894
R906 a_n8300_8799.n340 a_n8300_8799.n339 0.189894
R907 a_n8300_8799.n367 a_n8300_8799.n340 0.189894
R908 a_n8300_8799.n367 a_n8300_8799.n366 0.189894
R909 a_n8300_8799.n366 a_n8300_8799.n365 0.189894
R910 a_n8300_8799.n365 a_n8300_8799.n342 0.189894
R911 a_n8300_8799.n343 a_n8300_8799.n342 0.189894
R912 a_n8300_8799.n360 a_n8300_8799.n343 0.189894
R913 a_n8300_8799.n360 a_n8300_8799.n359 0.189894
R914 a_n8300_8799.n359 a_n8300_8799.n358 0.189894
R915 a_n8300_8799.n358 a_n8300_8799.n345 0.189894
R916 a_n8300_8799.n346 a_n8300_8799.n345 0.189894
R917 a_n8300_8799.n353 a_n8300_8799.n346 0.189894
R918 a_n8300_8799.n353 a_n8300_8799.n352 0.189894
R919 a_n8300_8799.n352 a_n8300_8799.n351 0.189894
R920 a_n8300_8799.n37 a_n8300_8799.n32 0.189894
R921 a_n8300_8799.n38 a_n8300_8799.n37 0.189894
R922 a_n8300_8799.n39 a_n8300_8799.n38 0.189894
R923 a_n8300_8799.n39 a_n8300_8799.n30 0.189894
R924 a_n8300_8799.n43 a_n8300_8799.n30 0.189894
R925 a_n8300_8799.n44 a_n8300_8799.n43 0.189894
R926 a_n8300_8799.n45 a_n8300_8799.n44 0.189894
R927 a_n8300_8799.n45 a_n8300_8799.n28 0.189894
R928 a_n8300_8799.n49 a_n8300_8799.n28 0.189894
R929 a_n8300_8799.n50 a_n8300_8799.n49 0.189894
R930 a_n8300_8799.n51 a_n8300_8799.n50 0.189894
R931 a_n8300_8799.n51 a_n8300_8799.n26 0.189894
R932 a_n8300_8799.n55 a_n8300_8799.n26 0.189894
R933 a_n8300_8799.n56 a_n8300_8799.n55 0.189894
R934 a_n8300_8799.n57 a_n8300_8799.n56 0.189894
R935 a_n8300_8799.n57 a_n8300_8799.n24 0.189894
R936 a_n8300_8799.n61 a_n8300_8799.n24 0.189894
R937 a_n8300_8799.n62 a_n8300_8799.n61 0.189894
R938 a_n8300_8799.n63 a_n8300_8799.n62 0.189894
R939 a_n8300_8799.n63 a_n8300_8799.n22 0.189894
R940 a_n8300_8799.n67 a_n8300_8799.n22 0.189894
R941 a_n8300_8799.n68 a_n8300_8799.n67 0.189894
R942 a_n8300_8799.n69 a_n8300_8799.n68 0.189894
R943 a_n8300_8799.n69 a_n8300_8799.n20 0.189894
R944 a_n8300_8799.n73 a_n8300_8799.n20 0.189894
R945 a_n8300_8799.n74 a_n8300_8799.n73 0.189894
R946 a_n8300_8799.n75 a_n8300_8799.n74 0.189894
R947 a_n8300_8799.n75 a_n8300_8799.n18 0.189894
R948 a_n8300_8799.n79 a_n8300_8799.n18 0.189894
R949 a_n8300_8799.n99 a_n8300_8799.n94 0.189894
R950 a_n8300_8799.n100 a_n8300_8799.n99 0.189894
R951 a_n8300_8799.n101 a_n8300_8799.n100 0.189894
R952 a_n8300_8799.n101 a_n8300_8799.n92 0.189894
R953 a_n8300_8799.n105 a_n8300_8799.n92 0.189894
R954 a_n8300_8799.n106 a_n8300_8799.n105 0.189894
R955 a_n8300_8799.n107 a_n8300_8799.n106 0.189894
R956 a_n8300_8799.n107 a_n8300_8799.n90 0.189894
R957 a_n8300_8799.n111 a_n8300_8799.n90 0.189894
R958 a_n8300_8799.n112 a_n8300_8799.n111 0.189894
R959 a_n8300_8799.n113 a_n8300_8799.n112 0.189894
R960 a_n8300_8799.n113 a_n8300_8799.n88 0.189894
R961 a_n8300_8799.n117 a_n8300_8799.n88 0.189894
R962 a_n8300_8799.n118 a_n8300_8799.n117 0.189894
R963 a_n8300_8799.n119 a_n8300_8799.n118 0.189894
R964 a_n8300_8799.n119 a_n8300_8799.n86 0.189894
R965 a_n8300_8799.n123 a_n8300_8799.n86 0.189894
R966 a_n8300_8799.n124 a_n8300_8799.n123 0.189894
R967 a_n8300_8799.n125 a_n8300_8799.n124 0.189894
R968 a_n8300_8799.n125 a_n8300_8799.n84 0.189894
R969 a_n8300_8799.n129 a_n8300_8799.n84 0.189894
R970 a_n8300_8799.n130 a_n8300_8799.n129 0.189894
R971 a_n8300_8799.n131 a_n8300_8799.n130 0.189894
R972 a_n8300_8799.n131 a_n8300_8799.n82 0.189894
R973 a_n8300_8799.n135 a_n8300_8799.n82 0.189894
R974 a_n8300_8799.n136 a_n8300_8799.n135 0.189894
R975 a_n8300_8799.n137 a_n8300_8799.n136 0.189894
R976 a_n8300_8799.n137 a_n8300_8799.n80 0.189894
R977 a_n8300_8799.n141 a_n8300_8799.n80 0.189894
R978 a_n8300_8799.n162 a_n8300_8799.n157 0.189894
R979 a_n8300_8799.n163 a_n8300_8799.n162 0.189894
R980 a_n8300_8799.n164 a_n8300_8799.n163 0.189894
R981 a_n8300_8799.n164 a_n8300_8799.n155 0.189894
R982 a_n8300_8799.n168 a_n8300_8799.n155 0.189894
R983 a_n8300_8799.n169 a_n8300_8799.n168 0.189894
R984 a_n8300_8799.n170 a_n8300_8799.n169 0.189894
R985 a_n8300_8799.n170 a_n8300_8799.n153 0.189894
R986 a_n8300_8799.n174 a_n8300_8799.n153 0.189894
R987 a_n8300_8799.n175 a_n8300_8799.n174 0.189894
R988 a_n8300_8799.n176 a_n8300_8799.n175 0.189894
R989 a_n8300_8799.n176 a_n8300_8799.n151 0.189894
R990 a_n8300_8799.n180 a_n8300_8799.n151 0.189894
R991 a_n8300_8799.n181 a_n8300_8799.n180 0.189894
R992 a_n8300_8799.n182 a_n8300_8799.n181 0.189894
R993 a_n8300_8799.n182 a_n8300_8799.n149 0.189894
R994 a_n8300_8799.n186 a_n8300_8799.n149 0.189894
R995 a_n8300_8799.n187 a_n8300_8799.n186 0.189894
R996 a_n8300_8799.n188 a_n8300_8799.n187 0.189894
R997 a_n8300_8799.n188 a_n8300_8799.n147 0.189894
R998 a_n8300_8799.n192 a_n8300_8799.n147 0.189894
R999 a_n8300_8799.n193 a_n8300_8799.n192 0.189894
R1000 a_n8300_8799.n194 a_n8300_8799.n193 0.189894
R1001 a_n8300_8799.n194 a_n8300_8799.n145 0.189894
R1002 a_n8300_8799.n198 a_n8300_8799.n145 0.189894
R1003 a_n8300_8799.n199 a_n8300_8799.n198 0.189894
R1004 a_n8300_8799.n200 a_n8300_8799.n199 0.189894
R1005 a_n8300_8799.n200 a_n8300_8799.n143 0.189894
R1006 a_n8300_8799.n204 a_n8300_8799.n143 0.189894
R1007 gnd.n6959 gnd.n454 1305.8
R1008 gnd.n4906 gnd.n4905 939.716
R1009 gnd.n7371 gnd.n107 795.207
R1010 gnd.n7535 gnd.n103 795.207
R1011 gnd.n1498 gnd.n1445 795.207
R1012 gnd.n4421 gnd.n1500 795.207
R1013 gnd.n4666 gnd.n1274 795.207
R1014 gnd.n3145 gnd.n1272 795.207
R1015 gnd.n2471 gnd.n960 795.207
R1016 gnd.n2533 gnd.n2472 795.207
R1017 gnd.n7533 gnd.n109 775.989
R1018 gnd.n177 gnd.n105 775.989
R1019 gnd.n4424 gnd.n4423 775.989
R1020 gnd.n4496 gnd.n1449 775.989
R1021 gnd.n4668 gnd.n1269 775.989
R1022 gnd.n2325 gnd.n1271 775.989
R1023 gnd.n4827 gnd.n4826 775.989
R1024 gnd.n4903 gnd.n964 775.989
R1025 gnd.n6311 gnd.n929 766.379
R1026 gnd.n6227 gnd.n931 766.379
R1027 gnd.n5415 gnd.n5318 766.379
R1028 gnd.n5411 gnd.n5316 766.379
R1029 gnd.n6308 gnd.n4908 756.769
R1030 gnd.n6277 gnd.n932 756.769
R1031 gnd.n5594 gnd.n5225 756.769
R1032 gnd.n5592 gnd.n5228 756.769
R1033 gnd.n3191 gnd.n1279 711.122
R1034 gnd.n4508 gnd.n1405 711.122
R1035 gnd.n3201 gnd.n2177 711.122
R1036 gnd.n4209 gnd.n1408 711.122
R1037 gnd.n6501 gnd.n727 670.282
R1038 gnd.n6958 gnd.n455 670.282
R1039 gnd.n7172 gnd.n7170 670.282
R1040 gnd.n2411 gnd.n895 670.282
R1041 gnd.n730 gnd.n727 585
R1042 gnd.n6499 gnd.n727 585
R1043 gnd.n6497 gnd.n6496 585
R1044 gnd.n6498 gnd.n6497 585
R1045 gnd.n6495 gnd.n729 585
R1046 gnd.n729 gnd.n728 585
R1047 gnd.n6494 gnd.n6493 585
R1048 gnd.n6493 gnd.n6492 585
R1049 gnd.n735 gnd.n734 585
R1050 gnd.n6491 gnd.n735 585
R1051 gnd.n6489 gnd.n6488 585
R1052 gnd.n6490 gnd.n6489 585
R1053 gnd.n6487 gnd.n737 585
R1054 gnd.n737 gnd.n736 585
R1055 gnd.n6486 gnd.n6485 585
R1056 gnd.n6485 gnd.n6484 585
R1057 gnd.n743 gnd.n742 585
R1058 gnd.n6483 gnd.n743 585
R1059 gnd.n6481 gnd.n6480 585
R1060 gnd.n6482 gnd.n6481 585
R1061 gnd.n6479 gnd.n745 585
R1062 gnd.n745 gnd.n744 585
R1063 gnd.n6478 gnd.n6477 585
R1064 gnd.n6477 gnd.n6476 585
R1065 gnd.n751 gnd.n750 585
R1066 gnd.n6475 gnd.n751 585
R1067 gnd.n6473 gnd.n6472 585
R1068 gnd.n6474 gnd.n6473 585
R1069 gnd.n6471 gnd.n753 585
R1070 gnd.n753 gnd.n752 585
R1071 gnd.n6470 gnd.n6469 585
R1072 gnd.n6469 gnd.n6468 585
R1073 gnd.n759 gnd.n758 585
R1074 gnd.n6467 gnd.n759 585
R1075 gnd.n6465 gnd.n6464 585
R1076 gnd.n6466 gnd.n6465 585
R1077 gnd.n6463 gnd.n761 585
R1078 gnd.n761 gnd.n760 585
R1079 gnd.n6462 gnd.n6461 585
R1080 gnd.n6461 gnd.n6460 585
R1081 gnd.n767 gnd.n766 585
R1082 gnd.n6459 gnd.n767 585
R1083 gnd.n6457 gnd.n6456 585
R1084 gnd.n6458 gnd.n6457 585
R1085 gnd.n6455 gnd.n769 585
R1086 gnd.n769 gnd.n768 585
R1087 gnd.n6454 gnd.n6453 585
R1088 gnd.n6453 gnd.n6452 585
R1089 gnd.n775 gnd.n774 585
R1090 gnd.n6451 gnd.n775 585
R1091 gnd.n6449 gnd.n6448 585
R1092 gnd.n6450 gnd.n6449 585
R1093 gnd.n6447 gnd.n777 585
R1094 gnd.n777 gnd.n776 585
R1095 gnd.n6446 gnd.n6445 585
R1096 gnd.n6445 gnd.n6444 585
R1097 gnd.n783 gnd.n782 585
R1098 gnd.n6443 gnd.n783 585
R1099 gnd.n6441 gnd.n6440 585
R1100 gnd.n6442 gnd.n6441 585
R1101 gnd.n6439 gnd.n785 585
R1102 gnd.n785 gnd.n784 585
R1103 gnd.n6438 gnd.n6437 585
R1104 gnd.n6437 gnd.n6436 585
R1105 gnd.n791 gnd.n790 585
R1106 gnd.n6435 gnd.n791 585
R1107 gnd.n6433 gnd.n6432 585
R1108 gnd.n6434 gnd.n6433 585
R1109 gnd.n6431 gnd.n793 585
R1110 gnd.n793 gnd.n792 585
R1111 gnd.n6430 gnd.n6429 585
R1112 gnd.n6429 gnd.n6428 585
R1113 gnd.n799 gnd.n798 585
R1114 gnd.n6427 gnd.n799 585
R1115 gnd.n6425 gnd.n6424 585
R1116 gnd.n6426 gnd.n6425 585
R1117 gnd.n6423 gnd.n801 585
R1118 gnd.n801 gnd.n800 585
R1119 gnd.n6422 gnd.n6421 585
R1120 gnd.n6421 gnd.n6420 585
R1121 gnd.n807 gnd.n806 585
R1122 gnd.n6419 gnd.n807 585
R1123 gnd.n6417 gnd.n6416 585
R1124 gnd.n6418 gnd.n6417 585
R1125 gnd.n6415 gnd.n809 585
R1126 gnd.n809 gnd.n808 585
R1127 gnd.n6414 gnd.n6413 585
R1128 gnd.n6413 gnd.n6412 585
R1129 gnd.n815 gnd.n814 585
R1130 gnd.n6411 gnd.n815 585
R1131 gnd.n6409 gnd.n6408 585
R1132 gnd.n6410 gnd.n6409 585
R1133 gnd.n6407 gnd.n817 585
R1134 gnd.n817 gnd.n816 585
R1135 gnd.n6406 gnd.n6405 585
R1136 gnd.n6405 gnd.n6404 585
R1137 gnd.n823 gnd.n822 585
R1138 gnd.n6403 gnd.n823 585
R1139 gnd.n6401 gnd.n6400 585
R1140 gnd.n6402 gnd.n6401 585
R1141 gnd.n6399 gnd.n825 585
R1142 gnd.n825 gnd.n824 585
R1143 gnd.n6398 gnd.n6397 585
R1144 gnd.n6397 gnd.n6396 585
R1145 gnd.n831 gnd.n830 585
R1146 gnd.n6395 gnd.n831 585
R1147 gnd.n6393 gnd.n6392 585
R1148 gnd.n6394 gnd.n6393 585
R1149 gnd.n6391 gnd.n833 585
R1150 gnd.n833 gnd.n832 585
R1151 gnd.n6390 gnd.n6389 585
R1152 gnd.n6389 gnd.n6388 585
R1153 gnd.n839 gnd.n838 585
R1154 gnd.n6387 gnd.n839 585
R1155 gnd.n6385 gnd.n6384 585
R1156 gnd.n6386 gnd.n6385 585
R1157 gnd.n6383 gnd.n841 585
R1158 gnd.n841 gnd.n840 585
R1159 gnd.n6382 gnd.n6381 585
R1160 gnd.n6381 gnd.n6380 585
R1161 gnd.n847 gnd.n846 585
R1162 gnd.n6379 gnd.n847 585
R1163 gnd.n6377 gnd.n6376 585
R1164 gnd.n6378 gnd.n6377 585
R1165 gnd.n6375 gnd.n849 585
R1166 gnd.n849 gnd.n848 585
R1167 gnd.n6374 gnd.n6373 585
R1168 gnd.n6373 gnd.n6372 585
R1169 gnd.n855 gnd.n854 585
R1170 gnd.n6371 gnd.n855 585
R1171 gnd.n6369 gnd.n6368 585
R1172 gnd.n6370 gnd.n6369 585
R1173 gnd.n6367 gnd.n857 585
R1174 gnd.n857 gnd.n856 585
R1175 gnd.n6366 gnd.n6365 585
R1176 gnd.n6365 gnd.n6364 585
R1177 gnd.n863 gnd.n862 585
R1178 gnd.n6363 gnd.n863 585
R1179 gnd.n6361 gnd.n6360 585
R1180 gnd.n6362 gnd.n6361 585
R1181 gnd.n6359 gnd.n865 585
R1182 gnd.n865 gnd.n864 585
R1183 gnd.n6358 gnd.n6357 585
R1184 gnd.n6357 gnd.n6356 585
R1185 gnd.n871 gnd.n870 585
R1186 gnd.n6355 gnd.n871 585
R1187 gnd.n6353 gnd.n6352 585
R1188 gnd.n6354 gnd.n6353 585
R1189 gnd.n6351 gnd.n873 585
R1190 gnd.n873 gnd.n872 585
R1191 gnd.n6350 gnd.n6349 585
R1192 gnd.n6349 gnd.n6348 585
R1193 gnd.n879 gnd.n878 585
R1194 gnd.n6347 gnd.n879 585
R1195 gnd.n6345 gnd.n6344 585
R1196 gnd.n6346 gnd.n6345 585
R1197 gnd.n6343 gnd.n881 585
R1198 gnd.n881 gnd.n880 585
R1199 gnd.n6342 gnd.n6341 585
R1200 gnd.n6341 gnd.n6340 585
R1201 gnd.n887 gnd.n886 585
R1202 gnd.n6339 gnd.n887 585
R1203 gnd.n6337 gnd.n6336 585
R1204 gnd.n6338 gnd.n6337 585
R1205 gnd.n6335 gnd.n889 585
R1206 gnd.n889 gnd.n888 585
R1207 gnd.n6334 gnd.n6333 585
R1208 gnd.n6333 gnd.n6332 585
R1209 gnd.n6502 gnd.n6501 585
R1210 gnd.n6501 gnd.n6500 585
R1211 gnd.n725 gnd.n724 585
R1212 gnd.n724 gnd.n723 585
R1213 gnd.n6507 gnd.n6506 585
R1214 gnd.n6508 gnd.n6507 585
R1215 gnd.n722 gnd.n721 585
R1216 gnd.n6509 gnd.n722 585
R1217 gnd.n6512 gnd.n6511 585
R1218 gnd.n6511 gnd.n6510 585
R1219 gnd.n719 gnd.n718 585
R1220 gnd.n718 gnd.n717 585
R1221 gnd.n6517 gnd.n6516 585
R1222 gnd.n6518 gnd.n6517 585
R1223 gnd.n716 gnd.n715 585
R1224 gnd.n6519 gnd.n716 585
R1225 gnd.n6522 gnd.n6521 585
R1226 gnd.n6521 gnd.n6520 585
R1227 gnd.n713 gnd.n712 585
R1228 gnd.n712 gnd.n711 585
R1229 gnd.n6527 gnd.n6526 585
R1230 gnd.n6528 gnd.n6527 585
R1231 gnd.n710 gnd.n709 585
R1232 gnd.n6529 gnd.n710 585
R1233 gnd.n6532 gnd.n6531 585
R1234 gnd.n6531 gnd.n6530 585
R1235 gnd.n707 gnd.n706 585
R1236 gnd.n706 gnd.n705 585
R1237 gnd.n6537 gnd.n6536 585
R1238 gnd.n6538 gnd.n6537 585
R1239 gnd.n704 gnd.n703 585
R1240 gnd.n6539 gnd.n704 585
R1241 gnd.n6542 gnd.n6541 585
R1242 gnd.n6541 gnd.n6540 585
R1243 gnd.n701 gnd.n700 585
R1244 gnd.n700 gnd.n699 585
R1245 gnd.n6547 gnd.n6546 585
R1246 gnd.n6548 gnd.n6547 585
R1247 gnd.n698 gnd.n697 585
R1248 gnd.n6549 gnd.n698 585
R1249 gnd.n6552 gnd.n6551 585
R1250 gnd.n6551 gnd.n6550 585
R1251 gnd.n695 gnd.n694 585
R1252 gnd.n694 gnd.n693 585
R1253 gnd.n6557 gnd.n6556 585
R1254 gnd.n6558 gnd.n6557 585
R1255 gnd.n692 gnd.n691 585
R1256 gnd.n6559 gnd.n692 585
R1257 gnd.n6562 gnd.n6561 585
R1258 gnd.n6561 gnd.n6560 585
R1259 gnd.n689 gnd.n688 585
R1260 gnd.n688 gnd.n687 585
R1261 gnd.n6567 gnd.n6566 585
R1262 gnd.n6568 gnd.n6567 585
R1263 gnd.n686 gnd.n685 585
R1264 gnd.n6569 gnd.n686 585
R1265 gnd.n6572 gnd.n6571 585
R1266 gnd.n6571 gnd.n6570 585
R1267 gnd.n683 gnd.n682 585
R1268 gnd.n682 gnd.n681 585
R1269 gnd.n6577 gnd.n6576 585
R1270 gnd.n6578 gnd.n6577 585
R1271 gnd.n680 gnd.n679 585
R1272 gnd.n6579 gnd.n680 585
R1273 gnd.n6582 gnd.n6581 585
R1274 gnd.n6581 gnd.n6580 585
R1275 gnd.n677 gnd.n676 585
R1276 gnd.n676 gnd.n675 585
R1277 gnd.n6587 gnd.n6586 585
R1278 gnd.n6588 gnd.n6587 585
R1279 gnd.n674 gnd.n673 585
R1280 gnd.n6589 gnd.n674 585
R1281 gnd.n6592 gnd.n6591 585
R1282 gnd.n6591 gnd.n6590 585
R1283 gnd.n671 gnd.n670 585
R1284 gnd.n670 gnd.n669 585
R1285 gnd.n6597 gnd.n6596 585
R1286 gnd.n6598 gnd.n6597 585
R1287 gnd.n668 gnd.n667 585
R1288 gnd.n6599 gnd.n668 585
R1289 gnd.n6602 gnd.n6601 585
R1290 gnd.n6601 gnd.n6600 585
R1291 gnd.n665 gnd.n664 585
R1292 gnd.n664 gnd.n663 585
R1293 gnd.n6607 gnd.n6606 585
R1294 gnd.n6608 gnd.n6607 585
R1295 gnd.n662 gnd.n661 585
R1296 gnd.n6609 gnd.n662 585
R1297 gnd.n6612 gnd.n6611 585
R1298 gnd.n6611 gnd.n6610 585
R1299 gnd.n659 gnd.n658 585
R1300 gnd.n658 gnd.n657 585
R1301 gnd.n6617 gnd.n6616 585
R1302 gnd.n6618 gnd.n6617 585
R1303 gnd.n656 gnd.n655 585
R1304 gnd.n6619 gnd.n656 585
R1305 gnd.n6622 gnd.n6621 585
R1306 gnd.n6621 gnd.n6620 585
R1307 gnd.n653 gnd.n652 585
R1308 gnd.n652 gnd.n651 585
R1309 gnd.n6627 gnd.n6626 585
R1310 gnd.n6628 gnd.n6627 585
R1311 gnd.n650 gnd.n649 585
R1312 gnd.n6629 gnd.n650 585
R1313 gnd.n6632 gnd.n6631 585
R1314 gnd.n6631 gnd.n6630 585
R1315 gnd.n647 gnd.n646 585
R1316 gnd.n646 gnd.n645 585
R1317 gnd.n6637 gnd.n6636 585
R1318 gnd.n6638 gnd.n6637 585
R1319 gnd.n644 gnd.n643 585
R1320 gnd.n6639 gnd.n644 585
R1321 gnd.n6642 gnd.n6641 585
R1322 gnd.n6641 gnd.n6640 585
R1323 gnd.n641 gnd.n640 585
R1324 gnd.n640 gnd.n639 585
R1325 gnd.n6647 gnd.n6646 585
R1326 gnd.n6648 gnd.n6647 585
R1327 gnd.n638 gnd.n637 585
R1328 gnd.n6649 gnd.n638 585
R1329 gnd.n6652 gnd.n6651 585
R1330 gnd.n6651 gnd.n6650 585
R1331 gnd.n635 gnd.n634 585
R1332 gnd.n634 gnd.n633 585
R1333 gnd.n6657 gnd.n6656 585
R1334 gnd.n6658 gnd.n6657 585
R1335 gnd.n632 gnd.n631 585
R1336 gnd.n6659 gnd.n632 585
R1337 gnd.n6662 gnd.n6661 585
R1338 gnd.n6661 gnd.n6660 585
R1339 gnd.n629 gnd.n628 585
R1340 gnd.n628 gnd.n627 585
R1341 gnd.n6667 gnd.n6666 585
R1342 gnd.n6668 gnd.n6667 585
R1343 gnd.n626 gnd.n625 585
R1344 gnd.n6669 gnd.n626 585
R1345 gnd.n6672 gnd.n6671 585
R1346 gnd.n6671 gnd.n6670 585
R1347 gnd.n623 gnd.n622 585
R1348 gnd.n622 gnd.n621 585
R1349 gnd.n6677 gnd.n6676 585
R1350 gnd.n6678 gnd.n6677 585
R1351 gnd.n620 gnd.n619 585
R1352 gnd.n6679 gnd.n620 585
R1353 gnd.n6682 gnd.n6681 585
R1354 gnd.n6681 gnd.n6680 585
R1355 gnd.n617 gnd.n616 585
R1356 gnd.n616 gnd.n615 585
R1357 gnd.n6687 gnd.n6686 585
R1358 gnd.n6688 gnd.n6687 585
R1359 gnd.n614 gnd.n613 585
R1360 gnd.n6689 gnd.n614 585
R1361 gnd.n6692 gnd.n6691 585
R1362 gnd.n6691 gnd.n6690 585
R1363 gnd.n611 gnd.n610 585
R1364 gnd.n610 gnd.n609 585
R1365 gnd.n6697 gnd.n6696 585
R1366 gnd.n6698 gnd.n6697 585
R1367 gnd.n608 gnd.n607 585
R1368 gnd.n6699 gnd.n608 585
R1369 gnd.n6702 gnd.n6701 585
R1370 gnd.n6701 gnd.n6700 585
R1371 gnd.n605 gnd.n604 585
R1372 gnd.n604 gnd.n603 585
R1373 gnd.n6707 gnd.n6706 585
R1374 gnd.n6708 gnd.n6707 585
R1375 gnd.n602 gnd.n601 585
R1376 gnd.n6709 gnd.n602 585
R1377 gnd.n6712 gnd.n6711 585
R1378 gnd.n6711 gnd.n6710 585
R1379 gnd.n599 gnd.n598 585
R1380 gnd.n598 gnd.n597 585
R1381 gnd.n6717 gnd.n6716 585
R1382 gnd.n6718 gnd.n6717 585
R1383 gnd.n596 gnd.n595 585
R1384 gnd.n6719 gnd.n596 585
R1385 gnd.n6722 gnd.n6721 585
R1386 gnd.n6721 gnd.n6720 585
R1387 gnd.n593 gnd.n592 585
R1388 gnd.n592 gnd.n591 585
R1389 gnd.n6727 gnd.n6726 585
R1390 gnd.n6728 gnd.n6727 585
R1391 gnd.n590 gnd.n589 585
R1392 gnd.n6729 gnd.n590 585
R1393 gnd.n6732 gnd.n6731 585
R1394 gnd.n6731 gnd.n6730 585
R1395 gnd.n587 gnd.n586 585
R1396 gnd.n586 gnd.n585 585
R1397 gnd.n6737 gnd.n6736 585
R1398 gnd.n6738 gnd.n6737 585
R1399 gnd.n584 gnd.n583 585
R1400 gnd.n6739 gnd.n584 585
R1401 gnd.n6742 gnd.n6741 585
R1402 gnd.n6741 gnd.n6740 585
R1403 gnd.n581 gnd.n580 585
R1404 gnd.n580 gnd.n579 585
R1405 gnd.n6747 gnd.n6746 585
R1406 gnd.n6748 gnd.n6747 585
R1407 gnd.n578 gnd.n577 585
R1408 gnd.n6749 gnd.n578 585
R1409 gnd.n6752 gnd.n6751 585
R1410 gnd.n6751 gnd.n6750 585
R1411 gnd.n575 gnd.n574 585
R1412 gnd.n574 gnd.n573 585
R1413 gnd.n6757 gnd.n6756 585
R1414 gnd.n6758 gnd.n6757 585
R1415 gnd.n572 gnd.n571 585
R1416 gnd.n6759 gnd.n572 585
R1417 gnd.n6762 gnd.n6761 585
R1418 gnd.n6761 gnd.n6760 585
R1419 gnd.n569 gnd.n568 585
R1420 gnd.n568 gnd.n567 585
R1421 gnd.n6767 gnd.n6766 585
R1422 gnd.n6768 gnd.n6767 585
R1423 gnd.n566 gnd.n565 585
R1424 gnd.n6769 gnd.n566 585
R1425 gnd.n6772 gnd.n6771 585
R1426 gnd.n6771 gnd.n6770 585
R1427 gnd.n563 gnd.n562 585
R1428 gnd.n562 gnd.n561 585
R1429 gnd.n6777 gnd.n6776 585
R1430 gnd.n6778 gnd.n6777 585
R1431 gnd.n560 gnd.n559 585
R1432 gnd.n6779 gnd.n560 585
R1433 gnd.n6782 gnd.n6781 585
R1434 gnd.n6781 gnd.n6780 585
R1435 gnd.n557 gnd.n556 585
R1436 gnd.n556 gnd.n555 585
R1437 gnd.n6787 gnd.n6786 585
R1438 gnd.n6788 gnd.n6787 585
R1439 gnd.n554 gnd.n553 585
R1440 gnd.n6789 gnd.n554 585
R1441 gnd.n6792 gnd.n6791 585
R1442 gnd.n6791 gnd.n6790 585
R1443 gnd.n551 gnd.n550 585
R1444 gnd.n550 gnd.n549 585
R1445 gnd.n6797 gnd.n6796 585
R1446 gnd.n6798 gnd.n6797 585
R1447 gnd.n548 gnd.n547 585
R1448 gnd.n6799 gnd.n548 585
R1449 gnd.n6802 gnd.n6801 585
R1450 gnd.n6801 gnd.n6800 585
R1451 gnd.n545 gnd.n544 585
R1452 gnd.n544 gnd.n543 585
R1453 gnd.n6807 gnd.n6806 585
R1454 gnd.n6808 gnd.n6807 585
R1455 gnd.n542 gnd.n541 585
R1456 gnd.n6809 gnd.n542 585
R1457 gnd.n6812 gnd.n6811 585
R1458 gnd.n6811 gnd.n6810 585
R1459 gnd.n539 gnd.n538 585
R1460 gnd.n538 gnd.n537 585
R1461 gnd.n6817 gnd.n6816 585
R1462 gnd.n6818 gnd.n6817 585
R1463 gnd.n536 gnd.n535 585
R1464 gnd.n6819 gnd.n536 585
R1465 gnd.n6822 gnd.n6821 585
R1466 gnd.n6821 gnd.n6820 585
R1467 gnd.n533 gnd.n532 585
R1468 gnd.n532 gnd.n531 585
R1469 gnd.n6827 gnd.n6826 585
R1470 gnd.n6828 gnd.n6827 585
R1471 gnd.n530 gnd.n529 585
R1472 gnd.n6829 gnd.n530 585
R1473 gnd.n6832 gnd.n6831 585
R1474 gnd.n6831 gnd.n6830 585
R1475 gnd.n527 gnd.n526 585
R1476 gnd.n526 gnd.n525 585
R1477 gnd.n6837 gnd.n6836 585
R1478 gnd.n6838 gnd.n6837 585
R1479 gnd.n524 gnd.n523 585
R1480 gnd.n6839 gnd.n524 585
R1481 gnd.n6842 gnd.n6841 585
R1482 gnd.n6841 gnd.n6840 585
R1483 gnd.n521 gnd.n520 585
R1484 gnd.n520 gnd.n519 585
R1485 gnd.n6847 gnd.n6846 585
R1486 gnd.n6848 gnd.n6847 585
R1487 gnd.n518 gnd.n517 585
R1488 gnd.n6849 gnd.n518 585
R1489 gnd.n6852 gnd.n6851 585
R1490 gnd.n6851 gnd.n6850 585
R1491 gnd.n515 gnd.n514 585
R1492 gnd.n514 gnd.n513 585
R1493 gnd.n6857 gnd.n6856 585
R1494 gnd.n6858 gnd.n6857 585
R1495 gnd.n512 gnd.n511 585
R1496 gnd.n6859 gnd.n512 585
R1497 gnd.n6862 gnd.n6861 585
R1498 gnd.n6861 gnd.n6860 585
R1499 gnd.n509 gnd.n508 585
R1500 gnd.n508 gnd.n507 585
R1501 gnd.n6867 gnd.n6866 585
R1502 gnd.n6868 gnd.n6867 585
R1503 gnd.n506 gnd.n505 585
R1504 gnd.n6869 gnd.n506 585
R1505 gnd.n6872 gnd.n6871 585
R1506 gnd.n6871 gnd.n6870 585
R1507 gnd.n503 gnd.n502 585
R1508 gnd.n502 gnd.n501 585
R1509 gnd.n6877 gnd.n6876 585
R1510 gnd.n6878 gnd.n6877 585
R1511 gnd.n500 gnd.n499 585
R1512 gnd.n6879 gnd.n500 585
R1513 gnd.n6882 gnd.n6881 585
R1514 gnd.n6881 gnd.n6880 585
R1515 gnd.n497 gnd.n496 585
R1516 gnd.n496 gnd.n495 585
R1517 gnd.n6887 gnd.n6886 585
R1518 gnd.n6888 gnd.n6887 585
R1519 gnd.n494 gnd.n493 585
R1520 gnd.n6889 gnd.n494 585
R1521 gnd.n6892 gnd.n6891 585
R1522 gnd.n6891 gnd.n6890 585
R1523 gnd.n491 gnd.n490 585
R1524 gnd.n490 gnd.n489 585
R1525 gnd.n6897 gnd.n6896 585
R1526 gnd.n6898 gnd.n6897 585
R1527 gnd.n488 gnd.n487 585
R1528 gnd.n6899 gnd.n488 585
R1529 gnd.n6902 gnd.n6901 585
R1530 gnd.n6901 gnd.n6900 585
R1531 gnd.n485 gnd.n484 585
R1532 gnd.n484 gnd.n483 585
R1533 gnd.n6907 gnd.n6906 585
R1534 gnd.n6908 gnd.n6907 585
R1535 gnd.n482 gnd.n481 585
R1536 gnd.n6909 gnd.n482 585
R1537 gnd.n6912 gnd.n6911 585
R1538 gnd.n6911 gnd.n6910 585
R1539 gnd.n479 gnd.n478 585
R1540 gnd.n478 gnd.n477 585
R1541 gnd.n6917 gnd.n6916 585
R1542 gnd.n6918 gnd.n6917 585
R1543 gnd.n476 gnd.n475 585
R1544 gnd.n6919 gnd.n476 585
R1545 gnd.n6922 gnd.n6921 585
R1546 gnd.n6921 gnd.n6920 585
R1547 gnd.n473 gnd.n472 585
R1548 gnd.n472 gnd.n471 585
R1549 gnd.n6927 gnd.n6926 585
R1550 gnd.n6928 gnd.n6927 585
R1551 gnd.n470 gnd.n469 585
R1552 gnd.n6929 gnd.n470 585
R1553 gnd.n6932 gnd.n6931 585
R1554 gnd.n6931 gnd.n6930 585
R1555 gnd.n467 gnd.n466 585
R1556 gnd.n466 gnd.n465 585
R1557 gnd.n6937 gnd.n6936 585
R1558 gnd.n6938 gnd.n6937 585
R1559 gnd.n464 gnd.n463 585
R1560 gnd.n6939 gnd.n464 585
R1561 gnd.n6942 gnd.n6941 585
R1562 gnd.n6941 gnd.n6940 585
R1563 gnd.n461 gnd.n460 585
R1564 gnd.n460 gnd.n459 585
R1565 gnd.n6948 gnd.n6947 585
R1566 gnd.n6949 gnd.n6948 585
R1567 gnd.n458 gnd.n457 585
R1568 gnd.n6950 gnd.n458 585
R1569 gnd.n6953 gnd.n6952 585
R1570 gnd.n6952 gnd.n6951 585
R1571 gnd.n6954 gnd.n455 585
R1572 gnd.n455 gnd.n454 585
R1573 gnd.n330 gnd.n329 585
R1574 gnd.n7161 gnd.n329 585
R1575 gnd.n7164 gnd.n7163 585
R1576 gnd.n7163 gnd.n7162 585
R1577 gnd.n333 gnd.n332 585
R1578 gnd.n7160 gnd.n333 585
R1579 gnd.n7158 gnd.n7157 585
R1580 gnd.n7159 gnd.n7158 585
R1581 gnd.n336 gnd.n335 585
R1582 gnd.n335 gnd.n334 585
R1583 gnd.n7153 gnd.n7152 585
R1584 gnd.n7152 gnd.n7151 585
R1585 gnd.n339 gnd.n338 585
R1586 gnd.n7150 gnd.n339 585
R1587 gnd.n7148 gnd.n7147 585
R1588 gnd.n7149 gnd.n7148 585
R1589 gnd.n342 gnd.n341 585
R1590 gnd.n341 gnd.n340 585
R1591 gnd.n7143 gnd.n7142 585
R1592 gnd.n7142 gnd.n7141 585
R1593 gnd.n345 gnd.n344 585
R1594 gnd.n7140 gnd.n345 585
R1595 gnd.n7138 gnd.n7137 585
R1596 gnd.n7139 gnd.n7138 585
R1597 gnd.n348 gnd.n347 585
R1598 gnd.n347 gnd.n346 585
R1599 gnd.n7133 gnd.n7132 585
R1600 gnd.n7132 gnd.n7131 585
R1601 gnd.n351 gnd.n350 585
R1602 gnd.n7130 gnd.n351 585
R1603 gnd.n7128 gnd.n7127 585
R1604 gnd.n7129 gnd.n7128 585
R1605 gnd.n354 gnd.n353 585
R1606 gnd.n353 gnd.n352 585
R1607 gnd.n7123 gnd.n7122 585
R1608 gnd.n7122 gnd.n7121 585
R1609 gnd.n357 gnd.n356 585
R1610 gnd.n7120 gnd.n357 585
R1611 gnd.n7118 gnd.n7117 585
R1612 gnd.n7119 gnd.n7118 585
R1613 gnd.n360 gnd.n359 585
R1614 gnd.n359 gnd.n358 585
R1615 gnd.n7113 gnd.n7112 585
R1616 gnd.n7112 gnd.n7111 585
R1617 gnd.n363 gnd.n362 585
R1618 gnd.n7110 gnd.n363 585
R1619 gnd.n7108 gnd.n7107 585
R1620 gnd.n7109 gnd.n7108 585
R1621 gnd.n366 gnd.n365 585
R1622 gnd.n365 gnd.n364 585
R1623 gnd.n7103 gnd.n7102 585
R1624 gnd.n7102 gnd.n7101 585
R1625 gnd.n369 gnd.n368 585
R1626 gnd.n7100 gnd.n369 585
R1627 gnd.n7098 gnd.n7097 585
R1628 gnd.n7099 gnd.n7098 585
R1629 gnd.n372 gnd.n371 585
R1630 gnd.n371 gnd.n370 585
R1631 gnd.n7093 gnd.n7092 585
R1632 gnd.n7092 gnd.n7091 585
R1633 gnd.n375 gnd.n374 585
R1634 gnd.n7090 gnd.n375 585
R1635 gnd.n7088 gnd.n7087 585
R1636 gnd.n7089 gnd.n7088 585
R1637 gnd.n378 gnd.n377 585
R1638 gnd.n377 gnd.n376 585
R1639 gnd.n7083 gnd.n7082 585
R1640 gnd.n7082 gnd.n7081 585
R1641 gnd.n381 gnd.n380 585
R1642 gnd.n7080 gnd.n381 585
R1643 gnd.n7078 gnd.n7077 585
R1644 gnd.n7079 gnd.n7078 585
R1645 gnd.n384 gnd.n383 585
R1646 gnd.n383 gnd.n382 585
R1647 gnd.n7073 gnd.n7072 585
R1648 gnd.n7072 gnd.n7071 585
R1649 gnd.n387 gnd.n386 585
R1650 gnd.n7070 gnd.n387 585
R1651 gnd.n7068 gnd.n7067 585
R1652 gnd.n7069 gnd.n7068 585
R1653 gnd.n390 gnd.n389 585
R1654 gnd.n389 gnd.n388 585
R1655 gnd.n7063 gnd.n7062 585
R1656 gnd.n7062 gnd.n7061 585
R1657 gnd.n393 gnd.n392 585
R1658 gnd.n7060 gnd.n393 585
R1659 gnd.n7058 gnd.n7057 585
R1660 gnd.n7059 gnd.n7058 585
R1661 gnd.n396 gnd.n395 585
R1662 gnd.n395 gnd.n394 585
R1663 gnd.n7053 gnd.n7052 585
R1664 gnd.n7052 gnd.n7051 585
R1665 gnd.n399 gnd.n398 585
R1666 gnd.n7050 gnd.n399 585
R1667 gnd.n7048 gnd.n7047 585
R1668 gnd.n7049 gnd.n7048 585
R1669 gnd.n402 gnd.n401 585
R1670 gnd.n401 gnd.n400 585
R1671 gnd.n7043 gnd.n7042 585
R1672 gnd.n7042 gnd.n7041 585
R1673 gnd.n405 gnd.n404 585
R1674 gnd.n7040 gnd.n405 585
R1675 gnd.n7038 gnd.n7037 585
R1676 gnd.n7039 gnd.n7038 585
R1677 gnd.n408 gnd.n407 585
R1678 gnd.n407 gnd.n406 585
R1679 gnd.n7033 gnd.n7032 585
R1680 gnd.n7032 gnd.n7031 585
R1681 gnd.n411 gnd.n410 585
R1682 gnd.n7030 gnd.n411 585
R1683 gnd.n7028 gnd.n7027 585
R1684 gnd.n7029 gnd.n7028 585
R1685 gnd.n414 gnd.n413 585
R1686 gnd.n413 gnd.n412 585
R1687 gnd.n7023 gnd.n7022 585
R1688 gnd.n7022 gnd.n7021 585
R1689 gnd.n417 gnd.n416 585
R1690 gnd.n7020 gnd.n417 585
R1691 gnd.n7018 gnd.n7017 585
R1692 gnd.n7019 gnd.n7018 585
R1693 gnd.n420 gnd.n419 585
R1694 gnd.n419 gnd.n418 585
R1695 gnd.n7013 gnd.n7012 585
R1696 gnd.n7012 gnd.n7011 585
R1697 gnd.n423 gnd.n422 585
R1698 gnd.n7010 gnd.n423 585
R1699 gnd.n7008 gnd.n7007 585
R1700 gnd.n7009 gnd.n7008 585
R1701 gnd.n426 gnd.n425 585
R1702 gnd.n425 gnd.n424 585
R1703 gnd.n7003 gnd.n7002 585
R1704 gnd.n7002 gnd.n7001 585
R1705 gnd.n429 gnd.n428 585
R1706 gnd.n7000 gnd.n429 585
R1707 gnd.n6998 gnd.n6997 585
R1708 gnd.n6999 gnd.n6998 585
R1709 gnd.n432 gnd.n431 585
R1710 gnd.n431 gnd.n430 585
R1711 gnd.n6993 gnd.n6992 585
R1712 gnd.n6992 gnd.n6991 585
R1713 gnd.n435 gnd.n434 585
R1714 gnd.n6990 gnd.n435 585
R1715 gnd.n6988 gnd.n6987 585
R1716 gnd.n6989 gnd.n6988 585
R1717 gnd.n438 gnd.n437 585
R1718 gnd.n437 gnd.n436 585
R1719 gnd.n6983 gnd.n6982 585
R1720 gnd.n6982 gnd.n6981 585
R1721 gnd.n441 gnd.n440 585
R1722 gnd.n6980 gnd.n441 585
R1723 gnd.n6978 gnd.n6977 585
R1724 gnd.n6979 gnd.n6978 585
R1725 gnd.n444 gnd.n443 585
R1726 gnd.n443 gnd.n442 585
R1727 gnd.n6973 gnd.n6972 585
R1728 gnd.n6972 gnd.n6971 585
R1729 gnd.n447 gnd.n446 585
R1730 gnd.n6970 gnd.n447 585
R1731 gnd.n6968 gnd.n6967 585
R1732 gnd.n6969 gnd.n6968 585
R1733 gnd.n450 gnd.n449 585
R1734 gnd.n449 gnd.n448 585
R1735 gnd.n6963 gnd.n6962 585
R1736 gnd.n6962 gnd.n6961 585
R1737 gnd.n453 gnd.n452 585
R1738 gnd.n6960 gnd.n453 585
R1739 gnd.n6958 gnd.n6957 585
R1740 gnd.n6959 gnd.n6958 585
R1741 gnd.n4666 gnd.n4665 585
R1742 gnd.n4667 gnd.n4666 585
R1743 gnd.n1260 gnd.n1259 585
R1744 gnd.n2831 gnd.n1260 585
R1745 gnd.n4675 gnd.n4674 585
R1746 gnd.n4674 gnd.n4673 585
R1747 gnd.n4676 gnd.n1254 585
R1748 gnd.n2793 gnd.n1254 585
R1749 gnd.n4678 gnd.n4677 585
R1750 gnd.n4679 gnd.n4678 585
R1751 gnd.n1239 gnd.n1238 585
R1752 gnd.n2784 gnd.n1239 585
R1753 gnd.n4687 gnd.n4686 585
R1754 gnd.n4686 gnd.n4685 585
R1755 gnd.n4688 gnd.n1233 585
R1756 gnd.n2776 gnd.n1233 585
R1757 gnd.n4690 gnd.n4689 585
R1758 gnd.n4691 gnd.n4690 585
R1759 gnd.n1217 gnd.n1216 585
R1760 gnd.n2709 gnd.n1217 585
R1761 gnd.n4699 gnd.n4698 585
R1762 gnd.n4698 gnd.n4697 585
R1763 gnd.n4700 gnd.n1211 585
R1764 gnd.n2697 gnd.n1211 585
R1765 gnd.n4702 gnd.n4701 585
R1766 gnd.n4703 gnd.n4702 585
R1767 gnd.n1197 gnd.n1196 585
R1768 gnd.n2692 gnd.n1197 585
R1769 gnd.n4711 gnd.n4710 585
R1770 gnd.n4710 gnd.n4709 585
R1771 gnd.n4712 gnd.n1191 585
R1772 gnd.n2723 gnd.n1191 585
R1773 gnd.n4714 gnd.n4713 585
R1774 gnd.n4715 gnd.n4714 585
R1775 gnd.n1175 gnd.n1174 585
R1776 gnd.n2684 gnd.n1175 585
R1777 gnd.n4723 gnd.n4722 585
R1778 gnd.n4722 gnd.n4721 585
R1779 gnd.n4724 gnd.n1169 585
R1780 gnd.n2676 gnd.n1169 585
R1781 gnd.n4726 gnd.n4725 585
R1782 gnd.n4727 gnd.n4726 585
R1783 gnd.n1156 gnd.n1155 585
R1784 gnd.n2667 gnd.n1156 585
R1785 gnd.n4735 gnd.n4734 585
R1786 gnd.n4734 gnd.n4733 585
R1787 gnd.n4736 gnd.n1150 585
R1788 gnd.n2659 gnd.n1150 585
R1789 gnd.n4738 gnd.n4737 585
R1790 gnd.n4739 gnd.n4738 585
R1791 gnd.n1137 gnd.n1136 585
R1792 gnd.n2627 gnd.n1137 585
R1793 gnd.n4748 gnd.n4747 585
R1794 gnd.n4747 gnd.n4746 585
R1795 gnd.n4749 gnd.n1131 585
R1796 gnd.n2636 gnd.n1131 585
R1797 gnd.n4751 gnd.n4750 585
R1798 gnd.n4752 gnd.n4751 585
R1799 gnd.n1119 gnd.n1118 585
R1800 gnd.n2642 gnd.n1119 585
R1801 gnd.n4760 gnd.n4759 585
R1802 gnd.n4759 gnd.n4758 585
R1803 gnd.n4761 gnd.n1113 585
R1804 gnd.n2648 gnd.n1113 585
R1805 gnd.n4763 gnd.n4762 585
R1806 gnd.n4764 gnd.n4763 585
R1807 gnd.n1096 gnd.n1095 585
R1808 gnd.n2592 gnd.n1096 585
R1809 gnd.n4772 gnd.n4771 585
R1810 gnd.n4771 gnd.n4770 585
R1811 gnd.n4773 gnd.n1090 585
R1812 gnd.n1098 gnd.n1090 585
R1813 gnd.n4775 gnd.n4774 585
R1814 gnd.n4776 gnd.n4775 585
R1815 gnd.n1077 gnd.n1076 585
R1816 gnd.n1080 gnd.n1077 585
R1817 gnd.n4784 gnd.n4783 585
R1818 gnd.n4783 gnd.n4782 585
R1819 gnd.n4785 gnd.n1071 585
R1820 gnd.n1071 gnd.n1070 585
R1821 gnd.n4787 gnd.n4786 585
R1822 gnd.n4788 gnd.n4787 585
R1823 gnd.n1056 gnd.n1055 585
R1824 gnd.n1067 gnd.n1056 585
R1825 gnd.n4796 gnd.n4795 585
R1826 gnd.n4795 gnd.n4794 585
R1827 gnd.n4797 gnd.n1050 585
R1828 gnd.n1057 gnd.n1050 585
R1829 gnd.n4799 gnd.n4798 585
R1830 gnd.n4800 gnd.n4799 585
R1831 gnd.n1037 gnd.n1036 585
R1832 gnd.n1040 gnd.n1037 585
R1833 gnd.n4808 gnd.n4807 585
R1834 gnd.n4807 gnd.n4806 585
R1835 gnd.n4809 gnd.n1031 585
R1836 gnd.n1031 gnd.n1029 585
R1837 gnd.n4811 gnd.n4810 585
R1838 gnd.n4812 gnd.n4811 585
R1839 gnd.n1032 gnd.n1030 585
R1840 gnd.n1030 gnd.n1017 585
R1841 gnd.n2538 gnd.n1018 585
R1842 gnd.n4818 gnd.n1018 585
R1843 gnd.n2475 gnd.n2473 585
R1844 gnd.n2473 gnd.n1015 585
R1845 gnd.n2543 gnd.n2542 585
R1846 gnd.n2550 gnd.n2543 585
R1847 gnd.n2474 gnd.n2472 585
R1848 gnd.n2472 gnd.n961 585
R1849 gnd.n2534 gnd.n2533 585
R1850 gnd.n2532 gnd.n2531 585
R1851 gnd.n2530 gnd.n2529 585
R1852 gnd.n2528 gnd.n2527 585
R1853 gnd.n2526 gnd.n2525 585
R1854 gnd.n2524 gnd.n2523 585
R1855 gnd.n2522 gnd.n2521 585
R1856 gnd.n2520 gnd.n2519 585
R1857 gnd.n2518 gnd.n2517 585
R1858 gnd.n2516 gnd.n2515 585
R1859 gnd.n2514 gnd.n2513 585
R1860 gnd.n2512 gnd.n2511 585
R1861 gnd.n2510 gnd.n2509 585
R1862 gnd.n2508 gnd.n2507 585
R1863 gnd.n2506 gnd.n2505 585
R1864 gnd.n2504 gnd.n2503 585
R1865 gnd.n2502 gnd.n2501 585
R1866 gnd.n2494 gnd.n2491 585
R1867 gnd.n2497 gnd.n960 585
R1868 gnd.n4905 gnd.n960 585
R1869 gnd.n3146 gnd.n3145 585
R1870 gnd.n2248 gnd.n2240 585
R1871 gnd.n3153 gnd.n2237 585
R1872 gnd.n3154 gnd.n2236 585
R1873 gnd.n2262 gnd.n2230 585
R1874 gnd.n3161 gnd.n2229 585
R1875 gnd.n3162 gnd.n2228 585
R1876 gnd.n2260 gnd.n2220 585
R1877 gnd.n3169 gnd.n2219 585
R1878 gnd.n3170 gnd.n2218 585
R1879 gnd.n2257 gnd.n2212 585
R1880 gnd.n3177 gnd.n2211 585
R1881 gnd.n3178 gnd.n2210 585
R1882 gnd.n2255 gnd.n2203 585
R1883 gnd.n3185 gnd.n2202 585
R1884 gnd.n3186 gnd.n2201 585
R1885 gnd.n2252 gnd.n2200 585
R1886 gnd.n2251 gnd.n2250 585
R1887 gnd.n1276 gnd.n1274 585
R1888 gnd.n3143 gnd.n1274 585
R1889 gnd.n2333 gnd.n1272 585
R1890 gnd.n4667 gnd.n1272 585
R1891 gnd.n2830 gnd.n2829 585
R1892 gnd.n2831 gnd.n2830 585
R1893 gnd.n2332 gnd.n1263 585
R1894 gnd.n4673 gnd.n1263 585
R1895 gnd.n2795 gnd.n2794 585
R1896 gnd.n2794 gnd.n2793 585
R1897 gnd.n2335 gnd.n1252 585
R1898 gnd.n4679 gnd.n1252 585
R1899 gnd.n2783 gnd.n2782 585
R1900 gnd.n2784 gnd.n2783 585
R1901 gnd.n2339 gnd.n1241 585
R1902 gnd.n4685 gnd.n1241 585
R1903 gnd.n2778 gnd.n2777 585
R1904 gnd.n2777 gnd.n2776 585
R1905 gnd.n2341 gnd.n1231 585
R1906 gnd.n4691 gnd.n1231 585
R1907 gnd.n2711 gnd.n2710 585
R1908 gnd.n2710 gnd.n2709 585
R1909 gnd.n2361 gnd.n1220 585
R1910 gnd.n4697 gnd.n1220 585
R1911 gnd.n2715 gnd.n2360 585
R1912 gnd.n2697 gnd.n2360 585
R1913 gnd.n2716 gnd.n1210 585
R1914 gnd.n4703 gnd.n1210 585
R1915 gnd.n2717 gnd.n2359 585
R1916 gnd.n2692 gnd.n2359 585
R1917 gnd.n2356 gnd.n1199 585
R1918 gnd.n4709 gnd.n1199 585
R1919 gnd.n2722 gnd.n2721 585
R1920 gnd.n2723 gnd.n2722 585
R1921 gnd.n2355 gnd.n1189 585
R1922 gnd.n4715 gnd.n1189 585
R1923 gnd.n2683 gnd.n2682 585
R1924 gnd.n2684 gnd.n2683 585
R1925 gnd.n2368 gnd.n1178 585
R1926 gnd.n4721 gnd.n1178 585
R1927 gnd.n2678 gnd.n2677 585
R1928 gnd.n2677 gnd.n2676 585
R1929 gnd.n2370 gnd.n1168 585
R1930 gnd.n4727 gnd.n1168 585
R1931 gnd.n2666 gnd.n2665 585
R1932 gnd.n2667 gnd.n2666 585
R1933 gnd.n2375 gnd.n1158 585
R1934 gnd.n4733 gnd.n1158 585
R1935 gnd.n2661 gnd.n2660 585
R1936 gnd.n2660 gnd.n2659 585
R1937 gnd.n2377 gnd.n1148 585
R1938 gnd.n4739 gnd.n1148 585
R1939 gnd.n2629 gnd.n2628 585
R1940 gnd.n2628 gnd.n2627 585
R1941 gnd.n2633 gnd.n1140 585
R1942 gnd.n4746 gnd.n1140 585
R1943 gnd.n2635 gnd.n2634 585
R1944 gnd.n2636 gnd.n2635 585
R1945 gnd.n2419 gnd.n1130 585
R1946 gnd.n4752 gnd.n1130 585
R1947 gnd.n2644 gnd.n2643 585
R1948 gnd.n2643 gnd.n2642 585
R1949 gnd.n2645 gnd.n1121 585
R1950 gnd.n4758 gnd.n1121 585
R1951 gnd.n2647 gnd.n2646 585
R1952 gnd.n2648 gnd.n2647 585
R1953 gnd.n2415 gnd.n1111 585
R1954 gnd.n4764 gnd.n1111 585
R1955 gnd.n2591 gnd.n2590 585
R1956 gnd.n2592 gnd.n2591 585
R1957 gnd.n2460 gnd.n1100 585
R1958 gnd.n4770 gnd.n1100 585
R1959 gnd.n2585 gnd.n2584 585
R1960 gnd.n2584 gnd.n1098 585
R1961 gnd.n2583 gnd.n1089 585
R1962 gnd.n4776 gnd.n1089 585
R1963 gnd.n2582 gnd.n2581 585
R1964 gnd.n2581 gnd.n1080 585
R1965 gnd.n2462 gnd.n1079 585
R1966 gnd.n4782 gnd.n1079 585
R1967 gnd.n2577 gnd.n2576 585
R1968 gnd.n2576 gnd.n1070 585
R1969 gnd.n2575 gnd.n1069 585
R1970 gnd.n4788 gnd.n1069 585
R1971 gnd.n2574 gnd.n2573 585
R1972 gnd.n2573 gnd.n1067 585
R1973 gnd.n2464 gnd.n1059 585
R1974 gnd.n4794 gnd.n1059 585
R1975 gnd.n2569 gnd.n2568 585
R1976 gnd.n2568 gnd.n1057 585
R1977 gnd.n2567 gnd.n1049 585
R1978 gnd.n4800 gnd.n1049 585
R1979 gnd.n2566 gnd.n2565 585
R1980 gnd.n2565 gnd.n1040 585
R1981 gnd.n2466 gnd.n1039 585
R1982 gnd.n4806 gnd.n1039 585
R1983 gnd.n2561 gnd.n2560 585
R1984 gnd.n2560 gnd.n1029 585
R1985 gnd.n2559 gnd.n1028 585
R1986 gnd.n4812 gnd.n1028 585
R1987 gnd.n2558 gnd.n2557 585
R1988 gnd.n2557 gnd.n1017 585
R1989 gnd.n2468 gnd.n1016 585
R1990 gnd.n4818 gnd.n1016 585
R1991 gnd.n2553 gnd.n2552 585
R1992 gnd.n2552 gnd.n1015 585
R1993 gnd.n2551 gnd.n2470 585
R1994 gnd.n2551 gnd.n2550 585
R1995 gnd.n2495 gnd.n2471 585
R1996 gnd.n2471 gnd.n961 585
R1997 gnd.n7438 gnd.n107 585
R1998 gnd.n7534 gnd.n107 585
R1999 gnd.n7439 gnd.n7369 585
R2000 gnd.n7369 gnd.n104 585
R2001 gnd.n7440 gnd.n187 585
R2002 gnd.n7454 gnd.n187 585
R2003 gnd.n198 gnd.n196 585
R2004 gnd.n196 gnd.n185 585
R2005 gnd.n7445 gnd.n7444 585
R2006 gnd.n7446 gnd.n7445 585
R2007 gnd.n197 gnd.n195 585
R2008 gnd.n195 gnd.n193 585
R2009 gnd.n7365 gnd.n7364 585
R2010 gnd.n7364 gnd.n7363 585
R2011 gnd.n201 gnd.n200 585
R2012 gnd.n211 gnd.n201 585
R2013 gnd.n7354 gnd.n7353 585
R2014 gnd.n7355 gnd.n7354 585
R2015 gnd.n213 gnd.n212 585
R2016 gnd.n212 gnd.n208 585
R2017 gnd.n7349 gnd.n7348 585
R2018 gnd.n7348 gnd.n7347 585
R2019 gnd.n216 gnd.n215 585
R2020 gnd.n218 gnd.n216 585
R2021 gnd.n7338 gnd.n7337 585
R2022 gnd.n7339 gnd.n7338 585
R2023 gnd.n228 gnd.n227 585
R2024 gnd.n227 gnd.n225 585
R2025 gnd.n7333 gnd.n7332 585
R2026 gnd.n7332 gnd.n7331 585
R2027 gnd.n231 gnd.n230 585
R2028 gnd.n241 gnd.n231 585
R2029 gnd.n7322 gnd.n7321 585
R2030 gnd.n7323 gnd.n7322 585
R2031 gnd.n243 gnd.n242 585
R2032 gnd.n242 gnd.n238 585
R2033 gnd.n7317 gnd.n7316 585
R2034 gnd.n7316 gnd.n7315 585
R2035 gnd.n246 gnd.n245 585
R2036 gnd.n248 gnd.n246 585
R2037 gnd.n7306 gnd.n7305 585
R2038 gnd.n7307 gnd.n7306 585
R2039 gnd.n259 gnd.n258 585
R2040 gnd.n7260 gnd.n258 585
R2041 gnd.n7301 gnd.n7300 585
R2042 gnd.n7300 gnd.n7299 585
R2043 gnd.n262 gnd.n261 585
R2044 gnd.n7265 gnd.n262 585
R2045 gnd.n7278 gnd.n7277 585
R2046 gnd.n7277 gnd.n7276 585
R2047 gnd.n7279 gnd.n293 585
R2048 gnd.n7271 gnd.n293 585
R2049 gnd.n319 gnd.n290 585
R2050 gnd.n320 gnd.n319 585
R2051 gnd.n7284 gnd.n289 585
R2052 gnd.n7205 gnd.n289 585
R2053 gnd.n7285 gnd.n288 585
R2054 gnd.n7200 gnd.n288 585
R2055 gnd.n7286 gnd.n287 585
R2056 gnd.n314 gnd.n287 585
R2057 gnd.n284 gnd.n282 585
R2058 gnd.n7192 gnd.n282 585
R2059 gnd.n7291 gnd.n7290 585
R2060 gnd.n7292 gnd.n7291 585
R2061 gnd.n283 gnd.n281 585
R2062 gnd.n4349 gnd.n281 585
R2063 gnd.n4390 gnd.n4388 585
R2064 gnd.n4388 gnd.n4387 585
R2065 gnd.n4391 gnd.n1526 585
R2066 gnd.n1538 gnd.n1526 585
R2067 gnd.n4392 gnd.n1525 585
R2068 gnd.n4379 gnd.n1525 585
R2069 gnd.n4360 gnd.n1523 585
R2070 gnd.n4361 gnd.n4360 585
R2071 gnd.n4396 gnd.n1522 585
R2072 gnd.n1546 gnd.n1522 585
R2073 gnd.n4397 gnd.n1521 585
R2074 gnd.n4326 gnd.n1521 585
R2075 gnd.n4398 gnd.n1520 585
R2076 gnd.n1573 gnd.n1520 585
R2077 gnd.n4315 gnd.n1518 585
R2078 gnd.n4316 gnd.n4315 585
R2079 gnd.n4402 gnd.n1517 585
R2080 gnd.n4303 gnd.n1517 585
R2081 gnd.n4403 gnd.n1516 585
R2082 gnd.n1580 gnd.n1516 585
R2083 gnd.n4404 gnd.n1515 585
R2084 gnd.n4289 gnd.n1515 585
R2085 gnd.n1600 gnd.n1513 585
R2086 gnd.n1601 gnd.n1600 585
R2087 gnd.n4408 gnd.n1512 585
R2088 gnd.n4279 gnd.n1512 585
R2089 gnd.n4409 gnd.n1511 585
R2090 gnd.n4267 gnd.n1511 585
R2091 gnd.n4410 gnd.n1510 585
R2092 gnd.n1671 gnd.n1510 585
R2093 gnd.n1618 gnd.n1508 585
R2094 gnd.n4258 gnd.n1618 585
R2095 gnd.n4414 gnd.n1507 585
R2096 gnd.n1628 gnd.n1507 585
R2097 gnd.n4415 gnd.n1506 585
R2098 gnd.n4248 gnd.n1506 585
R2099 gnd.n4416 gnd.n1505 585
R2100 gnd.n4236 gnd.n1505 585
R2101 gnd.n1502 gnd.n1501 585
R2102 gnd.n1647 gnd.n1501 585
R2103 gnd.n4421 gnd.n4420 585
R2104 gnd.n4422 gnd.n4421 585
R2105 gnd.n1722 gnd.n1500 585
R2106 gnd.n1727 gnd.n1726 585
R2107 gnd.n1729 gnd.n1728 585
R2108 gnd.n1732 gnd.n1731 585
R2109 gnd.n1730 gnd.n1715 585
R2110 gnd.n1746 gnd.n1745 585
R2111 gnd.n1748 gnd.n1747 585
R2112 gnd.n1751 gnd.n1750 585
R2113 gnd.n1749 gnd.n1708 585
R2114 gnd.n1765 gnd.n1764 585
R2115 gnd.n1767 gnd.n1766 585
R2116 gnd.n1770 gnd.n1769 585
R2117 gnd.n1768 gnd.n1701 585
R2118 gnd.n1783 gnd.n1782 585
R2119 gnd.n1785 gnd.n1784 585
R2120 gnd.n1694 gnd.n1693 585
R2121 gnd.n1798 gnd.n1695 585
R2122 gnd.n1799 gnd.n1690 585
R2123 gnd.n1800 gnd.n1445 585
R2124 gnd.n4498 gnd.n1445 585
R2125 gnd.n7409 gnd.n103 585
R2126 gnd.n7410 gnd.n7407 585
R2127 gnd.n7411 gnd.n7403 585
R2128 gnd.n7401 gnd.n7399 585
R2129 gnd.n7415 gnd.n7398 585
R2130 gnd.n7416 gnd.n7396 585
R2131 gnd.n7417 gnd.n7395 585
R2132 gnd.n7393 gnd.n7391 585
R2133 gnd.n7421 gnd.n7390 585
R2134 gnd.n7422 gnd.n7388 585
R2135 gnd.n7423 gnd.n7387 585
R2136 gnd.n7385 gnd.n7383 585
R2137 gnd.n7427 gnd.n7382 585
R2138 gnd.n7428 gnd.n7380 585
R2139 gnd.n7429 gnd.n7379 585
R2140 gnd.n7377 gnd.n7375 585
R2141 gnd.n7433 gnd.n7374 585
R2142 gnd.n7434 gnd.n7372 585
R2143 gnd.n7435 gnd.n7371 585
R2144 gnd.n7371 gnd.n106 585
R2145 gnd.n7536 gnd.n7535 585
R2146 gnd.n7535 gnd.n7534 585
R2147 gnd.n7537 gnd.n101 585
R2148 gnd.n104 gnd.n101 585
R2149 gnd.n7538 gnd.n100 585
R2150 gnd.n7454 gnd.n100 585
R2151 gnd.n184 gnd.n98 585
R2152 gnd.n185 gnd.n184 585
R2153 gnd.n7542 gnd.n97 585
R2154 gnd.n7446 gnd.n97 585
R2155 gnd.n7543 gnd.n96 585
R2156 gnd.n193 gnd.n96 585
R2157 gnd.n7544 gnd.n95 585
R2158 gnd.n7363 gnd.n95 585
R2159 gnd.n210 gnd.n93 585
R2160 gnd.n211 gnd.n210 585
R2161 gnd.n7548 gnd.n92 585
R2162 gnd.n7355 gnd.n92 585
R2163 gnd.n7549 gnd.n91 585
R2164 gnd.n208 gnd.n91 585
R2165 gnd.n7550 gnd.n90 585
R2166 gnd.n7347 gnd.n90 585
R2167 gnd.n217 gnd.n88 585
R2168 gnd.n218 gnd.n217 585
R2169 gnd.n7554 gnd.n87 585
R2170 gnd.n7339 gnd.n87 585
R2171 gnd.n7555 gnd.n86 585
R2172 gnd.n225 gnd.n86 585
R2173 gnd.n7556 gnd.n85 585
R2174 gnd.n7331 gnd.n85 585
R2175 gnd.n240 gnd.n83 585
R2176 gnd.n241 gnd.n240 585
R2177 gnd.n7560 gnd.n82 585
R2178 gnd.n7323 gnd.n82 585
R2179 gnd.n7561 gnd.n81 585
R2180 gnd.n238 gnd.n81 585
R2181 gnd.n7562 gnd.n80 585
R2182 gnd.n7315 gnd.n80 585
R2183 gnd.n247 gnd.n78 585
R2184 gnd.n248 gnd.n247 585
R2185 gnd.n7566 gnd.n77 585
R2186 gnd.n7307 gnd.n77 585
R2187 gnd.n7567 gnd.n76 585
R2188 gnd.n7260 gnd.n76 585
R2189 gnd.n7568 gnd.n75 585
R2190 gnd.n7299 gnd.n75 585
R2191 gnd.n7264 gnd.n73 585
R2192 gnd.n7265 gnd.n7264 585
R2193 gnd.n7572 gnd.n72 585
R2194 gnd.n7276 gnd.n72 585
R2195 gnd.n7573 gnd.n71 585
R2196 gnd.n7271 gnd.n71 585
R2197 gnd.n7574 gnd.n70 585
R2198 gnd.n320 gnd.n70 585
R2199 gnd.n303 gnd.n69 585
R2200 gnd.n7205 gnd.n303 585
R2201 gnd.n7199 gnd.n7198 585
R2202 gnd.n7200 gnd.n7199 585
R2203 gnd.n309 gnd.n308 585
R2204 gnd.n314 gnd.n308 585
R2205 gnd.n7194 gnd.n7193 585
R2206 gnd.n7193 gnd.n7192 585
R2207 gnd.n311 gnd.n280 585
R2208 gnd.n7292 gnd.n280 585
R2209 gnd.n4352 gnd.n4350 585
R2210 gnd.n4350 gnd.n4349 585
R2211 gnd.n4353 gnd.n1528 585
R2212 gnd.n4387 gnd.n1528 585
R2213 gnd.n4354 gnd.n1553 585
R2214 gnd.n1553 gnd.n1538 585
R2215 gnd.n1550 gnd.n1537 585
R2216 gnd.n4379 gnd.n1537 585
R2217 gnd.n4359 gnd.n4358 585
R2218 gnd.n4361 gnd.n4359 585
R2219 gnd.n1549 gnd.n1548 585
R2220 gnd.n1548 gnd.n1546 585
R2221 gnd.n4296 gnd.n1562 585
R2222 gnd.n4326 gnd.n1562 585
R2223 gnd.n4297 gnd.n4295 585
R2224 gnd.n4295 gnd.n1573 585
R2225 gnd.n1584 gnd.n1572 585
R2226 gnd.n4316 gnd.n1572 585
R2227 gnd.n4302 gnd.n4301 585
R2228 gnd.n4303 gnd.n4302 585
R2229 gnd.n1583 gnd.n1582 585
R2230 gnd.n1582 gnd.n1580 585
R2231 gnd.n4291 gnd.n4290 585
R2232 gnd.n4290 gnd.n4289 585
R2233 gnd.n1587 gnd.n1586 585
R2234 gnd.n1601 gnd.n1587 585
R2235 gnd.n1611 gnd.n1599 585
R2236 gnd.n4279 gnd.n1599 585
R2237 gnd.n4266 gnd.n4265 585
R2238 gnd.n4267 gnd.n4266 585
R2239 gnd.n1610 gnd.n1609 585
R2240 gnd.n1671 gnd.n1609 585
R2241 gnd.n4260 gnd.n4259 585
R2242 gnd.n4259 gnd.n4258 585
R2243 gnd.n1614 gnd.n1613 585
R2244 gnd.n1628 gnd.n1614 585
R2245 gnd.n1682 gnd.n1627 585
R2246 gnd.n4248 gnd.n1627 585
R2247 gnd.n4235 gnd.n4234 585
R2248 gnd.n4236 gnd.n4235 585
R2249 gnd.n1681 gnd.n1680 585
R2250 gnd.n1680 gnd.n1647 585
R2251 gnd.n4229 gnd.n1498 585
R2252 gnd.n4422 gnd.n1498 585
R2253 gnd.n6312 gnd.n6311 585
R2254 gnd.n6311 gnd.n6310 585
R2255 gnd.n6313 gnd.n924 585
R2256 gnd.n6220 gnd.n924 585
R2257 gnd.n6315 gnd.n6314 585
R2258 gnd.n6316 gnd.n6315 585
R2259 gnd.n925 gnd.n923 585
R2260 gnd.n923 gnd.n919 585
R2261 gnd.n906 gnd.n905 585
R2262 gnd.n910 gnd.n906 585
R2263 gnd.n6326 gnd.n6325 585
R2264 gnd.n6325 gnd.n6324 585
R2265 gnd.n6327 gnd.n900 585
R2266 gnd.n6209 gnd.n900 585
R2267 gnd.n6329 gnd.n6328 585
R2268 gnd.n6330 gnd.n6329 585
R2269 gnd.n901 gnd.n899 585
R2270 gnd.n6203 gnd.n899 585
R2271 gnd.n6184 gnd.n5009 585
R2272 gnd.n5009 gnd.n5008 585
R2273 gnd.n6186 gnd.n6185 585
R2274 gnd.n6187 gnd.n6186 585
R2275 gnd.n5010 gnd.n5007 585
R2276 gnd.n5007 gnd.n5003 585
R2277 gnd.n5891 gnd.n5890 585
R2278 gnd.n5890 gnd.n5889 585
R2279 gnd.n5017 gnd.n5016 585
R2280 gnd.n5026 gnd.n5017 585
R2281 gnd.n5880 gnd.n5879 585
R2282 gnd.n5879 gnd.n5878 585
R2283 gnd.n5024 gnd.n5023 585
R2284 gnd.n5866 gnd.n5024 585
R2285 gnd.n5841 gnd.n5041 585
R2286 gnd.n5834 gnd.n5041 585
R2287 gnd.n5843 gnd.n5842 585
R2288 gnd.n5844 gnd.n5843 585
R2289 gnd.n5042 gnd.n5040 585
R2290 gnd.n5050 gnd.n5040 585
R2291 gnd.n5817 gnd.n5062 585
R2292 gnd.n5062 gnd.n5049 585
R2293 gnd.n5819 gnd.n5818 585
R2294 gnd.n5820 gnd.n5819 585
R2295 gnd.n5063 gnd.n5061 585
R2296 gnd.n5061 gnd.n5057 585
R2297 gnd.n5805 gnd.n5804 585
R2298 gnd.n5804 gnd.n5803 585
R2299 gnd.n5068 gnd.n5067 585
R2300 gnd.n5072 gnd.n5068 585
R2301 gnd.n5789 gnd.n5788 585
R2302 gnd.n5790 gnd.n5789 585
R2303 gnd.n5082 gnd.n5081 585
R2304 gnd.n5780 gnd.n5081 585
R2305 gnd.n5754 gnd.n5097 585
R2306 gnd.n5097 gnd.n5089 585
R2307 gnd.n5756 gnd.n5755 585
R2308 gnd.n5757 gnd.n5756 585
R2309 gnd.n5098 gnd.n5096 585
R2310 gnd.n5102 gnd.n5096 585
R2311 gnd.n5735 gnd.n5734 585
R2312 gnd.n5736 gnd.n5735 585
R2313 gnd.n5114 gnd.n5113 585
R2314 gnd.n5113 gnd.n5109 585
R2315 gnd.n5725 gnd.n5724 585
R2316 gnd.n5726 gnd.n5725 585
R2317 gnd.n5122 gnd.n5121 585
R2318 gnd.n5126 gnd.n5121 585
R2319 gnd.n5703 gnd.n5138 585
R2320 gnd.n5482 gnd.n5138 585
R2321 gnd.n5705 gnd.n5704 585
R2322 gnd.n5706 gnd.n5705 585
R2323 gnd.n5139 gnd.n5137 585
R2324 gnd.n5137 gnd.n5133 585
R2325 gnd.n5694 gnd.n5693 585
R2326 gnd.n5695 gnd.n5694 585
R2327 gnd.n5147 gnd.n5146 585
R2328 gnd.n5152 gnd.n5146 585
R2329 gnd.n5672 gnd.n5164 585
R2330 gnd.n5164 gnd.n5151 585
R2331 gnd.n5674 gnd.n5673 585
R2332 gnd.n5675 gnd.n5674 585
R2333 gnd.n5165 gnd.n5163 585
R2334 gnd.n5163 gnd.n5159 585
R2335 gnd.n5663 gnd.n5662 585
R2336 gnd.n5664 gnd.n5663 585
R2337 gnd.n5173 gnd.n5172 585
R2338 gnd.n5547 gnd.n5172 585
R2339 gnd.n5641 gnd.n5189 585
R2340 gnd.n5189 gnd.n5177 585
R2341 gnd.n5643 gnd.n5642 585
R2342 gnd.n5644 gnd.n5643 585
R2343 gnd.n5190 gnd.n5188 585
R2344 gnd.n5188 gnd.n5184 585
R2345 gnd.n5632 gnd.n5631 585
R2346 gnd.n5633 gnd.n5632 585
R2347 gnd.n5197 gnd.n5196 585
R2348 gnd.n5202 gnd.n5196 585
R2349 gnd.n5610 gnd.n5215 585
R2350 gnd.n5215 gnd.n5201 585
R2351 gnd.n5612 gnd.n5611 585
R2352 gnd.n5613 gnd.n5612 585
R2353 gnd.n5216 gnd.n5214 585
R2354 gnd.n5214 gnd.n5210 585
R2355 gnd.n5601 gnd.n5600 585
R2356 gnd.n5602 gnd.n5601 585
R2357 gnd.n5223 gnd.n5222 585
R2358 gnd.n5227 gnd.n5222 585
R2359 gnd.n5578 gnd.n5244 585
R2360 gnd.n5244 gnd.n5226 585
R2361 gnd.n5580 gnd.n5579 585
R2362 gnd.n5581 gnd.n5580 585
R2363 gnd.n5245 gnd.n5243 585
R2364 gnd.n5243 gnd.n5234 585
R2365 gnd.n5573 gnd.n5572 585
R2366 gnd.n5572 gnd.n5571 585
R2367 gnd.n5292 gnd.n5291 585
R2368 gnd.n5293 gnd.n5292 585
R2369 gnd.n5446 gnd.n5445 585
R2370 gnd.n5447 gnd.n5446 585
R2371 gnd.n5302 gnd.n5301 585
R2372 gnd.n5301 gnd.n5300 585
R2373 gnd.n5441 gnd.n5440 585
R2374 gnd.n5440 gnd.n5439 585
R2375 gnd.n5305 gnd.n5304 585
R2376 gnd.n5306 gnd.n5305 585
R2377 gnd.n5430 gnd.n5429 585
R2378 gnd.n5431 gnd.n5430 585
R2379 gnd.n5313 gnd.n5312 585
R2380 gnd.n5422 gnd.n5312 585
R2381 gnd.n5425 gnd.n5424 585
R2382 gnd.n5424 gnd.n5423 585
R2383 gnd.n5316 gnd.n5315 585
R2384 gnd.n5317 gnd.n5316 585
R2385 gnd.n5411 gnd.n5410 585
R2386 gnd.n5409 gnd.n5335 585
R2387 gnd.n5408 gnd.n5334 585
R2388 gnd.n5413 gnd.n5334 585
R2389 gnd.n5407 gnd.n5406 585
R2390 gnd.n5405 gnd.n5404 585
R2391 gnd.n5403 gnd.n5402 585
R2392 gnd.n5401 gnd.n5400 585
R2393 gnd.n5399 gnd.n5398 585
R2394 gnd.n5397 gnd.n5396 585
R2395 gnd.n5395 gnd.n5394 585
R2396 gnd.n5393 gnd.n5392 585
R2397 gnd.n5391 gnd.n5390 585
R2398 gnd.n5389 gnd.n5388 585
R2399 gnd.n5387 gnd.n5386 585
R2400 gnd.n5385 gnd.n5384 585
R2401 gnd.n5383 gnd.n5382 585
R2402 gnd.n5381 gnd.n5380 585
R2403 gnd.n5379 gnd.n5378 585
R2404 gnd.n5377 gnd.n5376 585
R2405 gnd.n5375 gnd.n5374 585
R2406 gnd.n5373 gnd.n5372 585
R2407 gnd.n5371 gnd.n5370 585
R2408 gnd.n5369 gnd.n5368 585
R2409 gnd.n5367 gnd.n5366 585
R2410 gnd.n5365 gnd.n5364 585
R2411 gnd.n5322 gnd.n5321 585
R2412 gnd.n5416 gnd.n5415 585
R2413 gnd.n6228 gnd.n6227 585
R2414 gnd.n6229 gnd.n4985 585
R2415 gnd.n6231 gnd.n6230 585
R2416 gnd.n6233 gnd.n4984 585
R2417 gnd.n6235 gnd.n6234 585
R2418 gnd.n6236 gnd.n4975 585
R2419 gnd.n6238 gnd.n6237 585
R2420 gnd.n6240 gnd.n4973 585
R2421 gnd.n6242 gnd.n6241 585
R2422 gnd.n6243 gnd.n4968 585
R2423 gnd.n6245 gnd.n6244 585
R2424 gnd.n6247 gnd.n4966 585
R2425 gnd.n6249 gnd.n6248 585
R2426 gnd.n6250 gnd.n4961 585
R2427 gnd.n6252 gnd.n6251 585
R2428 gnd.n6254 gnd.n4959 585
R2429 gnd.n6256 gnd.n6255 585
R2430 gnd.n6257 gnd.n4954 585
R2431 gnd.n6259 gnd.n6258 585
R2432 gnd.n6261 gnd.n4952 585
R2433 gnd.n6263 gnd.n6262 585
R2434 gnd.n6264 gnd.n4947 585
R2435 gnd.n6266 gnd.n6265 585
R2436 gnd.n6268 gnd.n4945 585
R2437 gnd.n6270 gnd.n6269 585
R2438 gnd.n6271 gnd.n4943 585
R2439 gnd.n6272 gnd.n929 585
R2440 gnd.n4906 gnd.n929 585
R2441 gnd.n6223 gnd.n931 585
R2442 gnd.n6310 gnd.n931 585
R2443 gnd.n6222 gnd.n6221 585
R2444 gnd.n6221 gnd.n6220 585
R2445 gnd.n6219 gnd.n921 585
R2446 gnd.n6316 gnd.n921 585
R2447 gnd.n6213 gnd.n4990 585
R2448 gnd.n6213 gnd.n919 585
R2449 gnd.n6215 gnd.n6214 585
R2450 gnd.n6214 gnd.n910 585
R2451 gnd.n6212 gnd.n908 585
R2452 gnd.n6324 gnd.n908 585
R2453 gnd.n6211 gnd.n6210 585
R2454 gnd.n6210 gnd.n6209 585
R2455 gnd.n4992 gnd.n897 585
R2456 gnd.n6330 gnd.n897 585
R2457 gnd.n6205 gnd.n6204 585
R2458 gnd.n6204 gnd.n6203 585
R2459 gnd.n4995 gnd.n4994 585
R2460 gnd.n5008 gnd.n4995 585
R2461 gnd.n5855 gnd.n5005 585
R2462 gnd.n6187 gnd.n5005 585
R2463 gnd.n5857 gnd.n5856 585
R2464 gnd.n5856 gnd.n5003 585
R2465 gnd.n5858 gnd.n5019 585
R2466 gnd.n5889 gnd.n5019 585
R2467 gnd.n5860 gnd.n5859 585
R2468 gnd.n5859 gnd.n5026 585
R2469 gnd.n5861 gnd.n5025 585
R2470 gnd.n5878 gnd.n5025 585
R2471 gnd.n5863 gnd.n5862 585
R2472 gnd.n5866 gnd.n5863 585
R2473 gnd.n5035 gnd.n5034 585
R2474 gnd.n5834 gnd.n5034 585
R2475 gnd.n5846 gnd.n5845 585
R2476 gnd.n5845 gnd.n5844 585
R2477 gnd.n5038 gnd.n5037 585
R2478 gnd.n5050 gnd.n5038 585
R2479 gnd.n5770 gnd.n5769 585
R2480 gnd.n5769 gnd.n5049 585
R2481 gnd.n5771 gnd.n5059 585
R2482 gnd.n5820 gnd.n5059 585
R2483 gnd.n5773 gnd.n5772 585
R2484 gnd.n5772 gnd.n5057 585
R2485 gnd.n5774 gnd.n5069 585
R2486 gnd.n5803 gnd.n5069 585
R2487 gnd.n5776 gnd.n5775 585
R2488 gnd.n5775 gnd.n5072 585
R2489 gnd.n5777 gnd.n5079 585
R2490 gnd.n5790 gnd.n5079 585
R2491 gnd.n5779 gnd.n5778 585
R2492 gnd.n5780 gnd.n5779 585
R2493 gnd.n5091 gnd.n5090 585
R2494 gnd.n5090 gnd.n5089 585
R2495 gnd.n5759 gnd.n5758 585
R2496 gnd.n5758 gnd.n5757 585
R2497 gnd.n5094 gnd.n5093 585
R2498 gnd.n5102 gnd.n5094 585
R2499 gnd.n5474 gnd.n5111 585
R2500 gnd.n5736 gnd.n5111 585
R2501 gnd.n5477 gnd.n5476 585
R2502 gnd.n5476 gnd.n5109 585
R2503 gnd.n5478 gnd.n5120 585
R2504 gnd.n5726 gnd.n5120 585
R2505 gnd.n5481 gnd.n5480 585
R2506 gnd.n5481 gnd.n5126 585
R2507 gnd.n5484 gnd.n5483 585
R2508 gnd.n5483 gnd.n5482 585
R2509 gnd.n5485 gnd.n5135 585
R2510 gnd.n5706 gnd.n5135 585
R2511 gnd.n5473 gnd.n5472 585
R2512 gnd.n5472 gnd.n5133 585
R2513 gnd.n5537 gnd.n5145 585
R2514 gnd.n5695 gnd.n5145 585
R2515 gnd.n5539 gnd.n5538 585
R2516 gnd.n5539 gnd.n5152 585
R2517 gnd.n5541 gnd.n5540 585
R2518 gnd.n5540 gnd.n5151 585
R2519 gnd.n5542 gnd.n5161 585
R2520 gnd.n5675 gnd.n5161 585
R2521 gnd.n5544 gnd.n5543 585
R2522 gnd.n5543 gnd.n5159 585
R2523 gnd.n5545 gnd.n5171 585
R2524 gnd.n5664 gnd.n5171 585
R2525 gnd.n5548 gnd.n5546 585
R2526 gnd.n5548 gnd.n5547 585
R2527 gnd.n5550 gnd.n5549 585
R2528 gnd.n5549 gnd.n5177 585
R2529 gnd.n5551 gnd.n5186 585
R2530 gnd.n5644 gnd.n5186 585
R2531 gnd.n5553 gnd.n5552 585
R2532 gnd.n5552 gnd.n5184 585
R2533 gnd.n5554 gnd.n5195 585
R2534 gnd.n5633 gnd.n5195 585
R2535 gnd.n5556 gnd.n5555 585
R2536 gnd.n5556 gnd.n5202 585
R2537 gnd.n5558 gnd.n5557 585
R2538 gnd.n5557 gnd.n5201 585
R2539 gnd.n5559 gnd.n5212 585
R2540 gnd.n5613 gnd.n5212 585
R2541 gnd.n5561 gnd.n5560 585
R2542 gnd.n5560 gnd.n5210 585
R2543 gnd.n5562 gnd.n5221 585
R2544 gnd.n5602 gnd.n5221 585
R2545 gnd.n5564 gnd.n5563 585
R2546 gnd.n5564 gnd.n5227 585
R2547 gnd.n5566 gnd.n5565 585
R2548 gnd.n5565 gnd.n5226 585
R2549 gnd.n5567 gnd.n5242 585
R2550 gnd.n5581 gnd.n5242 585
R2551 gnd.n5568 gnd.n5295 585
R2552 gnd.n5295 gnd.n5234 585
R2553 gnd.n5570 gnd.n5569 585
R2554 gnd.n5571 gnd.n5570 585
R2555 gnd.n5296 gnd.n5294 585
R2556 gnd.n5294 gnd.n5293 585
R2557 gnd.n5449 gnd.n5448 585
R2558 gnd.n5448 gnd.n5447 585
R2559 gnd.n5299 gnd.n5298 585
R2560 gnd.n5300 gnd.n5299 585
R2561 gnd.n5438 gnd.n5437 585
R2562 gnd.n5439 gnd.n5438 585
R2563 gnd.n5308 gnd.n5307 585
R2564 gnd.n5307 gnd.n5306 585
R2565 gnd.n5433 gnd.n5432 585
R2566 gnd.n5432 gnd.n5431 585
R2567 gnd.n5311 gnd.n5310 585
R2568 gnd.n5422 gnd.n5311 585
R2569 gnd.n5421 gnd.n5420 585
R2570 gnd.n5423 gnd.n5421 585
R2571 gnd.n5319 gnd.n5318 585
R2572 gnd.n5318 gnd.n5317 585
R2573 gnd.n6308 gnd.n6307 585
R2574 gnd.n6309 gnd.n6308 585
R2575 gnd.n4909 gnd.n4907 585
R2576 gnd.n4907 gnd.n930 585
R2577 gnd.n918 gnd.n917 585
R2578 gnd.n922 gnd.n918 585
R2579 gnd.n6319 gnd.n6318 585
R2580 gnd.n6318 gnd.n6317 585
R2581 gnd.n6320 gnd.n912 585
R2582 gnd.n6172 gnd.n912 585
R2583 gnd.n6322 gnd.n6321 585
R2584 gnd.n6323 gnd.n6322 585
R2585 gnd.n913 gnd.n911 585
R2586 gnd.n911 gnd.n907 585
R2587 gnd.n6198 gnd.n6197 585
R2588 gnd.n6197 gnd.n898 585
R2589 gnd.n6199 gnd.n4998 585
R2590 gnd.n4998 gnd.n896 585
R2591 gnd.n6201 gnd.n6200 585
R2592 gnd.n6202 gnd.n6201 585
R2593 gnd.n4999 gnd.n4997 585
R2594 gnd.n5006 gnd.n4997 585
R2595 gnd.n6190 gnd.n6189 585
R2596 gnd.n6189 gnd.n6188 585
R2597 gnd.n5002 gnd.n5001 585
R2598 gnd.n5888 gnd.n5002 585
R2599 gnd.n5874 gnd.n5028 585
R2600 gnd.n5028 gnd.n5018 585
R2601 gnd.n5876 gnd.n5875 585
R2602 gnd.n5877 gnd.n5876 585
R2603 gnd.n5029 gnd.n5027 585
R2604 gnd.n5865 gnd.n5027 585
R2605 gnd.n5869 gnd.n5868 585
R2606 gnd.n5868 gnd.n5867 585
R2607 gnd.n5032 gnd.n5031 585
R2608 gnd.n5835 gnd.n5032 585
R2609 gnd.n5828 gnd.n5052 585
R2610 gnd.n5052 gnd.n5039 585
R2611 gnd.n5830 gnd.n5829 585
R2612 gnd.n5831 gnd.n5830 585
R2613 gnd.n5053 gnd.n5051 585
R2614 gnd.n5060 gnd.n5051 585
R2615 gnd.n5823 gnd.n5822 585
R2616 gnd.n5822 gnd.n5821 585
R2617 gnd.n5056 gnd.n5055 585
R2618 gnd.n5802 gnd.n5056 585
R2619 gnd.n5798 gnd.n5797 585
R2620 gnd.n5799 gnd.n5798 585
R2621 gnd.n5074 gnd.n5073 585
R2622 gnd.n5080 gnd.n5073 585
R2623 gnd.n5793 gnd.n5792 585
R2624 gnd.n5792 gnd.n5791 585
R2625 gnd.n5077 gnd.n5076 585
R2626 gnd.n5781 gnd.n5077 585
R2627 gnd.n5744 gnd.n5104 585
R2628 gnd.n5104 gnd.n5095 585
R2629 gnd.n5746 gnd.n5745 585
R2630 gnd.n5747 gnd.n5746 585
R2631 gnd.n5105 gnd.n5103 585
R2632 gnd.n5112 gnd.n5103 585
R2633 gnd.n5739 gnd.n5738 585
R2634 gnd.n5738 gnd.n5737 585
R2635 gnd.n5108 gnd.n5107 585
R2636 gnd.n5727 gnd.n5108 585
R2637 gnd.n5714 gnd.n5128 585
R2638 gnd.n5128 gnd.n5119 585
R2639 gnd.n5716 gnd.n5715 585
R2640 gnd.n5717 gnd.n5716 585
R2641 gnd.n5129 gnd.n5127 585
R2642 gnd.n5136 gnd.n5127 585
R2643 gnd.n5709 gnd.n5708 585
R2644 gnd.n5708 gnd.n5707 585
R2645 gnd.n5132 gnd.n5131 585
R2646 gnd.n5696 gnd.n5132 585
R2647 gnd.n5683 gnd.n5154 585
R2648 gnd.n5154 gnd.n5144 585
R2649 gnd.n5685 gnd.n5684 585
R2650 gnd.n5686 gnd.n5685 585
R2651 gnd.n5155 gnd.n5153 585
R2652 gnd.n5162 gnd.n5153 585
R2653 gnd.n5678 gnd.n5677 585
R2654 gnd.n5677 gnd.n5676 585
R2655 gnd.n5158 gnd.n5157 585
R2656 gnd.n5665 gnd.n5158 585
R2657 gnd.n5652 gnd.n5179 585
R2658 gnd.n5179 gnd.n5170 585
R2659 gnd.n5654 gnd.n5653 585
R2660 gnd.n5655 gnd.n5654 585
R2661 gnd.n5180 gnd.n5178 585
R2662 gnd.n5187 gnd.n5178 585
R2663 gnd.n5647 gnd.n5646 585
R2664 gnd.n5646 gnd.n5645 585
R2665 gnd.n5183 gnd.n5182 585
R2666 gnd.n5634 gnd.n5183 585
R2667 gnd.n5621 gnd.n5205 585
R2668 gnd.n5205 gnd.n5204 585
R2669 gnd.n5623 gnd.n5622 585
R2670 gnd.n5624 gnd.n5623 585
R2671 gnd.n5206 gnd.n5203 585
R2672 gnd.n5213 gnd.n5203 585
R2673 gnd.n5616 gnd.n5615 585
R2674 gnd.n5615 gnd.n5614 585
R2675 gnd.n5209 gnd.n5208 585
R2676 gnd.n5603 gnd.n5209 585
R2677 gnd.n5590 gnd.n5230 585
R2678 gnd.n5230 gnd.n5229 585
R2679 gnd.n5592 gnd.n5591 585
R2680 gnd.n5593 gnd.n5592 585
R2681 gnd.n5586 gnd.n5228 585
R2682 gnd.n5585 gnd.n5584 585
R2683 gnd.n5233 gnd.n5232 585
R2684 gnd.n5582 gnd.n5233 585
R2685 gnd.n5255 gnd.n5254 585
R2686 gnd.n5258 gnd.n5257 585
R2687 gnd.n5256 gnd.n5251 585
R2688 gnd.n5263 gnd.n5262 585
R2689 gnd.n5265 gnd.n5264 585
R2690 gnd.n5268 gnd.n5267 585
R2691 gnd.n5266 gnd.n5249 585
R2692 gnd.n5273 gnd.n5272 585
R2693 gnd.n5275 gnd.n5274 585
R2694 gnd.n5278 gnd.n5277 585
R2695 gnd.n5276 gnd.n5247 585
R2696 gnd.n5283 gnd.n5282 585
R2697 gnd.n5287 gnd.n5284 585
R2698 gnd.n5288 gnd.n5225 585
R2699 gnd.n6277 gnd.n6276 585
R2700 gnd.n6279 gnd.n4938 585
R2701 gnd.n6281 gnd.n6280 585
R2702 gnd.n6282 gnd.n4931 585
R2703 gnd.n6284 gnd.n6283 585
R2704 gnd.n6286 gnd.n4929 585
R2705 gnd.n6288 gnd.n6287 585
R2706 gnd.n6289 gnd.n4924 585
R2707 gnd.n6291 gnd.n6290 585
R2708 gnd.n6293 gnd.n4922 585
R2709 gnd.n6295 gnd.n6294 585
R2710 gnd.n6296 gnd.n4917 585
R2711 gnd.n6298 gnd.n6297 585
R2712 gnd.n6300 gnd.n4915 585
R2713 gnd.n6302 gnd.n6301 585
R2714 gnd.n6303 gnd.n4913 585
R2715 gnd.n6304 gnd.n4908 585
R2716 gnd.n4908 gnd.n4906 585
R2717 gnd.n6166 gnd.n932 585
R2718 gnd.n6309 gnd.n932 585
R2719 gnd.n6168 gnd.n6167 585
R2720 gnd.n6168 gnd.n930 585
R2721 gnd.n6170 gnd.n6169 585
R2722 gnd.n6169 gnd.n922 585
R2723 gnd.n6171 gnd.n920 585
R2724 gnd.n6317 gnd.n920 585
R2725 gnd.n6174 gnd.n6173 585
R2726 gnd.n6173 gnd.n6172 585
R2727 gnd.n6175 gnd.n909 585
R2728 gnd.n6323 gnd.n909 585
R2729 gnd.n6177 gnd.n6176 585
R2730 gnd.n6177 gnd.n907 585
R2731 gnd.n6178 gnd.n5901 585
R2732 gnd.n6178 gnd.n898 585
R2733 gnd.n6180 gnd.n6179 585
R2734 gnd.n6179 gnd.n896 585
R2735 gnd.n6181 gnd.n4996 585
R2736 gnd.n6202 gnd.n4996 585
R2737 gnd.n5898 gnd.n5897 585
R2738 gnd.n5897 gnd.n5006 585
R2739 gnd.n5896 gnd.n5004 585
R2740 gnd.n6188 gnd.n5004 585
R2741 gnd.n5887 gnd.n5014 585
R2742 gnd.n5888 gnd.n5887 585
R2743 gnd.n5886 gnd.n5885 585
R2744 gnd.n5886 gnd.n5018 585
R2745 gnd.n5884 gnd.n5020 585
R2746 gnd.n5877 gnd.n5020 585
R2747 gnd.n5864 gnd.n5021 585
R2748 gnd.n5865 gnd.n5864 585
R2749 gnd.n5838 gnd.n5033 585
R2750 gnd.n5867 gnd.n5033 585
R2751 gnd.n5837 gnd.n5836 585
R2752 gnd.n5836 gnd.n5835 585
R2753 gnd.n5833 gnd.n5046 585
R2754 gnd.n5833 gnd.n5039 585
R2755 gnd.n5832 gnd.n5048 585
R2756 gnd.n5832 gnd.n5831 585
R2757 gnd.n5811 gnd.n5047 585
R2758 gnd.n5060 gnd.n5047 585
R2759 gnd.n5810 gnd.n5058 585
R2760 gnd.n5821 gnd.n5058 585
R2761 gnd.n5801 gnd.n5065 585
R2762 gnd.n5802 gnd.n5801 585
R2763 gnd.n5800 gnd.n5071 585
R2764 gnd.n5800 gnd.n5799 585
R2765 gnd.n5785 gnd.n5070 585
R2766 gnd.n5080 gnd.n5070 585
R2767 gnd.n5784 gnd.n5078 585
R2768 gnd.n5791 gnd.n5078 585
R2769 gnd.n5783 gnd.n5782 585
R2770 gnd.n5782 gnd.n5781 585
R2771 gnd.n5088 gnd.n5085 585
R2772 gnd.n5095 gnd.n5088 585
R2773 gnd.n5749 gnd.n5748 585
R2774 gnd.n5748 gnd.n5747 585
R2775 gnd.n5101 gnd.n5100 585
R2776 gnd.n5112 gnd.n5101 585
R2777 gnd.n5730 gnd.n5110 585
R2778 gnd.n5737 gnd.n5110 585
R2779 gnd.n5729 gnd.n5728 585
R2780 gnd.n5728 gnd.n5727 585
R2781 gnd.n5118 gnd.n5116 585
R2782 gnd.n5119 gnd.n5118 585
R2783 gnd.n5719 gnd.n5718 585
R2784 gnd.n5718 gnd.n5717 585
R2785 gnd.n5125 gnd.n5124 585
R2786 gnd.n5136 gnd.n5125 585
R2787 gnd.n5699 gnd.n5134 585
R2788 gnd.n5707 gnd.n5134 585
R2789 gnd.n5698 gnd.n5697 585
R2790 gnd.n5697 gnd.n5696 585
R2791 gnd.n5143 gnd.n5141 585
R2792 gnd.n5144 gnd.n5143 585
R2793 gnd.n5688 gnd.n5687 585
R2794 gnd.n5687 gnd.n5686 585
R2795 gnd.n5150 gnd.n5149 585
R2796 gnd.n5162 gnd.n5150 585
R2797 gnd.n5668 gnd.n5160 585
R2798 gnd.n5676 gnd.n5160 585
R2799 gnd.n5667 gnd.n5666 585
R2800 gnd.n5666 gnd.n5665 585
R2801 gnd.n5169 gnd.n5167 585
R2802 gnd.n5170 gnd.n5169 585
R2803 gnd.n5657 gnd.n5656 585
R2804 gnd.n5656 gnd.n5655 585
R2805 gnd.n5176 gnd.n5175 585
R2806 gnd.n5187 gnd.n5176 585
R2807 gnd.n5637 gnd.n5185 585
R2808 gnd.n5645 gnd.n5185 585
R2809 gnd.n5636 gnd.n5635 585
R2810 gnd.n5635 gnd.n5634 585
R2811 gnd.n5194 gnd.n5192 585
R2812 gnd.n5204 gnd.n5194 585
R2813 gnd.n5626 gnd.n5625 585
R2814 gnd.n5625 gnd.n5624 585
R2815 gnd.n5200 gnd.n5199 585
R2816 gnd.n5213 gnd.n5200 585
R2817 gnd.n5606 gnd.n5211 585
R2818 gnd.n5614 gnd.n5211 585
R2819 gnd.n5605 gnd.n5604 585
R2820 gnd.n5604 gnd.n5603 585
R2821 gnd.n5220 gnd.n5218 585
R2822 gnd.n5229 gnd.n5220 585
R2823 gnd.n5595 gnd.n5594 585
R2824 gnd.n5594 gnd.n5593 585
R2825 gnd.n4669 gnd.n4668 585
R2826 gnd.n4668 gnd.n4667 585
R2827 gnd.n4670 gnd.n1264 585
R2828 gnd.n2831 gnd.n1264 585
R2829 gnd.n4672 gnd.n4671 585
R2830 gnd.n4673 gnd.n4672 585
R2831 gnd.n1249 gnd.n1248 585
R2832 gnd.n2793 gnd.n1249 585
R2833 gnd.n4681 gnd.n4680 585
R2834 gnd.n4680 gnd.n4679 585
R2835 gnd.n4682 gnd.n1243 585
R2836 gnd.n2784 gnd.n1243 585
R2837 gnd.n4684 gnd.n4683 585
R2838 gnd.n4685 gnd.n4684 585
R2839 gnd.n1228 gnd.n1227 585
R2840 gnd.n2776 gnd.n1228 585
R2841 gnd.n4693 gnd.n4692 585
R2842 gnd.n4692 gnd.n4691 585
R2843 gnd.n4694 gnd.n1222 585
R2844 gnd.n2709 gnd.n1222 585
R2845 gnd.n4696 gnd.n4695 585
R2846 gnd.n4697 gnd.n4696 585
R2847 gnd.n1207 gnd.n1206 585
R2848 gnd.n2697 gnd.n1207 585
R2849 gnd.n4705 gnd.n4704 585
R2850 gnd.n4704 gnd.n4703 585
R2851 gnd.n4706 gnd.n1201 585
R2852 gnd.n2692 gnd.n1201 585
R2853 gnd.n4708 gnd.n4707 585
R2854 gnd.n4709 gnd.n4708 585
R2855 gnd.n1186 gnd.n1185 585
R2856 gnd.n2723 gnd.n1186 585
R2857 gnd.n4717 gnd.n4716 585
R2858 gnd.n4716 gnd.n4715 585
R2859 gnd.n4718 gnd.n1180 585
R2860 gnd.n2684 gnd.n1180 585
R2861 gnd.n4720 gnd.n4719 585
R2862 gnd.n4721 gnd.n4720 585
R2863 gnd.n1165 gnd.n1164 585
R2864 gnd.n2676 gnd.n1165 585
R2865 gnd.n4729 gnd.n4728 585
R2866 gnd.n4728 gnd.n4727 585
R2867 gnd.n4730 gnd.n1160 585
R2868 gnd.n2667 gnd.n1160 585
R2869 gnd.n4732 gnd.n4731 585
R2870 gnd.n4733 gnd.n4732 585
R2871 gnd.n1161 gnd.n1145 585
R2872 gnd.n2659 gnd.n1145 585
R2873 gnd.n4741 gnd.n4740 585
R2874 gnd.n4740 gnd.n4739 585
R2875 gnd.n4742 gnd.n1142 585
R2876 gnd.n2627 gnd.n1142 585
R2877 gnd.n4745 gnd.n4744 585
R2878 gnd.n4746 gnd.n4745 585
R2879 gnd.n1143 gnd.n1127 585
R2880 gnd.n2636 gnd.n1127 585
R2881 gnd.n4754 gnd.n4753 585
R2882 gnd.n4753 gnd.n4752 585
R2883 gnd.n4755 gnd.n1123 585
R2884 gnd.n2642 gnd.n1123 585
R2885 gnd.n4757 gnd.n4756 585
R2886 gnd.n4758 gnd.n4757 585
R2887 gnd.n1108 gnd.n1107 585
R2888 gnd.n2648 gnd.n1108 585
R2889 gnd.n4766 gnd.n4765 585
R2890 gnd.n4765 gnd.n4764 585
R2891 gnd.n4767 gnd.n1102 585
R2892 gnd.n2592 gnd.n1102 585
R2893 gnd.n4769 gnd.n4768 585
R2894 gnd.n4770 gnd.n4769 585
R2895 gnd.n1087 gnd.n1086 585
R2896 gnd.n1098 gnd.n1087 585
R2897 gnd.n4778 gnd.n4777 585
R2898 gnd.n4777 gnd.n4776 585
R2899 gnd.n4779 gnd.n1081 585
R2900 gnd.n1081 gnd.n1080 585
R2901 gnd.n4781 gnd.n4780 585
R2902 gnd.n4782 gnd.n4781 585
R2903 gnd.n1066 gnd.n1065 585
R2904 gnd.n1070 gnd.n1066 585
R2905 gnd.n4790 gnd.n4789 585
R2906 gnd.n4789 gnd.n4788 585
R2907 gnd.n4791 gnd.n1060 585
R2908 gnd.n1067 gnd.n1060 585
R2909 gnd.n4793 gnd.n4792 585
R2910 gnd.n4794 gnd.n4793 585
R2911 gnd.n1047 gnd.n1046 585
R2912 gnd.n1057 gnd.n1047 585
R2913 gnd.n4802 gnd.n4801 585
R2914 gnd.n4801 gnd.n4800 585
R2915 gnd.n4803 gnd.n1041 585
R2916 gnd.n1041 gnd.n1040 585
R2917 gnd.n4805 gnd.n4804 585
R2918 gnd.n4806 gnd.n4805 585
R2919 gnd.n1026 gnd.n1025 585
R2920 gnd.n1029 gnd.n1026 585
R2921 gnd.n4814 gnd.n4813 585
R2922 gnd.n4813 gnd.n4812 585
R2923 gnd.n4815 gnd.n1020 585
R2924 gnd.n1020 gnd.n1017 585
R2925 gnd.n4817 gnd.n4816 585
R2926 gnd.n4818 gnd.n4817 585
R2927 gnd.n1021 gnd.n1019 585
R2928 gnd.n1019 gnd.n1015 585
R2929 gnd.n2549 gnd.n2548 585
R2930 gnd.n2550 gnd.n2549 585
R2931 gnd.n2544 gnd.n964 585
R2932 gnd.n964 gnd.n961 585
R2933 gnd.n4903 gnd.n4902 585
R2934 gnd.n4901 gnd.n963 585
R2935 gnd.n4900 gnd.n962 585
R2936 gnd.n4905 gnd.n962 585
R2937 gnd.n4899 gnd.n4898 585
R2938 gnd.n4897 gnd.n4896 585
R2939 gnd.n4895 gnd.n4894 585
R2940 gnd.n4893 gnd.n4892 585
R2941 gnd.n4891 gnd.n4890 585
R2942 gnd.n4889 gnd.n4888 585
R2943 gnd.n4887 gnd.n4886 585
R2944 gnd.n4885 gnd.n4884 585
R2945 gnd.n4883 gnd.n4882 585
R2946 gnd.n4881 gnd.n4880 585
R2947 gnd.n4879 gnd.n4878 585
R2948 gnd.n4877 gnd.n4876 585
R2949 gnd.n4875 gnd.n4874 585
R2950 gnd.n4873 gnd.n4872 585
R2951 gnd.n4871 gnd.n4870 585
R2952 gnd.n4868 gnd.n4867 585
R2953 gnd.n4866 gnd.n4865 585
R2954 gnd.n4864 gnd.n4863 585
R2955 gnd.n4862 gnd.n4861 585
R2956 gnd.n4860 gnd.n4859 585
R2957 gnd.n4858 gnd.n4857 585
R2958 gnd.n4856 gnd.n4855 585
R2959 gnd.n4854 gnd.n4853 585
R2960 gnd.n4852 gnd.n4851 585
R2961 gnd.n4850 gnd.n4849 585
R2962 gnd.n4848 gnd.n4847 585
R2963 gnd.n4846 gnd.n4845 585
R2964 gnd.n4844 gnd.n4843 585
R2965 gnd.n4842 gnd.n4841 585
R2966 gnd.n4840 gnd.n4839 585
R2967 gnd.n4838 gnd.n4837 585
R2968 gnd.n4836 gnd.n4835 585
R2969 gnd.n4834 gnd.n4833 585
R2970 gnd.n4832 gnd.n1003 585
R2971 gnd.n1007 gnd.n1004 585
R2972 gnd.n4828 gnd.n4827 585
R2973 gnd.n2326 gnd.n2325 585
R2974 gnd.n2839 gnd.n2838 585
R2975 gnd.n2841 gnd.n2840 585
R2976 gnd.n2843 gnd.n2842 585
R2977 gnd.n2845 gnd.n2844 585
R2978 gnd.n2847 gnd.n2846 585
R2979 gnd.n2849 gnd.n2848 585
R2980 gnd.n2851 gnd.n2850 585
R2981 gnd.n2853 gnd.n2852 585
R2982 gnd.n2855 gnd.n2854 585
R2983 gnd.n2857 gnd.n2856 585
R2984 gnd.n2859 gnd.n2858 585
R2985 gnd.n2861 gnd.n2860 585
R2986 gnd.n2863 gnd.n2862 585
R2987 gnd.n2865 gnd.n2864 585
R2988 gnd.n2867 gnd.n2866 585
R2989 gnd.n2869 gnd.n2868 585
R2990 gnd.n2871 gnd.n2870 585
R2991 gnd.n2873 gnd.n2872 585
R2992 gnd.n2876 gnd.n2875 585
R2993 gnd.n2874 gnd.n2304 585
R2994 gnd.n3116 gnd.n3115 585
R2995 gnd.n3118 gnd.n3117 585
R2996 gnd.n3120 gnd.n3119 585
R2997 gnd.n3122 gnd.n3121 585
R2998 gnd.n3124 gnd.n3123 585
R2999 gnd.n3126 gnd.n3125 585
R3000 gnd.n3128 gnd.n3127 585
R3001 gnd.n3130 gnd.n3129 585
R3002 gnd.n3132 gnd.n3131 585
R3003 gnd.n3134 gnd.n3133 585
R3004 gnd.n3136 gnd.n3135 585
R3005 gnd.n3138 gnd.n3137 585
R3006 gnd.n3139 gnd.n2285 585
R3007 gnd.n3141 gnd.n3140 585
R3008 gnd.n2286 gnd.n2284 585
R3009 gnd.n2287 gnd.n1269 585
R3010 gnd.n3143 gnd.n1269 585
R3011 gnd.n2834 gnd.n1271 585
R3012 gnd.n4667 gnd.n1271 585
R3013 gnd.n2833 gnd.n2832 585
R3014 gnd.n2832 gnd.n2831 585
R3015 gnd.n2330 gnd.n1262 585
R3016 gnd.n4673 gnd.n1262 585
R3017 gnd.n2792 gnd.n2791 585
R3018 gnd.n2793 gnd.n2792 585
R3019 gnd.n2336 gnd.n1251 585
R3020 gnd.n4679 gnd.n1251 585
R3021 gnd.n2786 gnd.n2785 585
R3022 gnd.n2785 gnd.n2784 585
R3023 gnd.n2338 gnd.n1240 585
R3024 gnd.n4685 gnd.n1240 585
R3025 gnd.n2705 gnd.n2342 585
R3026 gnd.n2776 gnd.n2342 585
R3027 gnd.n2706 gnd.n1230 585
R3028 gnd.n4691 gnd.n1230 585
R3029 gnd.n2708 gnd.n2707 585
R3030 gnd.n2709 gnd.n2708 585
R3031 gnd.n2362 gnd.n1219 585
R3032 gnd.n4697 gnd.n1219 585
R3033 gnd.n2699 gnd.n2698 585
R3034 gnd.n2698 gnd.n2697 585
R3035 gnd.n2695 gnd.n1209 585
R3036 gnd.n4703 gnd.n1209 585
R3037 gnd.n2694 gnd.n2693 585
R3038 gnd.n2693 gnd.n2692 585
R3039 gnd.n2364 gnd.n1198 585
R3040 gnd.n4709 gnd.n1198 585
R3041 gnd.n2688 gnd.n2354 585
R3042 gnd.n2723 gnd.n2354 585
R3043 gnd.n2687 gnd.n1188 585
R3044 gnd.n4715 gnd.n1188 585
R3045 gnd.n2686 gnd.n2685 585
R3046 gnd.n2685 gnd.n2684 585
R3047 gnd.n2366 gnd.n1177 585
R3048 gnd.n4721 gnd.n1177 585
R3049 gnd.n2675 gnd.n2674 585
R3050 gnd.n2676 gnd.n2675 585
R3051 gnd.n2372 gnd.n1167 585
R3052 gnd.n4727 gnd.n1167 585
R3053 gnd.n2669 gnd.n2668 585
R3054 gnd.n2668 gnd.n2667 585
R3055 gnd.n2374 gnd.n1157 585
R3056 gnd.n4733 gnd.n1157 585
R3057 gnd.n2623 gnd.n2378 585
R3058 gnd.n2659 gnd.n2378 585
R3059 gnd.n2624 gnd.n1147 585
R3060 gnd.n4739 gnd.n1147 585
R3061 gnd.n2626 gnd.n2625 585
R3062 gnd.n2627 gnd.n2626 585
R3063 gnd.n2602 gnd.n1139 585
R3064 gnd.n4746 gnd.n1139 585
R3065 gnd.n2638 gnd.n2637 585
R3066 gnd.n2637 gnd.n2636 585
R3067 gnd.n2639 gnd.n1129 585
R3068 gnd.n4752 gnd.n1129 585
R3069 gnd.n2641 gnd.n2640 585
R3070 gnd.n2642 gnd.n2641 585
R3071 gnd.n2420 gnd.n1120 585
R3072 gnd.n4758 gnd.n1120 585
R3073 gnd.n2596 gnd.n2414 585
R3074 gnd.n2648 gnd.n2414 585
R3075 gnd.n2595 gnd.n1110 585
R3076 gnd.n4764 gnd.n1110 585
R3077 gnd.n2594 gnd.n2593 585
R3078 gnd.n2593 gnd.n2592 585
R3079 gnd.n2422 gnd.n1099 585
R3080 gnd.n4770 gnd.n1099 585
R3081 gnd.n2456 gnd.n2455 585
R3082 gnd.n2455 gnd.n1098 585
R3083 gnd.n2454 gnd.n1088 585
R3084 gnd.n4776 gnd.n1088 585
R3085 gnd.n2453 gnd.n2452 585
R3086 gnd.n2452 gnd.n1080 585
R3087 gnd.n2424 gnd.n1078 585
R3088 gnd.n4782 gnd.n1078 585
R3089 gnd.n2448 gnd.n2447 585
R3090 gnd.n2447 gnd.n1070 585
R3091 gnd.n2446 gnd.n1068 585
R3092 gnd.n4788 gnd.n1068 585
R3093 gnd.n2445 gnd.n2444 585
R3094 gnd.n2444 gnd.n1067 585
R3095 gnd.n2426 gnd.n1058 585
R3096 gnd.n4794 gnd.n1058 585
R3097 gnd.n2440 gnd.n2439 585
R3098 gnd.n2439 gnd.n1057 585
R3099 gnd.n2438 gnd.n1048 585
R3100 gnd.n4800 gnd.n1048 585
R3101 gnd.n2437 gnd.n2436 585
R3102 gnd.n2436 gnd.n1040 585
R3103 gnd.n2428 gnd.n1038 585
R3104 gnd.n4806 gnd.n1038 585
R3105 gnd.n2432 gnd.n2431 585
R3106 gnd.n2431 gnd.n1029 585
R3107 gnd.n2430 gnd.n1027 585
R3108 gnd.n4812 gnd.n1027 585
R3109 gnd.n1014 gnd.n1012 585
R3110 gnd.n1017 gnd.n1014 585
R3111 gnd.n4820 gnd.n4819 585
R3112 gnd.n4819 gnd.n4818 585
R3113 gnd.n1013 gnd.n1010 585
R3114 gnd.n1015 gnd.n1013 585
R3115 gnd.n4824 gnd.n1009 585
R3116 gnd.n2550 gnd.n1009 585
R3117 gnd.n4826 gnd.n4825 585
R3118 gnd.n4826 gnd.n961 585
R3119 gnd.n7533 gnd.n7532 585
R3120 gnd.n7534 gnd.n7533 585
R3121 gnd.n110 gnd.n108 585
R3122 gnd.n108 gnd.n104 585
R3123 gnd.n7453 gnd.n7452 585
R3124 gnd.n7454 gnd.n7453 585
R3125 gnd.n189 gnd.n188 585
R3126 gnd.n188 gnd.n185 585
R3127 gnd.n7448 gnd.n7447 585
R3128 gnd.n7447 gnd.n7446 585
R3129 gnd.n192 gnd.n191 585
R3130 gnd.n193 gnd.n192 585
R3131 gnd.n7362 gnd.n7361 585
R3132 gnd.n7363 gnd.n7362 585
R3133 gnd.n204 gnd.n203 585
R3134 gnd.n211 gnd.n203 585
R3135 gnd.n7357 gnd.n7356 585
R3136 gnd.n7356 gnd.n7355 585
R3137 gnd.n207 gnd.n206 585
R3138 gnd.n208 gnd.n207 585
R3139 gnd.n7346 gnd.n7345 585
R3140 gnd.n7347 gnd.n7346 585
R3141 gnd.n221 gnd.n220 585
R3142 gnd.n220 gnd.n218 585
R3143 gnd.n7341 gnd.n7340 585
R3144 gnd.n7340 gnd.n7339 585
R3145 gnd.n224 gnd.n223 585
R3146 gnd.n225 gnd.n224 585
R3147 gnd.n7330 gnd.n7329 585
R3148 gnd.n7331 gnd.n7330 585
R3149 gnd.n234 gnd.n233 585
R3150 gnd.n241 gnd.n233 585
R3151 gnd.n7325 gnd.n7324 585
R3152 gnd.n7324 gnd.n7323 585
R3153 gnd.n237 gnd.n236 585
R3154 gnd.n238 gnd.n237 585
R3155 gnd.n7314 gnd.n7313 585
R3156 gnd.n7315 gnd.n7314 585
R3157 gnd.n252 gnd.n251 585
R3158 gnd.n251 gnd.n248 585
R3159 gnd.n7309 gnd.n7308 585
R3160 gnd.n7308 gnd.n7307 585
R3161 gnd.n255 gnd.n254 585
R3162 gnd.n7260 gnd.n255 585
R3163 gnd.n7298 gnd.n7297 585
R3164 gnd.n7299 gnd.n7298 585
R3165 gnd.n267 gnd.n266 585
R3166 gnd.n7265 gnd.n266 585
R3167 gnd.n7275 gnd.n7274 585
R3168 gnd.n7276 gnd.n7275 585
R3169 gnd.n7273 gnd.n7272 585
R3170 gnd.n7272 gnd.n7271 585
R3171 gnd.n7202 gnd.n297 585
R3172 gnd.n320 gnd.n297 585
R3173 gnd.n7204 gnd.n7203 585
R3174 gnd.n7205 gnd.n7204 585
R3175 gnd.n7201 gnd.n306 585
R3176 gnd.n7201 gnd.n7200 585
R3177 gnd.n305 gnd.n273 585
R3178 gnd.n314 gnd.n305 585
R3179 gnd.n277 gnd.n274 585
R3180 gnd.n7192 gnd.n277 585
R3181 gnd.n7294 gnd.n7293 585
R3182 gnd.n7293 gnd.n7292 585
R3183 gnd.n276 gnd.n275 585
R3184 gnd.n4349 gnd.n276 585
R3185 gnd.n4386 gnd.n4385 585
R3186 gnd.n4387 gnd.n4386 585
R3187 gnd.n1531 gnd.n1530 585
R3188 gnd.n1538 gnd.n1530 585
R3189 gnd.n4381 gnd.n4380 585
R3190 gnd.n4380 gnd.n4379 585
R3191 gnd.n1534 gnd.n1533 585
R3192 gnd.n4361 gnd.n1534 585
R3193 gnd.n4323 gnd.n1565 585
R3194 gnd.n1565 gnd.n1546 585
R3195 gnd.n4325 gnd.n4324 585
R3196 gnd.n4326 gnd.n4325 585
R3197 gnd.n1566 gnd.n1564 585
R3198 gnd.n1573 gnd.n1564 585
R3199 gnd.n4318 gnd.n4317 585
R3200 gnd.n4317 gnd.n4316 585
R3201 gnd.n1569 gnd.n1568 585
R3202 gnd.n4303 gnd.n1569 585
R3203 gnd.n4286 gnd.n1592 585
R3204 gnd.n1592 gnd.n1580 585
R3205 gnd.n4288 gnd.n4287 585
R3206 gnd.n4289 gnd.n4288 585
R3207 gnd.n1593 gnd.n1591 585
R3208 gnd.n1601 gnd.n1591 585
R3209 gnd.n4281 gnd.n4280 585
R3210 gnd.n4280 gnd.n4279 585
R3211 gnd.n1596 gnd.n1595 585
R3212 gnd.n4267 gnd.n1596 585
R3213 gnd.n4255 gnd.n1620 585
R3214 gnd.n1671 gnd.n1620 585
R3215 gnd.n4257 gnd.n4256 585
R3216 gnd.n4258 gnd.n4257 585
R3217 gnd.n1621 gnd.n1619 585
R3218 gnd.n1628 gnd.n1619 585
R3219 gnd.n4250 gnd.n4249 585
R3220 gnd.n4249 gnd.n4248 585
R3221 gnd.n1624 gnd.n1623 585
R3222 gnd.n4236 gnd.n1624 585
R3223 gnd.n1646 gnd.n1645 585
R3224 gnd.n1647 gnd.n1646 585
R3225 gnd.n1642 gnd.n1449 585
R3226 gnd.n4422 gnd.n1449 585
R3227 gnd.n4496 gnd.n4495 585
R3228 gnd.n4494 gnd.n1448 585
R3229 gnd.n4493 gnd.n1447 585
R3230 gnd.n4498 gnd.n1447 585
R3231 gnd.n4492 gnd.n4491 585
R3232 gnd.n4490 gnd.n4489 585
R3233 gnd.n4488 gnd.n4487 585
R3234 gnd.n4486 gnd.n4485 585
R3235 gnd.n4484 gnd.n4483 585
R3236 gnd.n4482 gnd.n4481 585
R3237 gnd.n4480 gnd.n4479 585
R3238 gnd.n4478 gnd.n4477 585
R3239 gnd.n4476 gnd.n4475 585
R3240 gnd.n4474 gnd.n4473 585
R3241 gnd.n4472 gnd.n4471 585
R3242 gnd.n4470 gnd.n4469 585
R3243 gnd.n4468 gnd.n4467 585
R3244 gnd.n4465 gnd.n4464 585
R3245 gnd.n4463 gnd.n4462 585
R3246 gnd.n4461 gnd.n4460 585
R3247 gnd.n4459 gnd.n4458 585
R3248 gnd.n4457 gnd.n4456 585
R3249 gnd.n4455 gnd.n4454 585
R3250 gnd.n4453 gnd.n4452 585
R3251 gnd.n4451 gnd.n4450 585
R3252 gnd.n4449 gnd.n4448 585
R3253 gnd.n4447 gnd.n4446 585
R3254 gnd.n4445 gnd.n4444 585
R3255 gnd.n4443 gnd.n4442 585
R3256 gnd.n4441 gnd.n4440 585
R3257 gnd.n4439 gnd.n4438 585
R3258 gnd.n4437 gnd.n4436 585
R3259 gnd.n4435 gnd.n4434 585
R3260 gnd.n4433 gnd.n4432 585
R3261 gnd.n4431 gnd.n4430 585
R3262 gnd.n4429 gnd.n1489 585
R3263 gnd.n1493 gnd.n1490 585
R3264 gnd.n4425 gnd.n4424 585
R3265 gnd.n178 gnd.n177 585
R3266 gnd.n7462 gnd.n173 585
R3267 gnd.n7464 gnd.n7463 585
R3268 gnd.n7466 gnd.n171 585
R3269 gnd.n7468 gnd.n7467 585
R3270 gnd.n7469 gnd.n166 585
R3271 gnd.n7471 gnd.n7470 585
R3272 gnd.n7473 gnd.n164 585
R3273 gnd.n7475 gnd.n7474 585
R3274 gnd.n7476 gnd.n159 585
R3275 gnd.n7478 gnd.n7477 585
R3276 gnd.n7480 gnd.n157 585
R3277 gnd.n7482 gnd.n7481 585
R3278 gnd.n7483 gnd.n152 585
R3279 gnd.n7485 gnd.n7484 585
R3280 gnd.n7487 gnd.n150 585
R3281 gnd.n7489 gnd.n7488 585
R3282 gnd.n7490 gnd.n145 585
R3283 gnd.n7492 gnd.n7491 585
R3284 gnd.n7494 gnd.n143 585
R3285 gnd.n7496 gnd.n7495 585
R3286 gnd.n7500 gnd.n138 585
R3287 gnd.n7502 gnd.n7501 585
R3288 gnd.n7504 gnd.n136 585
R3289 gnd.n7506 gnd.n7505 585
R3290 gnd.n7507 gnd.n131 585
R3291 gnd.n7509 gnd.n7508 585
R3292 gnd.n7511 gnd.n129 585
R3293 gnd.n7513 gnd.n7512 585
R3294 gnd.n7514 gnd.n124 585
R3295 gnd.n7516 gnd.n7515 585
R3296 gnd.n7518 gnd.n122 585
R3297 gnd.n7520 gnd.n7519 585
R3298 gnd.n7521 gnd.n117 585
R3299 gnd.n7523 gnd.n7522 585
R3300 gnd.n7525 gnd.n115 585
R3301 gnd.n7527 gnd.n7526 585
R3302 gnd.n7528 gnd.n113 585
R3303 gnd.n7529 gnd.n109 585
R3304 gnd.n109 gnd.n106 585
R3305 gnd.n7458 gnd.n105 585
R3306 gnd.n7534 gnd.n105 585
R3307 gnd.n7457 gnd.n7456 585
R3308 gnd.n7456 gnd.n104 585
R3309 gnd.n7455 gnd.n182 585
R3310 gnd.n7455 gnd.n7454 585
R3311 gnd.n7234 gnd.n183 585
R3312 gnd.n185 gnd.n183 585
R3313 gnd.n7235 gnd.n194 585
R3314 gnd.n7446 gnd.n194 585
R3315 gnd.n7237 gnd.n7236 585
R3316 gnd.n7236 gnd.n193 585
R3317 gnd.n7238 gnd.n202 585
R3318 gnd.n7363 gnd.n202 585
R3319 gnd.n7240 gnd.n7239 585
R3320 gnd.n7239 gnd.n211 585
R3321 gnd.n7241 gnd.n209 585
R3322 gnd.n7355 gnd.n209 585
R3323 gnd.n7243 gnd.n7242 585
R3324 gnd.n7242 gnd.n208 585
R3325 gnd.n7244 gnd.n219 585
R3326 gnd.n7347 gnd.n219 585
R3327 gnd.n7246 gnd.n7245 585
R3328 gnd.n7245 gnd.n218 585
R3329 gnd.n7247 gnd.n226 585
R3330 gnd.n7339 gnd.n226 585
R3331 gnd.n7249 gnd.n7248 585
R3332 gnd.n7248 gnd.n225 585
R3333 gnd.n7250 gnd.n232 585
R3334 gnd.n7331 gnd.n232 585
R3335 gnd.n7252 gnd.n7251 585
R3336 gnd.n7251 gnd.n241 585
R3337 gnd.n7253 gnd.n239 585
R3338 gnd.n7323 gnd.n239 585
R3339 gnd.n7255 gnd.n7254 585
R3340 gnd.n7254 gnd.n238 585
R3341 gnd.n7256 gnd.n249 585
R3342 gnd.n7315 gnd.n249 585
R3343 gnd.n7258 gnd.n7257 585
R3344 gnd.n7257 gnd.n248 585
R3345 gnd.n7259 gnd.n257 585
R3346 gnd.n7307 gnd.n257 585
R3347 gnd.n7262 gnd.n7261 585
R3348 gnd.n7261 gnd.n7260 585
R3349 gnd.n7263 gnd.n264 585
R3350 gnd.n7299 gnd.n264 585
R3351 gnd.n7267 gnd.n7266 585
R3352 gnd.n7266 gnd.n7265 585
R3353 gnd.n7268 gnd.n295 585
R3354 gnd.n7276 gnd.n295 585
R3355 gnd.n7270 gnd.n7269 585
R3356 gnd.n7271 gnd.n7270 585
R3357 gnd.n7208 gnd.n298 585
R3358 gnd.n320 gnd.n298 585
R3359 gnd.n7207 gnd.n7206 585
R3360 gnd.n7206 gnd.n7205 585
R3361 gnd.n301 gnd.n299 585
R3362 gnd.n7200 gnd.n301 585
R3363 gnd.n4344 gnd.n4343 585
R3364 gnd.n4343 gnd.n314 585
R3365 gnd.n4345 gnd.n313 585
R3366 gnd.n7192 gnd.n313 585
R3367 gnd.n4346 gnd.n279 585
R3368 gnd.n7292 gnd.n279 585
R3369 gnd.n4348 gnd.n4347 585
R3370 gnd.n4349 gnd.n4348 585
R3371 gnd.n1554 gnd.n1527 585
R3372 gnd.n4387 gnd.n1527 585
R3373 gnd.n4335 gnd.n4334 585
R3374 gnd.n4334 gnd.n1538 585
R3375 gnd.n4333 gnd.n1536 585
R3376 gnd.n4379 gnd.n1536 585
R3377 gnd.n4332 gnd.n1547 585
R3378 gnd.n4361 gnd.n1547 585
R3379 gnd.n1560 gnd.n1556 585
R3380 gnd.n1560 gnd.n1546 585
R3381 gnd.n4328 gnd.n4327 585
R3382 gnd.n4327 gnd.n4326 585
R3383 gnd.n1559 gnd.n1558 585
R3384 gnd.n1573 gnd.n1559 585
R3385 gnd.n1662 gnd.n1571 585
R3386 gnd.n4316 gnd.n1571 585
R3387 gnd.n1663 gnd.n1581 585
R3388 gnd.n4303 gnd.n1581 585
R3389 gnd.n1665 gnd.n1664 585
R3390 gnd.n1664 gnd.n1580 585
R3391 gnd.n1666 gnd.n1589 585
R3392 gnd.n4289 gnd.n1589 585
R3393 gnd.n1668 gnd.n1667 585
R3394 gnd.n1667 gnd.n1601 585
R3395 gnd.n1669 gnd.n1598 585
R3396 gnd.n4279 gnd.n1598 585
R3397 gnd.n1670 gnd.n1608 585
R3398 gnd.n4267 gnd.n1608 585
R3399 gnd.n1673 gnd.n1672 585
R3400 gnd.n1672 gnd.n1671 585
R3401 gnd.n1674 gnd.n1616 585
R3402 gnd.n4258 gnd.n1616 585
R3403 gnd.n1676 gnd.n1675 585
R3404 gnd.n1675 gnd.n1628 585
R3405 gnd.n1677 gnd.n1626 585
R3406 gnd.n4248 gnd.n1626 585
R3407 gnd.n1679 gnd.n1678 585
R3408 gnd.n4236 gnd.n1679 585
R3409 gnd.n1648 gnd.n1495 585
R3410 gnd.n1647 gnd.n1495 585
R3411 gnd.n4423 gnd.n1496 585
R3412 gnd.n4423 gnd.n4422 585
R3413 gnd.n3687 gnd.n3495 585
R3414 gnd.n3495 gnd.n1876 585
R3415 gnd.n3689 gnd.n3688 585
R3416 gnd.n3690 gnd.n3689 585
R3417 gnd.n3488 gnd.n3487 585
R3418 gnd.n3488 gnd.n1884 585
R3419 gnd.n3698 gnd.n3697 585
R3420 gnd.n3697 gnd.n3696 585
R3421 gnd.n3699 gnd.n3485 585
R3422 gnd.n3490 gnd.n3485 585
R3423 gnd.n3701 gnd.n3700 585
R3424 gnd.n3702 gnd.n3701 585
R3425 gnd.n3486 gnd.n3475 585
R3426 gnd.n3475 gnd.n1890 585
R3427 gnd.n3709 gnd.n3476 585
R3428 gnd.n3709 gnd.n3708 585
R3429 gnd.n3710 gnd.n3474 585
R3430 gnd.n3710 gnd.n1898 585
R3431 gnd.n3712 gnd.n3711 585
R3432 gnd.n3711 gnd.n1897 585
R3433 gnd.n3713 gnd.n3471 585
R3434 gnd.n3471 gnd.n3470 585
R3435 gnd.n3715 gnd.n3714 585
R3436 gnd.n3716 gnd.n3715 585
R3437 gnd.n3473 gnd.n3469 585
R3438 gnd.n3469 gnd.n1904 585
R3439 gnd.n3472 gnd.n3461 585
R3440 gnd.n3723 gnd.n3461 585
R3441 gnd.n3725 gnd.n3460 585
R3442 gnd.n3725 gnd.n3724 585
R3443 gnd.n3727 gnd.n3726 585
R3444 gnd.n3726 gnd.n1911 585
R3445 gnd.n3728 gnd.n3458 585
R3446 gnd.n3458 gnd.n3457 585
R3447 gnd.n3730 gnd.n3729 585
R3448 gnd.n3731 gnd.n3730 585
R3449 gnd.n3459 gnd.n3455 585
R3450 gnd.n3455 gnd.n1917 585
R3451 gnd.n3449 gnd.n3448 585
R3452 gnd.n3738 gnd.n3449 585
R3453 gnd.n3741 gnd.n3740 585
R3454 gnd.n3740 gnd.n3739 585
R3455 gnd.n3742 gnd.n3445 585
R3456 gnd.n3445 gnd.n1924 585
R3457 gnd.n3744 gnd.n3743 585
R3458 gnd.n3745 gnd.n3744 585
R3459 gnd.n3447 gnd.n3444 585
R3460 gnd.n3444 gnd.n3442 585
R3461 gnd.n3446 gnd.n3434 585
R3462 gnd.n3751 gnd.n3434 585
R3463 gnd.n3754 gnd.n3433 585
R3464 gnd.n3754 gnd.n3753 585
R3465 gnd.n3756 gnd.n3755 585
R3466 gnd.n3755 gnd.n1936 585
R3467 gnd.n3757 gnd.n3431 585
R3468 gnd.n3431 gnd.n3430 585
R3469 gnd.n3759 gnd.n3758 585
R3470 gnd.n3760 gnd.n3759 585
R3471 gnd.n3432 gnd.n3429 585
R3472 gnd.n3429 gnd.n1943 585
R3473 gnd.n3421 gnd.n3420 585
R3474 gnd.n3766 gnd.n3421 585
R3475 gnd.n3770 gnd.n3769 585
R3476 gnd.n3769 gnd.n3768 585
R3477 gnd.n3771 gnd.n3417 585
R3478 gnd.n3417 gnd.n1949 585
R3479 gnd.n3773 gnd.n3772 585
R3480 gnd.n3774 gnd.n3773 585
R3481 gnd.n3419 gnd.n3416 585
R3482 gnd.n3416 gnd.n1957 585
R3483 gnd.n3418 gnd.n1955 585
R3484 gnd.n4034 gnd.n1955 585
R3485 gnd.n3409 gnd.n3408 585
R3486 gnd.n3781 gnd.n3409 585
R3487 gnd.n3785 gnd.n3784 585
R3488 gnd.n3784 gnd.n3783 585
R3489 gnd.n3786 gnd.n3405 585
R3490 gnd.n3405 gnd.n1964 585
R3491 gnd.n3788 gnd.n3787 585
R3492 gnd.n3789 gnd.n3788 585
R3493 gnd.n3407 gnd.n3404 585
R3494 gnd.n3404 gnd.n1972 585
R3495 gnd.n3406 gnd.n3395 585
R3496 gnd.n3395 gnd.n1970 585
R3497 gnd.n3797 gnd.n3394 585
R3498 gnd.n3797 gnd.n3796 585
R3499 gnd.n3799 gnd.n3798 585
R3500 gnd.n3798 gnd.n1979 585
R3501 gnd.n3800 gnd.n3391 585
R3502 gnd.n3391 gnd.n1978 585
R3503 gnd.n3802 gnd.n3801 585
R3504 gnd.n3803 gnd.n3802 585
R3505 gnd.n3393 gnd.n3390 585
R3506 gnd.n3390 gnd.n1987 585
R3507 gnd.n3392 gnd.n3381 585
R3508 gnd.n3381 gnd.n1985 585
R3509 gnd.n3811 gnd.n3380 585
R3510 gnd.n3811 gnd.n3810 585
R3511 gnd.n3813 gnd.n3812 585
R3512 gnd.n3812 gnd.n1994 585
R3513 gnd.n3814 gnd.n3377 585
R3514 gnd.n3377 gnd.n1993 585
R3515 gnd.n3816 gnd.n3815 585
R3516 gnd.n3817 gnd.n3816 585
R3517 gnd.n3379 gnd.n3376 585
R3518 gnd.n3376 gnd.n2002 585
R3519 gnd.n3378 gnd.n3367 585
R3520 gnd.n3367 gnd.n2000 585
R3521 gnd.n3825 gnd.n3366 585
R3522 gnd.n3825 gnd.n3824 585
R3523 gnd.n3827 gnd.n3826 585
R3524 gnd.n3826 gnd.n2009 585
R3525 gnd.n3828 gnd.n3363 585
R3526 gnd.n3363 gnd.n2008 585
R3527 gnd.n3830 gnd.n3829 585
R3528 gnd.n3831 gnd.n3830 585
R3529 gnd.n3365 gnd.n3362 585
R3530 gnd.n3362 gnd.n2017 585
R3531 gnd.n3364 gnd.n3355 585
R3532 gnd.n3355 gnd.n2015 585
R3533 gnd.n3839 gnd.n3354 585
R3534 gnd.n3839 gnd.n3838 585
R3535 gnd.n3841 gnd.n3840 585
R3536 gnd.n3840 gnd.n2024 585
R3537 gnd.n3842 gnd.n3351 585
R3538 gnd.n3351 gnd.n2023 585
R3539 gnd.n3844 gnd.n3843 585
R3540 gnd.n3845 gnd.n3844 585
R3541 gnd.n3353 gnd.n3350 585
R3542 gnd.n3350 gnd.n2031 585
R3543 gnd.n3352 gnd.n3340 585
R3544 gnd.n3851 gnd.n3340 585
R3545 gnd.n3854 gnd.n3339 585
R3546 gnd.n3854 gnd.n3853 585
R3547 gnd.n3856 gnd.n3855 585
R3548 gnd.n3855 gnd.n2038 585
R3549 gnd.n3857 gnd.n3336 585
R3550 gnd.n3336 gnd.n2037 585
R3551 gnd.n3859 gnd.n3858 585
R3552 gnd.n3860 gnd.n3859 585
R3553 gnd.n3338 gnd.n3335 585
R3554 gnd.n3335 gnd.n2046 585
R3555 gnd.n3337 gnd.n3327 585
R3556 gnd.n3327 gnd.n2044 585
R3557 gnd.n3869 gnd.n3326 585
R3558 gnd.n3869 gnd.n3868 585
R3559 gnd.n3871 gnd.n3870 585
R3560 gnd.n3870 gnd.n2053 585
R3561 gnd.n3872 gnd.n3323 585
R3562 gnd.n3323 gnd.n2052 585
R3563 gnd.n3874 gnd.n3873 585
R3564 gnd.n3875 gnd.n3874 585
R3565 gnd.n3325 gnd.n3322 585
R3566 gnd.n3322 gnd.n2061 585
R3567 gnd.n3324 gnd.n3314 585
R3568 gnd.n3314 gnd.n2059 585
R3569 gnd.n3884 gnd.n3313 585
R3570 gnd.n3884 gnd.n3883 585
R3571 gnd.n3886 gnd.n3885 585
R3572 gnd.n3885 gnd.n2068 585
R3573 gnd.n3887 gnd.n2092 585
R3574 gnd.n2092 gnd.n2067 585
R3575 gnd.n3889 gnd.n3888 585
R3576 gnd.n3890 gnd.n3889 585
R3577 gnd.n3312 gnd.n2091 585
R3578 gnd.n2091 gnd.n2076 585
R3579 gnd.n3311 gnd.n3310 585
R3580 gnd.n3310 gnd.n2074 585
R3581 gnd.n3309 gnd.n3306 585
R3582 gnd.n3309 gnd.n3308 585
R3583 gnd.n3305 gnd.n2082 585
R3584 gnd.n3898 gnd.n2082 585
R3585 gnd.n3304 gnd.n3303 585
R3586 gnd.n3303 gnd.n3302 585
R3587 gnd.n2094 gnd.n2093 585
R3588 gnd.n2095 gnd.n2094 585
R3589 gnd.n3027 gnd.n3026 585
R3590 gnd.n3028 gnd.n3027 585
R3591 gnd.n3025 gnd.n3023 585
R3592 gnd.n3023 gnd.n2103 585
R3593 gnd.n3024 gnd.n3013 585
R3594 gnd.n3013 gnd.n2102 585
R3595 gnd.n3037 gnd.n3012 585
R3596 gnd.n3037 gnd.n3036 585
R3597 gnd.n3039 gnd.n3038 585
R3598 gnd.n3038 gnd.n2110 585
R3599 gnd.n3040 gnd.n2907 585
R3600 gnd.n2907 gnd.n2906 585
R3601 gnd.n3042 gnd.n3041 585
R3602 gnd.n3043 gnd.n3042 585
R3603 gnd.n3011 gnd.n2905 585
R3604 gnd.n2905 gnd.n2116 585
R3605 gnd.n3009 gnd.n3008 585
R3606 gnd.n3006 gnd.n2928 585
R3607 gnd.n3005 gnd.n3004 585
R3608 gnd.n3005 gnd.n2123 585
R3609 gnd.n3003 gnd.n2929 585
R3610 gnd.n3002 gnd.n3001 585
R3611 gnd.n2999 gnd.n2930 585
R3612 gnd.n2997 gnd.n2996 585
R3613 gnd.n2995 gnd.n2931 585
R3614 gnd.n2994 gnd.n2993 585
R3615 gnd.n2991 gnd.n2932 585
R3616 gnd.n2989 gnd.n2988 585
R3617 gnd.n2987 gnd.n2933 585
R3618 gnd.n2986 gnd.n2985 585
R3619 gnd.n2983 gnd.n2934 585
R3620 gnd.n2981 gnd.n2980 585
R3621 gnd.n2979 gnd.n2935 585
R3622 gnd.n2978 gnd.n2977 585
R3623 gnd.n2975 gnd.n2936 585
R3624 gnd.n2973 gnd.n2972 585
R3625 gnd.n2971 gnd.n2937 585
R3626 gnd.n2970 gnd.n2969 585
R3627 gnd.n2967 gnd.n2938 585
R3628 gnd.n2965 gnd.n2964 585
R3629 gnd.n2963 gnd.n2939 585
R3630 gnd.n2962 gnd.n2961 585
R3631 gnd.n2959 gnd.n2940 585
R3632 gnd.n2957 gnd.n2956 585
R3633 gnd.n2955 gnd.n2941 585
R3634 gnd.n2954 gnd.n2953 585
R3635 gnd.n2951 gnd.n2950 585
R3636 gnd.n2949 gnd.n2948 585
R3637 gnd.n2947 gnd.n2881 585
R3638 gnd.n3113 gnd.n3112 585
R3639 gnd.n3110 gnd.n2880 585
R3640 gnd.n3108 gnd.n3107 585
R3641 gnd.n3106 gnd.n2883 585
R3642 gnd.n3104 gnd.n3103 585
R3643 gnd.n3101 gnd.n2886 585
R3644 gnd.n3099 gnd.n3098 585
R3645 gnd.n3097 gnd.n2887 585
R3646 gnd.n3096 gnd.n3095 585
R3647 gnd.n3093 gnd.n2888 585
R3648 gnd.n3091 gnd.n3090 585
R3649 gnd.n3089 gnd.n2889 585
R3650 gnd.n3088 gnd.n3087 585
R3651 gnd.n3085 gnd.n2890 585
R3652 gnd.n3083 gnd.n3082 585
R3653 gnd.n3081 gnd.n2891 585
R3654 gnd.n3080 gnd.n3079 585
R3655 gnd.n3077 gnd.n2892 585
R3656 gnd.n3075 gnd.n3074 585
R3657 gnd.n3073 gnd.n2893 585
R3658 gnd.n3072 gnd.n3071 585
R3659 gnd.n3069 gnd.n2894 585
R3660 gnd.n3067 gnd.n3066 585
R3661 gnd.n3065 gnd.n2895 585
R3662 gnd.n3064 gnd.n3063 585
R3663 gnd.n3061 gnd.n2896 585
R3664 gnd.n3059 gnd.n3058 585
R3665 gnd.n3057 gnd.n2897 585
R3666 gnd.n3056 gnd.n3055 585
R3667 gnd.n3053 gnd.n2898 585
R3668 gnd.n3051 gnd.n3050 585
R3669 gnd.n3049 gnd.n2899 585
R3670 gnd.n3048 gnd.n3047 585
R3671 gnd.n3568 gnd.n3567 585
R3672 gnd.n3569 gnd.n3565 585
R3673 gnd.n3571 gnd.n3570 585
R3674 gnd.n3573 gnd.n3563 585
R3675 gnd.n3575 gnd.n3574 585
R3676 gnd.n3576 gnd.n3562 585
R3677 gnd.n3578 gnd.n3577 585
R3678 gnd.n3580 gnd.n3560 585
R3679 gnd.n3582 gnd.n3581 585
R3680 gnd.n3583 gnd.n3559 585
R3681 gnd.n3585 gnd.n3584 585
R3682 gnd.n3587 gnd.n3557 585
R3683 gnd.n3589 gnd.n3588 585
R3684 gnd.n3590 gnd.n3556 585
R3685 gnd.n3592 gnd.n3591 585
R3686 gnd.n3594 gnd.n3554 585
R3687 gnd.n3596 gnd.n3595 585
R3688 gnd.n3597 gnd.n3553 585
R3689 gnd.n3599 gnd.n3598 585
R3690 gnd.n3601 gnd.n3551 585
R3691 gnd.n3603 gnd.n3602 585
R3692 gnd.n3604 gnd.n3550 585
R3693 gnd.n3606 gnd.n3605 585
R3694 gnd.n3608 gnd.n3548 585
R3695 gnd.n3610 gnd.n3609 585
R3696 gnd.n3611 gnd.n3547 585
R3697 gnd.n3613 gnd.n3612 585
R3698 gnd.n3615 gnd.n3545 585
R3699 gnd.n3617 gnd.n3616 585
R3700 gnd.n3619 gnd.n3542 585
R3701 gnd.n3621 gnd.n3620 585
R3702 gnd.n3623 gnd.n3541 585
R3703 gnd.n3624 gnd.n3516 585
R3704 gnd.n3627 gnd.n1466 585
R3705 gnd.n3629 gnd.n3628 585
R3706 gnd.n3631 gnd.n3539 585
R3707 gnd.n3633 gnd.n3632 585
R3708 gnd.n3635 gnd.n3536 585
R3709 gnd.n3637 gnd.n3636 585
R3710 gnd.n3639 gnd.n3534 585
R3711 gnd.n3641 gnd.n3640 585
R3712 gnd.n3642 gnd.n3533 585
R3713 gnd.n3644 gnd.n3643 585
R3714 gnd.n3646 gnd.n3531 585
R3715 gnd.n3648 gnd.n3647 585
R3716 gnd.n3649 gnd.n3530 585
R3717 gnd.n3651 gnd.n3650 585
R3718 gnd.n3653 gnd.n3528 585
R3719 gnd.n3655 gnd.n3654 585
R3720 gnd.n3656 gnd.n3527 585
R3721 gnd.n3658 gnd.n3657 585
R3722 gnd.n3660 gnd.n3525 585
R3723 gnd.n3662 gnd.n3661 585
R3724 gnd.n3663 gnd.n3524 585
R3725 gnd.n3665 gnd.n3664 585
R3726 gnd.n3667 gnd.n3522 585
R3727 gnd.n3669 gnd.n3668 585
R3728 gnd.n3670 gnd.n3521 585
R3729 gnd.n3672 gnd.n3671 585
R3730 gnd.n3674 gnd.n3519 585
R3731 gnd.n3676 gnd.n3675 585
R3732 gnd.n3677 gnd.n3518 585
R3733 gnd.n3679 gnd.n3678 585
R3734 gnd.n3681 gnd.n3517 585
R3735 gnd.n3682 gnd.n3515 585
R3736 gnd.n3685 gnd.n3684 585
R3737 gnd.n3493 gnd.n3492 585
R3738 gnd.n3493 gnd.n1876 585
R3739 gnd.n3692 gnd.n3691 585
R3740 gnd.n3691 gnd.n3690 585
R3741 gnd.n3693 gnd.n3491 585
R3742 gnd.n3491 gnd.n1884 585
R3743 gnd.n3695 gnd.n3694 585
R3744 gnd.n3696 gnd.n3695 585
R3745 gnd.n3484 gnd.n3483 585
R3746 gnd.n3490 gnd.n3484 585
R3747 gnd.n3704 gnd.n3703 585
R3748 gnd.n3703 gnd.n3702 585
R3749 gnd.n3705 gnd.n3479 585
R3750 gnd.n3479 gnd.n1890 585
R3751 gnd.n3707 gnd.n3706 585
R3752 gnd.n3708 gnd.n3707 585
R3753 gnd.n3482 gnd.n3478 585
R3754 gnd.n3478 gnd.n1898 585
R3755 gnd.n3481 gnd.n3480 585
R3756 gnd.n3480 gnd.n1897 585
R3757 gnd.n3468 gnd.n3467 585
R3758 gnd.n3470 gnd.n3468 585
R3759 gnd.n3718 gnd.n3717 585
R3760 gnd.n3717 gnd.n3716 585
R3761 gnd.n3719 gnd.n3463 585
R3762 gnd.n3463 gnd.n1904 585
R3763 gnd.n3721 gnd.n3720 585
R3764 gnd.n3723 gnd.n3721 585
R3765 gnd.n3466 gnd.n3462 585
R3766 gnd.n3724 gnd.n3462 585
R3767 gnd.n3465 gnd.n3464 585
R3768 gnd.n3464 gnd.n1911 585
R3769 gnd.n3454 gnd.n3453 585
R3770 gnd.n3457 gnd.n3454 585
R3771 gnd.n3733 gnd.n3732 585
R3772 gnd.n3732 gnd.n3731 585
R3773 gnd.n3734 gnd.n3451 585
R3774 gnd.n3451 gnd.n1917 585
R3775 gnd.n3736 gnd.n3735 585
R3776 gnd.n3738 gnd.n3736 585
R3777 gnd.n3452 gnd.n3450 585
R3778 gnd.n3739 gnd.n3450 585
R3779 gnd.n3441 gnd.n3440 585
R3780 gnd.n3441 gnd.n1924 585
R3781 gnd.n3747 gnd.n3746 585
R3782 gnd.n3746 gnd.n3745 585
R3783 gnd.n3748 gnd.n3436 585
R3784 gnd.n3442 gnd.n3436 585
R3785 gnd.n3750 gnd.n3749 585
R3786 gnd.n3751 gnd.n3750 585
R3787 gnd.n3439 gnd.n3435 585
R3788 gnd.n3753 gnd.n3435 585
R3789 gnd.n3438 gnd.n3437 585
R3790 gnd.n3437 gnd.n1936 585
R3791 gnd.n3427 gnd.n3426 585
R3792 gnd.n3430 gnd.n3427 585
R3793 gnd.n3762 gnd.n3761 585
R3794 gnd.n3761 gnd.n3760 585
R3795 gnd.n3763 gnd.n3423 585
R3796 gnd.n3423 gnd.n1943 585
R3797 gnd.n3765 gnd.n3764 585
R3798 gnd.n3766 gnd.n3765 585
R3799 gnd.n3425 gnd.n3422 585
R3800 gnd.n3768 gnd.n3422 585
R3801 gnd.n3424 gnd.n3414 585
R3802 gnd.n3414 gnd.n1949 585
R3803 gnd.n3775 gnd.n3413 585
R3804 gnd.n3775 gnd.n3774 585
R3805 gnd.n3777 gnd.n3776 585
R3806 gnd.n3776 gnd.n1957 585
R3807 gnd.n3778 gnd.n1958 585
R3808 gnd.n4034 gnd.n1958 585
R3809 gnd.n3780 gnd.n3779 585
R3810 gnd.n3781 gnd.n3780 585
R3811 gnd.n3412 gnd.n3410 585
R3812 gnd.n3783 gnd.n3410 585
R3813 gnd.n3411 gnd.n3402 585
R3814 gnd.n3402 gnd.n1964 585
R3815 gnd.n3790 gnd.n3401 585
R3816 gnd.n3790 gnd.n3789 585
R3817 gnd.n3792 gnd.n3791 585
R3818 gnd.n3791 gnd.n1972 585
R3819 gnd.n3793 gnd.n3398 585
R3820 gnd.n3398 gnd.n1970 585
R3821 gnd.n3795 gnd.n3794 585
R3822 gnd.n3796 gnd.n3795 585
R3823 gnd.n3400 gnd.n3397 585
R3824 gnd.n3397 gnd.n1979 585
R3825 gnd.n3399 gnd.n3388 585
R3826 gnd.n3388 gnd.n1978 585
R3827 gnd.n3804 gnd.n3387 585
R3828 gnd.n3804 gnd.n3803 585
R3829 gnd.n3806 gnd.n3805 585
R3830 gnd.n3805 gnd.n1987 585
R3831 gnd.n3807 gnd.n3384 585
R3832 gnd.n3384 gnd.n1985 585
R3833 gnd.n3809 gnd.n3808 585
R3834 gnd.n3810 gnd.n3809 585
R3835 gnd.n3386 gnd.n3383 585
R3836 gnd.n3383 gnd.n1994 585
R3837 gnd.n3385 gnd.n3374 585
R3838 gnd.n3374 gnd.n1993 585
R3839 gnd.n3818 gnd.n3373 585
R3840 gnd.n3818 gnd.n3817 585
R3841 gnd.n3820 gnd.n3819 585
R3842 gnd.n3819 gnd.n2002 585
R3843 gnd.n3821 gnd.n3370 585
R3844 gnd.n3370 gnd.n2000 585
R3845 gnd.n3823 gnd.n3822 585
R3846 gnd.n3824 gnd.n3823 585
R3847 gnd.n3372 gnd.n3369 585
R3848 gnd.n3369 gnd.n2009 585
R3849 gnd.n3371 gnd.n3360 585
R3850 gnd.n3360 gnd.n2008 585
R3851 gnd.n3832 gnd.n3359 585
R3852 gnd.n3832 gnd.n3831 585
R3853 gnd.n3834 gnd.n3833 585
R3854 gnd.n3833 gnd.n2017 585
R3855 gnd.n3835 gnd.n3357 585
R3856 gnd.n3357 gnd.n2015 585
R3857 gnd.n3837 gnd.n3836 585
R3858 gnd.n3838 gnd.n3837 585
R3859 gnd.n3358 gnd.n3356 585
R3860 gnd.n3356 gnd.n2024 585
R3861 gnd.n3348 gnd.n3347 585
R3862 gnd.n3348 gnd.n2023 585
R3863 gnd.n3847 gnd.n3846 585
R3864 gnd.n3846 gnd.n3845 585
R3865 gnd.n3848 gnd.n3342 585
R3866 gnd.n3342 gnd.n2031 585
R3867 gnd.n3850 gnd.n3849 585
R3868 gnd.n3851 gnd.n3850 585
R3869 gnd.n3346 gnd.n3341 585
R3870 gnd.n3853 gnd.n3341 585
R3871 gnd.n3345 gnd.n3344 585
R3872 gnd.n3344 gnd.n2038 585
R3873 gnd.n3343 gnd.n3333 585
R3874 gnd.n3333 gnd.n2037 585
R3875 gnd.n3861 gnd.n3332 585
R3876 gnd.n3861 gnd.n3860 585
R3877 gnd.n3863 gnd.n3862 585
R3878 gnd.n3862 gnd.n2046 585
R3879 gnd.n3864 gnd.n3329 585
R3880 gnd.n3329 gnd.n2044 585
R3881 gnd.n3866 gnd.n3865 585
R3882 gnd.n3868 gnd.n3866 585
R3883 gnd.n3331 gnd.n3328 585
R3884 gnd.n3328 gnd.n2053 585
R3885 gnd.n3330 gnd.n3320 585
R3886 gnd.n3320 gnd.n2052 585
R3887 gnd.n3876 gnd.n3319 585
R3888 gnd.n3876 gnd.n3875 585
R3889 gnd.n3878 gnd.n3877 585
R3890 gnd.n3877 gnd.n2061 585
R3891 gnd.n3879 gnd.n3316 585
R3892 gnd.n3316 gnd.n2059 585
R3893 gnd.n3881 gnd.n3880 585
R3894 gnd.n3883 gnd.n3881 585
R3895 gnd.n3318 gnd.n3315 585
R3896 gnd.n3315 gnd.n2068 585
R3897 gnd.n3317 gnd.n2088 585
R3898 gnd.n2088 gnd.n2067 585
R3899 gnd.n3891 gnd.n2089 585
R3900 gnd.n3891 gnd.n3890 585
R3901 gnd.n3892 gnd.n2087 585
R3902 gnd.n3892 gnd.n2076 585
R3903 gnd.n3894 gnd.n3893 585
R3904 gnd.n3893 gnd.n2074 585
R3905 gnd.n3895 gnd.n2085 585
R3906 gnd.n3308 gnd.n2085 585
R3907 gnd.n3897 gnd.n3896 585
R3908 gnd.n3898 gnd.n3897 585
R3909 gnd.n2086 gnd.n2084 585
R3910 gnd.n3302 gnd.n2084 585
R3911 gnd.n3020 gnd.n3019 585
R3912 gnd.n3020 gnd.n2095 585
R3913 gnd.n3029 gnd.n3018 585
R3914 gnd.n3029 gnd.n3028 585
R3915 gnd.n3031 gnd.n3030 585
R3916 gnd.n3030 gnd.n2103 585
R3917 gnd.n3032 gnd.n3015 585
R3918 gnd.n3015 gnd.n2102 585
R3919 gnd.n3034 gnd.n3033 585
R3920 gnd.n3036 gnd.n3034 585
R3921 gnd.n3017 gnd.n3014 585
R3922 gnd.n3014 gnd.n2110 585
R3923 gnd.n3016 gnd.n2901 585
R3924 gnd.n2906 gnd.n2901 585
R3925 gnd.n3044 gnd.n2902 585
R3926 gnd.n3044 gnd.n3043 585
R3927 gnd.n3045 gnd.n2900 585
R3928 gnd.n3045 gnd.n2116 585
R3929 gnd.n895 gnd.n894 585
R3930 gnd.n1097 gnd.n895 585
R3931 gnd.n7170 gnd.n7169 585
R3932 gnd.n7170 gnd.n250 585
R3933 gnd.n7172 gnd.n328 585
R3934 gnd.n7172 gnd.n7171 585
R3935 gnd.n7174 gnd.n7173 585
R3936 gnd.n7173 gnd.n256 585
R3937 gnd.n7175 gnd.n324 585
R3938 gnd.n324 gnd.n265 585
R3939 gnd.n7177 gnd.n7176 585
R3940 gnd.n7177 gnd.n263 585
R3941 gnd.n7178 gnd.n323 585
R3942 gnd.n7178 gnd.n296 585
R3943 gnd.n7180 gnd.n7179 585
R3944 gnd.n7179 gnd.n294 585
R3945 gnd.n7182 gnd.n322 585
R3946 gnd.n322 gnd.n321 585
R3947 gnd.n7184 gnd.n7183 585
R3948 gnd.n7184 gnd.n304 585
R3949 gnd.n7186 gnd.n7185 585
R3950 gnd.n7185 gnd.n302 585
R3951 gnd.n7187 gnd.n316 585
R3952 gnd.n316 gnd.n307 585
R3953 gnd.n7190 gnd.n7189 585
R3954 gnd.n7191 gnd.n7190 585
R3955 gnd.n317 gnd.n315 585
R3956 gnd.n315 gnd.n312 585
R3957 gnd.n4372 gnd.n4371 585
R3958 gnd.n4372 gnd.n278 585
R3959 gnd.n4374 gnd.n4373 585
R3960 gnd.n4373 gnd.n1529 585
R3961 gnd.n4375 gnd.n1541 585
R3962 gnd.n1541 gnd.n1540 585
R3963 gnd.n4377 gnd.n4376 585
R3964 gnd.n4378 gnd.n4377 585
R3965 gnd.n1542 gnd.n1539 585
R3966 gnd.n1539 gnd.n1535 585
R3967 gnd.n4364 gnd.n4363 585
R3968 gnd.n4363 gnd.n4362 585
R3969 gnd.n1545 gnd.n1544 585
R3970 gnd.n1563 gnd.n1545 585
R3971 gnd.n4311 gnd.n1575 585
R3972 gnd.n1575 gnd.n1561 585
R3973 gnd.n4313 gnd.n4312 585
R3974 gnd.n4314 gnd.n4313 585
R3975 gnd.n1576 gnd.n1574 585
R3976 gnd.n1574 gnd.n1570 585
R3977 gnd.n4306 gnd.n4305 585
R3978 gnd.n4305 gnd.n4304 585
R3979 gnd.n1579 gnd.n1578 585
R3980 gnd.n1590 gnd.n1579 585
R3981 gnd.n4275 gnd.n1603 585
R3982 gnd.n1603 gnd.n1588 585
R3983 gnd.n4277 gnd.n4276 585
R3984 gnd.n4278 gnd.n4277 585
R3985 gnd.n1604 gnd.n1602 585
R3986 gnd.n1602 gnd.n1597 585
R3987 gnd.n4270 gnd.n4269 585
R3988 gnd.n4269 gnd.n4268 585
R3989 gnd.n1607 gnd.n1606 585
R3990 gnd.n1617 gnd.n1607 585
R3991 gnd.n4244 gnd.n1630 585
R3992 gnd.n1630 gnd.n1615 585
R3993 gnd.n4246 gnd.n4245 585
R3994 gnd.n4247 gnd.n4246 585
R3995 gnd.n1631 gnd.n1629 585
R3996 gnd.n1629 gnd.n1625 585
R3997 gnd.n4239 gnd.n4238 585
R3998 gnd.n4238 gnd.n4237 585
R3999 gnd.n1641 gnd.n1633 585
R4000 gnd.n1641 gnd.n1499 585
R4001 gnd.n1640 gnd.n1639 585
R4002 gnd.n1640 gnd.n1497 585
R4003 gnd.n1635 gnd.n1634 585
R4004 gnd.n1634 gnd.n1446 585
R4005 gnd.n1416 gnd.n1415 585
R4006 gnd.n4499 gnd.n1416 585
R4007 gnd.n4502 gnd.n4501 585
R4008 gnd.n4501 gnd.n4500 585
R4009 gnd.n4503 gnd.n1410 585
R4010 gnd.n1417 gnd.n1410 585
R4011 gnd.n4505 gnd.n4504 585
R4012 gnd.n4506 gnd.n4505 585
R4013 gnd.n1411 gnd.n1407 585
R4014 gnd.n4507 gnd.n1407 585
R4015 gnd.n4196 gnd.n1826 585
R4016 gnd.n1826 gnd.n1406 585
R4017 gnd.n4198 gnd.n4197 585
R4018 gnd.n4199 gnd.n4198 585
R4019 gnd.n1827 gnd.n1825 585
R4020 gnd.n1825 gnd.n1823 585
R4021 gnd.n4190 gnd.n4189 585
R4022 gnd.n4189 gnd.n4188 585
R4023 gnd.n1830 gnd.n1829 585
R4024 gnd.n1831 gnd.n1830 585
R4025 gnd.n4177 gnd.n4176 585
R4026 gnd.n4178 gnd.n4177 585
R4027 gnd.n1840 gnd.n1839 585
R4028 gnd.n1845 gnd.n1839 585
R4029 gnd.n4172 gnd.n4171 585
R4030 gnd.n4171 gnd.n4170 585
R4031 gnd.n1843 gnd.n1842 585
R4032 gnd.n1844 gnd.n1843 585
R4033 gnd.n4161 gnd.n4160 585
R4034 gnd.n4162 gnd.n4161 585
R4035 gnd.n1854 gnd.n1853 585
R4036 gnd.n1853 gnd.n1851 585
R4037 gnd.n4156 gnd.n4155 585
R4038 gnd.n4155 gnd.n4154 585
R4039 gnd.n1857 gnd.n1856 585
R4040 gnd.n1858 gnd.n1857 585
R4041 gnd.n4145 gnd.n4144 585
R4042 gnd.n4146 gnd.n4145 585
R4043 gnd.n1867 gnd.n1866 585
R4044 gnd.n1866 gnd.n1864 585
R4045 gnd.n4140 gnd.n4139 585
R4046 gnd.n4139 gnd.n4138 585
R4047 gnd.n1870 gnd.n1869 585
R4048 gnd.n1878 gnd.n1870 585
R4049 gnd.n4129 gnd.n4128 585
R4050 gnd.n4130 gnd.n4129 585
R4051 gnd.n1880 gnd.n1879 585
R4052 gnd.n3494 gnd.n1879 585
R4053 gnd.n4124 gnd.n4123 585
R4054 gnd.n4123 gnd.n4122 585
R4055 gnd.n1883 gnd.n1882 585
R4056 gnd.n3489 gnd.n1883 585
R4057 gnd.n4113 gnd.n4112 585
R4058 gnd.n4114 gnd.n4113 585
R4059 gnd.n1893 gnd.n1892 585
R4060 gnd.n3477 gnd.n1892 585
R4061 gnd.n4108 gnd.n4107 585
R4062 gnd.n4107 gnd.n4106 585
R4063 gnd.n1896 gnd.n1895 585
R4064 gnd.n3470 gnd.n1896 585
R4065 gnd.n4097 gnd.n4096 585
R4066 gnd.n4098 gnd.n4097 585
R4067 gnd.n1907 gnd.n1906 585
R4068 gnd.n3722 gnd.n1906 585
R4069 gnd.n4092 gnd.n4091 585
R4070 gnd.n4091 gnd.n4090 585
R4071 gnd.n1910 gnd.n1909 585
R4072 gnd.n3456 gnd.n1910 585
R4073 gnd.n4081 gnd.n4080 585
R4074 gnd.n4082 gnd.n4081 585
R4075 gnd.n1920 gnd.n1919 585
R4076 gnd.n3737 gnd.n1919 585
R4077 gnd.n4076 gnd.n4075 585
R4078 gnd.n4075 gnd.n4074 585
R4079 gnd.n1923 gnd.n1922 585
R4080 gnd.n3443 gnd.n1923 585
R4081 gnd.n4065 gnd.n4064 585
R4082 gnd.n4066 gnd.n4065 585
R4083 gnd.n1932 gnd.n1931 585
R4084 gnd.n3752 gnd.n1931 585
R4085 gnd.n4060 gnd.n4059 585
R4086 gnd.n4059 gnd.n4058 585
R4087 gnd.n1935 gnd.n1934 585
R4088 gnd.n3428 gnd.n1935 585
R4089 gnd.n4049 gnd.n4048 585
R4090 gnd.n4050 gnd.n4049 585
R4091 gnd.n1945 gnd.n1944 585
R4092 gnd.n3767 gnd.n1944 585
R4093 gnd.n4044 gnd.n4043 585
R4094 gnd.n4043 gnd.n4042 585
R4095 gnd.n1948 gnd.n1947 585
R4096 gnd.n3415 gnd.n1948 585
R4097 gnd.n4033 gnd.n4032 585
R4098 gnd.n4034 gnd.n4033 585
R4099 gnd.n1960 gnd.n1959 585
R4100 gnd.n3782 gnd.n1959 585
R4101 gnd.n4028 gnd.n4027 585
R4102 gnd.n4027 gnd.n4026 585
R4103 gnd.n1963 gnd.n1962 585
R4104 gnd.n3403 gnd.n1963 585
R4105 gnd.n4017 gnd.n4016 585
R4106 gnd.n4018 gnd.n4017 585
R4107 gnd.n1974 gnd.n1973 585
R4108 gnd.n3396 gnd.n1973 585
R4109 gnd.n4012 gnd.n4011 585
R4110 gnd.n4011 gnd.n4010 585
R4111 gnd.n1977 gnd.n1976 585
R4112 gnd.n3389 gnd.n1977 585
R4113 gnd.n4001 gnd.n4000 585
R4114 gnd.n4002 gnd.n4001 585
R4115 gnd.n1989 gnd.n1988 585
R4116 gnd.n3382 gnd.n1988 585
R4117 gnd.n3996 gnd.n3995 585
R4118 gnd.n3995 gnd.n3994 585
R4119 gnd.n1992 gnd.n1991 585
R4120 gnd.n3375 gnd.n1992 585
R4121 gnd.n3985 gnd.n3984 585
R4122 gnd.n3986 gnd.n3985 585
R4123 gnd.n2004 gnd.n2003 585
R4124 gnd.n3368 gnd.n2003 585
R4125 gnd.n3980 gnd.n3979 585
R4126 gnd.n3979 gnd.n3978 585
R4127 gnd.n2007 gnd.n2006 585
R4128 gnd.n3361 gnd.n2007 585
R4129 gnd.n3969 gnd.n3968 585
R4130 gnd.n3970 gnd.n3969 585
R4131 gnd.n2019 gnd.n2018 585
R4132 gnd.n3838 gnd.n2018 585
R4133 gnd.n3964 gnd.n3963 585
R4134 gnd.n3963 gnd.n3962 585
R4135 gnd.n2022 gnd.n2021 585
R4136 gnd.n3349 gnd.n2022 585
R4137 gnd.n3953 gnd.n3952 585
R4138 gnd.n3954 gnd.n3953 585
R4139 gnd.n2033 gnd.n2032 585
R4140 gnd.n3852 gnd.n2032 585
R4141 gnd.n3948 gnd.n3947 585
R4142 gnd.n3947 gnd.n3946 585
R4143 gnd.n2036 gnd.n2035 585
R4144 gnd.n3334 gnd.n2036 585
R4145 gnd.n3937 gnd.n3936 585
R4146 gnd.n3938 gnd.n3937 585
R4147 gnd.n2048 gnd.n2047 585
R4148 gnd.n3867 gnd.n2047 585
R4149 gnd.n3932 gnd.n3931 585
R4150 gnd.n3931 gnd.n3930 585
R4151 gnd.n2051 gnd.n2050 585
R4152 gnd.n3321 gnd.n2051 585
R4153 gnd.n3921 gnd.n3920 585
R4154 gnd.n3922 gnd.n3921 585
R4155 gnd.n2063 gnd.n2062 585
R4156 gnd.n3882 gnd.n2062 585
R4157 gnd.n3916 gnd.n3915 585
R4158 gnd.n3915 gnd.n3914 585
R4159 gnd.n2066 gnd.n2065 585
R4160 gnd.n2090 gnd.n2066 585
R4161 gnd.n3905 gnd.n3904 585
R4162 gnd.n3906 gnd.n3905 585
R4163 gnd.n2078 gnd.n2077 585
R4164 gnd.n3307 gnd.n2077 585
R4165 gnd.n3900 gnd.n3899 585
R4166 gnd.n3899 gnd.n3898 585
R4167 gnd.n2081 gnd.n2080 585
R4168 gnd.n3301 gnd.n2081 585
R4169 gnd.n3289 gnd.n2105 585
R4170 gnd.n3022 gnd.n2105 585
R4171 gnd.n3291 gnd.n3290 585
R4172 gnd.n3292 gnd.n3291 585
R4173 gnd.n2106 gnd.n2104 585
R4174 gnd.n3035 gnd.n2104 585
R4175 gnd.n3284 gnd.n3283 585
R4176 gnd.n3283 gnd.n3282 585
R4177 gnd.n2109 gnd.n2108 585
R4178 gnd.n2904 gnd.n2109 585
R4179 gnd.n3273 gnd.n3272 585
R4180 gnd.n3274 gnd.n3273 585
R4181 gnd.n2118 gnd.n2117 585
R4182 gnd.n2122 gnd.n2117 585
R4183 gnd.n3268 gnd.n3267 585
R4184 gnd.n3267 gnd.n3266 585
R4185 gnd.n2121 gnd.n2120 585
R4186 gnd.n2131 gnd.n2121 585
R4187 gnd.n3257 gnd.n3256 585
R4188 gnd.n3258 gnd.n3257 585
R4189 gnd.n2133 gnd.n2132 585
R4190 gnd.n2132 gnd.n2129 585
R4191 gnd.n3252 gnd.n3251 585
R4192 gnd.n3251 gnd.n3250 585
R4193 gnd.n2136 gnd.n2135 585
R4194 gnd.n2144 gnd.n2136 585
R4195 gnd.n3241 gnd.n3240 585
R4196 gnd.n3242 gnd.n3241 585
R4197 gnd.n2146 gnd.n2145 585
R4198 gnd.n2145 gnd.n2142 585
R4199 gnd.n3236 gnd.n3235 585
R4200 gnd.n3235 gnd.n3234 585
R4201 gnd.n2149 gnd.n2148 585
R4202 gnd.n2151 gnd.n2149 585
R4203 gnd.n3225 gnd.n3224 585
R4204 gnd.n3226 gnd.n3225 585
R4205 gnd.n2159 gnd.n2158 585
R4206 gnd.n2158 gnd.n2157 585
R4207 gnd.n3220 gnd.n3219 585
R4208 gnd.n3219 gnd.n3218 585
R4209 gnd.n2162 gnd.n2161 585
R4210 gnd.n2164 gnd.n2162 585
R4211 gnd.n3209 gnd.n3208 585
R4212 gnd.n3210 gnd.n3209 585
R4213 gnd.n2171 gnd.n2170 585
R4214 gnd.n2176 gnd.n2170 585
R4215 gnd.n3204 gnd.n3203 585
R4216 gnd.n3203 gnd.n3202 585
R4217 gnd.n2174 gnd.n2173 585
R4218 gnd.n2175 gnd.n2174 585
R4219 gnd.n2756 gnd.n2755 585
R4220 gnd.n2756 gnd.n2181 585
R4221 gnd.n2759 gnd.n2758 585
R4222 gnd.n2758 gnd.n2757 585
R4223 gnd.n2760 gnd.n2749 585
R4224 gnd.n2749 gnd.n2265 585
R4225 gnd.n2762 gnd.n2761 585
R4226 gnd.n2762 gnd.n2249 585
R4227 gnd.n2763 gnd.n2748 585
R4228 gnd.n2763 gnd.n1273 585
R4229 gnd.n2765 gnd.n2764 585
R4230 gnd.n2764 gnd.n1270 585
R4231 gnd.n2766 gnd.n2743 585
R4232 gnd.n2743 gnd.n2331 585
R4233 gnd.n2768 gnd.n2767 585
R4234 gnd.n2768 gnd.n1261 585
R4235 gnd.n2769 gnd.n2742 585
R4236 gnd.n2769 gnd.n1253 585
R4237 gnd.n2771 gnd.n2770 585
R4238 gnd.n2770 gnd.n1250 585
R4239 gnd.n2772 gnd.n2344 585
R4240 gnd.n2344 gnd.n1242 585
R4241 gnd.n2774 gnd.n2773 585
R4242 gnd.n2775 gnd.n2774 585
R4243 gnd.n2345 gnd.n2343 585
R4244 gnd.n2343 gnd.n1232 585
R4245 gnd.n2736 gnd.n2735 585
R4246 gnd.n2735 gnd.n1229 585
R4247 gnd.n2734 gnd.n2347 585
R4248 gnd.n2734 gnd.n1221 585
R4249 gnd.n2733 gnd.n2732 585
R4250 gnd.n2733 gnd.n1218 585
R4251 gnd.n2349 gnd.n2348 585
R4252 gnd.n2696 gnd.n2348 585
R4253 gnd.n2728 gnd.n2727 585
R4254 gnd.n2727 gnd.n1208 585
R4255 gnd.n2726 gnd.n2351 585
R4256 gnd.n2726 gnd.n1200 585
R4257 gnd.n2725 gnd.n2353 585
R4258 gnd.n2725 gnd.n2724 585
R4259 gnd.n2391 gnd.n2352 585
R4260 gnd.n2352 gnd.n1190 585
R4261 gnd.n2393 gnd.n2392 585
R4262 gnd.n2392 gnd.n1187 585
R4263 gnd.n2394 gnd.n2385 585
R4264 gnd.n2385 gnd.n1179 585
R4265 gnd.n2396 gnd.n2395 585
R4266 gnd.n2396 gnd.n1176 585
R4267 gnd.n2397 gnd.n2384 585
R4268 gnd.n2397 gnd.n2371 585
R4269 gnd.n2399 gnd.n2398 585
R4270 gnd.n2398 gnd.n1166 585
R4271 gnd.n2382 gnd.n2380 585
R4272 gnd.n2380 gnd.n1159 585
R4273 gnd.n2657 gnd.n2656 585
R4274 gnd.n2658 gnd.n2657 585
R4275 gnd.n2381 gnd.n2379 585
R4276 gnd.n2379 gnd.n1149 585
R4277 gnd.n2607 gnd.n2606 585
R4278 gnd.n2606 gnd.n1146 585
R4279 gnd.n2609 gnd.n2608 585
R4280 gnd.n2609 gnd.n1141 585
R4281 gnd.n2611 gnd.n2610 585
R4282 gnd.n2610 gnd.n1138 585
R4283 gnd.n2613 gnd.n2612 585
R4284 gnd.n2614 gnd.n2613 585
R4285 gnd.n2605 gnd.n2604 585
R4286 gnd.n2605 gnd.n1128 585
R4287 gnd.n2603 gnd.n2413 585
R4288 gnd.n2413 gnd.n1122 585
R4289 gnd.n2650 gnd.n2407 585
R4290 gnd.n2650 gnd.n2649 585
R4291 gnd.n2652 gnd.n2651 585
R4292 gnd.n2651 gnd.n1112 585
R4293 gnd.n2412 gnd.n2406 585
R4294 gnd.n2412 gnd.n1109 585
R4295 gnd.n2411 gnd.n2410 585
R4296 gnd.n2411 gnd.n1101 585
R4297 gnd.n4509 gnd.n4508 585
R4298 gnd.n4508 gnd.n4507 585
R4299 gnd.n4510 gnd.n1404 585
R4300 gnd.n1406 gnd.n1404 585
R4301 gnd.n1824 gnd.n1402 585
R4302 gnd.n4199 gnd.n1824 585
R4303 gnd.n4514 gnd.n1401 585
R4304 gnd.n1823 gnd.n1401 585
R4305 gnd.n4515 gnd.n1400 585
R4306 gnd.n4188 gnd.n1400 585
R4307 gnd.n4516 gnd.n1399 585
R4308 gnd.n1831 gnd.n1399 585
R4309 gnd.n1838 gnd.n1397 585
R4310 gnd.n4178 gnd.n1838 585
R4311 gnd.n4520 gnd.n1396 585
R4312 gnd.n1845 gnd.n1396 585
R4313 gnd.n4521 gnd.n1395 585
R4314 gnd.n4170 gnd.n1395 585
R4315 gnd.n4522 gnd.n1394 585
R4316 gnd.n1844 gnd.n1394 585
R4317 gnd.n1852 gnd.n1392 585
R4318 gnd.n4162 gnd.n1852 585
R4319 gnd.n4526 gnd.n1391 585
R4320 gnd.n1851 gnd.n1391 585
R4321 gnd.n4527 gnd.n1390 585
R4322 gnd.n4154 gnd.n1390 585
R4323 gnd.n4528 gnd.n1389 585
R4324 gnd.n1858 gnd.n1389 585
R4325 gnd.n1865 gnd.n1387 585
R4326 gnd.n4146 gnd.n1865 585
R4327 gnd.n4532 gnd.n1386 585
R4328 gnd.n1864 gnd.n1386 585
R4329 gnd.n4533 gnd.n1385 585
R4330 gnd.n4138 gnd.n1385 585
R4331 gnd.n4534 gnd.n1384 585
R4332 gnd.n1878 gnd.n1384 585
R4333 gnd.n1877 gnd.n1382 585
R4334 gnd.n4130 gnd.n1877 585
R4335 gnd.n4538 gnd.n1381 585
R4336 gnd.n3494 gnd.n1381 585
R4337 gnd.n4539 gnd.n1380 585
R4338 gnd.n4122 gnd.n1380 585
R4339 gnd.n4540 gnd.n1379 585
R4340 gnd.n3489 gnd.n1379 585
R4341 gnd.n1891 gnd.n1377 585
R4342 gnd.n4114 gnd.n1891 585
R4343 gnd.n4544 gnd.n1376 585
R4344 gnd.n3477 gnd.n1376 585
R4345 gnd.n4545 gnd.n1375 585
R4346 gnd.n4106 gnd.n1375 585
R4347 gnd.n4546 gnd.n1374 585
R4348 gnd.n3470 gnd.n1374 585
R4349 gnd.n1905 gnd.n1372 585
R4350 gnd.n4098 gnd.n1905 585
R4351 gnd.n4550 gnd.n1371 585
R4352 gnd.n3722 gnd.n1371 585
R4353 gnd.n4551 gnd.n1370 585
R4354 gnd.n4090 gnd.n1370 585
R4355 gnd.n4552 gnd.n1369 585
R4356 gnd.n3456 gnd.n1369 585
R4357 gnd.n1918 gnd.n1367 585
R4358 gnd.n4082 gnd.n1918 585
R4359 gnd.n4556 gnd.n1366 585
R4360 gnd.n3737 gnd.n1366 585
R4361 gnd.n4557 gnd.n1365 585
R4362 gnd.n4074 gnd.n1365 585
R4363 gnd.n4558 gnd.n1364 585
R4364 gnd.n3443 gnd.n1364 585
R4365 gnd.n1930 gnd.n1362 585
R4366 gnd.n4066 gnd.n1930 585
R4367 gnd.n4562 gnd.n1361 585
R4368 gnd.n3752 gnd.n1361 585
R4369 gnd.n4563 gnd.n1360 585
R4370 gnd.n4058 gnd.n1360 585
R4371 gnd.n4564 gnd.n1359 585
R4372 gnd.n3428 gnd.n1359 585
R4373 gnd.n1942 gnd.n1357 585
R4374 gnd.n4050 gnd.n1942 585
R4375 gnd.n4568 gnd.n1356 585
R4376 gnd.n3767 gnd.n1356 585
R4377 gnd.n4569 gnd.n1355 585
R4378 gnd.n4042 gnd.n1355 585
R4379 gnd.n4570 gnd.n1354 585
R4380 gnd.n3415 gnd.n1354 585
R4381 gnd.n1956 gnd.n1352 585
R4382 gnd.n4034 gnd.n1956 585
R4383 gnd.n4574 gnd.n1351 585
R4384 gnd.n3782 gnd.n1351 585
R4385 gnd.n4575 gnd.n1350 585
R4386 gnd.n4026 gnd.n1350 585
R4387 gnd.n4576 gnd.n1349 585
R4388 gnd.n3403 gnd.n1349 585
R4389 gnd.n1971 gnd.n1347 585
R4390 gnd.n4018 gnd.n1971 585
R4391 gnd.n4580 gnd.n1346 585
R4392 gnd.n3396 gnd.n1346 585
R4393 gnd.n4581 gnd.n1345 585
R4394 gnd.n4010 gnd.n1345 585
R4395 gnd.n4582 gnd.n1344 585
R4396 gnd.n3389 gnd.n1344 585
R4397 gnd.n1986 gnd.n1342 585
R4398 gnd.n4002 gnd.n1986 585
R4399 gnd.n4586 gnd.n1341 585
R4400 gnd.n3382 gnd.n1341 585
R4401 gnd.n4587 gnd.n1340 585
R4402 gnd.n3994 gnd.n1340 585
R4403 gnd.n4588 gnd.n1339 585
R4404 gnd.n3375 gnd.n1339 585
R4405 gnd.n2001 gnd.n1337 585
R4406 gnd.n3986 gnd.n2001 585
R4407 gnd.n4592 gnd.n1336 585
R4408 gnd.n3368 gnd.n1336 585
R4409 gnd.n4593 gnd.n1335 585
R4410 gnd.n3978 gnd.n1335 585
R4411 gnd.n4594 gnd.n1334 585
R4412 gnd.n3361 gnd.n1334 585
R4413 gnd.n2016 gnd.n1332 585
R4414 gnd.n3970 gnd.n2016 585
R4415 gnd.n4598 gnd.n1331 585
R4416 gnd.n3838 gnd.n1331 585
R4417 gnd.n4599 gnd.n1330 585
R4418 gnd.n3962 gnd.n1330 585
R4419 gnd.n4600 gnd.n1329 585
R4420 gnd.n3349 gnd.n1329 585
R4421 gnd.n2030 gnd.n1327 585
R4422 gnd.n3954 gnd.n2030 585
R4423 gnd.n4604 gnd.n1326 585
R4424 gnd.n3852 gnd.n1326 585
R4425 gnd.n4605 gnd.n1325 585
R4426 gnd.n3946 gnd.n1325 585
R4427 gnd.n4606 gnd.n1324 585
R4428 gnd.n3334 gnd.n1324 585
R4429 gnd.n2045 gnd.n1322 585
R4430 gnd.n3938 gnd.n2045 585
R4431 gnd.n4610 gnd.n1321 585
R4432 gnd.n3867 gnd.n1321 585
R4433 gnd.n4611 gnd.n1320 585
R4434 gnd.n3930 gnd.n1320 585
R4435 gnd.n4612 gnd.n1319 585
R4436 gnd.n3321 gnd.n1319 585
R4437 gnd.n2060 gnd.n1317 585
R4438 gnd.n3922 gnd.n2060 585
R4439 gnd.n4616 gnd.n1316 585
R4440 gnd.n3882 gnd.n1316 585
R4441 gnd.n4617 gnd.n1315 585
R4442 gnd.n3914 gnd.n1315 585
R4443 gnd.n4618 gnd.n1314 585
R4444 gnd.n2090 gnd.n1314 585
R4445 gnd.n2075 gnd.n1312 585
R4446 gnd.n3906 gnd.n2075 585
R4447 gnd.n4622 gnd.n1311 585
R4448 gnd.n3307 gnd.n1311 585
R4449 gnd.n4623 gnd.n1310 585
R4450 gnd.n3898 gnd.n1310 585
R4451 gnd.n4624 gnd.n1309 585
R4452 gnd.n3301 gnd.n1309 585
R4453 gnd.n3021 gnd.n1307 585
R4454 gnd.n3022 gnd.n3021 585
R4455 gnd.n4628 gnd.n1306 585
R4456 gnd.n3292 gnd.n1306 585
R4457 gnd.n4629 gnd.n1305 585
R4458 gnd.n3035 gnd.n1305 585
R4459 gnd.n4630 gnd.n1304 585
R4460 gnd.n3282 gnd.n1304 585
R4461 gnd.n2903 gnd.n1302 585
R4462 gnd.n2904 gnd.n2903 585
R4463 gnd.n4634 gnd.n1301 585
R4464 gnd.n3274 gnd.n1301 585
R4465 gnd.n4635 gnd.n1300 585
R4466 gnd.n2122 gnd.n1300 585
R4467 gnd.n4636 gnd.n1299 585
R4468 gnd.n3266 gnd.n1299 585
R4469 gnd.n2130 gnd.n1297 585
R4470 gnd.n2131 gnd.n2130 585
R4471 gnd.n4640 gnd.n1296 585
R4472 gnd.n3258 gnd.n1296 585
R4473 gnd.n4641 gnd.n1295 585
R4474 gnd.n2129 gnd.n1295 585
R4475 gnd.n4642 gnd.n1294 585
R4476 gnd.n3250 gnd.n1294 585
R4477 gnd.n2143 gnd.n1292 585
R4478 gnd.n2144 gnd.n2143 585
R4479 gnd.n4646 gnd.n1291 585
R4480 gnd.n3242 gnd.n1291 585
R4481 gnd.n4647 gnd.n1290 585
R4482 gnd.n2142 gnd.n1290 585
R4483 gnd.n4648 gnd.n1289 585
R4484 gnd.n3234 gnd.n1289 585
R4485 gnd.n2150 gnd.n1287 585
R4486 gnd.n2151 gnd.n2150 585
R4487 gnd.n4652 gnd.n1286 585
R4488 gnd.n3226 gnd.n1286 585
R4489 gnd.n4653 gnd.n1285 585
R4490 gnd.n2157 gnd.n1285 585
R4491 gnd.n4654 gnd.n1284 585
R4492 gnd.n3218 gnd.n1284 585
R4493 gnd.n2163 gnd.n1282 585
R4494 gnd.n2164 gnd.n2163 585
R4495 gnd.n4658 gnd.n1281 585
R4496 gnd.n3210 gnd.n1281 585
R4497 gnd.n4659 gnd.n1280 585
R4498 gnd.n2176 gnd.n1280 585
R4499 gnd.n4660 gnd.n1279 585
R4500 gnd.n3202 gnd.n1279 585
R4501 gnd.n3191 gnd.n3190 585
R4502 gnd.n3189 gnd.n2195 585
R4503 gnd.n2197 gnd.n2194 585
R4504 gnd.n3193 gnd.n2194 585
R4505 gnd.n3182 gnd.n2205 585
R4506 gnd.n3181 gnd.n2206 585
R4507 gnd.n2208 gnd.n2207 585
R4508 gnd.n3174 gnd.n2214 585
R4509 gnd.n3173 gnd.n2215 585
R4510 gnd.n2222 gnd.n2216 585
R4511 gnd.n3166 gnd.n2223 585
R4512 gnd.n3165 gnd.n2224 585
R4513 gnd.n2226 gnd.n2225 585
R4514 gnd.n3158 gnd.n2232 585
R4515 gnd.n3157 gnd.n2233 585
R4516 gnd.n2242 gnd.n2234 585
R4517 gnd.n3150 gnd.n2243 585
R4518 gnd.n3149 gnd.n2244 585
R4519 gnd.n2246 gnd.n2245 585
R4520 gnd.n2824 gnd.n2799 585
R4521 gnd.n2823 gnd.n2800 585
R4522 gnd.n2822 gnd.n2801 585
R4523 gnd.n2803 gnd.n2802 585
R4524 gnd.n2818 gnd.n2805 585
R4525 gnd.n2817 gnd.n2806 585
R4526 gnd.n2816 gnd.n2807 585
R4527 gnd.n2813 gnd.n2812 585
R4528 gnd.n2180 gnd.n2179 585
R4529 gnd.n3196 gnd.n3195 585
R4530 gnd.n3197 gnd.n2177 585
R4531 gnd.n4203 gnd.n1408 585
R4532 gnd.n4507 gnd.n1408 585
R4533 gnd.n4202 gnd.n4201 585
R4534 gnd.n4201 gnd.n1406 585
R4535 gnd.n4200 gnd.n1821 585
R4536 gnd.n4200 gnd.n4199 585
R4537 gnd.n1834 gnd.n1822 585
R4538 gnd.n1823 gnd.n1822 585
R4539 gnd.n4187 gnd.n4186 585
R4540 gnd.n4188 gnd.n4187 585
R4541 gnd.n1833 gnd.n1832 585
R4542 gnd.n1832 gnd.n1831 585
R4543 gnd.n4180 gnd.n4179 585
R4544 gnd.n4179 gnd.n4178 585
R4545 gnd.n1837 gnd.n1836 585
R4546 gnd.n1845 gnd.n1837 585
R4547 gnd.n4169 gnd.n4168 585
R4548 gnd.n4170 gnd.n4169 585
R4549 gnd.n1847 gnd.n1846 585
R4550 gnd.n1846 gnd.n1844 585
R4551 gnd.n4164 gnd.n4163 585
R4552 gnd.n4163 gnd.n4162 585
R4553 gnd.n1850 gnd.n1849 585
R4554 gnd.n1851 gnd.n1850 585
R4555 gnd.n4153 gnd.n4152 585
R4556 gnd.n4154 gnd.n4153 585
R4557 gnd.n1860 gnd.n1859 585
R4558 gnd.n1859 gnd.n1858 585
R4559 gnd.n4148 gnd.n4147 585
R4560 gnd.n4147 gnd.n4146 585
R4561 gnd.n1863 gnd.n1862 585
R4562 gnd.n1864 gnd.n1863 585
R4563 gnd.n4137 gnd.n4136 585
R4564 gnd.n4138 gnd.n4137 585
R4565 gnd.n1872 gnd.n1871 585
R4566 gnd.n1878 gnd.n1871 585
R4567 gnd.n4132 gnd.n4131 585
R4568 gnd.n4131 gnd.n4130 585
R4569 gnd.n1875 gnd.n1874 585
R4570 gnd.n3494 gnd.n1875 585
R4571 gnd.n4121 gnd.n4120 585
R4572 gnd.n4122 gnd.n4121 585
R4573 gnd.n1886 gnd.n1885 585
R4574 gnd.n3489 gnd.n1885 585
R4575 gnd.n4116 gnd.n4115 585
R4576 gnd.n4115 gnd.n4114 585
R4577 gnd.n1889 gnd.n1888 585
R4578 gnd.n3477 gnd.n1889 585
R4579 gnd.n4105 gnd.n4104 585
R4580 gnd.n4106 gnd.n4105 585
R4581 gnd.n1900 gnd.n1899 585
R4582 gnd.n3470 gnd.n1899 585
R4583 gnd.n4100 gnd.n4099 585
R4584 gnd.n4099 gnd.n4098 585
R4585 gnd.n1903 gnd.n1902 585
R4586 gnd.n3722 gnd.n1903 585
R4587 gnd.n4089 gnd.n4088 585
R4588 gnd.n4090 gnd.n4089 585
R4589 gnd.n1913 gnd.n1912 585
R4590 gnd.n3456 gnd.n1912 585
R4591 gnd.n4084 gnd.n4083 585
R4592 gnd.n4083 gnd.n4082 585
R4593 gnd.n1916 gnd.n1915 585
R4594 gnd.n3737 gnd.n1916 585
R4595 gnd.n4073 gnd.n4072 585
R4596 gnd.n4074 gnd.n4073 585
R4597 gnd.n1926 gnd.n1925 585
R4598 gnd.n3443 gnd.n1925 585
R4599 gnd.n4068 gnd.n4067 585
R4600 gnd.n4067 gnd.n4066 585
R4601 gnd.n1929 gnd.n1928 585
R4602 gnd.n3752 gnd.n1929 585
R4603 gnd.n4057 gnd.n4056 585
R4604 gnd.n4058 gnd.n4057 585
R4605 gnd.n1938 gnd.n1937 585
R4606 gnd.n3428 gnd.n1937 585
R4607 gnd.n4052 gnd.n4051 585
R4608 gnd.n4051 gnd.n4050 585
R4609 gnd.n1941 gnd.n1940 585
R4610 gnd.n3767 gnd.n1941 585
R4611 gnd.n4041 gnd.n4040 585
R4612 gnd.n4042 gnd.n4041 585
R4613 gnd.n1951 gnd.n1950 585
R4614 gnd.n3415 gnd.n1950 585
R4615 gnd.n4036 gnd.n4035 585
R4616 gnd.n4035 gnd.n4034 585
R4617 gnd.n1954 gnd.n1953 585
R4618 gnd.n3782 gnd.n1954 585
R4619 gnd.n4025 gnd.n4024 585
R4620 gnd.n4026 gnd.n4025 585
R4621 gnd.n1966 gnd.n1965 585
R4622 gnd.n3403 gnd.n1965 585
R4623 gnd.n4020 gnd.n4019 585
R4624 gnd.n4019 gnd.n4018 585
R4625 gnd.n1969 gnd.n1968 585
R4626 gnd.n3396 gnd.n1969 585
R4627 gnd.n4009 gnd.n4008 585
R4628 gnd.n4010 gnd.n4009 585
R4629 gnd.n1981 gnd.n1980 585
R4630 gnd.n3389 gnd.n1980 585
R4631 gnd.n4004 gnd.n4003 585
R4632 gnd.n4003 gnd.n4002 585
R4633 gnd.n1984 gnd.n1983 585
R4634 gnd.n3382 gnd.n1984 585
R4635 gnd.n3993 gnd.n3992 585
R4636 gnd.n3994 gnd.n3993 585
R4637 gnd.n1996 gnd.n1995 585
R4638 gnd.n3375 gnd.n1995 585
R4639 gnd.n3988 gnd.n3987 585
R4640 gnd.n3987 gnd.n3986 585
R4641 gnd.n1999 gnd.n1998 585
R4642 gnd.n3368 gnd.n1999 585
R4643 gnd.n3977 gnd.n3976 585
R4644 gnd.n3978 gnd.n3977 585
R4645 gnd.n2011 gnd.n2010 585
R4646 gnd.n3361 gnd.n2010 585
R4647 gnd.n3972 gnd.n3971 585
R4648 gnd.n3971 gnd.n3970 585
R4649 gnd.n2014 gnd.n2013 585
R4650 gnd.n3838 gnd.n2014 585
R4651 gnd.n3961 gnd.n3960 585
R4652 gnd.n3962 gnd.n3961 585
R4653 gnd.n2026 gnd.n2025 585
R4654 gnd.n3349 gnd.n2025 585
R4655 gnd.n3956 gnd.n3955 585
R4656 gnd.n3955 gnd.n3954 585
R4657 gnd.n2029 gnd.n2028 585
R4658 gnd.n3852 gnd.n2029 585
R4659 gnd.n3945 gnd.n3944 585
R4660 gnd.n3946 gnd.n3945 585
R4661 gnd.n2040 gnd.n2039 585
R4662 gnd.n3334 gnd.n2039 585
R4663 gnd.n3940 gnd.n3939 585
R4664 gnd.n3939 gnd.n3938 585
R4665 gnd.n2043 gnd.n2042 585
R4666 gnd.n3867 gnd.n2043 585
R4667 gnd.n3929 gnd.n3928 585
R4668 gnd.n3930 gnd.n3929 585
R4669 gnd.n2055 gnd.n2054 585
R4670 gnd.n3321 gnd.n2054 585
R4671 gnd.n3924 gnd.n3923 585
R4672 gnd.n3923 gnd.n3922 585
R4673 gnd.n2058 gnd.n2057 585
R4674 gnd.n3882 gnd.n2058 585
R4675 gnd.n3913 gnd.n3912 585
R4676 gnd.n3914 gnd.n3913 585
R4677 gnd.n2070 gnd.n2069 585
R4678 gnd.n2090 gnd.n2069 585
R4679 gnd.n3908 gnd.n3907 585
R4680 gnd.n3907 gnd.n3906 585
R4681 gnd.n2073 gnd.n2072 585
R4682 gnd.n3307 gnd.n2073 585
R4683 gnd.n2098 gnd.n2083 585
R4684 gnd.n3898 gnd.n2083 585
R4685 gnd.n3300 gnd.n3299 585
R4686 gnd.n3301 gnd.n3300 585
R4687 gnd.n2097 gnd.n2096 585
R4688 gnd.n3022 gnd.n2096 585
R4689 gnd.n3294 gnd.n3293 585
R4690 gnd.n3293 gnd.n3292 585
R4691 gnd.n2101 gnd.n2100 585
R4692 gnd.n3035 gnd.n2101 585
R4693 gnd.n3281 gnd.n3280 585
R4694 gnd.n3282 gnd.n3281 585
R4695 gnd.n2112 gnd.n2111 585
R4696 gnd.n2904 gnd.n2111 585
R4697 gnd.n3276 gnd.n3275 585
R4698 gnd.n3275 gnd.n3274 585
R4699 gnd.n2115 gnd.n2114 585
R4700 gnd.n2122 gnd.n2115 585
R4701 gnd.n3265 gnd.n3264 585
R4702 gnd.n3266 gnd.n3265 585
R4703 gnd.n2125 gnd.n2124 585
R4704 gnd.n2131 gnd.n2124 585
R4705 gnd.n3260 gnd.n3259 585
R4706 gnd.n3259 gnd.n3258 585
R4707 gnd.n2128 gnd.n2127 585
R4708 gnd.n2129 gnd.n2128 585
R4709 gnd.n3249 gnd.n3248 585
R4710 gnd.n3250 gnd.n3249 585
R4711 gnd.n2138 gnd.n2137 585
R4712 gnd.n2144 gnd.n2137 585
R4713 gnd.n3244 gnd.n3243 585
R4714 gnd.n3243 gnd.n3242 585
R4715 gnd.n2141 gnd.n2140 585
R4716 gnd.n2142 gnd.n2141 585
R4717 gnd.n3233 gnd.n3232 585
R4718 gnd.n3234 gnd.n3233 585
R4719 gnd.n2153 gnd.n2152 585
R4720 gnd.n2152 gnd.n2151 585
R4721 gnd.n3228 gnd.n3227 585
R4722 gnd.n3227 gnd.n3226 585
R4723 gnd.n2156 gnd.n2155 585
R4724 gnd.n2157 gnd.n2156 585
R4725 gnd.n3217 gnd.n3216 585
R4726 gnd.n3218 gnd.n3217 585
R4727 gnd.n2166 gnd.n2165 585
R4728 gnd.n2165 gnd.n2164 585
R4729 gnd.n3212 gnd.n3211 585
R4730 gnd.n3211 gnd.n3210 585
R4731 gnd.n2169 gnd.n2168 585
R4732 gnd.n2176 gnd.n2169 585
R4733 gnd.n3201 gnd.n3200 585
R4734 gnd.n3202 gnd.n3201 585
R4735 gnd.n4210 gnd.n4209 585
R4736 gnd.n4209 gnd.n1409 585
R4737 gnd.n4211 gnd.n4208 585
R4738 gnd.n4206 gnd.n1819 585
R4739 gnd.n4215 gnd.n1818 585
R4740 gnd.n4219 gnd.n1816 585
R4741 gnd.n4220 gnd.n1815 585
R4742 gnd.n1813 gnd.n1811 585
R4743 gnd.n4224 gnd.n1810 585
R4744 gnd.n4225 gnd.n1808 585
R4745 gnd.n4226 gnd.n1807 585
R4746 gnd.n1805 gnd.n1685 585
R4747 gnd.n1804 gnd.n1803 585
R4748 gnd.n1793 gnd.n1687 585
R4749 gnd.n1795 gnd.n1794 585
R4750 gnd.n1791 gnd.n1697 585
R4751 gnd.n1790 gnd.n1789 585
R4752 gnd.n1777 gnd.n1699 585
R4753 gnd.n1779 gnd.n1778 585
R4754 gnd.n1775 gnd.n1703 585
R4755 gnd.n1774 gnd.n1773 585
R4756 gnd.n1758 gnd.n1705 585
R4757 gnd.n1760 gnd.n1759 585
R4758 gnd.n1756 gnd.n1710 585
R4759 gnd.n1755 gnd.n1754 585
R4760 gnd.n1739 gnd.n1712 585
R4761 gnd.n1741 gnd.n1740 585
R4762 gnd.n1737 gnd.n1717 585
R4763 gnd.n1736 gnd.n1735 585
R4764 gnd.n1719 gnd.n1405 585
R4765 gnd.n3684 gnd.n3495 482.89
R4766 gnd.n3567 gnd.n3493 482.89
R4767 gnd.n3047 gnd.n3045 482.89
R4768 gnd.n3008 gnd.n2905 482.89
R4769 gnd.n2884 gnd.t124 443.966
R4770 gnd.n3543 gnd.t137 443.966
R4771 gnd.n2942 gnd.t165 443.966
R4772 gnd.n3537 gnd.t90 443.966
R4773 gnd.n6500 gnd.n6499 404.397
R4774 gnd.n2808 gnd.t114 371.625
R4775 gnd.n7404 gnd.t140 371.625
R4776 gnd.n1691 gnd.t131 371.625
R4777 gnd.n2238 gnd.t153 371.625
R4778 gnd.n1469 gnd.t101 371.625
R4779 gnd.n1491 gnd.t94 371.625
R4780 gnd.n179 gnd.t159 371.625
R4781 gnd.n7497 gnd.t83 371.625
R4782 gnd.n983 gnd.t63 371.625
R4783 gnd.n1005 gnd.t150 371.625
R4784 gnd.n2327 gnd.t156 371.625
R4785 gnd.n2305 gnd.t75 371.625
R4786 gnd.n2492 gnd.t104 371.625
R4787 gnd.n4216 gnd.t71 371.625
R4788 gnd.n5285 gnd.t146 323.425
R4789 gnd.n4936 gnd.t79 323.425
R4790 gnd.n6152 gnd.n6126 289.615
R4791 gnd.n6120 gnd.n6094 289.615
R4792 gnd.n6088 gnd.n6062 289.615
R4793 gnd.n6057 gnd.n6031 289.615
R4794 gnd.n6025 gnd.n5999 289.615
R4795 gnd.n5993 gnd.n5967 289.615
R4796 gnd.n5961 gnd.n5935 289.615
R4797 gnd.n5930 gnd.n5904 289.615
R4798 gnd.n5359 gnd.t107 279.217
R4799 gnd.n4980 gnd.t67 279.217
R4800 gnd.n2914 gnd.t145 260.649
R4801 gnd.n3507 gnd.t89 260.649
R4802 gnd.n3007 gnd.n2123 256.663
R4803 gnd.n3000 gnd.n2123 256.663
R4804 gnd.n2998 gnd.n2123 256.663
R4805 gnd.n2992 gnd.n2123 256.663
R4806 gnd.n2990 gnd.n2123 256.663
R4807 gnd.n2984 gnd.n2123 256.663
R4808 gnd.n2982 gnd.n2123 256.663
R4809 gnd.n2976 gnd.n2123 256.663
R4810 gnd.n2974 gnd.n2123 256.663
R4811 gnd.n2968 gnd.n2123 256.663
R4812 gnd.n2966 gnd.n2123 256.663
R4813 gnd.n2960 gnd.n2123 256.663
R4814 gnd.n2958 gnd.n2123 256.663
R4815 gnd.n2952 gnd.n2123 256.663
R4816 gnd.n2945 gnd.n2123 256.663
R4817 gnd.n2946 gnd.n2123 256.663
R4818 gnd.n3113 gnd.n2882 256.663
R4819 gnd.n3111 gnd.n2123 256.663
R4820 gnd.n3109 gnd.n2123 256.663
R4821 gnd.n3102 gnd.n2123 256.663
R4822 gnd.n3100 gnd.n2123 256.663
R4823 gnd.n3094 gnd.n2123 256.663
R4824 gnd.n3092 gnd.n2123 256.663
R4825 gnd.n3086 gnd.n2123 256.663
R4826 gnd.n3084 gnd.n2123 256.663
R4827 gnd.n3078 gnd.n2123 256.663
R4828 gnd.n3076 gnd.n2123 256.663
R4829 gnd.n3070 gnd.n2123 256.663
R4830 gnd.n3068 gnd.n2123 256.663
R4831 gnd.n3062 gnd.n2123 256.663
R4832 gnd.n3060 gnd.n2123 256.663
R4833 gnd.n3054 gnd.n2123 256.663
R4834 gnd.n3052 gnd.n2123 256.663
R4835 gnd.n3046 gnd.n2123 256.663
R4836 gnd.n3566 gnd.n3516 256.663
R4837 gnd.n3572 gnd.n3516 256.663
R4838 gnd.n3564 gnd.n3516 256.663
R4839 gnd.n3579 gnd.n3516 256.663
R4840 gnd.n3561 gnd.n3516 256.663
R4841 gnd.n3586 gnd.n3516 256.663
R4842 gnd.n3558 gnd.n3516 256.663
R4843 gnd.n3593 gnd.n3516 256.663
R4844 gnd.n3555 gnd.n3516 256.663
R4845 gnd.n3600 gnd.n3516 256.663
R4846 gnd.n3552 gnd.n3516 256.663
R4847 gnd.n3607 gnd.n3516 256.663
R4848 gnd.n3549 gnd.n3516 256.663
R4849 gnd.n3614 gnd.n3516 256.663
R4850 gnd.n3546 gnd.n3516 256.663
R4851 gnd.n3622 gnd.n3516 256.663
R4852 gnd.n3625 gnd.n1466 256.663
R4853 gnd.n3626 gnd.n3516 256.663
R4854 gnd.n3630 gnd.n3516 256.663
R4855 gnd.n3540 gnd.n3516 256.663
R4856 gnd.n3638 gnd.n3516 256.663
R4857 gnd.n3535 gnd.n3516 256.663
R4858 gnd.n3645 gnd.n3516 256.663
R4859 gnd.n3532 gnd.n3516 256.663
R4860 gnd.n3652 gnd.n3516 256.663
R4861 gnd.n3529 gnd.n3516 256.663
R4862 gnd.n3659 gnd.n3516 256.663
R4863 gnd.n3526 gnd.n3516 256.663
R4864 gnd.n3666 gnd.n3516 256.663
R4865 gnd.n3523 gnd.n3516 256.663
R4866 gnd.n3673 gnd.n3516 256.663
R4867 gnd.n3520 gnd.n3516 256.663
R4868 gnd.n3680 gnd.n3516 256.663
R4869 gnd.n3683 gnd.n3516 256.663
R4870 gnd.n4905 gnd.n951 242.672
R4871 gnd.n4905 gnd.n952 242.672
R4872 gnd.n4905 gnd.n953 242.672
R4873 gnd.n4905 gnd.n954 242.672
R4874 gnd.n4905 gnd.n955 242.672
R4875 gnd.n4905 gnd.n956 242.672
R4876 gnd.n4905 gnd.n957 242.672
R4877 gnd.n4905 gnd.n958 242.672
R4878 gnd.n4905 gnd.n959 242.672
R4879 gnd.n3144 gnd.n3143 242.672
R4880 gnd.n3143 gnd.n2264 242.672
R4881 gnd.n3143 gnd.n2263 242.672
R4882 gnd.n3143 gnd.n2261 242.672
R4883 gnd.n3143 gnd.n2259 242.672
R4884 gnd.n3143 gnd.n2258 242.672
R4885 gnd.n3143 gnd.n2256 242.672
R4886 gnd.n3143 gnd.n2254 242.672
R4887 gnd.n3143 gnd.n2253 242.672
R4888 gnd.n4498 gnd.n1436 242.672
R4889 gnd.n4498 gnd.n1437 242.672
R4890 gnd.n4498 gnd.n1438 242.672
R4891 gnd.n4498 gnd.n1439 242.672
R4892 gnd.n4498 gnd.n1440 242.672
R4893 gnd.n4498 gnd.n1441 242.672
R4894 gnd.n4498 gnd.n1442 242.672
R4895 gnd.n4498 gnd.n1443 242.672
R4896 gnd.n4498 gnd.n1444 242.672
R4897 gnd.n7406 gnd.n106 242.672
R4898 gnd.n7402 gnd.n106 242.672
R4899 gnd.n7397 gnd.n106 242.672
R4900 gnd.n7394 gnd.n106 242.672
R4901 gnd.n7389 gnd.n106 242.672
R4902 gnd.n7386 gnd.n106 242.672
R4903 gnd.n7381 gnd.n106 242.672
R4904 gnd.n7378 gnd.n106 242.672
R4905 gnd.n7373 gnd.n106 242.672
R4906 gnd.n5413 gnd.n5412 242.672
R4907 gnd.n5413 gnd.n5323 242.672
R4908 gnd.n5413 gnd.n5324 242.672
R4909 gnd.n5413 gnd.n5325 242.672
R4910 gnd.n5413 gnd.n5326 242.672
R4911 gnd.n5413 gnd.n5327 242.672
R4912 gnd.n5413 gnd.n5328 242.672
R4913 gnd.n5413 gnd.n5329 242.672
R4914 gnd.n5413 gnd.n5330 242.672
R4915 gnd.n5413 gnd.n5331 242.672
R4916 gnd.n5413 gnd.n5332 242.672
R4917 gnd.n5413 gnd.n5333 242.672
R4918 gnd.n5414 gnd.n5413 242.672
R4919 gnd.n6226 gnd.n4906 242.672
R4920 gnd.n6232 gnd.n4906 242.672
R4921 gnd.n4983 gnd.n4906 242.672
R4922 gnd.n6239 gnd.n4906 242.672
R4923 gnd.n4974 gnd.n4906 242.672
R4924 gnd.n6246 gnd.n4906 242.672
R4925 gnd.n4967 gnd.n4906 242.672
R4926 gnd.n6253 gnd.n4906 242.672
R4927 gnd.n4960 gnd.n4906 242.672
R4928 gnd.n6260 gnd.n4906 242.672
R4929 gnd.n4953 gnd.n4906 242.672
R4930 gnd.n6267 gnd.n4906 242.672
R4931 gnd.n4946 gnd.n4906 242.672
R4932 gnd.n5583 gnd.n5582 242.672
R4933 gnd.n5582 gnd.n5235 242.672
R4934 gnd.n5582 gnd.n5236 242.672
R4935 gnd.n5582 gnd.n5237 242.672
R4936 gnd.n5582 gnd.n5238 242.672
R4937 gnd.n5582 gnd.n5239 242.672
R4938 gnd.n5582 gnd.n5240 242.672
R4939 gnd.n5582 gnd.n5241 242.672
R4940 gnd.n6278 gnd.n4906 242.672
R4941 gnd.n4939 gnd.n4906 242.672
R4942 gnd.n6285 gnd.n4906 242.672
R4943 gnd.n4930 gnd.n4906 242.672
R4944 gnd.n6292 gnd.n4906 242.672
R4945 gnd.n4923 gnd.n4906 242.672
R4946 gnd.n6299 gnd.n4906 242.672
R4947 gnd.n4916 gnd.n4906 242.672
R4948 gnd.n4905 gnd.n4904 242.672
R4949 gnd.n4905 gnd.n933 242.672
R4950 gnd.n4905 gnd.n934 242.672
R4951 gnd.n4905 gnd.n935 242.672
R4952 gnd.n4905 gnd.n936 242.672
R4953 gnd.n4905 gnd.n937 242.672
R4954 gnd.n4905 gnd.n938 242.672
R4955 gnd.n4905 gnd.n939 242.672
R4956 gnd.n4905 gnd.n940 242.672
R4957 gnd.n4905 gnd.n941 242.672
R4958 gnd.n4905 gnd.n942 242.672
R4959 gnd.n4905 gnd.n943 242.672
R4960 gnd.n4905 gnd.n944 242.672
R4961 gnd.n4905 gnd.n945 242.672
R4962 gnd.n4905 gnd.n946 242.672
R4963 gnd.n4905 gnd.n947 242.672
R4964 gnd.n4905 gnd.n948 242.672
R4965 gnd.n4905 gnd.n949 242.672
R4966 gnd.n4905 gnd.n950 242.672
R4967 gnd.n3143 gnd.n2266 242.672
R4968 gnd.n3143 gnd.n2267 242.672
R4969 gnd.n3143 gnd.n2268 242.672
R4970 gnd.n3143 gnd.n2269 242.672
R4971 gnd.n3143 gnd.n2270 242.672
R4972 gnd.n3143 gnd.n2271 242.672
R4973 gnd.n3143 gnd.n2272 242.672
R4974 gnd.n3143 gnd.n2273 242.672
R4975 gnd.n3143 gnd.n2274 242.672
R4976 gnd.n3143 gnd.n2275 242.672
R4977 gnd.n3143 gnd.n2276 242.672
R4978 gnd.n3114 gnd.n2307 242.672
R4979 gnd.n3143 gnd.n2277 242.672
R4980 gnd.n3143 gnd.n2278 242.672
R4981 gnd.n3143 gnd.n2279 242.672
R4982 gnd.n3143 gnd.n2280 242.672
R4983 gnd.n3143 gnd.n2281 242.672
R4984 gnd.n3143 gnd.n2282 242.672
R4985 gnd.n3143 gnd.n2283 242.672
R4986 gnd.n3143 gnd.n3142 242.672
R4987 gnd.n4498 gnd.n4497 242.672
R4988 gnd.n4498 gnd.n1418 242.672
R4989 gnd.n4498 gnd.n1419 242.672
R4990 gnd.n4498 gnd.n1420 242.672
R4991 gnd.n4498 gnd.n1421 242.672
R4992 gnd.n4498 gnd.n1422 242.672
R4993 gnd.n4498 gnd.n1423 242.672
R4994 gnd.n4498 gnd.n1424 242.672
R4995 gnd.n4466 gnd.n1467 242.672
R4996 gnd.n4498 gnd.n1425 242.672
R4997 gnd.n4498 gnd.n1426 242.672
R4998 gnd.n4498 gnd.n1427 242.672
R4999 gnd.n4498 gnd.n1428 242.672
R5000 gnd.n4498 gnd.n1429 242.672
R5001 gnd.n4498 gnd.n1430 242.672
R5002 gnd.n4498 gnd.n1431 242.672
R5003 gnd.n4498 gnd.n1432 242.672
R5004 gnd.n4498 gnd.n1433 242.672
R5005 gnd.n4498 gnd.n1434 242.672
R5006 gnd.n4498 gnd.n1435 242.672
R5007 gnd.n176 gnd.n106 242.672
R5008 gnd.n7465 gnd.n106 242.672
R5009 gnd.n172 gnd.n106 242.672
R5010 gnd.n7472 gnd.n106 242.672
R5011 gnd.n165 gnd.n106 242.672
R5012 gnd.n7479 gnd.n106 242.672
R5013 gnd.n158 gnd.n106 242.672
R5014 gnd.n7486 gnd.n106 242.672
R5015 gnd.n151 gnd.n106 242.672
R5016 gnd.n7493 gnd.n106 242.672
R5017 gnd.n144 gnd.n106 242.672
R5018 gnd.n7503 gnd.n106 242.672
R5019 gnd.n137 gnd.n106 242.672
R5020 gnd.n7510 gnd.n106 242.672
R5021 gnd.n130 gnd.n106 242.672
R5022 gnd.n7517 gnd.n106 242.672
R5023 gnd.n123 gnd.n106 242.672
R5024 gnd.n7524 gnd.n106 242.672
R5025 gnd.n116 gnd.n106 242.672
R5026 gnd.n3193 gnd.n3192 242.672
R5027 gnd.n3193 gnd.n2182 242.672
R5028 gnd.n3193 gnd.n2183 242.672
R5029 gnd.n3193 gnd.n2184 242.672
R5030 gnd.n3193 gnd.n2185 242.672
R5031 gnd.n3193 gnd.n2186 242.672
R5032 gnd.n3193 gnd.n2187 242.672
R5033 gnd.n3193 gnd.n2188 242.672
R5034 gnd.n3193 gnd.n2189 242.672
R5035 gnd.n3193 gnd.n2190 242.672
R5036 gnd.n3193 gnd.n2191 242.672
R5037 gnd.n3193 gnd.n2192 242.672
R5038 gnd.n3193 gnd.n2193 242.672
R5039 gnd.n3194 gnd.n3193 242.672
R5040 gnd.n4207 gnd.n1409 242.672
R5041 gnd.n1817 gnd.n1409 242.672
R5042 gnd.n1814 gnd.n1409 242.672
R5043 gnd.n1809 gnd.n1409 242.672
R5044 gnd.n1806 gnd.n1409 242.672
R5045 gnd.n1686 gnd.n1409 242.672
R5046 gnd.n1792 gnd.n1409 242.672
R5047 gnd.n1698 gnd.n1409 242.672
R5048 gnd.n1776 gnd.n1409 242.672
R5049 gnd.n1704 gnd.n1409 242.672
R5050 gnd.n1757 gnd.n1409 242.672
R5051 gnd.n1711 gnd.n1409 242.672
R5052 gnd.n1738 gnd.n1409 242.672
R5053 gnd.n1718 gnd.n1409 242.672
R5054 gnd.n113 gnd.n109 240.244
R5055 gnd.n7526 gnd.n7525 240.244
R5056 gnd.n7523 gnd.n117 240.244
R5057 gnd.n7519 gnd.n7518 240.244
R5058 gnd.n7516 gnd.n124 240.244
R5059 gnd.n7512 gnd.n7511 240.244
R5060 gnd.n7509 gnd.n131 240.244
R5061 gnd.n7505 gnd.n7504 240.244
R5062 gnd.n7502 gnd.n138 240.244
R5063 gnd.n7495 gnd.n7494 240.244
R5064 gnd.n7492 gnd.n145 240.244
R5065 gnd.n7488 gnd.n7487 240.244
R5066 gnd.n7485 gnd.n152 240.244
R5067 gnd.n7481 gnd.n7480 240.244
R5068 gnd.n7478 gnd.n159 240.244
R5069 gnd.n7474 gnd.n7473 240.244
R5070 gnd.n7471 gnd.n166 240.244
R5071 gnd.n7467 gnd.n7466 240.244
R5072 gnd.n7464 gnd.n173 240.244
R5073 gnd.n4423 gnd.n1495 240.244
R5074 gnd.n1679 gnd.n1495 240.244
R5075 gnd.n1679 gnd.n1626 240.244
R5076 gnd.n1675 gnd.n1626 240.244
R5077 gnd.n1675 gnd.n1616 240.244
R5078 gnd.n1672 gnd.n1616 240.244
R5079 gnd.n1672 gnd.n1608 240.244
R5080 gnd.n1608 gnd.n1598 240.244
R5081 gnd.n1667 gnd.n1598 240.244
R5082 gnd.n1667 gnd.n1589 240.244
R5083 gnd.n1664 gnd.n1589 240.244
R5084 gnd.n1664 gnd.n1581 240.244
R5085 gnd.n1581 gnd.n1571 240.244
R5086 gnd.n1571 gnd.n1559 240.244
R5087 gnd.n4327 gnd.n1559 240.244
R5088 gnd.n4327 gnd.n1560 240.244
R5089 gnd.n1560 gnd.n1547 240.244
R5090 gnd.n1547 gnd.n1536 240.244
R5091 gnd.n4334 gnd.n1536 240.244
R5092 gnd.n4334 gnd.n1527 240.244
R5093 gnd.n4348 gnd.n1527 240.244
R5094 gnd.n4348 gnd.n279 240.244
R5095 gnd.n313 gnd.n279 240.244
R5096 gnd.n4343 gnd.n313 240.244
R5097 gnd.n4343 gnd.n301 240.244
R5098 gnd.n7206 gnd.n301 240.244
R5099 gnd.n7206 gnd.n298 240.244
R5100 gnd.n7270 gnd.n298 240.244
R5101 gnd.n7270 gnd.n295 240.244
R5102 gnd.n7266 gnd.n295 240.244
R5103 gnd.n7266 gnd.n264 240.244
R5104 gnd.n7261 gnd.n264 240.244
R5105 gnd.n7261 gnd.n257 240.244
R5106 gnd.n7257 gnd.n257 240.244
R5107 gnd.n7257 gnd.n249 240.244
R5108 gnd.n7254 gnd.n249 240.244
R5109 gnd.n7254 gnd.n239 240.244
R5110 gnd.n7251 gnd.n239 240.244
R5111 gnd.n7251 gnd.n232 240.244
R5112 gnd.n7248 gnd.n232 240.244
R5113 gnd.n7248 gnd.n226 240.244
R5114 gnd.n7245 gnd.n226 240.244
R5115 gnd.n7245 gnd.n219 240.244
R5116 gnd.n7242 gnd.n219 240.244
R5117 gnd.n7242 gnd.n209 240.244
R5118 gnd.n7239 gnd.n209 240.244
R5119 gnd.n7239 gnd.n202 240.244
R5120 gnd.n7236 gnd.n202 240.244
R5121 gnd.n7236 gnd.n194 240.244
R5122 gnd.n194 gnd.n183 240.244
R5123 gnd.n7455 gnd.n183 240.244
R5124 gnd.n7456 gnd.n7455 240.244
R5125 gnd.n7456 gnd.n105 240.244
R5126 gnd.n1448 gnd.n1447 240.244
R5127 gnd.n4491 gnd.n1447 240.244
R5128 gnd.n4489 gnd.n4488 240.244
R5129 gnd.n4485 gnd.n4484 240.244
R5130 gnd.n4481 gnd.n4480 240.244
R5131 gnd.n4477 gnd.n4476 240.244
R5132 gnd.n4473 gnd.n4472 240.244
R5133 gnd.n4469 gnd.n4468 240.244
R5134 gnd.n4464 gnd.n4463 240.244
R5135 gnd.n4460 gnd.n4459 240.244
R5136 gnd.n4456 gnd.n4455 240.244
R5137 gnd.n4452 gnd.n4451 240.244
R5138 gnd.n4448 gnd.n4447 240.244
R5139 gnd.n4444 gnd.n4443 240.244
R5140 gnd.n4440 gnd.n4439 240.244
R5141 gnd.n4436 gnd.n4435 240.244
R5142 gnd.n4432 gnd.n4431 240.244
R5143 gnd.n1490 gnd.n1489 240.244
R5144 gnd.n1646 gnd.n1449 240.244
R5145 gnd.n1646 gnd.n1624 240.244
R5146 gnd.n4249 gnd.n1624 240.244
R5147 gnd.n4249 gnd.n1619 240.244
R5148 gnd.n4257 gnd.n1619 240.244
R5149 gnd.n4257 gnd.n1620 240.244
R5150 gnd.n1620 gnd.n1596 240.244
R5151 gnd.n4280 gnd.n1596 240.244
R5152 gnd.n4280 gnd.n1591 240.244
R5153 gnd.n4288 gnd.n1591 240.244
R5154 gnd.n4288 gnd.n1592 240.244
R5155 gnd.n1592 gnd.n1569 240.244
R5156 gnd.n4317 gnd.n1569 240.244
R5157 gnd.n4317 gnd.n1564 240.244
R5158 gnd.n4325 gnd.n1564 240.244
R5159 gnd.n4325 gnd.n1565 240.244
R5160 gnd.n1565 gnd.n1534 240.244
R5161 gnd.n4380 gnd.n1534 240.244
R5162 gnd.n4380 gnd.n1530 240.244
R5163 gnd.n4386 gnd.n1530 240.244
R5164 gnd.n4386 gnd.n276 240.244
R5165 gnd.n7293 gnd.n276 240.244
R5166 gnd.n7293 gnd.n277 240.244
R5167 gnd.n305 gnd.n277 240.244
R5168 gnd.n7201 gnd.n305 240.244
R5169 gnd.n7204 gnd.n7201 240.244
R5170 gnd.n7204 gnd.n297 240.244
R5171 gnd.n7272 gnd.n297 240.244
R5172 gnd.n7275 gnd.n7272 240.244
R5173 gnd.n7275 gnd.n266 240.244
R5174 gnd.n7298 gnd.n266 240.244
R5175 gnd.n7298 gnd.n255 240.244
R5176 gnd.n7308 gnd.n255 240.244
R5177 gnd.n7308 gnd.n251 240.244
R5178 gnd.n7314 gnd.n251 240.244
R5179 gnd.n7314 gnd.n237 240.244
R5180 gnd.n7324 gnd.n237 240.244
R5181 gnd.n7324 gnd.n233 240.244
R5182 gnd.n7330 gnd.n233 240.244
R5183 gnd.n7330 gnd.n224 240.244
R5184 gnd.n7340 gnd.n224 240.244
R5185 gnd.n7340 gnd.n220 240.244
R5186 gnd.n7346 gnd.n220 240.244
R5187 gnd.n7346 gnd.n207 240.244
R5188 gnd.n7356 gnd.n207 240.244
R5189 gnd.n7356 gnd.n203 240.244
R5190 gnd.n7362 gnd.n203 240.244
R5191 gnd.n7362 gnd.n192 240.244
R5192 gnd.n7447 gnd.n192 240.244
R5193 gnd.n7447 gnd.n188 240.244
R5194 gnd.n7453 gnd.n188 240.244
R5195 gnd.n7453 gnd.n108 240.244
R5196 gnd.n7533 gnd.n108 240.244
R5197 gnd.n2284 gnd.n1269 240.244
R5198 gnd.n3141 gnd.n2285 240.244
R5199 gnd.n3137 gnd.n3136 240.244
R5200 gnd.n3133 gnd.n3132 240.244
R5201 gnd.n3129 gnd.n3128 240.244
R5202 gnd.n3125 gnd.n3124 240.244
R5203 gnd.n3121 gnd.n3120 240.244
R5204 gnd.n3117 gnd.n3116 240.244
R5205 gnd.n2875 gnd.n2874 240.244
R5206 gnd.n2872 gnd.n2871 240.244
R5207 gnd.n2868 gnd.n2867 240.244
R5208 gnd.n2864 gnd.n2863 240.244
R5209 gnd.n2860 gnd.n2859 240.244
R5210 gnd.n2856 gnd.n2855 240.244
R5211 gnd.n2852 gnd.n2851 240.244
R5212 gnd.n2848 gnd.n2847 240.244
R5213 gnd.n2844 gnd.n2843 240.244
R5214 gnd.n2840 gnd.n2839 240.244
R5215 gnd.n4826 gnd.n1009 240.244
R5216 gnd.n1013 gnd.n1009 240.244
R5217 gnd.n4819 gnd.n1013 240.244
R5218 gnd.n4819 gnd.n1014 240.244
R5219 gnd.n1027 gnd.n1014 240.244
R5220 gnd.n2431 gnd.n1027 240.244
R5221 gnd.n2431 gnd.n1038 240.244
R5222 gnd.n2436 gnd.n1038 240.244
R5223 gnd.n2436 gnd.n1048 240.244
R5224 gnd.n2439 gnd.n1048 240.244
R5225 gnd.n2439 gnd.n1058 240.244
R5226 gnd.n2444 gnd.n1058 240.244
R5227 gnd.n2444 gnd.n1068 240.244
R5228 gnd.n2447 gnd.n1068 240.244
R5229 gnd.n2447 gnd.n1078 240.244
R5230 gnd.n2452 gnd.n1078 240.244
R5231 gnd.n2452 gnd.n1088 240.244
R5232 gnd.n2455 gnd.n1088 240.244
R5233 gnd.n2455 gnd.n1099 240.244
R5234 gnd.n2593 gnd.n1099 240.244
R5235 gnd.n2593 gnd.n1110 240.244
R5236 gnd.n2414 gnd.n1110 240.244
R5237 gnd.n2414 gnd.n1120 240.244
R5238 gnd.n2641 gnd.n1120 240.244
R5239 gnd.n2641 gnd.n1129 240.244
R5240 gnd.n2637 gnd.n1129 240.244
R5241 gnd.n2637 gnd.n1139 240.244
R5242 gnd.n2626 gnd.n1139 240.244
R5243 gnd.n2626 gnd.n1147 240.244
R5244 gnd.n2378 gnd.n1147 240.244
R5245 gnd.n2378 gnd.n1157 240.244
R5246 gnd.n2668 gnd.n1157 240.244
R5247 gnd.n2668 gnd.n1167 240.244
R5248 gnd.n2675 gnd.n1167 240.244
R5249 gnd.n2675 gnd.n1177 240.244
R5250 gnd.n2685 gnd.n1177 240.244
R5251 gnd.n2685 gnd.n1188 240.244
R5252 gnd.n2354 gnd.n1188 240.244
R5253 gnd.n2354 gnd.n1198 240.244
R5254 gnd.n2693 gnd.n1198 240.244
R5255 gnd.n2693 gnd.n1209 240.244
R5256 gnd.n2698 gnd.n1209 240.244
R5257 gnd.n2698 gnd.n1219 240.244
R5258 gnd.n2708 gnd.n1219 240.244
R5259 gnd.n2708 gnd.n1230 240.244
R5260 gnd.n2342 gnd.n1230 240.244
R5261 gnd.n2342 gnd.n1240 240.244
R5262 gnd.n2785 gnd.n1240 240.244
R5263 gnd.n2785 gnd.n1251 240.244
R5264 gnd.n2792 gnd.n1251 240.244
R5265 gnd.n2792 gnd.n1262 240.244
R5266 gnd.n2832 gnd.n1262 240.244
R5267 gnd.n2832 gnd.n1271 240.244
R5268 gnd.n963 gnd.n962 240.244
R5269 gnd.n4898 gnd.n962 240.244
R5270 gnd.n4896 gnd.n4895 240.244
R5271 gnd.n4892 gnd.n4891 240.244
R5272 gnd.n4888 gnd.n4887 240.244
R5273 gnd.n4884 gnd.n4883 240.244
R5274 gnd.n4880 gnd.n4879 240.244
R5275 gnd.n4876 gnd.n4875 240.244
R5276 gnd.n4872 gnd.n4871 240.244
R5277 gnd.n4867 gnd.n4866 240.244
R5278 gnd.n4863 gnd.n4862 240.244
R5279 gnd.n4859 gnd.n4858 240.244
R5280 gnd.n4855 gnd.n4854 240.244
R5281 gnd.n4851 gnd.n4850 240.244
R5282 gnd.n4847 gnd.n4846 240.244
R5283 gnd.n4843 gnd.n4842 240.244
R5284 gnd.n4839 gnd.n4838 240.244
R5285 gnd.n4835 gnd.n4834 240.244
R5286 gnd.n1004 gnd.n1003 240.244
R5287 gnd.n2549 gnd.n964 240.244
R5288 gnd.n2549 gnd.n1019 240.244
R5289 gnd.n4817 gnd.n1019 240.244
R5290 gnd.n4817 gnd.n1020 240.244
R5291 gnd.n4813 gnd.n1020 240.244
R5292 gnd.n4813 gnd.n1026 240.244
R5293 gnd.n4805 gnd.n1026 240.244
R5294 gnd.n4805 gnd.n1041 240.244
R5295 gnd.n4801 gnd.n1041 240.244
R5296 gnd.n4801 gnd.n1047 240.244
R5297 gnd.n4793 gnd.n1047 240.244
R5298 gnd.n4793 gnd.n1060 240.244
R5299 gnd.n4789 gnd.n1060 240.244
R5300 gnd.n4789 gnd.n1066 240.244
R5301 gnd.n4781 gnd.n1066 240.244
R5302 gnd.n4781 gnd.n1081 240.244
R5303 gnd.n4777 gnd.n1081 240.244
R5304 gnd.n4777 gnd.n1087 240.244
R5305 gnd.n4769 gnd.n1087 240.244
R5306 gnd.n4769 gnd.n1102 240.244
R5307 gnd.n4765 gnd.n1102 240.244
R5308 gnd.n4765 gnd.n1108 240.244
R5309 gnd.n4757 gnd.n1108 240.244
R5310 gnd.n4757 gnd.n1123 240.244
R5311 gnd.n4753 gnd.n1123 240.244
R5312 gnd.n4753 gnd.n1127 240.244
R5313 gnd.n4745 gnd.n1127 240.244
R5314 gnd.n4745 gnd.n1142 240.244
R5315 gnd.n4740 gnd.n1142 240.244
R5316 gnd.n4740 gnd.n1145 240.244
R5317 gnd.n4732 gnd.n1145 240.244
R5318 gnd.n4732 gnd.n1160 240.244
R5319 gnd.n4728 gnd.n1160 240.244
R5320 gnd.n4728 gnd.n1165 240.244
R5321 gnd.n4720 gnd.n1165 240.244
R5322 gnd.n4720 gnd.n1180 240.244
R5323 gnd.n4716 gnd.n1180 240.244
R5324 gnd.n4716 gnd.n1186 240.244
R5325 gnd.n4708 gnd.n1186 240.244
R5326 gnd.n4708 gnd.n1201 240.244
R5327 gnd.n4704 gnd.n1201 240.244
R5328 gnd.n4704 gnd.n1207 240.244
R5329 gnd.n4696 gnd.n1207 240.244
R5330 gnd.n4696 gnd.n1222 240.244
R5331 gnd.n4692 gnd.n1222 240.244
R5332 gnd.n4692 gnd.n1228 240.244
R5333 gnd.n4684 gnd.n1228 240.244
R5334 gnd.n4684 gnd.n1243 240.244
R5335 gnd.n4680 gnd.n1243 240.244
R5336 gnd.n4680 gnd.n1249 240.244
R5337 gnd.n4672 gnd.n1249 240.244
R5338 gnd.n4672 gnd.n1264 240.244
R5339 gnd.n4668 gnd.n1264 240.244
R5340 gnd.n4913 gnd.n4908 240.244
R5341 gnd.n6301 gnd.n6300 240.244
R5342 gnd.n6298 gnd.n4917 240.244
R5343 gnd.n6294 gnd.n6293 240.244
R5344 gnd.n6291 gnd.n4924 240.244
R5345 gnd.n6287 gnd.n6286 240.244
R5346 gnd.n6284 gnd.n4931 240.244
R5347 gnd.n6280 gnd.n6279 240.244
R5348 gnd.n5594 gnd.n5220 240.244
R5349 gnd.n5604 gnd.n5220 240.244
R5350 gnd.n5604 gnd.n5211 240.244
R5351 gnd.n5211 gnd.n5200 240.244
R5352 gnd.n5625 gnd.n5200 240.244
R5353 gnd.n5625 gnd.n5194 240.244
R5354 gnd.n5635 gnd.n5194 240.244
R5355 gnd.n5635 gnd.n5185 240.244
R5356 gnd.n5185 gnd.n5176 240.244
R5357 gnd.n5656 gnd.n5176 240.244
R5358 gnd.n5656 gnd.n5169 240.244
R5359 gnd.n5666 gnd.n5169 240.244
R5360 gnd.n5666 gnd.n5160 240.244
R5361 gnd.n5160 gnd.n5150 240.244
R5362 gnd.n5687 gnd.n5150 240.244
R5363 gnd.n5687 gnd.n5143 240.244
R5364 gnd.n5697 gnd.n5143 240.244
R5365 gnd.n5697 gnd.n5134 240.244
R5366 gnd.n5134 gnd.n5125 240.244
R5367 gnd.n5718 gnd.n5125 240.244
R5368 gnd.n5718 gnd.n5118 240.244
R5369 gnd.n5728 gnd.n5118 240.244
R5370 gnd.n5728 gnd.n5110 240.244
R5371 gnd.n5110 gnd.n5101 240.244
R5372 gnd.n5748 gnd.n5101 240.244
R5373 gnd.n5748 gnd.n5088 240.244
R5374 gnd.n5782 gnd.n5088 240.244
R5375 gnd.n5782 gnd.n5078 240.244
R5376 gnd.n5078 gnd.n5070 240.244
R5377 gnd.n5800 gnd.n5070 240.244
R5378 gnd.n5801 gnd.n5800 240.244
R5379 gnd.n5801 gnd.n5058 240.244
R5380 gnd.n5058 gnd.n5047 240.244
R5381 gnd.n5832 gnd.n5047 240.244
R5382 gnd.n5833 gnd.n5832 240.244
R5383 gnd.n5836 gnd.n5833 240.244
R5384 gnd.n5836 gnd.n5033 240.244
R5385 gnd.n5864 gnd.n5033 240.244
R5386 gnd.n5864 gnd.n5020 240.244
R5387 gnd.n5886 gnd.n5020 240.244
R5388 gnd.n5887 gnd.n5886 240.244
R5389 gnd.n5887 gnd.n5004 240.244
R5390 gnd.n5897 gnd.n5004 240.244
R5391 gnd.n5897 gnd.n4996 240.244
R5392 gnd.n6179 gnd.n4996 240.244
R5393 gnd.n6179 gnd.n6178 240.244
R5394 gnd.n6178 gnd.n6177 240.244
R5395 gnd.n6177 gnd.n909 240.244
R5396 gnd.n6173 gnd.n909 240.244
R5397 gnd.n6173 gnd.n920 240.244
R5398 gnd.n6169 gnd.n920 240.244
R5399 gnd.n6169 gnd.n6168 240.244
R5400 gnd.n6168 gnd.n932 240.244
R5401 gnd.n5584 gnd.n5233 240.244
R5402 gnd.n5254 gnd.n5233 240.244
R5403 gnd.n5257 gnd.n5256 240.244
R5404 gnd.n5264 gnd.n5263 240.244
R5405 gnd.n5267 gnd.n5266 240.244
R5406 gnd.n5274 gnd.n5273 240.244
R5407 gnd.n5277 gnd.n5276 240.244
R5408 gnd.n5284 gnd.n5283 240.244
R5409 gnd.n5592 gnd.n5230 240.244
R5410 gnd.n5230 gnd.n5209 240.244
R5411 gnd.n5615 gnd.n5209 240.244
R5412 gnd.n5615 gnd.n5203 240.244
R5413 gnd.n5623 gnd.n5203 240.244
R5414 gnd.n5623 gnd.n5205 240.244
R5415 gnd.n5205 gnd.n5183 240.244
R5416 gnd.n5646 gnd.n5183 240.244
R5417 gnd.n5646 gnd.n5178 240.244
R5418 gnd.n5654 gnd.n5178 240.244
R5419 gnd.n5654 gnd.n5179 240.244
R5420 gnd.n5179 gnd.n5158 240.244
R5421 gnd.n5677 gnd.n5158 240.244
R5422 gnd.n5677 gnd.n5153 240.244
R5423 gnd.n5685 gnd.n5153 240.244
R5424 gnd.n5685 gnd.n5154 240.244
R5425 gnd.n5154 gnd.n5132 240.244
R5426 gnd.n5708 gnd.n5132 240.244
R5427 gnd.n5708 gnd.n5127 240.244
R5428 gnd.n5716 gnd.n5127 240.244
R5429 gnd.n5716 gnd.n5128 240.244
R5430 gnd.n5128 gnd.n5108 240.244
R5431 gnd.n5738 gnd.n5108 240.244
R5432 gnd.n5738 gnd.n5103 240.244
R5433 gnd.n5746 gnd.n5103 240.244
R5434 gnd.n5746 gnd.n5104 240.244
R5435 gnd.n5104 gnd.n5077 240.244
R5436 gnd.n5792 gnd.n5077 240.244
R5437 gnd.n5792 gnd.n5073 240.244
R5438 gnd.n5798 gnd.n5073 240.244
R5439 gnd.n5798 gnd.n5056 240.244
R5440 gnd.n5822 gnd.n5056 240.244
R5441 gnd.n5822 gnd.n5051 240.244
R5442 gnd.n5830 gnd.n5051 240.244
R5443 gnd.n5830 gnd.n5052 240.244
R5444 gnd.n5052 gnd.n5032 240.244
R5445 gnd.n5868 gnd.n5032 240.244
R5446 gnd.n5868 gnd.n5027 240.244
R5447 gnd.n5876 gnd.n5027 240.244
R5448 gnd.n5876 gnd.n5028 240.244
R5449 gnd.n5028 gnd.n5002 240.244
R5450 gnd.n6189 gnd.n5002 240.244
R5451 gnd.n6189 gnd.n4997 240.244
R5452 gnd.n6201 gnd.n4997 240.244
R5453 gnd.n6201 gnd.n4998 240.244
R5454 gnd.n6197 gnd.n4998 240.244
R5455 gnd.n6197 gnd.n911 240.244
R5456 gnd.n6322 gnd.n911 240.244
R5457 gnd.n6322 gnd.n912 240.244
R5458 gnd.n6318 gnd.n912 240.244
R5459 gnd.n6318 gnd.n918 240.244
R5460 gnd.n4907 gnd.n918 240.244
R5461 gnd.n6308 gnd.n4907 240.244
R5462 gnd.n4943 gnd.n929 240.244
R5463 gnd.n6269 gnd.n6268 240.244
R5464 gnd.n6266 gnd.n4947 240.244
R5465 gnd.n6262 gnd.n6261 240.244
R5466 gnd.n6259 gnd.n4954 240.244
R5467 gnd.n6255 gnd.n6254 240.244
R5468 gnd.n6252 gnd.n4961 240.244
R5469 gnd.n6248 gnd.n6247 240.244
R5470 gnd.n6245 gnd.n4968 240.244
R5471 gnd.n6241 gnd.n6240 240.244
R5472 gnd.n6238 gnd.n4975 240.244
R5473 gnd.n6234 gnd.n6233 240.244
R5474 gnd.n6231 gnd.n4985 240.244
R5475 gnd.n5421 gnd.n5318 240.244
R5476 gnd.n5421 gnd.n5311 240.244
R5477 gnd.n5432 gnd.n5311 240.244
R5478 gnd.n5432 gnd.n5307 240.244
R5479 gnd.n5438 gnd.n5307 240.244
R5480 gnd.n5438 gnd.n5299 240.244
R5481 gnd.n5448 gnd.n5299 240.244
R5482 gnd.n5448 gnd.n5294 240.244
R5483 gnd.n5570 gnd.n5294 240.244
R5484 gnd.n5570 gnd.n5295 240.244
R5485 gnd.n5295 gnd.n5242 240.244
R5486 gnd.n5565 gnd.n5242 240.244
R5487 gnd.n5565 gnd.n5564 240.244
R5488 gnd.n5564 gnd.n5221 240.244
R5489 gnd.n5560 gnd.n5221 240.244
R5490 gnd.n5560 gnd.n5212 240.244
R5491 gnd.n5557 gnd.n5212 240.244
R5492 gnd.n5557 gnd.n5556 240.244
R5493 gnd.n5556 gnd.n5195 240.244
R5494 gnd.n5552 gnd.n5195 240.244
R5495 gnd.n5552 gnd.n5186 240.244
R5496 gnd.n5549 gnd.n5186 240.244
R5497 gnd.n5549 gnd.n5548 240.244
R5498 gnd.n5548 gnd.n5171 240.244
R5499 gnd.n5543 gnd.n5171 240.244
R5500 gnd.n5543 gnd.n5161 240.244
R5501 gnd.n5540 gnd.n5161 240.244
R5502 gnd.n5540 gnd.n5539 240.244
R5503 gnd.n5539 gnd.n5145 240.244
R5504 gnd.n5472 gnd.n5145 240.244
R5505 gnd.n5472 gnd.n5135 240.244
R5506 gnd.n5483 gnd.n5135 240.244
R5507 gnd.n5483 gnd.n5481 240.244
R5508 gnd.n5481 gnd.n5120 240.244
R5509 gnd.n5476 gnd.n5120 240.244
R5510 gnd.n5476 gnd.n5111 240.244
R5511 gnd.n5111 gnd.n5094 240.244
R5512 gnd.n5758 gnd.n5094 240.244
R5513 gnd.n5758 gnd.n5090 240.244
R5514 gnd.n5779 gnd.n5090 240.244
R5515 gnd.n5779 gnd.n5079 240.244
R5516 gnd.n5775 gnd.n5079 240.244
R5517 gnd.n5775 gnd.n5069 240.244
R5518 gnd.n5772 gnd.n5069 240.244
R5519 gnd.n5772 gnd.n5059 240.244
R5520 gnd.n5769 gnd.n5059 240.244
R5521 gnd.n5769 gnd.n5038 240.244
R5522 gnd.n5845 gnd.n5038 240.244
R5523 gnd.n5845 gnd.n5034 240.244
R5524 gnd.n5863 gnd.n5034 240.244
R5525 gnd.n5863 gnd.n5025 240.244
R5526 gnd.n5859 gnd.n5025 240.244
R5527 gnd.n5859 gnd.n5019 240.244
R5528 gnd.n5856 gnd.n5019 240.244
R5529 gnd.n5856 gnd.n5005 240.244
R5530 gnd.n5005 gnd.n4995 240.244
R5531 gnd.n6204 gnd.n4995 240.244
R5532 gnd.n6204 gnd.n897 240.244
R5533 gnd.n6210 gnd.n897 240.244
R5534 gnd.n6210 gnd.n908 240.244
R5535 gnd.n6214 gnd.n908 240.244
R5536 gnd.n6214 gnd.n6213 240.244
R5537 gnd.n6213 gnd.n921 240.244
R5538 gnd.n6221 gnd.n921 240.244
R5539 gnd.n6221 gnd.n931 240.244
R5540 gnd.n5335 gnd.n5334 240.244
R5541 gnd.n5406 gnd.n5334 240.244
R5542 gnd.n5404 gnd.n5403 240.244
R5543 gnd.n5400 gnd.n5399 240.244
R5544 gnd.n5396 gnd.n5395 240.244
R5545 gnd.n5392 gnd.n5391 240.244
R5546 gnd.n5388 gnd.n5387 240.244
R5547 gnd.n5384 gnd.n5383 240.244
R5548 gnd.n5380 gnd.n5379 240.244
R5549 gnd.n5376 gnd.n5375 240.244
R5550 gnd.n5372 gnd.n5371 240.244
R5551 gnd.n5368 gnd.n5367 240.244
R5552 gnd.n5364 gnd.n5322 240.244
R5553 gnd.n5424 gnd.n5316 240.244
R5554 gnd.n5424 gnd.n5312 240.244
R5555 gnd.n5430 gnd.n5312 240.244
R5556 gnd.n5430 gnd.n5305 240.244
R5557 gnd.n5440 gnd.n5305 240.244
R5558 gnd.n5440 gnd.n5301 240.244
R5559 gnd.n5446 gnd.n5301 240.244
R5560 gnd.n5446 gnd.n5292 240.244
R5561 gnd.n5572 gnd.n5292 240.244
R5562 gnd.n5572 gnd.n5243 240.244
R5563 gnd.n5580 gnd.n5243 240.244
R5564 gnd.n5580 gnd.n5244 240.244
R5565 gnd.n5244 gnd.n5222 240.244
R5566 gnd.n5601 gnd.n5222 240.244
R5567 gnd.n5601 gnd.n5214 240.244
R5568 gnd.n5612 gnd.n5214 240.244
R5569 gnd.n5612 gnd.n5215 240.244
R5570 gnd.n5215 gnd.n5196 240.244
R5571 gnd.n5632 gnd.n5196 240.244
R5572 gnd.n5632 gnd.n5188 240.244
R5573 gnd.n5643 gnd.n5188 240.244
R5574 gnd.n5643 gnd.n5189 240.244
R5575 gnd.n5189 gnd.n5172 240.244
R5576 gnd.n5663 gnd.n5172 240.244
R5577 gnd.n5663 gnd.n5163 240.244
R5578 gnd.n5674 gnd.n5163 240.244
R5579 gnd.n5674 gnd.n5164 240.244
R5580 gnd.n5164 gnd.n5146 240.244
R5581 gnd.n5694 gnd.n5146 240.244
R5582 gnd.n5694 gnd.n5137 240.244
R5583 gnd.n5705 gnd.n5137 240.244
R5584 gnd.n5705 gnd.n5138 240.244
R5585 gnd.n5138 gnd.n5121 240.244
R5586 gnd.n5725 gnd.n5121 240.244
R5587 gnd.n5725 gnd.n5113 240.244
R5588 gnd.n5735 gnd.n5113 240.244
R5589 gnd.n5735 gnd.n5096 240.244
R5590 gnd.n5756 gnd.n5096 240.244
R5591 gnd.n5756 gnd.n5097 240.244
R5592 gnd.n5097 gnd.n5081 240.244
R5593 gnd.n5789 gnd.n5081 240.244
R5594 gnd.n5789 gnd.n5068 240.244
R5595 gnd.n5804 gnd.n5068 240.244
R5596 gnd.n5804 gnd.n5061 240.244
R5597 gnd.n5819 gnd.n5061 240.244
R5598 gnd.n5819 gnd.n5062 240.244
R5599 gnd.n5062 gnd.n5040 240.244
R5600 gnd.n5843 gnd.n5040 240.244
R5601 gnd.n5843 gnd.n5041 240.244
R5602 gnd.n5041 gnd.n5024 240.244
R5603 gnd.n5879 gnd.n5024 240.244
R5604 gnd.n5879 gnd.n5017 240.244
R5605 gnd.n5890 gnd.n5017 240.244
R5606 gnd.n5890 gnd.n5007 240.244
R5607 gnd.n6186 gnd.n5007 240.244
R5608 gnd.n6186 gnd.n5009 240.244
R5609 gnd.n5009 gnd.n899 240.244
R5610 gnd.n6329 gnd.n899 240.244
R5611 gnd.n6329 gnd.n900 240.244
R5612 gnd.n6325 gnd.n900 240.244
R5613 gnd.n6325 gnd.n906 240.244
R5614 gnd.n923 gnd.n906 240.244
R5615 gnd.n6315 gnd.n923 240.244
R5616 gnd.n6315 gnd.n924 240.244
R5617 gnd.n6311 gnd.n924 240.244
R5618 gnd.n7372 gnd.n7371 240.244
R5619 gnd.n7377 gnd.n7374 240.244
R5620 gnd.n7380 gnd.n7379 240.244
R5621 gnd.n7385 gnd.n7382 240.244
R5622 gnd.n7388 gnd.n7387 240.244
R5623 gnd.n7393 gnd.n7390 240.244
R5624 gnd.n7396 gnd.n7395 240.244
R5625 gnd.n7401 gnd.n7398 240.244
R5626 gnd.n7407 gnd.n7403 240.244
R5627 gnd.n1680 gnd.n1498 240.244
R5628 gnd.n4235 gnd.n1680 240.244
R5629 gnd.n4235 gnd.n1627 240.244
R5630 gnd.n1627 gnd.n1614 240.244
R5631 gnd.n4259 gnd.n1614 240.244
R5632 gnd.n4259 gnd.n1609 240.244
R5633 gnd.n4266 gnd.n1609 240.244
R5634 gnd.n4266 gnd.n1599 240.244
R5635 gnd.n1599 gnd.n1587 240.244
R5636 gnd.n4290 gnd.n1587 240.244
R5637 gnd.n4290 gnd.n1582 240.244
R5638 gnd.n4302 gnd.n1582 240.244
R5639 gnd.n4302 gnd.n1572 240.244
R5640 gnd.n4295 gnd.n1572 240.244
R5641 gnd.n4295 gnd.n1562 240.244
R5642 gnd.n1562 gnd.n1548 240.244
R5643 gnd.n4359 gnd.n1548 240.244
R5644 gnd.n4359 gnd.n1537 240.244
R5645 gnd.n1553 gnd.n1537 240.244
R5646 gnd.n1553 gnd.n1528 240.244
R5647 gnd.n4350 gnd.n1528 240.244
R5648 gnd.n4350 gnd.n280 240.244
R5649 gnd.n7193 gnd.n280 240.244
R5650 gnd.n7193 gnd.n308 240.244
R5651 gnd.n7199 gnd.n308 240.244
R5652 gnd.n7199 gnd.n303 240.244
R5653 gnd.n303 gnd.n70 240.244
R5654 gnd.n71 gnd.n70 240.244
R5655 gnd.n72 gnd.n71 240.244
R5656 gnd.n7264 gnd.n72 240.244
R5657 gnd.n7264 gnd.n75 240.244
R5658 gnd.n76 gnd.n75 240.244
R5659 gnd.n77 gnd.n76 240.244
R5660 gnd.n247 gnd.n77 240.244
R5661 gnd.n247 gnd.n80 240.244
R5662 gnd.n81 gnd.n80 240.244
R5663 gnd.n82 gnd.n81 240.244
R5664 gnd.n240 gnd.n82 240.244
R5665 gnd.n240 gnd.n85 240.244
R5666 gnd.n86 gnd.n85 240.244
R5667 gnd.n87 gnd.n86 240.244
R5668 gnd.n217 gnd.n87 240.244
R5669 gnd.n217 gnd.n90 240.244
R5670 gnd.n91 gnd.n90 240.244
R5671 gnd.n92 gnd.n91 240.244
R5672 gnd.n210 gnd.n92 240.244
R5673 gnd.n210 gnd.n95 240.244
R5674 gnd.n96 gnd.n95 240.244
R5675 gnd.n97 gnd.n96 240.244
R5676 gnd.n184 gnd.n97 240.244
R5677 gnd.n184 gnd.n100 240.244
R5678 gnd.n101 gnd.n100 240.244
R5679 gnd.n7535 gnd.n101 240.244
R5680 gnd.n1728 gnd.n1727 240.244
R5681 gnd.n1731 gnd.n1730 240.244
R5682 gnd.n1747 gnd.n1746 240.244
R5683 gnd.n1750 gnd.n1749 240.244
R5684 gnd.n1766 gnd.n1765 240.244
R5685 gnd.n1769 gnd.n1768 240.244
R5686 gnd.n1784 gnd.n1783 240.244
R5687 gnd.n1695 gnd.n1694 240.244
R5688 gnd.n1690 gnd.n1445 240.244
R5689 gnd.n4421 gnd.n1501 240.244
R5690 gnd.n1505 gnd.n1501 240.244
R5691 gnd.n1506 gnd.n1505 240.244
R5692 gnd.n1507 gnd.n1506 240.244
R5693 gnd.n1618 gnd.n1507 240.244
R5694 gnd.n1618 gnd.n1510 240.244
R5695 gnd.n1511 gnd.n1510 240.244
R5696 gnd.n1512 gnd.n1511 240.244
R5697 gnd.n1600 gnd.n1512 240.244
R5698 gnd.n1600 gnd.n1515 240.244
R5699 gnd.n1516 gnd.n1515 240.244
R5700 gnd.n1517 gnd.n1516 240.244
R5701 gnd.n4315 gnd.n1517 240.244
R5702 gnd.n4315 gnd.n1520 240.244
R5703 gnd.n1521 gnd.n1520 240.244
R5704 gnd.n1522 gnd.n1521 240.244
R5705 gnd.n4360 gnd.n1522 240.244
R5706 gnd.n4360 gnd.n1525 240.244
R5707 gnd.n1526 gnd.n1525 240.244
R5708 gnd.n4388 gnd.n1526 240.244
R5709 gnd.n4388 gnd.n281 240.244
R5710 gnd.n7291 gnd.n281 240.244
R5711 gnd.n7291 gnd.n282 240.244
R5712 gnd.n287 gnd.n282 240.244
R5713 gnd.n288 gnd.n287 240.244
R5714 gnd.n289 gnd.n288 240.244
R5715 gnd.n319 gnd.n289 240.244
R5716 gnd.n319 gnd.n293 240.244
R5717 gnd.n7277 gnd.n293 240.244
R5718 gnd.n7277 gnd.n262 240.244
R5719 gnd.n7300 gnd.n262 240.244
R5720 gnd.n7300 gnd.n258 240.244
R5721 gnd.n7306 gnd.n258 240.244
R5722 gnd.n7306 gnd.n246 240.244
R5723 gnd.n7316 gnd.n246 240.244
R5724 gnd.n7316 gnd.n242 240.244
R5725 gnd.n7322 gnd.n242 240.244
R5726 gnd.n7322 gnd.n231 240.244
R5727 gnd.n7332 gnd.n231 240.244
R5728 gnd.n7332 gnd.n227 240.244
R5729 gnd.n7338 gnd.n227 240.244
R5730 gnd.n7338 gnd.n216 240.244
R5731 gnd.n7348 gnd.n216 240.244
R5732 gnd.n7348 gnd.n212 240.244
R5733 gnd.n7354 gnd.n212 240.244
R5734 gnd.n7354 gnd.n201 240.244
R5735 gnd.n7364 gnd.n201 240.244
R5736 gnd.n7364 gnd.n195 240.244
R5737 gnd.n7445 gnd.n195 240.244
R5738 gnd.n7445 gnd.n196 240.244
R5739 gnd.n196 gnd.n187 240.244
R5740 gnd.n7369 gnd.n187 240.244
R5741 gnd.n7369 gnd.n107 240.244
R5742 gnd.n2251 gnd.n1274 240.244
R5743 gnd.n2252 gnd.n2201 240.244
R5744 gnd.n2255 gnd.n2202 240.244
R5745 gnd.n2211 gnd.n2210 240.244
R5746 gnd.n2257 gnd.n2218 240.244
R5747 gnd.n2260 gnd.n2219 240.244
R5748 gnd.n2229 gnd.n2228 240.244
R5749 gnd.n2262 gnd.n2236 240.244
R5750 gnd.n2248 gnd.n2237 240.244
R5751 gnd.n2551 gnd.n2471 240.244
R5752 gnd.n2552 gnd.n2551 240.244
R5753 gnd.n2552 gnd.n1016 240.244
R5754 gnd.n2557 gnd.n1016 240.244
R5755 gnd.n2557 gnd.n1028 240.244
R5756 gnd.n2560 gnd.n1028 240.244
R5757 gnd.n2560 gnd.n1039 240.244
R5758 gnd.n2565 gnd.n1039 240.244
R5759 gnd.n2565 gnd.n1049 240.244
R5760 gnd.n2568 gnd.n1049 240.244
R5761 gnd.n2568 gnd.n1059 240.244
R5762 gnd.n2573 gnd.n1059 240.244
R5763 gnd.n2573 gnd.n1069 240.244
R5764 gnd.n2576 gnd.n1069 240.244
R5765 gnd.n2576 gnd.n1079 240.244
R5766 gnd.n2581 gnd.n1079 240.244
R5767 gnd.n2581 gnd.n1089 240.244
R5768 gnd.n2584 gnd.n1089 240.244
R5769 gnd.n2584 gnd.n1100 240.244
R5770 gnd.n2591 gnd.n1100 240.244
R5771 gnd.n2591 gnd.n1111 240.244
R5772 gnd.n2647 gnd.n1111 240.244
R5773 gnd.n2647 gnd.n1121 240.244
R5774 gnd.n2643 gnd.n1121 240.244
R5775 gnd.n2643 gnd.n1130 240.244
R5776 gnd.n2635 gnd.n1130 240.244
R5777 gnd.n2635 gnd.n1140 240.244
R5778 gnd.n2628 gnd.n1140 240.244
R5779 gnd.n2628 gnd.n1148 240.244
R5780 gnd.n2660 gnd.n1148 240.244
R5781 gnd.n2660 gnd.n1158 240.244
R5782 gnd.n2666 gnd.n1158 240.244
R5783 gnd.n2666 gnd.n1168 240.244
R5784 gnd.n2677 gnd.n1168 240.244
R5785 gnd.n2677 gnd.n1178 240.244
R5786 gnd.n2683 gnd.n1178 240.244
R5787 gnd.n2683 gnd.n1189 240.244
R5788 gnd.n2722 gnd.n1189 240.244
R5789 gnd.n2722 gnd.n1199 240.244
R5790 gnd.n2359 gnd.n1199 240.244
R5791 gnd.n2359 gnd.n1210 240.244
R5792 gnd.n2360 gnd.n1210 240.244
R5793 gnd.n2360 gnd.n1220 240.244
R5794 gnd.n2710 gnd.n1220 240.244
R5795 gnd.n2710 gnd.n1231 240.244
R5796 gnd.n2777 gnd.n1231 240.244
R5797 gnd.n2777 gnd.n1241 240.244
R5798 gnd.n2783 gnd.n1241 240.244
R5799 gnd.n2783 gnd.n1252 240.244
R5800 gnd.n2794 gnd.n1252 240.244
R5801 gnd.n2794 gnd.n1263 240.244
R5802 gnd.n2830 gnd.n1263 240.244
R5803 gnd.n2830 gnd.n1272 240.244
R5804 gnd.n2531 gnd.n2530 240.244
R5805 gnd.n2527 gnd.n2526 240.244
R5806 gnd.n2523 gnd.n2522 240.244
R5807 gnd.n2519 gnd.n2518 240.244
R5808 gnd.n2515 gnd.n2514 240.244
R5809 gnd.n2511 gnd.n2510 240.244
R5810 gnd.n2507 gnd.n2506 240.244
R5811 gnd.n2503 gnd.n2502 240.244
R5812 gnd.n2491 gnd.n960 240.244
R5813 gnd.n2543 gnd.n2472 240.244
R5814 gnd.n2543 gnd.n2473 240.244
R5815 gnd.n2473 gnd.n1018 240.244
R5816 gnd.n1030 gnd.n1018 240.244
R5817 gnd.n4811 gnd.n1030 240.244
R5818 gnd.n4811 gnd.n1031 240.244
R5819 gnd.n4807 gnd.n1031 240.244
R5820 gnd.n4807 gnd.n1037 240.244
R5821 gnd.n4799 gnd.n1037 240.244
R5822 gnd.n4799 gnd.n1050 240.244
R5823 gnd.n4795 gnd.n1050 240.244
R5824 gnd.n4795 gnd.n1056 240.244
R5825 gnd.n4787 gnd.n1056 240.244
R5826 gnd.n4787 gnd.n1071 240.244
R5827 gnd.n4783 gnd.n1071 240.244
R5828 gnd.n4783 gnd.n1077 240.244
R5829 gnd.n4775 gnd.n1077 240.244
R5830 gnd.n4775 gnd.n1090 240.244
R5831 gnd.n4771 gnd.n1090 240.244
R5832 gnd.n4771 gnd.n1096 240.244
R5833 gnd.n4763 gnd.n1096 240.244
R5834 gnd.n4763 gnd.n1113 240.244
R5835 gnd.n4759 gnd.n1113 240.244
R5836 gnd.n4759 gnd.n1119 240.244
R5837 gnd.n4751 gnd.n1119 240.244
R5838 gnd.n4751 gnd.n1131 240.244
R5839 gnd.n4747 gnd.n1131 240.244
R5840 gnd.n4747 gnd.n1137 240.244
R5841 gnd.n4738 gnd.n1137 240.244
R5842 gnd.n4738 gnd.n1150 240.244
R5843 gnd.n4734 gnd.n1150 240.244
R5844 gnd.n4734 gnd.n1156 240.244
R5845 gnd.n4726 gnd.n1156 240.244
R5846 gnd.n4726 gnd.n1169 240.244
R5847 gnd.n4722 gnd.n1169 240.244
R5848 gnd.n4722 gnd.n1175 240.244
R5849 gnd.n4714 gnd.n1175 240.244
R5850 gnd.n4714 gnd.n1191 240.244
R5851 gnd.n4710 gnd.n1191 240.244
R5852 gnd.n4710 gnd.n1197 240.244
R5853 gnd.n4702 gnd.n1197 240.244
R5854 gnd.n4702 gnd.n1211 240.244
R5855 gnd.n4698 gnd.n1211 240.244
R5856 gnd.n4698 gnd.n1217 240.244
R5857 gnd.n4690 gnd.n1217 240.244
R5858 gnd.n4690 gnd.n1233 240.244
R5859 gnd.n4686 gnd.n1233 240.244
R5860 gnd.n4686 gnd.n1239 240.244
R5861 gnd.n4678 gnd.n1239 240.244
R5862 gnd.n4678 gnd.n1254 240.244
R5863 gnd.n4674 gnd.n1254 240.244
R5864 gnd.n4674 gnd.n1260 240.244
R5865 gnd.n4666 gnd.n1260 240.244
R5866 gnd.n6501 gnd.n724 240.244
R5867 gnd.n6507 gnd.n724 240.244
R5868 gnd.n6507 gnd.n722 240.244
R5869 gnd.n6511 gnd.n722 240.244
R5870 gnd.n6511 gnd.n718 240.244
R5871 gnd.n6517 gnd.n718 240.244
R5872 gnd.n6517 gnd.n716 240.244
R5873 gnd.n6521 gnd.n716 240.244
R5874 gnd.n6521 gnd.n712 240.244
R5875 gnd.n6527 gnd.n712 240.244
R5876 gnd.n6527 gnd.n710 240.244
R5877 gnd.n6531 gnd.n710 240.244
R5878 gnd.n6531 gnd.n706 240.244
R5879 gnd.n6537 gnd.n706 240.244
R5880 gnd.n6537 gnd.n704 240.244
R5881 gnd.n6541 gnd.n704 240.244
R5882 gnd.n6541 gnd.n700 240.244
R5883 gnd.n6547 gnd.n700 240.244
R5884 gnd.n6547 gnd.n698 240.244
R5885 gnd.n6551 gnd.n698 240.244
R5886 gnd.n6551 gnd.n694 240.244
R5887 gnd.n6557 gnd.n694 240.244
R5888 gnd.n6557 gnd.n692 240.244
R5889 gnd.n6561 gnd.n692 240.244
R5890 gnd.n6561 gnd.n688 240.244
R5891 gnd.n6567 gnd.n688 240.244
R5892 gnd.n6567 gnd.n686 240.244
R5893 gnd.n6571 gnd.n686 240.244
R5894 gnd.n6571 gnd.n682 240.244
R5895 gnd.n6577 gnd.n682 240.244
R5896 gnd.n6577 gnd.n680 240.244
R5897 gnd.n6581 gnd.n680 240.244
R5898 gnd.n6581 gnd.n676 240.244
R5899 gnd.n6587 gnd.n676 240.244
R5900 gnd.n6587 gnd.n674 240.244
R5901 gnd.n6591 gnd.n674 240.244
R5902 gnd.n6591 gnd.n670 240.244
R5903 gnd.n6597 gnd.n670 240.244
R5904 gnd.n6597 gnd.n668 240.244
R5905 gnd.n6601 gnd.n668 240.244
R5906 gnd.n6601 gnd.n664 240.244
R5907 gnd.n6607 gnd.n664 240.244
R5908 gnd.n6607 gnd.n662 240.244
R5909 gnd.n6611 gnd.n662 240.244
R5910 gnd.n6611 gnd.n658 240.244
R5911 gnd.n6617 gnd.n658 240.244
R5912 gnd.n6617 gnd.n656 240.244
R5913 gnd.n6621 gnd.n656 240.244
R5914 gnd.n6621 gnd.n652 240.244
R5915 gnd.n6627 gnd.n652 240.244
R5916 gnd.n6627 gnd.n650 240.244
R5917 gnd.n6631 gnd.n650 240.244
R5918 gnd.n6631 gnd.n646 240.244
R5919 gnd.n6637 gnd.n646 240.244
R5920 gnd.n6637 gnd.n644 240.244
R5921 gnd.n6641 gnd.n644 240.244
R5922 gnd.n6641 gnd.n640 240.244
R5923 gnd.n6647 gnd.n640 240.244
R5924 gnd.n6647 gnd.n638 240.244
R5925 gnd.n6651 gnd.n638 240.244
R5926 gnd.n6651 gnd.n634 240.244
R5927 gnd.n6657 gnd.n634 240.244
R5928 gnd.n6657 gnd.n632 240.244
R5929 gnd.n6661 gnd.n632 240.244
R5930 gnd.n6661 gnd.n628 240.244
R5931 gnd.n6667 gnd.n628 240.244
R5932 gnd.n6667 gnd.n626 240.244
R5933 gnd.n6671 gnd.n626 240.244
R5934 gnd.n6671 gnd.n622 240.244
R5935 gnd.n6677 gnd.n622 240.244
R5936 gnd.n6677 gnd.n620 240.244
R5937 gnd.n6681 gnd.n620 240.244
R5938 gnd.n6681 gnd.n616 240.244
R5939 gnd.n6687 gnd.n616 240.244
R5940 gnd.n6687 gnd.n614 240.244
R5941 gnd.n6691 gnd.n614 240.244
R5942 gnd.n6691 gnd.n610 240.244
R5943 gnd.n6697 gnd.n610 240.244
R5944 gnd.n6697 gnd.n608 240.244
R5945 gnd.n6701 gnd.n608 240.244
R5946 gnd.n6701 gnd.n604 240.244
R5947 gnd.n6707 gnd.n604 240.244
R5948 gnd.n6707 gnd.n602 240.244
R5949 gnd.n6711 gnd.n602 240.244
R5950 gnd.n6711 gnd.n598 240.244
R5951 gnd.n6717 gnd.n598 240.244
R5952 gnd.n6717 gnd.n596 240.244
R5953 gnd.n6721 gnd.n596 240.244
R5954 gnd.n6721 gnd.n592 240.244
R5955 gnd.n6727 gnd.n592 240.244
R5956 gnd.n6727 gnd.n590 240.244
R5957 gnd.n6731 gnd.n590 240.244
R5958 gnd.n6731 gnd.n586 240.244
R5959 gnd.n6737 gnd.n586 240.244
R5960 gnd.n6737 gnd.n584 240.244
R5961 gnd.n6741 gnd.n584 240.244
R5962 gnd.n6741 gnd.n580 240.244
R5963 gnd.n6747 gnd.n580 240.244
R5964 gnd.n6747 gnd.n578 240.244
R5965 gnd.n6751 gnd.n578 240.244
R5966 gnd.n6751 gnd.n574 240.244
R5967 gnd.n6757 gnd.n574 240.244
R5968 gnd.n6757 gnd.n572 240.244
R5969 gnd.n6761 gnd.n572 240.244
R5970 gnd.n6761 gnd.n568 240.244
R5971 gnd.n6767 gnd.n568 240.244
R5972 gnd.n6767 gnd.n566 240.244
R5973 gnd.n6771 gnd.n566 240.244
R5974 gnd.n6771 gnd.n562 240.244
R5975 gnd.n6777 gnd.n562 240.244
R5976 gnd.n6777 gnd.n560 240.244
R5977 gnd.n6781 gnd.n560 240.244
R5978 gnd.n6781 gnd.n556 240.244
R5979 gnd.n6787 gnd.n556 240.244
R5980 gnd.n6787 gnd.n554 240.244
R5981 gnd.n6791 gnd.n554 240.244
R5982 gnd.n6791 gnd.n550 240.244
R5983 gnd.n6797 gnd.n550 240.244
R5984 gnd.n6797 gnd.n548 240.244
R5985 gnd.n6801 gnd.n548 240.244
R5986 gnd.n6801 gnd.n544 240.244
R5987 gnd.n6807 gnd.n544 240.244
R5988 gnd.n6807 gnd.n542 240.244
R5989 gnd.n6811 gnd.n542 240.244
R5990 gnd.n6811 gnd.n538 240.244
R5991 gnd.n6817 gnd.n538 240.244
R5992 gnd.n6817 gnd.n536 240.244
R5993 gnd.n6821 gnd.n536 240.244
R5994 gnd.n6821 gnd.n532 240.244
R5995 gnd.n6827 gnd.n532 240.244
R5996 gnd.n6827 gnd.n530 240.244
R5997 gnd.n6831 gnd.n530 240.244
R5998 gnd.n6831 gnd.n526 240.244
R5999 gnd.n6837 gnd.n526 240.244
R6000 gnd.n6837 gnd.n524 240.244
R6001 gnd.n6841 gnd.n524 240.244
R6002 gnd.n6841 gnd.n520 240.244
R6003 gnd.n6847 gnd.n520 240.244
R6004 gnd.n6847 gnd.n518 240.244
R6005 gnd.n6851 gnd.n518 240.244
R6006 gnd.n6851 gnd.n514 240.244
R6007 gnd.n6857 gnd.n514 240.244
R6008 gnd.n6857 gnd.n512 240.244
R6009 gnd.n6861 gnd.n512 240.244
R6010 gnd.n6861 gnd.n508 240.244
R6011 gnd.n6867 gnd.n508 240.244
R6012 gnd.n6867 gnd.n506 240.244
R6013 gnd.n6871 gnd.n506 240.244
R6014 gnd.n6871 gnd.n502 240.244
R6015 gnd.n6877 gnd.n502 240.244
R6016 gnd.n6877 gnd.n500 240.244
R6017 gnd.n6881 gnd.n500 240.244
R6018 gnd.n6881 gnd.n496 240.244
R6019 gnd.n6887 gnd.n496 240.244
R6020 gnd.n6887 gnd.n494 240.244
R6021 gnd.n6891 gnd.n494 240.244
R6022 gnd.n6891 gnd.n490 240.244
R6023 gnd.n6897 gnd.n490 240.244
R6024 gnd.n6897 gnd.n488 240.244
R6025 gnd.n6901 gnd.n488 240.244
R6026 gnd.n6901 gnd.n484 240.244
R6027 gnd.n6907 gnd.n484 240.244
R6028 gnd.n6907 gnd.n482 240.244
R6029 gnd.n6911 gnd.n482 240.244
R6030 gnd.n6911 gnd.n478 240.244
R6031 gnd.n6917 gnd.n478 240.244
R6032 gnd.n6917 gnd.n476 240.244
R6033 gnd.n6921 gnd.n476 240.244
R6034 gnd.n6921 gnd.n472 240.244
R6035 gnd.n6927 gnd.n472 240.244
R6036 gnd.n6927 gnd.n470 240.244
R6037 gnd.n6931 gnd.n470 240.244
R6038 gnd.n6931 gnd.n466 240.244
R6039 gnd.n6937 gnd.n466 240.244
R6040 gnd.n6937 gnd.n464 240.244
R6041 gnd.n6941 gnd.n464 240.244
R6042 gnd.n6941 gnd.n460 240.244
R6043 gnd.n6948 gnd.n460 240.244
R6044 gnd.n6948 gnd.n458 240.244
R6045 gnd.n6952 gnd.n458 240.244
R6046 gnd.n6952 gnd.n455 240.244
R6047 gnd.n6958 gnd.n453 240.244
R6048 gnd.n6962 gnd.n453 240.244
R6049 gnd.n6962 gnd.n449 240.244
R6050 gnd.n6968 gnd.n449 240.244
R6051 gnd.n6968 gnd.n447 240.244
R6052 gnd.n6972 gnd.n447 240.244
R6053 gnd.n6972 gnd.n443 240.244
R6054 gnd.n6978 gnd.n443 240.244
R6055 gnd.n6978 gnd.n441 240.244
R6056 gnd.n6982 gnd.n441 240.244
R6057 gnd.n6982 gnd.n437 240.244
R6058 gnd.n6988 gnd.n437 240.244
R6059 gnd.n6988 gnd.n435 240.244
R6060 gnd.n6992 gnd.n435 240.244
R6061 gnd.n6992 gnd.n431 240.244
R6062 gnd.n6998 gnd.n431 240.244
R6063 gnd.n6998 gnd.n429 240.244
R6064 gnd.n7002 gnd.n429 240.244
R6065 gnd.n7002 gnd.n425 240.244
R6066 gnd.n7008 gnd.n425 240.244
R6067 gnd.n7008 gnd.n423 240.244
R6068 gnd.n7012 gnd.n423 240.244
R6069 gnd.n7012 gnd.n419 240.244
R6070 gnd.n7018 gnd.n419 240.244
R6071 gnd.n7018 gnd.n417 240.244
R6072 gnd.n7022 gnd.n417 240.244
R6073 gnd.n7022 gnd.n413 240.244
R6074 gnd.n7028 gnd.n413 240.244
R6075 gnd.n7028 gnd.n411 240.244
R6076 gnd.n7032 gnd.n411 240.244
R6077 gnd.n7032 gnd.n407 240.244
R6078 gnd.n7038 gnd.n407 240.244
R6079 gnd.n7038 gnd.n405 240.244
R6080 gnd.n7042 gnd.n405 240.244
R6081 gnd.n7042 gnd.n401 240.244
R6082 gnd.n7048 gnd.n401 240.244
R6083 gnd.n7048 gnd.n399 240.244
R6084 gnd.n7052 gnd.n399 240.244
R6085 gnd.n7052 gnd.n395 240.244
R6086 gnd.n7058 gnd.n395 240.244
R6087 gnd.n7058 gnd.n393 240.244
R6088 gnd.n7062 gnd.n393 240.244
R6089 gnd.n7062 gnd.n389 240.244
R6090 gnd.n7068 gnd.n389 240.244
R6091 gnd.n7068 gnd.n387 240.244
R6092 gnd.n7072 gnd.n387 240.244
R6093 gnd.n7072 gnd.n383 240.244
R6094 gnd.n7078 gnd.n383 240.244
R6095 gnd.n7078 gnd.n381 240.244
R6096 gnd.n7082 gnd.n381 240.244
R6097 gnd.n7082 gnd.n377 240.244
R6098 gnd.n7088 gnd.n377 240.244
R6099 gnd.n7088 gnd.n375 240.244
R6100 gnd.n7092 gnd.n375 240.244
R6101 gnd.n7092 gnd.n371 240.244
R6102 gnd.n7098 gnd.n371 240.244
R6103 gnd.n7098 gnd.n369 240.244
R6104 gnd.n7102 gnd.n369 240.244
R6105 gnd.n7102 gnd.n365 240.244
R6106 gnd.n7108 gnd.n365 240.244
R6107 gnd.n7108 gnd.n363 240.244
R6108 gnd.n7112 gnd.n363 240.244
R6109 gnd.n7112 gnd.n359 240.244
R6110 gnd.n7118 gnd.n359 240.244
R6111 gnd.n7118 gnd.n357 240.244
R6112 gnd.n7122 gnd.n357 240.244
R6113 gnd.n7122 gnd.n353 240.244
R6114 gnd.n7128 gnd.n353 240.244
R6115 gnd.n7128 gnd.n351 240.244
R6116 gnd.n7132 gnd.n351 240.244
R6117 gnd.n7132 gnd.n347 240.244
R6118 gnd.n7138 gnd.n347 240.244
R6119 gnd.n7138 gnd.n345 240.244
R6120 gnd.n7142 gnd.n345 240.244
R6121 gnd.n7142 gnd.n341 240.244
R6122 gnd.n7148 gnd.n341 240.244
R6123 gnd.n7148 gnd.n339 240.244
R6124 gnd.n7152 gnd.n339 240.244
R6125 gnd.n7152 gnd.n335 240.244
R6126 gnd.n7158 gnd.n335 240.244
R6127 gnd.n7158 gnd.n333 240.244
R6128 gnd.n7163 gnd.n333 240.244
R6129 gnd.n7163 gnd.n329 240.244
R6130 gnd.n7170 gnd.n329 240.244
R6131 gnd.n2412 gnd.n2411 240.244
R6132 gnd.n2651 gnd.n2412 240.244
R6133 gnd.n2651 gnd.n2650 240.244
R6134 gnd.n2650 gnd.n2413 240.244
R6135 gnd.n2605 gnd.n2413 240.244
R6136 gnd.n2613 gnd.n2605 240.244
R6137 gnd.n2613 gnd.n2610 240.244
R6138 gnd.n2610 gnd.n2609 240.244
R6139 gnd.n2609 gnd.n2606 240.244
R6140 gnd.n2606 gnd.n2379 240.244
R6141 gnd.n2657 gnd.n2379 240.244
R6142 gnd.n2657 gnd.n2380 240.244
R6143 gnd.n2398 gnd.n2380 240.244
R6144 gnd.n2398 gnd.n2397 240.244
R6145 gnd.n2397 gnd.n2396 240.244
R6146 gnd.n2396 gnd.n2385 240.244
R6147 gnd.n2392 gnd.n2385 240.244
R6148 gnd.n2392 gnd.n2352 240.244
R6149 gnd.n2725 gnd.n2352 240.244
R6150 gnd.n2726 gnd.n2725 240.244
R6151 gnd.n2727 gnd.n2726 240.244
R6152 gnd.n2727 gnd.n2348 240.244
R6153 gnd.n2733 gnd.n2348 240.244
R6154 gnd.n2734 gnd.n2733 240.244
R6155 gnd.n2735 gnd.n2734 240.244
R6156 gnd.n2735 gnd.n2343 240.244
R6157 gnd.n2774 gnd.n2343 240.244
R6158 gnd.n2774 gnd.n2344 240.244
R6159 gnd.n2770 gnd.n2344 240.244
R6160 gnd.n2770 gnd.n2769 240.244
R6161 gnd.n2769 gnd.n2768 240.244
R6162 gnd.n2768 gnd.n2743 240.244
R6163 gnd.n2764 gnd.n2743 240.244
R6164 gnd.n2764 gnd.n2763 240.244
R6165 gnd.n2763 gnd.n2762 240.244
R6166 gnd.n2762 gnd.n2749 240.244
R6167 gnd.n2758 gnd.n2749 240.244
R6168 gnd.n2758 gnd.n2756 240.244
R6169 gnd.n2756 gnd.n2174 240.244
R6170 gnd.n3203 gnd.n2174 240.244
R6171 gnd.n3203 gnd.n2170 240.244
R6172 gnd.n3209 gnd.n2170 240.244
R6173 gnd.n3209 gnd.n2162 240.244
R6174 gnd.n3219 gnd.n2162 240.244
R6175 gnd.n3219 gnd.n2158 240.244
R6176 gnd.n3225 gnd.n2158 240.244
R6177 gnd.n3225 gnd.n2149 240.244
R6178 gnd.n3235 gnd.n2149 240.244
R6179 gnd.n3235 gnd.n2145 240.244
R6180 gnd.n3241 gnd.n2145 240.244
R6181 gnd.n3241 gnd.n2136 240.244
R6182 gnd.n3251 gnd.n2136 240.244
R6183 gnd.n3251 gnd.n2132 240.244
R6184 gnd.n3257 gnd.n2132 240.244
R6185 gnd.n3257 gnd.n2121 240.244
R6186 gnd.n3267 gnd.n2121 240.244
R6187 gnd.n3267 gnd.n2117 240.244
R6188 gnd.n3273 gnd.n2117 240.244
R6189 gnd.n3273 gnd.n2109 240.244
R6190 gnd.n3283 gnd.n2109 240.244
R6191 gnd.n3283 gnd.n2104 240.244
R6192 gnd.n3291 gnd.n2104 240.244
R6193 gnd.n3291 gnd.n2105 240.244
R6194 gnd.n2105 gnd.n2081 240.244
R6195 gnd.n3899 gnd.n2081 240.244
R6196 gnd.n3899 gnd.n2077 240.244
R6197 gnd.n3905 gnd.n2077 240.244
R6198 gnd.n3905 gnd.n2066 240.244
R6199 gnd.n3915 gnd.n2066 240.244
R6200 gnd.n3915 gnd.n2062 240.244
R6201 gnd.n3921 gnd.n2062 240.244
R6202 gnd.n3921 gnd.n2051 240.244
R6203 gnd.n3931 gnd.n2051 240.244
R6204 gnd.n3931 gnd.n2047 240.244
R6205 gnd.n3937 gnd.n2047 240.244
R6206 gnd.n3937 gnd.n2036 240.244
R6207 gnd.n3947 gnd.n2036 240.244
R6208 gnd.n3947 gnd.n2032 240.244
R6209 gnd.n3953 gnd.n2032 240.244
R6210 gnd.n3953 gnd.n2022 240.244
R6211 gnd.n3963 gnd.n2022 240.244
R6212 gnd.n3963 gnd.n2018 240.244
R6213 gnd.n3969 gnd.n2018 240.244
R6214 gnd.n3969 gnd.n2007 240.244
R6215 gnd.n3979 gnd.n2007 240.244
R6216 gnd.n3979 gnd.n2003 240.244
R6217 gnd.n3985 gnd.n2003 240.244
R6218 gnd.n3985 gnd.n1992 240.244
R6219 gnd.n3995 gnd.n1992 240.244
R6220 gnd.n3995 gnd.n1988 240.244
R6221 gnd.n4001 gnd.n1988 240.244
R6222 gnd.n4001 gnd.n1977 240.244
R6223 gnd.n4011 gnd.n1977 240.244
R6224 gnd.n4011 gnd.n1973 240.244
R6225 gnd.n4017 gnd.n1973 240.244
R6226 gnd.n4017 gnd.n1963 240.244
R6227 gnd.n4027 gnd.n1963 240.244
R6228 gnd.n4027 gnd.n1959 240.244
R6229 gnd.n4033 gnd.n1959 240.244
R6230 gnd.n4033 gnd.n1948 240.244
R6231 gnd.n4043 gnd.n1948 240.244
R6232 gnd.n4043 gnd.n1944 240.244
R6233 gnd.n4049 gnd.n1944 240.244
R6234 gnd.n4049 gnd.n1935 240.244
R6235 gnd.n4059 gnd.n1935 240.244
R6236 gnd.n4059 gnd.n1931 240.244
R6237 gnd.n4065 gnd.n1931 240.244
R6238 gnd.n4065 gnd.n1923 240.244
R6239 gnd.n4075 gnd.n1923 240.244
R6240 gnd.n4075 gnd.n1919 240.244
R6241 gnd.n4081 gnd.n1919 240.244
R6242 gnd.n4081 gnd.n1910 240.244
R6243 gnd.n4091 gnd.n1910 240.244
R6244 gnd.n4091 gnd.n1906 240.244
R6245 gnd.n4097 gnd.n1906 240.244
R6246 gnd.n4097 gnd.n1896 240.244
R6247 gnd.n4107 gnd.n1896 240.244
R6248 gnd.n4107 gnd.n1892 240.244
R6249 gnd.n4113 gnd.n1892 240.244
R6250 gnd.n4113 gnd.n1883 240.244
R6251 gnd.n4123 gnd.n1883 240.244
R6252 gnd.n4123 gnd.n1879 240.244
R6253 gnd.n4129 gnd.n1879 240.244
R6254 gnd.n4129 gnd.n1870 240.244
R6255 gnd.n4139 gnd.n1870 240.244
R6256 gnd.n4139 gnd.n1866 240.244
R6257 gnd.n4145 gnd.n1866 240.244
R6258 gnd.n4145 gnd.n1857 240.244
R6259 gnd.n4155 gnd.n1857 240.244
R6260 gnd.n4155 gnd.n1853 240.244
R6261 gnd.n4161 gnd.n1853 240.244
R6262 gnd.n4161 gnd.n1843 240.244
R6263 gnd.n4171 gnd.n1843 240.244
R6264 gnd.n4171 gnd.n1839 240.244
R6265 gnd.n4177 gnd.n1839 240.244
R6266 gnd.n4177 gnd.n1830 240.244
R6267 gnd.n4189 gnd.n1830 240.244
R6268 gnd.n4189 gnd.n1825 240.244
R6269 gnd.n4198 gnd.n1825 240.244
R6270 gnd.n4198 gnd.n1826 240.244
R6271 gnd.n1826 gnd.n1407 240.244
R6272 gnd.n4505 gnd.n1407 240.244
R6273 gnd.n4505 gnd.n1410 240.244
R6274 gnd.n4501 gnd.n1410 240.244
R6275 gnd.n4501 gnd.n1416 240.244
R6276 gnd.n1634 gnd.n1416 240.244
R6277 gnd.n1640 gnd.n1634 240.244
R6278 gnd.n1641 gnd.n1640 240.244
R6279 gnd.n4238 gnd.n1641 240.244
R6280 gnd.n4238 gnd.n1629 240.244
R6281 gnd.n4246 gnd.n1629 240.244
R6282 gnd.n4246 gnd.n1630 240.244
R6283 gnd.n1630 gnd.n1607 240.244
R6284 gnd.n4269 gnd.n1607 240.244
R6285 gnd.n4269 gnd.n1602 240.244
R6286 gnd.n4277 gnd.n1602 240.244
R6287 gnd.n4277 gnd.n1603 240.244
R6288 gnd.n1603 gnd.n1579 240.244
R6289 gnd.n4305 gnd.n1579 240.244
R6290 gnd.n4305 gnd.n1574 240.244
R6291 gnd.n4313 gnd.n1574 240.244
R6292 gnd.n4313 gnd.n1575 240.244
R6293 gnd.n1575 gnd.n1545 240.244
R6294 gnd.n4363 gnd.n1545 240.244
R6295 gnd.n4363 gnd.n1539 240.244
R6296 gnd.n4377 gnd.n1539 240.244
R6297 gnd.n4377 gnd.n1541 240.244
R6298 gnd.n4373 gnd.n1541 240.244
R6299 gnd.n4373 gnd.n4372 240.244
R6300 gnd.n4372 gnd.n315 240.244
R6301 gnd.n7190 gnd.n315 240.244
R6302 gnd.n7190 gnd.n316 240.244
R6303 gnd.n7185 gnd.n316 240.244
R6304 gnd.n7185 gnd.n7184 240.244
R6305 gnd.n7184 gnd.n322 240.244
R6306 gnd.n7179 gnd.n322 240.244
R6307 gnd.n7179 gnd.n7178 240.244
R6308 gnd.n7178 gnd.n7177 240.244
R6309 gnd.n7177 gnd.n324 240.244
R6310 gnd.n7173 gnd.n324 240.244
R6311 gnd.n7173 gnd.n7172 240.244
R6312 gnd.n6497 gnd.n727 240.244
R6313 gnd.n6497 gnd.n729 240.244
R6314 gnd.n6493 gnd.n729 240.244
R6315 gnd.n6493 gnd.n735 240.244
R6316 gnd.n6489 gnd.n735 240.244
R6317 gnd.n6489 gnd.n737 240.244
R6318 gnd.n6485 gnd.n737 240.244
R6319 gnd.n6485 gnd.n743 240.244
R6320 gnd.n6481 gnd.n743 240.244
R6321 gnd.n6481 gnd.n745 240.244
R6322 gnd.n6477 gnd.n745 240.244
R6323 gnd.n6477 gnd.n751 240.244
R6324 gnd.n6473 gnd.n751 240.244
R6325 gnd.n6473 gnd.n753 240.244
R6326 gnd.n6469 gnd.n753 240.244
R6327 gnd.n6469 gnd.n759 240.244
R6328 gnd.n6465 gnd.n759 240.244
R6329 gnd.n6465 gnd.n761 240.244
R6330 gnd.n6461 gnd.n761 240.244
R6331 gnd.n6461 gnd.n767 240.244
R6332 gnd.n6457 gnd.n767 240.244
R6333 gnd.n6457 gnd.n769 240.244
R6334 gnd.n6453 gnd.n769 240.244
R6335 gnd.n6453 gnd.n775 240.244
R6336 gnd.n6449 gnd.n775 240.244
R6337 gnd.n6449 gnd.n777 240.244
R6338 gnd.n6445 gnd.n777 240.244
R6339 gnd.n6445 gnd.n783 240.244
R6340 gnd.n6441 gnd.n783 240.244
R6341 gnd.n6441 gnd.n785 240.244
R6342 gnd.n6437 gnd.n785 240.244
R6343 gnd.n6437 gnd.n791 240.244
R6344 gnd.n6433 gnd.n791 240.244
R6345 gnd.n6433 gnd.n793 240.244
R6346 gnd.n6429 gnd.n793 240.244
R6347 gnd.n6429 gnd.n799 240.244
R6348 gnd.n6425 gnd.n799 240.244
R6349 gnd.n6425 gnd.n801 240.244
R6350 gnd.n6421 gnd.n801 240.244
R6351 gnd.n6421 gnd.n807 240.244
R6352 gnd.n6417 gnd.n807 240.244
R6353 gnd.n6417 gnd.n809 240.244
R6354 gnd.n6413 gnd.n809 240.244
R6355 gnd.n6413 gnd.n815 240.244
R6356 gnd.n6409 gnd.n815 240.244
R6357 gnd.n6409 gnd.n817 240.244
R6358 gnd.n6405 gnd.n817 240.244
R6359 gnd.n6405 gnd.n823 240.244
R6360 gnd.n6401 gnd.n823 240.244
R6361 gnd.n6401 gnd.n825 240.244
R6362 gnd.n6397 gnd.n825 240.244
R6363 gnd.n6397 gnd.n831 240.244
R6364 gnd.n6393 gnd.n831 240.244
R6365 gnd.n6393 gnd.n833 240.244
R6366 gnd.n6389 gnd.n833 240.244
R6367 gnd.n6389 gnd.n839 240.244
R6368 gnd.n6385 gnd.n839 240.244
R6369 gnd.n6385 gnd.n841 240.244
R6370 gnd.n6381 gnd.n841 240.244
R6371 gnd.n6381 gnd.n847 240.244
R6372 gnd.n6377 gnd.n847 240.244
R6373 gnd.n6377 gnd.n849 240.244
R6374 gnd.n6373 gnd.n849 240.244
R6375 gnd.n6373 gnd.n855 240.244
R6376 gnd.n6369 gnd.n855 240.244
R6377 gnd.n6369 gnd.n857 240.244
R6378 gnd.n6365 gnd.n857 240.244
R6379 gnd.n6365 gnd.n863 240.244
R6380 gnd.n6361 gnd.n863 240.244
R6381 gnd.n6361 gnd.n865 240.244
R6382 gnd.n6357 gnd.n865 240.244
R6383 gnd.n6357 gnd.n871 240.244
R6384 gnd.n6353 gnd.n871 240.244
R6385 gnd.n6353 gnd.n873 240.244
R6386 gnd.n6349 gnd.n873 240.244
R6387 gnd.n6349 gnd.n879 240.244
R6388 gnd.n6345 gnd.n879 240.244
R6389 gnd.n6345 gnd.n881 240.244
R6390 gnd.n6341 gnd.n881 240.244
R6391 gnd.n6341 gnd.n887 240.244
R6392 gnd.n6337 gnd.n887 240.244
R6393 gnd.n6337 gnd.n889 240.244
R6394 gnd.n6333 gnd.n889 240.244
R6395 gnd.n6333 gnd.n895 240.244
R6396 gnd.n1280 gnd.n1279 240.244
R6397 gnd.n1281 gnd.n1280 240.244
R6398 gnd.n2163 gnd.n1281 240.244
R6399 gnd.n2163 gnd.n1284 240.244
R6400 gnd.n1285 gnd.n1284 240.244
R6401 gnd.n1286 gnd.n1285 240.244
R6402 gnd.n2150 gnd.n1286 240.244
R6403 gnd.n2150 gnd.n1289 240.244
R6404 gnd.n1290 gnd.n1289 240.244
R6405 gnd.n1291 gnd.n1290 240.244
R6406 gnd.n2143 gnd.n1291 240.244
R6407 gnd.n2143 gnd.n1294 240.244
R6408 gnd.n1295 gnd.n1294 240.244
R6409 gnd.n1296 gnd.n1295 240.244
R6410 gnd.n2130 gnd.n1296 240.244
R6411 gnd.n2130 gnd.n1299 240.244
R6412 gnd.n1300 gnd.n1299 240.244
R6413 gnd.n1301 gnd.n1300 240.244
R6414 gnd.n2903 gnd.n1301 240.244
R6415 gnd.n2903 gnd.n1304 240.244
R6416 gnd.n1305 gnd.n1304 240.244
R6417 gnd.n1306 gnd.n1305 240.244
R6418 gnd.n3021 gnd.n1306 240.244
R6419 gnd.n3021 gnd.n1309 240.244
R6420 gnd.n1310 gnd.n1309 240.244
R6421 gnd.n1311 gnd.n1310 240.244
R6422 gnd.n2075 gnd.n1311 240.244
R6423 gnd.n2075 gnd.n1314 240.244
R6424 gnd.n1315 gnd.n1314 240.244
R6425 gnd.n1316 gnd.n1315 240.244
R6426 gnd.n2060 gnd.n1316 240.244
R6427 gnd.n2060 gnd.n1319 240.244
R6428 gnd.n1320 gnd.n1319 240.244
R6429 gnd.n1321 gnd.n1320 240.244
R6430 gnd.n2045 gnd.n1321 240.244
R6431 gnd.n2045 gnd.n1324 240.244
R6432 gnd.n1325 gnd.n1324 240.244
R6433 gnd.n1326 gnd.n1325 240.244
R6434 gnd.n2030 gnd.n1326 240.244
R6435 gnd.n2030 gnd.n1329 240.244
R6436 gnd.n1330 gnd.n1329 240.244
R6437 gnd.n1331 gnd.n1330 240.244
R6438 gnd.n2016 gnd.n1331 240.244
R6439 gnd.n2016 gnd.n1334 240.244
R6440 gnd.n1335 gnd.n1334 240.244
R6441 gnd.n1336 gnd.n1335 240.244
R6442 gnd.n2001 gnd.n1336 240.244
R6443 gnd.n2001 gnd.n1339 240.244
R6444 gnd.n1340 gnd.n1339 240.244
R6445 gnd.n1341 gnd.n1340 240.244
R6446 gnd.n1986 gnd.n1341 240.244
R6447 gnd.n1986 gnd.n1344 240.244
R6448 gnd.n1345 gnd.n1344 240.244
R6449 gnd.n1346 gnd.n1345 240.244
R6450 gnd.n1971 gnd.n1346 240.244
R6451 gnd.n1971 gnd.n1349 240.244
R6452 gnd.n1350 gnd.n1349 240.244
R6453 gnd.n1351 gnd.n1350 240.244
R6454 gnd.n1956 gnd.n1351 240.244
R6455 gnd.n1956 gnd.n1354 240.244
R6456 gnd.n1355 gnd.n1354 240.244
R6457 gnd.n1356 gnd.n1355 240.244
R6458 gnd.n1942 gnd.n1356 240.244
R6459 gnd.n1942 gnd.n1359 240.244
R6460 gnd.n1360 gnd.n1359 240.244
R6461 gnd.n1361 gnd.n1360 240.244
R6462 gnd.n1930 gnd.n1361 240.244
R6463 gnd.n1930 gnd.n1364 240.244
R6464 gnd.n1365 gnd.n1364 240.244
R6465 gnd.n1366 gnd.n1365 240.244
R6466 gnd.n1918 gnd.n1366 240.244
R6467 gnd.n1918 gnd.n1369 240.244
R6468 gnd.n1370 gnd.n1369 240.244
R6469 gnd.n1371 gnd.n1370 240.244
R6470 gnd.n1905 gnd.n1371 240.244
R6471 gnd.n1905 gnd.n1374 240.244
R6472 gnd.n1375 gnd.n1374 240.244
R6473 gnd.n1376 gnd.n1375 240.244
R6474 gnd.n1891 gnd.n1376 240.244
R6475 gnd.n1891 gnd.n1379 240.244
R6476 gnd.n1380 gnd.n1379 240.244
R6477 gnd.n1381 gnd.n1380 240.244
R6478 gnd.n1877 gnd.n1381 240.244
R6479 gnd.n1877 gnd.n1384 240.244
R6480 gnd.n1385 gnd.n1384 240.244
R6481 gnd.n1386 gnd.n1385 240.244
R6482 gnd.n1865 gnd.n1386 240.244
R6483 gnd.n1865 gnd.n1389 240.244
R6484 gnd.n1390 gnd.n1389 240.244
R6485 gnd.n1391 gnd.n1390 240.244
R6486 gnd.n1852 gnd.n1391 240.244
R6487 gnd.n1852 gnd.n1394 240.244
R6488 gnd.n1395 gnd.n1394 240.244
R6489 gnd.n1396 gnd.n1395 240.244
R6490 gnd.n1838 gnd.n1396 240.244
R6491 gnd.n1838 gnd.n1399 240.244
R6492 gnd.n1400 gnd.n1399 240.244
R6493 gnd.n1401 gnd.n1400 240.244
R6494 gnd.n1824 gnd.n1401 240.244
R6495 gnd.n1824 gnd.n1404 240.244
R6496 gnd.n4508 gnd.n1404 240.244
R6497 gnd.n2195 gnd.n2194 240.244
R6498 gnd.n2205 gnd.n2194 240.244
R6499 gnd.n2207 gnd.n2206 240.244
R6500 gnd.n2215 gnd.n2214 240.244
R6501 gnd.n2223 gnd.n2222 240.244
R6502 gnd.n2225 gnd.n2224 240.244
R6503 gnd.n2233 gnd.n2232 240.244
R6504 gnd.n2243 gnd.n2242 240.244
R6505 gnd.n2245 gnd.n2244 240.244
R6506 gnd.n2800 gnd.n2799 240.244
R6507 gnd.n2802 gnd.n2801 240.244
R6508 gnd.n2806 gnd.n2805 240.244
R6509 gnd.n2812 gnd.n2807 240.244
R6510 gnd.n3195 gnd.n2180 240.244
R6511 gnd.n3201 gnd.n2169 240.244
R6512 gnd.n3211 gnd.n2169 240.244
R6513 gnd.n3211 gnd.n2165 240.244
R6514 gnd.n3217 gnd.n2165 240.244
R6515 gnd.n3217 gnd.n2156 240.244
R6516 gnd.n3227 gnd.n2156 240.244
R6517 gnd.n3227 gnd.n2152 240.244
R6518 gnd.n3233 gnd.n2152 240.244
R6519 gnd.n3233 gnd.n2141 240.244
R6520 gnd.n3243 gnd.n2141 240.244
R6521 gnd.n3243 gnd.n2137 240.244
R6522 gnd.n3249 gnd.n2137 240.244
R6523 gnd.n3249 gnd.n2128 240.244
R6524 gnd.n3259 gnd.n2128 240.244
R6525 gnd.n3259 gnd.n2124 240.244
R6526 gnd.n3265 gnd.n2124 240.244
R6527 gnd.n3265 gnd.n2115 240.244
R6528 gnd.n3275 gnd.n2115 240.244
R6529 gnd.n3275 gnd.n2111 240.244
R6530 gnd.n3281 gnd.n2111 240.244
R6531 gnd.n3281 gnd.n2101 240.244
R6532 gnd.n3293 gnd.n2101 240.244
R6533 gnd.n3293 gnd.n2096 240.244
R6534 gnd.n3300 gnd.n2096 240.244
R6535 gnd.n3300 gnd.n2083 240.244
R6536 gnd.n2083 gnd.n2073 240.244
R6537 gnd.n3907 gnd.n2073 240.244
R6538 gnd.n3907 gnd.n2069 240.244
R6539 gnd.n3913 gnd.n2069 240.244
R6540 gnd.n3913 gnd.n2058 240.244
R6541 gnd.n3923 gnd.n2058 240.244
R6542 gnd.n3923 gnd.n2054 240.244
R6543 gnd.n3929 gnd.n2054 240.244
R6544 gnd.n3929 gnd.n2043 240.244
R6545 gnd.n3939 gnd.n2043 240.244
R6546 gnd.n3939 gnd.n2039 240.244
R6547 gnd.n3945 gnd.n2039 240.244
R6548 gnd.n3945 gnd.n2029 240.244
R6549 gnd.n3955 gnd.n2029 240.244
R6550 gnd.n3955 gnd.n2025 240.244
R6551 gnd.n3961 gnd.n2025 240.244
R6552 gnd.n3961 gnd.n2014 240.244
R6553 gnd.n3971 gnd.n2014 240.244
R6554 gnd.n3971 gnd.n2010 240.244
R6555 gnd.n3977 gnd.n2010 240.244
R6556 gnd.n3977 gnd.n1999 240.244
R6557 gnd.n3987 gnd.n1999 240.244
R6558 gnd.n3987 gnd.n1995 240.244
R6559 gnd.n3993 gnd.n1995 240.244
R6560 gnd.n3993 gnd.n1984 240.244
R6561 gnd.n4003 gnd.n1984 240.244
R6562 gnd.n4003 gnd.n1980 240.244
R6563 gnd.n4009 gnd.n1980 240.244
R6564 gnd.n4009 gnd.n1969 240.244
R6565 gnd.n4019 gnd.n1969 240.244
R6566 gnd.n4019 gnd.n1965 240.244
R6567 gnd.n4025 gnd.n1965 240.244
R6568 gnd.n4025 gnd.n1954 240.244
R6569 gnd.n4035 gnd.n1954 240.244
R6570 gnd.n4035 gnd.n1950 240.244
R6571 gnd.n4041 gnd.n1950 240.244
R6572 gnd.n4041 gnd.n1941 240.244
R6573 gnd.n4051 gnd.n1941 240.244
R6574 gnd.n4051 gnd.n1937 240.244
R6575 gnd.n4057 gnd.n1937 240.244
R6576 gnd.n4057 gnd.n1929 240.244
R6577 gnd.n4067 gnd.n1929 240.244
R6578 gnd.n4067 gnd.n1925 240.244
R6579 gnd.n4073 gnd.n1925 240.244
R6580 gnd.n4073 gnd.n1916 240.244
R6581 gnd.n4083 gnd.n1916 240.244
R6582 gnd.n4083 gnd.n1912 240.244
R6583 gnd.n4089 gnd.n1912 240.244
R6584 gnd.n4089 gnd.n1903 240.244
R6585 gnd.n4099 gnd.n1903 240.244
R6586 gnd.n4099 gnd.n1899 240.244
R6587 gnd.n4105 gnd.n1899 240.244
R6588 gnd.n4105 gnd.n1889 240.244
R6589 gnd.n4115 gnd.n1889 240.244
R6590 gnd.n4115 gnd.n1885 240.244
R6591 gnd.n4121 gnd.n1885 240.244
R6592 gnd.n4121 gnd.n1875 240.244
R6593 gnd.n4131 gnd.n1875 240.244
R6594 gnd.n4131 gnd.n1871 240.244
R6595 gnd.n4137 gnd.n1871 240.244
R6596 gnd.n4137 gnd.n1863 240.244
R6597 gnd.n4147 gnd.n1863 240.244
R6598 gnd.n4147 gnd.n1859 240.244
R6599 gnd.n4153 gnd.n1859 240.244
R6600 gnd.n4153 gnd.n1850 240.244
R6601 gnd.n4163 gnd.n1850 240.244
R6602 gnd.n4163 gnd.n1846 240.244
R6603 gnd.n4169 gnd.n1846 240.244
R6604 gnd.n4169 gnd.n1837 240.244
R6605 gnd.n4179 gnd.n1837 240.244
R6606 gnd.n4179 gnd.n1832 240.244
R6607 gnd.n4187 gnd.n1832 240.244
R6608 gnd.n4187 gnd.n1822 240.244
R6609 gnd.n4200 gnd.n1822 240.244
R6610 gnd.n4201 gnd.n4200 240.244
R6611 gnd.n4201 gnd.n1408 240.244
R6612 gnd.n1737 gnd.n1736 240.244
R6613 gnd.n1740 gnd.n1739 240.244
R6614 gnd.n1756 gnd.n1755 240.244
R6615 gnd.n1759 gnd.n1758 240.244
R6616 gnd.n1775 gnd.n1774 240.244
R6617 gnd.n1778 gnd.n1777 240.244
R6618 gnd.n1791 gnd.n1790 240.244
R6619 gnd.n1794 gnd.n1793 240.244
R6620 gnd.n1805 gnd.n1804 240.244
R6621 gnd.n1808 gnd.n1807 240.244
R6622 gnd.n1813 gnd.n1810 240.244
R6623 gnd.n1816 gnd.n1815 240.244
R6624 gnd.n4206 gnd.n1818 240.244
R6625 gnd.n4209 gnd.n4208 240.244
R6626 gnd.n2914 gnd.n2913 240.132
R6627 gnd.n3507 gnd.n3506 240.132
R6628 gnd.n6500 gnd.n723 225.874
R6629 gnd.n6508 gnd.n723 225.874
R6630 gnd.n6509 gnd.n6508 225.874
R6631 gnd.n6510 gnd.n6509 225.874
R6632 gnd.n6510 gnd.n717 225.874
R6633 gnd.n6518 gnd.n717 225.874
R6634 gnd.n6519 gnd.n6518 225.874
R6635 gnd.n6520 gnd.n6519 225.874
R6636 gnd.n6520 gnd.n711 225.874
R6637 gnd.n6528 gnd.n711 225.874
R6638 gnd.n6529 gnd.n6528 225.874
R6639 gnd.n6530 gnd.n6529 225.874
R6640 gnd.n6530 gnd.n705 225.874
R6641 gnd.n6538 gnd.n705 225.874
R6642 gnd.n6539 gnd.n6538 225.874
R6643 gnd.n6540 gnd.n6539 225.874
R6644 gnd.n6540 gnd.n699 225.874
R6645 gnd.n6548 gnd.n699 225.874
R6646 gnd.n6549 gnd.n6548 225.874
R6647 gnd.n6550 gnd.n6549 225.874
R6648 gnd.n6550 gnd.n693 225.874
R6649 gnd.n6558 gnd.n693 225.874
R6650 gnd.n6559 gnd.n6558 225.874
R6651 gnd.n6560 gnd.n6559 225.874
R6652 gnd.n6560 gnd.n687 225.874
R6653 gnd.n6568 gnd.n687 225.874
R6654 gnd.n6569 gnd.n6568 225.874
R6655 gnd.n6570 gnd.n6569 225.874
R6656 gnd.n6570 gnd.n681 225.874
R6657 gnd.n6578 gnd.n681 225.874
R6658 gnd.n6579 gnd.n6578 225.874
R6659 gnd.n6580 gnd.n6579 225.874
R6660 gnd.n6580 gnd.n675 225.874
R6661 gnd.n6588 gnd.n675 225.874
R6662 gnd.n6589 gnd.n6588 225.874
R6663 gnd.n6590 gnd.n6589 225.874
R6664 gnd.n6590 gnd.n669 225.874
R6665 gnd.n6598 gnd.n669 225.874
R6666 gnd.n6599 gnd.n6598 225.874
R6667 gnd.n6600 gnd.n6599 225.874
R6668 gnd.n6600 gnd.n663 225.874
R6669 gnd.n6608 gnd.n663 225.874
R6670 gnd.n6609 gnd.n6608 225.874
R6671 gnd.n6610 gnd.n6609 225.874
R6672 gnd.n6610 gnd.n657 225.874
R6673 gnd.n6618 gnd.n657 225.874
R6674 gnd.n6619 gnd.n6618 225.874
R6675 gnd.n6620 gnd.n6619 225.874
R6676 gnd.n6620 gnd.n651 225.874
R6677 gnd.n6628 gnd.n651 225.874
R6678 gnd.n6629 gnd.n6628 225.874
R6679 gnd.n6630 gnd.n6629 225.874
R6680 gnd.n6630 gnd.n645 225.874
R6681 gnd.n6638 gnd.n645 225.874
R6682 gnd.n6639 gnd.n6638 225.874
R6683 gnd.n6640 gnd.n6639 225.874
R6684 gnd.n6640 gnd.n639 225.874
R6685 gnd.n6648 gnd.n639 225.874
R6686 gnd.n6649 gnd.n6648 225.874
R6687 gnd.n6650 gnd.n6649 225.874
R6688 gnd.n6650 gnd.n633 225.874
R6689 gnd.n6658 gnd.n633 225.874
R6690 gnd.n6659 gnd.n6658 225.874
R6691 gnd.n6660 gnd.n6659 225.874
R6692 gnd.n6660 gnd.n627 225.874
R6693 gnd.n6668 gnd.n627 225.874
R6694 gnd.n6669 gnd.n6668 225.874
R6695 gnd.n6670 gnd.n6669 225.874
R6696 gnd.n6670 gnd.n621 225.874
R6697 gnd.n6678 gnd.n621 225.874
R6698 gnd.n6679 gnd.n6678 225.874
R6699 gnd.n6680 gnd.n6679 225.874
R6700 gnd.n6680 gnd.n615 225.874
R6701 gnd.n6688 gnd.n615 225.874
R6702 gnd.n6689 gnd.n6688 225.874
R6703 gnd.n6690 gnd.n6689 225.874
R6704 gnd.n6690 gnd.n609 225.874
R6705 gnd.n6698 gnd.n609 225.874
R6706 gnd.n6699 gnd.n6698 225.874
R6707 gnd.n6700 gnd.n6699 225.874
R6708 gnd.n6700 gnd.n603 225.874
R6709 gnd.n6708 gnd.n603 225.874
R6710 gnd.n6709 gnd.n6708 225.874
R6711 gnd.n6710 gnd.n6709 225.874
R6712 gnd.n6710 gnd.n597 225.874
R6713 gnd.n6718 gnd.n597 225.874
R6714 gnd.n6719 gnd.n6718 225.874
R6715 gnd.n6720 gnd.n6719 225.874
R6716 gnd.n6720 gnd.n591 225.874
R6717 gnd.n6728 gnd.n591 225.874
R6718 gnd.n6729 gnd.n6728 225.874
R6719 gnd.n6730 gnd.n6729 225.874
R6720 gnd.n6730 gnd.n585 225.874
R6721 gnd.n6738 gnd.n585 225.874
R6722 gnd.n6739 gnd.n6738 225.874
R6723 gnd.n6740 gnd.n6739 225.874
R6724 gnd.n6740 gnd.n579 225.874
R6725 gnd.n6748 gnd.n579 225.874
R6726 gnd.n6749 gnd.n6748 225.874
R6727 gnd.n6750 gnd.n6749 225.874
R6728 gnd.n6750 gnd.n573 225.874
R6729 gnd.n6758 gnd.n573 225.874
R6730 gnd.n6759 gnd.n6758 225.874
R6731 gnd.n6760 gnd.n6759 225.874
R6732 gnd.n6760 gnd.n567 225.874
R6733 gnd.n6768 gnd.n567 225.874
R6734 gnd.n6769 gnd.n6768 225.874
R6735 gnd.n6770 gnd.n6769 225.874
R6736 gnd.n6770 gnd.n561 225.874
R6737 gnd.n6778 gnd.n561 225.874
R6738 gnd.n6779 gnd.n6778 225.874
R6739 gnd.n6780 gnd.n6779 225.874
R6740 gnd.n6780 gnd.n555 225.874
R6741 gnd.n6788 gnd.n555 225.874
R6742 gnd.n6789 gnd.n6788 225.874
R6743 gnd.n6790 gnd.n6789 225.874
R6744 gnd.n6790 gnd.n549 225.874
R6745 gnd.n6798 gnd.n549 225.874
R6746 gnd.n6799 gnd.n6798 225.874
R6747 gnd.n6800 gnd.n6799 225.874
R6748 gnd.n6800 gnd.n543 225.874
R6749 gnd.n6808 gnd.n543 225.874
R6750 gnd.n6809 gnd.n6808 225.874
R6751 gnd.n6810 gnd.n6809 225.874
R6752 gnd.n6810 gnd.n537 225.874
R6753 gnd.n6818 gnd.n537 225.874
R6754 gnd.n6819 gnd.n6818 225.874
R6755 gnd.n6820 gnd.n6819 225.874
R6756 gnd.n6820 gnd.n531 225.874
R6757 gnd.n6828 gnd.n531 225.874
R6758 gnd.n6829 gnd.n6828 225.874
R6759 gnd.n6830 gnd.n6829 225.874
R6760 gnd.n6830 gnd.n525 225.874
R6761 gnd.n6838 gnd.n525 225.874
R6762 gnd.n6839 gnd.n6838 225.874
R6763 gnd.n6840 gnd.n6839 225.874
R6764 gnd.n6840 gnd.n519 225.874
R6765 gnd.n6848 gnd.n519 225.874
R6766 gnd.n6849 gnd.n6848 225.874
R6767 gnd.n6850 gnd.n6849 225.874
R6768 gnd.n6850 gnd.n513 225.874
R6769 gnd.n6858 gnd.n513 225.874
R6770 gnd.n6859 gnd.n6858 225.874
R6771 gnd.n6860 gnd.n6859 225.874
R6772 gnd.n6860 gnd.n507 225.874
R6773 gnd.n6868 gnd.n507 225.874
R6774 gnd.n6869 gnd.n6868 225.874
R6775 gnd.n6870 gnd.n6869 225.874
R6776 gnd.n6870 gnd.n501 225.874
R6777 gnd.n6878 gnd.n501 225.874
R6778 gnd.n6879 gnd.n6878 225.874
R6779 gnd.n6880 gnd.n6879 225.874
R6780 gnd.n6880 gnd.n495 225.874
R6781 gnd.n6888 gnd.n495 225.874
R6782 gnd.n6889 gnd.n6888 225.874
R6783 gnd.n6890 gnd.n6889 225.874
R6784 gnd.n6890 gnd.n489 225.874
R6785 gnd.n6898 gnd.n489 225.874
R6786 gnd.n6899 gnd.n6898 225.874
R6787 gnd.n6900 gnd.n6899 225.874
R6788 gnd.n6900 gnd.n483 225.874
R6789 gnd.n6908 gnd.n483 225.874
R6790 gnd.n6909 gnd.n6908 225.874
R6791 gnd.n6910 gnd.n6909 225.874
R6792 gnd.n6910 gnd.n477 225.874
R6793 gnd.n6918 gnd.n477 225.874
R6794 gnd.n6919 gnd.n6918 225.874
R6795 gnd.n6920 gnd.n6919 225.874
R6796 gnd.n6920 gnd.n471 225.874
R6797 gnd.n6928 gnd.n471 225.874
R6798 gnd.n6929 gnd.n6928 225.874
R6799 gnd.n6930 gnd.n6929 225.874
R6800 gnd.n6930 gnd.n465 225.874
R6801 gnd.n6938 gnd.n465 225.874
R6802 gnd.n6939 gnd.n6938 225.874
R6803 gnd.n6940 gnd.n6939 225.874
R6804 gnd.n6940 gnd.n459 225.874
R6805 gnd.n6949 gnd.n459 225.874
R6806 gnd.n6950 gnd.n6949 225.874
R6807 gnd.n6951 gnd.n6950 225.874
R6808 gnd.n6951 gnd.n454 225.874
R6809 gnd.n5359 gnd.t110 224.174
R6810 gnd.n4980 gnd.t69 224.174
R6811 gnd.n1467 gnd.n1424 199.319
R6812 gnd.n1467 gnd.n1425 199.319
R6813 gnd.n2307 gnd.n2277 199.319
R6814 gnd.n2307 gnd.n2276 199.319
R6815 gnd.n2915 gnd.n2912 186.49
R6816 gnd.n3508 gnd.n3505 186.49
R6817 gnd.n6153 gnd.n6152 185
R6818 gnd.n6151 gnd.n6150 185
R6819 gnd.n6130 gnd.n6129 185
R6820 gnd.n6145 gnd.n6144 185
R6821 gnd.n6143 gnd.n6142 185
R6822 gnd.n6134 gnd.n6133 185
R6823 gnd.n6137 gnd.n6136 185
R6824 gnd.n6121 gnd.n6120 185
R6825 gnd.n6119 gnd.n6118 185
R6826 gnd.n6098 gnd.n6097 185
R6827 gnd.n6113 gnd.n6112 185
R6828 gnd.n6111 gnd.n6110 185
R6829 gnd.n6102 gnd.n6101 185
R6830 gnd.n6105 gnd.n6104 185
R6831 gnd.n6089 gnd.n6088 185
R6832 gnd.n6087 gnd.n6086 185
R6833 gnd.n6066 gnd.n6065 185
R6834 gnd.n6081 gnd.n6080 185
R6835 gnd.n6079 gnd.n6078 185
R6836 gnd.n6070 gnd.n6069 185
R6837 gnd.n6073 gnd.n6072 185
R6838 gnd.n6058 gnd.n6057 185
R6839 gnd.n6056 gnd.n6055 185
R6840 gnd.n6035 gnd.n6034 185
R6841 gnd.n6050 gnd.n6049 185
R6842 gnd.n6048 gnd.n6047 185
R6843 gnd.n6039 gnd.n6038 185
R6844 gnd.n6042 gnd.n6041 185
R6845 gnd.n6026 gnd.n6025 185
R6846 gnd.n6024 gnd.n6023 185
R6847 gnd.n6003 gnd.n6002 185
R6848 gnd.n6018 gnd.n6017 185
R6849 gnd.n6016 gnd.n6015 185
R6850 gnd.n6007 gnd.n6006 185
R6851 gnd.n6010 gnd.n6009 185
R6852 gnd.n5994 gnd.n5993 185
R6853 gnd.n5992 gnd.n5991 185
R6854 gnd.n5971 gnd.n5970 185
R6855 gnd.n5986 gnd.n5985 185
R6856 gnd.n5984 gnd.n5983 185
R6857 gnd.n5975 gnd.n5974 185
R6858 gnd.n5978 gnd.n5977 185
R6859 gnd.n5962 gnd.n5961 185
R6860 gnd.n5960 gnd.n5959 185
R6861 gnd.n5939 gnd.n5938 185
R6862 gnd.n5954 gnd.n5953 185
R6863 gnd.n5952 gnd.n5951 185
R6864 gnd.n5943 gnd.n5942 185
R6865 gnd.n5946 gnd.n5945 185
R6866 gnd.n5931 gnd.n5930 185
R6867 gnd.n5929 gnd.n5928 185
R6868 gnd.n5908 gnd.n5907 185
R6869 gnd.n5923 gnd.n5922 185
R6870 gnd.n5921 gnd.n5920 185
R6871 gnd.n5912 gnd.n5911 185
R6872 gnd.n5915 gnd.n5914 185
R6873 gnd.n5360 gnd.t109 178.987
R6874 gnd.n4981 gnd.t70 178.987
R6875 gnd.n1 gnd.t16 170.774
R6876 gnd.n9 gnd.t236 170.103
R6877 gnd.n8 gnd.t326 170.103
R6878 gnd.n7 gnd.t253 170.103
R6879 gnd.n6 gnd.t300 170.103
R6880 gnd.n5 gnd.t171 170.103
R6881 gnd.n4 gnd.t264 170.103
R6882 gnd.n3 gnd.t304 170.103
R6883 gnd.n2 gnd.t50 170.103
R6884 gnd.n1 gnd.t302 170.103
R6885 gnd.n3682 gnd.n3681 163.367
R6886 gnd.n3679 gnd.n3518 163.367
R6887 gnd.n3675 gnd.n3674 163.367
R6888 gnd.n3672 gnd.n3521 163.367
R6889 gnd.n3668 gnd.n3667 163.367
R6890 gnd.n3665 gnd.n3524 163.367
R6891 gnd.n3661 gnd.n3660 163.367
R6892 gnd.n3658 gnd.n3527 163.367
R6893 gnd.n3654 gnd.n3653 163.367
R6894 gnd.n3651 gnd.n3530 163.367
R6895 gnd.n3647 gnd.n3646 163.367
R6896 gnd.n3644 gnd.n3533 163.367
R6897 gnd.n3640 gnd.n3639 163.367
R6898 gnd.n3637 gnd.n3536 163.367
R6899 gnd.n3632 gnd.n3631 163.367
R6900 gnd.n3629 gnd.n3627 163.367
R6901 gnd.n3624 gnd.n3623 163.367
R6902 gnd.n3621 gnd.n3542 163.367
R6903 gnd.n3616 gnd.n3615 163.367
R6904 gnd.n3613 gnd.n3547 163.367
R6905 gnd.n3609 gnd.n3608 163.367
R6906 gnd.n3606 gnd.n3550 163.367
R6907 gnd.n3602 gnd.n3601 163.367
R6908 gnd.n3599 gnd.n3553 163.367
R6909 gnd.n3595 gnd.n3594 163.367
R6910 gnd.n3592 gnd.n3556 163.367
R6911 gnd.n3588 gnd.n3587 163.367
R6912 gnd.n3585 gnd.n3559 163.367
R6913 gnd.n3581 gnd.n3580 163.367
R6914 gnd.n3578 gnd.n3562 163.367
R6915 gnd.n3574 gnd.n3573 163.367
R6916 gnd.n3571 gnd.n3565 163.367
R6917 gnd.n3045 gnd.n3044 163.367
R6918 gnd.n3044 gnd.n2901 163.367
R6919 gnd.n3014 gnd.n2901 163.367
R6920 gnd.n3034 gnd.n3014 163.367
R6921 gnd.n3034 gnd.n3015 163.367
R6922 gnd.n3030 gnd.n3015 163.367
R6923 gnd.n3030 gnd.n3029 163.367
R6924 gnd.n3029 gnd.n3020 163.367
R6925 gnd.n3020 gnd.n2084 163.367
R6926 gnd.n3897 gnd.n2084 163.367
R6927 gnd.n3897 gnd.n2085 163.367
R6928 gnd.n3893 gnd.n2085 163.367
R6929 gnd.n3893 gnd.n3892 163.367
R6930 gnd.n3892 gnd.n3891 163.367
R6931 gnd.n3891 gnd.n2088 163.367
R6932 gnd.n3315 gnd.n2088 163.367
R6933 gnd.n3881 gnd.n3315 163.367
R6934 gnd.n3881 gnd.n3316 163.367
R6935 gnd.n3877 gnd.n3316 163.367
R6936 gnd.n3877 gnd.n3876 163.367
R6937 gnd.n3876 gnd.n3320 163.367
R6938 gnd.n3328 gnd.n3320 163.367
R6939 gnd.n3866 gnd.n3328 163.367
R6940 gnd.n3866 gnd.n3329 163.367
R6941 gnd.n3862 gnd.n3329 163.367
R6942 gnd.n3862 gnd.n3861 163.367
R6943 gnd.n3861 gnd.n3333 163.367
R6944 gnd.n3344 gnd.n3333 163.367
R6945 gnd.n3344 gnd.n3341 163.367
R6946 gnd.n3850 gnd.n3341 163.367
R6947 gnd.n3850 gnd.n3342 163.367
R6948 gnd.n3846 gnd.n3342 163.367
R6949 gnd.n3846 gnd.n3348 163.367
R6950 gnd.n3356 gnd.n3348 163.367
R6951 gnd.n3837 gnd.n3356 163.367
R6952 gnd.n3837 gnd.n3357 163.367
R6953 gnd.n3833 gnd.n3357 163.367
R6954 gnd.n3833 gnd.n3832 163.367
R6955 gnd.n3832 gnd.n3360 163.367
R6956 gnd.n3369 gnd.n3360 163.367
R6957 gnd.n3823 gnd.n3369 163.367
R6958 gnd.n3823 gnd.n3370 163.367
R6959 gnd.n3819 gnd.n3370 163.367
R6960 gnd.n3819 gnd.n3818 163.367
R6961 gnd.n3818 gnd.n3374 163.367
R6962 gnd.n3383 gnd.n3374 163.367
R6963 gnd.n3809 gnd.n3383 163.367
R6964 gnd.n3809 gnd.n3384 163.367
R6965 gnd.n3805 gnd.n3384 163.367
R6966 gnd.n3805 gnd.n3804 163.367
R6967 gnd.n3804 gnd.n3388 163.367
R6968 gnd.n3397 gnd.n3388 163.367
R6969 gnd.n3795 gnd.n3397 163.367
R6970 gnd.n3795 gnd.n3398 163.367
R6971 gnd.n3791 gnd.n3398 163.367
R6972 gnd.n3791 gnd.n3790 163.367
R6973 gnd.n3790 gnd.n3402 163.367
R6974 gnd.n3410 gnd.n3402 163.367
R6975 gnd.n3780 gnd.n3410 163.367
R6976 gnd.n3780 gnd.n1958 163.367
R6977 gnd.n3776 gnd.n1958 163.367
R6978 gnd.n3776 gnd.n3775 163.367
R6979 gnd.n3775 gnd.n3414 163.367
R6980 gnd.n3422 gnd.n3414 163.367
R6981 gnd.n3765 gnd.n3422 163.367
R6982 gnd.n3765 gnd.n3423 163.367
R6983 gnd.n3761 gnd.n3423 163.367
R6984 gnd.n3761 gnd.n3427 163.367
R6985 gnd.n3437 gnd.n3427 163.367
R6986 gnd.n3437 gnd.n3435 163.367
R6987 gnd.n3750 gnd.n3435 163.367
R6988 gnd.n3750 gnd.n3436 163.367
R6989 gnd.n3746 gnd.n3436 163.367
R6990 gnd.n3746 gnd.n3441 163.367
R6991 gnd.n3450 gnd.n3441 163.367
R6992 gnd.n3736 gnd.n3450 163.367
R6993 gnd.n3736 gnd.n3451 163.367
R6994 gnd.n3732 gnd.n3451 163.367
R6995 gnd.n3732 gnd.n3454 163.367
R6996 gnd.n3464 gnd.n3454 163.367
R6997 gnd.n3464 gnd.n3462 163.367
R6998 gnd.n3721 gnd.n3462 163.367
R6999 gnd.n3721 gnd.n3463 163.367
R7000 gnd.n3717 gnd.n3463 163.367
R7001 gnd.n3717 gnd.n3468 163.367
R7002 gnd.n3480 gnd.n3468 163.367
R7003 gnd.n3480 gnd.n3478 163.367
R7004 gnd.n3707 gnd.n3478 163.367
R7005 gnd.n3707 gnd.n3479 163.367
R7006 gnd.n3703 gnd.n3479 163.367
R7007 gnd.n3703 gnd.n3484 163.367
R7008 gnd.n3695 gnd.n3484 163.367
R7009 gnd.n3695 gnd.n3491 163.367
R7010 gnd.n3691 gnd.n3491 163.367
R7011 gnd.n3691 gnd.n3493 163.367
R7012 gnd.n3006 gnd.n3005 163.367
R7013 gnd.n3005 gnd.n2929 163.367
R7014 gnd.n3001 gnd.n2999 163.367
R7015 gnd.n2997 gnd.n2931 163.367
R7016 gnd.n2993 gnd.n2991 163.367
R7017 gnd.n2989 gnd.n2933 163.367
R7018 gnd.n2985 gnd.n2983 163.367
R7019 gnd.n2981 gnd.n2935 163.367
R7020 gnd.n2977 gnd.n2975 163.367
R7021 gnd.n2973 gnd.n2937 163.367
R7022 gnd.n2969 gnd.n2967 163.367
R7023 gnd.n2965 gnd.n2939 163.367
R7024 gnd.n2961 gnd.n2959 163.367
R7025 gnd.n2957 gnd.n2941 163.367
R7026 gnd.n2953 gnd.n2951 163.367
R7027 gnd.n2948 gnd.n2947 163.367
R7028 gnd.n3112 gnd.n3110 163.367
R7029 gnd.n3108 gnd.n2883 163.367
R7030 gnd.n3103 gnd.n3101 163.367
R7031 gnd.n3099 gnd.n2887 163.367
R7032 gnd.n3095 gnd.n3093 163.367
R7033 gnd.n3091 gnd.n2889 163.367
R7034 gnd.n3087 gnd.n3085 163.367
R7035 gnd.n3083 gnd.n2891 163.367
R7036 gnd.n3079 gnd.n3077 163.367
R7037 gnd.n3075 gnd.n2893 163.367
R7038 gnd.n3071 gnd.n3069 163.367
R7039 gnd.n3067 gnd.n2895 163.367
R7040 gnd.n3063 gnd.n3061 163.367
R7041 gnd.n3059 gnd.n2897 163.367
R7042 gnd.n3055 gnd.n3053 163.367
R7043 gnd.n3051 gnd.n2899 163.367
R7044 gnd.n3042 gnd.n2905 163.367
R7045 gnd.n3042 gnd.n2907 163.367
R7046 gnd.n3038 gnd.n2907 163.367
R7047 gnd.n3038 gnd.n3037 163.367
R7048 gnd.n3037 gnd.n3013 163.367
R7049 gnd.n3023 gnd.n3013 163.367
R7050 gnd.n3027 gnd.n3023 163.367
R7051 gnd.n3027 gnd.n2094 163.367
R7052 gnd.n3303 gnd.n2094 163.367
R7053 gnd.n3303 gnd.n2082 163.367
R7054 gnd.n3309 gnd.n2082 163.367
R7055 gnd.n3310 gnd.n3309 163.367
R7056 gnd.n3310 gnd.n2091 163.367
R7057 gnd.n3889 gnd.n2091 163.367
R7058 gnd.n3889 gnd.n2092 163.367
R7059 gnd.n3885 gnd.n2092 163.367
R7060 gnd.n3885 gnd.n3884 163.367
R7061 gnd.n3884 gnd.n3314 163.367
R7062 gnd.n3322 gnd.n3314 163.367
R7063 gnd.n3874 gnd.n3322 163.367
R7064 gnd.n3874 gnd.n3323 163.367
R7065 gnd.n3870 gnd.n3323 163.367
R7066 gnd.n3870 gnd.n3869 163.367
R7067 gnd.n3869 gnd.n3327 163.367
R7068 gnd.n3335 gnd.n3327 163.367
R7069 gnd.n3859 gnd.n3335 163.367
R7070 gnd.n3859 gnd.n3336 163.367
R7071 gnd.n3855 gnd.n3336 163.367
R7072 gnd.n3855 gnd.n3854 163.367
R7073 gnd.n3854 gnd.n3340 163.367
R7074 gnd.n3350 gnd.n3340 163.367
R7075 gnd.n3844 gnd.n3350 163.367
R7076 gnd.n3844 gnd.n3351 163.367
R7077 gnd.n3840 gnd.n3351 163.367
R7078 gnd.n3840 gnd.n3839 163.367
R7079 gnd.n3839 gnd.n3355 163.367
R7080 gnd.n3362 gnd.n3355 163.367
R7081 gnd.n3830 gnd.n3362 163.367
R7082 gnd.n3830 gnd.n3363 163.367
R7083 gnd.n3826 gnd.n3363 163.367
R7084 gnd.n3826 gnd.n3825 163.367
R7085 gnd.n3825 gnd.n3367 163.367
R7086 gnd.n3376 gnd.n3367 163.367
R7087 gnd.n3816 gnd.n3376 163.367
R7088 gnd.n3816 gnd.n3377 163.367
R7089 gnd.n3812 gnd.n3377 163.367
R7090 gnd.n3812 gnd.n3811 163.367
R7091 gnd.n3811 gnd.n3381 163.367
R7092 gnd.n3390 gnd.n3381 163.367
R7093 gnd.n3802 gnd.n3390 163.367
R7094 gnd.n3802 gnd.n3391 163.367
R7095 gnd.n3798 gnd.n3391 163.367
R7096 gnd.n3798 gnd.n3797 163.367
R7097 gnd.n3797 gnd.n3395 163.367
R7098 gnd.n3404 gnd.n3395 163.367
R7099 gnd.n3788 gnd.n3404 163.367
R7100 gnd.n3788 gnd.n3405 163.367
R7101 gnd.n3784 gnd.n3405 163.367
R7102 gnd.n3784 gnd.n3409 163.367
R7103 gnd.n3409 gnd.n1955 163.367
R7104 gnd.n3416 gnd.n1955 163.367
R7105 gnd.n3773 gnd.n3416 163.367
R7106 gnd.n3773 gnd.n3417 163.367
R7107 gnd.n3769 gnd.n3417 163.367
R7108 gnd.n3769 gnd.n3421 163.367
R7109 gnd.n3429 gnd.n3421 163.367
R7110 gnd.n3759 gnd.n3429 163.367
R7111 gnd.n3759 gnd.n3431 163.367
R7112 gnd.n3755 gnd.n3431 163.367
R7113 gnd.n3755 gnd.n3754 163.367
R7114 gnd.n3754 gnd.n3434 163.367
R7115 gnd.n3444 gnd.n3434 163.367
R7116 gnd.n3744 gnd.n3444 163.367
R7117 gnd.n3744 gnd.n3445 163.367
R7118 gnd.n3740 gnd.n3445 163.367
R7119 gnd.n3740 gnd.n3449 163.367
R7120 gnd.n3455 gnd.n3449 163.367
R7121 gnd.n3730 gnd.n3455 163.367
R7122 gnd.n3730 gnd.n3458 163.367
R7123 gnd.n3726 gnd.n3458 163.367
R7124 gnd.n3726 gnd.n3725 163.367
R7125 gnd.n3725 gnd.n3461 163.367
R7126 gnd.n3469 gnd.n3461 163.367
R7127 gnd.n3715 gnd.n3469 163.367
R7128 gnd.n3715 gnd.n3471 163.367
R7129 gnd.n3711 gnd.n3471 163.367
R7130 gnd.n3711 gnd.n3710 163.367
R7131 gnd.n3710 gnd.n3709 163.367
R7132 gnd.n3709 gnd.n3475 163.367
R7133 gnd.n3701 gnd.n3475 163.367
R7134 gnd.n3701 gnd.n3485 163.367
R7135 gnd.n3697 gnd.n3485 163.367
R7136 gnd.n3697 gnd.n3488 163.367
R7137 gnd.n3689 gnd.n3488 163.367
R7138 gnd.n3689 gnd.n3495 163.367
R7139 gnd.n3514 gnd.n3513 156.462
R7140 gnd.n6093 gnd.n6061 153.042
R7141 gnd.n6157 gnd.n6156 152.079
R7142 gnd.n6125 gnd.n6124 152.079
R7143 gnd.n6093 gnd.n6092 152.079
R7144 gnd.n2920 gnd.n2919 152
R7145 gnd.n2921 gnd.n2910 152
R7146 gnd.n2923 gnd.n2922 152
R7147 gnd.n2925 gnd.n2908 152
R7148 gnd.n2927 gnd.n2926 152
R7149 gnd.n3512 gnd.n3496 152
R7150 gnd.n3504 gnd.n3497 152
R7151 gnd.n3503 gnd.n3502 152
R7152 gnd.n3501 gnd.n3498 152
R7153 gnd.n3499 gnd.t87 150.546
R7154 gnd.t3 gnd.n6135 147.661
R7155 gnd.t269 gnd.n6103 147.661
R7156 gnd.t1 gnd.n6071 147.661
R7157 gnd.t18 gnd.n6040 147.661
R7158 gnd.t20 gnd.n6008 147.661
R7159 gnd.t321 gnd.n5976 147.661
R7160 gnd.t218 gnd.n5944 147.661
R7161 gnd.t313 gnd.n5913 147.661
R7162 gnd.n3626 gnd.n3625 143.351
R7163 gnd.n2946 gnd.n2882 143.351
R7164 gnd.n3111 gnd.n2882 143.351
R7165 gnd.n4466 gnd.n1466 138.177
R7166 gnd.n3114 gnd.n3113 138.177
R7167 gnd.n2917 gnd.t128 130.484
R7168 gnd.n6960 gnd.n6959 127.278
R7169 gnd.n6961 gnd.n6960 127.278
R7170 gnd.n6961 gnd.n448 127.278
R7171 gnd.n6969 gnd.n448 127.278
R7172 gnd.n6970 gnd.n6969 127.278
R7173 gnd.n6971 gnd.n6970 127.278
R7174 gnd.n6971 gnd.n442 127.278
R7175 gnd.n6979 gnd.n442 127.278
R7176 gnd.n6980 gnd.n6979 127.278
R7177 gnd.n6981 gnd.n6980 127.278
R7178 gnd.n6981 gnd.n436 127.278
R7179 gnd.n6989 gnd.n436 127.278
R7180 gnd.n6990 gnd.n6989 127.278
R7181 gnd.n6991 gnd.n6990 127.278
R7182 gnd.n6991 gnd.n430 127.278
R7183 gnd.n6999 gnd.n430 127.278
R7184 gnd.n7000 gnd.n6999 127.278
R7185 gnd.n7001 gnd.n7000 127.278
R7186 gnd.n7001 gnd.n424 127.278
R7187 gnd.n7009 gnd.n424 127.278
R7188 gnd.n7010 gnd.n7009 127.278
R7189 gnd.n7011 gnd.n7010 127.278
R7190 gnd.n7011 gnd.n418 127.278
R7191 gnd.n7019 gnd.n418 127.278
R7192 gnd.n7020 gnd.n7019 127.278
R7193 gnd.n7021 gnd.n7020 127.278
R7194 gnd.n7021 gnd.n412 127.278
R7195 gnd.n7029 gnd.n412 127.278
R7196 gnd.n7030 gnd.n7029 127.278
R7197 gnd.n7031 gnd.n7030 127.278
R7198 gnd.n7031 gnd.n406 127.278
R7199 gnd.n7039 gnd.n406 127.278
R7200 gnd.n7040 gnd.n7039 127.278
R7201 gnd.n7041 gnd.n7040 127.278
R7202 gnd.n7041 gnd.n400 127.278
R7203 gnd.n7049 gnd.n400 127.278
R7204 gnd.n7050 gnd.n7049 127.278
R7205 gnd.n7051 gnd.n7050 127.278
R7206 gnd.n7051 gnd.n394 127.278
R7207 gnd.n7059 gnd.n394 127.278
R7208 gnd.n7060 gnd.n7059 127.278
R7209 gnd.n7061 gnd.n7060 127.278
R7210 gnd.n7061 gnd.n388 127.278
R7211 gnd.n7069 gnd.n388 127.278
R7212 gnd.n7070 gnd.n7069 127.278
R7213 gnd.n7071 gnd.n7070 127.278
R7214 gnd.n7071 gnd.n382 127.278
R7215 gnd.n7079 gnd.n382 127.278
R7216 gnd.n7080 gnd.n7079 127.278
R7217 gnd.n7081 gnd.n7080 127.278
R7218 gnd.n7081 gnd.n376 127.278
R7219 gnd.n7089 gnd.n376 127.278
R7220 gnd.n7090 gnd.n7089 127.278
R7221 gnd.n7091 gnd.n7090 127.278
R7222 gnd.n7091 gnd.n370 127.278
R7223 gnd.n7099 gnd.n370 127.278
R7224 gnd.n7100 gnd.n7099 127.278
R7225 gnd.n7101 gnd.n7100 127.278
R7226 gnd.n7101 gnd.n364 127.278
R7227 gnd.n7109 gnd.n364 127.278
R7228 gnd.n7110 gnd.n7109 127.278
R7229 gnd.n7111 gnd.n7110 127.278
R7230 gnd.n7111 gnd.n358 127.278
R7231 gnd.n7119 gnd.n358 127.278
R7232 gnd.n7120 gnd.n7119 127.278
R7233 gnd.n7121 gnd.n7120 127.278
R7234 gnd.n7121 gnd.n352 127.278
R7235 gnd.n7129 gnd.n352 127.278
R7236 gnd.n7130 gnd.n7129 127.278
R7237 gnd.n7131 gnd.n7130 127.278
R7238 gnd.n7131 gnd.n346 127.278
R7239 gnd.n7139 gnd.n346 127.278
R7240 gnd.n7140 gnd.n7139 127.278
R7241 gnd.n7141 gnd.n7140 127.278
R7242 gnd.n7141 gnd.n340 127.278
R7243 gnd.n7149 gnd.n340 127.278
R7244 gnd.n7150 gnd.n7149 127.278
R7245 gnd.n7151 gnd.n7150 127.278
R7246 gnd.n7151 gnd.n334 127.278
R7247 gnd.n7159 gnd.n334 127.278
R7248 gnd.n7160 gnd.n7159 127.278
R7249 gnd.n7162 gnd.n7160 127.278
R7250 gnd.n7162 gnd.n7161 127.278
R7251 gnd.n2926 gnd.t143 126.766
R7252 gnd.n2924 gnd.t98 126.766
R7253 gnd.n2910 gnd.t134 126.766
R7254 gnd.n2918 gnd.t118 126.766
R7255 gnd.n3500 gnd.t60 126.766
R7256 gnd.n3502 gnd.t162 126.766
R7257 gnd.n3511 gnd.t121 126.766
R7258 gnd.n3513 gnd.t111 126.766
R7259 gnd.n6152 gnd.n6151 104.615
R7260 gnd.n6151 gnd.n6129 104.615
R7261 gnd.n6144 gnd.n6129 104.615
R7262 gnd.n6144 gnd.n6143 104.615
R7263 gnd.n6143 gnd.n6133 104.615
R7264 gnd.n6136 gnd.n6133 104.615
R7265 gnd.n6120 gnd.n6119 104.615
R7266 gnd.n6119 gnd.n6097 104.615
R7267 gnd.n6112 gnd.n6097 104.615
R7268 gnd.n6112 gnd.n6111 104.615
R7269 gnd.n6111 gnd.n6101 104.615
R7270 gnd.n6104 gnd.n6101 104.615
R7271 gnd.n6088 gnd.n6087 104.615
R7272 gnd.n6087 gnd.n6065 104.615
R7273 gnd.n6080 gnd.n6065 104.615
R7274 gnd.n6080 gnd.n6079 104.615
R7275 gnd.n6079 gnd.n6069 104.615
R7276 gnd.n6072 gnd.n6069 104.615
R7277 gnd.n6057 gnd.n6056 104.615
R7278 gnd.n6056 gnd.n6034 104.615
R7279 gnd.n6049 gnd.n6034 104.615
R7280 gnd.n6049 gnd.n6048 104.615
R7281 gnd.n6048 gnd.n6038 104.615
R7282 gnd.n6041 gnd.n6038 104.615
R7283 gnd.n6025 gnd.n6024 104.615
R7284 gnd.n6024 gnd.n6002 104.615
R7285 gnd.n6017 gnd.n6002 104.615
R7286 gnd.n6017 gnd.n6016 104.615
R7287 gnd.n6016 gnd.n6006 104.615
R7288 gnd.n6009 gnd.n6006 104.615
R7289 gnd.n5993 gnd.n5992 104.615
R7290 gnd.n5992 gnd.n5970 104.615
R7291 gnd.n5985 gnd.n5970 104.615
R7292 gnd.n5985 gnd.n5984 104.615
R7293 gnd.n5984 gnd.n5974 104.615
R7294 gnd.n5977 gnd.n5974 104.615
R7295 gnd.n5961 gnd.n5960 104.615
R7296 gnd.n5960 gnd.n5938 104.615
R7297 gnd.n5953 gnd.n5938 104.615
R7298 gnd.n5953 gnd.n5952 104.615
R7299 gnd.n5952 gnd.n5942 104.615
R7300 gnd.n5945 gnd.n5942 104.615
R7301 gnd.n5930 gnd.n5929 104.615
R7302 gnd.n5929 gnd.n5907 104.615
R7303 gnd.n5922 gnd.n5907 104.615
R7304 gnd.n5922 gnd.n5921 104.615
R7305 gnd.n5921 gnd.n5911 104.615
R7306 gnd.n5914 gnd.n5911 104.615
R7307 gnd.n5285 gnd.t149 100.632
R7308 gnd.n4936 gnd.t81 100.632
R7309 gnd.n7526 gnd.n116 99.6594
R7310 gnd.n7524 gnd.n7523 99.6594
R7311 gnd.n7519 gnd.n123 99.6594
R7312 gnd.n7517 gnd.n7516 99.6594
R7313 gnd.n7512 gnd.n130 99.6594
R7314 gnd.n7510 gnd.n7509 99.6594
R7315 gnd.n7505 gnd.n137 99.6594
R7316 gnd.n7503 gnd.n7502 99.6594
R7317 gnd.n7495 gnd.n144 99.6594
R7318 gnd.n7493 gnd.n7492 99.6594
R7319 gnd.n7488 gnd.n151 99.6594
R7320 gnd.n7486 gnd.n7485 99.6594
R7321 gnd.n7481 gnd.n158 99.6594
R7322 gnd.n7479 gnd.n7478 99.6594
R7323 gnd.n7474 gnd.n165 99.6594
R7324 gnd.n7472 gnd.n7471 99.6594
R7325 gnd.n7467 gnd.n172 99.6594
R7326 gnd.n7465 gnd.n7464 99.6594
R7327 gnd.n177 gnd.n176 99.6594
R7328 gnd.n4497 gnd.n4496 99.6594
R7329 gnd.n4491 gnd.n1418 99.6594
R7330 gnd.n4488 gnd.n1419 99.6594
R7331 gnd.n4484 gnd.n1420 99.6594
R7332 gnd.n4480 gnd.n1421 99.6594
R7333 gnd.n4476 gnd.n1422 99.6594
R7334 gnd.n4472 gnd.n1423 99.6594
R7335 gnd.n4468 gnd.n1424 99.6594
R7336 gnd.n4463 gnd.n1426 99.6594
R7337 gnd.n4459 gnd.n1427 99.6594
R7338 gnd.n4455 gnd.n1428 99.6594
R7339 gnd.n4451 gnd.n1429 99.6594
R7340 gnd.n4447 gnd.n1430 99.6594
R7341 gnd.n4443 gnd.n1431 99.6594
R7342 gnd.n4439 gnd.n1432 99.6594
R7343 gnd.n4435 gnd.n1433 99.6594
R7344 gnd.n4431 gnd.n1434 99.6594
R7345 gnd.n1490 gnd.n1435 99.6594
R7346 gnd.n3142 gnd.n3141 99.6594
R7347 gnd.n3137 gnd.n2283 99.6594
R7348 gnd.n3133 gnd.n2282 99.6594
R7349 gnd.n3129 gnd.n2281 99.6594
R7350 gnd.n3125 gnd.n2280 99.6594
R7351 gnd.n3121 gnd.n2279 99.6594
R7352 gnd.n3117 gnd.n2278 99.6594
R7353 gnd.n2874 gnd.n2276 99.6594
R7354 gnd.n2872 gnd.n2275 99.6594
R7355 gnd.n2868 gnd.n2274 99.6594
R7356 gnd.n2864 gnd.n2273 99.6594
R7357 gnd.n2860 gnd.n2272 99.6594
R7358 gnd.n2856 gnd.n2271 99.6594
R7359 gnd.n2852 gnd.n2270 99.6594
R7360 gnd.n2848 gnd.n2269 99.6594
R7361 gnd.n2844 gnd.n2268 99.6594
R7362 gnd.n2840 gnd.n2267 99.6594
R7363 gnd.n2325 gnd.n2266 99.6594
R7364 gnd.n4904 gnd.n4903 99.6594
R7365 gnd.n4898 gnd.n933 99.6594
R7366 gnd.n4895 gnd.n934 99.6594
R7367 gnd.n4891 gnd.n935 99.6594
R7368 gnd.n4887 gnd.n936 99.6594
R7369 gnd.n4883 gnd.n937 99.6594
R7370 gnd.n4879 gnd.n938 99.6594
R7371 gnd.n4875 gnd.n939 99.6594
R7372 gnd.n4871 gnd.n940 99.6594
R7373 gnd.n4866 gnd.n941 99.6594
R7374 gnd.n4862 gnd.n942 99.6594
R7375 gnd.n4858 gnd.n943 99.6594
R7376 gnd.n4854 gnd.n944 99.6594
R7377 gnd.n4850 gnd.n945 99.6594
R7378 gnd.n4846 gnd.n946 99.6594
R7379 gnd.n4842 gnd.n947 99.6594
R7380 gnd.n4838 gnd.n948 99.6594
R7381 gnd.n4834 gnd.n949 99.6594
R7382 gnd.n1004 gnd.n950 99.6594
R7383 gnd.n6301 gnd.n4916 99.6594
R7384 gnd.n6299 gnd.n6298 99.6594
R7385 gnd.n6294 gnd.n4923 99.6594
R7386 gnd.n6292 gnd.n6291 99.6594
R7387 gnd.n6287 gnd.n4930 99.6594
R7388 gnd.n6285 gnd.n6284 99.6594
R7389 gnd.n6280 gnd.n4939 99.6594
R7390 gnd.n6278 gnd.n6277 99.6594
R7391 gnd.n5583 gnd.n5228 99.6594
R7392 gnd.n5254 gnd.n5235 99.6594
R7393 gnd.n5256 gnd.n5236 99.6594
R7394 gnd.n5264 gnd.n5237 99.6594
R7395 gnd.n5266 gnd.n5238 99.6594
R7396 gnd.n5274 gnd.n5239 99.6594
R7397 gnd.n5276 gnd.n5240 99.6594
R7398 gnd.n5284 gnd.n5241 99.6594
R7399 gnd.n6269 gnd.n4946 99.6594
R7400 gnd.n6267 gnd.n6266 99.6594
R7401 gnd.n6262 gnd.n4953 99.6594
R7402 gnd.n6260 gnd.n6259 99.6594
R7403 gnd.n6255 gnd.n4960 99.6594
R7404 gnd.n6253 gnd.n6252 99.6594
R7405 gnd.n6248 gnd.n4967 99.6594
R7406 gnd.n6246 gnd.n6245 99.6594
R7407 gnd.n6241 gnd.n4974 99.6594
R7408 gnd.n6239 gnd.n6238 99.6594
R7409 gnd.n6234 gnd.n4983 99.6594
R7410 gnd.n6232 gnd.n6231 99.6594
R7411 gnd.n6227 gnd.n6226 99.6594
R7412 gnd.n5412 gnd.n5411 99.6594
R7413 gnd.n5406 gnd.n5323 99.6594
R7414 gnd.n5403 gnd.n5324 99.6594
R7415 gnd.n5399 gnd.n5325 99.6594
R7416 gnd.n5395 gnd.n5326 99.6594
R7417 gnd.n5391 gnd.n5327 99.6594
R7418 gnd.n5387 gnd.n5328 99.6594
R7419 gnd.n5383 gnd.n5329 99.6594
R7420 gnd.n5379 gnd.n5330 99.6594
R7421 gnd.n5375 gnd.n5331 99.6594
R7422 gnd.n5371 gnd.n5332 99.6594
R7423 gnd.n5367 gnd.n5333 99.6594
R7424 gnd.n5414 gnd.n5322 99.6594
R7425 gnd.n7374 gnd.n7373 99.6594
R7426 gnd.n7379 gnd.n7378 99.6594
R7427 gnd.n7382 gnd.n7381 99.6594
R7428 gnd.n7387 gnd.n7386 99.6594
R7429 gnd.n7390 gnd.n7389 99.6594
R7430 gnd.n7395 gnd.n7394 99.6594
R7431 gnd.n7398 gnd.n7397 99.6594
R7432 gnd.n7403 gnd.n7402 99.6594
R7433 gnd.n7406 gnd.n103 99.6594
R7434 gnd.n1500 gnd.n1436 99.6594
R7435 gnd.n1728 gnd.n1437 99.6594
R7436 gnd.n1730 gnd.n1438 99.6594
R7437 gnd.n1747 gnd.n1439 99.6594
R7438 gnd.n1749 gnd.n1440 99.6594
R7439 gnd.n1766 gnd.n1441 99.6594
R7440 gnd.n1768 gnd.n1442 99.6594
R7441 gnd.n1784 gnd.n1443 99.6594
R7442 gnd.n1695 gnd.n1444 99.6594
R7443 gnd.n2253 gnd.n2252 99.6594
R7444 gnd.n2254 gnd.n2202 99.6594
R7445 gnd.n2256 gnd.n2210 99.6594
R7446 gnd.n2258 gnd.n2257 99.6594
R7447 gnd.n2259 gnd.n2219 99.6594
R7448 gnd.n2261 gnd.n2228 99.6594
R7449 gnd.n2263 gnd.n2262 99.6594
R7450 gnd.n2264 gnd.n2237 99.6594
R7451 gnd.n3145 gnd.n3144 99.6594
R7452 gnd.n2533 gnd.n951 99.6594
R7453 gnd.n2530 gnd.n952 99.6594
R7454 gnd.n2526 gnd.n953 99.6594
R7455 gnd.n2522 gnd.n954 99.6594
R7456 gnd.n2518 gnd.n955 99.6594
R7457 gnd.n2514 gnd.n956 99.6594
R7458 gnd.n2510 gnd.n957 99.6594
R7459 gnd.n2506 gnd.n958 99.6594
R7460 gnd.n2502 gnd.n959 99.6594
R7461 gnd.n2531 gnd.n951 99.6594
R7462 gnd.n2527 gnd.n952 99.6594
R7463 gnd.n2523 gnd.n953 99.6594
R7464 gnd.n2519 gnd.n954 99.6594
R7465 gnd.n2515 gnd.n955 99.6594
R7466 gnd.n2511 gnd.n956 99.6594
R7467 gnd.n2507 gnd.n957 99.6594
R7468 gnd.n2503 gnd.n958 99.6594
R7469 gnd.n2491 gnd.n959 99.6594
R7470 gnd.n3144 gnd.n2248 99.6594
R7471 gnd.n2264 gnd.n2236 99.6594
R7472 gnd.n2263 gnd.n2229 99.6594
R7473 gnd.n2261 gnd.n2260 99.6594
R7474 gnd.n2259 gnd.n2218 99.6594
R7475 gnd.n2258 gnd.n2211 99.6594
R7476 gnd.n2256 gnd.n2255 99.6594
R7477 gnd.n2254 gnd.n2201 99.6594
R7478 gnd.n2253 gnd.n2251 99.6594
R7479 gnd.n1727 gnd.n1436 99.6594
R7480 gnd.n1731 gnd.n1437 99.6594
R7481 gnd.n1746 gnd.n1438 99.6594
R7482 gnd.n1750 gnd.n1439 99.6594
R7483 gnd.n1765 gnd.n1440 99.6594
R7484 gnd.n1769 gnd.n1441 99.6594
R7485 gnd.n1783 gnd.n1442 99.6594
R7486 gnd.n1694 gnd.n1443 99.6594
R7487 gnd.n1690 gnd.n1444 99.6594
R7488 gnd.n7407 gnd.n7406 99.6594
R7489 gnd.n7402 gnd.n7401 99.6594
R7490 gnd.n7397 gnd.n7396 99.6594
R7491 gnd.n7394 gnd.n7393 99.6594
R7492 gnd.n7389 gnd.n7388 99.6594
R7493 gnd.n7386 gnd.n7385 99.6594
R7494 gnd.n7381 gnd.n7380 99.6594
R7495 gnd.n7378 gnd.n7377 99.6594
R7496 gnd.n7373 gnd.n7372 99.6594
R7497 gnd.n5412 gnd.n5335 99.6594
R7498 gnd.n5404 gnd.n5323 99.6594
R7499 gnd.n5400 gnd.n5324 99.6594
R7500 gnd.n5396 gnd.n5325 99.6594
R7501 gnd.n5392 gnd.n5326 99.6594
R7502 gnd.n5388 gnd.n5327 99.6594
R7503 gnd.n5384 gnd.n5328 99.6594
R7504 gnd.n5380 gnd.n5329 99.6594
R7505 gnd.n5376 gnd.n5330 99.6594
R7506 gnd.n5372 gnd.n5331 99.6594
R7507 gnd.n5368 gnd.n5332 99.6594
R7508 gnd.n5364 gnd.n5333 99.6594
R7509 gnd.n5415 gnd.n5414 99.6594
R7510 gnd.n6226 gnd.n4985 99.6594
R7511 gnd.n6233 gnd.n6232 99.6594
R7512 gnd.n4983 gnd.n4975 99.6594
R7513 gnd.n6240 gnd.n6239 99.6594
R7514 gnd.n4974 gnd.n4968 99.6594
R7515 gnd.n6247 gnd.n6246 99.6594
R7516 gnd.n4967 gnd.n4961 99.6594
R7517 gnd.n6254 gnd.n6253 99.6594
R7518 gnd.n4960 gnd.n4954 99.6594
R7519 gnd.n6261 gnd.n6260 99.6594
R7520 gnd.n4953 gnd.n4947 99.6594
R7521 gnd.n6268 gnd.n6267 99.6594
R7522 gnd.n4946 gnd.n4943 99.6594
R7523 gnd.n5584 gnd.n5583 99.6594
R7524 gnd.n5257 gnd.n5235 99.6594
R7525 gnd.n5263 gnd.n5236 99.6594
R7526 gnd.n5267 gnd.n5237 99.6594
R7527 gnd.n5273 gnd.n5238 99.6594
R7528 gnd.n5277 gnd.n5239 99.6594
R7529 gnd.n5283 gnd.n5240 99.6594
R7530 gnd.n5241 gnd.n5225 99.6594
R7531 gnd.n6279 gnd.n6278 99.6594
R7532 gnd.n4939 gnd.n4931 99.6594
R7533 gnd.n6286 gnd.n6285 99.6594
R7534 gnd.n4930 gnd.n4924 99.6594
R7535 gnd.n6293 gnd.n6292 99.6594
R7536 gnd.n4923 gnd.n4917 99.6594
R7537 gnd.n6300 gnd.n6299 99.6594
R7538 gnd.n4916 gnd.n4913 99.6594
R7539 gnd.n4904 gnd.n963 99.6594
R7540 gnd.n4896 gnd.n933 99.6594
R7541 gnd.n4892 gnd.n934 99.6594
R7542 gnd.n4888 gnd.n935 99.6594
R7543 gnd.n4884 gnd.n936 99.6594
R7544 gnd.n4880 gnd.n937 99.6594
R7545 gnd.n4876 gnd.n938 99.6594
R7546 gnd.n4872 gnd.n939 99.6594
R7547 gnd.n4867 gnd.n940 99.6594
R7548 gnd.n4863 gnd.n941 99.6594
R7549 gnd.n4859 gnd.n942 99.6594
R7550 gnd.n4855 gnd.n943 99.6594
R7551 gnd.n4851 gnd.n944 99.6594
R7552 gnd.n4847 gnd.n945 99.6594
R7553 gnd.n4843 gnd.n946 99.6594
R7554 gnd.n4839 gnd.n947 99.6594
R7555 gnd.n4835 gnd.n948 99.6594
R7556 gnd.n1003 gnd.n949 99.6594
R7557 gnd.n4827 gnd.n950 99.6594
R7558 gnd.n2839 gnd.n2266 99.6594
R7559 gnd.n2843 gnd.n2267 99.6594
R7560 gnd.n2847 gnd.n2268 99.6594
R7561 gnd.n2851 gnd.n2269 99.6594
R7562 gnd.n2855 gnd.n2270 99.6594
R7563 gnd.n2859 gnd.n2271 99.6594
R7564 gnd.n2863 gnd.n2272 99.6594
R7565 gnd.n2867 gnd.n2273 99.6594
R7566 gnd.n2871 gnd.n2274 99.6594
R7567 gnd.n2875 gnd.n2275 99.6594
R7568 gnd.n3116 gnd.n2277 99.6594
R7569 gnd.n3120 gnd.n2278 99.6594
R7570 gnd.n3124 gnd.n2279 99.6594
R7571 gnd.n3128 gnd.n2280 99.6594
R7572 gnd.n3132 gnd.n2281 99.6594
R7573 gnd.n3136 gnd.n2282 99.6594
R7574 gnd.n2285 gnd.n2283 99.6594
R7575 gnd.n3142 gnd.n2284 99.6594
R7576 gnd.n4497 gnd.n1448 99.6594
R7577 gnd.n4489 gnd.n1418 99.6594
R7578 gnd.n4485 gnd.n1419 99.6594
R7579 gnd.n4481 gnd.n1420 99.6594
R7580 gnd.n4477 gnd.n1421 99.6594
R7581 gnd.n4473 gnd.n1422 99.6594
R7582 gnd.n4469 gnd.n1423 99.6594
R7583 gnd.n4464 gnd.n1425 99.6594
R7584 gnd.n4460 gnd.n1426 99.6594
R7585 gnd.n4456 gnd.n1427 99.6594
R7586 gnd.n4452 gnd.n1428 99.6594
R7587 gnd.n4448 gnd.n1429 99.6594
R7588 gnd.n4444 gnd.n1430 99.6594
R7589 gnd.n4440 gnd.n1431 99.6594
R7590 gnd.n4436 gnd.n1432 99.6594
R7591 gnd.n4432 gnd.n1433 99.6594
R7592 gnd.n1489 gnd.n1434 99.6594
R7593 gnd.n4424 gnd.n1435 99.6594
R7594 gnd.n176 gnd.n173 99.6594
R7595 gnd.n7466 gnd.n7465 99.6594
R7596 gnd.n172 gnd.n166 99.6594
R7597 gnd.n7473 gnd.n7472 99.6594
R7598 gnd.n165 gnd.n159 99.6594
R7599 gnd.n7480 gnd.n7479 99.6594
R7600 gnd.n158 gnd.n152 99.6594
R7601 gnd.n7487 gnd.n7486 99.6594
R7602 gnd.n151 gnd.n145 99.6594
R7603 gnd.n7494 gnd.n7493 99.6594
R7604 gnd.n144 gnd.n138 99.6594
R7605 gnd.n7504 gnd.n7503 99.6594
R7606 gnd.n137 gnd.n131 99.6594
R7607 gnd.n7511 gnd.n7510 99.6594
R7608 gnd.n130 gnd.n124 99.6594
R7609 gnd.n7518 gnd.n7517 99.6594
R7610 gnd.n123 gnd.n117 99.6594
R7611 gnd.n7525 gnd.n7524 99.6594
R7612 gnd.n116 gnd.n113 99.6594
R7613 gnd.n3192 gnd.n3191 99.6594
R7614 gnd.n2205 gnd.n2182 99.6594
R7615 gnd.n2207 gnd.n2183 99.6594
R7616 gnd.n2215 gnd.n2184 99.6594
R7617 gnd.n2223 gnd.n2185 99.6594
R7618 gnd.n2225 gnd.n2186 99.6594
R7619 gnd.n2233 gnd.n2187 99.6594
R7620 gnd.n2243 gnd.n2188 99.6594
R7621 gnd.n2245 gnd.n2189 99.6594
R7622 gnd.n2800 gnd.n2190 99.6594
R7623 gnd.n2802 gnd.n2191 99.6594
R7624 gnd.n2806 gnd.n2192 99.6594
R7625 gnd.n2812 gnd.n2193 99.6594
R7626 gnd.n3195 gnd.n3194 99.6594
R7627 gnd.n3192 gnd.n2195 99.6594
R7628 gnd.n2206 gnd.n2182 99.6594
R7629 gnd.n2214 gnd.n2183 99.6594
R7630 gnd.n2222 gnd.n2184 99.6594
R7631 gnd.n2224 gnd.n2185 99.6594
R7632 gnd.n2232 gnd.n2186 99.6594
R7633 gnd.n2242 gnd.n2187 99.6594
R7634 gnd.n2244 gnd.n2188 99.6594
R7635 gnd.n2799 gnd.n2189 99.6594
R7636 gnd.n2801 gnd.n2190 99.6594
R7637 gnd.n2805 gnd.n2191 99.6594
R7638 gnd.n2807 gnd.n2192 99.6594
R7639 gnd.n2193 gnd.n2180 99.6594
R7640 gnd.n3194 gnd.n2177 99.6594
R7641 gnd.n1736 gnd.n1718 99.6594
R7642 gnd.n1740 gnd.n1738 99.6594
R7643 gnd.n1755 gnd.n1711 99.6594
R7644 gnd.n1759 gnd.n1757 99.6594
R7645 gnd.n1774 gnd.n1704 99.6594
R7646 gnd.n1778 gnd.n1776 99.6594
R7647 gnd.n1790 gnd.n1698 99.6594
R7648 gnd.n1794 gnd.n1792 99.6594
R7649 gnd.n1804 gnd.n1686 99.6594
R7650 gnd.n1807 gnd.n1806 99.6594
R7651 gnd.n1810 gnd.n1809 99.6594
R7652 gnd.n1815 gnd.n1814 99.6594
R7653 gnd.n1818 gnd.n1817 99.6594
R7654 gnd.n4208 gnd.n4207 99.6594
R7655 gnd.n4207 gnd.n4206 99.6594
R7656 gnd.n1817 gnd.n1816 99.6594
R7657 gnd.n1814 gnd.n1813 99.6594
R7658 gnd.n1809 gnd.n1808 99.6594
R7659 gnd.n1806 gnd.n1805 99.6594
R7660 gnd.n1793 gnd.n1686 99.6594
R7661 gnd.n1792 gnd.n1791 99.6594
R7662 gnd.n1777 gnd.n1698 99.6594
R7663 gnd.n1776 gnd.n1775 99.6594
R7664 gnd.n1758 gnd.n1704 99.6594
R7665 gnd.n1757 gnd.n1756 99.6594
R7666 gnd.n1739 gnd.n1711 99.6594
R7667 gnd.n1738 gnd.n1737 99.6594
R7668 gnd.n1718 gnd.n1405 99.6594
R7669 gnd.n2808 gnd.t117 98.63
R7670 gnd.n7404 gnd.t141 98.63
R7671 gnd.n1691 gnd.t133 98.63
R7672 gnd.n2238 gnd.t154 98.63
R7673 gnd.n1469 gnd.t103 98.63
R7674 gnd.n1491 gnd.t97 98.63
R7675 gnd.n179 gnd.t160 98.63
R7676 gnd.n7497 gnd.t85 98.63
R7677 gnd.n983 gnd.t66 98.63
R7678 gnd.n1005 gnd.t152 98.63
R7679 gnd.n2327 gnd.t157 98.63
R7680 gnd.n2305 gnd.t77 98.63
R7681 gnd.n2492 gnd.t106 98.63
R7682 gnd.n4216 gnd.t73 98.63
R7683 gnd.n2884 gnd.t127 92.8196
R7684 gnd.n3543 gnd.t138 92.8196
R7685 gnd.n2942 gnd.t167 92.8118
R7686 gnd.n3537 gnd.t92 92.8118
R7687 gnd.n2917 gnd.n2916 81.8399
R7688 gnd.n7161 gnd.n186 76.3673
R7689 gnd.n5286 gnd.t148 74.8376
R7690 gnd.n4937 gnd.t82 74.8376
R7691 gnd.n2885 gnd.t126 72.8438
R7692 gnd.n3544 gnd.t139 72.8438
R7693 gnd.n2918 gnd.n2911 72.8411
R7694 gnd.n2924 gnd.n2909 72.8411
R7695 gnd.n3511 gnd.n3510 72.8411
R7696 gnd.n2809 gnd.t116 72.836
R7697 gnd.n2943 gnd.t166 72.836
R7698 gnd.n3538 gnd.t93 72.836
R7699 gnd.n7405 gnd.t142 72.836
R7700 gnd.n1692 gnd.t132 72.836
R7701 gnd.n2239 gnd.t155 72.836
R7702 gnd.n1470 gnd.t102 72.836
R7703 gnd.n1492 gnd.t96 72.836
R7704 gnd.n180 gnd.t161 72.836
R7705 gnd.n7498 gnd.t86 72.836
R7706 gnd.n984 gnd.t65 72.836
R7707 gnd.n1006 gnd.t151 72.836
R7708 gnd.n2328 gnd.t158 72.836
R7709 gnd.n2306 gnd.t78 72.836
R7710 gnd.n2493 gnd.t105 72.836
R7711 gnd.n4217 gnd.t74 72.836
R7712 gnd.n3683 gnd.n3682 71.676
R7713 gnd.n3680 gnd.n3679 71.676
R7714 gnd.n3675 gnd.n3520 71.676
R7715 gnd.n3673 gnd.n3672 71.676
R7716 gnd.n3668 gnd.n3523 71.676
R7717 gnd.n3666 gnd.n3665 71.676
R7718 gnd.n3661 gnd.n3526 71.676
R7719 gnd.n3659 gnd.n3658 71.676
R7720 gnd.n3654 gnd.n3529 71.676
R7721 gnd.n3652 gnd.n3651 71.676
R7722 gnd.n3647 gnd.n3532 71.676
R7723 gnd.n3645 gnd.n3644 71.676
R7724 gnd.n3640 gnd.n3535 71.676
R7725 gnd.n3638 gnd.n3637 71.676
R7726 gnd.n3632 gnd.n3540 71.676
R7727 gnd.n3630 gnd.n3629 71.676
R7728 gnd.n3625 gnd.n3624 71.676
R7729 gnd.n3622 gnd.n3621 71.676
R7730 gnd.n3616 gnd.n3546 71.676
R7731 gnd.n3614 gnd.n3613 71.676
R7732 gnd.n3609 gnd.n3549 71.676
R7733 gnd.n3607 gnd.n3606 71.676
R7734 gnd.n3602 gnd.n3552 71.676
R7735 gnd.n3600 gnd.n3599 71.676
R7736 gnd.n3595 gnd.n3555 71.676
R7737 gnd.n3593 gnd.n3592 71.676
R7738 gnd.n3588 gnd.n3558 71.676
R7739 gnd.n3586 gnd.n3585 71.676
R7740 gnd.n3581 gnd.n3561 71.676
R7741 gnd.n3579 gnd.n3578 71.676
R7742 gnd.n3574 gnd.n3564 71.676
R7743 gnd.n3572 gnd.n3571 71.676
R7744 gnd.n3567 gnd.n3566 71.676
R7745 gnd.n3008 gnd.n3007 71.676
R7746 gnd.n3000 gnd.n2929 71.676
R7747 gnd.n2999 gnd.n2998 71.676
R7748 gnd.n2992 gnd.n2931 71.676
R7749 gnd.n2991 gnd.n2990 71.676
R7750 gnd.n2984 gnd.n2933 71.676
R7751 gnd.n2983 gnd.n2982 71.676
R7752 gnd.n2976 gnd.n2935 71.676
R7753 gnd.n2975 gnd.n2974 71.676
R7754 gnd.n2968 gnd.n2937 71.676
R7755 gnd.n2967 gnd.n2966 71.676
R7756 gnd.n2960 gnd.n2939 71.676
R7757 gnd.n2959 gnd.n2958 71.676
R7758 gnd.n2952 gnd.n2941 71.676
R7759 gnd.n2951 gnd.n2945 71.676
R7760 gnd.n2947 gnd.n2946 71.676
R7761 gnd.n3110 gnd.n3109 71.676
R7762 gnd.n3102 gnd.n2883 71.676
R7763 gnd.n3101 gnd.n3100 71.676
R7764 gnd.n3094 gnd.n2887 71.676
R7765 gnd.n3093 gnd.n3092 71.676
R7766 gnd.n3086 gnd.n2889 71.676
R7767 gnd.n3085 gnd.n3084 71.676
R7768 gnd.n3078 gnd.n2891 71.676
R7769 gnd.n3077 gnd.n3076 71.676
R7770 gnd.n3070 gnd.n2893 71.676
R7771 gnd.n3069 gnd.n3068 71.676
R7772 gnd.n3062 gnd.n2895 71.676
R7773 gnd.n3061 gnd.n3060 71.676
R7774 gnd.n3054 gnd.n2897 71.676
R7775 gnd.n3053 gnd.n3052 71.676
R7776 gnd.n3046 gnd.n2899 71.676
R7777 gnd.n3007 gnd.n3006 71.676
R7778 gnd.n3001 gnd.n3000 71.676
R7779 gnd.n2998 gnd.n2997 71.676
R7780 gnd.n2993 gnd.n2992 71.676
R7781 gnd.n2990 gnd.n2989 71.676
R7782 gnd.n2985 gnd.n2984 71.676
R7783 gnd.n2982 gnd.n2981 71.676
R7784 gnd.n2977 gnd.n2976 71.676
R7785 gnd.n2974 gnd.n2973 71.676
R7786 gnd.n2969 gnd.n2968 71.676
R7787 gnd.n2966 gnd.n2965 71.676
R7788 gnd.n2961 gnd.n2960 71.676
R7789 gnd.n2958 gnd.n2957 71.676
R7790 gnd.n2953 gnd.n2952 71.676
R7791 gnd.n2948 gnd.n2945 71.676
R7792 gnd.n3112 gnd.n3111 71.676
R7793 gnd.n3109 gnd.n3108 71.676
R7794 gnd.n3103 gnd.n3102 71.676
R7795 gnd.n3100 gnd.n3099 71.676
R7796 gnd.n3095 gnd.n3094 71.676
R7797 gnd.n3092 gnd.n3091 71.676
R7798 gnd.n3087 gnd.n3086 71.676
R7799 gnd.n3084 gnd.n3083 71.676
R7800 gnd.n3079 gnd.n3078 71.676
R7801 gnd.n3076 gnd.n3075 71.676
R7802 gnd.n3071 gnd.n3070 71.676
R7803 gnd.n3068 gnd.n3067 71.676
R7804 gnd.n3063 gnd.n3062 71.676
R7805 gnd.n3060 gnd.n3059 71.676
R7806 gnd.n3055 gnd.n3054 71.676
R7807 gnd.n3052 gnd.n3051 71.676
R7808 gnd.n3047 gnd.n3046 71.676
R7809 gnd.n3566 gnd.n3565 71.676
R7810 gnd.n3573 gnd.n3572 71.676
R7811 gnd.n3564 gnd.n3562 71.676
R7812 gnd.n3580 gnd.n3579 71.676
R7813 gnd.n3561 gnd.n3559 71.676
R7814 gnd.n3587 gnd.n3586 71.676
R7815 gnd.n3558 gnd.n3556 71.676
R7816 gnd.n3594 gnd.n3593 71.676
R7817 gnd.n3555 gnd.n3553 71.676
R7818 gnd.n3601 gnd.n3600 71.676
R7819 gnd.n3552 gnd.n3550 71.676
R7820 gnd.n3608 gnd.n3607 71.676
R7821 gnd.n3549 gnd.n3547 71.676
R7822 gnd.n3615 gnd.n3614 71.676
R7823 gnd.n3546 gnd.n3542 71.676
R7824 gnd.n3623 gnd.n3622 71.676
R7825 gnd.n3627 gnd.n3626 71.676
R7826 gnd.n3631 gnd.n3630 71.676
R7827 gnd.n3540 gnd.n3536 71.676
R7828 gnd.n3639 gnd.n3638 71.676
R7829 gnd.n3535 gnd.n3533 71.676
R7830 gnd.n3646 gnd.n3645 71.676
R7831 gnd.n3532 gnd.n3530 71.676
R7832 gnd.n3653 gnd.n3652 71.676
R7833 gnd.n3529 gnd.n3527 71.676
R7834 gnd.n3660 gnd.n3659 71.676
R7835 gnd.n3526 gnd.n3524 71.676
R7836 gnd.n3667 gnd.n3666 71.676
R7837 gnd.n3523 gnd.n3521 71.676
R7838 gnd.n3674 gnd.n3673 71.676
R7839 gnd.n3520 gnd.n3518 71.676
R7840 gnd.n3681 gnd.n3680 71.676
R7841 gnd.n3684 gnd.n3683 71.676
R7842 gnd.n10 gnd.t5 69.1507
R7843 gnd.n18 gnd.t284 68.4792
R7844 gnd.n17 gnd.t214 68.4792
R7845 gnd.n16 gnd.t240 68.4792
R7846 gnd.n15 gnd.t188 68.4792
R7847 gnd.n14 gnd.t247 68.4792
R7848 gnd.n13 gnd.t216 68.4792
R7849 gnd.n12 gnd.t306 68.4792
R7850 gnd.n11 gnd.t26 68.4792
R7851 gnd.n10 gnd.t249 68.4792
R7852 gnd.n5413 gnd.n5317 64.369
R7853 gnd.n3105 gnd.n2885 59.5399
R7854 gnd.n3618 gnd.n3544 59.5399
R7855 gnd.n2944 gnd.n2943 59.5399
R7856 gnd.n3634 gnd.n3538 59.5399
R7857 gnd.n3010 gnd.n2927 59.1804
R7858 gnd.n6309 gnd.n4906 57.3586
R7859 gnd.n4905 gnd.n961 57.3586
R7860 gnd.n7534 gnd.n106 57.3586
R7861 gnd.n5519 gnd.t288 56.607
R7862 gnd.n52 gnd.t195 56.607
R7863 gnd.n5488 gnd.t40 56.407
R7864 gnd.n5503 gnd.t238 56.407
R7865 gnd.n21 gnd.t316 56.407
R7866 gnd.n36 gnd.t43 56.407
R7867 gnd.n5532 gnd.t281 55.8337
R7868 gnd.n5501 gnd.t297 55.8337
R7869 gnd.n5516 gnd.t8 55.8337
R7870 gnd.n65 gnd.t259 55.8337
R7871 gnd.n34 gnd.t169 55.8337
R7872 gnd.n49 gnd.t276 55.8337
R7873 gnd.n2915 gnd.n2914 54.358
R7874 gnd.n3508 gnd.n3507 54.358
R7875 gnd.n5519 gnd.n5518 53.0052
R7876 gnd.n5521 gnd.n5520 53.0052
R7877 gnd.n5523 gnd.n5522 53.0052
R7878 gnd.n5525 gnd.n5524 53.0052
R7879 gnd.n5527 gnd.n5526 53.0052
R7880 gnd.n5529 gnd.n5528 53.0052
R7881 gnd.n5531 gnd.n5530 53.0052
R7882 gnd.n5488 gnd.n5487 53.0052
R7883 gnd.n5490 gnd.n5489 53.0052
R7884 gnd.n5492 gnd.n5491 53.0052
R7885 gnd.n5494 gnd.n5493 53.0052
R7886 gnd.n5496 gnd.n5495 53.0052
R7887 gnd.n5498 gnd.n5497 53.0052
R7888 gnd.n5500 gnd.n5499 53.0052
R7889 gnd.n5503 gnd.n5502 53.0052
R7890 gnd.n5505 gnd.n5504 53.0052
R7891 gnd.n5507 gnd.n5506 53.0052
R7892 gnd.n5509 gnd.n5508 53.0052
R7893 gnd.n5511 gnd.n5510 53.0052
R7894 gnd.n5513 gnd.n5512 53.0052
R7895 gnd.n5515 gnd.n5514 53.0052
R7896 gnd.n64 gnd.n63 53.0052
R7897 gnd.n62 gnd.n61 53.0052
R7898 gnd.n60 gnd.n59 53.0052
R7899 gnd.n58 gnd.n57 53.0052
R7900 gnd.n56 gnd.n55 53.0052
R7901 gnd.n54 gnd.n53 53.0052
R7902 gnd.n52 gnd.n51 53.0052
R7903 gnd.n33 gnd.n32 53.0052
R7904 gnd.n31 gnd.n30 53.0052
R7905 gnd.n29 gnd.n28 53.0052
R7906 gnd.n27 gnd.n26 53.0052
R7907 gnd.n25 gnd.n24 53.0052
R7908 gnd.n23 gnd.n22 53.0052
R7909 gnd.n21 gnd.n20 53.0052
R7910 gnd.n48 gnd.n47 53.0052
R7911 gnd.n46 gnd.n45 53.0052
R7912 gnd.n44 gnd.n43 53.0052
R7913 gnd.n42 gnd.n41 53.0052
R7914 gnd.n40 gnd.n39 53.0052
R7915 gnd.n38 gnd.n37 53.0052
R7916 gnd.n36 gnd.n35 53.0052
R7917 gnd.n3499 gnd.n3498 52.4801
R7918 gnd.n6136 gnd.t3 52.3082
R7919 gnd.n6104 gnd.t269 52.3082
R7920 gnd.n6072 gnd.t1 52.3082
R7921 gnd.n6041 gnd.t18 52.3082
R7922 gnd.n6009 gnd.t20 52.3082
R7923 gnd.n5977 gnd.t321 52.3082
R7924 gnd.n5945 gnd.t218 52.3082
R7925 gnd.n5914 gnd.t313 52.3082
R7926 gnd.n5966 gnd.n5934 51.4173
R7927 gnd.n6030 gnd.n6029 50.455
R7928 gnd.n5998 gnd.n5997 50.455
R7929 gnd.n5966 gnd.n5965 50.455
R7930 gnd.n5360 gnd.n5359 45.1884
R7931 gnd.n4981 gnd.n4980 45.1884
R7932 gnd.n3686 gnd.n3514 44.3322
R7933 gnd.n2918 gnd.n2917 44.3189
R7934 gnd.n2810 gnd.n2809 42.4732
R7935 gnd.n4218 gnd.n4217 42.4732
R7936 gnd.n5361 gnd.n5360 42.2793
R7937 gnd.n4982 gnd.n4981 42.2793
R7938 gnd.n5287 gnd.n5286 42.2793
R7939 gnd.n4938 gnd.n4937 42.2793
R7940 gnd.n7410 gnd.n7405 42.2793
R7941 gnd.n1799 gnd.n1692 42.2793
R7942 gnd.n2240 gnd.n2239 42.2793
R7943 gnd.n1493 gnd.n1492 42.2793
R7944 gnd.n7462 gnd.n180 42.2793
R7945 gnd.n7499 gnd.n7498 42.2793
R7946 gnd.n4869 gnd.n984 42.2793
R7947 gnd.n1007 gnd.n1006 42.2793
R7948 gnd.n2838 gnd.n2328 42.2793
R7949 gnd.n2494 gnd.n2493 42.2793
R7950 gnd.n2916 gnd.n2915 41.6274
R7951 gnd.n3509 gnd.n3508 41.6274
R7952 gnd.n2925 gnd.n2924 40.8975
R7953 gnd.n3512 gnd.n3511 40.8975
R7954 gnd.n4466 gnd.n1470 36.9518
R7955 gnd.n3114 gnd.n2306 36.9518
R7956 gnd.n6499 gnd.n6498 36.594
R7957 gnd.n6498 gnd.n728 36.594
R7958 gnd.n6492 gnd.n728 36.594
R7959 gnd.n6492 gnd.n6491 36.594
R7960 gnd.n6491 gnd.n6490 36.594
R7961 gnd.n6490 gnd.n736 36.594
R7962 gnd.n6484 gnd.n736 36.594
R7963 gnd.n6484 gnd.n6483 36.594
R7964 gnd.n6483 gnd.n6482 36.594
R7965 gnd.n6482 gnd.n744 36.594
R7966 gnd.n6476 gnd.n744 36.594
R7967 gnd.n6476 gnd.n6475 36.594
R7968 gnd.n6475 gnd.n6474 36.594
R7969 gnd.n6474 gnd.n752 36.594
R7970 gnd.n6468 gnd.n752 36.594
R7971 gnd.n6468 gnd.n6467 36.594
R7972 gnd.n6467 gnd.n6466 36.594
R7973 gnd.n6466 gnd.n760 36.594
R7974 gnd.n6460 gnd.n760 36.594
R7975 gnd.n6460 gnd.n6459 36.594
R7976 gnd.n6459 gnd.n6458 36.594
R7977 gnd.n6458 gnd.n768 36.594
R7978 gnd.n6452 gnd.n768 36.594
R7979 gnd.n6452 gnd.n6451 36.594
R7980 gnd.n6451 gnd.n6450 36.594
R7981 gnd.n6450 gnd.n776 36.594
R7982 gnd.n6444 gnd.n776 36.594
R7983 gnd.n6444 gnd.n6443 36.594
R7984 gnd.n6443 gnd.n6442 36.594
R7985 gnd.n6442 gnd.n784 36.594
R7986 gnd.n6436 gnd.n784 36.594
R7987 gnd.n6436 gnd.n6435 36.594
R7988 gnd.n6435 gnd.n6434 36.594
R7989 gnd.n6434 gnd.n792 36.594
R7990 gnd.n6428 gnd.n792 36.594
R7991 gnd.n6428 gnd.n6427 36.594
R7992 gnd.n6427 gnd.n6426 36.594
R7993 gnd.n6426 gnd.n800 36.594
R7994 gnd.n6420 gnd.n800 36.594
R7995 gnd.n6420 gnd.n6419 36.594
R7996 gnd.n6419 gnd.n6418 36.594
R7997 gnd.n6418 gnd.n808 36.594
R7998 gnd.n6412 gnd.n808 36.594
R7999 gnd.n6412 gnd.n6411 36.594
R8000 gnd.n6411 gnd.n6410 36.594
R8001 gnd.n6410 gnd.n816 36.594
R8002 gnd.n6404 gnd.n816 36.594
R8003 gnd.n6404 gnd.n6403 36.594
R8004 gnd.n6403 gnd.n6402 36.594
R8005 gnd.n6402 gnd.n824 36.594
R8006 gnd.n6396 gnd.n824 36.594
R8007 gnd.n6396 gnd.n6395 36.594
R8008 gnd.n6395 gnd.n6394 36.594
R8009 gnd.n6394 gnd.n832 36.594
R8010 gnd.n6388 gnd.n832 36.594
R8011 gnd.n6388 gnd.n6387 36.594
R8012 gnd.n6387 gnd.n6386 36.594
R8013 gnd.n6386 gnd.n840 36.594
R8014 gnd.n6380 gnd.n840 36.594
R8015 gnd.n6380 gnd.n6379 36.594
R8016 gnd.n6379 gnd.n6378 36.594
R8017 gnd.n6378 gnd.n848 36.594
R8018 gnd.n6372 gnd.n848 36.594
R8019 gnd.n6372 gnd.n6371 36.594
R8020 gnd.n6371 gnd.n6370 36.594
R8021 gnd.n6370 gnd.n856 36.594
R8022 gnd.n6364 gnd.n856 36.594
R8023 gnd.n6364 gnd.n6363 36.594
R8024 gnd.n6363 gnd.n6362 36.594
R8025 gnd.n6362 gnd.n864 36.594
R8026 gnd.n6356 gnd.n864 36.594
R8027 gnd.n6356 gnd.n6355 36.594
R8028 gnd.n6355 gnd.n6354 36.594
R8029 gnd.n6354 gnd.n872 36.594
R8030 gnd.n6348 gnd.n872 36.594
R8031 gnd.n6348 gnd.n6347 36.594
R8032 gnd.n6347 gnd.n6346 36.594
R8033 gnd.n6346 gnd.n880 36.594
R8034 gnd.n6340 gnd.n880 36.594
R8035 gnd.n6340 gnd.n6339 36.594
R8036 gnd.n6339 gnd.n6338 36.594
R8037 gnd.n6338 gnd.n888 36.594
R8038 gnd.n6332 gnd.n888 36.594
R8039 gnd.n2924 gnd.n2923 35.055
R8040 gnd.n2919 gnd.n2918 35.055
R8041 gnd.n3501 gnd.n3500 35.055
R8042 gnd.n3511 gnd.n3497 35.055
R8043 gnd.n5423 gnd.n5317 31.8661
R8044 gnd.n5423 gnd.n5422 31.8661
R8045 gnd.n5431 gnd.n5306 31.8661
R8046 gnd.n5439 gnd.n5306 31.8661
R8047 gnd.n5439 gnd.n5300 31.8661
R8048 gnd.n5447 gnd.n5300 31.8661
R8049 gnd.n5447 gnd.n5293 31.8661
R8050 gnd.n5571 gnd.n5293 31.8661
R8051 gnd.n5581 gnd.n5226 31.8661
R8052 gnd.n2550 gnd.n961 31.8661
R8053 gnd.n4818 gnd.n1015 31.8661
R8054 gnd.n4818 gnd.n1017 31.8661
R8055 gnd.n4812 gnd.n1017 31.8661
R8056 gnd.n4812 gnd.n1029 31.8661
R8057 gnd.n4806 gnd.n1040 31.8661
R8058 gnd.n4800 gnd.n1040 31.8661
R8059 gnd.n4794 gnd.n1057 31.8661
R8060 gnd.n4788 gnd.n1067 31.8661
R8061 gnd.n4788 gnd.n1070 31.8661
R8062 gnd.n4782 gnd.n1080 31.8661
R8063 gnd.n4776 gnd.n1080 31.8661
R8064 gnd.n4770 gnd.n1098 31.8661
R8065 gnd.n2249 gnd.n1273 31.8661
R8066 gnd.n2757 gnd.n2265 31.8661
R8067 gnd.n2757 gnd.n2181 31.8661
R8068 gnd.n3202 gnd.n2175 31.8661
R8069 gnd.n3202 gnd.n2176 31.8661
R8070 gnd.n3210 gnd.n2164 31.8661
R8071 gnd.n3218 gnd.n2164 31.8661
R8072 gnd.n3218 gnd.n2157 31.8661
R8073 gnd.n3226 gnd.n2157 31.8661
R8074 gnd.n3234 gnd.n2151 31.8661
R8075 gnd.n3234 gnd.n2142 31.8661
R8076 gnd.n3242 gnd.n2142 31.8661
R8077 gnd.n3242 gnd.n2144 31.8661
R8078 gnd.n3250 gnd.n2129 31.8661
R8079 gnd.n3258 gnd.n2129 31.8661
R8080 gnd.n3258 gnd.n2131 31.8661
R8081 gnd.n4130 gnd.n1878 31.8661
R8082 gnd.n4146 gnd.n1864 31.8661
R8083 gnd.n4146 gnd.n1858 31.8661
R8084 gnd.n4154 gnd.n1858 31.8661
R8085 gnd.n4162 gnd.n1851 31.8661
R8086 gnd.n4162 gnd.n1844 31.8661
R8087 gnd.n4170 gnd.n1844 31.8661
R8088 gnd.n4170 gnd.n1845 31.8661
R8089 gnd.n4178 gnd.n1831 31.8661
R8090 gnd.n4188 gnd.n1831 31.8661
R8091 gnd.n4188 gnd.n1823 31.8661
R8092 gnd.n4199 gnd.n1823 31.8661
R8093 gnd.n4507 gnd.n1406 31.8661
R8094 gnd.n4507 gnd.n4506 31.8661
R8095 gnd.n4500 gnd.n1417 31.8661
R8096 gnd.n4500 gnd.n4499 31.8661
R8097 gnd.n1497 gnd.n1446 31.8661
R8098 gnd.n7315 gnd.n248 31.8661
R8099 gnd.n7323 gnd.n238 31.8661
R8100 gnd.n7323 gnd.n241 31.8661
R8101 gnd.n7331 gnd.n225 31.8661
R8102 gnd.n7339 gnd.n225 31.8661
R8103 gnd.n7347 gnd.n218 31.8661
R8104 gnd.n7355 gnd.n208 31.8661
R8105 gnd.n7355 gnd.n211 31.8661
R8106 gnd.n7363 gnd.n193 31.8661
R8107 gnd.n7446 gnd.n193 31.8661
R8108 gnd.n7446 gnd.n185 31.8661
R8109 gnd.n7454 gnd.n185 31.8661
R8110 gnd.n7534 gnd.n104 31.8661
R8111 gnd.n3568 gnd.n3492 31.3761
R8112 gnd.n3048 gnd.n2900 31.3761
R8113 gnd.n3266 gnd.n2123 30.9101
R8114 gnd.n2122 gnd.t144 30.5915
R8115 gnd.n4794 gnd.t177 27.7236
R8116 gnd.t179 gnd.n218 27.7236
R8117 gnd.n2131 gnd.t301 27.0862
R8118 gnd.t213 gnd.n1864 27.0862
R8119 gnd.n4138 gnd.t112 26.1303
R8120 gnd.n2809 gnd.n2808 25.7944
R8121 gnd.n5286 gnd.n5285 25.7944
R8122 gnd.n4937 gnd.n4936 25.7944
R8123 gnd.n7405 gnd.n7404 25.7944
R8124 gnd.n1692 gnd.n1691 25.7944
R8125 gnd.n2239 gnd.n2238 25.7944
R8126 gnd.n1470 gnd.n1469 25.7944
R8127 gnd.n1492 gnd.n1491 25.7944
R8128 gnd.n180 gnd.n179 25.7944
R8129 gnd.n7498 gnd.n7497 25.7944
R8130 gnd.n984 gnd.n983 25.7944
R8131 gnd.n1006 gnd.n1005 25.7944
R8132 gnd.n2328 gnd.n2327 25.7944
R8133 gnd.n2306 gnd.n2305 25.7944
R8134 gnd.n2493 gnd.n2492 25.7944
R8135 gnd.n4217 gnd.n4216 25.7944
R8136 gnd.n1057 gnd.t257 25.1743
R8137 gnd.n7347 gnd.t27 25.1743
R8138 gnd.n5593 gnd.n5227 24.8557
R8139 gnd.n5603 gnd.n5210 24.8557
R8140 gnd.n5213 gnd.n5201 24.8557
R8141 gnd.n5624 gnd.n5202 24.8557
R8142 gnd.n5634 gnd.n5184 24.8557
R8143 gnd.n5645 gnd.n5644 24.8557
R8144 gnd.n5664 gnd.n5170 24.8557
R8145 gnd.n5665 gnd.n5159 24.8557
R8146 gnd.n5676 gnd.n5675 24.8557
R8147 gnd.n5686 gnd.n5152 24.8557
R8148 gnd.n5695 gnd.n5144 24.8557
R8149 gnd.n5707 gnd.n5706 24.8557
R8150 gnd.n5482 gnd.n5136 24.8557
R8151 gnd.n5717 gnd.n5126 24.8557
R8152 gnd.n5726 gnd.n5119 24.8557
R8153 gnd.n5112 gnd.n5102 24.8557
R8154 gnd.n5095 gnd.n5089 24.8557
R8155 gnd.n5781 gnd.n5780 24.8557
R8156 gnd.n5791 gnd.n5790 24.8557
R8157 gnd.n5080 gnd.n5072 24.8557
R8158 gnd.n5802 gnd.n5057 24.8557
R8159 gnd.n5821 gnd.n5820 24.8557
R8160 gnd.n5831 gnd.n5050 24.8557
R8161 gnd.n5844 gnd.n5039 24.8557
R8162 gnd.n5835 gnd.n5834 24.8557
R8163 gnd.n5867 gnd.n5866 24.8557
R8164 gnd.n5877 gnd.n5026 24.8557
R8165 gnd.n5889 gnd.n5018 24.8557
R8166 gnd.n6188 gnd.n6187 24.8557
R8167 gnd.n6203 gnd.n6202 24.8557
R8168 gnd.n6324 gnd.n907 24.8557
R8169 gnd.n6323 gnd.n910 24.8557
R8170 gnd.n6172 gnd.n919 24.8557
R8171 gnd.n6310 gnd.n930 24.8557
R8172 gnd.n2176 gnd.t115 24.537
R8173 gnd.n3250 gnd.t4 24.537
R8174 gnd.n4154 gnd.t235 24.537
R8175 gnd.t72 gnd.n1406 24.537
R8176 gnd.n3193 gnd.n2175 23.8997
R8177 gnd.n4506 gnd.n1409 23.8997
R8178 gnd.n5614 gnd.t312 23.2624
R8179 gnd.n5229 gnd.t147 22.6251
R8180 gnd.n2550 gnd.t64 22.6251
R8181 gnd.t84 gnd.n104 22.6251
R8182 gnd.n6332 gnd.n6331 21.9566
R8183 gnd.n3043 gnd.n2116 21.6691
R8184 gnd.n3890 gnd.n2076 21.6691
R8185 gnd.n3875 gnd.n2061 21.6691
R8186 gnd.n3868 gnd.n2053 21.6691
R8187 gnd.n3860 gnd.n2046 21.6691
R8188 gnd.n3853 gnd.n2038 21.6691
R8189 gnd.n3845 gnd.n2031 21.6691
R8190 gnd.n3838 gnd.n2024 21.6691
R8191 gnd.n3810 gnd.n1985 21.6691
R8192 gnd.n4034 gnd.n1957 21.6691
R8193 gnd.n3768 gnd.n1949 21.6691
R8194 gnd.n3760 gnd.n1943 21.6691
R8195 gnd.n3753 gnd.n1936 21.6691
R8196 gnd.n3745 gnd.n3442 21.6691
R8197 gnd.n3739 gnd.n3738 21.6691
R8198 gnd.n3724 gnd.n3723 21.6691
R8199 gnd.n3470 gnd.n1897 21.6691
R8200 gnd.n3708 gnd.n1890 21.6691
R8201 gnd.t17 gnd.n5234 21.3504
R8202 gnd.t119 gnd.n2103 21.0318
R8203 gnd.t9 gnd.n5003 20.7131
R8204 gnd.n1097 gnd.t56 20.3945
R8205 gnd.n3022 gnd.n2095 20.3945
R8206 gnd.n3906 gnd.n2074 20.3945
R8207 gnd.n3722 gnd.n1904 20.3945
R8208 gnd.n250 gnd.t58 20.3945
R8209 gnd.t44 gnd.n5049 20.0758
R8210 gnd.t25 gnd.n2068 20.0758
R8211 gnd.n3457 gnd.t252 20.0758
R8212 gnd.n2885 gnd.n2884 19.9763
R8213 gnd.n3544 gnd.n3543 19.9763
R8214 gnd.n2943 gnd.n2942 19.9763
R8215 gnd.n3538 gnd.n3537 19.9763
R8216 gnd.n2912 gnd.t120 19.8005
R8217 gnd.n2912 gnd.t130 19.8005
R8218 gnd.n2913 gnd.t100 19.8005
R8219 gnd.n2913 gnd.t136 19.8005
R8220 gnd.n3505 gnd.t123 19.8005
R8221 gnd.n3505 gnd.t113 19.8005
R8222 gnd.n3506 gnd.t62 19.8005
R8223 gnd.n3506 gnd.t164 19.8005
R8224 gnd.n3143 gnd.n2265 19.7572
R8225 gnd.n4499 gnd.n4498 19.7572
R8226 gnd.n2909 gnd.n2908 19.5087
R8227 gnd.n2922 gnd.n2909 19.5087
R8228 gnd.n2920 gnd.n2911 19.5087
R8229 gnd.n3510 gnd.n3504 19.5087
R8230 gnd.n5757 gnd.t54 19.4385
R8231 gnd.n3226 gnd.t15 19.4385
R8232 gnd.n4178 gnd.t283 19.4385
R8233 gnd.n3200 gnd.n2168 19.3944
R8234 gnd.n3212 gnd.n2168 19.3944
R8235 gnd.n3212 gnd.n2166 19.3944
R8236 gnd.n3216 gnd.n2166 19.3944
R8237 gnd.n3216 gnd.n2155 19.3944
R8238 gnd.n3228 gnd.n2155 19.3944
R8239 gnd.n3228 gnd.n2153 19.3944
R8240 gnd.n3232 gnd.n2153 19.3944
R8241 gnd.n3232 gnd.n2140 19.3944
R8242 gnd.n3244 gnd.n2140 19.3944
R8243 gnd.n3244 gnd.n2138 19.3944
R8244 gnd.n3248 gnd.n2138 19.3944
R8245 gnd.n3248 gnd.n2127 19.3944
R8246 gnd.n3260 gnd.n2127 19.3944
R8247 gnd.n3260 gnd.n2125 19.3944
R8248 gnd.n3264 gnd.n2125 19.3944
R8249 gnd.n3264 gnd.n2114 19.3944
R8250 gnd.n3276 gnd.n2114 19.3944
R8251 gnd.n3276 gnd.n2112 19.3944
R8252 gnd.n3280 gnd.n2112 19.3944
R8253 gnd.n3280 gnd.n2100 19.3944
R8254 gnd.n3294 gnd.n2100 19.3944
R8255 gnd.n3294 gnd.n2097 19.3944
R8256 gnd.n3299 gnd.n2097 19.3944
R8257 gnd.n3299 gnd.n2098 19.3944
R8258 gnd.n2098 gnd.n2072 19.3944
R8259 gnd.n3908 gnd.n2072 19.3944
R8260 gnd.n3908 gnd.n2070 19.3944
R8261 gnd.n3912 gnd.n2070 19.3944
R8262 gnd.n3912 gnd.n2057 19.3944
R8263 gnd.n3924 gnd.n2057 19.3944
R8264 gnd.n3924 gnd.n2055 19.3944
R8265 gnd.n3928 gnd.n2055 19.3944
R8266 gnd.n3928 gnd.n2042 19.3944
R8267 gnd.n3940 gnd.n2042 19.3944
R8268 gnd.n3940 gnd.n2040 19.3944
R8269 gnd.n3944 gnd.n2040 19.3944
R8270 gnd.n3944 gnd.n2028 19.3944
R8271 gnd.n3956 gnd.n2028 19.3944
R8272 gnd.n3956 gnd.n2026 19.3944
R8273 gnd.n3960 gnd.n2026 19.3944
R8274 gnd.n3960 gnd.n2013 19.3944
R8275 gnd.n3972 gnd.n2013 19.3944
R8276 gnd.n3972 gnd.n2011 19.3944
R8277 gnd.n3976 gnd.n2011 19.3944
R8278 gnd.n3976 gnd.n1998 19.3944
R8279 gnd.n3988 gnd.n1998 19.3944
R8280 gnd.n3988 gnd.n1996 19.3944
R8281 gnd.n3992 gnd.n1996 19.3944
R8282 gnd.n3992 gnd.n1983 19.3944
R8283 gnd.n4004 gnd.n1983 19.3944
R8284 gnd.n4004 gnd.n1981 19.3944
R8285 gnd.n4008 gnd.n1981 19.3944
R8286 gnd.n4008 gnd.n1968 19.3944
R8287 gnd.n4020 gnd.n1968 19.3944
R8288 gnd.n4020 gnd.n1966 19.3944
R8289 gnd.n4024 gnd.n1966 19.3944
R8290 gnd.n4024 gnd.n1953 19.3944
R8291 gnd.n4036 gnd.n1953 19.3944
R8292 gnd.n4036 gnd.n1951 19.3944
R8293 gnd.n4040 gnd.n1951 19.3944
R8294 gnd.n4040 gnd.n1940 19.3944
R8295 gnd.n4052 gnd.n1940 19.3944
R8296 gnd.n4052 gnd.n1938 19.3944
R8297 gnd.n4056 gnd.n1938 19.3944
R8298 gnd.n4056 gnd.n1928 19.3944
R8299 gnd.n4068 gnd.n1928 19.3944
R8300 gnd.n4068 gnd.n1926 19.3944
R8301 gnd.n4072 gnd.n1926 19.3944
R8302 gnd.n4072 gnd.n1915 19.3944
R8303 gnd.n4084 gnd.n1915 19.3944
R8304 gnd.n4084 gnd.n1913 19.3944
R8305 gnd.n4088 gnd.n1913 19.3944
R8306 gnd.n4088 gnd.n1902 19.3944
R8307 gnd.n4100 gnd.n1902 19.3944
R8308 gnd.n4100 gnd.n1900 19.3944
R8309 gnd.n4104 gnd.n1900 19.3944
R8310 gnd.n4104 gnd.n1888 19.3944
R8311 gnd.n4116 gnd.n1888 19.3944
R8312 gnd.n4116 gnd.n1886 19.3944
R8313 gnd.n4120 gnd.n1886 19.3944
R8314 gnd.n4120 gnd.n1874 19.3944
R8315 gnd.n4132 gnd.n1874 19.3944
R8316 gnd.n4132 gnd.n1872 19.3944
R8317 gnd.n4136 gnd.n1872 19.3944
R8318 gnd.n4136 gnd.n1862 19.3944
R8319 gnd.n4148 gnd.n1862 19.3944
R8320 gnd.n4148 gnd.n1860 19.3944
R8321 gnd.n4152 gnd.n1860 19.3944
R8322 gnd.n4152 gnd.n1849 19.3944
R8323 gnd.n4164 gnd.n1849 19.3944
R8324 gnd.n4164 gnd.n1847 19.3944
R8325 gnd.n4168 gnd.n1847 19.3944
R8326 gnd.n4168 gnd.n1836 19.3944
R8327 gnd.n4180 gnd.n1836 19.3944
R8328 gnd.n4180 gnd.n1833 19.3944
R8329 gnd.n4186 gnd.n1833 19.3944
R8330 gnd.n4186 gnd.n1834 19.3944
R8331 gnd.n1834 gnd.n1821 19.3944
R8332 gnd.n4202 gnd.n1821 19.3944
R8333 gnd.n4203 gnd.n4202 19.3944
R8334 gnd.n2813 gnd.n2179 19.3944
R8335 gnd.n3196 gnd.n2179 19.3944
R8336 gnd.n3197 gnd.n3196 19.3944
R8337 gnd.n3190 gnd.n3189 19.3944
R8338 gnd.n3189 gnd.n2197 19.3944
R8339 gnd.n3182 gnd.n2197 19.3944
R8340 gnd.n3182 gnd.n3181 19.3944
R8341 gnd.n3181 gnd.n2208 19.3944
R8342 gnd.n3174 gnd.n2208 19.3944
R8343 gnd.n3174 gnd.n3173 19.3944
R8344 gnd.n3173 gnd.n2216 19.3944
R8345 gnd.n3166 gnd.n2216 19.3944
R8346 gnd.n3166 gnd.n3165 19.3944
R8347 gnd.n3165 gnd.n2226 19.3944
R8348 gnd.n3158 gnd.n2226 19.3944
R8349 gnd.n3158 gnd.n3157 19.3944
R8350 gnd.n3157 gnd.n2234 19.3944
R8351 gnd.n3150 gnd.n2234 19.3944
R8352 gnd.n3150 gnd.n3149 19.3944
R8353 gnd.n3149 gnd.n2246 19.3944
R8354 gnd.n2824 gnd.n2246 19.3944
R8355 gnd.n2824 gnd.n2823 19.3944
R8356 gnd.n2823 gnd.n2822 19.3944
R8357 gnd.n2822 gnd.n2803 19.3944
R8358 gnd.n2818 gnd.n2803 19.3944
R8359 gnd.n2818 gnd.n2817 19.3944
R8360 gnd.n2817 gnd.n2816 19.3944
R8361 gnd.n5410 gnd.n5409 19.3944
R8362 gnd.n5409 gnd.n5408 19.3944
R8363 gnd.n5408 gnd.n5407 19.3944
R8364 gnd.n5407 gnd.n5405 19.3944
R8365 gnd.n5405 gnd.n5402 19.3944
R8366 gnd.n5402 gnd.n5401 19.3944
R8367 gnd.n5401 gnd.n5398 19.3944
R8368 gnd.n5398 gnd.n5397 19.3944
R8369 gnd.n5397 gnd.n5394 19.3944
R8370 gnd.n5394 gnd.n5393 19.3944
R8371 gnd.n5393 gnd.n5390 19.3944
R8372 gnd.n5390 gnd.n5389 19.3944
R8373 gnd.n5389 gnd.n5386 19.3944
R8374 gnd.n5386 gnd.n5385 19.3944
R8375 gnd.n5385 gnd.n5382 19.3944
R8376 gnd.n5382 gnd.n5381 19.3944
R8377 gnd.n5381 gnd.n5378 19.3944
R8378 gnd.n5378 gnd.n5377 19.3944
R8379 gnd.n5377 gnd.n5374 19.3944
R8380 gnd.n5374 gnd.n5373 19.3944
R8381 gnd.n5373 gnd.n5370 19.3944
R8382 gnd.n5370 gnd.n5369 19.3944
R8383 gnd.n5366 gnd.n5365 19.3944
R8384 gnd.n5365 gnd.n5321 19.3944
R8385 gnd.n5416 gnd.n5321 19.3944
R8386 gnd.n6230 gnd.n4984 19.3944
R8387 gnd.n6230 gnd.n6229 19.3944
R8388 gnd.n6229 gnd.n6228 19.3944
R8389 gnd.n6272 gnd.n6271 19.3944
R8390 gnd.n6271 gnd.n6270 19.3944
R8391 gnd.n6270 gnd.n4945 19.3944
R8392 gnd.n6265 gnd.n4945 19.3944
R8393 gnd.n6265 gnd.n6264 19.3944
R8394 gnd.n6264 gnd.n6263 19.3944
R8395 gnd.n6263 gnd.n4952 19.3944
R8396 gnd.n6258 gnd.n4952 19.3944
R8397 gnd.n6258 gnd.n6257 19.3944
R8398 gnd.n6257 gnd.n6256 19.3944
R8399 gnd.n6256 gnd.n4959 19.3944
R8400 gnd.n6251 gnd.n4959 19.3944
R8401 gnd.n6251 gnd.n6250 19.3944
R8402 gnd.n6250 gnd.n6249 19.3944
R8403 gnd.n6249 gnd.n4966 19.3944
R8404 gnd.n6244 gnd.n4966 19.3944
R8405 gnd.n6244 gnd.n6243 19.3944
R8406 gnd.n6243 gnd.n6242 19.3944
R8407 gnd.n6242 gnd.n4973 19.3944
R8408 gnd.n6237 gnd.n4973 19.3944
R8409 gnd.n6237 gnd.n6236 19.3944
R8410 gnd.n6236 gnd.n6235 19.3944
R8411 gnd.n5595 gnd.n5218 19.3944
R8412 gnd.n5605 gnd.n5218 19.3944
R8413 gnd.n5606 gnd.n5605 19.3944
R8414 gnd.n5606 gnd.n5199 19.3944
R8415 gnd.n5626 gnd.n5199 19.3944
R8416 gnd.n5626 gnd.n5192 19.3944
R8417 gnd.n5636 gnd.n5192 19.3944
R8418 gnd.n5637 gnd.n5636 19.3944
R8419 gnd.n5637 gnd.n5175 19.3944
R8420 gnd.n5657 gnd.n5175 19.3944
R8421 gnd.n5657 gnd.n5167 19.3944
R8422 gnd.n5667 gnd.n5167 19.3944
R8423 gnd.n5668 gnd.n5667 19.3944
R8424 gnd.n5668 gnd.n5149 19.3944
R8425 gnd.n5688 gnd.n5149 19.3944
R8426 gnd.n5688 gnd.n5141 19.3944
R8427 gnd.n5698 gnd.n5141 19.3944
R8428 gnd.n5699 gnd.n5698 19.3944
R8429 gnd.n5699 gnd.n5124 19.3944
R8430 gnd.n5719 gnd.n5124 19.3944
R8431 gnd.n5719 gnd.n5116 19.3944
R8432 gnd.n5729 gnd.n5116 19.3944
R8433 gnd.n5730 gnd.n5729 19.3944
R8434 gnd.n5730 gnd.n5100 19.3944
R8435 gnd.n5749 gnd.n5100 19.3944
R8436 gnd.n5749 gnd.n5085 19.3944
R8437 gnd.n5783 gnd.n5085 19.3944
R8438 gnd.n5784 gnd.n5783 19.3944
R8439 gnd.n5785 gnd.n5784 19.3944
R8440 gnd.n5785 gnd.n5071 19.3944
R8441 gnd.n5071 gnd.n5065 19.3944
R8442 gnd.n5810 gnd.n5065 19.3944
R8443 gnd.n5811 gnd.n5810 19.3944
R8444 gnd.n5811 gnd.n5048 19.3944
R8445 gnd.n5048 gnd.n5046 19.3944
R8446 gnd.n5837 gnd.n5046 19.3944
R8447 gnd.n5838 gnd.n5837 19.3944
R8448 gnd.n5838 gnd.n5021 19.3944
R8449 gnd.n5884 gnd.n5021 19.3944
R8450 gnd.n5885 gnd.n5884 19.3944
R8451 gnd.n5885 gnd.n5014 19.3944
R8452 gnd.n5896 gnd.n5014 19.3944
R8453 gnd.n5898 gnd.n5896 19.3944
R8454 gnd.n6181 gnd.n5898 19.3944
R8455 gnd.n6181 gnd.n6180 19.3944
R8456 gnd.n6180 gnd.n5901 19.3944
R8457 gnd.n6176 gnd.n5901 19.3944
R8458 gnd.n6176 gnd.n6175 19.3944
R8459 gnd.n6175 gnd.n6174 19.3944
R8460 gnd.n6174 gnd.n6171 19.3944
R8461 gnd.n6171 gnd.n6170 19.3944
R8462 gnd.n6170 gnd.n6167 19.3944
R8463 gnd.n6167 gnd.n6166 19.3944
R8464 gnd.n5586 gnd.n5585 19.3944
R8465 gnd.n5585 gnd.n5232 19.3944
R8466 gnd.n5255 gnd.n5232 19.3944
R8467 gnd.n5258 gnd.n5255 19.3944
R8468 gnd.n5258 gnd.n5251 19.3944
R8469 gnd.n5262 gnd.n5251 19.3944
R8470 gnd.n5265 gnd.n5262 19.3944
R8471 gnd.n5268 gnd.n5265 19.3944
R8472 gnd.n5268 gnd.n5249 19.3944
R8473 gnd.n5272 gnd.n5249 19.3944
R8474 gnd.n5275 gnd.n5272 19.3944
R8475 gnd.n5278 gnd.n5275 19.3944
R8476 gnd.n5278 gnd.n5247 19.3944
R8477 gnd.n5282 gnd.n5247 19.3944
R8478 gnd.n5591 gnd.n5590 19.3944
R8479 gnd.n5590 gnd.n5208 19.3944
R8480 gnd.n5616 gnd.n5208 19.3944
R8481 gnd.n5616 gnd.n5206 19.3944
R8482 gnd.n5622 gnd.n5206 19.3944
R8483 gnd.n5622 gnd.n5621 19.3944
R8484 gnd.n5621 gnd.n5182 19.3944
R8485 gnd.n5647 gnd.n5182 19.3944
R8486 gnd.n5647 gnd.n5180 19.3944
R8487 gnd.n5653 gnd.n5180 19.3944
R8488 gnd.n5653 gnd.n5652 19.3944
R8489 gnd.n5652 gnd.n5157 19.3944
R8490 gnd.n5678 gnd.n5157 19.3944
R8491 gnd.n5678 gnd.n5155 19.3944
R8492 gnd.n5684 gnd.n5155 19.3944
R8493 gnd.n5684 gnd.n5683 19.3944
R8494 gnd.n5683 gnd.n5131 19.3944
R8495 gnd.n5709 gnd.n5131 19.3944
R8496 gnd.n5709 gnd.n5129 19.3944
R8497 gnd.n5715 gnd.n5129 19.3944
R8498 gnd.n5715 gnd.n5714 19.3944
R8499 gnd.n5714 gnd.n5107 19.3944
R8500 gnd.n5739 gnd.n5107 19.3944
R8501 gnd.n5739 gnd.n5105 19.3944
R8502 gnd.n5745 gnd.n5105 19.3944
R8503 gnd.n5745 gnd.n5744 19.3944
R8504 gnd.n5744 gnd.n5076 19.3944
R8505 gnd.n5793 gnd.n5076 19.3944
R8506 gnd.n5793 gnd.n5074 19.3944
R8507 gnd.n5797 gnd.n5074 19.3944
R8508 gnd.n5797 gnd.n5055 19.3944
R8509 gnd.n5823 gnd.n5055 19.3944
R8510 gnd.n5823 gnd.n5053 19.3944
R8511 gnd.n5829 gnd.n5053 19.3944
R8512 gnd.n5829 gnd.n5828 19.3944
R8513 gnd.n5828 gnd.n5031 19.3944
R8514 gnd.n5869 gnd.n5031 19.3944
R8515 gnd.n5869 gnd.n5029 19.3944
R8516 gnd.n5875 gnd.n5029 19.3944
R8517 gnd.n5875 gnd.n5874 19.3944
R8518 gnd.n5874 gnd.n5001 19.3944
R8519 gnd.n6190 gnd.n5001 19.3944
R8520 gnd.n6190 gnd.n4999 19.3944
R8521 gnd.n6200 gnd.n4999 19.3944
R8522 gnd.n6200 gnd.n6199 19.3944
R8523 gnd.n6199 gnd.n6198 19.3944
R8524 gnd.n6198 gnd.n913 19.3944
R8525 gnd.n6321 gnd.n913 19.3944
R8526 gnd.n6321 gnd.n6320 19.3944
R8527 gnd.n6320 gnd.n6319 19.3944
R8528 gnd.n6319 gnd.n917 19.3944
R8529 gnd.n4909 gnd.n917 19.3944
R8530 gnd.n6307 gnd.n4909 19.3944
R8531 gnd.n6304 gnd.n6303 19.3944
R8532 gnd.n6303 gnd.n6302 19.3944
R8533 gnd.n6302 gnd.n4915 19.3944
R8534 gnd.n6297 gnd.n4915 19.3944
R8535 gnd.n6297 gnd.n6296 19.3944
R8536 gnd.n6296 gnd.n6295 19.3944
R8537 gnd.n6295 gnd.n4922 19.3944
R8538 gnd.n6290 gnd.n4922 19.3944
R8539 gnd.n6290 gnd.n6289 19.3944
R8540 gnd.n6289 gnd.n6288 19.3944
R8541 gnd.n6288 gnd.n4929 19.3944
R8542 gnd.n6283 gnd.n4929 19.3944
R8543 gnd.n6283 gnd.n6282 19.3944
R8544 gnd.n6282 gnd.n6281 19.3944
R8545 gnd.n5420 gnd.n5319 19.3944
R8546 gnd.n5420 gnd.n5310 19.3944
R8547 gnd.n5433 gnd.n5310 19.3944
R8548 gnd.n5433 gnd.n5308 19.3944
R8549 gnd.n5437 gnd.n5308 19.3944
R8550 gnd.n5437 gnd.n5298 19.3944
R8551 gnd.n5449 gnd.n5298 19.3944
R8552 gnd.n5449 gnd.n5296 19.3944
R8553 gnd.n5569 gnd.n5296 19.3944
R8554 gnd.n5569 gnd.n5568 19.3944
R8555 gnd.n5568 gnd.n5567 19.3944
R8556 gnd.n5567 gnd.n5566 19.3944
R8557 gnd.n5566 gnd.n5563 19.3944
R8558 gnd.n5563 gnd.n5562 19.3944
R8559 gnd.n5562 gnd.n5561 19.3944
R8560 gnd.n5561 gnd.n5559 19.3944
R8561 gnd.n5559 gnd.n5558 19.3944
R8562 gnd.n5558 gnd.n5555 19.3944
R8563 gnd.n5555 gnd.n5554 19.3944
R8564 gnd.n5554 gnd.n5553 19.3944
R8565 gnd.n5553 gnd.n5551 19.3944
R8566 gnd.n5551 gnd.n5550 19.3944
R8567 gnd.n5550 gnd.n5546 19.3944
R8568 gnd.n5546 gnd.n5545 19.3944
R8569 gnd.n5545 gnd.n5544 19.3944
R8570 gnd.n5544 gnd.n5542 19.3944
R8571 gnd.n5542 gnd.n5541 19.3944
R8572 gnd.n5541 gnd.n5538 19.3944
R8573 gnd.n5538 gnd.n5537 19.3944
R8574 gnd.n5485 gnd.n5473 19.3944
R8575 gnd.n5484 gnd.n5480 19.3944
R8576 gnd.n5478 gnd.n5477 19.3944
R8577 gnd.n5474 gnd.n5093 19.3944
R8578 gnd.n5759 gnd.n5093 19.3944
R8579 gnd.n5759 gnd.n5091 19.3944
R8580 gnd.n5778 gnd.n5091 19.3944
R8581 gnd.n5778 gnd.n5777 19.3944
R8582 gnd.n5777 gnd.n5776 19.3944
R8583 gnd.n5776 gnd.n5774 19.3944
R8584 gnd.n5774 gnd.n5773 19.3944
R8585 gnd.n5773 gnd.n5771 19.3944
R8586 gnd.n5771 gnd.n5770 19.3944
R8587 gnd.n5770 gnd.n5037 19.3944
R8588 gnd.n5846 gnd.n5037 19.3944
R8589 gnd.n5846 gnd.n5035 19.3944
R8590 gnd.n5862 gnd.n5035 19.3944
R8591 gnd.n5862 gnd.n5861 19.3944
R8592 gnd.n5861 gnd.n5860 19.3944
R8593 gnd.n5860 gnd.n5858 19.3944
R8594 gnd.n5858 gnd.n5857 19.3944
R8595 gnd.n5857 gnd.n5855 19.3944
R8596 gnd.n5855 gnd.n4994 19.3944
R8597 gnd.n6205 gnd.n4994 19.3944
R8598 gnd.n6205 gnd.n4992 19.3944
R8599 gnd.n6211 gnd.n4992 19.3944
R8600 gnd.n6212 gnd.n6211 19.3944
R8601 gnd.n6215 gnd.n6212 19.3944
R8602 gnd.n6215 gnd.n4990 19.3944
R8603 gnd.n6219 gnd.n4990 19.3944
R8604 gnd.n6222 gnd.n6219 19.3944
R8605 gnd.n6223 gnd.n6222 19.3944
R8606 gnd.n5425 gnd.n5315 19.3944
R8607 gnd.n5425 gnd.n5313 19.3944
R8608 gnd.n5429 gnd.n5313 19.3944
R8609 gnd.n5429 gnd.n5304 19.3944
R8610 gnd.n5441 gnd.n5304 19.3944
R8611 gnd.n5441 gnd.n5302 19.3944
R8612 gnd.n5445 gnd.n5302 19.3944
R8613 gnd.n5445 gnd.n5291 19.3944
R8614 gnd.n5573 gnd.n5291 19.3944
R8615 gnd.n5573 gnd.n5245 19.3944
R8616 gnd.n5579 gnd.n5245 19.3944
R8617 gnd.n5579 gnd.n5578 19.3944
R8618 gnd.n5578 gnd.n5223 19.3944
R8619 gnd.n5600 gnd.n5223 19.3944
R8620 gnd.n5600 gnd.n5216 19.3944
R8621 gnd.n5611 gnd.n5216 19.3944
R8622 gnd.n5611 gnd.n5610 19.3944
R8623 gnd.n5610 gnd.n5197 19.3944
R8624 gnd.n5631 gnd.n5197 19.3944
R8625 gnd.n5631 gnd.n5190 19.3944
R8626 gnd.n5642 gnd.n5190 19.3944
R8627 gnd.n5642 gnd.n5641 19.3944
R8628 gnd.n5641 gnd.n5173 19.3944
R8629 gnd.n5662 gnd.n5173 19.3944
R8630 gnd.n5662 gnd.n5165 19.3944
R8631 gnd.n5673 gnd.n5165 19.3944
R8632 gnd.n5673 gnd.n5672 19.3944
R8633 gnd.n5672 gnd.n5147 19.3944
R8634 gnd.n5693 gnd.n5147 19.3944
R8635 gnd.n5693 gnd.n5139 19.3944
R8636 gnd.n5704 gnd.n5139 19.3944
R8637 gnd.n5704 gnd.n5703 19.3944
R8638 gnd.n5703 gnd.n5122 19.3944
R8639 gnd.n5724 gnd.n5122 19.3944
R8640 gnd.n5724 gnd.n5114 19.3944
R8641 gnd.n5734 gnd.n5114 19.3944
R8642 gnd.n5734 gnd.n5098 19.3944
R8643 gnd.n5755 gnd.n5098 19.3944
R8644 gnd.n5755 gnd.n5754 19.3944
R8645 gnd.n5754 gnd.n5082 19.3944
R8646 gnd.n5788 gnd.n5082 19.3944
R8647 gnd.n5788 gnd.n5067 19.3944
R8648 gnd.n5805 gnd.n5067 19.3944
R8649 gnd.n5805 gnd.n5063 19.3944
R8650 gnd.n5818 gnd.n5063 19.3944
R8651 gnd.n5818 gnd.n5817 19.3944
R8652 gnd.n5817 gnd.n5042 19.3944
R8653 gnd.n5842 gnd.n5042 19.3944
R8654 gnd.n5842 gnd.n5841 19.3944
R8655 gnd.n5841 gnd.n5023 19.3944
R8656 gnd.n5880 gnd.n5023 19.3944
R8657 gnd.n5880 gnd.n5016 19.3944
R8658 gnd.n5891 gnd.n5016 19.3944
R8659 gnd.n5891 gnd.n5010 19.3944
R8660 gnd.n6185 gnd.n5010 19.3944
R8661 gnd.n6185 gnd.n6184 19.3944
R8662 gnd.n6184 gnd.n901 19.3944
R8663 gnd.n6328 gnd.n901 19.3944
R8664 gnd.n6328 gnd.n6327 19.3944
R8665 gnd.n6327 gnd.n6326 19.3944
R8666 gnd.n6326 gnd.n905 19.3944
R8667 gnd.n925 gnd.n905 19.3944
R8668 gnd.n6314 gnd.n925 19.3944
R8669 gnd.n6314 gnd.n6313 19.3944
R8670 gnd.n6313 gnd.n6312 19.3944
R8671 gnd.n4229 gnd.n1681 19.3944
R8672 gnd.n4234 gnd.n1681 19.3944
R8673 gnd.n4234 gnd.n1682 19.3944
R8674 gnd.n1682 gnd.n1613 19.3944
R8675 gnd.n4260 gnd.n1613 19.3944
R8676 gnd.n4260 gnd.n1610 19.3944
R8677 gnd.n4265 gnd.n1610 19.3944
R8678 gnd.n4265 gnd.n1611 19.3944
R8679 gnd.n1611 gnd.n1586 19.3944
R8680 gnd.n4291 gnd.n1586 19.3944
R8681 gnd.n4291 gnd.n1583 19.3944
R8682 gnd.n4301 gnd.n1583 19.3944
R8683 gnd.n4301 gnd.n1584 19.3944
R8684 gnd.n4297 gnd.n1584 19.3944
R8685 gnd.n4297 gnd.n4296 19.3944
R8686 gnd.n4296 gnd.n1549 19.3944
R8687 gnd.n4358 gnd.n1549 19.3944
R8688 gnd.n4358 gnd.n1550 19.3944
R8689 gnd.n4354 gnd.n1550 19.3944
R8690 gnd.n4354 gnd.n4353 19.3944
R8691 gnd.n4353 gnd.n4352 19.3944
R8692 gnd.n4352 gnd.n311 19.3944
R8693 gnd.n7194 gnd.n311 19.3944
R8694 gnd.n7194 gnd.n309 19.3944
R8695 gnd.n7198 gnd.n309 19.3944
R8696 gnd.n7198 gnd.n69 19.3944
R8697 gnd.n7574 gnd.n69 19.3944
R8698 gnd.n7574 gnd.n7573 19.3944
R8699 gnd.n7573 gnd.n7572 19.3944
R8700 gnd.n7572 gnd.n73 19.3944
R8701 gnd.n7568 gnd.n73 19.3944
R8702 gnd.n7568 gnd.n7567 19.3944
R8703 gnd.n7567 gnd.n7566 19.3944
R8704 gnd.n7566 gnd.n78 19.3944
R8705 gnd.n7562 gnd.n78 19.3944
R8706 gnd.n7562 gnd.n7561 19.3944
R8707 gnd.n7561 gnd.n7560 19.3944
R8708 gnd.n7560 gnd.n83 19.3944
R8709 gnd.n7556 gnd.n83 19.3944
R8710 gnd.n7556 gnd.n7555 19.3944
R8711 gnd.n7555 gnd.n7554 19.3944
R8712 gnd.n7554 gnd.n88 19.3944
R8713 gnd.n7550 gnd.n88 19.3944
R8714 gnd.n7550 gnd.n7549 19.3944
R8715 gnd.n7549 gnd.n7548 19.3944
R8716 gnd.n7548 gnd.n93 19.3944
R8717 gnd.n7544 gnd.n93 19.3944
R8718 gnd.n7544 gnd.n7543 19.3944
R8719 gnd.n7543 gnd.n7542 19.3944
R8720 gnd.n7542 gnd.n98 19.3944
R8721 gnd.n7538 gnd.n98 19.3944
R8722 gnd.n7538 gnd.n7537 19.3944
R8723 gnd.n7537 gnd.n7536 19.3944
R8724 gnd.n7435 gnd.n7434 19.3944
R8725 gnd.n7434 gnd.n7433 19.3944
R8726 gnd.n7433 gnd.n7375 19.3944
R8727 gnd.n7429 gnd.n7375 19.3944
R8728 gnd.n7429 gnd.n7428 19.3944
R8729 gnd.n7428 gnd.n7427 19.3944
R8730 gnd.n7427 gnd.n7383 19.3944
R8731 gnd.n7423 gnd.n7383 19.3944
R8732 gnd.n7423 gnd.n7422 19.3944
R8733 gnd.n7422 gnd.n7421 19.3944
R8734 gnd.n7421 gnd.n7391 19.3944
R8735 gnd.n7417 gnd.n7391 19.3944
R8736 gnd.n7417 gnd.n7416 19.3944
R8737 gnd.n7416 gnd.n7415 19.3944
R8738 gnd.n7415 gnd.n7399 19.3944
R8739 gnd.n7411 gnd.n7399 19.3944
R8740 gnd.n1726 gnd.n1722 19.3944
R8741 gnd.n1729 gnd.n1726 19.3944
R8742 gnd.n1732 gnd.n1729 19.3944
R8743 gnd.n1732 gnd.n1715 19.3944
R8744 gnd.n1745 gnd.n1715 19.3944
R8745 gnd.n1748 gnd.n1745 19.3944
R8746 gnd.n1751 gnd.n1748 19.3944
R8747 gnd.n1751 gnd.n1708 19.3944
R8748 gnd.n1764 gnd.n1708 19.3944
R8749 gnd.n1767 gnd.n1764 19.3944
R8750 gnd.n1770 gnd.n1767 19.3944
R8751 gnd.n1770 gnd.n1701 19.3944
R8752 gnd.n1782 gnd.n1701 19.3944
R8753 gnd.n1785 gnd.n1782 19.3944
R8754 gnd.n1785 gnd.n1693 19.3944
R8755 gnd.n1798 gnd.n1693 19.3944
R8756 gnd.n4420 gnd.n1502 19.3944
R8757 gnd.n4416 gnd.n1502 19.3944
R8758 gnd.n4416 gnd.n4415 19.3944
R8759 gnd.n4415 gnd.n4414 19.3944
R8760 gnd.n4414 gnd.n1508 19.3944
R8761 gnd.n4410 gnd.n1508 19.3944
R8762 gnd.n4410 gnd.n4409 19.3944
R8763 gnd.n4409 gnd.n4408 19.3944
R8764 gnd.n4408 gnd.n1513 19.3944
R8765 gnd.n4404 gnd.n1513 19.3944
R8766 gnd.n4404 gnd.n4403 19.3944
R8767 gnd.n4403 gnd.n4402 19.3944
R8768 gnd.n4402 gnd.n1518 19.3944
R8769 gnd.n4398 gnd.n1518 19.3944
R8770 gnd.n4398 gnd.n4397 19.3944
R8771 gnd.n4397 gnd.n4396 19.3944
R8772 gnd.n4396 gnd.n1523 19.3944
R8773 gnd.n4392 gnd.n1523 19.3944
R8774 gnd.n4392 gnd.n4391 19.3944
R8775 gnd.n4391 gnd.n4390 19.3944
R8776 gnd.n4390 gnd.n283 19.3944
R8777 gnd.n7290 gnd.n283 19.3944
R8778 gnd.n7290 gnd.n284 19.3944
R8779 gnd.n7286 gnd.n284 19.3944
R8780 gnd.n7286 gnd.n7285 19.3944
R8781 gnd.n7285 gnd.n7284 19.3944
R8782 gnd.n7284 gnd.n290 19.3944
R8783 gnd.n7279 gnd.n290 19.3944
R8784 gnd.n7279 gnd.n7278 19.3944
R8785 gnd.n7278 gnd.n261 19.3944
R8786 gnd.n7301 gnd.n261 19.3944
R8787 gnd.n7301 gnd.n259 19.3944
R8788 gnd.n7305 gnd.n259 19.3944
R8789 gnd.n7305 gnd.n245 19.3944
R8790 gnd.n7317 gnd.n245 19.3944
R8791 gnd.n7317 gnd.n243 19.3944
R8792 gnd.n7321 gnd.n243 19.3944
R8793 gnd.n7321 gnd.n230 19.3944
R8794 gnd.n7333 gnd.n230 19.3944
R8795 gnd.n7333 gnd.n228 19.3944
R8796 gnd.n7337 gnd.n228 19.3944
R8797 gnd.n7337 gnd.n215 19.3944
R8798 gnd.n7349 gnd.n215 19.3944
R8799 gnd.n7349 gnd.n213 19.3944
R8800 gnd.n7353 gnd.n213 19.3944
R8801 gnd.n7353 gnd.n200 19.3944
R8802 gnd.n7365 gnd.n200 19.3944
R8803 gnd.n7365 gnd.n197 19.3944
R8804 gnd.n7444 gnd.n197 19.3944
R8805 gnd.n7444 gnd.n198 19.3944
R8806 gnd.n7440 gnd.n198 19.3944
R8807 gnd.n7440 gnd.n7439 19.3944
R8808 gnd.n7439 gnd.n7438 19.3944
R8809 gnd.n2250 gnd.n1276 19.3944
R8810 gnd.n2250 gnd.n2200 19.3944
R8811 gnd.n3186 gnd.n2200 19.3944
R8812 gnd.n3186 gnd.n3185 19.3944
R8813 gnd.n3185 gnd.n2203 19.3944
R8814 gnd.n3178 gnd.n2203 19.3944
R8815 gnd.n3178 gnd.n3177 19.3944
R8816 gnd.n3177 gnd.n2212 19.3944
R8817 gnd.n3170 gnd.n2212 19.3944
R8818 gnd.n3170 gnd.n3169 19.3944
R8819 gnd.n3169 gnd.n2220 19.3944
R8820 gnd.n3162 gnd.n2220 19.3944
R8821 gnd.n3162 gnd.n3161 19.3944
R8822 gnd.n3161 gnd.n2230 19.3944
R8823 gnd.n3154 gnd.n2230 19.3944
R8824 gnd.n3154 gnd.n3153 19.3944
R8825 gnd.n6957 gnd.n452 19.3944
R8826 gnd.n6963 gnd.n452 19.3944
R8827 gnd.n6963 gnd.n450 19.3944
R8828 gnd.n6967 gnd.n450 19.3944
R8829 gnd.n6967 gnd.n446 19.3944
R8830 gnd.n6973 gnd.n446 19.3944
R8831 gnd.n6973 gnd.n444 19.3944
R8832 gnd.n6977 gnd.n444 19.3944
R8833 gnd.n6977 gnd.n440 19.3944
R8834 gnd.n6983 gnd.n440 19.3944
R8835 gnd.n6983 gnd.n438 19.3944
R8836 gnd.n6987 gnd.n438 19.3944
R8837 gnd.n6987 gnd.n434 19.3944
R8838 gnd.n6993 gnd.n434 19.3944
R8839 gnd.n6993 gnd.n432 19.3944
R8840 gnd.n6997 gnd.n432 19.3944
R8841 gnd.n6997 gnd.n428 19.3944
R8842 gnd.n7003 gnd.n428 19.3944
R8843 gnd.n7003 gnd.n426 19.3944
R8844 gnd.n7007 gnd.n426 19.3944
R8845 gnd.n7007 gnd.n422 19.3944
R8846 gnd.n7013 gnd.n422 19.3944
R8847 gnd.n7013 gnd.n420 19.3944
R8848 gnd.n7017 gnd.n420 19.3944
R8849 gnd.n7017 gnd.n416 19.3944
R8850 gnd.n7023 gnd.n416 19.3944
R8851 gnd.n7023 gnd.n414 19.3944
R8852 gnd.n7027 gnd.n414 19.3944
R8853 gnd.n7027 gnd.n410 19.3944
R8854 gnd.n7033 gnd.n410 19.3944
R8855 gnd.n7033 gnd.n408 19.3944
R8856 gnd.n7037 gnd.n408 19.3944
R8857 gnd.n7037 gnd.n404 19.3944
R8858 gnd.n7043 gnd.n404 19.3944
R8859 gnd.n7043 gnd.n402 19.3944
R8860 gnd.n7047 gnd.n402 19.3944
R8861 gnd.n7047 gnd.n398 19.3944
R8862 gnd.n7053 gnd.n398 19.3944
R8863 gnd.n7053 gnd.n396 19.3944
R8864 gnd.n7057 gnd.n396 19.3944
R8865 gnd.n7057 gnd.n392 19.3944
R8866 gnd.n7063 gnd.n392 19.3944
R8867 gnd.n7063 gnd.n390 19.3944
R8868 gnd.n7067 gnd.n390 19.3944
R8869 gnd.n7067 gnd.n386 19.3944
R8870 gnd.n7073 gnd.n386 19.3944
R8871 gnd.n7073 gnd.n384 19.3944
R8872 gnd.n7077 gnd.n384 19.3944
R8873 gnd.n7077 gnd.n380 19.3944
R8874 gnd.n7083 gnd.n380 19.3944
R8875 gnd.n7083 gnd.n378 19.3944
R8876 gnd.n7087 gnd.n378 19.3944
R8877 gnd.n7087 gnd.n374 19.3944
R8878 gnd.n7093 gnd.n374 19.3944
R8879 gnd.n7093 gnd.n372 19.3944
R8880 gnd.n7097 gnd.n372 19.3944
R8881 gnd.n7097 gnd.n368 19.3944
R8882 gnd.n7103 gnd.n368 19.3944
R8883 gnd.n7103 gnd.n366 19.3944
R8884 gnd.n7107 gnd.n366 19.3944
R8885 gnd.n7107 gnd.n362 19.3944
R8886 gnd.n7113 gnd.n362 19.3944
R8887 gnd.n7113 gnd.n360 19.3944
R8888 gnd.n7117 gnd.n360 19.3944
R8889 gnd.n7117 gnd.n356 19.3944
R8890 gnd.n7123 gnd.n356 19.3944
R8891 gnd.n7123 gnd.n354 19.3944
R8892 gnd.n7127 gnd.n354 19.3944
R8893 gnd.n7127 gnd.n350 19.3944
R8894 gnd.n7133 gnd.n350 19.3944
R8895 gnd.n7133 gnd.n348 19.3944
R8896 gnd.n7137 gnd.n348 19.3944
R8897 gnd.n7137 gnd.n344 19.3944
R8898 gnd.n7143 gnd.n344 19.3944
R8899 gnd.n7143 gnd.n342 19.3944
R8900 gnd.n7147 gnd.n342 19.3944
R8901 gnd.n7147 gnd.n338 19.3944
R8902 gnd.n7153 gnd.n338 19.3944
R8903 gnd.n7153 gnd.n336 19.3944
R8904 gnd.n7157 gnd.n336 19.3944
R8905 gnd.n7157 gnd.n332 19.3944
R8906 gnd.n7164 gnd.n332 19.3944
R8907 gnd.n7164 gnd.n330 19.3944
R8908 gnd.n7169 gnd.n330 19.3944
R8909 gnd.n6502 gnd.n725 19.3944
R8910 gnd.n6506 gnd.n725 19.3944
R8911 gnd.n6506 gnd.n721 19.3944
R8912 gnd.n6512 gnd.n721 19.3944
R8913 gnd.n6512 gnd.n719 19.3944
R8914 gnd.n6516 gnd.n719 19.3944
R8915 gnd.n6516 gnd.n715 19.3944
R8916 gnd.n6522 gnd.n715 19.3944
R8917 gnd.n6522 gnd.n713 19.3944
R8918 gnd.n6526 gnd.n713 19.3944
R8919 gnd.n6526 gnd.n709 19.3944
R8920 gnd.n6532 gnd.n709 19.3944
R8921 gnd.n6532 gnd.n707 19.3944
R8922 gnd.n6536 gnd.n707 19.3944
R8923 gnd.n6536 gnd.n703 19.3944
R8924 gnd.n6542 gnd.n703 19.3944
R8925 gnd.n6542 gnd.n701 19.3944
R8926 gnd.n6546 gnd.n701 19.3944
R8927 gnd.n6546 gnd.n697 19.3944
R8928 gnd.n6552 gnd.n697 19.3944
R8929 gnd.n6552 gnd.n695 19.3944
R8930 gnd.n6556 gnd.n695 19.3944
R8931 gnd.n6556 gnd.n691 19.3944
R8932 gnd.n6562 gnd.n691 19.3944
R8933 gnd.n6562 gnd.n689 19.3944
R8934 gnd.n6566 gnd.n689 19.3944
R8935 gnd.n6566 gnd.n685 19.3944
R8936 gnd.n6572 gnd.n685 19.3944
R8937 gnd.n6572 gnd.n683 19.3944
R8938 gnd.n6576 gnd.n683 19.3944
R8939 gnd.n6576 gnd.n679 19.3944
R8940 gnd.n6582 gnd.n679 19.3944
R8941 gnd.n6582 gnd.n677 19.3944
R8942 gnd.n6586 gnd.n677 19.3944
R8943 gnd.n6586 gnd.n673 19.3944
R8944 gnd.n6592 gnd.n673 19.3944
R8945 gnd.n6592 gnd.n671 19.3944
R8946 gnd.n6596 gnd.n671 19.3944
R8947 gnd.n6596 gnd.n667 19.3944
R8948 gnd.n6602 gnd.n667 19.3944
R8949 gnd.n6602 gnd.n665 19.3944
R8950 gnd.n6606 gnd.n665 19.3944
R8951 gnd.n6606 gnd.n661 19.3944
R8952 gnd.n6612 gnd.n661 19.3944
R8953 gnd.n6612 gnd.n659 19.3944
R8954 gnd.n6616 gnd.n659 19.3944
R8955 gnd.n6616 gnd.n655 19.3944
R8956 gnd.n6622 gnd.n655 19.3944
R8957 gnd.n6622 gnd.n653 19.3944
R8958 gnd.n6626 gnd.n653 19.3944
R8959 gnd.n6626 gnd.n649 19.3944
R8960 gnd.n6632 gnd.n649 19.3944
R8961 gnd.n6632 gnd.n647 19.3944
R8962 gnd.n6636 gnd.n647 19.3944
R8963 gnd.n6636 gnd.n643 19.3944
R8964 gnd.n6642 gnd.n643 19.3944
R8965 gnd.n6642 gnd.n641 19.3944
R8966 gnd.n6646 gnd.n641 19.3944
R8967 gnd.n6646 gnd.n637 19.3944
R8968 gnd.n6652 gnd.n637 19.3944
R8969 gnd.n6652 gnd.n635 19.3944
R8970 gnd.n6656 gnd.n635 19.3944
R8971 gnd.n6656 gnd.n631 19.3944
R8972 gnd.n6662 gnd.n631 19.3944
R8973 gnd.n6662 gnd.n629 19.3944
R8974 gnd.n6666 gnd.n629 19.3944
R8975 gnd.n6666 gnd.n625 19.3944
R8976 gnd.n6672 gnd.n625 19.3944
R8977 gnd.n6672 gnd.n623 19.3944
R8978 gnd.n6676 gnd.n623 19.3944
R8979 gnd.n6676 gnd.n619 19.3944
R8980 gnd.n6682 gnd.n619 19.3944
R8981 gnd.n6682 gnd.n617 19.3944
R8982 gnd.n6686 gnd.n617 19.3944
R8983 gnd.n6686 gnd.n613 19.3944
R8984 gnd.n6692 gnd.n613 19.3944
R8985 gnd.n6692 gnd.n611 19.3944
R8986 gnd.n6696 gnd.n611 19.3944
R8987 gnd.n6696 gnd.n607 19.3944
R8988 gnd.n6702 gnd.n607 19.3944
R8989 gnd.n6702 gnd.n605 19.3944
R8990 gnd.n6706 gnd.n605 19.3944
R8991 gnd.n6706 gnd.n601 19.3944
R8992 gnd.n6712 gnd.n601 19.3944
R8993 gnd.n6712 gnd.n599 19.3944
R8994 gnd.n6716 gnd.n599 19.3944
R8995 gnd.n6716 gnd.n595 19.3944
R8996 gnd.n6722 gnd.n595 19.3944
R8997 gnd.n6722 gnd.n593 19.3944
R8998 gnd.n6726 gnd.n593 19.3944
R8999 gnd.n6726 gnd.n589 19.3944
R9000 gnd.n6732 gnd.n589 19.3944
R9001 gnd.n6732 gnd.n587 19.3944
R9002 gnd.n6736 gnd.n587 19.3944
R9003 gnd.n6736 gnd.n583 19.3944
R9004 gnd.n6742 gnd.n583 19.3944
R9005 gnd.n6742 gnd.n581 19.3944
R9006 gnd.n6746 gnd.n581 19.3944
R9007 gnd.n6746 gnd.n577 19.3944
R9008 gnd.n6752 gnd.n577 19.3944
R9009 gnd.n6752 gnd.n575 19.3944
R9010 gnd.n6756 gnd.n575 19.3944
R9011 gnd.n6756 gnd.n571 19.3944
R9012 gnd.n6762 gnd.n571 19.3944
R9013 gnd.n6762 gnd.n569 19.3944
R9014 gnd.n6766 gnd.n569 19.3944
R9015 gnd.n6766 gnd.n565 19.3944
R9016 gnd.n6772 gnd.n565 19.3944
R9017 gnd.n6772 gnd.n563 19.3944
R9018 gnd.n6776 gnd.n563 19.3944
R9019 gnd.n6776 gnd.n559 19.3944
R9020 gnd.n6782 gnd.n559 19.3944
R9021 gnd.n6782 gnd.n557 19.3944
R9022 gnd.n6786 gnd.n557 19.3944
R9023 gnd.n6786 gnd.n553 19.3944
R9024 gnd.n6792 gnd.n553 19.3944
R9025 gnd.n6792 gnd.n551 19.3944
R9026 gnd.n6796 gnd.n551 19.3944
R9027 gnd.n6796 gnd.n547 19.3944
R9028 gnd.n6802 gnd.n547 19.3944
R9029 gnd.n6802 gnd.n545 19.3944
R9030 gnd.n6806 gnd.n545 19.3944
R9031 gnd.n6806 gnd.n541 19.3944
R9032 gnd.n6812 gnd.n541 19.3944
R9033 gnd.n6812 gnd.n539 19.3944
R9034 gnd.n6816 gnd.n539 19.3944
R9035 gnd.n6816 gnd.n535 19.3944
R9036 gnd.n6822 gnd.n535 19.3944
R9037 gnd.n6822 gnd.n533 19.3944
R9038 gnd.n6826 gnd.n533 19.3944
R9039 gnd.n6826 gnd.n529 19.3944
R9040 gnd.n6832 gnd.n529 19.3944
R9041 gnd.n6832 gnd.n527 19.3944
R9042 gnd.n6836 gnd.n527 19.3944
R9043 gnd.n6836 gnd.n523 19.3944
R9044 gnd.n6842 gnd.n523 19.3944
R9045 gnd.n6842 gnd.n521 19.3944
R9046 gnd.n6846 gnd.n521 19.3944
R9047 gnd.n6846 gnd.n517 19.3944
R9048 gnd.n6852 gnd.n517 19.3944
R9049 gnd.n6852 gnd.n515 19.3944
R9050 gnd.n6856 gnd.n515 19.3944
R9051 gnd.n6856 gnd.n511 19.3944
R9052 gnd.n6862 gnd.n511 19.3944
R9053 gnd.n6862 gnd.n509 19.3944
R9054 gnd.n6866 gnd.n509 19.3944
R9055 gnd.n6866 gnd.n505 19.3944
R9056 gnd.n6872 gnd.n505 19.3944
R9057 gnd.n6872 gnd.n503 19.3944
R9058 gnd.n6876 gnd.n503 19.3944
R9059 gnd.n6876 gnd.n499 19.3944
R9060 gnd.n6882 gnd.n499 19.3944
R9061 gnd.n6882 gnd.n497 19.3944
R9062 gnd.n6886 gnd.n497 19.3944
R9063 gnd.n6886 gnd.n493 19.3944
R9064 gnd.n6892 gnd.n493 19.3944
R9065 gnd.n6892 gnd.n491 19.3944
R9066 gnd.n6896 gnd.n491 19.3944
R9067 gnd.n6896 gnd.n487 19.3944
R9068 gnd.n6902 gnd.n487 19.3944
R9069 gnd.n6902 gnd.n485 19.3944
R9070 gnd.n6906 gnd.n485 19.3944
R9071 gnd.n6906 gnd.n481 19.3944
R9072 gnd.n6912 gnd.n481 19.3944
R9073 gnd.n6912 gnd.n479 19.3944
R9074 gnd.n6916 gnd.n479 19.3944
R9075 gnd.n6916 gnd.n475 19.3944
R9076 gnd.n6922 gnd.n475 19.3944
R9077 gnd.n6922 gnd.n473 19.3944
R9078 gnd.n6926 gnd.n473 19.3944
R9079 gnd.n6926 gnd.n469 19.3944
R9080 gnd.n6932 gnd.n469 19.3944
R9081 gnd.n6932 gnd.n467 19.3944
R9082 gnd.n6936 gnd.n467 19.3944
R9083 gnd.n6936 gnd.n463 19.3944
R9084 gnd.n6942 gnd.n463 19.3944
R9085 gnd.n6942 gnd.n461 19.3944
R9086 gnd.n6947 gnd.n461 19.3944
R9087 gnd.n6947 gnd.n457 19.3944
R9088 gnd.n6953 gnd.n457 19.3944
R9089 gnd.n6954 gnd.n6953 19.3944
R9090 gnd.n4495 gnd.n4494 19.3944
R9091 gnd.n4494 gnd.n4493 19.3944
R9092 gnd.n4493 gnd.n4492 19.3944
R9093 gnd.n4492 gnd.n4490 19.3944
R9094 gnd.n4490 gnd.n4487 19.3944
R9095 gnd.n4487 gnd.n4486 19.3944
R9096 gnd.n4486 gnd.n4483 19.3944
R9097 gnd.n4483 gnd.n4482 19.3944
R9098 gnd.n4482 gnd.n4479 19.3944
R9099 gnd.n4479 gnd.n4478 19.3944
R9100 gnd.n4478 gnd.n4475 19.3944
R9101 gnd.n4475 gnd.n4474 19.3944
R9102 gnd.n4474 gnd.n4471 19.3944
R9103 gnd.n4471 gnd.n4470 19.3944
R9104 gnd.n4470 gnd.n4467 19.3944
R9105 gnd.n4465 gnd.n4462 19.3944
R9106 gnd.n4462 gnd.n4461 19.3944
R9107 gnd.n4461 gnd.n4458 19.3944
R9108 gnd.n4458 gnd.n4457 19.3944
R9109 gnd.n4457 gnd.n4454 19.3944
R9110 gnd.n4454 gnd.n4453 19.3944
R9111 gnd.n4453 gnd.n4450 19.3944
R9112 gnd.n4450 gnd.n4449 19.3944
R9113 gnd.n4449 gnd.n4446 19.3944
R9114 gnd.n4446 gnd.n4445 19.3944
R9115 gnd.n4445 gnd.n4442 19.3944
R9116 gnd.n4442 gnd.n4441 19.3944
R9117 gnd.n4441 gnd.n4438 19.3944
R9118 gnd.n4438 gnd.n4437 19.3944
R9119 gnd.n4437 gnd.n4434 19.3944
R9120 gnd.n4434 gnd.n4433 19.3944
R9121 gnd.n4433 gnd.n4430 19.3944
R9122 gnd.n4430 gnd.n4429 19.3944
R9123 gnd.n1648 gnd.n1496 19.3944
R9124 gnd.n1678 gnd.n1648 19.3944
R9125 gnd.n1678 gnd.n1677 19.3944
R9126 gnd.n1677 gnd.n1676 19.3944
R9127 gnd.n1676 gnd.n1674 19.3944
R9128 gnd.n1674 gnd.n1673 19.3944
R9129 gnd.n1673 gnd.n1670 19.3944
R9130 gnd.n1670 gnd.n1669 19.3944
R9131 gnd.n1669 gnd.n1668 19.3944
R9132 gnd.n1668 gnd.n1666 19.3944
R9133 gnd.n1666 gnd.n1665 19.3944
R9134 gnd.n1665 gnd.n1663 19.3944
R9135 gnd.n1663 gnd.n1662 19.3944
R9136 gnd.n1662 gnd.n1558 19.3944
R9137 gnd.n4328 gnd.n1558 19.3944
R9138 gnd.n4328 gnd.n1556 19.3944
R9139 gnd.n4332 gnd.n1556 19.3944
R9140 gnd.n4333 gnd.n4332 19.3944
R9141 gnd.n4335 gnd.n4333 19.3944
R9142 gnd.n4335 gnd.n1554 19.3944
R9143 gnd.n4347 gnd.n1554 19.3944
R9144 gnd.n4347 gnd.n4346 19.3944
R9145 gnd.n4346 gnd.n4345 19.3944
R9146 gnd.n4345 gnd.n4344 19.3944
R9147 gnd.n4344 gnd.n299 19.3944
R9148 gnd.n7207 gnd.n299 19.3944
R9149 gnd.n7208 gnd.n7207 19.3944
R9150 gnd.n7269 gnd.n7208 19.3944
R9151 gnd.n7269 gnd.n7268 19.3944
R9152 gnd.n7268 gnd.n7267 19.3944
R9153 gnd.n7267 gnd.n7263 19.3944
R9154 gnd.n7263 gnd.n7262 19.3944
R9155 gnd.n7262 gnd.n7259 19.3944
R9156 gnd.n7259 gnd.n7258 19.3944
R9157 gnd.n7258 gnd.n7256 19.3944
R9158 gnd.n7256 gnd.n7255 19.3944
R9159 gnd.n7255 gnd.n7253 19.3944
R9160 gnd.n7253 gnd.n7252 19.3944
R9161 gnd.n7252 gnd.n7250 19.3944
R9162 gnd.n7250 gnd.n7249 19.3944
R9163 gnd.n7249 gnd.n7247 19.3944
R9164 gnd.n7247 gnd.n7246 19.3944
R9165 gnd.n7246 gnd.n7244 19.3944
R9166 gnd.n7244 gnd.n7243 19.3944
R9167 gnd.n7243 gnd.n7241 19.3944
R9168 gnd.n7241 gnd.n7240 19.3944
R9169 gnd.n7240 gnd.n7238 19.3944
R9170 gnd.n7238 gnd.n7237 19.3944
R9171 gnd.n7237 gnd.n7235 19.3944
R9172 gnd.n7235 gnd.n7234 19.3944
R9173 gnd.n7234 gnd.n182 19.3944
R9174 gnd.n7457 gnd.n182 19.3944
R9175 gnd.n7458 gnd.n7457 19.3944
R9176 gnd.n7496 gnd.n143 19.3944
R9177 gnd.n7491 gnd.n143 19.3944
R9178 gnd.n7491 gnd.n7490 19.3944
R9179 gnd.n7490 gnd.n7489 19.3944
R9180 gnd.n7489 gnd.n150 19.3944
R9181 gnd.n7484 gnd.n150 19.3944
R9182 gnd.n7484 gnd.n7483 19.3944
R9183 gnd.n7483 gnd.n7482 19.3944
R9184 gnd.n7482 gnd.n157 19.3944
R9185 gnd.n7477 gnd.n157 19.3944
R9186 gnd.n7477 gnd.n7476 19.3944
R9187 gnd.n7476 gnd.n7475 19.3944
R9188 gnd.n7475 gnd.n164 19.3944
R9189 gnd.n7470 gnd.n164 19.3944
R9190 gnd.n7470 gnd.n7469 19.3944
R9191 gnd.n7469 gnd.n7468 19.3944
R9192 gnd.n7468 gnd.n171 19.3944
R9193 gnd.n7463 gnd.n171 19.3944
R9194 gnd.n7529 gnd.n7528 19.3944
R9195 gnd.n7528 gnd.n7527 19.3944
R9196 gnd.n7527 gnd.n115 19.3944
R9197 gnd.n7522 gnd.n115 19.3944
R9198 gnd.n7522 gnd.n7521 19.3944
R9199 gnd.n7521 gnd.n7520 19.3944
R9200 gnd.n7520 gnd.n122 19.3944
R9201 gnd.n7515 gnd.n122 19.3944
R9202 gnd.n7515 gnd.n7514 19.3944
R9203 gnd.n7514 gnd.n7513 19.3944
R9204 gnd.n7513 gnd.n129 19.3944
R9205 gnd.n7508 gnd.n129 19.3944
R9206 gnd.n7508 gnd.n7507 19.3944
R9207 gnd.n7507 gnd.n7506 19.3944
R9208 gnd.n7506 gnd.n136 19.3944
R9209 gnd.n7501 gnd.n136 19.3944
R9210 gnd.n7501 gnd.n7500 19.3944
R9211 gnd.n1645 gnd.n1642 19.3944
R9212 gnd.n1645 gnd.n1623 19.3944
R9213 gnd.n4250 gnd.n1623 19.3944
R9214 gnd.n4250 gnd.n1621 19.3944
R9215 gnd.n4256 gnd.n1621 19.3944
R9216 gnd.n4256 gnd.n4255 19.3944
R9217 gnd.n4255 gnd.n1595 19.3944
R9218 gnd.n4281 gnd.n1595 19.3944
R9219 gnd.n4281 gnd.n1593 19.3944
R9220 gnd.n4287 gnd.n1593 19.3944
R9221 gnd.n4287 gnd.n4286 19.3944
R9222 gnd.n4286 gnd.n1568 19.3944
R9223 gnd.n4318 gnd.n1568 19.3944
R9224 gnd.n4318 gnd.n1566 19.3944
R9225 gnd.n4324 gnd.n1566 19.3944
R9226 gnd.n4324 gnd.n4323 19.3944
R9227 gnd.n4323 gnd.n1533 19.3944
R9228 gnd.n4381 gnd.n1533 19.3944
R9229 gnd.n4381 gnd.n1531 19.3944
R9230 gnd.n4385 gnd.n1531 19.3944
R9231 gnd.n4385 gnd.n275 19.3944
R9232 gnd.n7294 gnd.n275 19.3944
R9233 gnd.n274 gnd.n273 19.3944
R9234 gnd.n306 gnd.n273 19.3944
R9235 gnd.n7203 gnd.n7202 19.3944
R9236 gnd.n7274 gnd.n7273 19.3944
R9237 gnd.n7297 gnd.n267 19.3944
R9238 gnd.n7297 gnd.n254 19.3944
R9239 gnd.n7309 gnd.n254 19.3944
R9240 gnd.n7309 gnd.n252 19.3944
R9241 gnd.n7313 gnd.n252 19.3944
R9242 gnd.n7313 gnd.n236 19.3944
R9243 gnd.n7325 gnd.n236 19.3944
R9244 gnd.n7325 gnd.n234 19.3944
R9245 gnd.n7329 gnd.n234 19.3944
R9246 gnd.n7329 gnd.n223 19.3944
R9247 gnd.n7341 gnd.n223 19.3944
R9248 gnd.n7341 gnd.n221 19.3944
R9249 gnd.n7345 gnd.n221 19.3944
R9250 gnd.n7345 gnd.n206 19.3944
R9251 gnd.n7357 gnd.n206 19.3944
R9252 gnd.n7357 gnd.n204 19.3944
R9253 gnd.n7361 gnd.n204 19.3944
R9254 gnd.n7361 gnd.n191 19.3944
R9255 gnd.n7448 gnd.n191 19.3944
R9256 gnd.n7448 gnd.n189 19.3944
R9257 gnd.n7452 gnd.n189 19.3944
R9258 gnd.n7452 gnd.n110 19.3944
R9259 gnd.n7532 gnd.n110 19.3944
R9260 gnd.n2410 gnd.n2406 19.3944
R9261 gnd.n2652 gnd.n2406 19.3944
R9262 gnd.n2652 gnd.n2407 19.3944
R9263 gnd.n2604 gnd.n2603 19.3944
R9264 gnd.n2612 gnd.n2611 19.3944
R9265 gnd.n2608 gnd.n2607 19.3944
R9266 gnd.n2656 gnd.n2381 19.3944
R9267 gnd.n2399 gnd.n2382 19.3944
R9268 gnd.n2399 gnd.n2384 19.3944
R9269 gnd.n2395 gnd.n2384 19.3944
R9270 gnd.n2395 gnd.n2394 19.3944
R9271 gnd.n2394 gnd.n2393 19.3944
R9272 gnd.n2393 gnd.n2391 19.3944
R9273 gnd.n2391 gnd.n2353 19.3944
R9274 gnd.n2353 gnd.n2351 19.3944
R9275 gnd.n2728 gnd.n2351 19.3944
R9276 gnd.n2728 gnd.n2349 19.3944
R9277 gnd.n2732 gnd.n2349 19.3944
R9278 gnd.n2732 gnd.n2347 19.3944
R9279 gnd.n2736 gnd.n2347 19.3944
R9280 gnd.n2736 gnd.n2345 19.3944
R9281 gnd.n2773 gnd.n2345 19.3944
R9282 gnd.n2773 gnd.n2772 19.3944
R9283 gnd.n2772 gnd.n2771 19.3944
R9284 gnd.n2771 gnd.n2742 19.3944
R9285 gnd.n2767 gnd.n2742 19.3944
R9286 gnd.n2767 gnd.n2766 19.3944
R9287 gnd.n2766 gnd.n2765 19.3944
R9288 gnd.n2765 gnd.n2748 19.3944
R9289 gnd.n2761 gnd.n2748 19.3944
R9290 gnd.n2761 gnd.n2760 19.3944
R9291 gnd.n2760 gnd.n2759 19.3944
R9292 gnd.n2759 gnd.n2755 19.3944
R9293 gnd.n2755 gnd.n2173 19.3944
R9294 gnd.n3204 gnd.n2173 19.3944
R9295 gnd.n3204 gnd.n2171 19.3944
R9296 gnd.n3208 gnd.n2171 19.3944
R9297 gnd.n3208 gnd.n2161 19.3944
R9298 gnd.n3220 gnd.n2161 19.3944
R9299 gnd.n3220 gnd.n2159 19.3944
R9300 gnd.n3224 gnd.n2159 19.3944
R9301 gnd.n3224 gnd.n2148 19.3944
R9302 gnd.n3236 gnd.n2148 19.3944
R9303 gnd.n3236 gnd.n2146 19.3944
R9304 gnd.n3240 gnd.n2146 19.3944
R9305 gnd.n3240 gnd.n2135 19.3944
R9306 gnd.n3252 gnd.n2135 19.3944
R9307 gnd.n3252 gnd.n2133 19.3944
R9308 gnd.n3256 gnd.n2133 19.3944
R9309 gnd.n3256 gnd.n2120 19.3944
R9310 gnd.n3268 gnd.n2120 19.3944
R9311 gnd.n3268 gnd.n2118 19.3944
R9312 gnd.n3272 gnd.n2118 19.3944
R9313 gnd.n3272 gnd.n2108 19.3944
R9314 gnd.n3284 gnd.n2108 19.3944
R9315 gnd.n3284 gnd.n2106 19.3944
R9316 gnd.n3290 gnd.n2106 19.3944
R9317 gnd.n3290 gnd.n3289 19.3944
R9318 gnd.n3289 gnd.n2080 19.3944
R9319 gnd.n3900 gnd.n2080 19.3944
R9320 gnd.n3900 gnd.n2078 19.3944
R9321 gnd.n3904 gnd.n2078 19.3944
R9322 gnd.n3904 gnd.n2065 19.3944
R9323 gnd.n3916 gnd.n2065 19.3944
R9324 gnd.n3916 gnd.n2063 19.3944
R9325 gnd.n3920 gnd.n2063 19.3944
R9326 gnd.n3920 gnd.n2050 19.3944
R9327 gnd.n3932 gnd.n2050 19.3944
R9328 gnd.n3932 gnd.n2048 19.3944
R9329 gnd.n3936 gnd.n2048 19.3944
R9330 gnd.n3936 gnd.n2035 19.3944
R9331 gnd.n3948 gnd.n2035 19.3944
R9332 gnd.n3948 gnd.n2033 19.3944
R9333 gnd.n3952 gnd.n2033 19.3944
R9334 gnd.n3952 gnd.n2021 19.3944
R9335 gnd.n3964 gnd.n2021 19.3944
R9336 gnd.n3964 gnd.n2019 19.3944
R9337 gnd.n3968 gnd.n2019 19.3944
R9338 gnd.n3968 gnd.n2006 19.3944
R9339 gnd.n3980 gnd.n2006 19.3944
R9340 gnd.n3980 gnd.n2004 19.3944
R9341 gnd.n3984 gnd.n2004 19.3944
R9342 gnd.n3984 gnd.n1991 19.3944
R9343 gnd.n3996 gnd.n1991 19.3944
R9344 gnd.n3996 gnd.n1989 19.3944
R9345 gnd.n4000 gnd.n1989 19.3944
R9346 gnd.n4000 gnd.n1976 19.3944
R9347 gnd.n4012 gnd.n1976 19.3944
R9348 gnd.n4012 gnd.n1974 19.3944
R9349 gnd.n4016 gnd.n1974 19.3944
R9350 gnd.n4016 gnd.n1962 19.3944
R9351 gnd.n4028 gnd.n1962 19.3944
R9352 gnd.n4028 gnd.n1960 19.3944
R9353 gnd.n4032 gnd.n1960 19.3944
R9354 gnd.n4032 gnd.n1947 19.3944
R9355 gnd.n4044 gnd.n1947 19.3944
R9356 gnd.n4044 gnd.n1945 19.3944
R9357 gnd.n4048 gnd.n1945 19.3944
R9358 gnd.n4048 gnd.n1934 19.3944
R9359 gnd.n4060 gnd.n1934 19.3944
R9360 gnd.n4060 gnd.n1932 19.3944
R9361 gnd.n4064 gnd.n1932 19.3944
R9362 gnd.n4064 gnd.n1922 19.3944
R9363 gnd.n4076 gnd.n1922 19.3944
R9364 gnd.n4076 gnd.n1920 19.3944
R9365 gnd.n4080 gnd.n1920 19.3944
R9366 gnd.n4080 gnd.n1909 19.3944
R9367 gnd.n4092 gnd.n1909 19.3944
R9368 gnd.n4092 gnd.n1907 19.3944
R9369 gnd.n4096 gnd.n1907 19.3944
R9370 gnd.n4096 gnd.n1895 19.3944
R9371 gnd.n4108 gnd.n1895 19.3944
R9372 gnd.n4108 gnd.n1893 19.3944
R9373 gnd.n4112 gnd.n1893 19.3944
R9374 gnd.n4112 gnd.n1882 19.3944
R9375 gnd.n4124 gnd.n1882 19.3944
R9376 gnd.n4124 gnd.n1880 19.3944
R9377 gnd.n4128 gnd.n1880 19.3944
R9378 gnd.n4128 gnd.n1869 19.3944
R9379 gnd.n4140 gnd.n1869 19.3944
R9380 gnd.n4140 gnd.n1867 19.3944
R9381 gnd.n4144 gnd.n1867 19.3944
R9382 gnd.n4144 gnd.n1856 19.3944
R9383 gnd.n4156 gnd.n1856 19.3944
R9384 gnd.n4156 gnd.n1854 19.3944
R9385 gnd.n4160 gnd.n1854 19.3944
R9386 gnd.n4160 gnd.n1842 19.3944
R9387 gnd.n4172 gnd.n1842 19.3944
R9388 gnd.n4172 gnd.n1840 19.3944
R9389 gnd.n4176 gnd.n1840 19.3944
R9390 gnd.n4176 gnd.n1829 19.3944
R9391 gnd.n4190 gnd.n1829 19.3944
R9392 gnd.n4190 gnd.n1827 19.3944
R9393 gnd.n4197 gnd.n1827 19.3944
R9394 gnd.n4197 gnd.n4196 19.3944
R9395 gnd.n4196 gnd.n1411 19.3944
R9396 gnd.n4504 gnd.n1411 19.3944
R9397 gnd.n4504 gnd.n4503 19.3944
R9398 gnd.n4503 gnd.n4502 19.3944
R9399 gnd.n4502 gnd.n1415 19.3944
R9400 gnd.n1635 gnd.n1415 19.3944
R9401 gnd.n1639 gnd.n1635 19.3944
R9402 gnd.n1639 gnd.n1633 19.3944
R9403 gnd.n4239 gnd.n1633 19.3944
R9404 gnd.n4239 gnd.n1631 19.3944
R9405 gnd.n4245 gnd.n1631 19.3944
R9406 gnd.n4245 gnd.n4244 19.3944
R9407 gnd.n4244 gnd.n1606 19.3944
R9408 gnd.n4270 gnd.n1606 19.3944
R9409 gnd.n4270 gnd.n1604 19.3944
R9410 gnd.n4276 gnd.n1604 19.3944
R9411 gnd.n4276 gnd.n4275 19.3944
R9412 gnd.n4275 gnd.n1578 19.3944
R9413 gnd.n4306 gnd.n1578 19.3944
R9414 gnd.n4306 gnd.n1576 19.3944
R9415 gnd.n4312 gnd.n1576 19.3944
R9416 gnd.n4312 gnd.n4311 19.3944
R9417 gnd.n4311 gnd.n1544 19.3944
R9418 gnd.n4364 gnd.n1544 19.3944
R9419 gnd.n4364 gnd.n1542 19.3944
R9420 gnd.n4376 gnd.n1542 19.3944
R9421 gnd.n4376 gnd.n4375 19.3944
R9422 gnd.n4375 gnd.n4374 19.3944
R9423 gnd.n4374 gnd.n4371 19.3944
R9424 gnd.n7189 gnd.n317 19.3944
R9425 gnd.n7187 gnd.n7186 19.3944
R9426 gnd.n7183 gnd.n7182 19.3944
R9427 gnd.n7180 gnd.n323 19.3944
R9428 gnd.n7176 gnd.n7175 19.3944
R9429 gnd.n7175 gnd.n7174 19.3944
R9430 gnd.n7174 gnd.n328 19.3944
R9431 gnd.n4902 gnd.n4901 19.3944
R9432 gnd.n4901 gnd.n4900 19.3944
R9433 gnd.n4900 gnd.n4899 19.3944
R9434 gnd.n4899 gnd.n4897 19.3944
R9435 gnd.n4897 gnd.n4894 19.3944
R9436 gnd.n4894 gnd.n4893 19.3944
R9437 gnd.n4893 gnd.n4890 19.3944
R9438 gnd.n4890 gnd.n4889 19.3944
R9439 gnd.n4889 gnd.n4886 19.3944
R9440 gnd.n4886 gnd.n4885 19.3944
R9441 gnd.n4885 gnd.n4882 19.3944
R9442 gnd.n4882 gnd.n4881 19.3944
R9443 gnd.n4881 gnd.n4878 19.3944
R9444 gnd.n4878 gnd.n4877 19.3944
R9445 gnd.n4877 gnd.n4874 19.3944
R9446 gnd.n4874 gnd.n4873 19.3944
R9447 gnd.n4873 gnd.n4870 19.3944
R9448 gnd.n4868 gnd.n4865 19.3944
R9449 gnd.n4865 gnd.n4864 19.3944
R9450 gnd.n4864 gnd.n4861 19.3944
R9451 gnd.n4861 gnd.n4860 19.3944
R9452 gnd.n4860 gnd.n4857 19.3944
R9453 gnd.n4857 gnd.n4856 19.3944
R9454 gnd.n4856 gnd.n4853 19.3944
R9455 gnd.n4853 gnd.n4852 19.3944
R9456 gnd.n4852 gnd.n4849 19.3944
R9457 gnd.n4849 gnd.n4848 19.3944
R9458 gnd.n4848 gnd.n4845 19.3944
R9459 gnd.n4845 gnd.n4844 19.3944
R9460 gnd.n4844 gnd.n4841 19.3944
R9461 gnd.n4841 gnd.n4840 19.3944
R9462 gnd.n4840 gnd.n4837 19.3944
R9463 gnd.n4837 gnd.n4836 19.3944
R9464 gnd.n4836 gnd.n4833 19.3944
R9465 gnd.n4833 gnd.n4832 19.3944
R9466 gnd.n4825 gnd.n4824 19.3944
R9467 gnd.n4824 gnd.n1010 19.3944
R9468 gnd.n4820 gnd.n1010 19.3944
R9469 gnd.n4820 gnd.n1012 19.3944
R9470 gnd.n2430 gnd.n1012 19.3944
R9471 gnd.n2432 gnd.n2430 19.3944
R9472 gnd.n2432 gnd.n2428 19.3944
R9473 gnd.n2437 gnd.n2428 19.3944
R9474 gnd.n2438 gnd.n2437 19.3944
R9475 gnd.n2440 gnd.n2438 19.3944
R9476 gnd.n2440 gnd.n2426 19.3944
R9477 gnd.n2445 gnd.n2426 19.3944
R9478 gnd.n2446 gnd.n2445 19.3944
R9479 gnd.n2448 gnd.n2446 19.3944
R9480 gnd.n2448 gnd.n2424 19.3944
R9481 gnd.n2453 gnd.n2424 19.3944
R9482 gnd.n2454 gnd.n2453 19.3944
R9483 gnd.n2456 gnd.n2454 19.3944
R9484 gnd.n2456 gnd.n2422 19.3944
R9485 gnd.n2594 gnd.n2422 19.3944
R9486 gnd.n2595 gnd.n2594 19.3944
R9487 gnd.n2596 gnd.n2595 19.3944
R9488 gnd.n2596 gnd.n2420 19.3944
R9489 gnd.n2640 gnd.n2420 19.3944
R9490 gnd.n2640 gnd.n2639 19.3944
R9491 gnd.n2639 gnd.n2638 19.3944
R9492 gnd.n2638 gnd.n2602 19.3944
R9493 gnd.n2625 gnd.n2602 19.3944
R9494 gnd.n2625 gnd.n2624 19.3944
R9495 gnd.n2624 gnd.n2623 19.3944
R9496 gnd.n2623 gnd.n2374 19.3944
R9497 gnd.n2669 gnd.n2374 19.3944
R9498 gnd.n2669 gnd.n2372 19.3944
R9499 gnd.n2674 gnd.n2372 19.3944
R9500 gnd.n2674 gnd.n2366 19.3944
R9501 gnd.n2686 gnd.n2366 19.3944
R9502 gnd.n2687 gnd.n2686 19.3944
R9503 gnd.n2688 gnd.n2687 19.3944
R9504 gnd.n2688 gnd.n2364 19.3944
R9505 gnd.n2694 gnd.n2364 19.3944
R9506 gnd.n2695 gnd.n2694 19.3944
R9507 gnd.n2699 gnd.n2695 19.3944
R9508 gnd.n2699 gnd.n2362 19.3944
R9509 gnd.n2707 gnd.n2362 19.3944
R9510 gnd.n2707 gnd.n2706 19.3944
R9511 gnd.n2706 gnd.n2705 19.3944
R9512 gnd.n2705 gnd.n2338 19.3944
R9513 gnd.n2786 gnd.n2338 19.3944
R9514 gnd.n2786 gnd.n2336 19.3944
R9515 gnd.n2791 gnd.n2336 19.3944
R9516 gnd.n2791 gnd.n2330 19.3944
R9517 gnd.n2833 gnd.n2330 19.3944
R9518 gnd.n2834 gnd.n2833 19.3944
R9519 gnd.n2876 gnd.n2304 19.3944
R9520 gnd.n2876 gnd.n2873 19.3944
R9521 gnd.n2873 gnd.n2870 19.3944
R9522 gnd.n2870 gnd.n2869 19.3944
R9523 gnd.n2869 gnd.n2866 19.3944
R9524 gnd.n2866 gnd.n2865 19.3944
R9525 gnd.n2865 gnd.n2862 19.3944
R9526 gnd.n2862 gnd.n2861 19.3944
R9527 gnd.n2861 gnd.n2858 19.3944
R9528 gnd.n2858 gnd.n2857 19.3944
R9529 gnd.n2857 gnd.n2854 19.3944
R9530 gnd.n2854 gnd.n2853 19.3944
R9531 gnd.n2853 gnd.n2850 19.3944
R9532 gnd.n2850 gnd.n2849 19.3944
R9533 gnd.n2849 gnd.n2846 19.3944
R9534 gnd.n2846 gnd.n2845 19.3944
R9535 gnd.n2845 gnd.n2842 19.3944
R9536 gnd.n2842 gnd.n2841 19.3944
R9537 gnd.n2287 gnd.n2286 19.3944
R9538 gnd.n3140 gnd.n2286 19.3944
R9539 gnd.n3140 gnd.n3139 19.3944
R9540 gnd.n3139 gnd.n3138 19.3944
R9541 gnd.n3138 gnd.n3135 19.3944
R9542 gnd.n3135 gnd.n3134 19.3944
R9543 gnd.n3134 gnd.n3131 19.3944
R9544 gnd.n3131 gnd.n3130 19.3944
R9545 gnd.n3130 gnd.n3127 19.3944
R9546 gnd.n3127 gnd.n3126 19.3944
R9547 gnd.n3126 gnd.n3123 19.3944
R9548 gnd.n3123 gnd.n3122 19.3944
R9549 gnd.n3122 gnd.n3119 19.3944
R9550 gnd.n3119 gnd.n3118 19.3944
R9551 gnd.n3118 gnd.n3115 19.3944
R9552 gnd.n2542 gnd.n2474 19.3944
R9553 gnd.n2542 gnd.n2475 19.3944
R9554 gnd.n2538 gnd.n2475 19.3944
R9555 gnd.n2538 gnd.n1032 19.3944
R9556 gnd.n4810 gnd.n1032 19.3944
R9557 gnd.n4810 gnd.n4809 19.3944
R9558 gnd.n4809 gnd.n4808 19.3944
R9559 gnd.n4808 gnd.n1036 19.3944
R9560 gnd.n4798 gnd.n1036 19.3944
R9561 gnd.n4798 gnd.n4797 19.3944
R9562 gnd.n4797 gnd.n4796 19.3944
R9563 gnd.n4796 gnd.n1055 19.3944
R9564 gnd.n4786 gnd.n1055 19.3944
R9565 gnd.n4786 gnd.n4785 19.3944
R9566 gnd.n4785 gnd.n4784 19.3944
R9567 gnd.n4784 gnd.n1076 19.3944
R9568 gnd.n4774 gnd.n1076 19.3944
R9569 gnd.n4774 gnd.n4773 19.3944
R9570 gnd.n4773 gnd.n4772 19.3944
R9571 gnd.n4772 gnd.n1095 19.3944
R9572 gnd.n4762 gnd.n1095 19.3944
R9573 gnd.n4762 gnd.n4761 19.3944
R9574 gnd.n4761 gnd.n4760 19.3944
R9575 gnd.n4760 gnd.n1118 19.3944
R9576 gnd.n4750 gnd.n1118 19.3944
R9577 gnd.n4750 gnd.n4749 19.3944
R9578 gnd.n4749 gnd.n4748 19.3944
R9579 gnd.n4748 gnd.n1136 19.3944
R9580 gnd.n4737 gnd.n1136 19.3944
R9581 gnd.n4737 gnd.n4736 19.3944
R9582 gnd.n4736 gnd.n4735 19.3944
R9583 gnd.n4735 gnd.n1155 19.3944
R9584 gnd.n4725 gnd.n1155 19.3944
R9585 gnd.n4725 gnd.n4724 19.3944
R9586 gnd.n4724 gnd.n4723 19.3944
R9587 gnd.n4723 gnd.n1174 19.3944
R9588 gnd.n4713 gnd.n1174 19.3944
R9589 gnd.n4713 gnd.n4712 19.3944
R9590 gnd.n4712 gnd.n4711 19.3944
R9591 gnd.n4711 gnd.n1196 19.3944
R9592 gnd.n4701 gnd.n1196 19.3944
R9593 gnd.n4701 gnd.n4700 19.3944
R9594 gnd.n4700 gnd.n4699 19.3944
R9595 gnd.n4699 gnd.n1216 19.3944
R9596 gnd.n4689 gnd.n1216 19.3944
R9597 gnd.n4689 gnd.n4688 19.3944
R9598 gnd.n4688 gnd.n4687 19.3944
R9599 gnd.n4687 gnd.n1238 19.3944
R9600 gnd.n4677 gnd.n1238 19.3944
R9601 gnd.n4677 gnd.n4676 19.3944
R9602 gnd.n4676 gnd.n4675 19.3944
R9603 gnd.n4675 gnd.n1259 19.3944
R9604 gnd.n4665 gnd.n1259 19.3944
R9605 gnd.n2534 gnd.n2532 19.3944
R9606 gnd.n2532 gnd.n2529 19.3944
R9607 gnd.n2529 gnd.n2528 19.3944
R9608 gnd.n2528 gnd.n2525 19.3944
R9609 gnd.n2525 gnd.n2524 19.3944
R9610 gnd.n2524 gnd.n2521 19.3944
R9611 gnd.n2521 gnd.n2520 19.3944
R9612 gnd.n2520 gnd.n2517 19.3944
R9613 gnd.n2517 gnd.n2516 19.3944
R9614 gnd.n2516 gnd.n2513 19.3944
R9615 gnd.n2513 gnd.n2512 19.3944
R9616 gnd.n2512 gnd.n2509 19.3944
R9617 gnd.n2509 gnd.n2508 19.3944
R9618 gnd.n2508 gnd.n2505 19.3944
R9619 gnd.n2505 gnd.n2504 19.3944
R9620 gnd.n2504 gnd.n2501 19.3944
R9621 gnd.n2495 gnd.n2470 19.3944
R9622 gnd.n2553 gnd.n2470 19.3944
R9623 gnd.n2553 gnd.n2468 19.3944
R9624 gnd.n2558 gnd.n2468 19.3944
R9625 gnd.n2559 gnd.n2558 19.3944
R9626 gnd.n2561 gnd.n2559 19.3944
R9627 gnd.n2561 gnd.n2466 19.3944
R9628 gnd.n2566 gnd.n2466 19.3944
R9629 gnd.n2567 gnd.n2566 19.3944
R9630 gnd.n2569 gnd.n2567 19.3944
R9631 gnd.n2569 gnd.n2464 19.3944
R9632 gnd.n2574 gnd.n2464 19.3944
R9633 gnd.n2575 gnd.n2574 19.3944
R9634 gnd.n2577 gnd.n2575 19.3944
R9635 gnd.n2577 gnd.n2462 19.3944
R9636 gnd.n2582 gnd.n2462 19.3944
R9637 gnd.n2583 gnd.n2582 19.3944
R9638 gnd.n2585 gnd.n2583 19.3944
R9639 gnd.n2585 gnd.n2460 19.3944
R9640 gnd.n2590 gnd.n2460 19.3944
R9641 gnd.n2590 gnd.n2415 19.3944
R9642 gnd.n2646 gnd.n2415 19.3944
R9643 gnd.n2646 gnd.n2645 19.3944
R9644 gnd.n2645 gnd.n2644 19.3944
R9645 gnd.n2644 gnd.n2419 19.3944
R9646 gnd.n2634 gnd.n2419 19.3944
R9647 gnd.n2634 gnd.n2633 19.3944
R9648 gnd.n2633 gnd.n2629 19.3944
R9649 gnd.n2629 gnd.n2377 19.3944
R9650 gnd.n2661 gnd.n2377 19.3944
R9651 gnd.n2661 gnd.n2375 19.3944
R9652 gnd.n2665 gnd.n2375 19.3944
R9653 gnd.n2665 gnd.n2370 19.3944
R9654 gnd.n2678 gnd.n2370 19.3944
R9655 gnd.n2678 gnd.n2368 19.3944
R9656 gnd.n2682 gnd.n2368 19.3944
R9657 gnd.n2682 gnd.n2355 19.3944
R9658 gnd.n2721 gnd.n2355 19.3944
R9659 gnd.n2721 gnd.n2356 19.3944
R9660 gnd.n2717 gnd.n2356 19.3944
R9661 gnd.n2717 gnd.n2716 19.3944
R9662 gnd.n2716 gnd.n2715 19.3944
R9663 gnd.n2715 gnd.n2361 19.3944
R9664 gnd.n2711 gnd.n2361 19.3944
R9665 gnd.n2711 gnd.n2341 19.3944
R9666 gnd.n2778 gnd.n2341 19.3944
R9667 gnd.n2778 gnd.n2339 19.3944
R9668 gnd.n2782 gnd.n2339 19.3944
R9669 gnd.n2782 gnd.n2335 19.3944
R9670 gnd.n2795 gnd.n2335 19.3944
R9671 gnd.n2795 gnd.n2332 19.3944
R9672 gnd.n2829 gnd.n2332 19.3944
R9673 gnd.n2829 gnd.n2333 19.3944
R9674 gnd.n2548 gnd.n2544 19.3944
R9675 gnd.n2548 gnd.n1021 19.3944
R9676 gnd.n4816 gnd.n1021 19.3944
R9677 gnd.n4816 gnd.n4815 19.3944
R9678 gnd.n4815 gnd.n4814 19.3944
R9679 gnd.n4814 gnd.n1025 19.3944
R9680 gnd.n4804 gnd.n1025 19.3944
R9681 gnd.n4804 gnd.n4803 19.3944
R9682 gnd.n4803 gnd.n4802 19.3944
R9683 gnd.n4802 gnd.n1046 19.3944
R9684 gnd.n4792 gnd.n1046 19.3944
R9685 gnd.n4792 gnd.n4791 19.3944
R9686 gnd.n4791 gnd.n4790 19.3944
R9687 gnd.n4790 gnd.n1065 19.3944
R9688 gnd.n4780 gnd.n1065 19.3944
R9689 gnd.n4780 gnd.n4779 19.3944
R9690 gnd.n4779 gnd.n4778 19.3944
R9691 gnd.n4778 gnd.n1086 19.3944
R9692 gnd.n4768 gnd.n1086 19.3944
R9693 gnd.n4768 gnd.n4767 19.3944
R9694 gnd.n4767 gnd.n4766 19.3944
R9695 gnd.n4766 gnd.n1107 19.3944
R9696 gnd.n4756 gnd.n4755 19.3944
R9697 gnd.n4755 gnd.n4754 19.3944
R9698 gnd.n4744 gnd.n1143 19.3944
R9699 gnd.n4742 gnd.n4741 19.3944
R9700 gnd.n4731 gnd.n1161 19.3944
R9701 gnd.n4731 gnd.n4730 19.3944
R9702 gnd.n4730 gnd.n4729 19.3944
R9703 gnd.n4729 gnd.n1164 19.3944
R9704 gnd.n4719 gnd.n1164 19.3944
R9705 gnd.n4719 gnd.n4718 19.3944
R9706 gnd.n4718 gnd.n4717 19.3944
R9707 gnd.n4717 gnd.n1185 19.3944
R9708 gnd.n4707 gnd.n1185 19.3944
R9709 gnd.n4707 gnd.n4706 19.3944
R9710 gnd.n4706 gnd.n4705 19.3944
R9711 gnd.n4705 gnd.n1206 19.3944
R9712 gnd.n4695 gnd.n1206 19.3944
R9713 gnd.n4695 gnd.n4694 19.3944
R9714 gnd.n4694 gnd.n4693 19.3944
R9715 gnd.n4693 gnd.n1227 19.3944
R9716 gnd.n4683 gnd.n1227 19.3944
R9717 gnd.n4683 gnd.n4682 19.3944
R9718 gnd.n4682 gnd.n4681 19.3944
R9719 gnd.n4681 gnd.n1248 19.3944
R9720 gnd.n4671 gnd.n1248 19.3944
R9721 gnd.n4671 gnd.n4670 19.3944
R9722 gnd.n4670 gnd.n4669 19.3944
R9723 gnd.n6496 gnd.n730 19.3944
R9724 gnd.n6496 gnd.n6495 19.3944
R9725 gnd.n6495 gnd.n6494 19.3944
R9726 gnd.n6494 gnd.n734 19.3944
R9727 gnd.n6488 gnd.n734 19.3944
R9728 gnd.n6488 gnd.n6487 19.3944
R9729 gnd.n6487 gnd.n6486 19.3944
R9730 gnd.n6486 gnd.n742 19.3944
R9731 gnd.n6480 gnd.n742 19.3944
R9732 gnd.n6480 gnd.n6479 19.3944
R9733 gnd.n6479 gnd.n6478 19.3944
R9734 gnd.n6478 gnd.n750 19.3944
R9735 gnd.n6472 gnd.n750 19.3944
R9736 gnd.n6472 gnd.n6471 19.3944
R9737 gnd.n6471 gnd.n6470 19.3944
R9738 gnd.n6470 gnd.n758 19.3944
R9739 gnd.n6464 gnd.n758 19.3944
R9740 gnd.n6464 gnd.n6463 19.3944
R9741 gnd.n6463 gnd.n6462 19.3944
R9742 gnd.n6462 gnd.n766 19.3944
R9743 gnd.n6456 gnd.n766 19.3944
R9744 gnd.n6456 gnd.n6455 19.3944
R9745 gnd.n6455 gnd.n6454 19.3944
R9746 gnd.n6454 gnd.n774 19.3944
R9747 gnd.n6448 gnd.n774 19.3944
R9748 gnd.n6448 gnd.n6447 19.3944
R9749 gnd.n6447 gnd.n6446 19.3944
R9750 gnd.n6446 gnd.n782 19.3944
R9751 gnd.n6440 gnd.n782 19.3944
R9752 gnd.n6440 gnd.n6439 19.3944
R9753 gnd.n6439 gnd.n6438 19.3944
R9754 gnd.n6438 gnd.n790 19.3944
R9755 gnd.n6432 gnd.n790 19.3944
R9756 gnd.n6432 gnd.n6431 19.3944
R9757 gnd.n6431 gnd.n6430 19.3944
R9758 gnd.n6430 gnd.n798 19.3944
R9759 gnd.n6424 gnd.n798 19.3944
R9760 gnd.n6424 gnd.n6423 19.3944
R9761 gnd.n6423 gnd.n6422 19.3944
R9762 gnd.n6422 gnd.n806 19.3944
R9763 gnd.n6416 gnd.n806 19.3944
R9764 gnd.n6416 gnd.n6415 19.3944
R9765 gnd.n6415 gnd.n6414 19.3944
R9766 gnd.n6414 gnd.n814 19.3944
R9767 gnd.n6408 gnd.n814 19.3944
R9768 gnd.n6408 gnd.n6407 19.3944
R9769 gnd.n6407 gnd.n6406 19.3944
R9770 gnd.n6406 gnd.n822 19.3944
R9771 gnd.n6400 gnd.n822 19.3944
R9772 gnd.n6400 gnd.n6399 19.3944
R9773 gnd.n6399 gnd.n6398 19.3944
R9774 gnd.n6398 gnd.n830 19.3944
R9775 gnd.n6392 gnd.n830 19.3944
R9776 gnd.n6392 gnd.n6391 19.3944
R9777 gnd.n6391 gnd.n6390 19.3944
R9778 gnd.n6390 gnd.n838 19.3944
R9779 gnd.n6384 gnd.n838 19.3944
R9780 gnd.n6384 gnd.n6383 19.3944
R9781 gnd.n6383 gnd.n6382 19.3944
R9782 gnd.n6382 gnd.n846 19.3944
R9783 gnd.n6376 gnd.n846 19.3944
R9784 gnd.n6376 gnd.n6375 19.3944
R9785 gnd.n6375 gnd.n6374 19.3944
R9786 gnd.n6374 gnd.n854 19.3944
R9787 gnd.n6368 gnd.n854 19.3944
R9788 gnd.n6368 gnd.n6367 19.3944
R9789 gnd.n6367 gnd.n6366 19.3944
R9790 gnd.n6366 gnd.n862 19.3944
R9791 gnd.n6360 gnd.n862 19.3944
R9792 gnd.n6360 gnd.n6359 19.3944
R9793 gnd.n6359 gnd.n6358 19.3944
R9794 gnd.n6358 gnd.n870 19.3944
R9795 gnd.n6352 gnd.n870 19.3944
R9796 gnd.n6352 gnd.n6351 19.3944
R9797 gnd.n6351 gnd.n6350 19.3944
R9798 gnd.n6350 gnd.n878 19.3944
R9799 gnd.n6344 gnd.n878 19.3944
R9800 gnd.n6344 gnd.n6343 19.3944
R9801 gnd.n6343 gnd.n6342 19.3944
R9802 gnd.n6342 gnd.n886 19.3944
R9803 gnd.n6336 gnd.n886 19.3944
R9804 gnd.n6336 gnd.n6335 19.3944
R9805 gnd.n6335 gnd.n6334 19.3944
R9806 gnd.n6334 gnd.n894 19.3944
R9807 gnd.n4660 gnd.n4659 19.3944
R9808 gnd.n4659 gnd.n4658 19.3944
R9809 gnd.n4658 gnd.n1282 19.3944
R9810 gnd.n4654 gnd.n1282 19.3944
R9811 gnd.n4654 gnd.n4653 19.3944
R9812 gnd.n4653 gnd.n4652 19.3944
R9813 gnd.n4652 gnd.n1287 19.3944
R9814 gnd.n4648 gnd.n1287 19.3944
R9815 gnd.n4648 gnd.n4647 19.3944
R9816 gnd.n4647 gnd.n4646 19.3944
R9817 gnd.n4646 gnd.n1292 19.3944
R9818 gnd.n4642 gnd.n1292 19.3944
R9819 gnd.n4642 gnd.n4641 19.3944
R9820 gnd.n4641 gnd.n4640 19.3944
R9821 gnd.n4640 gnd.n1297 19.3944
R9822 gnd.n4636 gnd.n1297 19.3944
R9823 gnd.n4636 gnd.n4635 19.3944
R9824 gnd.n4635 gnd.n4634 19.3944
R9825 gnd.n4634 gnd.n1302 19.3944
R9826 gnd.n4630 gnd.n1302 19.3944
R9827 gnd.n4630 gnd.n4629 19.3944
R9828 gnd.n4629 gnd.n4628 19.3944
R9829 gnd.n4628 gnd.n1307 19.3944
R9830 gnd.n4624 gnd.n1307 19.3944
R9831 gnd.n4624 gnd.n4623 19.3944
R9832 gnd.n4623 gnd.n4622 19.3944
R9833 gnd.n4622 gnd.n1312 19.3944
R9834 gnd.n4618 gnd.n1312 19.3944
R9835 gnd.n4618 gnd.n4617 19.3944
R9836 gnd.n4617 gnd.n4616 19.3944
R9837 gnd.n4616 gnd.n1317 19.3944
R9838 gnd.n4612 gnd.n1317 19.3944
R9839 gnd.n4612 gnd.n4611 19.3944
R9840 gnd.n4611 gnd.n4610 19.3944
R9841 gnd.n4610 gnd.n1322 19.3944
R9842 gnd.n4606 gnd.n1322 19.3944
R9843 gnd.n4606 gnd.n4605 19.3944
R9844 gnd.n4605 gnd.n4604 19.3944
R9845 gnd.n4604 gnd.n1327 19.3944
R9846 gnd.n4600 gnd.n1327 19.3944
R9847 gnd.n4600 gnd.n4599 19.3944
R9848 gnd.n4599 gnd.n4598 19.3944
R9849 gnd.n4598 gnd.n1332 19.3944
R9850 gnd.n4594 gnd.n1332 19.3944
R9851 gnd.n4594 gnd.n4593 19.3944
R9852 gnd.n4593 gnd.n4592 19.3944
R9853 gnd.n4592 gnd.n1337 19.3944
R9854 gnd.n4588 gnd.n1337 19.3944
R9855 gnd.n4588 gnd.n4587 19.3944
R9856 gnd.n4587 gnd.n4586 19.3944
R9857 gnd.n4586 gnd.n1342 19.3944
R9858 gnd.n4582 gnd.n1342 19.3944
R9859 gnd.n4582 gnd.n4581 19.3944
R9860 gnd.n4581 gnd.n4580 19.3944
R9861 gnd.n4580 gnd.n1347 19.3944
R9862 gnd.n4576 gnd.n1347 19.3944
R9863 gnd.n4576 gnd.n4575 19.3944
R9864 gnd.n4575 gnd.n4574 19.3944
R9865 gnd.n4574 gnd.n1352 19.3944
R9866 gnd.n4570 gnd.n1352 19.3944
R9867 gnd.n4570 gnd.n4569 19.3944
R9868 gnd.n4569 gnd.n4568 19.3944
R9869 gnd.n4568 gnd.n1357 19.3944
R9870 gnd.n4564 gnd.n1357 19.3944
R9871 gnd.n4564 gnd.n4563 19.3944
R9872 gnd.n4563 gnd.n4562 19.3944
R9873 gnd.n4562 gnd.n1362 19.3944
R9874 gnd.n4558 gnd.n1362 19.3944
R9875 gnd.n4558 gnd.n4557 19.3944
R9876 gnd.n4557 gnd.n4556 19.3944
R9877 gnd.n4556 gnd.n1367 19.3944
R9878 gnd.n4552 gnd.n1367 19.3944
R9879 gnd.n4552 gnd.n4551 19.3944
R9880 gnd.n4551 gnd.n4550 19.3944
R9881 gnd.n4550 gnd.n1372 19.3944
R9882 gnd.n4546 gnd.n1372 19.3944
R9883 gnd.n4546 gnd.n4545 19.3944
R9884 gnd.n4545 gnd.n4544 19.3944
R9885 gnd.n4544 gnd.n1377 19.3944
R9886 gnd.n4540 gnd.n1377 19.3944
R9887 gnd.n4540 gnd.n4539 19.3944
R9888 gnd.n4539 gnd.n4538 19.3944
R9889 gnd.n4538 gnd.n1382 19.3944
R9890 gnd.n4534 gnd.n1382 19.3944
R9891 gnd.n4534 gnd.n4533 19.3944
R9892 gnd.n4533 gnd.n4532 19.3944
R9893 gnd.n4532 gnd.n1387 19.3944
R9894 gnd.n4528 gnd.n1387 19.3944
R9895 gnd.n4528 gnd.n4527 19.3944
R9896 gnd.n4527 gnd.n4526 19.3944
R9897 gnd.n4526 gnd.n1392 19.3944
R9898 gnd.n4522 gnd.n1392 19.3944
R9899 gnd.n4522 gnd.n4521 19.3944
R9900 gnd.n4521 gnd.n4520 19.3944
R9901 gnd.n4520 gnd.n1397 19.3944
R9902 gnd.n4516 gnd.n1397 19.3944
R9903 gnd.n4516 gnd.n4515 19.3944
R9904 gnd.n4515 gnd.n4514 19.3944
R9905 gnd.n4514 gnd.n1402 19.3944
R9906 gnd.n4510 gnd.n1402 19.3944
R9907 gnd.n4510 gnd.n4509 19.3944
R9908 gnd.n4215 gnd.n1819 19.3944
R9909 gnd.n4211 gnd.n1819 19.3944
R9910 gnd.n4211 gnd.n4210 19.3944
R9911 gnd.n1735 gnd.n1719 19.3944
R9912 gnd.n1735 gnd.n1717 19.3944
R9913 gnd.n1741 gnd.n1717 19.3944
R9914 gnd.n1741 gnd.n1712 19.3944
R9915 gnd.n1754 gnd.n1712 19.3944
R9916 gnd.n1754 gnd.n1710 19.3944
R9917 gnd.n1760 gnd.n1710 19.3944
R9918 gnd.n1760 gnd.n1705 19.3944
R9919 gnd.n1773 gnd.n1705 19.3944
R9920 gnd.n1773 gnd.n1703 19.3944
R9921 gnd.n1779 gnd.n1703 19.3944
R9922 gnd.n1779 gnd.n1699 19.3944
R9923 gnd.n1789 gnd.n1699 19.3944
R9924 gnd.n1789 gnd.n1697 19.3944
R9925 gnd.n1795 gnd.n1697 19.3944
R9926 gnd.n1795 gnd.n1687 19.3944
R9927 gnd.n1803 gnd.n1687 19.3944
R9928 gnd.n1803 gnd.n1685 19.3944
R9929 gnd.n4226 gnd.n1685 19.3944
R9930 gnd.n4226 gnd.n4225 19.3944
R9931 gnd.n4225 gnd.n4224 19.3944
R9932 gnd.n4224 gnd.n1811 19.3944
R9933 gnd.n4220 gnd.n1811 19.3944
R9934 gnd.n4220 gnd.n4219 19.3944
R9935 gnd.n3011 gnd.n3010 19.2005
R9936 gnd.n3687 gnd.n3686 19.2005
R9937 gnd.n3914 gnd.n2067 19.1199
R9938 gnd.n3368 gnd.n2009 19.1199
R9939 gnd.n4018 gnd.n1972 19.1199
R9940 gnd.n3456 gnd.n1911 19.1199
R9941 gnd.t52 gnd.n5133 18.8012
R9942 gnd.n5737 gnd.t268 18.8012
R9943 gnd.n3308 gnd.t49 18.8012
R9944 gnd.n3716 gnd.t239 18.8012
R9945 gnd.n5582 gnd.n5581 18.4825
R9946 gnd.n4764 gnd.n1109 18.4825
R9947 gnd.n2648 gnd.n1112 18.4825
R9948 gnd.n2642 gnd.n1122 18.4825
R9949 gnd.n4752 gnd.n1128 18.4825
R9950 gnd.n2636 gnd.n2614 18.4825
R9951 gnd.n4746 gnd.n1138 18.4825
R9952 gnd.n4739 gnd.n1146 18.4825
R9953 gnd.n2659 gnd.n1149 18.4825
R9954 gnd.n2667 gnd.n1159 18.4825
R9955 gnd.n4727 gnd.n1166 18.4825
R9956 gnd.n2676 gnd.n2371 18.4825
R9957 gnd.n4721 gnd.n1176 18.4825
R9958 gnd.n4715 gnd.n1187 18.4825
R9959 gnd.n2723 gnd.n1190 18.4825
R9960 gnd.n2692 gnd.n1200 18.4825
R9961 gnd.n4703 gnd.n1208 18.4825
R9962 gnd.n2697 gnd.n2696 18.4825
R9963 gnd.n4697 gnd.n1218 18.4825
R9964 gnd.n4691 gnd.n1229 18.4825
R9965 gnd.n2776 gnd.n1232 18.4825
R9966 gnd.n2784 gnd.n1242 18.4825
R9967 gnd.n4679 gnd.n1250 18.4825
R9968 gnd.n2793 gnd.n1253 18.4825
R9969 gnd.n4673 gnd.n1261 18.4825
R9970 gnd.n2831 gnd.n2331 18.4825
R9971 gnd.n4667 gnd.n1270 18.4825
R9972 gnd.n4422 gnd.n1499 18.4825
R9973 gnd.n4237 gnd.n1647 18.4825
R9974 gnd.n4236 gnd.n1625 18.4825
R9975 gnd.n4248 gnd.n4247 18.4825
R9976 gnd.n1628 gnd.n1615 18.4825
R9977 gnd.n4258 gnd.n1617 18.4825
R9978 gnd.n4267 gnd.n1597 18.4825
R9979 gnd.n4279 gnd.n4278 18.4825
R9980 gnd.n4289 gnd.n1590 18.4825
R9981 gnd.n4304 gnd.n1580 18.4825
R9982 gnd.n4303 gnd.n1570 18.4825
R9983 gnd.n4316 gnd.n4314 18.4825
R9984 gnd.n4326 gnd.n1563 18.4825
R9985 gnd.n4362 gnd.n1546 18.4825
R9986 gnd.n4379 gnd.n4378 18.4825
R9987 gnd.n1540 gnd.n1538 18.4825
R9988 gnd.n4387 gnd.n1529 18.4825
R9989 gnd.n4349 gnd.n278 18.4825
R9990 gnd.n7192 gnd.n7191 18.4825
R9991 gnd.n314 gnd.n307 18.4825
R9992 gnd.n7205 gnd.n304 18.4825
R9993 gnd.n321 gnd.n320 18.4825
R9994 gnd.n7271 gnd.n294 18.4825
R9995 gnd.n7276 gnd.n296 18.4825
R9996 gnd.n7299 gnd.n265 18.4825
R9997 gnd.n7260 gnd.n256 18.4825
R9998 gnd.n4467 gnd.n4466 18.4247
R9999 gnd.n3115 gnd.n3114 18.4247
R10000 gnd.n7411 gnd.n7410 18.2308
R10001 gnd.n1799 gnd.n1798 18.2308
R10002 gnd.n3153 gnd.n2240 18.2308
R10003 gnd.n2501 gnd.n2494 18.2308
R10004 gnd.t14 gnd.n5177 18.1639
R10005 gnd.n6331 gnd.n6330 18.1639
R10006 gnd.n2906 gnd.n2904 17.8452
R10007 gnd.n3922 gnd.n2059 17.8452
R10008 gnd.n3375 gnd.n2002 17.8452
R10009 gnd.n4010 gnd.n1979 17.8452
R10010 gnd.n3737 gnd.n1917 17.8452
R10011 gnd.n3494 gnd.n1884 17.8452
R10012 gnd.n5204 gnd.t12 17.5266
R10013 gnd.t7 gnd.n1029 17.5266
R10014 gnd.n4685 gnd.t39 17.5266
R10015 gnd.n1671 gnd.t42 17.5266
R10016 gnd.n7363 gnd.t168 17.5266
R10017 gnd.t197 gnd.n2037 17.2079
R10018 gnd.n3430 gnd.t38 17.2079
R10019 gnd.n5162 gnd.t55 16.8893
R10020 gnd.t243 gnd.n1070 16.8893
R10021 gnd.n4709 gnd.t181 16.8893
R10022 gnd.n1573 gnd.t192 16.8893
R10023 gnd.n7331 gnd.t29 16.8893
R10024 gnd.n3930 gnd.n2052 16.5706
R10025 gnd.t267 gnd.n3851 16.5706
R10026 gnd.n3382 gnd.n1994 16.5706
R10027 gnd.n4002 gnd.n1987 16.5706
R10028 gnd.n3766 gnd.t262 16.5706
R10029 gnd.n3443 gnd.n1924 16.5706
R10030 gnd.n5431 gnd.t108 16.2519
R10031 gnd.n5727 gnd.t10 16.2519
R10032 gnd.n4733 gnd.t46 16.2519
R10033 gnd.n7292 gnd.t225 16.2519
R10034 gnd.t172 gnd.n2023 15.9333
R10035 gnd.n3774 gnd.t196 15.9333
R10036 gnd.n6137 gnd.n6135 15.6674
R10037 gnd.n6105 gnd.n6103 15.6674
R10038 gnd.n6073 gnd.n6071 15.6674
R10039 gnd.n6042 gnd.n6040 15.6674
R10040 gnd.n6010 gnd.n6008 15.6674
R10041 gnd.n5978 gnd.n5976 15.6674
R10042 gnd.n5946 gnd.n5944 15.6674
R10043 gnd.n5915 gnd.n5913 15.6674
R10044 gnd.n5422 gnd.t108 15.6146
R10045 gnd.t68 gnd.n6316 15.6146
R10046 gnd.n6220 gnd.t80 15.6146
R10047 gnd.n4758 gnd.t174 15.6146
R10048 gnd.n7265 gnd.t205 15.6146
R10049 gnd.n3321 gnd.n2052 15.296
R10050 gnd.n3938 gnd.n2044 15.296
R10051 gnd.t198 gnd.n2015 15.296
R10052 gnd.n3994 gnd.n1994 15.296
R10053 gnd.n3389 gnd.n1987 15.296
R10054 gnd.n3781 gnd.t51 15.296
R10055 gnd.n3752 gnd.n3751 15.296
R10056 gnd.n4074 gnd.n1924 15.296
R10057 gnd.n3489 gnd.t91 15.296
R10058 gnd.n3500 gnd.n3499 15.0827
R10059 gnd.n2916 gnd.n2911 15.0481
R10060 gnd.n3510 gnd.n3509 15.0481
R10061 gnd.n5865 gnd.t36 14.9773
R10062 gnd.n4782 gnd.t243 14.9773
R10063 gnd.n241 gnd.t29 14.9773
R10064 gnd.t292 gnd.n2008 14.6587
R10065 gnd.n3789 gnd.t266 14.6587
R10066 gnd.n3477 gnd.t88 14.6587
R10067 gnd.t19 gnd.n5006 14.34
R10068 gnd.t13 gnd.n898 14.34
R10069 gnd.n4806 gnd.t7 14.34
R10070 gnd.n3036 gnd.t248 14.34
R10071 gnd.t325 gnd.n3490 14.34
R10072 gnd.n211 gnd.t168 14.34
R10073 gnd.n3882 gnd.n2059 14.0214
R10074 gnd.n3946 gnd.n2037 14.0214
R10075 gnd.t294 gnd.n2000 14.0214
R10076 gnd.n3986 gnd.n2002 14.0214
R10077 gnd.n3396 gnd.n1979 14.0214
R10078 gnd.n3796 gnd.t219 14.0214
R10079 gnd.n3430 gnd.n3428 14.0214
R10080 gnd.n4082 gnd.n1917 14.0214
R10081 gnd.n4122 gnd.n1884 14.0214
R10082 gnd.n5547 gnd.t0 13.7027
R10083 gnd.t31 gnd.n1101 13.7027
R10084 gnd.n3361 gnd.t263 13.7027
R10085 gnd.n4026 gnd.t246 13.7027
R10086 gnd.n7171 gnd.t185 13.7027
R10087 gnd.n5288 gnd.n5287 13.5763
R10088 gnd.n6276 gnd.n4938 13.5763
R10089 gnd.n4429 gnd.n1493 13.5763
R10090 gnd.n7463 gnd.n7462 13.5763
R10091 gnd.n4832 gnd.n1007 13.5763
R10092 gnd.n2841 gnd.n2838 13.5763
R10093 gnd.n5582 gnd.n5234 13.384
R10094 gnd.n4770 gnd.n1101 13.384
R10095 gnd.n2592 gnd.n1109 13.384
R10096 gnd.n4764 gnd.n1112 13.384
R10097 gnd.n2649 gnd.n2648 13.384
R10098 gnd.n4758 gnd.n1122 13.384
R10099 gnd.n2642 gnd.n1128 13.384
R10100 gnd.n2636 gnd.n1138 13.384
R10101 gnd.n4746 gnd.n1141 13.384
R10102 gnd.n2627 gnd.n1146 13.384
R10103 gnd.n4739 gnd.n1149 13.384
R10104 gnd.n2659 gnd.n2658 13.384
R10105 gnd.n4733 gnd.n1159 13.384
R10106 gnd.n2667 gnd.n1166 13.384
R10107 gnd.n2676 gnd.n1176 13.384
R10108 gnd.n4721 gnd.n1179 13.384
R10109 gnd.n2684 gnd.n1187 13.384
R10110 gnd.n4715 gnd.n1190 13.384
R10111 gnd.n2724 gnd.n2723 13.384
R10112 gnd.n4709 gnd.n1200 13.384
R10113 gnd.n2692 gnd.n1208 13.384
R10114 gnd.n2697 gnd.n1218 13.384
R10115 gnd.n4697 gnd.n1221 13.384
R10116 gnd.n2709 gnd.n1229 13.384
R10117 gnd.n4691 gnd.n1232 13.384
R10118 gnd.n2776 gnd.n2775 13.384
R10119 gnd.n4685 gnd.n1242 13.384
R10120 gnd.n2784 gnd.n1250 13.384
R10121 gnd.n4679 gnd.n1253 13.384
R10122 gnd.n2793 gnd.n1261 13.384
R10123 gnd.n2831 gnd.n1270 13.384
R10124 gnd.n4667 gnd.n1273 13.384
R10125 gnd.t37 gnd.n1993 13.384
R10126 gnd.n3803 gnd.t291 13.384
R10127 gnd.n4422 gnd.n1497 13.384
R10128 gnd.n1647 gnd.n1499 13.384
R10129 gnd.n4248 gnd.n1625 13.384
R10130 gnd.n4247 gnd.n1628 13.384
R10131 gnd.n4258 gnd.n1615 13.384
R10132 gnd.n1671 gnd.n1617 13.384
R10133 gnd.n4268 gnd.n4267 13.384
R10134 gnd.n4279 gnd.n1597 13.384
R10135 gnd.n4278 gnd.n1601 13.384
R10136 gnd.n4289 gnd.n1588 13.384
R10137 gnd.n1590 gnd.n1580 13.384
R10138 gnd.n4316 gnd.n1570 13.384
R10139 gnd.n4314 gnd.n1573 13.384
R10140 gnd.n4326 gnd.n1561 13.384
R10141 gnd.n1563 gnd.n1546 13.384
R10142 gnd.n4362 gnd.n4361 13.384
R10143 gnd.n4379 gnd.n1535 13.384
R10144 gnd.n4378 gnd.n1538 13.384
R10145 gnd.n4349 gnd.n1529 13.384
R10146 gnd.n7292 gnd.n278 13.384
R10147 gnd.n7192 gnd.n312 13.384
R10148 gnd.n7191 gnd.n314 13.384
R10149 gnd.n7200 gnd.n307 13.384
R10150 gnd.n7205 gnd.n302 13.384
R10151 gnd.n320 gnd.n304 13.384
R10152 gnd.n7276 gnd.n294 13.384
R10153 gnd.n7265 gnd.n296 13.384
R10154 gnd.n7299 gnd.n263 13.384
R10155 gnd.n7260 gnd.n265 13.384
R10156 gnd.n7307 gnd.n256 13.384
R10157 gnd.n7171 gnd.n248 13.384
R10158 gnd.n2927 gnd.n2908 13.1884
R10159 gnd.n2922 gnd.n2921 13.1884
R10160 gnd.n2921 gnd.n2920 13.1884
R10161 gnd.n3503 gnd.n3498 13.1884
R10162 gnd.n3504 gnd.n3503 13.1884
R10163 gnd.n2923 gnd.n2910 13.146
R10164 gnd.n2919 gnd.n2910 13.146
R10165 gnd.n3502 gnd.n3501 13.146
R10166 gnd.n3502 gnd.n3497 13.146
R10167 gnd.t33 gnd.n1141 13.0654
R10168 gnd.t233 gnd.n302 13.0654
R10169 gnd.n6138 gnd.n6134 12.8005
R10170 gnd.n6106 gnd.n6102 12.8005
R10171 gnd.n6074 gnd.n6070 12.8005
R10172 gnd.n6043 gnd.n6039 12.8005
R10173 gnd.n6011 gnd.n6007 12.8005
R10174 gnd.n5979 gnd.n5975 12.8005
R10175 gnd.n5947 gnd.n5943 12.8005
R10176 gnd.n5916 gnd.n5912 12.8005
R10177 gnd.n3292 gnd.n2102 12.7467
R10178 gnd.n3898 gnd.t129 12.7467
R10179 gnd.n2090 gnd.n2067 12.7467
R10180 gnd.n3978 gnd.n2009 12.7467
R10181 gnd.n3403 gnd.n1972 12.7467
R10182 gnd.n4090 gnd.n1911 12.7467
R10183 gnd.n3690 gnd.t122 12.7467
R10184 gnd.t21 gnd.n1179 12.4281
R10185 gnd.t15 gnd.n2151 12.4281
R10186 gnd.n1845 gnd.t283 12.4281
R10187 gnd.t183 gnd.n1535 12.4281
R10188 gnd.n5287 gnd.n5282 12.4126
R10189 gnd.n6281 gnd.n4938 12.4126
R10190 gnd.n4425 gnd.n1493 12.4126
R10191 gnd.n7462 gnd.n178 12.4126
R10192 gnd.n4828 gnd.n1007 12.4126
R10193 gnd.n2838 gnd.n2326 12.4126
R10194 gnd.n3010 gnd.n3009 12.1761
R10195 gnd.n3686 gnd.n3685 12.1761
R10196 gnd.n3143 gnd.n2249 12.1094
R10197 gnd.n3282 gnd.t99 12.1094
R10198 gnd.n4498 gnd.n1446 12.1094
R10199 gnd.n6142 gnd.n6141 12.0247
R10200 gnd.n6110 gnd.n6109 12.0247
R10201 gnd.n6078 gnd.n6077 12.0247
R10202 gnd.n6047 gnd.n6046 12.0247
R10203 gnd.n6015 gnd.n6014 12.0247
R10204 gnd.n5983 gnd.n5982 12.0247
R10205 gnd.n5951 gnd.n5950 12.0247
R10206 gnd.n5920 gnd.n5919 12.0247
R10207 gnd.t272 gnd.n1221 11.7908
R10208 gnd.t23 gnd.n1588 11.7908
R10209 gnd.n3301 gnd.n2095 11.4721
R10210 gnd.n3307 gnd.n2074 11.4721
R10211 gnd.n3962 gnd.n2023 11.4721
R10212 gnd.n3970 gnd.n2017 11.4721
R10213 gnd.n3783 gnd.n3782 11.4721
R10214 gnd.n3774 gnd.n3415 11.4721
R10215 gnd.n4098 gnd.n1904 11.4721
R10216 gnd.n4106 gnd.n1898 11.4721
R10217 gnd.n6145 gnd.n6132 11.249
R10218 gnd.n6113 gnd.n6100 11.249
R10219 gnd.n6081 gnd.n6068 11.249
R10220 gnd.n6050 gnd.n6037 11.249
R10221 gnd.n6018 gnd.n6005 11.249
R10222 gnd.n5986 gnd.n5973 11.249
R10223 gnd.n5954 gnd.n5941 11.249
R10224 gnd.n5923 gnd.n5910 11.249
R10225 gnd.n5655 gnd.t0 11.1535
R10226 gnd.n3851 gnd.t305 11.1535
R10227 gnd.t299 gnd.n3766 11.1535
R10228 gnd.n3620 gnd.n3541 10.6151
R10229 gnd.n3620 gnd.n3619 10.6151
R10230 gnd.n3617 gnd.n3545 10.6151
R10231 gnd.n3612 gnd.n3545 10.6151
R10232 gnd.n3612 gnd.n3611 10.6151
R10233 gnd.n3611 gnd.n3610 10.6151
R10234 gnd.n3610 gnd.n3548 10.6151
R10235 gnd.n3605 gnd.n3548 10.6151
R10236 gnd.n3605 gnd.n3604 10.6151
R10237 gnd.n3604 gnd.n3603 10.6151
R10238 gnd.n3603 gnd.n3551 10.6151
R10239 gnd.n3598 gnd.n3551 10.6151
R10240 gnd.n3598 gnd.n3597 10.6151
R10241 gnd.n3597 gnd.n3596 10.6151
R10242 gnd.n3596 gnd.n3554 10.6151
R10243 gnd.n3591 gnd.n3554 10.6151
R10244 gnd.n3591 gnd.n3590 10.6151
R10245 gnd.n3590 gnd.n3589 10.6151
R10246 gnd.n3589 gnd.n3557 10.6151
R10247 gnd.n3584 gnd.n3557 10.6151
R10248 gnd.n3584 gnd.n3583 10.6151
R10249 gnd.n3583 gnd.n3582 10.6151
R10250 gnd.n3582 gnd.n3560 10.6151
R10251 gnd.n3577 gnd.n3560 10.6151
R10252 gnd.n3577 gnd.n3576 10.6151
R10253 gnd.n3576 gnd.n3575 10.6151
R10254 gnd.n3575 gnd.n3563 10.6151
R10255 gnd.n3570 gnd.n3563 10.6151
R10256 gnd.n3570 gnd.n3569 10.6151
R10257 gnd.n3569 gnd.n3568 10.6151
R10258 gnd.n2902 gnd.n2900 10.6151
R10259 gnd.n3016 gnd.n2902 10.6151
R10260 gnd.n3017 gnd.n3016 10.6151
R10261 gnd.n3033 gnd.n3017 10.6151
R10262 gnd.n3033 gnd.n3032 10.6151
R10263 gnd.n3032 gnd.n3031 10.6151
R10264 gnd.n3031 gnd.n3018 10.6151
R10265 gnd.n3019 gnd.n3018 10.6151
R10266 gnd.n3019 gnd.n2086 10.6151
R10267 gnd.n3896 gnd.n2086 10.6151
R10268 gnd.n3896 gnd.n3895 10.6151
R10269 gnd.n3895 gnd.n3894 10.6151
R10270 gnd.n3894 gnd.n2087 10.6151
R10271 gnd.n2089 gnd.n2087 10.6151
R10272 gnd.n3317 gnd.n2089 10.6151
R10273 gnd.n3318 gnd.n3317 10.6151
R10274 gnd.n3880 gnd.n3318 10.6151
R10275 gnd.n3880 gnd.n3879 10.6151
R10276 gnd.n3879 gnd.n3878 10.6151
R10277 gnd.n3878 gnd.n3319 10.6151
R10278 gnd.n3330 gnd.n3319 10.6151
R10279 gnd.n3331 gnd.n3330 10.6151
R10280 gnd.n3865 gnd.n3331 10.6151
R10281 gnd.n3865 gnd.n3864 10.6151
R10282 gnd.n3864 gnd.n3863 10.6151
R10283 gnd.n3863 gnd.n3332 10.6151
R10284 gnd.n3343 gnd.n3332 10.6151
R10285 gnd.n3345 gnd.n3343 10.6151
R10286 gnd.n3346 gnd.n3345 10.6151
R10287 gnd.n3849 gnd.n3346 10.6151
R10288 gnd.n3849 gnd.n3848 10.6151
R10289 gnd.n3848 gnd.n3847 10.6151
R10290 gnd.n3847 gnd.n3347 10.6151
R10291 gnd.n3358 gnd.n3347 10.6151
R10292 gnd.n3836 gnd.n3358 10.6151
R10293 gnd.n3836 gnd.n3835 10.6151
R10294 gnd.n3835 gnd.n3834 10.6151
R10295 gnd.n3834 gnd.n3359 10.6151
R10296 gnd.n3371 gnd.n3359 10.6151
R10297 gnd.n3372 gnd.n3371 10.6151
R10298 gnd.n3822 gnd.n3372 10.6151
R10299 gnd.n3822 gnd.n3821 10.6151
R10300 gnd.n3821 gnd.n3820 10.6151
R10301 gnd.n3820 gnd.n3373 10.6151
R10302 gnd.n3385 gnd.n3373 10.6151
R10303 gnd.n3386 gnd.n3385 10.6151
R10304 gnd.n3808 gnd.n3386 10.6151
R10305 gnd.n3808 gnd.n3807 10.6151
R10306 gnd.n3807 gnd.n3806 10.6151
R10307 gnd.n3806 gnd.n3387 10.6151
R10308 gnd.n3399 gnd.n3387 10.6151
R10309 gnd.n3400 gnd.n3399 10.6151
R10310 gnd.n3794 gnd.n3400 10.6151
R10311 gnd.n3794 gnd.n3793 10.6151
R10312 gnd.n3793 gnd.n3792 10.6151
R10313 gnd.n3792 gnd.n3401 10.6151
R10314 gnd.n3411 gnd.n3401 10.6151
R10315 gnd.n3412 gnd.n3411 10.6151
R10316 gnd.n3779 gnd.n3412 10.6151
R10317 gnd.n3779 gnd.n3778 10.6151
R10318 gnd.n3778 gnd.n3777 10.6151
R10319 gnd.n3777 gnd.n3413 10.6151
R10320 gnd.n3424 gnd.n3413 10.6151
R10321 gnd.n3425 gnd.n3424 10.6151
R10322 gnd.n3764 gnd.n3425 10.6151
R10323 gnd.n3764 gnd.n3763 10.6151
R10324 gnd.n3763 gnd.n3762 10.6151
R10325 gnd.n3762 gnd.n3426 10.6151
R10326 gnd.n3438 gnd.n3426 10.6151
R10327 gnd.n3439 gnd.n3438 10.6151
R10328 gnd.n3749 gnd.n3439 10.6151
R10329 gnd.n3749 gnd.n3748 10.6151
R10330 gnd.n3748 gnd.n3747 10.6151
R10331 gnd.n3747 gnd.n3440 10.6151
R10332 gnd.n3452 gnd.n3440 10.6151
R10333 gnd.n3735 gnd.n3452 10.6151
R10334 gnd.n3735 gnd.n3734 10.6151
R10335 gnd.n3734 gnd.n3733 10.6151
R10336 gnd.n3733 gnd.n3453 10.6151
R10337 gnd.n3465 gnd.n3453 10.6151
R10338 gnd.n3466 gnd.n3465 10.6151
R10339 gnd.n3720 gnd.n3466 10.6151
R10340 gnd.n3720 gnd.n3719 10.6151
R10341 gnd.n3719 gnd.n3718 10.6151
R10342 gnd.n3718 gnd.n3467 10.6151
R10343 gnd.n3481 gnd.n3467 10.6151
R10344 gnd.n3482 gnd.n3481 10.6151
R10345 gnd.n3706 gnd.n3482 10.6151
R10346 gnd.n3706 gnd.n3705 10.6151
R10347 gnd.n3705 gnd.n3704 10.6151
R10348 gnd.n3704 gnd.n3483 10.6151
R10349 gnd.n3694 gnd.n3483 10.6151
R10350 gnd.n3694 gnd.n3693 10.6151
R10351 gnd.n3693 gnd.n3692 10.6151
R10352 gnd.n3692 gnd.n3492 10.6151
R10353 gnd.n3107 gnd.n2880 10.6151
R10354 gnd.n3107 gnd.n3106 10.6151
R10355 gnd.n3104 gnd.n2886 10.6151
R10356 gnd.n3098 gnd.n2886 10.6151
R10357 gnd.n3098 gnd.n3097 10.6151
R10358 gnd.n3097 gnd.n3096 10.6151
R10359 gnd.n3096 gnd.n2888 10.6151
R10360 gnd.n3090 gnd.n2888 10.6151
R10361 gnd.n3090 gnd.n3089 10.6151
R10362 gnd.n3089 gnd.n3088 10.6151
R10363 gnd.n3088 gnd.n2890 10.6151
R10364 gnd.n3082 gnd.n2890 10.6151
R10365 gnd.n3082 gnd.n3081 10.6151
R10366 gnd.n3081 gnd.n3080 10.6151
R10367 gnd.n3080 gnd.n2892 10.6151
R10368 gnd.n3074 gnd.n2892 10.6151
R10369 gnd.n3074 gnd.n3073 10.6151
R10370 gnd.n3073 gnd.n3072 10.6151
R10371 gnd.n3072 gnd.n2894 10.6151
R10372 gnd.n3066 gnd.n2894 10.6151
R10373 gnd.n3066 gnd.n3065 10.6151
R10374 gnd.n3065 gnd.n3064 10.6151
R10375 gnd.n3064 gnd.n2896 10.6151
R10376 gnd.n3058 gnd.n2896 10.6151
R10377 gnd.n3058 gnd.n3057 10.6151
R10378 gnd.n3057 gnd.n3056 10.6151
R10379 gnd.n3056 gnd.n2898 10.6151
R10380 gnd.n3050 gnd.n2898 10.6151
R10381 gnd.n3050 gnd.n3049 10.6151
R10382 gnd.n3049 gnd.n3048 10.6151
R10383 gnd.n3009 gnd.n2928 10.6151
R10384 gnd.n3004 gnd.n2928 10.6151
R10385 gnd.n3004 gnd.n3003 10.6151
R10386 gnd.n3003 gnd.n3002 10.6151
R10387 gnd.n3002 gnd.n2930 10.6151
R10388 gnd.n2996 gnd.n2930 10.6151
R10389 gnd.n2996 gnd.n2995 10.6151
R10390 gnd.n2995 gnd.n2994 10.6151
R10391 gnd.n2994 gnd.n2932 10.6151
R10392 gnd.n2988 gnd.n2932 10.6151
R10393 gnd.n2988 gnd.n2987 10.6151
R10394 gnd.n2987 gnd.n2986 10.6151
R10395 gnd.n2986 gnd.n2934 10.6151
R10396 gnd.n2980 gnd.n2934 10.6151
R10397 gnd.n2980 gnd.n2979 10.6151
R10398 gnd.n2979 gnd.n2978 10.6151
R10399 gnd.n2978 gnd.n2936 10.6151
R10400 gnd.n2972 gnd.n2936 10.6151
R10401 gnd.n2972 gnd.n2971 10.6151
R10402 gnd.n2971 gnd.n2970 10.6151
R10403 gnd.n2970 gnd.n2938 10.6151
R10404 gnd.n2964 gnd.n2938 10.6151
R10405 gnd.n2964 gnd.n2963 10.6151
R10406 gnd.n2963 gnd.n2962 10.6151
R10407 gnd.n2962 gnd.n2940 10.6151
R10408 gnd.n2956 gnd.n2940 10.6151
R10409 gnd.n2956 gnd.n2955 10.6151
R10410 gnd.n2955 gnd.n2954 10.6151
R10411 gnd.n2950 gnd.n2949 10.6151
R10412 gnd.n2949 gnd.n2881 10.6151
R10413 gnd.n3685 gnd.n3515 10.6151
R10414 gnd.n3517 gnd.n3515 10.6151
R10415 gnd.n3678 gnd.n3517 10.6151
R10416 gnd.n3678 gnd.n3677 10.6151
R10417 gnd.n3677 gnd.n3676 10.6151
R10418 gnd.n3676 gnd.n3519 10.6151
R10419 gnd.n3671 gnd.n3519 10.6151
R10420 gnd.n3671 gnd.n3670 10.6151
R10421 gnd.n3670 gnd.n3669 10.6151
R10422 gnd.n3669 gnd.n3522 10.6151
R10423 gnd.n3664 gnd.n3522 10.6151
R10424 gnd.n3664 gnd.n3663 10.6151
R10425 gnd.n3663 gnd.n3662 10.6151
R10426 gnd.n3662 gnd.n3525 10.6151
R10427 gnd.n3657 gnd.n3525 10.6151
R10428 gnd.n3657 gnd.n3656 10.6151
R10429 gnd.n3656 gnd.n3655 10.6151
R10430 gnd.n3655 gnd.n3528 10.6151
R10431 gnd.n3650 gnd.n3528 10.6151
R10432 gnd.n3650 gnd.n3649 10.6151
R10433 gnd.n3649 gnd.n3648 10.6151
R10434 gnd.n3648 gnd.n3531 10.6151
R10435 gnd.n3643 gnd.n3531 10.6151
R10436 gnd.n3643 gnd.n3642 10.6151
R10437 gnd.n3642 gnd.n3641 10.6151
R10438 gnd.n3641 gnd.n3534 10.6151
R10439 gnd.n3636 gnd.n3534 10.6151
R10440 gnd.n3636 gnd.n3635 10.6151
R10441 gnd.n3633 gnd.n3539 10.6151
R10442 gnd.n3628 gnd.n3539 10.6151
R10443 gnd.n3041 gnd.n3011 10.6151
R10444 gnd.n3041 gnd.n3040 10.6151
R10445 gnd.n3040 gnd.n3039 10.6151
R10446 gnd.n3039 gnd.n3012 10.6151
R10447 gnd.n3024 gnd.n3012 10.6151
R10448 gnd.n3025 gnd.n3024 10.6151
R10449 gnd.n3026 gnd.n3025 10.6151
R10450 gnd.n3026 gnd.n2093 10.6151
R10451 gnd.n3304 gnd.n2093 10.6151
R10452 gnd.n3305 gnd.n3304 10.6151
R10453 gnd.n3306 gnd.n3305 10.6151
R10454 gnd.n3311 gnd.n3306 10.6151
R10455 gnd.n3312 gnd.n3311 10.6151
R10456 gnd.n3888 gnd.n3312 10.6151
R10457 gnd.n3888 gnd.n3887 10.6151
R10458 gnd.n3887 gnd.n3886 10.6151
R10459 gnd.n3886 gnd.n3313 10.6151
R10460 gnd.n3324 gnd.n3313 10.6151
R10461 gnd.n3325 gnd.n3324 10.6151
R10462 gnd.n3873 gnd.n3325 10.6151
R10463 gnd.n3873 gnd.n3872 10.6151
R10464 gnd.n3872 gnd.n3871 10.6151
R10465 gnd.n3871 gnd.n3326 10.6151
R10466 gnd.n3337 gnd.n3326 10.6151
R10467 gnd.n3338 gnd.n3337 10.6151
R10468 gnd.n3858 gnd.n3338 10.6151
R10469 gnd.n3858 gnd.n3857 10.6151
R10470 gnd.n3857 gnd.n3856 10.6151
R10471 gnd.n3856 gnd.n3339 10.6151
R10472 gnd.n3352 gnd.n3339 10.6151
R10473 gnd.n3353 gnd.n3352 10.6151
R10474 gnd.n3843 gnd.n3353 10.6151
R10475 gnd.n3843 gnd.n3842 10.6151
R10476 gnd.n3842 gnd.n3841 10.6151
R10477 gnd.n3841 gnd.n3354 10.6151
R10478 gnd.n3364 gnd.n3354 10.6151
R10479 gnd.n3365 gnd.n3364 10.6151
R10480 gnd.n3829 gnd.n3365 10.6151
R10481 gnd.n3829 gnd.n3828 10.6151
R10482 gnd.n3828 gnd.n3827 10.6151
R10483 gnd.n3827 gnd.n3366 10.6151
R10484 gnd.n3378 gnd.n3366 10.6151
R10485 gnd.n3379 gnd.n3378 10.6151
R10486 gnd.n3815 gnd.n3379 10.6151
R10487 gnd.n3815 gnd.n3814 10.6151
R10488 gnd.n3814 gnd.n3813 10.6151
R10489 gnd.n3813 gnd.n3380 10.6151
R10490 gnd.n3392 gnd.n3380 10.6151
R10491 gnd.n3393 gnd.n3392 10.6151
R10492 gnd.n3801 gnd.n3393 10.6151
R10493 gnd.n3801 gnd.n3800 10.6151
R10494 gnd.n3800 gnd.n3799 10.6151
R10495 gnd.n3799 gnd.n3394 10.6151
R10496 gnd.n3406 gnd.n3394 10.6151
R10497 gnd.n3407 gnd.n3406 10.6151
R10498 gnd.n3787 gnd.n3407 10.6151
R10499 gnd.n3787 gnd.n3786 10.6151
R10500 gnd.n3786 gnd.n3785 10.6151
R10501 gnd.n3785 gnd.n3408 10.6151
R10502 gnd.n3418 gnd.n3408 10.6151
R10503 gnd.n3419 gnd.n3418 10.6151
R10504 gnd.n3772 gnd.n3419 10.6151
R10505 gnd.n3772 gnd.n3771 10.6151
R10506 gnd.n3771 gnd.n3770 10.6151
R10507 gnd.n3770 gnd.n3420 10.6151
R10508 gnd.n3432 gnd.n3420 10.6151
R10509 gnd.n3758 gnd.n3432 10.6151
R10510 gnd.n3758 gnd.n3757 10.6151
R10511 gnd.n3757 gnd.n3756 10.6151
R10512 gnd.n3756 gnd.n3433 10.6151
R10513 gnd.n3446 gnd.n3433 10.6151
R10514 gnd.n3447 gnd.n3446 10.6151
R10515 gnd.n3743 gnd.n3447 10.6151
R10516 gnd.n3743 gnd.n3742 10.6151
R10517 gnd.n3742 gnd.n3741 10.6151
R10518 gnd.n3741 gnd.n3448 10.6151
R10519 gnd.n3459 gnd.n3448 10.6151
R10520 gnd.n3729 gnd.n3459 10.6151
R10521 gnd.n3729 gnd.n3728 10.6151
R10522 gnd.n3728 gnd.n3727 10.6151
R10523 gnd.n3727 gnd.n3460 10.6151
R10524 gnd.n3472 gnd.n3460 10.6151
R10525 gnd.n3473 gnd.n3472 10.6151
R10526 gnd.n3714 gnd.n3473 10.6151
R10527 gnd.n3714 gnd.n3713 10.6151
R10528 gnd.n3713 gnd.n3712 10.6151
R10529 gnd.n3712 gnd.n3474 10.6151
R10530 gnd.n3476 gnd.n3474 10.6151
R10531 gnd.n3486 gnd.n3476 10.6151
R10532 gnd.n3700 gnd.n3486 10.6151
R10533 gnd.n3700 gnd.n3699 10.6151
R10534 gnd.n3699 gnd.n3698 10.6151
R10535 gnd.n3698 gnd.n3487 10.6151
R10536 gnd.n3688 gnd.n3487 10.6151
R10537 gnd.n3688 gnd.n3687 10.6151
R10538 gnd.n5571 gnd.t17 10.5161
R10539 gnd.n5008 gnd.t19 10.5161
R10540 gnd.n6209 gnd.t13 10.5161
R10541 gnd.n3867 gnd.t303 10.5161
R10542 gnd.n4066 gnd.t187 10.5161
R10543 gnd.n6146 gnd.n6130 10.4732
R10544 gnd.n6114 gnd.n6098 10.4732
R10545 gnd.n6082 gnd.n6066 10.4732
R10546 gnd.n6051 gnd.n6035 10.4732
R10547 gnd.n6019 gnd.n6003 10.4732
R10548 gnd.n5987 gnd.n5971 10.4732
R10549 gnd.n5955 gnd.n5939 10.4732
R10550 gnd.n5924 gnd.n5908 10.4732
R10551 gnd.n3302 gnd.n3301 10.1975
R10552 gnd.n3962 gnd.n2024 10.1975
R10553 gnd.n3970 gnd.n2015 10.1975
R10554 gnd.n3782 gnd.n3781 10.1975
R10555 gnd.n3415 gnd.n1957 10.1975
R10556 gnd.n4106 gnd.n1897 10.1975
R10557 gnd.n5878 gnd.t36 9.87883
R10558 gnd.n7577 gnd.n66 9.73455
R10559 gnd.n6150 gnd.n6149 9.69747
R10560 gnd.n6118 gnd.n6117 9.69747
R10561 gnd.n6086 gnd.n6085 9.69747
R10562 gnd.n6055 gnd.n6054 9.69747
R10563 gnd.n6023 gnd.n6022 9.69747
R10564 gnd.n5991 gnd.n5990 9.69747
R10565 gnd.n5959 gnd.n5958 9.69747
R10566 gnd.n5928 gnd.n5927 9.69747
R10567 gnd.n4663 gnd.n1276 9.45751
R10568 gnd.n1722 gnd.n1503 9.45599
R10569 gnd.n6156 gnd.n6155 9.45567
R10570 gnd.n6124 gnd.n6123 9.45567
R10571 gnd.n6092 gnd.n6091 9.45567
R10572 gnd.n6061 gnd.n6060 9.45567
R10573 gnd.n6029 gnd.n6028 9.45567
R10574 gnd.n5997 gnd.n5996 9.45567
R10575 gnd.n5965 gnd.n5964 9.45567
R10576 gnd.n5934 gnd.n5933 9.45567
R10577 gnd.n5534 gnd.n5533 9.39724
R10578 gnd.n6155 gnd.n6154 9.3005
R10579 gnd.n6128 gnd.n6127 9.3005
R10580 gnd.n6149 gnd.n6148 9.3005
R10581 gnd.n6147 gnd.n6146 9.3005
R10582 gnd.n6132 gnd.n6131 9.3005
R10583 gnd.n6141 gnd.n6140 9.3005
R10584 gnd.n6139 gnd.n6138 9.3005
R10585 gnd.n6123 gnd.n6122 9.3005
R10586 gnd.n6096 gnd.n6095 9.3005
R10587 gnd.n6117 gnd.n6116 9.3005
R10588 gnd.n6115 gnd.n6114 9.3005
R10589 gnd.n6100 gnd.n6099 9.3005
R10590 gnd.n6109 gnd.n6108 9.3005
R10591 gnd.n6107 gnd.n6106 9.3005
R10592 gnd.n6091 gnd.n6090 9.3005
R10593 gnd.n6064 gnd.n6063 9.3005
R10594 gnd.n6085 gnd.n6084 9.3005
R10595 gnd.n6083 gnd.n6082 9.3005
R10596 gnd.n6068 gnd.n6067 9.3005
R10597 gnd.n6077 gnd.n6076 9.3005
R10598 gnd.n6075 gnd.n6074 9.3005
R10599 gnd.n6060 gnd.n6059 9.3005
R10600 gnd.n6033 gnd.n6032 9.3005
R10601 gnd.n6054 gnd.n6053 9.3005
R10602 gnd.n6052 gnd.n6051 9.3005
R10603 gnd.n6037 gnd.n6036 9.3005
R10604 gnd.n6046 gnd.n6045 9.3005
R10605 gnd.n6044 gnd.n6043 9.3005
R10606 gnd.n6028 gnd.n6027 9.3005
R10607 gnd.n6001 gnd.n6000 9.3005
R10608 gnd.n6022 gnd.n6021 9.3005
R10609 gnd.n6020 gnd.n6019 9.3005
R10610 gnd.n6005 gnd.n6004 9.3005
R10611 gnd.n6014 gnd.n6013 9.3005
R10612 gnd.n6012 gnd.n6011 9.3005
R10613 gnd.n5996 gnd.n5995 9.3005
R10614 gnd.n5969 gnd.n5968 9.3005
R10615 gnd.n5990 gnd.n5989 9.3005
R10616 gnd.n5988 gnd.n5987 9.3005
R10617 gnd.n5973 gnd.n5972 9.3005
R10618 gnd.n5982 gnd.n5981 9.3005
R10619 gnd.n5980 gnd.n5979 9.3005
R10620 gnd.n5964 gnd.n5963 9.3005
R10621 gnd.n5937 gnd.n5936 9.3005
R10622 gnd.n5958 gnd.n5957 9.3005
R10623 gnd.n5956 gnd.n5955 9.3005
R10624 gnd.n5941 gnd.n5940 9.3005
R10625 gnd.n5950 gnd.n5949 9.3005
R10626 gnd.n5948 gnd.n5947 9.3005
R10627 gnd.n5933 gnd.n5932 9.3005
R10628 gnd.n5906 gnd.n5905 9.3005
R10629 gnd.n5927 gnd.n5926 9.3005
R10630 gnd.n5925 gnd.n5924 9.3005
R10631 gnd.n5910 gnd.n5909 9.3005
R10632 gnd.n5919 gnd.n5918 9.3005
R10633 gnd.n5917 gnd.n5916 9.3005
R10634 gnd.n6303 gnd.n4912 9.3005
R10635 gnd.n6302 gnd.n4914 9.3005
R10636 gnd.n4918 gnd.n4915 9.3005
R10637 gnd.n6297 gnd.n4919 9.3005
R10638 gnd.n6296 gnd.n4920 9.3005
R10639 gnd.n6295 gnd.n4921 9.3005
R10640 gnd.n4925 gnd.n4922 9.3005
R10641 gnd.n6290 gnd.n4926 9.3005
R10642 gnd.n6289 gnd.n4927 9.3005
R10643 gnd.n6288 gnd.n4928 9.3005
R10644 gnd.n4932 gnd.n4929 9.3005
R10645 gnd.n6283 gnd.n4933 9.3005
R10646 gnd.n6282 gnd.n4934 9.3005
R10647 gnd.n6281 gnd.n4935 9.3005
R10648 gnd.n4940 gnd.n4938 9.3005
R10649 gnd.n6276 gnd.n6275 9.3005
R10650 gnd.n6305 gnd.n6304 9.3005
R10651 gnd.n5590 gnd.n5589 9.3005
R10652 gnd.n5208 gnd.n5207 9.3005
R10653 gnd.n5617 gnd.n5616 9.3005
R10654 gnd.n5618 gnd.n5206 9.3005
R10655 gnd.n5622 gnd.n5619 9.3005
R10656 gnd.n5621 gnd.n5620 9.3005
R10657 gnd.n5182 gnd.n5181 9.3005
R10658 gnd.n5648 gnd.n5647 9.3005
R10659 gnd.n5649 gnd.n5180 9.3005
R10660 gnd.n5653 gnd.n5650 9.3005
R10661 gnd.n5652 gnd.n5651 9.3005
R10662 gnd.n5157 gnd.n5156 9.3005
R10663 gnd.n5679 gnd.n5678 9.3005
R10664 gnd.n5680 gnd.n5155 9.3005
R10665 gnd.n5684 gnd.n5681 9.3005
R10666 gnd.n5683 gnd.n5682 9.3005
R10667 gnd.n5131 gnd.n5130 9.3005
R10668 gnd.n5710 gnd.n5709 9.3005
R10669 gnd.n5711 gnd.n5129 9.3005
R10670 gnd.n5715 gnd.n5712 9.3005
R10671 gnd.n5714 gnd.n5713 9.3005
R10672 gnd.n5107 gnd.n5106 9.3005
R10673 gnd.n5740 gnd.n5739 9.3005
R10674 gnd.n5741 gnd.n5105 9.3005
R10675 gnd.n5745 gnd.n5742 9.3005
R10676 gnd.n5744 gnd.n5743 9.3005
R10677 gnd.n5076 gnd.n5075 9.3005
R10678 gnd.n5794 gnd.n5793 9.3005
R10679 gnd.n5795 gnd.n5074 9.3005
R10680 gnd.n5797 gnd.n5796 9.3005
R10681 gnd.n5055 gnd.n5054 9.3005
R10682 gnd.n5824 gnd.n5823 9.3005
R10683 gnd.n5825 gnd.n5053 9.3005
R10684 gnd.n5829 gnd.n5826 9.3005
R10685 gnd.n5828 gnd.n5827 9.3005
R10686 gnd.n5031 gnd.n5030 9.3005
R10687 gnd.n5870 gnd.n5869 9.3005
R10688 gnd.n5871 gnd.n5029 9.3005
R10689 gnd.n5875 gnd.n5872 9.3005
R10690 gnd.n5874 gnd.n5873 9.3005
R10691 gnd.n5001 gnd.n5000 9.3005
R10692 gnd.n6191 gnd.n6190 9.3005
R10693 gnd.n6192 gnd.n4999 9.3005
R10694 gnd.n6200 gnd.n6193 9.3005
R10695 gnd.n6199 gnd.n6194 9.3005
R10696 gnd.n6198 gnd.n6196 9.3005
R10697 gnd.n6195 gnd.n913 9.3005
R10698 gnd.n6321 gnd.n914 9.3005
R10699 gnd.n6320 gnd.n915 9.3005
R10700 gnd.n6319 gnd.n916 9.3005
R10701 gnd.n4910 gnd.n917 9.3005
R10702 gnd.n4911 gnd.n4909 9.3005
R10703 gnd.n6307 gnd.n6306 9.3005
R10704 gnd.n5591 gnd.n5588 9.3005
R10705 gnd.n5287 gnd.n5246 9.3005
R10706 gnd.n5282 gnd.n5281 9.3005
R10707 gnd.n5280 gnd.n5247 9.3005
R10708 gnd.n5279 gnd.n5278 9.3005
R10709 gnd.n5275 gnd.n5248 9.3005
R10710 gnd.n5272 gnd.n5271 9.3005
R10711 gnd.n5270 gnd.n5249 9.3005
R10712 gnd.n5269 gnd.n5268 9.3005
R10713 gnd.n5265 gnd.n5250 9.3005
R10714 gnd.n5262 gnd.n5261 9.3005
R10715 gnd.n5260 gnd.n5251 9.3005
R10716 gnd.n5259 gnd.n5258 9.3005
R10717 gnd.n5255 gnd.n5253 9.3005
R10718 gnd.n5252 gnd.n5232 9.3005
R10719 gnd.n5585 gnd.n5231 9.3005
R10720 gnd.n5587 gnd.n5586 9.3005
R10721 gnd.n5289 gnd.n5288 9.3005
R10722 gnd.n5598 gnd.n5218 9.3005
R10723 gnd.n5605 gnd.n5219 9.3005
R10724 gnd.n5607 gnd.n5606 9.3005
R10725 gnd.n5608 gnd.n5199 9.3005
R10726 gnd.n5627 gnd.n5626 9.3005
R10727 gnd.n5629 gnd.n5192 9.3005
R10728 gnd.n5636 gnd.n5193 9.3005
R10729 gnd.n5638 gnd.n5637 9.3005
R10730 gnd.n5639 gnd.n5175 9.3005
R10731 gnd.n5658 gnd.n5657 9.3005
R10732 gnd.n5660 gnd.n5167 9.3005
R10733 gnd.n5667 gnd.n5168 9.3005
R10734 gnd.n5669 gnd.n5668 9.3005
R10735 gnd.n5670 gnd.n5149 9.3005
R10736 gnd.n5689 gnd.n5688 9.3005
R10737 gnd.n5691 gnd.n5141 9.3005
R10738 gnd.n5698 gnd.n5142 9.3005
R10739 gnd.n5700 gnd.n5699 9.3005
R10740 gnd.n5701 gnd.n5124 9.3005
R10741 gnd.n5720 gnd.n5719 9.3005
R10742 gnd.n5722 gnd.n5116 9.3005
R10743 gnd.n5729 gnd.n5117 9.3005
R10744 gnd.n5731 gnd.n5730 9.3005
R10745 gnd.n5732 gnd.n5100 9.3005
R10746 gnd.n5750 gnd.n5749 9.3005
R10747 gnd.n5752 gnd.n5085 9.3005
R10748 gnd.n5783 gnd.n5087 9.3005
R10749 gnd.n5784 gnd.n5083 9.3005
R10750 gnd.n5786 gnd.n5785 9.3005
R10751 gnd.n5071 gnd.n5066 9.3005
R10752 gnd.n5807 gnd.n5065 9.3005
R10753 gnd.n5810 gnd.n5809 9.3005
R10754 gnd.n5812 gnd.n5811 9.3005
R10755 gnd.n5815 gnd.n5048 9.3005
R10756 gnd.n5813 gnd.n5046 9.3005
R10757 gnd.n5837 gnd.n5044 9.3005
R10758 gnd.n5839 gnd.n5838 9.3005
R10759 gnd.n5022 gnd.n5021 9.3005
R10760 gnd.n5884 gnd.n5883 9.3005
R10761 gnd.n5885 gnd.n5015 9.3005
R10762 gnd.n5893 gnd.n5014 9.3005
R10763 gnd.n5896 gnd.n5895 9.3005
R10764 gnd.n5898 gnd.n5012 9.3005
R10765 gnd.n6182 gnd.n6181 9.3005
R10766 gnd.n6180 gnd.n5899 9.3005
R10767 gnd.n5901 gnd.n5900 9.3005
R10768 gnd.n6176 gnd.n5902 9.3005
R10769 gnd.n6175 gnd.n5903 9.3005
R10770 gnd.n6174 gnd.n6161 9.3005
R10771 gnd.n6171 gnd.n6163 9.3005
R10772 gnd.n6170 gnd.n6164 9.3005
R10773 gnd.n6167 gnd.n6165 9.3005
R10774 gnd.n6166 gnd.n4941 9.3005
R10775 gnd.n5596 gnd.n5595 9.3005
R10776 gnd.n6271 gnd.n4942 9.3005
R10777 gnd.n6270 gnd.n4944 9.3005
R10778 gnd.n4948 gnd.n4945 9.3005
R10779 gnd.n6265 gnd.n4949 9.3005
R10780 gnd.n6264 gnd.n4950 9.3005
R10781 gnd.n6263 gnd.n4951 9.3005
R10782 gnd.n4955 gnd.n4952 9.3005
R10783 gnd.n6258 gnd.n4956 9.3005
R10784 gnd.n6257 gnd.n4957 9.3005
R10785 gnd.n6256 gnd.n4958 9.3005
R10786 gnd.n4962 gnd.n4959 9.3005
R10787 gnd.n6251 gnd.n4963 9.3005
R10788 gnd.n6250 gnd.n4964 9.3005
R10789 gnd.n6249 gnd.n4965 9.3005
R10790 gnd.n4969 gnd.n4966 9.3005
R10791 gnd.n6244 gnd.n4970 9.3005
R10792 gnd.n6243 gnd.n4971 9.3005
R10793 gnd.n6242 gnd.n4972 9.3005
R10794 gnd.n4976 gnd.n4973 9.3005
R10795 gnd.n6237 gnd.n4977 9.3005
R10796 gnd.n6236 gnd.n4978 9.3005
R10797 gnd.n6235 gnd.n4979 9.3005
R10798 gnd.n4986 gnd.n4984 9.3005
R10799 gnd.n6230 gnd.n4987 9.3005
R10800 gnd.n6229 gnd.n4988 9.3005
R10801 gnd.n6228 gnd.n6225 9.3005
R10802 gnd.n6273 gnd.n6272 9.3005
R10803 gnd.n5093 gnd.n5092 9.3005
R10804 gnd.n5760 gnd.n5759 9.3005
R10805 gnd.n5761 gnd.n5091 9.3005
R10806 gnd.n5778 gnd.n5762 9.3005
R10807 gnd.n5777 gnd.n5763 9.3005
R10808 gnd.n5776 gnd.n5764 9.3005
R10809 gnd.n5774 gnd.n5765 9.3005
R10810 gnd.n5773 gnd.n5766 9.3005
R10811 gnd.n5771 gnd.n5767 9.3005
R10812 gnd.n5770 gnd.n5768 9.3005
R10813 gnd.n5037 gnd.n5036 9.3005
R10814 gnd.n5847 gnd.n5846 9.3005
R10815 gnd.n5848 gnd.n5035 9.3005
R10816 gnd.n5862 gnd.n5849 9.3005
R10817 gnd.n5861 gnd.n5850 9.3005
R10818 gnd.n5860 gnd.n5851 9.3005
R10819 gnd.n5858 gnd.n5852 9.3005
R10820 gnd.n5857 gnd.n5853 9.3005
R10821 gnd.n5855 gnd.n5854 9.3005
R10822 gnd.n4994 gnd.n4993 9.3005
R10823 gnd.n6206 gnd.n6205 9.3005
R10824 gnd.n6207 gnd.n4992 9.3005
R10825 gnd.n6211 gnd.n6208 9.3005
R10826 gnd.n6212 gnd.n4991 9.3005
R10827 gnd.n6216 gnd.n6215 9.3005
R10828 gnd.n6217 gnd.n4990 9.3005
R10829 gnd.n6219 gnd.n6218 9.3005
R10830 gnd.n6222 gnd.n4989 9.3005
R10831 gnd.n6224 gnd.n6223 9.3005
R10832 gnd.n5420 gnd.n5419 9.3005
R10833 gnd.n5310 gnd.n5309 9.3005
R10834 gnd.n5434 gnd.n5433 9.3005
R10835 gnd.n5435 gnd.n5308 9.3005
R10836 gnd.n5437 gnd.n5436 9.3005
R10837 gnd.n5298 gnd.n5297 9.3005
R10838 gnd.n5450 gnd.n5449 9.3005
R10839 gnd.n5451 gnd.n5296 9.3005
R10840 gnd.n5569 gnd.n5452 9.3005
R10841 gnd.n5568 gnd.n5453 9.3005
R10842 gnd.n5567 gnd.n5454 9.3005
R10843 gnd.n5566 gnd.n5455 9.3005
R10844 gnd.n5563 gnd.n5456 9.3005
R10845 gnd.n5562 gnd.n5457 9.3005
R10846 gnd.n5561 gnd.n5458 9.3005
R10847 gnd.n5559 gnd.n5459 9.3005
R10848 gnd.n5558 gnd.n5460 9.3005
R10849 gnd.n5555 gnd.n5461 9.3005
R10850 gnd.n5554 gnd.n5462 9.3005
R10851 gnd.n5553 gnd.n5463 9.3005
R10852 gnd.n5551 gnd.n5464 9.3005
R10853 gnd.n5550 gnd.n5465 9.3005
R10854 gnd.n5546 gnd.n5466 9.3005
R10855 gnd.n5545 gnd.n5467 9.3005
R10856 gnd.n5544 gnd.n5468 9.3005
R10857 gnd.n5542 gnd.n5469 9.3005
R10858 gnd.n5541 gnd.n5470 9.3005
R10859 gnd.n5538 gnd.n5471 9.3005
R10860 gnd.n5418 gnd.n5319 9.3005
R10861 gnd.n5321 gnd.n5320 9.3005
R10862 gnd.n5365 gnd.n5363 9.3005
R10863 gnd.n5366 gnd.n5362 9.3005
R10864 gnd.n5369 gnd.n5358 9.3005
R10865 gnd.n5370 gnd.n5357 9.3005
R10866 gnd.n5373 gnd.n5356 9.3005
R10867 gnd.n5374 gnd.n5355 9.3005
R10868 gnd.n5377 gnd.n5354 9.3005
R10869 gnd.n5378 gnd.n5353 9.3005
R10870 gnd.n5381 gnd.n5352 9.3005
R10871 gnd.n5382 gnd.n5351 9.3005
R10872 gnd.n5385 gnd.n5350 9.3005
R10873 gnd.n5386 gnd.n5349 9.3005
R10874 gnd.n5389 gnd.n5348 9.3005
R10875 gnd.n5390 gnd.n5347 9.3005
R10876 gnd.n5393 gnd.n5346 9.3005
R10877 gnd.n5394 gnd.n5345 9.3005
R10878 gnd.n5397 gnd.n5344 9.3005
R10879 gnd.n5398 gnd.n5343 9.3005
R10880 gnd.n5401 gnd.n5342 9.3005
R10881 gnd.n5402 gnd.n5341 9.3005
R10882 gnd.n5405 gnd.n5340 9.3005
R10883 gnd.n5407 gnd.n5339 9.3005
R10884 gnd.n5408 gnd.n5338 9.3005
R10885 gnd.n5409 gnd.n5337 9.3005
R10886 gnd.n5410 gnd.n5336 9.3005
R10887 gnd.n5417 gnd.n5416 9.3005
R10888 gnd.n5426 gnd.n5425 9.3005
R10889 gnd.n5427 gnd.n5313 9.3005
R10890 gnd.n5429 gnd.n5428 9.3005
R10891 gnd.n5304 gnd.n5303 9.3005
R10892 gnd.n5442 gnd.n5441 9.3005
R10893 gnd.n5443 gnd.n5302 9.3005
R10894 gnd.n5445 gnd.n5444 9.3005
R10895 gnd.n5291 gnd.n5290 9.3005
R10896 gnd.n5574 gnd.n5573 9.3005
R10897 gnd.n5575 gnd.n5245 9.3005
R10898 gnd.n5579 gnd.n5577 9.3005
R10899 gnd.n5578 gnd.n5224 9.3005
R10900 gnd.n5597 gnd.n5223 9.3005
R10901 gnd.n5600 gnd.n5599 9.3005
R10902 gnd.n5217 gnd.n5216 9.3005
R10903 gnd.n5611 gnd.n5609 9.3005
R10904 gnd.n5610 gnd.n5198 9.3005
R10905 gnd.n5628 gnd.n5197 9.3005
R10906 gnd.n5631 gnd.n5630 9.3005
R10907 gnd.n5191 gnd.n5190 9.3005
R10908 gnd.n5642 gnd.n5640 9.3005
R10909 gnd.n5641 gnd.n5174 9.3005
R10910 gnd.n5659 gnd.n5173 9.3005
R10911 gnd.n5662 gnd.n5661 9.3005
R10912 gnd.n5166 gnd.n5165 9.3005
R10913 gnd.n5673 gnd.n5671 9.3005
R10914 gnd.n5672 gnd.n5148 9.3005
R10915 gnd.n5690 gnd.n5147 9.3005
R10916 gnd.n5693 gnd.n5692 9.3005
R10917 gnd.n5140 gnd.n5139 9.3005
R10918 gnd.n5704 gnd.n5702 9.3005
R10919 gnd.n5703 gnd.n5123 9.3005
R10920 gnd.n5721 gnd.n5122 9.3005
R10921 gnd.n5724 gnd.n5723 9.3005
R10922 gnd.n5115 gnd.n5114 9.3005
R10923 gnd.n5734 gnd.n5733 9.3005
R10924 gnd.n5099 gnd.n5098 9.3005
R10925 gnd.n5755 gnd.n5751 9.3005
R10926 gnd.n5754 gnd.n5753 9.3005
R10927 gnd.n5086 gnd.n5082 9.3005
R10928 gnd.n5788 gnd.n5787 9.3005
R10929 gnd.n5084 gnd.n5067 9.3005
R10930 gnd.n5806 gnd.n5805 9.3005
R10931 gnd.n5808 gnd.n5063 9.3005
R10932 gnd.n5818 gnd.n5064 9.3005
R10933 gnd.n5817 gnd.n5816 9.3005
R10934 gnd.n5814 gnd.n5042 9.3005
R10935 gnd.n5842 gnd.n5043 9.3005
R10936 gnd.n5841 gnd.n5840 9.3005
R10937 gnd.n5045 gnd.n5023 9.3005
R10938 gnd.n5881 gnd.n5880 9.3005
R10939 gnd.n5882 gnd.n5016 9.3005
R10940 gnd.n5892 gnd.n5891 9.3005
R10941 gnd.n5894 gnd.n5010 9.3005
R10942 gnd.n6185 gnd.n5011 9.3005
R10943 gnd.n6184 gnd.n6183 9.3005
R10944 gnd.n5013 gnd.n901 9.3005
R10945 gnd.n6328 gnd.n902 9.3005
R10946 gnd.n6327 gnd.n903 9.3005
R10947 gnd.n6326 gnd.n904 9.3005
R10948 gnd.n6160 gnd.n905 9.3005
R10949 gnd.n6162 gnd.n925 9.3005
R10950 gnd.n6314 gnd.n926 9.3005
R10951 gnd.n6313 gnd.n927 9.3005
R10952 gnd.n6312 gnd.n928 9.3005
R10953 gnd.n5315 gnd.n5314 9.3005
R10954 gnd.n6503 gnd.n6502 9.3005
R10955 gnd.n6504 gnd.n725 9.3005
R10956 gnd.n6506 gnd.n6505 9.3005
R10957 gnd.n721 gnd.n720 9.3005
R10958 gnd.n6513 gnd.n6512 9.3005
R10959 gnd.n6514 gnd.n719 9.3005
R10960 gnd.n6516 gnd.n6515 9.3005
R10961 gnd.n715 gnd.n714 9.3005
R10962 gnd.n6523 gnd.n6522 9.3005
R10963 gnd.n6524 gnd.n713 9.3005
R10964 gnd.n6526 gnd.n6525 9.3005
R10965 gnd.n709 gnd.n708 9.3005
R10966 gnd.n6533 gnd.n6532 9.3005
R10967 gnd.n6534 gnd.n707 9.3005
R10968 gnd.n6536 gnd.n6535 9.3005
R10969 gnd.n703 gnd.n702 9.3005
R10970 gnd.n6543 gnd.n6542 9.3005
R10971 gnd.n6544 gnd.n701 9.3005
R10972 gnd.n6546 gnd.n6545 9.3005
R10973 gnd.n697 gnd.n696 9.3005
R10974 gnd.n6553 gnd.n6552 9.3005
R10975 gnd.n6554 gnd.n695 9.3005
R10976 gnd.n6556 gnd.n6555 9.3005
R10977 gnd.n691 gnd.n690 9.3005
R10978 gnd.n6563 gnd.n6562 9.3005
R10979 gnd.n6564 gnd.n689 9.3005
R10980 gnd.n6566 gnd.n6565 9.3005
R10981 gnd.n685 gnd.n684 9.3005
R10982 gnd.n6573 gnd.n6572 9.3005
R10983 gnd.n6574 gnd.n683 9.3005
R10984 gnd.n6576 gnd.n6575 9.3005
R10985 gnd.n679 gnd.n678 9.3005
R10986 gnd.n6583 gnd.n6582 9.3005
R10987 gnd.n6584 gnd.n677 9.3005
R10988 gnd.n6586 gnd.n6585 9.3005
R10989 gnd.n673 gnd.n672 9.3005
R10990 gnd.n6593 gnd.n6592 9.3005
R10991 gnd.n6594 gnd.n671 9.3005
R10992 gnd.n6596 gnd.n6595 9.3005
R10993 gnd.n667 gnd.n666 9.3005
R10994 gnd.n6603 gnd.n6602 9.3005
R10995 gnd.n6604 gnd.n665 9.3005
R10996 gnd.n6606 gnd.n6605 9.3005
R10997 gnd.n661 gnd.n660 9.3005
R10998 gnd.n6613 gnd.n6612 9.3005
R10999 gnd.n6614 gnd.n659 9.3005
R11000 gnd.n6616 gnd.n6615 9.3005
R11001 gnd.n655 gnd.n654 9.3005
R11002 gnd.n6623 gnd.n6622 9.3005
R11003 gnd.n6624 gnd.n653 9.3005
R11004 gnd.n6626 gnd.n6625 9.3005
R11005 gnd.n649 gnd.n648 9.3005
R11006 gnd.n6633 gnd.n6632 9.3005
R11007 gnd.n6634 gnd.n647 9.3005
R11008 gnd.n6636 gnd.n6635 9.3005
R11009 gnd.n643 gnd.n642 9.3005
R11010 gnd.n6643 gnd.n6642 9.3005
R11011 gnd.n6644 gnd.n641 9.3005
R11012 gnd.n6646 gnd.n6645 9.3005
R11013 gnd.n637 gnd.n636 9.3005
R11014 gnd.n6653 gnd.n6652 9.3005
R11015 gnd.n6654 gnd.n635 9.3005
R11016 gnd.n6656 gnd.n6655 9.3005
R11017 gnd.n631 gnd.n630 9.3005
R11018 gnd.n6663 gnd.n6662 9.3005
R11019 gnd.n6664 gnd.n629 9.3005
R11020 gnd.n6666 gnd.n6665 9.3005
R11021 gnd.n625 gnd.n624 9.3005
R11022 gnd.n6673 gnd.n6672 9.3005
R11023 gnd.n6674 gnd.n623 9.3005
R11024 gnd.n6676 gnd.n6675 9.3005
R11025 gnd.n619 gnd.n618 9.3005
R11026 gnd.n6683 gnd.n6682 9.3005
R11027 gnd.n6684 gnd.n617 9.3005
R11028 gnd.n6686 gnd.n6685 9.3005
R11029 gnd.n613 gnd.n612 9.3005
R11030 gnd.n6693 gnd.n6692 9.3005
R11031 gnd.n6694 gnd.n611 9.3005
R11032 gnd.n6696 gnd.n6695 9.3005
R11033 gnd.n607 gnd.n606 9.3005
R11034 gnd.n6703 gnd.n6702 9.3005
R11035 gnd.n6704 gnd.n605 9.3005
R11036 gnd.n6706 gnd.n6705 9.3005
R11037 gnd.n601 gnd.n600 9.3005
R11038 gnd.n6713 gnd.n6712 9.3005
R11039 gnd.n6714 gnd.n599 9.3005
R11040 gnd.n6716 gnd.n6715 9.3005
R11041 gnd.n595 gnd.n594 9.3005
R11042 gnd.n6723 gnd.n6722 9.3005
R11043 gnd.n6724 gnd.n593 9.3005
R11044 gnd.n6726 gnd.n6725 9.3005
R11045 gnd.n589 gnd.n588 9.3005
R11046 gnd.n6733 gnd.n6732 9.3005
R11047 gnd.n6734 gnd.n587 9.3005
R11048 gnd.n6736 gnd.n6735 9.3005
R11049 gnd.n583 gnd.n582 9.3005
R11050 gnd.n6743 gnd.n6742 9.3005
R11051 gnd.n6744 gnd.n581 9.3005
R11052 gnd.n6746 gnd.n6745 9.3005
R11053 gnd.n577 gnd.n576 9.3005
R11054 gnd.n6753 gnd.n6752 9.3005
R11055 gnd.n6754 gnd.n575 9.3005
R11056 gnd.n6756 gnd.n6755 9.3005
R11057 gnd.n571 gnd.n570 9.3005
R11058 gnd.n6763 gnd.n6762 9.3005
R11059 gnd.n6764 gnd.n569 9.3005
R11060 gnd.n6766 gnd.n6765 9.3005
R11061 gnd.n565 gnd.n564 9.3005
R11062 gnd.n6773 gnd.n6772 9.3005
R11063 gnd.n6774 gnd.n563 9.3005
R11064 gnd.n6776 gnd.n6775 9.3005
R11065 gnd.n559 gnd.n558 9.3005
R11066 gnd.n6783 gnd.n6782 9.3005
R11067 gnd.n6784 gnd.n557 9.3005
R11068 gnd.n6786 gnd.n6785 9.3005
R11069 gnd.n553 gnd.n552 9.3005
R11070 gnd.n6793 gnd.n6792 9.3005
R11071 gnd.n6794 gnd.n551 9.3005
R11072 gnd.n6796 gnd.n6795 9.3005
R11073 gnd.n547 gnd.n546 9.3005
R11074 gnd.n6803 gnd.n6802 9.3005
R11075 gnd.n6804 gnd.n545 9.3005
R11076 gnd.n6806 gnd.n6805 9.3005
R11077 gnd.n541 gnd.n540 9.3005
R11078 gnd.n6813 gnd.n6812 9.3005
R11079 gnd.n6814 gnd.n539 9.3005
R11080 gnd.n6816 gnd.n6815 9.3005
R11081 gnd.n535 gnd.n534 9.3005
R11082 gnd.n6823 gnd.n6822 9.3005
R11083 gnd.n6824 gnd.n533 9.3005
R11084 gnd.n6826 gnd.n6825 9.3005
R11085 gnd.n529 gnd.n528 9.3005
R11086 gnd.n6833 gnd.n6832 9.3005
R11087 gnd.n6834 gnd.n527 9.3005
R11088 gnd.n6836 gnd.n6835 9.3005
R11089 gnd.n523 gnd.n522 9.3005
R11090 gnd.n6843 gnd.n6842 9.3005
R11091 gnd.n6844 gnd.n521 9.3005
R11092 gnd.n6846 gnd.n6845 9.3005
R11093 gnd.n517 gnd.n516 9.3005
R11094 gnd.n6853 gnd.n6852 9.3005
R11095 gnd.n6854 gnd.n515 9.3005
R11096 gnd.n6856 gnd.n6855 9.3005
R11097 gnd.n511 gnd.n510 9.3005
R11098 gnd.n6863 gnd.n6862 9.3005
R11099 gnd.n6864 gnd.n509 9.3005
R11100 gnd.n6866 gnd.n6865 9.3005
R11101 gnd.n505 gnd.n504 9.3005
R11102 gnd.n6873 gnd.n6872 9.3005
R11103 gnd.n6874 gnd.n503 9.3005
R11104 gnd.n6876 gnd.n6875 9.3005
R11105 gnd.n499 gnd.n498 9.3005
R11106 gnd.n6883 gnd.n6882 9.3005
R11107 gnd.n6884 gnd.n497 9.3005
R11108 gnd.n6886 gnd.n6885 9.3005
R11109 gnd.n493 gnd.n492 9.3005
R11110 gnd.n6893 gnd.n6892 9.3005
R11111 gnd.n6894 gnd.n491 9.3005
R11112 gnd.n6896 gnd.n6895 9.3005
R11113 gnd.n487 gnd.n486 9.3005
R11114 gnd.n6903 gnd.n6902 9.3005
R11115 gnd.n6904 gnd.n485 9.3005
R11116 gnd.n6906 gnd.n6905 9.3005
R11117 gnd.n481 gnd.n480 9.3005
R11118 gnd.n6913 gnd.n6912 9.3005
R11119 gnd.n6914 gnd.n479 9.3005
R11120 gnd.n6916 gnd.n6915 9.3005
R11121 gnd.n475 gnd.n474 9.3005
R11122 gnd.n6923 gnd.n6922 9.3005
R11123 gnd.n6924 gnd.n473 9.3005
R11124 gnd.n6926 gnd.n6925 9.3005
R11125 gnd.n469 gnd.n468 9.3005
R11126 gnd.n6933 gnd.n6932 9.3005
R11127 gnd.n6934 gnd.n467 9.3005
R11128 gnd.n6936 gnd.n6935 9.3005
R11129 gnd.n463 gnd.n462 9.3005
R11130 gnd.n6943 gnd.n6942 9.3005
R11131 gnd.n6944 gnd.n461 9.3005
R11132 gnd.n6947 gnd.n6946 9.3005
R11133 gnd.n6945 gnd.n457 9.3005
R11134 gnd.n6953 gnd.n456 9.3005
R11135 gnd.n6955 gnd.n6954 9.3005
R11136 gnd.n452 gnd.n451 9.3005
R11137 gnd.n6964 gnd.n6963 9.3005
R11138 gnd.n6965 gnd.n450 9.3005
R11139 gnd.n6967 gnd.n6966 9.3005
R11140 gnd.n446 gnd.n445 9.3005
R11141 gnd.n6974 gnd.n6973 9.3005
R11142 gnd.n6975 gnd.n444 9.3005
R11143 gnd.n6977 gnd.n6976 9.3005
R11144 gnd.n440 gnd.n439 9.3005
R11145 gnd.n6984 gnd.n6983 9.3005
R11146 gnd.n6985 gnd.n438 9.3005
R11147 gnd.n6987 gnd.n6986 9.3005
R11148 gnd.n434 gnd.n433 9.3005
R11149 gnd.n6994 gnd.n6993 9.3005
R11150 gnd.n6995 gnd.n432 9.3005
R11151 gnd.n6997 gnd.n6996 9.3005
R11152 gnd.n428 gnd.n427 9.3005
R11153 gnd.n7004 gnd.n7003 9.3005
R11154 gnd.n7005 gnd.n426 9.3005
R11155 gnd.n7007 gnd.n7006 9.3005
R11156 gnd.n422 gnd.n421 9.3005
R11157 gnd.n7014 gnd.n7013 9.3005
R11158 gnd.n7015 gnd.n420 9.3005
R11159 gnd.n7017 gnd.n7016 9.3005
R11160 gnd.n416 gnd.n415 9.3005
R11161 gnd.n7024 gnd.n7023 9.3005
R11162 gnd.n7025 gnd.n414 9.3005
R11163 gnd.n7027 gnd.n7026 9.3005
R11164 gnd.n410 gnd.n409 9.3005
R11165 gnd.n7034 gnd.n7033 9.3005
R11166 gnd.n7035 gnd.n408 9.3005
R11167 gnd.n7037 gnd.n7036 9.3005
R11168 gnd.n404 gnd.n403 9.3005
R11169 gnd.n7044 gnd.n7043 9.3005
R11170 gnd.n7045 gnd.n402 9.3005
R11171 gnd.n7047 gnd.n7046 9.3005
R11172 gnd.n398 gnd.n397 9.3005
R11173 gnd.n7054 gnd.n7053 9.3005
R11174 gnd.n7055 gnd.n396 9.3005
R11175 gnd.n7057 gnd.n7056 9.3005
R11176 gnd.n392 gnd.n391 9.3005
R11177 gnd.n7064 gnd.n7063 9.3005
R11178 gnd.n7065 gnd.n390 9.3005
R11179 gnd.n7067 gnd.n7066 9.3005
R11180 gnd.n386 gnd.n385 9.3005
R11181 gnd.n7074 gnd.n7073 9.3005
R11182 gnd.n7075 gnd.n384 9.3005
R11183 gnd.n7077 gnd.n7076 9.3005
R11184 gnd.n380 gnd.n379 9.3005
R11185 gnd.n7084 gnd.n7083 9.3005
R11186 gnd.n7085 gnd.n378 9.3005
R11187 gnd.n7087 gnd.n7086 9.3005
R11188 gnd.n374 gnd.n373 9.3005
R11189 gnd.n7094 gnd.n7093 9.3005
R11190 gnd.n7095 gnd.n372 9.3005
R11191 gnd.n7097 gnd.n7096 9.3005
R11192 gnd.n368 gnd.n367 9.3005
R11193 gnd.n7104 gnd.n7103 9.3005
R11194 gnd.n7105 gnd.n366 9.3005
R11195 gnd.n7107 gnd.n7106 9.3005
R11196 gnd.n362 gnd.n361 9.3005
R11197 gnd.n7114 gnd.n7113 9.3005
R11198 gnd.n7115 gnd.n360 9.3005
R11199 gnd.n7117 gnd.n7116 9.3005
R11200 gnd.n356 gnd.n355 9.3005
R11201 gnd.n7124 gnd.n7123 9.3005
R11202 gnd.n7125 gnd.n354 9.3005
R11203 gnd.n7127 gnd.n7126 9.3005
R11204 gnd.n350 gnd.n349 9.3005
R11205 gnd.n7134 gnd.n7133 9.3005
R11206 gnd.n7135 gnd.n348 9.3005
R11207 gnd.n7137 gnd.n7136 9.3005
R11208 gnd.n344 gnd.n343 9.3005
R11209 gnd.n7144 gnd.n7143 9.3005
R11210 gnd.n7145 gnd.n342 9.3005
R11211 gnd.n7147 gnd.n7146 9.3005
R11212 gnd.n338 gnd.n337 9.3005
R11213 gnd.n7154 gnd.n7153 9.3005
R11214 gnd.n7155 gnd.n336 9.3005
R11215 gnd.n7157 gnd.n7156 9.3005
R11216 gnd.n332 gnd.n331 9.3005
R11217 gnd.n7165 gnd.n7164 9.3005
R11218 gnd.n7166 gnd.n330 9.3005
R11219 gnd.n7169 gnd.n7168 9.3005
R11220 gnd.n6957 gnd.n6956 9.3005
R11221 gnd.n7528 gnd.n112 9.3005
R11222 gnd.n7527 gnd.n114 9.3005
R11223 gnd.n118 gnd.n115 9.3005
R11224 gnd.n7522 gnd.n119 9.3005
R11225 gnd.n7521 gnd.n120 9.3005
R11226 gnd.n7520 gnd.n121 9.3005
R11227 gnd.n125 gnd.n122 9.3005
R11228 gnd.n7515 gnd.n126 9.3005
R11229 gnd.n7514 gnd.n127 9.3005
R11230 gnd.n7513 gnd.n128 9.3005
R11231 gnd.n132 gnd.n129 9.3005
R11232 gnd.n7508 gnd.n133 9.3005
R11233 gnd.n7507 gnd.n134 9.3005
R11234 gnd.n7506 gnd.n135 9.3005
R11235 gnd.n139 gnd.n136 9.3005
R11236 gnd.n7501 gnd.n140 9.3005
R11237 gnd.n7500 gnd.n141 9.3005
R11238 gnd.n7496 gnd.n142 9.3005
R11239 gnd.n146 gnd.n143 9.3005
R11240 gnd.n7491 gnd.n147 9.3005
R11241 gnd.n7490 gnd.n148 9.3005
R11242 gnd.n7489 gnd.n149 9.3005
R11243 gnd.n153 gnd.n150 9.3005
R11244 gnd.n7484 gnd.n154 9.3005
R11245 gnd.n7483 gnd.n155 9.3005
R11246 gnd.n7482 gnd.n156 9.3005
R11247 gnd.n160 gnd.n157 9.3005
R11248 gnd.n7477 gnd.n161 9.3005
R11249 gnd.n7476 gnd.n162 9.3005
R11250 gnd.n7475 gnd.n163 9.3005
R11251 gnd.n167 gnd.n164 9.3005
R11252 gnd.n7470 gnd.n168 9.3005
R11253 gnd.n7469 gnd.n169 9.3005
R11254 gnd.n7468 gnd.n170 9.3005
R11255 gnd.n174 gnd.n171 9.3005
R11256 gnd.n7463 gnd.n175 9.3005
R11257 gnd.n7462 gnd.n7461 9.3005
R11258 gnd.n7460 gnd.n178 9.3005
R11259 gnd.n7530 gnd.n7529 9.3005
R11260 gnd.n1649 gnd.n1648 9.3005
R11261 gnd.n1678 gnd.n1650 9.3005
R11262 gnd.n1677 gnd.n1651 9.3005
R11263 gnd.n1676 gnd.n1652 9.3005
R11264 gnd.n1674 gnd.n1653 9.3005
R11265 gnd.n1673 gnd.n1654 9.3005
R11266 gnd.n1670 gnd.n1655 9.3005
R11267 gnd.n1669 gnd.n1656 9.3005
R11268 gnd.n1668 gnd.n1657 9.3005
R11269 gnd.n1666 gnd.n1658 9.3005
R11270 gnd.n1665 gnd.n1659 9.3005
R11271 gnd.n1663 gnd.n1660 9.3005
R11272 gnd.n1662 gnd.n1661 9.3005
R11273 gnd.n1558 gnd.n1557 9.3005
R11274 gnd.n4329 gnd.n4328 9.3005
R11275 gnd.n4330 gnd.n1556 9.3005
R11276 gnd.n4332 gnd.n4331 9.3005
R11277 gnd.n4333 gnd.n1555 9.3005
R11278 gnd.n4336 gnd.n4335 9.3005
R11279 gnd.n4337 gnd.n1554 9.3005
R11280 gnd.n4347 gnd.n4338 9.3005
R11281 gnd.n4346 gnd.n4339 9.3005
R11282 gnd.n4345 gnd.n4340 9.3005
R11283 gnd.n4344 gnd.n4342 9.3005
R11284 gnd.n4341 gnd.n299 9.3005
R11285 gnd.n7207 gnd.n300 9.3005
R11286 gnd.n7209 gnd.n7208 9.3005
R11287 gnd.n7269 gnd.n7210 9.3005
R11288 gnd.n7268 gnd.n7211 9.3005
R11289 gnd.n7267 gnd.n7212 9.3005
R11290 gnd.n7263 gnd.n7213 9.3005
R11291 gnd.n7262 gnd.n7214 9.3005
R11292 gnd.n7259 gnd.n7215 9.3005
R11293 gnd.n7258 gnd.n7216 9.3005
R11294 gnd.n7256 gnd.n7217 9.3005
R11295 gnd.n7255 gnd.n7218 9.3005
R11296 gnd.n7253 gnd.n7219 9.3005
R11297 gnd.n7252 gnd.n7220 9.3005
R11298 gnd.n7250 gnd.n7221 9.3005
R11299 gnd.n7249 gnd.n7222 9.3005
R11300 gnd.n7247 gnd.n7223 9.3005
R11301 gnd.n7246 gnd.n7224 9.3005
R11302 gnd.n7244 gnd.n7225 9.3005
R11303 gnd.n7243 gnd.n7226 9.3005
R11304 gnd.n7241 gnd.n7227 9.3005
R11305 gnd.n7240 gnd.n7228 9.3005
R11306 gnd.n7238 gnd.n7229 9.3005
R11307 gnd.n7237 gnd.n7230 9.3005
R11308 gnd.n7235 gnd.n7231 9.3005
R11309 gnd.n7234 gnd.n7233 9.3005
R11310 gnd.n7232 gnd.n182 9.3005
R11311 gnd.n7457 gnd.n181 9.3005
R11312 gnd.n7459 gnd.n7458 9.3005
R11313 gnd.n1496 gnd.n1494 9.3005
R11314 gnd.n4429 gnd.n4428 9.3005
R11315 gnd.n4430 gnd.n1488 9.3005
R11316 gnd.n4433 gnd.n1487 9.3005
R11317 gnd.n4434 gnd.n1486 9.3005
R11318 gnd.n4437 gnd.n1485 9.3005
R11319 gnd.n4438 gnd.n1484 9.3005
R11320 gnd.n4441 gnd.n1483 9.3005
R11321 gnd.n4442 gnd.n1482 9.3005
R11322 gnd.n4445 gnd.n1481 9.3005
R11323 gnd.n4446 gnd.n1480 9.3005
R11324 gnd.n4449 gnd.n1479 9.3005
R11325 gnd.n4450 gnd.n1478 9.3005
R11326 gnd.n4453 gnd.n1477 9.3005
R11327 gnd.n4454 gnd.n1476 9.3005
R11328 gnd.n4457 gnd.n1475 9.3005
R11329 gnd.n4458 gnd.n1474 9.3005
R11330 gnd.n4461 gnd.n1473 9.3005
R11331 gnd.n4462 gnd.n1472 9.3005
R11332 gnd.n4465 gnd.n1471 9.3005
R11333 gnd.n4467 gnd.n1465 9.3005
R11334 gnd.n4470 gnd.n1464 9.3005
R11335 gnd.n4471 gnd.n1463 9.3005
R11336 gnd.n4474 gnd.n1462 9.3005
R11337 gnd.n4475 gnd.n1461 9.3005
R11338 gnd.n4478 gnd.n1460 9.3005
R11339 gnd.n4479 gnd.n1459 9.3005
R11340 gnd.n4482 gnd.n1458 9.3005
R11341 gnd.n4483 gnd.n1457 9.3005
R11342 gnd.n4486 gnd.n1456 9.3005
R11343 gnd.n4487 gnd.n1455 9.3005
R11344 gnd.n4490 gnd.n1454 9.3005
R11345 gnd.n4492 gnd.n1453 9.3005
R11346 gnd.n4493 gnd.n1452 9.3005
R11347 gnd.n4494 gnd.n1451 9.3005
R11348 gnd.n4495 gnd.n1450 9.3005
R11349 gnd.n4427 gnd.n1493 9.3005
R11350 gnd.n4426 gnd.n4425 9.3005
R11351 gnd.n1645 gnd.n1644 9.3005
R11352 gnd.n1623 gnd.n1622 9.3005
R11353 gnd.n4251 gnd.n4250 9.3005
R11354 gnd.n4252 gnd.n1621 9.3005
R11355 gnd.n4256 gnd.n4253 9.3005
R11356 gnd.n4255 gnd.n4254 9.3005
R11357 gnd.n1595 gnd.n1594 9.3005
R11358 gnd.n4282 gnd.n4281 9.3005
R11359 gnd.n4283 gnd.n1593 9.3005
R11360 gnd.n4287 gnd.n4284 9.3005
R11361 gnd.n4286 gnd.n4285 9.3005
R11362 gnd.n1568 gnd.n1567 9.3005
R11363 gnd.n4319 gnd.n4318 9.3005
R11364 gnd.n4320 gnd.n1566 9.3005
R11365 gnd.n4324 gnd.n4321 9.3005
R11366 gnd.n4323 gnd.n4322 9.3005
R11367 gnd.n1533 gnd.n1532 9.3005
R11368 gnd.n4382 gnd.n4381 9.3005
R11369 gnd.n4383 gnd.n1531 9.3005
R11370 gnd.n4385 gnd.n4384 9.3005
R11371 gnd.n275 gnd.n268 9.3005
R11372 gnd.n254 gnd.n253 9.3005
R11373 gnd.n7310 gnd.n7309 9.3005
R11374 gnd.n7311 gnd.n252 9.3005
R11375 gnd.n7313 gnd.n7312 9.3005
R11376 gnd.n236 gnd.n235 9.3005
R11377 gnd.n7326 gnd.n7325 9.3005
R11378 gnd.n7327 gnd.n234 9.3005
R11379 gnd.n7329 gnd.n7328 9.3005
R11380 gnd.n223 gnd.n222 9.3005
R11381 gnd.n7342 gnd.n7341 9.3005
R11382 gnd.n7343 gnd.n221 9.3005
R11383 gnd.n7345 gnd.n7344 9.3005
R11384 gnd.n206 gnd.n205 9.3005
R11385 gnd.n7358 gnd.n7357 9.3005
R11386 gnd.n7359 gnd.n204 9.3005
R11387 gnd.n7361 gnd.n7360 9.3005
R11388 gnd.n191 gnd.n190 9.3005
R11389 gnd.n7449 gnd.n7448 9.3005
R11390 gnd.n7450 gnd.n189 9.3005
R11391 gnd.n7452 gnd.n7451 9.3005
R11392 gnd.n111 gnd.n110 9.3005
R11393 gnd.n7532 gnd.n7531 9.3005
R11394 gnd.n1643 gnd.n1642 9.3005
R11395 gnd.n7296 gnd.n273 9.3005
R11396 gnd.n7297 gnd.n7296 9.3005
R11397 gnd.n2400 gnd.n2399 9.3005
R11398 gnd.n2384 gnd.n2383 9.3005
R11399 gnd.n2395 gnd.n2386 9.3005
R11400 gnd.n2394 gnd.n2387 9.3005
R11401 gnd.n2393 gnd.n2388 9.3005
R11402 gnd.n2391 gnd.n2390 9.3005
R11403 gnd.n2389 gnd.n2353 9.3005
R11404 gnd.n2351 gnd.n2350 9.3005
R11405 gnd.n2729 gnd.n2728 9.3005
R11406 gnd.n2730 gnd.n2349 9.3005
R11407 gnd.n2732 gnd.n2731 9.3005
R11408 gnd.n2347 gnd.n2346 9.3005
R11409 gnd.n2737 gnd.n2736 9.3005
R11410 gnd.n2738 gnd.n2345 9.3005
R11411 gnd.n2773 gnd.n2739 9.3005
R11412 gnd.n2772 gnd.n2740 9.3005
R11413 gnd.n2771 gnd.n2741 9.3005
R11414 gnd.n2744 gnd.n2742 9.3005
R11415 gnd.n2767 gnd.n2745 9.3005
R11416 gnd.n2766 gnd.n2746 9.3005
R11417 gnd.n2765 gnd.n2747 9.3005
R11418 gnd.n2750 gnd.n2748 9.3005
R11419 gnd.n2761 gnd.n2751 9.3005
R11420 gnd.n2760 gnd.n2752 9.3005
R11421 gnd.n2759 gnd.n2753 9.3005
R11422 gnd.n2755 gnd.n2754 9.3005
R11423 gnd.n2173 gnd.n2172 9.3005
R11424 gnd.n3205 gnd.n3204 9.3005
R11425 gnd.n3206 gnd.n2171 9.3005
R11426 gnd.n3208 gnd.n3207 9.3005
R11427 gnd.n2161 gnd.n2160 9.3005
R11428 gnd.n3221 gnd.n3220 9.3005
R11429 gnd.n3222 gnd.n2159 9.3005
R11430 gnd.n3224 gnd.n3223 9.3005
R11431 gnd.n2148 gnd.n2147 9.3005
R11432 gnd.n3237 gnd.n3236 9.3005
R11433 gnd.n3238 gnd.n2146 9.3005
R11434 gnd.n3240 gnd.n3239 9.3005
R11435 gnd.n2135 gnd.n2134 9.3005
R11436 gnd.n3253 gnd.n3252 9.3005
R11437 gnd.n3254 gnd.n2133 9.3005
R11438 gnd.n3256 gnd.n3255 9.3005
R11439 gnd.n2120 gnd.n2119 9.3005
R11440 gnd.n3269 gnd.n3268 9.3005
R11441 gnd.n3270 gnd.n2118 9.3005
R11442 gnd.n3272 gnd.n3271 9.3005
R11443 gnd.n2108 gnd.n2107 9.3005
R11444 gnd.n3285 gnd.n3284 9.3005
R11445 gnd.n3286 gnd.n2106 9.3005
R11446 gnd.n3290 gnd.n3287 9.3005
R11447 gnd.n3289 gnd.n3288 9.3005
R11448 gnd.n2080 gnd.n2079 9.3005
R11449 gnd.n3901 gnd.n3900 9.3005
R11450 gnd.n3902 gnd.n2078 9.3005
R11451 gnd.n3904 gnd.n3903 9.3005
R11452 gnd.n2065 gnd.n2064 9.3005
R11453 gnd.n3917 gnd.n3916 9.3005
R11454 gnd.n3918 gnd.n2063 9.3005
R11455 gnd.n3920 gnd.n3919 9.3005
R11456 gnd.n2050 gnd.n2049 9.3005
R11457 gnd.n3933 gnd.n3932 9.3005
R11458 gnd.n3934 gnd.n2048 9.3005
R11459 gnd.n3936 gnd.n3935 9.3005
R11460 gnd.n2035 gnd.n2034 9.3005
R11461 gnd.n3949 gnd.n3948 9.3005
R11462 gnd.n3950 gnd.n2033 9.3005
R11463 gnd.n3952 gnd.n3951 9.3005
R11464 gnd.n2021 gnd.n2020 9.3005
R11465 gnd.n3965 gnd.n3964 9.3005
R11466 gnd.n3966 gnd.n2019 9.3005
R11467 gnd.n3968 gnd.n3967 9.3005
R11468 gnd.n2006 gnd.n2005 9.3005
R11469 gnd.n3981 gnd.n3980 9.3005
R11470 gnd.n3982 gnd.n2004 9.3005
R11471 gnd.n3984 gnd.n3983 9.3005
R11472 gnd.n1991 gnd.n1990 9.3005
R11473 gnd.n3997 gnd.n3996 9.3005
R11474 gnd.n3998 gnd.n1989 9.3005
R11475 gnd.n4000 gnd.n3999 9.3005
R11476 gnd.n1976 gnd.n1975 9.3005
R11477 gnd.n4013 gnd.n4012 9.3005
R11478 gnd.n4014 gnd.n1974 9.3005
R11479 gnd.n4016 gnd.n4015 9.3005
R11480 gnd.n1962 gnd.n1961 9.3005
R11481 gnd.n4029 gnd.n4028 9.3005
R11482 gnd.n4030 gnd.n1960 9.3005
R11483 gnd.n4032 gnd.n4031 9.3005
R11484 gnd.n1947 gnd.n1946 9.3005
R11485 gnd.n4045 gnd.n4044 9.3005
R11486 gnd.n4046 gnd.n1945 9.3005
R11487 gnd.n4048 gnd.n4047 9.3005
R11488 gnd.n1934 gnd.n1933 9.3005
R11489 gnd.n4061 gnd.n4060 9.3005
R11490 gnd.n4062 gnd.n1932 9.3005
R11491 gnd.n4064 gnd.n4063 9.3005
R11492 gnd.n1922 gnd.n1921 9.3005
R11493 gnd.n4077 gnd.n4076 9.3005
R11494 gnd.n4078 gnd.n1920 9.3005
R11495 gnd.n4080 gnd.n4079 9.3005
R11496 gnd.n1909 gnd.n1908 9.3005
R11497 gnd.n4093 gnd.n4092 9.3005
R11498 gnd.n4094 gnd.n1907 9.3005
R11499 gnd.n4096 gnd.n4095 9.3005
R11500 gnd.n1895 gnd.n1894 9.3005
R11501 gnd.n4109 gnd.n4108 9.3005
R11502 gnd.n4110 gnd.n1893 9.3005
R11503 gnd.n4112 gnd.n4111 9.3005
R11504 gnd.n1882 gnd.n1881 9.3005
R11505 gnd.n4125 gnd.n4124 9.3005
R11506 gnd.n4126 gnd.n1880 9.3005
R11507 gnd.n4128 gnd.n4127 9.3005
R11508 gnd.n1869 gnd.n1868 9.3005
R11509 gnd.n4141 gnd.n4140 9.3005
R11510 gnd.n4142 gnd.n1867 9.3005
R11511 gnd.n4144 gnd.n4143 9.3005
R11512 gnd.n1856 gnd.n1855 9.3005
R11513 gnd.n4157 gnd.n4156 9.3005
R11514 gnd.n4158 gnd.n1854 9.3005
R11515 gnd.n4160 gnd.n4159 9.3005
R11516 gnd.n1842 gnd.n1841 9.3005
R11517 gnd.n4173 gnd.n4172 9.3005
R11518 gnd.n4174 gnd.n1840 9.3005
R11519 gnd.n4176 gnd.n4175 9.3005
R11520 gnd.n1829 gnd.n1828 9.3005
R11521 gnd.n4191 gnd.n4190 9.3005
R11522 gnd.n4192 gnd.n1827 9.3005
R11523 gnd.n4197 gnd.n4193 9.3005
R11524 gnd.n4196 gnd.n4195 9.3005
R11525 gnd.n4194 gnd.n1411 9.3005
R11526 gnd.n4504 gnd.n1412 9.3005
R11527 gnd.n4503 gnd.n1413 9.3005
R11528 gnd.n4502 gnd.n1414 9.3005
R11529 gnd.n1636 gnd.n1415 9.3005
R11530 gnd.n1637 gnd.n1635 9.3005
R11531 gnd.n1639 gnd.n1638 9.3005
R11532 gnd.n1633 gnd.n1632 9.3005
R11533 gnd.n4240 gnd.n4239 9.3005
R11534 gnd.n4241 gnd.n1631 9.3005
R11535 gnd.n4245 gnd.n4242 9.3005
R11536 gnd.n4244 gnd.n4243 9.3005
R11537 gnd.n1606 gnd.n1605 9.3005
R11538 gnd.n4271 gnd.n4270 9.3005
R11539 gnd.n4272 gnd.n1604 9.3005
R11540 gnd.n4276 gnd.n4273 9.3005
R11541 gnd.n4275 gnd.n4274 9.3005
R11542 gnd.n1578 gnd.n1577 9.3005
R11543 gnd.n4307 gnd.n4306 9.3005
R11544 gnd.n4308 gnd.n1576 9.3005
R11545 gnd.n4312 gnd.n4309 9.3005
R11546 gnd.n4311 gnd.n4310 9.3005
R11547 gnd.n1544 gnd.n1543 9.3005
R11548 gnd.n4365 gnd.n4364 9.3005
R11549 gnd.n4366 gnd.n1542 9.3005
R11550 gnd.n4376 gnd.n4367 9.3005
R11551 gnd.n4375 gnd.n4368 9.3005
R11552 gnd.n4374 gnd.n4369 9.3005
R11553 gnd.n7175 gnd.n326 9.3005
R11554 gnd.n7174 gnd.n327 9.3005
R11555 gnd.n7167 gnd.n328 9.3005
R11556 gnd.n3115 gnd.n2303 9.3005
R11557 gnd.n3118 gnd.n2302 9.3005
R11558 gnd.n3119 gnd.n2301 9.3005
R11559 gnd.n3122 gnd.n2300 9.3005
R11560 gnd.n3123 gnd.n2299 9.3005
R11561 gnd.n3126 gnd.n2298 9.3005
R11562 gnd.n3127 gnd.n2297 9.3005
R11563 gnd.n3130 gnd.n2296 9.3005
R11564 gnd.n3131 gnd.n2295 9.3005
R11565 gnd.n3134 gnd.n2294 9.3005
R11566 gnd.n3135 gnd.n2293 9.3005
R11567 gnd.n3138 gnd.n2292 9.3005
R11568 gnd.n3139 gnd.n2291 9.3005
R11569 gnd.n3140 gnd.n2290 9.3005
R11570 gnd.n2289 gnd.n2286 9.3005
R11571 gnd.n2288 gnd.n2287 9.3005
R11572 gnd.n2877 gnd.n2876 9.3005
R11573 gnd.n2873 gnd.n2308 9.3005
R11574 gnd.n2870 gnd.n2309 9.3005
R11575 gnd.n2869 gnd.n2310 9.3005
R11576 gnd.n2866 gnd.n2311 9.3005
R11577 gnd.n2865 gnd.n2312 9.3005
R11578 gnd.n2862 gnd.n2313 9.3005
R11579 gnd.n2861 gnd.n2314 9.3005
R11580 gnd.n2858 gnd.n2315 9.3005
R11581 gnd.n2857 gnd.n2316 9.3005
R11582 gnd.n2854 gnd.n2317 9.3005
R11583 gnd.n2853 gnd.n2318 9.3005
R11584 gnd.n2850 gnd.n2319 9.3005
R11585 gnd.n2849 gnd.n2320 9.3005
R11586 gnd.n2846 gnd.n2321 9.3005
R11587 gnd.n2845 gnd.n2322 9.3005
R11588 gnd.n2842 gnd.n2323 9.3005
R11589 gnd.n2841 gnd.n2324 9.3005
R11590 gnd.n2838 gnd.n2837 9.3005
R11591 gnd.n2836 gnd.n2326 9.3005
R11592 gnd.n2878 gnd.n2304 9.3005
R11593 gnd.n2470 gnd.n2469 9.3005
R11594 gnd.n2554 gnd.n2553 9.3005
R11595 gnd.n2555 gnd.n2468 9.3005
R11596 gnd.n2558 gnd.n2556 9.3005
R11597 gnd.n2559 gnd.n2467 9.3005
R11598 gnd.n2562 gnd.n2561 9.3005
R11599 gnd.n2563 gnd.n2466 9.3005
R11600 gnd.n2566 gnd.n2564 9.3005
R11601 gnd.n2567 gnd.n2465 9.3005
R11602 gnd.n2570 gnd.n2569 9.3005
R11603 gnd.n2571 gnd.n2464 9.3005
R11604 gnd.n2574 gnd.n2572 9.3005
R11605 gnd.n2575 gnd.n2463 9.3005
R11606 gnd.n2578 gnd.n2577 9.3005
R11607 gnd.n2579 gnd.n2462 9.3005
R11608 gnd.n2582 gnd.n2580 9.3005
R11609 gnd.n2583 gnd.n2461 9.3005
R11610 gnd.n2586 gnd.n2585 9.3005
R11611 gnd.n2587 gnd.n2460 9.3005
R11612 gnd.n2590 gnd.n2589 9.3005
R11613 gnd.n2588 gnd.n2415 9.3005
R11614 gnd.n2646 gnd.n2416 9.3005
R11615 gnd.n2645 gnd.n2417 9.3005
R11616 gnd.n2644 gnd.n2418 9.3005
R11617 gnd.n2615 gnd.n2419 9.3005
R11618 gnd.n2634 gnd.n2616 9.3005
R11619 gnd.n2496 gnd.n2495 9.3005
R11620 gnd.n2501 gnd.n2500 9.3005
R11621 gnd.n2504 gnd.n2490 9.3005
R11622 gnd.n2505 gnd.n2489 9.3005
R11623 gnd.n2508 gnd.n2488 9.3005
R11624 gnd.n2509 gnd.n2487 9.3005
R11625 gnd.n2512 gnd.n2486 9.3005
R11626 gnd.n2513 gnd.n2485 9.3005
R11627 gnd.n2516 gnd.n2484 9.3005
R11628 gnd.n2517 gnd.n2483 9.3005
R11629 gnd.n2520 gnd.n2482 9.3005
R11630 gnd.n2521 gnd.n2481 9.3005
R11631 gnd.n2524 gnd.n2480 9.3005
R11632 gnd.n2525 gnd.n2479 9.3005
R11633 gnd.n2528 gnd.n2478 9.3005
R11634 gnd.n2529 gnd.n2477 9.3005
R11635 gnd.n2532 gnd.n2476 9.3005
R11636 gnd.n2535 gnd.n2534 9.3005
R11637 gnd.n2499 gnd.n2494 9.3005
R11638 gnd.n2498 gnd.n2497 9.3005
R11639 gnd.n2542 gnd.n2541 9.3005
R11640 gnd.n2540 gnd.n2475 9.3005
R11641 gnd.n2539 gnd.n2538 9.3005
R11642 gnd.n2537 gnd.n1032 9.3005
R11643 gnd.n4810 gnd.n1033 9.3005
R11644 gnd.n4809 gnd.n1034 9.3005
R11645 gnd.n4808 gnd.n1035 9.3005
R11646 gnd.n1051 gnd.n1036 9.3005
R11647 gnd.n4798 gnd.n1052 9.3005
R11648 gnd.n4797 gnd.n1053 9.3005
R11649 gnd.n4796 gnd.n1054 9.3005
R11650 gnd.n1072 gnd.n1055 9.3005
R11651 gnd.n4786 gnd.n1073 9.3005
R11652 gnd.n4785 gnd.n1074 9.3005
R11653 gnd.n4784 gnd.n1075 9.3005
R11654 gnd.n1091 gnd.n1076 9.3005
R11655 gnd.n4774 gnd.n1092 9.3005
R11656 gnd.n4773 gnd.n1093 9.3005
R11657 gnd.n4772 gnd.n1094 9.3005
R11658 gnd.n1114 gnd.n1095 9.3005
R11659 gnd.n4762 gnd.n1115 9.3005
R11660 gnd.n4761 gnd.n1116 9.3005
R11661 gnd.n4760 gnd.n1117 9.3005
R11662 gnd.n1132 gnd.n1118 9.3005
R11663 gnd.n4750 gnd.n1133 9.3005
R11664 gnd.n4749 gnd.n1134 9.3005
R11665 gnd.n4748 gnd.n1135 9.3005
R11666 gnd.n1151 gnd.n1136 9.3005
R11667 gnd.n4737 gnd.n1152 9.3005
R11668 gnd.n4736 gnd.n1153 9.3005
R11669 gnd.n4735 gnd.n1154 9.3005
R11670 gnd.n1170 gnd.n1155 9.3005
R11671 gnd.n4725 gnd.n1171 9.3005
R11672 gnd.n4724 gnd.n1172 9.3005
R11673 gnd.n4723 gnd.n1173 9.3005
R11674 gnd.n1192 gnd.n1174 9.3005
R11675 gnd.n4713 gnd.n1193 9.3005
R11676 gnd.n4712 gnd.n1194 9.3005
R11677 gnd.n4711 gnd.n1195 9.3005
R11678 gnd.n1212 gnd.n1196 9.3005
R11679 gnd.n4701 gnd.n1213 9.3005
R11680 gnd.n4700 gnd.n1214 9.3005
R11681 gnd.n4699 gnd.n1215 9.3005
R11682 gnd.n1234 gnd.n1216 9.3005
R11683 gnd.n4689 gnd.n1235 9.3005
R11684 gnd.n4688 gnd.n1236 9.3005
R11685 gnd.n4687 gnd.n1237 9.3005
R11686 gnd.n1255 gnd.n1238 9.3005
R11687 gnd.n4677 gnd.n1256 9.3005
R11688 gnd.n4676 gnd.n1257 9.3005
R11689 gnd.n4675 gnd.n1258 9.3005
R11690 gnd.n1275 gnd.n1259 9.3005
R11691 gnd.n4665 gnd.n4664 9.3005
R11692 gnd.n2536 gnd.n2474 9.3005
R11693 gnd.n4824 gnd.n4823 9.3005
R11694 gnd.n4822 gnd.n1010 9.3005
R11695 gnd.n4821 gnd.n4820 9.3005
R11696 gnd.n1012 gnd.n1011 9.3005
R11697 gnd.n2430 gnd.n2429 9.3005
R11698 gnd.n2433 gnd.n2432 9.3005
R11699 gnd.n2434 gnd.n2428 9.3005
R11700 gnd.n2437 gnd.n2435 9.3005
R11701 gnd.n2438 gnd.n2427 9.3005
R11702 gnd.n2441 gnd.n2440 9.3005
R11703 gnd.n2442 gnd.n2426 9.3005
R11704 gnd.n2445 gnd.n2443 9.3005
R11705 gnd.n2446 gnd.n2425 9.3005
R11706 gnd.n2449 gnd.n2448 9.3005
R11707 gnd.n2450 gnd.n2424 9.3005
R11708 gnd.n2453 gnd.n2451 9.3005
R11709 gnd.n2454 gnd.n2423 9.3005
R11710 gnd.n2457 gnd.n2456 9.3005
R11711 gnd.n2458 gnd.n2422 9.3005
R11712 gnd.n2594 gnd.n2459 9.3005
R11713 gnd.n2595 gnd.n2421 9.3005
R11714 gnd.n2597 gnd.n2596 9.3005
R11715 gnd.n2598 gnd.n2420 9.3005
R11716 gnd.n2640 gnd.n2599 9.3005
R11717 gnd.n2639 gnd.n2600 9.3005
R11718 gnd.n2638 gnd.n2601 9.3005
R11719 gnd.n2619 gnd.n2602 9.3005
R11720 gnd.n2625 gnd.n2620 9.3005
R11721 gnd.n2624 gnd.n2621 9.3005
R11722 gnd.n2623 gnd.n2622 9.3005
R11723 gnd.n2374 gnd.n2373 9.3005
R11724 gnd.n2670 gnd.n2669 9.3005
R11725 gnd.n2671 gnd.n2372 9.3005
R11726 gnd.n2674 gnd.n2673 9.3005
R11727 gnd.n2672 gnd.n2366 9.3005
R11728 gnd.n2686 gnd.n2367 9.3005
R11729 gnd.n2687 gnd.n2365 9.3005
R11730 gnd.n2689 gnd.n2688 9.3005
R11731 gnd.n2690 gnd.n2364 9.3005
R11732 gnd.n2694 gnd.n2691 9.3005
R11733 gnd.n2695 gnd.n2363 9.3005
R11734 gnd.n2700 gnd.n2699 9.3005
R11735 gnd.n2701 gnd.n2362 9.3005
R11736 gnd.n2707 gnd.n2702 9.3005
R11737 gnd.n2706 gnd.n2703 9.3005
R11738 gnd.n2705 gnd.n2704 9.3005
R11739 gnd.n2338 gnd.n2337 9.3005
R11740 gnd.n2787 gnd.n2786 9.3005
R11741 gnd.n2788 gnd.n2336 9.3005
R11742 gnd.n2791 gnd.n2790 9.3005
R11743 gnd.n2789 gnd.n2330 9.3005
R11744 gnd.n2833 gnd.n2329 9.3005
R11745 gnd.n2835 gnd.n2834 9.3005
R11746 gnd.n4825 gnd.n1008 9.3005
R11747 gnd.n4832 gnd.n4831 9.3005
R11748 gnd.n4833 gnd.n1002 9.3005
R11749 gnd.n4836 gnd.n1001 9.3005
R11750 gnd.n4837 gnd.n1000 9.3005
R11751 gnd.n4840 gnd.n999 9.3005
R11752 gnd.n4841 gnd.n998 9.3005
R11753 gnd.n4844 gnd.n997 9.3005
R11754 gnd.n4845 gnd.n996 9.3005
R11755 gnd.n4848 gnd.n995 9.3005
R11756 gnd.n4849 gnd.n994 9.3005
R11757 gnd.n4852 gnd.n993 9.3005
R11758 gnd.n4853 gnd.n992 9.3005
R11759 gnd.n4856 gnd.n991 9.3005
R11760 gnd.n4857 gnd.n990 9.3005
R11761 gnd.n4860 gnd.n989 9.3005
R11762 gnd.n4861 gnd.n988 9.3005
R11763 gnd.n4864 gnd.n987 9.3005
R11764 gnd.n4865 gnd.n986 9.3005
R11765 gnd.n4868 gnd.n985 9.3005
R11766 gnd.n4870 gnd.n982 9.3005
R11767 gnd.n4873 gnd.n981 9.3005
R11768 gnd.n4874 gnd.n980 9.3005
R11769 gnd.n4877 gnd.n979 9.3005
R11770 gnd.n4878 gnd.n978 9.3005
R11771 gnd.n4881 gnd.n977 9.3005
R11772 gnd.n4882 gnd.n976 9.3005
R11773 gnd.n4885 gnd.n975 9.3005
R11774 gnd.n4886 gnd.n974 9.3005
R11775 gnd.n4889 gnd.n973 9.3005
R11776 gnd.n4890 gnd.n972 9.3005
R11777 gnd.n4893 gnd.n971 9.3005
R11778 gnd.n4894 gnd.n970 9.3005
R11779 gnd.n4897 gnd.n969 9.3005
R11780 gnd.n4899 gnd.n968 9.3005
R11781 gnd.n4900 gnd.n967 9.3005
R11782 gnd.n4901 gnd.n966 9.3005
R11783 gnd.n4902 gnd.n965 9.3005
R11784 gnd.n4830 gnd.n1007 9.3005
R11785 gnd.n4829 gnd.n4828 9.3005
R11786 gnd.n2548 gnd.n2547 9.3005
R11787 gnd.n2546 gnd.n1021 9.3005
R11788 gnd.n4816 gnd.n1022 9.3005
R11789 gnd.n4815 gnd.n1023 9.3005
R11790 gnd.n4814 gnd.n1024 9.3005
R11791 gnd.n1042 gnd.n1025 9.3005
R11792 gnd.n4804 gnd.n1043 9.3005
R11793 gnd.n4803 gnd.n1044 9.3005
R11794 gnd.n4802 gnd.n1045 9.3005
R11795 gnd.n1061 gnd.n1046 9.3005
R11796 gnd.n4792 gnd.n1062 9.3005
R11797 gnd.n4791 gnd.n1063 9.3005
R11798 gnd.n4790 gnd.n1064 9.3005
R11799 gnd.n1082 gnd.n1065 9.3005
R11800 gnd.n4780 gnd.n1083 9.3005
R11801 gnd.n4779 gnd.n1084 9.3005
R11802 gnd.n4778 gnd.n1085 9.3005
R11803 gnd.n1103 gnd.n1086 9.3005
R11804 gnd.n4768 gnd.n1104 9.3005
R11805 gnd.n4767 gnd.n1105 9.3005
R11806 gnd.n4766 gnd.n1106 9.3005
R11807 gnd.n4730 gnd.n1162 9.3005
R11808 gnd.n4729 gnd.n1163 9.3005
R11809 gnd.n1181 gnd.n1164 9.3005
R11810 gnd.n4719 gnd.n1182 9.3005
R11811 gnd.n4718 gnd.n1183 9.3005
R11812 gnd.n4717 gnd.n1184 9.3005
R11813 gnd.n1202 gnd.n1185 9.3005
R11814 gnd.n4707 gnd.n1203 9.3005
R11815 gnd.n4706 gnd.n1204 9.3005
R11816 gnd.n4705 gnd.n1205 9.3005
R11817 gnd.n1223 gnd.n1206 9.3005
R11818 gnd.n4695 gnd.n1224 9.3005
R11819 gnd.n4694 gnd.n1225 9.3005
R11820 gnd.n4693 gnd.n1226 9.3005
R11821 gnd.n1244 gnd.n1227 9.3005
R11822 gnd.n4683 gnd.n1245 9.3005
R11823 gnd.n4682 gnd.n1246 9.3005
R11824 gnd.n4681 gnd.n1247 9.3005
R11825 gnd.n1265 gnd.n1248 9.3005
R11826 gnd.n4671 gnd.n1266 9.3005
R11827 gnd.n4670 gnd.n1267 9.3005
R11828 gnd.n4669 gnd.n1268 9.3005
R11829 gnd.n2545 gnd.n2544 9.3005
R11830 gnd.n4755 gnd.n1125 9.3005
R11831 gnd.n4731 gnd.n1125 9.3005
R11832 gnd.n2406 gnd.n2405 9.3005
R11833 gnd.n2653 gnd.n2652 9.3005
R11834 gnd.n2410 gnd.n2409 9.3005
R11835 gnd.n6334 gnd.n893 9.3005
R11836 gnd.n6335 gnd.n892 9.3005
R11837 gnd.n6336 gnd.n891 9.3005
R11838 gnd.n890 gnd.n886 9.3005
R11839 gnd.n6342 gnd.n885 9.3005
R11840 gnd.n6343 gnd.n884 9.3005
R11841 gnd.n6344 gnd.n883 9.3005
R11842 gnd.n882 gnd.n878 9.3005
R11843 gnd.n6350 gnd.n877 9.3005
R11844 gnd.n6351 gnd.n876 9.3005
R11845 gnd.n6352 gnd.n875 9.3005
R11846 gnd.n874 gnd.n870 9.3005
R11847 gnd.n6358 gnd.n869 9.3005
R11848 gnd.n6359 gnd.n868 9.3005
R11849 gnd.n6360 gnd.n867 9.3005
R11850 gnd.n866 gnd.n862 9.3005
R11851 gnd.n6366 gnd.n861 9.3005
R11852 gnd.n6367 gnd.n860 9.3005
R11853 gnd.n6368 gnd.n859 9.3005
R11854 gnd.n858 gnd.n854 9.3005
R11855 gnd.n6374 gnd.n853 9.3005
R11856 gnd.n6375 gnd.n852 9.3005
R11857 gnd.n6376 gnd.n851 9.3005
R11858 gnd.n850 gnd.n846 9.3005
R11859 gnd.n6382 gnd.n845 9.3005
R11860 gnd.n6383 gnd.n844 9.3005
R11861 gnd.n6384 gnd.n843 9.3005
R11862 gnd.n842 gnd.n838 9.3005
R11863 gnd.n6390 gnd.n837 9.3005
R11864 gnd.n6391 gnd.n836 9.3005
R11865 gnd.n6392 gnd.n835 9.3005
R11866 gnd.n834 gnd.n830 9.3005
R11867 gnd.n6398 gnd.n829 9.3005
R11868 gnd.n6399 gnd.n828 9.3005
R11869 gnd.n6400 gnd.n827 9.3005
R11870 gnd.n826 gnd.n822 9.3005
R11871 gnd.n6406 gnd.n821 9.3005
R11872 gnd.n6407 gnd.n820 9.3005
R11873 gnd.n6408 gnd.n819 9.3005
R11874 gnd.n818 gnd.n814 9.3005
R11875 gnd.n6414 gnd.n813 9.3005
R11876 gnd.n6415 gnd.n812 9.3005
R11877 gnd.n6416 gnd.n811 9.3005
R11878 gnd.n810 gnd.n806 9.3005
R11879 gnd.n6422 gnd.n805 9.3005
R11880 gnd.n6423 gnd.n804 9.3005
R11881 gnd.n6424 gnd.n803 9.3005
R11882 gnd.n802 gnd.n798 9.3005
R11883 gnd.n6430 gnd.n797 9.3005
R11884 gnd.n6431 gnd.n796 9.3005
R11885 gnd.n6432 gnd.n795 9.3005
R11886 gnd.n794 gnd.n790 9.3005
R11887 gnd.n6438 gnd.n789 9.3005
R11888 gnd.n6439 gnd.n788 9.3005
R11889 gnd.n6440 gnd.n787 9.3005
R11890 gnd.n786 gnd.n782 9.3005
R11891 gnd.n6446 gnd.n781 9.3005
R11892 gnd.n6447 gnd.n780 9.3005
R11893 gnd.n6448 gnd.n779 9.3005
R11894 gnd.n778 gnd.n774 9.3005
R11895 gnd.n6454 gnd.n773 9.3005
R11896 gnd.n6455 gnd.n772 9.3005
R11897 gnd.n6456 gnd.n771 9.3005
R11898 gnd.n770 gnd.n766 9.3005
R11899 gnd.n6462 gnd.n765 9.3005
R11900 gnd.n6463 gnd.n764 9.3005
R11901 gnd.n6464 gnd.n763 9.3005
R11902 gnd.n762 gnd.n758 9.3005
R11903 gnd.n6470 gnd.n757 9.3005
R11904 gnd.n6471 gnd.n756 9.3005
R11905 gnd.n6472 gnd.n755 9.3005
R11906 gnd.n754 gnd.n750 9.3005
R11907 gnd.n6478 gnd.n749 9.3005
R11908 gnd.n6479 gnd.n748 9.3005
R11909 gnd.n6480 gnd.n747 9.3005
R11910 gnd.n746 gnd.n742 9.3005
R11911 gnd.n6486 gnd.n741 9.3005
R11912 gnd.n6487 gnd.n740 9.3005
R11913 gnd.n6488 gnd.n739 9.3005
R11914 gnd.n738 gnd.n734 9.3005
R11915 gnd.n6494 gnd.n733 9.3005
R11916 gnd.n6495 gnd.n732 9.3005
R11917 gnd.n6496 gnd.n731 9.3005
R11918 gnd.n730 gnd.n726 9.3005
R11919 gnd.n2408 gnd.n894 9.3005
R11920 gnd.n1735 gnd.n1734 9.3005
R11921 gnd.n1721 gnd.n1717 9.3005
R11922 gnd.n1742 gnd.n1741 9.3005
R11923 gnd.n1743 gnd.n1712 9.3005
R11924 gnd.n1754 gnd.n1753 9.3005
R11925 gnd.n1714 gnd.n1710 9.3005
R11926 gnd.n1761 gnd.n1760 9.3005
R11927 gnd.n1762 gnd.n1705 9.3005
R11928 gnd.n1773 gnd.n1772 9.3005
R11929 gnd.n1707 gnd.n1703 9.3005
R11930 gnd.n1780 gnd.n1779 9.3005
R11931 gnd.n1700 gnd.n1699 9.3005
R11932 gnd.n1789 gnd.n1788 9.3005
R11933 gnd.n1697 gnd.n1696 9.3005
R11934 gnd.n1796 gnd.n1795 9.3005
R11935 gnd.n1688 gnd.n1687 9.3005
R11936 gnd.n1803 gnd.n1802 9.3005
R11937 gnd.n1685 gnd.n1683 9.3005
R11938 gnd.n1724 gnd.n1719 9.3005
R11939 gnd.n1798 gnd.n1797 9.3005
R11940 gnd.n1787 gnd.n1693 9.3005
R11941 gnd.n1786 gnd.n1785 9.3005
R11942 gnd.n1782 gnd.n1781 9.3005
R11943 gnd.n1702 gnd.n1701 9.3005
R11944 gnd.n1771 gnd.n1770 9.3005
R11945 gnd.n1767 gnd.n1706 9.3005
R11946 gnd.n1764 gnd.n1763 9.3005
R11947 gnd.n1709 gnd.n1708 9.3005
R11948 gnd.n1752 gnd.n1751 9.3005
R11949 gnd.n1748 gnd.n1713 9.3005
R11950 gnd.n1745 gnd.n1744 9.3005
R11951 gnd.n1716 gnd.n1715 9.3005
R11952 gnd.n1733 gnd.n1732 9.3005
R11953 gnd.n1729 gnd.n1720 9.3005
R11954 gnd.n1726 gnd.n1725 9.3005
R11955 gnd.n1799 gnd.n1689 9.3005
R11956 gnd.n1801 gnd.n1800 9.3005
R11957 gnd.n4227 gnd.n4226 9.3005
R11958 gnd.n4225 gnd.n1684 9.3005
R11959 gnd.n4224 gnd.n4223 9.3005
R11960 gnd.n4222 gnd.n1811 9.3005
R11961 gnd.n4221 gnd.n4220 9.3005
R11962 gnd.n4219 gnd.n1812 9.3005
R11963 gnd.n4215 gnd.n4214 9.3005
R11964 gnd.n4213 gnd.n1819 9.3005
R11965 gnd.n4212 gnd.n4211 9.3005
R11966 gnd.n4210 gnd.n4205 9.3005
R11967 gnd.n2168 gnd.n2167 9.3005
R11968 gnd.n3213 gnd.n3212 9.3005
R11969 gnd.n3214 gnd.n2166 9.3005
R11970 gnd.n3216 gnd.n3215 9.3005
R11971 gnd.n2155 gnd.n2154 9.3005
R11972 gnd.n3229 gnd.n3228 9.3005
R11973 gnd.n3230 gnd.n2153 9.3005
R11974 gnd.n3232 gnd.n3231 9.3005
R11975 gnd.n2140 gnd.n2139 9.3005
R11976 gnd.n3245 gnd.n3244 9.3005
R11977 gnd.n3246 gnd.n2138 9.3005
R11978 gnd.n3248 gnd.n3247 9.3005
R11979 gnd.n2127 gnd.n2126 9.3005
R11980 gnd.n3261 gnd.n3260 9.3005
R11981 gnd.n3262 gnd.n2125 9.3005
R11982 gnd.n3264 gnd.n3263 9.3005
R11983 gnd.n2114 gnd.n2113 9.3005
R11984 gnd.n3277 gnd.n3276 9.3005
R11985 gnd.n3278 gnd.n2112 9.3005
R11986 gnd.n3280 gnd.n3279 9.3005
R11987 gnd.n2100 gnd.n2099 9.3005
R11988 gnd.n3295 gnd.n3294 9.3005
R11989 gnd.n3296 gnd.n2097 9.3005
R11990 gnd.n3299 gnd.n3298 9.3005
R11991 gnd.n3297 gnd.n2098 9.3005
R11992 gnd.n2072 gnd.n2071 9.3005
R11993 gnd.n3909 gnd.n3908 9.3005
R11994 gnd.n3910 gnd.n2070 9.3005
R11995 gnd.n3912 gnd.n3911 9.3005
R11996 gnd.n2057 gnd.n2056 9.3005
R11997 gnd.n3925 gnd.n3924 9.3005
R11998 gnd.n3926 gnd.n2055 9.3005
R11999 gnd.n3928 gnd.n3927 9.3005
R12000 gnd.n2042 gnd.n2041 9.3005
R12001 gnd.n3941 gnd.n3940 9.3005
R12002 gnd.n3942 gnd.n2040 9.3005
R12003 gnd.n3944 gnd.n3943 9.3005
R12004 gnd.n2028 gnd.n2027 9.3005
R12005 gnd.n3957 gnd.n3956 9.3005
R12006 gnd.n3958 gnd.n2026 9.3005
R12007 gnd.n3960 gnd.n3959 9.3005
R12008 gnd.n2013 gnd.n2012 9.3005
R12009 gnd.n3973 gnd.n3972 9.3005
R12010 gnd.n3974 gnd.n2011 9.3005
R12011 gnd.n3976 gnd.n3975 9.3005
R12012 gnd.n1998 gnd.n1997 9.3005
R12013 gnd.n3989 gnd.n3988 9.3005
R12014 gnd.n3990 gnd.n1996 9.3005
R12015 gnd.n3992 gnd.n3991 9.3005
R12016 gnd.n1983 gnd.n1982 9.3005
R12017 gnd.n4005 gnd.n4004 9.3005
R12018 gnd.n4006 gnd.n1981 9.3005
R12019 gnd.n4008 gnd.n4007 9.3005
R12020 gnd.n1968 gnd.n1967 9.3005
R12021 gnd.n4021 gnd.n4020 9.3005
R12022 gnd.n4022 gnd.n1966 9.3005
R12023 gnd.n4024 gnd.n4023 9.3005
R12024 gnd.n1953 gnd.n1952 9.3005
R12025 gnd.n4037 gnd.n4036 9.3005
R12026 gnd.n4038 gnd.n1951 9.3005
R12027 gnd.n4040 gnd.n4039 9.3005
R12028 gnd.n1940 gnd.n1939 9.3005
R12029 gnd.n4053 gnd.n4052 9.3005
R12030 gnd.n4054 gnd.n1938 9.3005
R12031 gnd.n4056 gnd.n4055 9.3005
R12032 gnd.n1928 gnd.n1927 9.3005
R12033 gnd.n4069 gnd.n4068 9.3005
R12034 gnd.n4070 gnd.n1926 9.3005
R12035 gnd.n4072 gnd.n4071 9.3005
R12036 gnd.n1915 gnd.n1914 9.3005
R12037 gnd.n4085 gnd.n4084 9.3005
R12038 gnd.n4086 gnd.n1913 9.3005
R12039 gnd.n4088 gnd.n4087 9.3005
R12040 gnd.n1902 gnd.n1901 9.3005
R12041 gnd.n4101 gnd.n4100 9.3005
R12042 gnd.n4102 gnd.n1900 9.3005
R12043 gnd.n4104 gnd.n4103 9.3005
R12044 gnd.n1888 gnd.n1887 9.3005
R12045 gnd.n4117 gnd.n4116 9.3005
R12046 gnd.n4118 gnd.n1886 9.3005
R12047 gnd.n4120 gnd.n4119 9.3005
R12048 gnd.n1874 gnd.n1873 9.3005
R12049 gnd.n4133 gnd.n4132 9.3005
R12050 gnd.n4134 gnd.n1872 9.3005
R12051 gnd.n4136 gnd.n4135 9.3005
R12052 gnd.n1862 gnd.n1861 9.3005
R12053 gnd.n4149 gnd.n4148 9.3005
R12054 gnd.n4150 gnd.n1860 9.3005
R12055 gnd.n4152 gnd.n4151 9.3005
R12056 gnd.n1849 gnd.n1848 9.3005
R12057 gnd.n4165 gnd.n4164 9.3005
R12058 gnd.n4166 gnd.n1847 9.3005
R12059 gnd.n4168 gnd.n4167 9.3005
R12060 gnd.n1836 gnd.n1835 9.3005
R12061 gnd.n4181 gnd.n4180 9.3005
R12062 gnd.n4182 gnd.n1833 9.3005
R12063 gnd.n4186 gnd.n4185 9.3005
R12064 gnd.n4184 gnd.n1834 9.3005
R12065 gnd.n4183 gnd.n1821 9.3005
R12066 gnd.n4202 gnd.n1820 9.3005
R12067 gnd.n4204 gnd.n4203 9.3005
R12068 gnd.n3200 gnd.n3199 9.3005
R12069 gnd.n3196 gnd.n2178 9.3005
R12070 gnd.n2811 gnd.n2179 9.3005
R12071 gnd.n2814 gnd.n2813 9.3005
R12072 gnd.n2816 gnd.n2815 9.3005
R12073 gnd.n2817 gnd.n2804 9.3005
R12074 gnd.n2819 gnd.n2818 9.3005
R12075 gnd.n2820 gnd.n2803 9.3005
R12076 gnd.n2822 gnd.n2821 9.3005
R12077 gnd.n2823 gnd.n2798 9.3005
R12078 gnd.n3198 gnd.n3197 9.3005
R12079 gnd.n2633 gnd.n2632 9.3005
R12080 gnd.n2631 gnd.n2629 9.3005
R12081 gnd.n2377 gnd.n2376 9.3005
R12082 gnd.n2662 gnd.n2661 9.3005
R12083 gnd.n2663 gnd.n2375 9.3005
R12084 gnd.n2665 gnd.n2664 9.3005
R12085 gnd.n2370 gnd.n2369 9.3005
R12086 gnd.n2679 gnd.n2678 9.3005
R12087 gnd.n2680 gnd.n2368 9.3005
R12088 gnd.n2682 gnd.n2681 9.3005
R12089 gnd.n2357 gnd.n2355 9.3005
R12090 gnd.n2721 gnd.n2720 9.3005
R12091 gnd.n2719 gnd.n2356 9.3005
R12092 gnd.n2718 gnd.n2717 9.3005
R12093 gnd.n2716 gnd.n2358 9.3005
R12094 gnd.n2715 gnd.n2714 9.3005
R12095 gnd.n2713 gnd.n2361 9.3005
R12096 gnd.n2712 gnd.n2711 9.3005
R12097 gnd.n2341 gnd.n2340 9.3005
R12098 gnd.n2779 gnd.n2778 9.3005
R12099 gnd.n2780 gnd.n2339 9.3005
R12100 gnd.n2782 gnd.n2781 9.3005
R12101 gnd.n2335 gnd.n2334 9.3005
R12102 gnd.n2796 gnd.n2795 9.3005
R12103 gnd.n2797 gnd.n2332 9.3005
R12104 gnd.n2829 gnd.n2828 9.3005
R12105 gnd.n2827 gnd.n2333 9.3005
R12106 gnd.n2825 gnd.n2824 9.3005
R12107 gnd.n2247 gnd.n2246 9.3005
R12108 gnd.n3149 gnd.n3148 9.3005
R12109 gnd.n3151 gnd.n3150 9.3005
R12110 gnd.n2235 gnd.n2234 9.3005
R12111 gnd.n3157 gnd.n3156 9.3005
R12112 gnd.n3159 gnd.n3158 9.3005
R12113 gnd.n2227 gnd.n2226 9.3005
R12114 gnd.n3165 gnd.n3164 9.3005
R12115 gnd.n3167 gnd.n3166 9.3005
R12116 gnd.n2217 gnd.n2216 9.3005
R12117 gnd.n3173 gnd.n3172 9.3005
R12118 gnd.n3175 gnd.n3174 9.3005
R12119 gnd.n2209 gnd.n2208 9.3005
R12120 gnd.n3181 gnd.n3180 9.3005
R12121 gnd.n3183 gnd.n3182 9.3005
R12122 gnd.n2199 gnd.n2197 9.3005
R12123 gnd.n3189 gnd.n3188 9.3005
R12124 gnd.n3190 gnd.n2196 9.3005
R12125 gnd.n2250 gnd.n1277 9.3005
R12126 gnd.n2200 gnd.n2198 9.3005
R12127 gnd.n3187 gnd.n3186 9.3005
R12128 gnd.n3185 gnd.n3184 9.3005
R12129 gnd.n2204 gnd.n2203 9.3005
R12130 gnd.n3179 gnd.n3178 9.3005
R12131 gnd.n3177 gnd.n3176 9.3005
R12132 gnd.n2213 gnd.n2212 9.3005
R12133 gnd.n3171 gnd.n3170 9.3005
R12134 gnd.n3169 gnd.n3168 9.3005
R12135 gnd.n2221 gnd.n2220 9.3005
R12136 gnd.n3163 gnd.n3162 9.3005
R12137 gnd.n3161 gnd.n3160 9.3005
R12138 gnd.n2231 gnd.n2230 9.3005
R12139 gnd.n3155 gnd.n3154 9.3005
R12140 gnd.n3153 gnd.n3152 9.3005
R12141 gnd.n2241 gnd.n2240 9.3005
R12142 gnd.n3147 gnd.n3146 9.3005
R12143 gnd.n4659 gnd.n1278 9.3005
R12144 gnd.n4658 gnd.n4657 9.3005
R12145 gnd.n4656 gnd.n1282 9.3005
R12146 gnd.n4655 gnd.n4654 9.3005
R12147 gnd.n4653 gnd.n1283 9.3005
R12148 gnd.n4652 gnd.n4651 9.3005
R12149 gnd.n4650 gnd.n1287 9.3005
R12150 gnd.n4649 gnd.n4648 9.3005
R12151 gnd.n4647 gnd.n1288 9.3005
R12152 gnd.n4646 gnd.n4645 9.3005
R12153 gnd.n4644 gnd.n1292 9.3005
R12154 gnd.n4643 gnd.n4642 9.3005
R12155 gnd.n4641 gnd.n1293 9.3005
R12156 gnd.n4640 gnd.n4639 9.3005
R12157 gnd.n4638 gnd.n1297 9.3005
R12158 gnd.n4637 gnd.n4636 9.3005
R12159 gnd.n4635 gnd.n1298 9.3005
R12160 gnd.n4634 gnd.n4633 9.3005
R12161 gnd.n4632 gnd.n1302 9.3005
R12162 gnd.n4631 gnd.n4630 9.3005
R12163 gnd.n4629 gnd.n1303 9.3005
R12164 gnd.n4628 gnd.n4627 9.3005
R12165 gnd.n4626 gnd.n1307 9.3005
R12166 gnd.n4625 gnd.n4624 9.3005
R12167 gnd.n4623 gnd.n1308 9.3005
R12168 gnd.n4622 gnd.n4621 9.3005
R12169 gnd.n4620 gnd.n1312 9.3005
R12170 gnd.n4619 gnd.n4618 9.3005
R12171 gnd.n4617 gnd.n1313 9.3005
R12172 gnd.n4616 gnd.n4615 9.3005
R12173 gnd.n4614 gnd.n1317 9.3005
R12174 gnd.n4613 gnd.n4612 9.3005
R12175 gnd.n4611 gnd.n1318 9.3005
R12176 gnd.n4610 gnd.n4609 9.3005
R12177 gnd.n4608 gnd.n1322 9.3005
R12178 gnd.n4607 gnd.n4606 9.3005
R12179 gnd.n4605 gnd.n1323 9.3005
R12180 gnd.n4604 gnd.n4603 9.3005
R12181 gnd.n4602 gnd.n1327 9.3005
R12182 gnd.n4601 gnd.n4600 9.3005
R12183 gnd.n4599 gnd.n1328 9.3005
R12184 gnd.n4598 gnd.n4597 9.3005
R12185 gnd.n4596 gnd.n1332 9.3005
R12186 gnd.n4595 gnd.n4594 9.3005
R12187 gnd.n4593 gnd.n1333 9.3005
R12188 gnd.n4592 gnd.n4591 9.3005
R12189 gnd.n4590 gnd.n1337 9.3005
R12190 gnd.n4589 gnd.n4588 9.3005
R12191 gnd.n4587 gnd.n1338 9.3005
R12192 gnd.n4586 gnd.n4585 9.3005
R12193 gnd.n4584 gnd.n1342 9.3005
R12194 gnd.n4583 gnd.n4582 9.3005
R12195 gnd.n4581 gnd.n1343 9.3005
R12196 gnd.n4580 gnd.n4579 9.3005
R12197 gnd.n4578 gnd.n1347 9.3005
R12198 gnd.n4577 gnd.n4576 9.3005
R12199 gnd.n4575 gnd.n1348 9.3005
R12200 gnd.n4574 gnd.n4573 9.3005
R12201 gnd.n4572 gnd.n1352 9.3005
R12202 gnd.n4571 gnd.n4570 9.3005
R12203 gnd.n4569 gnd.n1353 9.3005
R12204 gnd.n4568 gnd.n4567 9.3005
R12205 gnd.n4566 gnd.n1357 9.3005
R12206 gnd.n4565 gnd.n4564 9.3005
R12207 gnd.n4563 gnd.n1358 9.3005
R12208 gnd.n4562 gnd.n4561 9.3005
R12209 gnd.n4560 gnd.n1362 9.3005
R12210 gnd.n4559 gnd.n4558 9.3005
R12211 gnd.n4557 gnd.n1363 9.3005
R12212 gnd.n4556 gnd.n4555 9.3005
R12213 gnd.n4554 gnd.n1367 9.3005
R12214 gnd.n4553 gnd.n4552 9.3005
R12215 gnd.n4551 gnd.n1368 9.3005
R12216 gnd.n4550 gnd.n4549 9.3005
R12217 gnd.n4548 gnd.n1372 9.3005
R12218 gnd.n4547 gnd.n4546 9.3005
R12219 gnd.n4545 gnd.n1373 9.3005
R12220 gnd.n4544 gnd.n4543 9.3005
R12221 gnd.n4542 gnd.n1377 9.3005
R12222 gnd.n4541 gnd.n4540 9.3005
R12223 gnd.n4539 gnd.n1378 9.3005
R12224 gnd.n4538 gnd.n4537 9.3005
R12225 gnd.n4536 gnd.n1382 9.3005
R12226 gnd.n4535 gnd.n4534 9.3005
R12227 gnd.n4533 gnd.n1383 9.3005
R12228 gnd.n4532 gnd.n4531 9.3005
R12229 gnd.n4530 gnd.n1387 9.3005
R12230 gnd.n4529 gnd.n4528 9.3005
R12231 gnd.n4527 gnd.n1388 9.3005
R12232 gnd.n4526 gnd.n4525 9.3005
R12233 gnd.n4524 gnd.n1392 9.3005
R12234 gnd.n4523 gnd.n4522 9.3005
R12235 gnd.n4521 gnd.n1393 9.3005
R12236 gnd.n4520 gnd.n4519 9.3005
R12237 gnd.n4518 gnd.n1397 9.3005
R12238 gnd.n4517 gnd.n4516 9.3005
R12239 gnd.n4515 gnd.n1398 9.3005
R12240 gnd.n4514 gnd.n4513 9.3005
R12241 gnd.n4512 gnd.n1402 9.3005
R12242 gnd.n4511 gnd.n4510 9.3005
R12243 gnd.n4509 gnd.n1403 9.3005
R12244 gnd.n4661 gnd.n4660 9.3005
R12245 gnd.n4418 gnd.n1502 9.3005
R12246 gnd.n4417 gnd.n4416 9.3005
R12247 gnd.n4415 gnd.n1504 9.3005
R12248 gnd.n4414 gnd.n4413 9.3005
R12249 gnd.n4412 gnd.n1508 9.3005
R12250 gnd.n4411 gnd.n4410 9.3005
R12251 gnd.n4409 gnd.n1509 9.3005
R12252 gnd.n4408 gnd.n4407 9.3005
R12253 gnd.n4406 gnd.n1513 9.3005
R12254 gnd.n4405 gnd.n4404 9.3005
R12255 gnd.n4403 gnd.n1514 9.3005
R12256 gnd.n4402 gnd.n4401 9.3005
R12257 gnd.n4400 gnd.n1518 9.3005
R12258 gnd.n4399 gnd.n4398 9.3005
R12259 gnd.n4397 gnd.n1519 9.3005
R12260 gnd.n4396 gnd.n4395 9.3005
R12261 gnd.n4394 gnd.n1523 9.3005
R12262 gnd.n4393 gnd.n4392 9.3005
R12263 gnd.n4391 gnd.n1524 9.3005
R12264 gnd.n4390 gnd.n4389 9.3005
R12265 gnd.n285 gnd.n283 9.3005
R12266 gnd.n7290 gnd.n7289 9.3005
R12267 gnd.n7288 gnd.n284 9.3005
R12268 gnd.n7287 gnd.n7286 9.3005
R12269 gnd.n7285 gnd.n286 9.3005
R12270 gnd.n7284 gnd.n7283 9.3005
R12271 gnd.n7281 gnd.n290 9.3005
R12272 gnd.n7280 gnd.n7279 9.3005
R12273 gnd.n7278 gnd.n292 9.3005
R12274 gnd.n261 gnd.n260 9.3005
R12275 gnd.n7302 gnd.n7301 9.3005
R12276 gnd.n7303 gnd.n259 9.3005
R12277 gnd.n7305 gnd.n7304 9.3005
R12278 gnd.n245 gnd.n244 9.3005
R12279 gnd.n7318 gnd.n7317 9.3005
R12280 gnd.n7319 gnd.n243 9.3005
R12281 gnd.n7321 gnd.n7320 9.3005
R12282 gnd.n230 gnd.n229 9.3005
R12283 gnd.n7334 gnd.n7333 9.3005
R12284 gnd.n7335 gnd.n228 9.3005
R12285 gnd.n7337 gnd.n7336 9.3005
R12286 gnd.n215 gnd.n214 9.3005
R12287 gnd.n7350 gnd.n7349 9.3005
R12288 gnd.n7351 gnd.n213 9.3005
R12289 gnd.n7353 gnd.n7352 9.3005
R12290 gnd.n200 gnd.n199 9.3005
R12291 gnd.n7366 gnd.n7365 9.3005
R12292 gnd.n7367 gnd.n197 9.3005
R12293 gnd.n7444 gnd.n7443 9.3005
R12294 gnd.n7442 gnd.n198 9.3005
R12295 gnd.n7441 gnd.n7440 9.3005
R12296 gnd.n7439 gnd.n7368 9.3005
R12297 gnd.n7438 gnd.n7437 9.3005
R12298 gnd.n4420 gnd.n4419 9.3005
R12299 gnd.n7434 gnd.n7370 9.3005
R12300 gnd.n7433 gnd.n7432 9.3005
R12301 gnd.n7431 gnd.n7375 9.3005
R12302 gnd.n7430 gnd.n7429 9.3005
R12303 gnd.n7428 gnd.n7376 9.3005
R12304 gnd.n7427 gnd.n7426 9.3005
R12305 gnd.n7425 gnd.n7383 9.3005
R12306 gnd.n7424 gnd.n7423 9.3005
R12307 gnd.n7422 gnd.n7384 9.3005
R12308 gnd.n7421 gnd.n7420 9.3005
R12309 gnd.n7419 gnd.n7391 9.3005
R12310 gnd.n7418 gnd.n7417 9.3005
R12311 gnd.n7416 gnd.n7392 9.3005
R12312 gnd.n7415 gnd.n7414 9.3005
R12313 gnd.n7413 gnd.n7399 9.3005
R12314 gnd.n7412 gnd.n7411 9.3005
R12315 gnd.n7410 gnd.n7400 9.3005
R12316 gnd.n7409 gnd.n7408 9.3005
R12317 gnd.n7436 gnd.n7435 9.3005
R12318 gnd.n4231 gnd.n1681 9.3005
R12319 gnd.n4234 gnd.n4233 9.3005
R12320 gnd.n4232 gnd.n1682 9.3005
R12321 gnd.n1613 gnd.n1612 9.3005
R12322 gnd.n4261 gnd.n4260 9.3005
R12323 gnd.n4262 gnd.n1610 9.3005
R12324 gnd.n4265 gnd.n4264 9.3005
R12325 gnd.n4263 gnd.n1611 9.3005
R12326 gnd.n1586 gnd.n1585 9.3005
R12327 gnd.n4292 gnd.n4291 9.3005
R12328 gnd.n4293 gnd.n1583 9.3005
R12329 gnd.n4301 gnd.n4300 9.3005
R12330 gnd.n4299 gnd.n1584 9.3005
R12331 gnd.n4298 gnd.n4297 9.3005
R12332 gnd.n4296 gnd.n4294 9.3005
R12333 gnd.n1551 gnd.n1549 9.3005
R12334 gnd.n4358 gnd.n4357 9.3005
R12335 gnd.n4356 gnd.n1550 9.3005
R12336 gnd.n4355 gnd.n4354 9.3005
R12337 gnd.n4353 gnd.n1552 9.3005
R12338 gnd.n4352 gnd.n4351 9.3005
R12339 gnd.n311 gnd.n310 9.3005
R12340 gnd.n7195 gnd.n7194 9.3005
R12341 gnd.n7196 gnd.n309 9.3005
R12342 gnd.n7198 gnd.n7197 9.3005
R12343 gnd.n69 gnd.n67 9.3005
R12344 gnd.n7575 gnd.n7574 9.3005
R12345 gnd.n7573 gnd.n68 9.3005
R12346 gnd.n7572 gnd.n7571 9.3005
R12347 gnd.n7570 gnd.n73 9.3005
R12348 gnd.n7569 gnd.n7568 9.3005
R12349 gnd.n7567 gnd.n74 9.3005
R12350 gnd.n7566 gnd.n7565 9.3005
R12351 gnd.n7564 gnd.n78 9.3005
R12352 gnd.n7563 gnd.n7562 9.3005
R12353 gnd.n7561 gnd.n79 9.3005
R12354 gnd.n7560 gnd.n7559 9.3005
R12355 gnd.n7558 gnd.n83 9.3005
R12356 gnd.n7557 gnd.n7556 9.3005
R12357 gnd.n7555 gnd.n84 9.3005
R12358 gnd.n7554 gnd.n7553 9.3005
R12359 gnd.n7552 gnd.n88 9.3005
R12360 gnd.n7551 gnd.n7550 9.3005
R12361 gnd.n7549 gnd.n89 9.3005
R12362 gnd.n7548 gnd.n7547 9.3005
R12363 gnd.n7546 gnd.n93 9.3005
R12364 gnd.n7545 gnd.n7544 9.3005
R12365 gnd.n7543 gnd.n94 9.3005
R12366 gnd.n7542 gnd.n7541 9.3005
R12367 gnd.n7540 gnd.n98 9.3005
R12368 gnd.n7539 gnd.n7538 9.3005
R12369 gnd.n7537 gnd.n99 9.3005
R12370 gnd.n7536 gnd.n102 9.3005
R12371 gnd.n4230 gnd.n4229 9.3005
R12372 gnd.n5803 gnd.t35 9.24152
R12373 gnd.n6317 gnd.t68 9.24152
R12374 gnd.t80 gnd.n922 9.24152
R12375 gnd.t64 gnd.n1015 9.24152
R12376 gnd.n2696 gnd.t199 9.24152
R12377 gnd.n4673 gnd.t76 9.24152
R12378 gnd.t95 gnd.n4236 9.24152
R12379 gnd.n4304 gnd.t207 9.24152
R12380 gnd.t320 gnd.t35 8.92286
R12381 gnd.n3035 gnd.t135 8.92286
R12382 gnd.n3292 gnd.n2103 8.92286
R12383 gnd.n3302 gnd.t129 8.92286
R12384 gnd.t6 gnd.n3307 8.92286
R12385 gnd.n3954 gnd.n2031 8.92286
R12386 gnd.n3978 gnd.n2008 8.92286
R12387 gnd.n3789 gnd.n3403 8.92286
R12388 gnd.n3768 gnd.n3767 8.92286
R12389 gnd.n4098 gnd.t190 8.92286
R12390 gnd.n4114 gnd.n1890 8.92286
R12391 gnd.t122 gnd.n1876 8.92286
R12392 gnd.n6153 gnd.n6128 8.92171
R12393 gnd.n6121 gnd.n6096 8.92171
R12394 gnd.n6089 gnd.n6064 8.92171
R12395 gnd.n6058 gnd.n6033 8.92171
R12396 gnd.n6026 gnd.n6001 8.92171
R12397 gnd.n5994 gnd.n5969 8.92171
R12398 gnd.n5962 gnd.n5937 8.92171
R12399 gnd.n5931 gnd.n5906 8.92171
R12400 gnd.n3514 gnd.n3496 8.72777
R12401 gnd.t10 gnd.n5109 8.60421
R12402 gnd.n2371 gnd.t228 8.60421
R12403 gnd.n1540 gnd.t203 8.60421
R12404 gnd.n5517 gnd.n5501 8.43467
R12405 gnd.n50 gnd.n34 8.43467
R12406 gnd.n2630 gnd.n0 8.41456
R12407 gnd.n7577 gnd.n7576 8.41456
R12408 gnd.n6154 gnd.n6126 8.14595
R12409 gnd.n6122 gnd.n6094 8.14595
R12410 gnd.n6090 gnd.n6062 8.14595
R12411 gnd.n6059 gnd.n6031 8.14595
R12412 gnd.n6027 gnd.n5999 8.14595
R12413 gnd.n5995 gnd.n5967 8.14595
R12414 gnd.n5963 gnd.n5935 8.14595
R12415 gnd.n5932 gnd.n5904 8.14595
R12416 gnd.n6159 gnd.n6158 7.97301
R12417 gnd.t55 gnd.n5151 7.9669
R12418 gnd.n2614 gnd.t201 7.9669
R12419 gnd.n3193 gnd.n2181 7.9669
R12420 gnd.n1417 gnd.n1409 7.9669
R12421 gnd.n321 gnd.t289 7.9669
R12422 gnd.n7410 gnd.n7409 7.75808
R12423 gnd.n1800 gnd.n1799 7.75808
R12424 gnd.n3146 gnd.n2240 7.75808
R12425 gnd.n2497 gnd.n2494 7.75808
R12426 gnd.n3282 gnd.n2110 7.64824
R12427 gnd.n3946 gnd.n2038 7.64824
R12428 gnd.n3824 gnd.t294 7.64824
R12429 gnd.n3986 gnd.n2000 7.64824
R12430 gnd.n3796 gnd.n3396 7.64824
R12431 gnd.t219 gnd.n1970 7.64824
R12432 gnd.n3760 gnd.n3428 7.64824
R12433 gnd.n186 gnd.t84 7.64824
R12434 gnd.n5633 gnd.t12 7.32958
R12435 gnd.n3210 gnd.t115 7.32958
R12436 gnd.n2144 gnd.t4 7.32958
R12437 gnd.t248 gnd.n2110 7.32958
R12438 gnd.n3696 gnd.t325 7.32958
R12439 gnd.t235 gnd.n1851 7.32958
R12440 gnd.n4199 gnd.t72 7.32958
R12441 gnd.n2926 gnd.n2925 7.30353
R12442 gnd.n3513 gnd.n3512 7.30353
R12443 gnd.n5593 gnd.n5226 7.01093
R12444 gnd.n5229 gnd.n5227 7.01093
R12445 gnd.n5603 gnd.n5602 7.01093
R12446 gnd.n5614 gnd.n5210 7.01093
R12447 gnd.n5613 gnd.n5213 7.01093
R12448 gnd.n5624 gnd.n5201 7.01093
R12449 gnd.n5204 gnd.n5202 7.01093
R12450 gnd.n5634 gnd.n5633 7.01093
R12451 gnd.n5645 gnd.n5184 7.01093
R12452 gnd.n5644 gnd.n5187 7.01093
R12453 gnd.n5655 gnd.n5177 7.01093
R12454 gnd.n5547 gnd.n5170 7.01093
R12455 gnd.n5676 gnd.n5159 7.01093
R12456 gnd.n5675 gnd.n5162 7.01093
R12457 gnd.n5686 gnd.n5151 7.01093
R12458 gnd.n5152 gnd.n5144 7.01093
R12459 gnd.n5707 gnd.n5133 7.01093
R12460 gnd.n5706 gnd.n5136 7.01093
R12461 gnd.n5126 gnd.n5119 7.01093
R12462 gnd.n5727 gnd.n5726 7.01093
R12463 gnd.n5737 gnd.n5109 7.01093
R12464 gnd.n5736 gnd.n5112 7.01093
R12465 gnd.n5747 gnd.n5102 7.01093
R12466 gnd.n5757 gnd.n5095 7.01093
R12467 gnd.n5781 gnd.n5089 7.01093
R12468 gnd.n5790 gnd.n5080 7.01093
R12469 gnd.n5799 gnd.n5072 7.01093
R12470 gnd.n5803 gnd.n5802 7.01093
R12471 gnd.n5821 gnd.n5057 7.01093
R12472 gnd.n5820 gnd.n5060 7.01093
R12473 gnd.n5831 gnd.n5049 7.01093
R12474 gnd.n5050 gnd.n5039 7.01093
R12475 gnd.n5866 gnd.n5865 7.01093
R12476 gnd.n5878 gnd.n5877 7.01093
R12477 gnd.n5026 gnd.n5018 7.01093
R12478 gnd.n5889 gnd.n5888 7.01093
R12479 gnd.n6188 gnd.n5003 7.01093
R12480 gnd.n6187 gnd.n5006 7.01093
R12481 gnd.n6203 gnd.n896 7.01093
R12482 gnd.n6330 gnd.n898 7.01093
R12483 gnd.n6209 gnd.n907 7.01093
R12484 gnd.n6324 gnd.n6323 7.01093
R12485 gnd.n6172 gnd.n910 7.01093
R12486 gnd.n6317 gnd.n919 7.01093
R12487 gnd.n6316 gnd.n922 7.01093
R12488 gnd.n6220 gnd.n930 7.01093
R12489 gnd.n6310 gnd.n6309 7.01093
R12490 gnd.t173 gnd.n2090 7.01093
R12491 gnd.n3831 gnd.t292 7.01093
R12492 gnd.t266 gnd.n1964 7.01093
R12493 gnd.n4090 gnd.t254 7.01093
R12494 gnd.n5187 gnd.t14 6.69227
R12495 gnd.n5799 gnd.t320 6.69227
R12496 gnd.n6202 gnd.t211 6.69227
R12497 gnd.n6331 gnd.n896 6.69227
R12498 gnd.n4800 gnd.t257 6.69227
R12499 gnd.n2709 gnd.t272 6.69227
R12500 gnd.t263 gnd.n2017 6.69227
R12501 gnd.n3783 gnd.t246 6.69227
R12502 gnd.n1601 gnd.t23 6.69227
R12503 gnd.t27 gnd.n208 6.69227
R12504 gnd.n3619 gnd.n3618 6.5566
R12505 gnd.n3106 gnd.n3105 6.5566
R12506 gnd.n2950 gnd.n2944 6.5566
R12507 gnd.n3634 gnd.n3633 6.5566
R12508 gnd.n3274 gnd.n2116 6.37362
R12509 gnd.t135 gnd.t125 6.37362
R12510 gnd.n3938 gnd.n2046 6.37362
R12511 gnd.n3838 gnd.t198 6.37362
R12512 gnd.n3994 gnd.n1993 6.37362
R12513 gnd.n3803 gnd.n3389 6.37362
R12514 gnd.n4034 gnd.t51 6.37362
R12515 gnd.n3753 gnd.n3752 6.37362
R12516 gnd.n4114 gnd.t61 6.37362
R12517 gnd.n3702 gnd.t61 6.37362
R12518 gnd.n4130 gnd.n1876 6.37362
R12519 gnd.n2813 gnd.n2810 6.20656
R12520 gnd.n7499 gnd.n7496 6.20656
R12521 gnd.n4869 gnd.n4868 6.20656
R12522 gnd.n4218 gnd.n4215 6.20656
R12523 gnd.t217 gnd.n5695 6.05496
R12524 gnd.n5696 gnd.t52 6.05496
R12525 gnd.t268 gnd.n5736 6.05496
R12526 gnd.n5835 gnd.t53 6.05496
R12527 gnd.n4776 gnd.t56 6.05496
R12528 gnd.n2684 gnd.t21 6.05496
R12529 gnd.t303 gnd.n2044 6.05496
R12530 gnd.t215 gnd.t37 6.05496
R12531 gnd.t291 gnd.t170 6.05496
R12532 gnd.n3751 gnd.t187 6.05496
R12533 gnd.n4361 gnd.t183 6.05496
R12534 gnd.t58 gnd.n238 6.05496
R12535 gnd.n6156 gnd.n6126 5.81868
R12536 gnd.n6124 gnd.n6094 5.81868
R12537 gnd.n6092 gnd.n6062 5.81868
R12538 gnd.n6061 gnd.n6031 5.81868
R12539 gnd.n6029 gnd.n5999 5.81868
R12540 gnd.n5997 gnd.n5967 5.81868
R12541 gnd.n5965 gnd.n5935 5.81868
R12542 gnd.n5934 gnd.n5904 5.81868
R12543 gnd.t88 gnd.n1898 5.73631
R12544 gnd.n3541 gnd.n1466 5.62001
R12545 gnd.n3113 gnd.n2880 5.62001
R12546 gnd.n3113 gnd.n2881 5.62001
R12547 gnd.n3628 gnd.n1466 5.62001
R12548 gnd.n5366 gnd.n5361 5.4308
R12549 gnd.n4984 gnd.n4982 5.4308
R12550 gnd.n5747 gnd.t54 5.41765
R12551 gnd.n5791 gnd.t11 5.41765
R12552 gnd.n5867 gnd.t2 5.41765
R12553 gnd.n1098 gnd.n1097 5.41765
R12554 gnd.n4752 gnd.t201 5.41765
R12555 gnd.n2627 gnd.t33 5.41765
R12556 gnd.n7200 gnd.t233 5.41765
R12557 gnd.n7271 gnd.t289 5.41765
R12558 gnd.n7315 gnd.n250 5.41765
R12559 gnd.t48 gnd.n3882 5.09899
R12560 gnd.n3930 gnd.n2053 5.09899
R12561 gnd.n3810 gnd.n3382 5.09899
R12562 gnd.n4002 gnd.n1985 5.09899
R12563 gnd.n3745 gnd.n3443 5.09899
R12564 gnd.n4082 gnd.t222 5.09899
R12565 gnd.n6154 gnd.n6153 5.04292
R12566 gnd.n6122 gnd.n6121 5.04292
R12567 gnd.n6090 gnd.n6089 5.04292
R12568 gnd.n6059 gnd.n6058 5.04292
R12569 gnd.n6027 gnd.n6026 5.04292
R12570 gnd.n5995 gnd.n5994 5.04292
R12571 gnd.n5963 gnd.n5962 5.04292
R12572 gnd.n5932 gnd.n5931 5.04292
R12573 gnd.n5533 gnd.n5532 4.82753
R12574 gnd.n66 gnd.n65 4.82753
R12575 gnd.n5717 gnd.t45 4.78034
R12576 gnd.n5060 gnd.t44 4.78034
R12577 gnd.n2592 gnd.t31 4.78034
R12578 gnd.n4727 gnd.t228 4.78034
R12579 gnd.n3266 gnd.t301 4.78034
R12580 gnd.n3516 gnd.t112 4.78034
R12581 gnd.n4138 gnd.t213 4.78034
R12582 gnd.n4387 gnd.t203 4.78034
R12583 gnd.n7307 gnd.t185 4.78034
R12584 gnd.n5537 gnd.n5536 4.74817
R12585 gnd.n5486 gnd.n5484 4.74817
R12586 gnd.n5479 gnd.n5478 4.74817
R12587 gnd.n5475 gnd.n5474 4.74817
R12588 gnd.n5536 gnd.n5473 4.74817
R12589 gnd.n5486 gnd.n5485 4.74817
R12590 gnd.n5480 gnd.n5479 4.74817
R12591 gnd.n5477 gnd.n5475 4.74817
R12592 gnd.n7295 gnd.n7294 4.74817
R12593 gnd.n7203 gnd.n272 4.74817
R12594 gnd.n7273 gnd.n271 4.74817
R12595 gnd.n270 gnd.n267 4.74817
R12596 gnd.n7295 gnd.n274 4.74817
R12597 gnd.n306 gnd.n272 4.74817
R12598 gnd.n7202 gnd.n271 4.74817
R12599 gnd.n7274 gnd.n270 4.74817
R12600 gnd.n2407 gnd.n2404 4.74817
R12601 gnd.n2612 gnd.n2403 4.74817
R12602 gnd.n2608 gnd.n2402 4.74817
R12603 gnd.n2401 gnd.n2381 4.74817
R12604 gnd.n2655 gnd.n2382 4.74817
R12605 gnd.n4370 gnd.n317 4.74817
R12606 gnd.n7188 gnd.n7187 4.74817
R12607 gnd.n7183 gnd.n318 4.74817
R12608 gnd.n7181 gnd.n7180 4.74817
R12609 gnd.n7176 gnd.n325 4.74817
R12610 gnd.n4371 gnd.n4370 4.74817
R12611 gnd.n7189 gnd.n7188 4.74817
R12612 gnd.n7186 gnd.n318 4.74817
R12613 gnd.n7182 gnd.n7181 4.74817
R12614 gnd.n325 gnd.n323 4.74817
R12615 gnd.n1124 gnd.n1107 4.74817
R12616 gnd.n1143 gnd.n1126 4.74817
R12617 gnd.n4743 gnd.n4742 4.74817
R12618 gnd.n1161 gnd.n1144 4.74817
R12619 gnd.n4756 gnd.n1124 4.74817
R12620 gnd.n4754 gnd.n1126 4.74817
R12621 gnd.n4744 gnd.n4743 4.74817
R12622 gnd.n4741 gnd.n1144 4.74817
R12623 gnd.n2603 gnd.n2404 4.74817
R12624 gnd.n2604 gnd.n2403 4.74817
R12625 gnd.n2611 gnd.n2402 4.74817
R12626 gnd.n2607 gnd.n2401 4.74817
R12627 gnd.n2656 gnd.n2655 4.74817
R12628 gnd.n5517 gnd.n5516 4.7074
R12629 gnd.n50 gnd.n49 4.7074
R12630 gnd.n5533 gnd.n5517 4.65959
R12631 gnd.n66 gnd.n50 4.65959
R12632 gnd.n4466 gnd.n1468 4.6132
R12633 gnd.n3114 gnd.n2879 4.6132
R12634 gnd.n3349 gnd.t172 4.46168
R12635 gnd.n4042 gnd.t196 4.46168
R12636 gnd.n4122 gnd.t163 4.46168
R12637 gnd.n3509 gnd.n3496 4.46111
R12638 gnd.n6139 gnd.n6135 4.38594
R12639 gnd.n6107 gnd.n6103 4.38594
R12640 gnd.n6075 gnd.n6071 4.38594
R12641 gnd.n6044 gnd.n6040 4.38594
R12642 gnd.n6012 gnd.n6008 4.38594
R12643 gnd.n5980 gnd.n5976 4.38594
R12644 gnd.n5948 gnd.n5944 4.38594
R12645 gnd.n5917 gnd.n5913 4.38594
R12646 gnd.n6150 gnd.n6128 4.26717
R12647 gnd.n6118 gnd.n6096 4.26717
R12648 gnd.n6086 gnd.n6064 4.26717
R12649 gnd.n6055 gnd.n6033 4.26717
R12650 gnd.n6023 gnd.n6001 4.26717
R12651 gnd.n5991 gnd.n5969 4.26717
R12652 gnd.n5959 gnd.n5937 4.26717
R12653 gnd.n5928 gnd.n5906 4.26717
R12654 gnd.n5665 gnd.t212 4.14303
R12655 gnd.n5888 gnd.t9 4.14303
R12656 gnd.n1067 gnd.t177 4.14303
R12657 gnd.n4703 gnd.t199 4.14303
R12658 gnd.n2331 gnd.t76 4.14303
R12659 gnd.n4237 gnd.t95 4.14303
R12660 gnd.t207 gnd.n4303 4.14303
R12661 gnd.n7339 gnd.t179 4.14303
R12662 gnd.n6158 gnd.n6157 4.08274
R12663 gnd.n3618 gnd.n3617 4.05904
R12664 gnd.n3105 gnd.n3104 4.05904
R12665 gnd.n2954 gnd.n2944 4.05904
R12666 gnd.n3635 gnd.n3634 4.05904
R12667 gnd.n19 gnd.n9 3.99943
R12668 gnd.n3043 gnd.n2904 3.82437
R12669 gnd.t125 gnd.n2102 3.82437
R12670 gnd.n3922 gnd.n2061 3.82437
R12671 gnd.n3868 gnd.t189 3.82437
R12672 gnd.n3860 gnd.n3334 3.82437
R12673 gnd.n3817 gnd.n3375 3.82437
R12674 gnd.n4010 gnd.n1978 3.82437
R12675 gnd.n4058 gnd.n1936 3.82437
R12676 gnd.n3442 gnd.t293 3.82437
R12677 gnd.n3738 gnd.n3737 3.82437
R12678 gnd.n3702 gnd.t91 3.82437
R12679 gnd.n3690 gnd.n3494 3.82437
R12680 gnd.n6158 gnd.n6030 3.70378
R12681 gnd.n5535 gnd.n5534 3.65935
R12682 gnd.n19 gnd.n18 3.60163
R12683 gnd.n6149 gnd.n6130 3.49141
R12684 gnd.n6117 gnd.n6098 3.49141
R12685 gnd.n6085 gnd.n6066 3.49141
R12686 gnd.n6054 gnd.n6035 3.49141
R12687 gnd.n6022 gnd.n6003 3.49141
R12688 gnd.n5990 gnd.n5971 3.49141
R12689 gnd.n5958 gnd.n5939 3.49141
R12690 gnd.n5927 gnd.n5908 3.49141
R12691 gnd.n3875 gnd.t265 3.18706
R12692 gnd.t265 gnd.n3321 3.18706
R12693 gnd.n4074 gnd.t295 3.18706
R12694 gnd.n3739 gnd.t295 3.18706
R12695 gnd.n3696 gnd.t163 3.18706
R12696 gnd.t212 gnd.n5664 2.8684
R12697 gnd.n2649 gnd.t174 2.8684
R12698 gnd.n3898 gnd.t49 2.8684
R12699 gnd.n3470 gnd.t239 2.8684
R12700 gnd.t205 gnd.n263 2.8684
R12701 gnd.n5518 gnd.t230 2.82907
R12702 gnd.n5518 gnd.t324 2.82907
R12703 gnd.n5520 gnd.t245 2.82907
R12704 gnd.n5520 gnd.t232 2.82907
R12705 gnd.n5522 gnd.t309 2.82907
R12706 gnd.n5522 gnd.t287 2.82907
R12707 gnd.n5524 gnd.t331 2.82907
R12708 gnd.n5524 gnd.t308 2.82907
R12709 gnd.n5526 gnd.t251 2.82907
R12710 gnd.n5526 gnd.t242 2.82907
R12711 gnd.n5528 gnd.t244 2.82907
R12712 gnd.n5528 gnd.t310 2.82907
R12713 gnd.n5530 gnd.t307 2.82907
R12714 gnd.n5530 gnd.t227 2.82907
R12715 gnd.n5487 gnd.t200 2.82907
R12716 gnd.n5487 gnd.t275 2.82907
R12717 gnd.n5489 gnd.t314 2.82907
R12718 gnd.n5489 gnd.t182 2.82907
R12719 gnd.n5491 gnd.t47 2.82907
R12720 gnd.n5491 gnd.t229 2.82907
R12721 gnd.n5493 gnd.t250 2.82907
R12722 gnd.n5493 gnd.t210 2.82907
R12723 gnd.n5495 gnd.t32 2.82907
R12724 gnd.n5495 gnd.t175 2.82907
R12725 gnd.n5497 gnd.t298 2.82907
R12726 gnd.n5497 gnd.t57 2.82907
R12727 gnd.n5499 gnd.t322 2.82907
R12728 gnd.n5499 gnd.t178 2.82907
R12729 gnd.n5502 gnd.t279 2.82907
R12730 gnd.n5502 gnd.t273 2.82907
R12731 gnd.n5504 gnd.t22 2.82907
R12732 gnd.n5504 gnd.t282 2.82907
R12733 gnd.n5506 gnd.t194 2.82907
R12734 gnd.n5506 gnd.t286 2.82907
R12735 gnd.n5508 gnd.t202 2.82907
R12736 gnd.n5508 gnd.t34 2.82907
R12737 gnd.n5510 gnd.t41 2.82907
R12738 gnd.n5510 gnd.t221 2.82907
R12739 gnd.n5512 gnd.t274 2.82907
R12740 gnd.n5512 gnd.t176 2.82907
R12741 gnd.n5514 gnd.t258 2.82907
R12742 gnd.n5514 gnd.t271 2.82907
R12743 gnd.n63 gnd.t241 2.82907
R12744 gnd.n63 gnd.t317 2.82907
R12745 gnd.n61 gnd.t223 2.82907
R12746 gnd.n61 gnd.t328 2.82907
R12747 gnd.n59 gnd.t311 2.82907
R12748 gnd.n59 gnd.t323 2.82907
R12749 gnd.n57 gnd.t330 2.82907
R12750 gnd.n57 gnd.t290 2.82907
R12751 gnd.n55 gnd.t280 2.82907
R12752 gnd.n55 gnd.t226 2.82907
R12753 gnd.n53 gnd.t224 2.82907
R12754 gnd.n53 gnd.t329 2.82907
R12755 gnd.n51 gnd.t319 2.82907
R12756 gnd.n51 gnd.t327 2.82907
R12757 gnd.n32 gnd.t191 2.82907
R12758 gnd.n32 gnd.t237 2.82907
R12759 gnd.n30 gnd.t209 2.82907
R12760 gnd.n30 gnd.t30 2.82907
R12761 gnd.n28 gnd.t206 2.82907
R12762 gnd.n28 gnd.t270 2.82907
R12763 gnd.n26 gnd.t285 2.82907
R12764 gnd.n26 gnd.t315 2.82907
R12765 gnd.n24 gnd.t260 2.82907
R12766 gnd.n24 gnd.t278 2.82907
R12767 gnd.n22 gnd.t220 2.82907
R12768 gnd.n22 gnd.t184 2.82907
R12769 gnd.n20 gnd.t24 2.82907
R12770 gnd.n20 gnd.t208 2.82907
R12771 gnd.n47 gnd.t180 2.82907
R12772 gnd.n47 gnd.t28 2.82907
R12773 gnd.n45 gnd.t59 2.82907
R12774 gnd.n45 gnd.t256 2.82907
R12775 gnd.n43 gnd.t296 2.82907
R12776 gnd.n43 gnd.t186 2.82907
R12777 gnd.n41 gnd.t234 2.82907
R12778 gnd.n41 gnd.t318 2.82907
R12779 gnd.n39 gnd.t204 2.82907
R12780 gnd.n39 gnd.t277 2.82907
R12781 gnd.n37 gnd.t193 2.82907
R12782 gnd.n37 gnd.t261 2.82907
R12783 gnd.n35 gnd.t255 2.82907
R12784 gnd.n35 gnd.t231 2.82907
R12785 gnd.n6146 gnd.n6145 2.71565
R12786 gnd.n6114 gnd.n6113 2.71565
R12787 gnd.n6082 gnd.n6081 2.71565
R12788 gnd.n6051 gnd.n6050 2.71565
R12789 gnd.n6019 gnd.n6018 2.71565
R12790 gnd.n5987 gnd.n5986 2.71565
R12791 gnd.n5955 gnd.n5954 2.71565
R12792 gnd.n5924 gnd.n5923 2.71565
R12793 gnd.n3036 gnd.n3035 2.54975
R12794 gnd.n3914 gnd.n2068 2.54975
R12795 gnd.n3883 gnd.t48 2.54975
R12796 gnd.n3853 gnd.n3852 2.54975
R12797 gnd.n3852 gnd.t267 2.54975
R12798 gnd.n3824 gnd.n3368 2.54975
R12799 gnd.n4018 gnd.n1970 2.54975
R12800 gnd.n4050 gnd.t262 2.54975
R12801 gnd.n4050 gnd.n1943 2.54975
R12802 gnd.n3731 gnd.t222 2.54975
R12803 gnd.n3457 gnd.n3456 2.54975
R12804 gnd.n3490 gnd.n3489 2.54975
R12805 gnd.n5536 gnd.n5535 2.27742
R12806 gnd.n5535 gnd.n5486 2.27742
R12807 gnd.n5535 gnd.n5479 2.27742
R12808 gnd.n5535 gnd.n5475 2.27742
R12809 gnd.n7296 gnd.n7295 2.27742
R12810 gnd.n7296 gnd.n272 2.27742
R12811 gnd.n7296 gnd.n271 2.27742
R12812 gnd.n7296 gnd.n270 2.27742
R12813 gnd.n4370 gnd.n269 2.27742
R12814 gnd.n7188 gnd.n269 2.27742
R12815 gnd.n318 gnd.n269 2.27742
R12816 gnd.n7181 gnd.n269 2.27742
R12817 gnd.n325 gnd.n269 2.27742
R12818 gnd.n1125 gnd.n1124 2.27742
R12819 gnd.n1126 gnd.n1125 2.27742
R12820 gnd.n4743 gnd.n1125 2.27742
R12821 gnd.n1144 gnd.n1125 2.27742
R12822 gnd.n2654 gnd.n2404 2.27742
R12823 gnd.n2654 gnd.n2403 2.27742
R12824 gnd.n2654 gnd.n2402 2.27742
R12825 gnd.n2654 gnd.n2401 2.27742
R12826 gnd.n2655 gnd.n2654 2.27742
R12827 gnd.n5602 gnd.t147 2.23109
R12828 gnd.n5482 gnd.t45 2.23109
R12829 gnd.n2658 gnd.t46 2.23109
R12830 gnd.n3817 gnd.t215 2.23109
R12831 gnd.t170 gnd.n1978 2.23109
R12832 gnd.n312 gnd.t225 2.23109
R12833 gnd.n6142 gnd.n6132 1.93989
R12834 gnd.n6110 gnd.n6100 1.93989
R12835 gnd.n6078 gnd.n6068 1.93989
R12836 gnd.n6047 gnd.n6037 1.93989
R12837 gnd.n6015 gnd.n6005 1.93989
R12838 gnd.n5983 gnd.n5973 1.93989
R12839 gnd.n5951 gnd.n5941 1.93989
R12840 gnd.n5920 gnd.n5910 1.93989
R12841 gnd.n2906 gnd.t99 1.91244
R12842 gnd.n3890 gnd.t173 1.91244
R12843 gnd.n3724 gnd.t254 1.91244
R12844 gnd.t312 gnd.n5613 1.59378
R12845 gnd.n5780 gnd.t11 1.59378
R12846 gnd.n5834 gnd.t2 1.59378
R12847 gnd.n2724 gnd.t181 1.59378
R12848 gnd.n3883 gnd.t25 1.59378
R12849 gnd.n3954 gnd.t305 1.59378
R12850 gnd.n3767 gnd.t299 1.59378
R12851 gnd.n3731 gnd.t252 1.59378
R12852 gnd.t192 gnd.n1561 1.59378
R12853 gnd.n7454 gnd.n186 1.59378
R12854 gnd.n3274 gnd.t144 1.27512
R12855 gnd.n3028 gnd.n3022 1.27512
R12856 gnd.n3308 gnd.t6 1.27512
R12857 gnd.n3906 gnd.n2076 1.27512
R12858 gnd.t189 gnd.n3867 1.27512
R12859 gnd.n3845 gnd.n3349 1.27512
R12860 gnd.n3831 gnd.n3361 1.27512
R12861 gnd.n4026 gnd.n1964 1.27512
R12862 gnd.n4042 gnd.n1949 1.27512
R12863 gnd.n4066 gnd.t293 1.27512
R12864 gnd.n3723 gnd.n3722 1.27512
R12865 gnd.n3716 gnd.t190 1.27512
R12866 gnd.n3708 gnd.n3477 1.27512
R12867 gnd.n5369 gnd.n5361 1.16414
R12868 gnd.n6235 gnd.n4982 1.16414
R12869 gnd.n6141 gnd.n6134 1.16414
R12870 gnd.n6109 gnd.n6102 1.16414
R12871 gnd.n6077 gnd.n6070 1.16414
R12872 gnd.n6046 gnd.n6039 1.16414
R12873 gnd.n6014 gnd.n6007 1.16414
R12874 gnd.n5982 gnd.n5975 1.16414
R12875 gnd.n5950 gnd.n5943 1.16414
R12876 gnd.n5919 gnd.n5912 1.16414
R12877 gnd.n4466 gnd.n4465 0.970197
R12878 gnd.n3114 gnd.n2304 0.970197
R12879 gnd.n6125 gnd.n6093 0.962709
R12880 gnd.n6157 gnd.n6125 0.962709
R12881 gnd.n5998 gnd.n5966 0.962709
R12882 gnd.n6030 gnd.n5998 0.962709
R12883 gnd.n5696 gnd.t217 0.956468
R12884 gnd.n5844 gnd.t53 0.956468
R12885 gnd.n2775 gnd.t39 0.956468
R12886 gnd.n2123 gnd.n2122 0.956468
R12887 gnd.n3516 gnd.n1878 0.956468
R12888 gnd.n4268 gnd.t42 0.956468
R12889 gnd.n5527 gnd.n5525 0.773756
R12890 gnd.n60 gnd.n58 0.773756
R12891 gnd.n5532 gnd.n5531 0.773756
R12892 gnd.n5531 gnd.n5529 0.773756
R12893 gnd.n5529 gnd.n5527 0.773756
R12894 gnd.n5525 gnd.n5523 0.773756
R12895 gnd.n5523 gnd.n5521 0.773756
R12896 gnd.n5521 gnd.n5519 0.773756
R12897 gnd.n54 gnd.n52 0.773756
R12898 gnd.n56 gnd.n54 0.773756
R12899 gnd.n58 gnd.n56 0.773756
R12900 gnd.n62 gnd.n60 0.773756
R12901 gnd.n64 gnd.n62 0.773756
R12902 gnd.n65 gnd.n64 0.773756
R12903 gnd.n2 gnd.n1 0.672012
R12904 gnd.n3 gnd.n2 0.672012
R12905 gnd.n4 gnd.n3 0.672012
R12906 gnd.n5 gnd.n4 0.672012
R12907 gnd.n6 gnd.n5 0.672012
R12908 gnd.n7 gnd.n6 0.672012
R12909 gnd.n8 gnd.n7 0.672012
R12910 gnd.n9 gnd.n8 0.672012
R12911 gnd.n11 gnd.n10 0.672012
R12912 gnd.n12 gnd.n11 0.672012
R12913 gnd.n13 gnd.n12 0.672012
R12914 gnd.n14 gnd.n13 0.672012
R12915 gnd.n15 gnd.n14 0.672012
R12916 gnd.n16 gnd.n15 0.672012
R12917 gnd.n17 gnd.n16 0.672012
R12918 gnd.n18 gnd.n17 0.672012
R12919 gnd gnd.n0 0.665707
R12920 gnd.n3028 gnd.t119 0.637812
R12921 gnd.n3334 gnd.t197 0.637812
R12922 gnd.n4058 gnd.t38 0.637812
R12923 gnd.n5501 gnd.n5500 0.573776
R12924 gnd.n5500 gnd.n5498 0.573776
R12925 gnd.n5498 gnd.n5496 0.573776
R12926 gnd.n5496 gnd.n5494 0.573776
R12927 gnd.n5494 gnd.n5492 0.573776
R12928 gnd.n5492 gnd.n5490 0.573776
R12929 gnd.n5490 gnd.n5488 0.573776
R12930 gnd.n5516 gnd.n5515 0.573776
R12931 gnd.n5515 gnd.n5513 0.573776
R12932 gnd.n5513 gnd.n5511 0.573776
R12933 gnd.n5511 gnd.n5509 0.573776
R12934 gnd.n5509 gnd.n5507 0.573776
R12935 gnd.n5507 gnd.n5505 0.573776
R12936 gnd.n5505 gnd.n5503 0.573776
R12937 gnd.n23 gnd.n21 0.573776
R12938 gnd.n25 gnd.n23 0.573776
R12939 gnd.n27 gnd.n25 0.573776
R12940 gnd.n29 gnd.n27 0.573776
R12941 gnd.n31 gnd.n29 0.573776
R12942 gnd.n33 gnd.n31 0.573776
R12943 gnd.n34 gnd.n33 0.573776
R12944 gnd.n38 gnd.n36 0.573776
R12945 gnd.n40 gnd.n38 0.573776
R12946 gnd.n42 gnd.n40 0.573776
R12947 gnd.n44 gnd.n42 0.573776
R12948 gnd.n46 gnd.n44 0.573776
R12949 gnd.n48 gnd.n46 0.573776
R12950 gnd.n49 gnd.n48 0.573776
R12951 gnd.n7578 gnd.n7577 0.553847
R12952 gnd.n7296 gnd.n269 0.548625
R12953 gnd.n2654 gnd.n1125 0.548625
R12954 gnd.n2498 gnd.n2496 0.505073
R12955 gnd.n2536 gnd.n2535 0.505073
R12956 gnd.n7437 gnd.n7436 0.505073
R12957 gnd.n7408 gnd.n102 0.505073
R12958 gnd.n7531 gnd.n7530 0.492878
R12959 gnd.n7460 gnd.n7459 0.492878
R12960 gnd.n4426 gnd.n1494 0.492878
R12961 gnd.n1643 gnd.n1450 0.492878
R12962 gnd.n2288 gnd.n1268 0.492878
R12963 gnd.n2836 gnd.n2835 0.492878
R12964 gnd.n4829 gnd.n1008 0.492878
R12965 gnd.n2545 gnd.n965 0.492878
R12966 gnd.n6225 gnd.n6224 0.486781
R12967 gnd.n1723 gnd.n1403 0.486781
R12968 gnd.n5418 gnd.n5417 0.48678
R12969 gnd.n4662 gnd.n4661 0.485256
R12970 gnd.n6306 gnd.n6305 0.480683
R12971 gnd.n5588 gnd.n5587 0.480683
R12972 gnd.n4205 gnd.n4204 0.451719
R12973 gnd.n3199 gnd.n3198 0.451719
R12974 gnd.n6503 gnd.n726 0.425805
R12975 gnd.n6956 gnd.n6955 0.425805
R12976 gnd.n7168 gnd.n7167 0.425805
R12977 gnd.n2409 gnd.n2408 0.425805
R12978 gnd.n4664 gnd.n4663 0.406268
R12979 gnd.n4419 gnd.n1503 0.404992
R12980 gnd.n2816 gnd.n2810 0.388379
R12981 gnd.n6138 gnd.n6137 0.388379
R12982 gnd.n6106 gnd.n6105 0.388379
R12983 gnd.n6074 gnd.n6073 0.388379
R12984 gnd.n6043 gnd.n6042 0.388379
R12985 gnd.n6011 gnd.n6010 0.388379
R12986 gnd.n5979 gnd.n5978 0.388379
R12987 gnd.n5947 gnd.n5946 0.388379
R12988 gnd.n5916 gnd.n5915 0.388379
R12989 gnd.n7500 gnd.n7499 0.388379
R12990 gnd.n4870 gnd.n4869 0.388379
R12991 gnd.n4219 gnd.n4218 0.388379
R12992 gnd.n7578 gnd.n19 0.374463
R12993 gnd gnd.n7578 0.367492
R12994 gnd.n5008 gnd.t211 0.319156
R12995 gnd.n5336 gnd.n5314 0.311721
R12996 gnd.n2827 gnd.n2826 0.27489
R12997 gnd.n4230 gnd.n4228 0.27489
R12998 gnd.n6275 gnd.n6274 0.268793
R12999 gnd.n6274 gnd.n6273 0.241354
R13000 gnd.n1468 gnd.n1465 0.229039
R13001 gnd.n1471 gnd.n1468 0.229039
R13002 gnd.n2879 gnd.n2303 0.229039
R13003 gnd.n2879 gnd.n2878 0.229039
R13004 gnd.n5576 gnd.n5289 0.206293
R13005 gnd.n5534 gnd.n0 0.169152
R13006 gnd.n6155 gnd.n6127 0.155672
R13007 gnd.n6148 gnd.n6127 0.155672
R13008 gnd.n6148 gnd.n6147 0.155672
R13009 gnd.n6147 gnd.n6131 0.155672
R13010 gnd.n6140 gnd.n6131 0.155672
R13011 gnd.n6140 gnd.n6139 0.155672
R13012 gnd.n6123 gnd.n6095 0.155672
R13013 gnd.n6116 gnd.n6095 0.155672
R13014 gnd.n6116 gnd.n6115 0.155672
R13015 gnd.n6115 gnd.n6099 0.155672
R13016 gnd.n6108 gnd.n6099 0.155672
R13017 gnd.n6108 gnd.n6107 0.155672
R13018 gnd.n6091 gnd.n6063 0.155672
R13019 gnd.n6084 gnd.n6063 0.155672
R13020 gnd.n6084 gnd.n6083 0.155672
R13021 gnd.n6083 gnd.n6067 0.155672
R13022 gnd.n6076 gnd.n6067 0.155672
R13023 gnd.n6076 gnd.n6075 0.155672
R13024 gnd.n6060 gnd.n6032 0.155672
R13025 gnd.n6053 gnd.n6032 0.155672
R13026 gnd.n6053 gnd.n6052 0.155672
R13027 gnd.n6052 gnd.n6036 0.155672
R13028 gnd.n6045 gnd.n6036 0.155672
R13029 gnd.n6045 gnd.n6044 0.155672
R13030 gnd.n6028 gnd.n6000 0.155672
R13031 gnd.n6021 gnd.n6000 0.155672
R13032 gnd.n6021 gnd.n6020 0.155672
R13033 gnd.n6020 gnd.n6004 0.155672
R13034 gnd.n6013 gnd.n6004 0.155672
R13035 gnd.n6013 gnd.n6012 0.155672
R13036 gnd.n5996 gnd.n5968 0.155672
R13037 gnd.n5989 gnd.n5968 0.155672
R13038 gnd.n5989 gnd.n5988 0.155672
R13039 gnd.n5988 gnd.n5972 0.155672
R13040 gnd.n5981 gnd.n5972 0.155672
R13041 gnd.n5981 gnd.n5980 0.155672
R13042 gnd.n5964 gnd.n5936 0.155672
R13043 gnd.n5957 gnd.n5936 0.155672
R13044 gnd.n5957 gnd.n5956 0.155672
R13045 gnd.n5956 gnd.n5940 0.155672
R13046 gnd.n5949 gnd.n5940 0.155672
R13047 gnd.n5949 gnd.n5948 0.155672
R13048 gnd.n5933 gnd.n5905 0.155672
R13049 gnd.n5926 gnd.n5905 0.155672
R13050 gnd.n5926 gnd.n5925 0.155672
R13051 gnd.n5925 gnd.n5909 0.155672
R13052 gnd.n5918 gnd.n5909 0.155672
R13053 gnd.n5918 gnd.n5917 0.155672
R13054 gnd.n6305 gnd.n4912 0.152939
R13055 gnd.n4914 gnd.n4912 0.152939
R13056 gnd.n4918 gnd.n4914 0.152939
R13057 gnd.n4919 gnd.n4918 0.152939
R13058 gnd.n4920 gnd.n4919 0.152939
R13059 gnd.n4921 gnd.n4920 0.152939
R13060 gnd.n4925 gnd.n4921 0.152939
R13061 gnd.n4926 gnd.n4925 0.152939
R13062 gnd.n4927 gnd.n4926 0.152939
R13063 gnd.n4928 gnd.n4927 0.152939
R13064 gnd.n4932 gnd.n4928 0.152939
R13065 gnd.n4933 gnd.n4932 0.152939
R13066 gnd.n4934 gnd.n4933 0.152939
R13067 gnd.n4935 gnd.n4934 0.152939
R13068 gnd.n4940 gnd.n4935 0.152939
R13069 gnd.n6275 gnd.n4940 0.152939
R13070 gnd.n5589 gnd.n5588 0.152939
R13071 gnd.n5589 gnd.n5207 0.152939
R13072 gnd.n5617 gnd.n5207 0.152939
R13073 gnd.n5618 gnd.n5617 0.152939
R13074 gnd.n5619 gnd.n5618 0.152939
R13075 gnd.n5620 gnd.n5619 0.152939
R13076 gnd.n5620 gnd.n5181 0.152939
R13077 gnd.n5648 gnd.n5181 0.152939
R13078 gnd.n5649 gnd.n5648 0.152939
R13079 gnd.n5650 gnd.n5649 0.152939
R13080 gnd.n5651 gnd.n5650 0.152939
R13081 gnd.n5651 gnd.n5156 0.152939
R13082 gnd.n5679 gnd.n5156 0.152939
R13083 gnd.n5680 gnd.n5679 0.152939
R13084 gnd.n5681 gnd.n5680 0.152939
R13085 gnd.n5682 gnd.n5681 0.152939
R13086 gnd.n5682 gnd.n5130 0.152939
R13087 gnd.n5710 gnd.n5130 0.152939
R13088 gnd.n5711 gnd.n5710 0.152939
R13089 gnd.n5712 gnd.n5711 0.152939
R13090 gnd.n5713 gnd.n5712 0.152939
R13091 gnd.n5713 gnd.n5106 0.152939
R13092 gnd.n5740 gnd.n5106 0.152939
R13093 gnd.n5741 gnd.n5740 0.152939
R13094 gnd.n5742 gnd.n5741 0.152939
R13095 gnd.n5743 gnd.n5742 0.152939
R13096 gnd.n5743 gnd.n5075 0.152939
R13097 gnd.n5794 gnd.n5075 0.152939
R13098 gnd.n5795 gnd.n5794 0.152939
R13099 gnd.n5796 gnd.n5795 0.152939
R13100 gnd.n5796 gnd.n5054 0.152939
R13101 gnd.n5824 gnd.n5054 0.152939
R13102 gnd.n5825 gnd.n5824 0.152939
R13103 gnd.n5826 gnd.n5825 0.152939
R13104 gnd.n5827 gnd.n5826 0.152939
R13105 gnd.n5827 gnd.n5030 0.152939
R13106 gnd.n5870 gnd.n5030 0.152939
R13107 gnd.n5871 gnd.n5870 0.152939
R13108 gnd.n5872 gnd.n5871 0.152939
R13109 gnd.n5873 gnd.n5872 0.152939
R13110 gnd.n5873 gnd.n5000 0.152939
R13111 gnd.n6191 gnd.n5000 0.152939
R13112 gnd.n6192 gnd.n6191 0.152939
R13113 gnd.n6193 gnd.n6192 0.152939
R13114 gnd.n6194 gnd.n6193 0.152939
R13115 gnd.n6196 gnd.n6194 0.152939
R13116 gnd.n6196 gnd.n6195 0.152939
R13117 gnd.n6195 gnd.n914 0.152939
R13118 gnd.n915 gnd.n914 0.152939
R13119 gnd.n916 gnd.n915 0.152939
R13120 gnd.n4910 gnd.n916 0.152939
R13121 gnd.n4911 gnd.n4910 0.152939
R13122 gnd.n6306 gnd.n4911 0.152939
R13123 gnd.n5587 gnd.n5231 0.152939
R13124 gnd.n5252 gnd.n5231 0.152939
R13125 gnd.n5253 gnd.n5252 0.152939
R13126 gnd.n5259 gnd.n5253 0.152939
R13127 gnd.n5260 gnd.n5259 0.152939
R13128 gnd.n5261 gnd.n5260 0.152939
R13129 gnd.n5261 gnd.n5250 0.152939
R13130 gnd.n5269 gnd.n5250 0.152939
R13131 gnd.n5270 gnd.n5269 0.152939
R13132 gnd.n5271 gnd.n5270 0.152939
R13133 gnd.n5271 gnd.n5248 0.152939
R13134 gnd.n5279 gnd.n5248 0.152939
R13135 gnd.n5280 gnd.n5279 0.152939
R13136 gnd.n5281 gnd.n5280 0.152939
R13137 gnd.n5281 gnd.n5246 0.152939
R13138 gnd.n5289 gnd.n5246 0.152939
R13139 gnd.n6273 gnd.n4942 0.152939
R13140 gnd.n4944 gnd.n4942 0.152939
R13141 gnd.n4948 gnd.n4944 0.152939
R13142 gnd.n4949 gnd.n4948 0.152939
R13143 gnd.n4950 gnd.n4949 0.152939
R13144 gnd.n4951 gnd.n4950 0.152939
R13145 gnd.n4955 gnd.n4951 0.152939
R13146 gnd.n4956 gnd.n4955 0.152939
R13147 gnd.n4957 gnd.n4956 0.152939
R13148 gnd.n4958 gnd.n4957 0.152939
R13149 gnd.n4962 gnd.n4958 0.152939
R13150 gnd.n4963 gnd.n4962 0.152939
R13151 gnd.n4964 gnd.n4963 0.152939
R13152 gnd.n4965 gnd.n4964 0.152939
R13153 gnd.n4969 gnd.n4965 0.152939
R13154 gnd.n4970 gnd.n4969 0.152939
R13155 gnd.n4971 gnd.n4970 0.152939
R13156 gnd.n4972 gnd.n4971 0.152939
R13157 gnd.n4976 gnd.n4972 0.152939
R13158 gnd.n4977 gnd.n4976 0.152939
R13159 gnd.n4978 gnd.n4977 0.152939
R13160 gnd.n4979 gnd.n4978 0.152939
R13161 gnd.n4986 gnd.n4979 0.152939
R13162 gnd.n4987 gnd.n4986 0.152939
R13163 gnd.n4988 gnd.n4987 0.152939
R13164 gnd.n6225 gnd.n4988 0.152939
R13165 gnd.n5760 gnd.n5092 0.152939
R13166 gnd.n5761 gnd.n5760 0.152939
R13167 gnd.n5762 gnd.n5761 0.152939
R13168 gnd.n5763 gnd.n5762 0.152939
R13169 gnd.n5764 gnd.n5763 0.152939
R13170 gnd.n5765 gnd.n5764 0.152939
R13171 gnd.n5766 gnd.n5765 0.152939
R13172 gnd.n5767 gnd.n5766 0.152939
R13173 gnd.n5768 gnd.n5767 0.152939
R13174 gnd.n5768 gnd.n5036 0.152939
R13175 gnd.n5847 gnd.n5036 0.152939
R13176 gnd.n5848 gnd.n5847 0.152939
R13177 gnd.n5849 gnd.n5848 0.152939
R13178 gnd.n5850 gnd.n5849 0.152939
R13179 gnd.n5851 gnd.n5850 0.152939
R13180 gnd.n5852 gnd.n5851 0.152939
R13181 gnd.n5853 gnd.n5852 0.152939
R13182 gnd.n5854 gnd.n5853 0.152939
R13183 gnd.n5854 gnd.n4993 0.152939
R13184 gnd.n6206 gnd.n4993 0.152939
R13185 gnd.n6207 gnd.n6206 0.152939
R13186 gnd.n6208 gnd.n6207 0.152939
R13187 gnd.n6208 gnd.n4991 0.152939
R13188 gnd.n6216 gnd.n4991 0.152939
R13189 gnd.n6217 gnd.n6216 0.152939
R13190 gnd.n6218 gnd.n6217 0.152939
R13191 gnd.n6218 gnd.n4989 0.152939
R13192 gnd.n6224 gnd.n4989 0.152939
R13193 gnd.n5419 gnd.n5418 0.152939
R13194 gnd.n5419 gnd.n5309 0.152939
R13195 gnd.n5434 gnd.n5309 0.152939
R13196 gnd.n5435 gnd.n5434 0.152939
R13197 gnd.n5436 gnd.n5435 0.152939
R13198 gnd.n5436 gnd.n5297 0.152939
R13199 gnd.n5450 gnd.n5297 0.152939
R13200 gnd.n5451 gnd.n5450 0.152939
R13201 gnd.n5452 gnd.n5451 0.152939
R13202 gnd.n5453 gnd.n5452 0.152939
R13203 gnd.n5454 gnd.n5453 0.152939
R13204 gnd.n5455 gnd.n5454 0.152939
R13205 gnd.n5456 gnd.n5455 0.152939
R13206 gnd.n5457 gnd.n5456 0.152939
R13207 gnd.n5458 gnd.n5457 0.152939
R13208 gnd.n5459 gnd.n5458 0.152939
R13209 gnd.n5460 gnd.n5459 0.152939
R13210 gnd.n5461 gnd.n5460 0.152939
R13211 gnd.n5462 gnd.n5461 0.152939
R13212 gnd.n5463 gnd.n5462 0.152939
R13213 gnd.n5464 gnd.n5463 0.152939
R13214 gnd.n5465 gnd.n5464 0.152939
R13215 gnd.n5466 gnd.n5465 0.152939
R13216 gnd.n5467 gnd.n5466 0.152939
R13217 gnd.n5468 gnd.n5467 0.152939
R13218 gnd.n5469 gnd.n5468 0.152939
R13219 gnd.n5470 gnd.n5469 0.152939
R13220 gnd.n5471 gnd.n5470 0.152939
R13221 gnd.n5337 gnd.n5336 0.152939
R13222 gnd.n5338 gnd.n5337 0.152939
R13223 gnd.n5339 gnd.n5338 0.152939
R13224 gnd.n5340 gnd.n5339 0.152939
R13225 gnd.n5341 gnd.n5340 0.152939
R13226 gnd.n5342 gnd.n5341 0.152939
R13227 gnd.n5343 gnd.n5342 0.152939
R13228 gnd.n5344 gnd.n5343 0.152939
R13229 gnd.n5345 gnd.n5344 0.152939
R13230 gnd.n5346 gnd.n5345 0.152939
R13231 gnd.n5347 gnd.n5346 0.152939
R13232 gnd.n5348 gnd.n5347 0.152939
R13233 gnd.n5349 gnd.n5348 0.152939
R13234 gnd.n5350 gnd.n5349 0.152939
R13235 gnd.n5351 gnd.n5350 0.152939
R13236 gnd.n5352 gnd.n5351 0.152939
R13237 gnd.n5353 gnd.n5352 0.152939
R13238 gnd.n5354 gnd.n5353 0.152939
R13239 gnd.n5355 gnd.n5354 0.152939
R13240 gnd.n5356 gnd.n5355 0.152939
R13241 gnd.n5357 gnd.n5356 0.152939
R13242 gnd.n5358 gnd.n5357 0.152939
R13243 gnd.n5362 gnd.n5358 0.152939
R13244 gnd.n5363 gnd.n5362 0.152939
R13245 gnd.n5363 gnd.n5320 0.152939
R13246 gnd.n5417 gnd.n5320 0.152939
R13247 gnd.n6504 gnd.n6503 0.152939
R13248 gnd.n6505 gnd.n6504 0.152939
R13249 gnd.n6505 gnd.n720 0.152939
R13250 gnd.n6513 gnd.n720 0.152939
R13251 gnd.n6514 gnd.n6513 0.152939
R13252 gnd.n6515 gnd.n6514 0.152939
R13253 gnd.n6515 gnd.n714 0.152939
R13254 gnd.n6523 gnd.n714 0.152939
R13255 gnd.n6524 gnd.n6523 0.152939
R13256 gnd.n6525 gnd.n6524 0.152939
R13257 gnd.n6525 gnd.n708 0.152939
R13258 gnd.n6533 gnd.n708 0.152939
R13259 gnd.n6534 gnd.n6533 0.152939
R13260 gnd.n6535 gnd.n6534 0.152939
R13261 gnd.n6535 gnd.n702 0.152939
R13262 gnd.n6543 gnd.n702 0.152939
R13263 gnd.n6544 gnd.n6543 0.152939
R13264 gnd.n6545 gnd.n6544 0.152939
R13265 gnd.n6545 gnd.n696 0.152939
R13266 gnd.n6553 gnd.n696 0.152939
R13267 gnd.n6554 gnd.n6553 0.152939
R13268 gnd.n6555 gnd.n6554 0.152939
R13269 gnd.n6555 gnd.n690 0.152939
R13270 gnd.n6563 gnd.n690 0.152939
R13271 gnd.n6564 gnd.n6563 0.152939
R13272 gnd.n6565 gnd.n6564 0.152939
R13273 gnd.n6565 gnd.n684 0.152939
R13274 gnd.n6573 gnd.n684 0.152939
R13275 gnd.n6574 gnd.n6573 0.152939
R13276 gnd.n6575 gnd.n6574 0.152939
R13277 gnd.n6575 gnd.n678 0.152939
R13278 gnd.n6583 gnd.n678 0.152939
R13279 gnd.n6584 gnd.n6583 0.152939
R13280 gnd.n6585 gnd.n6584 0.152939
R13281 gnd.n6585 gnd.n672 0.152939
R13282 gnd.n6593 gnd.n672 0.152939
R13283 gnd.n6594 gnd.n6593 0.152939
R13284 gnd.n6595 gnd.n6594 0.152939
R13285 gnd.n6595 gnd.n666 0.152939
R13286 gnd.n6603 gnd.n666 0.152939
R13287 gnd.n6604 gnd.n6603 0.152939
R13288 gnd.n6605 gnd.n6604 0.152939
R13289 gnd.n6605 gnd.n660 0.152939
R13290 gnd.n6613 gnd.n660 0.152939
R13291 gnd.n6614 gnd.n6613 0.152939
R13292 gnd.n6615 gnd.n6614 0.152939
R13293 gnd.n6615 gnd.n654 0.152939
R13294 gnd.n6623 gnd.n654 0.152939
R13295 gnd.n6624 gnd.n6623 0.152939
R13296 gnd.n6625 gnd.n6624 0.152939
R13297 gnd.n6625 gnd.n648 0.152939
R13298 gnd.n6633 gnd.n648 0.152939
R13299 gnd.n6634 gnd.n6633 0.152939
R13300 gnd.n6635 gnd.n6634 0.152939
R13301 gnd.n6635 gnd.n642 0.152939
R13302 gnd.n6643 gnd.n642 0.152939
R13303 gnd.n6644 gnd.n6643 0.152939
R13304 gnd.n6645 gnd.n6644 0.152939
R13305 gnd.n6645 gnd.n636 0.152939
R13306 gnd.n6653 gnd.n636 0.152939
R13307 gnd.n6654 gnd.n6653 0.152939
R13308 gnd.n6655 gnd.n6654 0.152939
R13309 gnd.n6655 gnd.n630 0.152939
R13310 gnd.n6663 gnd.n630 0.152939
R13311 gnd.n6664 gnd.n6663 0.152939
R13312 gnd.n6665 gnd.n6664 0.152939
R13313 gnd.n6665 gnd.n624 0.152939
R13314 gnd.n6673 gnd.n624 0.152939
R13315 gnd.n6674 gnd.n6673 0.152939
R13316 gnd.n6675 gnd.n6674 0.152939
R13317 gnd.n6675 gnd.n618 0.152939
R13318 gnd.n6683 gnd.n618 0.152939
R13319 gnd.n6684 gnd.n6683 0.152939
R13320 gnd.n6685 gnd.n6684 0.152939
R13321 gnd.n6685 gnd.n612 0.152939
R13322 gnd.n6693 gnd.n612 0.152939
R13323 gnd.n6694 gnd.n6693 0.152939
R13324 gnd.n6695 gnd.n6694 0.152939
R13325 gnd.n6695 gnd.n606 0.152939
R13326 gnd.n6703 gnd.n606 0.152939
R13327 gnd.n6704 gnd.n6703 0.152939
R13328 gnd.n6705 gnd.n6704 0.152939
R13329 gnd.n6705 gnd.n600 0.152939
R13330 gnd.n6713 gnd.n600 0.152939
R13331 gnd.n6714 gnd.n6713 0.152939
R13332 gnd.n6715 gnd.n6714 0.152939
R13333 gnd.n6715 gnd.n594 0.152939
R13334 gnd.n6723 gnd.n594 0.152939
R13335 gnd.n6724 gnd.n6723 0.152939
R13336 gnd.n6725 gnd.n6724 0.152939
R13337 gnd.n6725 gnd.n588 0.152939
R13338 gnd.n6733 gnd.n588 0.152939
R13339 gnd.n6734 gnd.n6733 0.152939
R13340 gnd.n6735 gnd.n6734 0.152939
R13341 gnd.n6735 gnd.n582 0.152939
R13342 gnd.n6743 gnd.n582 0.152939
R13343 gnd.n6744 gnd.n6743 0.152939
R13344 gnd.n6745 gnd.n6744 0.152939
R13345 gnd.n6745 gnd.n576 0.152939
R13346 gnd.n6753 gnd.n576 0.152939
R13347 gnd.n6754 gnd.n6753 0.152939
R13348 gnd.n6755 gnd.n6754 0.152939
R13349 gnd.n6755 gnd.n570 0.152939
R13350 gnd.n6763 gnd.n570 0.152939
R13351 gnd.n6764 gnd.n6763 0.152939
R13352 gnd.n6765 gnd.n6764 0.152939
R13353 gnd.n6765 gnd.n564 0.152939
R13354 gnd.n6773 gnd.n564 0.152939
R13355 gnd.n6774 gnd.n6773 0.152939
R13356 gnd.n6775 gnd.n6774 0.152939
R13357 gnd.n6775 gnd.n558 0.152939
R13358 gnd.n6783 gnd.n558 0.152939
R13359 gnd.n6784 gnd.n6783 0.152939
R13360 gnd.n6785 gnd.n6784 0.152939
R13361 gnd.n6785 gnd.n552 0.152939
R13362 gnd.n6793 gnd.n552 0.152939
R13363 gnd.n6794 gnd.n6793 0.152939
R13364 gnd.n6795 gnd.n6794 0.152939
R13365 gnd.n6795 gnd.n546 0.152939
R13366 gnd.n6803 gnd.n546 0.152939
R13367 gnd.n6804 gnd.n6803 0.152939
R13368 gnd.n6805 gnd.n6804 0.152939
R13369 gnd.n6805 gnd.n540 0.152939
R13370 gnd.n6813 gnd.n540 0.152939
R13371 gnd.n6814 gnd.n6813 0.152939
R13372 gnd.n6815 gnd.n6814 0.152939
R13373 gnd.n6815 gnd.n534 0.152939
R13374 gnd.n6823 gnd.n534 0.152939
R13375 gnd.n6824 gnd.n6823 0.152939
R13376 gnd.n6825 gnd.n6824 0.152939
R13377 gnd.n6825 gnd.n528 0.152939
R13378 gnd.n6833 gnd.n528 0.152939
R13379 gnd.n6834 gnd.n6833 0.152939
R13380 gnd.n6835 gnd.n6834 0.152939
R13381 gnd.n6835 gnd.n522 0.152939
R13382 gnd.n6843 gnd.n522 0.152939
R13383 gnd.n6844 gnd.n6843 0.152939
R13384 gnd.n6845 gnd.n6844 0.152939
R13385 gnd.n6845 gnd.n516 0.152939
R13386 gnd.n6853 gnd.n516 0.152939
R13387 gnd.n6854 gnd.n6853 0.152939
R13388 gnd.n6855 gnd.n6854 0.152939
R13389 gnd.n6855 gnd.n510 0.152939
R13390 gnd.n6863 gnd.n510 0.152939
R13391 gnd.n6864 gnd.n6863 0.152939
R13392 gnd.n6865 gnd.n6864 0.152939
R13393 gnd.n6865 gnd.n504 0.152939
R13394 gnd.n6873 gnd.n504 0.152939
R13395 gnd.n6874 gnd.n6873 0.152939
R13396 gnd.n6875 gnd.n6874 0.152939
R13397 gnd.n6875 gnd.n498 0.152939
R13398 gnd.n6883 gnd.n498 0.152939
R13399 gnd.n6884 gnd.n6883 0.152939
R13400 gnd.n6885 gnd.n6884 0.152939
R13401 gnd.n6885 gnd.n492 0.152939
R13402 gnd.n6893 gnd.n492 0.152939
R13403 gnd.n6894 gnd.n6893 0.152939
R13404 gnd.n6895 gnd.n6894 0.152939
R13405 gnd.n6895 gnd.n486 0.152939
R13406 gnd.n6903 gnd.n486 0.152939
R13407 gnd.n6904 gnd.n6903 0.152939
R13408 gnd.n6905 gnd.n6904 0.152939
R13409 gnd.n6905 gnd.n480 0.152939
R13410 gnd.n6913 gnd.n480 0.152939
R13411 gnd.n6914 gnd.n6913 0.152939
R13412 gnd.n6915 gnd.n6914 0.152939
R13413 gnd.n6915 gnd.n474 0.152939
R13414 gnd.n6923 gnd.n474 0.152939
R13415 gnd.n6924 gnd.n6923 0.152939
R13416 gnd.n6925 gnd.n6924 0.152939
R13417 gnd.n6925 gnd.n468 0.152939
R13418 gnd.n6933 gnd.n468 0.152939
R13419 gnd.n6934 gnd.n6933 0.152939
R13420 gnd.n6935 gnd.n6934 0.152939
R13421 gnd.n6935 gnd.n462 0.152939
R13422 gnd.n6943 gnd.n462 0.152939
R13423 gnd.n6944 gnd.n6943 0.152939
R13424 gnd.n6946 gnd.n6944 0.152939
R13425 gnd.n6946 gnd.n6945 0.152939
R13426 gnd.n6945 gnd.n456 0.152939
R13427 gnd.n6955 gnd.n456 0.152939
R13428 gnd.n6956 gnd.n451 0.152939
R13429 gnd.n6964 gnd.n451 0.152939
R13430 gnd.n6965 gnd.n6964 0.152939
R13431 gnd.n6966 gnd.n6965 0.152939
R13432 gnd.n6966 gnd.n445 0.152939
R13433 gnd.n6974 gnd.n445 0.152939
R13434 gnd.n6975 gnd.n6974 0.152939
R13435 gnd.n6976 gnd.n6975 0.152939
R13436 gnd.n6976 gnd.n439 0.152939
R13437 gnd.n6984 gnd.n439 0.152939
R13438 gnd.n6985 gnd.n6984 0.152939
R13439 gnd.n6986 gnd.n6985 0.152939
R13440 gnd.n6986 gnd.n433 0.152939
R13441 gnd.n6994 gnd.n433 0.152939
R13442 gnd.n6995 gnd.n6994 0.152939
R13443 gnd.n6996 gnd.n6995 0.152939
R13444 gnd.n6996 gnd.n427 0.152939
R13445 gnd.n7004 gnd.n427 0.152939
R13446 gnd.n7005 gnd.n7004 0.152939
R13447 gnd.n7006 gnd.n7005 0.152939
R13448 gnd.n7006 gnd.n421 0.152939
R13449 gnd.n7014 gnd.n421 0.152939
R13450 gnd.n7015 gnd.n7014 0.152939
R13451 gnd.n7016 gnd.n7015 0.152939
R13452 gnd.n7016 gnd.n415 0.152939
R13453 gnd.n7024 gnd.n415 0.152939
R13454 gnd.n7025 gnd.n7024 0.152939
R13455 gnd.n7026 gnd.n7025 0.152939
R13456 gnd.n7026 gnd.n409 0.152939
R13457 gnd.n7034 gnd.n409 0.152939
R13458 gnd.n7035 gnd.n7034 0.152939
R13459 gnd.n7036 gnd.n7035 0.152939
R13460 gnd.n7036 gnd.n403 0.152939
R13461 gnd.n7044 gnd.n403 0.152939
R13462 gnd.n7045 gnd.n7044 0.152939
R13463 gnd.n7046 gnd.n7045 0.152939
R13464 gnd.n7046 gnd.n397 0.152939
R13465 gnd.n7054 gnd.n397 0.152939
R13466 gnd.n7055 gnd.n7054 0.152939
R13467 gnd.n7056 gnd.n7055 0.152939
R13468 gnd.n7056 gnd.n391 0.152939
R13469 gnd.n7064 gnd.n391 0.152939
R13470 gnd.n7065 gnd.n7064 0.152939
R13471 gnd.n7066 gnd.n7065 0.152939
R13472 gnd.n7066 gnd.n385 0.152939
R13473 gnd.n7074 gnd.n385 0.152939
R13474 gnd.n7075 gnd.n7074 0.152939
R13475 gnd.n7076 gnd.n7075 0.152939
R13476 gnd.n7076 gnd.n379 0.152939
R13477 gnd.n7084 gnd.n379 0.152939
R13478 gnd.n7085 gnd.n7084 0.152939
R13479 gnd.n7086 gnd.n7085 0.152939
R13480 gnd.n7086 gnd.n373 0.152939
R13481 gnd.n7094 gnd.n373 0.152939
R13482 gnd.n7095 gnd.n7094 0.152939
R13483 gnd.n7096 gnd.n7095 0.152939
R13484 gnd.n7096 gnd.n367 0.152939
R13485 gnd.n7104 gnd.n367 0.152939
R13486 gnd.n7105 gnd.n7104 0.152939
R13487 gnd.n7106 gnd.n7105 0.152939
R13488 gnd.n7106 gnd.n361 0.152939
R13489 gnd.n7114 gnd.n361 0.152939
R13490 gnd.n7115 gnd.n7114 0.152939
R13491 gnd.n7116 gnd.n7115 0.152939
R13492 gnd.n7116 gnd.n355 0.152939
R13493 gnd.n7124 gnd.n355 0.152939
R13494 gnd.n7125 gnd.n7124 0.152939
R13495 gnd.n7126 gnd.n7125 0.152939
R13496 gnd.n7126 gnd.n349 0.152939
R13497 gnd.n7134 gnd.n349 0.152939
R13498 gnd.n7135 gnd.n7134 0.152939
R13499 gnd.n7136 gnd.n7135 0.152939
R13500 gnd.n7136 gnd.n343 0.152939
R13501 gnd.n7144 gnd.n343 0.152939
R13502 gnd.n7145 gnd.n7144 0.152939
R13503 gnd.n7146 gnd.n7145 0.152939
R13504 gnd.n7146 gnd.n337 0.152939
R13505 gnd.n7154 gnd.n337 0.152939
R13506 gnd.n7155 gnd.n7154 0.152939
R13507 gnd.n7156 gnd.n7155 0.152939
R13508 gnd.n7156 gnd.n331 0.152939
R13509 gnd.n7165 gnd.n331 0.152939
R13510 gnd.n7166 gnd.n7165 0.152939
R13511 gnd.n7168 gnd.n7166 0.152939
R13512 gnd.n327 gnd.n326 0.152939
R13513 gnd.n7167 gnd.n327 0.152939
R13514 gnd.n7310 gnd.n253 0.152939
R13515 gnd.n7311 gnd.n7310 0.152939
R13516 gnd.n7312 gnd.n7311 0.152939
R13517 gnd.n7312 gnd.n235 0.152939
R13518 gnd.n7326 gnd.n235 0.152939
R13519 gnd.n7327 gnd.n7326 0.152939
R13520 gnd.n7328 gnd.n7327 0.152939
R13521 gnd.n7328 gnd.n222 0.152939
R13522 gnd.n7342 gnd.n222 0.152939
R13523 gnd.n7343 gnd.n7342 0.152939
R13524 gnd.n7344 gnd.n7343 0.152939
R13525 gnd.n7344 gnd.n205 0.152939
R13526 gnd.n7358 gnd.n205 0.152939
R13527 gnd.n7359 gnd.n7358 0.152939
R13528 gnd.n7360 gnd.n7359 0.152939
R13529 gnd.n7360 gnd.n190 0.152939
R13530 gnd.n7449 gnd.n190 0.152939
R13531 gnd.n7450 gnd.n7449 0.152939
R13532 gnd.n7451 gnd.n7450 0.152939
R13533 gnd.n7451 gnd.n111 0.152939
R13534 gnd.n7531 gnd.n111 0.152939
R13535 gnd.n7530 gnd.n112 0.152939
R13536 gnd.n114 gnd.n112 0.152939
R13537 gnd.n118 gnd.n114 0.152939
R13538 gnd.n119 gnd.n118 0.152939
R13539 gnd.n120 gnd.n119 0.152939
R13540 gnd.n121 gnd.n120 0.152939
R13541 gnd.n125 gnd.n121 0.152939
R13542 gnd.n126 gnd.n125 0.152939
R13543 gnd.n127 gnd.n126 0.152939
R13544 gnd.n128 gnd.n127 0.152939
R13545 gnd.n132 gnd.n128 0.152939
R13546 gnd.n133 gnd.n132 0.152939
R13547 gnd.n134 gnd.n133 0.152939
R13548 gnd.n135 gnd.n134 0.152939
R13549 gnd.n139 gnd.n135 0.152939
R13550 gnd.n140 gnd.n139 0.152939
R13551 gnd.n141 gnd.n140 0.152939
R13552 gnd.n142 gnd.n141 0.152939
R13553 gnd.n146 gnd.n142 0.152939
R13554 gnd.n147 gnd.n146 0.152939
R13555 gnd.n148 gnd.n147 0.152939
R13556 gnd.n149 gnd.n148 0.152939
R13557 gnd.n153 gnd.n149 0.152939
R13558 gnd.n154 gnd.n153 0.152939
R13559 gnd.n155 gnd.n154 0.152939
R13560 gnd.n156 gnd.n155 0.152939
R13561 gnd.n160 gnd.n156 0.152939
R13562 gnd.n161 gnd.n160 0.152939
R13563 gnd.n162 gnd.n161 0.152939
R13564 gnd.n163 gnd.n162 0.152939
R13565 gnd.n167 gnd.n163 0.152939
R13566 gnd.n168 gnd.n167 0.152939
R13567 gnd.n169 gnd.n168 0.152939
R13568 gnd.n170 gnd.n169 0.152939
R13569 gnd.n174 gnd.n170 0.152939
R13570 gnd.n175 gnd.n174 0.152939
R13571 gnd.n7461 gnd.n175 0.152939
R13572 gnd.n7461 gnd.n7460 0.152939
R13573 gnd.n1649 gnd.n1494 0.152939
R13574 gnd.n1650 gnd.n1649 0.152939
R13575 gnd.n1651 gnd.n1650 0.152939
R13576 gnd.n1652 gnd.n1651 0.152939
R13577 gnd.n1653 gnd.n1652 0.152939
R13578 gnd.n1654 gnd.n1653 0.152939
R13579 gnd.n1655 gnd.n1654 0.152939
R13580 gnd.n1656 gnd.n1655 0.152939
R13581 gnd.n1657 gnd.n1656 0.152939
R13582 gnd.n1658 gnd.n1657 0.152939
R13583 gnd.n1659 gnd.n1658 0.152939
R13584 gnd.n1660 gnd.n1659 0.152939
R13585 gnd.n1661 gnd.n1660 0.152939
R13586 gnd.n1661 gnd.n1557 0.152939
R13587 gnd.n4329 gnd.n1557 0.152939
R13588 gnd.n4330 gnd.n4329 0.152939
R13589 gnd.n4331 gnd.n4330 0.152939
R13590 gnd.n4331 gnd.n1555 0.152939
R13591 gnd.n4336 gnd.n1555 0.152939
R13592 gnd.n4337 gnd.n4336 0.152939
R13593 gnd.n4338 gnd.n4337 0.152939
R13594 gnd.n4339 gnd.n4338 0.152939
R13595 gnd.n4340 gnd.n4339 0.152939
R13596 gnd.n4342 gnd.n4340 0.152939
R13597 gnd.n4342 gnd.n4341 0.152939
R13598 gnd.n4341 gnd.n300 0.152939
R13599 gnd.n7210 gnd.n7209 0.152939
R13600 gnd.n7211 gnd.n7210 0.152939
R13601 gnd.n7212 gnd.n7211 0.152939
R13602 gnd.n7213 gnd.n7212 0.152939
R13603 gnd.n7214 gnd.n7213 0.152939
R13604 gnd.n7215 gnd.n7214 0.152939
R13605 gnd.n7216 gnd.n7215 0.152939
R13606 gnd.n7217 gnd.n7216 0.152939
R13607 gnd.n7218 gnd.n7217 0.152939
R13608 gnd.n7219 gnd.n7218 0.152939
R13609 gnd.n7220 gnd.n7219 0.152939
R13610 gnd.n7221 gnd.n7220 0.152939
R13611 gnd.n7222 gnd.n7221 0.152939
R13612 gnd.n7223 gnd.n7222 0.152939
R13613 gnd.n7224 gnd.n7223 0.152939
R13614 gnd.n7225 gnd.n7224 0.152939
R13615 gnd.n7226 gnd.n7225 0.152939
R13616 gnd.n7227 gnd.n7226 0.152939
R13617 gnd.n7228 gnd.n7227 0.152939
R13618 gnd.n7229 gnd.n7228 0.152939
R13619 gnd.n7230 gnd.n7229 0.152939
R13620 gnd.n7231 gnd.n7230 0.152939
R13621 gnd.n7233 gnd.n7231 0.152939
R13622 gnd.n7233 gnd.n7232 0.152939
R13623 gnd.n7232 gnd.n181 0.152939
R13624 gnd.n7459 gnd.n181 0.152939
R13625 gnd.n1451 gnd.n1450 0.152939
R13626 gnd.n1452 gnd.n1451 0.152939
R13627 gnd.n1453 gnd.n1452 0.152939
R13628 gnd.n1454 gnd.n1453 0.152939
R13629 gnd.n1455 gnd.n1454 0.152939
R13630 gnd.n1456 gnd.n1455 0.152939
R13631 gnd.n1457 gnd.n1456 0.152939
R13632 gnd.n1458 gnd.n1457 0.152939
R13633 gnd.n1459 gnd.n1458 0.152939
R13634 gnd.n1460 gnd.n1459 0.152939
R13635 gnd.n1461 gnd.n1460 0.152939
R13636 gnd.n1462 gnd.n1461 0.152939
R13637 gnd.n1463 gnd.n1462 0.152939
R13638 gnd.n1464 gnd.n1463 0.152939
R13639 gnd.n1465 gnd.n1464 0.152939
R13640 gnd.n1472 gnd.n1471 0.152939
R13641 gnd.n1473 gnd.n1472 0.152939
R13642 gnd.n1474 gnd.n1473 0.152939
R13643 gnd.n1475 gnd.n1474 0.152939
R13644 gnd.n1476 gnd.n1475 0.152939
R13645 gnd.n1477 gnd.n1476 0.152939
R13646 gnd.n1478 gnd.n1477 0.152939
R13647 gnd.n1479 gnd.n1478 0.152939
R13648 gnd.n1480 gnd.n1479 0.152939
R13649 gnd.n1481 gnd.n1480 0.152939
R13650 gnd.n1482 gnd.n1481 0.152939
R13651 gnd.n1483 gnd.n1482 0.152939
R13652 gnd.n1484 gnd.n1483 0.152939
R13653 gnd.n1485 gnd.n1484 0.152939
R13654 gnd.n1486 gnd.n1485 0.152939
R13655 gnd.n1487 gnd.n1486 0.152939
R13656 gnd.n1488 gnd.n1487 0.152939
R13657 gnd.n4428 gnd.n1488 0.152939
R13658 gnd.n4428 gnd.n4427 0.152939
R13659 gnd.n4427 gnd.n4426 0.152939
R13660 gnd.n1644 gnd.n1643 0.152939
R13661 gnd.n1644 gnd.n1622 0.152939
R13662 gnd.n4251 gnd.n1622 0.152939
R13663 gnd.n4252 gnd.n4251 0.152939
R13664 gnd.n4253 gnd.n4252 0.152939
R13665 gnd.n4254 gnd.n4253 0.152939
R13666 gnd.n4254 gnd.n1594 0.152939
R13667 gnd.n4282 gnd.n1594 0.152939
R13668 gnd.n4283 gnd.n4282 0.152939
R13669 gnd.n4284 gnd.n4283 0.152939
R13670 gnd.n4285 gnd.n4284 0.152939
R13671 gnd.n4285 gnd.n1567 0.152939
R13672 gnd.n4319 gnd.n1567 0.152939
R13673 gnd.n4320 gnd.n4319 0.152939
R13674 gnd.n4321 gnd.n4320 0.152939
R13675 gnd.n4322 gnd.n4321 0.152939
R13676 gnd.n4322 gnd.n1532 0.152939
R13677 gnd.n4382 gnd.n1532 0.152939
R13678 gnd.n4383 gnd.n4382 0.152939
R13679 gnd.n4384 gnd.n4383 0.152939
R13680 gnd.n4384 gnd.n268 0.152939
R13681 gnd.n2400 gnd.n2383 0.152939
R13682 gnd.n2386 gnd.n2383 0.152939
R13683 gnd.n2387 gnd.n2386 0.152939
R13684 gnd.n2388 gnd.n2387 0.152939
R13685 gnd.n2390 gnd.n2388 0.152939
R13686 gnd.n2390 gnd.n2389 0.152939
R13687 gnd.n2389 gnd.n2350 0.152939
R13688 gnd.n2729 gnd.n2350 0.152939
R13689 gnd.n2730 gnd.n2729 0.152939
R13690 gnd.n2731 gnd.n2730 0.152939
R13691 gnd.n2731 gnd.n2346 0.152939
R13692 gnd.n2737 gnd.n2346 0.152939
R13693 gnd.n2738 gnd.n2737 0.152939
R13694 gnd.n2739 gnd.n2738 0.152939
R13695 gnd.n2740 gnd.n2739 0.152939
R13696 gnd.n2741 gnd.n2740 0.152939
R13697 gnd.n2744 gnd.n2741 0.152939
R13698 gnd.n2745 gnd.n2744 0.152939
R13699 gnd.n2746 gnd.n2745 0.152939
R13700 gnd.n2747 gnd.n2746 0.152939
R13701 gnd.n2750 gnd.n2747 0.152939
R13702 gnd.n2751 gnd.n2750 0.152939
R13703 gnd.n2752 gnd.n2751 0.152939
R13704 gnd.n2753 gnd.n2752 0.152939
R13705 gnd.n2754 gnd.n2753 0.152939
R13706 gnd.n2754 gnd.n2172 0.152939
R13707 gnd.n3205 gnd.n2172 0.152939
R13708 gnd.n3206 gnd.n3205 0.152939
R13709 gnd.n3207 gnd.n3206 0.152939
R13710 gnd.n3207 gnd.n2160 0.152939
R13711 gnd.n3221 gnd.n2160 0.152939
R13712 gnd.n3222 gnd.n3221 0.152939
R13713 gnd.n3223 gnd.n3222 0.152939
R13714 gnd.n3223 gnd.n2147 0.152939
R13715 gnd.n3237 gnd.n2147 0.152939
R13716 gnd.n3238 gnd.n3237 0.152939
R13717 gnd.n3239 gnd.n3238 0.152939
R13718 gnd.n3239 gnd.n2134 0.152939
R13719 gnd.n3253 gnd.n2134 0.152939
R13720 gnd.n3254 gnd.n3253 0.152939
R13721 gnd.n3255 gnd.n3254 0.152939
R13722 gnd.n3255 gnd.n2119 0.152939
R13723 gnd.n3269 gnd.n2119 0.152939
R13724 gnd.n3270 gnd.n3269 0.152939
R13725 gnd.n3271 gnd.n3270 0.152939
R13726 gnd.n3271 gnd.n2107 0.152939
R13727 gnd.n3285 gnd.n2107 0.152939
R13728 gnd.n3286 gnd.n3285 0.152939
R13729 gnd.n3287 gnd.n3286 0.152939
R13730 gnd.n3288 gnd.n3287 0.152939
R13731 gnd.n3288 gnd.n2079 0.152939
R13732 gnd.n3901 gnd.n2079 0.152939
R13733 gnd.n3902 gnd.n3901 0.152939
R13734 gnd.n3903 gnd.n3902 0.152939
R13735 gnd.n3903 gnd.n2064 0.152939
R13736 gnd.n3917 gnd.n2064 0.152939
R13737 gnd.n3918 gnd.n3917 0.152939
R13738 gnd.n3919 gnd.n3918 0.152939
R13739 gnd.n3919 gnd.n2049 0.152939
R13740 gnd.n3933 gnd.n2049 0.152939
R13741 gnd.n3934 gnd.n3933 0.152939
R13742 gnd.n3935 gnd.n3934 0.152939
R13743 gnd.n3935 gnd.n2034 0.152939
R13744 gnd.n3949 gnd.n2034 0.152939
R13745 gnd.n3950 gnd.n3949 0.152939
R13746 gnd.n3951 gnd.n3950 0.152939
R13747 gnd.n3951 gnd.n2020 0.152939
R13748 gnd.n3965 gnd.n2020 0.152939
R13749 gnd.n3966 gnd.n3965 0.152939
R13750 gnd.n3967 gnd.n3966 0.152939
R13751 gnd.n3967 gnd.n2005 0.152939
R13752 gnd.n3981 gnd.n2005 0.152939
R13753 gnd.n3982 gnd.n3981 0.152939
R13754 gnd.n3983 gnd.n3982 0.152939
R13755 gnd.n3983 gnd.n1990 0.152939
R13756 gnd.n3997 gnd.n1990 0.152939
R13757 gnd.n3998 gnd.n3997 0.152939
R13758 gnd.n3999 gnd.n3998 0.152939
R13759 gnd.n3999 gnd.n1975 0.152939
R13760 gnd.n4013 gnd.n1975 0.152939
R13761 gnd.n4014 gnd.n4013 0.152939
R13762 gnd.n4015 gnd.n4014 0.152939
R13763 gnd.n4015 gnd.n1961 0.152939
R13764 gnd.n4029 gnd.n1961 0.152939
R13765 gnd.n4030 gnd.n4029 0.152939
R13766 gnd.n4031 gnd.n4030 0.152939
R13767 gnd.n4031 gnd.n1946 0.152939
R13768 gnd.n4045 gnd.n1946 0.152939
R13769 gnd.n4046 gnd.n4045 0.152939
R13770 gnd.n4047 gnd.n4046 0.152939
R13771 gnd.n4047 gnd.n1933 0.152939
R13772 gnd.n4061 gnd.n1933 0.152939
R13773 gnd.n4062 gnd.n4061 0.152939
R13774 gnd.n4063 gnd.n4062 0.152939
R13775 gnd.n4063 gnd.n1921 0.152939
R13776 gnd.n4077 gnd.n1921 0.152939
R13777 gnd.n4078 gnd.n4077 0.152939
R13778 gnd.n4079 gnd.n4078 0.152939
R13779 gnd.n4079 gnd.n1908 0.152939
R13780 gnd.n4093 gnd.n1908 0.152939
R13781 gnd.n4094 gnd.n4093 0.152939
R13782 gnd.n4095 gnd.n4094 0.152939
R13783 gnd.n4095 gnd.n1894 0.152939
R13784 gnd.n4109 gnd.n1894 0.152939
R13785 gnd.n4110 gnd.n4109 0.152939
R13786 gnd.n4111 gnd.n4110 0.152939
R13787 gnd.n4111 gnd.n1881 0.152939
R13788 gnd.n4125 gnd.n1881 0.152939
R13789 gnd.n4126 gnd.n4125 0.152939
R13790 gnd.n4127 gnd.n4126 0.152939
R13791 gnd.n4127 gnd.n1868 0.152939
R13792 gnd.n4141 gnd.n1868 0.152939
R13793 gnd.n4142 gnd.n4141 0.152939
R13794 gnd.n4143 gnd.n4142 0.152939
R13795 gnd.n4143 gnd.n1855 0.152939
R13796 gnd.n4157 gnd.n1855 0.152939
R13797 gnd.n4158 gnd.n4157 0.152939
R13798 gnd.n4159 gnd.n4158 0.152939
R13799 gnd.n4159 gnd.n1841 0.152939
R13800 gnd.n4173 gnd.n1841 0.152939
R13801 gnd.n4174 gnd.n4173 0.152939
R13802 gnd.n4175 gnd.n4174 0.152939
R13803 gnd.n4175 gnd.n1828 0.152939
R13804 gnd.n4191 gnd.n1828 0.152939
R13805 gnd.n4192 gnd.n4191 0.152939
R13806 gnd.n4193 gnd.n4192 0.152939
R13807 gnd.n4195 gnd.n4193 0.152939
R13808 gnd.n4195 gnd.n4194 0.152939
R13809 gnd.n4194 gnd.n1412 0.152939
R13810 gnd.n1413 gnd.n1412 0.152939
R13811 gnd.n1414 gnd.n1413 0.152939
R13812 gnd.n1636 gnd.n1414 0.152939
R13813 gnd.n1637 gnd.n1636 0.152939
R13814 gnd.n1638 gnd.n1637 0.152939
R13815 gnd.n1638 gnd.n1632 0.152939
R13816 gnd.n4240 gnd.n1632 0.152939
R13817 gnd.n4241 gnd.n4240 0.152939
R13818 gnd.n4242 gnd.n4241 0.152939
R13819 gnd.n4243 gnd.n4242 0.152939
R13820 gnd.n4243 gnd.n1605 0.152939
R13821 gnd.n4271 gnd.n1605 0.152939
R13822 gnd.n4272 gnd.n4271 0.152939
R13823 gnd.n4273 gnd.n4272 0.152939
R13824 gnd.n4274 gnd.n4273 0.152939
R13825 gnd.n4274 gnd.n1577 0.152939
R13826 gnd.n4307 gnd.n1577 0.152939
R13827 gnd.n4308 gnd.n4307 0.152939
R13828 gnd.n4309 gnd.n4308 0.152939
R13829 gnd.n4310 gnd.n4309 0.152939
R13830 gnd.n4310 gnd.n1543 0.152939
R13831 gnd.n4365 gnd.n1543 0.152939
R13832 gnd.n4366 gnd.n4365 0.152939
R13833 gnd.n4367 gnd.n4366 0.152939
R13834 gnd.n4368 gnd.n4367 0.152939
R13835 gnd.n4369 gnd.n4368 0.152939
R13836 gnd.n1163 gnd.n1162 0.152939
R13837 gnd.n1181 gnd.n1163 0.152939
R13838 gnd.n1182 gnd.n1181 0.152939
R13839 gnd.n1183 gnd.n1182 0.152939
R13840 gnd.n1184 gnd.n1183 0.152939
R13841 gnd.n1202 gnd.n1184 0.152939
R13842 gnd.n1203 gnd.n1202 0.152939
R13843 gnd.n1204 gnd.n1203 0.152939
R13844 gnd.n1205 gnd.n1204 0.152939
R13845 gnd.n1223 gnd.n1205 0.152939
R13846 gnd.n1224 gnd.n1223 0.152939
R13847 gnd.n1225 gnd.n1224 0.152939
R13848 gnd.n1226 gnd.n1225 0.152939
R13849 gnd.n1244 gnd.n1226 0.152939
R13850 gnd.n1245 gnd.n1244 0.152939
R13851 gnd.n1246 gnd.n1245 0.152939
R13852 gnd.n1247 gnd.n1246 0.152939
R13853 gnd.n1265 gnd.n1247 0.152939
R13854 gnd.n1266 gnd.n1265 0.152939
R13855 gnd.n1267 gnd.n1266 0.152939
R13856 gnd.n1268 gnd.n1267 0.152939
R13857 gnd.n2289 gnd.n2288 0.152939
R13858 gnd.n2290 gnd.n2289 0.152939
R13859 gnd.n2291 gnd.n2290 0.152939
R13860 gnd.n2292 gnd.n2291 0.152939
R13861 gnd.n2293 gnd.n2292 0.152939
R13862 gnd.n2294 gnd.n2293 0.152939
R13863 gnd.n2295 gnd.n2294 0.152939
R13864 gnd.n2296 gnd.n2295 0.152939
R13865 gnd.n2297 gnd.n2296 0.152939
R13866 gnd.n2298 gnd.n2297 0.152939
R13867 gnd.n2299 gnd.n2298 0.152939
R13868 gnd.n2300 gnd.n2299 0.152939
R13869 gnd.n2301 gnd.n2300 0.152939
R13870 gnd.n2302 gnd.n2301 0.152939
R13871 gnd.n2303 gnd.n2302 0.152939
R13872 gnd.n2878 gnd.n2877 0.152939
R13873 gnd.n2877 gnd.n2308 0.152939
R13874 gnd.n2309 gnd.n2308 0.152939
R13875 gnd.n2310 gnd.n2309 0.152939
R13876 gnd.n2311 gnd.n2310 0.152939
R13877 gnd.n2312 gnd.n2311 0.152939
R13878 gnd.n2313 gnd.n2312 0.152939
R13879 gnd.n2314 gnd.n2313 0.152939
R13880 gnd.n2315 gnd.n2314 0.152939
R13881 gnd.n2316 gnd.n2315 0.152939
R13882 gnd.n2317 gnd.n2316 0.152939
R13883 gnd.n2318 gnd.n2317 0.152939
R13884 gnd.n2319 gnd.n2318 0.152939
R13885 gnd.n2320 gnd.n2319 0.152939
R13886 gnd.n2321 gnd.n2320 0.152939
R13887 gnd.n2322 gnd.n2321 0.152939
R13888 gnd.n2323 gnd.n2322 0.152939
R13889 gnd.n2324 gnd.n2323 0.152939
R13890 gnd.n2837 gnd.n2324 0.152939
R13891 gnd.n2837 gnd.n2836 0.152939
R13892 gnd.n2496 gnd.n2469 0.152939
R13893 gnd.n2554 gnd.n2469 0.152939
R13894 gnd.n2555 gnd.n2554 0.152939
R13895 gnd.n2556 gnd.n2555 0.152939
R13896 gnd.n2556 gnd.n2467 0.152939
R13897 gnd.n2562 gnd.n2467 0.152939
R13898 gnd.n2563 gnd.n2562 0.152939
R13899 gnd.n2564 gnd.n2563 0.152939
R13900 gnd.n2564 gnd.n2465 0.152939
R13901 gnd.n2570 gnd.n2465 0.152939
R13902 gnd.n2571 gnd.n2570 0.152939
R13903 gnd.n2572 gnd.n2571 0.152939
R13904 gnd.n2572 gnd.n2463 0.152939
R13905 gnd.n2578 gnd.n2463 0.152939
R13906 gnd.n2579 gnd.n2578 0.152939
R13907 gnd.n2580 gnd.n2579 0.152939
R13908 gnd.n2580 gnd.n2461 0.152939
R13909 gnd.n2586 gnd.n2461 0.152939
R13910 gnd.n2587 gnd.n2586 0.152939
R13911 gnd.n2589 gnd.n2587 0.152939
R13912 gnd.n2589 gnd.n2588 0.152939
R13913 gnd.n2588 gnd.n2416 0.152939
R13914 gnd.n2417 gnd.n2416 0.152939
R13915 gnd.n2418 gnd.n2417 0.152939
R13916 gnd.n2615 gnd.n2418 0.152939
R13917 gnd.n2616 gnd.n2615 0.152939
R13918 gnd.n2535 gnd.n2476 0.152939
R13919 gnd.n2477 gnd.n2476 0.152939
R13920 gnd.n2478 gnd.n2477 0.152939
R13921 gnd.n2479 gnd.n2478 0.152939
R13922 gnd.n2480 gnd.n2479 0.152939
R13923 gnd.n2481 gnd.n2480 0.152939
R13924 gnd.n2482 gnd.n2481 0.152939
R13925 gnd.n2483 gnd.n2482 0.152939
R13926 gnd.n2484 gnd.n2483 0.152939
R13927 gnd.n2485 gnd.n2484 0.152939
R13928 gnd.n2486 gnd.n2485 0.152939
R13929 gnd.n2487 gnd.n2486 0.152939
R13930 gnd.n2488 gnd.n2487 0.152939
R13931 gnd.n2489 gnd.n2488 0.152939
R13932 gnd.n2490 gnd.n2489 0.152939
R13933 gnd.n2500 gnd.n2490 0.152939
R13934 gnd.n2500 gnd.n2499 0.152939
R13935 gnd.n2499 gnd.n2498 0.152939
R13936 gnd.n2541 gnd.n2536 0.152939
R13937 gnd.n2541 gnd.n2540 0.152939
R13938 gnd.n2540 gnd.n2539 0.152939
R13939 gnd.n2539 gnd.n2537 0.152939
R13940 gnd.n2537 gnd.n1033 0.152939
R13941 gnd.n1034 gnd.n1033 0.152939
R13942 gnd.n1035 gnd.n1034 0.152939
R13943 gnd.n1051 gnd.n1035 0.152939
R13944 gnd.n1052 gnd.n1051 0.152939
R13945 gnd.n1053 gnd.n1052 0.152939
R13946 gnd.n1054 gnd.n1053 0.152939
R13947 gnd.n1072 gnd.n1054 0.152939
R13948 gnd.n1073 gnd.n1072 0.152939
R13949 gnd.n1074 gnd.n1073 0.152939
R13950 gnd.n1075 gnd.n1074 0.152939
R13951 gnd.n1091 gnd.n1075 0.152939
R13952 gnd.n1092 gnd.n1091 0.152939
R13953 gnd.n1093 gnd.n1092 0.152939
R13954 gnd.n1094 gnd.n1093 0.152939
R13955 gnd.n1114 gnd.n1094 0.152939
R13956 gnd.n1115 gnd.n1114 0.152939
R13957 gnd.n1116 gnd.n1115 0.152939
R13958 gnd.n1117 gnd.n1116 0.152939
R13959 gnd.n1132 gnd.n1117 0.152939
R13960 gnd.n1133 gnd.n1132 0.152939
R13961 gnd.n1134 gnd.n1133 0.152939
R13962 gnd.n1151 gnd.n1135 0.152939
R13963 gnd.n1152 gnd.n1151 0.152939
R13964 gnd.n1153 gnd.n1152 0.152939
R13965 gnd.n1154 gnd.n1153 0.152939
R13966 gnd.n1170 gnd.n1154 0.152939
R13967 gnd.n1171 gnd.n1170 0.152939
R13968 gnd.n1172 gnd.n1171 0.152939
R13969 gnd.n1173 gnd.n1172 0.152939
R13970 gnd.n1192 gnd.n1173 0.152939
R13971 gnd.n1193 gnd.n1192 0.152939
R13972 gnd.n1194 gnd.n1193 0.152939
R13973 gnd.n1195 gnd.n1194 0.152939
R13974 gnd.n1212 gnd.n1195 0.152939
R13975 gnd.n1213 gnd.n1212 0.152939
R13976 gnd.n1214 gnd.n1213 0.152939
R13977 gnd.n1215 gnd.n1214 0.152939
R13978 gnd.n1234 gnd.n1215 0.152939
R13979 gnd.n1235 gnd.n1234 0.152939
R13980 gnd.n1236 gnd.n1235 0.152939
R13981 gnd.n1237 gnd.n1236 0.152939
R13982 gnd.n1255 gnd.n1237 0.152939
R13983 gnd.n1256 gnd.n1255 0.152939
R13984 gnd.n1257 gnd.n1256 0.152939
R13985 gnd.n1258 gnd.n1257 0.152939
R13986 gnd.n1275 gnd.n1258 0.152939
R13987 gnd.n4664 gnd.n1275 0.152939
R13988 gnd.n4823 gnd.n1008 0.152939
R13989 gnd.n4823 gnd.n4822 0.152939
R13990 gnd.n4822 gnd.n4821 0.152939
R13991 gnd.n4821 gnd.n1011 0.152939
R13992 gnd.n2429 gnd.n1011 0.152939
R13993 gnd.n2433 gnd.n2429 0.152939
R13994 gnd.n2434 gnd.n2433 0.152939
R13995 gnd.n2435 gnd.n2434 0.152939
R13996 gnd.n2435 gnd.n2427 0.152939
R13997 gnd.n2441 gnd.n2427 0.152939
R13998 gnd.n2442 gnd.n2441 0.152939
R13999 gnd.n2443 gnd.n2442 0.152939
R14000 gnd.n2443 gnd.n2425 0.152939
R14001 gnd.n2449 gnd.n2425 0.152939
R14002 gnd.n2450 gnd.n2449 0.152939
R14003 gnd.n2451 gnd.n2450 0.152939
R14004 gnd.n2451 gnd.n2423 0.152939
R14005 gnd.n2457 gnd.n2423 0.152939
R14006 gnd.n2458 gnd.n2457 0.152939
R14007 gnd.n2459 gnd.n2458 0.152939
R14008 gnd.n2459 gnd.n2421 0.152939
R14009 gnd.n2597 gnd.n2421 0.152939
R14010 gnd.n2598 gnd.n2597 0.152939
R14011 gnd.n2599 gnd.n2598 0.152939
R14012 gnd.n2600 gnd.n2599 0.152939
R14013 gnd.n2601 gnd.n2600 0.152939
R14014 gnd.n2620 gnd.n2619 0.152939
R14015 gnd.n2621 gnd.n2620 0.152939
R14016 gnd.n2622 gnd.n2621 0.152939
R14017 gnd.n2622 gnd.n2373 0.152939
R14018 gnd.n2670 gnd.n2373 0.152939
R14019 gnd.n2671 gnd.n2670 0.152939
R14020 gnd.n2673 gnd.n2671 0.152939
R14021 gnd.n2673 gnd.n2672 0.152939
R14022 gnd.n2672 gnd.n2367 0.152939
R14023 gnd.n2367 gnd.n2365 0.152939
R14024 gnd.n2689 gnd.n2365 0.152939
R14025 gnd.n2690 gnd.n2689 0.152939
R14026 gnd.n2691 gnd.n2690 0.152939
R14027 gnd.n2691 gnd.n2363 0.152939
R14028 gnd.n2700 gnd.n2363 0.152939
R14029 gnd.n2701 gnd.n2700 0.152939
R14030 gnd.n2702 gnd.n2701 0.152939
R14031 gnd.n2703 gnd.n2702 0.152939
R14032 gnd.n2704 gnd.n2703 0.152939
R14033 gnd.n2704 gnd.n2337 0.152939
R14034 gnd.n2787 gnd.n2337 0.152939
R14035 gnd.n2788 gnd.n2787 0.152939
R14036 gnd.n2790 gnd.n2788 0.152939
R14037 gnd.n2790 gnd.n2789 0.152939
R14038 gnd.n2789 gnd.n2329 0.152939
R14039 gnd.n2835 gnd.n2329 0.152939
R14040 gnd.n966 gnd.n965 0.152939
R14041 gnd.n967 gnd.n966 0.152939
R14042 gnd.n968 gnd.n967 0.152939
R14043 gnd.n969 gnd.n968 0.152939
R14044 gnd.n970 gnd.n969 0.152939
R14045 gnd.n971 gnd.n970 0.152939
R14046 gnd.n972 gnd.n971 0.152939
R14047 gnd.n973 gnd.n972 0.152939
R14048 gnd.n974 gnd.n973 0.152939
R14049 gnd.n975 gnd.n974 0.152939
R14050 gnd.n976 gnd.n975 0.152939
R14051 gnd.n977 gnd.n976 0.152939
R14052 gnd.n978 gnd.n977 0.152939
R14053 gnd.n979 gnd.n978 0.152939
R14054 gnd.n980 gnd.n979 0.152939
R14055 gnd.n981 gnd.n980 0.152939
R14056 gnd.n982 gnd.n981 0.152939
R14057 gnd.n985 gnd.n982 0.152939
R14058 gnd.n986 gnd.n985 0.152939
R14059 gnd.n987 gnd.n986 0.152939
R14060 gnd.n988 gnd.n987 0.152939
R14061 gnd.n989 gnd.n988 0.152939
R14062 gnd.n990 gnd.n989 0.152939
R14063 gnd.n991 gnd.n990 0.152939
R14064 gnd.n992 gnd.n991 0.152939
R14065 gnd.n993 gnd.n992 0.152939
R14066 gnd.n994 gnd.n993 0.152939
R14067 gnd.n995 gnd.n994 0.152939
R14068 gnd.n996 gnd.n995 0.152939
R14069 gnd.n997 gnd.n996 0.152939
R14070 gnd.n998 gnd.n997 0.152939
R14071 gnd.n999 gnd.n998 0.152939
R14072 gnd.n1000 gnd.n999 0.152939
R14073 gnd.n1001 gnd.n1000 0.152939
R14074 gnd.n1002 gnd.n1001 0.152939
R14075 gnd.n4831 gnd.n1002 0.152939
R14076 gnd.n4831 gnd.n4830 0.152939
R14077 gnd.n4830 gnd.n4829 0.152939
R14078 gnd.n2547 gnd.n2545 0.152939
R14079 gnd.n2547 gnd.n2546 0.152939
R14080 gnd.n2546 gnd.n1022 0.152939
R14081 gnd.n1023 gnd.n1022 0.152939
R14082 gnd.n1024 gnd.n1023 0.152939
R14083 gnd.n1042 gnd.n1024 0.152939
R14084 gnd.n1043 gnd.n1042 0.152939
R14085 gnd.n1044 gnd.n1043 0.152939
R14086 gnd.n1045 gnd.n1044 0.152939
R14087 gnd.n1061 gnd.n1045 0.152939
R14088 gnd.n1062 gnd.n1061 0.152939
R14089 gnd.n1063 gnd.n1062 0.152939
R14090 gnd.n1064 gnd.n1063 0.152939
R14091 gnd.n1082 gnd.n1064 0.152939
R14092 gnd.n1083 gnd.n1082 0.152939
R14093 gnd.n1084 gnd.n1083 0.152939
R14094 gnd.n1085 gnd.n1084 0.152939
R14095 gnd.n1103 gnd.n1085 0.152939
R14096 gnd.n1104 gnd.n1103 0.152939
R14097 gnd.n1105 gnd.n1104 0.152939
R14098 gnd.n1106 gnd.n1105 0.152939
R14099 gnd.n2409 gnd.n2405 0.152939
R14100 gnd.n2653 gnd.n2405 0.152939
R14101 gnd.n731 gnd.n726 0.152939
R14102 gnd.n732 gnd.n731 0.152939
R14103 gnd.n733 gnd.n732 0.152939
R14104 gnd.n738 gnd.n733 0.152939
R14105 gnd.n739 gnd.n738 0.152939
R14106 gnd.n740 gnd.n739 0.152939
R14107 gnd.n741 gnd.n740 0.152939
R14108 gnd.n746 gnd.n741 0.152939
R14109 gnd.n747 gnd.n746 0.152939
R14110 gnd.n748 gnd.n747 0.152939
R14111 gnd.n749 gnd.n748 0.152939
R14112 gnd.n754 gnd.n749 0.152939
R14113 gnd.n755 gnd.n754 0.152939
R14114 gnd.n756 gnd.n755 0.152939
R14115 gnd.n757 gnd.n756 0.152939
R14116 gnd.n762 gnd.n757 0.152939
R14117 gnd.n763 gnd.n762 0.152939
R14118 gnd.n764 gnd.n763 0.152939
R14119 gnd.n765 gnd.n764 0.152939
R14120 gnd.n770 gnd.n765 0.152939
R14121 gnd.n771 gnd.n770 0.152939
R14122 gnd.n772 gnd.n771 0.152939
R14123 gnd.n773 gnd.n772 0.152939
R14124 gnd.n778 gnd.n773 0.152939
R14125 gnd.n779 gnd.n778 0.152939
R14126 gnd.n780 gnd.n779 0.152939
R14127 gnd.n781 gnd.n780 0.152939
R14128 gnd.n786 gnd.n781 0.152939
R14129 gnd.n787 gnd.n786 0.152939
R14130 gnd.n788 gnd.n787 0.152939
R14131 gnd.n789 gnd.n788 0.152939
R14132 gnd.n794 gnd.n789 0.152939
R14133 gnd.n795 gnd.n794 0.152939
R14134 gnd.n796 gnd.n795 0.152939
R14135 gnd.n797 gnd.n796 0.152939
R14136 gnd.n802 gnd.n797 0.152939
R14137 gnd.n803 gnd.n802 0.152939
R14138 gnd.n804 gnd.n803 0.152939
R14139 gnd.n805 gnd.n804 0.152939
R14140 gnd.n810 gnd.n805 0.152939
R14141 gnd.n811 gnd.n810 0.152939
R14142 gnd.n812 gnd.n811 0.152939
R14143 gnd.n813 gnd.n812 0.152939
R14144 gnd.n818 gnd.n813 0.152939
R14145 gnd.n819 gnd.n818 0.152939
R14146 gnd.n820 gnd.n819 0.152939
R14147 gnd.n821 gnd.n820 0.152939
R14148 gnd.n826 gnd.n821 0.152939
R14149 gnd.n827 gnd.n826 0.152939
R14150 gnd.n828 gnd.n827 0.152939
R14151 gnd.n829 gnd.n828 0.152939
R14152 gnd.n834 gnd.n829 0.152939
R14153 gnd.n835 gnd.n834 0.152939
R14154 gnd.n836 gnd.n835 0.152939
R14155 gnd.n837 gnd.n836 0.152939
R14156 gnd.n842 gnd.n837 0.152939
R14157 gnd.n843 gnd.n842 0.152939
R14158 gnd.n844 gnd.n843 0.152939
R14159 gnd.n845 gnd.n844 0.152939
R14160 gnd.n850 gnd.n845 0.152939
R14161 gnd.n851 gnd.n850 0.152939
R14162 gnd.n852 gnd.n851 0.152939
R14163 gnd.n853 gnd.n852 0.152939
R14164 gnd.n858 gnd.n853 0.152939
R14165 gnd.n859 gnd.n858 0.152939
R14166 gnd.n860 gnd.n859 0.152939
R14167 gnd.n861 gnd.n860 0.152939
R14168 gnd.n866 gnd.n861 0.152939
R14169 gnd.n867 gnd.n866 0.152939
R14170 gnd.n868 gnd.n867 0.152939
R14171 gnd.n869 gnd.n868 0.152939
R14172 gnd.n874 gnd.n869 0.152939
R14173 gnd.n875 gnd.n874 0.152939
R14174 gnd.n876 gnd.n875 0.152939
R14175 gnd.n877 gnd.n876 0.152939
R14176 gnd.n882 gnd.n877 0.152939
R14177 gnd.n883 gnd.n882 0.152939
R14178 gnd.n884 gnd.n883 0.152939
R14179 gnd.n885 gnd.n884 0.152939
R14180 gnd.n890 gnd.n885 0.152939
R14181 gnd.n891 gnd.n890 0.152939
R14182 gnd.n892 gnd.n891 0.152939
R14183 gnd.n893 gnd.n892 0.152939
R14184 gnd.n2408 gnd.n893 0.152939
R14185 gnd.n4227 gnd.n1684 0.152939
R14186 gnd.n4223 gnd.n1684 0.152939
R14187 gnd.n4223 gnd.n4222 0.152939
R14188 gnd.n4222 gnd.n4221 0.152939
R14189 gnd.n4221 gnd.n1812 0.152939
R14190 gnd.n4214 gnd.n1812 0.152939
R14191 gnd.n4214 gnd.n4213 0.152939
R14192 gnd.n4213 gnd.n4212 0.152939
R14193 gnd.n4212 gnd.n4205 0.152939
R14194 gnd.n3199 gnd.n2167 0.152939
R14195 gnd.n3213 gnd.n2167 0.152939
R14196 gnd.n3214 gnd.n3213 0.152939
R14197 gnd.n3215 gnd.n3214 0.152939
R14198 gnd.n3215 gnd.n2154 0.152939
R14199 gnd.n3229 gnd.n2154 0.152939
R14200 gnd.n3230 gnd.n3229 0.152939
R14201 gnd.n3231 gnd.n3230 0.152939
R14202 gnd.n3231 gnd.n2139 0.152939
R14203 gnd.n3245 gnd.n2139 0.152939
R14204 gnd.n3246 gnd.n3245 0.152939
R14205 gnd.n3247 gnd.n3246 0.152939
R14206 gnd.n3247 gnd.n2126 0.152939
R14207 gnd.n3261 gnd.n2126 0.152939
R14208 gnd.n3262 gnd.n3261 0.152939
R14209 gnd.n3263 gnd.n3262 0.152939
R14210 gnd.n3263 gnd.n2113 0.152939
R14211 gnd.n3277 gnd.n2113 0.152939
R14212 gnd.n3278 gnd.n3277 0.152939
R14213 gnd.n3279 gnd.n3278 0.152939
R14214 gnd.n3279 gnd.n2099 0.152939
R14215 gnd.n3295 gnd.n2099 0.152939
R14216 gnd.n3296 gnd.n3295 0.152939
R14217 gnd.n3298 gnd.n3296 0.152939
R14218 gnd.n3298 gnd.n3297 0.152939
R14219 gnd.n3297 gnd.n2071 0.152939
R14220 gnd.n3909 gnd.n2071 0.152939
R14221 gnd.n3910 gnd.n3909 0.152939
R14222 gnd.n3911 gnd.n3910 0.152939
R14223 gnd.n3911 gnd.n2056 0.152939
R14224 gnd.n3925 gnd.n2056 0.152939
R14225 gnd.n3926 gnd.n3925 0.152939
R14226 gnd.n3927 gnd.n3926 0.152939
R14227 gnd.n3927 gnd.n2041 0.152939
R14228 gnd.n3941 gnd.n2041 0.152939
R14229 gnd.n3942 gnd.n3941 0.152939
R14230 gnd.n3943 gnd.n3942 0.152939
R14231 gnd.n3943 gnd.n2027 0.152939
R14232 gnd.n3957 gnd.n2027 0.152939
R14233 gnd.n3958 gnd.n3957 0.152939
R14234 gnd.n3959 gnd.n3958 0.152939
R14235 gnd.n3959 gnd.n2012 0.152939
R14236 gnd.n3973 gnd.n2012 0.152939
R14237 gnd.n3974 gnd.n3973 0.152939
R14238 gnd.n3975 gnd.n3974 0.152939
R14239 gnd.n3975 gnd.n1997 0.152939
R14240 gnd.n3989 gnd.n1997 0.152939
R14241 gnd.n3990 gnd.n3989 0.152939
R14242 gnd.n3991 gnd.n3990 0.152939
R14243 gnd.n3991 gnd.n1982 0.152939
R14244 gnd.n4005 gnd.n1982 0.152939
R14245 gnd.n4006 gnd.n4005 0.152939
R14246 gnd.n4007 gnd.n4006 0.152939
R14247 gnd.n4007 gnd.n1967 0.152939
R14248 gnd.n4021 gnd.n1967 0.152939
R14249 gnd.n4022 gnd.n4021 0.152939
R14250 gnd.n4023 gnd.n4022 0.152939
R14251 gnd.n4023 gnd.n1952 0.152939
R14252 gnd.n4037 gnd.n1952 0.152939
R14253 gnd.n4038 gnd.n4037 0.152939
R14254 gnd.n4039 gnd.n4038 0.152939
R14255 gnd.n4039 gnd.n1939 0.152939
R14256 gnd.n4053 gnd.n1939 0.152939
R14257 gnd.n4054 gnd.n4053 0.152939
R14258 gnd.n4055 gnd.n4054 0.152939
R14259 gnd.n4055 gnd.n1927 0.152939
R14260 gnd.n4069 gnd.n1927 0.152939
R14261 gnd.n4070 gnd.n4069 0.152939
R14262 gnd.n4071 gnd.n4070 0.152939
R14263 gnd.n4071 gnd.n1914 0.152939
R14264 gnd.n4085 gnd.n1914 0.152939
R14265 gnd.n4086 gnd.n4085 0.152939
R14266 gnd.n4087 gnd.n4086 0.152939
R14267 gnd.n4087 gnd.n1901 0.152939
R14268 gnd.n4101 gnd.n1901 0.152939
R14269 gnd.n4102 gnd.n4101 0.152939
R14270 gnd.n4103 gnd.n4102 0.152939
R14271 gnd.n4103 gnd.n1887 0.152939
R14272 gnd.n4117 gnd.n1887 0.152939
R14273 gnd.n4118 gnd.n4117 0.152939
R14274 gnd.n4119 gnd.n4118 0.152939
R14275 gnd.n4119 gnd.n1873 0.152939
R14276 gnd.n4133 gnd.n1873 0.152939
R14277 gnd.n4134 gnd.n4133 0.152939
R14278 gnd.n4135 gnd.n4134 0.152939
R14279 gnd.n4135 gnd.n1861 0.152939
R14280 gnd.n4149 gnd.n1861 0.152939
R14281 gnd.n4150 gnd.n4149 0.152939
R14282 gnd.n4151 gnd.n4150 0.152939
R14283 gnd.n4151 gnd.n1848 0.152939
R14284 gnd.n4165 gnd.n1848 0.152939
R14285 gnd.n4166 gnd.n4165 0.152939
R14286 gnd.n4167 gnd.n4166 0.152939
R14287 gnd.n4167 gnd.n1835 0.152939
R14288 gnd.n4181 gnd.n1835 0.152939
R14289 gnd.n4182 gnd.n4181 0.152939
R14290 gnd.n4185 gnd.n4182 0.152939
R14291 gnd.n4185 gnd.n4184 0.152939
R14292 gnd.n4184 gnd.n4183 0.152939
R14293 gnd.n4183 gnd.n1820 0.152939
R14294 gnd.n4204 gnd.n1820 0.152939
R14295 gnd.n2821 gnd.n2798 0.152939
R14296 gnd.n2821 gnd.n2820 0.152939
R14297 gnd.n2820 gnd.n2819 0.152939
R14298 gnd.n2819 gnd.n2804 0.152939
R14299 gnd.n2815 gnd.n2804 0.152939
R14300 gnd.n2815 gnd.n2814 0.152939
R14301 gnd.n2814 gnd.n2811 0.152939
R14302 gnd.n2811 gnd.n2178 0.152939
R14303 gnd.n3198 gnd.n2178 0.152939
R14304 gnd.n2632 gnd.n2631 0.152939
R14305 gnd.n2631 gnd.n2376 0.152939
R14306 gnd.n2662 gnd.n2376 0.152939
R14307 gnd.n2663 gnd.n2662 0.152939
R14308 gnd.n2664 gnd.n2663 0.152939
R14309 gnd.n2664 gnd.n2369 0.152939
R14310 gnd.n2679 gnd.n2369 0.152939
R14311 gnd.n2680 gnd.n2679 0.152939
R14312 gnd.n2681 gnd.n2680 0.152939
R14313 gnd.n2681 gnd.n2357 0.152939
R14314 gnd.n2720 gnd.n2357 0.152939
R14315 gnd.n2720 gnd.n2719 0.152939
R14316 gnd.n2719 gnd.n2718 0.152939
R14317 gnd.n2718 gnd.n2358 0.152939
R14318 gnd.n2714 gnd.n2358 0.152939
R14319 gnd.n2714 gnd.n2713 0.152939
R14320 gnd.n2713 gnd.n2712 0.152939
R14321 gnd.n2712 gnd.n2340 0.152939
R14322 gnd.n2779 gnd.n2340 0.152939
R14323 gnd.n2780 gnd.n2779 0.152939
R14324 gnd.n2781 gnd.n2780 0.152939
R14325 gnd.n2781 gnd.n2334 0.152939
R14326 gnd.n2796 gnd.n2334 0.152939
R14327 gnd.n2797 gnd.n2796 0.152939
R14328 gnd.n2828 gnd.n2797 0.152939
R14329 gnd.n2828 gnd.n2827 0.152939
R14330 gnd.n4661 gnd.n1278 0.152939
R14331 gnd.n4657 gnd.n1278 0.152939
R14332 gnd.n4657 gnd.n4656 0.152939
R14333 gnd.n4656 gnd.n4655 0.152939
R14334 gnd.n4655 gnd.n1283 0.152939
R14335 gnd.n4651 gnd.n1283 0.152939
R14336 gnd.n4651 gnd.n4650 0.152939
R14337 gnd.n4650 gnd.n4649 0.152939
R14338 gnd.n4649 gnd.n1288 0.152939
R14339 gnd.n4645 gnd.n1288 0.152939
R14340 gnd.n4645 gnd.n4644 0.152939
R14341 gnd.n4644 gnd.n4643 0.152939
R14342 gnd.n4643 gnd.n1293 0.152939
R14343 gnd.n4639 gnd.n1293 0.152939
R14344 gnd.n4639 gnd.n4638 0.152939
R14345 gnd.n4638 gnd.n4637 0.152939
R14346 gnd.n4637 gnd.n1298 0.152939
R14347 gnd.n4633 gnd.n1298 0.152939
R14348 gnd.n4633 gnd.n4632 0.152939
R14349 gnd.n4632 gnd.n4631 0.152939
R14350 gnd.n4631 gnd.n1303 0.152939
R14351 gnd.n4627 gnd.n1303 0.152939
R14352 gnd.n4627 gnd.n4626 0.152939
R14353 gnd.n4626 gnd.n4625 0.152939
R14354 gnd.n4625 gnd.n1308 0.152939
R14355 gnd.n4621 gnd.n1308 0.152939
R14356 gnd.n4621 gnd.n4620 0.152939
R14357 gnd.n4620 gnd.n4619 0.152939
R14358 gnd.n4619 gnd.n1313 0.152939
R14359 gnd.n4615 gnd.n1313 0.152939
R14360 gnd.n4615 gnd.n4614 0.152939
R14361 gnd.n4614 gnd.n4613 0.152939
R14362 gnd.n4613 gnd.n1318 0.152939
R14363 gnd.n4609 gnd.n1318 0.152939
R14364 gnd.n4609 gnd.n4608 0.152939
R14365 gnd.n4608 gnd.n4607 0.152939
R14366 gnd.n4607 gnd.n1323 0.152939
R14367 gnd.n4603 gnd.n1323 0.152939
R14368 gnd.n4603 gnd.n4602 0.152939
R14369 gnd.n4602 gnd.n4601 0.152939
R14370 gnd.n4601 gnd.n1328 0.152939
R14371 gnd.n4597 gnd.n1328 0.152939
R14372 gnd.n4597 gnd.n4596 0.152939
R14373 gnd.n4596 gnd.n4595 0.152939
R14374 gnd.n4595 gnd.n1333 0.152939
R14375 gnd.n4591 gnd.n1333 0.152939
R14376 gnd.n4591 gnd.n4590 0.152939
R14377 gnd.n4590 gnd.n4589 0.152939
R14378 gnd.n4589 gnd.n1338 0.152939
R14379 gnd.n4585 gnd.n1338 0.152939
R14380 gnd.n4585 gnd.n4584 0.152939
R14381 gnd.n4584 gnd.n4583 0.152939
R14382 gnd.n4583 gnd.n1343 0.152939
R14383 gnd.n4579 gnd.n1343 0.152939
R14384 gnd.n4579 gnd.n4578 0.152939
R14385 gnd.n4578 gnd.n4577 0.152939
R14386 gnd.n4577 gnd.n1348 0.152939
R14387 gnd.n4573 gnd.n1348 0.152939
R14388 gnd.n4573 gnd.n4572 0.152939
R14389 gnd.n4572 gnd.n4571 0.152939
R14390 gnd.n4571 gnd.n1353 0.152939
R14391 gnd.n4567 gnd.n1353 0.152939
R14392 gnd.n4567 gnd.n4566 0.152939
R14393 gnd.n4566 gnd.n4565 0.152939
R14394 gnd.n4565 gnd.n1358 0.152939
R14395 gnd.n4561 gnd.n1358 0.152939
R14396 gnd.n4561 gnd.n4560 0.152939
R14397 gnd.n4560 gnd.n4559 0.152939
R14398 gnd.n4559 gnd.n1363 0.152939
R14399 gnd.n4555 gnd.n1363 0.152939
R14400 gnd.n4555 gnd.n4554 0.152939
R14401 gnd.n4554 gnd.n4553 0.152939
R14402 gnd.n4553 gnd.n1368 0.152939
R14403 gnd.n4549 gnd.n1368 0.152939
R14404 gnd.n4549 gnd.n4548 0.152939
R14405 gnd.n4548 gnd.n4547 0.152939
R14406 gnd.n4547 gnd.n1373 0.152939
R14407 gnd.n4543 gnd.n1373 0.152939
R14408 gnd.n4543 gnd.n4542 0.152939
R14409 gnd.n4542 gnd.n4541 0.152939
R14410 gnd.n4541 gnd.n1378 0.152939
R14411 gnd.n4537 gnd.n1378 0.152939
R14412 gnd.n4537 gnd.n4536 0.152939
R14413 gnd.n4536 gnd.n4535 0.152939
R14414 gnd.n4535 gnd.n1383 0.152939
R14415 gnd.n4531 gnd.n1383 0.152939
R14416 gnd.n4531 gnd.n4530 0.152939
R14417 gnd.n4530 gnd.n4529 0.152939
R14418 gnd.n4529 gnd.n1388 0.152939
R14419 gnd.n4525 gnd.n1388 0.152939
R14420 gnd.n4525 gnd.n4524 0.152939
R14421 gnd.n4524 gnd.n4523 0.152939
R14422 gnd.n4523 gnd.n1393 0.152939
R14423 gnd.n4519 gnd.n1393 0.152939
R14424 gnd.n4519 gnd.n4518 0.152939
R14425 gnd.n4518 gnd.n4517 0.152939
R14426 gnd.n4517 gnd.n1398 0.152939
R14427 gnd.n4513 gnd.n1398 0.152939
R14428 gnd.n4513 gnd.n4512 0.152939
R14429 gnd.n4512 gnd.n4511 0.152939
R14430 gnd.n4511 gnd.n1403 0.152939
R14431 gnd.n4419 gnd.n4418 0.152939
R14432 gnd.n4418 gnd.n4417 0.152939
R14433 gnd.n4417 gnd.n1504 0.152939
R14434 gnd.n4413 gnd.n1504 0.152939
R14435 gnd.n4413 gnd.n4412 0.152939
R14436 gnd.n4412 gnd.n4411 0.152939
R14437 gnd.n4411 gnd.n1509 0.152939
R14438 gnd.n4407 gnd.n1509 0.152939
R14439 gnd.n4407 gnd.n4406 0.152939
R14440 gnd.n4406 gnd.n4405 0.152939
R14441 gnd.n4405 gnd.n1514 0.152939
R14442 gnd.n4401 gnd.n1514 0.152939
R14443 gnd.n4401 gnd.n4400 0.152939
R14444 gnd.n4400 gnd.n4399 0.152939
R14445 gnd.n4399 gnd.n1519 0.152939
R14446 gnd.n4395 gnd.n1519 0.152939
R14447 gnd.n4395 gnd.n4394 0.152939
R14448 gnd.n4394 gnd.n4393 0.152939
R14449 gnd.n4393 gnd.n1524 0.152939
R14450 gnd.n4389 gnd.n1524 0.152939
R14451 gnd.n4389 gnd.n285 0.152939
R14452 gnd.n7289 gnd.n285 0.152939
R14453 gnd.n7289 gnd.n7288 0.152939
R14454 gnd.n7288 gnd.n7287 0.152939
R14455 gnd.n7287 gnd.n286 0.152939
R14456 gnd.n7283 gnd.n286 0.152939
R14457 gnd.n7281 gnd.n7280 0.152939
R14458 gnd.n7280 gnd.n292 0.152939
R14459 gnd.n292 gnd.n260 0.152939
R14460 gnd.n7302 gnd.n260 0.152939
R14461 gnd.n7303 gnd.n7302 0.152939
R14462 gnd.n7304 gnd.n7303 0.152939
R14463 gnd.n7304 gnd.n244 0.152939
R14464 gnd.n7318 gnd.n244 0.152939
R14465 gnd.n7319 gnd.n7318 0.152939
R14466 gnd.n7320 gnd.n7319 0.152939
R14467 gnd.n7320 gnd.n229 0.152939
R14468 gnd.n7334 gnd.n229 0.152939
R14469 gnd.n7335 gnd.n7334 0.152939
R14470 gnd.n7336 gnd.n7335 0.152939
R14471 gnd.n7336 gnd.n214 0.152939
R14472 gnd.n7350 gnd.n214 0.152939
R14473 gnd.n7351 gnd.n7350 0.152939
R14474 gnd.n7352 gnd.n7351 0.152939
R14475 gnd.n7352 gnd.n199 0.152939
R14476 gnd.n7366 gnd.n199 0.152939
R14477 gnd.n7367 gnd.n7366 0.152939
R14478 gnd.n7443 gnd.n7367 0.152939
R14479 gnd.n7443 gnd.n7442 0.152939
R14480 gnd.n7442 gnd.n7441 0.152939
R14481 gnd.n7441 gnd.n7368 0.152939
R14482 gnd.n7437 gnd.n7368 0.152939
R14483 gnd.n7436 gnd.n7370 0.152939
R14484 gnd.n7432 gnd.n7370 0.152939
R14485 gnd.n7432 gnd.n7431 0.152939
R14486 gnd.n7431 gnd.n7430 0.152939
R14487 gnd.n7430 gnd.n7376 0.152939
R14488 gnd.n7426 gnd.n7376 0.152939
R14489 gnd.n7426 gnd.n7425 0.152939
R14490 gnd.n7425 gnd.n7424 0.152939
R14491 gnd.n7424 gnd.n7384 0.152939
R14492 gnd.n7420 gnd.n7384 0.152939
R14493 gnd.n7420 gnd.n7419 0.152939
R14494 gnd.n7419 gnd.n7418 0.152939
R14495 gnd.n7418 gnd.n7392 0.152939
R14496 gnd.n7414 gnd.n7392 0.152939
R14497 gnd.n7414 gnd.n7413 0.152939
R14498 gnd.n7413 gnd.n7412 0.152939
R14499 gnd.n7412 gnd.n7400 0.152939
R14500 gnd.n7408 gnd.n7400 0.152939
R14501 gnd.n4231 gnd.n4230 0.152939
R14502 gnd.n4233 gnd.n4231 0.152939
R14503 gnd.n4233 gnd.n4232 0.152939
R14504 gnd.n4232 gnd.n1612 0.152939
R14505 gnd.n4261 gnd.n1612 0.152939
R14506 gnd.n4262 gnd.n4261 0.152939
R14507 gnd.n4264 gnd.n4262 0.152939
R14508 gnd.n4264 gnd.n4263 0.152939
R14509 gnd.n4263 gnd.n1585 0.152939
R14510 gnd.n4292 gnd.n1585 0.152939
R14511 gnd.n4293 gnd.n4292 0.152939
R14512 gnd.n4300 gnd.n4293 0.152939
R14513 gnd.n4300 gnd.n4299 0.152939
R14514 gnd.n4299 gnd.n4298 0.152939
R14515 gnd.n4298 gnd.n4294 0.152939
R14516 gnd.n4294 gnd.n1551 0.152939
R14517 gnd.n4357 gnd.n1551 0.152939
R14518 gnd.n4357 gnd.n4356 0.152939
R14519 gnd.n4356 gnd.n4355 0.152939
R14520 gnd.n4355 gnd.n1552 0.152939
R14521 gnd.n4351 gnd.n1552 0.152939
R14522 gnd.n4351 gnd.n310 0.152939
R14523 gnd.n7195 gnd.n310 0.152939
R14524 gnd.n7196 gnd.n7195 0.152939
R14525 gnd.n7197 gnd.n7196 0.152939
R14526 gnd.n7197 gnd.n67 0.152939
R14527 gnd.n7575 gnd.n68 0.152939
R14528 gnd.n7571 gnd.n68 0.152939
R14529 gnd.n7571 gnd.n7570 0.152939
R14530 gnd.n7570 gnd.n7569 0.152939
R14531 gnd.n7569 gnd.n74 0.152939
R14532 gnd.n7565 gnd.n74 0.152939
R14533 gnd.n7565 gnd.n7564 0.152939
R14534 gnd.n7564 gnd.n7563 0.152939
R14535 gnd.n7563 gnd.n79 0.152939
R14536 gnd.n7559 gnd.n79 0.152939
R14537 gnd.n7559 gnd.n7558 0.152939
R14538 gnd.n7558 gnd.n7557 0.152939
R14539 gnd.n7557 gnd.n84 0.152939
R14540 gnd.n7553 gnd.n84 0.152939
R14541 gnd.n7553 gnd.n7552 0.152939
R14542 gnd.n7552 gnd.n7551 0.152939
R14543 gnd.n7551 gnd.n89 0.152939
R14544 gnd.n7547 gnd.n89 0.152939
R14545 gnd.n7547 gnd.n7546 0.152939
R14546 gnd.n7546 gnd.n7545 0.152939
R14547 gnd.n7545 gnd.n94 0.152939
R14548 gnd.n7541 gnd.n94 0.152939
R14549 gnd.n7541 gnd.n7540 0.152939
R14550 gnd.n7540 gnd.n7539 0.152939
R14551 gnd.n7539 gnd.n99 0.152939
R14552 gnd.n102 gnd.n99 0.152939
R14553 gnd.n4228 gnd.n4227 0.151415
R14554 gnd.n2826 gnd.n2798 0.151415
R14555 gnd.n2654 gnd.n2400 0.140744
R14556 gnd.n4369 gnd.n269 0.140744
R14557 gnd.n5535 gnd.n5092 0.0767195
R14558 gnd.n5535 gnd.n5471 0.0767195
R14559 gnd.n7296 gnd.n253 0.0767195
R14560 gnd.n300 gnd.n291 0.0767195
R14561 gnd.n7209 gnd.n291 0.0767195
R14562 gnd.n7296 gnd.n268 0.0767195
R14563 gnd.n1162 gnd.n1125 0.0767195
R14564 gnd.n2617 gnd.n1134 0.0767195
R14565 gnd.n2617 gnd.n1135 0.0767195
R14566 gnd.n2618 gnd.n2601 0.0767195
R14567 gnd.n2619 gnd.n2618 0.0767195
R14568 gnd.n1125 gnd.n1106 0.0767195
R14569 gnd.n7283 gnd.n7282 0.0767195
R14570 gnd.n7282 gnd.n7281 0.0767195
R14571 gnd.n7576 gnd.n67 0.0767195
R14572 gnd.n7576 gnd.n7575 0.0767195
R14573 gnd.n2630 gnd.n2616 0.0695946
R14574 gnd.n2632 gnd.n2630 0.0695946
R14575 gnd.n4663 gnd.n4662 0.063
R14576 gnd.n1723 gnd.n1503 0.063
R14577 gnd.n6274 gnd.n4941 0.0477147
R14578 gnd.n5426 gnd.n5314 0.0442063
R14579 gnd.n5427 gnd.n5426 0.0442063
R14580 gnd.n5428 gnd.n5427 0.0442063
R14581 gnd.n5428 gnd.n5303 0.0442063
R14582 gnd.n5442 gnd.n5303 0.0442063
R14583 gnd.n5443 gnd.n5442 0.0442063
R14584 gnd.n5444 gnd.n5443 0.0442063
R14585 gnd.n5444 gnd.n5290 0.0442063
R14586 gnd.n5574 gnd.n5290 0.0442063
R14587 gnd.n5575 gnd.n5574 0.0442063
R14588 gnd.n5577 gnd.n5224 0.0344674
R14589 gnd.n1802 gnd.n1683 0.0343753
R14590 gnd.n2825 gnd.n2247 0.0343753
R14591 gnd.n5597 gnd.n5596 0.0269946
R14592 gnd.n5599 gnd.n5598 0.0269946
R14593 gnd.n5219 gnd.n5217 0.0269946
R14594 gnd.n5609 gnd.n5607 0.0269946
R14595 gnd.n5608 gnd.n5198 0.0269946
R14596 gnd.n5628 gnd.n5627 0.0269946
R14597 gnd.n5630 gnd.n5629 0.0269946
R14598 gnd.n5193 gnd.n5191 0.0269946
R14599 gnd.n5640 gnd.n5638 0.0269946
R14600 gnd.n5639 gnd.n5174 0.0269946
R14601 gnd.n5659 gnd.n5658 0.0269946
R14602 gnd.n5661 gnd.n5660 0.0269946
R14603 gnd.n5168 gnd.n5166 0.0269946
R14604 gnd.n5671 gnd.n5669 0.0269946
R14605 gnd.n5670 gnd.n5148 0.0269946
R14606 gnd.n5690 gnd.n5689 0.0269946
R14607 gnd.n5692 gnd.n5691 0.0269946
R14608 gnd.n5142 gnd.n5140 0.0269946
R14609 gnd.n5702 gnd.n5700 0.0269946
R14610 gnd.n5701 gnd.n5123 0.0269946
R14611 gnd.n5721 gnd.n5720 0.0269946
R14612 gnd.n5723 gnd.n5722 0.0269946
R14613 gnd.n5117 gnd.n5115 0.0269946
R14614 gnd.n5733 gnd.n5731 0.0269946
R14615 gnd.n5732 gnd.n5099 0.0269946
R14616 gnd.n5751 gnd.n5750 0.0269946
R14617 gnd.n5753 gnd.n5752 0.0269946
R14618 gnd.n5087 gnd.n5086 0.0269946
R14619 gnd.n5787 gnd.n5083 0.0269946
R14620 gnd.n5786 gnd.n5084 0.0269946
R14621 gnd.n5806 gnd.n5066 0.0269946
R14622 gnd.n5808 gnd.n5807 0.0269946
R14623 gnd.n5809 gnd.n5064 0.0269946
R14624 gnd.n5816 gnd.n5812 0.0269946
R14625 gnd.n5815 gnd.n5814 0.0269946
R14626 gnd.n5813 gnd.n5043 0.0269946
R14627 gnd.n5840 gnd.n5044 0.0269946
R14628 gnd.n5839 gnd.n5045 0.0269946
R14629 gnd.n5881 gnd.n5022 0.0269946
R14630 gnd.n5883 gnd.n5882 0.0269946
R14631 gnd.n5892 gnd.n5015 0.0269946
R14632 gnd.n5894 gnd.n5893 0.0269946
R14633 gnd.n5895 gnd.n5011 0.0269946
R14634 gnd.n6183 gnd.n5012 0.0269946
R14635 gnd.n6182 gnd.n5013 0.0269946
R14636 gnd.n5899 gnd.n902 0.0269946
R14637 gnd.n5900 gnd.n903 0.0269946
R14638 gnd.n5902 gnd.n904 0.0269946
R14639 gnd.n6162 gnd.n6161 0.0269946
R14640 gnd.n6163 gnd.n926 0.0269946
R14641 gnd.n6164 gnd.n927 0.0269946
R14642 gnd.n6165 gnd.n928 0.0269946
R14643 gnd.n1725 gnd.n1723 0.0245515
R14644 gnd.n4662 gnd.n1277 0.0245515
R14645 gnd.n5577 gnd.n5576 0.0202011
R14646 gnd.n1725 gnd.n1724 0.0174377
R14647 gnd.n1724 gnd.n1720 0.0174377
R14648 gnd.n1734 gnd.n1720 0.0174377
R14649 gnd.n1734 gnd.n1733 0.0174377
R14650 gnd.n1733 gnd.n1721 0.0174377
R14651 gnd.n1721 gnd.n1716 0.0174377
R14652 gnd.n1742 gnd.n1716 0.0174377
R14653 gnd.n1744 gnd.n1742 0.0174377
R14654 gnd.n1744 gnd.n1743 0.0174377
R14655 gnd.n1743 gnd.n1713 0.0174377
R14656 gnd.n1753 gnd.n1713 0.0174377
R14657 gnd.n1753 gnd.n1752 0.0174377
R14658 gnd.n1752 gnd.n1714 0.0174377
R14659 gnd.n1714 gnd.n1709 0.0174377
R14660 gnd.n1761 gnd.n1709 0.0174377
R14661 gnd.n1763 gnd.n1761 0.0174377
R14662 gnd.n1763 gnd.n1762 0.0174377
R14663 gnd.n1762 gnd.n1706 0.0174377
R14664 gnd.n1772 gnd.n1706 0.0174377
R14665 gnd.n1772 gnd.n1771 0.0174377
R14666 gnd.n1771 gnd.n1707 0.0174377
R14667 gnd.n1707 gnd.n1702 0.0174377
R14668 gnd.n1780 gnd.n1702 0.0174377
R14669 gnd.n1781 gnd.n1780 0.0174377
R14670 gnd.n1781 gnd.n1700 0.0174377
R14671 gnd.n1786 gnd.n1700 0.0174377
R14672 gnd.n1788 gnd.n1786 0.0174377
R14673 gnd.n1788 gnd.n1787 0.0174377
R14674 gnd.n1787 gnd.n1696 0.0174377
R14675 gnd.n1797 gnd.n1696 0.0174377
R14676 gnd.n1797 gnd.n1796 0.0174377
R14677 gnd.n1796 gnd.n1689 0.0174377
R14678 gnd.n1689 gnd.n1688 0.0174377
R14679 gnd.n1801 gnd.n1688 0.0174377
R14680 gnd.n1802 gnd.n1801 0.0174377
R14681 gnd.n2196 gnd.n1277 0.0174377
R14682 gnd.n2198 gnd.n2196 0.0174377
R14683 gnd.n3188 gnd.n2198 0.0174377
R14684 gnd.n3188 gnd.n3187 0.0174377
R14685 gnd.n3187 gnd.n2199 0.0174377
R14686 gnd.n3184 gnd.n2199 0.0174377
R14687 gnd.n3184 gnd.n3183 0.0174377
R14688 gnd.n3183 gnd.n2204 0.0174377
R14689 gnd.n3180 gnd.n2204 0.0174377
R14690 gnd.n3180 gnd.n3179 0.0174377
R14691 gnd.n3179 gnd.n2209 0.0174377
R14692 gnd.n3176 gnd.n2209 0.0174377
R14693 gnd.n3176 gnd.n3175 0.0174377
R14694 gnd.n3175 gnd.n2213 0.0174377
R14695 gnd.n3172 gnd.n2213 0.0174377
R14696 gnd.n3172 gnd.n3171 0.0174377
R14697 gnd.n3171 gnd.n2217 0.0174377
R14698 gnd.n3168 gnd.n2217 0.0174377
R14699 gnd.n3168 gnd.n3167 0.0174377
R14700 gnd.n3167 gnd.n2221 0.0174377
R14701 gnd.n3164 gnd.n2221 0.0174377
R14702 gnd.n3164 gnd.n3163 0.0174377
R14703 gnd.n3163 gnd.n2227 0.0174377
R14704 gnd.n3160 gnd.n2227 0.0174377
R14705 gnd.n3160 gnd.n3159 0.0174377
R14706 gnd.n3159 gnd.n2231 0.0174377
R14707 gnd.n3156 gnd.n2231 0.0174377
R14708 gnd.n3156 gnd.n3155 0.0174377
R14709 gnd.n3155 gnd.n2235 0.0174377
R14710 gnd.n3152 gnd.n2235 0.0174377
R14711 gnd.n3152 gnd.n3151 0.0174377
R14712 gnd.n3151 gnd.n2241 0.0174377
R14713 gnd.n3148 gnd.n2241 0.0174377
R14714 gnd.n3148 gnd.n3147 0.0174377
R14715 gnd.n3147 gnd.n2247 0.0174377
R14716 gnd.n5576 gnd.n5575 0.0148637
R14717 gnd.n6159 gnd.n5903 0.0144266
R14718 gnd.n6160 gnd.n6159 0.0130679
R14719 gnd.n326 gnd.n269 0.0126951
R14720 gnd.n2654 gnd.n2653 0.0126951
R14721 gnd.n5596 gnd.n5224 0.00797283
R14722 gnd.n5598 gnd.n5597 0.00797283
R14723 gnd.n5599 gnd.n5219 0.00797283
R14724 gnd.n5607 gnd.n5217 0.00797283
R14725 gnd.n5609 gnd.n5608 0.00797283
R14726 gnd.n5627 gnd.n5198 0.00797283
R14727 gnd.n5629 gnd.n5628 0.00797283
R14728 gnd.n5630 gnd.n5193 0.00797283
R14729 gnd.n5638 gnd.n5191 0.00797283
R14730 gnd.n5640 gnd.n5639 0.00797283
R14731 gnd.n5658 gnd.n5174 0.00797283
R14732 gnd.n5660 gnd.n5659 0.00797283
R14733 gnd.n5661 gnd.n5168 0.00797283
R14734 gnd.n5669 gnd.n5166 0.00797283
R14735 gnd.n5671 gnd.n5670 0.00797283
R14736 gnd.n5689 gnd.n5148 0.00797283
R14737 gnd.n5691 gnd.n5690 0.00797283
R14738 gnd.n5692 gnd.n5142 0.00797283
R14739 gnd.n5700 gnd.n5140 0.00797283
R14740 gnd.n5702 gnd.n5701 0.00797283
R14741 gnd.n5720 gnd.n5123 0.00797283
R14742 gnd.n5722 gnd.n5721 0.00797283
R14743 gnd.n5723 gnd.n5117 0.00797283
R14744 gnd.n5731 gnd.n5115 0.00797283
R14745 gnd.n5733 gnd.n5732 0.00797283
R14746 gnd.n5750 gnd.n5099 0.00797283
R14747 gnd.n5752 gnd.n5751 0.00797283
R14748 gnd.n5753 gnd.n5087 0.00797283
R14749 gnd.n5086 gnd.n5083 0.00797283
R14750 gnd.n5787 gnd.n5786 0.00797283
R14751 gnd.n5084 gnd.n5066 0.00797283
R14752 gnd.n5807 gnd.n5806 0.00797283
R14753 gnd.n5809 gnd.n5808 0.00797283
R14754 gnd.n5812 gnd.n5064 0.00797283
R14755 gnd.n5816 gnd.n5815 0.00797283
R14756 gnd.n5814 gnd.n5813 0.00797283
R14757 gnd.n5044 gnd.n5043 0.00797283
R14758 gnd.n5840 gnd.n5839 0.00797283
R14759 gnd.n5045 gnd.n5022 0.00797283
R14760 gnd.n5883 gnd.n5881 0.00797283
R14761 gnd.n5882 gnd.n5015 0.00797283
R14762 gnd.n5893 gnd.n5892 0.00797283
R14763 gnd.n5895 gnd.n5894 0.00797283
R14764 gnd.n5012 gnd.n5011 0.00797283
R14765 gnd.n6183 gnd.n6182 0.00797283
R14766 gnd.n5899 gnd.n5013 0.00797283
R14767 gnd.n5900 gnd.n902 0.00797283
R14768 gnd.n5902 gnd.n903 0.00797283
R14769 gnd.n5903 gnd.n904 0.00797283
R14770 gnd.n6161 gnd.n6160 0.00797283
R14771 gnd.n6163 gnd.n6162 0.00797283
R14772 gnd.n6164 gnd.n926 0.00797283
R14773 gnd.n6165 gnd.n927 0.00797283
R14774 gnd.n4941 gnd.n928 0.00797283
R14775 gnd.n7282 gnd.n291 0.00507153
R14776 gnd.n2618 gnd.n2617 0.00507153
R14777 gnd.n4228 gnd.n1683 0.000838753
R14778 gnd.n2826 gnd.n2825 0.000838753
R14779 vdd.n327 vdd.n291 756.745
R14780 vdd.n268 vdd.n232 756.745
R14781 vdd.n225 vdd.n189 756.745
R14782 vdd.n166 vdd.n130 756.745
R14783 vdd.n124 vdd.n88 756.745
R14784 vdd.n65 vdd.n29 756.745
R14785 vdd.n2108 vdd.n2072 756.745
R14786 vdd.n2167 vdd.n2131 756.745
R14787 vdd.n2006 vdd.n1970 756.745
R14788 vdd.n2065 vdd.n2029 756.745
R14789 vdd.n1905 vdd.n1869 756.745
R14790 vdd.n1964 vdd.n1928 756.745
R14791 vdd.n1253 vdd.t221 640.208
R14792 vdd.n981 vdd.t263 640.208
R14793 vdd.n1273 vdd.t236 640.208
R14794 vdd.n972 vdd.t287 640.208
R14795 vdd.n872 vdd.t243 640.208
R14796 vdd.n2704 vdd.t281 640.208
R14797 vdd.n832 vdd.t290 640.208
R14798 vdd.n2701 vdd.t267 640.208
R14799 vdd.n799 vdd.t217 640.208
R14800 vdd.n1043 vdd.t274 640.208
R14801 vdd.n1679 vdd.t253 592.009
R14802 vdd.n1717 vdd.t271 592.009
R14803 vdd.n1613 vdd.t284 592.009
R14804 vdd.n2269 vdd.t229 592.009
R14805 vdd.n1190 vdd.t260 592.009
R14806 vdd.n1150 vdd.t278 592.009
R14807 vdd.n426 vdd.t250 592.009
R14808 vdd.n440 vdd.t239 592.009
R14809 vdd.n452 vdd.t257 592.009
R14810 vdd.n768 vdd.t233 592.009
R14811 vdd.n3276 vdd.t247 592.009
R14812 vdd.n688 vdd.t225 592.009
R14813 vdd.n328 vdd.n327 585
R14814 vdd.n326 vdd.n293 585
R14815 vdd.n325 vdd.n324 585
R14816 vdd.n296 vdd.n294 585
R14817 vdd.n319 vdd.n318 585
R14818 vdd.n317 vdd.n316 585
R14819 vdd.n300 vdd.n299 585
R14820 vdd.n311 vdd.n310 585
R14821 vdd.n309 vdd.n308 585
R14822 vdd.n304 vdd.n303 585
R14823 vdd.n269 vdd.n268 585
R14824 vdd.n267 vdd.n234 585
R14825 vdd.n266 vdd.n265 585
R14826 vdd.n237 vdd.n235 585
R14827 vdd.n260 vdd.n259 585
R14828 vdd.n258 vdd.n257 585
R14829 vdd.n241 vdd.n240 585
R14830 vdd.n252 vdd.n251 585
R14831 vdd.n250 vdd.n249 585
R14832 vdd.n245 vdd.n244 585
R14833 vdd.n226 vdd.n225 585
R14834 vdd.n224 vdd.n191 585
R14835 vdd.n223 vdd.n222 585
R14836 vdd.n194 vdd.n192 585
R14837 vdd.n217 vdd.n216 585
R14838 vdd.n215 vdd.n214 585
R14839 vdd.n198 vdd.n197 585
R14840 vdd.n209 vdd.n208 585
R14841 vdd.n207 vdd.n206 585
R14842 vdd.n202 vdd.n201 585
R14843 vdd.n167 vdd.n166 585
R14844 vdd.n165 vdd.n132 585
R14845 vdd.n164 vdd.n163 585
R14846 vdd.n135 vdd.n133 585
R14847 vdd.n158 vdd.n157 585
R14848 vdd.n156 vdd.n155 585
R14849 vdd.n139 vdd.n138 585
R14850 vdd.n150 vdd.n149 585
R14851 vdd.n148 vdd.n147 585
R14852 vdd.n143 vdd.n142 585
R14853 vdd.n125 vdd.n124 585
R14854 vdd.n123 vdd.n90 585
R14855 vdd.n122 vdd.n121 585
R14856 vdd.n93 vdd.n91 585
R14857 vdd.n116 vdd.n115 585
R14858 vdd.n114 vdd.n113 585
R14859 vdd.n97 vdd.n96 585
R14860 vdd.n108 vdd.n107 585
R14861 vdd.n106 vdd.n105 585
R14862 vdd.n101 vdd.n100 585
R14863 vdd.n66 vdd.n65 585
R14864 vdd.n64 vdd.n31 585
R14865 vdd.n63 vdd.n62 585
R14866 vdd.n34 vdd.n32 585
R14867 vdd.n57 vdd.n56 585
R14868 vdd.n55 vdd.n54 585
R14869 vdd.n38 vdd.n37 585
R14870 vdd.n49 vdd.n48 585
R14871 vdd.n47 vdd.n46 585
R14872 vdd.n42 vdd.n41 585
R14873 vdd.n2109 vdd.n2108 585
R14874 vdd.n2107 vdd.n2074 585
R14875 vdd.n2106 vdd.n2105 585
R14876 vdd.n2077 vdd.n2075 585
R14877 vdd.n2100 vdd.n2099 585
R14878 vdd.n2098 vdd.n2097 585
R14879 vdd.n2081 vdd.n2080 585
R14880 vdd.n2092 vdd.n2091 585
R14881 vdd.n2090 vdd.n2089 585
R14882 vdd.n2085 vdd.n2084 585
R14883 vdd.n2168 vdd.n2167 585
R14884 vdd.n2166 vdd.n2133 585
R14885 vdd.n2165 vdd.n2164 585
R14886 vdd.n2136 vdd.n2134 585
R14887 vdd.n2159 vdd.n2158 585
R14888 vdd.n2157 vdd.n2156 585
R14889 vdd.n2140 vdd.n2139 585
R14890 vdd.n2151 vdd.n2150 585
R14891 vdd.n2149 vdd.n2148 585
R14892 vdd.n2144 vdd.n2143 585
R14893 vdd.n2007 vdd.n2006 585
R14894 vdd.n2005 vdd.n1972 585
R14895 vdd.n2004 vdd.n2003 585
R14896 vdd.n1975 vdd.n1973 585
R14897 vdd.n1998 vdd.n1997 585
R14898 vdd.n1996 vdd.n1995 585
R14899 vdd.n1979 vdd.n1978 585
R14900 vdd.n1990 vdd.n1989 585
R14901 vdd.n1988 vdd.n1987 585
R14902 vdd.n1983 vdd.n1982 585
R14903 vdd.n2066 vdd.n2065 585
R14904 vdd.n2064 vdd.n2031 585
R14905 vdd.n2063 vdd.n2062 585
R14906 vdd.n2034 vdd.n2032 585
R14907 vdd.n2057 vdd.n2056 585
R14908 vdd.n2055 vdd.n2054 585
R14909 vdd.n2038 vdd.n2037 585
R14910 vdd.n2049 vdd.n2048 585
R14911 vdd.n2047 vdd.n2046 585
R14912 vdd.n2042 vdd.n2041 585
R14913 vdd.n1906 vdd.n1905 585
R14914 vdd.n1904 vdd.n1871 585
R14915 vdd.n1903 vdd.n1902 585
R14916 vdd.n1874 vdd.n1872 585
R14917 vdd.n1897 vdd.n1896 585
R14918 vdd.n1895 vdd.n1894 585
R14919 vdd.n1878 vdd.n1877 585
R14920 vdd.n1889 vdd.n1888 585
R14921 vdd.n1887 vdd.n1886 585
R14922 vdd.n1882 vdd.n1881 585
R14923 vdd.n1965 vdd.n1964 585
R14924 vdd.n1963 vdd.n1930 585
R14925 vdd.n1962 vdd.n1961 585
R14926 vdd.n1933 vdd.n1931 585
R14927 vdd.n1956 vdd.n1955 585
R14928 vdd.n1954 vdd.n1953 585
R14929 vdd.n1937 vdd.n1936 585
R14930 vdd.n1948 vdd.n1947 585
R14931 vdd.n1946 vdd.n1945 585
R14932 vdd.n1941 vdd.n1940 585
R14933 vdd.n3448 vdd.n392 509.269
R14934 vdd.n3444 vdd.n393 509.269
R14935 vdd.n3316 vdd.n685 509.269
R14936 vdd.n3313 vdd.n684 509.269
R14937 vdd.n2264 vdd.n1437 509.269
R14938 vdd.n2267 vdd.n2266 509.269
R14939 vdd.n1586 vdd.n1550 509.269
R14940 vdd.n1782 vdd.n1551 509.269
R14941 vdd.n305 vdd.t38 329.043
R14942 vdd.n246 vdd.t124 329.043
R14943 vdd.n203 vdd.t174 329.043
R14944 vdd.n144 vdd.t107 329.043
R14945 vdd.n102 vdd.t75 329.043
R14946 vdd.n43 vdd.t64 329.043
R14947 vdd.n2086 vdd.t165 329.043
R14948 vdd.n2145 vdd.t99 329.043
R14949 vdd.n1984 vdd.t153 329.043
R14950 vdd.n2043 vdd.t76 329.043
R14951 vdd.n1883 vdd.t66 329.043
R14952 vdd.n1942 vdd.t74 329.043
R14953 vdd.n1679 vdd.t256 319.788
R14954 vdd.n1717 vdd.t273 319.788
R14955 vdd.n1613 vdd.t286 319.788
R14956 vdd.n2269 vdd.t231 319.788
R14957 vdd.n1190 vdd.t261 319.788
R14958 vdd.n1150 vdd.t279 319.788
R14959 vdd.n426 vdd.t251 319.788
R14960 vdd.n440 vdd.t241 319.788
R14961 vdd.n452 vdd.t258 319.788
R14962 vdd.n768 vdd.t235 319.788
R14963 vdd.n3276 vdd.t249 319.788
R14964 vdd.n688 vdd.t228 319.788
R14965 vdd.n1680 vdd.t255 303.69
R14966 vdd.n1718 vdd.t272 303.69
R14967 vdd.n1614 vdd.t285 303.69
R14968 vdd.n2270 vdd.t232 303.69
R14969 vdd.n1191 vdd.t262 303.69
R14970 vdd.n1151 vdd.t280 303.69
R14971 vdd.n427 vdd.t252 303.69
R14972 vdd.n441 vdd.t242 303.69
R14973 vdd.n453 vdd.t259 303.69
R14974 vdd.n769 vdd.t234 303.69
R14975 vdd.n3277 vdd.t248 303.69
R14976 vdd.n689 vdd.t227 303.69
R14977 vdd.n2936 vdd.n927 291.221
R14978 vdd.n3150 vdd.n809 291.221
R14979 vdd.n3087 vdd.n806 291.221
R14980 vdd.n2868 vdd.n2867 291.221
R14981 vdd.n2664 vdd.n969 291.221
R14982 vdd.n2595 vdd.n2594 291.221
R14983 vdd.n1309 vdd.n1308 291.221
R14984 vdd.n2415 vdd.n1075 291.221
R14985 vdd.n3066 vdd.n807 291.221
R14986 vdd.n3153 vdd.n3152 291.221
R14987 vdd.n2772 vdd.n2698 291.221
R14988 vdd.n2940 vdd.n931 291.221
R14989 vdd.n2592 vdd.n979 291.221
R14990 vdd.n977 vdd.n951 291.221
R14991 vdd.n1387 vdd.n1116 291.221
R14992 vdd.n2419 vdd.n1080 291.221
R14993 vdd.n3068 vdd.n807 185
R14994 vdd.n3151 vdd.n807 185
R14995 vdd.n3070 vdd.n3069 185
R14996 vdd.n3069 vdd.n805 185
R14997 vdd.n3071 vdd.n839 185
R14998 vdd.n3081 vdd.n839 185
R14999 vdd.n3072 vdd.n848 185
R15000 vdd.n848 vdd.n846 185
R15001 vdd.n3074 vdd.n3073 185
R15002 vdd.n3075 vdd.n3074 185
R15003 vdd.n3027 vdd.n847 185
R15004 vdd.n847 vdd.n843 185
R15005 vdd.n3026 vdd.n3025 185
R15006 vdd.n3025 vdd.n3024 185
R15007 vdd.n850 vdd.n849 185
R15008 vdd.n851 vdd.n850 185
R15009 vdd.n3017 vdd.n3016 185
R15010 vdd.n3018 vdd.n3017 185
R15011 vdd.n3015 vdd.n860 185
R15012 vdd.n860 vdd.n857 185
R15013 vdd.n3014 vdd.n3013 185
R15014 vdd.n3013 vdd.n3012 185
R15015 vdd.n862 vdd.n861 185
R15016 vdd.n870 vdd.n862 185
R15017 vdd.n3005 vdd.n3004 185
R15018 vdd.n3006 vdd.n3005 185
R15019 vdd.n3002 vdd.n871 185
R15020 vdd.n878 vdd.n871 185
R15021 vdd.n3001 vdd.n3000 185
R15022 vdd.n3000 vdd.n2999 185
R15023 vdd.n874 vdd.n873 185
R15024 vdd.n875 vdd.n874 185
R15025 vdd.n2992 vdd.n2991 185
R15026 vdd.n2993 vdd.n2992 185
R15027 vdd.n2990 vdd.n885 185
R15028 vdd.n885 vdd.n882 185
R15029 vdd.n2989 vdd.n2988 185
R15030 vdd.n2988 vdd.n2987 185
R15031 vdd.n887 vdd.n886 185
R15032 vdd.n895 vdd.n887 185
R15033 vdd.n2980 vdd.n2979 185
R15034 vdd.n2981 vdd.n2980 185
R15035 vdd.n2978 vdd.n896 185
R15036 vdd.n901 vdd.n896 185
R15037 vdd.n2977 vdd.n2976 185
R15038 vdd.n2976 vdd.n2975 185
R15039 vdd.n898 vdd.n897 185
R15040 vdd.n2847 vdd.n898 185
R15041 vdd.n2968 vdd.n2967 185
R15042 vdd.n2969 vdd.n2968 185
R15043 vdd.n2966 vdd.n908 185
R15044 vdd.n908 vdd.n905 185
R15045 vdd.n2965 vdd.n2964 185
R15046 vdd.n2964 vdd.n2963 185
R15047 vdd.n910 vdd.n909 185
R15048 vdd.n911 vdd.n910 185
R15049 vdd.n2956 vdd.n2955 185
R15050 vdd.n2957 vdd.n2956 185
R15051 vdd.n2954 vdd.n920 185
R15052 vdd.n920 vdd.n917 185
R15053 vdd.n2953 vdd.n2952 185
R15054 vdd.n2952 vdd.n2951 185
R15055 vdd.n922 vdd.n921 185
R15056 vdd.n2862 vdd.n922 185
R15057 vdd.n2944 vdd.n2943 185
R15058 vdd.n2945 vdd.n2944 185
R15059 vdd.n2942 vdd.n931 185
R15060 vdd.n931 vdd.n928 185
R15061 vdd.n2941 vdd.n2940 185
R15062 vdd.n933 vdd.n932 185
R15063 vdd.n2708 vdd.n2707 185
R15064 vdd.n2710 vdd.n2709 185
R15065 vdd.n2712 vdd.n2711 185
R15066 vdd.n2714 vdd.n2713 185
R15067 vdd.n2716 vdd.n2715 185
R15068 vdd.n2718 vdd.n2717 185
R15069 vdd.n2720 vdd.n2719 185
R15070 vdd.n2722 vdd.n2721 185
R15071 vdd.n2724 vdd.n2723 185
R15072 vdd.n2726 vdd.n2725 185
R15073 vdd.n2728 vdd.n2727 185
R15074 vdd.n2730 vdd.n2729 185
R15075 vdd.n2732 vdd.n2731 185
R15076 vdd.n2734 vdd.n2733 185
R15077 vdd.n2736 vdd.n2735 185
R15078 vdd.n2738 vdd.n2737 185
R15079 vdd.n2740 vdd.n2739 185
R15080 vdd.n2742 vdd.n2741 185
R15081 vdd.n2744 vdd.n2743 185
R15082 vdd.n2746 vdd.n2745 185
R15083 vdd.n2748 vdd.n2747 185
R15084 vdd.n2750 vdd.n2749 185
R15085 vdd.n2752 vdd.n2751 185
R15086 vdd.n2754 vdd.n2753 185
R15087 vdd.n2756 vdd.n2755 185
R15088 vdd.n2758 vdd.n2757 185
R15089 vdd.n2760 vdd.n2759 185
R15090 vdd.n2762 vdd.n2761 185
R15091 vdd.n2764 vdd.n2763 185
R15092 vdd.n2766 vdd.n2765 185
R15093 vdd.n2768 vdd.n2767 185
R15094 vdd.n2770 vdd.n2769 185
R15095 vdd.n2771 vdd.n2698 185
R15096 vdd.n2938 vdd.n2698 185
R15097 vdd.n3154 vdd.n3153 185
R15098 vdd.n3155 vdd.n798 185
R15099 vdd.n3157 vdd.n3156 185
R15100 vdd.n3159 vdd.n796 185
R15101 vdd.n3161 vdd.n3160 185
R15102 vdd.n3162 vdd.n795 185
R15103 vdd.n3164 vdd.n3163 185
R15104 vdd.n3166 vdd.n793 185
R15105 vdd.n3168 vdd.n3167 185
R15106 vdd.n3169 vdd.n792 185
R15107 vdd.n3171 vdd.n3170 185
R15108 vdd.n3173 vdd.n790 185
R15109 vdd.n3175 vdd.n3174 185
R15110 vdd.n3176 vdd.n789 185
R15111 vdd.n3178 vdd.n3177 185
R15112 vdd.n3180 vdd.n788 185
R15113 vdd.n3181 vdd.n786 185
R15114 vdd.n3184 vdd.n3183 185
R15115 vdd.n787 vdd.n785 185
R15116 vdd.n3040 vdd.n3039 185
R15117 vdd.n3042 vdd.n3041 185
R15118 vdd.n3044 vdd.n3036 185
R15119 vdd.n3046 vdd.n3045 185
R15120 vdd.n3047 vdd.n3035 185
R15121 vdd.n3049 vdd.n3048 185
R15122 vdd.n3051 vdd.n3033 185
R15123 vdd.n3053 vdd.n3052 185
R15124 vdd.n3054 vdd.n3032 185
R15125 vdd.n3056 vdd.n3055 185
R15126 vdd.n3058 vdd.n3030 185
R15127 vdd.n3060 vdd.n3059 185
R15128 vdd.n3061 vdd.n3029 185
R15129 vdd.n3063 vdd.n3062 185
R15130 vdd.n3065 vdd.n3028 185
R15131 vdd.n3067 vdd.n3066 185
R15132 vdd.n3066 vdd.n692 185
R15133 vdd.n3152 vdd.n802 185
R15134 vdd.n3152 vdd.n3151 185
R15135 vdd.n2775 vdd.n804 185
R15136 vdd.n805 vdd.n804 185
R15137 vdd.n2776 vdd.n838 185
R15138 vdd.n3081 vdd.n838 185
R15139 vdd.n2778 vdd.n2777 185
R15140 vdd.n2777 vdd.n846 185
R15141 vdd.n2779 vdd.n845 185
R15142 vdd.n3075 vdd.n845 185
R15143 vdd.n2781 vdd.n2780 185
R15144 vdd.n2780 vdd.n843 185
R15145 vdd.n2782 vdd.n853 185
R15146 vdd.n3024 vdd.n853 185
R15147 vdd.n2784 vdd.n2783 185
R15148 vdd.n2783 vdd.n851 185
R15149 vdd.n2785 vdd.n859 185
R15150 vdd.n3018 vdd.n859 185
R15151 vdd.n2787 vdd.n2786 185
R15152 vdd.n2786 vdd.n857 185
R15153 vdd.n2788 vdd.n864 185
R15154 vdd.n3012 vdd.n864 185
R15155 vdd.n2790 vdd.n2789 185
R15156 vdd.n2789 vdd.n870 185
R15157 vdd.n2791 vdd.n869 185
R15158 vdd.n3006 vdd.n869 185
R15159 vdd.n2793 vdd.n2792 185
R15160 vdd.n2792 vdd.n878 185
R15161 vdd.n2794 vdd.n877 185
R15162 vdd.n2999 vdd.n877 185
R15163 vdd.n2796 vdd.n2795 185
R15164 vdd.n2795 vdd.n875 185
R15165 vdd.n2797 vdd.n884 185
R15166 vdd.n2993 vdd.n884 185
R15167 vdd.n2799 vdd.n2798 185
R15168 vdd.n2798 vdd.n882 185
R15169 vdd.n2800 vdd.n889 185
R15170 vdd.n2987 vdd.n889 185
R15171 vdd.n2802 vdd.n2801 185
R15172 vdd.n2801 vdd.n895 185
R15173 vdd.n2803 vdd.n894 185
R15174 vdd.n2981 vdd.n894 185
R15175 vdd.n2805 vdd.n2804 185
R15176 vdd.n2804 vdd.n901 185
R15177 vdd.n2806 vdd.n900 185
R15178 vdd.n2975 vdd.n900 185
R15179 vdd.n2849 vdd.n2848 185
R15180 vdd.n2848 vdd.n2847 185
R15181 vdd.n2850 vdd.n907 185
R15182 vdd.n2969 vdd.n907 185
R15183 vdd.n2852 vdd.n2851 185
R15184 vdd.n2851 vdd.n905 185
R15185 vdd.n2853 vdd.n913 185
R15186 vdd.n2963 vdd.n913 185
R15187 vdd.n2855 vdd.n2854 185
R15188 vdd.n2854 vdd.n911 185
R15189 vdd.n2856 vdd.n919 185
R15190 vdd.n2957 vdd.n919 185
R15191 vdd.n2858 vdd.n2857 185
R15192 vdd.n2857 vdd.n917 185
R15193 vdd.n2859 vdd.n924 185
R15194 vdd.n2951 vdd.n924 185
R15195 vdd.n2861 vdd.n2860 185
R15196 vdd.n2862 vdd.n2861 185
R15197 vdd.n2774 vdd.n930 185
R15198 vdd.n2945 vdd.n930 185
R15199 vdd.n2773 vdd.n2772 185
R15200 vdd.n2772 vdd.n928 185
R15201 vdd.n2264 vdd.n2263 185
R15202 vdd.n2265 vdd.n2264 185
R15203 vdd.n1438 vdd.n1436 185
R15204 vdd.n2256 vdd.n1436 185
R15205 vdd.n2259 vdd.n2258 185
R15206 vdd.n2258 vdd.n2257 185
R15207 vdd.n1441 vdd.n1440 185
R15208 vdd.n1442 vdd.n1441 185
R15209 vdd.n2245 vdd.n2244 185
R15210 vdd.n2246 vdd.n2245 185
R15211 vdd.n1450 vdd.n1449 185
R15212 vdd.n2237 vdd.n1449 185
R15213 vdd.n2240 vdd.n2239 185
R15214 vdd.n2239 vdd.n2238 185
R15215 vdd.n1453 vdd.n1452 185
R15216 vdd.n1460 vdd.n1453 185
R15217 vdd.n2228 vdd.n2227 185
R15218 vdd.n2229 vdd.n2228 185
R15219 vdd.n1462 vdd.n1461 185
R15220 vdd.n1461 vdd.n1459 185
R15221 vdd.n2223 vdd.n2222 185
R15222 vdd.n2222 vdd.n2221 185
R15223 vdd.n1465 vdd.n1464 185
R15224 vdd.n1466 vdd.n1465 185
R15225 vdd.n2212 vdd.n2211 185
R15226 vdd.n2213 vdd.n2212 185
R15227 vdd.n1473 vdd.n1472 185
R15228 vdd.n2204 vdd.n1472 185
R15229 vdd.n2207 vdd.n2206 185
R15230 vdd.n2206 vdd.n2205 185
R15231 vdd.n1476 vdd.n1475 185
R15232 vdd.n1482 vdd.n1476 185
R15233 vdd.n2195 vdd.n2194 185
R15234 vdd.n2196 vdd.n2195 185
R15235 vdd.n1484 vdd.n1483 185
R15236 vdd.n2187 vdd.n1483 185
R15237 vdd.n2190 vdd.n2189 185
R15238 vdd.n2189 vdd.n2188 185
R15239 vdd.n1487 vdd.n1486 185
R15240 vdd.n1488 vdd.n1487 185
R15241 vdd.n2178 vdd.n2177 185
R15242 vdd.n2179 vdd.n2178 185
R15243 vdd.n1496 vdd.n1495 185
R15244 vdd.n1495 vdd.n1494 185
R15245 vdd.n1866 vdd.n1865 185
R15246 vdd.n1865 vdd.n1864 185
R15247 vdd.n1499 vdd.n1498 185
R15248 vdd.n1505 vdd.n1499 185
R15249 vdd.n1855 vdd.n1854 185
R15250 vdd.n1856 vdd.n1855 185
R15251 vdd.n1507 vdd.n1506 185
R15252 vdd.n1847 vdd.n1506 185
R15253 vdd.n1850 vdd.n1849 185
R15254 vdd.n1849 vdd.n1848 185
R15255 vdd.n1510 vdd.n1509 185
R15256 vdd.n1517 vdd.n1510 185
R15257 vdd.n1838 vdd.n1837 185
R15258 vdd.n1839 vdd.n1838 185
R15259 vdd.n1519 vdd.n1518 185
R15260 vdd.n1518 vdd.n1516 185
R15261 vdd.n1833 vdd.n1832 185
R15262 vdd.n1832 vdd.n1831 185
R15263 vdd.n1522 vdd.n1521 185
R15264 vdd.n1523 vdd.n1522 185
R15265 vdd.n1822 vdd.n1821 185
R15266 vdd.n1823 vdd.n1822 185
R15267 vdd.n1530 vdd.n1529 185
R15268 vdd.n1814 vdd.n1529 185
R15269 vdd.n1817 vdd.n1816 185
R15270 vdd.n1816 vdd.n1815 185
R15271 vdd.n1533 vdd.n1532 185
R15272 vdd.n1539 vdd.n1533 185
R15273 vdd.n1805 vdd.n1804 185
R15274 vdd.n1806 vdd.n1805 185
R15275 vdd.n1541 vdd.n1540 185
R15276 vdd.n1797 vdd.n1540 185
R15277 vdd.n1800 vdd.n1799 185
R15278 vdd.n1799 vdd.n1798 185
R15279 vdd.n1544 vdd.n1543 185
R15280 vdd.n1545 vdd.n1544 185
R15281 vdd.n1788 vdd.n1787 185
R15282 vdd.n1789 vdd.n1788 185
R15283 vdd.n1552 vdd.n1551 185
R15284 vdd.n1587 vdd.n1551 185
R15285 vdd.n1783 vdd.n1782 185
R15286 vdd.n1555 vdd.n1554 185
R15287 vdd.n1779 vdd.n1778 185
R15288 vdd.n1780 vdd.n1779 185
R15289 vdd.n1589 vdd.n1588 185
R15290 vdd.n1774 vdd.n1591 185
R15291 vdd.n1773 vdd.n1592 185
R15292 vdd.n1772 vdd.n1593 185
R15293 vdd.n1595 vdd.n1594 185
R15294 vdd.n1768 vdd.n1597 185
R15295 vdd.n1767 vdd.n1598 185
R15296 vdd.n1766 vdd.n1599 185
R15297 vdd.n1601 vdd.n1600 185
R15298 vdd.n1762 vdd.n1603 185
R15299 vdd.n1761 vdd.n1604 185
R15300 vdd.n1760 vdd.n1605 185
R15301 vdd.n1607 vdd.n1606 185
R15302 vdd.n1756 vdd.n1609 185
R15303 vdd.n1755 vdd.n1610 185
R15304 vdd.n1754 vdd.n1611 185
R15305 vdd.n1615 vdd.n1612 185
R15306 vdd.n1750 vdd.n1617 185
R15307 vdd.n1749 vdd.n1618 185
R15308 vdd.n1748 vdd.n1619 185
R15309 vdd.n1621 vdd.n1620 185
R15310 vdd.n1744 vdd.n1623 185
R15311 vdd.n1743 vdd.n1624 185
R15312 vdd.n1742 vdd.n1625 185
R15313 vdd.n1627 vdd.n1626 185
R15314 vdd.n1738 vdd.n1629 185
R15315 vdd.n1737 vdd.n1630 185
R15316 vdd.n1736 vdd.n1631 185
R15317 vdd.n1633 vdd.n1632 185
R15318 vdd.n1732 vdd.n1635 185
R15319 vdd.n1731 vdd.n1636 185
R15320 vdd.n1730 vdd.n1637 185
R15321 vdd.n1639 vdd.n1638 185
R15322 vdd.n1726 vdd.n1641 185
R15323 vdd.n1725 vdd.n1642 185
R15324 vdd.n1724 vdd.n1643 185
R15325 vdd.n1645 vdd.n1644 185
R15326 vdd.n1720 vdd.n1647 185
R15327 vdd.n1719 vdd.n1716 185
R15328 vdd.n1715 vdd.n1648 185
R15329 vdd.n1650 vdd.n1649 185
R15330 vdd.n1711 vdd.n1652 185
R15331 vdd.n1710 vdd.n1653 185
R15332 vdd.n1709 vdd.n1654 185
R15333 vdd.n1656 vdd.n1655 185
R15334 vdd.n1705 vdd.n1658 185
R15335 vdd.n1704 vdd.n1659 185
R15336 vdd.n1703 vdd.n1660 185
R15337 vdd.n1662 vdd.n1661 185
R15338 vdd.n1699 vdd.n1664 185
R15339 vdd.n1698 vdd.n1665 185
R15340 vdd.n1697 vdd.n1666 185
R15341 vdd.n1668 vdd.n1667 185
R15342 vdd.n1693 vdd.n1670 185
R15343 vdd.n1692 vdd.n1671 185
R15344 vdd.n1691 vdd.n1672 185
R15345 vdd.n1674 vdd.n1673 185
R15346 vdd.n1687 vdd.n1676 185
R15347 vdd.n1686 vdd.n1677 185
R15348 vdd.n1685 vdd.n1678 185
R15349 vdd.n1682 vdd.n1586 185
R15350 vdd.n1780 vdd.n1586 185
R15351 vdd.n2268 vdd.n2267 185
R15352 vdd.n2272 vdd.n1432 185
R15353 vdd.n1431 vdd.n1425 185
R15354 vdd.n1429 vdd.n1428 185
R15355 vdd.n1427 vdd.n1221 185
R15356 vdd.n2276 vdd.n1218 185
R15357 vdd.n2278 vdd.n2277 185
R15358 vdd.n2280 vdd.n1216 185
R15359 vdd.n2282 vdd.n2281 185
R15360 vdd.n2283 vdd.n1211 185
R15361 vdd.n2285 vdd.n2284 185
R15362 vdd.n2287 vdd.n1209 185
R15363 vdd.n2289 vdd.n2288 185
R15364 vdd.n2290 vdd.n1204 185
R15365 vdd.n2292 vdd.n2291 185
R15366 vdd.n2294 vdd.n1202 185
R15367 vdd.n2296 vdd.n2295 185
R15368 vdd.n2297 vdd.n1198 185
R15369 vdd.n2299 vdd.n2298 185
R15370 vdd.n2301 vdd.n1195 185
R15371 vdd.n2303 vdd.n2302 185
R15372 vdd.n1196 vdd.n1189 185
R15373 vdd.n2307 vdd.n1193 185
R15374 vdd.n2308 vdd.n1185 185
R15375 vdd.n2310 vdd.n2309 185
R15376 vdd.n2312 vdd.n1183 185
R15377 vdd.n2314 vdd.n2313 185
R15378 vdd.n2315 vdd.n1178 185
R15379 vdd.n2317 vdd.n2316 185
R15380 vdd.n2319 vdd.n1176 185
R15381 vdd.n2321 vdd.n2320 185
R15382 vdd.n2322 vdd.n1171 185
R15383 vdd.n2324 vdd.n2323 185
R15384 vdd.n2326 vdd.n1169 185
R15385 vdd.n2328 vdd.n2327 185
R15386 vdd.n2329 vdd.n1164 185
R15387 vdd.n2331 vdd.n2330 185
R15388 vdd.n2333 vdd.n1162 185
R15389 vdd.n2335 vdd.n2334 185
R15390 vdd.n2336 vdd.n1158 185
R15391 vdd.n2338 vdd.n2337 185
R15392 vdd.n2340 vdd.n1155 185
R15393 vdd.n2342 vdd.n2341 185
R15394 vdd.n1156 vdd.n1149 185
R15395 vdd.n2346 vdd.n1153 185
R15396 vdd.n2347 vdd.n1145 185
R15397 vdd.n2349 vdd.n2348 185
R15398 vdd.n2351 vdd.n1143 185
R15399 vdd.n2353 vdd.n2352 185
R15400 vdd.n2354 vdd.n1138 185
R15401 vdd.n2356 vdd.n2355 185
R15402 vdd.n2358 vdd.n1136 185
R15403 vdd.n2360 vdd.n2359 185
R15404 vdd.n2361 vdd.n1131 185
R15405 vdd.n2363 vdd.n2362 185
R15406 vdd.n2365 vdd.n1129 185
R15407 vdd.n2367 vdd.n2366 185
R15408 vdd.n2368 vdd.n1127 185
R15409 vdd.n2370 vdd.n2369 185
R15410 vdd.n2373 vdd.n2372 185
R15411 vdd.n2375 vdd.n2374 185
R15412 vdd.n2377 vdd.n1125 185
R15413 vdd.n2379 vdd.n2378 185
R15414 vdd.n1437 vdd.n1124 185
R15415 vdd.n2266 vdd.n1435 185
R15416 vdd.n2266 vdd.n2265 185
R15417 vdd.n1445 vdd.n1434 185
R15418 vdd.n2256 vdd.n1434 185
R15419 vdd.n2255 vdd.n2254 185
R15420 vdd.n2257 vdd.n2255 185
R15421 vdd.n1444 vdd.n1443 185
R15422 vdd.n1443 vdd.n1442 185
R15423 vdd.n2248 vdd.n2247 185
R15424 vdd.n2247 vdd.n2246 185
R15425 vdd.n1448 vdd.n1447 185
R15426 vdd.n2237 vdd.n1448 185
R15427 vdd.n2236 vdd.n2235 185
R15428 vdd.n2238 vdd.n2236 185
R15429 vdd.n1455 vdd.n1454 185
R15430 vdd.n1460 vdd.n1454 185
R15431 vdd.n2231 vdd.n2230 185
R15432 vdd.n2230 vdd.n2229 185
R15433 vdd.n1458 vdd.n1457 185
R15434 vdd.n1459 vdd.n1458 185
R15435 vdd.n2220 vdd.n2219 185
R15436 vdd.n2221 vdd.n2220 185
R15437 vdd.n1468 vdd.n1467 185
R15438 vdd.n1467 vdd.n1466 185
R15439 vdd.n2215 vdd.n2214 185
R15440 vdd.n2214 vdd.n2213 185
R15441 vdd.n1471 vdd.n1470 185
R15442 vdd.n2204 vdd.n1471 185
R15443 vdd.n2203 vdd.n2202 185
R15444 vdd.n2205 vdd.n2203 185
R15445 vdd.n1478 vdd.n1477 185
R15446 vdd.n1482 vdd.n1477 185
R15447 vdd.n2198 vdd.n2197 185
R15448 vdd.n2197 vdd.n2196 185
R15449 vdd.n1481 vdd.n1480 185
R15450 vdd.n2187 vdd.n1481 185
R15451 vdd.n2186 vdd.n2185 185
R15452 vdd.n2188 vdd.n2186 185
R15453 vdd.n1490 vdd.n1489 185
R15454 vdd.n1489 vdd.n1488 185
R15455 vdd.n2181 vdd.n2180 185
R15456 vdd.n2180 vdd.n2179 185
R15457 vdd.n1493 vdd.n1492 185
R15458 vdd.n1494 vdd.n1493 185
R15459 vdd.n1863 vdd.n1862 185
R15460 vdd.n1864 vdd.n1863 185
R15461 vdd.n1501 vdd.n1500 185
R15462 vdd.n1505 vdd.n1500 185
R15463 vdd.n1858 vdd.n1857 185
R15464 vdd.n1857 vdd.n1856 185
R15465 vdd.n1504 vdd.n1503 185
R15466 vdd.n1847 vdd.n1504 185
R15467 vdd.n1846 vdd.n1845 185
R15468 vdd.n1848 vdd.n1846 185
R15469 vdd.n1512 vdd.n1511 185
R15470 vdd.n1517 vdd.n1511 185
R15471 vdd.n1841 vdd.n1840 185
R15472 vdd.n1840 vdd.n1839 185
R15473 vdd.n1515 vdd.n1514 185
R15474 vdd.n1516 vdd.n1515 185
R15475 vdd.n1830 vdd.n1829 185
R15476 vdd.n1831 vdd.n1830 185
R15477 vdd.n1525 vdd.n1524 185
R15478 vdd.n1524 vdd.n1523 185
R15479 vdd.n1825 vdd.n1824 185
R15480 vdd.n1824 vdd.n1823 185
R15481 vdd.n1528 vdd.n1527 185
R15482 vdd.n1814 vdd.n1528 185
R15483 vdd.n1813 vdd.n1812 185
R15484 vdd.n1815 vdd.n1813 185
R15485 vdd.n1535 vdd.n1534 185
R15486 vdd.n1539 vdd.n1534 185
R15487 vdd.n1808 vdd.n1807 185
R15488 vdd.n1807 vdd.n1806 185
R15489 vdd.n1538 vdd.n1537 185
R15490 vdd.n1797 vdd.n1538 185
R15491 vdd.n1796 vdd.n1795 185
R15492 vdd.n1798 vdd.n1796 185
R15493 vdd.n1547 vdd.n1546 185
R15494 vdd.n1546 vdd.n1545 185
R15495 vdd.n1791 vdd.n1790 185
R15496 vdd.n1790 vdd.n1789 185
R15497 vdd.n1550 vdd.n1549 185
R15498 vdd.n1587 vdd.n1550 185
R15499 vdd.n971 vdd.n969 185
R15500 vdd.n2593 vdd.n969 185
R15501 vdd.n2515 vdd.n989 185
R15502 vdd.n989 vdd.n976 185
R15503 vdd.n2517 vdd.n2516 185
R15504 vdd.n2518 vdd.n2517 185
R15505 vdd.n2514 vdd.n988 185
R15506 vdd.n1338 vdd.n988 185
R15507 vdd.n2513 vdd.n2512 185
R15508 vdd.n2512 vdd.n2511 185
R15509 vdd.n991 vdd.n990 185
R15510 vdd.n992 vdd.n991 185
R15511 vdd.n2502 vdd.n2501 185
R15512 vdd.n2503 vdd.n2502 185
R15513 vdd.n2500 vdd.n1002 185
R15514 vdd.n1002 vdd.n999 185
R15515 vdd.n2499 vdd.n2498 185
R15516 vdd.n2498 vdd.n2497 185
R15517 vdd.n1004 vdd.n1003 185
R15518 vdd.n1005 vdd.n1004 185
R15519 vdd.n2490 vdd.n2489 185
R15520 vdd.n2491 vdd.n2490 185
R15521 vdd.n2488 vdd.n1013 185
R15522 vdd.n1018 vdd.n1013 185
R15523 vdd.n2487 vdd.n2486 185
R15524 vdd.n2486 vdd.n2485 185
R15525 vdd.n1015 vdd.n1014 185
R15526 vdd.n1024 vdd.n1015 185
R15527 vdd.n2478 vdd.n2477 185
R15528 vdd.n2479 vdd.n2478 185
R15529 vdd.n2476 vdd.n1025 185
R15530 vdd.n1359 vdd.n1025 185
R15531 vdd.n2475 vdd.n2474 185
R15532 vdd.n2474 vdd.n2473 185
R15533 vdd.n1027 vdd.n1026 185
R15534 vdd.n1028 vdd.n1027 185
R15535 vdd.n2466 vdd.n2465 185
R15536 vdd.n2467 vdd.n2466 185
R15537 vdd.n2464 vdd.n1037 185
R15538 vdd.n1037 vdd.n1034 185
R15539 vdd.n2463 vdd.n2462 185
R15540 vdd.n2462 vdd.n2461 185
R15541 vdd.n1039 vdd.n1038 185
R15542 vdd.n1048 vdd.n1039 185
R15543 vdd.n2453 vdd.n2452 185
R15544 vdd.n2454 vdd.n2453 185
R15545 vdd.n2451 vdd.n1049 185
R15546 vdd.n1055 vdd.n1049 185
R15547 vdd.n2450 vdd.n2449 185
R15548 vdd.n2449 vdd.n2448 185
R15549 vdd.n1051 vdd.n1050 185
R15550 vdd.n1052 vdd.n1051 185
R15551 vdd.n2441 vdd.n2440 185
R15552 vdd.n2442 vdd.n2441 185
R15553 vdd.n2439 vdd.n1062 185
R15554 vdd.n1062 vdd.n1059 185
R15555 vdd.n2438 vdd.n2437 185
R15556 vdd.n2437 vdd.n2436 185
R15557 vdd.n1064 vdd.n1063 185
R15558 vdd.n1065 vdd.n1064 185
R15559 vdd.n2429 vdd.n2428 185
R15560 vdd.n2430 vdd.n2429 185
R15561 vdd.n2427 vdd.n1073 185
R15562 vdd.n1079 vdd.n1073 185
R15563 vdd.n2426 vdd.n2425 185
R15564 vdd.n2425 vdd.n2424 185
R15565 vdd.n1075 vdd.n1074 185
R15566 vdd.n1076 vdd.n1075 185
R15567 vdd.n2415 vdd.n2414 185
R15568 vdd.n2413 vdd.n1118 185
R15569 vdd.n2412 vdd.n1117 185
R15570 vdd.n2417 vdd.n1117 185
R15571 vdd.n2411 vdd.n2410 185
R15572 vdd.n2409 vdd.n2408 185
R15573 vdd.n2407 vdd.n2406 185
R15574 vdd.n2405 vdd.n2404 185
R15575 vdd.n2403 vdd.n2402 185
R15576 vdd.n2401 vdd.n2400 185
R15577 vdd.n2399 vdd.n2398 185
R15578 vdd.n2397 vdd.n2396 185
R15579 vdd.n2395 vdd.n2394 185
R15580 vdd.n2393 vdd.n2392 185
R15581 vdd.n2391 vdd.n2390 185
R15582 vdd.n2389 vdd.n2388 185
R15583 vdd.n2387 vdd.n2386 185
R15584 vdd.n2385 vdd.n2384 185
R15585 vdd.n2383 vdd.n2382 185
R15586 vdd.n1275 vdd.n1119 185
R15587 vdd.n1277 vdd.n1276 185
R15588 vdd.n1279 vdd.n1278 185
R15589 vdd.n1281 vdd.n1280 185
R15590 vdd.n1283 vdd.n1282 185
R15591 vdd.n1285 vdd.n1284 185
R15592 vdd.n1287 vdd.n1286 185
R15593 vdd.n1289 vdd.n1288 185
R15594 vdd.n1291 vdd.n1290 185
R15595 vdd.n1293 vdd.n1292 185
R15596 vdd.n1295 vdd.n1294 185
R15597 vdd.n1297 vdd.n1296 185
R15598 vdd.n1299 vdd.n1298 185
R15599 vdd.n1301 vdd.n1300 185
R15600 vdd.n1304 vdd.n1303 185
R15601 vdd.n1306 vdd.n1305 185
R15602 vdd.n1308 vdd.n1307 185
R15603 vdd.n2596 vdd.n2595 185
R15604 vdd.n2598 vdd.n2597 185
R15605 vdd.n2600 vdd.n2599 185
R15606 vdd.n2603 vdd.n2602 185
R15607 vdd.n2605 vdd.n2604 185
R15608 vdd.n2607 vdd.n2606 185
R15609 vdd.n2609 vdd.n2608 185
R15610 vdd.n2611 vdd.n2610 185
R15611 vdd.n2613 vdd.n2612 185
R15612 vdd.n2615 vdd.n2614 185
R15613 vdd.n2617 vdd.n2616 185
R15614 vdd.n2619 vdd.n2618 185
R15615 vdd.n2621 vdd.n2620 185
R15616 vdd.n2623 vdd.n2622 185
R15617 vdd.n2625 vdd.n2624 185
R15618 vdd.n2627 vdd.n2626 185
R15619 vdd.n2629 vdd.n2628 185
R15620 vdd.n2631 vdd.n2630 185
R15621 vdd.n2633 vdd.n2632 185
R15622 vdd.n2635 vdd.n2634 185
R15623 vdd.n2637 vdd.n2636 185
R15624 vdd.n2639 vdd.n2638 185
R15625 vdd.n2641 vdd.n2640 185
R15626 vdd.n2643 vdd.n2642 185
R15627 vdd.n2645 vdd.n2644 185
R15628 vdd.n2647 vdd.n2646 185
R15629 vdd.n2649 vdd.n2648 185
R15630 vdd.n2651 vdd.n2650 185
R15631 vdd.n2653 vdd.n2652 185
R15632 vdd.n2655 vdd.n2654 185
R15633 vdd.n2657 vdd.n2656 185
R15634 vdd.n2659 vdd.n2658 185
R15635 vdd.n2661 vdd.n2660 185
R15636 vdd.n2662 vdd.n970 185
R15637 vdd.n2664 vdd.n2663 185
R15638 vdd.n2665 vdd.n2664 185
R15639 vdd.n2594 vdd.n974 185
R15640 vdd.n2594 vdd.n2593 185
R15641 vdd.n1336 vdd.n975 185
R15642 vdd.n976 vdd.n975 185
R15643 vdd.n1337 vdd.n986 185
R15644 vdd.n2518 vdd.n986 185
R15645 vdd.n1340 vdd.n1339 185
R15646 vdd.n1339 vdd.n1338 185
R15647 vdd.n1341 vdd.n993 185
R15648 vdd.n2511 vdd.n993 185
R15649 vdd.n1343 vdd.n1342 185
R15650 vdd.n1342 vdd.n992 185
R15651 vdd.n1344 vdd.n1000 185
R15652 vdd.n2503 vdd.n1000 185
R15653 vdd.n1346 vdd.n1345 185
R15654 vdd.n1345 vdd.n999 185
R15655 vdd.n1347 vdd.n1006 185
R15656 vdd.n2497 vdd.n1006 185
R15657 vdd.n1349 vdd.n1348 185
R15658 vdd.n1348 vdd.n1005 185
R15659 vdd.n1350 vdd.n1011 185
R15660 vdd.n2491 vdd.n1011 185
R15661 vdd.n1352 vdd.n1351 185
R15662 vdd.n1351 vdd.n1018 185
R15663 vdd.n1353 vdd.n1016 185
R15664 vdd.n2485 vdd.n1016 185
R15665 vdd.n1355 vdd.n1354 185
R15666 vdd.n1354 vdd.n1024 185
R15667 vdd.n1356 vdd.n1022 185
R15668 vdd.n2479 vdd.n1022 185
R15669 vdd.n1358 vdd.n1357 185
R15670 vdd.n1359 vdd.n1358 185
R15671 vdd.n1335 vdd.n1029 185
R15672 vdd.n2473 vdd.n1029 185
R15673 vdd.n1334 vdd.n1333 185
R15674 vdd.n1333 vdd.n1028 185
R15675 vdd.n1332 vdd.n1035 185
R15676 vdd.n2467 vdd.n1035 185
R15677 vdd.n1331 vdd.n1330 185
R15678 vdd.n1330 vdd.n1034 185
R15679 vdd.n1329 vdd.n1040 185
R15680 vdd.n2461 vdd.n1040 185
R15681 vdd.n1328 vdd.n1327 185
R15682 vdd.n1327 vdd.n1048 185
R15683 vdd.n1326 vdd.n1046 185
R15684 vdd.n2454 vdd.n1046 185
R15685 vdd.n1325 vdd.n1324 185
R15686 vdd.n1324 vdd.n1055 185
R15687 vdd.n1323 vdd.n1053 185
R15688 vdd.n2448 vdd.n1053 185
R15689 vdd.n1322 vdd.n1321 185
R15690 vdd.n1321 vdd.n1052 185
R15691 vdd.n1320 vdd.n1060 185
R15692 vdd.n2442 vdd.n1060 185
R15693 vdd.n1319 vdd.n1318 185
R15694 vdd.n1318 vdd.n1059 185
R15695 vdd.n1317 vdd.n1066 185
R15696 vdd.n2436 vdd.n1066 185
R15697 vdd.n1316 vdd.n1315 185
R15698 vdd.n1315 vdd.n1065 185
R15699 vdd.n1314 vdd.n1071 185
R15700 vdd.n2430 vdd.n1071 185
R15701 vdd.n1313 vdd.n1312 185
R15702 vdd.n1312 vdd.n1079 185
R15703 vdd.n1311 vdd.n1077 185
R15704 vdd.n2424 vdd.n1077 185
R15705 vdd.n1310 vdd.n1309 185
R15706 vdd.n1309 vdd.n1076 185
R15707 vdd.n3449 vdd.n3448 185
R15708 vdd.n3448 vdd.n3447 185
R15709 vdd.n3450 vdd.n387 185
R15710 vdd.n387 vdd.n386 185
R15711 vdd.n3452 vdd.n3451 185
R15712 vdd.n3453 vdd.n3452 185
R15713 vdd.n382 vdd.n381 185
R15714 vdd.n3454 vdd.n382 185
R15715 vdd.n3457 vdd.n3456 185
R15716 vdd.n3456 vdd.n3455 185
R15717 vdd.n3458 vdd.n376 185
R15718 vdd.n376 vdd.n375 185
R15719 vdd.n3460 vdd.n3459 185
R15720 vdd.n3461 vdd.n3460 185
R15721 vdd.n371 vdd.n370 185
R15722 vdd.n3462 vdd.n371 185
R15723 vdd.n3465 vdd.n3464 185
R15724 vdd.n3464 vdd.n3463 185
R15725 vdd.n3466 vdd.n365 185
R15726 vdd.n3423 vdd.n365 185
R15727 vdd.n3468 vdd.n3467 185
R15728 vdd.n3469 vdd.n3468 185
R15729 vdd.n360 vdd.n359 185
R15730 vdd.n3470 vdd.n360 185
R15731 vdd.n3473 vdd.n3472 185
R15732 vdd.n3472 vdd.n3471 185
R15733 vdd.n3474 vdd.n354 185
R15734 vdd.n361 vdd.n354 185
R15735 vdd.n3476 vdd.n3475 185
R15736 vdd.n3477 vdd.n3476 185
R15737 vdd.n350 vdd.n349 185
R15738 vdd.n3478 vdd.n350 185
R15739 vdd.n3481 vdd.n3480 185
R15740 vdd.n3480 vdd.n3479 185
R15741 vdd.n3482 vdd.n345 185
R15742 vdd.n345 vdd.n344 185
R15743 vdd.n3484 vdd.n3483 185
R15744 vdd.n3485 vdd.n3484 185
R15745 vdd.n339 vdd.n337 185
R15746 vdd.n3486 vdd.n339 185
R15747 vdd.n3489 vdd.n3488 185
R15748 vdd.n3488 vdd.n3487 185
R15749 vdd.n338 vdd.n336 185
R15750 vdd.n340 vdd.n338 185
R15751 vdd.n3399 vdd.n3398 185
R15752 vdd.n3400 vdd.n3399 185
R15753 vdd.n635 vdd.n634 185
R15754 vdd.n634 vdd.n633 185
R15755 vdd.n3394 vdd.n3393 185
R15756 vdd.n3393 vdd.n3392 185
R15757 vdd.n638 vdd.n637 185
R15758 vdd.n644 vdd.n638 185
R15759 vdd.n3380 vdd.n3379 185
R15760 vdd.n3381 vdd.n3380 185
R15761 vdd.n646 vdd.n645 185
R15762 vdd.n3372 vdd.n645 185
R15763 vdd.n3375 vdd.n3374 185
R15764 vdd.n3374 vdd.n3373 185
R15765 vdd.n649 vdd.n648 185
R15766 vdd.n656 vdd.n649 185
R15767 vdd.n3363 vdd.n3362 185
R15768 vdd.n3364 vdd.n3363 185
R15769 vdd.n658 vdd.n657 185
R15770 vdd.n657 vdd.n655 185
R15771 vdd.n3358 vdd.n3357 185
R15772 vdd.n3357 vdd.n3356 185
R15773 vdd.n661 vdd.n660 185
R15774 vdd.n662 vdd.n661 185
R15775 vdd.n3347 vdd.n3346 185
R15776 vdd.n3348 vdd.n3347 185
R15777 vdd.n669 vdd.n668 185
R15778 vdd.n3339 vdd.n668 185
R15779 vdd.n3342 vdd.n3341 185
R15780 vdd.n3341 vdd.n3340 185
R15781 vdd.n672 vdd.n671 185
R15782 vdd.n679 vdd.n672 185
R15783 vdd.n3330 vdd.n3329 185
R15784 vdd.n3331 vdd.n3330 185
R15785 vdd.n681 vdd.n680 185
R15786 vdd.n680 vdd.n678 185
R15787 vdd.n3325 vdd.n3324 185
R15788 vdd.n3324 vdd.n3323 185
R15789 vdd.n684 vdd.n683 185
R15790 vdd.n723 vdd.n684 185
R15791 vdd.n3313 vdd.n3312 185
R15792 vdd.n3311 vdd.n725 185
R15793 vdd.n3310 vdd.n724 185
R15794 vdd.n3315 vdd.n724 185
R15795 vdd.n729 vdd.n728 185
R15796 vdd.n733 vdd.n732 185
R15797 vdd.n3306 vdd.n734 185
R15798 vdd.n3305 vdd.n3304 185
R15799 vdd.n3303 vdd.n3302 185
R15800 vdd.n3301 vdd.n3300 185
R15801 vdd.n3299 vdd.n3298 185
R15802 vdd.n3297 vdd.n3296 185
R15803 vdd.n3295 vdd.n3294 185
R15804 vdd.n3293 vdd.n3292 185
R15805 vdd.n3291 vdd.n3290 185
R15806 vdd.n3289 vdd.n3288 185
R15807 vdd.n3287 vdd.n3286 185
R15808 vdd.n3285 vdd.n3284 185
R15809 vdd.n3283 vdd.n3282 185
R15810 vdd.n3281 vdd.n3280 185
R15811 vdd.n3279 vdd.n3278 185
R15812 vdd.n3270 vdd.n747 185
R15813 vdd.n3272 vdd.n3271 185
R15814 vdd.n3269 vdd.n3268 185
R15815 vdd.n3267 vdd.n3266 185
R15816 vdd.n3265 vdd.n3264 185
R15817 vdd.n3263 vdd.n3262 185
R15818 vdd.n3261 vdd.n3260 185
R15819 vdd.n3259 vdd.n3258 185
R15820 vdd.n3257 vdd.n3256 185
R15821 vdd.n3255 vdd.n3254 185
R15822 vdd.n3253 vdd.n3252 185
R15823 vdd.n3251 vdd.n3250 185
R15824 vdd.n3249 vdd.n3248 185
R15825 vdd.n3247 vdd.n3246 185
R15826 vdd.n3245 vdd.n3244 185
R15827 vdd.n3243 vdd.n3242 185
R15828 vdd.n3241 vdd.n3240 185
R15829 vdd.n3239 vdd.n3238 185
R15830 vdd.n3237 vdd.n3236 185
R15831 vdd.n3235 vdd.n3234 185
R15832 vdd.n3233 vdd.n3232 185
R15833 vdd.n3231 vdd.n3230 185
R15834 vdd.n3224 vdd.n767 185
R15835 vdd.n3226 vdd.n3225 185
R15836 vdd.n3223 vdd.n3222 185
R15837 vdd.n3221 vdd.n3220 185
R15838 vdd.n3219 vdd.n3218 185
R15839 vdd.n3217 vdd.n3216 185
R15840 vdd.n3215 vdd.n3214 185
R15841 vdd.n3213 vdd.n3212 185
R15842 vdd.n3211 vdd.n3210 185
R15843 vdd.n3209 vdd.n3208 185
R15844 vdd.n3207 vdd.n3206 185
R15845 vdd.n3205 vdd.n3204 185
R15846 vdd.n3203 vdd.n3202 185
R15847 vdd.n3201 vdd.n3200 185
R15848 vdd.n3199 vdd.n3198 185
R15849 vdd.n3197 vdd.n3196 185
R15850 vdd.n3195 vdd.n3194 185
R15851 vdd.n3193 vdd.n3192 185
R15852 vdd.n3191 vdd.n3190 185
R15853 vdd.n3189 vdd.n3188 185
R15854 vdd.n3187 vdd.n691 185
R15855 vdd.n3317 vdd.n3316 185
R15856 vdd.n3316 vdd.n3315 185
R15857 vdd.n3444 vdd.n3443 185
R15858 vdd.n618 vdd.n425 185
R15859 vdd.n617 vdd.n616 185
R15860 vdd.n615 vdd.n614 185
R15861 vdd.n613 vdd.n430 185
R15862 vdd.n609 vdd.n608 185
R15863 vdd.n607 vdd.n606 185
R15864 vdd.n605 vdd.n604 185
R15865 vdd.n603 vdd.n432 185
R15866 vdd.n599 vdd.n598 185
R15867 vdd.n597 vdd.n596 185
R15868 vdd.n595 vdd.n594 185
R15869 vdd.n593 vdd.n434 185
R15870 vdd.n589 vdd.n588 185
R15871 vdd.n587 vdd.n586 185
R15872 vdd.n585 vdd.n584 185
R15873 vdd.n583 vdd.n436 185
R15874 vdd.n579 vdd.n578 185
R15875 vdd.n577 vdd.n576 185
R15876 vdd.n575 vdd.n574 185
R15877 vdd.n573 vdd.n438 185
R15878 vdd.n569 vdd.n568 185
R15879 vdd.n567 vdd.n566 185
R15880 vdd.n565 vdd.n564 185
R15881 vdd.n563 vdd.n442 185
R15882 vdd.n559 vdd.n558 185
R15883 vdd.n557 vdd.n556 185
R15884 vdd.n555 vdd.n554 185
R15885 vdd.n553 vdd.n444 185
R15886 vdd.n549 vdd.n548 185
R15887 vdd.n547 vdd.n546 185
R15888 vdd.n545 vdd.n544 185
R15889 vdd.n543 vdd.n446 185
R15890 vdd.n539 vdd.n538 185
R15891 vdd.n537 vdd.n536 185
R15892 vdd.n535 vdd.n534 185
R15893 vdd.n533 vdd.n448 185
R15894 vdd.n529 vdd.n528 185
R15895 vdd.n527 vdd.n526 185
R15896 vdd.n525 vdd.n524 185
R15897 vdd.n523 vdd.n450 185
R15898 vdd.n519 vdd.n518 185
R15899 vdd.n517 vdd.n516 185
R15900 vdd.n515 vdd.n514 185
R15901 vdd.n513 vdd.n454 185
R15902 vdd.n509 vdd.n508 185
R15903 vdd.n507 vdd.n506 185
R15904 vdd.n505 vdd.n504 185
R15905 vdd.n503 vdd.n456 185
R15906 vdd.n499 vdd.n498 185
R15907 vdd.n497 vdd.n496 185
R15908 vdd.n495 vdd.n494 185
R15909 vdd.n493 vdd.n458 185
R15910 vdd.n489 vdd.n488 185
R15911 vdd.n487 vdd.n486 185
R15912 vdd.n485 vdd.n484 185
R15913 vdd.n483 vdd.n460 185
R15914 vdd.n479 vdd.n478 185
R15915 vdd.n477 vdd.n476 185
R15916 vdd.n475 vdd.n474 185
R15917 vdd.n473 vdd.n462 185
R15918 vdd.n469 vdd.n468 185
R15919 vdd.n467 vdd.n466 185
R15920 vdd.n465 vdd.n392 185
R15921 vdd.n3440 vdd.n393 185
R15922 vdd.n3447 vdd.n393 185
R15923 vdd.n3439 vdd.n3438 185
R15924 vdd.n3438 vdd.n386 185
R15925 vdd.n3437 vdd.n385 185
R15926 vdd.n3453 vdd.n385 185
R15927 vdd.n621 vdd.n384 185
R15928 vdd.n3454 vdd.n384 185
R15929 vdd.n3433 vdd.n383 185
R15930 vdd.n3455 vdd.n383 185
R15931 vdd.n3432 vdd.n3431 185
R15932 vdd.n3431 vdd.n375 185
R15933 vdd.n3430 vdd.n374 185
R15934 vdd.n3461 vdd.n374 185
R15935 vdd.n623 vdd.n373 185
R15936 vdd.n3462 vdd.n373 185
R15937 vdd.n3426 vdd.n372 185
R15938 vdd.n3463 vdd.n372 185
R15939 vdd.n3425 vdd.n3424 185
R15940 vdd.n3424 vdd.n3423 185
R15941 vdd.n3422 vdd.n364 185
R15942 vdd.n3469 vdd.n364 185
R15943 vdd.n625 vdd.n363 185
R15944 vdd.n3470 vdd.n363 185
R15945 vdd.n3418 vdd.n362 185
R15946 vdd.n3471 vdd.n362 185
R15947 vdd.n3417 vdd.n3416 185
R15948 vdd.n3416 vdd.n361 185
R15949 vdd.n3415 vdd.n353 185
R15950 vdd.n3477 vdd.n353 185
R15951 vdd.n627 vdd.n352 185
R15952 vdd.n3478 vdd.n352 185
R15953 vdd.n3411 vdd.n351 185
R15954 vdd.n3479 vdd.n351 185
R15955 vdd.n3410 vdd.n3409 185
R15956 vdd.n3409 vdd.n344 185
R15957 vdd.n3408 vdd.n343 185
R15958 vdd.n3485 vdd.n343 185
R15959 vdd.n629 vdd.n342 185
R15960 vdd.n3486 vdd.n342 185
R15961 vdd.n3404 vdd.n341 185
R15962 vdd.n3487 vdd.n341 185
R15963 vdd.n3403 vdd.n3402 185
R15964 vdd.n3402 vdd.n340 185
R15965 vdd.n3401 vdd.n631 185
R15966 vdd.n3401 vdd.n3400 185
R15967 vdd.n3389 vdd.n632 185
R15968 vdd.n633 vdd.n632 185
R15969 vdd.n3391 vdd.n3390 185
R15970 vdd.n3392 vdd.n3391 185
R15971 vdd.n640 vdd.n639 185
R15972 vdd.n644 vdd.n639 185
R15973 vdd.n3383 vdd.n3382 185
R15974 vdd.n3382 vdd.n3381 185
R15975 vdd.n643 vdd.n642 185
R15976 vdd.n3372 vdd.n643 185
R15977 vdd.n3371 vdd.n3370 185
R15978 vdd.n3373 vdd.n3371 185
R15979 vdd.n651 vdd.n650 185
R15980 vdd.n656 vdd.n650 185
R15981 vdd.n3366 vdd.n3365 185
R15982 vdd.n3365 vdd.n3364 185
R15983 vdd.n654 vdd.n653 185
R15984 vdd.n655 vdd.n654 185
R15985 vdd.n3355 vdd.n3354 185
R15986 vdd.n3356 vdd.n3355 185
R15987 vdd.n664 vdd.n663 185
R15988 vdd.n663 vdd.n662 185
R15989 vdd.n3350 vdd.n3349 185
R15990 vdd.n3349 vdd.n3348 185
R15991 vdd.n667 vdd.n666 185
R15992 vdd.n3339 vdd.n667 185
R15993 vdd.n3338 vdd.n3337 185
R15994 vdd.n3340 vdd.n3338 185
R15995 vdd.n674 vdd.n673 185
R15996 vdd.n679 vdd.n673 185
R15997 vdd.n3333 vdd.n3332 185
R15998 vdd.n3332 vdd.n3331 185
R15999 vdd.n677 vdd.n676 185
R16000 vdd.n678 vdd.n677 185
R16001 vdd.n3322 vdd.n3321 185
R16002 vdd.n3323 vdd.n3322 185
R16003 vdd.n686 vdd.n685 185
R16004 vdd.n723 vdd.n685 185
R16005 vdd.n2936 vdd.n2935 185
R16006 vdd.n2934 vdd.n2700 185
R16007 vdd.n2933 vdd.n2699 185
R16008 vdd.n2938 vdd.n2699 185
R16009 vdd.n2932 vdd.n2931 185
R16010 vdd.n2930 vdd.n2929 185
R16011 vdd.n2928 vdd.n2927 185
R16012 vdd.n2926 vdd.n2925 185
R16013 vdd.n2924 vdd.n2923 185
R16014 vdd.n2922 vdd.n2921 185
R16015 vdd.n2920 vdd.n2919 185
R16016 vdd.n2918 vdd.n2917 185
R16017 vdd.n2916 vdd.n2915 185
R16018 vdd.n2914 vdd.n2913 185
R16019 vdd.n2912 vdd.n2911 185
R16020 vdd.n2910 vdd.n2909 185
R16021 vdd.n2908 vdd.n2907 185
R16022 vdd.n2906 vdd.n2905 185
R16023 vdd.n2904 vdd.n2903 185
R16024 vdd.n2902 vdd.n2901 185
R16025 vdd.n2900 vdd.n2899 185
R16026 vdd.n2898 vdd.n2897 185
R16027 vdd.n2896 vdd.n2895 185
R16028 vdd.n2894 vdd.n2893 185
R16029 vdd.n2892 vdd.n2891 185
R16030 vdd.n2890 vdd.n2889 185
R16031 vdd.n2888 vdd.n2887 185
R16032 vdd.n2886 vdd.n2885 185
R16033 vdd.n2884 vdd.n2883 185
R16034 vdd.n2882 vdd.n2881 185
R16035 vdd.n2880 vdd.n2879 185
R16036 vdd.n2878 vdd.n2877 185
R16037 vdd.n2876 vdd.n2875 185
R16038 vdd.n2873 vdd.n2872 185
R16039 vdd.n2871 vdd.n2870 185
R16040 vdd.n2869 vdd.n2868 185
R16041 vdd.n3087 vdd.n3086 185
R16042 vdd.n3089 vdd.n834 185
R16043 vdd.n3091 vdd.n3090 185
R16044 vdd.n3093 vdd.n831 185
R16045 vdd.n3095 vdd.n3094 185
R16046 vdd.n3097 vdd.n829 185
R16047 vdd.n3099 vdd.n3098 185
R16048 vdd.n3100 vdd.n828 185
R16049 vdd.n3102 vdd.n3101 185
R16050 vdd.n3104 vdd.n826 185
R16051 vdd.n3106 vdd.n3105 185
R16052 vdd.n3107 vdd.n825 185
R16053 vdd.n3109 vdd.n3108 185
R16054 vdd.n3111 vdd.n823 185
R16055 vdd.n3113 vdd.n3112 185
R16056 vdd.n3114 vdd.n822 185
R16057 vdd.n3116 vdd.n3115 185
R16058 vdd.n3118 vdd.n731 185
R16059 vdd.n3120 vdd.n3119 185
R16060 vdd.n3122 vdd.n820 185
R16061 vdd.n3124 vdd.n3123 185
R16062 vdd.n3125 vdd.n819 185
R16063 vdd.n3127 vdd.n3126 185
R16064 vdd.n3129 vdd.n817 185
R16065 vdd.n3131 vdd.n3130 185
R16066 vdd.n3132 vdd.n816 185
R16067 vdd.n3134 vdd.n3133 185
R16068 vdd.n3136 vdd.n814 185
R16069 vdd.n3138 vdd.n3137 185
R16070 vdd.n3139 vdd.n813 185
R16071 vdd.n3141 vdd.n3140 185
R16072 vdd.n3143 vdd.n812 185
R16073 vdd.n3144 vdd.n811 185
R16074 vdd.n3147 vdd.n3146 185
R16075 vdd.n3148 vdd.n809 185
R16076 vdd.n809 vdd.n692 185
R16077 vdd.n3085 vdd.n806 185
R16078 vdd.n3151 vdd.n806 185
R16079 vdd.n3084 vdd.n3083 185
R16080 vdd.n3083 vdd.n805 185
R16081 vdd.n3082 vdd.n836 185
R16082 vdd.n3082 vdd.n3081 185
R16083 vdd.n2816 vdd.n837 185
R16084 vdd.n846 vdd.n837 185
R16085 vdd.n2817 vdd.n844 185
R16086 vdd.n3075 vdd.n844 185
R16087 vdd.n2819 vdd.n2818 185
R16088 vdd.n2818 vdd.n843 185
R16089 vdd.n2820 vdd.n852 185
R16090 vdd.n3024 vdd.n852 185
R16091 vdd.n2822 vdd.n2821 185
R16092 vdd.n2821 vdd.n851 185
R16093 vdd.n2823 vdd.n858 185
R16094 vdd.n3018 vdd.n858 185
R16095 vdd.n2825 vdd.n2824 185
R16096 vdd.n2824 vdd.n857 185
R16097 vdd.n2826 vdd.n863 185
R16098 vdd.n3012 vdd.n863 185
R16099 vdd.n2828 vdd.n2827 185
R16100 vdd.n2827 vdd.n870 185
R16101 vdd.n2829 vdd.n868 185
R16102 vdd.n3006 vdd.n868 185
R16103 vdd.n2831 vdd.n2830 185
R16104 vdd.n2830 vdd.n878 185
R16105 vdd.n2832 vdd.n876 185
R16106 vdd.n2999 vdd.n876 185
R16107 vdd.n2834 vdd.n2833 185
R16108 vdd.n2833 vdd.n875 185
R16109 vdd.n2835 vdd.n883 185
R16110 vdd.n2993 vdd.n883 185
R16111 vdd.n2837 vdd.n2836 185
R16112 vdd.n2836 vdd.n882 185
R16113 vdd.n2838 vdd.n888 185
R16114 vdd.n2987 vdd.n888 185
R16115 vdd.n2840 vdd.n2839 185
R16116 vdd.n2839 vdd.n895 185
R16117 vdd.n2841 vdd.n893 185
R16118 vdd.n2981 vdd.n893 185
R16119 vdd.n2843 vdd.n2842 185
R16120 vdd.n2842 vdd.n901 185
R16121 vdd.n2844 vdd.n899 185
R16122 vdd.n2975 vdd.n899 185
R16123 vdd.n2846 vdd.n2845 185
R16124 vdd.n2847 vdd.n2846 185
R16125 vdd.n2815 vdd.n906 185
R16126 vdd.n2969 vdd.n906 185
R16127 vdd.n2814 vdd.n2813 185
R16128 vdd.n2813 vdd.n905 185
R16129 vdd.n2812 vdd.n912 185
R16130 vdd.n2963 vdd.n912 185
R16131 vdd.n2811 vdd.n2810 185
R16132 vdd.n2810 vdd.n911 185
R16133 vdd.n2809 vdd.n918 185
R16134 vdd.n2957 vdd.n918 185
R16135 vdd.n2808 vdd.n2807 185
R16136 vdd.n2807 vdd.n917 185
R16137 vdd.n2703 vdd.n923 185
R16138 vdd.n2951 vdd.n923 185
R16139 vdd.n2864 vdd.n2863 185
R16140 vdd.n2863 vdd.n2862 185
R16141 vdd.n2865 vdd.n929 185
R16142 vdd.n2945 vdd.n929 185
R16143 vdd.n2867 vdd.n2866 185
R16144 vdd.n2867 vdd.n928 185
R16145 vdd.n927 vdd.n926 185
R16146 vdd.n928 vdd.n927 185
R16147 vdd.n2947 vdd.n2946 185
R16148 vdd.n2946 vdd.n2945 185
R16149 vdd.n2948 vdd.n925 185
R16150 vdd.n2862 vdd.n925 185
R16151 vdd.n2950 vdd.n2949 185
R16152 vdd.n2951 vdd.n2950 185
R16153 vdd.n916 vdd.n915 185
R16154 vdd.n917 vdd.n916 185
R16155 vdd.n2959 vdd.n2958 185
R16156 vdd.n2958 vdd.n2957 185
R16157 vdd.n2960 vdd.n914 185
R16158 vdd.n914 vdd.n911 185
R16159 vdd.n2962 vdd.n2961 185
R16160 vdd.n2963 vdd.n2962 185
R16161 vdd.n904 vdd.n903 185
R16162 vdd.n905 vdd.n904 185
R16163 vdd.n2971 vdd.n2970 185
R16164 vdd.n2970 vdd.n2969 185
R16165 vdd.n2972 vdd.n902 185
R16166 vdd.n2847 vdd.n902 185
R16167 vdd.n2974 vdd.n2973 185
R16168 vdd.n2975 vdd.n2974 185
R16169 vdd.n892 vdd.n891 185
R16170 vdd.n901 vdd.n892 185
R16171 vdd.n2983 vdd.n2982 185
R16172 vdd.n2982 vdd.n2981 185
R16173 vdd.n2984 vdd.n890 185
R16174 vdd.n895 vdd.n890 185
R16175 vdd.n2986 vdd.n2985 185
R16176 vdd.n2987 vdd.n2986 185
R16177 vdd.n881 vdd.n880 185
R16178 vdd.n882 vdd.n881 185
R16179 vdd.n2995 vdd.n2994 185
R16180 vdd.n2994 vdd.n2993 185
R16181 vdd.n2996 vdd.n879 185
R16182 vdd.n879 vdd.n875 185
R16183 vdd.n2998 vdd.n2997 185
R16184 vdd.n2999 vdd.n2998 185
R16185 vdd.n867 vdd.n866 185
R16186 vdd.n878 vdd.n867 185
R16187 vdd.n3008 vdd.n3007 185
R16188 vdd.n3007 vdd.n3006 185
R16189 vdd.n3009 vdd.n865 185
R16190 vdd.n870 vdd.n865 185
R16191 vdd.n3011 vdd.n3010 185
R16192 vdd.n3012 vdd.n3011 185
R16193 vdd.n856 vdd.n855 185
R16194 vdd.n857 vdd.n856 185
R16195 vdd.n3020 vdd.n3019 185
R16196 vdd.n3019 vdd.n3018 185
R16197 vdd.n3021 vdd.n854 185
R16198 vdd.n854 vdd.n851 185
R16199 vdd.n3023 vdd.n3022 185
R16200 vdd.n3024 vdd.n3023 185
R16201 vdd.n842 vdd.n841 185
R16202 vdd.n843 vdd.n842 185
R16203 vdd.n3077 vdd.n3076 185
R16204 vdd.n3076 vdd.n3075 185
R16205 vdd.n3078 vdd.n840 185
R16206 vdd.n846 vdd.n840 185
R16207 vdd.n3080 vdd.n3079 185
R16208 vdd.n3081 vdd.n3080 185
R16209 vdd.n810 vdd.n808 185
R16210 vdd.n808 vdd.n805 185
R16211 vdd.n3150 vdd.n3149 185
R16212 vdd.n3151 vdd.n3150 185
R16213 vdd.n2592 vdd.n2591 185
R16214 vdd.n2593 vdd.n2592 185
R16215 vdd.n980 vdd.n978 185
R16216 vdd.n978 vdd.n976 185
R16217 vdd.n2507 vdd.n987 185
R16218 vdd.n2518 vdd.n987 185
R16219 vdd.n2508 vdd.n996 185
R16220 vdd.n1338 vdd.n996 185
R16221 vdd.n2510 vdd.n2509 185
R16222 vdd.n2511 vdd.n2510 185
R16223 vdd.n2506 vdd.n995 185
R16224 vdd.n995 vdd.n992 185
R16225 vdd.n2505 vdd.n2504 185
R16226 vdd.n2504 vdd.n2503 185
R16227 vdd.n998 vdd.n997 185
R16228 vdd.n999 vdd.n998 185
R16229 vdd.n2496 vdd.n2495 185
R16230 vdd.n2497 vdd.n2496 185
R16231 vdd.n2494 vdd.n1008 185
R16232 vdd.n1008 vdd.n1005 185
R16233 vdd.n2493 vdd.n2492 185
R16234 vdd.n2492 vdd.n2491 185
R16235 vdd.n1010 vdd.n1009 185
R16236 vdd.n1018 vdd.n1010 185
R16237 vdd.n2484 vdd.n2483 185
R16238 vdd.n2485 vdd.n2484 185
R16239 vdd.n2482 vdd.n1019 185
R16240 vdd.n1024 vdd.n1019 185
R16241 vdd.n2481 vdd.n2480 185
R16242 vdd.n2480 vdd.n2479 185
R16243 vdd.n1021 vdd.n1020 185
R16244 vdd.n1359 vdd.n1021 185
R16245 vdd.n2472 vdd.n2471 185
R16246 vdd.n2473 vdd.n2472 185
R16247 vdd.n2470 vdd.n1031 185
R16248 vdd.n1031 vdd.n1028 185
R16249 vdd.n2469 vdd.n2468 185
R16250 vdd.n2468 vdd.n2467 185
R16251 vdd.n1033 vdd.n1032 185
R16252 vdd.n1034 vdd.n1033 185
R16253 vdd.n2460 vdd.n2459 185
R16254 vdd.n2461 vdd.n2460 185
R16255 vdd.n2457 vdd.n1042 185
R16256 vdd.n1048 vdd.n1042 185
R16257 vdd.n2456 vdd.n2455 185
R16258 vdd.n2455 vdd.n2454 185
R16259 vdd.n1045 vdd.n1044 185
R16260 vdd.n1055 vdd.n1045 185
R16261 vdd.n2447 vdd.n2446 185
R16262 vdd.n2448 vdd.n2447 185
R16263 vdd.n2445 vdd.n1056 185
R16264 vdd.n1056 vdd.n1052 185
R16265 vdd.n2444 vdd.n2443 185
R16266 vdd.n2443 vdd.n2442 185
R16267 vdd.n1058 vdd.n1057 185
R16268 vdd.n1059 vdd.n1058 185
R16269 vdd.n2435 vdd.n2434 185
R16270 vdd.n2436 vdd.n2435 185
R16271 vdd.n2433 vdd.n1068 185
R16272 vdd.n1068 vdd.n1065 185
R16273 vdd.n2432 vdd.n2431 185
R16274 vdd.n2431 vdd.n2430 185
R16275 vdd.n1070 vdd.n1069 185
R16276 vdd.n1079 vdd.n1070 185
R16277 vdd.n2423 vdd.n2422 185
R16278 vdd.n2424 vdd.n2423 185
R16279 vdd.n2421 vdd.n1080 185
R16280 vdd.n1080 vdd.n1076 185
R16281 vdd.n2523 vdd.n951 185
R16282 vdd.n2665 vdd.n951 185
R16283 vdd.n2525 vdd.n2524 185
R16284 vdd.n2527 vdd.n2526 185
R16285 vdd.n2529 vdd.n2528 185
R16286 vdd.n2531 vdd.n2530 185
R16287 vdd.n2533 vdd.n2532 185
R16288 vdd.n2535 vdd.n2534 185
R16289 vdd.n2537 vdd.n2536 185
R16290 vdd.n2539 vdd.n2538 185
R16291 vdd.n2541 vdd.n2540 185
R16292 vdd.n2543 vdd.n2542 185
R16293 vdd.n2545 vdd.n2544 185
R16294 vdd.n2547 vdd.n2546 185
R16295 vdd.n2549 vdd.n2548 185
R16296 vdd.n2551 vdd.n2550 185
R16297 vdd.n2553 vdd.n2552 185
R16298 vdd.n2555 vdd.n2554 185
R16299 vdd.n2557 vdd.n2556 185
R16300 vdd.n2559 vdd.n2558 185
R16301 vdd.n2561 vdd.n2560 185
R16302 vdd.n2563 vdd.n2562 185
R16303 vdd.n2565 vdd.n2564 185
R16304 vdd.n2567 vdd.n2566 185
R16305 vdd.n2569 vdd.n2568 185
R16306 vdd.n2571 vdd.n2570 185
R16307 vdd.n2573 vdd.n2572 185
R16308 vdd.n2575 vdd.n2574 185
R16309 vdd.n2577 vdd.n2576 185
R16310 vdd.n2579 vdd.n2578 185
R16311 vdd.n2581 vdd.n2580 185
R16312 vdd.n2583 vdd.n2582 185
R16313 vdd.n2585 vdd.n2584 185
R16314 vdd.n2587 vdd.n2586 185
R16315 vdd.n2589 vdd.n2588 185
R16316 vdd.n2590 vdd.n979 185
R16317 vdd.n2522 vdd.n977 185
R16318 vdd.n2593 vdd.n977 185
R16319 vdd.n2521 vdd.n2520 185
R16320 vdd.n2520 vdd.n976 185
R16321 vdd.n2519 vdd.n984 185
R16322 vdd.n2519 vdd.n2518 185
R16323 vdd.n1256 vdd.n985 185
R16324 vdd.n1338 vdd.n985 185
R16325 vdd.n1257 vdd.n994 185
R16326 vdd.n2511 vdd.n994 185
R16327 vdd.n1259 vdd.n1258 185
R16328 vdd.n1258 vdd.n992 185
R16329 vdd.n1260 vdd.n1001 185
R16330 vdd.n2503 vdd.n1001 185
R16331 vdd.n1262 vdd.n1261 185
R16332 vdd.n1261 vdd.n999 185
R16333 vdd.n1263 vdd.n1007 185
R16334 vdd.n2497 vdd.n1007 185
R16335 vdd.n1265 vdd.n1264 185
R16336 vdd.n1264 vdd.n1005 185
R16337 vdd.n1266 vdd.n1012 185
R16338 vdd.n2491 vdd.n1012 185
R16339 vdd.n1268 vdd.n1267 185
R16340 vdd.n1267 vdd.n1018 185
R16341 vdd.n1269 vdd.n1017 185
R16342 vdd.n2485 vdd.n1017 185
R16343 vdd.n1271 vdd.n1270 185
R16344 vdd.n1270 vdd.n1024 185
R16345 vdd.n1272 vdd.n1023 185
R16346 vdd.n2479 vdd.n1023 185
R16347 vdd.n1361 vdd.n1360 185
R16348 vdd.n1360 vdd.n1359 185
R16349 vdd.n1362 vdd.n1030 185
R16350 vdd.n2473 vdd.n1030 185
R16351 vdd.n1364 vdd.n1363 185
R16352 vdd.n1363 vdd.n1028 185
R16353 vdd.n1365 vdd.n1036 185
R16354 vdd.n2467 vdd.n1036 185
R16355 vdd.n1367 vdd.n1366 185
R16356 vdd.n1366 vdd.n1034 185
R16357 vdd.n1368 vdd.n1041 185
R16358 vdd.n2461 vdd.n1041 185
R16359 vdd.n1370 vdd.n1369 185
R16360 vdd.n1369 vdd.n1048 185
R16361 vdd.n1371 vdd.n1047 185
R16362 vdd.n2454 vdd.n1047 185
R16363 vdd.n1373 vdd.n1372 185
R16364 vdd.n1372 vdd.n1055 185
R16365 vdd.n1374 vdd.n1054 185
R16366 vdd.n2448 vdd.n1054 185
R16367 vdd.n1376 vdd.n1375 185
R16368 vdd.n1375 vdd.n1052 185
R16369 vdd.n1377 vdd.n1061 185
R16370 vdd.n2442 vdd.n1061 185
R16371 vdd.n1379 vdd.n1378 185
R16372 vdd.n1378 vdd.n1059 185
R16373 vdd.n1380 vdd.n1067 185
R16374 vdd.n2436 vdd.n1067 185
R16375 vdd.n1382 vdd.n1381 185
R16376 vdd.n1381 vdd.n1065 185
R16377 vdd.n1383 vdd.n1072 185
R16378 vdd.n2430 vdd.n1072 185
R16379 vdd.n1385 vdd.n1384 185
R16380 vdd.n1384 vdd.n1079 185
R16381 vdd.n1386 vdd.n1078 185
R16382 vdd.n2424 vdd.n1078 185
R16383 vdd.n1388 vdd.n1387 185
R16384 vdd.n1387 vdd.n1076 185
R16385 vdd.n2420 vdd.n2419 185
R16386 vdd.n1082 vdd.n1081 185
R16387 vdd.n1223 vdd.n1222 185
R16388 vdd.n1225 vdd.n1224 185
R16389 vdd.n1227 vdd.n1226 185
R16390 vdd.n1229 vdd.n1228 185
R16391 vdd.n1231 vdd.n1230 185
R16392 vdd.n1233 vdd.n1232 185
R16393 vdd.n1235 vdd.n1234 185
R16394 vdd.n1237 vdd.n1236 185
R16395 vdd.n1239 vdd.n1238 185
R16396 vdd.n1241 vdd.n1240 185
R16397 vdd.n1243 vdd.n1242 185
R16398 vdd.n1245 vdd.n1244 185
R16399 vdd.n1247 vdd.n1246 185
R16400 vdd.n1249 vdd.n1248 185
R16401 vdd.n1251 vdd.n1250 185
R16402 vdd.n1422 vdd.n1252 185
R16403 vdd.n1421 vdd.n1420 185
R16404 vdd.n1419 vdd.n1418 185
R16405 vdd.n1417 vdd.n1416 185
R16406 vdd.n1415 vdd.n1414 185
R16407 vdd.n1413 vdd.n1412 185
R16408 vdd.n1411 vdd.n1410 185
R16409 vdd.n1409 vdd.n1408 185
R16410 vdd.n1407 vdd.n1406 185
R16411 vdd.n1405 vdd.n1404 185
R16412 vdd.n1403 vdd.n1402 185
R16413 vdd.n1401 vdd.n1400 185
R16414 vdd.n1399 vdd.n1398 185
R16415 vdd.n1397 vdd.n1396 185
R16416 vdd.n1395 vdd.n1394 185
R16417 vdd.n1393 vdd.n1392 185
R16418 vdd.n1391 vdd.n1390 185
R16419 vdd.n1389 vdd.n1116 185
R16420 vdd.n2417 vdd.n1116 185
R16421 vdd.n2417 vdd.n1083 179.345
R16422 vdd.n3315 vdd.n692 179.345
R16423 vdd.n327 vdd.n326 171.744
R16424 vdd.n326 vdd.n325 171.744
R16425 vdd.n325 vdd.n294 171.744
R16426 vdd.n318 vdd.n294 171.744
R16427 vdd.n318 vdd.n317 171.744
R16428 vdd.n317 vdd.n299 171.744
R16429 vdd.n310 vdd.n299 171.744
R16430 vdd.n310 vdd.n309 171.744
R16431 vdd.n309 vdd.n303 171.744
R16432 vdd.n268 vdd.n267 171.744
R16433 vdd.n267 vdd.n266 171.744
R16434 vdd.n266 vdd.n235 171.744
R16435 vdd.n259 vdd.n235 171.744
R16436 vdd.n259 vdd.n258 171.744
R16437 vdd.n258 vdd.n240 171.744
R16438 vdd.n251 vdd.n240 171.744
R16439 vdd.n251 vdd.n250 171.744
R16440 vdd.n250 vdd.n244 171.744
R16441 vdd.n225 vdd.n224 171.744
R16442 vdd.n224 vdd.n223 171.744
R16443 vdd.n223 vdd.n192 171.744
R16444 vdd.n216 vdd.n192 171.744
R16445 vdd.n216 vdd.n215 171.744
R16446 vdd.n215 vdd.n197 171.744
R16447 vdd.n208 vdd.n197 171.744
R16448 vdd.n208 vdd.n207 171.744
R16449 vdd.n207 vdd.n201 171.744
R16450 vdd.n166 vdd.n165 171.744
R16451 vdd.n165 vdd.n164 171.744
R16452 vdd.n164 vdd.n133 171.744
R16453 vdd.n157 vdd.n133 171.744
R16454 vdd.n157 vdd.n156 171.744
R16455 vdd.n156 vdd.n138 171.744
R16456 vdd.n149 vdd.n138 171.744
R16457 vdd.n149 vdd.n148 171.744
R16458 vdd.n148 vdd.n142 171.744
R16459 vdd.n124 vdd.n123 171.744
R16460 vdd.n123 vdd.n122 171.744
R16461 vdd.n122 vdd.n91 171.744
R16462 vdd.n115 vdd.n91 171.744
R16463 vdd.n115 vdd.n114 171.744
R16464 vdd.n114 vdd.n96 171.744
R16465 vdd.n107 vdd.n96 171.744
R16466 vdd.n107 vdd.n106 171.744
R16467 vdd.n106 vdd.n100 171.744
R16468 vdd.n65 vdd.n64 171.744
R16469 vdd.n64 vdd.n63 171.744
R16470 vdd.n63 vdd.n32 171.744
R16471 vdd.n56 vdd.n32 171.744
R16472 vdd.n56 vdd.n55 171.744
R16473 vdd.n55 vdd.n37 171.744
R16474 vdd.n48 vdd.n37 171.744
R16475 vdd.n48 vdd.n47 171.744
R16476 vdd.n47 vdd.n41 171.744
R16477 vdd.n2108 vdd.n2107 171.744
R16478 vdd.n2107 vdd.n2106 171.744
R16479 vdd.n2106 vdd.n2075 171.744
R16480 vdd.n2099 vdd.n2075 171.744
R16481 vdd.n2099 vdd.n2098 171.744
R16482 vdd.n2098 vdd.n2080 171.744
R16483 vdd.n2091 vdd.n2080 171.744
R16484 vdd.n2091 vdd.n2090 171.744
R16485 vdd.n2090 vdd.n2084 171.744
R16486 vdd.n2167 vdd.n2166 171.744
R16487 vdd.n2166 vdd.n2165 171.744
R16488 vdd.n2165 vdd.n2134 171.744
R16489 vdd.n2158 vdd.n2134 171.744
R16490 vdd.n2158 vdd.n2157 171.744
R16491 vdd.n2157 vdd.n2139 171.744
R16492 vdd.n2150 vdd.n2139 171.744
R16493 vdd.n2150 vdd.n2149 171.744
R16494 vdd.n2149 vdd.n2143 171.744
R16495 vdd.n2006 vdd.n2005 171.744
R16496 vdd.n2005 vdd.n2004 171.744
R16497 vdd.n2004 vdd.n1973 171.744
R16498 vdd.n1997 vdd.n1973 171.744
R16499 vdd.n1997 vdd.n1996 171.744
R16500 vdd.n1996 vdd.n1978 171.744
R16501 vdd.n1989 vdd.n1978 171.744
R16502 vdd.n1989 vdd.n1988 171.744
R16503 vdd.n1988 vdd.n1982 171.744
R16504 vdd.n2065 vdd.n2064 171.744
R16505 vdd.n2064 vdd.n2063 171.744
R16506 vdd.n2063 vdd.n2032 171.744
R16507 vdd.n2056 vdd.n2032 171.744
R16508 vdd.n2056 vdd.n2055 171.744
R16509 vdd.n2055 vdd.n2037 171.744
R16510 vdd.n2048 vdd.n2037 171.744
R16511 vdd.n2048 vdd.n2047 171.744
R16512 vdd.n2047 vdd.n2041 171.744
R16513 vdd.n1905 vdd.n1904 171.744
R16514 vdd.n1904 vdd.n1903 171.744
R16515 vdd.n1903 vdd.n1872 171.744
R16516 vdd.n1896 vdd.n1872 171.744
R16517 vdd.n1896 vdd.n1895 171.744
R16518 vdd.n1895 vdd.n1877 171.744
R16519 vdd.n1888 vdd.n1877 171.744
R16520 vdd.n1888 vdd.n1887 171.744
R16521 vdd.n1887 vdd.n1881 171.744
R16522 vdd.n1964 vdd.n1963 171.744
R16523 vdd.n1963 vdd.n1962 171.744
R16524 vdd.n1962 vdd.n1931 171.744
R16525 vdd.n1955 vdd.n1931 171.744
R16526 vdd.n1955 vdd.n1954 171.744
R16527 vdd.n1954 vdd.n1936 171.744
R16528 vdd.n1947 vdd.n1936 171.744
R16529 vdd.n1947 vdd.n1946 171.744
R16530 vdd.n1946 vdd.n1940 171.744
R16531 vdd.n468 vdd.n467 146.341
R16532 vdd.n474 vdd.n473 146.341
R16533 vdd.n478 vdd.n477 146.341
R16534 vdd.n484 vdd.n483 146.341
R16535 vdd.n488 vdd.n487 146.341
R16536 vdd.n494 vdd.n493 146.341
R16537 vdd.n498 vdd.n497 146.341
R16538 vdd.n504 vdd.n503 146.341
R16539 vdd.n508 vdd.n507 146.341
R16540 vdd.n514 vdd.n513 146.341
R16541 vdd.n518 vdd.n517 146.341
R16542 vdd.n524 vdd.n523 146.341
R16543 vdd.n528 vdd.n527 146.341
R16544 vdd.n534 vdd.n533 146.341
R16545 vdd.n538 vdd.n537 146.341
R16546 vdd.n544 vdd.n543 146.341
R16547 vdd.n548 vdd.n547 146.341
R16548 vdd.n554 vdd.n553 146.341
R16549 vdd.n558 vdd.n557 146.341
R16550 vdd.n564 vdd.n563 146.341
R16551 vdd.n568 vdd.n567 146.341
R16552 vdd.n574 vdd.n573 146.341
R16553 vdd.n578 vdd.n577 146.341
R16554 vdd.n584 vdd.n583 146.341
R16555 vdd.n588 vdd.n587 146.341
R16556 vdd.n594 vdd.n593 146.341
R16557 vdd.n598 vdd.n597 146.341
R16558 vdd.n604 vdd.n603 146.341
R16559 vdd.n608 vdd.n607 146.341
R16560 vdd.n614 vdd.n613 146.341
R16561 vdd.n616 vdd.n425 146.341
R16562 vdd.n3322 vdd.n685 146.341
R16563 vdd.n3322 vdd.n677 146.341
R16564 vdd.n3332 vdd.n677 146.341
R16565 vdd.n3332 vdd.n673 146.341
R16566 vdd.n3338 vdd.n673 146.341
R16567 vdd.n3338 vdd.n667 146.341
R16568 vdd.n3349 vdd.n667 146.341
R16569 vdd.n3349 vdd.n663 146.341
R16570 vdd.n3355 vdd.n663 146.341
R16571 vdd.n3355 vdd.n654 146.341
R16572 vdd.n3365 vdd.n654 146.341
R16573 vdd.n3365 vdd.n650 146.341
R16574 vdd.n3371 vdd.n650 146.341
R16575 vdd.n3371 vdd.n643 146.341
R16576 vdd.n3382 vdd.n643 146.341
R16577 vdd.n3382 vdd.n639 146.341
R16578 vdd.n3391 vdd.n639 146.341
R16579 vdd.n3391 vdd.n632 146.341
R16580 vdd.n3401 vdd.n632 146.341
R16581 vdd.n3402 vdd.n3401 146.341
R16582 vdd.n3402 vdd.n341 146.341
R16583 vdd.n342 vdd.n341 146.341
R16584 vdd.n343 vdd.n342 146.341
R16585 vdd.n3409 vdd.n343 146.341
R16586 vdd.n3409 vdd.n351 146.341
R16587 vdd.n352 vdd.n351 146.341
R16588 vdd.n353 vdd.n352 146.341
R16589 vdd.n3416 vdd.n353 146.341
R16590 vdd.n3416 vdd.n362 146.341
R16591 vdd.n363 vdd.n362 146.341
R16592 vdd.n364 vdd.n363 146.341
R16593 vdd.n3424 vdd.n364 146.341
R16594 vdd.n3424 vdd.n372 146.341
R16595 vdd.n373 vdd.n372 146.341
R16596 vdd.n374 vdd.n373 146.341
R16597 vdd.n3431 vdd.n374 146.341
R16598 vdd.n3431 vdd.n383 146.341
R16599 vdd.n384 vdd.n383 146.341
R16600 vdd.n385 vdd.n384 146.341
R16601 vdd.n3438 vdd.n385 146.341
R16602 vdd.n3438 vdd.n393 146.341
R16603 vdd.n725 vdd.n724 146.341
R16604 vdd.n728 vdd.n724 146.341
R16605 vdd.n734 vdd.n733 146.341
R16606 vdd.n3304 vdd.n3303 146.341
R16607 vdd.n3300 vdd.n3299 146.341
R16608 vdd.n3296 vdd.n3295 146.341
R16609 vdd.n3292 vdd.n3291 146.341
R16610 vdd.n3288 vdd.n3287 146.341
R16611 vdd.n3284 vdd.n3283 146.341
R16612 vdd.n3280 vdd.n3279 146.341
R16613 vdd.n3271 vdd.n3270 146.341
R16614 vdd.n3268 vdd.n3267 146.341
R16615 vdd.n3264 vdd.n3263 146.341
R16616 vdd.n3260 vdd.n3259 146.341
R16617 vdd.n3256 vdd.n3255 146.341
R16618 vdd.n3252 vdd.n3251 146.341
R16619 vdd.n3248 vdd.n3247 146.341
R16620 vdd.n3244 vdd.n3243 146.341
R16621 vdd.n3240 vdd.n3239 146.341
R16622 vdd.n3236 vdd.n3235 146.341
R16623 vdd.n3232 vdd.n3231 146.341
R16624 vdd.n3225 vdd.n3224 146.341
R16625 vdd.n3222 vdd.n3221 146.341
R16626 vdd.n3218 vdd.n3217 146.341
R16627 vdd.n3214 vdd.n3213 146.341
R16628 vdd.n3210 vdd.n3209 146.341
R16629 vdd.n3206 vdd.n3205 146.341
R16630 vdd.n3202 vdd.n3201 146.341
R16631 vdd.n3198 vdd.n3197 146.341
R16632 vdd.n3194 vdd.n3193 146.341
R16633 vdd.n3190 vdd.n3189 146.341
R16634 vdd.n3316 vdd.n691 146.341
R16635 vdd.n3324 vdd.n684 146.341
R16636 vdd.n3324 vdd.n680 146.341
R16637 vdd.n3330 vdd.n680 146.341
R16638 vdd.n3330 vdd.n672 146.341
R16639 vdd.n3341 vdd.n672 146.341
R16640 vdd.n3341 vdd.n668 146.341
R16641 vdd.n3347 vdd.n668 146.341
R16642 vdd.n3347 vdd.n661 146.341
R16643 vdd.n3357 vdd.n661 146.341
R16644 vdd.n3357 vdd.n657 146.341
R16645 vdd.n3363 vdd.n657 146.341
R16646 vdd.n3363 vdd.n649 146.341
R16647 vdd.n3374 vdd.n649 146.341
R16648 vdd.n3374 vdd.n645 146.341
R16649 vdd.n3380 vdd.n645 146.341
R16650 vdd.n3380 vdd.n638 146.341
R16651 vdd.n3393 vdd.n638 146.341
R16652 vdd.n3393 vdd.n634 146.341
R16653 vdd.n3399 vdd.n634 146.341
R16654 vdd.n3399 vdd.n338 146.341
R16655 vdd.n3488 vdd.n338 146.341
R16656 vdd.n3488 vdd.n339 146.341
R16657 vdd.n3484 vdd.n339 146.341
R16658 vdd.n3484 vdd.n345 146.341
R16659 vdd.n3480 vdd.n345 146.341
R16660 vdd.n3480 vdd.n350 146.341
R16661 vdd.n3476 vdd.n350 146.341
R16662 vdd.n3476 vdd.n354 146.341
R16663 vdd.n3472 vdd.n354 146.341
R16664 vdd.n3472 vdd.n360 146.341
R16665 vdd.n3468 vdd.n360 146.341
R16666 vdd.n3468 vdd.n365 146.341
R16667 vdd.n3464 vdd.n365 146.341
R16668 vdd.n3464 vdd.n371 146.341
R16669 vdd.n3460 vdd.n371 146.341
R16670 vdd.n3460 vdd.n376 146.341
R16671 vdd.n3456 vdd.n376 146.341
R16672 vdd.n3456 vdd.n382 146.341
R16673 vdd.n3452 vdd.n382 146.341
R16674 vdd.n3452 vdd.n387 146.341
R16675 vdd.n3448 vdd.n387 146.341
R16676 vdd.n2378 vdd.n2377 146.341
R16677 vdd.n2375 vdd.n2372 146.341
R16678 vdd.n2370 vdd.n1127 146.341
R16679 vdd.n2366 vdd.n2365 146.341
R16680 vdd.n2363 vdd.n1131 146.341
R16681 vdd.n2359 vdd.n2358 146.341
R16682 vdd.n2356 vdd.n1138 146.341
R16683 vdd.n2352 vdd.n2351 146.341
R16684 vdd.n2349 vdd.n1145 146.341
R16685 vdd.n1156 vdd.n1153 146.341
R16686 vdd.n2341 vdd.n2340 146.341
R16687 vdd.n2338 vdd.n1158 146.341
R16688 vdd.n2334 vdd.n2333 146.341
R16689 vdd.n2331 vdd.n1164 146.341
R16690 vdd.n2327 vdd.n2326 146.341
R16691 vdd.n2324 vdd.n1171 146.341
R16692 vdd.n2320 vdd.n2319 146.341
R16693 vdd.n2317 vdd.n1178 146.341
R16694 vdd.n2313 vdd.n2312 146.341
R16695 vdd.n2310 vdd.n1185 146.341
R16696 vdd.n1196 vdd.n1193 146.341
R16697 vdd.n2302 vdd.n2301 146.341
R16698 vdd.n2299 vdd.n1198 146.341
R16699 vdd.n2295 vdd.n2294 146.341
R16700 vdd.n2292 vdd.n1204 146.341
R16701 vdd.n2288 vdd.n2287 146.341
R16702 vdd.n2285 vdd.n1211 146.341
R16703 vdd.n2281 vdd.n2280 146.341
R16704 vdd.n2278 vdd.n1218 146.341
R16705 vdd.n1429 vdd.n1427 146.341
R16706 vdd.n1432 vdd.n1431 146.341
R16707 vdd.n1790 vdd.n1550 146.341
R16708 vdd.n1790 vdd.n1546 146.341
R16709 vdd.n1796 vdd.n1546 146.341
R16710 vdd.n1796 vdd.n1538 146.341
R16711 vdd.n1807 vdd.n1538 146.341
R16712 vdd.n1807 vdd.n1534 146.341
R16713 vdd.n1813 vdd.n1534 146.341
R16714 vdd.n1813 vdd.n1528 146.341
R16715 vdd.n1824 vdd.n1528 146.341
R16716 vdd.n1824 vdd.n1524 146.341
R16717 vdd.n1830 vdd.n1524 146.341
R16718 vdd.n1830 vdd.n1515 146.341
R16719 vdd.n1840 vdd.n1515 146.341
R16720 vdd.n1840 vdd.n1511 146.341
R16721 vdd.n1846 vdd.n1511 146.341
R16722 vdd.n1846 vdd.n1504 146.341
R16723 vdd.n1857 vdd.n1504 146.341
R16724 vdd.n1857 vdd.n1500 146.341
R16725 vdd.n1863 vdd.n1500 146.341
R16726 vdd.n1863 vdd.n1493 146.341
R16727 vdd.n2180 vdd.n1493 146.341
R16728 vdd.n2180 vdd.n1489 146.341
R16729 vdd.n2186 vdd.n1489 146.341
R16730 vdd.n2186 vdd.n1481 146.341
R16731 vdd.n2197 vdd.n1481 146.341
R16732 vdd.n2197 vdd.n1477 146.341
R16733 vdd.n2203 vdd.n1477 146.341
R16734 vdd.n2203 vdd.n1471 146.341
R16735 vdd.n2214 vdd.n1471 146.341
R16736 vdd.n2214 vdd.n1467 146.341
R16737 vdd.n2220 vdd.n1467 146.341
R16738 vdd.n2220 vdd.n1458 146.341
R16739 vdd.n2230 vdd.n1458 146.341
R16740 vdd.n2230 vdd.n1454 146.341
R16741 vdd.n2236 vdd.n1454 146.341
R16742 vdd.n2236 vdd.n1448 146.341
R16743 vdd.n2247 vdd.n1448 146.341
R16744 vdd.n2247 vdd.n1443 146.341
R16745 vdd.n2255 vdd.n1443 146.341
R16746 vdd.n2255 vdd.n1434 146.341
R16747 vdd.n2266 vdd.n1434 146.341
R16748 vdd.n1779 vdd.n1555 146.341
R16749 vdd.n1779 vdd.n1588 146.341
R16750 vdd.n1592 vdd.n1591 146.341
R16751 vdd.n1594 vdd.n1593 146.341
R16752 vdd.n1598 vdd.n1597 146.341
R16753 vdd.n1600 vdd.n1599 146.341
R16754 vdd.n1604 vdd.n1603 146.341
R16755 vdd.n1606 vdd.n1605 146.341
R16756 vdd.n1610 vdd.n1609 146.341
R16757 vdd.n1612 vdd.n1611 146.341
R16758 vdd.n1618 vdd.n1617 146.341
R16759 vdd.n1620 vdd.n1619 146.341
R16760 vdd.n1624 vdd.n1623 146.341
R16761 vdd.n1626 vdd.n1625 146.341
R16762 vdd.n1630 vdd.n1629 146.341
R16763 vdd.n1632 vdd.n1631 146.341
R16764 vdd.n1636 vdd.n1635 146.341
R16765 vdd.n1638 vdd.n1637 146.341
R16766 vdd.n1642 vdd.n1641 146.341
R16767 vdd.n1644 vdd.n1643 146.341
R16768 vdd.n1716 vdd.n1647 146.341
R16769 vdd.n1649 vdd.n1648 146.341
R16770 vdd.n1653 vdd.n1652 146.341
R16771 vdd.n1655 vdd.n1654 146.341
R16772 vdd.n1659 vdd.n1658 146.341
R16773 vdd.n1661 vdd.n1660 146.341
R16774 vdd.n1665 vdd.n1664 146.341
R16775 vdd.n1667 vdd.n1666 146.341
R16776 vdd.n1671 vdd.n1670 146.341
R16777 vdd.n1673 vdd.n1672 146.341
R16778 vdd.n1677 vdd.n1676 146.341
R16779 vdd.n1678 vdd.n1586 146.341
R16780 vdd.n1788 vdd.n1551 146.341
R16781 vdd.n1788 vdd.n1544 146.341
R16782 vdd.n1799 vdd.n1544 146.341
R16783 vdd.n1799 vdd.n1540 146.341
R16784 vdd.n1805 vdd.n1540 146.341
R16785 vdd.n1805 vdd.n1533 146.341
R16786 vdd.n1816 vdd.n1533 146.341
R16787 vdd.n1816 vdd.n1529 146.341
R16788 vdd.n1822 vdd.n1529 146.341
R16789 vdd.n1822 vdd.n1522 146.341
R16790 vdd.n1832 vdd.n1522 146.341
R16791 vdd.n1832 vdd.n1518 146.341
R16792 vdd.n1838 vdd.n1518 146.341
R16793 vdd.n1838 vdd.n1510 146.341
R16794 vdd.n1849 vdd.n1510 146.341
R16795 vdd.n1849 vdd.n1506 146.341
R16796 vdd.n1855 vdd.n1506 146.341
R16797 vdd.n1855 vdd.n1499 146.341
R16798 vdd.n1865 vdd.n1499 146.341
R16799 vdd.n1865 vdd.n1495 146.341
R16800 vdd.n2178 vdd.n1495 146.341
R16801 vdd.n2178 vdd.n1487 146.341
R16802 vdd.n2189 vdd.n1487 146.341
R16803 vdd.n2189 vdd.n1483 146.341
R16804 vdd.n2195 vdd.n1483 146.341
R16805 vdd.n2195 vdd.n1476 146.341
R16806 vdd.n2206 vdd.n1476 146.341
R16807 vdd.n2206 vdd.n1472 146.341
R16808 vdd.n2212 vdd.n1472 146.341
R16809 vdd.n2212 vdd.n1465 146.341
R16810 vdd.n2222 vdd.n1465 146.341
R16811 vdd.n2222 vdd.n1461 146.341
R16812 vdd.n2228 vdd.n1461 146.341
R16813 vdd.n2228 vdd.n1453 146.341
R16814 vdd.n2239 vdd.n1453 146.341
R16815 vdd.n2239 vdd.n1449 146.341
R16816 vdd.n2245 vdd.n1449 146.341
R16817 vdd.n2245 vdd.n1441 146.341
R16818 vdd.n2258 vdd.n1441 146.341
R16819 vdd.n2258 vdd.n1436 146.341
R16820 vdd.n2264 vdd.n1436 146.341
R16821 vdd.n1253 vdd.t224 127.284
R16822 vdd.n981 vdd.t265 127.284
R16823 vdd.n1273 vdd.t238 127.284
R16824 vdd.n972 vdd.t288 127.284
R16825 vdd.n872 vdd.t245 127.284
R16826 vdd.n872 vdd.t246 127.284
R16827 vdd.n2704 vdd.t283 127.284
R16828 vdd.n832 vdd.t291 127.284
R16829 vdd.n2701 vdd.t270 127.284
R16830 vdd.n799 vdd.t219 127.284
R16831 vdd.n1043 vdd.t276 127.284
R16832 vdd.n1043 vdd.t277 127.284
R16833 vdd.n22 vdd.n20 117.314
R16834 vdd.n17 vdd.n15 117.314
R16835 vdd.n27 vdd.n26 116.927
R16836 vdd.n24 vdd.n23 116.927
R16837 vdd.n22 vdd.n21 116.927
R16838 vdd.n17 vdd.n16 116.927
R16839 vdd.n19 vdd.n18 116.927
R16840 vdd.n27 vdd.n25 116.927
R16841 vdd.n1254 vdd.t223 111.188
R16842 vdd.n982 vdd.t266 111.188
R16843 vdd.n1274 vdd.t237 111.188
R16844 vdd.n973 vdd.t289 111.188
R16845 vdd.n2705 vdd.t282 111.188
R16846 vdd.n833 vdd.t292 111.188
R16847 vdd.n2702 vdd.t269 111.188
R16848 vdd.n800 vdd.t220 111.188
R16849 vdd.n2946 vdd.n927 99.5127
R16850 vdd.n2946 vdd.n925 99.5127
R16851 vdd.n2950 vdd.n925 99.5127
R16852 vdd.n2950 vdd.n916 99.5127
R16853 vdd.n2958 vdd.n916 99.5127
R16854 vdd.n2958 vdd.n914 99.5127
R16855 vdd.n2962 vdd.n914 99.5127
R16856 vdd.n2962 vdd.n904 99.5127
R16857 vdd.n2970 vdd.n904 99.5127
R16858 vdd.n2970 vdd.n902 99.5127
R16859 vdd.n2974 vdd.n902 99.5127
R16860 vdd.n2974 vdd.n892 99.5127
R16861 vdd.n2982 vdd.n892 99.5127
R16862 vdd.n2982 vdd.n890 99.5127
R16863 vdd.n2986 vdd.n890 99.5127
R16864 vdd.n2986 vdd.n881 99.5127
R16865 vdd.n2994 vdd.n881 99.5127
R16866 vdd.n2994 vdd.n879 99.5127
R16867 vdd.n2998 vdd.n879 99.5127
R16868 vdd.n2998 vdd.n867 99.5127
R16869 vdd.n3007 vdd.n867 99.5127
R16870 vdd.n3007 vdd.n865 99.5127
R16871 vdd.n3011 vdd.n865 99.5127
R16872 vdd.n3011 vdd.n856 99.5127
R16873 vdd.n3019 vdd.n856 99.5127
R16874 vdd.n3019 vdd.n854 99.5127
R16875 vdd.n3023 vdd.n854 99.5127
R16876 vdd.n3023 vdd.n842 99.5127
R16877 vdd.n3076 vdd.n842 99.5127
R16878 vdd.n3076 vdd.n840 99.5127
R16879 vdd.n3080 vdd.n840 99.5127
R16880 vdd.n3080 vdd.n808 99.5127
R16881 vdd.n3150 vdd.n808 99.5127
R16882 vdd.n3146 vdd.n809 99.5127
R16883 vdd.n3144 vdd.n3143 99.5127
R16884 vdd.n3141 vdd.n813 99.5127
R16885 vdd.n3137 vdd.n3136 99.5127
R16886 vdd.n3134 vdd.n816 99.5127
R16887 vdd.n3130 vdd.n3129 99.5127
R16888 vdd.n3127 vdd.n819 99.5127
R16889 vdd.n3123 vdd.n3122 99.5127
R16890 vdd.n3120 vdd.n3118 99.5127
R16891 vdd.n3116 vdd.n822 99.5127
R16892 vdd.n3112 vdd.n3111 99.5127
R16893 vdd.n3109 vdd.n825 99.5127
R16894 vdd.n3105 vdd.n3104 99.5127
R16895 vdd.n3102 vdd.n828 99.5127
R16896 vdd.n3098 vdd.n3097 99.5127
R16897 vdd.n3095 vdd.n831 99.5127
R16898 vdd.n3090 vdd.n3089 99.5127
R16899 vdd.n2867 vdd.n929 99.5127
R16900 vdd.n2863 vdd.n929 99.5127
R16901 vdd.n2863 vdd.n923 99.5127
R16902 vdd.n2807 vdd.n923 99.5127
R16903 vdd.n2807 vdd.n918 99.5127
R16904 vdd.n2810 vdd.n918 99.5127
R16905 vdd.n2810 vdd.n912 99.5127
R16906 vdd.n2813 vdd.n912 99.5127
R16907 vdd.n2813 vdd.n906 99.5127
R16908 vdd.n2846 vdd.n906 99.5127
R16909 vdd.n2846 vdd.n899 99.5127
R16910 vdd.n2842 vdd.n899 99.5127
R16911 vdd.n2842 vdd.n893 99.5127
R16912 vdd.n2839 vdd.n893 99.5127
R16913 vdd.n2839 vdd.n888 99.5127
R16914 vdd.n2836 vdd.n888 99.5127
R16915 vdd.n2836 vdd.n883 99.5127
R16916 vdd.n2833 vdd.n883 99.5127
R16917 vdd.n2833 vdd.n876 99.5127
R16918 vdd.n2830 vdd.n876 99.5127
R16919 vdd.n2830 vdd.n868 99.5127
R16920 vdd.n2827 vdd.n868 99.5127
R16921 vdd.n2827 vdd.n863 99.5127
R16922 vdd.n2824 vdd.n863 99.5127
R16923 vdd.n2824 vdd.n858 99.5127
R16924 vdd.n2821 vdd.n858 99.5127
R16925 vdd.n2821 vdd.n852 99.5127
R16926 vdd.n2818 vdd.n852 99.5127
R16927 vdd.n2818 vdd.n844 99.5127
R16928 vdd.n844 vdd.n837 99.5127
R16929 vdd.n3082 vdd.n837 99.5127
R16930 vdd.n3083 vdd.n3082 99.5127
R16931 vdd.n3083 vdd.n806 99.5127
R16932 vdd.n2700 vdd.n2699 99.5127
R16933 vdd.n2931 vdd.n2699 99.5127
R16934 vdd.n2929 vdd.n2928 99.5127
R16935 vdd.n2925 vdd.n2924 99.5127
R16936 vdd.n2921 vdd.n2920 99.5127
R16937 vdd.n2917 vdd.n2916 99.5127
R16938 vdd.n2913 vdd.n2912 99.5127
R16939 vdd.n2909 vdd.n2908 99.5127
R16940 vdd.n2905 vdd.n2904 99.5127
R16941 vdd.n2901 vdd.n2900 99.5127
R16942 vdd.n2897 vdd.n2896 99.5127
R16943 vdd.n2893 vdd.n2892 99.5127
R16944 vdd.n2889 vdd.n2888 99.5127
R16945 vdd.n2885 vdd.n2884 99.5127
R16946 vdd.n2881 vdd.n2880 99.5127
R16947 vdd.n2877 vdd.n2876 99.5127
R16948 vdd.n2872 vdd.n2871 99.5127
R16949 vdd.n2664 vdd.n970 99.5127
R16950 vdd.n2660 vdd.n2659 99.5127
R16951 vdd.n2656 vdd.n2655 99.5127
R16952 vdd.n2652 vdd.n2651 99.5127
R16953 vdd.n2648 vdd.n2647 99.5127
R16954 vdd.n2644 vdd.n2643 99.5127
R16955 vdd.n2640 vdd.n2639 99.5127
R16956 vdd.n2636 vdd.n2635 99.5127
R16957 vdd.n2632 vdd.n2631 99.5127
R16958 vdd.n2628 vdd.n2627 99.5127
R16959 vdd.n2624 vdd.n2623 99.5127
R16960 vdd.n2620 vdd.n2619 99.5127
R16961 vdd.n2616 vdd.n2615 99.5127
R16962 vdd.n2612 vdd.n2611 99.5127
R16963 vdd.n2608 vdd.n2607 99.5127
R16964 vdd.n2604 vdd.n2603 99.5127
R16965 vdd.n2599 vdd.n2598 99.5127
R16966 vdd.n1309 vdd.n1077 99.5127
R16967 vdd.n1312 vdd.n1077 99.5127
R16968 vdd.n1312 vdd.n1071 99.5127
R16969 vdd.n1315 vdd.n1071 99.5127
R16970 vdd.n1315 vdd.n1066 99.5127
R16971 vdd.n1318 vdd.n1066 99.5127
R16972 vdd.n1318 vdd.n1060 99.5127
R16973 vdd.n1321 vdd.n1060 99.5127
R16974 vdd.n1321 vdd.n1053 99.5127
R16975 vdd.n1324 vdd.n1053 99.5127
R16976 vdd.n1324 vdd.n1046 99.5127
R16977 vdd.n1327 vdd.n1046 99.5127
R16978 vdd.n1327 vdd.n1040 99.5127
R16979 vdd.n1330 vdd.n1040 99.5127
R16980 vdd.n1330 vdd.n1035 99.5127
R16981 vdd.n1333 vdd.n1035 99.5127
R16982 vdd.n1333 vdd.n1029 99.5127
R16983 vdd.n1358 vdd.n1029 99.5127
R16984 vdd.n1358 vdd.n1022 99.5127
R16985 vdd.n1354 vdd.n1022 99.5127
R16986 vdd.n1354 vdd.n1016 99.5127
R16987 vdd.n1351 vdd.n1016 99.5127
R16988 vdd.n1351 vdd.n1011 99.5127
R16989 vdd.n1348 vdd.n1011 99.5127
R16990 vdd.n1348 vdd.n1006 99.5127
R16991 vdd.n1345 vdd.n1006 99.5127
R16992 vdd.n1345 vdd.n1000 99.5127
R16993 vdd.n1342 vdd.n1000 99.5127
R16994 vdd.n1342 vdd.n993 99.5127
R16995 vdd.n1339 vdd.n993 99.5127
R16996 vdd.n1339 vdd.n986 99.5127
R16997 vdd.n986 vdd.n975 99.5127
R16998 vdd.n2594 vdd.n975 99.5127
R16999 vdd.n1118 vdd.n1117 99.5127
R17000 vdd.n2410 vdd.n1117 99.5127
R17001 vdd.n2408 vdd.n2407 99.5127
R17002 vdd.n2404 vdd.n2403 99.5127
R17003 vdd.n2400 vdd.n2399 99.5127
R17004 vdd.n2396 vdd.n2395 99.5127
R17005 vdd.n2392 vdd.n2391 99.5127
R17006 vdd.n2388 vdd.n2387 99.5127
R17007 vdd.n2384 vdd.n2383 99.5127
R17008 vdd.n1276 vdd.n1275 99.5127
R17009 vdd.n1280 vdd.n1279 99.5127
R17010 vdd.n1284 vdd.n1283 99.5127
R17011 vdd.n1288 vdd.n1287 99.5127
R17012 vdd.n1292 vdd.n1291 99.5127
R17013 vdd.n1296 vdd.n1295 99.5127
R17014 vdd.n1300 vdd.n1299 99.5127
R17015 vdd.n1305 vdd.n1304 99.5127
R17016 vdd.n2425 vdd.n1075 99.5127
R17017 vdd.n2425 vdd.n1073 99.5127
R17018 vdd.n2429 vdd.n1073 99.5127
R17019 vdd.n2429 vdd.n1064 99.5127
R17020 vdd.n2437 vdd.n1064 99.5127
R17021 vdd.n2437 vdd.n1062 99.5127
R17022 vdd.n2441 vdd.n1062 99.5127
R17023 vdd.n2441 vdd.n1051 99.5127
R17024 vdd.n2449 vdd.n1051 99.5127
R17025 vdd.n2449 vdd.n1049 99.5127
R17026 vdd.n2453 vdd.n1049 99.5127
R17027 vdd.n2453 vdd.n1039 99.5127
R17028 vdd.n2462 vdd.n1039 99.5127
R17029 vdd.n2462 vdd.n1037 99.5127
R17030 vdd.n2466 vdd.n1037 99.5127
R17031 vdd.n2466 vdd.n1027 99.5127
R17032 vdd.n2474 vdd.n1027 99.5127
R17033 vdd.n2474 vdd.n1025 99.5127
R17034 vdd.n2478 vdd.n1025 99.5127
R17035 vdd.n2478 vdd.n1015 99.5127
R17036 vdd.n2486 vdd.n1015 99.5127
R17037 vdd.n2486 vdd.n1013 99.5127
R17038 vdd.n2490 vdd.n1013 99.5127
R17039 vdd.n2490 vdd.n1004 99.5127
R17040 vdd.n2498 vdd.n1004 99.5127
R17041 vdd.n2498 vdd.n1002 99.5127
R17042 vdd.n2502 vdd.n1002 99.5127
R17043 vdd.n2502 vdd.n991 99.5127
R17044 vdd.n2512 vdd.n991 99.5127
R17045 vdd.n2512 vdd.n988 99.5127
R17046 vdd.n2517 vdd.n988 99.5127
R17047 vdd.n2517 vdd.n989 99.5127
R17048 vdd.n989 vdd.n969 99.5127
R17049 vdd.n3066 vdd.n3065 99.5127
R17050 vdd.n3063 vdd.n3029 99.5127
R17051 vdd.n3059 vdd.n3058 99.5127
R17052 vdd.n3056 vdd.n3032 99.5127
R17053 vdd.n3052 vdd.n3051 99.5127
R17054 vdd.n3049 vdd.n3035 99.5127
R17055 vdd.n3045 vdd.n3044 99.5127
R17056 vdd.n3042 vdd.n3039 99.5127
R17057 vdd.n3183 vdd.n787 99.5127
R17058 vdd.n3181 vdd.n3180 99.5127
R17059 vdd.n3178 vdd.n789 99.5127
R17060 vdd.n3174 vdd.n3173 99.5127
R17061 vdd.n3171 vdd.n792 99.5127
R17062 vdd.n3167 vdd.n3166 99.5127
R17063 vdd.n3164 vdd.n795 99.5127
R17064 vdd.n3160 vdd.n3159 99.5127
R17065 vdd.n3157 vdd.n798 99.5127
R17066 vdd.n2772 vdd.n930 99.5127
R17067 vdd.n2861 vdd.n930 99.5127
R17068 vdd.n2861 vdd.n924 99.5127
R17069 vdd.n2857 vdd.n924 99.5127
R17070 vdd.n2857 vdd.n919 99.5127
R17071 vdd.n2854 vdd.n919 99.5127
R17072 vdd.n2854 vdd.n913 99.5127
R17073 vdd.n2851 vdd.n913 99.5127
R17074 vdd.n2851 vdd.n907 99.5127
R17075 vdd.n2848 vdd.n907 99.5127
R17076 vdd.n2848 vdd.n900 99.5127
R17077 vdd.n2804 vdd.n900 99.5127
R17078 vdd.n2804 vdd.n894 99.5127
R17079 vdd.n2801 vdd.n894 99.5127
R17080 vdd.n2801 vdd.n889 99.5127
R17081 vdd.n2798 vdd.n889 99.5127
R17082 vdd.n2798 vdd.n884 99.5127
R17083 vdd.n2795 vdd.n884 99.5127
R17084 vdd.n2795 vdd.n877 99.5127
R17085 vdd.n2792 vdd.n877 99.5127
R17086 vdd.n2792 vdd.n869 99.5127
R17087 vdd.n2789 vdd.n869 99.5127
R17088 vdd.n2789 vdd.n864 99.5127
R17089 vdd.n2786 vdd.n864 99.5127
R17090 vdd.n2786 vdd.n859 99.5127
R17091 vdd.n2783 vdd.n859 99.5127
R17092 vdd.n2783 vdd.n853 99.5127
R17093 vdd.n2780 vdd.n853 99.5127
R17094 vdd.n2780 vdd.n845 99.5127
R17095 vdd.n2777 vdd.n845 99.5127
R17096 vdd.n2777 vdd.n838 99.5127
R17097 vdd.n838 vdd.n804 99.5127
R17098 vdd.n3152 vdd.n804 99.5127
R17099 vdd.n2707 vdd.n933 99.5127
R17100 vdd.n2711 vdd.n2710 99.5127
R17101 vdd.n2715 vdd.n2714 99.5127
R17102 vdd.n2719 vdd.n2718 99.5127
R17103 vdd.n2723 vdd.n2722 99.5127
R17104 vdd.n2727 vdd.n2726 99.5127
R17105 vdd.n2731 vdd.n2730 99.5127
R17106 vdd.n2735 vdd.n2734 99.5127
R17107 vdd.n2739 vdd.n2738 99.5127
R17108 vdd.n2743 vdd.n2742 99.5127
R17109 vdd.n2747 vdd.n2746 99.5127
R17110 vdd.n2751 vdd.n2750 99.5127
R17111 vdd.n2755 vdd.n2754 99.5127
R17112 vdd.n2759 vdd.n2758 99.5127
R17113 vdd.n2763 vdd.n2762 99.5127
R17114 vdd.n2767 vdd.n2766 99.5127
R17115 vdd.n2769 vdd.n2698 99.5127
R17116 vdd.n2944 vdd.n931 99.5127
R17117 vdd.n2944 vdd.n922 99.5127
R17118 vdd.n2952 vdd.n922 99.5127
R17119 vdd.n2952 vdd.n920 99.5127
R17120 vdd.n2956 vdd.n920 99.5127
R17121 vdd.n2956 vdd.n910 99.5127
R17122 vdd.n2964 vdd.n910 99.5127
R17123 vdd.n2964 vdd.n908 99.5127
R17124 vdd.n2968 vdd.n908 99.5127
R17125 vdd.n2968 vdd.n898 99.5127
R17126 vdd.n2976 vdd.n898 99.5127
R17127 vdd.n2976 vdd.n896 99.5127
R17128 vdd.n2980 vdd.n896 99.5127
R17129 vdd.n2980 vdd.n887 99.5127
R17130 vdd.n2988 vdd.n887 99.5127
R17131 vdd.n2988 vdd.n885 99.5127
R17132 vdd.n2992 vdd.n885 99.5127
R17133 vdd.n2992 vdd.n874 99.5127
R17134 vdd.n3000 vdd.n874 99.5127
R17135 vdd.n3000 vdd.n871 99.5127
R17136 vdd.n3005 vdd.n871 99.5127
R17137 vdd.n3005 vdd.n862 99.5127
R17138 vdd.n3013 vdd.n862 99.5127
R17139 vdd.n3013 vdd.n860 99.5127
R17140 vdd.n3017 vdd.n860 99.5127
R17141 vdd.n3017 vdd.n850 99.5127
R17142 vdd.n3025 vdd.n850 99.5127
R17143 vdd.n3025 vdd.n847 99.5127
R17144 vdd.n3074 vdd.n847 99.5127
R17145 vdd.n3074 vdd.n848 99.5127
R17146 vdd.n848 vdd.n839 99.5127
R17147 vdd.n3069 vdd.n839 99.5127
R17148 vdd.n3069 vdd.n807 99.5127
R17149 vdd.n2588 vdd.n2587 99.5127
R17150 vdd.n2584 vdd.n2583 99.5127
R17151 vdd.n2580 vdd.n2579 99.5127
R17152 vdd.n2576 vdd.n2575 99.5127
R17153 vdd.n2572 vdd.n2571 99.5127
R17154 vdd.n2568 vdd.n2567 99.5127
R17155 vdd.n2564 vdd.n2563 99.5127
R17156 vdd.n2560 vdd.n2559 99.5127
R17157 vdd.n2556 vdd.n2555 99.5127
R17158 vdd.n2552 vdd.n2551 99.5127
R17159 vdd.n2548 vdd.n2547 99.5127
R17160 vdd.n2544 vdd.n2543 99.5127
R17161 vdd.n2540 vdd.n2539 99.5127
R17162 vdd.n2536 vdd.n2535 99.5127
R17163 vdd.n2532 vdd.n2531 99.5127
R17164 vdd.n2528 vdd.n2527 99.5127
R17165 vdd.n2524 vdd.n951 99.5127
R17166 vdd.n1387 vdd.n1078 99.5127
R17167 vdd.n1384 vdd.n1078 99.5127
R17168 vdd.n1384 vdd.n1072 99.5127
R17169 vdd.n1381 vdd.n1072 99.5127
R17170 vdd.n1381 vdd.n1067 99.5127
R17171 vdd.n1378 vdd.n1067 99.5127
R17172 vdd.n1378 vdd.n1061 99.5127
R17173 vdd.n1375 vdd.n1061 99.5127
R17174 vdd.n1375 vdd.n1054 99.5127
R17175 vdd.n1372 vdd.n1054 99.5127
R17176 vdd.n1372 vdd.n1047 99.5127
R17177 vdd.n1369 vdd.n1047 99.5127
R17178 vdd.n1369 vdd.n1041 99.5127
R17179 vdd.n1366 vdd.n1041 99.5127
R17180 vdd.n1366 vdd.n1036 99.5127
R17181 vdd.n1363 vdd.n1036 99.5127
R17182 vdd.n1363 vdd.n1030 99.5127
R17183 vdd.n1360 vdd.n1030 99.5127
R17184 vdd.n1360 vdd.n1023 99.5127
R17185 vdd.n1270 vdd.n1023 99.5127
R17186 vdd.n1270 vdd.n1017 99.5127
R17187 vdd.n1267 vdd.n1017 99.5127
R17188 vdd.n1267 vdd.n1012 99.5127
R17189 vdd.n1264 vdd.n1012 99.5127
R17190 vdd.n1264 vdd.n1007 99.5127
R17191 vdd.n1261 vdd.n1007 99.5127
R17192 vdd.n1261 vdd.n1001 99.5127
R17193 vdd.n1258 vdd.n1001 99.5127
R17194 vdd.n1258 vdd.n994 99.5127
R17195 vdd.n994 vdd.n985 99.5127
R17196 vdd.n2519 vdd.n985 99.5127
R17197 vdd.n2520 vdd.n2519 99.5127
R17198 vdd.n2520 vdd.n977 99.5127
R17199 vdd.n1222 vdd.n1082 99.5127
R17200 vdd.n1226 vdd.n1225 99.5127
R17201 vdd.n1230 vdd.n1229 99.5127
R17202 vdd.n1234 vdd.n1233 99.5127
R17203 vdd.n1238 vdd.n1237 99.5127
R17204 vdd.n1242 vdd.n1241 99.5127
R17205 vdd.n1246 vdd.n1245 99.5127
R17206 vdd.n1250 vdd.n1249 99.5127
R17207 vdd.n1420 vdd.n1252 99.5127
R17208 vdd.n1418 vdd.n1417 99.5127
R17209 vdd.n1414 vdd.n1413 99.5127
R17210 vdd.n1410 vdd.n1409 99.5127
R17211 vdd.n1406 vdd.n1405 99.5127
R17212 vdd.n1402 vdd.n1401 99.5127
R17213 vdd.n1398 vdd.n1397 99.5127
R17214 vdd.n1394 vdd.n1393 99.5127
R17215 vdd.n1390 vdd.n1116 99.5127
R17216 vdd.n2423 vdd.n1080 99.5127
R17217 vdd.n2423 vdd.n1070 99.5127
R17218 vdd.n2431 vdd.n1070 99.5127
R17219 vdd.n2431 vdd.n1068 99.5127
R17220 vdd.n2435 vdd.n1068 99.5127
R17221 vdd.n2435 vdd.n1058 99.5127
R17222 vdd.n2443 vdd.n1058 99.5127
R17223 vdd.n2443 vdd.n1056 99.5127
R17224 vdd.n2447 vdd.n1056 99.5127
R17225 vdd.n2447 vdd.n1045 99.5127
R17226 vdd.n2455 vdd.n1045 99.5127
R17227 vdd.n2455 vdd.n1042 99.5127
R17228 vdd.n2460 vdd.n1042 99.5127
R17229 vdd.n2460 vdd.n1033 99.5127
R17230 vdd.n2468 vdd.n1033 99.5127
R17231 vdd.n2468 vdd.n1031 99.5127
R17232 vdd.n2472 vdd.n1031 99.5127
R17233 vdd.n2472 vdd.n1021 99.5127
R17234 vdd.n2480 vdd.n1021 99.5127
R17235 vdd.n2480 vdd.n1019 99.5127
R17236 vdd.n2484 vdd.n1019 99.5127
R17237 vdd.n2484 vdd.n1010 99.5127
R17238 vdd.n2492 vdd.n1010 99.5127
R17239 vdd.n2492 vdd.n1008 99.5127
R17240 vdd.n2496 vdd.n1008 99.5127
R17241 vdd.n2496 vdd.n998 99.5127
R17242 vdd.n2504 vdd.n998 99.5127
R17243 vdd.n2504 vdd.n995 99.5127
R17244 vdd.n2510 vdd.n995 99.5127
R17245 vdd.n2510 vdd.n996 99.5127
R17246 vdd.n996 vdd.n987 99.5127
R17247 vdd.n987 vdd.n978 99.5127
R17248 vdd.n2592 vdd.n978 99.5127
R17249 vdd.n9 vdd.n7 98.9633
R17250 vdd.n2 vdd.n0 98.9633
R17251 vdd.n9 vdd.n8 98.6055
R17252 vdd.n11 vdd.n10 98.6055
R17253 vdd.n13 vdd.n12 98.6055
R17254 vdd.n6 vdd.n5 98.6055
R17255 vdd.n4 vdd.n3 98.6055
R17256 vdd.n2 vdd.n1 98.6055
R17257 vdd.t38 vdd.n303 85.8723
R17258 vdd.t124 vdd.n244 85.8723
R17259 vdd.t174 vdd.n201 85.8723
R17260 vdd.t107 vdd.n142 85.8723
R17261 vdd.t75 vdd.n100 85.8723
R17262 vdd.t64 vdd.n41 85.8723
R17263 vdd.t165 vdd.n2084 85.8723
R17264 vdd.t99 vdd.n2143 85.8723
R17265 vdd.t153 vdd.n1982 85.8723
R17266 vdd.t76 vdd.n2041 85.8723
R17267 vdd.t66 vdd.n1881 85.8723
R17268 vdd.t74 vdd.n1940 85.8723
R17269 vdd.n3003 vdd.n872 78.546
R17270 vdd.n2458 vdd.n1043 78.546
R17271 vdd.n290 vdd.n289 75.1835
R17272 vdd.n288 vdd.n287 75.1835
R17273 vdd.n286 vdd.n285 75.1835
R17274 vdd.n284 vdd.n283 75.1835
R17275 vdd.n282 vdd.n281 75.1835
R17276 vdd.n280 vdd.n279 75.1835
R17277 vdd.n278 vdd.n277 75.1835
R17278 vdd.n276 vdd.n275 75.1835
R17279 vdd.n274 vdd.n273 75.1835
R17280 vdd.n188 vdd.n187 75.1835
R17281 vdd.n186 vdd.n185 75.1835
R17282 vdd.n184 vdd.n183 75.1835
R17283 vdd.n182 vdd.n181 75.1835
R17284 vdd.n180 vdd.n179 75.1835
R17285 vdd.n178 vdd.n177 75.1835
R17286 vdd.n176 vdd.n175 75.1835
R17287 vdd.n174 vdd.n173 75.1835
R17288 vdd.n172 vdd.n171 75.1835
R17289 vdd.n87 vdd.n86 75.1835
R17290 vdd.n85 vdd.n84 75.1835
R17291 vdd.n83 vdd.n82 75.1835
R17292 vdd.n81 vdd.n80 75.1835
R17293 vdd.n79 vdd.n78 75.1835
R17294 vdd.n77 vdd.n76 75.1835
R17295 vdd.n75 vdd.n74 75.1835
R17296 vdd.n73 vdd.n72 75.1835
R17297 vdd.n71 vdd.n70 75.1835
R17298 vdd.n2114 vdd.n2113 75.1835
R17299 vdd.n2116 vdd.n2115 75.1835
R17300 vdd.n2118 vdd.n2117 75.1835
R17301 vdd.n2120 vdd.n2119 75.1835
R17302 vdd.n2122 vdd.n2121 75.1835
R17303 vdd.n2124 vdd.n2123 75.1835
R17304 vdd.n2126 vdd.n2125 75.1835
R17305 vdd.n2128 vdd.n2127 75.1835
R17306 vdd.n2130 vdd.n2129 75.1835
R17307 vdd.n2012 vdd.n2011 75.1835
R17308 vdd.n2014 vdd.n2013 75.1835
R17309 vdd.n2016 vdd.n2015 75.1835
R17310 vdd.n2018 vdd.n2017 75.1835
R17311 vdd.n2020 vdd.n2019 75.1835
R17312 vdd.n2022 vdd.n2021 75.1835
R17313 vdd.n2024 vdd.n2023 75.1835
R17314 vdd.n2026 vdd.n2025 75.1835
R17315 vdd.n2028 vdd.n2027 75.1835
R17316 vdd.n1911 vdd.n1910 75.1835
R17317 vdd.n1913 vdd.n1912 75.1835
R17318 vdd.n1915 vdd.n1914 75.1835
R17319 vdd.n1917 vdd.n1916 75.1835
R17320 vdd.n1919 vdd.n1918 75.1835
R17321 vdd.n1921 vdd.n1920 75.1835
R17322 vdd.n1923 vdd.n1922 75.1835
R17323 vdd.n1925 vdd.n1924 75.1835
R17324 vdd.n1927 vdd.n1926 75.1835
R17325 vdd.n2939 vdd.n2938 72.8958
R17326 vdd.n2938 vdd.n2682 72.8958
R17327 vdd.n2938 vdd.n2683 72.8958
R17328 vdd.n2938 vdd.n2684 72.8958
R17329 vdd.n2938 vdd.n2685 72.8958
R17330 vdd.n2938 vdd.n2686 72.8958
R17331 vdd.n2938 vdd.n2687 72.8958
R17332 vdd.n2938 vdd.n2688 72.8958
R17333 vdd.n2938 vdd.n2689 72.8958
R17334 vdd.n2938 vdd.n2690 72.8958
R17335 vdd.n2938 vdd.n2691 72.8958
R17336 vdd.n2938 vdd.n2692 72.8958
R17337 vdd.n2938 vdd.n2693 72.8958
R17338 vdd.n2938 vdd.n2694 72.8958
R17339 vdd.n2938 vdd.n2695 72.8958
R17340 vdd.n2938 vdd.n2696 72.8958
R17341 vdd.n2938 vdd.n2697 72.8958
R17342 vdd.n803 vdd.n692 72.8958
R17343 vdd.n3158 vdd.n692 72.8958
R17344 vdd.n797 vdd.n692 72.8958
R17345 vdd.n3165 vdd.n692 72.8958
R17346 vdd.n794 vdd.n692 72.8958
R17347 vdd.n3172 vdd.n692 72.8958
R17348 vdd.n791 vdd.n692 72.8958
R17349 vdd.n3179 vdd.n692 72.8958
R17350 vdd.n3182 vdd.n692 72.8958
R17351 vdd.n3038 vdd.n692 72.8958
R17352 vdd.n3043 vdd.n692 72.8958
R17353 vdd.n3037 vdd.n692 72.8958
R17354 vdd.n3050 vdd.n692 72.8958
R17355 vdd.n3034 vdd.n692 72.8958
R17356 vdd.n3057 vdd.n692 72.8958
R17357 vdd.n3031 vdd.n692 72.8958
R17358 vdd.n3064 vdd.n692 72.8958
R17359 vdd.n2417 vdd.n2416 72.8958
R17360 vdd.n2417 vdd.n1084 72.8958
R17361 vdd.n2417 vdd.n1085 72.8958
R17362 vdd.n2417 vdd.n1086 72.8958
R17363 vdd.n2417 vdd.n1087 72.8958
R17364 vdd.n2417 vdd.n1088 72.8958
R17365 vdd.n2417 vdd.n1089 72.8958
R17366 vdd.n2417 vdd.n1090 72.8958
R17367 vdd.n2417 vdd.n1091 72.8958
R17368 vdd.n2417 vdd.n1092 72.8958
R17369 vdd.n2417 vdd.n1093 72.8958
R17370 vdd.n2417 vdd.n1094 72.8958
R17371 vdd.n2417 vdd.n1095 72.8958
R17372 vdd.n2417 vdd.n1096 72.8958
R17373 vdd.n2417 vdd.n1097 72.8958
R17374 vdd.n2417 vdd.n1098 72.8958
R17375 vdd.n2417 vdd.n1099 72.8958
R17376 vdd.n2665 vdd.n952 72.8958
R17377 vdd.n2665 vdd.n953 72.8958
R17378 vdd.n2665 vdd.n954 72.8958
R17379 vdd.n2665 vdd.n955 72.8958
R17380 vdd.n2665 vdd.n956 72.8958
R17381 vdd.n2665 vdd.n957 72.8958
R17382 vdd.n2665 vdd.n958 72.8958
R17383 vdd.n2665 vdd.n959 72.8958
R17384 vdd.n2665 vdd.n960 72.8958
R17385 vdd.n2665 vdd.n961 72.8958
R17386 vdd.n2665 vdd.n962 72.8958
R17387 vdd.n2665 vdd.n963 72.8958
R17388 vdd.n2665 vdd.n964 72.8958
R17389 vdd.n2665 vdd.n965 72.8958
R17390 vdd.n2665 vdd.n966 72.8958
R17391 vdd.n2665 vdd.n967 72.8958
R17392 vdd.n2665 vdd.n968 72.8958
R17393 vdd.n2938 vdd.n2937 72.8958
R17394 vdd.n2938 vdd.n2666 72.8958
R17395 vdd.n2938 vdd.n2667 72.8958
R17396 vdd.n2938 vdd.n2668 72.8958
R17397 vdd.n2938 vdd.n2669 72.8958
R17398 vdd.n2938 vdd.n2670 72.8958
R17399 vdd.n2938 vdd.n2671 72.8958
R17400 vdd.n2938 vdd.n2672 72.8958
R17401 vdd.n2938 vdd.n2673 72.8958
R17402 vdd.n2938 vdd.n2674 72.8958
R17403 vdd.n2938 vdd.n2675 72.8958
R17404 vdd.n2938 vdd.n2676 72.8958
R17405 vdd.n2938 vdd.n2677 72.8958
R17406 vdd.n2938 vdd.n2678 72.8958
R17407 vdd.n2938 vdd.n2679 72.8958
R17408 vdd.n2938 vdd.n2680 72.8958
R17409 vdd.n2938 vdd.n2681 72.8958
R17410 vdd.n3088 vdd.n692 72.8958
R17411 vdd.n835 vdd.n692 72.8958
R17412 vdd.n3096 vdd.n692 72.8958
R17413 vdd.n830 vdd.n692 72.8958
R17414 vdd.n3103 vdd.n692 72.8958
R17415 vdd.n827 vdd.n692 72.8958
R17416 vdd.n3110 vdd.n692 72.8958
R17417 vdd.n824 vdd.n692 72.8958
R17418 vdd.n3117 vdd.n692 72.8958
R17419 vdd.n3121 vdd.n692 72.8958
R17420 vdd.n821 vdd.n692 72.8958
R17421 vdd.n3128 vdd.n692 72.8958
R17422 vdd.n818 vdd.n692 72.8958
R17423 vdd.n3135 vdd.n692 72.8958
R17424 vdd.n815 vdd.n692 72.8958
R17425 vdd.n3142 vdd.n692 72.8958
R17426 vdd.n3145 vdd.n692 72.8958
R17427 vdd.n2665 vdd.n950 72.8958
R17428 vdd.n2665 vdd.n949 72.8958
R17429 vdd.n2665 vdd.n948 72.8958
R17430 vdd.n2665 vdd.n947 72.8958
R17431 vdd.n2665 vdd.n946 72.8958
R17432 vdd.n2665 vdd.n945 72.8958
R17433 vdd.n2665 vdd.n944 72.8958
R17434 vdd.n2665 vdd.n943 72.8958
R17435 vdd.n2665 vdd.n942 72.8958
R17436 vdd.n2665 vdd.n941 72.8958
R17437 vdd.n2665 vdd.n940 72.8958
R17438 vdd.n2665 vdd.n939 72.8958
R17439 vdd.n2665 vdd.n938 72.8958
R17440 vdd.n2665 vdd.n937 72.8958
R17441 vdd.n2665 vdd.n936 72.8958
R17442 vdd.n2665 vdd.n935 72.8958
R17443 vdd.n2665 vdd.n934 72.8958
R17444 vdd.n2418 vdd.n2417 72.8958
R17445 vdd.n2417 vdd.n1100 72.8958
R17446 vdd.n2417 vdd.n1101 72.8958
R17447 vdd.n2417 vdd.n1102 72.8958
R17448 vdd.n2417 vdd.n1103 72.8958
R17449 vdd.n2417 vdd.n1104 72.8958
R17450 vdd.n2417 vdd.n1105 72.8958
R17451 vdd.n2417 vdd.n1106 72.8958
R17452 vdd.n2417 vdd.n1107 72.8958
R17453 vdd.n2417 vdd.n1108 72.8958
R17454 vdd.n2417 vdd.n1109 72.8958
R17455 vdd.n2417 vdd.n1110 72.8958
R17456 vdd.n2417 vdd.n1111 72.8958
R17457 vdd.n2417 vdd.n1112 72.8958
R17458 vdd.n2417 vdd.n1113 72.8958
R17459 vdd.n2417 vdd.n1114 72.8958
R17460 vdd.n2417 vdd.n1115 72.8958
R17461 vdd.n1781 vdd.n1780 66.2847
R17462 vdd.n1780 vdd.n1556 66.2847
R17463 vdd.n1780 vdd.n1557 66.2847
R17464 vdd.n1780 vdd.n1558 66.2847
R17465 vdd.n1780 vdd.n1559 66.2847
R17466 vdd.n1780 vdd.n1560 66.2847
R17467 vdd.n1780 vdd.n1561 66.2847
R17468 vdd.n1780 vdd.n1562 66.2847
R17469 vdd.n1780 vdd.n1563 66.2847
R17470 vdd.n1780 vdd.n1564 66.2847
R17471 vdd.n1780 vdd.n1565 66.2847
R17472 vdd.n1780 vdd.n1566 66.2847
R17473 vdd.n1780 vdd.n1567 66.2847
R17474 vdd.n1780 vdd.n1568 66.2847
R17475 vdd.n1780 vdd.n1569 66.2847
R17476 vdd.n1780 vdd.n1570 66.2847
R17477 vdd.n1780 vdd.n1571 66.2847
R17478 vdd.n1780 vdd.n1572 66.2847
R17479 vdd.n1780 vdd.n1573 66.2847
R17480 vdd.n1780 vdd.n1574 66.2847
R17481 vdd.n1780 vdd.n1575 66.2847
R17482 vdd.n1780 vdd.n1576 66.2847
R17483 vdd.n1780 vdd.n1577 66.2847
R17484 vdd.n1780 vdd.n1578 66.2847
R17485 vdd.n1780 vdd.n1579 66.2847
R17486 vdd.n1780 vdd.n1580 66.2847
R17487 vdd.n1780 vdd.n1581 66.2847
R17488 vdd.n1780 vdd.n1582 66.2847
R17489 vdd.n1780 vdd.n1583 66.2847
R17490 vdd.n1780 vdd.n1584 66.2847
R17491 vdd.n1780 vdd.n1585 66.2847
R17492 vdd.n1433 vdd.n1083 66.2847
R17493 vdd.n1430 vdd.n1083 66.2847
R17494 vdd.n1426 vdd.n1083 66.2847
R17495 vdd.n2279 vdd.n1083 66.2847
R17496 vdd.n1217 vdd.n1083 66.2847
R17497 vdd.n2286 vdd.n1083 66.2847
R17498 vdd.n1210 vdd.n1083 66.2847
R17499 vdd.n2293 vdd.n1083 66.2847
R17500 vdd.n1203 vdd.n1083 66.2847
R17501 vdd.n2300 vdd.n1083 66.2847
R17502 vdd.n1197 vdd.n1083 66.2847
R17503 vdd.n1192 vdd.n1083 66.2847
R17504 vdd.n2311 vdd.n1083 66.2847
R17505 vdd.n1184 vdd.n1083 66.2847
R17506 vdd.n2318 vdd.n1083 66.2847
R17507 vdd.n1177 vdd.n1083 66.2847
R17508 vdd.n2325 vdd.n1083 66.2847
R17509 vdd.n1170 vdd.n1083 66.2847
R17510 vdd.n2332 vdd.n1083 66.2847
R17511 vdd.n1163 vdd.n1083 66.2847
R17512 vdd.n2339 vdd.n1083 66.2847
R17513 vdd.n1157 vdd.n1083 66.2847
R17514 vdd.n1152 vdd.n1083 66.2847
R17515 vdd.n2350 vdd.n1083 66.2847
R17516 vdd.n1144 vdd.n1083 66.2847
R17517 vdd.n2357 vdd.n1083 66.2847
R17518 vdd.n1137 vdd.n1083 66.2847
R17519 vdd.n2364 vdd.n1083 66.2847
R17520 vdd.n1130 vdd.n1083 66.2847
R17521 vdd.n2371 vdd.n1083 66.2847
R17522 vdd.n2376 vdd.n1083 66.2847
R17523 vdd.n1126 vdd.n1083 66.2847
R17524 vdd.n3315 vdd.n3314 66.2847
R17525 vdd.n3315 vdd.n693 66.2847
R17526 vdd.n3315 vdd.n694 66.2847
R17527 vdd.n3315 vdd.n695 66.2847
R17528 vdd.n3315 vdd.n696 66.2847
R17529 vdd.n3315 vdd.n697 66.2847
R17530 vdd.n3315 vdd.n698 66.2847
R17531 vdd.n3315 vdd.n699 66.2847
R17532 vdd.n3315 vdd.n700 66.2847
R17533 vdd.n3315 vdd.n701 66.2847
R17534 vdd.n3315 vdd.n702 66.2847
R17535 vdd.n3315 vdd.n703 66.2847
R17536 vdd.n3315 vdd.n704 66.2847
R17537 vdd.n3315 vdd.n705 66.2847
R17538 vdd.n3315 vdd.n706 66.2847
R17539 vdd.n3315 vdd.n707 66.2847
R17540 vdd.n3315 vdd.n708 66.2847
R17541 vdd.n3315 vdd.n709 66.2847
R17542 vdd.n3315 vdd.n710 66.2847
R17543 vdd.n3315 vdd.n711 66.2847
R17544 vdd.n3315 vdd.n712 66.2847
R17545 vdd.n3315 vdd.n713 66.2847
R17546 vdd.n3315 vdd.n714 66.2847
R17547 vdd.n3315 vdd.n715 66.2847
R17548 vdd.n3315 vdd.n716 66.2847
R17549 vdd.n3315 vdd.n717 66.2847
R17550 vdd.n3315 vdd.n718 66.2847
R17551 vdd.n3315 vdd.n719 66.2847
R17552 vdd.n3315 vdd.n720 66.2847
R17553 vdd.n3315 vdd.n721 66.2847
R17554 vdd.n3315 vdd.n722 66.2847
R17555 vdd.n3446 vdd.n3445 66.2847
R17556 vdd.n3446 vdd.n424 66.2847
R17557 vdd.n3446 vdd.n423 66.2847
R17558 vdd.n3446 vdd.n422 66.2847
R17559 vdd.n3446 vdd.n421 66.2847
R17560 vdd.n3446 vdd.n420 66.2847
R17561 vdd.n3446 vdd.n419 66.2847
R17562 vdd.n3446 vdd.n418 66.2847
R17563 vdd.n3446 vdd.n417 66.2847
R17564 vdd.n3446 vdd.n416 66.2847
R17565 vdd.n3446 vdd.n415 66.2847
R17566 vdd.n3446 vdd.n414 66.2847
R17567 vdd.n3446 vdd.n413 66.2847
R17568 vdd.n3446 vdd.n412 66.2847
R17569 vdd.n3446 vdd.n411 66.2847
R17570 vdd.n3446 vdd.n410 66.2847
R17571 vdd.n3446 vdd.n409 66.2847
R17572 vdd.n3446 vdd.n408 66.2847
R17573 vdd.n3446 vdd.n407 66.2847
R17574 vdd.n3446 vdd.n406 66.2847
R17575 vdd.n3446 vdd.n405 66.2847
R17576 vdd.n3446 vdd.n404 66.2847
R17577 vdd.n3446 vdd.n403 66.2847
R17578 vdd.n3446 vdd.n402 66.2847
R17579 vdd.n3446 vdd.n401 66.2847
R17580 vdd.n3446 vdd.n400 66.2847
R17581 vdd.n3446 vdd.n399 66.2847
R17582 vdd.n3446 vdd.n398 66.2847
R17583 vdd.n3446 vdd.n397 66.2847
R17584 vdd.n3446 vdd.n396 66.2847
R17585 vdd.n3446 vdd.n395 66.2847
R17586 vdd.n3446 vdd.n394 66.2847
R17587 vdd.n467 vdd.n394 52.4337
R17588 vdd.n473 vdd.n395 52.4337
R17589 vdd.n477 vdd.n396 52.4337
R17590 vdd.n483 vdd.n397 52.4337
R17591 vdd.n487 vdd.n398 52.4337
R17592 vdd.n493 vdd.n399 52.4337
R17593 vdd.n497 vdd.n400 52.4337
R17594 vdd.n503 vdd.n401 52.4337
R17595 vdd.n507 vdd.n402 52.4337
R17596 vdd.n513 vdd.n403 52.4337
R17597 vdd.n517 vdd.n404 52.4337
R17598 vdd.n523 vdd.n405 52.4337
R17599 vdd.n527 vdd.n406 52.4337
R17600 vdd.n533 vdd.n407 52.4337
R17601 vdd.n537 vdd.n408 52.4337
R17602 vdd.n543 vdd.n409 52.4337
R17603 vdd.n547 vdd.n410 52.4337
R17604 vdd.n553 vdd.n411 52.4337
R17605 vdd.n557 vdd.n412 52.4337
R17606 vdd.n563 vdd.n413 52.4337
R17607 vdd.n567 vdd.n414 52.4337
R17608 vdd.n573 vdd.n415 52.4337
R17609 vdd.n577 vdd.n416 52.4337
R17610 vdd.n583 vdd.n417 52.4337
R17611 vdd.n587 vdd.n418 52.4337
R17612 vdd.n593 vdd.n419 52.4337
R17613 vdd.n597 vdd.n420 52.4337
R17614 vdd.n603 vdd.n421 52.4337
R17615 vdd.n607 vdd.n422 52.4337
R17616 vdd.n613 vdd.n423 52.4337
R17617 vdd.n616 vdd.n424 52.4337
R17618 vdd.n3445 vdd.n3444 52.4337
R17619 vdd.n3314 vdd.n3313 52.4337
R17620 vdd.n728 vdd.n693 52.4337
R17621 vdd.n734 vdd.n694 52.4337
R17622 vdd.n3303 vdd.n695 52.4337
R17623 vdd.n3299 vdd.n696 52.4337
R17624 vdd.n3295 vdd.n697 52.4337
R17625 vdd.n3291 vdd.n698 52.4337
R17626 vdd.n3287 vdd.n699 52.4337
R17627 vdd.n3283 vdd.n700 52.4337
R17628 vdd.n3279 vdd.n701 52.4337
R17629 vdd.n3271 vdd.n702 52.4337
R17630 vdd.n3267 vdd.n703 52.4337
R17631 vdd.n3263 vdd.n704 52.4337
R17632 vdd.n3259 vdd.n705 52.4337
R17633 vdd.n3255 vdd.n706 52.4337
R17634 vdd.n3251 vdd.n707 52.4337
R17635 vdd.n3247 vdd.n708 52.4337
R17636 vdd.n3243 vdd.n709 52.4337
R17637 vdd.n3239 vdd.n710 52.4337
R17638 vdd.n3235 vdd.n711 52.4337
R17639 vdd.n3231 vdd.n712 52.4337
R17640 vdd.n3225 vdd.n713 52.4337
R17641 vdd.n3221 vdd.n714 52.4337
R17642 vdd.n3217 vdd.n715 52.4337
R17643 vdd.n3213 vdd.n716 52.4337
R17644 vdd.n3209 vdd.n717 52.4337
R17645 vdd.n3205 vdd.n718 52.4337
R17646 vdd.n3201 vdd.n719 52.4337
R17647 vdd.n3197 vdd.n720 52.4337
R17648 vdd.n3193 vdd.n721 52.4337
R17649 vdd.n3189 vdd.n722 52.4337
R17650 vdd.n2378 vdd.n1126 52.4337
R17651 vdd.n2376 vdd.n2375 52.4337
R17652 vdd.n2371 vdd.n2370 52.4337
R17653 vdd.n2366 vdd.n1130 52.4337
R17654 vdd.n2364 vdd.n2363 52.4337
R17655 vdd.n2359 vdd.n1137 52.4337
R17656 vdd.n2357 vdd.n2356 52.4337
R17657 vdd.n2352 vdd.n1144 52.4337
R17658 vdd.n2350 vdd.n2349 52.4337
R17659 vdd.n1153 vdd.n1152 52.4337
R17660 vdd.n2341 vdd.n1157 52.4337
R17661 vdd.n2339 vdd.n2338 52.4337
R17662 vdd.n2334 vdd.n1163 52.4337
R17663 vdd.n2332 vdd.n2331 52.4337
R17664 vdd.n2327 vdd.n1170 52.4337
R17665 vdd.n2325 vdd.n2324 52.4337
R17666 vdd.n2320 vdd.n1177 52.4337
R17667 vdd.n2318 vdd.n2317 52.4337
R17668 vdd.n2313 vdd.n1184 52.4337
R17669 vdd.n2311 vdd.n2310 52.4337
R17670 vdd.n1193 vdd.n1192 52.4337
R17671 vdd.n2302 vdd.n1197 52.4337
R17672 vdd.n2300 vdd.n2299 52.4337
R17673 vdd.n2295 vdd.n1203 52.4337
R17674 vdd.n2293 vdd.n2292 52.4337
R17675 vdd.n2288 vdd.n1210 52.4337
R17676 vdd.n2286 vdd.n2285 52.4337
R17677 vdd.n2281 vdd.n1217 52.4337
R17678 vdd.n2279 vdd.n2278 52.4337
R17679 vdd.n1427 vdd.n1426 52.4337
R17680 vdd.n1431 vdd.n1430 52.4337
R17681 vdd.n2267 vdd.n1433 52.4337
R17682 vdd.n1782 vdd.n1781 52.4337
R17683 vdd.n1588 vdd.n1556 52.4337
R17684 vdd.n1592 vdd.n1557 52.4337
R17685 vdd.n1594 vdd.n1558 52.4337
R17686 vdd.n1598 vdd.n1559 52.4337
R17687 vdd.n1600 vdd.n1560 52.4337
R17688 vdd.n1604 vdd.n1561 52.4337
R17689 vdd.n1606 vdd.n1562 52.4337
R17690 vdd.n1610 vdd.n1563 52.4337
R17691 vdd.n1612 vdd.n1564 52.4337
R17692 vdd.n1618 vdd.n1565 52.4337
R17693 vdd.n1620 vdd.n1566 52.4337
R17694 vdd.n1624 vdd.n1567 52.4337
R17695 vdd.n1626 vdd.n1568 52.4337
R17696 vdd.n1630 vdd.n1569 52.4337
R17697 vdd.n1632 vdd.n1570 52.4337
R17698 vdd.n1636 vdd.n1571 52.4337
R17699 vdd.n1638 vdd.n1572 52.4337
R17700 vdd.n1642 vdd.n1573 52.4337
R17701 vdd.n1644 vdd.n1574 52.4337
R17702 vdd.n1716 vdd.n1575 52.4337
R17703 vdd.n1649 vdd.n1576 52.4337
R17704 vdd.n1653 vdd.n1577 52.4337
R17705 vdd.n1655 vdd.n1578 52.4337
R17706 vdd.n1659 vdd.n1579 52.4337
R17707 vdd.n1661 vdd.n1580 52.4337
R17708 vdd.n1665 vdd.n1581 52.4337
R17709 vdd.n1667 vdd.n1582 52.4337
R17710 vdd.n1671 vdd.n1583 52.4337
R17711 vdd.n1673 vdd.n1584 52.4337
R17712 vdd.n1677 vdd.n1585 52.4337
R17713 vdd.n1781 vdd.n1555 52.4337
R17714 vdd.n1591 vdd.n1556 52.4337
R17715 vdd.n1593 vdd.n1557 52.4337
R17716 vdd.n1597 vdd.n1558 52.4337
R17717 vdd.n1599 vdd.n1559 52.4337
R17718 vdd.n1603 vdd.n1560 52.4337
R17719 vdd.n1605 vdd.n1561 52.4337
R17720 vdd.n1609 vdd.n1562 52.4337
R17721 vdd.n1611 vdd.n1563 52.4337
R17722 vdd.n1617 vdd.n1564 52.4337
R17723 vdd.n1619 vdd.n1565 52.4337
R17724 vdd.n1623 vdd.n1566 52.4337
R17725 vdd.n1625 vdd.n1567 52.4337
R17726 vdd.n1629 vdd.n1568 52.4337
R17727 vdd.n1631 vdd.n1569 52.4337
R17728 vdd.n1635 vdd.n1570 52.4337
R17729 vdd.n1637 vdd.n1571 52.4337
R17730 vdd.n1641 vdd.n1572 52.4337
R17731 vdd.n1643 vdd.n1573 52.4337
R17732 vdd.n1647 vdd.n1574 52.4337
R17733 vdd.n1648 vdd.n1575 52.4337
R17734 vdd.n1652 vdd.n1576 52.4337
R17735 vdd.n1654 vdd.n1577 52.4337
R17736 vdd.n1658 vdd.n1578 52.4337
R17737 vdd.n1660 vdd.n1579 52.4337
R17738 vdd.n1664 vdd.n1580 52.4337
R17739 vdd.n1666 vdd.n1581 52.4337
R17740 vdd.n1670 vdd.n1582 52.4337
R17741 vdd.n1672 vdd.n1583 52.4337
R17742 vdd.n1676 vdd.n1584 52.4337
R17743 vdd.n1678 vdd.n1585 52.4337
R17744 vdd.n1433 vdd.n1432 52.4337
R17745 vdd.n1430 vdd.n1429 52.4337
R17746 vdd.n1426 vdd.n1218 52.4337
R17747 vdd.n2280 vdd.n2279 52.4337
R17748 vdd.n1217 vdd.n1211 52.4337
R17749 vdd.n2287 vdd.n2286 52.4337
R17750 vdd.n1210 vdd.n1204 52.4337
R17751 vdd.n2294 vdd.n2293 52.4337
R17752 vdd.n1203 vdd.n1198 52.4337
R17753 vdd.n2301 vdd.n2300 52.4337
R17754 vdd.n1197 vdd.n1196 52.4337
R17755 vdd.n1192 vdd.n1185 52.4337
R17756 vdd.n2312 vdd.n2311 52.4337
R17757 vdd.n1184 vdd.n1178 52.4337
R17758 vdd.n2319 vdd.n2318 52.4337
R17759 vdd.n1177 vdd.n1171 52.4337
R17760 vdd.n2326 vdd.n2325 52.4337
R17761 vdd.n1170 vdd.n1164 52.4337
R17762 vdd.n2333 vdd.n2332 52.4337
R17763 vdd.n1163 vdd.n1158 52.4337
R17764 vdd.n2340 vdd.n2339 52.4337
R17765 vdd.n1157 vdd.n1156 52.4337
R17766 vdd.n1152 vdd.n1145 52.4337
R17767 vdd.n2351 vdd.n2350 52.4337
R17768 vdd.n1144 vdd.n1138 52.4337
R17769 vdd.n2358 vdd.n2357 52.4337
R17770 vdd.n1137 vdd.n1131 52.4337
R17771 vdd.n2365 vdd.n2364 52.4337
R17772 vdd.n1130 vdd.n1127 52.4337
R17773 vdd.n2372 vdd.n2371 52.4337
R17774 vdd.n2377 vdd.n2376 52.4337
R17775 vdd.n1437 vdd.n1126 52.4337
R17776 vdd.n3314 vdd.n725 52.4337
R17777 vdd.n733 vdd.n693 52.4337
R17778 vdd.n3304 vdd.n694 52.4337
R17779 vdd.n3300 vdd.n695 52.4337
R17780 vdd.n3296 vdd.n696 52.4337
R17781 vdd.n3292 vdd.n697 52.4337
R17782 vdd.n3288 vdd.n698 52.4337
R17783 vdd.n3284 vdd.n699 52.4337
R17784 vdd.n3280 vdd.n700 52.4337
R17785 vdd.n3270 vdd.n701 52.4337
R17786 vdd.n3268 vdd.n702 52.4337
R17787 vdd.n3264 vdd.n703 52.4337
R17788 vdd.n3260 vdd.n704 52.4337
R17789 vdd.n3256 vdd.n705 52.4337
R17790 vdd.n3252 vdd.n706 52.4337
R17791 vdd.n3248 vdd.n707 52.4337
R17792 vdd.n3244 vdd.n708 52.4337
R17793 vdd.n3240 vdd.n709 52.4337
R17794 vdd.n3236 vdd.n710 52.4337
R17795 vdd.n3232 vdd.n711 52.4337
R17796 vdd.n3224 vdd.n712 52.4337
R17797 vdd.n3222 vdd.n713 52.4337
R17798 vdd.n3218 vdd.n714 52.4337
R17799 vdd.n3214 vdd.n715 52.4337
R17800 vdd.n3210 vdd.n716 52.4337
R17801 vdd.n3206 vdd.n717 52.4337
R17802 vdd.n3202 vdd.n718 52.4337
R17803 vdd.n3198 vdd.n719 52.4337
R17804 vdd.n3194 vdd.n720 52.4337
R17805 vdd.n3190 vdd.n721 52.4337
R17806 vdd.n722 vdd.n691 52.4337
R17807 vdd.n3445 vdd.n425 52.4337
R17808 vdd.n614 vdd.n424 52.4337
R17809 vdd.n608 vdd.n423 52.4337
R17810 vdd.n604 vdd.n422 52.4337
R17811 vdd.n598 vdd.n421 52.4337
R17812 vdd.n594 vdd.n420 52.4337
R17813 vdd.n588 vdd.n419 52.4337
R17814 vdd.n584 vdd.n418 52.4337
R17815 vdd.n578 vdd.n417 52.4337
R17816 vdd.n574 vdd.n416 52.4337
R17817 vdd.n568 vdd.n415 52.4337
R17818 vdd.n564 vdd.n414 52.4337
R17819 vdd.n558 vdd.n413 52.4337
R17820 vdd.n554 vdd.n412 52.4337
R17821 vdd.n548 vdd.n411 52.4337
R17822 vdd.n544 vdd.n410 52.4337
R17823 vdd.n538 vdd.n409 52.4337
R17824 vdd.n534 vdd.n408 52.4337
R17825 vdd.n528 vdd.n407 52.4337
R17826 vdd.n524 vdd.n406 52.4337
R17827 vdd.n518 vdd.n405 52.4337
R17828 vdd.n514 vdd.n404 52.4337
R17829 vdd.n508 vdd.n403 52.4337
R17830 vdd.n504 vdd.n402 52.4337
R17831 vdd.n498 vdd.n401 52.4337
R17832 vdd.n494 vdd.n400 52.4337
R17833 vdd.n488 vdd.n399 52.4337
R17834 vdd.n484 vdd.n398 52.4337
R17835 vdd.n478 vdd.n397 52.4337
R17836 vdd.n474 vdd.n396 52.4337
R17837 vdd.n468 vdd.n395 52.4337
R17838 vdd.n394 vdd.n392 52.4337
R17839 vdd.t293 vdd.t209 51.4683
R17840 vdd.n274 vdd.n272 42.0461
R17841 vdd.n172 vdd.n170 42.0461
R17842 vdd.n71 vdd.n69 42.0461
R17843 vdd.n2114 vdd.n2112 42.0461
R17844 vdd.n2012 vdd.n2010 42.0461
R17845 vdd.n1911 vdd.n1909 42.0461
R17846 vdd.n332 vdd.n331 41.6884
R17847 vdd.n230 vdd.n229 41.6884
R17848 vdd.n129 vdd.n128 41.6884
R17849 vdd.n2172 vdd.n2171 41.6884
R17850 vdd.n2070 vdd.n2069 41.6884
R17851 vdd.n1969 vdd.n1968 41.6884
R17852 vdd.n1681 vdd.n1680 41.1157
R17853 vdd.n1719 vdd.n1718 41.1157
R17854 vdd.n1615 vdd.n1614 41.1157
R17855 vdd.n428 vdd.n427 41.1157
R17856 vdd.n566 vdd.n441 41.1157
R17857 vdd.n454 vdd.n453 41.1157
R17858 vdd.n3145 vdd.n3144 39.2114
R17859 vdd.n3142 vdd.n3141 39.2114
R17860 vdd.n3137 vdd.n815 39.2114
R17861 vdd.n3135 vdd.n3134 39.2114
R17862 vdd.n3130 vdd.n818 39.2114
R17863 vdd.n3128 vdd.n3127 39.2114
R17864 vdd.n3123 vdd.n821 39.2114
R17865 vdd.n3121 vdd.n3120 39.2114
R17866 vdd.n3117 vdd.n3116 39.2114
R17867 vdd.n3112 vdd.n824 39.2114
R17868 vdd.n3110 vdd.n3109 39.2114
R17869 vdd.n3105 vdd.n827 39.2114
R17870 vdd.n3103 vdd.n3102 39.2114
R17871 vdd.n3098 vdd.n830 39.2114
R17872 vdd.n3096 vdd.n3095 39.2114
R17873 vdd.n3090 vdd.n835 39.2114
R17874 vdd.n3088 vdd.n3087 39.2114
R17875 vdd.n2937 vdd.n2936 39.2114
R17876 vdd.n2931 vdd.n2666 39.2114
R17877 vdd.n2928 vdd.n2667 39.2114
R17878 vdd.n2924 vdd.n2668 39.2114
R17879 vdd.n2920 vdd.n2669 39.2114
R17880 vdd.n2916 vdd.n2670 39.2114
R17881 vdd.n2912 vdd.n2671 39.2114
R17882 vdd.n2908 vdd.n2672 39.2114
R17883 vdd.n2904 vdd.n2673 39.2114
R17884 vdd.n2900 vdd.n2674 39.2114
R17885 vdd.n2896 vdd.n2675 39.2114
R17886 vdd.n2892 vdd.n2676 39.2114
R17887 vdd.n2888 vdd.n2677 39.2114
R17888 vdd.n2884 vdd.n2678 39.2114
R17889 vdd.n2880 vdd.n2679 39.2114
R17890 vdd.n2876 vdd.n2680 39.2114
R17891 vdd.n2871 vdd.n2681 39.2114
R17892 vdd.n2660 vdd.n968 39.2114
R17893 vdd.n2656 vdd.n967 39.2114
R17894 vdd.n2652 vdd.n966 39.2114
R17895 vdd.n2648 vdd.n965 39.2114
R17896 vdd.n2644 vdd.n964 39.2114
R17897 vdd.n2640 vdd.n963 39.2114
R17898 vdd.n2636 vdd.n962 39.2114
R17899 vdd.n2632 vdd.n961 39.2114
R17900 vdd.n2628 vdd.n960 39.2114
R17901 vdd.n2624 vdd.n959 39.2114
R17902 vdd.n2620 vdd.n958 39.2114
R17903 vdd.n2616 vdd.n957 39.2114
R17904 vdd.n2612 vdd.n956 39.2114
R17905 vdd.n2608 vdd.n955 39.2114
R17906 vdd.n2604 vdd.n954 39.2114
R17907 vdd.n2599 vdd.n953 39.2114
R17908 vdd.n2595 vdd.n952 39.2114
R17909 vdd.n2416 vdd.n2415 39.2114
R17910 vdd.n2410 vdd.n1084 39.2114
R17911 vdd.n2407 vdd.n1085 39.2114
R17912 vdd.n2403 vdd.n1086 39.2114
R17913 vdd.n2399 vdd.n1087 39.2114
R17914 vdd.n2395 vdd.n1088 39.2114
R17915 vdd.n2391 vdd.n1089 39.2114
R17916 vdd.n2387 vdd.n1090 39.2114
R17917 vdd.n2383 vdd.n1091 39.2114
R17918 vdd.n1276 vdd.n1092 39.2114
R17919 vdd.n1280 vdd.n1093 39.2114
R17920 vdd.n1284 vdd.n1094 39.2114
R17921 vdd.n1288 vdd.n1095 39.2114
R17922 vdd.n1292 vdd.n1096 39.2114
R17923 vdd.n1296 vdd.n1097 39.2114
R17924 vdd.n1300 vdd.n1098 39.2114
R17925 vdd.n1305 vdd.n1099 39.2114
R17926 vdd.n3064 vdd.n3063 39.2114
R17927 vdd.n3059 vdd.n3031 39.2114
R17928 vdd.n3057 vdd.n3056 39.2114
R17929 vdd.n3052 vdd.n3034 39.2114
R17930 vdd.n3050 vdd.n3049 39.2114
R17931 vdd.n3045 vdd.n3037 39.2114
R17932 vdd.n3043 vdd.n3042 39.2114
R17933 vdd.n3038 vdd.n787 39.2114
R17934 vdd.n3182 vdd.n3181 39.2114
R17935 vdd.n3179 vdd.n3178 39.2114
R17936 vdd.n3174 vdd.n791 39.2114
R17937 vdd.n3172 vdd.n3171 39.2114
R17938 vdd.n3167 vdd.n794 39.2114
R17939 vdd.n3165 vdd.n3164 39.2114
R17940 vdd.n3160 vdd.n797 39.2114
R17941 vdd.n3158 vdd.n3157 39.2114
R17942 vdd.n3153 vdd.n803 39.2114
R17943 vdd.n2940 vdd.n2939 39.2114
R17944 vdd.n2707 vdd.n2682 39.2114
R17945 vdd.n2711 vdd.n2683 39.2114
R17946 vdd.n2715 vdd.n2684 39.2114
R17947 vdd.n2719 vdd.n2685 39.2114
R17948 vdd.n2723 vdd.n2686 39.2114
R17949 vdd.n2727 vdd.n2687 39.2114
R17950 vdd.n2731 vdd.n2688 39.2114
R17951 vdd.n2735 vdd.n2689 39.2114
R17952 vdd.n2739 vdd.n2690 39.2114
R17953 vdd.n2743 vdd.n2691 39.2114
R17954 vdd.n2747 vdd.n2692 39.2114
R17955 vdd.n2751 vdd.n2693 39.2114
R17956 vdd.n2755 vdd.n2694 39.2114
R17957 vdd.n2759 vdd.n2695 39.2114
R17958 vdd.n2763 vdd.n2696 39.2114
R17959 vdd.n2767 vdd.n2697 39.2114
R17960 vdd.n2939 vdd.n933 39.2114
R17961 vdd.n2710 vdd.n2682 39.2114
R17962 vdd.n2714 vdd.n2683 39.2114
R17963 vdd.n2718 vdd.n2684 39.2114
R17964 vdd.n2722 vdd.n2685 39.2114
R17965 vdd.n2726 vdd.n2686 39.2114
R17966 vdd.n2730 vdd.n2687 39.2114
R17967 vdd.n2734 vdd.n2688 39.2114
R17968 vdd.n2738 vdd.n2689 39.2114
R17969 vdd.n2742 vdd.n2690 39.2114
R17970 vdd.n2746 vdd.n2691 39.2114
R17971 vdd.n2750 vdd.n2692 39.2114
R17972 vdd.n2754 vdd.n2693 39.2114
R17973 vdd.n2758 vdd.n2694 39.2114
R17974 vdd.n2762 vdd.n2695 39.2114
R17975 vdd.n2766 vdd.n2696 39.2114
R17976 vdd.n2769 vdd.n2697 39.2114
R17977 vdd.n803 vdd.n798 39.2114
R17978 vdd.n3159 vdd.n3158 39.2114
R17979 vdd.n797 vdd.n795 39.2114
R17980 vdd.n3166 vdd.n3165 39.2114
R17981 vdd.n794 vdd.n792 39.2114
R17982 vdd.n3173 vdd.n3172 39.2114
R17983 vdd.n791 vdd.n789 39.2114
R17984 vdd.n3180 vdd.n3179 39.2114
R17985 vdd.n3183 vdd.n3182 39.2114
R17986 vdd.n3039 vdd.n3038 39.2114
R17987 vdd.n3044 vdd.n3043 39.2114
R17988 vdd.n3037 vdd.n3035 39.2114
R17989 vdd.n3051 vdd.n3050 39.2114
R17990 vdd.n3034 vdd.n3032 39.2114
R17991 vdd.n3058 vdd.n3057 39.2114
R17992 vdd.n3031 vdd.n3029 39.2114
R17993 vdd.n3065 vdd.n3064 39.2114
R17994 vdd.n2416 vdd.n1118 39.2114
R17995 vdd.n2408 vdd.n1084 39.2114
R17996 vdd.n2404 vdd.n1085 39.2114
R17997 vdd.n2400 vdd.n1086 39.2114
R17998 vdd.n2396 vdd.n1087 39.2114
R17999 vdd.n2392 vdd.n1088 39.2114
R18000 vdd.n2388 vdd.n1089 39.2114
R18001 vdd.n2384 vdd.n1090 39.2114
R18002 vdd.n1275 vdd.n1091 39.2114
R18003 vdd.n1279 vdd.n1092 39.2114
R18004 vdd.n1283 vdd.n1093 39.2114
R18005 vdd.n1287 vdd.n1094 39.2114
R18006 vdd.n1291 vdd.n1095 39.2114
R18007 vdd.n1295 vdd.n1096 39.2114
R18008 vdd.n1299 vdd.n1097 39.2114
R18009 vdd.n1304 vdd.n1098 39.2114
R18010 vdd.n1308 vdd.n1099 39.2114
R18011 vdd.n2598 vdd.n952 39.2114
R18012 vdd.n2603 vdd.n953 39.2114
R18013 vdd.n2607 vdd.n954 39.2114
R18014 vdd.n2611 vdd.n955 39.2114
R18015 vdd.n2615 vdd.n956 39.2114
R18016 vdd.n2619 vdd.n957 39.2114
R18017 vdd.n2623 vdd.n958 39.2114
R18018 vdd.n2627 vdd.n959 39.2114
R18019 vdd.n2631 vdd.n960 39.2114
R18020 vdd.n2635 vdd.n961 39.2114
R18021 vdd.n2639 vdd.n962 39.2114
R18022 vdd.n2643 vdd.n963 39.2114
R18023 vdd.n2647 vdd.n964 39.2114
R18024 vdd.n2651 vdd.n965 39.2114
R18025 vdd.n2655 vdd.n966 39.2114
R18026 vdd.n2659 vdd.n967 39.2114
R18027 vdd.n970 vdd.n968 39.2114
R18028 vdd.n2937 vdd.n2700 39.2114
R18029 vdd.n2929 vdd.n2666 39.2114
R18030 vdd.n2925 vdd.n2667 39.2114
R18031 vdd.n2921 vdd.n2668 39.2114
R18032 vdd.n2917 vdd.n2669 39.2114
R18033 vdd.n2913 vdd.n2670 39.2114
R18034 vdd.n2909 vdd.n2671 39.2114
R18035 vdd.n2905 vdd.n2672 39.2114
R18036 vdd.n2901 vdd.n2673 39.2114
R18037 vdd.n2897 vdd.n2674 39.2114
R18038 vdd.n2893 vdd.n2675 39.2114
R18039 vdd.n2889 vdd.n2676 39.2114
R18040 vdd.n2885 vdd.n2677 39.2114
R18041 vdd.n2881 vdd.n2678 39.2114
R18042 vdd.n2877 vdd.n2679 39.2114
R18043 vdd.n2872 vdd.n2680 39.2114
R18044 vdd.n2868 vdd.n2681 39.2114
R18045 vdd.n3089 vdd.n3088 39.2114
R18046 vdd.n835 vdd.n831 39.2114
R18047 vdd.n3097 vdd.n3096 39.2114
R18048 vdd.n830 vdd.n828 39.2114
R18049 vdd.n3104 vdd.n3103 39.2114
R18050 vdd.n827 vdd.n825 39.2114
R18051 vdd.n3111 vdd.n3110 39.2114
R18052 vdd.n824 vdd.n822 39.2114
R18053 vdd.n3118 vdd.n3117 39.2114
R18054 vdd.n3122 vdd.n3121 39.2114
R18055 vdd.n821 vdd.n819 39.2114
R18056 vdd.n3129 vdd.n3128 39.2114
R18057 vdd.n818 vdd.n816 39.2114
R18058 vdd.n3136 vdd.n3135 39.2114
R18059 vdd.n815 vdd.n813 39.2114
R18060 vdd.n3143 vdd.n3142 39.2114
R18061 vdd.n3146 vdd.n3145 39.2114
R18062 vdd.n979 vdd.n934 39.2114
R18063 vdd.n2587 vdd.n935 39.2114
R18064 vdd.n2583 vdd.n936 39.2114
R18065 vdd.n2579 vdd.n937 39.2114
R18066 vdd.n2575 vdd.n938 39.2114
R18067 vdd.n2571 vdd.n939 39.2114
R18068 vdd.n2567 vdd.n940 39.2114
R18069 vdd.n2563 vdd.n941 39.2114
R18070 vdd.n2559 vdd.n942 39.2114
R18071 vdd.n2555 vdd.n943 39.2114
R18072 vdd.n2551 vdd.n944 39.2114
R18073 vdd.n2547 vdd.n945 39.2114
R18074 vdd.n2543 vdd.n946 39.2114
R18075 vdd.n2539 vdd.n947 39.2114
R18076 vdd.n2535 vdd.n948 39.2114
R18077 vdd.n2531 vdd.n949 39.2114
R18078 vdd.n2527 vdd.n950 39.2114
R18079 vdd.n2419 vdd.n2418 39.2114
R18080 vdd.n1222 vdd.n1100 39.2114
R18081 vdd.n1226 vdd.n1101 39.2114
R18082 vdd.n1230 vdd.n1102 39.2114
R18083 vdd.n1234 vdd.n1103 39.2114
R18084 vdd.n1238 vdd.n1104 39.2114
R18085 vdd.n1242 vdd.n1105 39.2114
R18086 vdd.n1246 vdd.n1106 39.2114
R18087 vdd.n1250 vdd.n1107 39.2114
R18088 vdd.n1420 vdd.n1108 39.2114
R18089 vdd.n1417 vdd.n1109 39.2114
R18090 vdd.n1413 vdd.n1110 39.2114
R18091 vdd.n1409 vdd.n1111 39.2114
R18092 vdd.n1405 vdd.n1112 39.2114
R18093 vdd.n1401 vdd.n1113 39.2114
R18094 vdd.n1397 vdd.n1114 39.2114
R18095 vdd.n1393 vdd.n1115 39.2114
R18096 vdd.n2524 vdd.n950 39.2114
R18097 vdd.n2528 vdd.n949 39.2114
R18098 vdd.n2532 vdd.n948 39.2114
R18099 vdd.n2536 vdd.n947 39.2114
R18100 vdd.n2540 vdd.n946 39.2114
R18101 vdd.n2544 vdd.n945 39.2114
R18102 vdd.n2548 vdd.n944 39.2114
R18103 vdd.n2552 vdd.n943 39.2114
R18104 vdd.n2556 vdd.n942 39.2114
R18105 vdd.n2560 vdd.n941 39.2114
R18106 vdd.n2564 vdd.n940 39.2114
R18107 vdd.n2568 vdd.n939 39.2114
R18108 vdd.n2572 vdd.n938 39.2114
R18109 vdd.n2576 vdd.n937 39.2114
R18110 vdd.n2580 vdd.n936 39.2114
R18111 vdd.n2584 vdd.n935 39.2114
R18112 vdd.n2588 vdd.n934 39.2114
R18113 vdd.n2418 vdd.n1082 39.2114
R18114 vdd.n1225 vdd.n1100 39.2114
R18115 vdd.n1229 vdd.n1101 39.2114
R18116 vdd.n1233 vdd.n1102 39.2114
R18117 vdd.n1237 vdd.n1103 39.2114
R18118 vdd.n1241 vdd.n1104 39.2114
R18119 vdd.n1245 vdd.n1105 39.2114
R18120 vdd.n1249 vdd.n1106 39.2114
R18121 vdd.n1252 vdd.n1107 39.2114
R18122 vdd.n1418 vdd.n1108 39.2114
R18123 vdd.n1414 vdd.n1109 39.2114
R18124 vdd.n1410 vdd.n1110 39.2114
R18125 vdd.n1406 vdd.n1111 39.2114
R18126 vdd.n1402 vdd.n1112 39.2114
R18127 vdd.n1398 vdd.n1113 39.2114
R18128 vdd.n1394 vdd.n1114 39.2114
R18129 vdd.n1390 vdd.n1115 39.2114
R18130 vdd.n2271 vdd.n2270 37.2369
R18131 vdd.n2307 vdd.n1191 37.2369
R18132 vdd.n2346 vdd.n1151 37.2369
R18133 vdd.n3230 vdd.n769 37.2369
R18134 vdd.n3278 vdd.n3277 37.2369
R18135 vdd.n690 vdd.n689 37.2369
R18136 vdd.n2414 vdd.n1074 31.0639
R18137 vdd.n2663 vdd.n971 31.0639
R18138 vdd.n2596 vdd.n974 31.0639
R18139 vdd.n1310 vdd.n1307 31.0639
R18140 vdd.n2869 vdd.n2866 31.0639
R18141 vdd.n3086 vdd.n3085 31.0639
R18142 vdd.n2935 vdd.n926 31.0639
R18143 vdd.n3149 vdd.n3148 31.0639
R18144 vdd.n3068 vdd.n3067 31.0639
R18145 vdd.n3154 vdd.n802 31.0639
R18146 vdd.n2773 vdd.n2771 31.0639
R18147 vdd.n2942 vdd.n2941 31.0639
R18148 vdd.n2421 vdd.n2420 31.0639
R18149 vdd.n2591 vdd.n2590 31.0639
R18150 vdd.n2523 vdd.n2522 31.0639
R18151 vdd.n1389 vdd.n1388 31.0639
R18152 vdd.n1255 vdd.n1254 30.449
R18153 vdd.n983 vdd.n982 30.449
R18154 vdd.n1302 vdd.n1274 30.449
R18155 vdd.n2601 vdd.n973 30.449
R18156 vdd.n2706 vdd.n2705 30.449
R18157 vdd.n3092 vdd.n833 30.449
R18158 vdd.n2874 vdd.n2702 30.449
R18159 vdd.n801 vdd.n800 30.449
R18160 vdd.n1780 vdd.n1587 22.2201
R18161 vdd.n2265 vdd.n1083 22.2201
R18162 vdd.n3315 vdd.n723 22.2201
R18163 vdd.n3447 vdd.n3446 22.2201
R18164 vdd.n1791 vdd.n1549 19.3944
R18165 vdd.n1791 vdd.n1547 19.3944
R18166 vdd.n1795 vdd.n1547 19.3944
R18167 vdd.n1795 vdd.n1537 19.3944
R18168 vdd.n1808 vdd.n1537 19.3944
R18169 vdd.n1808 vdd.n1535 19.3944
R18170 vdd.n1812 vdd.n1535 19.3944
R18171 vdd.n1812 vdd.n1527 19.3944
R18172 vdd.n1825 vdd.n1527 19.3944
R18173 vdd.n1825 vdd.n1525 19.3944
R18174 vdd.n1829 vdd.n1525 19.3944
R18175 vdd.n1829 vdd.n1514 19.3944
R18176 vdd.n1841 vdd.n1514 19.3944
R18177 vdd.n1841 vdd.n1512 19.3944
R18178 vdd.n1845 vdd.n1512 19.3944
R18179 vdd.n1845 vdd.n1503 19.3944
R18180 vdd.n1858 vdd.n1503 19.3944
R18181 vdd.n1858 vdd.n1501 19.3944
R18182 vdd.n1862 vdd.n1501 19.3944
R18183 vdd.n1862 vdd.n1492 19.3944
R18184 vdd.n2181 vdd.n1492 19.3944
R18185 vdd.n2181 vdd.n1490 19.3944
R18186 vdd.n2185 vdd.n1490 19.3944
R18187 vdd.n2185 vdd.n1480 19.3944
R18188 vdd.n2198 vdd.n1480 19.3944
R18189 vdd.n2198 vdd.n1478 19.3944
R18190 vdd.n2202 vdd.n1478 19.3944
R18191 vdd.n2202 vdd.n1470 19.3944
R18192 vdd.n2215 vdd.n1470 19.3944
R18193 vdd.n2215 vdd.n1468 19.3944
R18194 vdd.n2219 vdd.n1468 19.3944
R18195 vdd.n2219 vdd.n1457 19.3944
R18196 vdd.n2231 vdd.n1457 19.3944
R18197 vdd.n2231 vdd.n1455 19.3944
R18198 vdd.n2235 vdd.n1455 19.3944
R18199 vdd.n2235 vdd.n1447 19.3944
R18200 vdd.n2248 vdd.n1447 19.3944
R18201 vdd.n2248 vdd.n1444 19.3944
R18202 vdd.n2254 vdd.n1444 19.3944
R18203 vdd.n2254 vdd.n1445 19.3944
R18204 vdd.n1445 vdd.n1435 19.3944
R18205 vdd.n1715 vdd.n1650 19.3944
R18206 vdd.n1711 vdd.n1650 19.3944
R18207 vdd.n1711 vdd.n1710 19.3944
R18208 vdd.n1710 vdd.n1709 19.3944
R18209 vdd.n1709 vdd.n1656 19.3944
R18210 vdd.n1705 vdd.n1656 19.3944
R18211 vdd.n1705 vdd.n1704 19.3944
R18212 vdd.n1704 vdd.n1703 19.3944
R18213 vdd.n1703 vdd.n1662 19.3944
R18214 vdd.n1699 vdd.n1662 19.3944
R18215 vdd.n1699 vdd.n1698 19.3944
R18216 vdd.n1698 vdd.n1697 19.3944
R18217 vdd.n1697 vdd.n1668 19.3944
R18218 vdd.n1693 vdd.n1668 19.3944
R18219 vdd.n1693 vdd.n1692 19.3944
R18220 vdd.n1692 vdd.n1691 19.3944
R18221 vdd.n1691 vdd.n1674 19.3944
R18222 vdd.n1687 vdd.n1674 19.3944
R18223 vdd.n1687 vdd.n1686 19.3944
R18224 vdd.n1686 vdd.n1685 19.3944
R18225 vdd.n1750 vdd.n1749 19.3944
R18226 vdd.n1749 vdd.n1748 19.3944
R18227 vdd.n1748 vdd.n1621 19.3944
R18228 vdd.n1744 vdd.n1621 19.3944
R18229 vdd.n1744 vdd.n1743 19.3944
R18230 vdd.n1743 vdd.n1742 19.3944
R18231 vdd.n1742 vdd.n1627 19.3944
R18232 vdd.n1738 vdd.n1627 19.3944
R18233 vdd.n1738 vdd.n1737 19.3944
R18234 vdd.n1737 vdd.n1736 19.3944
R18235 vdd.n1736 vdd.n1633 19.3944
R18236 vdd.n1732 vdd.n1633 19.3944
R18237 vdd.n1732 vdd.n1731 19.3944
R18238 vdd.n1731 vdd.n1730 19.3944
R18239 vdd.n1730 vdd.n1639 19.3944
R18240 vdd.n1726 vdd.n1639 19.3944
R18241 vdd.n1726 vdd.n1725 19.3944
R18242 vdd.n1725 vdd.n1724 19.3944
R18243 vdd.n1724 vdd.n1645 19.3944
R18244 vdd.n1720 vdd.n1645 19.3944
R18245 vdd.n1783 vdd.n1554 19.3944
R18246 vdd.n1778 vdd.n1554 19.3944
R18247 vdd.n1778 vdd.n1589 19.3944
R18248 vdd.n1774 vdd.n1589 19.3944
R18249 vdd.n1774 vdd.n1773 19.3944
R18250 vdd.n1773 vdd.n1772 19.3944
R18251 vdd.n1772 vdd.n1595 19.3944
R18252 vdd.n1768 vdd.n1595 19.3944
R18253 vdd.n1768 vdd.n1767 19.3944
R18254 vdd.n1767 vdd.n1766 19.3944
R18255 vdd.n1766 vdd.n1601 19.3944
R18256 vdd.n1762 vdd.n1601 19.3944
R18257 vdd.n1762 vdd.n1761 19.3944
R18258 vdd.n1761 vdd.n1760 19.3944
R18259 vdd.n1760 vdd.n1607 19.3944
R18260 vdd.n1756 vdd.n1607 19.3944
R18261 vdd.n1756 vdd.n1755 19.3944
R18262 vdd.n1755 vdd.n1754 19.3944
R18263 vdd.n2303 vdd.n1189 19.3944
R18264 vdd.n2303 vdd.n1195 19.3944
R18265 vdd.n2298 vdd.n1195 19.3944
R18266 vdd.n2298 vdd.n2297 19.3944
R18267 vdd.n2297 vdd.n2296 19.3944
R18268 vdd.n2296 vdd.n1202 19.3944
R18269 vdd.n2291 vdd.n1202 19.3944
R18270 vdd.n2291 vdd.n2290 19.3944
R18271 vdd.n2290 vdd.n2289 19.3944
R18272 vdd.n2289 vdd.n1209 19.3944
R18273 vdd.n2284 vdd.n1209 19.3944
R18274 vdd.n2284 vdd.n2283 19.3944
R18275 vdd.n2283 vdd.n2282 19.3944
R18276 vdd.n2282 vdd.n1216 19.3944
R18277 vdd.n2277 vdd.n1216 19.3944
R18278 vdd.n2277 vdd.n2276 19.3944
R18279 vdd.n1428 vdd.n1221 19.3944
R18280 vdd.n2272 vdd.n1425 19.3944
R18281 vdd.n2342 vdd.n1149 19.3944
R18282 vdd.n2342 vdd.n1155 19.3944
R18283 vdd.n2337 vdd.n1155 19.3944
R18284 vdd.n2337 vdd.n2336 19.3944
R18285 vdd.n2336 vdd.n2335 19.3944
R18286 vdd.n2335 vdd.n1162 19.3944
R18287 vdd.n2330 vdd.n1162 19.3944
R18288 vdd.n2330 vdd.n2329 19.3944
R18289 vdd.n2329 vdd.n2328 19.3944
R18290 vdd.n2328 vdd.n1169 19.3944
R18291 vdd.n2323 vdd.n1169 19.3944
R18292 vdd.n2323 vdd.n2322 19.3944
R18293 vdd.n2322 vdd.n2321 19.3944
R18294 vdd.n2321 vdd.n1176 19.3944
R18295 vdd.n2316 vdd.n1176 19.3944
R18296 vdd.n2316 vdd.n2315 19.3944
R18297 vdd.n2315 vdd.n2314 19.3944
R18298 vdd.n2314 vdd.n1183 19.3944
R18299 vdd.n2309 vdd.n1183 19.3944
R18300 vdd.n2309 vdd.n2308 19.3944
R18301 vdd.n2379 vdd.n1124 19.3944
R18302 vdd.n2379 vdd.n1125 19.3944
R18303 vdd.n2374 vdd.n2373 19.3944
R18304 vdd.n2369 vdd.n2368 19.3944
R18305 vdd.n2368 vdd.n2367 19.3944
R18306 vdd.n2367 vdd.n1129 19.3944
R18307 vdd.n2362 vdd.n1129 19.3944
R18308 vdd.n2362 vdd.n2361 19.3944
R18309 vdd.n2361 vdd.n2360 19.3944
R18310 vdd.n2360 vdd.n1136 19.3944
R18311 vdd.n2355 vdd.n1136 19.3944
R18312 vdd.n2355 vdd.n2354 19.3944
R18313 vdd.n2354 vdd.n2353 19.3944
R18314 vdd.n2353 vdd.n1143 19.3944
R18315 vdd.n2348 vdd.n1143 19.3944
R18316 vdd.n2348 vdd.n2347 19.3944
R18317 vdd.n1787 vdd.n1552 19.3944
R18318 vdd.n1787 vdd.n1543 19.3944
R18319 vdd.n1800 vdd.n1543 19.3944
R18320 vdd.n1800 vdd.n1541 19.3944
R18321 vdd.n1804 vdd.n1541 19.3944
R18322 vdd.n1804 vdd.n1532 19.3944
R18323 vdd.n1817 vdd.n1532 19.3944
R18324 vdd.n1817 vdd.n1530 19.3944
R18325 vdd.n1821 vdd.n1530 19.3944
R18326 vdd.n1821 vdd.n1521 19.3944
R18327 vdd.n1833 vdd.n1521 19.3944
R18328 vdd.n1833 vdd.n1519 19.3944
R18329 vdd.n1837 vdd.n1519 19.3944
R18330 vdd.n1837 vdd.n1509 19.3944
R18331 vdd.n1850 vdd.n1509 19.3944
R18332 vdd.n1850 vdd.n1507 19.3944
R18333 vdd.n1854 vdd.n1507 19.3944
R18334 vdd.n1854 vdd.n1498 19.3944
R18335 vdd.n1866 vdd.n1498 19.3944
R18336 vdd.n1866 vdd.n1496 19.3944
R18337 vdd.n2177 vdd.n1496 19.3944
R18338 vdd.n2177 vdd.n1486 19.3944
R18339 vdd.n2190 vdd.n1486 19.3944
R18340 vdd.n2190 vdd.n1484 19.3944
R18341 vdd.n2194 vdd.n1484 19.3944
R18342 vdd.n2194 vdd.n1475 19.3944
R18343 vdd.n2207 vdd.n1475 19.3944
R18344 vdd.n2207 vdd.n1473 19.3944
R18345 vdd.n2211 vdd.n1473 19.3944
R18346 vdd.n2211 vdd.n1464 19.3944
R18347 vdd.n2223 vdd.n1464 19.3944
R18348 vdd.n2223 vdd.n1462 19.3944
R18349 vdd.n2227 vdd.n1462 19.3944
R18350 vdd.n2227 vdd.n1452 19.3944
R18351 vdd.n2240 vdd.n1452 19.3944
R18352 vdd.n2240 vdd.n1450 19.3944
R18353 vdd.n2244 vdd.n1450 19.3944
R18354 vdd.n2244 vdd.n1440 19.3944
R18355 vdd.n2259 vdd.n1440 19.3944
R18356 vdd.n2259 vdd.n1438 19.3944
R18357 vdd.n2263 vdd.n1438 19.3944
R18358 vdd.n3321 vdd.n686 19.3944
R18359 vdd.n3321 vdd.n676 19.3944
R18360 vdd.n3333 vdd.n676 19.3944
R18361 vdd.n3333 vdd.n674 19.3944
R18362 vdd.n3337 vdd.n674 19.3944
R18363 vdd.n3337 vdd.n666 19.3944
R18364 vdd.n3350 vdd.n666 19.3944
R18365 vdd.n3350 vdd.n664 19.3944
R18366 vdd.n3354 vdd.n664 19.3944
R18367 vdd.n3354 vdd.n653 19.3944
R18368 vdd.n3366 vdd.n653 19.3944
R18369 vdd.n3366 vdd.n651 19.3944
R18370 vdd.n3370 vdd.n651 19.3944
R18371 vdd.n3370 vdd.n642 19.3944
R18372 vdd.n3383 vdd.n642 19.3944
R18373 vdd.n3383 vdd.n640 19.3944
R18374 vdd.n3390 vdd.n640 19.3944
R18375 vdd.n3390 vdd.n3389 19.3944
R18376 vdd.n3389 vdd.n631 19.3944
R18377 vdd.n3403 vdd.n631 19.3944
R18378 vdd.n3404 vdd.n3403 19.3944
R18379 vdd.n3404 vdd.n629 19.3944
R18380 vdd.n3408 vdd.n629 19.3944
R18381 vdd.n3410 vdd.n3408 19.3944
R18382 vdd.n3411 vdd.n3410 19.3944
R18383 vdd.n3411 vdd.n627 19.3944
R18384 vdd.n3415 vdd.n627 19.3944
R18385 vdd.n3417 vdd.n3415 19.3944
R18386 vdd.n3418 vdd.n3417 19.3944
R18387 vdd.n3418 vdd.n625 19.3944
R18388 vdd.n3422 vdd.n625 19.3944
R18389 vdd.n3425 vdd.n3422 19.3944
R18390 vdd.n3426 vdd.n3425 19.3944
R18391 vdd.n3426 vdd.n623 19.3944
R18392 vdd.n3430 vdd.n623 19.3944
R18393 vdd.n3432 vdd.n3430 19.3944
R18394 vdd.n3433 vdd.n3432 19.3944
R18395 vdd.n3433 vdd.n621 19.3944
R18396 vdd.n3437 vdd.n621 19.3944
R18397 vdd.n3439 vdd.n3437 19.3944
R18398 vdd.n3440 vdd.n3439 19.3944
R18399 vdd.n569 vdd.n438 19.3944
R18400 vdd.n575 vdd.n438 19.3944
R18401 vdd.n576 vdd.n575 19.3944
R18402 vdd.n579 vdd.n576 19.3944
R18403 vdd.n579 vdd.n436 19.3944
R18404 vdd.n585 vdd.n436 19.3944
R18405 vdd.n586 vdd.n585 19.3944
R18406 vdd.n589 vdd.n586 19.3944
R18407 vdd.n589 vdd.n434 19.3944
R18408 vdd.n595 vdd.n434 19.3944
R18409 vdd.n596 vdd.n595 19.3944
R18410 vdd.n599 vdd.n596 19.3944
R18411 vdd.n599 vdd.n432 19.3944
R18412 vdd.n605 vdd.n432 19.3944
R18413 vdd.n606 vdd.n605 19.3944
R18414 vdd.n609 vdd.n606 19.3944
R18415 vdd.n609 vdd.n430 19.3944
R18416 vdd.n615 vdd.n430 19.3944
R18417 vdd.n617 vdd.n615 19.3944
R18418 vdd.n618 vdd.n617 19.3944
R18419 vdd.n516 vdd.n515 19.3944
R18420 vdd.n519 vdd.n516 19.3944
R18421 vdd.n519 vdd.n450 19.3944
R18422 vdd.n525 vdd.n450 19.3944
R18423 vdd.n526 vdd.n525 19.3944
R18424 vdd.n529 vdd.n526 19.3944
R18425 vdd.n529 vdd.n448 19.3944
R18426 vdd.n535 vdd.n448 19.3944
R18427 vdd.n536 vdd.n535 19.3944
R18428 vdd.n539 vdd.n536 19.3944
R18429 vdd.n539 vdd.n446 19.3944
R18430 vdd.n545 vdd.n446 19.3944
R18431 vdd.n546 vdd.n545 19.3944
R18432 vdd.n549 vdd.n546 19.3944
R18433 vdd.n549 vdd.n444 19.3944
R18434 vdd.n555 vdd.n444 19.3944
R18435 vdd.n556 vdd.n555 19.3944
R18436 vdd.n559 vdd.n556 19.3944
R18437 vdd.n559 vdd.n442 19.3944
R18438 vdd.n565 vdd.n442 19.3944
R18439 vdd.n466 vdd.n465 19.3944
R18440 vdd.n469 vdd.n466 19.3944
R18441 vdd.n469 vdd.n462 19.3944
R18442 vdd.n475 vdd.n462 19.3944
R18443 vdd.n476 vdd.n475 19.3944
R18444 vdd.n479 vdd.n476 19.3944
R18445 vdd.n479 vdd.n460 19.3944
R18446 vdd.n485 vdd.n460 19.3944
R18447 vdd.n486 vdd.n485 19.3944
R18448 vdd.n489 vdd.n486 19.3944
R18449 vdd.n489 vdd.n458 19.3944
R18450 vdd.n495 vdd.n458 19.3944
R18451 vdd.n496 vdd.n495 19.3944
R18452 vdd.n499 vdd.n496 19.3944
R18453 vdd.n499 vdd.n456 19.3944
R18454 vdd.n505 vdd.n456 19.3944
R18455 vdd.n506 vdd.n505 19.3944
R18456 vdd.n509 vdd.n506 19.3944
R18457 vdd.n3325 vdd.n683 19.3944
R18458 vdd.n3325 vdd.n681 19.3944
R18459 vdd.n3329 vdd.n681 19.3944
R18460 vdd.n3329 vdd.n671 19.3944
R18461 vdd.n3342 vdd.n671 19.3944
R18462 vdd.n3342 vdd.n669 19.3944
R18463 vdd.n3346 vdd.n669 19.3944
R18464 vdd.n3346 vdd.n660 19.3944
R18465 vdd.n3358 vdd.n660 19.3944
R18466 vdd.n3358 vdd.n658 19.3944
R18467 vdd.n3362 vdd.n658 19.3944
R18468 vdd.n3362 vdd.n648 19.3944
R18469 vdd.n3375 vdd.n648 19.3944
R18470 vdd.n3375 vdd.n646 19.3944
R18471 vdd.n3379 vdd.n646 19.3944
R18472 vdd.n3379 vdd.n637 19.3944
R18473 vdd.n3394 vdd.n637 19.3944
R18474 vdd.n3394 vdd.n635 19.3944
R18475 vdd.n3398 vdd.n635 19.3944
R18476 vdd.n3398 vdd.n336 19.3944
R18477 vdd.n3489 vdd.n336 19.3944
R18478 vdd.n3489 vdd.n337 19.3944
R18479 vdd.n3483 vdd.n337 19.3944
R18480 vdd.n3483 vdd.n3482 19.3944
R18481 vdd.n3482 vdd.n3481 19.3944
R18482 vdd.n3481 vdd.n349 19.3944
R18483 vdd.n3475 vdd.n349 19.3944
R18484 vdd.n3475 vdd.n3474 19.3944
R18485 vdd.n3474 vdd.n3473 19.3944
R18486 vdd.n3473 vdd.n359 19.3944
R18487 vdd.n3467 vdd.n359 19.3944
R18488 vdd.n3467 vdd.n3466 19.3944
R18489 vdd.n3466 vdd.n3465 19.3944
R18490 vdd.n3465 vdd.n370 19.3944
R18491 vdd.n3459 vdd.n370 19.3944
R18492 vdd.n3459 vdd.n3458 19.3944
R18493 vdd.n3458 vdd.n3457 19.3944
R18494 vdd.n3457 vdd.n381 19.3944
R18495 vdd.n3451 vdd.n381 19.3944
R18496 vdd.n3451 vdd.n3450 19.3944
R18497 vdd.n3450 vdd.n3449 19.3944
R18498 vdd.n3272 vdd.n747 19.3944
R18499 vdd.n3272 vdd.n3269 19.3944
R18500 vdd.n3269 vdd.n3266 19.3944
R18501 vdd.n3266 vdd.n3265 19.3944
R18502 vdd.n3265 vdd.n3262 19.3944
R18503 vdd.n3262 vdd.n3261 19.3944
R18504 vdd.n3261 vdd.n3258 19.3944
R18505 vdd.n3258 vdd.n3257 19.3944
R18506 vdd.n3257 vdd.n3254 19.3944
R18507 vdd.n3254 vdd.n3253 19.3944
R18508 vdd.n3253 vdd.n3250 19.3944
R18509 vdd.n3250 vdd.n3249 19.3944
R18510 vdd.n3249 vdd.n3246 19.3944
R18511 vdd.n3246 vdd.n3245 19.3944
R18512 vdd.n3245 vdd.n3242 19.3944
R18513 vdd.n3242 vdd.n3241 19.3944
R18514 vdd.n3241 vdd.n3238 19.3944
R18515 vdd.n3238 vdd.n3237 19.3944
R18516 vdd.n3237 vdd.n3234 19.3944
R18517 vdd.n3234 vdd.n3233 19.3944
R18518 vdd.n3312 vdd.n3311 19.3944
R18519 vdd.n3311 vdd.n3310 19.3944
R18520 vdd.n732 vdd.n729 19.3944
R18521 vdd.n3306 vdd.n3305 19.3944
R18522 vdd.n3305 vdd.n3302 19.3944
R18523 vdd.n3302 vdd.n3301 19.3944
R18524 vdd.n3301 vdd.n3298 19.3944
R18525 vdd.n3298 vdd.n3297 19.3944
R18526 vdd.n3297 vdd.n3294 19.3944
R18527 vdd.n3294 vdd.n3293 19.3944
R18528 vdd.n3293 vdd.n3290 19.3944
R18529 vdd.n3290 vdd.n3289 19.3944
R18530 vdd.n3289 vdd.n3286 19.3944
R18531 vdd.n3286 vdd.n3285 19.3944
R18532 vdd.n3285 vdd.n3282 19.3944
R18533 vdd.n3282 vdd.n3281 19.3944
R18534 vdd.n3226 vdd.n767 19.3944
R18535 vdd.n3226 vdd.n3223 19.3944
R18536 vdd.n3223 vdd.n3220 19.3944
R18537 vdd.n3220 vdd.n3219 19.3944
R18538 vdd.n3219 vdd.n3216 19.3944
R18539 vdd.n3216 vdd.n3215 19.3944
R18540 vdd.n3215 vdd.n3212 19.3944
R18541 vdd.n3212 vdd.n3211 19.3944
R18542 vdd.n3211 vdd.n3208 19.3944
R18543 vdd.n3208 vdd.n3207 19.3944
R18544 vdd.n3207 vdd.n3204 19.3944
R18545 vdd.n3204 vdd.n3203 19.3944
R18546 vdd.n3203 vdd.n3200 19.3944
R18547 vdd.n3200 vdd.n3199 19.3944
R18548 vdd.n3199 vdd.n3196 19.3944
R18549 vdd.n3196 vdd.n3195 19.3944
R18550 vdd.n3192 vdd.n3191 19.3944
R18551 vdd.n3188 vdd.n3187 19.3944
R18552 vdd.n1719 vdd.n1715 19.0066
R18553 vdd.n2307 vdd.n1189 19.0066
R18554 vdd.n569 vdd.n566 19.0066
R18555 vdd.n3230 vdd.n767 19.0066
R18556 vdd.n1254 vdd.n1253 16.0975
R18557 vdd.n982 vdd.n981 16.0975
R18558 vdd.n1680 vdd.n1679 16.0975
R18559 vdd.n1718 vdd.n1717 16.0975
R18560 vdd.n1614 vdd.n1613 16.0975
R18561 vdd.n2270 vdd.n2269 16.0975
R18562 vdd.n1191 vdd.n1190 16.0975
R18563 vdd.n1151 vdd.n1150 16.0975
R18564 vdd.n1274 vdd.n1273 16.0975
R18565 vdd.n973 vdd.n972 16.0975
R18566 vdd.n2705 vdd.n2704 16.0975
R18567 vdd.n427 vdd.n426 16.0975
R18568 vdd.n441 vdd.n440 16.0975
R18569 vdd.n453 vdd.n452 16.0975
R18570 vdd.n769 vdd.n768 16.0975
R18571 vdd.n3277 vdd.n3276 16.0975
R18572 vdd.n833 vdd.n832 16.0975
R18573 vdd.n2702 vdd.n2701 16.0975
R18574 vdd.n689 vdd.n688 16.0975
R18575 vdd.n800 vdd.n799 16.0975
R18576 vdd.t209 vdd.n2665 15.4182
R18577 vdd.n2938 vdd.t293 15.4182
R18578 vdd.n28 vdd.n27 14.8356
R18579 vdd.n2417 vdd.n1076 14.0578
R18580 vdd.n3151 vdd.n692 14.0578
R18581 vdd.n328 vdd.n293 13.1884
R18582 vdd.n269 vdd.n234 13.1884
R18583 vdd.n226 vdd.n191 13.1884
R18584 vdd.n167 vdd.n132 13.1884
R18585 vdd.n125 vdd.n90 13.1884
R18586 vdd.n66 vdd.n31 13.1884
R18587 vdd.n2109 vdd.n2074 13.1884
R18588 vdd.n2168 vdd.n2133 13.1884
R18589 vdd.n2007 vdd.n1972 13.1884
R18590 vdd.n2066 vdd.n2031 13.1884
R18591 vdd.n1906 vdd.n1871 13.1884
R18592 vdd.n1965 vdd.n1930 13.1884
R18593 vdd.n1750 vdd.n1615 12.9944
R18594 vdd.n1754 vdd.n1615 12.9944
R18595 vdd.n2346 vdd.n1149 12.9944
R18596 vdd.n2347 vdd.n2346 12.9944
R18597 vdd.n515 vdd.n454 12.9944
R18598 vdd.n509 vdd.n454 12.9944
R18599 vdd.n3278 vdd.n747 12.9944
R18600 vdd.n3281 vdd.n3278 12.9944
R18601 vdd.n329 vdd.n291 12.8005
R18602 vdd.n324 vdd.n295 12.8005
R18603 vdd.n270 vdd.n232 12.8005
R18604 vdd.n265 vdd.n236 12.8005
R18605 vdd.n227 vdd.n189 12.8005
R18606 vdd.n222 vdd.n193 12.8005
R18607 vdd.n168 vdd.n130 12.8005
R18608 vdd.n163 vdd.n134 12.8005
R18609 vdd.n126 vdd.n88 12.8005
R18610 vdd.n121 vdd.n92 12.8005
R18611 vdd.n67 vdd.n29 12.8005
R18612 vdd.n62 vdd.n33 12.8005
R18613 vdd.n2110 vdd.n2072 12.8005
R18614 vdd.n2105 vdd.n2076 12.8005
R18615 vdd.n2169 vdd.n2131 12.8005
R18616 vdd.n2164 vdd.n2135 12.8005
R18617 vdd.n2008 vdd.n1970 12.8005
R18618 vdd.n2003 vdd.n1974 12.8005
R18619 vdd.n2067 vdd.n2029 12.8005
R18620 vdd.n2062 vdd.n2033 12.8005
R18621 vdd.n1907 vdd.n1869 12.8005
R18622 vdd.n1902 vdd.n1873 12.8005
R18623 vdd.n1966 vdd.n1928 12.8005
R18624 vdd.n1961 vdd.n1932 12.8005
R18625 vdd.n323 vdd.n296 12.0247
R18626 vdd.n264 vdd.n237 12.0247
R18627 vdd.n221 vdd.n194 12.0247
R18628 vdd.n162 vdd.n135 12.0247
R18629 vdd.n120 vdd.n93 12.0247
R18630 vdd.n61 vdd.n34 12.0247
R18631 vdd.n2104 vdd.n2077 12.0247
R18632 vdd.n2163 vdd.n2136 12.0247
R18633 vdd.n2002 vdd.n1975 12.0247
R18634 vdd.n2061 vdd.n2034 12.0247
R18635 vdd.n1901 vdd.n1874 12.0247
R18636 vdd.n1960 vdd.n1933 12.0247
R18637 vdd.n1789 vdd.n1545 11.337
R18638 vdd.n1798 vdd.n1545 11.337
R18639 vdd.n1798 vdd.n1797 11.337
R18640 vdd.n1806 vdd.n1539 11.337
R18641 vdd.n1815 vdd.n1814 11.337
R18642 vdd.n1831 vdd.n1523 11.337
R18643 vdd.n1839 vdd.n1516 11.337
R18644 vdd.n1848 vdd.n1847 11.337
R18645 vdd.n1856 vdd.n1505 11.337
R18646 vdd.n2179 vdd.n1494 11.337
R18647 vdd.n2188 vdd.n1488 11.337
R18648 vdd.n2196 vdd.n1482 11.337
R18649 vdd.n2205 vdd.n2204 11.337
R18650 vdd.n2221 vdd.n1466 11.337
R18651 vdd.n2229 vdd.n1459 11.337
R18652 vdd.n2238 vdd.n2237 11.337
R18653 vdd.n2246 vdd.n1442 11.337
R18654 vdd.n2257 vdd.n1442 11.337
R18655 vdd.n2257 vdd.n2256 11.337
R18656 vdd.n3323 vdd.n678 11.337
R18657 vdd.n3331 vdd.n678 11.337
R18658 vdd.n3331 vdd.n679 11.337
R18659 vdd.n3340 vdd.n3339 11.337
R18660 vdd.n3356 vdd.n662 11.337
R18661 vdd.n3364 vdd.n655 11.337
R18662 vdd.n3373 vdd.n3372 11.337
R18663 vdd.n3381 vdd.n644 11.337
R18664 vdd.n3400 vdd.n633 11.337
R18665 vdd.n3487 vdd.n340 11.337
R18666 vdd.n3485 vdd.n344 11.337
R18667 vdd.n3479 vdd.n3478 11.337
R18668 vdd.n3471 vdd.n361 11.337
R18669 vdd.n3470 vdd.n3469 11.337
R18670 vdd.n3463 vdd.n3462 11.337
R18671 vdd.n3461 vdd.n375 11.337
R18672 vdd.n3455 vdd.n3454 11.337
R18673 vdd.n3454 vdd.n3453 11.337
R18674 vdd.n3453 vdd.n386 11.337
R18675 vdd.n320 vdd.n319 11.249
R18676 vdd.n261 vdd.n260 11.249
R18677 vdd.n218 vdd.n217 11.249
R18678 vdd.n159 vdd.n158 11.249
R18679 vdd.n117 vdd.n116 11.249
R18680 vdd.n58 vdd.n57 11.249
R18681 vdd.n2101 vdd.n2100 11.249
R18682 vdd.n2160 vdd.n2159 11.249
R18683 vdd.n1999 vdd.n1998 11.249
R18684 vdd.n2058 vdd.n2057 11.249
R18685 vdd.n1898 vdd.n1897 11.249
R18686 vdd.n1957 vdd.n1956 11.249
R18687 vdd.n1587 vdd.t254 11.2237
R18688 vdd.n3447 vdd.t240 11.2237
R18689 vdd.t97 vdd.n1460 10.7702
R18690 vdd.n3348 vdd.t21 10.7702
R18691 vdd.n305 vdd.n304 10.7238
R18692 vdd.n246 vdd.n245 10.7238
R18693 vdd.n203 vdd.n202 10.7238
R18694 vdd.n144 vdd.n143 10.7238
R18695 vdd.n102 vdd.n101 10.7238
R18696 vdd.n43 vdd.n42 10.7238
R18697 vdd.n2086 vdd.n2085 10.7238
R18698 vdd.n2145 vdd.n2144 10.7238
R18699 vdd.n1984 vdd.n1983 10.7238
R18700 vdd.n2043 vdd.n2042 10.7238
R18701 vdd.n1883 vdd.n1882 10.7238
R18702 vdd.n1942 vdd.n1941 10.7238
R18703 vdd.n2593 vdd.t199 10.6568
R18704 vdd.t196 vdd.n928 10.6568
R18705 vdd.n2426 vdd.n1074 10.6151
R18706 vdd.n2427 vdd.n2426 10.6151
R18707 vdd.n2428 vdd.n2427 10.6151
R18708 vdd.n2428 vdd.n1063 10.6151
R18709 vdd.n2438 vdd.n1063 10.6151
R18710 vdd.n2439 vdd.n2438 10.6151
R18711 vdd.n2440 vdd.n2439 10.6151
R18712 vdd.n2440 vdd.n1050 10.6151
R18713 vdd.n2450 vdd.n1050 10.6151
R18714 vdd.n2451 vdd.n2450 10.6151
R18715 vdd.n2452 vdd.n2451 10.6151
R18716 vdd.n2452 vdd.n1038 10.6151
R18717 vdd.n2463 vdd.n1038 10.6151
R18718 vdd.n2464 vdd.n2463 10.6151
R18719 vdd.n2465 vdd.n2464 10.6151
R18720 vdd.n2465 vdd.n1026 10.6151
R18721 vdd.n2475 vdd.n1026 10.6151
R18722 vdd.n2476 vdd.n2475 10.6151
R18723 vdd.n2477 vdd.n2476 10.6151
R18724 vdd.n2477 vdd.n1014 10.6151
R18725 vdd.n2487 vdd.n1014 10.6151
R18726 vdd.n2488 vdd.n2487 10.6151
R18727 vdd.n2489 vdd.n2488 10.6151
R18728 vdd.n2489 vdd.n1003 10.6151
R18729 vdd.n2499 vdd.n1003 10.6151
R18730 vdd.n2500 vdd.n2499 10.6151
R18731 vdd.n2501 vdd.n2500 10.6151
R18732 vdd.n2501 vdd.n990 10.6151
R18733 vdd.n2513 vdd.n990 10.6151
R18734 vdd.n2514 vdd.n2513 10.6151
R18735 vdd.n2516 vdd.n2514 10.6151
R18736 vdd.n2516 vdd.n2515 10.6151
R18737 vdd.n2515 vdd.n971 10.6151
R18738 vdd.n2663 vdd.n2662 10.6151
R18739 vdd.n2662 vdd.n2661 10.6151
R18740 vdd.n2661 vdd.n2658 10.6151
R18741 vdd.n2658 vdd.n2657 10.6151
R18742 vdd.n2657 vdd.n2654 10.6151
R18743 vdd.n2654 vdd.n2653 10.6151
R18744 vdd.n2653 vdd.n2650 10.6151
R18745 vdd.n2650 vdd.n2649 10.6151
R18746 vdd.n2649 vdd.n2646 10.6151
R18747 vdd.n2646 vdd.n2645 10.6151
R18748 vdd.n2645 vdd.n2642 10.6151
R18749 vdd.n2642 vdd.n2641 10.6151
R18750 vdd.n2641 vdd.n2638 10.6151
R18751 vdd.n2638 vdd.n2637 10.6151
R18752 vdd.n2637 vdd.n2634 10.6151
R18753 vdd.n2634 vdd.n2633 10.6151
R18754 vdd.n2633 vdd.n2630 10.6151
R18755 vdd.n2630 vdd.n2629 10.6151
R18756 vdd.n2629 vdd.n2626 10.6151
R18757 vdd.n2626 vdd.n2625 10.6151
R18758 vdd.n2625 vdd.n2622 10.6151
R18759 vdd.n2622 vdd.n2621 10.6151
R18760 vdd.n2621 vdd.n2618 10.6151
R18761 vdd.n2618 vdd.n2617 10.6151
R18762 vdd.n2617 vdd.n2614 10.6151
R18763 vdd.n2614 vdd.n2613 10.6151
R18764 vdd.n2613 vdd.n2610 10.6151
R18765 vdd.n2610 vdd.n2609 10.6151
R18766 vdd.n2609 vdd.n2606 10.6151
R18767 vdd.n2606 vdd.n2605 10.6151
R18768 vdd.n2605 vdd.n2602 10.6151
R18769 vdd.n2600 vdd.n2597 10.6151
R18770 vdd.n2597 vdd.n2596 10.6151
R18771 vdd.n1311 vdd.n1310 10.6151
R18772 vdd.n1313 vdd.n1311 10.6151
R18773 vdd.n1314 vdd.n1313 10.6151
R18774 vdd.n1316 vdd.n1314 10.6151
R18775 vdd.n1317 vdd.n1316 10.6151
R18776 vdd.n1319 vdd.n1317 10.6151
R18777 vdd.n1320 vdd.n1319 10.6151
R18778 vdd.n1322 vdd.n1320 10.6151
R18779 vdd.n1323 vdd.n1322 10.6151
R18780 vdd.n1325 vdd.n1323 10.6151
R18781 vdd.n1326 vdd.n1325 10.6151
R18782 vdd.n1328 vdd.n1326 10.6151
R18783 vdd.n1329 vdd.n1328 10.6151
R18784 vdd.n1331 vdd.n1329 10.6151
R18785 vdd.n1332 vdd.n1331 10.6151
R18786 vdd.n1334 vdd.n1332 10.6151
R18787 vdd.n1335 vdd.n1334 10.6151
R18788 vdd.n1357 vdd.n1335 10.6151
R18789 vdd.n1357 vdd.n1356 10.6151
R18790 vdd.n1356 vdd.n1355 10.6151
R18791 vdd.n1355 vdd.n1353 10.6151
R18792 vdd.n1353 vdd.n1352 10.6151
R18793 vdd.n1352 vdd.n1350 10.6151
R18794 vdd.n1350 vdd.n1349 10.6151
R18795 vdd.n1349 vdd.n1347 10.6151
R18796 vdd.n1347 vdd.n1346 10.6151
R18797 vdd.n1346 vdd.n1344 10.6151
R18798 vdd.n1344 vdd.n1343 10.6151
R18799 vdd.n1343 vdd.n1341 10.6151
R18800 vdd.n1341 vdd.n1340 10.6151
R18801 vdd.n1340 vdd.n1337 10.6151
R18802 vdd.n1337 vdd.n1336 10.6151
R18803 vdd.n1336 vdd.n974 10.6151
R18804 vdd.n2414 vdd.n2413 10.6151
R18805 vdd.n2413 vdd.n2412 10.6151
R18806 vdd.n2412 vdd.n2411 10.6151
R18807 vdd.n2411 vdd.n2409 10.6151
R18808 vdd.n2409 vdd.n2406 10.6151
R18809 vdd.n2406 vdd.n2405 10.6151
R18810 vdd.n2405 vdd.n2402 10.6151
R18811 vdd.n2402 vdd.n2401 10.6151
R18812 vdd.n2401 vdd.n2398 10.6151
R18813 vdd.n2398 vdd.n2397 10.6151
R18814 vdd.n2397 vdd.n2394 10.6151
R18815 vdd.n2394 vdd.n2393 10.6151
R18816 vdd.n2393 vdd.n2390 10.6151
R18817 vdd.n2390 vdd.n2389 10.6151
R18818 vdd.n2389 vdd.n2386 10.6151
R18819 vdd.n2386 vdd.n2385 10.6151
R18820 vdd.n2385 vdd.n2382 10.6151
R18821 vdd.n2382 vdd.n1119 10.6151
R18822 vdd.n1277 vdd.n1119 10.6151
R18823 vdd.n1278 vdd.n1277 10.6151
R18824 vdd.n1281 vdd.n1278 10.6151
R18825 vdd.n1282 vdd.n1281 10.6151
R18826 vdd.n1285 vdd.n1282 10.6151
R18827 vdd.n1286 vdd.n1285 10.6151
R18828 vdd.n1289 vdd.n1286 10.6151
R18829 vdd.n1290 vdd.n1289 10.6151
R18830 vdd.n1293 vdd.n1290 10.6151
R18831 vdd.n1294 vdd.n1293 10.6151
R18832 vdd.n1297 vdd.n1294 10.6151
R18833 vdd.n1298 vdd.n1297 10.6151
R18834 vdd.n1301 vdd.n1298 10.6151
R18835 vdd.n1306 vdd.n1303 10.6151
R18836 vdd.n1307 vdd.n1306 10.6151
R18837 vdd.n2866 vdd.n2865 10.6151
R18838 vdd.n2865 vdd.n2864 10.6151
R18839 vdd.n2864 vdd.n2703 10.6151
R18840 vdd.n2808 vdd.n2703 10.6151
R18841 vdd.n2809 vdd.n2808 10.6151
R18842 vdd.n2811 vdd.n2809 10.6151
R18843 vdd.n2812 vdd.n2811 10.6151
R18844 vdd.n2814 vdd.n2812 10.6151
R18845 vdd.n2815 vdd.n2814 10.6151
R18846 vdd.n2845 vdd.n2815 10.6151
R18847 vdd.n2845 vdd.n2844 10.6151
R18848 vdd.n2844 vdd.n2843 10.6151
R18849 vdd.n2843 vdd.n2841 10.6151
R18850 vdd.n2841 vdd.n2840 10.6151
R18851 vdd.n2840 vdd.n2838 10.6151
R18852 vdd.n2838 vdd.n2837 10.6151
R18853 vdd.n2837 vdd.n2835 10.6151
R18854 vdd.n2835 vdd.n2834 10.6151
R18855 vdd.n2834 vdd.n2832 10.6151
R18856 vdd.n2832 vdd.n2831 10.6151
R18857 vdd.n2831 vdd.n2829 10.6151
R18858 vdd.n2829 vdd.n2828 10.6151
R18859 vdd.n2828 vdd.n2826 10.6151
R18860 vdd.n2826 vdd.n2825 10.6151
R18861 vdd.n2825 vdd.n2823 10.6151
R18862 vdd.n2823 vdd.n2822 10.6151
R18863 vdd.n2822 vdd.n2820 10.6151
R18864 vdd.n2820 vdd.n2819 10.6151
R18865 vdd.n2819 vdd.n2817 10.6151
R18866 vdd.n2817 vdd.n2816 10.6151
R18867 vdd.n2816 vdd.n836 10.6151
R18868 vdd.n3084 vdd.n836 10.6151
R18869 vdd.n3085 vdd.n3084 10.6151
R18870 vdd.n2935 vdd.n2934 10.6151
R18871 vdd.n2934 vdd.n2933 10.6151
R18872 vdd.n2933 vdd.n2932 10.6151
R18873 vdd.n2932 vdd.n2930 10.6151
R18874 vdd.n2930 vdd.n2927 10.6151
R18875 vdd.n2927 vdd.n2926 10.6151
R18876 vdd.n2926 vdd.n2923 10.6151
R18877 vdd.n2923 vdd.n2922 10.6151
R18878 vdd.n2922 vdd.n2919 10.6151
R18879 vdd.n2919 vdd.n2918 10.6151
R18880 vdd.n2918 vdd.n2915 10.6151
R18881 vdd.n2915 vdd.n2914 10.6151
R18882 vdd.n2914 vdd.n2911 10.6151
R18883 vdd.n2911 vdd.n2910 10.6151
R18884 vdd.n2910 vdd.n2907 10.6151
R18885 vdd.n2907 vdd.n2906 10.6151
R18886 vdd.n2906 vdd.n2903 10.6151
R18887 vdd.n2903 vdd.n2902 10.6151
R18888 vdd.n2902 vdd.n2899 10.6151
R18889 vdd.n2899 vdd.n2898 10.6151
R18890 vdd.n2898 vdd.n2895 10.6151
R18891 vdd.n2895 vdd.n2894 10.6151
R18892 vdd.n2894 vdd.n2891 10.6151
R18893 vdd.n2891 vdd.n2890 10.6151
R18894 vdd.n2890 vdd.n2887 10.6151
R18895 vdd.n2887 vdd.n2886 10.6151
R18896 vdd.n2886 vdd.n2883 10.6151
R18897 vdd.n2883 vdd.n2882 10.6151
R18898 vdd.n2882 vdd.n2879 10.6151
R18899 vdd.n2879 vdd.n2878 10.6151
R18900 vdd.n2878 vdd.n2875 10.6151
R18901 vdd.n2873 vdd.n2870 10.6151
R18902 vdd.n2870 vdd.n2869 10.6151
R18903 vdd.n2947 vdd.n926 10.6151
R18904 vdd.n2948 vdd.n2947 10.6151
R18905 vdd.n2949 vdd.n2948 10.6151
R18906 vdd.n2949 vdd.n915 10.6151
R18907 vdd.n2959 vdd.n915 10.6151
R18908 vdd.n2960 vdd.n2959 10.6151
R18909 vdd.n2961 vdd.n2960 10.6151
R18910 vdd.n2961 vdd.n903 10.6151
R18911 vdd.n2971 vdd.n903 10.6151
R18912 vdd.n2972 vdd.n2971 10.6151
R18913 vdd.n2973 vdd.n2972 10.6151
R18914 vdd.n2973 vdd.n891 10.6151
R18915 vdd.n2983 vdd.n891 10.6151
R18916 vdd.n2984 vdd.n2983 10.6151
R18917 vdd.n2985 vdd.n2984 10.6151
R18918 vdd.n2985 vdd.n880 10.6151
R18919 vdd.n2995 vdd.n880 10.6151
R18920 vdd.n2996 vdd.n2995 10.6151
R18921 vdd.n2997 vdd.n2996 10.6151
R18922 vdd.n2997 vdd.n866 10.6151
R18923 vdd.n3008 vdd.n866 10.6151
R18924 vdd.n3009 vdd.n3008 10.6151
R18925 vdd.n3010 vdd.n3009 10.6151
R18926 vdd.n3010 vdd.n855 10.6151
R18927 vdd.n3020 vdd.n855 10.6151
R18928 vdd.n3021 vdd.n3020 10.6151
R18929 vdd.n3022 vdd.n3021 10.6151
R18930 vdd.n3022 vdd.n841 10.6151
R18931 vdd.n3077 vdd.n841 10.6151
R18932 vdd.n3078 vdd.n3077 10.6151
R18933 vdd.n3079 vdd.n3078 10.6151
R18934 vdd.n3079 vdd.n810 10.6151
R18935 vdd.n3149 vdd.n810 10.6151
R18936 vdd.n3148 vdd.n3147 10.6151
R18937 vdd.n3147 vdd.n811 10.6151
R18938 vdd.n812 vdd.n811 10.6151
R18939 vdd.n3140 vdd.n812 10.6151
R18940 vdd.n3140 vdd.n3139 10.6151
R18941 vdd.n3139 vdd.n3138 10.6151
R18942 vdd.n3138 vdd.n814 10.6151
R18943 vdd.n3133 vdd.n814 10.6151
R18944 vdd.n3133 vdd.n3132 10.6151
R18945 vdd.n3132 vdd.n3131 10.6151
R18946 vdd.n3131 vdd.n817 10.6151
R18947 vdd.n3126 vdd.n817 10.6151
R18948 vdd.n3126 vdd.n3125 10.6151
R18949 vdd.n3125 vdd.n3124 10.6151
R18950 vdd.n3124 vdd.n820 10.6151
R18951 vdd.n3119 vdd.n820 10.6151
R18952 vdd.n3119 vdd.n731 10.6151
R18953 vdd.n3115 vdd.n731 10.6151
R18954 vdd.n3115 vdd.n3114 10.6151
R18955 vdd.n3114 vdd.n3113 10.6151
R18956 vdd.n3113 vdd.n823 10.6151
R18957 vdd.n3108 vdd.n823 10.6151
R18958 vdd.n3108 vdd.n3107 10.6151
R18959 vdd.n3107 vdd.n3106 10.6151
R18960 vdd.n3106 vdd.n826 10.6151
R18961 vdd.n3101 vdd.n826 10.6151
R18962 vdd.n3101 vdd.n3100 10.6151
R18963 vdd.n3100 vdd.n3099 10.6151
R18964 vdd.n3099 vdd.n829 10.6151
R18965 vdd.n3094 vdd.n829 10.6151
R18966 vdd.n3094 vdd.n3093 10.6151
R18967 vdd.n3091 vdd.n834 10.6151
R18968 vdd.n3086 vdd.n834 10.6151
R18969 vdd.n3067 vdd.n3028 10.6151
R18970 vdd.n3062 vdd.n3028 10.6151
R18971 vdd.n3062 vdd.n3061 10.6151
R18972 vdd.n3061 vdd.n3060 10.6151
R18973 vdd.n3060 vdd.n3030 10.6151
R18974 vdd.n3055 vdd.n3030 10.6151
R18975 vdd.n3055 vdd.n3054 10.6151
R18976 vdd.n3054 vdd.n3053 10.6151
R18977 vdd.n3053 vdd.n3033 10.6151
R18978 vdd.n3048 vdd.n3033 10.6151
R18979 vdd.n3048 vdd.n3047 10.6151
R18980 vdd.n3047 vdd.n3046 10.6151
R18981 vdd.n3046 vdd.n3036 10.6151
R18982 vdd.n3041 vdd.n3036 10.6151
R18983 vdd.n3041 vdd.n3040 10.6151
R18984 vdd.n3040 vdd.n785 10.6151
R18985 vdd.n3184 vdd.n785 10.6151
R18986 vdd.n3184 vdd.n786 10.6151
R18987 vdd.n788 vdd.n786 10.6151
R18988 vdd.n3177 vdd.n788 10.6151
R18989 vdd.n3177 vdd.n3176 10.6151
R18990 vdd.n3176 vdd.n3175 10.6151
R18991 vdd.n3175 vdd.n790 10.6151
R18992 vdd.n3170 vdd.n790 10.6151
R18993 vdd.n3170 vdd.n3169 10.6151
R18994 vdd.n3169 vdd.n3168 10.6151
R18995 vdd.n3168 vdd.n793 10.6151
R18996 vdd.n3163 vdd.n793 10.6151
R18997 vdd.n3163 vdd.n3162 10.6151
R18998 vdd.n3162 vdd.n3161 10.6151
R18999 vdd.n3161 vdd.n796 10.6151
R19000 vdd.n3156 vdd.n3155 10.6151
R19001 vdd.n3155 vdd.n3154 10.6151
R19002 vdd.n2774 vdd.n2773 10.6151
R19003 vdd.n2860 vdd.n2774 10.6151
R19004 vdd.n2860 vdd.n2859 10.6151
R19005 vdd.n2859 vdd.n2858 10.6151
R19006 vdd.n2858 vdd.n2856 10.6151
R19007 vdd.n2856 vdd.n2855 10.6151
R19008 vdd.n2855 vdd.n2853 10.6151
R19009 vdd.n2853 vdd.n2852 10.6151
R19010 vdd.n2852 vdd.n2850 10.6151
R19011 vdd.n2850 vdd.n2849 10.6151
R19012 vdd.n2849 vdd.n2806 10.6151
R19013 vdd.n2806 vdd.n2805 10.6151
R19014 vdd.n2805 vdd.n2803 10.6151
R19015 vdd.n2803 vdd.n2802 10.6151
R19016 vdd.n2802 vdd.n2800 10.6151
R19017 vdd.n2800 vdd.n2799 10.6151
R19018 vdd.n2799 vdd.n2797 10.6151
R19019 vdd.n2797 vdd.n2796 10.6151
R19020 vdd.n2796 vdd.n2794 10.6151
R19021 vdd.n2794 vdd.n2793 10.6151
R19022 vdd.n2793 vdd.n2791 10.6151
R19023 vdd.n2791 vdd.n2790 10.6151
R19024 vdd.n2790 vdd.n2788 10.6151
R19025 vdd.n2788 vdd.n2787 10.6151
R19026 vdd.n2787 vdd.n2785 10.6151
R19027 vdd.n2785 vdd.n2784 10.6151
R19028 vdd.n2784 vdd.n2782 10.6151
R19029 vdd.n2782 vdd.n2781 10.6151
R19030 vdd.n2781 vdd.n2779 10.6151
R19031 vdd.n2779 vdd.n2778 10.6151
R19032 vdd.n2778 vdd.n2776 10.6151
R19033 vdd.n2776 vdd.n2775 10.6151
R19034 vdd.n2775 vdd.n802 10.6151
R19035 vdd.n2941 vdd.n932 10.6151
R19036 vdd.n2708 vdd.n932 10.6151
R19037 vdd.n2709 vdd.n2708 10.6151
R19038 vdd.n2712 vdd.n2709 10.6151
R19039 vdd.n2713 vdd.n2712 10.6151
R19040 vdd.n2716 vdd.n2713 10.6151
R19041 vdd.n2717 vdd.n2716 10.6151
R19042 vdd.n2720 vdd.n2717 10.6151
R19043 vdd.n2721 vdd.n2720 10.6151
R19044 vdd.n2724 vdd.n2721 10.6151
R19045 vdd.n2725 vdd.n2724 10.6151
R19046 vdd.n2728 vdd.n2725 10.6151
R19047 vdd.n2729 vdd.n2728 10.6151
R19048 vdd.n2732 vdd.n2729 10.6151
R19049 vdd.n2733 vdd.n2732 10.6151
R19050 vdd.n2736 vdd.n2733 10.6151
R19051 vdd.n2737 vdd.n2736 10.6151
R19052 vdd.n2740 vdd.n2737 10.6151
R19053 vdd.n2741 vdd.n2740 10.6151
R19054 vdd.n2744 vdd.n2741 10.6151
R19055 vdd.n2745 vdd.n2744 10.6151
R19056 vdd.n2748 vdd.n2745 10.6151
R19057 vdd.n2749 vdd.n2748 10.6151
R19058 vdd.n2752 vdd.n2749 10.6151
R19059 vdd.n2753 vdd.n2752 10.6151
R19060 vdd.n2756 vdd.n2753 10.6151
R19061 vdd.n2757 vdd.n2756 10.6151
R19062 vdd.n2760 vdd.n2757 10.6151
R19063 vdd.n2761 vdd.n2760 10.6151
R19064 vdd.n2764 vdd.n2761 10.6151
R19065 vdd.n2765 vdd.n2764 10.6151
R19066 vdd.n2770 vdd.n2768 10.6151
R19067 vdd.n2771 vdd.n2770 10.6151
R19068 vdd.n2943 vdd.n2942 10.6151
R19069 vdd.n2943 vdd.n921 10.6151
R19070 vdd.n2953 vdd.n921 10.6151
R19071 vdd.n2954 vdd.n2953 10.6151
R19072 vdd.n2955 vdd.n2954 10.6151
R19073 vdd.n2955 vdd.n909 10.6151
R19074 vdd.n2965 vdd.n909 10.6151
R19075 vdd.n2966 vdd.n2965 10.6151
R19076 vdd.n2967 vdd.n2966 10.6151
R19077 vdd.n2967 vdd.n897 10.6151
R19078 vdd.n2977 vdd.n897 10.6151
R19079 vdd.n2978 vdd.n2977 10.6151
R19080 vdd.n2979 vdd.n2978 10.6151
R19081 vdd.n2979 vdd.n886 10.6151
R19082 vdd.n2989 vdd.n886 10.6151
R19083 vdd.n2990 vdd.n2989 10.6151
R19084 vdd.n2991 vdd.n2990 10.6151
R19085 vdd.n2991 vdd.n873 10.6151
R19086 vdd.n3001 vdd.n873 10.6151
R19087 vdd.n3002 vdd.n3001 10.6151
R19088 vdd.n3004 vdd.n861 10.6151
R19089 vdd.n3014 vdd.n861 10.6151
R19090 vdd.n3015 vdd.n3014 10.6151
R19091 vdd.n3016 vdd.n3015 10.6151
R19092 vdd.n3016 vdd.n849 10.6151
R19093 vdd.n3026 vdd.n849 10.6151
R19094 vdd.n3027 vdd.n3026 10.6151
R19095 vdd.n3073 vdd.n3027 10.6151
R19096 vdd.n3073 vdd.n3072 10.6151
R19097 vdd.n3072 vdd.n3071 10.6151
R19098 vdd.n3071 vdd.n3070 10.6151
R19099 vdd.n3070 vdd.n3068 10.6151
R19100 vdd.n2422 vdd.n2421 10.6151
R19101 vdd.n2422 vdd.n1069 10.6151
R19102 vdd.n2432 vdd.n1069 10.6151
R19103 vdd.n2433 vdd.n2432 10.6151
R19104 vdd.n2434 vdd.n2433 10.6151
R19105 vdd.n2434 vdd.n1057 10.6151
R19106 vdd.n2444 vdd.n1057 10.6151
R19107 vdd.n2445 vdd.n2444 10.6151
R19108 vdd.n2446 vdd.n2445 10.6151
R19109 vdd.n2446 vdd.n1044 10.6151
R19110 vdd.n2456 vdd.n1044 10.6151
R19111 vdd.n2457 vdd.n2456 10.6151
R19112 vdd.n2459 vdd.n1032 10.6151
R19113 vdd.n2469 vdd.n1032 10.6151
R19114 vdd.n2470 vdd.n2469 10.6151
R19115 vdd.n2471 vdd.n2470 10.6151
R19116 vdd.n2471 vdd.n1020 10.6151
R19117 vdd.n2481 vdd.n1020 10.6151
R19118 vdd.n2482 vdd.n2481 10.6151
R19119 vdd.n2483 vdd.n2482 10.6151
R19120 vdd.n2483 vdd.n1009 10.6151
R19121 vdd.n2493 vdd.n1009 10.6151
R19122 vdd.n2494 vdd.n2493 10.6151
R19123 vdd.n2495 vdd.n2494 10.6151
R19124 vdd.n2495 vdd.n997 10.6151
R19125 vdd.n2505 vdd.n997 10.6151
R19126 vdd.n2506 vdd.n2505 10.6151
R19127 vdd.n2509 vdd.n2506 10.6151
R19128 vdd.n2509 vdd.n2508 10.6151
R19129 vdd.n2508 vdd.n2507 10.6151
R19130 vdd.n2507 vdd.n980 10.6151
R19131 vdd.n2591 vdd.n980 10.6151
R19132 vdd.n2590 vdd.n2589 10.6151
R19133 vdd.n2589 vdd.n2586 10.6151
R19134 vdd.n2586 vdd.n2585 10.6151
R19135 vdd.n2585 vdd.n2582 10.6151
R19136 vdd.n2582 vdd.n2581 10.6151
R19137 vdd.n2581 vdd.n2578 10.6151
R19138 vdd.n2578 vdd.n2577 10.6151
R19139 vdd.n2577 vdd.n2574 10.6151
R19140 vdd.n2574 vdd.n2573 10.6151
R19141 vdd.n2573 vdd.n2570 10.6151
R19142 vdd.n2570 vdd.n2569 10.6151
R19143 vdd.n2569 vdd.n2566 10.6151
R19144 vdd.n2566 vdd.n2565 10.6151
R19145 vdd.n2565 vdd.n2562 10.6151
R19146 vdd.n2562 vdd.n2561 10.6151
R19147 vdd.n2561 vdd.n2558 10.6151
R19148 vdd.n2558 vdd.n2557 10.6151
R19149 vdd.n2557 vdd.n2554 10.6151
R19150 vdd.n2554 vdd.n2553 10.6151
R19151 vdd.n2553 vdd.n2550 10.6151
R19152 vdd.n2550 vdd.n2549 10.6151
R19153 vdd.n2549 vdd.n2546 10.6151
R19154 vdd.n2546 vdd.n2545 10.6151
R19155 vdd.n2545 vdd.n2542 10.6151
R19156 vdd.n2542 vdd.n2541 10.6151
R19157 vdd.n2541 vdd.n2538 10.6151
R19158 vdd.n2538 vdd.n2537 10.6151
R19159 vdd.n2537 vdd.n2534 10.6151
R19160 vdd.n2534 vdd.n2533 10.6151
R19161 vdd.n2533 vdd.n2530 10.6151
R19162 vdd.n2530 vdd.n2529 10.6151
R19163 vdd.n2526 vdd.n2525 10.6151
R19164 vdd.n2525 vdd.n2523 10.6151
R19165 vdd.n1388 vdd.n1386 10.6151
R19166 vdd.n1386 vdd.n1385 10.6151
R19167 vdd.n1385 vdd.n1383 10.6151
R19168 vdd.n1383 vdd.n1382 10.6151
R19169 vdd.n1382 vdd.n1380 10.6151
R19170 vdd.n1380 vdd.n1379 10.6151
R19171 vdd.n1379 vdd.n1377 10.6151
R19172 vdd.n1377 vdd.n1376 10.6151
R19173 vdd.n1376 vdd.n1374 10.6151
R19174 vdd.n1374 vdd.n1373 10.6151
R19175 vdd.n1373 vdd.n1371 10.6151
R19176 vdd.n1371 vdd.n1370 10.6151
R19177 vdd.n1370 vdd.n1368 10.6151
R19178 vdd.n1368 vdd.n1367 10.6151
R19179 vdd.n1367 vdd.n1365 10.6151
R19180 vdd.n1365 vdd.n1364 10.6151
R19181 vdd.n1364 vdd.n1362 10.6151
R19182 vdd.n1362 vdd.n1361 10.6151
R19183 vdd.n1361 vdd.n1272 10.6151
R19184 vdd.n1272 vdd.n1271 10.6151
R19185 vdd.n1271 vdd.n1269 10.6151
R19186 vdd.n1269 vdd.n1268 10.6151
R19187 vdd.n1268 vdd.n1266 10.6151
R19188 vdd.n1266 vdd.n1265 10.6151
R19189 vdd.n1265 vdd.n1263 10.6151
R19190 vdd.n1263 vdd.n1262 10.6151
R19191 vdd.n1262 vdd.n1260 10.6151
R19192 vdd.n1260 vdd.n1259 10.6151
R19193 vdd.n1259 vdd.n1257 10.6151
R19194 vdd.n1257 vdd.n1256 10.6151
R19195 vdd.n1256 vdd.n984 10.6151
R19196 vdd.n2521 vdd.n984 10.6151
R19197 vdd.n2522 vdd.n2521 10.6151
R19198 vdd.n2420 vdd.n1081 10.6151
R19199 vdd.n1223 vdd.n1081 10.6151
R19200 vdd.n1224 vdd.n1223 10.6151
R19201 vdd.n1227 vdd.n1224 10.6151
R19202 vdd.n1228 vdd.n1227 10.6151
R19203 vdd.n1231 vdd.n1228 10.6151
R19204 vdd.n1232 vdd.n1231 10.6151
R19205 vdd.n1235 vdd.n1232 10.6151
R19206 vdd.n1236 vdd.n1235 10.6151
R19207 vdd.n1239 vdd.n1236 10.6151
R19208 vdd.n1240 vdd.n1239 10.6151
R19209 vdd.n1243 vdd.n1240 10.6151
R19210 vdd.n1244 vdd.n1243 10.6151
R19211 vdd.n1247 vdd.n1244 10.6151
R19212 vdd.n1248 vdd.n1247 10.6151
R19213 vdd.n1251 vdd.n1248 10.6151
R19214 vdd.n1422 vdd.n1251 10.6151
R19215 vdd.n1422 vdd.n1421 10.6151
R19216 vdd.n1421 vdd.n1419 10.6151
R19217 vdd.n1419 vdd.n1416 10.6151
R19218 vdd.n1416 vdd.n1415 10.6151
R19219 vdd.n1415 vdd.n1412 10.6151
R19220 vdd.n1412 vdd.n1411 10.6151
R19221 vdd.n1411 vdd.n1408 10.6151
R19222 vdd.n1408 vdd.n1407 10.6151
R19223 vdd.n1407 vdd.n1404 10.6151
R19224 vdd.n1404 vdd.n1403 10.6151
R19225 vdd.n1403 vdd.n1400 10.6151
R19226 vdd.n1400 vdd.n1399 10.6151
R19227 vdd.n1399 vdd.n1396 10.6151
R19228 vdd.n1396 vdd.n1395 10.6151
R19229 vdd.n1392 vdd.n1391 10.6151
R19230 vdd.n1391 vdd.n1389 10.6151
R19231 vdd.n2213 vdd.t33 10.5435
R19232 vdd.n656 vdd.t29 10.5435
R19233 vdd.n316 vdd.n298 10.4732
R19234 vdd.n257 vdd.n239 10.4732
R19235 vdd.n214 vdd.n196 10.4732
R19236 vdd.n155 vdd.n137 10.4732
R19237 vdd.n113 vdd.n95 10.4732
R19238 vdd.n54 vdd.n36 10.4732
R19239 vdd.n2097 vdd.n2079 10.4732
R19240 vdd.n2156 vdd.n2138 10.4732
R19241 vdd.n1995 vdd.n1977 10.4732
R19242 vdd.n2054 vdd.n2036 10.4732
R19243 vdd.n1894 vdd.n1876 10.4732
R19244 vdd.n1953 vdd.n1935 10.4732
R19245 vdd.t60 vdd.n2187 10.3167
R19246 vdd.n3392 vdd.t108 10.3167
R19247 vdd.n1864 vdd.t31 10.09
R19248 vdd.n3486 vdd.t47 10.09
R19249 vdd.t23 vdd.n1517 9.86327
R19250 vdd.n3477 vdd.t105 9.86327
R19251 vdd.n2382 vdd.n2381 9.78206
R19252 vdd.n3308 vdd.n731 9.78206
R19253 vdd.n3185 vdd.n3184 9.78206
R19254 vdd.n2274 vdd.n1422 9.78206
R19255 vdd.n315 vdd.n300 9.69747
R19256 vdd.n256 vdd.n241 9.69747
R19257 vdd.n213 vdd.n198 9.69747
R19258 vdd.n154 vdd.n139 9.69747
R19259 vdd.n112 vdd.n97 9.69747
R19260 vdd.n53 vdd.n38 9.69747
R19261 vdd.n2096 vdd.n2081 9.69747
R19262 vdd.n2155 vdd.n2140 9.69747
R19263 vdd.n1994 vdd.n1979 9.69747
R19264 vdd.n2053 vdd.n2038 9.69747
R19265 vdd.n1893 vdd.n1878 9.69747
R19266 vdd.n1952 vdd.n1937 9.69747
R19267 vdd.n1823 vdd.t111 9.63654
R19268 vdd.n3423 vdd.t77 9.63654
R19269 vdd.n331 vdd.n330 9.45567
R19270 vdd.n272 vdd.n271 9.45567
R19271 vdd.n229 vdd.n228 9.45567
R19272 vdd.n170 vdd.n169 9.45567
R19273 vdd.n128 vdd.n127 9.45567
R19274 vdd.n69 vdd.n68 9.45567
R19275 vdd.n2112 vdd.n2111 9.45567
R19276 vdd.n2171 vdd.n2170 9.45567
R19277 vdd.n2010 vdd.n2009 9.45567
R19278 vdd.n2069 vdd.n2068 9.45567
R19279 vdd.n1909 vdd.n1908 9.45567
R19280 vdd.n1968 vdd.n1967 9.45567
R19281 vdd.n1797 vdd.t73 9.40981
R19282 vdd.n3455 vdd.t37 9.40981
R19283 vdd.n2344 vdd.n1149 9.3005
R19284 vdd.n2343 vdd.n2342 9.3005
R19285 vdd.n1155 vdd.n1154 9.3005
R19286 vdd.n2337 vdd.n1159 9.3005
R19287 vdd.n2336 vdd.n1160 9.3005
R19288 vdd.n2335 vdd.n1161 9.3005
R19289 vdd.n1165 vdd.n1162 9.3005
R19290 vdd.n2330 vdd.n1166 9.3005
R19291 vdd.n2329 vdd.n1167 9.3005
R19292 vdd.n2328 vdd.n1168 9.3005
R19293 vdd.n1172 vdd.n1169 9.3005
R19294 vdd.n2323 vdd.n1173 9.3005
R19295 vdd.n2322 vdd.n1174 9.3005
R19296 vdd.n2321 vdd.n1175 9.3005
R19297 vdd.n1179 vdd.n1176 9.3005
R19298 vdd.n2316 vdd.n1180 9.3005
R19299 vdd.n2315 vdd.n1181 9.3005
R19300 vdd.n2314 vdd.n1182 9.3005
R19301 vdd.n1186 vdd.n1183 9.3005
R19302 vdd.n2309 vdd.n1187 9.3005
R19303 vdd.n2308 vdd.n1188 9.3005
R19304 vdd.n2307 vdd.n2306 9.3005
R19305 vdd.n2305 vdd.n1189 9.3005
R19306 vdd.n2304 vdd.n2303 9.3005
R19307 vdd.n1195 vdd.n1194 9.3005
R19308 vdd.n2298 vdd.n1199 9.3005
R19309 vdd.n2297 vdd.n1200 9.3005
R19310 vdd.n2296 vdd.n1201 9.3005
R19311 vdd.n1205 vdd.n1202 9.3005
R19312 vdd.n2291 vdd.n1206 9.3005
R19313 vdd.n2290 vdd.n1207 9.3005
R19314 vdd.n2289 vdd.n1208 9.3005
R19315 vdd.n1212 vdd.n1209 9.3005
R19316 vdd.n2284 vdd.n1213 9.3005
R19317 vdd.n2283 vdd.n1214 9.3005
R19318 vdd.n2282 vdd.n1215 9.3005
R19319 vdd.n1219 vdd.n1216 9.3005
R19320 vdd.n2277 vdd.n1220 9.3005
R19321 vdd.n2346 vdd.n2345 9.3005
R19322 vdd.n2368 vdd.n1120 9.3005
R19323 vdd.n2367 vdd.n1128 9.3005
R19324 vdd.n1132 vdd.n1129 9.3005
R19325 vdd.n2362 vdd.n1133 9.3005
R19326 vdd.n2361 vdd.n1134 9.3005
R19327 vdd.n2360 vdd.n1135 9.3005
R19328 vdd.n1139 vdd.n1136 9.3005
R19329 vdd.n2355 vdd.n1140 9.3005
R19330 vdd.n2354 vdd.n1141 9.3005
R19331 vdd.n2353 vdd.n1142 9.3005
R19332 vdd.n1146 vdd.n1143 9.3005
R19333 vdd.n2348 vdd.n1147 9.3005
R19334 vdd.n2347 vdd.n1148 9.3005
R19335 vdd.n2380 vdd.n2379 9.3005
R19336 vdd.n1124 vdd.n1123 9.3005
R19337 vdd.n2177 vdd.n2176 9.3005
R19338 vdd.n1486 vdd.n1485 9.3005
R19339 vdd.n2191 vdd.n2190 9.3005
R19340 vdd.n2192 vdd.n1484 9.3005
R19341 vdd.n2194 vdd.n2193 9.3005
R19342 vdd.n1475 vdd.n1474 9.3005
R19343 vdd.n2208 vdd.n2207 9.3005
R19344 vdd.n2209 vdd.n1473 9.3005
R19345 vdd.n2211 vdd.n2210 9.3005
R19346 vdd.n1464 vdd.n1463 9.3005
R19347 vdd.n2224 vdd.n2223 9.3005
R19348 vdd.n2225 vdd.n1462 9.3005
R19349 vdd.n2227 vdd.n2226 9.3005
R19350 vdd.n1452 vdd.n1451 9.3005
R19351 vdd.n2241 vdd.n2240 9.3005
R19352 vdd.n2242 vdd.n1450 9.3005
R19353 vdd.n2244 vdd.n2243 9.3005
R19354 vdd.n1440 vdd.n1439 9.3005
R19355 vdd.n2260 vdd.n2259 9.3005
R19356 vdd.n2261 vdd.n1438 9.3005
R19357 vdd.n2263 vdd.n2262 9.3005
R19358 vdd.n307 vdd.n306 9.3005
R19359 vdd.n302 vdd.n301 9.3005
R19360 vdd.n313 vdd.n312 9.3005
R19361 vdd.n315 vdd.n314 9.3005
R19362 vdd.n298 vdd.n297 9.3005
R19363 vdd.n321 vdd.n320 9.3005
R19364 vdd.n323 vdd.n322 9.3005
R19365 vdd.n295 vdd.n292 9.3005
R19366 vdd.n330 vdd.n329 9.3005
R19367 vdd.n248 vdd.n247 9.3005
R19368 vdd.n243 vdd.n242 9.3005
R19369 vdd.n254 vdd.n253 9.3005
R19370 vdd.n256 vdd.n255 9.3005
R19371 vdd.n239 vdd.n238 9.3005
R19372 vdd.n262 vdd.n261 9.3005
R19373 vdd.n264 vdd.n263 9.3005
R19374 vdd.n236 vdd.n233 9.3005
R19375 vdd.n271 vdd.n270 9.3005
R19376 vdd.n205 vdd.n204 9.3005
R19377 vdd.n200 vdd.n199 9.3005
R19378 vdd.n211 vdd.n210 9.3005
R19379 vdd.n213 vdd.n212 9.3005
R19380 vdd.n196 vdd.n195 9.3005
R19381 vdd.n219 vdd.n218 9.3005
R19382 vdd.n221 vdd.n220 9.3005
R19383 vdd.n193 vdd.n190 9.3005
R19384 vdd.n228 vdd.n227 9.3005
R19385 vdd.n146 vdd.n145 9.3005
R19386 vdd.n141 vdd.n140 9.3005
R19387 vdd.n152 vdd.n151 9.3005
R19388 vdd.n154 vdd.n153 9.3005
R19389 vdd.n137 vdd.n136 9.3005
R19390 vdd.n160 vdd.n159 9.3005
R19391 vdd.n162 vdd.n161 9.3005
R19392 vdd.n134 vdd.n131 9.3005
R19393 vdd.n169 vdd.n168 9.3005
R19394 vdd.n104 vdd.n103 9.3005
R19395 vdd.n99 vdd.n98 9.3005
R19396 vdd.n110 vdd.n109 9.3005
R19397 vdd.n112 vdd.n111 9.3005
R19398 vdd.n95 vdd.n94 9.3005
R19399 vdd.n118 vdd.n117 9.3005
R19400 vdd.n120 vdd.n119 9.3005
R19401 vdd.n92 vdd.n89 9.3005
R19402 vdd.n127 vdd.n126 9.3005
R19403 vdd.n45 vdd.n44 9.3005
R19404 vdd.n40 vdd.n39 9.3005
R19405 vdd.n51 vdd.n50 9.3005
R19406 vdd.n53 vdd.n52 9.3005
R19407 vdd.n36 vdd.n35 9.3005
R19408 vdd.n59 vdd.n58 9.3005
R19409 vdd.n61 vdd.n60 9.3005
R19410 vdd.n33 vdd.n30 9.3005
R19411 vdd.n68 vdd.n67 9.3005
R19412 vdd.n3230 vdd.n3229 9.3005
R19413 vdd.n3233 vdd.n766 9.3005
R19414 vdd.n3234 vdd.n765 9.3005
R19415 vdd.n3237 vdd.n764 9.3005
R19416 vdd.n3238 vdd.n763 9.3005
R19417 vdd.n3241 vdd.n762 9.3005
R19418 vdd.n3242 vdd.n761 9.3005
R19419 vdd.n3245 vdd.n760 9.3005
R19420 vdd.n3246 vdd.n759 9.3005
R19421 vdd.n3249 vdd.n758 9.3005
R19422 vdd.n3250 vdd.n757 9.3005
R19423 vdd.n3253 vdd.n756 9.3005
R19424 vdd.n3254 vdd.n755 9.3005
R19425 vdd.n3257 vdd.n754 9.3005
R19426 vdd.n3258 vdd.n753 9.3005
R19427 vdd.n3261 vdd.n752 9.3005
R19428 vdd.n3262 vdd.n751 9.3005
R19429 vdd.n3265 vdd.n750 9.3005
R19430 vdd.n3266 vdd.n749 9.3005
R19431 vdd.n3269 vdd.n748 9.3005
R19432 vdd.n3273 vdd.n3272 9.3005
R19433 vdd.n3274 vdd.n747 9.3005
R19434 vdd.n3278 vdd.n3275 9.3005
R19435 vdd.n3281 vdd.n746 9.3005
R19436 vdd.n3282 vdd.n745 9.3005
R19437 vdd.n3285 vdd.n744 9.3005
R19438 vdd.n3286 vdd.n743 9.3005
R19439 vdd.n3289 vdd.n742 9.3005
R19440 vdd.n3290 vdd.n741 9.3005
R19441 vdd.n3293 vdd.n740 9.3005
R19442 vdd.n3294 vdd.n739 9.3005
R19443 vdd.n3297 vdd.n738 9.3005
R19444 vdd.n3298 vdd.n737 9.3005
R19445 vdd.n3301 vdd.n736 9.3005
R19446 vdd.n3302 vdd.n735 9.3005
R19447 vdd.n3305 vdd.n730 9.3005
R19448 vdd.n3311 vdd.n727 9.3005
R19449 vdd.n3312 vdd.n726 9.3005
R19450 vdd.n3326 vdd.n3325 9.3005
R19451 vdd.n3327 vdd.n681 9.3005
R19452 vdd.n3329 vdd.n3328 9.3005
R19453 vdd.n671 vdd.n670 9.3005
R19454 vdd.n3343 vdd.n3342 9.3005
R19455 vdd.n3344 vdd.n669 9.3005
R19456 vdd.n3346 vdd.n3345 9.3005
R19457 vdd.n660 vdd.n659 9.3005
R19458 vdd.n3359 vdd.n3358 9.3005
R19459 vdd.n3360 vdd.n658 9.3005
R19460 vdd.n3362 vdd.n3361 9.3005
R19461 vdd.n648 vdd.n647 9.3005
R19462 vdd.n3376 vdd.n3375 9.3005
R19463 vdd.n3377 vdd.n646 9.3005
R19464 vdd.n3379 vdd.n3378 9.3005
R19465 vdd.n637 vdd.n636 9.3005
R19466 vdd.n3395 vdd.n3394 9.3005
R19467 vdd.n3396 vdd.n635 9.3005
R19468 vdd.n3398 vdd.n3397 9.3005
R19469 vdd.n336 vdd.n334 9.3005
R19470 vdd.n683 vdd.n682 9.3005
R19471 vdd.n3490 vdd.n3489 9.3005
R19472 vdd.n337 vdd.n335 9.3005
R19473 vdd.n3483 vdd.n346 9.3005
R19474 vdd.n3482 vdd.n347 9.3005
R19475 vdd.n3481 vdd.n348 9.3005
R19476 vdd.n355 vdd.n349 9.3005
R19477 vdd.n3475 vdd.n356 9.3005
R19478 vdd.n3474 vdd.n357 9.3005
R19479 vdd.n3473 vdd.n358 9.3005
R19480 vdd.n366 vdd.n359 9.3005
R19481 vdd.n3467 vdd.n367 9.3005
R19482 vdd.n3466 vdd.n368 9.3005
R19483 vdd.n3465 vdd.n369 9.3005
R19484 vdd.n377 vdd.n370 9.3005
R19485 vdd.n3459 vdd.n378 9.3005
R19486 vdd.n3458 vdd.n379 9.3005
R19487 vdd.n3457 vdd.n380 9.3005
R19488 vdd.n388 vdd.n381 9.3005
R19489 vdd.n3451 vdd.n389 9.3005
R19490 vdd.n3450 vdd.n390 9.3005
R19491 vdd.n3449 vdd.n391 9.3005
R19492 vdd.n466 vdd.n463 9.3005
R19493 vdd.n470 vdd.n469 9.3005
R19494 vdd.n471 vdd.n462 9.3005
R19495 vdd.n475 vdd.n472 9.3005
R19496 vdd.n476 vdd.n461 9.3005
R19497 vdd.n480 vdd.n479 9.3005
R19498 vdd.n481 vdd.n460 9.3005
R19499 vdd.n485 vdd.n482 9.3005
R19500 vdd.n486 vdd.n459 9.3005
R19501 vdd.n490 vdd.n489 9.3005
R19502 vdd.n491 vdd.n458 9.3005
R19503 vdd.n495 vdd.n492 9.3005
R19504 vdd.n496 vdd.n457 9.3005
R19505 vdd.n500 vdd.n499 9.3005
R19506 vdd.n501 vdd.n456 9.3005
R19507 vdd.n505 vdd.n502 9.3005
R19508 vdd.n506 vdd.n455 9.3005
R19509 vdd.n510 vdd.n509 9.3005
R19510 vdd.n511 vdd.n454 9.3005
R19511 vdd.n515 vdd.n512 9.3005
R19512 vdd.n516 vdd.n451 9.3005
R19513 vdd.n520 vdd.n519 9.3005
R19514 vdd.n521 vdd.n450 9.3005
R19515 vdd.n525 vdd.n522 9.3005
R19516 vdd.n526 vdd.n449 9.3005
R19517 vdd.n530 vdd.n529 9.3005
R19518 vdd.n531 vdd.n448 9.3005
R19519 vdd.n535 vdd.n532 9.3005
R19520 vdd.n536 vdd.n447 9.3005
R19521 vdd.n540 vdd.n539 9.3005
R19522 vdd.n541 vdd.n446 9.3005
R19523 vdd.n545 vdd.n542 9.3005
R19524 vdd.n546 vdd.n445 9.3005
R19525 vdd.n550 vdd.n549 9.3005
R19526 vdd.n551 vdd.n444 9.3005
R19527 vdd.n555 vdd.n552 9.3005
R19528 vdd.n556 vdd.n443 9.3005
R19529 vdd.n560 vdd.n559 9.3005
R19530 vdd.n561 vdd.n442 9.3005
R19531 vdd.n565 vdd.n562 9.3005
R19532 vdd.n566 vdd.n439 9.3005
R19533 vdd.n570 vdd.n569 9.3005
R19534 vdd.n571 vdd.n438 9.3005
R19535 vdd.n575 vdd.n572 9.3005
R19536 vdd.n576 vdd.n437 9.3005
R19537 vdd.n580 vdd.n579 9.3005
R19538 vdd.n581 vdd.n436 9.3005
R19539 vdd.n585 vdd.n582 9.3005
R19540 vdd.n586 vdd.n435 9.3005
R19541 vdd.n590 vdd.n589 9.3005
R19542 vdd.n591 vdd.n434 9.3005
R19543 vdd.n595 vdd.n592 9.3005
R19544 vdd.n596 vdd.n433 9.3005
R19545 vdd.n600 vdd.n599 9.3005
R19546 vdd.n601 vdd.n432 9.3005
R19547 vdd.n605 vdd.n602 9.3005
R19548 vdd.n606 vdd.n431 9.3005
R19549 vdd.n610 vdd.n609 9.3005
R19550 vdd.n611 vdd.n430 9.3005
R19551 vdd.n615 vdd.n612 9.3005
R19552 vdd.n617 vdd.n429 9.3005
R19553 vdd.n619 vdd.n618 9.3005
R19554 vdd.n3443 vdd.n3442 9.3005
R19555 vdd.n465 vdd.n464 9.3005
R19556 vdd.n3321 vdd.n3320 9.3005
R19557 vdd.n676 vdd.n675 9.3005
R19558 vdd.n3334 vdd.n3333 9.3005
R19559 vdd.n3335 vdd.n674 9.3005
R19560 vdd.n3337 vdd.n3336 9.3005
R19561 vdd.n666 vdd.n665 9.3005
R19562 vdd.n3351 vdd.n3350 9.3005
R19563 vdd.n3352 vdd.n664 9.3005
R19564 vdd.n3354 vdd.n3353 9.3005
R19565 vdd.n653 vdd.n652 9.3005
R19566 vdd.n3367 vdd.n3366 9.3005
R19567 vdd.n3368 vdd.n651 9.3005
R19568 vdd.n3370 vdd.n3369 9.3005
R19569 vdd.n642 vdd.n641 9.3005
R19570 vdd.n3384 vdd.n3383 9.3005
R19571 vdd.n3385 vdd.n640 9.3005
R19572 vdd.n3390 vdd.n3386 9.3005
R19573 vdd.n3389 vdd.n3388 9.3005
R19574 vdd.n3387 vdd.n631 9.3005
R19575 vdd.n3403 vdd.n630 9.3005
R19576 vdd.n3405 vdd.n3404 9.3005
R19577 vdd.n3406 vdd.n629 9.3005
R19578 vdd.n3408 vdd.n3407 9.3005
R19579 vdd.n3410 vdd.n628 9.3005
R19580 vdd.n3412 vdd.n3411 9.3005
R19581 vdd.n3413 vdd.n627 9.3005
R19582 vdd.n3415 vdd.n3414 9.3005
R19583 vdd.n3417 vdd.n626 9.3005
R19584 vdd.n3419 vdd.n3418 9.3005
R19585 vdd.n3420 vdd.n625 9.3005
R19586 vdd.n3422 vdd.n3421 9.3005
R19587 vdd.n3425 vdd.n624 9.3005
R19588 vdd.n3427 vdd.n3426 9.3005
R19589 vdd.n3428 vdd.n623 9.3005
R19590 vdd.n3430 vdd.n3429 9.3005
R19591 vdd.n3432 vdd.n622 9.3005
R19592 vdd.n3434 vdd.n3433 9.3005
R19593 vdd.n3435 vdd.n621 9.3005
R19594 vdd.n3437 vdd.n3436 9.3005
R19595 vdd.n3439 vdd.n620 9.3005
R19596 vdd.n3441 vdd.n3440 9.3005
R19597 vdd.n3319 vdd.n686 9.3005
R19598 vdd.n3318 vdd.n3317 9.3005
R19599 vdd.n3187 vdd.n687 9.3005
R19600 vdd.n3196 vdd.n783 9.3005
R19601 vdd.n3199 vdd.n782 9.3005
R19602 vdd.n3200 vdd.n781 9.3005
R19603 vdd.n3203 vdd.n780 9.3005
R19604 vdd.n3204 vdd.n779 9.3005
R19605 vdd.n3207 vdd.n778 9.3005
R19606 vdd.n3208 vdd.n777 9.3005
R19607 vdd.n3211 vdd.n776 9.3005
R19608 vdd.n3212 vdd.n775 9.3005
R19609 vdd.n3215 vdd.n774 9.3005
R19610 vdd.n3216 vdd.n773 9.3005
R19611 vdd.n3219 vdd.n772 9.3005
R19612 vdd.n3220 vdd.n771 9.3005
R19613 vdd.n3223 vdd.n770 9.3005
R19614 vdd.n3227 vdd.n3226 9.3005
R19615 vdd.n3228 vdd.n767 9.3005
R19616 vdd.n2273 vdd.n2272 9.3005
R19617 vdd.n2268 vdd.n1424 9.3005
R19618 vdd.n1792 vdd.n1791 9.3005
R19619 vdd.n1793 vdd.n1547 9.3005
R19620 vdd.n1795 vdd.n1794 9.3005
R19621 vdd.n1537 vdd.n1536 9.3005
R19622 vdd.n1809 vdd.n1808 9.3005
R19623 vdd.n1810 vdd.n1535 9.3005
R19624 vdd.n1812 vdd.n1811 9.3005
R19625 vdd.n1527 vdd.n1526 9.3005
R19626 vdd.n1826 vdd.n1825 9.3005
R19627 vdd.n1827 vdd.n1525 9.3005
R19628 vdd.n1829 vdd.n1828 9.3005
R19629 vdd.n1514 vdd.n1513 9.3005
R19630 vdd.n1842 vdd.n1841 9.3005
R19631 vdd.n1843 vdd.n1512 9.3005
R19632 vdd.n1845 vdd.n1844 9.3005
R19633 vdd.n1503 vdd.n1502 9.3005
R19634 vdd.n1859 vdd.n1858 9.3005
R19635 vdd.n1860 vdd.n1501 9.3005
R19636 vdd.n1862 vdd.n1861 9.3005
R19637 vdd.n1492 vdd.n1491 9.3005
R19638 vdd.n2182 vdd.n2181 9.3005
R19639 vdd.n2183 vdd.n1490 9.3005
R19640 vdd.n2185 vdd.n2184 9.3005
R19641 vdd.n1480 vdd.n1479 9.3005
R19642 vdd.n2199 vdd.n2198 9.3005
R19643 vdd.n2200 vdd.n1478 9.3005
R19644 vdd.n2202 vdd.n2201 9.3005
R19645 vdd.n1470 vdd.n1469 9.3005
R19646 vdd.n2216 vdd.n2215 9.3005
R19647 vdd.n2217 vdd.n1468 9.3005
R19648 vdd.n2219 vdd.n2218 9.3005
R19649 vdd.n1457 vdd.n1456 9.3005
R19650 vdd.n2232 vdd.n2231 9.3005
R19651 vdd.n2233 vdd.n1455 9.3005
R19652 vdd.n2235 vdd.n2234 9.3005
R19653 vdd.n1447 vdd.n1446 9.3005
R19654 vdd.n2249 vdd.n2248 9.3005
R19655 vdd.n2250 vdd.n1444 9.3005
R19656 vdd.n2254 vdd.n2253 9.3005
R19657 vdd.n2252 vdd.n1445 9.3005
R19658 vdd.n2251 vdd.n1435 9.3005
R19659 vdd.n1549 vdd.n1548 9.3005
R19660 vdd.n1685 vdd.n1684 9.3005
R19661 vdd.n1686 vdd.n1675 9.3005
R19662 vdd.n1688 vdd.n1687 9.3005
R19663 vdd.n1689 vdd.n1674 9.3005
R19664 vdd.n1691 vdd.n1690 9.3005
R19665 vdd.n1692 vdd.n1669 9.3005
R19666 vdd.n1694 vdd.n1693 9.3005
R19667 vdd.n1695 vdd.n1668 9.3005
R19668 vdd.n1697 vdd.n1696 9.3005
R19669 vdd.n1698 vdd.n1663 9.3005
R19670 vdd.n1700 vdd.n1699 9.3005
R19671 vdd.n1701 vdd.n1662 9.3005
R19672 vdd.n1703 vdd.n1702 9.3005
R19673 vdd.n1704 vdd.n1657 9.3005
R19674 vdd.n1706 vdd.n1705 9.3005
R19675 vdd.n1707 vdd.n1656 9.3005
R19676 vdd.n1709 vdd.n1708 9.3005
R19677 vdd.n1710 vdd.n1651 9.3005
R19678 vdd.n1712 vdd.n1711 9.3005
R19679 vdd.n1713 vdd.n1650 9.3005
R19680 vdd.n1715 vdd.n1714 9.3005
R19681 vdd.n1719 vdd.n1646 9.3005
R19682 vdd.n1721 vdd.n1720 9.3005
R19683 vdd.n1722 vdd.n1645 9.3005
R19684 vdd.n1724 vdd.n1723 9.3005
R19685 vdd.n1725 vdd.n1640 9.3005
R19686 vdd.n1727 vdd.n1726 9.3005
R19687 vdd.n1728 vdd.n1639 9.3005
R19688 vdd.n1730 vdd.n1729 9.3005
R19689 vdd.n1731 vdd.n1634 9.3005
R19690 vdd.n1733 vdd.n1732 9.3005
R19691 vdd.n1734 vdd.n1633 9.3005
R19692 vdd.n1736 vdd.n1735 9.3005
R19693 vdd.n1737 vdd.n1628 9.3005
R19694 vdd.n1739 vdd.n1738 9.3005
R19695 vdd.n1740 vdd.n1627 9.3005
R19696 vdd.n1742 vdd.n1741 9.3005
R19697 vdd.n1743 vdd.n1622 9.3005
R19698 vdd.n1745 vdd.n1744 9.3005
R19699 vdd.n1746 vdd.n1621 9.3005
R19700 vdd.n1748 vdd.n1747 9.3005
R19701 vdd.n1749 vdd.n1616 9.3005
R19702 vdd.n1751 vdd.n1750 9.3005
R19703 vdd.n1752 vdd.n1615 9.3005
R19704 vdd.n1754 vdd.n1753 9.3005
R19705 vdd.n1755 vdd.n1608 9.3005
R19706 vdd.n1757 vdd.n1756 9.3005
R19707 vdd.n1758 vdd.n1607 9.3005
R19708 vdd.n1760 vdd.n1759 9.3005
R19709 vdd.n1761 vdd.n1602 9.3005
R19710 vdd.n1763 vdd.n1762 9.3005
R19711 vdd.n1764 vdd.n1601 9.3005
R19712 vdd.n1766 vdd.n1765 9.3005
R19713 vdd.n1767 vdd.n1596 9.3005
R19714 vdd.n1769 vdd.n1768 9.3005
R19715 vdd.n1770 vdd.n1595 9.3005
R19716 vdd.n1772 vdd.n1771 9.3005
R19717 vdd.n1773 vdd.n1590 9.3005
R19718 vdd.n1775 vdd.n1774 9.3005
R19719 vdd.n1776 vdd.n1589 9.3005
R19720 vdd.n1778 vdd.n1777 9.3005
R19721 vdd.n1554 vdd.n1553 9.3005
R19722 vdd.n1784 vdd.n1783 9.3005
R19723 vdd.n1683 vdd.n1682 9.3005
R19724 vdd.n1787 vdd.n1786 9.3005
R19725 vdd.n1543 vdd.n1542 9.3005
R19726 vdd.n1801 vdd.n1800 9.3005
R19727 vdd.n1802 vdd.n1541 9.3005
R19728 vdd.n1804 vdd.n1803 9.3005
R19729 vdd.n1532 vdd.n1531 9.3005
R19730 vdd.n1818 vdd.n1817 9.3005
R19731 vdd.n1819 vdd.n1530 9.3005
R19732 vdd.n1821 vdd.n1820 9.3005
R19733 vdd.n1521 vdd.n1520 9.3005
R19734 vdd.n1834 vdd.n1833 9.3005
R19735 vdd.n1835 vdd.n1519 9.3005
R19736 vdd.n1837 vdd.n1836 9.3005
R19737 vdd.n1509 vdd.n1508 9.3005
R19738 vdd.n1851 vdd.n1850 9.3005
R19739 vdd.n1852 vdd.n1507 9.3005
R19740 vdd.n1854 vdd.n1853 9.3005
R19741 vdd.n1498 vdd.n1497 9.3005
R19742 vdd.n1867 vdd.n1866 9.3005
R19743 vdd.n1868 vdd.n1496 9.3005
R19744 vdd.n1785 vdd.n1552 9.3005
R19745 vdd.n2088 vdd.n2087 9.3005
R19746 vdd.n2083 vdd.n2082 9.3005
R19747 vdd.n2094 vdd.n2093 9.3005
R19748 vdd.n2096 vdd.n2095 9.3005
R19749 vdd.n2079 vdd.n2078 9.3005
R19750 vdd.n2102 vdd.n2101 9.3005
R19751 vdd.n2104 vdd.n2103 9.3005
R19752 vdd.n2076 vdd.n2073 9.3005
R19753 vdd.n2111 vdd.n2110 9.3005
R19754 vdd.n2147 vdd.n2146 9.3005
R19755 vdd.n2142 vdd.n2141 9.3005
R19756 vdd.n2153 vdd.n2152 9.3005
R19757 vdd.n2155 vdd.n2154 9.3005
R19758 vdd.n2138 vdd.n2137 9.3005
R19759 vdd.n2161 vdd.n2160 9.3005
R19760 vdd.n2163 vdd.n2162 9.3005
R19761 vdd.n2135 vdd.n2132 9.3005
R19762 vdd.n2170 vdd.n2169 9.3005
R19763 vdd.n1986 vdd.n1985 9.3005
R19764 vdd.n1981 vdd.n1980 9.3005
R19765 vdd.n1992 vdd.n1991 9.3005
R19766 vdd.n1994 vdd.n1993 9.3005
R19767 vdd.n1977 vdd.n1976 9.3005
R19768 vdd.n2000 vdd.n1999 9.3005
R19769 vdd.n2002 vdd.n2001 9.3005
R19770 vdd.n1974 vdd.n1971 9.3005
R19771 vdd.n2009 vdd.n2008 9.3005
R19772 vdd.n2045 vdd.n2044 9.3005
R19773 vdd.n2040 vdd.n2039 9.3005
R19774 vdd.n2051 vdd.n2050 9.3005
R19775 vdd.n2053 vdd.n2052 9.3005
R19776 vdd.n2036 vdd.n2035 9.3005
R19777 vdd.n2059 vdd.n2058 9.3005
R19778 vdd.n2061 vdd.n2060 9.3005
R19779 vdd.n2033 vdd.n2030 9.3005
R19780 vdd.n2068 vdd.n2067 9.3005
R19781 vdd.n1885 vdd.n1884 9.3005
R19782 vdd.n1880 vdd.n1879 9.3005
R19783 vdd.n1891 vdd.n1890 9.3005
R19784 vdd.n1893 vdd.n1892 9.3005
R19785 vdd.n1876 vdd.n1875 9.3005
R19786 vdd.n1899 vdd.n1898 9.3005
R19787 vdd.n1901 vdd.n1900 9.3005
R19788 vdd.n1873 vdd.n1870 9.3005
R19789 vdd.n1908 vdd.n1907 9.3005
R19790 vdd.n1944 vdd.n1943 9.3005
R19791 vdd.n1939 vdd.n1938 9.3005
R19792 vdd.n1950 vdd.n1949 9.3005
R19793 vdd.n1952 vdd.n1951 9.3005
R19794 vdd.n1935 vdd.n1934 9.3005
R19795 vdd.n1958 vdd.n1957 9.3005
R19796 vdd.n1960 vdd.n1959 9.3005
R19797 vdd.n1932 vdd.n1929 9.3005
R19798 vdd.n1967 vdd.n1966 9.3005
R19799 vdd.n1823 vdd.t87 9.18308
R19800 vdd.n3423 vdd.t19 9.18308
R19801 vdd.n1517 vdd.t58 8.95635
R19802 vdd.n2265 vdd.t230 8.95635
R19803 vdd.n723 vdd.t226 8.95635
R19804 vdd.t35 vdd.n3477 8.95635
R19805 vdd.n312 vdd.n311 8.92171
R19806 vdd.n253 vdd.n252 8.92171
R19807 vdd.n210 vdd.n209 8.92171
R19808 vdd.n151 vdd.n150 8.92171
R19809 vdd.n109 vdd.n108 8.92171
R19810 vdd.n50 vdd.n49 8.92171
R19811 vdd.n2093 vdd.n2092 8.92171
R19812 vdd.n2152 vdd.n2151 8.92171
R19813 vdd.n1991 vdd.n1990 8.92171
R19814 vdd.n2050 vdd.n2049 8.92171
R19815 vdd.n1890 vdd.n1889 8.92171
R19816 vdd.n1949 vdd.n1948 8.92171
R19817 vdd.n231 vdd.n129 8.81535
R19818 vdd.n2071 vdd.n1969 8.81535
R19819 vdd.n1864 vdd.t118 8.72962
R19820 vdd.t39 vdd.n3486 8.72962
R19821 vdd.n2187 vdd.t44 8.50289
R19822 vdd.n3392 vdd.t41 8.50289
R19823 vdd.n28 vdd.n14 8.42249
R19824 vdd.n2213 vdd.t121 8.27616
R19825 vdd.t81 vdd.n656 8.27616
R19826 vdd.n3492 vdd.n3491 8.16225
R19827 vdd.n2175 vdd.n2174 8.16225
R19828 vdd.n308 vdd.n302 8.14595
R19829 vdd.n249 vdd.n243 8.14595
R19830 vdd.n206 vdd.n200 8.14595
R19831 vdd.n147 vdd.n141 8.14595
R19832 vdd.n105 vdd.n99 8.14595
R19833 vdd.n46 vdd.n40 8.14595
R19834 vdd.n2089 vdd.n2083 8.14595
R19835 vdd.n2148 vdd.n2142 8.14595
R19836 vdd.n1987 vdd.n1981 8.14595
R19837 vdd.n2046 vdd.n2040 8.14595
R19838 vdd.n1886 vdd.n1880 8.14595
R19839 vdd.n1945 vdd.n1939 8.14595
R19840 vdd.n1460 vdd.t25 8.04943
R19841 vdd.n3348 vdd.t139 8.04943
R19842 vdd.n2424 vdd.n1076 7.70933
R19843 vdd.n2424 vdd.n1079 7.70933
R19844 vdd.n2430 vdd.n1065 7.70933
R19845 vdd.n2436 vdd.n1065 7.70933
R19846 vdd.n2436 vdd.n1059 7.70933
R19847 vdd.n2442 vdd.n1059 7.70933
R19848 vdd.n2448 vdd.n1052 7.70933
R19849 vdd.n2448 vdd.n1055 7.70933
R19850 vdd.n2454 vdd.n1048 7.70933
R19851 vdd.n2461 vdd.n1034 7.70933
R19852 vdd.n2467 vdd.n1034 7.70933
R19853 vdd.n2473 vdd.n1028 7.70933
R19854 vdd.n2479 vdd.n1024 7.70933
R19855 vdd.n2485 vdd.n1018 7.70933
R19856 vdd.n2497 vdd.n1005 7.70933
R19857 vdd.n2503 vdd.n999 7.70933
R19858 vdd.n2503 vdd.n992 7.70933
R19859 vdd.n2511 vdd.n992 7.70933
R19860 vdd.n2593 vdd.n976 7.70933
R19861 vdd.n2945 vdd.n928 7.70933
R19862 vdd.n2957 vdd.n917 7.70933
R19863 vdd.n2957 vdd.n911 7.70933
R19864 vdd.n2963 vdd.n911 7.70933
R19865 vdd.n2969 vdd.n905 7.70933
R19866 vdd.n2975 vdd.n901 7.70933
R19867 vdd.n2981 vdd.n895 7.70933
R19868 vdd.n2993 vdd.n882 7.70933
R19869 vdd.n2999 vdd.n875 7.70933
R19870 vdd.n2999 vdd.n878 7.70933
R19871 vdd.n3006 vdd.n870 7.70933
R19872 vdd.n3012 vdd.n857 7.70933
R19873 vdd.n3018 vdd.n857 7.70933
R19874 vdd.n3024 vdd.n851 7.70933
R19875 vdd.n3024 vdd.n843 7.70933
R19876 vdd.n3075 vdd.n843 7.70933
R19877 vdd.n3075 vdd.n846 7.70933
R19878 vdd.n3081 vdd.n805 7.70933
R19879 vdd.n3151 vdd.n805 7.70933
R19880 vdd.n3004 vdd.n3003 7.49318
R19881 vdd.n2458 vdd.n2457 7.49318
R19882 vdd.n307 vdd.n304 7.3702
R19883 vdd.n248 vdd.n245 7.3702
R19884 vdd.n205 vdd.n202 7.3702
R19885 vdd.n146 vdd.n143 7.3702
R19886 vdd.n104 vdd.n101 7.3702
R19887 vdd.n45 vdd.n42 7.3702
R19888 vdd.n2088 vdd.n2085 7.3702
R19889 vdd.n2147 vdd.n2144 7.3702
R19890 vdd.n1986 vdd.n1983 7.3702
R19891 vdd.n2045 vdd.n2042 7.3702
R19892 vdd.n1885 vdd.n1882 7.3702
R19893 vdd.n1944 vdd.n1941 7.3702
R19894 vdd.n2442 vdd.t295 7.36923
R19895 vdd.t11 vdd.n851 7.36923
R19896 vdd.n2518 vdd.t206 7.25587
R19897 vdd.n2862 vdd.t194 7.25587
R19898 vdd.n2246 vdd.t65 7.1425
R19899 vdd.n679 vdd.t63 7.1425
R19900 vdd.n1720 vdd.n1719 6.98232
R19901 vdd.n2308 vdd.n2307 6.98232
R19902 vdd.n566 vdd.n565 6.98232
R19903 vdd.n3233 vdd.n3230 6.98232
R19904 vdd.t133 vdd.n1459 6.91577
R19905 vdd.n3356 vdd.t79 6.91577
R19906 vdd.n2205 vdd.t85 6.68904
R19907 vdd.n3372 vdd.t68 6.68904
R19908 vdd.t116 vdd.n1488 6.46231
R19909 vdd.n3400 vdd.t71 6.46231
R19910 vdd.n3492 vdd.n333 6.38151
R19911 vdd.n2174 vdd.n2173 6.38151
R19912 vdd.n1856 vdd.t56 6.23558
R19913 vdd.t130 vdd.n344 6.23558
R19914 vdd.t27 vdd.n1516 6.00885
R19915 vdd.n3471 vdd.t90 6.00885
R19916 vdd.t296 vdd.n1005 5.89549
R19917 vdd.n2969 vdd.t201 5.89549
R19918 vdd.n308 vdd.n307 5.81868
R19919 vdd.n249 vdd.n248 5.81868
R19920 vdd.n206 vdd.n205 5.81868
R19921 vdd.n147 vdd.n146 5.81868
R19922 vdd.n105 vdd.n104 5.81868
R19923 vdd.n46 vdd.n45 5.81868
R19924 vdd.n2089 vdd.n2088 5.81868
R19925 vdd.n2148 vdd.n2147 5.81868
R19926 vdd.n1987 vdd.n1986 5.81868
R19927 vdd.n2046 vdd.n2045 5.81868
R19928 vdd.n1886 vdd.n1885 5.81868
R19929 vdd.n1945 vdd.n1944 5.81868
R19930 vdd.n1815 vdd.t17 5.78212
R19931 vdd.n3462 vdd.t136 5.78212
R19932 vdd.n2601 vdd.n2600 5.77611
R19933 vdd.n1303 vdd.n1302 5.77611
R19934 vdd.n2874 vdd.n2873 5.77611
R19935 vdd.n3092 vdd.n3091 5.77611
R19936 vdd.n3156 vdd.n801 5.77611
R19937 vdd.n2768 vdd.n2706 5.77611
R19938 vdd.n2526 vdd.n983 5.77611
R19939 vdd.n1392 vdd.n1255 5.77611
R19940 vdd.n1682 vdd.n1681 5.62474
R19941 vdd.n2271 vdd.n2268 5.62474
R19942 vdd.n3443 vdd.n428 5.62474
R19943 vdd.n3317 vdd.n690 5.62474
R19944 vdd.n1539 vdd.t17 5.55539
R19945 vdd.t191 vdd.n1028 5.55539
R19946 vdd.n2473 vdd.t10 5.55539
R19947 vdd.t205 vdd.n882 5.55539
R19948 vdd.n2993 vdd.t1 5.55539
R19949 vdd.t136 vdd.n3461 5.55539
R19950 vdd.n1048 vdd.t275 5.44203
R19951 vdd.n3006 vdd.t244 5.44203
R19952 vdd.n1831 vdd.t27 5.32866
R19953 vdd.n2430 vdd.t222 5.32866
R19954 vdd.n1338 vdd.t264 5.32866
R19955 vdd.n2951 vdd.t268 5.32866
R19956 vdd.n846 vdd.t218 5.32866
R19957 vdd.t90 vdd.n3470 5.32866
R19958 vdd.n1847 vdd.t56 5.10193
R19959 vdd.n3479 vdd.t130 5.10193
R19960 vdd.n311 vdd.n302 5.04292
R19961 vdd.n252 vdd.n243 5.04292
R19962 vdd.n209 vdd.n200 5.04292
R19963 vdd.n150 vdd.n141 5.04292
R19964 vdd.n108 vdd.n99 5.04292
R19965 vdd.n49 vdd.n40 5.04292
R19966 vdd.n2092 vdd.n2083 5.04292
R19967 vdd.n2151 vdd.n2142 5.04292
R19968 vdd.n1990 vdd.n1981 5.04292
R19969 vdd.n2049 vdd.n2040 5.04292
R19970 vdd.n1889 vdd.n1880 5.04292
R19971 vdd.n1948 vdd.n1939 5.04292
R19972 vdd.n2479 vdd.t203 4.98857
R19973 vdd.n895 vdd.t189 4.98857
R19974 vdd.n2179 vdd.t116 4.8752
R19975 vdd.t13 vdd.t213 4.8752
R19976 vdd.t12 vdd.t15 4.8752
R19977 vdd.t211 vdd.t216 4.8752
R19978 vdd.t187 vdd.t198 4.8752
R19979 vdd.t71 vdd.n340 4.8752
R19980 vdd.n2602 vdd.n2601 4.83952
R19981 vdd.n1302 vdd.n1301 4.83952
R19982 vdd.n2875 vdd.n2874 4.83952
R19983 vdd.n3093 vdd.n3092 4.83952
R19984 vdd.n801 vdd.n796 4.83952
R19985 vdd.n2765 vdd.n2706 4.83952
R19986 vdd.n2529 vdd.n983 4.83952
R19987 vdd.n1395 vdd.n1255 4.83952
R19988 vdd.n2276 vdd.n2275 4.74817
R19989 vdd.n1428 vdd.n1423 4.74817
R19990 vdd.n1125 vdd.n1122 4.74817
R19991 vdd.n2369 vdd.n1121 4.74817
R19992 vdd.n2374 vdd.n1122 4.74817
R19993 vdd.n2373 vdd.n1121 4.74817
R19994 vdd.n3310 vdd.n3309 4.74817
R19995 vdd.n3307 vdd.n3306 4.74817
R19996 vdd.n3307 vdd.n732 4.74817
R19997 vdd.n3309 vdd.n729 4.74817
R19998 vdd.n3192 vdd.n784 4.74817
R19999 vdd.n3188 vdd.n3186 4.74817
R20000 vdd.n3191 vdd.n3186 4.74817
R20001 vdd.n3195 vdd.n784 4.74817
R20002 vdd.n2275 vdd.n1221 4.74817
R20003 vdd.n1425 vdd.n1423 4.74817
R20004 vdd.n333 vdd.n332 4.7074
R20005 vdd.n231 vdd.n230 4.7074
R20006 vdd.n2173 vdd.n2172 4.7074
R20007 vdd.n2071 vdd.n2070 4.7074
R20008 vdd.n1482 vdd.t85 4.64847
R20009 vdd.n2454 vdd.t180 4.64847
R20010 vdd.n1018 vdd.t0 4.64847
R20011 vdd.n2975 vdd.t14 4.64847
R20012 vdd.n870 vdd.t208 4.64847
R20013 vdd.n3381 vdd.t68 4.64847
R20014 vdd.n2221 vdd.t133 4.42174
R20015 vdd.t79 vdd.n655 4.42174
R20016 vdd.n312 vdd.n300 4.26717
R20017 vdd.n253 vdd.n241 4.26717
R20018 vdd.n210 vdd.n198 4.26717
R20019 vdd.n151 vdd.n139 4.26717
R20020 vdd.n109 vdd.n97 4.26717
R20021 vdd.n50 vdd.n38 4.26717
R20022 vdd.n2093 vdd.n2081 4.26717
R20023 vdd.n2152 vdd.n2140 4.26717
R20024 vdd.n1991 vdd.n1979 4.26717
R20025 vdd.n2050 vdd.n2038 4.26717
R20026 vdd.n1890 vdd.n1878 4.26717
R20027 vdd.n1949 vdd.n1937 4.26717
R20028 vdd.n2237 vdd.t65 4.19501
R20029 vdd.n3340 vdd.t63 4.19501
R20030 vdd.n333 vdd.n231 4.10845
R20031 vdd.n2173 vdd.n2071 4.10845
R20032 vdd.n289 vdd.t101 4.06363
R20033 vdd.n289 vdd.t149 4.06363
R20034 vdd.n287 vdd.t152 4.06363
R20035 vdd.n287 vdd.t20 4.06363
R20036 vdd.n285 vdd.t55 4.06363
R20037 vdd.n285 vdd.t125 4.06363
R20038 vdd.n283 vdd.t156 4.06363
R20039 vdd.n283 vdd.t167 4.06363
R20040 vdd.n281 vdd.t172 4.06363
R20041 vdd.n281 vdd.t62 4.06363
R20042 vdd.n279 vdd.t95 4.06363
R20043 vdd.n279 vdd.t171 4.06363
R20044 vdd.n277 vdd.t173 4.06363
R20045 vdd.n277 vdd.t94 4.06363
R20046 vdd.n275 vdd.t100 4.06363
R20047 vdd.n275 vdd.t103 4.06363
R20048 vdd.n273 vdd.t151 4.06363
R20049 vdd.n273 vdd.t46 4.06363
R20050 vdd.n187 vdd.t78 4.06363
R20051 vdd.n187 vdd.t137 4.06363
R20052 vdd.n185 vdd.t138 4.06363
R20053 vdd.n185 vdd.t169 4.06363
R20054 vdd.n183 vdd.t36 4.06363
R20055 vdd.n183 vdd.t106 4.06363
R20056 vdd.n181 vdd.t143 4.06363
R20057 vdd.n181 vdd.t157 4.06363
R20058 vdd.n179 vdd.t161 4.06363
R20059 vdd.n179 vdd.t40 4.06363
R20060 vdd.n177 vdd.t70 4.06363
R20061 vdd.n177 vdd.t160 4.06363
R20062 vdd.n175 vdd.t162 4.06363
R20063 vdd.n175 vdd.t69 4.06363
R20064 vdd.n173 vdd.t80 4.06363
R20065 vdd.n173 vdd.t82 4.06363
R20066 vdd.n171 vdd.t140 4.06363
R20067 vdd.n171 vdd.t22 4.06363
R20068 vdd.n86 vdd.t115 4.06363
R20069 vdd.n86 vdd.t141 4.06363
R20070 vdd.n84 vdd.t91 4.06363
R20071 vdd.n84 vdd.t163 4.06363
R20072 vdd.n82 vdd.t54 4.06363
R20073 vdd.n82 vdd.t150 4.06363
R20074 vdd.n80 vdd.t48 4.06363
R20075 vdd.n80 vdd.t131 4.06363
R20076 vdd.n78 vdd.t72 4.06363
R20077 vdd.n78 vdd.t158 4.06363
R20078 vdd.n76 vdd.t42 4.06363
R20079 vdd.n76 vdd.t109 4.06363
R20080 vdd.n74 vdd.t30 4.06363
R20081 vdd.n74 vdd.t83 4.06363
R20082 vdd.n72 vdd.t168 4.06363
R20083 vdd.n72 vdd.t147 4.06363
R20084 vdd.n70 vdd.t154 4.06363
R20085 vdd.n70 vdd.t96 4.06363
R20086 vdd.n2113 vdd.t120 4.06363
R20087 vdd.n2113 vdd.t52 4.06363
R20088 vdd.n2115 vdd.t176 4.06363
R20089 vdd.n2115 vdd.t146 4.06363
R20090 vdd.n2117 vdd.t144 4.06363
R20091 vdd.n2117 vdd.t93 4.06363
R20092 vdd.n2119 vdd.t89 4.06363
R20093 vdd.n2119 vdd.t145 4.06363
R20094 vdd.n2121 vdd.t128 4.06363
R20095 vdd.n2121 vdd.t127 4.06363
R20096 vdd.n2123 vdd.t84 4.06363
R20097 vdd.n2123 vdd.t53 4.06363
R20098 vdd.n2125 vdd.t51 4.06363
R20099 vdd.n2125 vdd.t126 4.06363
R20100 vdd.n2127 vdd.t104 4.06363
R20101 vdd.n2127 vdd.t49 4.06363
R20102 vdd.n2129 vdd.t43 4.06363
R20103 vdd.n2129 vdd.t148 4.06363
R20104 vdd.n2011 vdd.t102 4.06363
R20105 vdd.n2011 vdd.t26 4.06363
R20106 vdd.n2013 vdd.t166 4.06363
R20107 vdd.n2013 vdd.t134 4.06363
R20108 vdd.n2015 vdd.t129 4.06363
R20109 vdd.n2015 vdd.t67 4.06363
R20110 vdd.n2017 vdd.t61 4.06363
R20111 vdd.n2017 vdd.t110 4.06363
R20112 vdd.n2019 vdd.t119 4.06363
R20113 vdd.n2019 vdd.t117 4.06363
R20114 vdd.n2021 vdd.t57 4.06363
R20115 vdd.n2021 vdd.t32 4.06363
R20116 vdd.n2023 vdd.t24 4.06363
R20117 vdd.n2023 vdd.t114 4.06363
R20118 vdd.n2025 vdd.t88 4.06363
R20119 vdd.n2025 vdd.t28 4.06363
R20120 vdd.n2027 vdd.t18 4.06363
R20121 vdd.n2027 vdd.t135 4.06363
R20122 vdd.n1910 vdd.t98 4.06363
R20123 vdd.n1910 vdd.t155 4.06363
R20124 vdd.n1912 vdd.t122 4.06363
R20125 vdd.n1912 vdd.t170 4.06363
R20126 vdd.n1914 vdd.t86 4.06363
R20127 vdd.n1914 vdd.t34 4.06363
R20128 vdd.n1916 vdd.t113 4.06363
R20129 vdd.n1916 vdd.t45 4.06363
R20130 vdd.n1918 vdd.t159 4.06363
R20131 vdd.n1918 vdd.t175 4.06363
R20132 vdd.n1920 vdd.t132 4.06363
R20133 vdd.n1920 vdd.t50 4.06363
R20134 vdd.n1922 vdd.t123 4.06363
R20135 vdd.n1922 vdd.t59 4.06363
R20136 vdd.n1924 vdd.t164 4.06363
R20137 vdd.n1924 vdd.t92 4.06363
R20138 vdd.n1926 vdd.t142 4.06363
R20139 vdd.n1926 vdd.t112 4.06363
R20140 vdd.n26 vdd.t6 3.9605
R20141 vdd.n26 vdd.t177 3.9605
R20142 vdd.n23 vdd.t183 3.9605
R20143 vdd.n23 vdd.t182 3.9605
R20144 vdd.n21 vdd.t193 3.9605
R20145 vdd.n21 vdd.t186 3.9605
R20146 vdd.n20 vdd.t7 3.9605
R20147 vdd.n20 vdd.t9 3.9605
R20148 vdd.n15 vdd.t192 3.9605
R20149 vdd.n15 vdd.t8 3.9605
R20150 vdd.n16 vdd.t178 3.9605
R20151 vdd.n16 vdd.t4 3.9605
R20152 vdd.n18 vdd.t181 3.9605
R20153 vdd.n18 vdd.t184 3.9605
R20154 vdd.n25 vdd.t5 3.9605
R20155 vdd.n25 vdd.t185 3.9605
R20156 vdd.n2511 vdd.t2 3.85492
R20157 vdd.n1338 vdd.t2 3.85492
R20158 vdd.n2951 vdd.t298 3.85492
R20159 vdd.t298 vdd.n917 3.85492
R20160 vdd.n7 vdd.t188 3.61217
R20161 vdd.n7 vdd.t190 3.61217
R20162 vdd.n8 vdd.t212 3.61217
R20163 vdd.n8 vdd.t202 3.61217
R20164 vdd.n10 vdd.t195 3.61217
R20165 vdd.n10 vdd.t299 3.61217
R20166 vdd.n12 vdd.t294 3.61217
R20167 vdd.n12 vdd.t197 3.61217
R20168 vdd.n5 vdd.t200 3.61217
R20169 vdd.n5 vdd.t210 3.61217
R20170 vdd.n3 vdd.t3 3.61217
R20171 vdd.n3 vdd.t207 3.61217
R20172 vdd.n1 vdd.t297 3.61217
R20173 vdd.n1 vdd.t16 3.61217
R20174 vdd.n0 vdd.t204 3.61217
R20175 vdd.n0 vdd.t214 3.61217
R20176 vdd.n316 vdd.n315 3.49141
R20177 vdd.n257 vdd.n256 3.49141
R20178 vdd.n214 vdd.n213 3.49141
R20179 vdd.n155 vdd.n154 3.49141
R20180 vdd.n113 vdd.n112 3.49141
R20181 vdd.n54 vdd.n53 3.49141
R20182 vdd.n2097 vdd.n2096 3.49141
R20183 vdd.n2156 vdd.n2155 3.49141
R20184 vdd.n1995 vdd.n1994 3.49141
R20185 vdd.n2054 vdd.n2053 3.49141
R20186 vdd.n1894 vdd.n1893 3.49141
R20187 vdd.n1953 vdd.n1952 3.49141
R20188 vdd.n2665 vdd.t199 3.40145
R20189 vdd.n2938 vdd.t196 3.40145
R20190 vdd.n2238 vdd.t25 3.28809
R20191 vdd.n3339 vdd.t139 3.28809
R20192 vdd.n3003 vdd.n3002 3.12245
R20193 vdd.n2459 vdd.n2458 3.12245
R20194 vdd.t121 vdd.n1466 3.06136
R20195 vdd.n1055 vdd.t180 3.06136
R20196 vdd.n2491 vdd.t0 3.06136
R20197 vdd.n2847 vdd.t14 3.06136
R20198 vdd.n3012 vdd.t208 3.06136
R20199 vdd.n3364 vdd.t81 3.06136
R20200 vdd.n2196 vdd.t44 2.83463
R20201 vdd.n644 vdd.t41 2.83463
R20202 vdd.n1359 vdd.t203 2.72126
R20203 vdd.n2987 vdd.t189 2.72126
R20204 vdd.n319 vdd.n298 2.71565
R20205 vdd.n260 vdd.n239 2.71565
R20206 vdd.n217 vdd.n196 2.71565
R20207 vdd.n158 vdd.n137 2.71565
R20208 vdd.n116 vdd.n95 2.71565
R20209 vdd.n57 vdd.n36 2.71565
R20210 vdd.n2100 vdd.n2079 2.71565
R20211 vdd.n2159 vdd.n2138 2.71565
R20212 vdd.n1998 vdd.n1977 2.71565
R20213 vdd.n2057 vdd.n2036 2.71565
R20214 vdd.n1897 vdd.n1876 2.71565
R20215 vdd.n1956 vdd.n1935 2.71565
R20216 vdd.t118 vdd.n1494 2.6079
R20217 vdd.n3487 vdd.t39 2.6079
R20218 vdd.t15 vdd.n999 2.49453
R20219 vdd.n2963 vdd.t211 2.49453
R20220 vdd.n306 vdd.n305 2.4129
R20221 vdd.n247 vdd.n246 2.4129
R20222 vdd.n204 vdd.n203 2.4129
R20223 vdd.n145 vdd.n144 2.4129
R20224 vdd.n103 vdd.n102 2.4129
R20225 vdd.n44 vdd.n43 2.4129
R20226 vdd.n2087 vdd.n2086 2.4129
R20227 vdd.n2146 vdd.n2145 2.4129
R20228 vdd.n1985 vdd.n1984 2.4129
R20229 vdd.n2044 vdd.n2043 2.4129
R20230 vdd.n1884 vdd.n1883 2.4129
R20231 vdd.n1943 vdd.n1942 2.4129
R20232 vdd.n1848 vdd.t58 2.38117
R20233 vdd.n2256 vdd.t230 2.38117
R20234 vdd.n1079 vdd.t222 2.38117
R20235 vdd.n2518 vdd.t264 2.38117
R20236 vdd.n2862 vdd.t268 2.38117
R20237 vdd.n3081 vdd.t218 2.38117
R20238 vdd.n3323 vdd.t226 2.38117
R20239 vdd.n3478 vdd.t35 2.38117
R20240 vdd.n2381 vdd.n1122 2.27742
R20241 vdd.n2381 vdd.n1121 2.27742
R20242 vdd.n3308 vdd.n3307 2.27742
R20243 vdd.n3309 vdd.n3308 2.27742
R20244 vdd.n3186 vdd.n3185 2.27742
R20245 vdd.n3185 vdd.n784 2.27742
R20246 vdd.n2275 vdd.n2274 2.27742
R20247 vdd.n2274 vdd.n1423 2.27742
R20248 vdd.t87 vdd.n1523 2.15444
R20249 vdd.n2467 vdd.t191 2.15444
R20250 vdd.n1359 vdd.t10 2.15444
R20251 vdd.n2987 vdd.t205 2.15444
R20252 vdd.t1 vdd.n875 2.15444
R20253 vdd.n3469 vdd.t19 2.15444
R20254 vdd.n320 vdd.n296 1.93989
R20255 vdd.n261 vdd.n237 1.93989
R20256 vdd.n218 vdd.n194 1.93989
R20257 vdd.n159 vdd.n135 1.93989
R20258 vdd.n117 vdd.n93 1.93989
R20259 vdd.n58 vdd.n34 1.93989
R20260 vdd.n2101 vdd.n2077 1.93989
R20261 vdd.n2160 vdd.n2136 1.93989
R20262 vdd.n1999 vdd.n1975 1.93989
R20263 vdd.n2058 vdd.n2034 1.93989
R20264 vdd.n1898 vdd.n1874 1.93989
R20265 vdd.n1957 vdd.n1933 1.93989
R20266 vdd.n1806 vdd.t73 1.92771
R20267 vdd.t37 vdd.n375 1.92771
R20268 vdd.n2491 vdd.t296 1.81434
R20269 vdd.n2847 vdd.t201 1.81434
R20270 vdd.n1814 vdd.t111 1.70098
R20271 vdd.n3463 vdd.t77 1.70098
R20272 vdd.n2485 vdd.t213 1.58761
R20273 vdd.n901 vdd.t187 1.58761
R20274 vdd.n1839 vdd.t23 1.47425
R20275 vdd.n361 vdd.t105 1.47425
R20276 vdd.n1505 vdd.t31 1.24752
R20277 vdd.n2461 vdd.t179 1.24752
R20278 vdd.n1024 vdd.t13 1.24752
R20279 vdd.n2981 vdd.t198 1.24752
R20280 vdd.n878 vdd.t215 1.24752
R20281 vdd.t47 vdd.n3485 1.24752
R20282 vdd.n331 vdd.n291 1.16414
R20283 vdd.n324 vdd.n323 1.16414
R20284 vdd.n272 vdd.n232 1.16414
R20285 vdd.n265 vdd.n264 1.16414
R20286 vdd.n229 vdd.n189 1.16414
R20287 vdd.n222 vdd.n221 1.16414
R20288 vdd.n170 vdd.n130 1.16414
R20289 vdd.n163 vdd.n162 1.16414
R20290 vdd.n128 vdd.n88 1.16414
R20291 vdd.n121 vdd.n120 1.16414
R20292 vdd.n69 vdd.n29 1.16414
R20293 vdd.n62 vdd.n61 1.16414
R20294 vdd.n2112 vdd.n2072 1.16414
R20295 vdd.n2105 vdd.n2104 1.16414
R20296 vdd.n2171 vdd.n2131 1.16414
R20297 vdd.n2164 vdd.n2163 1.16414
R20298 vdd.n2010 vdd.n1970 1.16414
R20299 vdd.n2003 vdd.n2002 1.16414
R20300 vdd.n2069 vdd.n2029 1.16414
R20301 vdd.n2062 vdd.n2061 1.16414
R20302 vdd.n1909 vdd.n1869 1.16414
R20303 vdd.n1902 vdd.n1901 1.16414
R20304 vdd.n1968 vdd.n1928 1.16414
R20305 vdd.n1961 vdd.n1960 1.16414
R20306 vdd.n2188 vdd.t60 1.02079
R20307 vdd.t275 vdd.t179 1.02079
R20308 vdd.t215 vdd.t244 1.02079
R20309 vdd.t108 vdd.n633 1.02079
R20310 vdd.n2174 vdd.n28 1.00834
R20311 vdd vdd.n3492 1.0005
R20312 vdd.n1685 vdd.n1681 0.970197
R20313 vdd.n2272 vdd.n2271 0.970197
R20314 vdd.n618 vdd.n428 0.970197
R20315 vdd.n3187 vdd.n690 0.970197
R20316 vdd.n2204 vdd.t33 0.794056
R20317 vdd.n3373 vdd.t29 0.794056
R20318 vdd.n2229 vdd.t97 0.567326
R20319 vdd.t21 vdd.n662 0.567326
R20320 vdd.n2262 vdd.n1123 0.530988
R20321 vdd.n726 vdd.n682 0.530988
R20322 vdd.n464 vdd.n391 0.530988
R20323 vdd.n3442 vdd.n3441 0.530988
R20324 vdd.n3319 vdd.n3318 0.530988
R20325 vdd.n2251 vdd.n1424 0.530988
R20326 vdd.n1683 vdd.n1548 0.530988
R20327 vdd.n1785 vdd.n1784 0.530988
R20328 vdd.n4 vdd.n2 0.459552
R20329 vdd.n11 vdd.n9 0.459552
R20330 vdd.t206 vdd.n976 0.453961
R20331 vdd.n2945 vdd.t194 0.453961
R20332 vdd.n329 vdd.n328 0.388379
R20333 vdd.n295 vdd.n293 0.388379
R20334 vdd.n270 vdd.n269 0.388379
R20335 vdd.n236 vdd.n234 0.388379
R20336 vdd.n227 vdd.n226 0.388379
R20337 vdd.n193 vdd.n191 0.388379
R20338 vdd.n168 vdd.n167 0.388379
R20339 vdd.n134 vdd.n132 0.388379
R20340 vdd.n126 vdd.n125 0.388379
R20341 vdd.n92 vdd.n90 0.388379
R20342 vdd.n67 vdd.n66 0.388379
R20343 vdd.n33 vdd.n31 0.388379
R20344 vdd.n2110 vdd.n2109 0.388379
R20345 vdd.n2076 vdd.n2074 0.388379
R20346 vdd.n2169 vdd.n2168 0.388379
R20347 vdd.n2135 vdd.n2133 0.388379
R20348 vdd.n2008 vdd.n2007 0.388379
R20349 vdd.n1974 vdd.n1972 0.388379
R20350 vdd.n2067 vdd.n2066 0.388379
R20351 vdd.n2033 vdd.n2031 0.388379
R20352 vdd.n1907 vdd.n1906 0.388379
R20353 vdd.n1873 vdd.n1871 0.388379
R20354 vdd.n1966 vdd.n1965 0.388379
R20355 vdd.n1932 vdd.n1930 0.388379
R20356 vdd.n19 vdd.n17 0.387128
R20357 vdd.n24 vdd.n22 0.387128
R20358 vdd.n6 vdd.n4 0.358259
R20359 vdd.n13 vdd.n11 0.358259
R20360 vdd.n276 vdd.n274 0.358259
R20361 vdd.n278 vdd.n276 0.358259
R20362 vdd.n280 vdd.n278 0.358259
R20363 vdd.n282 vdd.n280 0.358259
R20364 vdd.n284 vdd.n282 0.358259
R20365 vdd.n286 vdd.n284 0.358259
R20366 vdd.n288 vdd.n286 0.358259
R20367 vdd.n290 vdd.n288 0.358259
R20368 vdd.n332 vdd.n290 0.358259
R20369 vdd.n174 vdd.n172 0.358259
R20370 vdd.n176 vdd.n174 0.358259
R20371 vdd.n178 vdd.n176 0.358259
R20372 vdd.n180 vdd.n178 0.358259
R20373 vdd.n182 vdd.n180 0.358259
R20374 vdd.n184 vdd.n182 0.358259
R20375 vdd.n186 vdd.n184 0.358259
R20376 vdd.n188 vdd.n186 0.358259
R20377 vdd.n230 vdd.n188 0.358259
R20378 vdd.n73 vdd.n71 0.358259
R20379 vdd.n75 vdd.n73 0.358259
R20380 vdd.n77 vdd.n75 0.358259
R20381 vdd.n79 vdd.n77 0.358259
R20382 vdd.n81 vdd.n79 0.358259
R20383 vdd.n83 vdd.n81 0.358259
R20384 vdd.n85 vdd.n83 0.358259
R20385 vdd.n87 vdd.n85 0.358259
R20386 vdd.n129 vdd.n87 0.358259
R20387 vdd.n2172 vdd.n2130 0.358259
R20388 vdd.n2130 vdd.n2128 0.358259
R20389 vdd.n2128 vdd.n2126 0.358259
R20390 vdd.n2126 vdd.n2124 0.358259
R20391 vdd.n2124 vdd.n2122 0.358259
R20392 vdd.n2122 vdd.n2120 0.358259
R20393 vdd.n2120 vdd.n2118 0.358259
R20394 vdd.n2118 vdd.n2116 0.358259
R20395 vdd.n2116 vdd.n2114 0.358259
R20396 vdd.n2070 vdd.n2028 0.358259
R20397 vdd.n2028 vdd.n2026 0.358259
R20398 vdd.n2026 vdd.n2024 0.358259
R20399 vdd.n2024 vdd.n2022 0.358259
R20400 vdd.n2022 vdd.n2020 0.358259
R20401 vdd.n2020 vdd.n2018 0.358259
R20402 vdd.n2018 vdd.n2016 0.358259
R20403 vdd.n2016 vdd.n2014 0.358259
R20404 vdd.n2014 vdd.n2012 0.358259
R20405 vdd.n1969 vdd.n1927 0.358259
R20406 vdd.n1927 vdd.n1925 0.358259
R20407 vdd.n1925 vdd.n1923 0.358259
R20408 vdd.n1923 vdd.n1921 0.358259
R20409 vdd.n1921 vdd.n1919 0.358259
R20410 vdd.n1919 vdd.n1917 0.358259
R20411 vdd.n1917 vdd.n1915 0.358259
R20412 vdd.n1915 vdd.n1913 0.358259
R20413 vdd.n1913 vdd.n1911 0.358259
R20414 vdd.t295 vdd.n1052 0.340595
R20415 vdd.n2497 vdd.t12 0.340595
R20416 vdd.t216 vdd.n905 0.340595
R20417 vdd.n3018 vdd.t11 0.340595
R20418 vdd.n14 vdd.n6 0.334552
R20419 vdd.n14 vdd.n13 0.334552
R20420 vdd.n27 vdd.n19 0.21707
R20421 vdd.n27 vdd.n24 0.21707
R20422 vdd.n330 vdd.n292 0.155672
R20423 vdd.n322 vdd.n292 0.155672
R20424 vdd.n322 vdd.n321 0.155672
R20425 vdd.n321 vdd.n297 0.155672
R20426 vdd.n314 vdd.n297 0.155672
R20427 vdd.n314 vdd.n313 0.155672
R20428 vdd.n313 vdd.n301 0.155672
R20429 vdd.n306 vdd.n301 0.155672
R20430 vdd.n271 vdd.n233 0.155672
R20431 vdd.n263 vdd.n233 0.155672
R20432 vdd.n263 vdd.n262 0.155672
R20433 vdd.n262 vdd.n238 0.155672
R20434 vdd.n255 vdd.n238 0.155672
R20435 vdd.n255 vdd.n254 0.155672
R20436 vdd.n254 vdd.n242 0.155672
R20437 vdd.n247 vdd.n242 0.155672
R20438 vdd.n228 vdd.n190 0.155672
R20439 vdd.n220 vdd.n190 0.155672
R20440 vdd.n220 vdd.n219 0.155672
R20441 vdd.n219 vdd.n195 0.155672
R20442 vdd.n212 vdd.n195 0.155672
R20443 vdd.n212 vdd.n211 0.155672
R20444 vdd.n211 vdd.n199 0.155672
R20445 vdd.n204 vdd.n199 0.155672
R20446 vdd.n169 vdd.n131 0.155672
R20447 vdd.n161 vdd.n131 0.155672
R20448 vdd.n161 vdd.n160 0.155672
R20449 vdd.n160 vdd.n136 0.155672
R20450 vdd.n153 vdd.n136 0.155672
R20451 vdd.n153 vdd.n152 0.155672
R20452 vdd.n152 vdd.n140 0.155672
R20453 vdd.n145 vdd.n140 0.155672
R20454 vdd.n127 vdd.n89 0.155672
R20455 vdd.n119 vdd.n89 0.155672
R20456 vdd.n119 vdd.n118 0.155672
R20457 vdd.n118 vdd.n94 0.155672
R20458 vdd.n111 vdd.n94 0.155672
R20459 vdd.n111 vdd.n110 0.155672
R20460 vdd.n110 vdd.n98 0.155672
R20461 vdd.n103 vdd.n98 0.155672
R20462 vdd.n68 vdd.n30 0.155672
R20463 vdd.n60 vdd.n30 0.155672
R20464 vdd.n60 vdd.n59 0.155672
R20465 vdd.n59 vdd.n35 0.155672
R20466 vdd.n52 vdd.n35 0.155672
R20467 vdd.n52 vdd.n51 0.155672
R20468 vdd.n51 vdd.n39 0.155672
R20469 vdd.n44 vdd.n39 0.155672
R20470 vdd.n2111 vdd.n2073 0.155672
R20471 vdd.n2103 vdd.n2073 0.155672
R20472 vdd.n2103 vdd.n2102 0.155672
R20473 vdd.n2102 vdd.n2078 0.155672
R20474 vdd.n2095 vdd.n2078 0.155672
R20475 vdd.n2095 vdd.n2094 0.155672
R20476 vdd.n2094 vdd.n2082 0.155672
R20477 vdd.n2087 vdd.n2082 0.155672
R20478 vdd.n2170 vdd.n2132 0.155672
R20479 vdd.n2162 vdd.n2132 0.155672
R20480 vdd.n2162 vdd.n2161 0.155672
R20481 vdd.n2161 vdd.n2137 0.155672
R20482 vdd.n2154 vdd.n2137 0.155672
R20483 vdd.n2154 vdd.n2153 0.155672
R20484 vdd.n2153 vdd.n2141 0.155672
R20485 vdd.n2146 vdd.n2141 0.155672
R20486 vdd.n2009 vdd.n1971 0.155672
R20487 vdd.n2001 vdd.n1971 0.155672
R20488 vdd.n2001 vdd.n2000 0.155672
R20489 vdd.n2000 vdd.n1976 0.155672
R20490 vdd.n1993 vdd.n1976 0.155672
R20491 vdd.n1993 vdd.n1992 0.155672
R20492 vdd.n1992 vdd.n1980 0.155672
R20493 vdd.n1985 vdd.n1980 0.155672
R20494 vdd.n2068 vdd.n2030 0.155672
R20495 vdd.n2060 vdd.n2030 0.155672
R20496 vdd.n2060 vdd.n2059 0.155672
R20497 vdd.n2059 vdd.n2035 0.155672
R20498 vdd.n2052 vdd.n2035 0.155672
R20499 vdd.n2052 vdd.n2051 0.155672
R20500 vdd.n2051 vdd.n2039 0.155672
R20501 vdd.n2044 vdd.n2039 0.155672
R20502 vdd.n1908 vdd.n1870 0.155672
R20503 vdd.n1900 vdd.n1870 0.155672
R20504 vdd.n1900 vdd.n1899 0.155672
R20505 vdd.n1899 vdd.n1875 0.155672
R20506 vdd.n1892 vdd.n1875 0.155672
R20507 vdd.n1892 vdd.n1891 0.155672
R20508 vdd.n1891 vdd.n1879 0.155672
R20509 vdd.n1884 vdd.n1879 0.155672
R20510 vdd.n1967 vdd.n1929 0.155672
R20511 vdd.n1959 vdd.n1929 0.155672
R20512 vdd.n1959 vdd.n1958 0.155672
R20513 vdd.n1958 vdd.n1934 0.155672
R20514 vdd.n1951 vdd.n1934 0.155672
R20515 vdd.n1951 vdd.n1950 0.155672
R20516 vdd.n1950 vdd.n1938 0.155672
R20517 vdd.n1943 vdd.n1938 0.155672
R20518 vdd.n1128 vdd.n1120 0.152939
R20519 vdd.n1132 vdd.n1128 0.152939
R20520 vdd.n1133 vdd.n1132 0.152939
R20521 vdd.n1134 vdd.n1133 0.152939
R20522 vdd.n1135 vdd.n1134 0.152939
R20523 vdd.n1139 vdd.n1135 0.152939
R20524 vdd.n1140 vdd.n1139 0.152939
R20525 vdd.n1141 vdd.n1140 0.152939
R20526 vdd.n1142 vdd.n1141 0.152939
R20527 vdd.n1146 vdd.n1142 0.152939
R20528 vdd.n1147 vdd.n1146 0.152939
R20529 vdd.n1148 vdd.n1147 0.152939
R20530 vdd.n2345 vdd.n1148 0.152939
R20531 vdd.n2345 vdd.n2344 0.152939
R20532 vdd.n2344 vdd.n2343 0.152939
R20533 vdd.n2343 vdd.n1154 0.152939
R20534 vdd.n1159 vdd.n1154 0.152939
R20535 vdd.n1160 vdd.n1159 0.152939
R20536 vdd.n1161 vdd.n1160 0.152939
R20537 vdd.n1165 vdd.n1161 0.152939
R20538 vdd.n1166 vdd.n1165 0.152939
R20539 vdd.n1167 vdd.n1166 0.152939
R20540 vdd.n1168 vdd.n1167 0.152939
R20541 vdd.n1172 vdd.n1168 0.152939
R20542 vdd.n1173 vdd.n1172 0.152939
R20543 vdd.n1174 vdd.n1173 0.152939
R20544 vdd.n1175 vdd.n1174 0.152939
R20545 vdd.n1179 vdd.n1175 0.152939
R20546 vdd.n1180 vdd.n1179 0.152939
R20547 vdd.n1181 vdd.n1180 0.152939
R20548 vdd.n1182 vdd.n1181 0.152939
R20549 vdd.n1186 vdd.n1182 0.152939
R20550 vdd.n1187 vdd.n1186 0.152939
R20551 vdd.n1188 vdd.n1187 0.152939
R20552 vdd.n2306 vdd.n1188 0.152939
R20553 vdd.n2306 vdd.n2305 0.152939
R20554 vdd.n2305 vdd.n2304 0.152939
R20555 vdd.n2304 vdd.n1194 0.152939
R20556 vdd.n1199 vdd.n1194 0.152939
R20557 vdd.n1200 vdd.n1199 0.152939
R20558 vdd.n1201 vdd.n1200 0.152939
R20559 vdd.n1205 vdd.n1201 0.152939
R20560 vdd.n1206 vdd.n1205 0.152939
R20561 vdd.n1207 vdd.n1206 0.152939
R20562 vdd.n1208 vdd.n1207 0.152939
R20563 vdd.n1212 vdd.n1208 0.152939
R20564 vdd.n1213 vdd.n1212 0.152939
R20565 vdd.n1214 vdd.n1213 0.152939
R20566 vdd.n1215 vdd.n1214 0.152939
R20567 vdd.n1219 vdd.n1215 0.152939
R20568 vdd.n1220 vdd.n1219 0.152939
R20569 vdd.n2380 vdd.n1123 0.152939
R20570 vdd.n2176 vdd.n1485 0.152939
R20571 vdd.n2191 vdd.n1485 0.152939
R20572 vdd.n2192 vdd.n2191 0.152939
R20573 vdd.n2193 vdd.n2192 0.152939
R20574 vdd.n2193 vdd.n1474 0.152939
R20575 vdd.n2208 vdd.n1474 0.152939
R20576 vdd.n2209 vdd.n2208 0.152939
R20577 vdd.n2210 vdd.n2209 0.152939
R20578 vdd.n2210 vdd.n1463 0.152939
R20579 vdd.n2224 vdd.n1463 0.152939
R20580 vdd.n2225 vdd.n2224 0.152939
R20581 vdd.n2226 vdd.n2225 0.152939
R20582 vdd.n2226 vdd.n1451 0.152939
R20583 vdd.n2241 vdd.n1451 0.152939
R20584 vdd.n2242 vdd.n2241 0.152939
R20585 vdd.n2243 vdd.n2242 0.152939
R20586 vdd.n2243 vdd.n1439 0.152939
R20587 vdd.n2260 vdd.n1439 0.152939
R20588 vdd.n2261 vdd.n2260 0.152939
R20589 vdd.n2262 vdd.n2261 0.152939
R20590 vdd.n735 vdd.n730 0.152939
R20591 vdd.n736 vdd.n735 0.152939
R20592 vdd.n737 vdd.n736 0.152939
R20593 vdd.n738 vdd.n737 0.152939
R20594 vdd.n739 vdd.n738 0.152939
R20595 vdd.n740 vdd.n739 0.152939
R20596 vdd.n741 vdd.n740 0.152939
R20597 vdd.n742 vdd.n741 0.152939
R20598 vdd.n743 vdd.n742 0.152939
R20599 vdd.n744 vdd.n743 0.152939
R20600 vdd.n745 vdd.n744 0.152939
R20601 vdd.n746 vdd.n745 0.152939
R20602 vdd.n3275 vdd.n746 0.152939
R20603 vdd.n3275 vdd.n3274 0.152939
R20604 vdd.n3274 vdd.n3273 0.152939
R20605 vdd.n3273 vdd.n748 0.152939
R20606 vdd.n749 vdd.n748 0.152939
R20607 vdd.n750 vdd.n749 0.152939
R20608 vdd.n751 vdd.n750 0.152939
R20609 vdd.n752 vdd.n751 0.152939
R20610 vdd.n753 vdd.n752 0.152939
R20611 vdd.n754 vdd.n753 0.152939
R20612 vdd.n755 vdd.n754 0.152939
R20613 vdd.n756 vdd.n755 0.152939
R20614 vdd.n757 vdd.n756 0.152939
R20615 vdd.n758 vdd.n757 0.152939
R20616 vdd.n759 vdd.n758 0.152939
R20617 vdd.n760 vdd.n759 0.152939
R20618 vdd.n761 vdd.n760 0.152939
R20619 vdd.n762 vdd.n761 0.152939
R20620 vdd.n763 vdd.n762 0.152939
R20621 vdd.n764 vdd.n763 0.152939
R20622 vdd.n765 vdd.n764 0.152939
R20623 vdd.n766 vdd.n765 0.152939
R20624 vdd.n3229 vdd.n766 0.152939
R20625 vdd.n3229 vdd.n3228 0.152939
R20626 vdd.n3228 vdd.n3227 0.152939
R20627 vdd.n3227 vdd.n770 0.152939
R20628 vdd.n771 vdd.n770 0.152939
R20629 vdd.n772 vdd.n771 0.152939
R20630 vdd.n773 vdd.n772 0.152939
R20631 vdd.n774 vdd.n773 0.152939
R20632 vdd.n775 vdd.n774 0.152939
R20633 vdd.n776 vdd.n775 0.152939
R20634 vdd.n777 vdd.n776 0.152939
R20635 vdd.n778 vdd.n777 0.152939
R20636 vdd.n779 vdd.n778 0.152939
R20637 vdd.n780 vdd.n779 0.152939
R20638 vdd.n781 vdd.n780 0.152939
R20639 vdd.n782 vdd.n781 0.152939
R20640 vdd.n783 vdd.n782 0.152939
R20641 vdd.n727 vdd.n726 0.152939
R20642 vdd.n3326 vdd.n682 0.152939
R20643 vdd.n3327 vdd.n3326 0.152939
R20644 vdd.n3328 vdd.n3327 0.152939
R20645 vdd.n3328 vdd.n670 0.152939
R20646 vdd.n3343 vdd.n670 0.152939
R20647 vdd.n3344 vdd.n3343 0.152939
R20648 vdd.n3345 vdd.n3344 0.152939
R20649 vdd.n3345 vdd.n659 0.152939
R20650 vdd.n3359 vdd.n659 0.152939
R20651 vdd.n3360 vdd.n3359 0.152939
R20652 vdd.n3361 vdd.n3360 0.152939
R20653 vdd.n3361 vdd.n647 0.152939
R20654 vdd.n3376 vdd.n647 0.152939
R20655 vdd.n3377 vdd.n3376 0.152939
R20656 vdd.n3378 vdd.n3377 0.152939
R20657 vdd.n3378 vdd.n636 0.152939
R20658 vdd.n3395 vdd.n636 0.152939
R20659 vdd.n3396 vdd.n3395 0.152939
R20660 vdd.n3397 vdd.n3396 0.152939
R20661 vdd.n3397 vdd.n334 0.152939
R20662 vdd.n3490 vdd.n335 0.152939
R20663 vdd.n346 vdd.n335 0.152939
R20664 vdd.n347 vdd.n346 0.152939
R20665 vdd.n348 vdd.n347 0.152939
R20666 vdd.n355 vdd.n348 0.152939
R20667 vdd.n356 vdd.n355 0.152939
R20668 vdd.n357 vdd.n356 0.152939
R20669 vdd.n358 vdd.n357 0.152939
R20670 vdd.n366 vdd.n358 0.152939
R20671 vdd.n367 vdd.n366 0.152939
R20672 vdd.n368 vdd.n367 0.152939
R20673 vdd.n369 vdd.n368 0.152939
R20674 vdd.n377 vdd.n369 0.152939
R20675 vdd.n378 vdd.n377 0.152939
R20676 vdd.n379 vdd.n378 0.152939
R20677 vdd.n380 vdd.n379 0.152939
R20678 vdd.n388 vdd.n380 0.152939
R20679 vdd.n389 vdd.n388 0.152939
R20680 vdd.n390 vdd.n389 0.152939
R20681 vdd.n391 vdd.n390 0.152939
R20682 vdd.n464 vdd.n463 0.152939
R20683 vdd.n470 vdd.n463 0.152939
R20684 vdd.n471 vdd.n470 0.152939
R20685 vdd.n472 vdd.n471 0.152939
R20686 vdd.n472 vdd.n461 0.152939
R20687 vdd.n480 vdd.n461 0.152939
R20688 vdd.n481 vdd.n480 0.152939
R20689 vdd.n482 vdd.n481 0.152939
R20690 vdd.n482 vdd.n459 0.152939
R20691 vdd.n490 vdd.n459 0.152939
R20692 vdd.n491 vdd.n490 0.152939
R20693 vdd.n492 vdd.n491 0.152939
R20694 vdd.n492 vdd.n457 0.152939
R20695 vdd.n500 vdd.n457 0.152939
R20696 vdd.n501 vdd.n500 0.152939
R20697 vdd.n502 vdd.n501 0.152939
R20698 vdd.n502 vdd.n455 0.152939
R20699 vdd.n510 vdd.n455 0.152939
R20700 vdd.n511 vdd.n510 0.152939
R20701 vdd.n512 vdd.n511 0.152939
R20702 vdd.n512 vdd.n451 0.152939
R20703 vdd.n520 vdd.n451 0.152939
R20704 vdd.n521 vdd.n520 0.152939
R20705 vdd.n522 vdd.n521 0.152939
R20706 vdd.n522 vdd.n449 0.152939
R20707 vdd.n530 vdd.n449 0.152939
R20708 vdd.n531 vdd.n530 0.152939
R20709 vdd.n532 vdd.n531 0.152939
R20710 vdd.n532 vdd.n447 0.152939
R20711 vdd.n540 vdd.n447 0.152939
R20712 vdd.n541 vdd.n540 0.152939
R20713 vdd.n542 vdd.n541 0.152939
R20714 vdd.n542 vdd.n445 0.152939
R20715 vdd.n550 vdd.n445 0.152939
R20716 vdd.n551 vdd.n550 0.152939
R20717 vdd.n552 vdd.n551 0.152939
R20718 vdd.n552 vdd.n443 0.152939
R20719 vdd.n560 vdd.n443 0.152939
R20720 vdd.n561 vdd.n560 0.152939
R20721 vdd.n562 vdd.n561 0.152939
R20722 vdd.n562 vdd.n439 0.152939
R20723 vdd.n570 vdd.n439 0.152939
R20724 vdd.n571 vdd.n570 0.152939
R20725 vdd.n572 vdd.n571 0.152939
R20726 vdd.n572 vdd.n437 0.152939
R20727 vdd.n580 vdd.n437 0.152939
R20728 vdd.n581 vdd.n580 0.152939
R20729 vdd.n582 vdd.n581 0.152939
R20730 vdd.n582 vdd.n435 0.152939
R20731 vdd.n590 vdd.n435 0.152939
R20732 vdd.n591 vdd.n590 0.152939
R20733 vdd.n592 vdd.n591 0.152939
R20734 vdd.n592 vdd.n433 0.152939
R20735 vdd.n600 vdd.n433 0.152939
R20736 vdd.n601 vdd.n600 0.152939
R20737 vdd.n602 vdd.n601 0.152939
R20738 vdd.n602 vdd.n431 0.152939
R20739 vdd.n610 vdd.n431 0.152939
R20740 vdd.n611 vdd.n610 0.152939
R20741 vdd.n612 vdd.n611 0.152939
R20742 vdd.n612 vdd.n429 0.152939
R20743 vdd.n619 vdd.n429 0.152939
R20744 vdd.n3442 vdd.n619 0.152939
R20745 vdd.n3320 vdd.n3319 0.152939
R20746 vdd.n3320 vdd.n675 0.152939
R20747 vdd.n3334 vdd.n675 0.152939
R20748 vdd.n3335 vdd.n3334 0.152939
R20749 vdd.n3336 vdd.n3335 0.152939
R20750 vdd.n3336 vdd.n665 0.152939
R20751 vdd.n3351 vdd.n665 0.152939
R20752 vdd.n3352 vdd.n3351 0.152939
R20753 vdd.n3353 vdd.n3352 0.152939
R20754 vdd.n3353 vdd.n652 0.152939
R20755 vdd.n3367 vdd.n652 0.152939
R20756 vdd.n3368 vdd.n3367 0.152939
R20757 vdd.n3369 vdd.n3368 0.152939
R20758 vdd.n3369 vdd.n641 0.152939
R20759 vdd.n3384 vdd.n641 0.152939
R20760 vdd.n3385 vdd.n3384 0.152939
R20761 vdd.n3386 vdd.n3385 0.152939
R20762 vdd.n3388 vdd.n3386 0.152939
R20763 vdd.n3388 vdd.n3387 0.152939
R20764 vdd.n3387 vdd.n630 0.152939
R20765 vdd.n3405 vdd.n630 0.152939
R20766 vdd.n3406 vdd.n3405 0.152939
R20767 vdd.n3407 vdd.n3406 0.152939
R20768 vdd.n3407 vdd.n628 0.152939
R20769 vdd.n3412 vdd.n628 0.152939
R20770 vdd.n3413 vdd.n3412 0.152939
R20771 vdd.n3414 vdd.n3413 0.152939
R20772 vdd.n3414 vdd.n626 0.152939
R20773 vdd.n3419 vdd.n626 0.152939
R20774 vdd.n3420 vdd.n3419 0.152939
R20775 vdd.n3421 vdd.n3420 0.152939
R20776 vdd.n3421 vdd.n624 0.152939
R20777 vdd.n3427 vdd.n624 0.152939
R20778 vdd.n3428 vdd.n3427 0.152939
R20779 vdd.n3429 vdd.n3428 0.152939
R20780 vdd.n3429 vdd.n622 0.152939
R20781 vdd.n3434 vdd.n622 0.152939
R20782 vdd.n3435 vdd.n3434 0.152939
R20783 vdd.n3436 vdd.n3435 0.152939
R20784 vdd.n3436 vdd.n620 0.152939
R20785 vdd.n3441 vdd.n620 0.152939
R20786 vdd.n3318 vdd.n687 0.152939
R20787 vdd.n2273 vdd.n1424 0.152939
R20788 vdd.n1792 vdd.n1548 0.152939
R20789 vdd.n1793 vdd.n1792 0.152939
R20790 vdd.n1794 vdd.n1793 0.152939
R20791 vdd.n1794 vdd.n1536 0.152939
R20792 vdd.n1809 vdd.n1536 0.152939
R20793 vdd.n1810 vdd.n1809 0.152939
R20794 vdd.n1811 vdd.n1810 0.152939
R20795 vdd.n1811 vdd.n1526 0.152939
R20796 vdd.n1826 vdd.n1526 0.152939
R20797 vdd.n1827 vdd.n1826 0.152939
R20798 vdd.n1828 vdd.n1827 0.152939
R20799 vdd.n1828 vdd.n1513 0.152939
R20800 vdd.n1842 vdd.n1513 0.152939
R20801 vdd.n1843 vdd.n1842 0.152939
R20802 vdd.n1844 vdd.n1843 0.152939
R20803 vdd.n1844 vdd.n1502 0.152939
R20804 vdd.n1859 vdd.n1502 0.152939
R20805 vdd.n1860 vdd.n1859 0.152939
R20806 vdd.n1861 vdd.n1860 0.152939
R20807 vdd.n1861 vdd.n1491 0.152939
R20808 vdd.n2182 vdd.n1491 0.152939
R20809 vdd.n2183 vdd.n2182 0.152939
R20810 vdd.n2184 vdd.n2183 0.152939
R20811 vdd.n2184 vdd.n1479 0.152939
R20812 vdd.n2199 vdd.n1479 0.152939
R20813 vdd.n2200 vdd.n2199 0.152939
R20814 vdd.n2201 vdd.n2200 0.152939
R20815 vdd.n2201 vdd.n1469 0.152939
R20816 vdd.n2216 vdd.n1469 0.152939
R20817 vdd.n2217 vdd.n2216 0.152939
R20818 vdd.n2218 vdd.n2217 0.152939
R20819 vdd.n2218 vdd.n1456 0.152939
R20820 vdd.n2232 vdd.n1456 0.152939
R20821 vdd.n2233 vdd.n2232 0.152939
R20822 vdd.n2234 vdd.n2233 0.152939
R20823 vdd.n2234 vdd.n1446 0.152939
R20824 vdd.n2249 vdd.n1446 0.152939
R20825 vdd.n2250 vdd.n2249 0.152939
R20826 vdd.n2253 vdd.n2250 0.152939
R20827 vdd.n2253 vdd.n2252 0.152939
R20828 vdd.n2252 vdd.n2251 0.152939
R20829 vdd.n1784 vdd.n1553 0.152939
R20830 vdd.n1777 vdd.n1553 0.152939
R20831 vdd.n1777 vdd.n1776 0.152939
R20832 vdd.n1776 vdd.n1775 0.152939
R20833 vdd.n1775 vdd.n1590 0.152939
R20834 vdd.n1771 vdd.n1590 0.152939
R20835 vdd.n1771 vdd.n1770 0.152939
R20836 vdd.n1770 vdd.n1769 0.152939
R20837 vdd.n1769 vdd.n1596 0.152939
R20838 vdd.n1765 vdd.n1596 0.152939
R20839 vdd.n1765 vdd.n1764 0.152939
R20840 vdd.n1764 vdd.n1763 0.152939
R20841 vdd.n1763 vdd.n1602 0.152939
R20842 vdd.n1759 vdd.n1602 0.152939
R20843 vdd.n1759 vdd.n1758 0.152939
R20844 vdd.n1758 vdd.n1757 0.152939
R20845 vdd.n1757 vdd.n1608 0.152939
R20846 vdd.n1753 vdd.n1608 0.152939
R20847 vdd.n1753 vdd.n1752 0.152939
R20848 vdd.n1752 vdd.n1751 0.152939
R20849 vdd.n1751 vdd.n1616 0.152939
R20850 vdd.n1747 vdd.n1616 0.152939
R20851 vdd.n1747 vdd.n1746 0.152939
R20852 vdd.n1746 vdd.n1745 0.152939
R20853 vdd.n1745 vdd.n1622 0.152939
R20854 vdd.n1741 vdd.n1622 0.152939
R20855 vdd.n1741 vdd.n1740 0.152939
R20856 vdd.n1740 vdd.n1739 0.152939
R20857 vdd.n1739 vdd.n1628 0.152939
R20858 vdd.n1735 vdd.n1628 0.152939
R20859 vdd.n1735 vdd.n1734 0.152939
R20860 vdd.n1734 vdd.n1733 0.152939
R20861 vdd.n1733 vdd.n1634 0.152939
R20862 vdd.n1729 vdd.n1634 0.152939
R20863 vdd.n1729 vdd.n1728 0.152939
R20864 vdd.n1728 vdd.n1727 0.152939
R20865 vdd.n1727 vdd.n1640 0.152939
R20866 vdd.n1723 vdd.n1640 0.152939
R20867 vdd.n1723 vdd.n1722 0.152939
R20868 vdd.n1722 vdd.n1721 0.152939
R20869 vdd.n1721 vdd.n1646 0.152939
R20870 vdd.n1714 vdd.n1646 0.152939
R20871 vdd.n1714 vdd.n1713 0.152939
R20872 vdd.n1713 vdd.n1712 0.152939
R20873 vdd.n1712 vdd.n1651 0.152939
R20874 vdd.n1708 vdd.n1651 0.152939
R20875 vdd.n1708 vdd.n1707 0.152939
R20876 vdd.n1707 vdd.n1706 0.152939
R20877 vdd.n1706 vdd.n1657 0.152939
R20878 vdd.n1702 vdd.n1657 0.152939
R20879 vdd.n1702 vdd.n1701 0.152939
R20880 vdd.n1701 vdd.n1700 0.152939
R20881 vdd.n1700 vdd.n1663 0.152939
R20882 vdd.n1696 vdd.n1663 0.152939
R20883 vdd.n1696 vdd.n1695 0.152939
R20884 vdd.n1695 vdd.n1694 0.152939
R20885 vdd.n1694 vdd.n1669 0.152939
R20886 vdd.n1690 vdd.n1669 0.152939
R20887 vdd.n1690 vdd.n1689 0.152939
R20888 vdd.n1689 vdd.n1688 0.152939
R20889 vdd.n1688 vdd.n1675 0.152939
R20890 vdd.n1684 vdd.n1675 0.152939
R20891 vdd.n1684 vdd.n1683 0.152939
R20892 vdd.n1786 vdd.n1785 0.152939
R20893 vdd.n1786 vdd.n1542 0.152939
R20894 vdd.n1801 vdd.n1542 0.152939
R20895 vdd.n1802 vdd.n1801 0.152939
R20896 vdd.n1803 vdd.n1802 0.152939
R20897 vdd.n1803 vdd.n1531 0.152939
R20898 vdd.n1818 vdd.n1531 0.152939
R20899 vdd.n1819 vdd.n1818 0.152939
R20900 vdd.n1820 vdd.n1819 0.152939
R20901 vdd.n1820 vdd.n1520 0.152939
R20902 vdd.n1834 vdd.n1520 0.152939
R20903 vdd.n1835 vdd.n1834 0.152939
R20904 vdd.n1836 vdd.n1835 0.152939
R20905 vdd.n1836 vdd.n1508 0.152939
R20906 vdd.n1851 vdd.n1508 0.152939
R20907 vdd.n1852 vdd.n1851 0.152939
R20908 vdd.n1853 vdd.n1852 0.152939
R20909 vdd.n1853 vdd.n1497 0.152939
R20910 vdd.n1867 vdd.n1497 0.152939
R20911 vdd.n1868 vdd.n1867 0.152939
R20912 vdd.n1789 vdd.t254 0.113865
R20913 vdd.t240 vdd.n386 0.113865
R20914 vdd.n2381 vdd.n2380 0.110256
R20915 vdd.n3308 vdd.n727 0.110256
R20916 vdd.n3185 vdd.n687 0.110256
R20917 vdd.n2274 vdd.n2273 0.110256
R20918 vdd.n2176 vdd.n2175 0.0695946
R20919 vdd.n3491 vdd.n334 0.0695946
R20920 vdd.n3491 vdd.n3490 0.0695946
R20921 vdd.n2175 vdd.n1868 0.0695946
R20922 vdd.n2381 vdd.n1120 0.0431829
R20923 vdd.n2274 vdd.n1220 0.0431829
R20924 vdd.n3308 vdd.n730 0.0431829
R20925 vdd.n3185 vdd.n783 0.0431829
R20926 vdd vdd.n28 0.00833333
R20927 CSoutput.n19 CSoutput.t188 184.661
R20928 CSoutput.n78 CSoutput.n77 165.8
R20929 CSoutput.n76 CSoutput.n0 165.8
R20930 CSoutput.n75 CSoutput.n74 165.8
R20931 CSoutput.n73 CSoutput.n72 165.8
R20932 CSoutput.n71 CSoutput.n2 165.8
R20933 CSoutput.n69 CSoutput.n68 165.8
R20934 CSoutput.n67 CSoutput.n3 165.8
R20935 CSoutput.n66 CSoutput.n65 165.8
R20936 CSoutput.n63 CSoutput.n4 165.8
R20937 CSoutput.n61 CSoutput.n60 165.8
R20938 CSoutput.n59 CSoutput.n5 165.8
R20939 CSoutput.n58 CSoutput.n57 165.8
R20940 CSoutput.n55 CSoutput.n6 165.8
R20941 CSoutput.n54 CSoutput.n53 165.8
R20942 CSoutput.n52 CSoutput.n51 165.8
R20943 CSoutput.n50 CSoutput.n8 165.8
R20944 CSoutput.n48 CSoutput.n47 165.8
R20945 CSoutput.n46 CSoutput.n9 165.8
R20946 CSoutput.n45 CSoutput.n44 165.8
R20947 CSoutput.n42 CSoutput.n10 165.8
R20948 CSoutput.n41 CSoutput.n40 165.8
R20949 CSoutput.n39 CSoutput.n38 165.8
R20950 CSoutput.n37 CSoutput.n12 165.8
R20951 CSoutput.n35 CSoutput.n34 165.8
R20952 CSoutput.n33 CSoutput.n13 165.8
R20953 CSoutput.n32 CSoutput.n31 165.8
R20954 CSoutput.n29 CSoutput.n14 165.8
R20955 CSoutput.n28 CSoutput.n27 165.8
R20956 CSoutput.n26 CSoutput.n25 165.8
R20957 CSoutput.n24 CSoutput.n16 165.8
R20958 CSoutput.n22 CSoutput.n21 165.8
R20959 CSoutput.n20 CSoutput.n17 165.8
R20960 CSoutput.n77 CSoutput.t189 162.194
R20961 CSoutput.n18 CSoutput.t190 120.501
R20962 CSoutput.n23 CSoutput.t198 120.501
R20963 CSoutput.n15 CSoutput.t194 120.501
R20964 CSoutput.n30 CSoutput.t191 120.501
R20965 CSoutput.n36 CSoutput.t201 120.501
R20966 CSoutput.n11 CSoutput.t204 120.501
R20967 CSoutput.n43 CSoutput.t193 120.501
R20968 CSoutput.n49 CSoutput.t205 120.501
R20969 CSoutput.n7 CSoutput.t184 120.501
R20970 CSoutput.n56 CSoutput.t200 120.501
R20971 CSoutput.n62 CSoutput.t192 120.501
R20972 CSoutput.n64 CSoutput.t186 120.501
R20973 CSoutput.n70 CSoutput.t203 120.501
R20974 CSoutput.n1 CSoutput.t197 120.501
R20975 CSoutput.n330 CSoutput.n328 103.469
R20976 CSoutput.n310 CSoutput.n308 103.469
R20977 CSoutput.n291 CSoutput.n289 103.469
R20978 CSoutput.n120 CSoutput.n118 103.469
R20979 CSoutput.n100 CSoutput.n98 103.469
R20980 CSoutput.n81 CSoutput.n79 103.469
R20981 CSoutput.n344 CSoutput.n343 103.111
R20982 CSoutput.n342 CSoutput.n341 103.111
R20983 CSoutput.n340 CSoutput.n339 103.111
R20984 CSoutput.n338 CSoutput.n337 103.111
R20985 CSoutput.n336 CSoutput.n335 103.111
R20986 CSoutput.n334 CSoutput.n333 103.111
R20987 CSoutput.n332 CSoutput.n331 103.111
R20988 CSoutput.n330 CSoutput.n329 103.111
R20989 CSoutput.n326 CSoutput.n325 103.111
R20990 CSoutput.n324 CSoutput.n323 103.111
R20991 CSoutput.n322 CSoutput.n321 103.111
R20992 CSoutput.n320 CSoutput.n319 103.111
R20993 CSoutput.n318 CSoutput.n317 103.111
R20994 CSoutput.n316 CSoutput.n315 103.111
R20995 CSoutput.n314 CSoutput.n313 103.111
R20996 CSoutput.n312 CSoutput.n311 103.111
R20997 CSoutput.n310 CSoutput.n309 103.111
R20998 CSoutput.n307 CSoutput.n306 103.111
R20999 CSoutput.n305 CSoutput.n304 103.111
R21000 CSoutput.n303 CSoutput.n302 103.111
R21001 CSoutput.n301 CSoutput.n300 103.111
R21002 CSoutput.n299 CSoutput.n298 103.111
R21003 CSoutput.n297 CSoutput.n296 103.111
R21004 CSoutput.n295 CSoutput.n294 103.111
R21005 CSoutput.n293 CSoutput.n292 103.111
R21006 CSoutput.n291 CSoutput.n290 103.111
R21007 CSoutput.n120 CSoutput.n119 103.111
R21008 CSoutput.n122 CSoutput.n121 103.111
R21009 CSoutput.n124 CSoutput.n123 103.111
R21010 CSoutput.n126 CSoutput.n125 103.111
R21011 CSoutput.n128 CSoutput.n127 103.111
R21012 CSoutput.n130 CSoutput.n129 103.111
R21013 CSoutput.n132 CSoutput.n131 103.111
R21014 CSoutput.n134 CSoutput.n133 103.111
R21015 CSoutput.n136 CSoutput.n135 103.111
R21016 CSoutput.n100 CSoutput.n99 103.111
R21017 CSoutput.n102 CSoutput.n101 103.111
R21018 CSoutput.n104 CSoutput.n103 103.111
R21019 CSoutput.n106 CSoutput.n105 103.111
R21020 CSoutput.n108 CSoutput.n107 103.111
R21021 CSoutput.n110 CSoutput.n109 103.111
R21022 CSoutput.n112 CSoutput.n111 103.111
R21023 CSoutput.n114 CSoutput.n113 103.111
R21024 CSoutput.n116 CSoutput.n115 103.111
R21025 CSoutput.n81 CSoutput.n80 103.111
R21026 CSoutput.n83 CSoutput.n82 103.111
R21027 CSoutput.n85 CSoutput.n84 103.111
R21028 CSoutput.n87 CSoutput.n86 103.111
R21029 CSoutput.n89 CSoutput.n88 103.111
R21030 CSoutput.n91 CSoutput.n90 103.111
R21031 CSoutput.n93 CSoutput.n92 103.111
R21032 CSoutput.n95 CSoutput.n94 103.111
R21033 CSoutput.n97 CSoutput.n96 103.111
R21034 CSoutput.n346 CSoutput.n345 103.111
R21035 CSoutput.n366 CSoutput.n364 81.5057
R21036 CSoutput.n351 CSoutput.n349 81.5057
R21037 CSoutput.n398 CSoutput.n396 81.5057
R21038 CSoutput.n383 CSoutput.n381 81.5057
R21039 CSoutput.n378 CSoutput.n377 80.9324
R21040 CSoutput.n376 CSoutput.n375 80.9324
R21041 CSoutput.n374 CSoutput.n373 80.9324
R21042 CSoutput.n372 CSoutput.n371 80.9324
R21043 CSoutput.n370 CSoutput.n369 80.9324
R21044 CSoutput.n368 CSoutput.n367 80.9324
R21045 CSoutput.n366 CSoutput.n365 80.9324
R21046 CSoutput.n363 CSoutput.n362 80.9324
R21047 CSoutput.n361 CSoutput.n360 80.9324
R21048 CSoutput.n359 CSoutput.n358 80.9324
R21049 CSoutput.n357 CSoutput.n356 80.9324
R21050 CSoutput.n355 CSoutput.n354 80.9324
R21051 CSoutput.n353 CSoutput.n352 80.9324
R21052 CSoutput.n351 CSoutput.n350 80.9324
R21053 CSoutput.n398 CSoutput.n397 80.9324
R21054 CSoutput.n400 CSoutput.n399 80.9324
R21055 CSoutput.n402 CSoutput.n401 80.9324
R21056 CSoutput.n404 CSoutput.n403 80.9324
R21057 CSoutput.n406 CSoutput.n405 80.9324
R21058 CSoutput.n408 CSoutput.n407 80.9324
R21059 CSoutput.n410 CSoutput.n409 80.9324
R21060 CSoutput.n383 CSoutput.n382 80.9324
R21061 CSoutput.n385 CSoutput.n384 80.9324
R21062 CSoutput.n387 CSoutput.n386 80.9324
R21063 CSoutput.n389 CSoutput.n388 80.9324
R21064 CSoutput.n391 CSoutput.n390 80.9324
R21065 CSoutput.n393 CSoutput.n392 80.9324
R21066 CSoutput.n395 CSoutput.n394 80.9324
R21067 CSoutput.n25 CSoutput.n24 48.1486
R21068 CSoutput.n69 CSoutput.n3 48.1486
R21069 CSoutput.n38 CSoutput.n37 48.1486
R21070 CSoutput.n42 CSoutput.n41 48.1486
R21071 CSoutput.n51 CSoutput.n50 48.1486
R21072 CSoutput.n55 CSoutput.n54 48.1486
R21073 CSoutput.n22 CSoutput.n17 46.462
R21074 CSoutput.n72 CSoutput.n71 46.462
R21075 CSoutput.n20 CSoutput.n19 44.9055
R21076 CSoutput.n29 CSoutput.n28 43.7635
R21077 CSoutput.n65 CSoutput.n63 43.7635
R21078 CSoutput.n35 CSoutput.n13 41.7396
R21079 CSoutput.n57 CSoutput.n5 41.7396
R21080 CSoutput.n44 CSoutput.n9 37.0171
R21081 CSoutput.n48 CSoutput.n9 37.0171
R21082 CSoutput.n76 CSoutput.n75 34.9932
R21083 CSoutput.n31 CSoutput.n13 32.2947
R21084 CSoutput.n61 CSoutput.n5 32.2947
R21085 CSoutput.n30 CSoutput.n29 29.6014
R21086 CSoutput.n63 CSoutput.n62 29.6014
R21087 CSoutput.n19 CSoutput.n18 28.4085
R21088 CSoutput.n18 CSoutput.n17 25.1176
R21089 CSoutput.n72 CSoutput.n1 25.1176
R21090 CSoutput.n43 CSoutput.n42 22.0922
R21091 CSoutput.n50 CSoutput.n49 22.0922
R21092 CSoutput.n77 CSoutput.n76 21.8586
R21093 CSoutput.n37 CSoutput.n36 18.9681
R21094 CSoutput.n56 CSoutput.n55 18.9681
R21095 CSoutput.n25 CSoutput.n15 17.6292
R21096 CSoutput.n64 CSoutput.n3 17.6292
R21097 CSoutput.n24 CSoutput.n23 15.844
R21098 CSoutput.n70 CSoutput.n69 15.844
R21099 CSoutput.n38 CSoutput.n11 14.5051
R21100 CSoutput.n54 CSoutput.n7 14.5051
R21101 CSoutput.n413 CSoutput.n78 11.6139
R21102 CSoutput.n41 CSoutput.n11 11.3811
R21103 CSoutput.n51 CSoutput.n7 11.3811
R21104 CSoutput.n23 CSoutput.n22 10.0422
R21105 CSoutput.n71 CSoutput.n70 10.0422
R21106 CSoutput.n327 CSoutput.n307 9.25285
R21107 CSoutput.n117 CSoutput.n97 9.25285
R21108 CSoutput.n379 CSoutput.n363 8.97993
R21109 CSoutput.n411 CSoutput.n395 8.97993
R21110 CSoutput.n380 CSoutput.n348 8.82395
R21111 CSoutput.n28 CSoutput.n15 8.25698
R21112 CSoutput.n65 CSoutput.n64 8.25698
R21113 CSoutput.n380 CSoutput.n379 7.89345
R21114 CSoutput.n412 CSoutput.n411 7.89345
R21115 CSoutput.n348 CSoutput.n347 7.12641
R21116 CSoutput.n138 CSoutput.n137 7.12641
R21117 CSoutput.n36 CSoutput.n35 6.91809
R21118 CSoutput.n57 CSoutput.n56 6.91809
R21119 CSoutput.n379 CSoutput.n378 5.25266
R21120 CSoutput.n411 CSoutput.n410 5.25266
R21121 CSoutput.n413 CSoutput.n138 5.23151
R21122 CSoutput.n347 CSoutput.n346 5.1449
R21123 CSoutput.n327 CSoutput.n326 5.1449
R21124 CSoutput.n137 CSoutput.n136 5.1449
R21125 CSoutput.n117 CSoutput.n116 5.1449
R21126 CSoutput.n229 CSoutput.n182 4.5005
R21127 CSoutput.n198 CSoutput.n182 4.5005
R21128 CSoutput.n193 CSoutput.n177 4.5005
R21129 CSoutput.n193 CSoutput.n179 4.5005
R21130 CSoutput.n193 CSoutput.n176 4.5005
R21131 CSoutput.n193 CSoutput.n180 4.5005
R21132 CSoutput.n193 CSoutput.n175 4.5005
R21133 CSoutput.n193 CSoutput.t199 4.5005
R21134 CSoutput.n193 CSoutput.n174 4.5005
R21135 CSoutput.n193 CSoutput.n181 4.5005
R21136 CSoutput.n193 CSoutput.n182 4.5005
R21137 CSoutput.n191 CSoutput.n177 4.5005
R21138 CSoutput.n191 CSoutput.n179 4.5005
R21139 CSoutput.n191 CSoutput.n176 4.5005
R21140 CSoutput.n191 CSoutput.n180 4.5005
R21141 CSoutput.n191 CSoutput.n175 4.5005
R21142 CSoutput.n191 CSoutput.t199 4.5005
R21143 CSoutput.n191 CSoutput.n174 4.5005
R21144 CSoutput.n191 CSoutput.n181 4.5005
R21145 CSoutput.n191 CSoutput.n182 4.5005
R21146 CSoutput.n190 CSoutput.n177 4.5005
R21147 CSoutput.n190 CSoutput.n179 4.5005
R21148 CSoutput.n190 CSoutput.n176 4.5005
R21149 CSoutput.n190 CSoutput.n180 4.5005
R21150 CSoutput.n190 CSoutput.n175 4.5005
R21151 CSoutput.n190 CSoutput.t199 4.5005
R21152 CSoutput.n190 CSoutput.n174 4.5005
R21153 CSoutput.n190 CSoutput.n181 4.5005
R21154 CSoutput.n190 CSoutput.n182 4.5005
R21155 CSoutput.n275 CSoutput.n177 4.5005
R21156 CSoutput.n275 CSoutput.n179 4.5005
R21157 CSoutput.n275 CSoutput.n176 4.5005
R21158 CSoutput.n275 CSoutput.n180 4.5005
R21159 CSoutput.n275 CSoutput.n175 4.5005
R21160 CSoutput.n275 CSoutput.t199 4.5005
R21161 CSoutput.n275 CSoutput.n174 4.5005
R21162 CSoutput.n275 CSoutput.n181 4.5005
R21163 CSoutput.n275 CSoutput.n182 4.5005
R21164 CSoutput.n273 CSoutput.n177 4.5005
R21165 CSoutput.n273 CSoutput.n179 4.5005
R21166 CSoutput.n273 CSoutput.n176 4.5005
R21167 CSoutput.n273 CSoutput.n180 4.5005
R21168 CSoutput.n273 CSoutput.n175 4.5005
R21169 CSoutput.n273 CSoutput.t199 4.5005
R21170 CSoutput.n273 CSoutput.n174 4.5005
R21171 CSoutput.n273 CSoutput.n181 4.5005
R21172 CSoutput.n271 CSoutput.n177 4.5005
R21173 CSoutput.n271 CSoutput.n179 4.5005
R21174 CSoutput.n271 CSoutput.n176 4.5005
R21175 CSoutput.n271 CSoutput.n180 4.5005
R21176 CSoutput.n271 CSoutput.n175 4.5005
R21177 CSoutput.n271 CSoutput.t199 4.5005
R21178 CSoutput.n271 CSoutput.n174 4.5005
R21179 CSoutput.n271 CSoutput.n181 4.5005
R21180 CSoutput.n201 CSoutput.n177 4.5005
R21181 CSoutput.n201 CSoutput.n179 4.5005
R21182 CSoutput.n201 CSoutput.n176 4.5005
R21183 CSoutput.n201 CSoutput.n180 4.5005
R21184 CSoutput.n201 CSoutput.n175 4.5005
R21185 CSoutput.n201 CSoutput.t199 4.5005
R21186 CSoutput.n201 CSoutput.n174 4.5005
R21187 CSoutput.n201 CSoutput.n181 4.5005
R21188 CSoutput.n201 CSoutput.n182 4.5005
R21189 CSoutput.n200 CSoutput.n177 4.5005
R21190 CSoutput.n200 CSoutput.n179 4.5005
R21191 CSoutput.n200 CSoutput.n176 4.5005
R21192 CSoutput.n200 CSoutput.n180 4.5005
R21193 CSoutput.n200 CSoutput.n175 4.5005
R21194 CSoutput.n200 CSoutput.t199 4.5005
R21195 CSoutput.n200 CSoutput.n174 4.5005
R21196 CSoutput.n200 CSoutput.n181 4.5005
R21197 CSoutput.n200 CSoutput.n182 4.5005
R21198 CSoutput.n204 CSoutput.n177 4.5005
R21199 CSoutput.n204 CSoutput.n179 4.5005
R21200 CSoutput.n204 CSoutput.n176 4.5005
R21201 CSoutput.n204 CSoutput.n180 4.5005
R21202 CSoutput.n204 CSoutput.n175 4.5005
R21203 CSoutput.n204 CSoutput.t199 4.5005
R21204 CSoutput.n204 CSoutput.n174 4.5005
R21205 CSoutput.n204 CSoutput.n181 4.5005
R21206 CSoutput.n204 CSoutput.n182 4.5005
R21207 CSoutput.n203 CSoutput.n177 4.5005
R21208 CSoutput.n203 CSoutput.n179 4.5005
R21209 CSoutput.n203 CSoutput.n176 4.5005
R21210 CSoutput.n203 CSoutput.n180 4.5005
R21211 CSoutput.n203 CSoutput.n175 4.5005
R21212 CSoutput.n203 CSoutput.t199 4.5005
R21213 CSoutput.n203 CSoutput.n174 4.5005
R21214 CSoutput.n203 CSoutput.n181 4.5005
R21215 CSoutput.n203 CSoutput.n182 4.5005
R21216 CSoutput.n186 CSoutput.n177 4.5005
R21217 CSoutput.n186 CSoutput.n179 4.5005
R21218 CSoutput.n186 CSoutput.n176 4.5005
R21219 CSoutput.n186 CSoutput.n180 4.5005
R21220 CSoutput.n186 CSoutput.n175 4.5005
R21221 CSoutput.n186 CSoutput.t199 4.5005
R21222 CSoutput.n186 CSoutput.n174 4.5005
R21223 CSoutput.n186 CSoutput.n181 4.5005
R21224 CSoutput.n186 CSoutput.n182 4.5005
R21225 CSoutput.n278 CSoutput.n177 4.5005
R21226 CSoutput.n278 CSoutput.n179 4.5005
R21227 CSoutput.n278 CSoutput.n176 4.5005
R21228 CSoutput.n278 CSoutput.n180 4.5005
R21229 CSoutput.n278 CSoutput.n175 4.5005
R21230 CSoutput.n278 CSoutput.t199 4.5005
R21231 CSoutput.n278 CSoutput.n174 4.5005
R21232 CSoutput.n278 CSoutput.n181 4.5005
R21233 CSoutput.n278 CSoutput.n182 4.5005
R21234 CSoutput.n265 CSoutput.n236 4.5005
R21235 CSoutput.n265 CSoutput.n242 4.5005
R21236 CSoutput.n223 CSoutput.n212 4.5005
R21237 CSoutput.n223 CSoutput.n214 4.5005
R21238 CSoutput.n223 CSoutput.n211 4.5005
R21239 CSoutput.n223 CSoutput.n215 4.5005
R21240 CSoutput.n223 CSoutput.n210 4.5005
R21241 CSoutput.n223 CSoutput.t195 4.5005
R21242 CSoutput.n223 CSoutput.n209 4.5005
R21243 CSoutput.n223 CSoutput.n216 4.5005
R21244 CSoutput.n265 CSoutput.n223 4.5005
R21245 CSoutput.n244 CSoutput.n212 4.5005
R21246 CSoutput.n244 CSoutput.n214 4.5005
R21247 CSoutput.n244 CSoutput.n211 4.5005
R21248 CSoutput.n244 CSoutput.n215 4.5005
R21249 CSoutput.n244 CSoutput.n210 4.5005
R21250 CSoutput.n244 CSoutput.t195 4.5005
R21251 CSoutput.n244 CSoutput.n209 4.5005
R21252 CSoutput.n244 CSoutput.n216 4.5005
R21253 CSoutput.n265 CSoutput.n244 4.5005
R21254 CSoutput.n222 CSoutput.n212 4.5005
R21255 CSoutput.n222 CSoutput.n214 4.5005
R21256 CSoutput.n222 CSoutput.n211 4.5005
R21257 CSoutput.n222 CSoutput.n215 4.5005
R21258 CSoutput.n222 CSoutput.n210 4.5005
R21259 CSoutput.n222 CSoutput.t195 4.5005
R21260 CSoutput.n222 CSoutput.n209 4.5005
R21261 CSoutput.n222 CSoutput.n216 4.5005
R21262 CSoutput.n265 CSoutput.n222 4.5005
R21263 CSoutput.n246 CSoutput.n212 4.5005
R21264 CSoutput.n246 CSoutput.n214 4.5005
R21265 CSoutput.n246 CSoutput.n211 4.5005
R21266 CSoutput.n246 CSoutput.n215 4.5005
R21267 CSoutput.n246 CSoutput.n210 4.5005
R21268 CSoutput.n246 CSoutput.t195 4.5005
R21269 CSoutput.n246 CSoutput.n209 4.5005
R21270 CSoutput.n246 CSoutput.n216 4.5005
R21271 CSoutput.n265 CSoutput.n246 4.5005
R21272 CSoutput.n212 CSoutput.n207 4.5005
R21273 CSoutput.n214 CSoutput.n207 4.5005
R21274 CSoutput.n211 CSoutput.n207 4.5005
R21275 CSoutput.n215 CSoutput.n207 4.5005
R21276 CSoutput.n210 CSoutput.n207 4.5005
R21277 CSoutput.t195 CSoutput.n207 4.5005
R21278 CSoutput.n209 CSoutput.n207 4.5005
R21279 CSoutput.n216 CSoutput.n207 4.5005
R21280 CSoutput.n268 CSoutput.n212 4.5005
R21281 CSoutput.n268 CSoutput.n214 4.5005
R21282 CSoutput.n268 CSoutput.n211 4.5005
R21283 CSoutput.n268 CSoutput.n215 4.5005
R21284 CSoutput.n268 CSoutput.n210 4.5005
R21285 CSoutput.n268 CSoutput.t195 4.5005
R21286 CSoutput.n268 CSoutput.n209 4.5005
R21287 CSoutput.n268 CSoutput.n216 4.5005
R21288 CSoutput.n266 CSoutput.n212 4.5005
R21289 CSoutput.n266 CSoutput.n214 4.5005
R21290 CSoutput.n266 CSoutput.n211 4.5005
R21291 CSoutput.n266 CSoutput.n215 4.5005
R21292 CSoutput.n266 CSoutput.n210 4.5005
R21293 CSoutput.n266 CSoutput.t195 4.5005
R21294 CSoutput.n266 CSoutput.n209 4.5005
R21295 CSoutput.n266 CSoutput.n216 4.5005
R21296 CSoutput.n266 CSoutput.n265 4.5005
R21297 CSoutput.n248 CSoutput.n212 4.5005
R21298 CSoutput.n248 CSoutput.n214 4.5005
R21299 CSoutput.n248 CSoutput.n211 4.5005
R21300 CSoutput.n248 CSoutput.n215 4.5005
R21301 CSoutput.n248 CSoutput.n210 4.5005
R21302 CSoutput.n248 CSoutput.t195 4.5005
R21303 CSoutput.n248 CSoutput.n209 4.5005
R21304 CSoutput.n248 CSoutput.n216 4.5005
R21305 CSoutput.n265 CSoutput.n248 4.5005
R21306 CSoutput.n220 CSoutput.n212 4.5005
R21307 CSoutput.n220 CSoutput.n214 4.5005
R21308 CSoutput.n220 CSoutput.n211 4.5005
R21309 CSoutput.n220 CSoutput.n215 4.5005
R21310 CSoutput.n220 CSoutput.n210 4.5005
R21311 CSoutput.n220 CSoutput.t195 4.5005
R21312 CSoutput.n220 CSoutput.n209 4.5005
R21313 CSoutput.n220 CSoutput.n216 4.5005
R21314 CSoutput.n265 CSoutput.n220 4.5005
R21315 CSoutput.n250 CSoutput.n212 4.5005
R21316 CSoutput.n250 CSoutput.n214 4.5005
R21317 CSoutput.n250 CSoutput.n211 4.5005
R21318 CSoutput.n250 CSoutput.n215 4.5005
R21319 CSoutput.n250 CSoutput.n210 4.5005
R21320 CSoutput.n250 CSoutput.t195 4.5005
R21321 CSoutput.n250 CSoutput.n209 4.5005
R21322 CSoutput.n250 CSoutput.n216 4.5005
R21323 CSoutput.n265 CSoutput.n250 4.5005
R21324 CSoutput.n219 CSoutput.n212 4.5005
R21325 CSoutput.n219 CSoutput.n214 4.5005
R21326 CSoutput.n219 CSoutput.n211 4.5005
R21327 CSoutput.n219 CSoutput.n215 4.5005
R21328 CSoutput.n219 CSoutput.n210 4.5005
R21329 CSoutput.n219 CSoutput.t195 4.5005
R21330 CSoutput.n219 CSoutput.n209 4.5005
R21331 CSoutput.n219 CSoutput.n216 4.5005
R21332 CSoutput.n265 CSoutput.n219 4.5005
R21333 CSoutput.n264 CSoutput.n212 4.5005
R21334 CSoutput.n264 CSoutput.n214 4.5005
R21335 CSoutput.n264 CSoutput.n211 4.5005
R21336 CSoutput.n264 CSoutput.n215 4.5005
R21337 CSoutput.n264 CSoutput.n210 4.5005
R21338 CSoutput.n264 CSoutput.t195 4.5005
R21339 CSoutput.n264 CSoutput.n209 4.5005
R21340 CSoutput.n264 CSoutput.n216 4.5005
R21341 CSoutput.n265 CSoutput.n264 4.5005
R21342 CSoutput.n263 CSoutput.n148 4.5005
R21343 CSoutput.n164 CSoutput.n148 4.5005
R21344 CSoutput.n159 CSoutput.n143 4.5005
R21345 CSoutput.n159 CSoutput.n145 4.5005
R21346 CSoutput.n159 CSoutput.n142 4.5005
R21347 CSoutput.n159 CSoutput.n146 4.5005
R21348 CSoutput.n159 CSoutput.n141 4.5005
R21349 CSoutput.n159 CSoutput.t185 4.5005
R21350 CSoutput.n159 CSoutput.n140 4.5005
R21351 CSoutput.n159 CSoutput.n147 4.5005
R21352 CSoutput.n159 CSoutput.n148 4.5005
R21353 CSoutput.n157 CSoutput.n143 4.5005
R21354 CSoutput.n157 CSoutput.n145 4.5005
R21355 CSoutput.n157 CSoutput.n142 4.5005
R21356 CSoutput.n157 CSoutput.n146 4.5005
R21357 CSoutput.n157 CSoutput.n141 4.5005
R21358 CSoutput.n157 CSoutput.t185 4.5005
R21359 CSoutput.n157 CSoutput.n140 4.5005
R21360 CSoutput.n157 CSoutput.n147 4.5005
R21361 CSoutput.n157 CSoutput.n148 4.5005
R21362 CSoutput.n156 CSoutput.n143 4.5005
R21363 CSoutput.n156 CSoutput.n145 4.5005
R21364 CSoutput.n156 CSoutput.n142 4.5005
R21365 CSoutput.n156 CSoutput.n146 4.5005
R21366 CSoutput.n156 CSoutput.n141 4.5005
R21367 CSoutput.n156 CSoutput.t185 4.5005
R21368 CSoutput.n156 CSoutput.n140 4.5005
R21369 CSoutput.n156 CSoutput.n147 4.5005
R21370 CSoutput.n156 CSoutput.n148 4.5005
R21371 CSoutput.n285 CSoutput.n143 4.5005
R21372 CSoutput.n285 CSoutput.n145 4.5005
R21373 CSoutput.n285 CSoutput.n142 4.5005
R21374 CSoutput.n285 CSoutput.n146 4.5005
R21375 CSoutput.n285 CSoutput.n141 4.5005
R21376 CSoutput.n285 CSoutput.t185 4.5005
R21377 CSoutput.n285 CSoutput.n140 4.5005
R21378 CSoutput.n285 CSoutput.n147 4.5005
R21379 CSoutput.n285 CSoutput.n148 4.5005
R21380 CSoutput.n283 CSoutput.n143 4.5005
R21381 CSoutput.n283 CSoutput.n145 4.5005
R21382 CSoutput.n283 CSoutput.n142 4.5005
R21383 CSoutput.n283 CSoutput.n146 4.5005
R21384 CSoutput.n283 CSoutput.n141 4.5005
R21385 CSoutput.n283 CSoutput.t185 4.5005
R21386 CSoutput.n283 CSoutput.n140 4.5005
R21387 CSoutput.n283 CSoutput.n147 4.5005
R21388 CSoutput.n281 CSoutput.n143 4.5005
R21389 CSoutput.n281 CSoutput.n145 4.5005
R21390 CSoutput.n281 CSoutput.n142 4.5005
R21391 CSoutput.n281 CSoutput.n146 4.5005
R21392 CSoutput.n281 CSoutput.n141 4.5005
R21393 CSoutput.n281 CSoutput.t185 4.5005
R21394 CSoutput.n281 CSoutput.n140 4.5005
R21395 CSoutput.n281 CSoutput.n147 4.5005
R21396 CSoutput.n167 CSoutput.n143 4.5005
R21397 CSoutput.n167 CSoutput.n145 4.5005
R21398 CSoutput.n167 CSoutput.n142 4.5005
R21399 CSoutput.n167 CSoutput.n146 4.5005
R21400 CSoutput.n167 CSoutput.n141 4.5005
R21401 CSoutput.n167 CSoutput.t185 4.5005
R21402 CSoutput.n167 CSoutput.n140 4.5005
R21403 CSoutput.n167 CSoutput.n147 4.5005
R21404 CSoutput.n167 CSoutput.n148 4.5005
R21405 CSoutput.n166 CSoutput.n143 4.5005
R21406 CSoutput.n166 CSoutput.n145 4.5005
R21407 CSoutput.n166 CSoutput.n142 4.5005
R21408 CSoutput.n166 CSoutput.n146 4.5005
R21409 CSoutput.n166 CSoutput.n141 4.5005
R21410 CSoutput.n166 CSoutput.t185 4.5005
R21411 CSoutput.n166 CSoutput.n140 4.5005
R21412 CSoutput.n166 CSoutput.n147 4.5005
R21413 CSoutput.n166 CSoutput.n148 4.5005
R21414 CSoutput.n170 CSoutput.n143 4.5005
R21415 CSoutput.n170 CSoutput.n145 4.5005
R21416 CSoutput.n170 CSoutput.n142 4.5005
R21417 CSoutput.n170 CSoutput.n146 4.5005
R21418 CSoutput.n170 CSoutput.n141 4.5005
R21419 CSoutput.n170 CSoutput.t185 4.5005
R21420 CSoutput.n170 CSoutput.n140 4.5005
R21421 CSoutput.n170 CSoutput.n147 4.5005
R21422 CSoutput.n170 CSoutput.n148 4.5005
R21423 CSoutput.n169 CSoutput.n143 4.5005
R21424 CSoutput.n169 CSoutput.n145 4.5005
R21425 CSoutput.n169 CSoutput.n142 4.5005
R21426 CSoutput.n169 CSoutput.n146 4.5005
R21427 CSoutput.n169 CSoutput.n141 4.5005
R21428 CSoutput.n169 CSoutput.t185 4.5005
R21429 CSoutput.n169 CSoutput.n140 4.5005
R21430 CSoutput.n169 CSoutput.n147 4.5005
R21431 CSoutput.n169 CSoutput.n148 4.5005
R21432 CSoutput.n152 CSoutput.n143 4.5005
R21433 CSoutput.n152 CSoutput.n145 4.5005
R21434 CSoutput.n152 CSoutput.n142 4.5005
R21435 CSoutput.n152 CSoutput.n146 4.5005
R21436 CSoutput.n152 CSoutput.n141 4.5005
R21437 CSoutput.n152 CSoutput.t185 4.5005
R21438 CSoutput.n152 CSoutput.n140 4.5005
R21439 CSoutput.n152 CSoutput.n147 4.5005
R21440 CSoutput.n152 CSoutput.n148 4.5005
R21441 CSoutput.n288 CSoutput.n143 4.5005
R21442 CSoutput.n288 CSoutput.n145 4.5005
R21443 CSoutput.n288 CSoutput.n142 4.5005
R21444 CSoutput.n288 CSoutput.n146 4.5005
R21445 CSoutput.n288 CSoutput.n141 4.5005
R21446 CSoutput.n288 CSoutput.t185 4.5005
R21447 CSoutput.n288 CSoutput.n140 4.5005
R21448 CSoutput.n288 CSoutput.n147 4.5005
R21449 CSoutput.n288 CSoutput.n148 4.5005
R21450 CSoutput.n347 CSoutput.n327 4.10845
R21451 CSoutput.n137 CSoutput.n117 4.10845
R21452 CSoutput.n345 CSoutput.t97 4.06363
R21453 CSoutput.n345 CSoutput.t15 4.06363
R21454 CSoutput.n343 CSoutput.t8 4.06363
R21455 CSoutput.n343 CSoutput.t59 4.06363
R21456 CSoutput.n341 CSoutput.t76 4.06363
R21457 CSoutput.n341 CSoutput.t100 4.06363
R21458 CSoutput.n339 CSoutput.t115 4.06363
R21459 CSoutput.n339 CSoutput.t28 4.06363
R21460 CSoutput.n337 CSoutput.t32 4.06363
R21461 CSoutput.n337 CSoutput.t104 4.06363
R21462 CSoutput.n335 CSoutput.t119 4.06363
R21463 CSoutput.n335 CSoutput.t120 4.06363
R21464 CSoutput.n333 CSoutput.t53 4.06363
R21465 CSoutput.n333 CSoutput.t54 4.06363
R21466 CSoutput.n331 CSoutput.t61 4.06363
R21467 CSoutput.n331 CSoutput.t121 4.06363
R21468 CSoutput.n329 CSoutput.t20 4.06363
R21469 CSoutput.n329 CSoutput.t58 4.06363
R21470 CSoutput.n328 CSoutput.t75 4.06363
R21471 CSoutput.n328 CSoutput.t99 4.06363
R21472 CSoutput.n325 CSoutput.t86 4.06363
R21473 CSoutput.n325 CSoutput.t122 4.06363
R21474 CSoutput.n323 CSoutput.t117 4.06363
R21475 CSoutput.n323 CSoutput.t42 4.06363
R21476 CSoutput.n321 CSoutput.t63 4.06363
R21477 CSoutput.n321 CSoutput.t87 4.06363
R21478 CSoutput.n319 CSoutput.t105 4.06363
R21479 CSoutput.n319 CSoutput.t14 4.06363
R21480 CSoutput.n317 CSoutput.t16 4.06363
R21481 CSoutput.n317 CSoutput.t91 4.06363
R21482 CSoutput.n315 CSoutput.t108 4.06363
R21483 CSoutput.n315 CSoutput.t109 4.06363
R21484 CSoutput.n313 CSoutput.t36 4.06363
R21485 CSoutput.n313 CSoutput.t37 4.06363
R21486 CSoutput.n311 CSoutput.t44 4.06363
R21487 CSoutput.n311 CSoutput.t110 4.06363
R21488 CSoutput.n309 CSoutput.t6 4.06363
R21489 CSoutput.n309 CSoutput.t43 4.06363
R21490 CSoutput.n308 CSoutput.t64 4.06363
R21491 CSoutput.n308 CSoutput.t88 4.06363
R21492 CSoutput.n306 CSoutput.t89 4.06363
R21493 CSoutput.n306 CSoutput.t40 4.06363
R21494 CSoutput.n304 CSoutput.t111 4.06363
R21495 CSoutput.n304 CSoutput.t68 4.06363
R21496 CSoutput.n302 CSoutput.t98 4.06363
R21497 CSoutput.n302 CSoutput.t50 4.06363
R21498 CSoutput.n300 CSoutput.t82 4.06363
R21499 CSoutput.n300 CSoutput.t27 4.06363
R21500 CSoutput.n298 CSoutput.t106 4.06363
R21501 CSoutput.n298 CSoutput.t21 4.06363
R21502 CSoutput.n296 CSoutput.t65 4.06363
R21503 CSoutput.n296 CSoutput.t38 4.06363
R21504 CSoutput.n294 CSoutput.t45 4.06363
R21505 CSoutput.n294 CSoutput.t17 4.06363
R21506 CSoutput.n292 CSoutput.t96 4.06363
R21507 CSoutput.n292 CSoutput.t11 4.06363
R21508 CSoutput.n290 CSoutput.t55 4.06363
R21509 CSoutput.n290 CSoutput.t116 4.06363
R21510 CSoutput.n289 CSoutput.t33 4.06363
R21511 CSoutput.n289 CSoutput.t102 4.06363
R21512 CSoutput.n118 CSoutput.t24 4.06363
R21513 CSoutput.n118 CSoutput.t113 4.06363
R21514 CSoutput.n119 CSoutput.t94 4.06363
R21515 CSoutput.n119 CSoutput.t72 4.06363
R21516 CSoutput.n121 CSoutput.t52 4.06363
R21517 CSoutput.n121 CSoutput.t124 4.06363
R21518 CSoutput.n123 CSoutput.t93 4.06363
R21519 CSoutput.n123 CSoutput.t92 4.06363
R21520 CSoutput.n125 CSoutput.t78 4.06363
R21521 CSoutput.n125 CSoutput.t49 4.06363
R21522 CSoutput.n127 CSoutput.t26 4.06363
R21523 CSoutput.n127 CSoutput.t79 4.06363
R21524 CSoutput.n129 CSoutput.t77 4.06363
R21525 CSoutput.n129 CSoutput.t46 4.06363
R21526 CSoutput.n131 CSoutput.t25 4.06363
R21527 CSoutput.n131 CSoutput.t23 4.06363
R21528 CSoutput.n133 CSoutput.t95 4.06363
R21529 CSoutput.n133 CSoutput.t62 4.06363
R21530 CSoutput.n135 CSoutput.t57 4.06363
R21531 CSoutput.n135 CSoutput.t18 4.06363
R21532 CSoutput.n98 CSoutput.t9 4.06363
R21533 CSoutput.n98 CSoutput.t101 4.06363
R21534 CSoutput.n99 CSoutput.t84 4.06363
R21535 CSoutput.n99 CSoutput.t60 4.06363
R21536 CSoutput.n101 CSoutput.t35 4.06363
R21537 CSoutput.n101 CSoutput.t114 4.06363
R21538 CSoutput.n103 CSoutput.t81 4.06363
R21539 CSoutput.n103 CSoutput.t80 4.06363
R21540 CSoutput.n105 CSoutput.t70 4.06363
R21541 CSoutput.n105 CSoutput.t31 4.06363
R21542 CSoutput.n107 CSoutput.t12 4.06363
R21543 CSoutput.n107 CSoutput.t71 4.06363
R21544 CSoutput.n109 CSoutput.t67 4.06363
R21545 CSoutput.n109 CSoutput.t29 4.06363
R21546 CSoutput.n111 CSoutput.t10 4.06363
R21547 CSoutput.n111 CSoutput.t7 4.06363
R21548 CSoutput.n113 CSoutput.t85 4.06363
R21549 CSoutput.n113 CSoutput.t48 4.06363
R21550 CSoutput.n115 CSoutput.t41 4.06363
R21551 CSoutput.n115 CSoutput.t5 4.06363
R21552 CSoutput.n79 CSoutput.t103 4.06363
R21553 CSoutput.n79 CSoutput.t34 4.06363
R21554 CSoutput.n80 CSoutput.t118 4.06363
R21555 CSoutput.n80 CSoutput.t56 4.06363
R21556 CSoutput.n82 CSoutput.t13 4.06363
R21557 CSoutput.n82 CSoutput.t73 4.06363
R21558 CSoutput.n84 CSoutput.t19 4.06363
R21559 CSoutput.n84 CSoutput.t47 4.06363
R21560 CSoutput.n86 CSoutput.t123 4.06363
R21561 CSoutput.n86 CSoutput.t66 4.06363
R21562 CSoutput.n88 CSoutput.t22 4.06363
R21563 CSoutput.n88 CSoutput.t107 4.06363
R21564 CSoutput.n90 CSoutput.t30 4.06363
R21565 CSoutput.n90 CSoutput.t83 4.06363
R21566 CSoutput.n92 CSoutput.t51 4.06363
R21567 CSoutput.n92 CSoutput.t74 4.06363
R21568 CSoutput.n94 CSoutput.t69 4.06363
R21569 CSoutput.n94 CSoutput.t112 4.06363
R21570 CSoutput.n96 CSoutput.t39 4.06363
R21571 CSoutput.n96 CSoutput.t90 4.06363
R21572 CSoutput.n44 CSoutput.n43 3.79402
R21573 CSoutput.n49 CSoutput.n48 3.79402
R21574 CSoutput.n413 CSoutput.n412 3.57343
R21575 CSoutput.n412 CSoutput.n380 3.3798
R21576 CSoutput.n377 CSoutput.t156 2.82907
R21577 CSoutput.n377 CSoutput.t133 2.82907
R21578 CSoutput.n375 CSoutput.t4 2.82907
R21579 CSoutput.n375 CSoutput.t141 2.82907
R21580 CSoutput.n373 CSoutput.t164 2.82907
R21581 CSoutput.n373 CSoutput.t149 2.82907
R21582 CSoutput.n371 CSoutput.t180 2.82907
R21583 CSoutput.n371 CSoutput.t147 2.82907
R21584 CSoutput.n369 CSoutput.t171 2.82907
R21585 CSoutput.n369 CSoutput.t174 2.82907
R21586 CSoutput.n367 CSoutput.t139 2.82907
R21587 CSoutput.n367 CSoutput.t162 2.82907
R21588 CSoutput.n365 CSoutput.t148 2.82907
R21589 CSoutput.n365 CSoutput.t151 2.82907
R21590 CSoutput.n364 CSoutput.t181 2.82907
R21591 CSoutput.n364 CSoutput.t2 2.82907
R21592 CSoutput.n362 CSoutput.t3 2.82907
R21593 CSoutput.n362 CSoutput.t169 2.82907
R21594 CSoutput.n360 CSoutput.t160 2.82907
R21595 CSoutput.n360 CSoutput.t137 2.82907
R21596 CSoutput.n358 CSoutput.t140 2.82907
R21597 CSoutput.n358 CSoutput.t132 2.82907
R21598 CSoutput.n356 CSoutput.t182 2.82907
R21599 CSoutput.n356 CSoutput.t176 2.82907
R21600 CSoutput.n354 CSoutput.t170 2.82907
R21601 CSoutput.n354 CSoutput.t155 2.82907
R21602 CSoutput.n352 CSoutput.t163 2.82907
R21603 CSoutput.n352 CSoutput.t146 2.82907
R21604 CSoutput.n350 CSoutput.t154 2.82907
R21605 CSoutput.n350 CSoutput.t142 2.82907
R21606 CSoutput.n349 CSoutput.t129 2.82907
R21607 CSoutput.n349 CSoutput.t159 2.82907
R21608 CSoutput.n396 CSoutput.t168 2.82907
R21609 CSoutput.n396 CSoutput.t127 2.82907
R21610 CSoutput.n397 CSoutput.t138 2.82907
R21611 CSoutput.n397 CSoutput.t144 2.82907
R21612 CSoutput.n399 CSoutput.t153 2.82907
R21613 CSoutput.n399 CSoutput.t179 2.82907
R21614 CSoutput.n401 CSoutput.t150 2.82907
R21615 CSoutput.n401 CSoutput.t130 2.82907
R21616 CSoutput.n403 CSoutput.t134 2.82907
R21617 CSoutput.n403 CSoutput.t158 2.82907
R21618 CSoutput.n405 CSoutput.t131 2.82907
R21619 CSoutput.n405 CSoutput.t125 2.82907
R21620 CSoutput.n407 CSoutput.t136 2.82907
R21621 CSoutput.n407 CSoutput.t178 2.82907
R21622 CSoutput.n409 CSoutput.t177 2.82907
R21623 CSoutput.n409 CSoutput.t183 2.82907
R21624 CSoutput.n381 CSoutput.t166 2.82907
R21625 CSoutput.n381 CSoutput.t157 2.82907
R21626 CSoutput.n382 CSoutput.t173 2.82907
R21627 CSoutput.n382 CSoutput.t172 2.82907
R21628 CSoutput.n384 CSoutput.t175 2.82907
R21629 CSoutput.n384 CSoutput.t1 2.82907
R21630 CSoutput.n386 CSoutput.t126 2.82907
R21631 CSoutput.n386 CSoutput.t143 2.82907
R21632 CSoutput.n388 CSoutput.t152 2.82907
R21633 CSoutput.n388 CSoutput.t145 2.82907
R21634 CSoutput.n390 CSoutput.t135 2.82907
R21635 CSoutput.n390 CSoutput.t128 2.82907
R21636 CSoutput.n392 CSoutput.t165 2.82907
R21637 CSoutput.n392 CSoutput.t167 2.82907
R21638 CSoutput.n394 CSoutput.t0 2.82907
R21639 CSoutput.n394 CSoutput.t161 2.82907
R21640 CSoutput.n348 CSoutput.n138 2.78353
R21641 CSoutput.n75 CSoutput.n1 2.45513
R21642 CSoutput.n229 CSoutput.n227 2.251
R21643 CSoutput.n229 CSoutput.n226 2.251
R21644 CSoutput.n229 CSoutput.n225 2.251
R21645 CSoutput.n229 CSoutput.n224 2.251
R21646 CSoutput.n198 CSoutput.n197 2.251
R21647 CSoutput.n198 CSoutput.n196 2.251
R21648 CSoutput.n198 CSoutput.n195 2.251
R21649 CSoutput.n198 CSoutput.n194 2.251
R21650 CSoutput.n271 CSoutput.n270 2.251
R21651 CSoutput.n236 CSoutput.n234 2.251
R21652 CSoutput.n236 CSoutput.n233 2.251
R21653 CSoutput.n236 CSoutput.n232 2.251
R21654 CSoutput.n254 CSoutput.n236 2.251
R21655 CSoutput.n242 CSoutput.n241 2.251
R21656 CSoutput.n242 CSoutput.n240 2.251
R21657 CSoutput.n242 CSoutput.n239 2.251
R21658 CSoutput.n242 CSoutput.n238 2.251
R21659 CSoutput.n268 CSoutput.n208 2.251
R21660 CSoutput.n263 CSoutput.n261 2.251
R21661 CSoutput.n263 CSoutput.n260 2.251
R21662 CSoutput.n263 CSoutput.n259 2.251
R21663 CSoutput.n263 CSoutput.n258 2.251
R21664 CSoutput.n164 CSoutput.n163 2.251
R21665 CSoutput.n164 CSoutput.n162 2.251
R21666 CSoutput.n164 CSoutput.n161 2.251
R21667 CSoutput.n164 CSoutput.n160 2.251
R21668 CSoutput.n281 CSoutput.n280 2.251
R21669 CSoutput.n198 CSoutput.n178 2.2505
R21670 CSoutput.n193 CSoutput.n178 2.2505
R21671 CSoutput.n191 CSoutput.n178 2.2505
R21672 CSoutput.n190 CSoutput.n178 2.2505
R21673 CSoutput.n275 CSoutput.n178 2.2505
R21674 CSoutput.n273 CSoutput.n178 2.2505
R21675 CSoutput.n271 CSoutput.n178 2.2505
R21676 CSoutput.n201 CSoutput.n178 2.2505
R21677 CSoutput.n200 CSoutput.n178 2.2505
R21678 CSoutput.n204 CSoutput.n178 2.2505
R21679 CSoutput.n203 CSoutput.n178 2.2505
R21680 CSoutput.n186 CSoutput.n178 2.2505
R21681 CSoutput.n278 CSoutput.n178 2.2505
R21682 CSoutput.n278 CSoutput.n277 2.2505
R21683 CSoutput.n242 CSoutput.n213 2.2505
R21684 CSoutput.n223 CSoutput.n213 2.2505
R21685 CSoutput.n244 CSoutput.n213 2.2505
R21686 CSoutput.n222 CSoutput.n213 2.2505
R21687 CSoutput.n246 CSoutput.n213 2.2505
R21688 CSoutput.n213 CSoutput.n207 2.2505
R21689 CSoutput.n268 CSoutput.n213 2.2505
R21690 CSoutput.n266 CSoutput.n213 2.2505
R21691 CSoutput.n248 CSoutput.n213 2.2505
R21692 CSoutput.n220 CSoutput.n213 2.2505
R21693 CSoutput.n250 CSoutput.n213 2.2505
R21694 CSoutput.n219 CSoutput.n213 2.2505
R21695 CSoutput.n264 CSoutput.n213 2.2505
R21696 CSoutput.n264 CSoutput.n217 2.2505
R21697 CSoutput.n164 CSoutput.n144 2.2505
R21698 CSoutput.n159 CSoutput.n144 2.2505
R21699 CSoutput.n157 CSoutput.n144 2.2505
R21700 CSoutput.n156 CSoutput.n144 2.2505
R21701 CSoutput.n285 CSoutput.n144 2.2505
R21702 CSoutput.n283 CSoutput.n144 2.2505
R21703 CSoutput.n281 CSoutput.n144 2.2505
R21704 CSoutput.n167 CSoutput.n144 2.2505
R21705 CSoutput.n166 CSoutput.n144 2.2505
R21706 CSoutput.n170 CSoutput.n144 2.2505
R21707 CSoutput.n169 CSoutput.n144 2.2505
R21708 CSoutput.n152 CSoutput.n144 2.2505
R21709 CSoutput.n288 CSoutput.n144 2.2505
R21710 CSoutput.n288 CSoutput.n287 2.2505
R21711 CSoutput.n206 CSoutput.n199 2.25024
R21712 CSoutput.n206 CSoutput.n192 2.25024
R21713 CSoutput.n274 CSoutput.n206 2.25024
R21714 CSoutput.n206 CSoutput.n202 2.25024
R21715 CSoutput.n206 CSoutput.n205 2.25024
R21716 CSoutput.n206 CSoutput.n173 2.25024
R21717 CSoutput.n256 CSoutput.n253 2.25024
R21718 CSoutput.n256 CSoutput.n252 2.25024
R21719 CSoutput.n256 CSoutput.n251 2.25024
R21720 CSoutput.n256 CSoutput.n218 2.25024
R21721 CSoutput.n256 CSoutput.n255 2.25024
R21722 CSoutput.n257 CSoutput.n256 2.25024
R21723 CSoutput.n172 CSoutput.n165 2.25024
R21724 CSoutput.n172 CSoutput.n158 2.25024
R21725 CSoutput.n284 CSoutput.n172 2.25024
R21726 CSoutput.n172 CSoutput.n168 2.25024
R21727 CSoutput.n172 CSoutput.n171 2.25024
R21728 CSoutput.n172 CSoutput.n139 2.25024
R21729 CSoutput.n273 CSoutput.n183 1.50111
R21730 CSoutput.n221 CSoutput.n207 1.50111
R21731 CSoutput.n283 CSoutput.n149 1.50111
R21732 CSoutput.n229 CSoutput.n228 1.501
R21733 CSoutput.n236 CSoutput.n235 1.501
R21734 CSoutput.n263 CSoutput.n262 1.501
R21735 CSoutput.n277 CSoutput.n188 1.12536
R21736 CSoutput.n277 CSoutput.n189 1.12536
R21737 CSoutput.n277 CSoutput.n276 1.12536
R21738 CSoutput.n237 CSoutput.n217 1.12536
R21739 CSoutput.n243 CSoutput.n217 1.12536
R21740 CSoutput.n245 CSoutput.n217 1.12536
R21741 CSoutput.n287 CSoutput.n154 1.12536
R21742 CSoutput.n287 CSoutput.n155 1.12536
R21743 CSoutput.n287 CSoutput.n286 1.12536
R21744 CSoutput.n277 CSoutput.n184 1.12536
R21745 CSoutput.n277 CSoutput.n185 1.12536
R21746 CSoutput.n277 CSoutput.n187 1.12536
R21747 CSoutput.n267 CSoutput.n217 1.12536
R21748 CSoutput.n247 CSoutput.n217 1.12536
R21749 CSoutput.n249 CSoutput.n217 1.12536
R21750 CSoutput.n287 CSoutput.n150 1.12536
R21751 CSoutput.n287 CSoutput.n151 1.12536
R21752 CSoutput.n287 CSoutput.n153 1.12536
R21753 CSoutput.n31 CSoutput.n30 0.669944
R21754 CSoutput.n62 CSoutput.n61 0.669944
R21755 CSoutput.n368 CSoutput.n366 0.573776
R21756 CSoutput.n370 CSoutput.n368 0.573776
R21757 CSoutput.n372 CSoutput.n370 0.573776
R21758 CSoutput.n374 CSoutput.n372 0.573776
R21759 CSoutput.n376 CSoutput.n374 0.573776
R21760 CSoutput.n378 CSoutput.n376 0.573776
R21761 CSoutput.n353 CSoutput.n351 0.573776
R21762 CSoutput.n355 CSoutput.n353 0.573776
R21763 CSoutput.n357 CSoutput.n355 0.573776
R21764 CSoutput.n359 CSoutput.n357 0.573776
R21765 CSoutput.n361 CSoutput.n359 0.573776
R21766 CSoutput.n363 CSoutput.n361 0.573776
R21767 CSoutput.n410 CSoutput.n408 0.573776
R21768 CSoutput.n408 CSoutput.n406 0.573776
R21769 CSoutput.n406 CSoutput.n404 0.573776
R21770 CSoutput.n404 CSoutput.n402 0.573776
R21771 CSoutput.n402 CSoutput.n400 0.573776
R21772 CSoutput.n400 CSoutput.n398 0.573776
R21773 CSoutput.n395 CSoutput.n393 0.573776
R21774 CSoutput.n393 CSoutput.n391 0.573776
R21775 CSoutput.n391 CSoutput.n389 0.573776
R21776 CSoutput.n389 CSoutput.n387 0.573776
R21777 CSoutput.n387 CSoutput.n385 0.573776
R21778 CSoutput.n385 CSoutput.n383 0.573776
R21779 CSoutput.n413 CSoutput.n288 0.53442
R21780 CSoutput.n332 CSoutput.n330 0.358259
R21781 CSoutput.n334 CSoutput.n332 0.358259
R21782 CSoutput.n336 CSoutput.n334 0.358259
R21783 CSoutput.n338 CSoutput.n336 0.358259
R21784 CSoutput.n340 CSoutput.n338 0.358259
R21785 CSoutput.n342 CSoutput.n340 0.358259
R21786 CSoutput.n344 CSoutput.n342 0.358259
R21787 CSoutput.n346 CSoutput.n344 0.358259
R21788 CSoutput.n312 CSoutput.n310 0.358259
R21789 CSoutput.n314 CSoutput.n312 0.358259
R21790 CSoutput.n316 CSoutput.n314 0.358259
R21791 CSoutput.n318 CSoutput.n316 0.358259
R21792 CSoutput.n320 CSoutput.n318 0.358259
R21793 CSoutput.n322 CSoutput.n320 0.358259
R21794 CSoutput.n324 CSoutput.n322 0.358259
R21795 CSoutput.n326 CSoutput.n324 0.358259
R21796 CSoutput.n293 CSoutput.n291 0.358259
R21797 CSoutput.n295 CSoutput.n293 0.358259
R21798 CSoutput.n297 CSoutput.n295 0.358259
R21799 CSoutput.n299 CSoutput.n297 0.358259
R21800 CSoutput.n301 CSoutput.n299 0.358259
R21801 CSoutput.n303 CSoutput.n301 0.358259
R21802 CSoutput.n305 CSoutput.n303 0.358259
R21803 CSoutput.n307 CSoutput.n305 0.358259
R21804 CSoutput.n136 CSoutput.n134 0.358259
R21805 CSoutput.n134 CSoutput.n132 0.358259
R21806 CSoutput.n132 CSoutput.n130 0.358259
R21807 CSoutput.n130 CSoutput.n128 0.358259
R21808 CSoutput.n128 CSoutput.n126 0.358259
R21809 CSoutput.n126 CSoutput.n124 0.358259
R21810 CSoutput.n124 CSoutput.n122 0.358259
R21811 CSoutput.n122 CSoutput.n120 0.358259
R21812 CSoutput.n116 CSoutput.n114 0.358259
R21813 CSoutput.n114 CSoutput.n112 0.358259
R21814 CSoutput.n112 CSoutput.n110 0.358259
R21815 CSoutput.n110 CSoutput.n108 0.358259
R21816 CSoutput.n108 CSoutput.n106 0.358259
R21817 CSoutput.n106 CSoutput.n104 0.358259
R21818 CSoutput.n104 CSoutput.n102 0.358259
R21819 CSoutput.n102 CSoutput.n100 0.358259
R21820 CSoutput.n97 CSoutput.n95 0.358259
R21821 CSoutput.n95 CSoutput.n93 0.358259
R21822 CSoutput.n93 CSoutput.n91 0.358259
R21823 CSoutput.n91 CSoutput.n89 0.358259
R21824 CSoutput.n89 CSoutput.n87 0.358259
R21825 CSoutput.n87 CSoutput.n85 0.358259
R21826 CSoutput.n85 CSoutput.n83 0.358259
R21827 CSoutput.n83 CSoutput.n81 0.358259
R21828 CSoutput.n21 CSoutput.n20 0.169105
R21829 CSoutput.n21 CSoutput.n16 0.169105
R21830 CSoutput.n26 CSoutput.n16 0.169105
R21831 CSoutput.n27 CSoutput.n26 0.169105
R21832 CSoutput.n27 CSoutput.n14 0.169105
R21833 CSoutput.n32 CSoutput.n14 0.169105
R21834 CSoutput.n33 CSoutput.n32 0.169105
R21835 CSoutput.n34 CSoutput.n33 0.169105
R21836 CSoutput.n34 CSoutput.n12 0.169105
R21837 CSoutput.n39 CSoutput.n12 0.169105
R21838 CSoutput.n40 CSoutput.n39 0.169105
R21839 CSoutput.n40 CSoutput.n10 0.169105
R21840 CSoutput.n45 CSoutput.n10 0.169105
R21841 CSoutput.n46 CSoutput.n45 0.169105
R21842 CSoutput.n47 CSoutput.n46 0.169105
R21843 CSoutput.n47 CSoutput.n8 0.169105
R21844 CSoutput.n52 CSoutput.n8 0.169105
R21845 CSoutput.n53 CSoutput.n52 0.169105
R21846 CSoutput.n53 CSoutput.n6 0.169105
R21847 CSoutput.n58 CSoutput.n6 0.169105
R21848 CSoutput.n59 CSoutput.n58 0.169105
R21849 CSoutput.n60 CSoutput.n59 0.169105
R21850 CSoutput.n60 CSoutput.n4 0.169105
R21851 CSoutput.n66 CSoutput.n4 0.169105
R21852 CSoutput.n67 CSoutput.n66 0.169105
R21853 CSoutput.n68 CSoutput.n67 0.169105
R21854 CSoutput.n68 CSoutput.n2 0.169105
R21855 CSoutput.n73 CSoutput.n2 0.169105
R21856 CSoutput.n74 CSoutput.n73 0.169105
R21857 CSoutput.n74 CSoutput.n0 0.169105
R21858 CSoutput.n78 CSoutput.n0 0.169105
R21859 CSoutput.n231 CSoutput.n230 0.0910737
R21860 CSoutput.n282 CSoutput.n279 0.0723685
R21861 CSoutput.n236 CSoutput.n231 0.0522944
R21862 CSoutput.n279 CSoutput.n278 0.0499135
R21863 CSoutput.n230 CSoutput.n229 0.0499135
R21864 CSoutput.n264 CSoutput.n263 0.0464294
R21865 CSoutput.n272 CSoutput.n269 0.0391444
R21866 CSoutput.n231 CSoutput.t202 0.023435
R21867 CSoutput.n279 CSoutput.t196 0.02262
R21868 CSoutput.n230 CSoutput.t187 0.02262
R21869 CSoutput CSoutput.n413 0.0052
R21870 CSoutput.n201 CSoutput.n184 0.00365111
R21871 CSoutput.n204 CSoutput.n185 0.00365111
R21872 CSoutput.n187 CSoutput.n186 0.00365111
R21873 CSoutput.n229 CSoutput.n188 0.00365111
R21874 CSoutput.n193 CSoutput.n189 0.00365111
R21875 CSoutput.n276 CSoutput.n190 0.00365111
R21876 CSoutput.n267 CSoutput.n266 0.00365111
R21877 CSoutput.n247 CSoutput.n220 0.00365111
R21878 CSoutput.n249 CSoutput.n219 0.00365111
R21879 CSoutput.n237 CSoutput.n236 0.00365111
R21880 CSoutput.n243 CSoutput.n223 0.00365111
R21881 CSoutput.n245 CSoutput.n222 0.00365111
R21882 CSoutput.n167 CSoutput.n150 0.00365111
R21883 CSoutput.n170 CSoutput.n151 0.00365111
R21884 CSoutput.n153 CSoutput.n152 0.00365111
R21885 CSoutput.n263 CSoutput.n154 0.00365111
R21886 CSoutput.n159 CSoutput.n155 0.00365111
R21887 CSoutput.n286 CSoutput.n156 0.00365111
R21888 CSoutput.n198 CSoutput.n188 0.00340054
R21889 CSoutput.n191 CSoutput.n189 0.00340054
R21890 CSoutput.n276 CSoutput.n275 0.00340054
R21891 CSoutput.n271 CSoutput.n184 0.00340054
R21892 CSoutput.n200 CSoutput.n185 0.00340054
R21893 CSoutput.n203 CSoutput.n187 0.00340054
R21894 CSoutput.n242 CSoutput.n237 0.00340054
R21895 CSoutput.n244 CSoutput.n243 0.00340054
R21896 CSoutput.n246 CSoutput.n245 0.00340054
R21897 CSoutput.n268 CSoutput.n267 0.00340054
R21898 CSoutput.n248 CSoutput.n247 0.00340054
R21899 CSoutput.n250 CSoutput.n249 0.00340054
R21900 CSoutput.n164 CSoutput.n154 0.00340054
R21901 CSoutput.n157 CSoutput.n155 0.00340054
R21902 CSoutput.n286 CSoutput.n285 0.00340054
R21903 CSoutput.n281 CSoutput.n150 0.00340054
R21904 CSoutput.n166 CSoutput.n151 0.00340054
R21905 CSoutput.n169 CSoutput.n153 0.00340054
R21906 CSoutput.n199 CSoutput.n193 0.00252698
R21907 CSoutput.n192 CSoutput.n190 0.00252698
R21908 CSoutput.n274 CSoutput.n273 0.00252698
R21909 CSoutput.n202 CSoutput.n200 0.00252698
R21910 CSoutput.n205 CSoutput.n203 0.00252698
R21911 CSoutput.n278 CSoutput.n173 0.00252698
R21912 CSoutput.n199 CSoutput.n198 0.00252698
R21913 CSoutput.n192 CSoutput.n191 0.00252698
R21914 CSoutput.n275 CSoutput.n274 0.00252698
R21915 CSoutput.n202 CSoutput.n201 0.00252698
R21916 CSoutput.n205 CSoutput.n204 0.00252698
R21917 CSoutput.n186 CSoutput.n173 0.00252698
R21918 CSoutput.n253 CSoutput.n223 0.00252698
R21919 CSoutput.n252 CSoutput.n222 0.00252698
R21920 CSoutput.n251 CSoutput.n207 0.00252698
R21921 CSoutput.n248 CSoutput.n218 0.00252698
R21922 CSoutput.n255 CSoutput.n250 0.00252698
R21923 CSoutput.n264 CSoutput.n257 0.00252698
R21924 CSoutput.n253 CSoutput.n242 0.00252698
R21925 CSoutput.n252 CSoutput.n244 0.00252698
R21926 CSoutput.n251 CSoutput.n246 0.00252698
R21927 CSoutput.n266 CSoutput.n218 0.00252698
R21928 CSoutput.n255 CSoutput.n220 0.00252698
R21929 CSoutput.n257 CSoutput.n219 0.00252698
R21930 CSoutput.n165 CSoutput.n159 0.00252698
R21931 CSoutput.n158 CSoutput.n156 0.00252698
R21932 CSoutput.n284 CSoutput.n283 0.00252698
R21933 CSoutput.n168 CSoutput.n166 0.00252698
R21934 CSoutput.n171 CSoutput.n169 0.00252698
R21935 CSoutput.n288 CSoutput.n139 0.00252698
R21936 CSoutput.n165 CSoutput.n164 0.00252698
R21937 CSoutput.n158 CSoutput.n157 0.00252698
R21938 CSoutput.n285 CSoutput.n284 0.00252698
R21939 CSoutput.n168 CSoutput.n167 0.00252698
R21940 CSoutput.n171 CSoutput.n170 0.00252698
R21941 CSoutput.n152 CSoutput.n139 0.00252698
R21942 CSoutput.n273 CSoutput.n272 0.0020275
R21943 CSoutput.n272 CSoutput.n271 0.0020275
R21944 CSoutput.n269 CSoutput.n207 0.0020275
R21945 CSoutput.n269 CSoutput.n268 0.0020275
R21946 CSoutput.n283 CSoutput.n282 0.0020275
R21947 CSoutput.n282 CSoutput.n281 0.0020275
R21948 CSoutput.n183 CSoutput.n182 0.00166668
R21949 CSoutput.n265 CSoutput.n221 0.00166668
R21950 CSoutput.n149 CSoutput.n148 0.00166668
R21951 CSoutput.n287 CSoutput.n149 0.00133328
R21952 CSoutput.n221 CSoutput.n217 0.00133328
R21953 CSoutput.n277 CSoutput.n183 0.00133328
R21954 CSoutput.n280 CSoutput.n172 0.001
R21955 CSoutput.n258 CSoutput.n172 0.001
R21956 CSoutput.n160 CSoutput.n140 0.001
R21957 CSoutput.n259 CSoutput.n140 0.001
R21958 CSoutput.n161 CSoutput.n141 0.001
R21959 CSoutput.n260 CSoutput.n141 0.001
R21960 CSoutput.n162 CSoutput.n142 0.001
R21961 CSoutput.n261 CSoutput.n142 0.001
R21962 CSoutput.n163 CSoutput.n143 0.001
R21963 CSoutput.n262 CSoutput.n143 0.001
R21964 CSoutput.n256 CSoutput.n208 0.001
R21965 CSoutput.n256 CSoutput.n254 0.001
R21966 CSoutput.n238 CSoutput.n209 0.001
R21967 CSoutput.n232 CSoutput.n209 0.001
R21968 CSoutput.n239 CSoutput.n210 0.001
R21969 CSoutput.n233 CSoutput.n210 0.001
R21970 CSoutput.n240 CSoutput.n211 0.001
R21971 CSoutput.n234 CSoutput.n211 0.001
R21972 CSoutput.n241 CSoutput.n212 0.001
R21973 CSoutput.n235 CSoutput.n212 0.001
R21974 CSoutput.n270 CSoutput.n206 0.001
R21975 CSoutput.n224 CSoutput.n206 0.001
R21976 CSoutput.n194 CSoutput.n174 0.001
R21977 CSoutput.n225 CSoutput.n174 0.001
R21978 CSoutput.n195 CSoutput.n175 0.001
R21979 CSoutput.n226 CSoutput.n175 0.001
R21980 CSoutput.n196 CSoutput.n176 0.001
R21981 CSoutput.n227 CSoutput.n176 0.001
R21982 CSoutput.n197 CSoutput.n177 0.001
R21983 CSoutput.n228 CSoutput.n177 0.001
R21984 CSoutput.n228 CSoutput.n178 0.001
R21985 CSoutput.n227 CSoutput.n179 0.001
R21986 CSoutput.n226 CSoutput.n180 0.001
R21987 CSoutput.n225 CSoutput.t199 0.001
R21988 CSoutput.n224 CSoutput.n181 0.001
R21989 CSoutput.n197 CSoutput.n179 0.001
R21990 CSoutput.n196 CSoutput.n180 0.001
R21991 CSoutput.n195 CSoutput.t199 0.001
R21992 CSoutput.n194 CSoutput.n181 0.001
R21993 CSoutput.n270 CSoutput.n182 0.001
R21994 CSoutput.n235 CSoutput.n213 0.001
R21995 CSoutput.n234 CSoutput.n214 0.001
R21996 CSoutput.n233 CSoutput.n215 0.001
R21997 CSoutput.n232 CSoutput.t195 0.001
R21998 CSoutput.n254 CSoutput.n216 0.001
R21999 CSoutput.n241 CSoutput.n214 0.001
R22000 CSoutput.n240 CSoutput.n215 0.001
R22001 CSoutput.n239 CSoutput.t195 0.001
R22002 CSoutput.n238 CSoutput.n216 0.001
R22003 CSoutput.n265 CSoutput.n208 0.001
R22004 CSoutput.n262 CSoutput.n144 0.001
R22005 CSoutput.n261 CSoutput.n145 0.001
R22006 CSoutput.n260 CSoutput.n146 0.001
R22007 CSoutput.n259 CSoutput.t185 0.001
R22008 CSoutput.n258 CSoutput.n147 0.001
R22009 CSoutput.n163 CSoutput.n145 0.001
R22010 CSoutput.n162 CSoutput.n146 0.001
R22011 CSoutput.n161 CSoutput.t185 0.001
R22012 CSoutput.n160 CSoutput.n147 0.001
R22013 CSoutput.n280 CSoutput.n148 0.001
R22014 a_n2408_n452.n102 a_n2408_n452.t73 512.366
R22015 a_n2408_n452.n101 a_n2408_n452.t64 512.366
R22016 a_n2408_n452.n100 a_n2408_n452.t56 512.366
R22017 a_n2408_n452.n104 a_n2408_n452.t81 512.366
R22018 a_n2408_n452.n103 a_n2408_n452.t70 512.366
R22019 a_n2408_n452.n99 a_n2408_n452.t69 512.366
R22020 a_n2408_n452.n106 a_n2408_n452.t77 512.366
R22021 a_n2408_n452.n105 a_n2408_n452.t62 512.366
R22022 a_n2408_n452.n98 a_n2408_n452.t63 512.366
R22023 a_n2408_n452.n108 a_n2408_n452.t65 512.366
R22024 a_n2408_n452.n107 a_n2408_n452.t74 512.366
R22025 a_n2408_n452.n97 a_n2408_n452.t87 512.366
R22026 a_n2408_n452.n31 a_n2408_n452.t86 533.335
R22027 a_n2408_n452.n76 a_n2408_n452.t67 512.366
R22028 a_n2408_n452.n71 a_n2408_n452.t71 512.366
R22029 a_n2408_n452.n75 a_n2408_n452.t61 512.366
R22030 a_n2408_n452.n74 a_n2408_n452.t76 512.366
R22031 a_n2408_n452.n72 a_n2408_n452.t83 512.366
R22032 a_n2408_n452.n73 a_n2408_n452.t84 512.366
R22033 a_n2408_n452.n38 a_n2408_n452.t13 533.335
R22034 a_n2408_n452.n92 a_n2408_n452.t29 512.366
R22035 a_n2408_n452.n70 a_n2408_n452.t27 512.366
R22036 a_n2408_n452.n91 a_n2408_n452.t37 512.366
R22037 a_n2408_n452.n90 a_n2408_n452.t33 512.366
R22038 a_n2408_n452.n65 a_n2408_n452.t21 512.366
R22039 a_n2408_n452.n77 a_n2408_n452.t31 512.366
R22040 a_n2408_n452.n49 a_n2408_n452.t11 533.335
R22041 a_n2408_n452.n115 a_n2408_n452.t19 512.366
R22042 a_n2408_n452.n116 a_n2408_n452.t15 512.366
R22043 a_n2408_n452.n117 a_n2408_n452.t35 512.366
R22044 a_n2408_n452.n118 a_n2408_n452.t39 512.366
R22045 a_n2408_n452.n68 a_n2408_n452.t9 512.366
R22046 a_n2408_n452.n119 a_n2408_n452.t23 512.366
R22047 a_n2408_n452.n42 a_n2408_n452.t82 533.335
R22048 a_n2408_n452.n110 a_n2408_n452.t60 512.366
R22049 a_n2408_n452.n111 a_n2408_n452.t79 512.366
R22050 a_n2408_n452.n112 a_n2408_n452.t80 512.366
R22051 a_n2408_n452.n113 a_n2408_n452.t57 512.366
R22052 a_n2408_n452.n69 a_n2408_n452.t66 512.366
R22053 a_n2408_n452.n114 a_n2408_n452.t75 512.366
R22054 a_n2408_n452.n5 a_n2408_n452.n63 70.1674
R22055 a_n2408_n452.n7 a_n2408_n452.n61 70.1674
R22056 a_n2408_n452.n9 a_n2408_n452.n59 70.1674
R22057 a_n2408_n452.n11 a_n2408_n452.n57 70.1674
R22058 a_n2408_n452.n37 a_n2408_n452.n22 70.1674
R22059 a_n2408_n452.n30 a_n2408_n452.n25 70.1674
R22060 a_n2408_n452.n77 a_n2408_n452.n30 20.9683
R22061 a_n2408_n452.n25 a_n2408_n452.n64 72.3034
R22062 a_n2408_n452.n73 a_n2408_n452.n37 20.9683
R22063 a_n2408_n452.n23 a_n2408_n452.n35 72.3034
R22064 a_n2408_n452.n35 a_n2408_n452.n72 16.6962
R22065 a_n2408_n452.n34 a_n2408_n452.n23 77.6622
R22066 a_n2408_n452.n74 a_n2408_n452.n34 5.97853
R22067 a_n2408_n452.n33 a_n2408_n452.n21 77.6622
R22068 a_n2408_n452.n21 a_n2408_n452.n32 72.3034
R22069 a_n2408_n452.n76 a_n2408_n452.n31 20.9683
R22070 a_n2408_n452.n24 a_n2408_n452.n31 70.1674
R22071 a_n2408_n452.n64 a_n2408_n452.n65 16.6962
R22072 a_n2408_n452.n41 a_n2408_n452.n25 77.6622
R22073 a_n2408_n452.n90 a_n2408_n452.n41 5.97853
R22074 a_n2408_n452.n40 a_n2408_n452.n20 77.6622
R22075 a_n2408_n452.n20 a_n2408_n452.n39 72.3034
R22076 a_n2408_n452.n92 a_n2408_n452.n38 20.9683
R22077 a_n2408_n452.n19 a_n2408_n452.n38 70.1674
R22078 a_n2408_n452.n13 a_n2408_n452.n55 70.1674
R22079 a_n2408_n452.n16 a_n2408_n452.n48 70.1674
R22080 a_n2408_n452.n114 a_n2408_n452.n48 20.9683
R22081 a_n2408_n452.n47 a_n2408_n452.n17 72.3034
R22082 a_n2408_n452.n47 a_n2408_n452.n69 16.6962
R22083 a_n2408_n452.n17 a_n2408_n452.n46 77.6622
R22084 a_n2408_n452.n113 a_n2408_n452.n46 5.97853
R22085 a_n2408_n452.n45 a_n2408_n452.n18 77.6622
R22086 a_n2408_n452.n18 a_n2408_n452.n44 72.3034
R22087 a_n2408_n452.n110 a_n2408_n452.n42 20.9683
R22088 a_n2408_n452.n43 a_n2408_n452.n42 70.1674
R22089 a_n2408_n452.n119 a_n2408_n452.n55 20.9683
R22090 a_n2408_n452.n54 a_n2408_n452.n14 72.3034
R22091 a_n2408_n452.n54 a_n2408_n452.n68 16.6962
R22092 a_n2408_n452.n14 a_n2408_n452.n53 77.6622
R22093 a_n2408_n452.n118 a_n2408_n452.n53 5.97853
R22094 a_n2408_n452.n52 a_n2408_n452.n15 77.6622
R22095 a_n2408_n452.n15 a_n2408_n452.n51 72.3034
R22096 a_n2408_n452.n115 a_n2408_n452.n49 20.9683
R22097 a_n2408_n452.n50 a_n2408_n452.n49 70.1674
R22098 a_n2408_n452.n57 a_n2408_n452.n97 20.9683
R22099 a_n2408_n452.n56 a_n2408_n452.n12 75.0448
R22100 a_n2408_n452.n107 a_n2408_n452.n56 11.2134
R22101 a_n2408_n452.n12 a_n2408_n452.n108 161.3
R22102 a_n2408_n452.n59 a_n2408_n452.n98 20.9683
R22103 a_n2408_n452.n58 a_n2408_n452.n10 75.0448
R22104 a_n2408_n452.n105 a_n2408_n452.n58 11.2134
R22105 a_n2408_n452.n10 a_n2408_n452.n106 161.3
R22106 a_n2408_n452.n61 a_n2408_n452.n99 20.9683
R22107 a_n2408_n452.n60 a_n2408_n452.n8 75.0448
R22108 a_n2408_n452.n103 a_n2408_n452.n60 11.2134
R22109 a_n2408_n452.n8 a_n2408_n452.n104 161.3
R22110 a_n2408_n452.n63 a_n2408_n452.n100 20.9683
R22111 a_n2408_n452.n62 a_n2408_n452.n6 75.0448
R22112 a_n2408_n452.n101 a_n2408_n452.n62 11.2134
R22113 a_n2408_n452.n6 a_n2408_n452.n102 161.3
R22114 a_n2408_n452.n3 a_n2408_n452.n87 81.3764
R22115 a_n2408_n452.n4 a_n2408_n452.n81 81.3764
R22116 a_n2408_n452.n0 a_n2408_n452.n78 81.3764
R22117 a_n2408_n452.n3 a_n2408_n452.n88 80.9324
R22118 a_n2408_n452.n2 a_n2408_n452.n89 80.9324
R22119 a_n2408_n452.n2 a_n2408_n452.n86 80.9324
R22120 a_n2408_n452.n2 a_n2408_n452.n85 80.9324
R22121 a_n2408_n452.n1 a_n2408_n452.n84 80.9324
R22122 a_n2408_n452.n4 a_n2408_n452.n82 80.9324
R22123 a_n2408_n452.n0 a_n2408_n452.n83 80.9324
R22124 a_n2408_n452.n0 a_n2408_n452.n80 80.9324
R22125 a_n2408_n452.n0 a_n2408_n452.n79 80.9324
R22126 a_n2408_n452.n28 a_n2408_n452.t12 74.6477
R22127 a_n2408_n452.n26 a_n2408_n452.t18 74.6477
R22128 a_n2408_n452.n27 a_n2408_n452.t14 74.2899
R22129 a_n2408_n452.n29 a_n2408_n452.t26 74.2897
R22130 a_n2408_n452.n28 a_n2408_n452.n67 70.6783
R22131 a_n2408_n452.n28 a_n2408_n452.n66 70.6783
R22132 a_n2408_n452.n26 a_n2408_n452.n93 70.6783
R22133 a_n2408_n452.n26 a_n2408_n452.n94 70.6783
R22134 a_n2408_n452.n27 a_n2408_n452.n95 70.6783
R22135 a_n2408_n452.n121 a_n2408_n452.n29 70.6782
R22136 a_n2408_n452.n102 a_n2408_n452.n101 48.2005
R22137 a_n2408_n452.t78 a_n2408_n452.n63 533.335
R22138 a_n2408_n452.n104 a_n2408_n452.n103 48.2005
R22139 a_n2408_n452.t85 a_n2408_n452.n61 533.335
R22140 a_n2408_n452.n106 a_n2408_n452.n105 48.2005
R22141 a_n2408_n452.t72 a_n2408_n452.n59 533.335
R22142 a_n2408_n452.n108 a_n2408_n452.n107 48.2005
R22143 a_n2408_n452.t68 a_n2408_n452.n57 533.335
R22144 a_n2408_n452.n75 a_n2408_n452.n74 48.2005
R22145 a_n2408_n452.n37 a_n2408_n452.t58 533.335
R22146 a_n2408_n452.n91 a_n2408_n452.n90 48.2005
R22147 a_n2408_n452.n30 a_n2408_n452.t17 533.335
R22148 a_n2408_n452.n118 a_n2408_n452.n117 48.2005
R22149 a_n2408_n452.t25 a_n2408_n452.n55 533.335
R22150 a_n2408_n452.n113 a_n2408_n452.n112 48.2005
R22151 a_n2408_n452.t59 a_n2408_n452.n48 533.335
R22152 a_n2408_n452.n32 a_n2408_n452.n71 16.6962
R22153 a_n2408_n452.n73 a_n2408_n452.n35 27.6507
R22154 a_n2408_n452.n39 a_n2408_n452.n70 16.6962
R22155 a_n2408_n452.n77 a_n2408_n452.n64 27.6507
R22156 a_n2408_n452.n116 a_n2408_n452.n51 16.6962
R22157 a_n2408_n452.n119 a_n2408_n452.n54 27.6507
R22158 a_n2408_n452.n111 a_n2408_n452.n44 16.6962
R22159 a_n2408_n452.n114 a_n2408_n452.n47 27.6507
R22160 a_n2408_n452.n33 a_n2408_n452.n71 41.7634
R22161 a_n2408_n452.n40 a_n2408_n452.n70 41.7634
R22162 a_n2408_n452.n116 a_n2408_n452.n52 41.7634
R22163 a_n2408_n452.n111 a_n2408_n452.n45 41.7634
R22164 a_n2408_n452.n1 a_n2408_n452.n0 32.6799
R22165 a_n2408_n452.n62 a_n2408_n452.n100 35.3134
R22166 a_n2408_n452.n60 a_n2408_n452.n99 35.3134
R22167 a_n2408_n452.n58 a_n2408_n452.n98 35.3134
R22168 a_n2408_n452.n56 a_n2408_n452.n97 35.3134
R22169 a_n2408_n452.n25 a_n2408_n452.n2 23.891
R22170 a_n2408_n452.n43 a_n2408_n452.n109 12.705
R22171 a_n2408_n452.n22 a_n2408_n452.n36 12.5005
R22172 a_n2408_n452.n33 a_n2408_n452.n75 5.97853
R22173 a_n2408_n452.n34 a_n2408_n452.n72 41.7634
R22174 a_n2408_n452.n40 a_n2408_n452.n91 5.97853
R22175 a_n2408_n452.n41 a_n2408_n452.n65 41.7634
R22176 a_n2408_n452.n117 a_n2408_n452.n52 5.97853
R22177 a_n2408_n452.n68 a_n2408_n452.n53 41.7634
R22178 a_n2408_n452.n112 a_n2408_n452.n45 5.97853
R22179 a_n2408_n452.n69 a_n2408_n452.n46 41.7634
R22180 a_n2408_n452.n96 a_n2408_n452.n19 11.1956
R22181 a_n2408_n452.n76 a_n2408_n452.n32 27.6507
R22182 a_n2408_n452.n92 a_n2408_n452.n39 27.6507
R22183 a_n2408_n452.n51 a_n2408_n452.n115 27.6507
R22184 a_n2408_n452.n44 a_n2408_n452.n110 27.6507
R22185 a_n2408_n452.n29 a_n2408_n452.n120 9.85898
R22186 a_n2408_n452.n109 a_n2408_n452.n12 8.73345
R22187 a_n2408_n452.n5 a_n2408_n452.n36 8.73345
R22188 a_n2408_n452.n120 a_n2408_n452.n13 7.36035
R22189 a_n2408_n452.n96 a_n2408_n452.n27 6.01559
R22190 a_n2408_n452.n120 a_n2408_n452.n36 5.3452
R22191 a_n2408_n452.n25 a_n2408_n452.n24 4.01186
R22192 a_n2408_n452.n50 a_n2408_n452.n16 4.01186
R22193 a_n2408_n452.n67 a_n2408_n452.t36 3.61217
R22194 a_n2408_n452.n67 a_n2408_n452.t40 3.61217
R22195 a_n2408_n452.n66 a_n2408_n452.t20 3.61217
R22196 a_n2408_n452.n66 a_n2408_n452.t16 3.61217
R22197 a_n2408_n452.n93 a_n2408_n452.t22 3.61217
R22198 a_n2408_n452.n93 a_n2408_n452.t32 3.61217
R22199 a_n2408_n452.n94 a_n2408_n452.t38 3.61217
R22200 a_n2408_n452.n94 a_n2408_n452.t34 3.61217
R22201 a_n2408_n452.n95 a_n2408_n452.t30 3.61217
R22202 a_n2408_n452.n95 a_n2408_n452.t28 3.61217
R22203 a_n2408_n452.t10 a_n2408_n452.n121 3.61217
R22204 a_n2408_n452.n121 a_n2408_n452.t24 3.61217
R22205 a_n2408_n452.n87 a_n2408_n452.t54 2.82907
R22206 a_n2408_n452.n87 a_n2408_n452.t1 2.82907
R22207 a_n2408_n452.n88 a_n2408_n452.t43 2.82907
R22208 a_n2408_n452.n88 a_n2408_n452.t51 2.82907
R22209 a_n2408_n452.n89 a_n2408_n452.t50 2.82907
R22210 a_n2408_n452.n89 a_n2408_n452.t5 2.82907
R22211 a_n2408_n452.n86 a_n2408_n452.t7 2.82907
R22212 a_n2408_n452.n86 a_n2408_n452.t42 2.82907
R22213 a_n2408_n452.n85 a_n2408_n452.t3 2.82907
R22214 a_n2408_n452.n85 a_n2408_n452.t48 2.82907
R22215 a_n2408_n452.n84 a_n2408_n452.t0 2.82907
R22216 a_n2408_n452.n84 a_n2408_n452.t6 2.82907
R22217 a_n2408_n452.n81 a_n2408_n452.t46 2.82907
R22218 a_n2408_n452.n81 a_n2408_n452.t8 2.82907
R22219 a_n2408_n452.n82 a_n2408_n452.t52 2.82907
R22220 a_n2408_n452.n82 a_n2408_n452.t45 2.82907
R22221 a_n2408_n452.n83 a_n2408_n452.t2 2.82907
R22222 a_n2408_n452.n83 a_n2408_n452.t53 2.82907
R22223 a_n2408_n452.n80 a_n2408_n452.t41 2.82907
R22224 a_n2408_n452.n80 a_n2408_n452.t47 2.82907
R22225 a_n2408_n452.n79 a_n2408_n452.t49 2.82907
R22226 a_n2408_n452.n79 a_n2408_n452.t4 2.82907
R22227 a_n2408_n452.n78 a_n2408_n452.t55 2.82907
R22228 a_n2408_n452.n78 a_n2408_n452.t44 2.82907
R22229 a_n2408_n452.n0 a_n2408_n452.n4 1.3324
R22230 a_n2408_n452.n109 a_n2408_n452.n96 1.30542
R22231 a_n2408_n452.n25 a_n2408_n452.n20 1.09898
R22232 a_n2408_n452.n29 a_n2408_n452.n28 1.07378
R22233 a_n2408_n452.n27 a_n2408_n452.n26 1.07378
R22234 a_n2408_n452.n9 a_n2408_n452.n8 1.04595
R22235 a_n2408_n452.n20 a_n2408_n452.n19 0.94747
R22236 a_n2408_n452.n2 a_n2408_n452.n3 0.888431
R22237 a_n2408_n452.n2 a_n2408_n452.n1 0.888431
R22238 a_n2408_n452.n23 a_n2408_n452.n21 0.758076
R22239 a_n2408_n452.n23 a_n2408_n452.n22 0.758076
R22240 a_n2408_n452.n18 a_n2408_n452.n17 0.758076
R22241 a_n2408_n452.n17 a_n2408_n452.n16 0.758076
R22242 a_n2408_n452.n15 a_n2408_n452.n14 0.758076
R22243 a_n2408_n452.n14 a_n2408_n452.n13 0.758076
R22244 a_n2408_n452.n12 a_n2408_n452.n11 0.758076
R22245 a_n2408_n452.n10 a_n2408_n452.n9 0.758076
R22246 a_n2408_n452.n8 a_n2408_n452.n7 0.758076
R22247 a_n2408_n452.n6 a_n2408_n452.n5 0.758076
R22248 a_n2408_n452.n11 a_n2408_n452.n10 0.67853
R22249 a_n2408_n452.n7 a_n2408_n452.n6 0.67853
R22250 a_n2408_n452.n50 a_n2408_n452.n15 0.568682
R22251 a_n2408_n452.n43 a_n2408_n452.n18 0.568682
R22252 a_n2408_n452.n21 a_n2408_n452.n24 0.568682
R22253 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R22254 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R22255 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R22256 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R22257 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R22258 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R22259 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R22260 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R22261 a_n2140_13878.n8 a_n2140_13878.t17 74.6477
R22262 a_n2140_13878.n13 a_n2140_13878.t18 74.2899
R22263 a_n2140_13878.n10 a_n2140_13878.t19 74.2899
R22264 a_n2140_13878.n9 a_n2140_13878.t16 74.2899
R22265 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R22266 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R22267 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R22268 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R22269 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R22270 a_n2140_13878.n15 a_n2140_13878.t6 3.61217
R22271 a_n2140_13878.n15 a_n2140_13878.t7 3.61217
R22272 a_n2140_13878.n17 a_n2140_13878.t13 3.61217
R22273 a_n2140_13878.n17 a_n2140_13878.t14 3.61217
R22274 a_n2140_13878.n19 a_n2140_13878.t0 3.61217
R22275 a_n2140_13878.n19 a_n2140_13878.t8 3.61217
R22276 a_n2140_13878.n11 a_n2140_13878.t22 3.61217
R22277 a_n2140_13878.n11 a_n2140_13878.t23 3.61217
R22278 a_n2140_13878.n7 a_n2140_13878.t20 3.61217
R22279 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R22280 a_n2140_13878.n5 a_n2140_13878.t9 3.61217
R22281 a_n2140_13878.n5 a_n2140_13878.t1 3.61217
R22282 a_n2140_13878.n3 a_n2140_13878.t12 3.61217
R22283 a_n2140_13878.n3 a_n2140_13878.t3 3.61217
R22284 a_n2140_13878.n1 a_n2140_13878.t2 3.61217
R22285 a_n2140_13878.n1 a_n2140_13878.t4 3.61217
R22286 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R22287 a_n2140_13878.n0 a_n2140_13878.t5 3.61217
R22288 a_n2140_13878.n21 a_n2140_13878.t11 3.61217
R22289 a_n2140_13878.t15 a_n2140_13878.n21 3.61217
R22290 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R22291 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R22292 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R22293 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R22294 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R22295 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R22296 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R22297 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R22298 minus.n53 minus.t28 323.478
R22299 minus.n11 minus.t8 323.478
R22300 minus.n82 minus.t13 297.12
R22301 minus.n80 minus.t15 297.12
R22302 minus.n44 minus.t5 297.12
R22303 minus.n74 minus.t6 297.12
R22304 minus.n46 minus.t26 297.12
R22305 minus.n68 minus.t21 297.12
R22306 minus.n48 minus.t23 297.12
R22307 minus.n62 minus.t16 297.12
R22308 minus.n50 minus.t17 297.12
R22309 minus.n56 minus.t9 297.12
R22310 minus.n52 minus.t27 297.12
R22311 minus.n10 minus.t7 297.12
R22312 minus.n14 minus.t11 297.12
R22313 minus.n16 minus.t10 297.12
R22314 minus.n20 minus.t12 297.12
R22315 minus.n22 minus.t20 297.12
R22316 minus.n26 minus.t18 297.12
R22317 minus.n28 minus.t25 297.12
R22318 minus.n32 minus.t24 297.12
R22319 minus.n34 minus.t14 297.12
R22320 minus.n38 minus.t22 297.12
R22321 minus.n40 minus.t19 297.12
R22322 minus.n88 minus.t2 243.255
R22323 minus.n87 minus.n85 224.169
R22324 minus.n87 minus.n86 223.454
R22325 minus.n55 minus.n54 161.3
R22326 minus.n56 minus.n51 161.3
R22327 minus.n58 minus.n57 161.3
R22328 minus.n59 minus.n50 161.3
R22329 minus.n61 minus.n60 161.3
R22330 minus.n62 minus.n49 161.3
R22331 minus.n64 minus.n63 161.3
R22332 minus.n65 minus.n48 161.3
R22333 minus.n67 minus.n66 161.3
R22334 minus.n68 minus.n47 161.3
R22335 minus.n70 minus.n69 161.3
R22336 minus.n71 minus.n46 161.3
R22337 minus.n73 minus.n72 161.3
R22338 minus.n74 minus.n45 161.3
R22339 minus.n76 minus.n75 161.3
R22340 minus.n77 minus.n44 161.3
R22341 minus.n79 minus.n78 161.3
R22342 minus.n80 minus.n43 161.3
R22343 minus.n81 minus.n42 161.3
R22344 minus.n83 minus.n82 161.3
R22345 minus.n41 minus.n40 161.3
R22346 minus.n39 minus.n0 161.3
R22347 minus.n38 minus.n37 161.3
R22348 minus.n36 minus.n1 161.3
R22349 minus.n35 minus.n34 161.3
R22350 minus.n33 minus.n2 161.3
R22351 minus.n32 minus.n31 161.3
R22352 minus.n30 minus.n3 161.3
R22353 minus.n29 minus.n28 161.3
R22354 minus.n27 minus.n4 161.3
R22355 minus.n26 minus.n25 161.3
R22356 minus.n24 minus.n5 161.3
R22357 minus.n23 minus.n22 161.3
R22358 minus.n21 minus.n6 161.3
R22359 minus.n20 minus.n19 161.3
R22360 minus.n18 minus.n7 161.3
R22361 minus.n17 minus.n16 161.3
R22362 minus.n15 minus.n8 161.3
R22363 minus.n14 minus.n13 161.3
R22364 minus.n12 minus.n9 161.3
R22365 minus.n82 minus.n81 46.0096
R22366 minus.n40 minus.n39 46.0096
R22367 minus.n12 minus.n11 45.0871
R22368 minus.n54 minus.n53 45.0871
R22369 minus.n80 minus.n79 41.6278
R22370 minus.n55 minus.n52 41.6278
R22371 minus.n10 minus.n9 41.6278
R22372 minus.n38 minus.n1 41.6278
R22373 minus.n75 minus.n44 37.246
R22374 minus.n57 minus.n56 37.246
R22375 minus.n15 minus.n14 37.246
R22376 minus.n34 minus.n33 37.246
R22377 minus.n84 minus.n83 33.3925
R22378 minus.n74 minus.n73 32.8641
R22379 minus.n61 minus.n50 32.8641
R22380 minus.n16 minus.n7 32.8641
R22381 minus.n32 minus.n3 32.8641
R22382 minus.n69 minus.n46 28.4823
R22383 minus.n63 minus.n62 28.4823
R22384 minus.n21 minus.n20 28.4823
R22385 minus.n28 minus.n27 28.4823
R22386 minus.n68 minus.n67 24.1005
R22387 minus.n67 minus.n48 24.1005
R22388 minus.n22 minus.n5 24.1005
R22389 minus.n26 minus.n5 24.1005
R22390 minus.n86 minus.t4 19.8005
R22391 minus.n86 minus.t3 19.8005
R22392 minus.n85 minus.t1 19.8005
R22393 minus.n85 minus.t0 19.8005
R22394 minus.n69 minus.n68 19.7187
R22395 minus.n63 minus.n48 19.7187
R22396 minus.n22 minus.n21 19.7187
R22397 minus.n27 minus.n26 19.7187
R22398 minus.n73 minus.n46 15.3369
R22399 minus.n62 minus.n61 15.3369
R22400 minus.n20 minus.n7 15.3369
R22401 minus.n28 minus.n3 15.3369
R22402 minus.n53 minus.n52 14.1472
R22403 minus.n11 minus.n10 14.1472
R22404 minus.n84 minus.n41 12.0933
R22405 minus minus.n89 11.7006
R22406 minus.n75 minus.n74 10.955
R22407 minus.n57 minus.n50 10.955
R22408 minus.n16 minus.n15 10.955
R22409 minus.n33 minus.n32 10.955
R22410 minus.n79 minus.n44 6.57323
R22411 minus.n56 minus.n55 6.57323
R22412 minus.n14 minus.n9 6.57323
R22413 minus.n34 minus.n1 6.57323
R22414 minus.n89 minus.n88 4.80222
R22415 minus.n81 minus.n80 2.19141
R22416 minus.n39 minus.n38 2.19141
R22417 minus.n89 minus.n84 0.972091
R22418 minus.n88 minus.n87 0.716017
R22419 minus.n83 minus.n42 0.189894
R22420 minus.n43 minus.n42 0.189894
R22421 minus.n78 minus.n43 0.189894
R22422 minus.n78 minus.n77 0.189894
R22423 minus.n77 minus.n76 0.189894
R22424 minus.n76 minus.n45 0.189894
R22425 minus.n72 minus.n45 0.189894
R22426 minus.n72 minus.n71 0.189894
R22427 minus.n71 minus.n70 0.189894
R22428 minus.n70 minus.n47 0.189894
R22429 minus.n66 minus.n47 0.189894
R22430 minus.n66 minus.n65 0.189894
R22431 minus.n65 minus.n64 0.189894
R22432 minus.n64 minus.n49 0.189894
R22433 minus.n60 minus.n49 0.189894
R22434 minus.n60 minus.n59 0.189894
R22435 minus.n59 minus.n58 0.189894
R22436 minus.n58 minus.n51 0.189894
R22437 minus.n54 minus.n51 0.189894
R22438 minus.n13 minus.n12 0.189894
R22439 minus.n13 minus.n8 0.189894
R22440 minus.n17 minus.n8 0.189894
R22441 minus.n18 minus.n17 0.189894
R22442 minus.n19 minus.n18 0.189894
R22443 minus.n19 minus.n6 0.189894
R22444 minus.n23 minus.n6 0.189894
R22445 minus.n24 minus.n23 0.189894
R22446 minus.n25 minus.n24 0.189894
R22447 minus.n25 minus.n4 0.189894
R22448 minus.n29 minus.n4 0.189894
R22449 minus.n30 minus.n29 0.189894
R22450 minus.n31 minus.n30 0.189894
R22451 minus.n31 minus.n2 0.189894
R22452 minus.n35 minus.n2 0.189894
R22453 minus.n36 minus.n35 0.189894
R22454 minus.n37 minus.n36 0.189894
R22455 minus.n37 minus.n0 0.189894
R22456 minus.n41 minus.n0 0.189894
R22457 commonsourceibias.n35 commonsourceibias.t16 223.028
R22458 commonsourceibias.n128 commonsourceibias.t85 223.028
R22459 commonsourceibias.n217 commonsourceibias.t75 223.028
R22460 commonsourceibias.n364 commonsourceibias.t54 223.028
R22461 commonsourceibias.n305 commonsourceibias.t91 223.028
R22462 commonsourceibias.n499 commonsourceibias.t78 223.028
R22463 commonsourceibias.n99 commonsourceibias.t60 207.983
R22464 commonsourceibias.n192 commonsourceibias.t92 207.983
R22465 commonsourceibias.n281 commonsourceibias.t81 207.983
R22466 commonsourceibias.n430 commonsourceibias.t8 207.983
R22467 commonsourceibias.n476 commonsourceibias.t110 207.983
R22468 commonsourceibias.n565 commonsourceibias.t97 207.983
R22469 commonsourceibias.n97 commonsourceibias.t14 168.701
R22470 commonsourceibias.n91 commonsourceibias.t38 168.701
R22471 commonsourceibias.n17 commonsourceibias.t4 168.701
R22472 commonsourceibias.n83 commonsourceibias.t28 168.701
R22473 commonsourceibias.n77 commonsourceibias.t62 168.701
R22474 commonsourceibias.n22 commonsourceibias.t18 168.701
R22475 commonsourceibias.n69 commonsourceibias.t26 168.701
R22476 commonsourceibias.n63 commonsourceibias.t6 168.701
R22477 commonsourceibias.n25 commonsourceibias.t32 168.701
R22478 commonsourceibias.n27 commonsourceibias.t42 168.701
R22479 commonsourceibias.n29 commonsourceibias.t20 168.701
R22480 commonsourceibias.n46 commonsourceibias.t30 168.701
R22481 commonsourceibias.n40 commonsourceibias.t56 168.701
R22482 commonsourceibias.n34 commonsourceibias.t12 168.701
R22483 commonsourceibias.n190 commonsourceibias.t106 168.701
R22484 commonsourceibias.n184 commonsourceibias.t119 168.701
R22485 commonsourceibias.n5 commonsourceibias.t84 168.701
R22486 commonsourceibias.n176 commonsourceibias.t100 168.701
R22487 commonsourceibias.n170 commonsourceibias.t114 168.701
R22488 commonsourceibias.n10 commonsourceibias.t80 168.701
R22489 commonsourceibias.n162 commonsourceibias.t76 168.701
R22490 commonsourceibias.n156 commonsourceibias.t105 168.701
R22491 commonsourceibias.n118 commonsourceibias.t121 168.701
R22492 commonsourceibias.n120 commonsourceibias.t71 168.701
R22493 commonsourceibias.n122 commonsourceibias.t99 168.701
R22494 commonsourceibias.n139 commonsourceibias.t95 168.701
R22495 commonsourceibias.n133 commonsourceibias.t109 168.701
R22496 commonsourceibias.n127 commonsourceibias.t89 168.701
R22497 commonsourceibias.n216 commonsourceibias.t77 168.701
R22498 commonsourceibias.n222 commonsourceibias.t96 168.701
R22499 commonsourceibias.n228 commonsourceibias.t82 168.701
R22500 commonsourceibias.n211 commonsourceibias.t86 168.701
R22501 commonsourceibias.n209 commonsourceibias.t127 168.701
R22502 commonsourceibias.n207 commonsourceibias.t108 168.701
R22503 commonsourceibias.n245 commonsourceibias.t93 168.701
R22504 commonsourceibias.n251 commonsourceibias.t67 168.701
R22505 commonsourceibias.n204 commonsourceibias.t70 168.701
R22506 commonsourceibias.n259 commonsourceibias.t101 168.701
R22507 commonsourceibias.n265 commonsourceibias.t87 168.701
R22508 commonsourceibias.n199 commonsourceibias.t74 168.701
R22509 commonsourceibias.n273 commonsourceibias.t107 168.701
R22510 commonsourceibias.n279 commonsourceibias.t94 168.701
R22511 commonsourceibias.n363 commonsourceibias.t52 168.701
R22512 commonsourceibias.n369 commonsourceibias.t2 168.701
R22513 commonsourceibias.n375 commonsourceibias.t48 168.701
R22514 commonsourceibias.n358 commonsourceibias.t40 168.701
R22515 commonsourceibias.n356 commonsourceibias.t58 168.701
R22516 commonsourceibias.n354 commonsourceibias.t50 168.701
R22517 commonsourceibias.n392 commonsourceibias.t24 168.701
R22518 commonsourceibias.n398 commonsourceibias.t44 168.701
R22519 commonsourceibias.n400 commonsourceibias.t36 168.701
R22520 commonsourceibias.n407 commonsourceibias.t10 168.701
R22521 commonsourceibias.n413 commonsourceibias.t46 168.701
R22522 commonsourceibias.n415 commonsourceibias.t22 168.701
R22523 commonsourceibias.n422 commonsourceibias.t0 168.701
R22524 commonsourceibias.n428 commonsourceibias.t34 168.701
R22525 commonsourceibias.n474 commonsourceibias.t123 168.701
R22526 commonsourceibias.n468 commonsourceibias.t68 168.701
R22527 commonsourceibias.n461 commonsourceibias.t102 168.701
R22528 commonsourceibias.n459 commonsourceibias.t117 168.701
R22529 commonsourceibias.n453 commonsourceibias.t64 168.701
R22530 commonsourceibias.n446 commonsourceibias.t72 168.701
R22531 commonsourceibias.n444 commonsourceibias.t90 168.701
R22532 commonsourceibias.n304 commonsourceibias.t83 168.701
R22533 commonsourceibias.n310 commonsourceibias.t126 168.701
R22534 commonsourceibias.n316 commonsourceibias.t113 168.701
R22535 commonsourceibias.n299 commonsourceibias.t116 168.701
R22536 commonsourceibias.n297 commonsourceibias.t66 168.701
R22537 commonsourceibias.n295 commonsourceibias.t69 168.701
R22538 commonsourceibias.n333 commonsourceibias.t122 168.701
R22539 commonsourceibias.n498 commonsourceibias.t73 168.701
R22540 commonsourceibias.n504 commonsourceibias.t115 168.701
R22541 commonsourceibias.n510 commonsourceibias.t98 168.701
R22542 commonsourceibias.n493 commonsourceibias.t103 168.701
R22543 commonsourceibias.n491 commonsourceibias.t120 168.701
R22544 commonsourceibias.n489 commonsourceibias.t125 168.701
R22545 commonsourceibias.n527 commonsourceibias.t111 168.701
R22546 commonsourceibias.n533 commonsourceibias.t79 168.701
R22547 commonsourceibias.n535 commonsourceibias.t65 168.701
R22548 commonsourceibias.n542 commonsourceibias.t118 168.701
R22549 commonsourceibias.n548 commonsourceibias.t104 168.701
R22550 commonsourceibias.n550 commonsourceibias.t88 168.701
R22551 commonsourceibias.n557 commonsourceibias.t124 168.701
R22552 commonsourceibias.n563 commonsourceibias.t112 168.701
R22553 commonsourceibias.n36 commonsourceibias.n33 161.3
R22554 commonsourceibias.n38 commonsourceibias.n37 161.3
R22555 commonsourceibias.n39 commonsourceibias.n32 161.3
R22556 commonsourceibias.n42 commonsourceibias.n41 161.3
R22557 commonsourceibias.n43 commonsourceibias.n31 161.3
R22558 commonsourceibias.n45 commonsourceibias.n44 161.3
R22559 commonsourceibias.n47 commonsourceibias.n30 161.3
R22560 commonsourceibias.n49 commonsourceibias.n48 161.3
R22561 commonsourceibias.n51 commonsourceibias.n50 161.3
R22562 commonsourceibias.n52 commonsourceibias.n28 161.3
R22563 commonsourceibias.n54 commonsourceibias.n53 161.3
R22564 commonsourceibias.n56 commonsourceibias.n55 161.3
R22565 commonsourceibias.n57 commonsourceibias.n26 161.3
R22566 commonsourceibias.n59 commonsourceibias.n58 161.3
R22567 commonsourceibias.n61 commonsourceibias.n60 161.3
R22568 commonsourceibias.n62 commonsourceibias.n24 161.3
R22569 commonsourceibias.n65 commonsourceibias.n64 161.3
R22570 commonsourceibias.n66 commonsourceibias.n23 161.3
R22571 commonsourceibias.n68 commonsourceibias.n67 161.3
R22572 commonsourceibias.n70 commonsourceibias.n21 161.3
R22573 commonsourceibias.n72 commonsourceibias.n71 161.3
R22574 commonsourceibias.n73 commonsourceibias.n20 161.3
R22575 commonsourceibias.n75 commonsourceibias.n74 161.3
R22576 commonsourceibias.n76 commonsourceibias.n19 161.3
R22577 commonsourceibias.n79 commonsourceibias.n78 161.3
R22578 commonsourceibias.n80 commonsourceibias.n18 161.3
R22579 commonsourceibias.n82 commonsourceibias.n81 161.3
R22580 commonsourceibias.n84 commonsourceibias.n16 161.3
R22581 commonsourceibias.n86 commonsourceibias.n85 161.3
R22582 commonsourceibias.n87 commonsourceibias.n15 161.3
R22583 commonsourceibias.n89 commonsourceibias.n88 161.3
R22584 commonsourceibias.n90 commonsourceibias.n14 161.3
R22585 commonsourceibias.n93 commonsourceibias.n92 161.3
R22586 commonsourceibias.n94 commonsourceibias.n13 161.3
R22587 commonsourceibias.n96 commonsourceibias.n95 161.3
R22588 commonsourceibias.n98 commonsourceibias.n12 161.3
R22589 commonsourceibias.n129 commonsourceibias.n126 161.3
R22590 commonsourceibias.n131 commonsourceibias.n130 161.3
R22591 commonsourceibias.n132 commonsourceibias.n125 161.3
R22592 commonsourceibias.n135 commonsourceibias.n134 161.3
R22593 commonsourceibias.n136 commonsourceibias.n124 161.3
R22594 commonsourceibias.n138 commonsourceibias.n137 161.3
R22595 commonsourceibias.n140 commonsourceibias.n123 161.3
R22596 commonsourceibias.n142 commonsourceibias.n141 161.3
R22597 commonsourceibias.n144 commonsourceibias.n143 161.3
R22598 commonsourceibias.n145 commonsourceibias.n121 161.3
R22599 commonsourceibias.n147 commonsourceibias.n146 161.3
R22600 commonsourceibias.n149 commonsourceibias.n148 161.3
R22601 commonsourceibias.n150 commonsourceibias.n119 161.3
R22602 commonsourceibias.n152 commonsourceibias.n151 161.3
R22603 commonsourceibias.n154 commonsourceibias.n153 161.3
R22604 commonsourceibias.n155 commonsourceibias.n117 161.3
R22605 commonsourceibias.n158 commonsourceibias.n157 161.3
R22606 commonsourceibias.n159 commonsourceibias.n11 161.3
R22607 commonsourceibias.n161 commonsourceibias.n160 161.3
R22608 commonsourceibias.n163 commonsourceibias.n9 161.3
R22609 commonsourceibias.n165 commonsourceibias.n164 161.3
R22610 commonsourceibias.n166 commonsourceibias.n8 161.3
R22611 commonsourceibias.n168 commonsourceibias.n167 161.3
R22612 commonsourceibias.n169 commonsourceibias.n7 161.3
R22613 commonsourceibias.n172 commonsourceibias.n171 161.3
R22614 commonsourceibias.n173 commonsourceibias.n6 161.3
R22615 commonsourceibias.n175 commonsourceibias.n174 161.3
R22616 commonsourceibias.n177 commonsourceibias.n4 161.3
R22617 commonsourceibias.n179 commonsourceibias.n178 161.3
R22618 commonsourceibias.n180 commonsourceibias.n3 161.3
R22619 commonsourceibias.n182 commonsourceibias.n181 161.3
R22620 commonsourceibias.n183 commonsourceibias.n2 161.3
R22621 commonsourceibias.n186 commonsourceibias.n185 161.3
R22622 commonsourceibias.n187 commonsourceibias.n1 161.3
R22623 commonsourceibias.n189 commonsourceibias.n188 161.3
R22624 commonsourceibias.n191 commonsourceibias.n0 161.3
R22625 commonsourceibias.n280 commonsourceibias.n194 161.3
R22626 commonsourceibias.n278 commonsourceibias.n277 161.3
R22627 commonsourceibias.n276 commonsourceibias.n195 161.3
R22628 commonsourceibias.n275 commonsourceibias.n274 161.3
R22629 commonsourceibias.n272 commonsourceibias.n196 161.3
R22630 commonsourceibias.n271 commonsourceibias.n270 161.3
R22631 commonsourceibias.n269 commonsourceibias.n197 161.3
R22632 commonsourceibias.n268 commonsourceibias.n267 161.3
R22633 commonsourceibias.n266 commonsourceibias.n198 161.3
R22634 commonsourceibias.n264 commonsourceibias.n263 161.3
R22635 commonsourceibias.n262 commonsourceibias.n200 161.3
R22636 commonsourceibias.n261 commonsourceibias.n260 161.3
R22637 commonsourceibias.n258 commonsourceibias.n201 161.3
R22638 commonsourceibias.n257 commonsourceibias.n256 161.3
R22639 commonsourceibias.n255 commonsourceibias.n202 161.3
R22640 commonsourceibias.n254 commonsourceibias.n253 161.3
R22641 commonsourceibias.n252 commonsourceibias.n203 161.3
R22642 commonsourceibias.n250 commonsourceibias.n249 161.3
R22643 commonsourceibias.n248 commonsourceibias.n205 161.3
R22644 commonsourceibias.n247 commonsourceibias.n246 161.3
R22645 commonsourceibias.n244 commonsourceibias.n206 161.3
R22646 commonsourceibias.n243 commonsourceibias.n242 161.3
R22647 commonsourceibias.n241 commonsourceibias.n240 161.3
R22648 commonsourceibias.n239 commonsourceibias.n208 161.3
R22649 commonsourceibias.n238 commonsourceibias.n237 161.3
R22650 commonsourceibias.n236 commonsourceibias.n235 161.3
R22651 commonsourceibias.n234 commonsourceibias.n210 161.3
R22652 commonsourceibias.n233 commonsourceibias.n232 161.3
R22653 commonsourceibias.n231 commonsourceibias.n230 161.3
R22654 commonsourceibias.n229 commonsourceibias.n212 161.3
R22655 commonsourceibias.n227 commonsourceibias.n226 161.3
R22656 commonsourceibias.n225 commonsourceibias.n213 161.3
R22657 commonsourceibias.n224 commonsourceibias.n223 161.3
R22658 commonsourceibias.n221 commonsourceibias.n214 161.3
R22659 commonsourceibias.n220 commonsourceibias.n219 161.3
R22660 commonsourceibias.n218 commonsourceibias.n215 161.3
R22661 commonsourceibias.n429 commonsourceibias.n343 161.3
R22662 commonsourceibias.n427 commonsourceibias.n426 161.3
R22663 commonsourceibias.n425 commonsourceibias.n344 161.3
R22664 commonsourceibias.n424 commonsourceibias.n423 161.3
R22665 commonsourceibias.n421 commonsourceibias.n345 161.3
R22666 commonsourceibias.n420 commonsourceibias.n419 161.3
R22667 commonsourceibias.n418 commonsourceibias.n346 161.3
R22668 commonsourceibias.n417 commonsourceibias.n416 161.3
R22669 commonsourceibias.n414 commonsourceibias.n347 161.3
R22670 commonsourceibias.n412 commonsourceibias.n411 161.3
R22671 commonsourceibias.n410 commonsourceibias.n348 161.3
R22672 commonsourceibias.n409 commonsourceibias.n408 161.3
R22673 commonsourceibias.n406 commonsourceibias.n349 161.3
R22674 commonsourceibias.n405 commonsourceibias.n404 161.3
R22675 commonsourceibias.n403 commonsourceibias.n350 161.3
R22676 commonsourceibias.n402 commonsourceibias.n401 161.3
R22677 commonsourceibias.n399 commonsourceibias.n351 161.3
R22678 commonsourceibias.n397 commonsourceibias.n396 161.3
R22679 commonsourceibias.n395 commonsourceibias.n352 161.3
R22680 commonsourceibias.n394 commonsourceibias.n393 161.3
R22681 commonsourceibias.n391 commonsourceibias.n353 161.3
R22682 commonsourceibias.n390 commonsourceibias.n389 161.3
R22683 commonsourceibias.n388 commonsourceibias.n387 161.3
R22684 commonsourceibias.n386 commonsourceibias.n355 161.3
R22685 commonsourceibias.n385 commonsourceibias.n384 161.3
R22686 commonsourceibias.n383 commonsourceibias.n382 161.3
R22687 commonsourceibias.n381 commonsourceibias.n357 161.3
R22688 commonsourceibias.n380 commonsourceibias.n379 161.3
R22689 commonsourceibias.n378 commonsourceibias.n377 161.3
R22690 commonsourceibias.n376 commonsourceibias.n359 161.3
R22691 commonsourceibias.n374 commonsourceibias.n373 161.3
R22692 commonsourceibias.n372 commonsourceibias.n360 161.3
R22693 commonsourceibias.n371 commonsourceibias.n370 161.3
R22694 commonsourceibias.n368 commonsourceibias.n361 161.3
R22695 commonsourceibias.n367 commonsourceibias.n366 161.3
R22696 commonsourceibias.n365 commonsourceibias.n362 161.3
R22697 commonsourceibias.n335 commonsourceibias.n334 161.3
R22698 commonsourceibias.n332 commonsourceibias.n294 161.3
R22699 commonsourceibias.n331 commonsourceibias.n330 161.3
R22700 commonsourceibias.n329 commonsourceibias.n328 161.3
R22701 commonsourceibias.n327 commonsourceibias.n296 161.3
R22702 commonsourceibias.n326 commonsourceibias.n325 161.3
R22703 commonsourceibias.n324 commonsourceibias.n323 161.3
R22704 commonsourceibias.n322 commonsourceibias.n298 161.3
R22705 commonsourceibias.n321 commonsourceibias.n320 161.3
R22706 commonsourceibias.n319 commonsourceibias.n318 161.3
R22707 commonsourceibias.n317 commonsourceibias.n300 161.3
R22708 commonsourceibias.n315 commonsourceibias.n314 161.3
R22709 commonsourceibias.n313 commonsourceibias.n301 161.3
R22710 commonsourceibias.n312 commonsourceibias.n311 161.3
R22711 commonsourceibias.n309 commonsourceibias.n302 161.3
R22712 commonsourceibias.n308 commonsourceibias.n307 161.3
R22713 commonsourceibias.n306 commonsourceibias.n303 161.3
R22714 commonsourceibias.n441 commonsourceibias.n293 161.3
R22715 commonsourceibias.n475 commonsourceibias.n284 161.3
R22716 commonsourceibias.n473 commonsourceibias.n472 161.3
R22717 commonsourceibias.n471 commonsourceibias.n285 161.3
R22718 commonsourceibias.n470 commonsourceibias.n469 161.3
R22719 commonsourceibias.n467 commonsourceibias.n286 161.3
R22720 commonsourceibias.n466 commonsourceibias.n465 161.3
R22721 commonsourceibias.n464 commonsourceibias.n287 161.3
R22722 commonsourceibias.n463 commonsourceibias.n462 161.3
R22723 commonsourceibias.n460 commonsourceibias.n288 161.3
R22724 commonsourceibias.n458 commonsourceibias.n457 161.3
R22725 commonsourceibias.n456 commonsourceibias.n289 161.3
R22726 commonsourceibias.n455 commonsourceibias.n454 161.3
R22727 commonsourceibias.n452 commonsourceibias.n290 161.3
R22728 commonsourceibias.n451 commonsourceibias.n450 161.3
R22729 commonsourceibias.n449 commonsourceibias.n291 161.3
R22730 commonsourceibias.n448 commonsourceibias.n447 161.3
R22731 commonsourceibias.n445 commonsourceibias.n292 161.3
R22732 commonsourceibias.n443 commonsourceibias.n442 161.3
R22733 commonsourceibias.n564 commonsourceibias.n478 161.3
R22734 commonsourceibias.n562 commonsourceibias.n561 161.3
R22735 commonsourceibias.n560 commonsourceibias.n479 161.3
R22736 commonsourceibias.n559 commonsourceibias.n558 161.3
R22737 commonsourceibias.n556 commonsourceibias.n480 161.3
R22738 commonsourceibias.n555 commonsourceibias.n554 161.3
R22739 commonsourceibias.n553 commonsourceibias.n481 161.3
R22740 commonsourceibias.n552 commonsourceibias.n551 161.3
R22741 commonsourceibias.n549 commonsourceibias.n482 161.3
R22742 commonsourceibias.n547 commonsourceibias.n546 161.3
R22743 commonsourceibias.n545 commonsourceibias.n483 161.3
R22744 commonsourceibias.n544 commonsourceibias.n543 161.3
R22745 commonsourceibias.n541 commonsourceibias.n484 161.3
R22746 commonsourceibias.n540 commonsourceibias.n539 161.3
R22747 commonsourceibias.n538 commonsourceibias.n485 161.3
R22748 commonsourceibias.n537 commonsourceibias.n536 161.3
R22749 commonsourceibias.n534 commonsourceibias.n486 161.3
R22750 commonsourceibias.n532 commonsourceibias.n531 161.3
R22751 commonsourceibias.n530 commonsourceibias.n487 161.3
R22752 commonsourceibias.n529 commonsourceibias.n528 161.3
R22753 commonsourceibias.n526 commonsourceibias.n488 161.3
R22754 commonsourceibias.n525 commonsourceibias.n524 161.3
R22755 commonsourceibias.n523 commonsourceibias.n522 161.3
R22756 commonsourceibias.n521 commonsourceibias.n490 161.3
R22757 commonsourceibias.n520 commonsourceibias.n519 161.3
R22758 commonsourceibias.n518 commonsourceibias.n517 161.3
R22759 commonsourceibias.n516 commonsourceibias.n492 161.3
R22760 commonsourceibias.n515 commonsourceibias.n514 161.3
R22761 commonsourceibias.n513 commonsourceibias.n512 161.3
R22762 commonsourceibias.n511 commonsourceibias.n494 161.3
R22763 commonsourceibias.n509 commonsourceibias.n508 161.3
R22764 commonsourceibias.n507 commonsourceibias.n495 161.3
R22765 commonsourceibias.n506 commonsourceibias.n505 161.3
R22766 commonsourceibias.n503 commonsourceibias.n496 161.3
R22767 commonsourceibias.n502 commonsourceibias.n501 161.3
R22768 commonsourceibias.n500 commonsourceibias.n497 161.3
R22769 commonsourceibias.n111 commonsourceibias.n109 81.5057
R22770 commonsourceibias.n338 commonsourceibias.n336 81.5057
R22771 commonsourceibias.n111 commonsourceibias.n110 80.9324
R22772 commonsourceibias.n113 commonsourceibias.n112 80.9324
R22773 commonsourceibias.n115 commonsourceibias.n114 80.9324
R22774 commonsourceibias.n108 commonsourceibias.n107 80.9324
R22775 commonsourceibias.n106 commonsourceibias.n105 80.9324
R22776 commonsourceibias.n104 commonsourceibias.n103 80.9324
R22777 commonsourceibias.n102 commonsourceibias.n101 80.9324
R22778 commonsourceibias.n433 commonsourceibias.n432 80.9324
R22779 commonsourceibias.n435 commonsourceibias.n434 80.9324
R22780 commonsourceibias.n437 commonsourceibias.n436 80.9324
R22781 commonsourceibias.n439 commonsourceibias.n438 80.9324
R22782 commonsourceibias.n342 commonsourceibias.n341 80.9324
R22783 commonsourceibias.n340 commonsourceibias.n339 80.9324
R22784 commonsourceibias.n338 commonsourceibias.n337 80.9324
R22785 commonsourceibias.n100 commonsourceibias.n99 80.6037
R22786 commonsourceibias.n193 commonsourceibias.n192 80.6037
R22787 commonsourceibias.n282 commonsourceibias.n281 80.6037
R22788 commonsourceibias.n431 commonsourceibias.n430 80.6037
R22789 commonsourceibias.n477 commonsourceibias.n476 80.6037
R22790 commonsourceibias.n566 commonsourceibias.n565 80.6037
R22791 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22792 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22793 commonsourceibias.n62 commonsourceibias.n61 56.5617
R22794 commonsourceibias.n48 commonsourceibias.n47 56.5617
R22795 commonsourceibias.n178 commonsourceibias.n177 56.5617
R22796 commonsourceibias.n164 commonsourceibias.n163 56.5617
R22797 commonsourceibias.n155 commonsourceibias.n154 56.5617
R22798 commonsourceibias.n141 commonsourceibias.n140 56.5617
R22799 commonsourceibias.n230 commonsourceibias.n229 56.5617
R22800 commonsourceibias.n244 commonsourceibias.n243 56.5617
R22801 commonsourceibias.n253 commonsourceibias.n252 56.5617
R22802 commonsourceibias.n267 commonsourceibias.n266 56.5617
R22803 commonsourceibias.n377 commonsourceibias.n376 56.5617
R22804 commonsourceibias.n391 commonsourceibias.n390 56.5617
R22805 commonsourceibias.n401 commonsourceibias.n399 56.5617
R22806 commonsourceibias.n416 commonsourceibias.n414 56.5617
R22807 commonsourceibias.n462 commonsourceibias.n460 56.5617
R22808 commonsourceibias.n447 commonsourceibias.n445 56.5617
R22809 commonsourceibias.n318 commonsourceibias.n317 56.5617
R22810 commonsourceibias.n332 commonsourceibias.n331 56.5617
R22811 commonsourceibias.n512 commonsourceibias.n511 56.5617
R22812 commonsourceibias.n526 commonsourceibias.n525 56.5617
R22813 commonsourceibias.n536 commonsourceibias.n534 56.5617
R22814 commonsourceibias.n551 commonsourceibias.n549 56.5617
R22815 commonsourceibias.n76 commonsourceibias.n75 56.0773
R22816 commonsourceibias.n57 commonsourceibias.n56 56.0773
R22817 commonsourceibias.n169 commonsourceibias.n168 56.0773
R22818 commonsourceibias.n150 commonsourceibias.n149 56.0773
R22819 commonsourceibias.n239 commonsourceibias.n238 56.0773
R22820 commonsourceibias.n258 commonsourceibias.n257 56.0773
R22821 commonsourceibias.n386 commonsourceibias.n385 56.0773
R22822 commonsourceibias.n406 commonsourceibias.n405 56.0773
R22823 commonsourceibias.n452 commonsourceibias.n451 56.0773
R22824 commonsourceibias.n327 commonsourceibias.n326 56.0773
R22825 commonsourceibias.n521 commonsourceibias.n520 56.0773
R22826 commonsourceibias.n541 commonsourceibias.n540 56.0773
R22827 commonsourceibias.n99 commonsourceibias.n98 55.3321
R22828 commonsourceibias.n192 commonsourceibias.n191 55.3321
R22829 commonsourceibias.n281 commonsourceibias.n280 55.3321
R22830 commonsourceibias.n430 commonsourceibias.n429 55.3321
R22831 commonsourceibias.n476 commonsourceibias.n475 55.3321
R22832 commonsourceibias.n565 commonsourceibias.n564 55.3321
R22833 commonsourceibias.n90 commonsourceibias.n89 55.1086
R22834 commonsourceibias.n41 commonsourceibias.n31 55.1086
R22835 commonsourceibias.n183 commonsourceibias.n182 55.1086
R22836 commonsourceibias.n134 commonsourceibias.n124 55.1086
R22837 commonsourceibias.n223 commonsourceibias.n213 55.1086
R22838 commonsourceibias.n272 commonsourceibias.n271 55.1086
R22839 commonsourceibias.n370 commonsourceibias.n360 55.1086
R22840 commonsourceibias.n421 commonsourceibias.n420 55.1086
R22841 commonsourceibias.n467 commonsourceibias.n466 55.1086
R22842 commonsourceibias.n311 commonsourceibias.n301 55.1086
R22843 commonsourceibias.n505 commonsourceibias.n495 55.1086
R22844 commonsourceibias.n556 commonsourceibias.n555 55.1086
R22845 commonsourceibias.n35 commonsourceibias.n34 47.4592
R22846 commonsourceibias.n128 commonsourceibias.n127 47.4592
R22847 commonsourceibias.n217 commonsourceibias.n216 47.4592
R22848 commonsourceibias.n364 commonsourceibias.n363 47.4592
R22849 commonsourceibias.n305 commonsourceibias.n304 47.4592
R22850 commonsourceibias.n499 commonsourceibias.n498 47.4592
R22851 commonsourceibias.n218 commonsourceibias.n217 44.0436
R22852 commonsourceibias.n365 commonsourceibias.n364 44.0436
R22853 commonsourceibias.n306 commonsourceibias.n305 44.0436
R22854 commonsourceibias.n500 commonsourceibias.n499 44.0436
R22855 commonsourceibias.n36 commonsourceibias.n35 44.0436
R22856 commonsourceibias.n129 commonsourceibias.n128 44.0436
R22857 commonsourceibias.n92 commonsourceibias.n13 42.5146
R22858 commonsourceibias.n39 commonsourceibias.n38 42.5146
R22859 commonsourceibias.n185 commonsourceibias.n1 42.5146
R22860 commonsourceibias.n132 commonsourceibias.n131 42.5146
R22861 commonsourceibias.n221 commonsourceibias.n220 42.5146
R22862 commonsourceibias.n274 commonsourceibias.n195 42.5146
R22863 commonsourceibias.n368 commonsourceibias.n367 42.5146
R22864 commonsourceibias.n423 commonsourceibias.n344 42.5146
R22865 commonsourceibias.n469 commonsourceibias.n285 42.5146
R22866 commonsourceibias.n309 commonsourceibias.n308 42.5146
R22867 commonsourceibias.n503 commonsourceibias.n502 42.5146
R22868 commonsourceibias.n558 commonsourceibias.n479 42.5146
R22869 commonsourceibias.n78 commonsourceibias.n18 41.5458
R22870 commonsourceibias.n53 commonsourceibias.n52 41.5458
R22871 commonsourceibias.n171 commonsourceibias.n6 41.5458
R22872 commonsourceibias.n146 commonsourceibias.n145 41.5458
R22873 commonsourceibias.n235 commonsourceibias.n234 41.5458
R22874 commonsourceibias.n260 commonsourceibias.n200 41.5458
R22875 commonsourceibias.n382 commonsourceibias.n381 41.5458
R22876 commonsourceibias.n408 commonsourceibias.n348 41.5458
R22877 commonsourceibias.n454 commonsourceibias.n289 41.5458
R22878 commonsourceibias.n323 commonsourceibias.n322 41.5458
R22879 commonsourceibias.n517 commonsourceibias.n516 41.5458
R22880 commonsourceibias.n543 commonsourceibias.n483 41.5458
R22881 commonsourceibias.n68 commonsourceibias.n23 40.577
R22882 commonsourceibias.n64 commonsourceibias.n23 40.577
R22883 commonsourceibias.n161 commonsourceibias.n11 40.577
R22884 commonsourceibias.n157 commonsourceibias.n11 40.577
R22885 commonsourceibias.n246 commonsourceibias.n205 40.577
R22886 commonsourceibias.n250 commonsourceibias.n205 40.577
R22887 commonsourceibias.n393 commonsourceibias.n352 40.577
R22888 commonsourceibias.n397 commonsourceibias.n352 40.577
R22889 commonsourceibias.n443 commonsourceibias.n293 40.577
R22890 commonsourceibias.n334 commonsourceibias.n293 40.577
R22891 commonsourceibias.n528 commonsourceibias.n487 40.577
R22892 commonsourceibias.n532 commonsourceibias.n487 40.577
R22893 commonsourceibias.n82 commonsourceibias.n18 39.6083
R22894 commonsourceibias.n52 commonsourceibias.n51 39.6083
R22895 commonsourceibias.n175 commonsourceibias.n6 39.6083
R22896 commonsourceibias.n145 commonsourceibias.n144 39.6083
R22897 commonsourceibias.n234 commonsourceibias.n233 39.6083
R22898 commonsourceibias.n264 commonsourceibias.n200 39.6083
R22899 commonsourceibias.n381 commonsourceibias.n380 39.6083
R22900 commonsourceibias.n412 commonsourceibias.n348 39.6083
R22901 commonsourceibias.n458 commonsourceibias.n289 39.6083
R22902 commonsourceibias.n322 commonsourceibias.n321 39.6083
R22903 commonsourceibias.n516 commonsourceibias.n515 39.6083
R22904 commonsourceibias.n547 commonsourceibias.n483 39.6083
R22905 commonsourceibias.n96 commonsourceibias.n13 38.6395
R22906 commonsourceibias.n38 commonsourceibias.n33 38.6395
R22907 commonsourceibias.n189 commonsourceibias.n1 38.6395
R22908 commonsourceibias.n131 commonsourceibias.n126 38.6395
R22909 commonsourceibias.n220 commonsourceibias.n215 38.6395
R22910 commonsourceibias.n278 commonsourceibias.n195 38.6395
R22911 commonsourceibias.n367 commonsourceibias.n362 38.6395
R22912 commonsourceibias.n427 commonsourceibias.n344 38.6395
R22913 commonsourceibias.n473 commonsourceibias.n285 38.6395
R22914 commonsourceibias.n308 commonsourceibias.n303 38.6395
R22915 commonsourceibias.n502 commonsourceibias.n497 38.6395
R22916 commonsourceibias.n562 commonsourceibias.n479 38.6395
R22917 commonsourceibias.n89 commonsourceibias.n15 26.0455
R22918 commonsourceibias.n45 commonsourceibias.n31 26.0455
R22919 commonsourceibias.n182 commonsourceibias.n3 26.0455
R22920 commonsourceibias.n138 commonsourceibias.n124 26.0455
R22921 commonsourceibias.n227 commonsourceibias.n213 26.0455
R22922 commonsourceibias.n271 commonsourceibias.n197 26.0455
R22923 commonsourceibias.n374 commonsourceibias.n360 26.0455
R22924 commonsourceibias.n420 commonsourceibias.n346 26.0455
R22925 commonsourceibias.n466 commonsourceibias.n287 26.0455
R22926 commonsourceibias.n315 commonsourceibias.n301 26.0455
R22927 commonsourceibias.n509 commonsourceibias.n495 26.0455
R22928 commonsourceibias.n555 commonsourceibias.n481 26.0455
R22929 commonsourceibias.n75 commonsourceibias.n20 25.0767
R22930 commonsourceibias.n58 commonsourceibias.n57 25.0767
R22931 commonsourceibias.n168 commonsourceibias.n8 25.0767
R22932 commonsourceibias.n151 commonsourceibias.n150 25.0767
R22933 commonsourceibias.n240 commonsourceibias.n239 25.0767
R22934 commonsourceibias.n257 commonsourceibias.n202 25.0767
R22935 commonsourceibias.n387 commonsourceibias.n386 25.0767
R22936 commonsourceibias.n405 commonsourceibias.n350 25.0767
R22937 commonsourceibias.n451 commonsourceibias.n291 25.0767
R22938 commonsourceibias.n328 commonsourceibias.n327 25.0767
R22939 commonsourceibias.n522 commonsourceibias.n521 25.0767
R22940 commonsourceibias.n540 commonsourceibias.n485 25.0767
R22941 commonsourceibias.n71 commonsourceibias.n22 24.3464
R22942 commonsourceibias.n61 commonsourceibias.n25 24.3464
R22943 commonsourceibias.n164 commonsourceibias.n10 24.3464
R22944 commonsourceibias.n154 commonsourceibias.n118 24.3464
R22945 commonsourceibias.n243 commonsourceibias.n207 24.3464
R22946 commonsourceibias.n253 commonsourceibias.n204 24.3464
R22947 commonsourceibias.n390 commonsourceibias.n354 24.3464
R22948 commonsourceibias.n401 commonsourceibias.n400 24.3464
R22949 commonsourceibias.n447 commonsourceibias.n446 24.3464
R22950 commonsourceibias.n331 commonsourceibias.n295 24.3464
R22951 commonsourceibias.n525 commonsourceibias.n489 24.3464
R22952 commonsourceibias.n536 commonsourceibias.n535 24.3464
R22953 commonsourceibias.n85 commonsourceibias.n17 23.8546
R22954 commonsourceibias.n47 commonsourceibias.n46 23.8546
R22955 commonsourceibias.n178 commonsourceibias.n5 23.8546
R22956 commonsourceibias.n140 commonsourceibias.n139 23.8546
R22957 commonsourceibias.n229 commonsourceibias.n228 23.8546
R22958 commonsourceibias.n267 commonsourceibias.n199 23.8546
R22959 commonsourceibias.n376 commonsourceibias.n375 23.8546
R22960 commonsourceibias.n416 commonsourceibias.n415 23.8546
R22961 commonsourceibias.n462 commonsourceibias.n461 23.8546
R22962 commonsourceibias.n317 commonsourceibias.n316 23.8546
R22963 commonsourceibias.n511 commonsourceibias.n510 23.8546
R22964 commonsourceibias.n551 commonsourceibias.n550 23.8546
R22965 commonsourceibias.n98 commonsourceibias.n97 17.4607
R22966 commonsourceibias.n191 commonsourceibias.n190 17.4607
R22967 commonsourceibias.n280 commonsourceibias.n279 17.4607
R22968 commonsourceibias.n429 commonsourceibias.n428 17.4607
R22969 commonsourceibias.n475 commonsourceibias.n474 17.4607
R22970 commonsourceibias.n564 commonsourceibias.n563 17.4607
R22971 commonsourceibias.n84 commonsourceibias.n83 16.9689
R22972 commonsourceibias.n48 commonsourceibias.n29 16.9689
R22973 commonsourceibias.n177 commonsourceibias.n176 16.9689
R22974 commonsourceibias.n141 commonsourceibias.n122 16.9689
R22975 commonsourceibias.n230 commonsourceibias.n211 16.9689
R22976 commonsourceibias.n266 commonsourceibias.n265 16.9689
R22977 commonsourceibias.n377 commonsourceibias.n358 16.9689
R22978 commonsourceibias.n414 commonsourceibias.n413 16.9689
R22979 commonsourceibias.n460 commonsourceibias.n459 16.9689
R22980 commonsourceibias.n318 commonsourceibias.n299 16.9689
R22981 commonsourceibias.n512 commonsourceibias.n493 16.9689
R22982 commonsourceibias.n549 commonsourceibias.n548 16.9689
R22983 commonsourceibias.n70 commonsourceibias.n69 16.477
R22984 commonsourceibias.n63 commonsourceibias.n62 16.477
R22985 commonsourceibias.n163 commonsourceibias.n162 16.477
R22986 commonsourceibias.n156 commonsourceibias.n155 16.477
R22987 commonsourceibias.n245 commonsourceibias.n244 16.477
R22988 commonsourceibias.n252 commonsourceibias.n251 16.477
R22989 commonsourceibias.n392 commonsourceibias.n391 16.477
R22990 commonsourceibias.n399 commonsourceibias.n398 16.477
R22991 commonsourceibias.n445 commonsourceibias.n444 16.477
R22992 commonsourceibias.n333 commonsourceibias.n332 16.477
R22993 commonsourceibias.n527 commonsourceibias.n526 16.477
R22994 commonsourceibias.n534 commonsourceibias.n533 16.477
R22995 commonsourceibias.n77 commonsourceibias.n76 15.9852
R22996 commonsourceibias.n56 commonsourceibias.n27 15.9852
R22997 commonsourceibias.n170 commonsourceibias.n169 15.9852
R22998 commonsourceibias.n149 commonsourceibias.n120 15.9852
R22999 commonsourceibias.n238 commonsourceibias.n209 15.9852
R23000 commonsourceibias.n259 commonsourceibias.n258 15.9852
R23001 commonsourceibias.n385 commonsourceibias.n356 15.9852
R23002 commonsourceibias.n407 commonsourceibias.n406 15.9852
R23003 commonsourceibias.n453 commonsourceibias.n452 15.9852
R23004 commonsourceibias.n326 commonsourceibias.n297 15.9852
R23005 commonsourceibias.n520 commonsourceibias.n491 15.9852
R23006 commonsourceibias.n542 commonsourceibias.n541 15.9852
R23007 commonsourceibias.n91 commonsourceibias.n90 15.4934
R23008 commonsourceibias.n41 commonsourceibias.n40 15.4934
R23009 commonsourceibias.n184 commonsourceibias.n183 15.4934
R23010 commonsourceibias.n134 commonsourceibias.n133 15.4934
R23011 commonsourceibias.n223 commonsourceibias.n222 15.4934
R23012 commonsourceibias.n273 commonsourceibias.n272 15.4934
R23013 commonsourceibias.n370 commonsourceibias.n369 15.4934
R23014 commonsourceibias.n422 commonsourceibias.n421 15.4934
R23015 commonsourceibias.n468 commonsourceibias.n467 15.4934
R23016 commonsourceibias.n311 commonsourceibias.n310 15.4934
R23017 commonsourceibias.n505 commonsourceibias.n504 15.4934
R23018 commonsourceibias.n557 commonsourceibias.n556 15.4934
R23019 commonsourceibias.n102 commonsourceibias.n100 13.2663
R23020 commonsourceibias.n433 commonsourceibias.n431 13.2663
R23021 commonsourceibias.n568 commonsourceibias.n283 12.2777
R23022 commonsourceibias.n568 commonsourceibias.n567 10.3347
R23023 commonsourceibias.n159 commonsourceibias.n116 9.50363
R23024 commonsourceibias.n441 commonsourceibias.n440 9.50363
R23025 commonsourceibias.n92 commonsourceibias.n91 9.09948
R23026 commonsourceibias.n40 commonsourceibias.n39 9.09948
R23027 commonsourceibias.n185 commonsourceibias.n184 9.09948
R23028 commonsourceibias.n133 commonsourceibias.n132 9.09948
R23029 commonsourceibias.n222 commonsourceibias.n221 9.09948
R23030 commonsourceibias.n274 commonsourceibias.n273 9.09948
R23031 commonsourceibias.n369 commonsourceibias.n368 9.09948
R23032 commonsourceibias.n423 commonsourceibias.n422 9.09948
R23033 commonsourceibias.n469 commonsourceibias.n468 9.09948
R23034 commonsourceibias.n310 commonsourceibias.n309 9.09948
R23035 commonsourceibias.n504 commonsourceibias.n503 9.09948
R23036 commonsourceibias.n558 commonsourceibias.n557 9.09948
R23037 commonsourceibias.n283 commonsourceibias.n193 8.79261
R23038 commonsourceibias.n567 commonsourceibias.n477 8.79261
R23039 commonsourceibias.n78 commonsourceibias.n77 8.60764
R23040 commonsourceibias.n53 commonsourceibias.n27 8.60764
R23041 commonsourceibias.n171 commonsourceibias.n170 8.60764
R23042 commonsourceibias.n146 commonsourceibias.n120 8.60764
R23043 commonsourceibias.n235 commonsourceibias.n209 8.60764
R23044 commonsourceibias.n260 commonsourceibias.n259 8.60764
R23045 commonsourceibias.n382 commonsourceibias.n356 8.60764
R23046 commonsourceibias.n408 commonsourceibias.n407 8.60764
R23047 commonsourceibias.n454 commonsourceibias.n453 8.60764
R23048 commonsourceibias.n323 commonsourceibias.n297 8.60764
R23049 commonsourceibias.n517 commonsourceibias.n491 8.60764
R23050 commonsourceibias.n543 commonsourceibias.n542 8.60764
R23051 commonsourceibias.n69 commonsourceibias.n68 8.11581
R23052 commonsourceibias.n64 commonsourceibias.n63 8.11581
R23053 commonsourceibias.n162 commonsourceibias.n161 8.11581
R23054 commonsourceibias.n157 commonsourceibias.n156 8.11581
R23055 commonsourceibias.n246 commonsourceibias.n245 8.11581
R23056 commonsourceibias.n251 commonsourceibias.n250 8.11581
R23057 commonsourceibias.n393 commonsourceibias.n392 8.11581
R23058 commonsourceibias.n398 commonsourceibias.n397 8.11581
R23059 commonsourceibias.n444 commonsourceibias.n443 8.11581
R23060 commonsourceibias.n334 commonsourceibias.n333 8.11581
R23061 commonsourceibias.n528 commonsourceibias.n527 8.11581
R23062 commonsourceibias.n533 commonsourceibias.n532 8.11581
R23063 commonsourceibias.n83 commonsourceibias.n82 7.62397
R23064 commonsourceibias.n51 commonsourceibias.n29 7.62397
R23065 commonsourceibias.n176 commonsourceibias.n175 7.62397
R23066 commonsourceibias.n144 commonsourceibias.n122 7.62397
R23067 commonsourceibias.n233 commonsourceibias.n211 7.62397
R23068 commonsourceibias.n265 commonsourceibias.n264 7.62397
R23069 commonsourceibias.n380 commonsourceibias.n358 7.62397
R23070 commonsourceibias.n413 commonsourceibias.n412 7.62397
R23071 commonsourceibias.n459 commonsourceibias.n458 7.62397
R23072 commonsourceibias.n321 commonsourceibias.n299 7.62397
R23073 commonsourceibias.n515 commonsourceibias.n493 7.62397
R23074 commonsourceibias.n548 commonsourceibias.n547 7.62397
R23075 commonsourceibias.n97 commonsourceibias.n96 7.13213
R23076 commonsourceibias.n34 commonsourceibias.n33 7.13213
R23077 commonsourceibias.n190 commonsourceibias.n189 7.13213
R23078 commonsourceibias.n127 commonsourceibias.n126 7.13213
R23079 commonsourceibias.n216 commonsourceibias.n215 7.13213
R23080 commonsourceibias.n279 commonsourceibias.n278 7.13213
R23081 commonsourceibias.n363 commonsourceibias.n362 7.13213
R23082 commonsourceibias.n428 commonsourceibias.n427 7.13213
R23083 commonsourceibias.n474 commonsourceibias.n473 7.13213
R23084 commonsourceibias.n304 commonsourceibias.n303 7.13213
R23085 commonsourceibias.n498 commonsourceibias.n497 7.13213
R23086 commonsourceibias.n563 commonsourceibias.n562 7.13213
R23087 commonsourceibias.n283 commonsourceibias.n282 5.06534
R23088 commonsourceibias.n567 commonsourceibias.n566 5.06534
R23089 commonsourceibias commonsourceibias.n568 4.04308
R23090 commonsourceibias.n109 commonsourceibias.t13 2.82907
R23091 commonsourceibias.n109 commonsourceibias.t17 2.82907
R23092 commonsourceibias.n110 commonsourceibias.t31 2.82907
R23093 commonsourceibias.n110 commonsourceibias.t57 2.82907
R23094 commonsourceibias.n112 commonsourceibias.t43 2.82907
R23095 commonsourceibias.n112 commonsourceibias.t21 2.82907
R23096 commonsourceibias.n114 commonsourceibias.t7 2.82907
R23097 commonsourceibias.n114 commonsourceibias.t33 2.82907
R23098 commonsourceibias.n107 commonsourceibias.t19 2.82907
R23099 commonsourceibias.n107 commonsourceibias.t27 2.82907
R23100 commonsourceibias.n105 commonsourceibias.t29 2.82907
R23101 commonsourceibias.n105 commonsourceibias.t63 2.82907
R23102 commonsourceibias.n103 commonsourceibias.t39 2.82907
R23103 commonsourceibias.n103 commonsourceibias.t5 2.82907
R23104 commonsourceibias.n101 commonsourceibias.t61 2.82907
R23105 commonsourceibias.n101 commonsourceibias.t15 2.82907
R23106 commonsourceibias.n432 commonsourceibias.t35 2.82907
R23107 commonsourceibias.n432 commonsourceibias.t9 2.82907
R23108 commonsourceibias.n434 commonsourceibias.t23 2.82907
R23109 commonsourceibias.n434 commonsourceibias.t1 2.82907
R23110 commonsourceibias.n436 commonsourceibias.t11 2.82907
R23111 commonsourceibias.n436 commonsourceibias.t47 2.82907
R23112 commonsourceibias.n438 commonsourceibias.t45 2.82907
R23113 commonsourceibias.n438 commonsourceibias.t37 2.82907
R23114 commonsourceibias.n341 commonsourceibias.t51 2.82907
R23115 commonsourceibias.n341 commonsourceibias.t25 2.82907
R23116 commonsourceibias.n339 commonsourceibias.t41 2.82907
R23117 commonsourceibias.n339 commonsourceibias.t59 2.82907
R23118 commonsourceibias.n337 commonsourceibias.t3 2.82907
R23119 commonsourceibias.n337 commonsourceibias.t49 2.82907
R23120 commonsourceibias.n336 commonsourceibias.t55 2.82907
R23121 commonsourceibias.n336 commonsourceibias.t53 2.82907
R23122 commonsourceibias.n17 commonsourceibias.n15 0.738255
R23123 commonsourceibias.n46 commonsourceibias.n45 0.738255
R23124 commonsourceibias.n5 commonsourceibias.n3 0.738255
R23125 commonsourceibias.n139 commonsourceibias.n138 0.738255
R23126 commonsourceibias.n228 commonsourceibias.n227 0.738255
R23127 commonsourceibias.n199 commonsourceibias.n197 0.738255
R23128 commonsourceibias.n375 commonsourceibias.n374 0.738255
R23129 commonsourceibias.n415 commonsourceibias.n346 0.738255
R23130 commonsourceibias.n461 commonsourceibias.n287 0.738255
R23131 commonsourceibias.n316 commonsourceibias.n315 0.738255
R23132 commonsourceibias.n510 commonsourceibias.n509 0.738255
R23133 commonsourceibias.n550 commonsourceibias.n481 0.738255
R23134 commonsourceibias.n104 commonsourceibias.n102 0.573776
R23135 commonsourceibias.n106 commonsourceibias.n104 0.573776
R23136 commonsourceibias.n108 commonsourceibias.n106 0.573776
R23137 commonsourceibias.n115 commonsourceibias.n113 0.573776
R23138 commonsourceibias.n113 commonsourceibias.n111 0.573776
R23139 commonsourceibias.n340 commonsourceibias.n338 0.573776
R23140 commonsourceibias.n342 commonsourceibias.n340 0.573776
R23141 commonsourceibias.n439 commonsourceibias.n437 0.573776
R23142 commonsourceibias.n437 commonsourceibias.n435 0.573776
R23143 commonsourceibias.n435 commonsourceibias.n433 0.573776
R23144 commonsourceibias.n116 commonsourceibias.n108 0.287138
R23145 commonsourceibias.n116 commonsourceibias.n115 0.287138
R23146 commonsourceibias.n440 commonsourceibias.n342 0.287138
R23147 commonsourceibias.n440 commonsourceibias.n439 0.287138
R23148 commonsourceibias.n100 commonsourceibias.n12 0.285035
R23149 commonsourceibias.n193 commonsourceibias.n0 0.285035
R23150 commonsourceibias.n282 commonsourceibias.n194 0.285035
R23151 commonsourceibias.n431 commonsourceibias.n343 0.285035
R23152 commonsourceibias.n477 commonsourceibias.n284 0.285035
R23153 commonsourceibias.n566 commonsourceibias.n478 0.285035
R23154 commonsourceibias.n22 commonsourceibias.n20 0.246418
R23155 commonsourceibias.n58 commonsourceibias.n25 0.246418
R23156 commonsourceibias.n10 commonsourceibias.n8 0.246418
R23157 commonsourceibias.n151 commonsourceibias.n118 0.246418
R23158 commonsourceibias.n240 commonsourceibias.n207 0.246418
R23159 commonsourceibias.n204 commonsourceibias.n202 0.246418
R23160 commonsourceibias.n387 commonsourceibias.n354 0.246418
R23161 commonsourceibias.n400 commonsourceibias.n350 0.246418
R23162 commonsourceibias.n446 commonsourceibias.n291 0.246418
R23163 commonsourceibias.n328 commonsourceibias.n295 0.246418
R23164 commonsourceibias.n522 commonsourceibias.n489 0.246418
R23165 commonsourceibias.n535 commonsourceibias.n485 0.246418
R23166 commonsourceibias.n95 commonsourceibias.n12 0.189894
R23167 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23168 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23169 commonsourceibias.n93 commonsourceibias.n14 0.189894
R23170 commonsourceibias.n88 commonsourceibias.n14 0.189894
R23171 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23172 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23173 commonsourceibias.n86 commonsourceibias.n16 0.189894
R23174 commonsourceibias.n81 commonsourceibias.n16 0.189894
R23175 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23176 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23177 commonsourceibias.n79 commonsourceibias.n19 0.189894
R23178 commonsourceibias.n74 commonsourceibias.n19 0.189894
R23179 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23180 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23181 commonsourceibias.n72 commonsourceibias.n21 0.189894
R23182 commonsourceibias.n67 commonsourceibias.n21 0.189894
R23183 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23184 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23185 commonsourceibias.n65 commonsourceibias.n24 0.189894
R23186 commonsourceibias.n60 commonsourceibias.n24 0.189894
R23187 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23188 commonsourceibias.n59 commonsourceibias.n26 0.189894
R23189 commonsourceibias.n55 commonsourceibias.n26 0.189894
R23190 commonsourceibias.n55 commonsourceibias.n54 0.189894
R23191 commonsourceibias.n54 commonsourceibias.n28 0.189894
R23192 commonsourceibias.n50 commonsourceibias.n28 0.189894
R23193 commonsourceibias.n50 commonsourceibias.n49 0.189894
R23194 commonsourceibias.n49 commonsourceibias.n30 0.189894
R23195 commonsourceibias.n44 commonsourceibias.n30 0.189894
R23196 commonsourceibias.n44 commonsourceibias.n43 0.189894
R23197 commonsourceibias.n43 commonsourceibias.n42 0.189894
R23198 commonsourceibias.n42 commonsourceibias.n32 0.189894
R23199 commonsourceibias.n37 commonsourceibias.n32 0.189894
R23200 commonsourceibias.n37 commonsourceibias.n36 0.189894
R23201 commonsourceibias.n158 commonsourceibias.n117 0.189894
R23202 commonsourceibias.n153 commonsourceibias.n117 0.189894
R23203 commonsourceibias.n153 commonsourceibias.n152 0.189894
R23204 commonsourceibias.n152 commonsourceibias.n119 0.189894
R23205 commonsourceibias.n148 commonsourceibias.n119 0.189894
R23206 commonsourceibias.n148 commonsourceibias.n147 0.189894
R23207 commonsourceibias.n147 commonsourceibias.n121 0.189894
R23208 commonsourceibias.n143 commonsourceibias.n121 0.189894
R23209 commonsourceibias.n143 commonsourceibias.n142 0.189894
R23210 commonsourceibias.n142 commonsourceibias.n123 0.189894
R23211 commonsourceibias.n137 commonsourceibias.n123 0.189894
R23212 commonsourceibias.n137 commonsourceibias.n136 0.189894
R23213 commonsourceibias.n136 commonsourceibias.n135 0.189894
R23214 commonsourceibias.n135 commonsourceibias.n125 0.189894
R23215 commonsourceibias.n130 commonsourceibias.n125 0.189894
R23216 commonsourceibias.n130 commonsourceibias.n129 0.189894
R23217 commonsourceibias.n188 commonsourceibias.n0 0.189894
R23218 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23219 commonsourceibias.n187 commonsourceibias.n186 0.189894
R23220 commonsourceibias.n186 commonsourceibias.n2 0.189894
R23221 commonsourceibias.n181 commonsourceibias.n2 0.189894
R23222 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23223 commonsourceibias.n180 commonsourceibias.n179 0.189894
R23224 commonsourceibias.n179 commonsourceibias.n4 0.189894
R23225 commonsourceibias.n174 commonsourceibias.n4 0.189894
R23226 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23227 commonsourceibias.n173 commonsourceibias.n172 0.189894
R23228 commonsourceibias.n172 commonsourceibias.n7 0.189894
R23229 commonsourceibias.n167 commonsourceibias.n7 0.189894
R23230 commonsourceibias.n167 commonsourceibias.n166 0.189894
R23231 commonsourceibias.n166 commonsourceibias.n165 0.189894
R23232 commonsourceibias.n165 commonsourceibias.n9 0.189894
R23233 commonsourceibias.n160 commonsourceibias.n9 0.189894
R23234 commonsourceibias.n277 commonsourceibias.n194 0.189894
R23235 commonsourceibias.n277 commonsourceibias.n276 0.189894
R23236 commonsourceibias.n276 commonsourceibias.n275 0.189894
R23237 commonsourceibias.n275 commonsourceibias.n196 0.189894
R23238 commonsourceibias.n270 commonsourceibias.n196 0.189894
R23239 commonsourceibias.n270 commonsourceibias.n269 0.189894
R23240 commonsourceibias.n269 commonsourceibias.n268 0.189894
R23241 commonsourceibias.n268 commonsourceibias.n198 0.189894
R23242 commonsourceibias.n263 commonsourceibias.n198 0.189894
R23243 commonsourceibias.n263 commonsourceibias.n262 0.189894
R23244 commonsourceibias.n262 commonsourceibias.n261 0.189894
R23245 commonsourceibias.n261 commonsourceibias.n201 0.189894
R23246 commonsourceibias.n256 commonsourceibias.n201 0.189894
R23247 commonsourceibias.n256 commonsourceibias.n255 0.189894
R23248 commonsourceibias.n255 commonsourceibias.n254 0.189894
R23249 commonsourceibias.n254 commonsourceibias.n203 0.189894
R23250 commonsourceibias.n249 commonsourceibias.n203 0.189894
R23251 commonsourceibias.n249 commonsourceibias.n248 0.189894
R23252 commonsourceibias.n248 commonsourceibias.n247 0.189894
R23253 commonsourceibias.n247 commonsourceibias.n206 0.189894
R23254 commonsourceibias.n242 commonsourceibias.n206 0.189894
R23255 commonsourceibias.n242 commonsourceibias.n241 0.189894
R23256 commonsourceibias.n241 commonsourceibias.n208 0.189894
R23257 commonsourceibias.n237 commonsourceibias.n208 0.189894
R23258 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23259 commonsourceibias.n236 commonsourceibias.n210 0.189894
R23260 commonsourceibias.n232 commonsourceibias.n210 0.189894
R23261 commonsourceibias.n232 commonsourceibias.n231 0.189894
R23262 commonsourceibias.n231 commonsourceibias.n212 0.189894
R23263 commonsourceibias.n226 commonsourceibias.n212 0.189894
R23264 commonsourceibias.n226 commonsourceibias.n225 0.189894
R23265 commonsourceibias.n225 commonsourceibias.n224 0.189894
R23266 commonsourceibias.n224 commonsourceibias.n214 0.189894
R23267 commonsourceibias.n219 commonsourceibias.n214 0.189894
R23268 commonsourceibias.n219 commonsourceibias.n218 0.189894
R23269 commonsourceibias.n366 commonsourceibias.n365 0.189894
R23270 commonsourceibias.n366 commonsourceibias.n361 0.189894
R23271 commonsourceibias.n371 commonsourceibias.n361 0.189894
R23272 commonsourceibias.n372 commonsourceibias.n371 0.189894
R23273 commonsourceibias.n373 commonsourceibias.n372 0.189894
R23274 commonsourceibias.n373 commonsourceibias.n359 0.189894
R23275 commonsourceibias.n378 commonsourceibias.n359 0.189894
R23276 commonsourceibias.n379 commonsourceibias.n378 0.189894
R23277 commonsourceibias.n379 commonsourceibias.n357 0.189894
R23278 commonsourceibias.n383 commonsourceibias.n357 0.189894
R23279 commonsourceibias.n384 commonsourceibias.n383 0.189894
R23280 commonsourceibias.n384 commonsourceibias.n355 0.189894
R23281 commonsourceibias.n388 commonsourceibias.n355 0.189894
R23282 commonsourceibias.n389 commonsourceibias.n388 0.189894
R23283 commonsourceibias.n389 commonsourceibias.n353 0.189894
R23284 commonsourceibias.n394 commonsourceibias.n353 0.189894
R23285 commonsourceibias.n395 commonsourceibias.n394 0.189894
R23286 commonsourceibias.n396 commonsourceibias.n395 0.189894
R23287 commonsourceibias.n396 commonsourceibias.n351 0.189894
R23288 commonsourceibias.n402 commonsourceibias.n351 0.189894
R23289 commonsourceibias.n403 commonsourceibias.n402 0.189894
R23290 commonsourceibias.n404 commonsourceibias.n403 0.189894
R23291 commonsourceibias.n404 commonsourceibias.n349 0.189894
R23292 commonsourceibias.n409 commonsourceibias.n349 0.189894
R23293 commonsourceibias.n410 commonsourceibias.n409 0.189894
R23294 commonsourceibias.n411 commonsourceibias.n410 0.189894
R23295 commonsourceibias.n411 commonsourceibias.n347 0.189894
R23296 commonsourceibias.n417 commonsourceibias.n347 0.189894
R23297 commonsourceibias.n418 commonsourceibias.n417 0.189894
R23298 commonsourceibias.n419 commonsourceibias.n418 0.189894
R23299 commonsourceibias.n419 commonsourceibias.n345 0.189894
R23300 commonsourceibias.n424 commonsourceibias.n345 0.189894
R23301 commonsourceibias.n425 commonsourceibias.n424 0.189894
R23302 commonsourceibias.n426 commonsourceibias.n425 0.189894
R23303 commonsourceibias.n426 commonsourceibias.n343 0.189894
R23304 commonsourceibias.n307 commonsourceibias.n306 0.189894
R23305 commonsourceibias.n307 commonsourceibias.n302 0.189894
R23306 commonsourceibias.n312 commonsourceibias.n302 0.189894
R23307 commonsourceibias.n313 commonsourceibias.n312 0.189894
R23308 commonsourceibias.n314 commonsourceibias.n313 0.189894
R23309 commonsourceibias.n314 commonsourceibias.n300 0.189894
R23310 commonsourceibias.n319 commonsourceibias.n300 0.189894
R23311 commonsourceibias.n320 commonsourceibias.n319 0.189894
R23312 commonsourceibias.n320 commonsourceibias.n298 0.189894
R23313 commonsourceibias.n324 commonsourceibias.n298 0.189894
R23314 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23315 commonsourceibias.n325 commonsourceibias.n296 0.189894
R23316 commonsourceibias.n329 commonsourceibias.n296 0.189894
R23317 commonsourceibias.n330 commonsourceibias.n329 0.189894
R23318 commonsourceibias.n330 commonsourceibias.n294 0.189894
R23319 commonsourceibias.n335 commonsourceibias.n294 0.189894
R23320 commonsourceibias.n442 commonsourceibias.n292 0.189894
R23321 commonsourceibias.n448 commonsourceibias.n292 0.189894
R23322 commonsourceibias.n449 commonsourceibias.n448 0.189894
R23323 commonsourceibias.n450 commonsourceibias.n449 0.189894
R23324 commonsourceibias.n450 commonsourceibias.n290 0.189894
R23325 commonsourceibias.n455 commonsourceibias.n290 0.189894
R23326 commonsourceibias.n456 commonsourceibias.n455 0.189894
R23327 commonsourceibias.n457 commonsourceibias.n456 0.189894
R23328 commonsourceibias.n457 commonsourceibias.n288 0.189894
R23329 commonsourceibias.n463 commonsourceibias.n288 0.189894
R23330 commonsourceibias.n464 commonsourceibias.n463 0.189894
R23331 commonsourceibias.n465 commonsourceibias.n464 0.189894
R23332 commonsourceibias.n465 commonsourceibias.n286 0.189894
R23333 commonsourceibias.n470 commonsourceibias.n286 0.189894
R23334 commonsourceibias.n471 commonsourceibias.n470 0.189894
R23335 commonsourceibias.n472 commonsourceibias.n471 0.189894
R23336 commonsourceibias.n472 commonsourceibias.n284 0.189894
R23337 commonsourceibias.n501 commonsourceibias.n500 0.189894
R23338 commonsourceibias.n501 commonsourceibias.n496 0.189894
R23339 commonsourceibias.n506 commonsourceibias.n496 0.189894
R23340 commonsourceibias.n507 commonsourceibias.n506 0.189894
R23341 commonsourceibias.n508 commonsourceibias.n507 0.189894
R23342 commonsourceibias.n508 commonsourceibias.n494 0.189894
R23343 commonsourceibias.n513 commonsourceibias.n494 0.189894
R23344 commonsourceibias.n514 commonsourceibias.n513 0.189894
R23345 commonsourceibias.n514 commonsourceibias.n492 0.189894
R23346 commonsourceibias.n518 commonsourceibias.n492 0.189894
R23347 commonsourceibias.n519 commonsourceibias.n518 0.189894
R23348 commonsourceibias.n519 commonsourceibias.n490 0.189894
R23349 commonsourceibias.n523 commonsourceibias.n490 0.189894
R23350 commonsourceibias.n524 commonsourceibias.n523 0.189894
R23351 commonsourceibias.n524 commonsourceibias.n488 0.189894
R23352 commonsourceibias.n529 commonsourceibias.n488 0.189894
R23353 commonsourceibias.n530 commonsourceibias.n529 0.189894
R23354 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23355 commonsourceibias.n531 commonsourceibias.n486 0.189894
R23356 commonsourceibias.n537 commonsourceibias.n486 0.189894
R23357 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23358 commonsourceibias.n539 commonsourceibias.n538 0.189894
R23359 commonsourceibias.n539 commonsourceibias.n484 0.189894
R23360 commonsourceibias.n544 commonsourceibias.n484 0.189894
R23361 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23362 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23363 commonsourceibias.n546 commonsourceibias.n482 0.189894
R23364 commonsourceibias.n552 commonsourceibias.n482 0.189894
R23365 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23366 commonsourceibias.n554 commonsourceibias.n553 0.189894
R23367 commonsourceibias.n554 commonsourceibias.n480 0.189894
R23368 commonsourceibias.n559 commonsourceibias.n480 0.189894
R23369 commonsourceibias.n560 commonsourceibias.n559 0.189894
R23370 commonsourceibias.n561 commonsourceibias.n560 0.189894
R23371 commonsourceibias.n561 commonsourceibias.n478 0.189894
R23372 commonsourceibias.n159 commonsourceibias.n158 0.170955
R23373 commonsourceibias.n160 commonsourceibias.n159 0.170955
R23374 commonsourceibias.n441 commonsourceibias.n335 0.170955
R23375 commonsourceibias.n442 commonsourceibias.n441 0.170955
R23376 diffpairibias.n0 diffpairibias.t27 436.822
R23377 diffpairibias.n27 diffpairibias.t24 435.479
R23378 diffpairibias.n26 diffpairibias.t21 435.479
R23379 diffpairibias.n25 diffpairibias.t22 435.479
R23380 diffpairibias.n24 diffpairibias.t26 435.479
R23381 diffpairibias.n23 diffpairibias.t20 435.479
R23382 diffpairibias.n0 diffpairibias.t23 435.479
R23383 diffpairibias.n1 diffpairibias.t28 435.479
R23384 diffpairibias.n2 diffpairibias.t25 435.479
R23385 diffpairibias.n3 diffpairibias.t29 435.479
R23386 diffpairibias.n13 diffpairibias.t14 377.536
R23387 diffpairibias.n13 diffpairibias.t0 376.193
R23388 diffpairibias.n14 diffpairibias.t10 376.193
R23389 diffpairibias.n15 diffpairibias.t12 376.193
R23390 diffpairibias.n16 diffpairibias.t6 376.193
R23391 diffpairibias.n17 diffpairibias.t2 376.193
R23392 diffpairibias.n18 diffpairibias.t16 376.193
R23393 diffpairibias.n19 diffpairibias.t4 376.193
R23394 diffpairibias.n20 diffpairibias.t18 376.193
R23395 diffpairibias.n21 diffpairibias.t8 376.193
R23396 diffpairibias.n4 diffpairibias.t15 113.368
R23397 diffpairibias.n4 diffpairibias.t1 112.698
R23398 diffpairibias.n5 diffpairibias.t11 112.698
R23399 diffpairibias.n6 diffpairibias.t13 112.698
R23400 diffpairibias.n7 diffpairibias.t7 112.698
R23401 diffpairibias.n8 diffpairibias.t3 112.698
R23402 diffpairibias.n9 diffpairibias.t17 112.698
R23403 diffpairibias.n10 diffpairibias.t5 112.698
R23404 diffpairibias.n11 diffpairibias.t19 112.698
R23405 diffpairibias.n12 diffpairibias.t9 112.698
R23406 diffpairibias.n22 diffpairibias.n21 4.77242
R23407 diffpairibias.n22 diffpairibias.n12 4.30807
R23408 diffpairibias.n23 diffpairibias.n22 4.13945
R23409 diffpairibias.n21 diffpairibias.n20 1.34352
R23410 diffpairibias.n20 diffpairibias.n19 1.34352
R23411 diffpairibias.n19 diffpairibias.n18 1.34352
R23412 diffpairibias.n18 diffpairibias.n17 1.34352
R23413 diffpairibias.n17 diffpairibias.n16 1.34352
R23414 diffpairibias.n16 diffpairibias.n15 1.34352
R23415 diffpairibias.n15 diffpairibias.n14 1.34352
R23416 diffpairibias.n14 diffpairibias.n13 1.34352
R23417 diffpairibias.n3 diffpairibias.n2 1.34352
R23418 diffpairibias.n2 diffpairibias.n1 1.34352
R23419 diffpairibias.n1 diffpairibias.n0 1.34352
R23420 diffpairibias.n24 diffpairibias.n23 1.34352
R23421 diffpairibias.n25 diffpairibias.n24 1.34352
R23422 diffpairibias.n26 diffpairibias.n25 1.34352
R23423 diffpairibias.n27 diffpairibias.n26 1.34352
R23424 diffpairibias.n28 diffpairibias.n27 0.862419
R23425 diffpairibias diffpairibias.n28 0.684875
R23426 diffpairibias.n12 diffpairibias.n11 0.672012
R23427 diffpairibias.n11 diffpairibias.n10 0.672012
R23428 diffpairibias.n10 diffpairibias.n9 0.672012
R23429 diffpairibias.n9 diffpairibias.n8 0.672012
R23430 diffpairibias.n8 diffpairibias.n7 0.672012
R23431 diffpairibias.n7 diffpairibias.n6 0.672012
R23432 diffpairibias.n6 diffpairibias.n5 0.672012
R23433 diffpairibias.n5 diffpairibias.n4 0.672012
R23434 diffpairibias.n28 diffpairibias.n3 0.190907
R23435 output.n41 output.n15 289.615
R23436 output.n72 output.n46 289.615
R23437 output.n104 output.n78 289.615
R23438 output.n136 output.n110 289.615
R23439 output.n77 output.n45 197.26
R23440 output.n77 output.n76 196.298
R23441 output.n109 output.n108 196.298
R23442 output.n141 output.n140 196.298
R23443 output.n42 output.n41 185
R23444 output.n40 output.n39 185
R23445 output.n19 output.n18 185
R23446 output.n34 output.n33 185
R23447 output.n32 output.n31 185
R23448 output.n23 output.n22 185
R23449 output.n26 output.n25 185
R23450 output.n73 output.n72 185
R23451 output.n71 output.n70 185
R23452 output.n50 output.n49 185
R23453 output.n65 output.n64 185
R23454 output.n63 output.n62 185
R23455 output.n54 output.n53 185
R23456 output.n57 output.n56 185
R23457 output.n105 output.n104 185
R23458 output.n103 output.n102 185
R23459 output.n82 output.n81 185
R23460 output.n97 output.n96 185
R23461 output.n95 output.n94 185
R23462 output.n86 output.n85 185
R23463 output.n89 output.n88 185
R23464 output.n137 output.n136 185
R23465 output.n135 output.n134 185
R23466 output.n114 output.n113 185
R23467 output.n129 output.n128 185
R23468 output.n127 output.n126 185
R23469 output.n118 output.n117 185
R23470 output.n121 output.n120 185
R23471 output.t1 output.n24 147.661
R23472 output.t19 output.n55 147.661
R23473 output.t0 output.n87 147.661
R23474 output.t2 output.n119 147.661
R23475 output.n41 output.n40 104.615
R23476 output.n40 output.n18 104.615
R23477 output.n33 output.n18 104.615
R23478 output.n33 output.n32 104.615
R23479 output.n32 output.n22 104.615
R23480 output.n25 output.n22 104.615
R23481 output.n72 output.n71 104.615
R23482 output.n71 output.n49 104.615
R23483 output.n64 output.n49 104.615
R23484 output.n64 output.n63 104.615
R23485 output.n63 output.n53 104.615
R23486 output.n56 output.n53 104.615
R23487 output.n104 output.n103 104.615
R23488 output.n103 output.n81 104.615
R23489 output.n96 output.n81 104.615
R23490 output.n96 output.n95 104.615
R23491 output.n95 output.n85 104.615
R23492 output.n88 output.n85 104.615
R23493 output.n136 output.n135 104.615
R23494 output.n135 output.n113 104.615
R23495 output.n128 output.n113 104.615
R23496 output.n128 output.n127 104.615
R23497 output.n127 output.n117 104.615
R23498 output.n120 output.n117 104.615
R23499 output.n1 output.t15 77.056
R23500 output.n14 output.t16 76.6694
R23501 output.n1 output.n0 72.7095
R23502 output.n3 output.n2 72.7095
R23503 output.n5 output.n4 72.7095
R23504 output.n7 output.n6 72.7095
R23505 output.n9 output.n8 72.7095
R23506 output.n11 output.n10 72.7095
R23507 output.n13 output.n12 72.7095
R23508 output.n25 output.t1 52.3082
R23509 output.n56 output.t19 52.3082
R23510 output.n88 output.t0 52.3082
R23511 output.n120 output.t2 52.3082
R23512 output.n26 output.n24 15.6674
R23513 output.n57 output.n55 15.6674
R23514 output.n89 output.n87 15.6674
R23515 output.n121 output.n119 15.6674
R23516 output.n27 output.n23 12.8005
R23517 output.n58 output.n54 12.8005
R23518 output.n90 output.n86 12.8005
R23519 output.n122 output.n118 12.8005
R23520 output.n31 output.n30 12.0247
R23521 output.n62 output.n61 12.0247
R23522 output.n94 output.n93 12.0247
R23523 output.n126 output.n125 12.0247
R23524 output.n34 output.n21 11.249
R23525 output.n65 output.n52 11.249
R23526 output.n97 output.n84 11.249
R23527 output.n129 output.n116 11.249
R23528 output.n35 output.n19 10.4732
R23529 output.n66 output.n50 10.4732
R23530 output.n98 output.n82 10.4732
R23531 output.n130 output.n114 10.4732
R23532 output.n39 output.n38 9.69747
R23533 output.n70 output.n69 9.69747
R23534 output.n102 output.n101 9.69747
R23535 output.n134 output.n133 9.69747
R23536 output.n45 output.n44 9.45567
R23537 output.n76 output.n75 9.45567
R23538 output.n108 output.n107 9.45567
R23539 output.n140 output.n139 9.45567
R23540 output.n44 output.n43 9.3005
R23541 output.n17 output.n16 9.3005
R23542 output.n38 output.n37 9.3005
R23543 output.n36 output.n35 9.3005
R23544 output.n21 output.n20 9.3005
R23545 output.n30 output.n29 9.3005
R23546 output.n28 output.n27 9.3005
R23547 output.n75 output.n74 9.3005
R23548 output.n48 output.n47 9.3005
R23549 output.n69 output.n68 9.3005
R23550 output.n67 output.n66 9.3005
R23551 output.n52 output.n51 9.3005
R23552 output.n61 output.n60 9.3005
R23553 output.n59 output.n58 9.3005
R23554 output.n107 output.n106 9.3005
R23555 output.n80 output.n79 9.3005
R23556 output.n101 output.n100 9.3005
R23557 output.n99 output.n98 9.3005
R23558 output.n84 output.n83 9.3005
R23559 output.n93 output.n92 9.3005
R23560 output.n91 output.n90 9.3005
R23561 output.n139 output.n138 9.3005
R23562 output.n112 output.n111 9.3005
R23563 output.n133 output.n132 9.3005
R23564 output.n131 output.n130 9.3005
R23565 output.n116 output.n115 9.3005
R23566 output.n125 output.n124 9.3005
R23567 output.n123 output.n122 9.3005
R23568 output.n42 output.n17 8.92171
R23569 output.n73 output.n48 8.92171
R23570 output.n105 output.n80 8.92171
R23571 output.n137 output.n112 8.92171
R23572 output output.n141 8.15037
R23573 output.n43 output.n15 8.14595
R23574 output.n74 output.n46 8.14595
R23575 output.n106 output.n78 8.14595
R23576 output.n138 output.n110 8.14595
R23577 output.n45 output.n15 5.81868
R23578 output.n76 output.n46 5.81868
R23579 output.n108 output.n78 5.81868
R23580 output.n140 output.n110 5.81868
R23581 output.n43 output.n42 5.04292
R23582 output.n74 output.n73 5.04292
R23583 output.n106 output.n105 5.04292
R23584 output.n138 output.n137 5.04292
R23585 output.n28 output.n24 4.38594
R23586 output.n59 output.n55 4.38594
R23587 output.n91 output.n87 4.38594
R23588 output.n123 output.n119 4.38594
R23589 output.n39 output.n17 4.26717
R23590 output.n70 output.n48 4.26717
R23591 output.n102 output.n80 4.26717
R23592 output.n134 output.n112 4.26717
R23593 output.n0 output.t5 3.9605
R23594 output.n0 output.t9 3.9605
R23595 output.n2 output.t12 3.9605
R23596 output.n2 output.t17 3.9605
R23597 output.n4 output.t18 3.9605
R23598 output.n4 output.t7 3.9605
R23599 output.n6 output.t11 3.9605
R23600 output.n6 output.t3 3.9605
R23601 output.n8 output.t6 3.9605
R23602 output.n8 output.t4 3.9605
R23603 output.n10 output.t10 3.9605
R23604 output.n10 output.t13 3.9605
R23605 output.n12 output.t14 3.9605
R23606 output.n12 output.t8 3.9605
R23607 output.n38 output.n19 3.49141
R23608 output.n69 output.n50 3.49141
R23609 output.n101 output.n82 3.49141
R23610 output.n133 output.n114 3.49141
R23611 output.n35 output.n34 2.71565
R23612 output.n66 output.n65 2.71565
R23613 output.n98 output.n97 2.71565
R23614 output.n130 output.n129 2.71565
R23615 output.n31 output.n21 1.93989
R23616 output.n62 output.n52 1.93989
R23617 output.n94 output.n84 1.93989
R23618 output.n126 output.n116 1.93989
R23619 output.n30 output.n23 1.16414
R23620 output.n61 output.n54 1.16414
R23621 output.n93 output.n86 1.16414
R23622 output.n125 output.n118 1.16414
R23623 output.n141 output.n109 0.962709
R23624 output.n109 output.n77 0.962709
R23625 output.n27 output.n26 0.388379
R23626 output.n58 output.n57 0.388379
R23627 output.n90 output.n89 0.388379
R23628 output.n122 output.n121 0.388379
R23629 output.n14 output.n13 0.387128
R23630 output.n13 output.n11 0.387128
R23631 output.n11 output.n9 0.387128
R23632 output.n9 output.n7 0.387128
R23633 output.n7 output.n5 0.387128
R23634 output.n5 output.n3 0.387128
R23635 output.n3 output.n1 0.387128
R23636 output.n44 output.n16 0.155672
R23637 output.n37 output.n16 0.155672
R23638 output.n37 output.n36 0.155672
R23639 output.n36 output.n20 0.155672
R23640 output.n29 output.n20 0.155672
R23641 output.n29 output.n28 0.155672
R23642 output.n75 output.n47 0.155672
R23643 output.n68 output.n47 0.155672
R23644 output.n68 output.n67 0.155672
R23645 output.n67 output.n51 0.155672
R23646 output.n60 output.n51 0.155672
R23647 output.n60 output.n59 0.155672
R23648 output.n107 output.n79 0.155672
R23649 output.n100 output.n79 0.155672
R23650 output.n100 output.n99 0.155672
R23651 output.n99 output.n83 0.155672
R23652 output.n92 output.n83 0.155672
R23653 output.n92 output.n91 0.155672
R23654 output.n139 output.n111 0.155672
R23655 output.n132 output.n111 0.155672
R23656 output.n132 output.n131 0.155672
R23657 output.n131 output.n115 0.155672
R23658 output.n124 output.n115 0.155672
R23659 output.n124 output.n123 0.155672
R23660 output output.n14 0.126227
R23661 a_n2318_8322.n8 a_n2318_8322.t19 74.6477
R23662 a_n2318_8322.n1 a_n2318_8322.t14 74.6477
R23663 a_n2318_8322.n20 a_n2318_8322.t13 74.6474
R23664 a_n2318_8322.n16 a_n2318_8322.t3 74.2899
R23665 a_n2318_8322.n9 a_n2318_8322.t17 74.2899
R23666 a_n2318_8322.n10 a_n2318_8322.t20 74.2899
R23667 a_n2318_8322.n13 a_n2318_8322.t21 74.2899
R23668 a_n2318_8322.n6 a_n2318_8322.t0 74.2899
R23669 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23670 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23671 a_n2318_8322.n8 a_n2318_8322.n7 70.6783
R23672 a_n2318_8322.n12 a_n2318_8322.n11 70.6783
R23673 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23674 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23675 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23676 a_n2318_8322.n22 a_n2318_8322.n21 70.6782
R23677 a_n2318_8322.n14 a_n2318_8322.n6 23.4712
R23678 a_n2318_8322.n15 a_n2318_8322.t24 10.0049
R23679 a_n2318_8322.n14 a_n2318_8322.n13 6.95632
R23680 a_n2318_8322.n16 a_n2318_8322.n15 6.19447
R23681 a_n2318_8322.n15 a_n2318_8322.n14 5.3452
R23682 a_n2318_8322.n19 a_n2318_8322.t10 3.61217
R23683 a_n2318_8322.n19 a_n2318_8322.t7 3.61217
R23684 a_n2318_8322.n17 a_n2318_8322.t12 3.61217
R23685 a_n2318_8322.n17 a_n2318_8322.t5 3.61217
R23686 a_n2318_8322.n7 a_n2318_8322.t23 3.61217
R23687 a_n2318_8322.n7 a_n2318_8322.t22 3.61217
R23688 a_n2318_8322.n11 a_n2318_8322.t18 3.61217
R23689 a_n2318_8322.n11 a_n2318_8322.t16 3.61217
R23690 a_n2318_8322.n0 a_n2318_8322.t2 3.61217
R23691 a_n2318_8322.n0 a_n2318_8322.t1 3.61217
R23692 a_n2318_8322.n2 a_n2318_8322.t11 3.61217
R23693 a_n2318_8322.n2 a_n2318_8322.t6 3.61217
R23694 a_n2318_8322.n4 a_n2318_8322.t9 3.61217
R23695 a_n2318_8322.n4 a_n2318_8322.t8 3.61217
R23696 a_n2318_8322.n22 a_n2318_8322.t4 3.61217
R23697 a_n2318_8322.t15 a_n2318_8322.n22 3.61217
R23698 a_n2318_8322.n13 a_n2318_8322.n12 0.358259
R23699 a_n2318_8322.n12 a_n2318_8322.n10 0.358259
R23700 a_n2318_8322.n9 a_n2318_8322.n8 0.358259
R23701 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23702 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23703 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23704 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23705 a_n2318_8322.n21 a_n2318_8322.n18 0.358259
R23706 a_n2318_8322.n21 a_n2318_8322.n20 0.358259
R23707 a_n2318_8322.n10 a_n2318_8322.n9 0.101793
R23708 a_n2318_8322.t26 a_n2318_8322.t27 0.0788333
R23709 a_n2318_8322.t25 a_n2318_8322.t26 0.0631667
R23710 a_n2318_8322.t24 a_n2318_8322.t25 0.0471944
R23711 a_n2318_8322.t24 a_n2318_8322.t27 0.0453889
R23712 outputibias.n27 outputibias.n1 289.615
R23713 outputibias.n58 outputibias.n32 289.615
R23714 outputibias.n90 outputibias.n64 289.615
R23715 outputibias.n122 outputibias.n96 289.615
R23716 outputibias.n28 outputibias.n27 185
R23717 outputibias.n26 outputibias.n25 185
R23718 outputibias.n5 outputibias.n4 185
R23719 outputibias.n20 outputibias.n19 185
R23720 outputibias.n18 outputibias.n17 185
R23721 outputibias.n9 outputibias.n8 185
R23722 outputibias.n12 outputibias.n11 185
R23723 outputibias.n59 outputibias.n58 185
R23724 outputibias.n57 outputibias.n56 185
R23725 outputibias.n36 outputibias.n35 185
R23726 outputibias.n51 outputibias.n50 185
R23727 outputibias.n49 outputibias.n48 185
R23728 outputibias.n40 outputibias.n39 185
R23729 outputibias.n43 outputibias.n42 185
R23730 outputibias.n91 outputibias.n90 185
R23731 outputibias.n89 outputibias.n88 185
R23732 outputibias.n68 outputibias.n67 185
R23733 outputibias.n83 outputibias.n82 185
R23734 outputibias.n81 outputibias.n80 185
R23735 outputibias.n72 outputibias.n71 185
R23736 outputibias.n75 outputibias.n74 185
R23737 outputibias.n123 outputibias.n122 185
R23738 outputibias.n121 outputibias.n120 185
R23739 outputibias.n100 outputibias.n99 185
R23740 outputibias.n115 outputibias.n114 185
R23741 outputibias.n113 outputibias.n112 185
R23742 outputibias.n104 outputibias.n103 185
R23743 outputibias.n107 outputibias.n106 185
R23744 outputibias.n0 outputibias.t8 178.945
R23745 outputibias.n133 outputibias.t11 177.018
R23746 outputibias.n132 outputibias.t9 177.018
R23747 outputibias.n0 outputibias.t10 177.018
R23748 outputibias.t5 outputibias.n10 147.661
R23749 outputibias.t7 outputibias.n41 147.661
R23750 outputibias.t1 outputibias.n73 147.661
R23751 outputibias.t3 outputibias.n105 147.661
R23752 outputibias.n128 outputibias.t4 132.363
R23753 outputibias.n128 outputibias.t6 130.436
R23754 outputibias.n129 outputibias.t0 130.436
R23755 outputibias.n130 outputibias.t2 130.436
R23756 outputibias.n27 outputibias.n26 104.615
R23757 outputibias.n26 outputibias.n4 104.615
R23758 outputibias.n19 outputibias.n4 104.615
R23759 outputibias.n19 outputibias.n18 104.615
R23760 outputibias.n18 outputibias.n8 104.615
R23761 outputibias.n11 outputibias.n8 104.615
R23762 outputibias.n58 outputibias.n57 104.615
R23763 outputibias.n57 outputibias.n35 104.615
R23764 outputibias.n50 outputibias.n35 104.615
R23765 outputibias.n50 outputibias.n49 104.615
R23766 outputibias.n49 outputibias.n39 104.615
R23767 outputibias.n42 outputibias.n39 104.615
R23768 outputibias.n90 outputibias.n89 104.615
R23769 outputibias.n89 outputibias.n67 104.615
R23770 outputibias.n82 outputibias.n67 104.615
R23771 outputibias.n82 outputibias.n81 104.615
R23772 outputibias.n81 outputibias.n71 104.615
R23773 outputibias.n74 outputibias.n71 104.615
R23774 outputibias.n122 outputibias.n121 104.615
R23775 outputibias.n121 outputibias.n99 104.615
R23776 outputibias.n114 outputibias.n99 104.615
R23777 outputibias.n114 outputibias.n113 104.615
R23778 outputibias.n113 outputibias.n103 104.615
R23779 outputibias.n106 outputibias.n103 104.615
R23780 outputibias.n63 outputibias.n31 95.6354
R23781 outputibias.n63 outputibias.n62 94.6732
R23782 outputibias.n95 outputibias.n94 94.6732
R23783 outputibias.n127 outputibias.n126 94.6732
R23784 outputibias.n11 outputibias.t5 52.3082
R23785 outputibias.n42 outputibias.t7 52.3082
R23786 outputibias.n74 outputibias.t1 52.3082
R23787 outputibias.n106 outputibias.t3 52.3082
R23788 outputibias.n12 outputibias.n10 15.6674
R23789 outputibias.n43 outputibias.n41 15.6674
R23790 outputibias.n75 outputibias.n73 15.6674
R23791 outputibias.n107 outputibias.n105 15.6674
R23792 outputibias.n13 outputibias.n9 12.8005
R23793 outputibias.n44 outputibias.n40 12.8005
R23794 outputibias.n76 outputibias.n72 12.8005
R23795 outputibias.n108 outputibias.n104 12.8005
R23796 outputibias.n17 outputibias.n16 12.0247
R23797 outputibias.n48 outputibias.n47 12.0247
R23798 outputibias.n80 outputibias.n79 12.0247
R23799 outputibias.n112 outputibias.n111 12.0247
R23800 outputibias.n20 outputibias.n7 11.249
R23801 outputibias.n51 outputibias.n38 11.249
R23802 outputibias.n83 outputibias.n70 11.249
R23803 outputibias.n115 outputibias.n102 11.249
R23804 outputibias.n21 outputibias.n5 10.4732
R23805 outputibias.n52 outputibias.n36 10.4732
R23806 outputibias.n84 outputibias.n68 10.4732
R23807 outputibias.n116 outputibias.n100 10.4732
R23808 outputibias.n25 outputibias.n24 9.69747
R23809 outputibias.n56 outputibias.n55 9.69747
R23810 outputibias.n88 outputibias.n87 9.69747
R23811 outputibias.n120 outputibias.n119 9.69747
R23812 outputibias.n31 outputibias.n30 9.45567
R23813 outputibias.n62 outputibias.n61 9.45567
R23814 outputibias.n94 outputibias.n93 9.45567
R23815 outputibias.n126 outputibias.n125 9.45567
R23816 outputibias.n30 outputibias.n29 9.3005
R23817 outputibias.n3 outputibias.n2 9.3005
R23818 outputibias.n24 outputibias.n23 9.3005
R23819 outputibias.n22 outputibias.n21 9.3005
R23820 outputibias.n7 outputibias.n6 9.3005
R23821 outputibias.n16 outputibias.n15 9.3005
R23822 outputibias.n14 outputibias.n13 9.3005
R23823 outputibias.n61 outputibias.n60 9.3005
R23824 outputibias.n34 outputibias.n33 9.3005
R23825 outputibias.n55 outputibias.n54 9.3005
R23826 outputibias.n53 outputibias.n52 9.3005
R23827 outputibias.n38 outputibias.n37 9.3005
R23828 outputibias.n47 outputibias.n46 9.3005
R23829 outputibias.n45 outputibias.n44 9.3005
R23830 outputibias.n93 outputibias.n92 9.3005
R23831 outputibias.n66 outputibias.n65 9.3005
R23832 outputibias.n87 outputibias.n86 9.3005
R23833 outputibias.n85 outputibias.n84 9.3005
R23834 outputibias.n70 outputibias.n69 9.3005
R23835 outputibias.n79 outputibias.n78 9.3005
R23836 outputibias.n77 outputibias.n76 9.3005
R23837 outputibias.n125 outputibias.n124 9.3005
R23838 outputibias.n98 outputibias.n97 9.3005
R23839 outputibias.n119 outputibias.n118 9.3005
R23840 outputibias.n117 outputibias.n116 9.3005
R23841 outputibias.n102 outputibias.n101 9.3005
R23842 outputibias.n111 outputibias.n110 9.3005
R23843 outputibias.n109 outputibias.n108 9.3005
R23844 outputibias.n28 outputibias.n3 8.92171
R23845 outputibias.n59 outputibias.n34 8.92171
R23846 outputibias.n91 outputibias.n66 8.92171
R23847 outputibias.n123 outputibias.n98 8.92171
R23848 outputibias.n29 outputibias.n1 8.14595
R23849 outputibias.n60 outputibias.n32 8.14595
R23850 outputibias.n92 outputibias.n64 8.14595
R23851 outputibias.n124 outputibias.n96 8.14595
R23852 outputibias.n31 outputibias.n1 5.81868
R23853 outputibias.n62 outputibias.n32 5.81868
R23854 outputibias.n94 outputibias.n64 5.81868
R23855 outputibias.n126 outputibias.n96 5.81868
R23856 outputibias.n131 outputibias.n130 5.20947
R23857 outputibias.n29 outputibias.n28 5.04292
R23858 outputibias.n60 outputibias.n59 5.04292
R23859 outputibias.n92 outputibias.n91 5.04292
R23860 outputibias.n124 outputibias.n123 5.04292
R23861 outputibias.n131 outputibias.n127 4.42209
R23862 outputibias.n14 outputibias.n10 4.38594
R23863 outputibias.n45 outputibias.n41 4.38594
R23864 outputibias.n77 outputibias.n73 4.38594
R23865 outputibias.n109 outputibias.n105 4.38594
R23866 outputibias.n132 outputibias.n131 4.28454
R23867 outputibias.n25 outputibias.n3 4.26717
R23868 outputibias.n56 outputibias.n34 4.26717
R23869 outputibias.n88 outputibias.n66 4.26717
R23870 outputibias.n120 outputibias.n98 4.26717
R23871 outputibias.n24 outputibias.n5 3.49141
R23872 outputibias.n55 outputibias.n36 3.49141
R23873 outputibias.n87 outputibias.n68 3.49141
R23874 outputibias.n119 outputibias.n100 3.49141
R23875 outputibias.n21 outputibias.n20 2.71565
R23876 outputibias.n52 outputibias.n51 2.71565
R23877 outputibias.n84 outputibias.n83 2.71565
R23878 outputibias.n116 outputibias.n115 2.71565
R23879 outputibias.n17 outputibias.n7 1.93989
R23880 outputibias.n48 outputibias.n38 1.93989
R23881 outputibias.n80 outputibias.n70 1.93989
R23882 outputibias.n112 outputibias.n102 1.93989
R23883 outputibias.n130 outputibias.n129 1.9266
R23884 outputibias.n129 outputibias.n128 1.9266
R23885 outputibias.n133 outputibias.n132 1.92658
R23886 outputibias.n134 outputibias.n133 1.29913
R23887 outputibias.n16 outputibias.n9 1.16414
R23888 outputibias.n47 outputibias.n40 1.16414
R23889 outputibias.n79 outputibias.n72 1.16414
R23890 outputibias.n111 outputibias.n104 1.16414
R23891 outputibias.n127 outputibias.n95 0.962709
R23892 outputibias.n95 outputibias.n63 0.962709
R23893 outputibias.n13 outputibias.n12 0.388379
R23894 outputibias.n44 outputibias.n43 0.388379
R23895 outputibias.n76 outputibias.n75 0.388379
R23896 outputibias.n108 outputibias.n107 0.388379
R23897 outputibias.n134 outputibias.n0 0.337251
R23898 outputibias outputibias.n134 0.302375
R23899 outputibias.n30 outputibias.n2 0.155672
R23900 outputibias.n23 outputibias.n2 0.155672
R23901 outputibias.n23 outputibias.n22 0.155672
R23902 outputibias.n22 outputibias.n6 0.155672
R23903 outputibias.n15 outputibias.n6 0.155672
R23904 outputibias.n15 outputibias.n14 0.155672
R23905 outputibias.n61 outputibias.n33 0.155672
R23906 outputibias.n54 outputibias.n33 0.155672
R23907 outputibias.n54 outputibias.n53 0.155672
R23908 outputibias.n53 outputibias.n37 0.155672
R23909 outputibias.n46 outputibias.n37 0.155672
R23910 outputibias.n46 outputibias.n45 0.155672
R23911 outputibias.n93 outputibias.n65 0.155672
R23912 outputibias.n86 outputibias.n65 0.155672
R23913 outputibias.n86 outputibias.n85 0.155672
R23914 outputibias.n85 outputibias.n69 0.155672
R23915 outputibias.n78 outputibias.n69 0.155672
R23916 outputibias.n78 outputibias.n77 0.155672
R23917 outputibias.n125 outputibias.n97 0.155672
R23918 outputibias.n118 outputibias.n97 0.155672
R23919 outputibias.n118 outputibias.n117 0.155672
R23920 outputibias.n117 outputibias.n101 0.155672
R23921 outputibias.n110 outputibias.n101 0.155672
R23922 outputibias.n110 outputibias.n109 0.155672
C0 commonsourceibias outputibias 0.003832f
C1 plus diffpairibias 4.56e-19
C2 vdd commonsourceibias 0.004218f
C3 CSoutput plus 0.892085f
C4 commonsourceibias diffpairibias 0.052527f
C5 CSoutput commonsourceibias 37.4715f
C6 minus plus 9.92364f
C7 minus commonsourceibias 0.337549f
C8 plus commonsourceibias 0.283677f
C9 output outputibias 2.34152f
C10 vdd output 7.23429f
C11 CSoutput output 6.13571f
C12 CSoutput outputibias 0.032386f
C13 vdd CSoutput 0.140911p
C14 minus diffpairibias 4.33e-19
C15 commonsourceibias output 0.006808f
C16 CSoutput minus 2.89653f
C17 vdd plus 0.095768f
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150736p
C22 plus gnd 36.8535f
C23 minus gnd 30.064781f
C24 CSoutput gnd 0.102341p
C25 vdd gnd 0.474239p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t5 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t7 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t3 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t2 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t6 gnd 0.108319f
C163 outputibias.t4 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 a_n2318_8322.t27 gnd 39.5861f
C174 a_n2318_8322.t24 gnd 29.0796f
C175 a_n2318_8322.t26 gnd 19.7234f
C176 a_n2318_8322.t25 gnd 39.5861f
C177 a_n2318_8322.t4 gnd 0.095743f
C178 a_n2318_8322.t14 gnd 0.896485f
C179 a_n2318_8322.t2 gnd 0.095743f
C180 a_n2318_8322.t1 gnd 0.095743f
C181 a_n2318_8322.n0 gnd 0.674411f
C182 a_n2318_8322.n1 gnd 0.753555f
C183 a_n2318_8322.t11 gnd 0.095743f
C184 a_n2318_8322.t6 gnd 0.095743f
C185 a_n2318_8322.n2 gnd 0.674411f
C186 a_n2318_8322.n3 gnd 0.382872f
C187 a_n2318_8322.t9 gnd 0.095743f
C188 a_n2318_8322.t8 gnd 0.095743f
C189 a_n2318_8322.n4 gnd 0.674411f
C190 a_n2318_8322.n5 gnd 0.382872f
C191 a_n2318_8322.t0 gnd 0.8947f
C192 a_n2318_8322.n6 gnd 1.55065f
C193 a_n2318_8322.t19 gnd 0.896485f
C194 a_n2318_8322.t23 gnd 0.095743f
C195 a_n2318_8322.t22 gnd 0.095743f
C196 a_n2318_8322.n7 gnd 0.674411f
C197 a_n2318_8322.n8 gnd 0.753555f
C198 a_n2318_8322.t17 gnd 0.8947f
C199 a_n2318_8322.n9 gnd 0.379199f
C200 a_n2318_8322.t20 gnd 0.8947f
C201 a_n2318_8322.n10 gnd 0.379199f
C202 a_n2318_8322.t18 gnd 0.095743f
C203 a_n2318_8322.t16 gnd 0.095743f
C204 a_n2318_8322.n11 gnd 0.674411f
C205 a_n2318_8322.n12 gnd 0.382872f
C206 a_n2318_8322.t21 gnd 0.8947f
C207 a_n2318_8322.n13 gnd 1.0738f
C208 a_n2318_8322.n14 gnd 1.82539f
C209 a_n2318_8322.n15 gnd 3.67064f
C210 a_n2318_8322.t3 gnd 0.8947f
C211 a_n2318_8322.n16 gnd 0.880763f
C212 a_n2318_8322.t12 gnd 0.095743f
C213 a_n2318_8322.t5 gnd 0.095743f
C214 a_n2318_8322.n17 gnd 0.674411f
C215 a_n2318_8322.n18 gnd 0.382872f
C216 a_n2318_8322.t13 gnd 0.896483f
C217 a_n2318_8322.t10 gnd 0.095743f
C218 a_n2318_8322.t7 gnd 0.095743f
C219 a_n2318_8322.n19 gnd 0.674411f
C220 a_n2318_8322.n20 gnd 0.753557f
C221 a_n2318_8322.n21 gnd 0.38287f
C222 a_n2318_8322.n22 gnd 0.674413f
C223 a_n2318_8322.t15 gnd 0.095743f
C224 output.t15 gnd 0.464308f
C225 output.t5 gnd 0.044422f
C226 output.t9 gnd 0.044422f
C227 output.n0 gnd 0.364624f
C228 output.n1 gnd 0.614102f
C229 output.t12 gnd 0.044422f
C230 output.t17 gnd 0.044422f
C231 output.n2 gnd 0.364624f
C232 output.n3 gnd 0.350265f
C233 output.t18 gnd 0.044422f
C234 output.t7 gnd 0.044422f
C235 output.n4 gnd 0.364624f
C236 output.n5 gnd 0.350265f
C237 output.t11 gnd 0.044422f
C238 output.t3 gnd 0.044422f
C239 output.n6 gnd 0.364624f
C240 output.n7 gnd 0.350265f
C241 output.t6 gnd 0.044422f
C242 output.t4 gnd 0.044422f
C243 output.n8 gnd 0.364624f
C244 output.n9 gnd 0.350265f
C245 output.t10 gnd 0.044422f
C246 output.t13 gnd 0.044422f
C247 output.n10 gnd 0.364624f
C248 output.n11 gnd 0.350265f
C249 output.t14 gnd 0.044422f
C250 output.t8 gnd 0.044422f
C251 output.n12 gnd 0.364624f
C252 output.n13 gnd 0.350265f
C253 output.t16 gnd 0.462979f
C254 output.n14 gnd 0.28994f
C255 output.n15 gnd 0.015803f
C256 output.n16 gnd 0.011243f
C257 output.n17 gnd 0.006041f
C258 output.n18 gnd 0.01428f
C259 output.n19 gnd 0.006397f
C260 output.n20 gnd 0.011243f
C261 output.n21 gnd 0.006041f
C262 output.n22 gnd 0.01428f
C263 output.n23 gnd 0.006397f
C264 output.n24 gnd 0.048111f
C265 output.t1 gnd 0.023274f
C266 output.n25 gnd 0.01071f
C267 output.n26 gnd 0.008435f
C268 output.n27 gnd 0.006041f
C269 output.n28 gnd 0.267512f
C270 output.n29 gnd 0.011243f
C271 output.n30 gnd 0.006041f
C272 output.n31 gnd 0.006397f
C273 output.n32 gnd 0.01428f
C274 output.n33 gnd 0.01428f
C275 output.n34 gnd 0.006397f
C276 output.n35 gnd 0.006041f
C277 output.n36 gnd 0.011243f
C278 output.n37 gnd 0.011243f
C279 output.n38 gnd 0.006041f
C280 output.n39 gnd 0.006397f
C281 output.n40 gnd 0.01428f
C282 output.n41 gnd 0.030913f
C283 output.n42 gnd 0.006397f
C284 output.n43 gnd 0.006041f
C285 output.n44 gnd 0.025987f
C286 output.n45 gnd 0.097665f
C287 output.n46 gnd 0.015803f
C288 output.n47 gnd 0.011243f
C289 output.n48 gnd 0.006041f
C290 output.n49 gnd 0.01428f
C291 output.n50 gnd 0.006397f
C292 output.n51 gnd 0.011243f
C293 output.n52 gnd 0.006041f
C294 output.n53 gnd 0.01428f
C295 output.n54 gnd 0.006397f
C296 output.n55 gnd 0.048111f
C297 output.t19 gnd 0.023274f
C298 output.n56 gnd 0.01071f
C299 output.n57 gnd 0.008435f
C300 output.n58 gnd 0.006041f
C301 output.n59 gnd 0.267512f
C302 output.n60 gnd 0.011243f
C303 output.n61 gnd 0.006041f
C304 output.n62 gnd 0.006397f
C305 output.n63 gnd 0.01428f
C306 output.n64 gnd 0.01428f
C307 output.n65 gnd 0.006397f
C308 output.n66 gnd 0.006041f
C309 output.n67 gnd 0.011243f
C310 output.n68 gnd 0.011243f
C311 output.n69 gnd 0.006041f
C312 output.n70 gnd 0.006397f
C313 output.n71 gnd 0.01428f
C314 output.n72 gnd 0.030913f
C315 output.n73 gnd 0.006397f
C316 output.n74 gnd 0.006041f
C317 output.n75 gnd 0.025987f
C318 output.n76 gnd 0.09306f
C319 output.n77 gnd 1.65264f
C320 output.n78 gnd 0.015803f
C321 output.n79 gnd 0.011243f
C322 output.n80 gnd 0.006041f
C323 output.n81 gnd 0.01428f
C324 output.n82 gnd 0.006397f
C325 output.n83 gnd 0.011243f
C326 output.n84 gnd 0.006041f
C327 output.n85 gnd 0.01428f
C328 output.n86 gnd 0.006397f
C329 output.n87 gnd 0.048111f
C330 output.t0 gnd 0.023274f
C331 output.n88 gnd 0.01071f
C332 output.n89 gnd 0.008435f
C333 output.n90 gnd 0.006041f
C334 output.n91 gnd 0.267512f
C335 output.n92 gnd 0.011243f
C336 output.n93 gnd 0.006041f
C337 output.n94 gnd 0.006397f
C338 output.n95 gnd 0.01428f
C339 output.n96 gnd 0.01428f
C340 output.n97 gnd 0.006397f
C341 output.n98 gnd 0.006041f
C342 output.n99 gnd 0.011243f
C343 output.n100 gnd 0.011243f
C344 output.n101 gnd 0.006041f
C345 output.n102 gnd 0.006397f
C346 output.n103 gnd 0.01428f
C347 output.n104 gnd 0.030913f
C348 output.n105 gnd 0.006397f
C349 output.n106 gnd 0.006041f
C350 output.n107 gnd 0.025987f
C351 output.n108 gnd 0.09306f
C352 output.n109 gnd 0.713089f
C353 output.n110 gnd 0.015803f
C354 output.n111 gnd 0.011243f
C355 output.n112 gnd 0.006041f
C356 output.n113 gnd 0.01428f
C357 output.n114 gnd 0.006397f
C358 output.n115 gnd 0.011243f
C359 output.n116 gnd 0.006041f
C360 output.n117 gnd 0.01428f
C361 output.n118 gnd 0.006397f
C362 output.n119 gnd 0.048111f
C363 output.t2 gnd 0.023274f
C364 output.n120 gnd 0.01071f
C365 output.n121 gnd 0.008435f
C366 output.n122 gnd 0.006041f
C367 output.n123 gnd 0.267512f
C368 output.n124 gnd 0.011243f
C369 output.n125 gnd 0.006041f
C370 output.n126 gnd 0.006397f
C371 output.n127 gnd 0.01428f
C372 output.n128 gnd 0.01428f
C373 output.n129 gnd 0.006397f
C374 output.n130 gnd 0.006041f
C375 output.n131 gnd 0.011243f
C376 output.n132 gnd 0.011243f
C377 output.n133 gnd 0.006041f
C378 output.n134 gnd 0.006397f
C379 output.n135 gnd 0.01428f
C380 output.n136 gnd 0.030913f
C381 output.n137 gnd 0.006397f
C382 output.n138 gnd 0.006041f
C383 output.n139 gnd 0.025987f
C384 output.n140 gnd 0.09306f
C385 output.n141 gnd 1.67353f
C386 diffpairibias.t27 gnd 0.090128f
C387 diffpairibias.t23 gnd 0.08996f
C388 diffpairibias.n0 gnd 0.105991f
C389 diffpairibias.t28 gnd 0.08996f
C390 diffpairibias.n1 gnd 0.051736f
C391 diffpairibias.t25 gnd 0.08996f
C392 diffpairibias.n2 gnd 0.051736f
C393 diffpairibias.t29 gnd 0.08996f
C394 diffpairibias.n3 gnd 0.041084f
C395 diffpairibias.t15 gnd 0.086371f
C396 diffpairibias.t1 gnd 0.085993f
C397 diffpairibias.n4 gnd 0.13579f
C398 diffpairibias.t11 gnd 0.085993f
C399 diffpairibias.n5 gnd 0.072463f
C400 diffpairibias.t13 gnd 0.085993f
C401 diffpairibias.n6 gnd 0.072463f
C402 diffpairibias.t7 gnd 0.085993f
C403 diffpairibias.n7 gnd 0.072463f
C404 diffpairibias.t3 gnd 0.085993f
C405 diffpairibias.n8 gnd 0.072463f
C406 diffpairibias.t17 gnd 0.085993f
C407 diffpairibias.n9 gnd 0.072463f
C408 diffpairibias.t5 gnd 0.085993f
C409 diffpairibias.n10 gnd 0.072463f
C410 diffpairibias.t19 gnd 0.085993f
C411 diffpairibias.n11 gnd 0.072463f
C412 diffpairibias.t9 gnd 0.085993f
C413 diffpairibias.n12 gnd 0.102883f
C414 diffpairibias.t14 gnd 0.086899f
C415 diffpairibias.t0 gnd 0.086748f
C416 diffpairibias.n13 gnd 0.094648f
C417 diffpairibias.t10 gnd 0.086748f
C418 diffpairibias.n14 gnd 0.052262f
C419 diffpairibias.t12 gnd 0.086748f
C420 diffpairibias.n15 gnd 0.052262f
C421 diffpairibias.t6 gnd 0.086748f
C422 diffpairibias.n16 gnd 0.052262f
C423 diffpairibias.t2 gnd 0.086748f
C424 diffpairibias.n17 gnd 0.052262f
C425 diffpairibias.t16 gnd 0.086748f
C426 diffpairibias.n18 gnd 0.052262f
C427 diffpairibias.t4 gnd 0.086748f
C428 diffpairibias.n19 gnd 0.052262f
C429 diffpairibias.t18 gnd 0.086748f
C430 diffpairibias.n20 gnd 0.052262f
C431 diffpairibias.t8 gnd 0.086748f
C432 diffpairibias.n21 gnd 0.061849f
C433 diffpairibias.n22 gnd 0.233513f
C434 diffpairibias.t20 gnd 0.08996f
C435 diffpairibias.n23 gnd 0.051747f
C436 diffpairibias.t26 gnd 0.08996f
C437 diffpairibias.n24 gnd 0.051736f
C438 diffpairibias.t22 gnd 0.08996f
C439 diffpairibias.n25 gnd 0.051736f
C440 diffpairibias.t21 gnd 0.08996f
C441 diffpairibias.n26 gnd 0.051736f
C442 diffpairibias.t24 gnd 0.08996f
C443 diffpairibias.n27 gnd 0.04729f
C444 diffpairibias.n28 gnd 0.047711f
C445 commonsourceibias.n0 gnd 0.010571f
C446 commonsourceibias.t92 gnd 0.160069f
C447 commonsourceibias.t106 gnd 0.148006f
C448 commonsourceibias.n1 gnd 0.006439f
C449 commonsourceibias.n2 gnd 0.007922f
C450 commonsourceibias.t119 gnd 0.148006f
C451 commonsourceibias.n3 gnd 0.008036f
C452 commonsourceibias.n4 gnd 0.007922f
C453 commonsourceibias.t84 gnd 0.148006f
C454 commonsourceibias.n5 gnd 0.059054f
C455 commonsourceibias.t100 gnd 0.148006f
C456 commonsourceibias.n6 gnd 0.006408f
C457 commonsourceibias.n7 gnd 0.007922f
C458 commonsourceibias.t114 gnd 0.148006f
C459 commonsourceibias.n8 gnd 0.007648f
C460 commonsourceibias.n9 gnd 0.007922f
C461 commonsourceibias.t80 gnd 0.148006f
C462 commonsourceibias.n10 gnd 0.059054f
C463 commonsourceibias.t76 gnd 0.148006f
C464 commonsourceibias.n11 gnd 0.006398f
C465 commonsourceibias.n12 gnd 0.010571f
C466 commonsourceibias.t60 gnd 0.160069f
C467 commonsourceibias.t14 gnd 0.148006f
C468 commonsourceibias.n13 gnd 0.006439f
C469 commonsourceibias.n14 gnd 0.007922f
C470 commonsourceibias.t38 gnd 0.148006f
C471 commonsourceibias.n15 gnd 0.008036f
C472 commonsourceibias.n16 gnd 0.007922f
C473 commonsourceibias.t4 gnd 0.148006f
C474 commonsourceibias.n17 gnd 0.059054f
C475 commonsourceibias.t28 gnd 0.148006f
C476 commonsourceibias.n18 gnd 0.006408f
C477 commonsourceibias.n19 gnd 0.007922f
C478 commonsourceibias.t62 gnd 0.148006f
C479 commonsourceibias.n20 gnd 0.007648f
C480 commonsourceibias.n21 gnd 0.007922f
C481 commonsourceibias.t18 gnd 0.148006f
C482 commonsourceibias.n22 gnd 0.059054f
C483 commonsourceibias.t26 gnd 0.148006f
C484 commonsourceibias.n23 gnd 0.006398f
C485 commonsourceibias.n24 gnd 0.007922f
C486 commonsourceibias.t6 gnd 0.148006f
C487 commonsourceibias.t32 gnd 0.148006f
C488 commonsourceibias.n25 gnd 0.059054f
C489 commonsourceibias.n26 gnd 0.007922f
C490 commonsourceibias.t42 gnd 0.148006f
C491 commonsourceibias.n27 gnd 0.059054f
C492 commonsourceibias.n28 gnd 0.007922f
C493 commonsourceibias.t20 gnd 0.148006f
C494 commonsourceibias.n29 gnd 0.059054f
C495 commonsourceibias.n30 gnd 0.007922f
C496 commonsourceibias.t30 gnd 0.148006f
C497 commonsourceibias.n31 gnd 0.009005f
C498 commonsourceibias.n32 gnd 0.007922f
C499 commonsourceibias.t56 gnd 0.148006f
C500 commonsourceibias.n33 gnd 0.010649f
C501 commonsourceibias.t16 gnd 0.164876f
C502 commonsourceibias.t12 gnd 0.148006f
C503 commonsourceibias.n34 gnd 0.065802f
C504 commonsourceibias.n35 gnd 0.070497f
C505 commonsourceibias.n36 gnd 0.03372f
C506 commonsourceibias.n37 gnd 0.007922f
C507 commonsourceibias.n38 gnd 0.006439f
C508 commonsourceibias.n39 gnd 0.010916f
C509 commonsourceibias.n40 gnd 0.059054f
C510 commonsourceibias.n41 gnd 0.010963f
C511 commonsourceibias.n42 gnd 0.007922f
C512 commonsourceibias.n43 gnd 0.007922f
C513 commonsourceibias.n44 gnd 0.007922f
C514 commonsourceibias.n45 gnd 0.008036f
C515 commonsourceibias.n46 gnd 0.059054f
C516 commonsourceibias.n47 gnd 0.009764f
C517 commonsourceibias.n48 gnd 0.010802f
C518 commonsourceibias.n49 gnd 0.007922f
C519 commonsourceibias.n50 gnd 0.007922f
C520 commonsourceibias.n51 gnd 0.010731f
C521 commonsourceibias.n52 gnd 0.006408f
C522 commonsourceibias.n53 gnd 0.010864f
C523 commonsourceibias.n54 gnd 0.007922f
C524 commonsourceibias.n55 gnd 0.007922f
C525 commonsourceibias.n56 gnd 0.010931f
C526 commonsourceibias.n57 gnd 0.009425f
C527 commonsourceibias.n58 gnd 0.007648f
C528 commonsourceibias.n59 gnd 0.007922f
C529 commonsourceibias.n60 gnd 0.007922f
C530 commonsourceibias.n61 gnd 0.00969f
C531 commonsourceibias.n62 gnd 0.010876f
C532 commonsourceibias.n63 gnd 0.059054f
C533 commonsourceibias.n64 gnd 0.010803f
C534 commonsourceibias.n65 gnd 0.007922f
C535 commonsourceibias.n66 gnd 0.007922f
C536 commonsourceibias.n67 gnd 0.007922f
C537 commonsourceibias.n68 gnd 0.010803f
C538 commonsourceibias.n69 gnd 0.059054f
C539 commonsourceibias.n70 gnd 0.010876f
C540 commonsourceibias.n71 gnd 0.00969f
C541 commonsourceibias.n72 gnd 0.007922f
C542 commonsourceibias.n73 gnd 0.007922f
C543 commonsourceibias.n74 gnd 0.007922f
C544 commonsourceibias.n75 gnd 0.009425f
C545 commonsourceibias.n76 gnd 0.010931f
C546 commonsourceibias.n77 gnd 0.059054f
C547 commonsourceibias.n78 gnd 0.010864f
C548 commonsourceibias.n79 gnd 0.007922f
C549 commonsourceibias.n80 gnd 0.007922f
C550 commonsourceibias.n81 gnd 0.007922f
C551 commonsourceibias.n82 gnd 0.010731f
C552 commonsourceibias.n83 gnd 0.059054f
C553 commonsourceibias.n84 gnd 0.010802f
C554 commonsourceibias.n85 gnd 0.009764f
C555 commonsourceibias.n86 gnd 0.007922f
C556 commonsourceibias.n87 gnd 0.007922f
C557 commonsourceibias.n88 gnd 0.007922f
C558 commonsourceibias.n89 gnd 0.009005f
C559 commonsourceibias.n90 gnd 0.010963f
C560 commonsourceibias.n91 gnd 0.059054f
C561 commonsourceibias.n92 gnd 0.010916f
C562 commonsourceibias.n93 gnd 0.007922f
C563 commonsourceibias.n94 gnd 0.007922f
C564 commonsourceibias.n95 gnd 0.007922f
C565 commonsourceibias.n96 gnd 0.010649f
C566 commonsourceibias.n97 gnd 0.059054f
C567 commonsourceibias.n98 gnd 0.010674f
C568 commonsourceibias.n99 gnd 0.071211f
C569 commonsourceibias.n100 gnd 0.079625f
C570 commonsourceibias.t61 gnd 0.017095f
C571 commonsourceibias.t15 gnd 0.017095f
C572 commonsourceibias.n101 gnd 0.151055f
C573 commonsourceibias.n102 gnd 0.130846f
C574 commonsourceibias.t39 gnd 0.017095f
C575 commonsourceibias.t5 gnd 0.017095f
C576 commonsourceibias.n103 gnd 0.151055f
C577 commonsourceibias.n104 gnd 0.069385f
C578 commonsourceibias.t29 gnd 0.017095f
C579 commonsourceibias.t63 gnd 0.017095f
C580 commonsourceibias.n105 gnd 0.151055f
C581 commonsourceibias.n106 gnd 0.069385f
C582 commonsourceibias.t19 gnd 0.017095f
C583 commonsourceibias.t27 gnd 0.017095f
C584 commonsourceibias.n107 gnd 0.151055f
C585 commonsourceibias.n108 gnd 0.057968f
C586 commonsourceibias.t13 gnd 0.017095f
C587 commonsourceibias.t17 gnd 0.017095f
C588 commonsourceibias.n109 gnd 0.15156f
C589 commonsourceibias.t31 gnd 0.017095f
C590 commonsourceibias.t57 gnd 0.017095f
C591 commonsourceibias.n110 gnd 0.151055f
C592 commonsourceibias.n111 gnd 0.140755f
C593 commonsourceibias.t43 gnd 0.017095f
C594 commonsourceibias.t21 gnd 0.017095f
C595 commonsourceibias.n112 gnd 0.151055f
C596 commonsourceibias.n113 gnd 0.069385f
C597 commonsourceibias.t7 gnd 0.017095f
C598 commonsourceibias.t33 gnd 0.017095f
C599 commonsourceibias.n114 gnd 0.151055f
C600 commonsourceibias.n115 gnd 0.057968f
C601 commonsourceibias.n116 gnd 0.070193f
C602 commonsourceibias.n117 gnd 0.007922f
C603 commonsourceibias.t105 gnd 0.148006f
C604 commonsourceibias.t121 gnd 0.148006f
C605 commonsourceibias.n118 gnd 0.059054f
C606 commonsourceibias.n119 gnd 0.007922f
C607 commonsourceibias.t71 gnd 0.148006f
C608 commonsourceibias.n120 gnd 0.059054f
C609 commonsourceibias.n121 gnd 0.007922f
C610 commonsourceibias.t99 gnd 0.148006f
C611 commonsourceibias.n122 gnd 0.059054f
C612 commonsourceibias.n123 gnd 0.007922f
C613 commonsourceibias.t95 gnd 0.148006f
C614 commonsourceibias.n124 gnd 0.009005f
C615 commonsourceibias.n125 gnd 0.007922f
C616 commonsourceibias.t109 gnd 0.148006f
C617 commonsourceibias.n126 gnd 0.010649f
C618 commonsourceibias.t85 gnd 0.164876f
C619 commonsourceibias.t89 gnd 0.148006f
C620 commonsourceibias.n127 gnd 0.065802f
C621 commonsourceibias.n128 gnd 0.070497f
C622 commonsourceibias.n129 gnd 0.03372f
C623 commonsourceibias.n130 gnd 0.007922f
C624 commonsourceibias.n131 gnd 0.006439f
C625 commonsourceibias.n132 gnd 0.010916f
C626 commonsourceibias.n133 gnd 0.059054f
C627 commonsourceibias.n134 gnd 0.010963f
C628 commonsourceibias.n135 gnd 0.007922f
C629 commonsourceibias.n136 gnd 0.007922f
C630 commonsourceibias.n137 gnd 0.007922f
C631 commonsourceibias.n138 gnd 0.008036f
C632 commonsourceibias.n139 gnd 0.059054f
C633 commonsourceibias.n140 gnd 0.009764f
C634 commonsourceibias.n141 gnd 0.010802f
C635 commonsourceibias.n142 gnd 0.007922f
C636 commonsourceibias.n143 gnd 0.007922f
C637 commonsourceibias.n144 gnd 0.010731f
C638 commonsourceibias.n145 gnd 0.006408f
C639 commonsourceibias.n146 gnd 0.010864f
C640 commonsourceibias.n147 gnd 0.007922f
C641 commonsourceibias.n148 gnd 0.007922f
C642 commonsourceibias.n149 gnd 0.010931f
C643 commonsourceibias.n150 gnd 0.009425f
C644 commonsourceibias.n151 gnd 0.007648f
C645 commonsourceibias.n152 gnd 0.007922f
C646 commonsourceibias.n153 gnd 0.007922f
C647 commonsourceibias.n154 gnd 0.00969f
C648 commonsourceibias.n155 gnd 0.010876f
C649 commonsourceibias.n156 gnd 0.059054f
C650 commonsourceibias.n157 gnd 0.010803f
C651 commonsourceibias.n158 gnd 0.007884f
C652 commonsourceibias.n159 gnd 0.057266f
C653 commonsourceibias.n160 gnd 0.007884f
C654 commonsourceibias.n161 gnd 0.010803f
C655 commonsourceibias.n162 gnd 0.059054f
C656 commonsourceibias.n163 gnd 0.010876f
C657 commonsourceibias.n164 gnd 0.00969f
C658 commonsourceibias.n165 gnd 0.007922f
C659 commonsourceibias.n166 gnd 0.007922f
C660 commonsourceibias.n167 gnd 0.007922f
C661 commonsourceibias.n168 gnd 0.009425f
C662 commonsourceibias.n169 gnd 0.010931f
C663 commonsourceibias.n170 gnd 0.059054f
C664 commonsourceibias.n171 gnd 0.010864f
C665 commonsourceibias.n172 gnd 0.007922f
C666 commonsourceibias.n173 gnd 0.007922f
C667 commonsourceibias.n174 gnd 0.007922f
C668 commonsourceibias.n175 gnd 0.010731f
C669 commonsourceibias.n176 gnd 0.059054f
C670 commonsourceibias.n177 gnd 0.010802f
C671 commonsourceibias.n178 gnd 0.009764f
C672 commonsourceibias.n179 gnd 0.007922f
C673 commonsourceibias.n180 gnd 0.007922f
C674 commonsourceibias.n181 gnd 0.007922f
C675 commonsourceibias.n182 gnd 0.009005f
C676 commonsourceibias.n183 gnd 0.010963f
C677 commonsourceibias.n184 gnd 0.059054f
C678 commonsourceibias.n185 gnd 0.010916f
C679 commonsourceibias.n186 gnd 0.007922f
C680 commonsourceibias.n187 gnd 0.007922f
C681 commonsourceibias.n188 gnd 0.007922f
C682 commonsourceibias.n189 gnd 0.010649f
C683 commonsourceibias.n190 gnd 0.059054f
C684 commonsourceibias.n191 gnd 0.010674f
C685 commonsourceibias.n192 gnd 0.071211f
C686 commonsourceibias.n193 gnd 0.047027f
C687 commonsourceibias.n194 gnd 0.010571f
C688 commonsourceibias.t94 gnd 0.148006f
C689 commonsourceibias.n195 gnd 0.006439f
C690 commonsourceibias.n196 gnd 0.007922f
C691 commonsourceibias.t107 gnd 0.148006f
C692 commonsourceibias.n197 gnd 0.008036f
C693 commonsourceibias.n198 gnd 0.007922f
C694 commonsourceibias.t74 gnd 0.148006f
C695 commonsourceibias.n199 gnd 0.059054f
C696 commonsourceibias.t87 gnd 0.148006f
C697 commonsourceibias.n200 gnd 0.006408f
C698 commonsourceibias.n201 gnd 0.007922f
C699 commonsourceibias.t101 gnd 0.148006f
C700 commonsourceibias.n202 gnd 0.007648f
C701 commonsourceibias.n203 gnd 0.007922f
C702 commonsourceibias.t70 gnd 0.148006f
C703 commonsourceibias.n204 gnd 0.059054f
C704 commonsourceibias.t67 gnd 0.148006f
C705 commonsourceibias.n205 gnd 0.006398f
C706 commonsourceibias.n206 gnd 0.007922f
C707 commonsourceibias.t93 gnd 0.148006f
C708 commonsourceibias.t108 gnd 0.148006f
C709 commonsourceibias.n207 gnd 0.059054f
C710 commonsourceibias.n208 gnd 0.007922f
C711 commonsourceibias.t127 gnd 0.148006f
C712 commonsourceibias.n209 gnd 0.059054f
C713 commonsourceibias.n210 gnd 0.007922f
C714 commonsourceibias.t86 gnd 0.148006f
C715 commonsourceibias.n211 gnd 0.059054f
C716 commonsourceibias.n212 gnd 0.007922f
C717 commonsourceibias.t82 gnd 0.148006f
C718 commonsourceibias.n213 gnd 0.009005f
C719 commonsourceibias.n214 gnd 0.007922f
C720 commonsourceibias.t96 gnd 0.148006f
C721 commonsourceibias.n215 gnd 0.010649f
C722 commonsourceibias.t75 gnd 0.164876f
C723 commonsourceibias.t77 gnd 0.148006f
C724 commonsourceibias.n216 gnd 0.065802f
C725 commonsourceibias.n217 gnd 0.070497f
C726 commonsourceibias.n218 gnd 0.03372f
C727 commonsourceibias.n219 gnd 0.007922f
C728 commonsourceibias.n220 gnd 0.006439f
C729 commonsourceibias.n221 gnd 0.010916f
C730 commonsourceibias.n222 gnd 0.059054f
C731 commonsourceibias.n223 gnd 0.010963f
C732 commonsourceibias.n224 gnd 0.007922f
C733 commonsourceibias.n225 gnd 0.007922f
C734 commonsourceibias.n226 gnd 0.007922f
C735 commonsourceibias.n227 gnd 0.008036f
C736 commonsourceibias.n228 gnd 0.059054f
C737 commonsourceibias.n229 gnd 0.009764f
C738 commonsourceibias.n230 gnd 0.010802f
C739 commonsourceibias.n231 gnd 0.007922f
C740 commonsourceibias.n232 gnd 0.007922f
C741 commonsourceibias.n233 gnd 0.010731f
C742 commonsourceibias.n234 gnd 0.006408f
C743 commonsourceibias.n235 gnd 0.010864f
C744 commonsourceibias.n236 gnd 0.007922f
C745 commonsourceibias.n237 gnd 0.007922f
C746 commonsourceibias.n238 gnd 0.010931f
C747 commonsourceibias.n239 gnd 0.009425f
C748 commonsourceibias.n240 gnd 0.007648f
C749 commonsourceibias.n241 gnd 0.007922f
C750 commonsourceibias.n242 gnd 0.007922f
C751 commonsourceibias.n243 gnd 0.00969f
C752 commonsourceibias.n244 gnd 0.010876f
C753 commonsourceibias.n245 gnd 0.059054f
C754 commonsourceibias.n246 gnd 0.010803f
C755 commonsourceibias.n247 gnd 0.007922f
C756 commonsourceibias.n248 gnd 0.007922f
C757 commonsourceibias.n249 gnd 0.007922f
C758 commonsourceibias.n250 gnd 0.010803f
C759 commonsourceibias.n251 gnd 0.059054f
C760 commonsourceibias.n252 gnd 0.010876f
C761 commonsourceibias.n253 gnd 0.00969f
C762 commonsourceibias.n254 gnd 0.007922f
C763 commonsourceibias.n255 gnd 0.007922f
C764 commonsourceibias.n256 gnd 0.007922f
C765 commonsourceibias.n257 gnd 0.009425f
C766 commonsourceibias.n258 gnd 0.010931f
C767 commonsourceibias.n259 gnd 0.059054f
C768 commonsourceibias.n260 gnd 0.010864f
C769 commonsourceibias.n261 gnd 0.007922f
C770 commonsourceibias.n262 gnd 0.007922f
C771 commonsourceibias.n263 gnd 0.007922f
C772 commonsourceibias.n264 gnd 0.010731f
C773 commonsourceibias.n265 gnd 0.059054f
C774 commonsourceibias.n266 gnd 0.010802f
C775 commonsourceibias.n267 gnd 0.009764f
C776 commonsourceibias.n268 gnd 0.007922f
C777 commonsourceibias.n269 gnd 0.007922f
C778 commonsourceibias.n270 gnd 0.007922f
C779 commonsourceibias.n271 gnd 0.009005f
C780 commonsourceibias.n272 gnd 0.010963f
C781 commonsourceibias.n273 gnd 0.059054f
C782 commonsourceibias.n274 gnd 0.010916f
C783 commonsourceibias.n275 gnd 0.007922f
C784 commonsourceibias.n276 gnd 0.007922f
C785 commonsourceibias.n277 gnd 0.007922f
C786 commonsourceibias.n278 gnd 0.010649f
C787 commonsourceibias.n279 gnd 0.059054f
C788 commonsourceibias.n280 gnd 0.010674f
C789 commonsourceibias.t81 gnd 0.160069f
C790 commonsourceibias.n281 gnd 0.071211f
C791 commonsourceibias.n282 gnd 0.025411f
C792 commonsourceibias.n283 gnd 0.458519f
C793 commonsourceibias.n284 gnd 0.010571f
C794 commonsourceibias.t110 gnd 0.160069f
C795 commonsourceibias.t123 gnd 0.148006f
C796 commonsourceibias.n285 gnd 0.006439f
C797 commonsourceibias.n286 gnd 0.007922f
C798 commonsourceibias.t68 gnd 0.148006f
C799 commonsourceibias.n287 gnd 0.008036f
C800 commonsourceibias.n288 gnd 0.007922f
C801 commonsourceibias.t117 gnd 0.148006f
C802 commonsourceibias.n289 gnd 0.006408f
C803 commonsourceibias.n290 gnd 0.007922f
C804 commonsourceibias.t64 gnd 0.148006f
C805 commonsourceibias.n291 gnd 0.007648f
C806 commonsourceibias.n292 gnd 0.007922f
C807 commonsourceibias.t90 gnd 0.148006f
C808 commonsourceibias.n293 gnd 0.006398f
C809 commonsourceibias.n294 gnd 0.007922f
C810 commonsourceibias.t122 gnd 0.148006f
C811 commonsourceibias.t69 gnd 0.148006f
C812 commonsourceibias.n295 gnd 0.059054f
C813 commonsourceibias.n296 gnd 0.007922f
C814 commonsourceibias.t66 gnd 0.148006f
C815 commonsourceibias.n297 gnd 0.059054f
C816 commonsourceibias.n298 gnd 0.007922f
C817 commonsourceibias.t116 gnd 0.148006f
C818 commonsourceibias.n299 gnd 0.059054f
C819 commonsourceibias.n300 gnd 0.007922f
C820 commonsourceibias.t113 gnd 0.148006f
C821 commonsourceibias.n301 gnd 0.009005f
C822 commonsourceibias.n302 gnd 0.007922f
C823 commonsourceibias.t126 gnd 0.148006f
C824 commonsourceibias.n303 gnd 0.010649f
C825 commonsourceibias.t91 gnd 0.164876f
C826 commonsourceibias.t83 gnd 0.148006f
C827 commonsourceibias.n304 gnd 0.065802f
C828 commonsourceibias.n305 gnd 0.070497f
C829 commonsourceibias.n306 gnd 0.03372f
C830 commonsourceibias.n307 gnd 0.007922f
C831 commonsourceibias.n308 gnd 0.006439f
C832 commonsourceibias.n309 gnd 0.010916f
C833 commonsourceibias.n310 gnd 0.059054f
C834 commonsourceibias.n311 gnd 0.010963f
C835 commonsourceibias.n312 gnd 0.007922f
C836 commonsourceibias.n313 gnd 0.007922f
C837 commonsourceibias.n314 gnd 0.007922f
C838 commonsourceibias.n315 gnd 0.008036f
C839 commonsourceibias.n316 gnd 0.059054f
C840 commonsourceibias.n317 gnd 0.009764f
C841 commonsourceibias.n318 gnd 0.010802f
C842 commonsourceibias.n319 gnd 0.007922f
C843 commonsourceibias.n320 gnd 0.007922f
C844 commonsourceibias.n321 gnd 0.010731f
C845 commonsourceibias.n322 gnd 0.006408f
C846 commonsourceibias.n323 gnd 0.010864f
C847 commonsourceibias.n324 gnd 0.007922f
C848 commonsourceibias.n325 gnd 0.007922f
C849 commonsourceibias.n326 gnd 0.010931f
C850 commonsourceibias.n327 gnd 0.009425f
C851 commonsourceibias.n328 gnd 0.007648f
C852 commonsourceibias.n329 gnd 0.007922f
C853 commonsourceibias.n330 gnd 0.007922f
C854 commonsourceibias.n331 gnd 0.00969f
C855 commonsourceibias.n332 gnd 0.010876f
C856 commonsourceibias.n333 gnd 0.059054f
C857 commonsourceibias.n334 gnd 0.010803f
C858 commonsourceibias.n335 gnd 0.007884f
C859 commonsourceibias.t55 gnd 0.017095f
C860 commonsourceibias.t53 gnd 0.017095f
C861 commonsourceibias.n336 gnd 0.15156f
C862 commonsourceibias.t3 gnd 0.017095f
C863 commonsourceibias.t49 gnd 0.017095f
C864 commonsourceibias.n337 gnd 0.151055f
C865 commonsourceibias.n338 gnd 0.140755f
C866 commonsourceibias.t41 gnd 0.017095f
C867 commonsourceibias.t59 gnd 0.017095f
C868 commonsourceibias.n339 gnd 0.151055f
C869 commonsourceibias.n340 gnd 0.069385f
C870 commonsourceibias.t51 gnd 0.017095f
C871 commonsourceibias.t25 gnd 0.017095f
C872 commonsourceibias.n341 gnd 0.151055f
C873 commonsourceibias.n342 gnd 0.057968f
C874 commonsourceibias.n343 gnd 0.010571f
C875 commonsourceibias.t34 gnd 0.148006f
C876 commonsourceibias.n344 gnd 0.006439f
C877 commonsourceibias.n345 gnd 0.007922f
C878 commonsourceibias.t0 gnd 0.148006f
C879 commonsourceibias.n346 gnd 0.008036f
C880 commonsourceibias.n347 gnd 0.007922f
C881 commonsourceibias.t46 gnd 0.148006f
C882 commonsourceibias.n348 gnd 0.006408f
C883 commonsourceibias.n349 gnd 0.007922f
C884 commonsourceibias.t10 gnd 0.148006f
C885 commonsourceibias.n350 gnd 0.007648f
C886 commonsourceibias.n351 gnd 0.007922f
C887 commonsourceibias.t44 gnd 0.148006f
C888 commonsourceibias.n352 gnd 0.006398f
C889 commonsourceibias.n353 gnd 0.007922f
C890 commonsourceibias.t24 gnd 0.148006f
C891 commonsourceibias.t50 gnd 0.148006f
C892 commonsourceibias.n354 gnd 0.059054f
C893 commonsourceibias.n355 gnd 0.007922f
C894 commonsourceibias.t58 gnd 0.148006f
C895 commonsourceibias.n356 gnd 0.059054f
C896 commonsourceibias.n357 gnd 0.007922f
C897 commonsourceibias.t40 gnd 0.148006f
C898 commonsourceibias.n358 gnd 0.059054f
C899 commonsourceibias.n359 gnd 0.007922f
C900 commonsourceibias.t48 gnd 0.148006f
C901 commonsourceibias.n360 gnd 0.009005f
C902 commonsourceibias.n361 gnd 0.007922f
C903 commonsourceibias.t2 gnd 0.148006f
C904 commonsourceibias.n362 gnd 0.010649f
C905 commonsourceibias.t54 gnd 0.164876f
C906 commonsourceibias.t52 gnd 0.148006f
C907 commonsourceibias.n363 gnd 0.065802f
C908 commonsourceibias.n364 gnd 0.070497f
C909 commonsourceibias.n365 gnd 0.03372f
C910 commonsourceibias.n366 gnd 0.007922f
C911 commonsourceibias.n367 gnd 0.006439f
C912 commonsourceibias.n368 gnd 0.010916f
C913 commonsourceibias.n369 gnd 0.059054f
C914 commonsourceibias.n370 gnd 0.010963f
C915 commonsourceibias.n371 gnd 0.007922f
C916 commonsourceibias.n372 gnd 0.007922f
C917 commonsourceibias.n373 gnd 0.007922f
C918 commonsourceibias.n374 gnd 0.008036f
C919 commonsourceibias.n375 gnd 0.059054f
C920 commonsourceibias.n376 gnd 0.009764f
C921 commonsourceibias.n377 gnd 0.010802f
C922 commonsourceibias.n378 gnd 0.007922f
C923 commonsourceibias.n379 gnd 0.007922f
C924 commonsourceibias.n380 gnd 0.010731f
C925 commonsourceibias.n381 gnd 0.006408f
C926 commonsourceibias.n382 gnd 0.010864f
C927 commonsourceibias.n383 gnd 0.007922f
C928 commonsourceibias.n384 gnd 0.007922f
C929 commonsourceibias.n385 gnd 0.010931f
C930 commonsourceibias.n386 gnd 0.009425f
C931 commonsourceibias.n387 gnd 0.007648f
C932 commonsourceibias.n388 gnd 0.007922f
C933 commonsourceibias.n389 gnd 0.007922f
C934 commonsourceibias.n390 gnd 0.00969f
C935 commonsourceibias.n391 gnd 0.010876f
C936 commonsourceibias.n392 gnd 0.059054f
C937 commonsourceibias.n393 gnd 0.010803f
C938 commonsourceibias.n394 gnd 0.007922f
C939 commonsourceibias.n395 gnd 0.007922f
C940 commonsourceibias.n396 gnd 0.007922f
C941 commonsourceibias.n397 gnd 0.010803f
C942 commonsourceibias.n398 gnd 0.059054f
C943 commonsourceibias.n399 gnd 0.010876f
C944 commonsourceibias.t36 gnd 0.148006f
C945 commonsourceibias.n400 gnd 0.059054f
C946 commonsourceibias.n401 gnd 0.00969f
C947 commonsourceibias.n402 gnd 0.007922f
C948 commonsourceibias.n403 gnd 0.007922f
C949 commonsourceibias.n404 gnd 0.007922f
C950 commonsourceibias.n405 gnd 0.009425f
C951 commonsourceibias.n406 gnd 0.010931f
C952 commonsourceibias.n407 gnd 0.059054f
C953 commonsourceibias.n408 gnd 0.010864f
C954 commonsourceibias.n409 gnd 0.007922f
C955 commonsourceibias.n410 gnd 0.007922f
C956 commonsourceibias.n411 gnd 0.007922f
C957 commonsourceibias.n412 gnd 0.010731f
C958 commonsourceibias.n413 gnd 0.059054f
C959 commonsourceibias.n414 gnd 0.010802f
C960 commonsourceibias.t22 gnd 0.148006f
C961 commonsourceibias.n415 gnd 0.059054f
C962 commonsourceibias.n416 gnd 0.009764f
C963 commonsourceibias.n417 gnd 0.007922f
C964 commonsourceibias.n418 gnd 0.007922f
C965 commonsourceibias.n419 gnd 0.007922f
C966 commonsourceibias.n420 gnd 0.009005f
C967 commonsourceibias.n421 gnd 0.010963f
C968 commonsourceibias.n422 gnd 0.059054f
C969 commonsourceibias.n423 gnd 0.010916f
C970 commonsourceibias.n424 gnd 0.007922f
C971 commonsourceibias.n425 gnd 0.007922f
C972 commonsourceibias.n426 gnd 0.007922f
C973 commonsourceibias.n427 gnd 0.010649f
C974 commonsourceibias.n428 gnd 0.059054f
C975 commonsourceibias.n429 gnd 0.010674f
C976 commonsourceibias.t8 gnd 0.160069f
C977 commonsourceibias.n430 gnd 0.071211f
C978 commonsourceibias.n431 gnd 0.079625f
C979 commonsourceibias.t35 gnd 0.017095f
C980 commonsourceibias.t9 gnd 0.017095f
C981 commonsourceibias.n432 gnd 0.151055f
C982 commonsourceibias.n433 gnd 0.130846f
C983 commonsourceibias.t23 gnd 0.017095f
C984 commonsourceibias.t1 gnd 0.017095f
C985 commonsourceibias.n434 gnd 0.151055f
C986 commonsourceibias.n435 gnd 0.069385f
C987 commonsourceibias.t11 gnd 0.017095f
C988 commonsourceibias.t47 gnd 0.017095f
C989 commonsourceibias.n436 gnd 0.151055f
C990 commonsourceibias.n437 gnd 0.069385f
C991 commonsourceibias.t45 gnd 0.017095f
C992 commonsourceibias.t37 gnd 0.017095f
C993 commonsourceibias.n438 gnd 0.151055f
C994 commonsourceibias.n439 gnd 0.057968f
C995 commonsourceibias.n440 gnd 0.070193f
C996 commonsourceibias.n441 gnd 0.057266f
C997 commonsourceibias.n442 gnd 0.007884f
C998 commonsourceibias.n443 gnd 0.010803f
C999 commonsourceibias.n444 gnd 0.059054f
C1000 commonsourceibias.n445 gnd 0.010876f
C1001 commonsourceibias.t72 gnd 0.148006f
C1002 commonsourceibias.n446 gnd 0.059054f
C1003 commonsourceibias.n447 gnd 0.00969f
C1004 commonsourceibias.n448 gnd 0.007922f
C1005 commonsourceibias.n449 gnd 0.007922f
C1006 commonsourceibias.n450 gnd 0.007922f
C1007 commonsourceibias.n451 gnd 0.009425f
C1008 commonsourceibias.n452 gnd 0.010931f
C1009 commonsourceibias.n453 gnd 0.059054f
C1010 commonsourceibias.n454 gnd 0.010864f
C1011 commonsourceibias.n455 gnd 0.007922f
C1012 commonsourceibias.n456 gnd 0.007922f
C1013 commonsourceibias.n457 gnd 0.007922f
C1014 commonsourceibias.n458 gnd 0.010731f
C1015 commonsourceibias.n459 gnd 0.059054f
C1016 commonsourceibias.n460 gnd 0.010802f
C1017 commonsourceibias.t102 gnd 0.148006f
C1018 commonsourceibias.n461 gnd 0.059054f
C1019 commonsourceibias.n462 gnd 0.009764f
C1020 commonsourceibias.n463 gnd 0.007922f
C1021 commonsourceibias.n464 gnd 0.007922f
C1022 commonsourceibias.n465 gnd 0.007922f
C1023 commonsourceibias.n466 gnd 0.009005f
C1024 commonsourceibias.n467 gnd 0.010963f
C1025 commonsourceibias.n468 gnd 0.059054f
C1026 commonsourceibias.n469 gnd 0.010916f
C1027 commonsourceibias.n470 gnd 0.007922f
C1028 commonsourceibias.n471 gnd 0.007922f
C1029 commonsourceibias.n472 gnd 0.007922f
C1030 commonsourceibias.n473 gnd 0.010649f
C1031 commonsourceibias.n474 gnd 0.059054f
C1032 commonsourceibias.n475 gnd 0.010674f
C1033 commonsourceibias.n476 gnd 0.071211f
C1034 commonsourceibias.n477 gnd 0.047027f
C1035 commonsourceibias.n478 gnd 0.010571f
C1036 commonsourceibias.t112 gnd 0.148006f
C1037 commonsourceibias.n479 gnd 0.006439f
C1038 commonsourceibias.n480 gnd 0.007922f
C1039 commonsourceibias.t124 gnd 0.148006f
C1040 commonsourceibias.n481 gnd 0.008036f
C1041 commonsourceibias.n482 gnd 0.007922f
C1042 commonsourceibias.t104 gnd 0.148006f
C1043 commonsourceibias.n483 gnd 0.006408f
C1044 commonsourceibias.n484 gnd 0.007922f
C1045 commonsourceibias.t118 gnd 0.148006f
C1046 commonsourceibias.n485 gnd 0.007648f
C1047 commonsourceibias.n486 gnd 0.007922f
C1048 commonsourceibias.t79 gnd 0.148006f
C1049 commonsourceibias.n487 gnd 0.006398f
C1050 commonsourceibias.n488 gnd 0.007922f
C1051 commonsourceibias.t111 gnd 0.148006f
C1052 commonsourceibias.t125 gnd 0.148006f
C1053 commonsourceibias.n489 gnd 0.059054f
C1054 commonsourceibias.n490 gnd 0.007922f
C1055 commonsourceibias.t120 gnd 0.148006f
C1056 commonsourceibias.n491 gnd 0.059054f
C1057 commonsourceibias.n492 gnd 0.007922f
C1058 commonsourceibias.t103 gnd 0.148006f
C1059 commonsourceibias.n493 gnd 0.059054f
C1060 commonsourceibias.n494 gnd 0.007922f
C1061 commonsourceibias.t98 gnd 0.148006f
C1062 commonsourceibias.n495 gnd 0.009005f
C1063 commonsourceibias.n496 gnd 0.007922f
C1064 commonsourceibias.t115 gnd 0.148006f
C1065 commonsourceibias.n497 gnd 0.010649f
C1066 commonsourceibias.t78 gnd 0.164876f
C1067 commonsourceibias.t73 gnd 0.148006f
C1068 commonsourceibias.n498 gnd 0.065802f
C1069 commonsourceibias.n499 gnd 0.070497f
C1070 commonsourceibias.n500 gnd 0.03372f
C1071 commonsourceibias.n501 gnd 0.007922f
C1072 commonsourceibias.n502 gnd 0.006439f
C1073 commonsourceibias.n503 gnd 0.010916f
C1074 commonsourceibias.n504 gnd 0.059054f
C1075 commonsourceibias.n505 gnd 0.010963f
C1076 commonsourceibias.n506 gnd 0.007922f
C1077 commonsourceibias.n507 gnd 0.007922f
C1078 commonsourceibias.n508 gnd 0.007922f
C1079 commonsourceibias.n509 gnd 0.008036f
C1080 commonsourceibias.n510 gnd 0.059054f
C1081 commonsourceibias.n511 gnd 0.009764f
C1082 commonsourceibias.n512 gnd 0.010802f
C1083 commonsourceibias.n513 gnd 0.007922f
C1084 commonsourceibias.n514 gnd 0.007922f
C1085 commonsourceibias.n515 gnd 0.010731f
C1086 commonsourceibias.n516 gnd 0.006408f
C1087 commonsourceibias.n517 gnd 0.010864f
C1088 commonsourceibias.n518 gnd 0.007922f
C1089 commonsourceibias.n519 gnd 0.007922f
C1090 commonsourceibias.n520 gnd 0.010931f
C1091 commonsourceibias.n521 gnd 0.009425f
C1092 commonsourceibias.n522 gnd 0.007648f
C1093 commonsourceibias.n523 gnd 0.007922f
C1094 commonsourceibias.n524 gnd 0.007922f
C1095 commonsourceibias.n525 gnd 0.00969f
C1096 commonsourceibias.n526 gnd 0.010876f
C1097 commonsourceibias.n527 gnd 0.059054f
C1098 commonsourceibias.n528 gnd 0.010803f
C1099 commonsourceibias.n529 gnd 0.007922f
C1100 commonsourceibias.n530 gnd 0.007922f
C1101 commonsourceibias.n531 gnd 0.007922f
C1102 commonsourceibias.n532 gnd 0.010803f
C1103 commonsourceibias.n533 gnd 0.059054f
C1104 commonsourceibias.n534 gnd 0.010876f
C1105 commonsourceibias.t65 gnd 0.148006f
C1106 commonsourceibias.n535 gnd 0.059054f
C1107 commonsourceibias.n536 gnd 0.00969f
C1108 commonsourceibias.n537 gnd 0.007922f
C1109 commonsourceibias.n538 gnd 0.007922f
C1110 commonsourceibias.n539 gnd 0.007922f
C1111 commonsourceibias.n540 gnd 0.009425f
C1112 commonsourceibias.n541 gnd 0.010931f
C1113 commonsourceibias.n542 gnd 0.059054f
C1114 commonsourceibias.n543 gnd 0.010864f
C1115 commonsourceibias.n544 gnd 0.007922f
C1116 commonsourceibias.n545 gnd 0.007922f
C1117 commonsourceibias.n546 gnd 0.007922f
C1118 commonsourceibias.n547 gnd 0.010731f
C1119 commonsourceibias.n548 gnd 0.059054f
C1120 commonsourceibias.n549 gnd 0.010802f
C1121 commonsourceibias.t88 gnd 0.148006f
C1122 commonsourceibias.n550 gnd 0.059054f
C1123 commonsourceibias.n551 gnd 0.009764f
C1124 commonsourceibias.n552 gnd 0.007922f
C1125 commonsourceibias.n553 gnd 0.007922f
C1126 commonsourceibias.n554 gnd 0.007922f
C1127 commonsourceibias.n555 gnd 0.009005f
C1128 commonsourceibias.n556 gnd 0.010963f
C1129 commonsourceibias.n557 gnd 0.059054f
C1130 commonsourceibias.n558 gnd 0.010916f
C1131 commonsourceibias.n559 gnd 0.007922f
C1132 commonsourceibias.n560 gnd 0.007922f
C1133 commonsourceibias.n561 gnd 0.007922f
C1134 commonsourceibias.n562 gnd 0.010649f
C1135 commonsourceibias.n563 gnd 0.059054f
C1136 commonsourceibias.n564 gnd 0.010674f
C1137 commonsourceibias.t97 gnd 0.160069f
C1138 commonsourceibias.n565 gnd 0.071211f
C1139 commonsourceibias.n566 gnd 0.025411f
C1140 commonsourceibias.n567 gnd 0.219034f
C1141 commonsourceibias.n568 gnd 4.63083f
C1142 minus.n0 gnd 0.031797f
C1143 minus.n1 gnd 0.007215f
C1144 minus.n2 gnd 0.031797f
C1145 minus.n3 gnd 0.007215f
C1146 minus.n4 gnd 0.031797f
C1147 minus.n5 gnd 0.007215f
C1148 minus.n6 gnd 0.031797f
C1149 minus.n7 gnd 0.007215f
C1150 minus.n8 gnd 0.031797f
C1151 minus.n9 gnd 0.007215f
C1152 minus.t8 gnd 0.466068f
C1153 minus.t7 gnd 0.449743f
C1154 minus.n10 gnd 0.206297f
C1155 minus.n11 gnd 0.185158f
C1156 minus.n12 gnd 0.136889f
C1157 minus.n13 gnd 0.031797f
C1158 minus.t11 gnd 0.449743f
C1159 minus.n14 gnd 0.19979f
C1160 minus.n15 gnd 0.007215f
C1161 minus.t10 gnd 0.449743f
C1162 minus.n16 gnd 0.19979f
C1163 minus.n17 gnd 0.031797f
C1164 minus.n18 gnd 0.031797f
C1165 minus.n19 gnd 0.031797f
C1166 minus.t12 gnd 0.449743f
C1167 minus.n20 gnd 0.19979f
C1168 minus.n21 gnd 0.007215f
C1169 minus.t20 gnd 0.449743f
C1170 minus.n22 gnd 0.19979f
C1171 minus.n23 gnd 0.031797f
C1172 minus.n24 gnd 0.031797f
C1173 minus.n25 gnd 0.031797f
C1174 minus.t18 gnd 0.449743f
C1175 minus.n26 gnd 0.19979f
C1176 minus.n27 gnd 0.007215f
C1177 minus.t25 gnd 0.449743f
C1178 minus.n28 gnd 0.19979f
C1179 minus.n29 gnd 0.031797f
C1180 minus.n30 gnd 0.031797f
C1181 minus.n31 gnd 0.031797f
C1182 minus.t24 gnd 0.449743f
C1183 minus.n32 gnd 0.19979f
C1184 minus.n33 gnd 0.007215f
C1185 minus.t14 gnd 0.449743f
C1186 minus.n34 gnd 0.19979f
C1187 minus.n35 gnd 0.031797f
C1188 minus.n36 gnd 0.031797f
C1189 minus.n37 gnd 0.031797f
C1190 minus.t22 gnd 0.449743f
C1191 minus.n38 gnd 0.19979f
C1192 minus.n39 gnd 0.007215f
C1193 minus.t19 gnd 0.449743f
C1194 minus.n40 gnd 0.200084f
C1195 minus.n41 gnd 0.368244f
C1196 minus.n42 gnd 0.031797f
C1197 minus.t13 gnd 0.449743f
C1198 minus.t15 gnd 0.449743f
C1199 minus.n43 gnd 0.031797f
C1200 minus.t5 gnd 0.449743f
C1201 minus.n44 gnd 0.19979f
C1202 minus.n45 gnd 0.031797f
C1203 minus.t6 gnd 0.449743f
C1204 minus.t26 gnd 0.449743f
C1205 minus.n46 gnd 0.19979f
C1206 minus.n47 gnd 0.031797f
C1207 minus.t21 gnd 0.449743f
C1208 minus.t23 gnd 0.449743f
C1209 minus.n48 gnd 0.19979f
C1210 minus.n49 gnd 0.031797f
C1211 minus.t16 gnd 0.449743f
C1212 minus.t17 gnd 0.449743f
C1213 minus.n50 gnd 0.19979f
C1214 minus.n51 gnd 0.031797f
C1215 minus.t9 gnd 0.449743f
C1216 minus.t27 gnd 0.449743f
C1217 minus.n52 gnd 0.206297f
C1218 minus.t28 gnd 0.466068f
C1219 minus.n53 gnd 0.185158f
C1220 minus.n54 gnd 0.136889f
C1221 minus.n55 gnd 0.007215f
C1222 minus.n56 gnd 0.19979f
C1223 minus.n57 gnd 0.007215f
C1224 minus.n58 gnd 0.031797f
C1225 minus.n59 gnd 0.031797f
C1226 minus.n60 gnd 0.031797f
C1227 minus.n61 gnd 0.007215f
C1228 minus.n62 gnd 0.19979f
C1229 minus.n63 gnd 0.007215f
C1230 minus.n64 gnd 0.031797f
C1231 minus.n65 gnd 0.031797f
C1232 minus.n66 gnd 0.031797f
C1233 minus.n67 gnd 0.007215f
C1234 minus.n68 gnd 0.19979f
C1235 minus.n69 gnd 0.007215f
C1236 minus.n70 gnd 0.031797f
C1237 minus.n71 gnd 0.031797f
C1238 minus.n72 gnd 0.031797f
C1239 minus.n73 gnd 0.007215f
C1240 minus.n74 gnd 0.19979f
C1241 minus.n75 gnd 0.007215f
C1242 minus.n76 gnd 0.031797f
C1243 minus.n77 gnd 0.031797f
C1244 minus.n78 gnd 0.031797f
C1245 minus.n79 gnd 0.007215f
C1246 minus.n80 gnd 0.19979f
C1247 minus.n81 gnd 0.007215f
C1248 minus.n82 gnd 0.200084f
C1249 minus.n83 gnd 1.06524f
C1250 minus.n84 gnd 1.58719f
C1251 minus.t1 gnd 0.009802f
C1252 minus.t0 gnd 0.009802f
C1253 minus.n85 gnd 0.032232f
C1254 minus.t4 gnd 0.009802f
C1255 minus.t3 gnd 0.009802f
C1256 minus.n86 gnd 0.03179f
C1257 minus.n87 gnd 0.271314f
C1258 minus.t2 gnd 0.054558f
C1259 minus.n88 gnd 0.148054f
C1260 minus.n89 gnd 2.10933f
C1261 a_n2140_13878.t11 gnd 0.186868f
C1262 a_n2140_13878.t10 gnd 0.186868f
C1263 a_n2140_13878.t5 gnd 0.186868f
C1264 a_n2140_13878.n0 gnd 1.47299f
C1265 a_n2140_13878.t2 gnd 0.186868f
C1266 a_n2140_13878.t4 gnd 0.186868f
C1267 a_n2140_13878.n1 gnd 1.47143f
C1268 a_n2140_13878.n2 gnd 2.05603f
C1269 a_n2140_13878.t12 gnd 0.186868f
C1270 a_n2140_13878.t3 gnd 0.186868f
C1271 a_n2140_13878.n3 gnd 1.47143f
C1272 a_n2140_13878.n4 gnd 1.00289f
C1273 a_n2140_13878.t9 gnd 0.186868f
C1274 a_n2140_13878.t1 gnd 0.186868f
C1275 a_n2140_13878.n5 gnd 1.47143f
C1276 a_n2140_13878.n6 gnd 4.06212f
C1277 a_n2140_13878.t17 gnd 1.74974f
C1278 a_n2140_13878.t20 gnd 0.186868f
C1279 a_n2140_13878.t21 gnd 0.186868f
C1280 a_n2140_13878.n7 gnd 1.3163f
C1281 a_n2140_13878.n8 gnd 1.47077f
C1282 a_n2140_13878.t16 gnd 1.74626f
C1283 a_n2140_13878.n9 gnd 0.740113f
C1284 a_n2140_13878.t19 gnd 1.74626f
C1285 a_n2140_13878.n10 gnd 0.740113f
C1286 a_n2140_13878.t22 gnd 0.186868f
C1287 a_n2140_13878.t23 gnd 0.186868f
C1288 a_n2140_13878.n11 gnd 1.3163f
C1289 a_n2140_13878.n12 gnd 0.74728f
C1290 a_n2140_13878.t18 gnd 1.74626f
C1291 a_n2140_13878.n13 gnd 2.09583f
C1292 a_n2140_13878.n14 gnd 2.85974f
C1293 a_n2140_13878.t6 gnd 0.186868f
C1294 a_n2140_13878.t7 gnd 0.186868f
C1295 a_n2140_13878.n15 gnd 1.47142f
C1296 a_n2140_13878.n16 gnd 2.01665f
C1297 a_n2140_13878.t13 gnd 0.186868f
C1298 a_n2140_13878.t14 gnd 0.186868f
C1299 a_n2140_13878.n17 gnd 1.47143f
C1300 a_n2140_13878.n18 gnd 0.651951f
C1301 a_n2140_13878.t0 gnd 0.186868f
C1302 a_n2140_13878.t8 gnd 0.186868f
C1303 a_n2140_13878.n19 gnd 1.47143f
C1304 a_n2140_13878.n20 gnd 1.32263f
C1305 a_n2140_13878.n21 gnd 1.47386f
C1306 a_n2140_13878.t15 gnd 0.186868f
C1307 a_n2408_n452.n0 gnd 3.95093f
C1308 a_n2408_n452.n1 gnd 2.90522f
C1309 a_n2408_n452.n2 gnd 3.88871f
C1310 a_n2408_n452.n3 gnd 0.820088f
C1311 a_n2408_n452.n4 gnd 0.82009f
C1312 a_n2408_n452.n5 gnd 0.668638f
C1313 a_n2408_n452.n6 gnd 0.204926f
C1314 a_n2408_n452.n7 gnd 0.150932f
C1315 a_n2408_n452.n8 gnd 0.237216f
C1316 a_n2408_n452.n9 gnd 0.183223f
C1317 a_n2408_n452.n10 gnd 0.204926f
C1318 a_n2408_n452.n11 gnd 0.150932f
C1319 a_n2408_n452.n12 gnd 0.722632f
C1320 a_n2408_n452.n13 gnd 0.512478f
C1321 a_n2408_n452.n14 gnd 0.215976f
C1322 a_n2408_n452.n15 gnd 0.215976f
C1323 a_n2408_n452.n16 gnd 0.44388f
C1324 a_n2408_n452.n17 gnd 0.215976f
C1325 a_n2408_n452.n18 gnd 0.215976f
C1326 a_n2408_n452.n19 gnd 0.668661f
C1327 a_n2408_n452.n20 gnd 0.215976f
C1328 a_n2408_n452.n21 gnd 0.215976f
C1329 a_n2408_n452.n22 gnd 0.747109f
C1330 a_n2408_n452.n23 gnd 0.215976f
C1331 a_n2408_n452.n24 gnd 0.44388f
C1332 a_n2408_n452.n25 gnd 3.3281f
C1333 a_n2408_n452.n26 gnd 1.7781f
C1334 a_n2408_n452.n27 gnd 1.89786f
C1335 a_n2408_n452.n28 gnd 1.7781f
C1336 a_n2408_n452.n29 gnd 2.07944f
C1337 a_n2408_n452.n30 gnd 0.285304f
C1338 a_n2408_n452.n31 gnd 0.285304f
C1339 a_n2408_n452.n32 gnd 0.004854f
C1340 a_n2408_n452.n33 gnd 0.010499f
C1341 a_n2408_n452.n34 gnd 0.010499f
C1342 a_n2408_n452.n35 gnd 0.004854f
C1343 a_n2408_n452.n36 gnd 1.45046f
C1344 a_n2408_n452.n37 gnd 0.285304f
C1345 a_n2408_n452.n38 gnd 0.285304f
C1346 a_n2408_n452.n39 gnd 0.004854f
C1347 a_n2408_n452.n40 gnd 0.010499f
C1348 a_n2408_n452.n41 gnd 0.010499f
C1349 a_n2408_n452.n42 gnd 0.285304f
C1350 a_n2408_n452.n43 gnd 0.76008f
C1351 a_n2408_n452.n44 gnd 0.004854f
C1352 a_n2408_n452.n45 gnd 0.010499f
C1353 a_n2408_n452.n46 gnd 0.010499f
C1354 a_n2408_n452.n47 gnd 0.004854f
C1355 a_n2408_n452.n48 gnd 0.285304f
C1356 a_n2408_n452.n49 gnd 0.285304f
C1357 a_n2408_n452.n50 gnd 0.44388f
C1358 a_n2408_n452.n51 gnd 0.004854f
C1359 a_n2408_n452.n52 gnd 0.010499f
C1360 a_n2408_n452.n53 gnd 0.010499f
C1361 a_n2408_n452.n54 gnd 0.004854f
C1362 a_n2408_n452.n55 gnd 0.285304f
C1363 a_n2408_n452.n56 gnd 0.008362f
C1364 a_n2408_n452.n57 gnd 0.285304f
C1365 a_n2408_n452.n58 gnd 0.008362f
C1366 a_n2408_n452.n59 gnd 0.285304f
C1367 a_n2408_n452.n60 gnd 0.008362f
C1368 a_n2408_n452.n61 gnd 0.285304f
C1369 a_n2408_n452.n62 gnd 0.008362f
C1370 a_n2408_n452.n63 gnd 0.285304f
C1371 a_n2408_n452.n64 gnd 0.004854f
C1372 a_n2408_n452.n65 gnd 0.304393f
C1373 a_n2408_n452.t24 gnd 0.149803f
C1374 a_n2408_n452.t12 gnd 1.40268f
C1375 a_n2408_n452.t20 gnd 0.149803f
C1376 a_n2408_n452.t16 gnd 0.149803f
C1377 a_n2408_n452.n66 gnd 1.05521f
C1378 a_n2408_n452.t36 gnd 0.149803f
C1379 a_n2408_n452.t40 gnd 0.149803f
C1380 a_n2408_n452.n67 gnd 1.05521f
C1381 a_n2408_n452.t9 gnd 0.696812f
C1382 a_n2408_n452.n68 gnd 0.304393f
C1383 a_n2408_n452.t35 gnd 0.696812f
C1384 a_n2408_n452.t11 gnd 0.708488f
C1385 a_n2408_n452.t19 gnd 0.696812f
C1386 a_n2408_n452.t66 gnd 0.696812f
C1387 a_n2408_n452.n69 gnd 0.304393f
C1388 a_n2408_n452.t80 gnd 0.696812f
C1389 a_n2408_n452.t82 gnd 0.708488f
C1390 a_n2408_n452.t60 gnd 0.696812f
C1391 a_n2408_n452.t13 gnd 0.708488f
C1392 a_n2408_n452.t29 gnd 0.696812f
C1393 a_n2408_n452.t27 gnd 0.696812f
C1394 a_n2408_n452.n70 gnd 0.304393f
C1395 a_n2408_n452.t37 gnd 0.696812f
C1396 a_n2408_n452.t33 gnd 0.696812f
C1397 a_n2408_n452.t21 gnd 0.696812f
C1398 a_n2408_n452.t31 gnd 0.696812f
C1399 a_n2408_n452.t17 gnd 0.708488f
C1400 a_n2408_n452.t86 gnd 0.708488f
C1401 a_n2408_n452.t67 gnd 0.696812f
C1402 a_n2408_n452.t71 gnd 0.696812f
C1403 a_n2408_n452.n71 gnd 0.304393f
C1404 a_n2408_n452.t61 gnd 0.696812f
C1405 a_n2408_n452.t76 gnd 0.696812f
C1406 a_n2408_n452.t83 gnd 0.696812f
C1407 a_n2408_n452.n72 gnd 0.304393f
C1408 a_n2408_n452.t84 gnd 0.696812f
C1409 a_n2408_n452.t58 gnd 0.708488f
C1410 a_n2408_n452.n73 gnd 0.306874f
C1411 a_n2408_n452.n74 gnd 0.299809f
C1412 a_n2408_n452.n75 gnd 0.299809f
C1413 a_n2408_n452.n76 gnd 0.306874f
C1414 a_n2408_n452.n77 gnd 0.306874f
C1415 a_n2408_n452.t55 gnd 0.116514f
C1416 a_n2408_n452.t44 gnd 0.116514f
C1417 a_n2408_n452.n78 gnd 1.03184f
C1418 a_n2408_n452.t49 gnd 0.116514f
C1419 a_n2408_n452.t4 gnd 0.116514f
C1420 a_n2408_n452.n79 gnd 1.02955f
C1421 a_n2408_n452.t41 gnd 0.116514f
C1422 a_n2408_n452.t47 gnd 0.116514f
C1423 a_n2408_n452.n80 gnd 1.02955f
C1424 a_n2408_n452.t46 gnd 0.116514f
C1425 a_n2408_n452.t8 gnd 0.116514f
C1426 a_n2408_n452.n81 gnd 1.03184f
C1427 a_n2408_n452.t52 gnd 0.116514f
C1428 a_n2408_n452.t45 gnd 0.116514f
C1429 a_n2408_n452.n82 gnd 1.02955f
C1430 a_n2408_n452.t2 gnd 0.116514f
C1431 a_n2408_n452.t53 gnd 0.116514f
C1432 a_n2408_n452.n83 gnd 1.02955f
C1433 a_n2408_n452.t0 gnd 0.116514f
C1434 a_n2408_n452.t6 gnd 0.116514f
C1435 a_n2408_n452.n84 gnd 1.02956f
C1436 a_n2408_n452.t3 gnd 0.116514f
C1437 a_n2408_n452.t48 gnd 0.116514f
C1438 a_n2408_n452.n85 gnd 1.02956f
C1439 a_n2408_n452.t7 gnd 0.116514f
C1440 a_n2408_n452.t42 gnd 0.116514f
C1441 a_n2408_n452.n86 gnd 1.02956f
C1442 a_n2408_n452.t54 gnd 0.116514f
C1443 a_n2408_n452.t1 gnd 0.116514f
C1444 a_n2408_n452.n87 gnd 1.03185f
C1445 a_n2408_n452.t43 gnd 0.116514f
C1446 a_n2408_n452.t51 gnd 0.116514f
C1447 a_n2408_n452.n88 gnd 1.02956f
C1448 a_n2408_n452.t50 gnd 0.116514f
C1449 a_n2408_n452.t5 gnd 0.116514f
C1450 a_n2408_n452.n89 gnd 1.02956f
C1451 a_n2408_n452.n90 gnd 0.299809f
C1452 a_n2408_n452.n91 gnd 0.299809f
C1453 a_n2408_n452.n92 gnd 0.306874f
C1454 a_n2408_n452.t18 gnd 1.40268f
C1455 a_n2408_n452.t22 gnd 0.149803f
C1456 a_n2408_n452.t32 gnd 0.149803f
C1457 a_n2408_n452.n93 gnd 1.05521f
C1458 a_n2408_n452.t38 gnd 0.149803f
C1459 a_n2408_n452.t34 gnd 0.149803f
C1460 a_n2408_n452.n94 gnd 1.05521f
C1461 a_n2408_n452.t30 gnd 0.149803f
C1462 a_n2408_n452.t28 gnd 0.149803f
C1463 a_n2408_n452.n95 gnd 1.05521f
C1464 a_n2408_n452.t14 gnd 1.39989f
C1465 a_n2408_n452.n96 gnd 0.859759f
C1466 a_n2408_n452.t65 gnd 0.696812f
C1467 a_n2408_n452.t74 gnd 0.696812f
C1468 a_n2408_n452.t87 gnd 0.696812f
C1469 a_n2408_n452.n97 gnd 0.306363f
C1470 a_n2408_n452.t77 gnd 0.696812f
C1471 a_n2408_n452.t62 gnd 0.696812f
C1472 a_n2408_n452.t63 gnd 0.696812f
C1473 a_n2408_n452.n98 gnd 0.306363f
C1474 a_n2408_n452.t81 gnd 0.696812f
C1475 a_n2408_n452.t70 gnd 0.696812f
C1476 a_n2408_n452.t69 gnd 0.696812f
C1477 a_n2408_n452.n99 gnd 0.306363f
C1478 a_n2408_n452.t73 gnd 0.696812f
C1479 a_n2408_n452.t64 gnd 0.696812f
C1480 a_n2408_n452.t56 gnd 0.696812f
C1481 a_n2408_n452.n100 gnd 0.306363f
C1482 a_n2408_n452.t78 gnd 0.708488f
C1483 a_n2408_n452.n101 gnd 0.302472f
C1484 a_n2408_n452.n102 gnd 0.296979f
C1485 a_n2408_n452.t85 gnd 0.708488f
C1486 a_n2408_n452.n103 gnd 0.302472f
C1487 a_n2408_n452.n104 gnd 0.296979f
C1488 a_n2408_n452.t72 gnd 0.708488f
C1489 a_n2408_n452.n105 gnd 0.302472f
C1490 a_n2408_n452.n106 gnd 0.296979f
C1491 a_n2408_n452.t68 gnd 0.708488f
C1492 a_n2408_n452.n107 gnd 0.302472f
C1493 a_n2408_n452.n108 gnd 0.296979f
C1494 a_n2408_n452.n109 gnd 1.1184f
C1495 a_n2408_n452.n110 gnd 0.306874f
C1496 a_n2408_n452.t79 gnd 0.696812f
C1497 a_n2408_n452.n111 gnd 0.304393f
C1498 a_n2408_n452.n112 gnd 0.299809f
C1499 a_n2408_n452.t57 gnd 0.696812f
C1500 a_n2408_n452.n113 gnd 0.299809f
C1501 a_n2408_n452.t75 gnd 0.696812f
C1502 a_n2408_n452.n114 gnd 0.306874f
C1503 a_n2408_n452.t59 gnd 0.708488f
C1504 a_n2408_n452.n115 gnd 0.306874f
C1505 a_n2408_n452.t15 gnd 0.696812f
C1506 a_n2408_n452.n116 gnd 0.304393f
C1507 a_n2408_n452.n117 gnd 0.299809f
C1508 a_n2408_n452.t39 gnd 0.696812f
C1509 a_n2408_n452.n118 gnd 0.299809f
C1510 a_n2408_n452.t23 gnd 0.696812f
C1511 a_n2408_n452.n119 gnd 0.306874f
C1512 a_n2408_n452.t25 gnd 0.708488f
C1513 a_n2408_n452.n120 gnd 1.19872f
C1514 a_n2408_n452.t26 gnd 1.39988f
C1515 a_n2408_n452.n121 gnd 1.05522f
C1516 a_n2408_n452.t10 gnd 0.149803f
C1517 CSoutput.n0 gnd 0.048261f
C1518 CSoutput.t197 gnd 0.319238f
C1519 CSoutput.n1 gnd 0.144152f
C1520 CSoutput.n2 gnd 0.048261f
C1521 CSoutput.t203 gnd 0.319238f
C1522 CSoutput.n3 gnd 0.038251f
C1523 CSoutput.n4 gnd 0.048261f
C1524 CSoutput.t192 gnd 0.319238f
C1525 CSoutput.n5 gnd 0.032984f
C1526 CSoutput.n6 gnd 0.048261f
C1527 CSoutput.t200 gnd 0.319238f
C1528 CSoutput.t184 gnd 0.319238f
C1529 CSoutput.n7 gnd 0.142581f
C1530 CSoutput.n8 gnd 0.048261f
C1531 CSoutput.t205 gnd 0.319238f
C1532 CSoutput.n9 gnd 0.031449f
C1533 CSoutput.n10 gnd 0.048261f
C1534 CSoutput.t193 gnd 0.319238f
C1535 CSoutput.t204 gnd 0.319238f
C1536 CSoutput.n11 gnd 0.142581f
C1537 CSoutput.n12 gnd 0.048261f
C1538 CSoutput.t201 gnd 0.319238f
C1539 CSoutput.n13 gnd 0.032984f
C1540 CSoutput.n14 gnd 0.048261f
C1541 CSoutput.t191 gnd 0.319238f
C1542 CSoutput.t194 gnd 0.319238f
C1543 CSoutput.n15 gnd 0.142581f
C1544 CSoutput.n16 gnd 0.048261f
C1545 CSoutput.t198 gnd 0.319238f
C1546 CSoutput.n17 gnd 0.035229f
C1547 CSoutput.t188 gnd 0.381497f
C1548 CSoutput.t190 gnd 0.319238f
C1549 CSoutput.n18 gnd 0.18202f
C1550 CSoutput.n19 gnd 0.176622f
C1551 CSoutput.n20 gnd 0.204903f
C1552 CSoutput.n21 gnd 0.048261f
C1553 CSoutput.n22 gnd 0.040279f
C1554 CSoutput.n23 gnd 0.142581f
C1555 CSoutput.n24 gnd 0.038828f
C1556 CSoutput.n25 gnd 0.038251f
C1557 CSoutput.n26 gnd 0.048261f
C1558 CSoutput.n27 gnd 0.048261f
C1559 CSoutput.n28 gnd 0.03997f
C1560 CSoutput.n29 gnd 0.033935f
C1561 CSoutput.n30 gnd 0.145755f
C1562 CSoutput.n31 gnd 0.034403f
C1563 CSoutput.n32 gnd 0.048261f
C1564 CSoutput.n33 gnd 0.048261f
C1565 CSoutput.n34 gnd 0.048261f
C1566 CSoutput.n35 gnd 0.039544f
C1567 CSoutput.n36 gnd 0.142581f
C1568 CSoutput.n37 gnd 0.037818f
C1569 CSoutput.n38 gnd 0.039261f
C1570 CSoutput.n39 gnd 0.048261f
C1571 CSoutput.n40 gnd 0.048261f
C1572 CSoutput.n41 gnd 0.040271f
C1573 CSoutput.n42 gnd 0.036808f
C1574 CSoutput.n43 gnd 0.142581f
C1575 CSoutput.n44 gnd 0.037741f
C1576 CSoutput.n45 gnd 0.048261f
C1577 CSoutput.n46 gnd 0.048261f
C1578 CSoutput.n47 gnd 0.048261f
C1579 CSoutput.n48 gnd 0.037741f
C1580 CSoutput.n49 gnd 0.142581f
C1581 CSoutput.n50 gnd 0.036808f
C1582 CSoutput.n51 gnd 0.040271f
C1583 CSoutput.n52 gnd 0.048261f
C1584 CSoutput.n53 gnd 0.048261f
C1585 CSoutput.n54 gnd 0.039261f
C1586 CSoutput.n55 gnd 0.037818f
C1587 CSoutput.n56 gnd 0.142581f
C1588 CSoutput.n57 gnd 0.039544f
C1589 CSoutput.n58 gnd 0.048261f
C1590 CSoutput.n59 gnd 0.048261f
C1591 CSoutput.n60 gnd 0.048261f
C1592 CSoutput.n61 gnd 0.034403f
C1593 CSoutput.n62 gnd 0.145755f
C1594 CSoutput.n63 gnd 0.033935f
C1595 CSoutput.t186 gnd 0.319238f
C1596 CSoutput.n64 gnd 0.142581f
C1597 CSoutput.n65 gnd 0.03997f
C1598 CSoutput.n66 gnd 0.048261f
C1599 CSoutput.n67 gnd 0.048261f
C1600 CSoutput.n68 gnd 0.048261f
C1601 CSoutput.n69 gnd 0.038828f
C1602 CSoutput.n70 gnd 0.142581f
C1603 CSoutput.n71 gnd 0.040279f
C1604 CSoutput.n72 gnd 0.035229f
C1605 CSoutput.n73 gnd 0.048261f
C1606 CSoutput.n74 gnd 0.048261f
C1607 CSoutput.n75 gnd 0.036535f
C1608 CSoutput.n76 gnd 0.021698f
C1609 CSoutput.t189 gnd 0.358686f
C1610 CSoutput.n77 gnd 0.178181f
C1611 CSoutput.n78 gnd 0.76242f
C1612 CSoutput.t103 gnd 0.060199f
C1613 CSoutput.t34 gnd 0.060199f
C1614 CSoutput.n79 gnd 0.466081f
C1615 CSoutput.t118 gnd 0.060199f
C1616 CSoutput.t56 gnd 0.060199f
C1617 CSoutput.n80 gnd 0.46525f
C1618 CSoutput.n81 gnd 0.472228f
C1619 CSoutput.t13 gnd 0.060199f
C1620 CSoutput.t73 gnd 0.060199f
C1621 CSoutput.n82 gnd 0.46525f
C1622 CSoutput.n83 gnd 0.232694f
C1623 CSoutput.t19 gnd 0.060199f
C1624 CSoutput.t47 gnd 0.060199f
C1625 CSoutput.n84 gnd 0.46525f
C1626 CSoutput.n85 gnd 0.232694f
C1627 CSoutput.t123 gnd 0.060199f
C1628 CSoutput.t66 gnd 0.060199f
C1629 CSoutput.n86 gnd 0.46525f
C1630 CSoutput.n87 gnd 0.232694f
C1631 CSoutput.t22 gnd 0.060199f
C1632 CSoutput.t107 gnd 0.060199f
C1633 CSoutput.n88 gnd 0.46525f
C1634 CSoutput.n89 gnd 0.232694f
C1635 CSoutput.t30 gnd 0.060199f
C1636 CSoutput.t83 gnd 0.060199f
C1637 CSoutput.n90 gnd 0.46525f
C1638 CSoutput.n91 gnd 0.232694f
C1639 CSoutput.t51 gnd 0.060199f
C1640 CSoutput.t74 gnd 0.060199f
C1641 CSoutput.n92 gnd 0.46525f
C1642 CSoutput.n93 gnd 0.232694f
C1643 CSoutput.t69 gnd 0.060199f
C1644 CSoutput.t112 gnd 0.060199f
C1645 CSoutput.n94 gnd 0.46525f
C1646 CSoutput.n95 gnd 0.232694f
C1647 CSoutput.t39 gnd 0.060199f
C1648 CSoutput.t90 gnd 0.060199f
C1649 CSoutput.n96 gnd 0.46525f
C1650 CSoutput.n97 gnd 0.426707f
C1651 CSoutput.t9 gnd 0.060199f
C1652 CSoutput.t101 gnd 0.060199f
C1653 CSoutput.n98 gnd 0.466081f
C1654 CSoutput.t84 gnd 0.060199f
C1655 CSoutput.t60 gnd 0.060199f
C1656 CSoutput.n99 gnd 0.46525f
C1657 CSoutput.n100 gnd 0.472228f
C1658 CSoutput.t35 gnd 0.060199f
C1659 CSoutput.t114 gnd 0.060199f
C1660 CSoutput.n101 gnd 0.46525f
C1661 CSoutput.n102 gnd 0.232694f
C1662 CSoutput.t81 gnd 0.060199f
C1663 CSoutput.t80 gnd 0.060199f
C1664 CSoutput.n103 gnd 0.46525f
C1665 CSoutput.n104 gnd 0.232694f
C1666 CSoutput.t70 gnd 0.060199f
C1667 CSoutput.t31 gnd 0.060199f
C1668 CSoutput.n105 gnd 0.46525f
C1669 CSoutput.n106 gnd 0.232694f
C1670 CSoutput.t12 gnd 0.060199f
C1671 CSoutput.t71 gnd 0.060199f
C1672 CSoutput.n107 gnd 0.46525f
C1673 CSoutput.n108 gnd 0.232694f
C1674 CSoutput.t67 gnd 0.060199f
C1675 CSoutput.t29 gnd 0.060199f
C1676 CSoutput.n109 gnd 0.46525f
C1677 CSoutput.n110 gnd 0.232694f
C1678 CSoutput.t10 gnd 0.060199f
C1679 CSoutput.t7 gnd 0.060199f
C1680 CSoutput.n111 gnd 0.46525f
C1681 CSoutput.n112 gnd 0.232694f
C1682 CSoutput.t85 gnd 0.060199f
C1683 CSoutput.t48 gnd 0.060199f
C1684 CSoutput.n113 gnd 0.46525f
C1685 CSoutput.n114 gnd 0.232694f
C1686 CSoutput.t41 gnd 0.060199f
C1687 CSoutput.t5 gnd 0.060199f
C1688 CSoutput.n115 gnd 0.46525f
C1689 CSoutput.n116 gnd 0.347005f
C1690 CSoutput.n117 gnd 0.437572f
C1691 CSoutput.t24 gnd 0.060199f
C1692 CSoutput.t113 gnd 0.060199f
C1693 CSoutput.n118 gnd 0.466081f
C1694 CSoutput.t94 gnd 0.060199f
C1695 CSoutput.t72 gnd 0.060199f
C1696 CSoutput.n119 gnd 0.46525f
C1697 CSoutput.n120 gnd 0.472228f
C1698 CSoutput.t52 gnd 0.060199f
C1699 CSoutput.t124 gnd 0.060199f
C1700 CSoutput.n121 gnd 0.46525f
C1701 CSoutput.n122 gnd 0.232694f
C1702 CSoutput.t93 gnd 0.060199f
C1703 CSoutput.t92 gnd 0.060199f
C1704 CSoutput.n123 gnd 0.46525f
C1705 CSoutput.n124 gnd 0.232694f
C1706 CSoutput.t78 gnd 0.060199f
C1707 CSoutput.t49 gnd 0.060199f
C1708 CSoutput.n125 gnd 0.46525f
C1709 CSoutput.n126 gnd 0.232694f
C1710 CSoutput.t26 gnd 0.060199f
C1711 CSoutput.t79 gnd 0.060199f
C1712 CSoutput.n127 gnd 0.46525f
C1713 CSoutput.n128 gnd 0.232694f
C1714 CSoutput.t77 gnd 0.060199f
C1715 CSoutput.t46 gnd 0.060199f
C1716 CSoutput.n129 gnd 0.46525f
C1717 CSoutput.n130 gnd 0.232694f
C1718 CSoutput.t25 gnd 0.060199f
C1719 CSoutput.t23 gnd 0.060199f
C1720 CSoutput.n131 gnd 0.46525f
C1721 CSoutput.n132 gnd 0.232694f
C1722 CSoutput.t95 gnd 0.060199f
C1723 CSoutput.t62 gnd 0.060199f
C1724 CSoutput.n133 gnd 0.46525f
C1725 CSoutput.n134 gnd 0.232694f
C1726 CSoutput.t57 gnd 0.060199f
C1727 CSoutput.t18 gnd 0.060199f
C1728 CSoutput.n135 gnd 0.46525f
C1729 CSoutput.n136 gnd 0.347005f
C1730 CSoutput.n137 gnd 0.489093f
C1731 CSoutput.n138 gnd 9.6554f
C1732 CSoutput.n140 gnd 0.853732f
C1733 CSoutput.n141 gnd 0.640299f
C1734 CSoutput.n142 gnd 0.853732f
C1735 CSoutput.n143 gnd 0.853732f
C1736 CSoutput.n144 gnd 2.29851f
C1737 CSoutput.n145 gnd 0.853732f
C1738 CSoutput.n146 gnd 0.853732f
C1739 CSoutput.t185 gnd 1.06717f
C1740 CSoutput.n147 gnd 0.853732f
C1741 CSoutput.n148 gnd 0.853732f
C1742 CSoutput.n152 gnd 0.853732f
C1743 CSoutput.n156 gnd 0.853732f
C1744 CSoutput.n157 gnd 0.853732f
C1745 CSoutput.n159 gnd 0.853732f
C1746 CSoutput.n164 gnd 0.853732f
C1747 CSoutput.n166 gnd 0.853732f
C1748 CSoutput.n167 gnd 0.853732f
C1749 CSoutput.n169 gnd 0.853732f
C1750 CSoutput.n170 gnd 0.853732f
C1751 CSoutput.n172 gnd 0.853732f
C1752 CSoutput.t196 gnd 14.2658f
C1753 CSoutput.n174 gnd 0.853732f
C1754 CSoutput.n175 gnd 0.640299f
C1755 CSoutput.n176 gnd 0.853732f
C1756 CSoutput.n177 gnd 0.853732f
C1757 CSoutput.n178 gnd 2.29851f
C1758 CSoutput.n179 gnd 0.853732f
C1759 CSoutput.n180 gnd 0.853732f
C1760 CSoutput.t199 gnd 1.06717f
C1761 CSoutput.n181 gnd 0.853732f
C1762 CSoutput.n182 gnd 0.853732f
C1763 CSoutput.n186 gnd 0.853732f
C1764 CSoutput.n190 gnd 0.853732f
C1765 CSoutput.n191 gnd 0.853732f
C1766 CSoutput.n193 gnd 0.853732f
C1767 CSoutput.n198 gnd 0.853732f
C1768 CSoutput.n200 gnd 0.853732f
C1769 CSoutput.n201 gnd 0.853732f
C1770 CSoutput.n203 gnd 0.853732f
C1771 CSoutput.n204 gnd 0.853732f
C1772 CSoutput.n206 gnd 0.853732f
C1773 CSoutput.n207 gnd 0.640299f
C1774 CSoutput.n209 gnd 0.853732f
C1775 CSoutput.n210 gnd 0.640299f
C1776 CSoutput.n211 gnd 0.853732f
C1777 CSoutput.n212 gnd 0.853732f
C1778 CSoutput.n213 gnd 2.29851f
C1779 CSoutput.n214 gnd 0.853732f
C1780 CSoutput.n215 gnd 0.853732f
C1781 CSoutput.t195 gnd 1.06717f
C1782 CSoutput.n216 gnd 0.853732f
C1783 CSoutput.n217 gnd 2.29851f
C1784 CSoutput.n219 gnd 0.853732f
C1785 CSoutput.n220 gnd 0.853732f
C1786 CSoutput.n222 gnd 0.853732f
C1787 CSoutput.n223 gnd 0.853732f
C1788 CSoutput.t202 gnd 14.033299f
C1789 CSoutput.t187 gnd 14.2658f
C1790 CSoutput.n229 gnd 2.67828f
C1791 CSoutput.n230 gnd 10.9104f
C1792 CSoutput.n231 gnd 11.3669f
C1793 CSoutput.n236 gnd 2.9013f
C1794 CSoutput.n242 gnd 0.853732f
C1795 CSoutput.n244 gnd 0.853732f
C1796 CSoutput.n246 gnd 0.853732f
C1797 CSoutput.n248 gnd 0.853732f
C1798 CSoutput.n250 gnd 0.853732f
C1799 CSoutput.n256 gnd 0.853732f
C1800 CSoutput.n263 gnd 1.56627f
C1801 CSoutput.n264 gnd 1.56627f
C1802 CSoutput.n265 gnd 0.853732f
C1803 CSoutput.n266 gnd 0.853732f
C1804 CSoutput.n268 gnd 0.640299f
C1805 CSoutput.n269 gnd 0.548359f
C1806 CSoutput.n271 gnd 0.640299f
C1807 CSoutput.n272 gnd 0.548359f
C1808 CSoutput.n273 gnd 0.640299f
C1809 CSoutput.n275 gnd 0.853732f
C1810 CSoutput.n277 gnd 2.29851f
C1811 CSoutput.n278 gnd 2.67828f
C1812 CSoutput.n279 gnd 10.0347f
C1813 CSoutput.n281 gnd 0.640299f
C1814 CSoutput.n282 gnd 1.64753f
C1815 CSoutput.n283 gnd 0.640299f
C1816 CSoutput.n285 gnd 0.853732f
C1817 CSoutput.n287 gnd 2.29851f
C1818 CSoutput.n288 gnd 5.00653f
C1819 CSoutput.t33 gnd 0.060199f
C1820 CSoutput.t102 gnd 0.060199f
C1821 CSoutput.n289 gnd 0.466081f
C1822 CSoutput.t55 gnd 0.060199f
C1823 CSoutput.t116 gnd 0.060199f
C1824 CSoutput.n290 gnd 0.46525f
C1825 CSoutput.n291 gnd 0.472228f
C1826 CSoutput.t96 gnd 0.060199f
C1827 CSoutput.t11 gnd 0.060199f
C1828 CSoutput.n292 gnd 0.46525f
C1829 CSoutput.n293 gnd 0.232694f
C1830 CSoutput.t45 gnd 0.060199f
C1831 CSoutput.t17 gnd 0.060199f
C1832 CSoutput.n294 gnd 0.46525f
C1833 CSoutput.n295 gnd 0.232694f
C1834 CSoutput.t65 gnd 0.060199f
C1835 CSoutput.t38 gnd 0.060199f
C1836 CSoutput.n296 gnd 0.46525f
C1837 CSoutput.n297 gnd 0.232694f
C1838 CSoutput.t106 gnd 0.060199f
C1839 CSoutput.t21 gnd 0.060199f
C1840 CSoutput.n298 gnd 0.46525f
C1841 CSoutput.n299 gnd 0.232694f
C1842 CSoutput.t82 gnd 0.060199f
C1843 CSoutput.t27 gnd 0.060199f
C1844 CSoutput.n300 gnd 0.46525f
C1845 CSoutput.n301 gnd 0.232694f
C1846 CSoutput.t98 gnd 0.060199f
C1847 CSoutput.t50 gnd 0.060199f
C1848 CSoutput.n302 gnd 0.46525f
C1849 CSoutput.n303 gnd 0.232694f
C1850 CSoutput.t111 gnd 0.060199f
C1851 CSoutput.t68 gnd 0.060199f
C1852 CSoutput.n304 gnd 0.46525f
C1853 CSoutput.n305 gnd 0.232694f
C1854 CSoutput.t89 gnd 0.060199f
C1855 CSoutput.t40 gnd 0.060199f
C1856 CSoutput.n306 gnd 0.46525f
C1857 CSoutput.n307 gnd 0.426707f
C1858 CSoutput.t64 gnd 0.060199f
C1859 CSoutput.t88 gnd 0.060199f
C1860 CSoutput.n308 gnd 0.466081f
C1861 CSoutput.t6 gnd 0.060199f
C1862 CSoutput.t43 gnd 0.060199f
C1863 CSoutput.n309 gnd 0.46525f
C1864 CSoutput.n310 gnd 0.472228f
C1865 CSoutput.t44 gnd 0.060199f
C1866 CSoutput.t110 gnd 0.060199f
C1867 CSoutput.n311 gnd 0.46525f
C1868 CSoutput.n312 gnd 0.232694f
C1869 CSoutput.t36 gnd 0.060199f
C1870 CSoutput.t37 gnd 0.060199f
C1871 CSoutput.n313 gnd 0.46525f
C1872 CSoutput.n314 gnd 0.232694f
C1873 CSoutput.t108 gnd 0.060199f
C1874 CSoutput.t109 gnd 0.060199f
C1875 CSoutput.n315 gnd 0.46525f
C1876 CSoutput.n316 gnd 0.232694f
C1877 CSoutput.t16 gnd 0.060199f
C1878 CSoutput.t91 gnd 0.060199f
C1879 CSoutput.n317 gnd 0.46525f
C1880 CSoutput.n318 gnd 0.232694f
C1881 CSoutput.t105 gnd 0.060199f
C1882 CSoutput.t14 gnd 0.060199f
C1883 CSoutput.n319 gnd 0.46525f
C1884 CSoutput.n320 gnd 0.232694f
C1885 CSoutput.t63 gnd 0.060199f
C1886 CSoutput.t87 gnd 0.060199f
C1887 CSoutput.n321 gnd 0.46525f
C1888 CSoutput.n322 gnd 0.232694f
C1889 CSoutput.t117 gnd 0.060199f
C1890 CSoutput.t42 gnd 0.060199f
C1891 CSoutput.n323 gnd 0.46525f
C1892 CSoutput.n324 gnd 0.232694f
C1893 CSoutput.t86 gnd 0.060199f
C1894 CSoutput.t122 gnd 0.060199f
C1895 CSoutput.n325 gnd 0.46525f
C1896 CSoutput.n326 gnd 0.347005f
C1897 CSoutput.n327 gnd 0.437572f
C1898 CSoutput.t75 gnd 0.060199f
C1899 CSoutput.t99 gnd 0.060199f
C1900 CSoutput.n328 gnd 0.466081f
C1901 CSoutput.t20 gnd 0.060199f
C1902 CSoutput.t58 gnd 0.060199f
C1903 CSoutput.n329 gnd 0.46525f
C1904 CSoutput.n330 gnd 0.472228f
C1905 CSoutput.t61 gnd 0.060199f
C1906 CSoutput.t121 gnd 0.060199f
C1907 CSoutput.n331 gnd 0.46525f
C1908 CSoutput.n332 gnd 0.232694f
C1909 CSoutput.t53 gnd 0.060199f
C1910 CSoutput.t54 gnd 0.060199f
C1911 CSoutput.n333 gnd 0.46525f
C1912 CSoutput.n334 gnd 0.232694f
C1913 CSoutput.t119 gnd 0.060199f
C1914 CSoutput.t120 gnd 0.060199f
C1915 CSoutput.n335 gnd 0.46525f
C1916 CSoutput.n336 gnd 0.232694f
C1917 CSoutput.t32 gnd 0.060199f
C1918 CSoutput.t104 gnd 0.060199f
C1919 CSoutput.n337 gnd 0.46525f
C1920 CSoutput.n338 gnd 0.232694f
C1921 CSoutput.t115 gnd 0.060199f
C1922 CSoutput.t28 gnd 0.060199f
C1923 CSoutput.n339 gnd 0.46525f
C1924 CSoutput.n340 gnd 0.232694f
C1925 CSoutput.t76 gnd 0.060199f
C1926 CSoutput.t100 gnd 0.060199f
C1927 CSoutput.n341 gnd 0.46525f
C1928 CSoutput.n342 gnd 0.232694f
C1929 CSoutput.t8 gnd 0.060199f
C1930 CSoutput.t59 gnd 0.060199f
C1931 CSoutput.n343 gnd 0.46525f
C1932 CSoutput.n344 gnd 0.232694f
C1933 CSoutput.t97 gnd 0.060199f
C1934 CSoutput.t15 gnd 0.060199f
C1935 CSoutput.n345 gnd 0.465248f
C1936 CSoutput.n346 gnd 0.347007f
C1937 CSoutput.n347 gnd 0.489093f
C1938 CSoutput.n348 gnd 13.526501f
C1939 CSoutput.t129 gnd 0.052674f
C1940 CSoutput.t159 gnd 0.052674f
C1941 CSoutput.n349 gnd 0.467005f
C1942 CSoutput.t154 gnd 0.052674f
C1943 CSoutput.t142 gnd 0.052674f
C1944 CSoutput.n350 gnd 0.465448f
C1945 CSoutput.n351 gnd 0.43371f
C1946 CSoutput.t163 gnd 0.052674f
C1947 CSoutput.t146 gnd 0.052674f
C1948 CSoutput.n352 gnd 0.465448f
C1949 CSoutput.n353 gnd 0.213799f
C1950 CSoutput.t170 gnd 0.052674f
C1951 CSoutput.t155 gnd 0.052674f
C1952 CSoutput.n354 gnd 0.465448f
C1953 CSoutput.n355 gnd 0.213799f
C1954 CSoutput.t182 gnd 0.052674f
C1955 CSoutput.t176 gnd 0.052674f
C1956 CSoutput.n356 gnd 0.465448f
C1957 CSoutput.n357 gnd 0.213799f
C1958 CSoutput.t140 gnd 0.052674f
C1959 CSoutput.t132 gnd 0.052674f
C1960 CSoutput.n358 gnd 0.465448f
C1961 CSoutput.n359 gnd 0.213799f
C1962 CSoutput.t160 gnd 0.052674f
C1963 CSoutput.t137 gnd 0.052674f
C1964 CSoutput.n360 gnd 0.465448f
C1965 CSoutput.n361 gnd 0.213799f
C1966 CSoutput.t3 gnd 0.052674f
C1967 CSoutput.t169 gnd 0.052674f
C1968 CSoutput.n362 gnd 0.465448f
C1969 CSoutput.n363 gnd 0.394288f
C1970 CSoutput.t181 gnd 0.052674f
C1971 CSoutput.t2 gnd 0.052674f
C1972 CSoutput.n364 gnd 0.467005f
C1973 CSoutput.t148 gnd 0.052674f
C1974 CSoutput.t151 gnd 0.052674f
C1975 CSoutput.n365 gnd 0.465448f
C1976 CSoutput.n366 gnd 0.43371f
C1977 CSoutput.t139 gnd 0.052674f
C1978 CSoutput.t162 gnd 0.052674f
C1979 CSoutput.n367 gnd 0.465448f
C1980 CSoutput.n368 gnd 0.213799f
C1981 CSoutput.t171 gnd 0.052674f
C1982 CSoutput.t174 gnd 0.052674f
C1983 CSoutput.n369 gnd 0.465448f
C1984 CSoutput.n370 gnd 0.213799f
C1985 CSoutput.t180 gnd 0.052674f
C1986 CSoutput.t147 gnd 0.052674f
C1987 CSoutput.n371 gnd 0.465448f
C1988 CSoutput.n372 gnd 0.213799f
C1989 CSoutput.t164 gnd 0.052674f
C1990 CSoutput.t149 gnd 0.052674f
C1991 CSoutput.n373 gnd 0.465448f
C1992 CSoutput.n374 gnd 0.213799f
C1993 CSoutput.t4 gnd 0.052674f
C1994 CSoutput.t141 gnd 0.052674f
C1995 CSoutput.n375 gnd 0.465448f
C1996 CSoutput.n376 gnd 0.213799f
C1997 CSoutput.t156 gnd 0.052674f
C1998 CSoutput.t133 gnd 0.052674f
C1999 CSoutput.n377 gnd 0.465448f
C2000 CSoutput.n378 gnd 0.324592f
C2001 CSoutput.n379 gnd 0.603117f
C2002 CSoutput.n380 gnd 14.022901f
C2003 CSoutput.t166 gnd 0.052674f
C2004 CSoutput.t157 gnd 0.052674f
C2005 CSoutput.n381 gnd 0.467005f
C2006 CSoutput.t173 gnd 0.052674f
C2007 CSoutput.t172 gnd 0.052674f
C2008 CSoutput.n382 gnd 0.465448f
C2009 CSoutput.n383 gnd 0.43371f
C2010 CSoutput.t175 gnd 0.052674f
C2011 CSoutput.t1 gnd 0.052674f
C2012 CSoutput.n384 gnd 0.465448f
C2013 CSoutput.n385 gnd 0.213799f
C2014 CSoutput.t126 gnd 0.052674f
C2015 CSoutput.t143 gnd 0.052674f
C2016 CSoutput.n386 gnd 0.465448f
C2017 CSoutput.n387 gnd 0.213799f
C2018 CSoutput.t152 gnd 0.052674f
C2019 CSoutput.t145 gnd 0.052674f
C2020 CSoutput.n388 gnd 0.465448f
C2021 CSoutput.n389 gnd 0.213799f
C2022 CSoutput.t135 gnd 0.052674f
C2023 CSoutput.t128 gnd 0.052674f
C2024 CSoutput.n390 gnd 0.465448f
C2025 CSoutput.n391 gnd 0.213799f
C2026 CSoutput.t165 gnd 0.052674f
C2027 CSoutput.t167 gnd 0.052674f
C2028 CSoutput.n392 gnd 0.465448f
C2029 CSoutput.n393 gnd 0.213799f
C2030 CSoutput.t0 gnd 0.052674f
C2031 CSoutput.t161 gnd 0.052674f
C2032 CSoutput.n394 gnd 0.465448f
C2033 CSoutput.n395 gnd 0.394288f
C2034 CSoutput.t168 gnd 0.052674f
C2035 CSoutput.t127 gnd 0.052674f
C2036 CSoutput.n396 gnd 0.467005f
C2037 CSoutput.t138 gnd 0.052674f
C2038 CSoutput.t144 gnd 0.052674f
C2039 CSoutput.n397 gnd 0.465448f
C2040 CSoutput.n398 gnd 0.43371f
C2041 CSoutput.t153 gnd 0.052674f
C2042 CSoutput.t179 gnd 0.052674f
C2043 CSoutput.n399 gnd 0.465448f
C2044 CSoutput.n400 gnd 0.213799f
C2045 CSoutput.t150 gnd 0.052674f
C2046 CSoutput.t130 gnd 0.052674f
C2047 CSoutput.n401 gnd 0.465448f
C2048 CSoutput.n402 gnd 0.213799f
C2049 CSoutput.t134 gnd 0.052674f
C2050 CSoutput.t158 gnd 0.052674f
C2051 CSoutput.n403 gnd 0.465448f
C2052 CSoutput.n404 gnd 0.213799f
C2053 CSoutput.t131 gnd 0.052674f
C2054 CSoutput.t125 gnd 0.052674f
C2055 CSoutput.n405 gnd 0.465448f
C2056 CSoutput.n406 gnd 0.213799f
C2057 CSoutput.t136 gnd 0.052674f
C2058 CSoutput.t178 gnd 0.052674f
C2059 CSoutput.n407 gnd 0.465448f
C2060 CSoutput.n408 gnd 0.213799f
C2061 CSoutput.t177 gnd 0.052674f
C2062 CSoutput.t183 gnd 0.052674f
C2063 CSoutput.n409 gnd 0.465448f
C2064 CSoutput.n410 gnd 0.324592f
C2065 CSoutput.n411 gnd 0.603117f
C2066 CSoutput.n412 gnd 8.385481f
C2067 CSoutput.n413 gnd 15.5359f
C2068 vdd.t204 gnd 0.039211f
C2069 vdd.t214 gnd 0.039211f
C2070 vdd.n0 gnd 0.309267f
C2071 vdd.t297 gnd 0.039211f
C2072 vdd.t16 gnd 0.039211f
C2073 vdd.n1 gnd 0.308756f
C2074 vdd.n2 gnd 0.284732f
C2075 vdd.t3 gnd 0.039211f
C2076 vdd.t207 gnd 0.039211f
C2077 vdd.n3 gnd 0.308756f
C2078 vdd.n4 gnd 0.144f
C2079 vdd.t200 gnd 0.039211f
C2080 vdd.t210 gnd 0.039211f
C2081 vdd.n5 gnd 0.308756f
C2082 vdd.n6 gnd 0.135117f
C2083 vdd.t188 gnd 0.039211f
C2084 vdd.t190 gnd 0.039211f
C2085 vdd.n7 gnd 0.309267f
C2086 vdd.t212 gnd 0.039211f
C2087 vdd.t202 gnd 0.039211f
C2088 vdd.n8 gnd 0.308756f
C2089 vdd.n9 gnd 0.284732f
C2090 vdd.t195 gnd 0.039211f
C2091 vdd.t299 gnd 0.039211f
C2092 vdd.n10 gnd 0.308756f
C2093 vdd.n11 gnd 0.144f
C2094 vdd.t294 gnd 0.039211f
C2095 vdd.t197 gnd 0.039211f
C2096 vdd.n12 gnd 0.308756f
C2097 vdd.n13 gnd 0.135117f
C2098 vdd.n14 gnd 0.095525f
C2099 vdd.t192 gnd 0.021784f
C2100 vdd.t8 gnd 0.021784f
C2101 vdd.n15 gnd 0.200514f
C2102 vdd.t178 gnd 0.021784f
C2103 vdd.t4 gnd 0.021784f
C2104 vdd.n16 gnd 0.199927f
C2105 vdd.n17 gnd 0.347935f
C2106 vdd.t181 gnd 0.021784f
C2107 vdd.t184 gnd 0.021784f
C2108 vdd.n18 gnd 0.199927f
C2109 vdd.n19 gnd 0.143945f
C2110 vdd.t7 gnd 0.021784f
C2111 vdd.t9 gnd 0.021784f
C2112 vdd.n20 gnd 0.200514f
C2113 vdd.t193 gnd 0.021784f
C2114 vdd.t186 gnd 0.021784f
C2115 vdd.n21 gnd 0.199927f
C2116 vdd.n22 gnd 0.347935f
C2117 vdd.t183 gnd 0.021784f
C2118 vdd.t182 gnd 0.021784f
C2119 vdd.n23 gnd 0.199927f
C2120 vdd.n24 gnd 0.143945f
C2121 vdd.t5 gnd 0.021784f
C2122 vdd.t185 gnd 0.021784f
C2123 vdd.n25 gnd 0.199927f
C2124 vdd.t6 gnd 0.021784f
C2125 vdd.t177 gnd 0.021784f
C2126 vdd.n26 gnd 0.199927f
C2127 vdd.n27 gnd 23.2416f
C2128 vdd.n28 gnd 8.862241f
C2129 vdd.n29 gnd 0.005941f
C2130 vdd.n30 gnd 0.005513f
C2131 vdd.n31 gnd 0.00305f
C2132 vdd.n32 gnd 0.007003f
C2133 vdd.n33 gnd 0.002963f
C2134 vdd.n34 gnd 0.003137f
C2135 vdd.n35 gnd 0.005513f
C2136 vdd.n36 gnd 0.002963f
C2137 vdd.n37 gnd 0.007003f
C2138 vdd.n38 gnd 0.003137f
C2139 vdd.n39 gnd 0.005513f
C2140 vdd.n40 gnd 0.002963f
C2141 vdd.n41 gnd 0.005252f
C2142 vdd.n42 gnd 0.005268f
C2143 vdd.t64 gnd 0.015044f
C2144 vdd.n43 gnd 0.033474f
C2145 vdd.n44 gnd 0.174205f
C2146 vdd.n45 gnd 0.002963f
C2147 vdd.n46 gnd 0.003137f
C2148 vdd.n47 gnd 0.007003f
C2149 vdd.n48 gnd 0.007003f
C2150 vdd.n49 gnd 0.003137f
C2151 vdd.n50 gnd 0.002963f
C2152 vdd.n51 gnd 0.005513f
C2153 vdd.n52 gnd 0.005513f
C2154 vdd.n53 gnd 0.002963f
C2155 vdd.n54 gnd 0.003137f
C2156 vdd.n55 gnd 0.007003f
C2157 vdd.n56 gnd 0.007003f
C2158 vdd.n57 gnd 0.003137f
C2159 vdd.n58 gnd 0.002963f
C2160 vdd.n59 gnd 0.005513f
C2161 vdd.n60 gnd 0.005513f
C2162 vdd.n61 gnd 0.002963f
C2163 vdd.n62 gnd 0.003137f
C2164 vdd.n63 gnd 0.007003f
C2165 vdd.n64 gnd 0.007003f
C2166 vdd.n65 gnd 0.016556f
C2167 vdd.n66 gnd 0.00305f
C2168 vdd.n67 gnd 0.002963f
C2169 vdd.n68 gnd 0.01425f
C2170 vdd.n69 gnd 0.009949f
C2171 vdd.t154 gnd 0.034855f
C2172 vdd.t96 gnd 0.034855f
C2173 vdd.n70 gnd 0.239545f
C2174 vdd.n71 gnd 0.188365f
C2175 vdd.t168 gnd 0.034855f
C2176 vdd.t147 gnd 0.034855f
C2177 vdd.n72 gnd 0.239545f
C2178 vdd.n73 gnd 0.15201f
C2179 vdd.t30 gnd 0.034855f
C2180 vdd.t83 gnd 0.034855f
C2181 vdd.n74 gnd 0.239545f
C2182 vdd.n75 gnd 0.15201f
C2183 vdd.t42 gnd 0.034855f
C2184 vdd.t109 gnd 0.034855f
C2185 vdd.n76 gnd 0.239545f
C2186 vdd.n77 gnd 0.15201f
C2187 vdd.t72 gnd 0.034855f
C2188 vdd.t158 gnd 0.034855f
C2189 vdd.n78 gnd 0.239545f
C2190 vdd.n79 gnd 0.15201f
C2191 vdd.t48 gnd 0.034855f
C2192 vdd.t131 gnd 0.034855f
C2193 vdd.n80 gnd 0.239545f
C2194 vdd.n81 gnd 0.15201f
C2195 vdd.t54 gnd 0.034855f
C2196 vdd.t150 gnd 0.034855f
C2197 vdd.n82 gnd 0.239545f
C2198 vdd.n83 gnd 0.15201f
C2199 vdd.t91 gnd 0.034855f
C2200 vdd.t163 gnd 0.034855f
C2201 vdd.n84 gnd 0.239545f
C2202 vdd.n85 gnd 0.15201f
C2203 vdd.t115 gnd 0.034855f
C2204 vdd.t141 gnd 0.034855f
C2205 vdd.n86 gnd 0.239545f
C2206 vdd.n87 gnd 0.15201f
C2207 vdd.n88 gnd 0.005941f
C2208 vdd.n89 gnd 0.005513f
C2209 vdd.n90 gnd 0.00305f
C2210 vdd.n91 gnd 0.007003f
C2211 vdd.n92 gnd 0.002963f
C2212 vdd.n93 gnd 0.003137f
C2213 vdd.n94 gnd 0.005513f
C2214 vdd.n95 gnd 0.002963f
C2215 vdd.n96 gnd 0.007003f
C2216 vdd.n97 gnd 0.003137f
C2217 vdd.n98 gnd 0.005513f
C2218 vdd.n99 gnd 0.002963f
C2219 vdd.n100 gnd 0.005252f
C2220 vdd.n101 gnd 0.005268f
C2221 vdd.t75 gnd 0.015044f
C2222 vdd.n102 gnd 0.033474f
C2223 vdd.n103 gnd 0.174205f
C2224 vdd.n104 gnd 0.002963f
C2225 vdd.n105 gnd 0.003137f
C2226 vdd.n106 gnd 0.007003f
C2227 vdd.n107 gnd 0.007003f
C2228 vdd.n108 gnd 0.003137f
C2229 vdd.n109 gnd 0.002963f
C2230 vdd.n110 gnd 0.005513f
C2231 vdd.n111 gnd 0.005513f
C2232 vdd.n112 gnd 0.002963f
C2233 vdd.n113 gnd 0.003137f
C2234 vdd.n114 gnd 0.007003f
C2235 vdd.n115 gnd 0.007003f
C2236 vdd.n116 gnd 0.003137f
C2237 vdd.n117 gnd 0.002963f
C2238 vdd.n118 gnd 0.005513f
C2239 vdd.n119 gnd 0.005513f
C2240 vdd.n120 gnd 0.002963f
C2241 vdd.n121 gnd 0.003137f
C2242 vdd.n122 gnd 0.007003f
C2243 vdd.n123 gnd 0.007003f
C2244 vdd.n124 gnd 0.016556f
C2245 vdd.n125 gnd 0.00305f
C2246 vdd.n126 gnd 0.002963f
C2247 vdd.n127 gnd 0.01425f
C2248 vdd.n128 gnd 0.009637f
C2249 vdd.n129 gnd 0.113096f
C2250 vdd.n130 gnd 0.005941f
C2251 vdd.n131 gnd 0.005513f
C2252 vdd.n132 gnd 0.00305f
C2253 vdd.n133 gnd 0.007003f
C2254 vdd.n134 gnd 0.002963f
C2255 vdd.n135 gnd 0.003137f
C2256 vdd.n136 gnd 0.005513f
C2257 vdd.n137 gnd 0.002963f
C2258 vdd.n138 gnd 0.007003f
C2259 vdd.n139 gnd 0.003137f
C2260 vdd.n140 gnd 0.005513f
C2261 vdd.n141 gnd 0.002963f
C2262 vdd.n142 gnd 0.005252f
C2263 vdd.n143 gnd 0.005268f
C2264 vdd.t107 gnd 0.015044f
C2265 vdd.n144 gnd 0.033474f
C2266 vdd.n145 gnd 0.174205f
C2267 vdd.n146 gnd 0.002963f
C2268 vdd.n147 gnd 0.003137f
C2269 vdd.n148 gnd 0.007003f
C2270 vdd.n149 gnd 0.007003f
C2271 vdd.n150 gnd 0.003137f
C2272 vdd.n151 gnd 0.002963f
C2273 vdd.n152 gnd 0.005513f
C2274 vdd.n153 gnd 0.005513f
C2275 vdd.n154 gnd 0.002963f
C2276 vdd.n155 gnd 0.003137f
C2277 vdd.n156 gnd 0.007003f
C2278 vdd.n157 gnd 0.007003f
C2279 vdd.n158 gnd 0.003137f
C2280 vdd.n159 gnd 0.002963f
C2281 vdd.n160 gnd 0.005513f
C2282 vdd.n161 gnd 0.005513f
C2283 vdd.n162 gnd 0.002963f
C2284 vdd.n163 gnd 0.003137f
C2285 vdd.n164 gnd 0.007003f
C2286 vdd.n165 gnd 0.007003f
C2287 vdd.n166 gnd 0.016556f
C2288 vdd.n167 gnd 0.00305f
C2289 vdd.n168 gnd 0.002963f
C2290 vdd.n169 gnd 0.01425f
C2291 vdd.n170 gnd 0.009949f
C2292 vdd.t140 gnd 0.034855f
C2293 vdd.t22 gnd 0.034855f
C2294 vdd.n171 gnd 0.239545f
C2295 vdd.n172 gnd 0.188365f
C2296 vdd.t80 gnd 0.034855f
C2297 vdd.t82 gnd 0.034855f
C2298 vdd.n173 gnd 0.239545f
C2299 vdd.n174 gnd 0.15201f
C2300 vdd.t162 gnd 0.034855f
C2301 vdd.t69 gnd 0.034855f
C2302 vdd.n175 gnd 0.239545f
C2303 vdd.n176 gnd 0.15201f
C2304 vdd.t70 gnd 0.034855f
C2305 vdd.t160 gnd 0.034855f
C2306 vdd.n177 gnd 0.239545f
C2307 vdd.n178 gnd 0.15201f
C2308 vdd.t161 gnd 0.034855f
C2309 vdd.t40 gnd 0.034855f
C2310 vdd.n179 gnd 0.239545f
C2311 vdd.n180 gnd 0.15201f
C2312 vdd.t143 gnd 0.034855f
C2313 vdd.t157 gnd 0.034855f
C2314 vdd.n181 gnd 0.239545f
C2315 vdd.n182 gnd 0.15201f
C2316 vdd.t36 gnd 0.034855f
C2317 vdd.t106 gnd 0.034855f
C2318 vdd.n183 gnd 0.239545f
C2319 vdd.n184 gnd 0.15201f
C2320 vdd.t138 gnd 0.034855f
C2321 vdd.t169 gnd 0.034855f
C2322 vdd.n185 gnd 0.239545f
C2323 vdd.n186 gnd 0.15201f
C2324 vdd.t78 gnd 0.034855f
C2325 vdd.t137 gnd 0.034855f
C2326 vdd.n187 gnd 0.239545f
C2327 vdd.n188 gnd 0.15201f
C2328 vdd.n189 gnd 0.005941f
C2329 vdd.n190 gnd 0.005513f
C2330 vdd.n191 gnd 0.00305f
C2331 vdd.n192 gnd 0.007003f
C2332 vdd.n193 gnd 0.002963f
C2333 vdd.n194 gnd 0.003137f
C2334 vdd.n195 gnd 0.005513f
C2335 vdd.n196 gnd 0.002963f
C2336 vdd.n197 gnd 0.007003f
C2337 vdd.n198 gnd 0.003137f
C2338 vdd.n199 gnd 0.005513f
C2339 vdd.n200 gnd 0.002963f
C2340 vdd.n201 gnd 0.005252f
C2341 vdd.n202 gnd 0.005268f
C2342 vdd.t174 gnd 0.015044f
C2343 vdd.n203 gnd 0.033474f
C2344 vdd.n204 gnd 0.174205f
C2345 vdd.n205 gnd 0.002963f
C2346 vdd.n206 gnd 0.003137f
C2347 vdd.n207 gnd 0.007003f
C2348 vdd.n208 gnd 0.007003f
C2349 vdd.n209 gnd 0.003137f
C2350 vdd.n210 gnd 0.002963f
C2351 vdd.n211 gnd 0.005513f
C2352 vdd.n212 gnd 0.005513f
C2353 vdd.n213 gnd 0.002963f
C2354 vdd.n214 gnd 0.003137f
C2355 vdd.n215 gnd 0.007003f
C2356 vdd.n216 gnd 0.007003f
C2357 vdd.n217 gnd 0.003137f
C2358 vdd.n218 gnd 0.002963f
C2359 vdd.n219 gnd 0.005513f
C2360 vdd.n220 gnd 0.005513f
C2361 vdd.n221 gnd 0.002963f
C2362 vdd.n222 gnd 0.003137f
C2363 vdd.n223 gnd 0.007003f
C2364 vdd.n224 gnd 0.007003f
C2365 vdd.n225 gnd 0.016556f
C2366 vdd.n226 gnd 0.00305f
C2367 vdd.n227 gnd 0.002963f
C2368 vdd.n228 gnd 0.01425f
C2369 vdd.n229 gnd 0.009637f
C2370 vdd.n230 gnd 0.067281f
C2371 vdd.n231 gnd 0.24243f
C2372 vdd.n232 gnd 0.005941f
C2373 vdd.n233 gnd 0.005513f
C2374 vdd.n234 gnd 0.00305f
C2375 vdd.n235 gnd 0.007003f
C2376 vdd.n236 gnd 0.002963f
C2377 vdd.n237 gnd 0.003137f
C2378 vdd.n238 gnd 0.005513f
C2379 vdd.n239 gnd 0.002963f
C2380 vdd.n240 gnd 0.007003f
C2381 vdd.n241 gnd 0.003137f
C2382 vdd.n242 gnd 0.005513f
C2383 vdd.n243 gnd 0.002963f
C2384 vdd.n244 gnd 0.005252f
C2385 vdd.n245 gnd 0.005268f
C2386 vdd.t124 gnd 0.015044f
C2387 vdd.n246 gnd 0.033474f
C2388 vdd.n247 gnd 0.174205f
C2389 vdd.n248 gnd 0.002963f
C2390 vdd.n249 gnd 0.003137f
C2391 vdd.n250 gnd 0.007003f
C2392 vdd.n251 gnd 0.007003f
C2393 vdd.n252 gnd 0.003137f
C2394 vdd.n253 gnd 0.002963f
C2395 vdd.n254 gnd 0.005513f
C2396 vdd.n255 gnd 0.005513f
C2397 vdd.n256 gnd 0.002963f
C2398 vdd.n257 gnd 0.003137f
C2399 vdd.n258 gnd 0.007003f
C2400 vdd.n259 gnd 0.007003f
C2401 vdd.n260 gnd 0.003137f
C2402 vdd.n261 gnd 0.002963f
C2403 vdd.n262 gnd 0.005513f
C2404 vdd.n263 gnd 0.005513f
C2405 vdd.n264 gnd 0.002963f
C2406 vdd.n265 gnd 0.003137f
C2407 vdd.n266 gnd 0.007003f
C2408 vdd.n267 gnd 0.007003f
C2409 vdd.n268 gnd 0.016556f
C2410 vdd.n269 gnd 0.00305f
C2411 vdd.n270 gnd 0.002963f
C2412 vdd.n271 gnd 0.01425f
C2413 vdd.n272 gnd 0.009949f
C2414 vdd.t151 gnd 0.034855f
C2415 vdd.t46 gnd 0.034855f
C2416 vdd.n273 gnd 0.239545f
C2417 vdd.n274 gnd 0.188365f
C2418 vdd.t100 gnd 0.034855f
C2419 vdd.t103 gnd 0.034855f
C2420 vdd.n275 gnd 0.239545f
C2421 vdd.n276 gnd 0.15201f
C2422 vdd.t173 gnd 0.034855f
C2423 vdd.t94 gnd 0.034855f
C2424 vdd.n277 gnd 0.239545f
C2425 vdd.n278 gnd 0.15201f
C2426 vdd.t95 gnd 0.034855f
C2427 vdd.t171 gnd 0.034855f
C2428 vdd.n279 gnd 0.239545f
C2429 vdd.n280 gnd 0.15201f
C2430 vdd.t172 gnd 0.034855f
C2431 vdd.t62 gnd 0.034855f
C2432 vdd.n281 gnd 0.239545f
C2433 vdd.n282 gnd 0.15201f
C2434 vdd.t156 gnd 0.034855f
C2435 vdd.t167 gnd 0.034855f
C2436 vdd.n283 gnd 0.239545f
C2437 vdd.n284 gnd 0.15201f
C2438 vdd.t55 gnd 0.034855f
C2439 vdd.t125 gnd 0.034855f
C2440 vdd.n285 gnd 0.239545f
C2441 vdd.n286 gnd 0.15201f
C2442 vdd.t152 gnd 0.034855f
C2443 vdd.t20 gnd 0.034855f
C2444 vdd.n287 gnd 0.239545f
C2445 vdd.n288 gnd 0.15201f
C2446 vdd.t101 gnd 0.034855f
C2447 vdd.t149 gnd 0.034855f
C2448 vdd.n289 gnd 0.239545f
C2449 vdd.n290 gnd 0.15201f
C2450 vdd.n291 gnd 0.005941f
C2451 vdd.n292 gnd 0.005513f
C2452 vdd.n293 gnd 0.00305f
C2453 vdd.n294 gnd 0.007003f
C2454 vdd.n295 gnd 0.002963f
C2455 vdd.n296 gnd 0.003137f
C2456 vdd.n297 gnd 0.005513f
C2457 vdd.n298 gnd 0.002963f
C2458 vdd.n299 gnd 0.007003f
C2459 vdd.n300 gnd 0.003137f
C2460 vdd.n301 gnd 0.005513f
C2461 vdd.n302 gnd 0.002963f
C2462 vdd.n303 gnd 0.005252f
C2463 vdd.n304 gnd 0.005268f
C2464 vdd.t38 gnd 0.015044f
C2465 vdd.n305 gnd 0.033474f
C2466 vdd.n306 gnd 0.174205f
C2467 vdd.n307 gnd 0.002963f
C2468 vdd.n308 gnd 0.003137f
C2469 vdd.n309 gnd 0.007003f
C2470 vdd.n310 gnd 0.007003f
C2471 vdd.n311 gnd 0.003137f
C2472 vdd.n312 gnd 0.002963f
C2473 vdd.n313 gnd 0.005513f
C2474 vdd.n314 gnd 0.005513f
C2475 vdd.n315 gnd 0.002963f
C2476 vdd.n316 gnd 0.003137f
C2477 vdd.n317 gnd 0.007003f
C2478 vdd.n318 gnd 0.007003f
C2479 vdd.n319 gnd 0.003137f
C2480 vdd.n320 gnd 0.002963f
C2481 vdd.n321 gnd 0.005513f
C2482 vdd.n322 gnd 0.005513f
C2483 vdd.n323 gnd 0.002963f
C2484 vdd.n324 gnd 0.003137f
C2485 vdd.n325 gnd 0.007003f
C2486 vdd.n326 gnd 0.007003f
C2487 vdd.n327 gnd 0.016556f
C2488 vdd.n328 gnd 0.00305f
C2489 vdd.n329 gnd 0.002963f
C2490 vdd.n330 gnd 0.01425f
C2491 vdd.n331 gnd 0.009637f
C2492 vdd.n332 gnd 0.067281f
C2493 vdd.n333 gnd 0.27753f
C2494 vdd.n334 gnd 0.00832f
C2495 vdd.n335 gnd 0.010826f
C2496 vdd.n336 gnd 0.008714f
C2497 vdd.n337 gnd 0.008714f
C2498 vdd.n338 gnd 0.010826f
C2499 vdd.n339 gnd 0.010826f
C2500 vdd.n340 gnd 0.791054f
C2501 vdd.n341 gnd 0.010826f
C2502 vdd.n342 gnd 0.010826f
C2503 vdd.n343 gnd 0.010826f
C2504 vdd.n344 gnd 0.857436f
C2505 vdd.n345 gnd 0.010826f
C2506 vdd.n346 gnd 0.010826f
C2507 vdd.n347 gnd 0.010826f
C2508 vdd.n348 gnd 0.010826f
C2509 vdd.n349 gnd 0.008714f
C2510 vdd.n350 gnd 0.010826f
C2511 vdd.t130 gnd 0.553185f
C2512 vdd.n351 gnd 0.010826f
C2513 vdd.n352 gnd 0.010826f
C2514 vdd.n353 gnd 0.010826f
C2515 vdd.t105 gnd 0.553185f
C2516 vdd.n354 gnd 0.010826f
C2517 vdd.n355 gnd 0.010826f
C2518 vdd.n356 gnd 0.010826f
C2519 vdd.n357 gnd 0.010826f
C2520 vdd.n358 gnd 0.010826f
C2521 vdd.n359 gnd 0.008714f
C2522 vdd.n360 gnd 0.010826f
C2523 vdd.n361 gnd 0.625099f
C2524 vdd.n362 gnd 0.010826f
C2525 vdd.n363 gnd 0.010826f
C2526 vdd.n364 gnd 0.010826f
C2527 vdd.t19 gnd 0.553185f
C2528 vdd.n365 gnd 0.010826f
C2529 vdd.n366 gnd 0.010826f
C2530 vdd.n367 gnd 0.010826f
C2531 vdd.n368 gnd 0.010826f
C2532 vdd.n369 gnd 0.010826f
C2533 vdd.n370 gnd 0.008714f
C2534 vdd.n371 gnd 0.010826f
C2535 vdd.t77 gnd 0.553185f
C2536 vdd.n372 gnd 0.010826f
C2537 vdd.n373 gnd 0.010826f
C2538 vdd.n374 gnd 0.010826f
C2539 vdd.n375 gnd 0.647226f
C2540 vdd.n376 gnd 0.010826f
C2541 vdd.n377 gnd 0.010826f
C2542 vdd.n378 gnd 0.010826f
C2543 vdd.n379 gnd 0.010826f
C2544 vdd.n380 gnd 0.010826f
C2545 vdd.n381 gnd 0.008714f
C2546 vdd.n382 gnd 0.010826f
C2547 vdd.t37 gnd 0.553185f
C2548 vdd.n383 gnd 0.010826f
C2549 vdd.n384 gnd 0.010826f
C2550 vdd.n385 gnd 0.010826f
C2551 vdd.n386 gnd 0.558717f
C2552 vdd.n387 gnd 0.010826f
C2553 vdd.n388 gnd 0.010826f
C2554 vdd.n389 gnd 0.010826f
C2555 vdd.n390 gnd 0.010826f
C2556 vdd.n391 gnd 0.026189f
C2557 vdd.n392 gnd 0.02675f
C2558 vdd.t240 gnd 0.553185f
C2559 vdd.n393 gnd 0.026189f
C2560 vdd.n425 gnd 0.010826f
C2561 vdd.t252 gnd 0.133189f
C2562 vdd.t251 gnd 0.142342f
C2563 vdd.t250 gnd 0.173943f
C2564 vdd.n426 gnd 0.22297f
C2565 vdd.n427 gnd 0.188206f
C2566 vdd.n428 gnd 0.01429f
C2567 vdd.n429 gnd 0.010826f
C2568 vdd.n430 gnd 0.008714f
C2569 vdd.n431 gnd 0.010826f
C2570 vdd.n432 gnd 0.008714f
C2571 vdd.n433 gnd 0.010826f
C2572 vdd.n434 gnd 0.008714f
C2573 vdd.n435 gnd 0.010826f
C2574 vdd.n436 gnd 0.008714f
C2575 vdd.n437 gnd 0.010826f
C2576 vdd.n438 gnd 0.008714f
C2577 vdd.n439 gnd 0.010826f
C2578 vdd.t242 gnd 0.133189f
C2579 vdd.t241 gnd 0.142342f
C2580 vdd.t239 gnd 0.173943f
C2581 vdd.n440 gnd 0.22297f
C2582 vdd.n441 gnd 0.188206f
C2583 vdd.n442 gnd 0.008714f
C2584 vdd.n443 gnd 0.010826f
C2585 vdd.n444 gnd 0.008714f
C2586 vdd.n445 gnd 0.010826f
C2587 vdd.n446 gnd 0.008714f
C2588 vdd.n447 gnd 0.010826f
C2589 vdd.n448 gnd 0.008714f
C2590 vdd.n449 gnd 0.010826f
C2591 vdd.n450 gnd 0.008714f
C2592 vdd.n451 gnd 0.010826f
C2593 vdd.t259 gnd 0.133189f
C2594 vdd.t258 gnd 0.142342f
C2595 vdd.t257 gnd 0.173943f
C2596 vdd.n452 gnd 0.22297f
C2597 vdd.n453 gnd 0.188206f
C2598 vdd.n454 gnd 0.018647f
C2599 vdd.n455 gnd 0.010826f
C2600 vdd.n456 gnd 0.008714f
C2601 vdd.n457 gnd 0.010826f
C2602 vdd.n458 gnd 0.008714f
C2603 vdd.n459 gnd 0.010826f
C2604 vdd.n460 gnd 0.008714f
C2605 vdd.n461 gnd 0.010826f
C2606 vdd.n462 gnd 0.008714f
C2607 vdd.n463 gnd 0.010826f
C2608 vdd.n464 gnd 0.02675f
C2609 vdd.n465 gnd 0.007232f
C2610 vdd.n466 gnd 0.008714f
C2611 vdd.n467 gnd 0.010826f
C2612 vdd.n468 gnd 0.010826f
C2613 vdd.n469 gnd 0.008714f
C2614 vdd.n470 gnd 0.010826f
C2615 vdd.n471 gnd 0.010826f
C2616 vdd.n472 gnd 0.010826f
C2617 vdd.n473 gnd 0.010826f
C2618 vdd.n474 gnd 0.010826f
C2619 vdd.n475 gnd 0.008714f
C2620 vdd.n476 gnd 0.008714f
C2621 vdd.n477 gnd 0.010826f
C2622 vdd.n478 gnd 0.010826f
C2623 vdd.n479 gnd 0.008714f
C2624 vdd.n480 gnd 0.010826f
C2625 vdd.n481 gnd 0.010826f
C2626 vdd.n482 gnd 0.010826f
C2627 vdd.n483 gnd 0.010826f
C2628 vdd.n484 gnd 0.010826f
C2629 vdd.n485 gnd 0.008714f
C2630 vdd.n486 gnd 0.008714f
C2631 vdd.n487 gnd 0.010826f
C2632 vdd.n488 gnd 0.010826f
C2633 vdd.n489 gnd 0.008714f
C2634 vdd.n490 gnd 0.010826f
C2635 vdd.n491 gnd 0.010826f
C2636 vdd.n492 gnd 0.010826f
C2637 vdd.n493 gnd 0.010826f
C2638 vdd.n494 gnd 0.010826f
C2639 vdd.n495 gnd 0.008714f
C2640 vdd.n496 gnd 0.008714f
C2641 vdd.n497 gnd 0.010826f
C2642 vdd.n498 gnd 0.010826f
C2643 vdd.n499 gnd 0.008714f
C2644 vdd.n500 gnd 0.010826f
C2645 vdd.n501 gnd 0.010826f
C2646 vdd.n502 gnd 0.010826f
C2647 vdd.n503 gnd 0.010826f
C2648 vdd.n504 gnd 0.010826f
C2649 vdd.n505 gnd 0.008714f
C2650 vdd.n506 gnd 0.008714f
C2651 vdd.n507 gnd 0.010826f
C2652 vdd.n508 gnd 0.010826f
C2653 vdd.n509 gnd 0.007276f
C2654 vdd.n510 gnd 0.010826f
C2655 vdd.n511 gnd 0.010826f
C2656 vdd.n512 gnd 0.010826f
C2657 vdd.n513 gnd 0.010826f
C2658 vdd.n514 gnd 0.010826f
C2659 vdd.n515 gnd 0.007276f
C2660 vdd.n516 gnd 0.008714f
C2661 vdd.n517 gnd 0.010826f
C2662 vdd.n518 gnd 0.010826f
C2663 vdd.n519 gnd 0.008714f
C2664 vdd.n520 gnd 0.010826f
C2665 vdd.n521 gnd 0.010826f
C2666 vdd.n522 gnd 0.010826f
C2667 vdd.n523 gnd 0.010826f
C2668 vdd.n524 gnd 0.010826f
C2669 vdd.n525 gnd 0.008714f
C2670 vdd.n526 gnd 0.008714f
C2671 vdd.n527 gnd 0.010826f
C2672 vdd.n528 gnd 0.010826f
C2673 vdd.n529 gnd 0.008714f
C2674 vdd.n530 gnd 0.010826f
C2675 vdd.n531 gnd 0.010826f
C2676 vdd.n532 gnd 0.010826f
C2677 vdd.n533 gnd 0.010826f
C2678 vdd.n534 gnd 0.010826f
C2679 vdd.n535 gnd 0.008714f
C2680 vdd.n536 gnd 0.008714f
C2681 vdd.n537 gnd 0.010826f
C2682 vdd.n538 gnd 0.010826f
C2683 vdd.n539 gnd 0.008714f
C2684 vdd.n540 gnd 0.010826f
C2685 vdd.n541 gnd 0.010826f
C2686 vdd.n542 gnd 0.010826f
C2687 vdd.n543 gnd 0.010826f
C2688 vdd.n544 gnd 0.010826f
C2689 vdd.n545 gnd 0.008714f
C2690 vdd.n546 gnd 0.008714f
C2691 vdd.n547 gnd 0.010826f
C2692 vdd.n548 gnd 0.010826f
C2693 vdd.n549 gnd 0.008714f
C2694 vdd.n550 gnd 0.010826f
C2695 vdd.n551 gnd 0.010826f
C2696 vdd.n552 gnd 0.010826f
C2697 vdd.n553 gnd 0.010826f
C2698 vdd.n554 gnd 0.010826f
C2699 vdd.n555 gnd 0.008714f
C2700 vdd.n556 gnd 0.008714f
C2701 vdd.n557 gnd 0.010826f
C2702 vdd.n558 gnd 0.010826f
C2703 vdd.n559 gnd 0.008714f
C2704 vdd.n560 gnd 0.010826f
C2705 vdd.n561 gnd 0.010826f
C2706 vdd.n562 gnd 0.010826f
C2707 vdd.n563 gnd 0.010826f
C2708 vdd.n564 gnd 0.010826f
C2709 vdd.n565 gnd 0.005925f
C2710 vdd.n566 gnd 0.018647f
C2711 vdd.n567 gnd 0.010826f
C2712 vdd.n568 gnd 0.010826f
C2713 vdd.n569 gnd 0.008627f
C2714 vdd.n570 gnd 0.010826f
C2715 vdd.n571 gnd 0.010826f
C2716 vdd.n572 gnd 0.010826f
C2717 vdd.n573 gnd 0.010826f
C2718 vdd.n574 gnd 0.010826f
C2719 vdd.n575 gnd 0.008714f
C2720 vdd.n576 gnd 0.008714f
C2721 vdd.n577 gnd 0.010826f
C2722 vdd.n578 gnd 0.010826f
C2723 vdd.n579 gnd 0.008714f
C2724 vdd.n580 gnd 0.010826f
C2725 vdd.n581 gnd 0.010826f
C2726 vdd.n582 gnd 0.010826f
C2727 vdd.n583 gnd 0.010826f
C2728 vdd.n584 gnd 0.010826f
C2729 vdd.n585 gnd 0.008714f
C2730 vdd.n586 gnd 0.008714f
C2731 vdd.n587 gnd 0.010826f
C2732 vdd.n588 gnd 0.010826f
C2733 vdd.n589 gnd 0.008714f
C2734 vdd.n590 gnd 0.010826f
C2735 vdd.n591 gnd 0.010826f
C2736 vdd.n592 gnd 0.010826f
C2737 vdd.n593 gnd 0.010826f
C2738 vdd.n594 gnd 0.010826f
C2739 vdd.n595 gnd 0.008714f
C2740 vdd.n596 gnd 0.008714f
C2741 vdd.n597 gnd 0.010826f
C2742 vdd.n598 gnd 0.010826f
C2743 vdd.n599 gnd 0.008714f
C2744 vdd.n600 gnd 0.010826f
C2745 vdd.n601 gnd 0.010826f
C2746 vdd.n602 gnd 0.010826f
C2747 vdd.n603 gnd 0.010826f
C2748 vdd.n604 gnd 0.010826f
C2749 vdd.n605 gnd 0.008714f
C2750 vdd.n606 gnd 0.008714f
C2751 vdd.n607 gnd 0.010826f
C2752 vdd.n608 gnd 0.010826f
C2753 vdd.n609 gnd 0.008714f
C2754 vdd.n610 gnd 0.010826f
C2755 vdd.n611 gnd 0.010826f
C2756 vdd.n612 gnd 0.010826f
C2757 vdd.n613 gnd 0.010826f
C2758 vdd.n614 gnd 0.010826f
C2759 vdd.n615 gnd 0.008714f
C2760 vdd.n616 gnd 0.010826f
C2761 vdd.n617 gnd 0.008714f
C2762 vdd.n618 gnd 0.004575f
C2763 vdd.n619 gnd 0.010826f
C2764 vdd.n620 gnd 0.010826f
C2765 vdd.n621 gnd 0.008714f
C2766 vdd.n622 gnd 0.010826f
C2767 vdd.n623 gnd 0.008714f
C2768 vdd.n624 gnd 0.010826f
C2769 vdd.n625 gnd 0.008714f
C2770 vdd.n626 gnd 0.010826f
C2771 vdd.n627 gnd 0.008714f
C2772 vdd.n628 gnd 0.010826f
C2773 vdd.n629 gnd 0.008714f
C2774 vdd.n630 gnd 0.010826f
C2775 vdd.n631 gnd 0.008714f
C2776 vdd.n632 gnd 0.010826f
C2777 vdd.n633 gnd 0.602971f
C2778 vdd.t71 gnd 0.553185f
C2779 vdd.n634 gnd 0.010826f
C2780 vdd.n635 gnd 0.008714f
C2781 vdd.n636 gnd 0.010826f
C2782 vdd.n637 gnd 0.008714f
C2783 vdd.n638 gnd 0.010826f
C2784 vdd.t41 gnd 0.553185f
C2785 vdd.n639 gnd 0.010826f
C2786 vdd.n640 gnd 0.008714f
C2787 vdd.n641 gnd 0.010826f
C2788 vdd.n642 gnd 0.008714f
C2789 vdd.n643 gnd 0.010826f
C2790 vdd.t68 gnd 0.553185f
C2791 vdd.n644 gnd 0.691481f
C2792 vdd.n645 gnd 0.010826f
C2793 vdd.n646 gnd 0.008714f
C2794 vdd.n647 gnd 0.010826f
C2795 vdd.n648 gnd 0.008714f
C2796 vdd.n649 gnd 0.010826f
C2797 vdd.t29 gnd 0.553185f
C2798 vdd.n650 gnd 0.010826f
C2799 vdd.n651 gnd 0.008714f
C2800 vdd.n652 gnd 0.010826f
C2801 vdd.n653 gnd 0.008714f
C2802 vdd.n654 gnd 0.010826f
C2803 vdd.n655 gnd 0.768927f
C2804 vdd.n656 gnd 0.918287f
C2805 vdd.t81 gnd 0.553185f
C2806 vdd.n657 gnd 0.010826f
C2807 vdd.n658 gnd 0.008714f
C2808 vdd.n659 gnd 0.010826f
C2809 vdd.n660 gnd 0.008714f
C2810 vdd.n661 gnd 0.010826f
C2811 vdd.n662 gnd 0.580844f
C2812 vdd.n663 gnd 0.010826f
C2813 vdd.n664 gnd 0.008714f
C2814 vdd.n665 gnd 0.010826f
C2815 vdd.n666 gnd 0.008714f
C2816 vdd.n667 gnd 0.010826f
C2817 vdd.t139 gnd 0.553185f
C2818 vdd.t21 gnd 0.553185f
C2819 vdd.n668 gnd 0.010826f
C2820 vdd.n669 gnd 0.008714f
C2821 vdd.n670 gnd 0.010826f
C2822 vdd.n671 gnd 0.008714f
C2823 vdd.n672 gnd 0.010826f
C2824 vdd.t63 gnd 0.553185f
C2825 vdd.n673 gnd 0.010826f
C2826 vdd.n674 gnd 0.008714f
C2827 vdd.n675 gnd 0.010826f
C2828 vdd.n676 gnd 0.008714f
C2829 vdd.n677 gnd 0.010826f
C2830 vdd.n678 gnd 1.10637f
C2831 vdd.n679 gnd 0.901691f
C2832 vdd.n680 gnd 0.010826f
C2833 vdd.n681 gnd 0.008714f
C2834 vdd.n682 gnd 0.026189f
C2835 vdd.n683 gnd 0.007232f
C2836 vdd.n684 gnd 0.026189f
C2837 vdd.t226 gnd 0.553185f
C2838 vdd.n685 gnd 0.026189f
C2839 vdd.n686 gnd 0.007232f
C2840 vdd.n687 gnd 0.00931f
C2841 vdd.t227 gnd 0.133189f
C2842 vdd.t228 gnd 0.142342f
C2843 vdd.t225 gnd 0.173943f
C2844 vdd.n688 gnd 0.22297f
C2845 vdd.n689 gnd 0.187335f
C2846 vdd.n690 gnd 0.013419f
C2847 vdd.n691 gnd 0.010826f
C2848 vdd.n692 gnd 9.43733f
C2849 vdd.n723 gnd 1.52126f
C2850 vdd.n724 gnd 0.010826f
C2851 vdd.n725 gnd 0.010826f
C2852 vdd.n726 gnd 0.02675f
C2853 vdd.n727 gnd 0.00931f
C2854 vdd.n728 gnd 0.010826f
C2855 vdd.n729 gnd 0.008714f
C2856 vdd.n730 gnd 0.006929f
C2857 vdd.n731 gnd 0.025283f
C2858 vdd.n732 gnd 0.008714f
C2859 vdd.n733 gnd 0.010826f
C2860 vdd.n734 gnd 0.010826f
C2861 vdd.n735 gnd 0.010826f
C2862 vdd.n736 gnd 0.010826f
C2863 vdd.n737 gnd 0.010826f
C2864 vdd.n738 gnd 0.010826f
C2865 vdd.n739 gnd 0.010826f
C2866 vdd.n740 gnd 0.010826f
C2867 vdd.n741 gnd 0.010826f
C2868 vdd.n742 gnd 0.010826f
C2869 vdd.n743 gnd 0.010826f
C2870 vdd.n744 gnd 0.010826f
C2871 vdd.n745 gnd 0.010826f
C2872 vdd.n746 gnd 0.010826f
C2873 vdd.n747 gnd 0.007276f
C2874 vdd.n748 gnd 0.010826f
C2875 vdd.n749 gnd 0.010826f
C2876 vdd.n750 gnd 0.010826f
C2877 vdd.n751 gnd 0.010826f
C2878 vdd.n752 gnd 0.010826f
C2879 vdd.n753 gnd 0.010826f
C2880 vdd.n754 gnd 0.010826f
C2881 vdd.n755 gnd 0.010826f
C2882 vdd.n756 gnd 0.010826f
C2883 vdd.n757 gnd 0.010826f
C2884 vdd.n758 gnd 0.010826f
C2885 vdd.n759 gnd 0.010826f
C2886 vdd.n760 gnd 0.010826f
C2887 vdd.n761 gnd 0.010826f
C2888 vdd.n762 gnd 0.010826f
C2889 vdd.n763 gnd 0.010826f
C2890 vdd.n764 gnd 0.010826f
C2891 vdd.n765 gnd 0.010826f
C2892 vdd.n766 gnd 0.010826f
C2893 vdd.n767 gnd 0.008627f
C2894 vdd.t234 gnd 0.133189f
C2895 vdd.t235 gnd 0.142342f
C2896 vdd.t233 gnd 0.173943f
C2897 vdd.n768 gnd 0.22297f
C2898 vdd.n769 gnd 0.187335f
C2899 vdd.n770 gnd 0.010826f
C2900 vdd.n771 gnd 0.010826f
C2901 vdd.n772 gnd 0.010826f
C2902 vdd.n773 gnd 0.010826f
C2903 vdd.n774 gnd 0.010826f
C2904 vdd.n775 gnd 0.010826f
C2905 vdd.n776 gnd 0.010826f
C2906 vdd.n777 gnd 0.010826f
C2907 vdd.n778 gnd 0.010826f
C2908 vdd.n779 gnd 0.010826f
C2909 vdd.n780 gnd 0.010826f
C2910 vdd.n781 gnd 0.010826f
C2911 vdd.n782 gnd 0.010826f
C2912 vdd.n783 gnd 0.006929f
C2913 vdd.n785 gnd 0.007362f
C2914 vdd.n786 gnd 0.007362f
C2915 vdd.n787 gnd 0.007362f
C2916 vdd.n788 gnd 0.007362f
C2917 vdd.n789 gnd 0.007362f
C2918 vdd.n790 gnd 0.007362f
C2919 vdd.n792 gnd 0.007362f
C2920 vdd.n793 gnd 0.007362f
C2921 vdd.n795 gnd 0.007362f
C2922 vdd.n796 gnd 0.005359f
C2923 vdd.n798 gnd 0.007362f
C2924 vdd.t220 gnd 0.297485f
C2925 vdd.t219 gnd 0.304513f
C2926 vdd.t217 gnd 0.19421f
C2927 vdd.n799 gnd 0.10496f
C2928 vdd.n800 gnd 0.059537f
C2929 vdd.n801 gnd 0.010521f
C2930 vdd.n802 gnd 0.01704f
C2931 vdd.n804 gnd 0.007362f
C2932 vdd.n805 gnd 0.752331f
C2933 vdd.n806 gnd 0.016126f
C2934 vdd.n807 gnd 0.016126f
C2935 vdd.n808 gnd 0.007362f
C2936 vdd.n809 gnd 0.017219f
C2937 vdd.n810 gnd 0.007362f
C2938 vdd.n811 gnd 0.007362f
C2939 vdd.n812 gnd 0.007362f
C2940 vdd.n813 gnd 0.007362f
C2941 vdd.n814 gnd 0.007362f
C2942 vdd.n816 gnd 0.007362f
C2943 vdd.n817 gnd 0.007362f
C2944 vdd.n819 gnd 0.007362f
C2945 vdd.n820 gnd 0.007362f
C2946 vdd.n822 gnd 0.007362f
C2947 vdd.n823 gnd 0.007362f
C2948 vdd.n825 gnd 0.007362f
C2949 vdd.n826 gnd 0.007362f
C2950 vdd.n828 gnd 0.007362f
C2951 vdd.n829 gnd 0.007362f
C2952 vdd.n831 gnd 0.007362f
C2953 vdd.t292 gnd 0.297485f
C2954 vdd.t291 gnd 0.304513f
C2955 vdd.t290 gnd 0.19421f
C2956 vdd.n832 gnd 0.10496f
C2957 vdd.n833 gnd 0.059537f
C2958 vdd.n834 gnd 0.007362f
C2959 vdd.n836 gnd 0.007362f
C2960 vdd.n837 gnd 0.007362f
C2961 vdd.t218 gnd 0.376166f
C2962 vdd.n838 gnd 0.007362f
C2963 vdd.n839 gnd 0.007362f
C2964 vdd.n840 gnd 0.007362f
C2965 vdd.n841 gnd 0.007362f
C2966 vdd.n842 gnd 0.007362f
C2967 vdd.n843 gnd 0.752331f
C2968 vdd.n844 gnd 0.007362f
C2969 vdd.n845 gnd 0.007362f
C2970 vdd.n846 gnd 0.636162f
C2971 vdd.n847 gnd 0.007362f
C2972 vdd.n848 gnd 0.007362f
C2973 vdd.n849 gnd 0.007362f
C2974 vdd.n850 gnd 0.007362f
C2975 vdd.n851 gnd 0.735736f
C2976 vdd.n852 gnd 0.007362f
C2977 vdd.n853 gnd 0.007362f
C2978 vdd.n854 gnd 0.007362f
C2979 vdd.n855 gnd 0.007362f
C2980 vdd.n856 gnd 0.007362f
C2981 vdd.n857 gnd 0.752331f
C2982 vdd.n858 gnd 0.007362f
C2983 vdd.n859 gnd 0.007362f
C2984 vdd.t11 gnd 0.376166f
C2985 vdd.n860 gnd 0.007362f
C2986 vdd.n861 gnd 0.007362f
C2987 vdd.n862 gnd 0.007362f
C2988 vdd.t208 gnd 0.376166f
C2989 vdd.n863 gnd 0.007362f
C2990 vdd.n864 gnd 0.007362f
C2991 vdd.n865 gnd 0.007362f
C2992 vdd.n866 gnd 0.007362f
C2993 vdd.n867 gnd 0.007362f
C2994 vdd.t244 gnd 0.315315f
C2995 vdd.n868 gnd 0.007362f
C2996 vdd.n869 gnd 0.007362f
C2997 vdd.n870 gnd 0.602971f
C2998 vdd.n871 gnd 0.007362f
C2999 vdd.t245 gnd 0.304513f
C3000 vdd.t243 gnd 0.19421f
C3001 vdd.t246 gnd 0.304513f
C3002 vdd.n872 gnd 0.171149f
C3003 vdd.n873 gnd 0.007362f
C3004 vdd.n874 gnd 0.007362f
C3005 vdd.n875 gnd 0.481271f
C3006 vdd.n876 gnd 0.007362f
C3007 vdd.n877 gnd 0.007362f
C3008 vdd.t215 gnd 0.110637f
C3009 vdd.n878 gnd 0.437016f
C3010 vdd.n879 gnd 0.007362f
C3011 vdd.n880 gnd 0.007362f
C3012 vdd.n881 gnd 0.007362f
C3013 vdd.n882 gnd 0.647226f
C3014 vdd.n883 gnd 0.007362f
C3015 vdd.n884 gnd 0.007362f
C3016 vdd.t1 gnd 0.376166f
C3017 vdd.n885 gnd 0.007362f
C3018 vdd.n886 gnd 0.007362f
C3019 vdd.n887 gnd 0.007362f
C3020 vdd.t189 gnd 0.376166f
C3021 vdd.n888 gnd 0.007362f
C3022 vdd.n889 gnd 0.007362f
C3023 vdd.t205 gnd 0.376166f
C3024 vdd.n890 gnd 0.007362f
C3025 vdd.n891 gnd 0.007362f
C3026 vdd.n892 gnd 0.007362f
C3027 vdd.t198 gnd 0.29872f
C3028 vdd.n893 gnd 0.007362f
C3029 vdd.n894 gnd 0.007362f
C3030 vdd.n895 gnd 0.619567f
C3031 vdd.n896 gnd 0.007362f
C3032 vdd.n897 gnd 0.007362f
C3033 vdd.n898 gnd 0.007362f
C3034 vdd.t14 gnd 0.376166f
C3035 vdd.n899 gnd 0.007362f
C3036 vdd.n900 gnd 0.007362f
C3037 vdd.t187 gnd 0.315315f
C3038 vdd.n901 gnd 0.453611f
C3039 vdd.n902 gnd 0.007362f
C3040 vdd.n903 gnd 0.007362f
C3041 vdd.n904 gnd 0.007362f
C3042 vdd.n905 gnd 0.392761f
C3043 vdd.n906 gnd 0.007362f
C3044 vdd.n907 gnd 0.007362f
C3045 vdd.t201 gnd 0.376166f
C3046 vdd.n908 gnd 0.007362f
C3047 vdd.n909 gnd 0.007362f
C3048 vdd.n910 gnd 0.007362f
C3049 vdd.n911 gnd 0.752331f
C3050 vdd.n912 gnd 0.007362f
C3051 vdd.n913 gnd 0.007362f
C3052 vdd.t216 gnd 0.254465f
C3053 vdd.t211 gnd 0.35957f
C3054 vdd.n914 gnd 0.007362f
C3055 vdd.n915 gnd 0.007362f
C3056 vdd.n916 gnd 0.007362f
C3057 vdd.n917 gnd 0.564248f
C3058 vdd.n918 gnd 0.007362f
C3059 vdd.n919 gnd 0.007362f
C3060 vdd.n920 gnd 0.007362f
C3061 vdd.n921 gnd 0.007362f
C3062 vdd.n922 gnd 0.007362f
C3063 vdd.t268 gnd 0.376166f
C3064 vdd.n923 gnd 0.007362f
C3065 vdd.n924 gnd 0.007362f
C3066 vdd.t298 gnd 0.376166f
C3067 vdd.n925 gnd 0.007362f
C3068 vdd.n926 gnd 0.016126f
C3069 vdd.n927 gnd 0.016126f
C3070 vdd.n928 gnd 0.896159f
C3071 vdd.n929 gnd 0.007362f
C3072 vdd.n930 gnd 0.007362f
C3073 vdd.t194 gnd 0.376166f
C3074 vdd.n931 gnd 0.016126f
C3075 vdd.n932 gnd 0.007362f
C3076 vdd.n933 gnd 0.007362f
C3077 vdd.t199 gnd 0.685949f
C3078 vdd.n951 gnd 0.017219f
C3079 vdd.n969 gnd 0.016126f
C3080 vdd.n970 gnd 0.007362f
C3081 vdd.n971 gnd 0.016126f
C3082 vdd.t289 gnd 0.297485f
C3083 vdd.t288 gnd 0.304513f
C3084 vdd.t287 gnd 0.19421f
C3085 vdd.n972 gnd 0.10496f
C3086 vdd.n973 gnd 0.059537f
C3087 vdd.n974 gnd 0.01704f
C3088 vdd.n975 gnd 0.007362f
C3089 vdd.n976 gnd 0.398293f
C3090 vdd.n977 gnd 0.016126f
C3091 vdd.n978 gnd 0.007362f
C3092 vdd.n979 gnd 0.017219f
C3093 vdd.n980 gnd 0.007362f
C3094 vdd.t266 gnd 0.297485f
C3095 vdd.t265 gnd 0.304513f
C3096 vdd.t263 gnd 0.19421f
C3097 vdd.n981 gnd 0.10496f
C3098 vdd.n982 gnd 0.059537f
C3099 vdd.n983 gnd 0.010521f
C3100 vdd.n984 gnd 0.007362f
C3101 vdd.n985 gnd 0.007362f
C3102 vdd.t264 gnd 0.376166f
C3103 vdd.n986 gnd 0.007362f
C3104 vdd.t206 gnd 0.376166f
C3105 vdd.n987 gnd 0.007362f
C3106 vdd.n988 gnd 0.007362f
C3107 vdd.n989 gnd 0.007362f
C3108 vdd.n990 gnd 0.007362f
C3109 vdd.n991 gnd 0.007362f
C3110 vdd.n992 gnd 0.752331f
C3111 vdd.n993 gnd 0.007362f
C3112 vdd.n994 gnd 0.007362f
C3113 vdd.t2 gnd 0.376166f
C3114 vdd.n995 gnd 0.007362f
C3115 vdd.n996 gnd 0.007362f
C3116 vdd.n997 gnd 0.007362f
C3117 vdd.n998 gnd 0.007362f
C3118 vdd.n999 gnd 0.497866f
C3119 vdd.n1000 gnd 0.007362f
C3120 vdd.n1001 gnd 0.007362f
C3121 vdd.n1002 gnd 0.007362f
C3122 vdd.n1003 gnd 0.007362f
C3123 vdd.n1004 gnd 0.007362f
C3124 vdd.n1005 gnd 0.663822f
C3125 vdd.n1006 gnd 0.007362f
C3126 vdd.n1007 gnd 0.007362f
C3127 vdd.t15 gnd 0.35957f
C3128 vdd.t12 gnd 0.254465f
C3129 vdd.n1008 gnd 0.007362f
C3130 vdd.n1009 gnd 0.007362f
C3131 vdd.n1010 gnd 0.007362f
C3132 vdd.t0 gnd 0.376166f
C3133 vdd.n1011 gnd 0.007362f
C3134 vdd.n1012 gnd 0.007362f
C3135 vdd.t296 gnd 0.376166f
C3136 vdd.n1013 gnd 0.007362f
C3137 vdd.n1014 gnd 0.007362f
C3138 vdd.n1015 gnd 0.007362f
C3139 vdd.t213 gnd 0.315315f
C3140 vdd.n1016 gnd 0.007362f
C3141 vdd.n1017 gnd 0.007362f
C3142 vdd.n1018 gnd 0.602971f
C3143 vdd.n1019 gnd 0.007362f
C3144 vdd.n1020 gnd 0.007362f
C3145 vdd.n1021 gnd 0.007362f
C3146 vdd.t203 gnd 0.376166f
C3147 vdd.n1022 gnd 0.007362f
C3148 vdd.n1023 gnd 0.007362f
C3149 vdd.t13 gnd 0.29872f
C3150 vdd.n1024 gnd 0.437016f
C3151 vdd.n1025 gnd 0.007362f
C3152 vdd.n1026 gnd 0.007362f
C3153 vdd.n1027 gnd 0.007362f
C3154 vdd.n1028 gnd 0.647226f
C3155 vdd.n1029 gnd 0.007362f
C3156 vdd.n1030 gnd 0.007362f
C3157 vdd.t10 gnd 0.376166f
C3158 vdd.n1031 gnd 0.007362f
C3159 vdd.n1032 gnd 0.007362f
C3160 vdd.n1033 gnd 0.007362f
C3161 vdd.n1034 gnd 0.752331f
C3162 vdd.n1035 gnd 0.007362f
C3163 vdd.n1036 gnd 0.007362f
C3164 vdd.t191 gnd 0.376166f
C3165 vdd.n1037 gnd 0.007362f
C3166 vdd.n1038 gnd 0.007362f
C3167 vdd.n1039 gnd 0.007362f
C3168 vdd.t179 gnd 0.110637f
C3169 vdd.n1040 gnd 0.007362f
C3170 vdd.n1041 gnd 0.007362f
C3171 vdd.n1042 gnd 0.007362f
C3172 vdd.t276 gnd 0.304513f
C3173 vdd.t274 gnd 0.19421f
C3174 vdd.t277 gnd 0.304513f
C3175 vdd.n1043 gnd 0.171149f
C3176 vdd.n1044 gnd 0.007362f
C3177 vdd.n1045 gnd 0.007362f
C3178 vdd.t180 gnd 0.376166f
C3179 vdd.n1046 gnd 0.007362f
C3180 vdd.n1047 gnd 0.007362f
C3181 vdd.t275 gnd 0.315315f
C3182 vdd.n1048 gnd 0.641694f
C3183 vdd.n1049 gnd 0.007362f
C3184 vdd.n1050 gnd 0.007362f
C3185 vdd.n1051 gnd 0.007362f
C3186 vdd.n1052 gnd 0.392761f
C3187 vdd.n1053 gnd 0.007362f
C3188 vdd.n1054 gnd 0.007362f
C3189 vdd.n1055 gnd 0.525526f
C3190 vdd.n1056 gnd 0.007362f
C3191 vdd.n1057 gnd 0.007362f
C3192 vdd.n1058 gnd 0.007362f
C3193 vdd.n1059 gnd 0.752331f
C3194 vdd.n1060 gnd 0.007362f
C3195 vdd.n1061 gnd 0.007362f
C3196 vdd.t295 gnd 0.376166f
C3197 vdd.n1062 gnd 0.007362f
C3198 vdd.n1063 gnd 0.007362f
C3199 vdd.n1064 gnd 0.007362f
C3200 vdd.n1065 gnd 0.752331f
C3201 vdd.n1066 gnd 0.007362f
C3202 vdd.n1067 gnd 0.007362f
C3203 vdd.n1068 gnd 0.007362f
C3204 vdd.n1069 gnd 0.007362f
C3205 vdd.n1070 gnd 0.007362f
C3206 vdd.t222 gnd 0.376166f
C3207 vdd.n1071 gnd 0.007362f
C3208 vdd.n1072 gnd 0.007362f
C3209 vdd.n1073 gnd 0.007362f
C3210 vdd.n1074 gnd 0.016126f
C3211 vdd.n1075 gnd 0.016126f
C3212 vdd.n1076 gnd 1.06211f
C3213 vdd.n1077 gnd 0.007362f
C3214 vdd.n1078 gnd 0.007362f
C3215 vdd.n1079 gnd 0.492334f
C3216 vdd.n1080 gnd 0.016126f
C3217 vdd.n1081 gnd 0.007362f
C3218 vdd.n1082 gnd 0.007362f
C3219 vdd.n1083 gnd 9.83562f
C3220 vdd.n1116 gnd 0.017219f
C3221 vdd.n1117 gnd 0.007362f
C3222 vdd.n1118 gnd 0.007362f
C3223 vdd.n1119 gnd 0.007362f
C3224 vdd.n1120 gnd 0.006929f
C3225 vdd.n1123 gnd 0.02675f
C3226 vdd.n1124 gnd 0.007232f
C3227 vdd.n1125 gnd 0.008714f
C3228 vdd.n1127 gnd 0.010826f
C3229 vdd.n1128 gnd 0.010826f
C3230 vdd.n1129 gnd 0.008714f
C3231 vdd.n1131 gnd 0.010826f
C3232 vdd.n1132 gnd 0.010826f
C3233 vdd.n1133 gnd 0.010826f
C3234 vdd.n1134 gnd 0.010826f
C3235 vdd.n1135 gnd 0.010826f
C3236 vdd.n1136 gnd 0.008714f
C3237 vdd.n1138 gnd 0.010826f
C3238 vdd.n1139 gnd 0.010826f
C3239 vdd.n1140 gnd 0.010826f
C3240 vdd.n1141 gnd 0.010826f
C3241 vdd.n1142 gnd 0.010826f
C3242 vdd.n1143 gnd 0.008714f
C3243 vdd.n1145 gnd 0.010826f
C3244 vdd.n1146 gnd 0.010826f
C3245 vdd.n1147 gnd 0.010826f
C3246 vdd.n1148 gnd 0.010826f
C3247 vdd.n1149 gnd 0.007276f
C3248 vdd.t280 gnd 0.133189f
C3249 vdd.t279 gnd 0.142342f
C3250 vdd.t278 gnd 0.173943f
C3251 vdd.n1150 gnd 0.22297f
C3252 vdd.n1151 gnd 0.187335f
C3253 vdd.n1153 gnd 0.010826f
C3254 vdd.n1154 gnd 0.010826f
C3255 vdd.n1155 gnd 0.008714f
C3256 vdd.n1156 gnd 0.010826f
C3257 vdd.n1158 gnd 0.010826f
C3258 vdd.n1159 gnd 0.010826f
C3259 vdd.n1160 gnd 0.010826f
C3260 vdd.n1161 gnd 0.010826f
C3261 vdd.n1162 gnd 0.008714f
C3262 vdd.n1164 gnd 0.010826f
C3263 vdd.n1165 gnd 0.010826f
C3264 vdd.n1166 gnd 0.010826f
C3265 vdd.n1167 gnd 0.010826f
C3266 vdd.n1168 gnd 0.010826f
C3267 vdd.n1169 gnd 0.008714f
C3268 vdd.n1171 gnd 0.010826f
C3269 vdd.n1172 gnd 0.010826f
C3270 vdd.n1173 gnd 0.010826f
C3271 vdd.n1174 gnd 0.010826f
C3272 vdd.n1175 gnd 0.010826f
C3273 vdd.n1176 gnd 0.008714f
C3274 vdd.n1178 gnd 0.010826f
C3275 vdd.n1179 gnd 0.010826f
C3276 vdd.n1180 gnd 0.010826f
C3277 vdd.n1181 gnd 0.010826f
C3278 vdd.n1182 gnd 0.010826f
C3279 vdd.n1183 gnd 0.008714f
C3280 vdd.n1185 gnd 0.010826f
C3281 vdd.n1186 gnd 0.010826f
C3282 vdd.n1187 gnd 0.010826f
C3283 vdd.n1188 gnd 0.010826f
C3284 vdd.n1189 gnd 0.008627f
C3285 vdd.t262 gnd 0.133189f
C3286 vdd.t261 gnd 0.142342f
C3287 vdd.t260 gnd 0.173943f
C3288 vdd.n1190 gnd 0.22297f
C3289 vdd.n1191 gnd 0.187335f
C3290 vdd.n1193 gnd 0.010826f
C3291 vdd.n1194 gnd 0.010826f
C3292 vdd.n1195 gnd 0.008714f
C3293 vdd.n1196 gnd 0.010826f
C3294 vdd.n1198 gnd 0.010826f
C3295 vdd.n1199 gnd 0.010826f
C3296 vdd.n1200 gnd 0.010826f
C3297 vdd.n1201 gnd 0.010826f
C3298 vdd.n1202 gnd 0.008714f
C3299 vdd.n1204 gnd 0.010826f
C3300 vdd.n1205 gnd 0.010826f
C3301 vdd.n1206 gnd 0.010826f
C3302 vdd.n1207 gnd 0.010826f
C3303 vdd.n1208 gnd 0.010826f
C3304 vdd.n1209 gnd 0.008714f
C3305 vdd.n1211 gnd 0.010826f
C3306 vdd.n1212 gnd 0.010826f
C3307 vdd.n1213 gnd 0.010826f
C3308 vdd.n1214 gnd 0.010826f
C3309 vdd.n1215 gnd 0.010826f
C3310 vdd.n1216 gnd 0.008714f
C3311 vdd.n1218 gnd 0.010826f
C3312 vdd.n1219 gnd 0.010826f
C3313 vdd.n1220 gnd 0.006929f
C3314 vdd.n1221 gnd 0.008714f
C3315 vdd.n1222 gnd 0.007362f
C3316 vdd.n1223 gnd 0.007362f
C3317 vdd.n1224 gnd 0.007362f
C3318 vdd.n1225 gnd 0.007362f
C3319 vdd.n1226 gnd 0.007362f
C3320 vdd.n1227 gnd 0.007362f
C3321 vdd.n1228 gnd 0.007362f
C3322 vdd.n1229 gnd 0.007362f
C3323 vdd.n1230 gnd 0.007362f
C3324 vdd.n1231 gnd 0.007362f
C3325 vdd.n1232 gnd 0.007362f
C3326 vdd.n1233 gnd 0.007362f
C3327 vdd.n1234 gnd 0.007362f
C3328 vdd.n1235 gnd 0.007362f
C3329 vdd.n1236 gnd 0.007362f
C3330 vdd.n1237 gnd 0.007362f
C3331 vdd.n1238 gnd 0.007362f
C3332 vdd.n1239 gnd 0.007362f
C3333 vdd.n1240 gnd 0.007362f
C3334 vdd.n1241 gnd 0.007362f
C3335 vdd.n1242 gnd 0.007362f
C3336 vdd.n1243 gnd 0.007362f
C3337 vdd.n1244 gnd 0.007362f
C3338 vdd.n1245 gnd 0.007362f
C3339 vdd.n1246 gnd 0.007362f
C3340 vdd.n1247 gnd 0.007362f
C3341 vdd.n1248 gnd 0.007362f
C3342 vdd.n1249 gnd 0.007362f
C3343 vdd.n1250 gnd 0.007362f
C3344 vdd.n1251 gnd 0.007362f
C3345 vdd.n1252 gnd 0.007362f
C3346 vdd.t223 gnd 0.297485f
C3347 vdd.t224 gnd 0.304513f
C3348 vdd.t221 gnd 0.19421f
C3349 vdd.n1253 gnd 0.10496f
C3350 vdd.n1254 gnd 0.059537f
C3351 vdd.n1255 gnd 0.010521f
C3352 vdd.n1256 gnd 0.007362f
C3353 vdd.n1257 gnd 0.007362f
C3354 vdd.n1258 gnd 0.007362f
C3355 vdd.n1259 gnd 0.007362f
C3356 vdd.n1260 gnd 0.007362f
C3357 vdd.n1261 gnd 0.007362f
C3358 vdd.n1262 gnd 0.007362f
C3359 vdd.n1263 gnd 0.007362f
C3360 vdd.n1264 gnd 0.007362f
C3361 vdd.n1265 gnd 0.007362f
C3362 vdd.n1266 gnd 0.007362f
C3363 vdd.n1267 gnd 0.007362f
C3364 vdd.n1268 gnd 0.007362f
C3365 vdd.n1269 gnd 0.007362f
C3366 vdd.n1270 gnd 0.007362f
C3367 vdd.n1271 gnd 0.007362f
C3368 vdd.n1272 gnd 0.007362f
C3369 vdd.t237 gnd 0.297485f
C3370 vdd.t238 gnd 0.304513f
C3371 vdd.t236 gnd 0.19421f
C3372 vdd.n1273 gnd 0.10496f
C3373 vdd.n1274 gnd 0.059537f
C3374 vdd.n1275 gnd 0.007362f
C3375 vdd.n1276 gnd 0.007362f
C3376 vdd.n1277 gnd 0.007362f
C3377 vdd.n1278 gnd 0.007362f
C3378 vdd.n1279 gnd 0.007362f
C3379 vdd.n1280 gnd 0.007362f
C3380 vdd.n1281 gnd 0.007362f
C3381 vdd.n1282 gnd 0.007362f
C3382 vdd.n1283 gnd 0.007362f
C3383 vdd.n1284 gnd 0.007362f
C3384 vdd.n1285 gnd 0.007362f
C3385 vdd.n1286 gnd 0.007362f
C3386 vdd.n1287 gnd 0.007362f
C3387 vdd.n1288 gnd 0.007362f
C3388 vdd.n1289 gnd 0.007362f
C3389 vdd.n1290 gnd 0.007362f
C3390 vdd.n1291 gnd 0.007362f
C3391 vdd.n1292 gnd 0.007362f
C3392 vdd.n1293 gnd 0.007362f
C3393 vdd.n1294 gnd 0.007362f
C3394 vdd.n1295 gnd 0.007362f
C3395 vdd.n1296 gnd 0.007362f
C3396 vdd.n1297 gnd 0.007362f
C3397 vdd.n1298 gnd 0.007362f
C3398 vdd.n1299 gnd 0.007362f
C3399 vdd.n1300 gnd 0.007362f
C3400 vdd.n1301 gnd 0.005359f
C3401 vdd.n1302 gnd 0.010521f
C3402 vdd.n1303 gnd 0.005684f
C3403 vdd.n1304 gnd 0.007362f
C3404 vdd.n1305 gnd 0.007362f
C3405 vdd.n1306 gnd 0.007362f
C3406 vdd.n1307 gnd 0.017219f
C3407 vdd.n1308 gnd 0.017219f
C3408 vdd.n1309 gnd 0.016126f
C3409 vdd.n1310 gnd 0.016126f
C3410 vdd.n1311 gnd 0.007362f
C3411 vdd.n1312 gnd 0.007362f
C3412 vdd.n1313 gnd 0.007362f
C3413 vdd.n1314 gnd 0.007362f
C3414 vdd.n1315 gnd 0.007362f
C3415 vdd.n1316 gnd 0.007362f
C3416 vdd.n1317 gnd 0.007362f
C3417 vdd.n1318 gnd 0.007362f
C3418 vdd.n1319 gnd 0.007362f
C3419 vdd.n1320 gnd 0.007362f
C3420 vdd.n1321 gnd 0.007362f
C3421 vdd.n1322 gnd 0.007362f
C3422 vdd.n1323 gnd 0.007362f
C3423 vdd.n1324 gnd 0.007362f
C3424 vdd.n1325 gnd 0.007362f
C3425 vdd.n1326 gnd 0.007362f
C3426 vdd.n1327 gnd 0.007362f
C3427 vdd.n1328 gnd 0.007362f
C3428 vdd.n1329 gnd 0.007362f
C3429 vdd.n1330 gnd 0.007362f
C3430 vdd.n1331 gnd 0.007362f
C3431 vdd.n1332 gnd 0.007362f
C3432 vdd.n1333 gnd 0.007362f
C3433 vdd.n1334 gnd 0.007362f
C3434 vdd.n1335 gnd 0.007362f
C3435 vdd.n1336 gnd 0.007362f
C3436 vdd.n1337 gnd 0.007362f
C3437 vdd.n1338 gnd 0.44808f
C3438 vdd.n1339 gnd 0.007362f
C3439 vdd.n1340 gnd 0.007362f
C3440 vdd.n1341 gnd 0.007362f
C3441 vdd.n1342 gnd 0.007362f
C3442 vdd.n1343 gnd 0.007362f
C3443 vdd.n1344 gnd 0.007362f
C3444 vdd.n1345 gnd 0.007362f
C3445 vdd.n1346 gnd 0.007362f
C3446 vdd.n1347 gnd 0.007362f
C3447 vdd.n1348 gnd 0.007362f
C3448 vdd.n1349 gnd 0.007362f
C3449 vdd.n1350 gnd 0.007362f
C3450 vdd.n1351 gnd 0.007362f
C3451 vdd.n1352 gnd 0.007362f
C3452 vdd.n1353 gnd 0.007362f
C3453 vdd.n1354 gnd 0.007362f
C3454 vdd.n1355 gnd 0.007362f
C3455 vdd.n1356 gnd 0.007362f
C3456 vdd.n1357 gnd 0.007362f
C3457 vdd.n1358 gnd 0.007362f
C3458 vdd.n1359 gnd 0.237869f
C3459 vdd.n1360 gnd 0.007362f
C3460 vdd.n1361 gnd 0.007362f
C3461 vdd.n1362 gnd 0.007362f
C3462 vdd.n1363 gnd 0.007362f
C3463 vdd.n1364 gnd 0.007362f
C3464 vdd.n1365 gnd 0.007362f
C3465 vdd.n1366 gnd 0.007362f
C3466 vdd.n1367 gnd 0.007362f
C3467 vdd.n1368 gnd 0.007362f
C3468 vdd.n1369 gnd 0.007362f
C3469 vdd.n1370 gnd 0.007362f
C3470 vdd.n1371 gnd 0.007362f
C3471 vdd.n1372 gnd 0.007362f
C3472 vdd.n1373 gnd 0.007362f
C3473 vdd.n1374 gnd 0.007362f
C3474 vdd.n1375 gnd 0.007362f
C3475 vdd.n1376 gnd 0.007362f
C3476 vdd.n1377 gnd 0.007362f
C3477 vdd.n1378 gnd 0.007362f
C3478 vdd.n1379 gnd 0.007362f
C3479 vdd.n1380 gnd 0.007362f
C3480 vdd.n1381 gnd 0.007362f
C3481 vdd.n1382 gnd 0.007362f
C3482 vdd.n1383 gnd 0.007362f
C3483 vdd.n1384 gnd 0.007362f
C3484 vdd.n1385 gnd 0.007362f
C3485 vdd.n1386 gnd 0.007362f
C3486 vdd.n1387 gnd 0.016126f
C3487 vdd.n1388 gnd 0.016126f
C3488 vdd.n1389 gnd 0.017219f
C3489 vdd.n1390 gnd 0.007362f
C3490 vdd.n1391 gnd 0.007362f
C3491 vdd.n1392 gnd 0.005684f
C3492 vdd.n1393 gnd 0.007362f
C3493 vdd.n1394 gnd 0.007362f
C3494 vdd.n1395 gnd 0.005359f
C3495 vdd.n1396 gnd 0.007362f
C3496 vdd.n1397 gnd 0.007362f
C3497 vdd.n1398 gnd 0.007362f
C3498 vdd.n1399 gnd 0.007362f
C3499 vdd.n1400 gnd 0.007362f
C3500 vdd.n1401 gnd 0.007362f
C3501 vdd.n1402 gnd 0.007362f
C3502 vdd.n1403 gnd 0.007362f
C3503 vdd.n1404 gnd 0.007362f
C3504 vdd.n1405 gnd 0.007362f
C3505 vdd.n1406 gnd 0.007362f
C3506 vdd.n1407 gnd 0.007362f
C3507 vdd.n1408 gnd 0.007362f
C3508 vdd.n1409 gnd 0.007362f
C3509 vdd.n1410 gnd 0.007362f
C3510 vdd.n1411 gnd 0.007362f
C3511 vdd.n1412 gnd 0.007362f
C3512 vdd.n1413 gnd 0.007362f
C3513 vdd.n1414 gnd 0.007362f
C3514 vdd.n1415 gnd 0.007362f
C3515 vdd.n1416 gnd 0.007362f
C3516 vdd.n1417 gnd 0.007362f
C3517 vdd.n1418 gnd 0.007362f
C3518 vdd.n1419 gnd 0.007362f
C3519 vdd.n1420 gnd 0.007362f
C3520 vdd.n1421 gnd 0.007362f
C3521 vdd.n1422 gnd 0.029505f
C3522 vdd.n1424 gnd 0.02675f
C3523 vdd.n1425 gnd 0.008714f
C3524 vdd.n1427 gnd 0.010826f
C3525 vdd.n1428 gnd 0.008714f
C3526 vdd.n1429 gnd 0.010826f
C3527 vdd.n1431 gnd 0.010826f
C3528 vdd.n1432 gnd 0.010826f
C3529 vdd.n1434 gnd 0.010826f
C3530 vdd.n1435 gnd 0.007232f
C3531 vdd.t230 gnd 0.553185f
C3532 vdd.n1436 gnd 0.010826f
C3533 vdd.n1437 gnd 0.02675f
C3534 vdd.n1438 gnd 0.008714f
C3535 vdd.n1439 gnd 0.010826f
C3536 vdd.n1440 gnd 0.008714f
C3537 vdd.n1441 gnd 0.010826f
C3538 vdd.n1442 gnd 1.10637f
C3539 vdd.n1443 gnd 0.010826f
C3540 vdd.n1444 gnd 0.008714f
C3541 vdd.n1445 gnd 0.008714f
C3542 vdd.n1446 gnd 0.010826f
C3543 vdd.n1447 gnd 0.008714f
C3544 vdd.n1448 gnd 0.010826f
C3545 vdd.t65 gnd 0.553185f
C3546 vdd.n1449 gnd 0.010826f
C3547 vdd.n1450 gnd 0.008714f
C3548 vdd.n1451 gnd 0.010826f
C3549 vdd.n1452 gnd 0.008714f
C3550 vdd.n1453 gnd 0.010826f
C3551 vdd.t25 gnd 0.553185f
C3552 vdd.n1454 gnd 0.010826f
C3553 vdd.n1455 gnd 0.008714f
C3554 vdd.n1456 gnd 0.010826f
C3555 vdd.n1457 gnd 0.008714f
C3556 vdd.n1458 gnd 0.010826f
C3557 vdd.n1459 gnd 0.890627f
C3558 vdd.n1460 gnd 0.918287f
C3559 vdd.t97 gnd 0.553185f
C3560 vdd.n1461 gnd 0.010826f
C3561 vdd.n1462 gnd 0.008714f
C3562 vdd.n1463 gnd 0.010826f
C3563 vdd.n1464 gnd 0.008714f
C3564 vdd.n1465 gnd 0.010826f
C3565 vdd.n1466 gnd 0.702545f
C3566 vdd.n1467 gnd 0.010826f
C3567 vdd.n1468 gnd 0.008714f
C3568 vdd.n1469 gnd 0.010826f
C3569 vdd.n1470 gnd 0.008714f
C3570 vdd.n1471 gnd 0.010826f
C3571 vdd.t33 gnd 0.553185f
C3572 vdd.t121 gnd 0.553185f
C3573 vdd.n1472 gnd 0.010826f
C3574 vdd.n1473 gnd 0.008714f
C3575 vdd.n1474 gnd 0.010826f
C3576 vdd.n1475 gnd 0.008714f
C3577 vdd.n1476 gnd 0.010826f
C3578 vdd.t85 gnd 0.553185f
C3579 vdd.n1477 gnd 0.010826f
C3580 vdd.n1478 gnd 0.008714f
C3581 vdd.n1479 gnd 0.010826f
C3582 vdd.n1480 gnd 0.008714f
C3583 vdd.n1481 gnd 0.010826f
C3584 vdd.t44 gnd 0.553185f
C3585 vdd.n1482 gnd 0.77999f
C3586 vdd.n1483 gnd 0.010826f
C3587 vdd.n1484 gnd 0.008714f
C3588 vdd.n1485 gnd 0.010826f
C3589 vdd.n1486 gnd 0.008714f
C3590 vdd.n1487 gnd 0.010826f
C3591 vdd.n1488 gnd 0.8685f
C3592 vdd.n1489 gnd 0.010826f
C3593 vdd.n1490 gnd 0.008714f
C3594 vdd.n1491 gnd 0.010826f
C3595 vdd.n1492 gnd 0.008714f
C3596 vdd.n1493 gnd 0.010826f
C3597 vdd.n1494 gnd 0.680417f
C3598 vdd.t116 gnd 0.553185f
C3599 vdd.n1495 gnd 0.010826f
C3600 vdd.n1496 gnd 0.008714f
C3601 vdd.n1497 gnd 0.010826f
C3602 vdd.n1498 gnd 0.008714f
C3603 vdd.n1499 gnd 0.010826f
C3604 vdd.t31 gnd 0.553185f
C3605 vdd.n1500 gnd 0.010826f
C3606 vdd.n1501 gnd 0.008714f
C3607 vdd.n1502 gnd 0.010826f
C3608 vdd.n1503 gnd 0.008714f
C3609 vdd.n1504 gnd 0.010826f
C3610 vdd.t56 gnd 0.553185f
C3611 vdd.n1505 gnd 0.614035f
C3612 vdd.n1506 gnd 0.010826f
C3613 vdd.n1507 gnd 0.008714f
C3614 vdd.n1508 gnd 0.010826f
C3615 vdd.n1509 gnd 0.008714f
C3616 vdd.n1510 gnd 0.010826f
C3617 vdd.t58 gnd 0.553185f
C3618 vdd.n1511 gnd 0.010826f
C3619 vdd.n1512 gnd 0.008714f
C3620 vdd.n1513 gnd 0.010826f
C3621 vdd.n1514 gnd 0.008714f
C3622 vdd.n1515 gnd 0.010826f
C3623 vdd.n1516 gnd 0.846373f
C3624 vdd.n1517 gnd 0.918287f
C3625 vdd.t23 gnd 0.553185f
C3626 vdd.n1518 gnd 0.010826f
C3627 vdd.n1519 gnd 0.008714f
C3628 vdd.n1520 gnd 0.010826f
C3629 vdd.n1521 gnd 0.008714f
C3630 vdd.n1522 gnd 0.010826f
C3631 vdd.n1523 gnd 0.65829f
C3632 vdd.n1524 gnd 0.010826f
C3633 vdd.n1525 gnd 0.008714f
C3634 vdd.n1526 gnd 0.010826f
C3635 vdd.n1527 gnd 0.008714f
C3636 vdd.n1528 gnd 0.010826f
C3637 vdd.t111 gnd 0.553185f
C3638 vdd.t87 gnd 0.553185f
C3639 vdd.n1529 gnd 0.010826f
C3640 vdd.n1530 gnd 0.008714f
C3641 vdd.n1531 gnd 0.010826f
C3642 vdd.n1532 gnd 0.008714f
C3643 vdd.n1533 gnd 0.010826f
C3644 vdd.t17 gnd 0.553185f
C3645 vdd.n1534 gnd 0.010826f
C3646 vdd.n1535 gnd 0.008714f
C3647 vdd.n1536 gnd 0.010826f
C3648 vdd.n1537 gnd 0.008714f
C3649 vdd.n1538 gnd 0.010826f
C3650 vdd.t73 gnd 0.553185f
C3651 vdd.n1539 gnd 0.824245f
C3652 vdd.n1540 gnd 0.010826f
C3653 vdd.n1541 gnd 0.008714f
C3654 vdd.n1542 gnd 0.010826f
C3655 vdd.n1543 gnd 0.008714f
C3656 vdd.n1544 gnd 0.010826f
C3657 vdd.n1545 gnd 1.10637f
C3658 vdd.n1546 gnd 0.010826f
C3659 vdd.n1547 gnd 0.008714f
C3660 vdd.n1548 gnd 0.026189f
C3661 vdd.n1549 gnd 0.007232f
C3662 vdd.n1550 gnd 0.026189f
C3663 vdd.t254 gnd 0.553185f
C3664 vdd.n1551 gnd 0.026189f
C3665 vdd.n1552 gnd 0.007232f
C3666 vdd.n1553 gnd 0.010826f
C3667 vdd.n1554 gnd 0.008714f
C3668 vdd.n1555 gnd 0.010826f
C3669 vdd.n1586 gnd 0.02675f
C3670 vdd.n1587 gnd 1.6319f
C3671 vdd.n1588 gnd 0.010826f
C3672 vdd.n1589 gnd 0.008714f
C3673 vdd.n1590 gnd 0.010826f
C3674 vdd.n1591 gnd 0.010826f
C3675 vdd.n1592 gnd 0.010826f
C3676 vdd.n1593 gnd 0.010826f
C3677 vdd.n1594 gnd 0.010826f
C3678 vdd.n1595 gnd 0.008714f
C3679 vdd.n1596 gnd 0.010826f
C3680 vdd.n1597 gnd 0.010826f
C3681 vdd.n1598 gnd 0.010826f
C3682 vdd.n1599 gnd 0.010826f
C3683 vdd.n1600 gnd 0.010826f
C3684 vdd.n1601 gnd 0.008714f
C3685 vdd.n1602 gnd 0.010826f
C3686 vdd.n1603 gnd 0.010826f
C3687 vdd.n1604 gnd 0.010826f
C3688 vdd.n1605 gnd 0.010826f
C3689 vdd.n1606 gnd 0.010826f
C3690 vdd.n1607 gnd 0.008714f
C3691 vdd.n1608 gnd 0.010826f
C3692 vdd.n1609 gnd 0.010826f
C3693 vdd.n1610 gnd 0.010826f
C3694 vdd.n1611 gnd 0.010826f
C3695 vdd.n1612 gnd 0.010826f
C3696 vdd.t285 gnd 0.133189f
C3697 vdd.t286 gnd 0.142342f
C3698 vdd.t284 gnd 0.173943f
C3699 vdd.n1613 gnd 0.22297f
C3700 vdd.n1614 gnd 0.188206f
C3701 vdd.n1615 gnd 0.018647f
C3702 vdd.n1616 gnd 0.010826f
C3703 vdd.n1617 gnd 0.010826f
C3704 vdd.n1618 gnd 0.010826f
C3705 vdd.n1619 gnd 0.010826f
C3706 vdd.n1620 gnd 0.010826f
C3707 vdd.n1621 gnd 0.008714f
C3708 vdd.n1622 gnd 0.010826f
C3709 vdd.n1623 gnd 0.010826f
C3710 vdd.n1624 gnd 0.010826f
C3711 vdd.n1625 gnd 0.010826f
C3712 vdd.n1626 gnd 0.010826f
C3713 vdd.n1627 gnd 0.008714f
C3714 vdd.n1628 gnd 0.010826f
C3715 vdd.n1629 gnd 0.010826f
C3716 vdd.n1630 gnd 0.010826f
C3717 vdd.n1631 gnd 0.010826f
C3718 vdd.n1632 gnd 0.010826f
C3719 vdd.n1633 gnd 0.008714f
C3720 vdd.n1634 gnd 0.010826f
C3721 vdd.n1635 gnd 0.010826f
C3722 vdd.n1636 gnd 0.010826f
C3723 vdd.n1637 gnd 0.010826f
C3724 vdd.n1638 gnd 0.010826f
C3725 vdd.n1639 gnd 0.008714f
C3726 vdd.n1640 gnd 0.010826f
C3727 vdd.n1641 gnd 0.010826f
C3728 vdd.n1642 gnd 0.010826f
C3729 vdd.n1643 gnd 0.010826f
C3730 vdd.n1644 gnd 0.010826f
C3731 vdd.n1645 gnd 0.008714f
C3732 vdd.n1646 gnd 0.010826f
C3733 vdd.n1647 gnd 0.010826f
C3734 vdd.n1648 gnd 0.010826f
C3735 vdd.n1649 gnd 0.010826f
C3736 vdd.n1650 gnd 0.008714f
C3737 vdd.n1651 gnd 0.010826f
C3738 vdd.n1652 gnd 0.010826f
C3739 vdd.n1653 gnd 0.010826f
C3740 vdd.n1654 gnd 0.010826f
C3741 vdd.n1655 gnd 0.010826f
C3742 vdd.n1656 gnd 0.008714f
C3743 vdd.n1657 gnd 0.010826f
C3744 vdd.n1658 gnd 0.010826f
C3745 vdd.n1659 gnd 0.010826f
C3746 vdd.n1660 gnd 0.010826f
C3747 vdd.n1661 gnd 0.010826f
C3748 vdd.n1662 gnd 0.008714f
C3749 vdd.n1663 gnd 0.010826f
C3750 vdd.n1664 gnd 0.010826f
C3751 vdd.n1665 gnd 0.010826f
C3752 vdd.n1666 gnd 0.010826f
C3753 vdd.n1667 gnd 0.010826f
C3754 vdd.n1668 gnd 0.008714f
C3755 vdd.n1669 gnd 0.010826f
C3756 vdd.n1670 gnd 0.010826f
C3757 vdd.n1671 gnd 0.010826f
C3758 vdd.n1672 gnd 0.010826f
C3759 vdd.n1673 gnd 0.010826f
C3760 vdd.n1674 gnd 0.008714f
C3761 vdd.n1675 gnd 0.010826f
C3762 vdd.n1676 gnd 0.010826f
C3763 vdd.n1677 gnd 0.010826f
C3764 vdd.n1678 gnd 0.010826f
C3765 vdd.t255 gnd 0.133189f
C3766 vdd.t256 gnd 0.142342f
C3767 vdd.t253 gnd 0.173943f
C3768 vdd.n1679 gnd 0.22297f
C3769 vdd.n1680 gnd 0.188206f
C3770 vdd.n1681 gnd 0.01429f
C3771 vdd.n1682 gnd 0.004139f
C3772 vdd.n1683 gnd 0.02675f
C3773 vdd.n1684 gnd 0.010826f
C3774 vdd.n1685 gnd 0.004575f
C3775 vdd.n1686 gnd 0.008714f
C3776 vdd.n1687 gnd 0.008714f
C3777 vdd.n1688 gnd 0.010826f
C3778 vdd.n1689 gnd 0.010826f
C3779 vdd.n1690 gnd 0.010826f
C3780 vdd.n1691 gnd 0.008714f
C3781 vdd.n1692 gnd 0.008714f
C3782 vdd.n1693 gnd 0.008714f
C3783 vdd.n1694 gnd 0.010826f
C3784 vdd.n1695 gnd 0.010826f
C3785 vdd.n1696 gnd 0.010826f
C3786 vdd.n1697 gnd 0.008714f
C3787 vdd.n1698 gnd 0.008714f
C3788 vdd.n1699 gnd 0.008714f
C3789 vdd.n1700 gnd 0.010826f
C3790 vdd.n1701 gnd 0.010826f
C3791 vdd.n1702 gnd 0.010826f
C3792 vdd.n1703 gnd 0.008714f
C3793 vdd.n1704 gnd 0.008714f
C3794 vdd.n1705 gnd 0.008714f
C3795 vdd.n1706 gnd 0.010826f
C3796 vdd.n1707 gnd 0.010826f
C3797 vdd.n1708 gnd 0.010826f
C3798 vdd.n1709 gnd 0.008714f
C3799 vdd.n1710 gnd 0.008714f
C3800 vdd.n1711 gnd 0.008714f
C3801 vdd.n1712 gnd 0.010826f
C3802 vdd.n1713 gnd 0.010826f
C3803 vdd.n1714 gnd 0.010826f
C3804 vdd.n1715 gnd 0.008627f
C3805 vdd.n1716 gnd 0.010826f
C3806 vdd.t272 gnd 0.133189f
C3807 vdd.t273 gnd 0.142342f
C3808 vdd.t271 gnd 0.173943f
C3809 vdd.n1717 gnd 0.22297f
C3810 vdd.n1718 gnd 0.188206f
C3811 vdd.n1719 gnd 0.018647f
C3812 vdd.n1720 gnd 0.005925f
C3813 vdd.n1721 gnd 0.010826f
C3814 vdd.n1722 gnd 0.010826f
C3815 vdd.n1723 gnd 0.010826f
C3816 vdd.n1724 gnd 0.008714f
C3817 vdd.n1725 gnd 0.008714f
C3818 vdd.n1726 gnd 0.008714f
C3819 vdd.n1727 gnd 0.010826f
C3820 vdd.n1728 gnd 0.010826f
C3821 vdd.n1729 gnd 0.010826f
C3822 vdd.n1730 gnd 0.008714f
C3823 vdd.n1731 gnd 0.008714f
C3824 vdd.n1732 gnd 0.008714f
C3825 vdd.n1733 gnd 0.010826f
C3826 vdd.n1734 gnd 0.010826f
C3827 vdd.n1735 gnd 0.010826f
C3828 vdd.n1736 gnd 0.008714f
C3829 vdd.n1737 gnd 0.008714f
C3830 vdd.n1738 gnd 0.008714f
C3831 vdd.n1739 gnd 0.010826f
C3832 vdd.n1740 gnd 0.010826f
C3833 vdd.n1741 gnd 0.010826f
C3834 vdd.n1742 gnd 0.008714f
C3835 vdd.n1743 gnd 0.008714f
C3836 vdd.n1744 gnd 0.008714f
C3837 vdd.n1745 gnd 0.010826f
C3838 vdd.n1746 gnd 0.010826f
C3839 vdd.n1747 gnd 0.010826f
C3840 vdd.n1748 gnd 0.008714f
C3841 vdd.n1749 gnd 0.008714f
C3842 vdd.n1750 gnd 0.007276f
C3843 vdd.n1751 gnd 0.010826f
C3844 vdd.n1752 gnd 0.010826f
C3845 vdd.n1753 gnd 0.010826f
C3846 vdd.n1754 gnd 0.007276f
C3847 vdd.n1755 gnd 0.008714f
C3848 vdd.n1756 gnd 0.008714f
C3849 vdd.n1757 gnd 0.010826f
C3850 vdd.n1758 gnd 0.010826f
C3851 vdd.n1759 gnd 0.010826f
C3852 vdd.n1760 gnd 0.008714f
C3853 vdd.n1761 gnd 0.008714f
C3854 vdd.n1762 gnd 0.008714f
C3855 vdd.n1763 gnd 0.010826f
C3856 vdd.n1764 gnd 0.010826f
C3857 vdd.n1765 gnd 0.010826f
C3858 vdd.n1766 gnd 0.008714f
C3859 vdd.n1767 gnd 0.008714f
C3860 vdd.n1768 gnd 0.008714f
C3861 vdd.n1769 gnd 0.010826f
C3862 vdd.n1770 gnd 0.010826f
C3863 vdd.n1771 gnd 0.010826f
C3864 vdd.n1772 gnd 0.008714f
C3865 vdd.n1773 gnd 0.008714f
C3866 vdd.n1774 gnd 0.008714f
C3867 vdd.n1775 gnd 0.010826f
C3868 vdd.n1776 gnd 0.010826f
C3869 vdd.n1777 gnd 0.010826f
C3870 vdd.n1778 gnd 0.008714f
C3871 vdd.n1779 gnd 0.010826f
C3872 vdd.n1780 gnd 2.6221f
C3873 vdd.n1782 gnd 0.02675f
C3874 vdd.n1783 gnd 0.007232f
C3875 vdd.n1784 gnd 0.02675f
C3876 vdd.n1785 gnd 0.026189f
C3877 vdd.n1786 gnd 0.010826f
C3878 vdd.n1787 gnd 0.008714f
C3879 vdd.n1788 gnd 0.010826f
C3880 vdd.n1789 gnd 0.558717f
C3881 vdd.n1790 gnd 0.010826f
C3882 vdd.n1791 gnd 0.008714f
C3883 vdd.n1792 gnd 0.010826f
C3884 vdd.n1793 gnd 0.010826f
C3885 vdd.n1794 gnd 0.010826f
C3886 vdd.n1795 gnd 0.008714f
C3887 vdd.n1796 gnd 0.010826f
C3888 vdd.n1797 gnd 1.01233f
C3889 vdd.n1798 gnd 1.10637f
C3890 vdd.n1799 gnd 0.010826f
C3891 vdd.n1800 gnd 0.008714f
C3892 vdd.n1801 gnd 0.010826f
C3893 vdd.n1802 gnd 0.010826f
C3894 vdd.n1803 gnd 0.010826f
C3895 vdd.n1804 gnd 0.008714f
C3896 vdd.n1805 gnd 0.010826f
C3897 vdd.n1806 gnd 0.647226f
C3898 vdd.n1807 gnd 0.010826f
C3899 vdd.n1808 gnd 0.008714f
C3900 vdd.n1809 gnd 0.010826f
C3901 vdd.n1810 gnd 0.010826f
C3902 vdd.n1811 gnd 0.010826f
C3903 vdd.n1812 gnd 0.008714f
C3904 vdd.n1813 gnd 0.010826f
C3905 vdd.n1814 gnd 0.636162f
C3906 vdd.n1815 gnd 0.835309f
C3907 vdd.n1816 gnd 0.010826f
C3908 vdd.n1817 gnd 0.008714f
C3909 vdd.n1818 gnd 0.010826f
C3910 vdd.n1819 gnd 0.010826f
C3911 vdd.n1820 gnd 0.010826f
C3912 vdd.n1821 gnd 0.008714f
C3913 vdd.n1822 gnd 0.010826f
C3914 vdd.n1823 gnd 0.918287f
C3915 vdd.n1824 gnd 0.010826f
C3916 vdd.n1825 gnd 0.008714f
C3917 vdd.n1826 gnd 0.010826f
C3918 vdd.n1827 gnd 0.010826f
C3919 vdd.n1828 gnd 0.010826f
C3920 vdd.n1829 gnd 0.008714f
C3921 vdd.n1830 gnd 0.010826f
C3922 vdd.t27 gnd 0.553185f
C3923 vdd.n1831 gnd 0.813182f
C3924 vdd.n1832 gnd 0.010826f
C3925 vdd.n1833 gnd 0.008714f
C3926 vdd.n1834 gnd 0.010826f
C3927 vdd.n1835 gnd 0.010826f
C3928 vdd.n1836 gnd 0.010826f
C3929 vdd.n1837 gnd 0.008714f
C3930 vdd.n1838 gnd 0.010826f
C3931 vdd.n1839 gnd 0.625099f
C3932 vdd.n1840 gnd 0.010826f
C3933 vdd.n1841 gnd 0.008714f
C3934 vdd.n1842 gnd 0.010826f
C3935 vdd.n1843 gnd 0.010826f
C3936 vdd.n1844 gnd 0.010826f
C3937 vdd.n1845 gnd 0.008714f
C3938 vdd.n1846 gnd 0.010826f
C3939 vdd.n1847 gnd 0.802118f
C3940 vdd.n1848 gnd 0.669354f
C3941 vdd.n1849 gnd 0.010826f
C3942 vdd.n1850 gnd 0.008714f
C3943 vdd.n1851 gnd 0.010826f
C3944 vdd.n1852 gnd 0.010826f
C3945 vdd.n1853 gnd 0.010826f
C3946 vdd.n1854 gnd 0.008714f
C3947 vdd.n1855 gnd 0.010826f
C3948 vdd.n1856 gnd 0.857436f
C3949 vdd.n1857 gnd 0.010826f
C3950 vdd.n1858 gnd 0.008714f
C3951 vdd.n1859 gnd 0.010826f
C3952 vdd.n1860 gnd 0.010826f
C3953 vdd.n1861 gnd 0.010826f
C3954 vdd.n1862 gnd 0.008714f
C3955 vdd.n1863 gnd 0.010826f
C3956 vdd.t118 gnd 0.553185f
C3957 vdd.n1864 gnd 0.918287f
C3958 vdd.n1865 gnd 0.010826f
C3959 vdd.n1866 gnd 0.008714f
C3960 vdd.n1867 gnd 0.010826f
C3961 vdd.n1868 gnd 0.00832f
C3962 vdd.n1869 gnd 0.005941f
C3963 vdd.n1870 gnd 0.005513f
C3964 vdd.n1871 gnd 0.00305f
C3965 vdd.n1872 gnd 0.007003f
C3966 vdd.n1873 gnd 0.002963f
C3967 vdd.n1874 gnd 0.003137f
C3968 vdd.n1875 gnd 0.005513f
C3969 vdd.n1876 gnd 0.002963f
C3970 vdd.n1877 gnd 0.007003f
C3971 vdd.n1878 gnd 0.003137f
C3972 vdd.n1879 gnd 0.005513f
C3973 vdd.n1880 gnd 0.002963f
C3974 vdd.n1881 gnd 0.005252f
C3975 vdd.n1882 gnd 0.005268f
C3976 vdd.t66 gnd 0.015044f
C3977 vdd.n1883 gnd 0.033474f
C3978 vdd.n1884 gnd 0.174205f
C3979 vdd.n1885 gnd 0.002963f
C3980 vdd.n1886 gnd 0.003137f
C3981 vdd.n1887 gnd 0.007003f
C3982 vdd.n1888 gnd 0.007003f
C3983 vdd.n1889 gnd 0.003137f
C3984 vdd.n1890 gnd 0.002963f
C3985 vdd.n1891 gnd 0.005513f
C3986 vdd.n1892 gnd 0.005513f
C3987 vdd.n1893 gnd 0.002963f
C3988 vdd.n1894 gnd 0.003137f
C3989 vdd.n1895 gnd 0.007003f
C3990 vdd.n1896 gnd 0.007003f
C3991 vdd.n1897 gnd 0.003137f
C3992 vdd.n1898 gnd 0.002963f
C3993 vdd.n1899 gnd 0.005513f
C3994 vdd.n1900 gnd 0.005513f
C3995 vdd.n1901 gnd 0.002963f
C3996 vdd.n1902 gnd 0.003137f
C3997 vdd.n1903 gnd 0.007003f
C3998 vdd.n1904 gnd 0.007003f
C3999 vdd.n1905 gnd 0.016556f
C4000 vdd.n1906 gnd 0.00305f
C4001 vdd.n1907 gnd 0.002963f
C4002 vdd.n1908 gnd 0.01425f
C4003 vdd.n1909 gnd 0.009949f
C4004 vdd.t98 gnd 0.034855f
C4005 vdd.t155 gnd 0.034855f
C4006 vdd.n1910 gnd 0.239545f
C4007 vdd.n1911 gnd 0.188365f
C4008 vdd.t122 gnd 0.034855f
C4009 vdd.t170 gnd 0.034855f
C4010 vdd.n1912 gnd 0.239545f
C4011 vdd.n1913 gnd 0.15201f
C4012 vdd.t86 gnd 0.034855f
C4013 vdd.t34 gnd 0.034855f
C4014 vdd.n1914 gnd 0.239545f
C4015 vdd.n1915 gnd 0.15201f
C4016 vdd.t113 gnd 0.034855f
C4017 vdd.t45 gnd 0.034855f
C4018 vdd.n1916 gnd 0.239545f
C4019 vdd.n1917 gnd 0.15201f
C4020 vdd.t159 gnd 0.034855f
C4021 vdd.t175 gnd 0.034855f
C4022 vdd.n1918 gnd 0.239545f
C4023 vdd.n1919 gnd 0.15201f
C4024 vdd.t132 gnd 0.034855f
C4025 vdd.t50 gnd 0.034855f
C4026 vdd.n1920 gnd 0.239545f
C4027 vdd.n1921 gnd 0.15201f
C4028 vdd.t123 gnd 0.034855f
C4029 vdd.t59 gnd 0.034855f
C4030 vdd.n1922 gnd 0.239545f
C4031 vdd.n1923 gnd 0.15201f
C4032 vdd.t164 gnd 0.034855f
C4033 vdd.t92 gnd 0.034855f
C4034 vdd.n1924 gnd 0.239545f
C4035 vdd.n1925 gnd 0.15201f
C4036 vdd.t142 gnd 0.034855f
C4037 vdd.t112 gnd 0.034855f
C4038 vdd.n1926 gnd 0.239545f
C4039 vdd.n1927 gnd 0.15201f
C4040 vdd.n1928 gnd 0.005941f
C4041 vdd.n1929 gnd 0.005513f
C4042 vdd.n1930 gnd 0.00305f
C4043 vdd.n1931 gnd 0.007003f
C4044 vdd.n1932 gnd 0.002963f
C4045 vdd.n1933 gnd 0.003137f
C4046 vdd.n1934 gnd 0.005513f
C4047 vdd.n1935 gnd 0.002963f
C4048 vdd.n1936 gnd 0.007003f
C4049 vdd.n1937 gnd 0.003137f
C4050 vdd.n1938 gnd 0.005513f
C4051 vdd.n1939 gnd 0.002963f
C4052 vdd.n1940 gnd 0.005252f
C4053 vdd.n1941 gnd 0.005268f
C4054 vdd.t74 gnd 0.015044f
C4055 vdd.n1942 gnd 0.033474f
C4056 vdd.n1943 gnd 0.174205f
C4057 vdd.n1944 gnd 0.002963f
C4058 vdd.n1945 gnd 0.003137f
C4059 vdd.n1946 gnd 0.007003f
C4060 vdd.n1947 gnd 0.007003f
C4061 vdd.n1948 gnd 0.003137f
C4062 vdd.n1949 gnd 0.002963f
C4063 vdd.n1950 gnd 0.005513f
C4064 vdd.n1951 gnd 0.005513f
C4065 vdd.n1952 gnd 0.002963f
C4066 vdd.n1953 gnd 0.003137f
C4067 vdd.n1954 gnd 0.007003f
C4068 vdd.n1955 gnd 0.007003f
C4069 vdd.n1956 gnd 0.003137f
C4070 vdd.n1957 gnd 0.002963f
C4071 vdd.n1958 gnd 0.005513f
C4072 vdd.n1959 gnd 0.005513f
C4073 vdd.n1960 gnd 0.002963f
C4074 vdd.n1961 gnd 0.003137f
C4075 vdd.n1962 gnd 0.007003f
C4076 vdd.n1963 gnd 0.007003f
C4077 vdd.n1964 gnd 0.016556f
C4078 vdd.n1965 gnd 0.00305f
C4079 vdd.n1966 gnd 0.002963f
C4080 vdd.n1967 gnd 0.01425f
C4081 vdd.n1968 gnd 0.009637f
C4082 vdd.n1969 gnd 0.113096f
C4083 vdd.n1970 gnd 0.005941f
C4084 vdd.n1971 gnd 0.005513f
C4085 vdd.n1972 gnd 0.00305f
C4086 vdd.n1973 gnd 0.007003f
C4087 vdd.n1974 gnd 0.002963f
C4088 vdd.n1975 gnd 0.003137f
C4089 vdd.n1976 gnd 0.005513f
C4090 vdd.n1977 gnd 0.002963f
C4091 vdd.n1978 gnd 0.007003f
C4092 vdd.n1979 gnd 0.003137f
C4093 vdd.n1980 gnd 0.005513f
C4094 vdd.n1981 gnd 0.002963f
C4095 vdd.n1982 gnd 0.005252f
C4096 vdd.n1983 gnd 0.005268f
C4097 vdd.t153 gnd 0.015044f
C4098 vdd.n1984 gnd 0.033474f
C4099 vdd.n1985 gnd 0.174205f
C4100 vdd.n1986 gnd 0.002963f
C4101 vdd.n1987 gnd 0.003137f
C4102 vdd.n1988 gnd 0.007003f
C4103 vdd.n1989 gnd 0.007003f
C4104 vdd.n1990 gnd 0.003137f
C4105 vdd.n1991 gnd 0.002963f
C4106 vdd.n1992 gnd 0.005513f
C4107 vdd.n1993 gnd 0.005513f
C4108 vdd.n1994 gnd 0.002963f
C4109 vdd.n1995 gnd 0.003137f
C4110 vdd.n1996 gnd 0.007003f
C4111 vdd.n1997 gnd 0.007003f
C4112 vdd.n1998 gnd 0.003137f
C4113 vdd.n1999 gnd 0.002963f
C4114 vdd.n2000 gnd 0.005513f
C4115 vdd.n2001 gnd 0.005513f
C4116 vdd.n2002 gnd 0.002963f
C4117 vdd.n2003 gnd 0.003137f
C4118 vdd.n2004 gnd 0.007003f
C4119 vdd.n2005 gnd 0.007003f
C4120 vdd.n2006 gnd 0.016556f
C4121 vdd.n2007 gnd 0.00305f
C4122 vdd.n2008 gnd 0.002963f
C4123 vdd.n2009 gnd 0.01425f
C4124 vdd.n2010 gnd 0.009949f
C4125 vdd.t102 gnd 0.034855f
C4126 vdd.t26 gnd 0.034855f
C4127 vdd.n2011 gnd 0.239545f
C4128 vdd.n2012 gnd 0.188365f
C4129 vdd.t166 gnd 0.034855f
C4130 vdd.t134 gnd 0.034855f
C4131 vdd.n2013 gnd 0.239545f
C4132 vdd.n2014 gnd 0.15201f
C4133 vdd.t129 gnd 0.034855f
C4134 vdd.t67 gnd 0.034855f
C4135 vdd.n2015 gnd 0.239545f
C4136 vdd.n2016 gnd 0.15201f
C4137 vdd.t61 gnd 0.034855f
C4138 vdd.t110 gnd 0.034855f
C4139 vdd.n2017 gnd 0.239545f
C4140 vdd.n2018 gnd 0.15201f
C4141 vdd.t119 gnd 0.034855f
C4142 vdd.t117 gnd 0.034855f
C4143 vdd.n2019 gnd 0.239545f
C4144 vdd.n2020 gnd 0.15201f
C4145 vdd.t57 gnd 0.034855f
C4146 vdd.t32 gnd 0.034855f
C4147 vdd.n2021 gnd 0.239545f
C4148 vdd.n2022 gnd 0.15201f
C4149 vdd.t24 gnd 0.034855f
C4150 vdd.t114 gnd 0.034855f
C4151 vdd.n2023 gnd 0.239545f
C4152 vdd.n2024 gnd 0.15201f
C4153 vdd.t88 gnd 0.034855f
C4154 vdd.t28 gnd 0.034855f
C4155 vdd.n2025 gnd 0.239545f
C4156 vdd.n2026 gnd 0.15201f
C4157 vdd.t18 gnd 0.034855f
C4158 vdd.t135 gnd 0.034855f
C4159 vdd.n2027 gnd 0.239545f
C4160 vdd.n2028 gnd 0.15201f
C4161 vdd.n2029 gnd 0.005941f
C4162 vdd.n2030 gnd 0.005513f
C4163 vdd.n2031 gnd 0.00305f
C4164 vdd.n2032 gnd 0.007003f
C4165 vdd.n2033 gnd 0.002963f
C4166 vdd.n2034 gnd 0.003137f
C4167 vdd.n2035 gnd 0.005513f
C4168 vdd.n2036 gnd 0.002963f
C4169 vdd.n2037 gnd 0.007003f
C4170 vdd.n2038 gnd 0.003137f
C4171 vdd.n2039 gnd 0.005513f
C4172 vdd.n2040 gnd 0.002963f
C4173 vdd.n2041 gnd 0.005252f
C4174 vdd.n2042 gnd 0.005268f
C4175 vdd.t76 gnd 0.015044f
C4176 vdd.n2043 gnd 0.033474f
C4177 vdd.n2044 gnd 0.174205f
C4178 vdd.n2045 gnd 0.002963f
C4179 vdd.n2046 gnd 0.003137f
C4180 vdd.n2047 gnd 0.007003f
C4181 vdd.n2048 gnd 0.007003f
C4182 vdd.n2049 gnd 0.003137f
C4183 vdd.n2050 gnd 0.002963f
C4184 vdd.n2051 gnd 0.005513f
C4185 vdd.n2052 gnd 0.005513f
C4186 vdd.n2053 gnd 0.002963f
C4187 vdd.n2054 gnd 0.003137f
C4188 vdd.n2055 gnd 0.007003f
C4189 vdd.n2056 gnd 0.007003f
C4190 vdd.n2057 gnd 0.003137f
C4191 vdd.n2058 gnd 0.002963f
C4192 vdd.n2059 gnd 0.005513f
C4193 vdd.n2060 gnd 0.005513f
C4194 vdd.n2061 gnd 0.002963f
C4195 vdd.n2062 gnd 0.003137f
C4196 vdd.n2063 gnd 0.007003f
C4197 vdd.n2064 gnd 0.007003f
C4198 vdd.n2065 gnd 0.016556f
C4199 vdd.n2066 gnd 0.00305f
C4200 vdd.n2067 gnd 0.002963f
C4201 vdd.n2068 gnd 0.01425f
C4202 vdd.n2069 gnd 0.009637f
C4203 vdd.n2070 gnd 0.067281f
C4204 vdd.n2071 gnd 0.24243f
C4205 vdd.n2072 gnd 0.005941f
C4206 vdd.n2073 gnd 0.005513f
C4207 vdd.n2074 gnd 0.00305f
C4208 vdd.n2075 gnd 0.007003f
C4209 vdd.n2076 gnd 0.002963f
C4210 vdd.n2077 gnd 0.003137f
C4211 vdd.n2078 gnd 0.005513f
C4212 vdd.n2079 gnd 0.002963f
C4213 vdd.n2080 gnd 0.007003f
C4214 vdd.n2081 gnd 0.003137f
C4215 vdd.n2082 gnd 0.005513f
C4216 vdd.n2083 gnd 0.002963f
C4217 vdd.n2084 gnd 0.005252f
C4218 vdd.n2085 gnd 0.005268f
C4219 vdd.t165 gnd 0.015044f
C4220 vdd.n2086 gnd 0.033474f
C4221 vdd.n2087 gnd 0.174205f
C4222 vdd.n2088 gnd 0.002963f
C4223 vdd.n2089 gnd 0.003137f
C4224 vdd.n2090 gnd 0.007003f
C4225 vdd.n2091 gnd 0.007003f
C4226 vdd.n2092 gnd 0.003137f
C4227 vdd.n2093 gnd 0.002963f
C4228 vdd.n2094 gnd 0.005513f
C4229 vdd.n2095 gnd 0.005513f
C4230 vdd.n2096 gnd 0.002963f
C4231 vdd.n2097 gnd 0.003137f
C4232 vdd.n2098 gnd 0.007003f
C4233 vdd.n2099 gnd 0.007003f
C4234 vdd.n2100 gnd 0.003137f
C4235 vdd.n2101 gnd 0.002963f
C4236 vdd.n2102 gnd 0.005513f
C4237 vdd.n2103 gnd 0.005513f
C4238 vdd.n2104 gnd 0.002963f
C4239 vdd.n2105 gnd 0.003137f
C4240 vdd.n2106 gnd 0.007003f
C4241 vdd.n2107 gnd 0.007003f
C4242 vdd.n2108 gnd 0.016556f
C4243 vdd.n2109 gnd 0.00305f
C4244 vdd.n2110 gnd 0.002963f
C4245 vdd.n2111 gnd 0.01425f
C4246 vdd.n2112 gnd 0.009949f
C4247 vdd.t120 gnd 0.034855f
C4248 vdd.t52 gnd 0.034855f
C4249 vdd.n2113 gnd 0.239545f
C4250 vdd.n2114 gnd 0.188365f
C4251 vdd.t176 gnd 0.034855f
C4252 vdd.t146 gnd 0.034855f
C4253 vdd.n2115 gnd 0.239545f
C4254 vdd.n2116 gnd 0.15201f
C4255 vdd.t144 gnd 0.034855f
C4256 vdd.t93 gnd 0.034855f
C4257 vdd.n2117 gnd 0.239545f
C4258 vdd.n2118 gnd 0.15201f
C4259 vdd.t89 gnd 0.034855f
C4260 vdd.t145 gnd 0.034855f
C4261 vdd.n2119 gnd 0.239545f
C4262 vdd.n2120 gnd 0.15201f
C4263 vdd.t128 gnd 0.034855f
C4264 vdd.t127 gnd 0.034855f
C4265 vdd.n2121 gnd 0.239545f
C4266 vdd.n2122 gnd 0.15201f
C4267 vdd.t84 gnd 0.034855f
C4268 vdd.t53 gnd 0.034855f
C4269 vdd.n2123 gnd 0.239545f
C4270 vdd.n2124 gnd 0.15201f
C4271 vdd.t51 gnd 0.034855f
C4272 vdd.t126 gnd 0.034855f
C4273 vdd.n2125 gnd 0.239545f
C4274 vdd.n2126 gnd 0.15201f
C4275 vdd.t104 gnd 0.034855f
C4276 vdd.t49 gnd 0.034855f
C4277 vdd.n2127 gnd 0.239545f
C4278 vdd.n2128 gnd 0.15201f
C4279 vdd.t43 gnd 0.034855f
C4280 vdd.t148 gnd 0.034855f
C4281 vdd.n2129 gnd 0.239545f
C4282 vdd.n2130 gnd 0.15201f
C4283 vdd.n2131 gnd 0.005941f
C4284 vdd.n2132 gnd 0.005513f
C4285 vdd.n2133 gnd 0.00305f
C4286 vdd.n2134 gnd 0.007003f
C4287 vdd.n2135 gnd 0.002963f
C4288 vdd.n2136 gnd 0.003137f
C4289 vdd.n2137 gnd 0.005513f
C4290 vdd.n2138 gnd 0.002963f
C4291 vdd.n2139 gnd 0.007003f
C4292 vdd.n2140 gnd 0.003137f
C4293 vdd.n2141 gnd 0.005513f
C4294 vdd.n2142 gnd 0.002963f
C4295 vdd.n2143 gnd 0.005252f
C4296 vdd.n2144 gnd 0.005268f
C4297 vdd.t99 gnd 0.015044f
C4298 vdd.n2145 gnd 0.033474f
C4299 vdd.n2146 gnd 0.174205f
C4300 vdd.n2147 gnd 0.002963f
C4301 vdd.n2148 gnd 0.003137f
C4302 vdd.n2149 gnd 0.007003f
C4303 vdd.n2150 gnd 0.007003f
C4304 vdd.n2151 gnd 0.003137f
C4305 vdd.n2152 gnd 0.002963f
C4306 vdd.n2153 gnd 0.005513f
C4307 vdd.n2154 gnd 0.005513f
C4308 vdd.n2155 gnd 0.002963f
C4309 vdd.n2156 gnd 0.003137f
C4310 vdd.n2157 gnd 0.007003f
C4311 vdd.n2158 gnd 0.007003f
C4312 vdd.n2159 gnd 0.003137f
C4313 vdd.n2160 gnd 0.002963f
C4314 vdd.n2161 gnd 0.005513f
C4315 vdd.n2162 gnd 0.005513f
C4316 vdd.n2163 gnd 0.002963f
C4317 vdd.n2164 gnd 0.003137f
C4318 vdd.n2165 gnd 0.007003f
C4319 vdd.n2166 gnd 0.007003f
C4320 vdd.n2167 gnd 0.016556f
C4321 vdd.n2168 gnd 0.00305f
C4322 vdd.n2169 gnd 0.002963f
C4323 vdd.n2170 gnd 0.01425f
C4324 vdd.n2171 gnd 0.009637f
C4325 vdd.n2172 gnd 0.067281f
C4326 vdd.n2173 gnd 0.27753f
C4327 vdd.n2174 gnd 2.91139f
C4328 vdd.n2175 gnd 0.638561f
C4329 vdd.n2176 gnd 0.00832f
C4330 vdd.n2177 gnd 0.008714f
C4331 vdd.n2178 gnd 0.010826f
C4332 vdd.n2179 gnd 0.791054f
C4333 vdd.n2180 gnd 0.010826f
C4334 vdd.n2181 gnd 0.008714f
C4335 vdd.n2182 gnd 0.010826f
C4336 vdd.n2183 gnd 0.010826f
C4337 vdd.n2184 gnd 0.010826f
C4338 vdd.n2185 gnd 0.008714f
C4339 vdd.n2186 gnd 0.010826f
C4340 vdd.n2187 gnd 0.918287f
C4341 vdd.t60 gnd 0.553185f
C4342 vdd.n2188 gnd 0.602971f
C4343 vdd.n2189 gnd 0.010826f
C4344 vdd.n2190 gnd 0.008714f
C4345 vdd.n2191 gnd 0.010826f
C4346 vdd.n2192 gnd 0.010826f
C4347 vdd.n2193 gnd 0.010826f
C4348 vdd.n2194 gnd 0.008714f
C4349 vdd.n2195 gnd 0.010826f
C4350 vdd.n2196 gnd 0.691481f
C4351 vdd.n2197 gnd 0.010826f
C4352 vdd.n2198 gnd 0.008714f
C4353 vdd.n2199 gnd 0.010826f
C4354 vdd.n2200 gnd 0.010826f
C4355 vdd.n2201 gnd 0.010826f
C4356 vdd.n2202 gnd 0.008714f
C4357 vdd.n2203 gnd 0.010826f
C4358 vdd.n2204 gnd 0.591908f
C4359 vdd.n2205 gnd 0.879564f
C4360 vdd.n2206 gnd 0.010826f
C4361 vdd.n2207 gnd 0.008714f
C4362 vdd.n2208 gnd 0.010826f
C4363 vdd.n2209 gnd 0.010826f
C4364 vdd.n2210 gnd 0.010826f
C4365 vdd.n2211 gnd 0.008714f
C4366 vdd.n2212 gnd 0.010826f
C4367 vdd.n2213 gnd 0.918287f
C4368 vdd.n2214 gnd 0.010826f
C4369 vdd.n2215 gnd 0.008714f
C4370 vdd.n2216 gnd 0.010826f
C4371 vdd.n2217 gnd 0.010826f
C4372 vdd.n2218 gnd 0.010826f
C4373 vdd.n2219 gnd 0.008714f
C4374 vdd.n2220 gnd 0.010826f
C4375 vdd.t133 gnd 0.553185f
C4376 vdd.n2221 gnd 0.768927f
C4377 vdd.n2222 gnd 0.010826f
C4378 vdd.n2223 gnd 0.008714f
C4379 vdd.n2224 gnd 0.010826f
C4380 vdd.n2225 gnd 0.010826f
C4381 vdd.n2226 gnd 0.010826f
C4382 vdd.n2227 gnd 0.008714f
C4383 vdd.n2228 gnd 0.010826f
C4384 vdd.n2229 gnd 0.580844f
C4385 vdd.n2230 gnd 0.010826f
C4386 vdd.n2231 gnd 0.008714f
C4387 vdd.n2232 gnd 0.010826f
C4388 vdd.n2233 gnd 0.010826f
C4389 vdd.n2234 gnd 0.010826f
C4390 vdd.n2235 gnd 0.008714f
C4391 vdd.n2236 gnd 0.010826f
C4392 vdd.n2237 gnd 0.757863f
C4393 vdd.n2238 gnd 0.713608f
C4394 vdd.n2239 gnd 0.010826f
C4395 vdd.n2240 gnd 0.008714f
C4396 vdd.n2241 gnd 0.010826f
C4397 vdd.n2242 gnd 0.010826f
C4398 vdd.n2243 gnd 0.010826f
C4399 vdd.n2244 gnd 0.008714f
C4400 vdd.n2245 gnd 0.010826f
C4401 vdd.n2246 gnd 0.901691f
C4402 vdd.n2247 gnd 0.010826f
C4403 vdd.n2248 gnd 0.008714f
C4404 vdd.n2249 gnd 0.010826f
C4405 vdd.n2250 gnd 0.010826f
C4406 vdd.n2251 gnd 0.026189f
C4407 vdd.n2252 gnd 0.010826f
C4408 vdd.n2253 gnd 0.010826f
C4409 vdd.n2254 gnd 0.008714f
C4410 vdd.n2255 gnd 0.010826f
C4411 vdd.n2256 gnd 0.669354f
C4412 vdd.n2257 gnd 1.10637f
C4413 vdd.n2258 gnd 0.010826f
C4414 vdd.n2259 gnd 0.008714f
C4415 vdd.n2260 gnd 0.010826f
C4416 vdd.n2261 gnd 0.010826f
C4417 vdd.n2262 gnd 0.026189f
C4418 vdd.n2263 gnd 0.007232f
C4419 vdd.n2264 gnd 0.026189f
C4420 vdd.n2265 gnd 1.52126f
C4421 vdd.n2266 gnd 0.026189f
C4422 vdd.n2267 gnd 0.02675f
C4423 vdd.n2268 gnd 0.004139f
C4424 vdd.t232 gnd 0.133189f
C4425 vdd.t231 gnd 0.142342f
C4426 vdd.t229 gnd 0.173943f
C4427 vdd.n2269 gnd 0.22297f
C4428 vdd.n2270 gnd 0.187335f
C4429 vdd.n2271 gnd 0.013419f
C4430 vdd.n2272 gnd 0.004575f
C4431 vdd.n2273 gnd 0.00931f
C4432 vdd.n2274 gnd 0.818724f
C4433 vdd.n2276 gnd 0.008714f
C4434 vdd.n2277 gnd 0.008714f
C4435 vdd.n2278 gnd 0.010826f
C4436 vdd.n2280 gnd 0.010826f
C4437 vdd.n2281 gnd 0.010826f
C4438 vdd.n2282 gnd 0.008714f
C4439 vdd.n2283 gnd 0.008714f
C4440 vdd.n2284 gnd 0.008714f
C4441 vdd.n2285 gnd 0.010826f
C4442 vdd.n2287 gnd 0.010826f
C4443 vdd.n2288 gnd 0.010826f
C4444 vdd.n2289 gnd 0.008714f
C4445 vdd.n2290 gnd 0.008714f
C4446 vdd.n2291 gnd 0.008714f
C4447 vdd.n2292 gnd 0.010826f
C4448 vdd.n2294 gnd 0.010826f
C4449 vdd.n2295 gnd 0.010826f
C4450 vdd.n2296 gnd 0.008714f
C4451 vdd.n2297 gnd 0.008714f
C4452 vdd.n2298 gnd 0.008714f
C4453 vdd.n2299 gnd 0.010826f
C4454 vdd.n2301 gnd 0.010826f
C4455 vdd.n2302 gnd 0.010826f
C4456 vdd.n2303 gnd 0.008714f
C4457 vdd.n2304 gnd 0.010826f
C4458 vdd.n2305 gnd 0.010826f
C4459 vdd.n2306 gnd 0.010826f
C4460 vdd.n2307 gnd 0.017776f
C4461 vdd.n2308 gnd 0.005925f
C4462 vdd.n2309 gnd 0.008714f
C4463 vdd.n2310 gnd 0.010826f
C4464 vdd.n2312 gnd 0.010826f
C4465 vdd.n2313 gnd 0.010826f
C4466 vdd.n2314 gnd 0.008714f
C4467 vdd.n2315 gnd 0.008714f
C4468 vdd.n2316 gnd 0.008714f
C4469 vdd.n2317 gnd 0.010826f
C4470 vdd.n2319 gnd 0.010826f
C4471 vdd.n2320 gnd 0.010826f
C4472 vdd.n2321 gnd 0.008714f
C4473 vdd.n2322 gnd 0.008714f
C4474 vdd.n2323 gnd 0.008714f
C4475 vdd.n2324 gnd 0.010826f
C4476 vdd.n2326 gnd 0.010826f
C4477 vdd.n2327 gnd 0.010826f
C4478 vdd.n2328 gnd 0.008714f
C4479 vdd.n2329 gnd 0.008714f
C4480 vdd.n2330 gnd 0.008714f
C4481 vdd.n2331 gnd 0.010826f
C4482 vdd.n2333 gnd 0.010826f
C4483 vdd.n2334 gnd 0.010826f
C4484 vdd.n2335 gnd 0.008714f
C4485 vdd.n2336 gnd 0.008714f
C4486 vdd.n2337 gnd 0.008714f
C4487 vdd.n2338 gnd 0.010826f
C4488 vdd.n2340 gnd 0.010826f
C4489 vdd.n2341 gnd 0.010826f
C4490 vdd.n2342 gnd 0.008714f
C4491 vdd.n2343 gnd 0.010826f
C4492 vdd.n2344 gnd 0.010826f
C4493 vdd.n2345 gnd 0.010826f
C4494 vdd.n2346 gnd 0.017776f
C4495 vdd.n2347 gnd 0.007276f
C4496 vdd.n2348 gnd 0.008714f
C4497 vdd.n2349 gnd 0.010826f
C4498 vdd.n2351 gnd 0.010826f
C4499 vdd.n2352 gnd 0.010826f
C4500 vdd.n2353 gnd 0.008714f
C4501 vdd.n2354 gnd 0.008714f
C4502 vdd.n2355 gnd 0.008714f
C4503 vdd.n2356 gnd 0.010826f
C4504 vdd.n2358 gnd 0.010826f
C4505 vdd.n2359 gnd 0.010826f
C4506 vdd.n2360 gnd 0.008714f
C4507 vdd.n2361 gnd 0.008714f
C4508 vdd.n2362 gnd 0.008714f
C4509 vdd.n2363 gnd 0.010826f
C4510 vdd.n2365 gnd 0.010826f
C4511 vdd.n2366 gnd 0.010826f
C4512 vdd.n2367 gnd 0.008714f
C4513 vdd.n2368 gnd 0.008714f
C4514 vdd.n2369 gnd 0.008714f
C4515 vdd.n2370 gnd 0.010826f
C4516 vdd.n2372 gnd 0.010826f
C4517 vdd.n2373 gnd 0.008714f
C4518 vdd.n2374 gnd 0.008714f
C4519 vdd.n2375 gnd 0.010826f
C4520 vdd.n2377 gnd 0.010826f
C4521 vdd.n2378 gnd 0.010826f
C4522 vdd.n2379 gnd 0.008714f
C4523 vdd.n2380 gnd 0.00931f
C4524 vdd.n2381 gnd 0.818724f
C4525 vdd.n2382 gnd 0.029505f
C4526 vdd.n2383 gnd 0.007362f
C4527 vdd.n2384 gnd 0.007362f
C4528 vdd.n2385 gnd 0.007362f
C4529 vdd.n2386 gnd 0.007362f
C4530 vdd.n2387 gnd 0.007362f
C4531 vdd.n2388 gnd 0.007362f
C4532 vdd.n2389 gnd 0.007362f
C4533 vdd.n2390 gnd 0.007362f
C4534 vdd.n2391 gnd 0.007362f
C4535 vdd.n2392 gnd 0.007362f
C4536 vdd.n2393 gnd 0.007362f
C4537 vdd.n2394 gnd 0.007362f
C4538 vdd.n2395 gnd 0.007362f
C4539 vdd.n2396 gnd 0.007362f
C4540 vdd.n2397 gnd 0.007362f
C4541 vdd.n2398 gnd 0.007362f
C4542 vdd.n2399 gnd 0.007362f
C4543 vdd.n2400 gnd 0.007362f
C4544 vdd.n2401 gnd 0.007362f
C4545 vdd.n2402 gnd 0.007362f
C4546 vdd.n2403 gnd 0.007362f
C4547 vdd.n2404 gnd 0.007362f
C4548 vdd.n2405 gnd 0.007362f
C4549 vdd.n2406 gnd 0.007362f
C4550 vdd.n2407 gnd 0.007362f
C4551 vdd.n2408 gnd 0.007362f
C4552 vdd.n2409 gnd 0.007362f
C4553 vdd.n2410 gnd 0.007362f
C4554 vdd.n2411 gnd 0.007362f
C4555 vdd.n2412 gnd 0.007362f
C4556 vdd.n2413 gnd 0.007362f
C4557 vdd.n2414 gnd 0.017219f
C4558 vdd.n2415 gnd 0.017219f
C4559 vdd.n2417 gnd 9.43733f
C4560 vdd.n2419 gnd 0.017219f
C4561 vdd.n2420 gnd 0.017219f
C4562 vdd.n2421 gnd 0.016126f
C4563 vdd.n2422 gnd 0.007362f
C4564 vdd.n2423 gnd 0.007362f
C4565 vdd.n2424 gnd 0.752331f
C4566 vdd.n2425 gnd 0.007362f
C4567 vdd.n2426 gnd 0.007362f
C4568 vdd.n2427 gnd 0.007362f
C4569 vdd.n2428 gnd 0.007362f
C4570 vdd.n2429 gnd 0.007362f
C4571 vdd.n2430 gnd 0.636162f
C4572 vdd.n2431 gnd 0.007362f
C4573 vdd.n2432 gnd 0.007362f
C4574 vdd.n2433 gnd 0.007362f
C4575 vdd.n2434 gnd 0.007362f
C4576 vdd.n2435 gnd 0.007362f
C4577 vdd.n2436 gnd 0.752331f
C4578 vdd.n2437 gnd 0.007362f
C4579 vdd.n2438 gnd 0.007362f
C4580 vdd.n2439 gnd 0.007362f
C4581 vdd.n2440 gnd 0.007362f
C4582 vdd.n2441 gnd 0.007362f
C4583 vdd.n2442 gnd 0.735736f
C4584 vdd.n2443 gnd 0.007362f
C4585 vdd.n2444 gnd 0.007362f
C4586 vdd.n2445 gnd 0.007362f
C4587 vdd.n2446 gnd 0.007362f
C4588 vdd.n2447 gnd 0.007362f
C4589 vdd.n2448 gnd 0.752331f
C4590 vdd.n2449 gnd 0.007362f
C4591 vdd.n2450 gnd 0.007362f
C4592 vdd.n2451 gnd 0.007362f
C4593 vdd.n2452 gnd 0.007362f
C4594 vdd.n2453 gnd 0.007362f
C4595 vdd.n2454 gnd 0.602971f
C4596 vdd.n2455 gnd 0.007362f
C4597 vdd.n2456 gnd 0.007362f
C4598 vdd.n2457 gnd 0.006279f
C4599 vdd.n2458 gnd 0.021326f
C4600 vdd.n2459 gnd 0.004763f
C4601 vdd.n2460 gnd 0.007362f
C4602 vdd.n2461 gnd 0.437016f
C4603 vdd.n2462 gnd 0.007362f
C4604 vdd.n2463 gnd 0.007362f
C4605 vdd.n2464 gnd 0.007362f
C4606 vdd.n2465 gnd 0.007362f
C4607 vdd.n2466 gnd 0.007362f
C4608 vdd.n2467 gnd 0.481271f
C4609 vdd.n2468 gnd 0.007362f
C4610 vdd.n2469 gnd 0.007362f
C4611 vdd.n2470 gnd 0.007362f
C4612 vdd.n2471 gnd 0.007362f
C4613 vdd.n2472 gnd 0.007362f
C4614 vdd.n2473 gnd 0.647226f
C4615 vdd.n2474 gnd 0.007362f
C4616 vdd.n2475 gnd 0.007362f
C4617 vdd.n2476 gnd 0.007362f
C4618 vdd.n2477 gnd 0.007362f
C4619 vdd.n2478 gnd 0.007362f
C4620 vdd.n2479 gnd 0.619567f
C4621 vdd.n2480 gnd 0.007362f
C4622 vdd.n2481 gnd 0.007362f
C4623 vdd.n2482 gnd 0.007362f
C4624 vdd.n2483 gnd 0.007362f
C4625 vdd.n2484 gnd 0.007362f
C4626 vdd.n2485 gnd 0.453611f
C4627 vdd.n2486 gnd 0.007362f
C4628 vdd.n2487 gnd 0.007362f
C4629 vdd.n2488 gnd 0.007362f
C4630 vdd.n2489 gnd 0.007362f
C4631 vdd.n2490 gnd 0.007362f
C4632 vdd.n2491 gnd 0.237869f
C4633 vdd.n2492 gnd 0.007362f
C4634 vdd.n2493 gnd 0.007362f
C4635 vdd.n2494 gnd 0.007362f
C4636 vdd.n2495 gnd 0.007362f
C4637 vdd.n2496 gnd 0.007362f
C4638 vdd.n2497 gnd 0.392761f
C4639 vdd.n2498 gnd 0.007362f
C4640 vdd.n2499 gnd 0.007362f
C4641 vdd.n2500 gnd 0.007362f
C4642 vdd.n2501 gnd 0.007362f
C4643 vdd.n2502 gnd 0.007362f
C4644 vdd.n2503 gnd 0.752331f
C4645 vdd.n2504 gnd 0.007362f
C4646 vdd.n2505 gnd 0.007362f
C4647 vdd.n2506 gnd 0.007362f
C4648 vdd.n2507 gnd 0.007362f
C4649 vdd.n2508 gnd 0.007362f
C4650 vdd.n2509 gnd 0.007362f
C4651 vdd.n2510 gnd 0.007362f
C4652 vdd.n2511 gnd 0.564248f
C4653 vdd.n2512 gnd 0.007362f
C4654 vdd.n2513 gnd 0.007362f
C4655 vdd.n2514 gnd 0.007362f
C4656 vdd.n2515 gnd 0.007362f
C4657 vdd.n2516 gnd 0.007362f
C4658 vdd.n2517 gnd 0.007362f
C4659 vdd.n2518 gnd 0.470207f
C4660 vdd.n2519 gnd 0.007362f
C4661 vdd.n2520 gnd 0.007362f
C4662 vdd.n2521 gnd 0.007362f
C4663 vdd.n2522 gnd 0.01704f
C4664 vdd.n2523 gnd 0.016304f
C4665 vdd.n2524 gnd 0.007362f
C4666 vdd.n2525 gnd 0.007362f
C4667 vdd.n2526 gnd 0.005684f
C4668 vdd.n2527 gnd 0.007362f
C4669 vdd.n2528 gnd 0.007362f
C4670 vdd.n2529 gnd 0.005359f
C4671 vdd.n2530 gnd 0.007362f
C4672 vdd.n2531 gnd 0.007362f
C4673 vdd.n2532 gnd 0.007362f
C4674 vdd.n2533 gnd 0.007362f
C4675 vdd.n2534 gnd 0.007362f
C4676 vdd.n2535 gnd 0.007362f
C4677 vdd.n2536 gnd 0.007362f
C4678 vdd.n2537 gnd 0.007362f
C4679 vdd.n2538 gnd 0.007362f
C4680 vdd.n2539 gnd 0.007362f
C4681 vdd.n2540 gnd 0.007362f
C4682 vdd.n2541 gnd 0.007362f
C4683 vdd.n2542 gnd 0.007362f
C4684 vdd.n2543 gnd 0.007362f
C4685 vdd.n2544 gnd 0.007362f
C4686 vdd.n2545 gnd 0.007362f
C4687 vdd.n2546 gnd 0.007362f
C4688 vdd.n2547 gnd 0.007362f
C4689 vdd.n2548 gnd 0.007362f
C4690 vdd.n2549 gnd 0.007362f
C4691 vdd.n2550 gnd 0.007362f
C4692 vdd.n2551 gnd 0.007362f
C4693 vdd.n2552 gnd 0.007362f
C4694 vdd.n2553 gnd 0.007362f
C4695 vdd.n2554 gnd 0.007362f
C4696 vdd.n2555 gnd 0.007362f
C4697 vdd.n2556 gnd 0.007362f
C4698 vdd.n2557 gnd 0.007362f
C4699 vdd.n2558 gnd 0.007362f
C4700 vdd.n2559 gnd 0.007362f
C4701 vdd.n2560 gnd 0.007362f
C4702 vdd.n2561 gnd 0.007362f
C4703 vdd.n2562 gnd 0.007362f
C4704 vdd.n2563 gnd 0.007362f
C4705 vdd.n2564 gnd 0.007362f
C4706 vdd.n2565 gnd 0.007362f
C4707 vdd.n2566 gnd 0.007362f
C4708 vdd.n2567 gnd 0.007362f
C4709 vdd.n2568 gnd 0.007362f
C4710 vdd.n2569 gnd 0.007362f
C4711 vdd.n2570 gnd 0.007362f
C4712 vdd.n2571 gnd 0.007362f
C4713 vdd.n2572 gnd 0.007362f
C4714 vdd.n2573 gnd 0.007362f
C4715 vdd.n2574 gnd 0.007362f
C4716 vdd.n2575 gnd 0.007362f
C4717 vdd.n2576 gnd 0.007362f
C4718 vdd.n2577 gnd 0.007362f
C4719 vdd.n2578 gnd 0.007362f
C4720 vdd.n2579 gnd 0.007362f
C4721 vdd.n2580 gnd 0.007362f
C4722 vdd.n2581 gnd 0.007362f
C4723 vdd.n2582 gnd 0.007362f
C4724 vdd.n2583 gnd 0.007362f
C4725 vdd.n2584 gnd 0.007362f
C4726 vdd.n2585 gnd 0.007362f
C4727 vdd.n2586 gnd 0.007362f
C4728 vdd.n2587 gnd 0.007362f
C4729 vdd.n2588 gnd 0.007362f
C4730 vdd.n2589 gnd 0.007362f
C4731 vdd.n2590 gnd 0.017219f
C4732 vdd.n2591 gnd 0.016126f
C4733 vdd.n2592 gnd 0.016126f
C4734 vdd.n2593 gnd 0.896159f
C4735 vdd.n2594 gnd 0.016126f
C4736 vdd.n2595 gnd 0.017219f
C4737 vdd.n2596 gnd 0.016304f
C4738 vdd.n2597 gnd 0.007362f
C4739 vdd.n2598 gnd 0.007362f
C4740 vdd.n2599 gnd 0.007362f
C4741 vdd.n2600 gnd 0.005684f
C4742 vdd.n2601 gnd 0.010521f
C4743 vdd.n2602 gnd 0.005359f
C4744 vdd.n2603 gnd 0.007362f
C4745 vdd.n2604 gnd 0.007362f
C4746 vdd.n2605 gnd 0.007362f
C4747 vdd.n2606 gnd 0.007362f
C4748 vdd.n2607 gnd 0.007362f
C4749 vdd.n2608 gnd 0.007362f
C4750 vdd.n2609 gnd 0.007362f
C4751 vdd.n2610 gnd 0.007362f
C4752 vdd.n2611 gnd 0.007362f
C4753 vdd.n2612 gnd 0.007362f
C4754 vdd.n2613 gnd 0.007362f
C4755 vdd.n2614 gnd 0.007362f
C4756 vdd.n2615 gnd 0.007362f
C4757 vdd.n2616 gnd 0.007362f
C4758 vdd.n2617 gnd 0.007362f
C4759 vdd.n2618 gnd 0.007362f
C4760 vdd.n2619 gnd 0.007362f
C4761 vdd.n2620 gnd 0.007362f
C4762 vdd.n2621 gnd 0.007362f
C4763 vdd.n2622 gnd 0.007362f
C4764 vdd.n2623 gnd 0.007362f
C4765 vdd.n2624 gnd 0.007362f
C4766 vdd.n2625 gnd 0.007362f
C4767 vdd.n2626 gnd 0.007362f
C4768 vdd.n2627 gnd 0.007362f
C4769 vdd.n2628 gnd 0.007362f
C4770 vdd.n2629 gnd 0.007362f
C4771 vdd.n2630 gnd 0.007362f
C4772 vdd.n2631 gnd 0.007362f
C4773 vdd.n2632 gnd 0.007362f
C4774 vdd.n2633 gnd 0.007362f
C4775 vdd.n2634 gnd 0.007362f
C4776 vdd.n2635 gnd 0.007362f
C4777 vdd.n2636 gnd 0.007362f
C4778 vdd.n2637 gnd 0.007362f
C4779 vdd.n2638 gnd 0.007362f
C4780 vdd.n2639 gnd 0.007362f
C4781 vdd.n2640 gnd 0.007362f
C4782 vdd.n2641 gnd 0.007362f
C4783 vdd.n2642 gnd 0.007362f
C4784 vdd.n2643 gnd 0.007362f
C4785 vdd.n2644 gnd 0.007362f
C4786 vdd.n2645 gnd 0.007362f
C4787 vdd.n2646 gnd 0.007362f
C4788 vdd.n2647 gnd 0.007362f
C4789 vdd.n2648 gnd 0.007362f
C4790 vdd.n2649 gnd 0.007362f
C4791 vdd.n2650 gnd 0.007362f
C4792 vdd.n2651 gnd 0.007362f
C4793 vdd.n2652 gnd 0.007362f
C4794 vdd.n2653 gnd 0.007362f
C4795 vdd.n2654 gnd 0.007362f
C4796 vdd.n2655 gnd 0.007362f
C4797 vdd.n2656 gnd 0.007362f
C4798 vdd.n2657 gnd 0.007362f
C4799 vdd.n2658 gnd 0.007362f
C4800 vdd.n2659 gnd 0.007362f
C4801 vdd.n2660 gnd 0.007362f
C4802 vdd.n2661 gnd 0.007362f
C4803 vdd.n2662 gnd 0.007362f
C4804 vdd.n2663 gnd 0.017219f
C4805 vdd.n2664 gnd 0.017219f
C4806 vdd.n2665 gnd 0.918287f
C4807 vdd.t209 gnd 3.26379f
C4808 vdd.t293 gnd 3.26379f
C4809 vdd.n2698 gnd 0.017219f
C4810 vdd.t196 gnd 0.685949f
C4811 vdd.n2699 gnd 0.007362f
C4812 vdd.n2700 gnd 0.007362f
C4813 vdd.t269 gnd 0.297485f
C4814 vdd.t270 gnd 0.304513f
C4815 vdd.t267 gnd 0.19421f
C4816 vdd.n2701 gnd 0.10496f
C4817 vdd.n2702 gnd 0.059537f
C4818 vdd.n2703 gnd 0.007362f
C4819 vdd.t282 gnd 0.297485f
C4820 vdd.t283 gnd 0.304513f
C4821 vdd.t281 gnd 0.19421f
C4822 vdd.n2704 gnd 0.10496f
C4823 vdd.n2705 gnd 0.059537f
C4824 vdd.n2706 gnd 0.010521f
C4825 vdd.n2707 gnd 0.007362f
C4826 vdd.n2708 gnd 0.007362f
C4827 vdd.n2709 gnd 0.007362f
C4828 vdd.n2710 gnd 0.007362f
C4829 vdd.n2711 gnd 0.007362f
C4830 vdd.n2712 gnd 0.007362f
C4831 vdd.n2713 gnd 0.007362f
C4832 vdd.n2714 gnd 0.007362f
C4833 vdd.n2715 gnd 0.007362f
C4834 vdd.n2716 gnd 0.007362f
C4835 vdd.n2717 gnd 0.007362f
C4836 vdd.n2718 gnd 0.007362f
C4837 vdd.n2719 gnd 0.007362f
C4838 vdd.n2720 gnd 0.007362f
C4839 vdd.n2721 gnd 0.007362f
C4840 vdd.n2722 gnd 0.007362f
C4841 vdd.n2723 gnd 0.007362f
C4842 vdd.n2724 gnd 0.007362f
C4843 vdd.n2725 gnd 0.007362f
C4844 vdd.n2726 gnd 0.007362f
C4845 vdd.n2727 gnd 0.007362f
C4846 vdd.n2728 gnd 0.007362f
C4847 vdd.n2729 gnd 0.007362f
C4848 vdd.n2730 gnd 0.007362f
C4849 vdd.n2731 gnd 0.007362f
C4850 vdd.n2732 gnd 0.007362f
C4851 vdd.n2733 gnd 0.007362f
C4852 vdd.n2734 gnd 0.007362f
C4853 vdd.n2735 gnd 0.007362f
C4854 vdd.n2736 gnd 0.007362f
C4855 vdd.n2737 gnd 0.007362f
C4856 vdd.n2738 gnd 0.007362f
C4857 vdd.n2739 gnd 0.007362f
C4858 vdd.n2740 gnd 0.007362f
C4859 vdd.n2741 gnd 0.007362f
C4860 vdd.n2742 gnd 0.007362f
C4861 vdd.n2743 gnd 0.007362f
C4862 vdd.n2744 gnd 0.007362f
C4863 vdd.n2745 gnd 0.007362f
C4864 vdd.n2746 gnd 0.007362f
C4865 vdd.n2747 gnd 0.007362f
C4866 vdd.n2748 gnd 0.007362f
C4867 vdd.n2749 gnd 0.007362f
C4868 vdd.n2750 gnd 0.007362f
C4869 vdd.n2751 gnd 0.007362f
C4870 vdd.n2752 gnd 0.007362f
C4871 vdd.n2753 gnd 0.007362f
C4872 vdd.n2754 gnd 0.007362f
C4873 vdd.n2755 gnd 0.007362f
C4874 vdd.n2756 gnd 0.007362f
C4875 vdd.n2757 gnd 0.007362f
C4876 vdd.n2758 gnd 0.007362f
C4877 vdd.n2759 gnd 0.007362f
C4878 vdd.n2760 gnd 0.007362f
C4879 vdd.n2761 gnd 0.007362f
C4880 vdd.n2762 gnd 0.007362f
C4881 vdd.n2763 gnd 0.007362f
C4882 vdd.n2764 gnd 0.007362f
C4883 vdd.n2765 gnd 0.005359f
C4884 vdd.n2766 gnd 0.007362f
C4885 vdd.n2767 gnd 0.007362f
C4886 vdd.n2768 gnd 0.005684f
C4887 vdd.n2769 gnd 0.007362f
C4888 vdd.n2770 gnd 0.007362f
C4889 vdd.n2771 gnd 0.017219f
C4890 vdd.n2772 gnd 0.016126f
C4891 vdd.n2773 gnd 0.016126f
C4892 vdd.n2774 gnd 0.007362f
C4893 vdd.n2775 gnd 0.007362f
C4894 vdd.n2776 gnd 0.007362f
C4895 vdd.n2777 gnd 0.007362f
C4896 vdd.n2778 gnd 0.007362f
C4897 vdd.n2779 gnd 0.007362f
C4898 vdd.n2780 gnd 0.007362f
C4899 vdd.n2781 gnd 0.007362f
C4900 vdd.n2782 gnd 0.007362f
C4901 vdd.n2783 gnd 0.007362f
C4902 vdd.n2784 gnd 0.007362f
C4903 vdd.n2785 gnd 0.007362f
C4904 vdd.n2786 gnd 0.007362f
C4905 vdd.n2787 gnd 0.007362f
C4906 vdd.n2788 gnd 0.007362f
C4907 vdd.n2789 gnd 0.007362f
C4908 vdd.n2790 gnd 0.007362f
C4909 vdd.n2791 gnd 0.007362f
C4910 vdd.n2792 gnd 0.007362f
C4911 vdd.n2793 gnd 0.007362f
C4912 vdd.n2794 gnd 0.007362f
C4913 vdd.n2795 gnd 0.007362f
C4914 vdd.n2796 gnd 0.007362f
C4915 vdd.n2797 gnd 0.007362f
C4916 vdd.n2798 gnd 0.007362f
C4917 vdd.n2799 gnd 0.007362f
C4918 vdd.n2800 gnd 0.007362f
C4919 vdd.n2801 gnd 0.007362f
C4920 vdd.n2802 gnd 0.007362f
C4921 vdd.n2803 gnd 0.007362f
C4922 vdd.n2804 gnd 0.007362f
C4923 vdd.n2805 gnd 0.007362f
C4924 vdd.n2806 gnd 0.007362f
C4925 vdd.n2807 gnd 0.007362f
C4926 vdd.n2808 gnd 0.007362f
C4927 vdd.n2809 gnd 0.007362f
C4928 vdd.n2810 gnd 0.007362f
C4929 vdd.n2811 gnd 0.007362f
C4930 vdd.n2812 gnd 0.007362f
C4931 vdd.n2813 gnd 0.007362f
C4932 vdd.n2814 gnd 0.007362f
C4933 vdd.n2815 gnd 0.007362f
C4934 vdd.n2816 gnd 0.007362f
C4935 vdd.n2817 gnd 0.007362f
C4936 vdd.n2818 gnd 0.007362f
C4937 vdd.n2819 gnd 0.007362f
C4938 vdd.n2820 gnd 0.007362f
C4939 vdd.n2821 gnd 0.007362f
C4940 vdd.n2822 gnd 0.007362f
C4941 vdd.n2823 gnd 0.007362f
C4942 vdd.n2824 gnd 0.007362f
C4943 vdd.n2825 gnd 0.007362f
C4944 vdd.n2826 gnd 0.007362f
C4945 vdd.n2827 gnd 0.007362f
C4946 vdd.n2828 gnd 0.007362f
C4947 vdd.n2829 gnd 0.007362f
C4948 vdd.n2830 gnd 0.007362f
C4949 vdd.n2831 gnd 0.007362f
C4950 vdd.n2832 gnd 0.007362f
C4951 vdd.n2833 gnd 0.007362f
C4952 vdd.n2834 gnd 0.007362f
C4953 vdd.n2835 gnd 0.007362f
C4954 vdd.n2836 gnd 0.007362f
C4955 vdd.n2837 gnd 0.007362f
C4956 vdd.n2838 gnd 0.007362f
C4957 vdd.n2839 gnd 0.007362f
C4958 vdd.n2840 gnd 0.007362f
C4959 vdd.n2841 gnd 0.007362f
C4960 vdd.n2842 gnd 0.007362f
C4961 vdd.n2843 gnd 0.007362f
C4962 vdd.n2844 gnd 0.007362f
C4963 vdd.n2845 gnd 0.007362f
C4964 vdd.n2846 gnd 0.007362f
C4965 vdd.n2847 gnd 0.237869f
C4966 vdd.n2848 gnd 0.007362f
C4967 vdd.n2849 gnd 0.007362f
C4968 vdd.n2850 gnd 0.007362f
C4969 vdd.n2851 gnd 0.007362f
C4970 vdd.n2852 gnd 0.007362f
C4971 vdd.n2853 gnd 0.007362f
C4972 vdd.n2854 gnd 0.007362f
C4973 vdd.n2855 gnd 0.007362f
C4974 vdd.n2856 gnd 0.007362f
C4975 vdd.n2857 gnd 0.007362f
C4976 vdd.n2858 gnd 0.007362f
C4977 vdd.n2859 gnd 0.007362f
C4978 vdd.n2860 gnd 0.007362f
C4979 vdd.n2861 gnd 0.007362f
C4980 vdd.n2862 gnd 0.470207f
C4981 vdd.n2863 gnd 0.007362f
C4982 vdd.n2864 gnd 0.007362f
C4983 vdd.n2865 gnd 0.007362f
C4984 vdd.n2866 gnd 0.016126f
C4985 vdd.n2867 gnd 0.016126f
C4986 vdd.n2868 gnd 0.017219f
C4987 vdd.n2869 gnd 0.017219f
C4988 vdd.n2870 gnd 0.007362f
C4989 vdd.n2871 gnd 0.007362f
C4990 vdd.n2872 gnd 0.007362f
C4991 vdd.n2873 gnd 0.005684f
C4992 vdd.n2874 gnd 0.010521f
C4993 vdd.n2875 gnd 0.005359f
C4994 vdd.n2876 gnd 0.007362f
C4995 vdd.n2877 gnd 0.007362f
C4996 vdd.n2878 gnd 0.007362f
C4997 vdd.n2879 gnd 0.007362f
C4998 vdd.n2880 gnd 0.007362f
C4999 vdd.n2881 gnd 0.007362f
C5000 vdd.n2882 gnd 0.007362f
C5001 vdd.n2883 gnd 0.007362f
C5002 vdd.n2884 gnd 0.007362f
C5003 vdd.n2885 gnd 0.007362f
C5004 vdd.n2886 gnd 0.007362f
C5005 vdd.n2887 gnd 0.007362f
C5006 vdd.n2888 gnd 0.007362f
C5007 vdd.n2889 gnd 0.007362f
C5008 vdd.n2890 gnd 0.007362f
C5009 vdd.n2891 gnd 0.007362f
C5010 vdd.n2892 gnd 0.007362f
C5011 vdd.n2893 gnd 0.007362f
C5012 vdd.n2894 gnd 0.007362f
C5013 vdd.n2895 gnd 0.007362f
C5014 vdd.n2896 gnd 0.007362f
C5015 vdd.n2897 gnd 0.007362f
C5016 vdd.n2898 gnd 0.007362f
C5017 vdd.n2899 gnd 0.007362f
C5018 vdd.n2900 gnd 0.007362f
C5019 vdd.n2901 gnd 0.007362f
C5020 vdd.n2902 gnd 0.007362f
C5021 vdd.n2903 gnd 0.007362f
C5022 vdd.n2904 gnd 0.007362f
C5023 vdd.n2905 gnd 0.007362f
C5024 vdd.n2906 gnd 0.007362f
C5025 vdd.n2907 gnd 0.007362f
C5026 vdd.n2908 gnd 0.007362f
C5027 vdd.n2909 gnd 0.007362f
C5028 vdd.n2910 gnd 0.007362f
C5029 vdd.n2911 gnd 0.007362f
C5030 vdd.n2912 gnd 0.007362f
C5031 vdd.n2913 gnd 0.007362f
C5032 vdd.n2914 gnd 0.007362f
C5033 vdd.n2915 gnd 0.007362f
C5034 vdd.n2916 gnd 0.007362f
C5035 vdd.n2917 gnd 0.007362f
C5036 vdd.n2918 gnd 0.007362f
C5037 vdd.n2919 gnd 0.007362f
C5038 vdd.n2920 gnd 0.007362f
C5039 vdd.n2921 gnd 0.007362f
C5040 vdd.n2922 gnd 0.007362f
C5041 vdd.n2923 gnd 0.007362f
C5042 vdd.n2924 gnd 0.007362f
C5043 vdd.n2925 gnd 0.007362f
C5044 vdd.n2926 gnd 0.007362f
C5045 vdd.n2927 gnd 0.007362f
C5046 vdd.n2928 gnd 0.007362f
C5047 vdd.n2929 gnd 0.007362f
C5048 vdd.n2930 gnd 0.007362f
C5049 vdd.n2931 gnd 0.007362f
C5050 vdd.n2932 gnd 0.007362f
C5051 vdd.n2933 gnd 0.007362f
C5052 vdd.n2934 gnd 0.007362f
C5053 vdd.n2935 gnd 0.017219f
C5054 vdd.n2936 gnd 0.017219f
C5055 vdd.n2938 gnd 0.918287f
C5056 vdd.n2940 gnd 0.017219f
C5057 vdd.n2941 gnd 0.017219f
C5058 vdd.n2942 gnd 0.016126f
C5059 vdd.n2943 gnd 0.007362f
C5060 vdd.n2944 gnd 0.007362f
C5061 vdd.n2945 gnd 0.398293f
C5062 vdd.n2946 gnd 0.007362f
C5063 vdd.n2947 gnd 0.007362f
C5064 vdd.n2948 gnd 0.007362f
C5065 vdd.n2949 gnd 0.007362f
C5066 vdd.n2950 gnd 0.007362f
C5067 vdd.n2951 gnd 0.44808f
C5068 vdd.n2952 gnd 0.007362f
C5069 vdd.n2953 gnd 0.007362f
C5070 vdd.n2954 gnd 0.007362f
C5071 vdd.n2955 gnd 0.007362f
C5072 vdd.n2956 gnd 0.007362f
C5073 vdd.n2957 gnd 0.752331f
C5074 vdd.n2958 gnd 0.007362f
C5075 vdd.n2959 gnd 0.007362f
C5076 vdd.n2960 gnd 0.007362f
C5077 vdd.n2961 gnd 0.007362f
C5078 vdd.n2962 gnd 0.007362f
C5079 vdd.n2963 gnd 0.497866f
C5080 vdd.n2964 gnd 0.007362f
C5081 vdd.n2965 gnd 0.007362f
C5082 vdd.n2966 gnd 0.007362f
C5083 vdd.n2967 gnd 0.007362f
C5084 vdd.n2968 gnd 0.007362f
C5085 vdd.n2969 gnd 0.663822f
C5086 vdd.n2970 gnd 0.007362f
C5087 vdd.n2971 gnd 0.007362f
C5088 vdd.n2972 gnd 0.007362f
C5089 vdd.n2973 gnd 0.007362f
C5090 vdd.n2974 gnd 0.007362f
C5091 vdd.n2975 gnd 0.602971f
C5092 vdd.n2976 gnd 0.007362f
C5093 vdd.n2977 gnd 0.007362f
C5094 vdd.n2978 gnd 0.007362f
C5095 vdd.n2979 gnd 0.007362f
C5096 vdd.n2980 gnd 0.007362f
C5097 vdd.n2981 gnd 0.437016f
C5098 vdd.n2982 gnd 0.007362f
C5099 vdd.n2983 gnd 0.007362f
C5100 vdd.n2984 gnd 0.007362f
C5101 vdd.n2985 gnd 0.007362f
C5102 vdd.n2986 gnd 0.007362f
C5103 vdd.n2987 gnd 0.237869f
C5104 vdd.n2988 gnd 0.007362f
C5105 vdd.n2989 gnd 0.007362f
C5106 vdd.n2990 gnd 0.007362f
C5107 vdd.n2991 gnd 0.007362f
C5108 vdd.n2992 gnd 0.007362f
C5109 vdd.n2993 gnd 0.647226f
C5110 vdd.n2994 gnd 0.007362f
C5111 vdd.n2995 gnd 0.007362f
C5112 vdd.n2996 gnd 0.007362f
C5113 vdd.n2997 gnd 0.007362f
C5114 vdd.n2998 gnd 0.007362f
C5115 vdd.n2999 gnd 0.752331f
C5116 vdd.n3000 gnd 0.007362f
C5117 vdd.n3001 gnd 0.007362f
C5118 vdd.n3002 gnd 0.004763f
C5119 vdd.n3003 gnd 0.021326f
C5120 vdd.n3004 gnd 0.006279f
C5121 vdd.n3005 gnd 0.007362f
C5122 vdd.n3006 gnd 0.641694f
C5123 vdd.n3007 gnd 0.007362f
C5124 vdd.n3008 gnd 0.007362f
C5125 vdd.n3009 gnd 0.007362f
C5126 vdd.n3010 gnd 0.007362f
C5127 vdd.n3011 gnd 0.007362f
C5128 vdd.n3012 gnd 0.525526f
C5129 vdd.n3013 gnd 0.007362f
C5130 vdd.n3014 gnd 0.007362f
C5131 vdd.n3015 gnd 0.007362f
C5132 vdd.n3016 gnd 0.007362f
C5133 vdd.n3017 gnd 0.007362f
C5134 vdd.n3018 gnd 0.392761f
C5135 vdd.n3019 gnd 0.007362f
C5136 vdd.n3020 gnd 0.007362f
C5137 vdd.n3021 gnd 0.007362f
C5138 vdd.n3022 gnd 0.007362f
C5139 vdd.n3023 gnd 0.007362f
C5140 vdd.n3024 gnd 0.752331f
C5141 vdd.n3025 gnd 0.007362f
C5142 vdd.n3026 gnd 0.007362f
C5143 vdd.n3027 gnd 0.007362f
C5144 vdd.n3028 gnd 0.007362f
C5145 vdd.n3029 gnd 0.007362f
C5146 vdd.n3030 gnd 0.007362f
C5147 vdd.n3032 gnd 0.007362f
C5148 vdd.n3033 gnd 0.007362f
C5149 vdd.n3035 gnd 0.007362f
C5150 vdd.n3036 gnd 0.007362f
C5151 vdd.n3039 gnd 0.007362f
C5152 vdd.n3040 gnd 0.007362f
C5153 vdd.n3041 gnd 0.007362f
C5154 vdd.n3042 gnd 0.007362f
C5155 vdd.n3044 gnd 0.007362f
C5156 vdd.n3045 gnd 0.007362f
C5157 vdd.n3046 gnd 0.007362f
C5158 vdd.n3047 gnd 0.007362f
C5159 vdd.n3048 gnd 0.007362f
C5160 vdd.n3049 gnd 0.007362f
C5161 vdd.n3051 gnd 0.007362f
C5162 vdd.n3052 gnd 0.007362f
C5163 vdd.n3053 gnd 0.007362f
C5164 vdd.n3054 gnd 0.007362f
C5165 vdd.n3055 gnd 0.007362f
C5166 vdd.n3056 gnd 0.007362f
C5167 vdd.n3058 gnd 0.007362f
C5168 vdd.n3059 gnd 0.007362f
C5169 vdd.n3060 gnd 0.007362f
C5170 vdd.n3061 gnd 0.007362f
C5171 vdd.n3062 gnd 0.007362f
C5172 vdd.n3063 gnd 0.007362f
C5173 vdd.n3065 gnd 0.007362f
C5174 vdd.n3066 gnd 0.017219f
C5175 vdd.n3067 gnd 0.017219f
C5176 vdd.n3068 gnd 0.016126f
C5177 vdd.n3069 gnd 0.007362f
C5178 vdd.n3070 gnd 0.007362f
C5179 vdd.n3071 gnd 0.007362f
C5180 vdd.n3072 gnd 0.007362f
C5181 vdd.n3073 gnd 0.007362f
C5182 vdd.n3074 gnd 0.007362f
C5183 vdd.n3075 gnd 0.752331f
C5184 vdd.n3076 gnd 0.007362f
C5185 vdd.n3077 gnd 0.007362f
C5186 vdd.n3078 gnd 0.007362f
C5187 vdd.n3079 gnd 0.007362f
C5188 vdd.n3080 gnd 0.007362f
C5189 vdd.n3081 gnd 0.492334f
C5190 vdd.n3082 gnd 0.007362f
C5191 vdd.n3083 gnd 0.007362f
C5192 vdd.n3084 gnd 0.007362f
C5193 vdd.n3085 gnd 0.01704f
C5194 vdd.n3086 gnd 0.016304f
C5195 vdd.n3087 gnd 0.017219f
C5196 vdd.n3089 gnd 0.007362f
C5197 vdd.n3090 gnd 0.007362f
C5198 vdd.n3091 gnd 0.005684f
C5199 vdd.n3092 gnd 0.010521f
C5200 vdd.n3093 gnd 0.005359f
C5201 vdd.n3094 gnd 0.007362f
C5202 vdd.n3095 gnd 0.007362f
C5203 vdd.n3097 gnd 0.007362f
C5204 vdd.n3098 gnd 0.007362f
C5205 vdd.n3099 gnd 0.007362f
C5206 vdd.n3100 gnd 0.007362f
C5207 vdd.n3101 gnd 0.007362f
C5208 vdd.n3102 gnd 0.007362f
C5209 vdd.n3104 gnd 0.007362f
C5210 vdd.n3105 gnd 0.007362f
C5211 vdd.n3106 gnd 0.007362f
C5212 vdd.n3107 gnd 0.007362f
C5213 vdd.n3108 gnd 0.007362f
C5214 vdd.n3109 gnd 0.007362f
C5215 vdd.n3111 gnd 0.007362f
C5216 vdd.n3112 gnd 0.007362f
C5217 vdd.n3113 gnd 0.007362f
C5218 vdd.n3114 gnd 0.007362f
C5219 vdd.n3115 gnd 0.007362f
C5220 vdd.n3116 gnd 0.007362f
C5221 vdd.n3118 gnd 0.007362f
C5222 vdd.n3119 gnd 0.007362f
C5223 vdd.n3120 gnd 0.007362f
C5224 vdd.n3122 gnd 0.007362f
C5225 vdd.n3123 gnd 0.007362f
C5226 vdd.n3124 gnd 0.007362f
C5227 vdd.n3125 gnd 0.007362f
C5228 vdd.n3126 gnd 0.007362f
C5229 vdd.n3127 gnd 0.007362f
C5230 vdd.n3129 gnd 0.007362f
C5231 vdd.n3130 gnd 0.007362f
C5232 vdd.n3131 gnd 0.007362f
C5233 vdd.n3132 gnd 0.007362f
C5234 vdd.n3133 gnd 0.007362f
C5235 vdd.n3134 gnd 0.007362f
C5236 vdd.n3136 gnd 0.007362f
C5237 vdd.n3137 gnd 0.007362f
C5238 vdd.n3138 gnd 0.007362f
C5239 vdd.n3139 gnd 0.007362f
C5240 vdd.n3140 gnd 0.007362f
C5241 vdd.n3141 gnd 0.007362f
C5242 vdd.n3143 gnd 0.007362f
C5243 vdd.n3144 gnd 0.007362f
C5244 vdd.n3146 gnd 0.007362f
C5245 vdd.n3147 gnd 0.007362f
C5246 vdd.n3148 gnd 0.017219f
C5247 vdd.n3149 gnd 0.016126f
C5248 vdd.n3150 gnd 0.016126f
C5249 vdd.n3151 gnd 1.06211f
C5250 vdd.n3152 gnd 0.016126f
C5251 vdd.n3153 gnd 0.017219f
C5252 vdd.n3154 gnd 0.016304f
C5253 vdd.n3155 gnd 0.007362f
C5254 vdd.n3156 gnd 0.005684f
C5255 vdd.n3157 gnd 0.007362f
C5256 vdd.n3159 gnd 0.007362f
C5257 vdd.n3160 gnd 0.007362f
C5258 vdd.n3161 gnd 0.007362f
C5259 vdd.n3162 gnd 0.007362f
C5260 vdd.n3163 gnd 0.007362f
C5261 vdd.n3164 gnd 0.007362f
C5262 vdd.n3166 gnd 0.007362f
C5263 vdd.n3167 gnd 0.007362f
C5264 vdd.n3168 gnd 0.007362f
C5265 vdd.n3169 gnd 0.007362f
C5266 vdd.n3170 gnd 0.007362f
C5267 vdd.n3171 gnd 0.007362f
C5268 vdd.n3173 gnd 0.007362f
C5269 vdd.n3174 gnd 0.007362f
C5270 vdd.n3175 gnd 0.007362f
C5271 vdd.n3176 gnd 0.007362f
C5272 vdd.n3177 gnd 0.007362f
C5273 vdd.n3178 gnd 0.007362f
C5274 vdd.n3180 gnd 0.007362f
C5275 vdd.n3181 gnd 0.007362f
C5276 vdd.n3183 gnd 0.007362f
C5277 vdd.n3184 gnd 0.025283f
C5278 vdd.n3185 gnd 0.822946f
C5279 vdd.n3187 gnd 0.004575f
C5280 vdd.n3188 gnd 0.008714f
C5281 vdd.n3189 gnd 0.010826f
C5282 vdd.n3190 gnd 0.010826f
C5283 vdd.n3191 gnd 0.008714f
C5284 vdd.n3192 gnd 0.008714f
C5285 vdd.n3193 gnd 0.010826f
C5286 vdd.n3194 gnd 0.010826f
C5287 vdd.n3195 gnd 0.008714f
C5288 vdd.n3196 gnd 0.008714f
C5289 vdd.n3197 gnd 0.010826f
C5290 vdd.n3198 gnd 0.010826f
C5291 vdd.n3199 gnd 0.008714f
C5292 vdd.n3200 gnd 0.008714f
C5293 vdd.n3201 gnd 0.010826f
C5294 vdd.n3202 gnd 0.010826f
C5295 vdd.n3203 gnd 0.008714f
C5296 vdd.n3204 gnd 0.008714f
C5297 vdd.n3205 gnd 0.010826f
C5298 vdd.n3206 gnd 0.010826f
C5299 vdd.n3207 gnd 0.008714f
C5300 vdd.n3208 gnd 0.008714f
C5301 vdd.n3209 gnd 0.010826f
C5302 vdd.n3210 gnd 0.010826f
C5303 vdd.n3211 gnd 0.008714f
C5304 vdd.n3212 gnd 0.008714f
C5305 vdd.n3213 gnd 0.010826f
C5306 vdd.n3214 gnd 0.010826f
C5307 vdd.n3215 gnd 0.008714f
C5308 vdd.n3216 gnd 0.008714f
C5309 vdd.n3217 gnd 0.010826f
C5310 vdd.n3218 gnd 0.010826f
C5311 vdd.n3219 gnd 0.008714f
C5312 vdd.n3220 gnd 0.008714f
C5313 vdd.n3221 gnd 0.010826f
C5314 vdd.n3222 gnd 0.010826f
C5315 vdd.n3223 gnd 0.008714f
C5316 vdd.n3224 gnd 0.010826f
C5317 vdd.n3225 gnd 0.010826f
C5318 vdd.n3226 gnd 0.008714f
C5319 vdd.n3227 gnd 0.010826f
C5320 vdd.n3228 gnd 0.010826f
C5321 vdd.n3229 gnd 0.010826f
C5322 vdd.n3230 gnd 0.017776f
C5323 vdd.n3231 gnd 0.010826f
C5324 vdd.n3232 gnd 0.010826f
C5325 vdd.n3233 gnd 0.005925f
C5326 vdd.n3234 gnd 0.008714f
C5327 vdd.n3235 gnd 0.010826f
C5328 vdd.n3236 gnd 0.010826f
C5329 vdd.n3237 gnd 0.008714f
C5330 vdd.n3238 gnd 0.008714f
C5331 vdd.n3239 gnd 0.010826f
C5332 vdd.n3240 gnd 0.010826f
C5333 vdd.n3241 gnd 0.008714f
C5334 vdd.n3242 gnd 0.008714f
C5335 vdd.n3243 gnd 0.010826f
C5336 vdd.n3244 gnd 0.010826f
C5337 vdd.n3245 gnd 0.008714f
C5338 vdd.n3246 gnd 0.008714f
C5339 vdd.n3247 gnd 0.010826f
C5340 vdd.n3248 gnd 0.010826f
C5341 vdd.n3249 gnd 0.008714f
C5342 vdd.n3250 gnd 0.008714f
C5343 vdd.n3251 gnd 0.010826f
C5344 vdd.n3252 gnd 0.010826f
C5345 vdd.n3253 gnd 0.008714f
C5346 vdd.n3254 gnd 0.008714f
C5347 vdd.n3255 gnd 0.010826f
C5348 vdd.n3256 gnd 0.010826f
C5349 vdd.n3257 gnd 0.008714f
C5350 vdd.n3258 gnd 0.008714f
C5351 vdd.n3259 gnd 0.010826f
C5352 vdd.n3260 gnd 0.010826f
C5353 vdd.n3261 gnd 0.008714f
C5354 vdd.n3262 gnd 0.008714f
C5355 vdd.n3263 gnd 0.010826f
C5356 vdd.n3264 gnd 0.010826f
C5357 vdd.n3265 gnd 0.008714f
C5358 vdd.n3266 gnd 0.008714f
C5359 vdd.n3267 gnd 0.010826f
C5360 vdd.n3268 gnd 0.010826f
C5361 vdd.n3269 gnd 0.008714f
C5362 vdd.n3270 gnd 0.010826f
C5363 vdd.n3271 gnd 0.010826f
C5364 vdd.n3272 gnd 0.008714f
C5365 vdd.n3273 gnd 0.010826f
C5366 vdd.n3274 gnd 0.010826f
C5367 vdd.n3275 gnd 0.010826f
C5368 vdd.t248 gnd 0.133189f
C5369 vdd.t249 gnd 0.142342f
C5370 vdd.t247 gnd 0.173943f
C5371 vdd.n3276 gnd 0.22297f
C5372 vdd.n3277 gnd 0.187335f
C5373 vdd.n3278 gnd 0.017776f
C5374 vdd.n3279 gnd 0.010826f
C5375 vdd.n3280 gnd 0.010826f
C5376 vdd.n3281 gnd 0.007276f
C5377 vdd.n3282 gnd 0.008714f
C5378 vdd.n3283 gnd 0.010826f
C5379 vdd.n3284 gnd 0.010826f
C5380 vdd.n3285 gnd 0.008714f
C5381 vdd.n3286 gnd 0.008714f
C5382 vdd.n3287 gnd 0.010826f
C5383 vdd.n3288 gnd 0.010826f
C5384 vdd.n3289 gnd 0.008714f
C5385 vdd.n3290 gnd 0.008714f
C5386 vdd.n3291 gnd 0.010826f
C5387 vdd.n3292 gnd 0.010826f
C5388 vdd.n3293 gnd 0.008714f
C5389 vdd.n3294 gnd 0.008714f
C5390 vdd.n3295 gnd 0.010826f
C5391 vdd.n3296 gnd 0.010826f
C5392 vdd.n3297 gnd 0.008714f
C5393 vdd.n3298 gnd 0.008714f
C5394 vdd.n3299 gnd 0.010826f
C5395 vdd.n3300 gnd 0.010826f
C5396 vdd.n3301 gnd 0.008714f
C5397 vdd.n3302 gnd 0.008714f
C5398 vdd.n3303 gnd 0.010826f
C5399 vdd.n3304 gnd 0.010826f
C5400 vdd.n3305 gnd 0.008714f
C5401 vdd.n3306 gnd 0.008714f
C5402 vdd.n3308 gnd 0.822946f
C5403 vdd.n3310 gnd 0.008714f
C5404 vdd.n3311 gnd 0.008714f
C5405 vdd.n3312 gnd 0.007232f
C5406 vdd.n3313 gnd 0.02675f
C5407 vdd.n3315 gnd 9.83562f
C5408 vdd.n3316 gnd 0.02675f
C5409 vdd.n3317 gnd 0.004139f
C5410 vdd.n3318 gnd 0.02675f
C5411 vdd.n3319 gnd 0.026189f
C5412 vdd.n3320 gnd 0.010826f
C5413 vdd.n3321 gnd 0.008714f
C5414 vdd.n3322 gnd 0.010826f
C5415 vdd.n3323 gnd 0.669354f
C5416 vdd.n3324 gnd 0.010826f
C5417 vdd.n3325 gnd 0.008714f
C5418 vdd.n3326 gnd 0.010826f
C5419 vdd.n3327 gnd 0.010826f
C5420 vdd.n3328 gnd 0.010826f
C5421 vdd.n3329 gnd 0.008714f
C5422 vdd.n3330 gnd 0.010826f
C5423 vdd.n3331 gnd 1.10637f
C5424 vdd.n3332 gnd 0.010826f
C5425 vdd.n3333 gnd 0.008714f
C5426 vdd.n3334 gnd 0.010826f
C5427 vdd.n3335 gnd 0.010826f
C5428 vdd.n3336 gnd 0.010826f
C5429 vdd.n3337 gnd 0.008714f
C5430 vdd.n3338 gnd 0.010826f
C5431 vdd.n3339 gnd 0.713608f
C5432 vdd.n3340 gnd 0.757863f
C5433 vdd.n3341 gnd 0.010826f
C5434 vdd.n3342 gnd 0.008714f
C5435 vdd.n3343 gnd 0.010826f
C5436 vdd.n3344 gnd 0.010826f
C5437 vdd.n3345 gnd 0.010826f
C5438 vdd.n3346 gnd 0.008714f
C5439 vdd.n3347 gnd 0.010826f
C5440 vdd.n3348 gnd 0.918287f
C5441 vdd.n3349 gnd 0.010826f
C5442 vdd.n3350 gnd 0.008714f
C5443 vdd.n3351 gnd 0.010826f
C5444 vdd.n3352 gnd 0.010826f
C5445 vdd.n3353 gnd 0.010826f
C5446 vdd.n3354 gnd 0.008714f
C5447 vdd.n3355 gnd 0.010826f
C5448 vdd.t79 gnd 0.553185f
C5449 vdd.n3356 gnd 0.890627f
C5450 vdd.n3357 gnd 0.010826f
C5451 vdd.n3358 gnd 0.008714f
C5452 vdd.n3359 gnd 0.010826f
C5453 vdd.n3360 gnd 0.010826f
C5454 vdd.n3361 gnd 0.010826f
C5455 vdd.n3362 gnd 0.008714f
C5456 vdd.n3363 gnd 0.010826f
C5457 vdd.n3364 gnd 0.702545f
C5458 vdd.n3365 gnd 0.010826f
C5459 vdd.n3366 gnd 0.008714f
C5460 vdd.n3367 gnd 0.010826f
C5461 vdd.n3368 gnd 0.010826f
C5462 vdd.n3369 gnd 0.010826f
C5463 vdd.n3370 gnd 0.008714f
C5464 vdd.n3371 gnd 0.010826f
C5465 vdd.n3372 gnd 0.879564f
C5466 vdd.n3373 gnd 0.591908f
C5467 vdd.n3374 gnd 0.010826f
C5468 vdd.n3375 gnd 0.008714f
C5469 vdd.n3376 gnd 0.010826f
C5470 vdd.n3377 gnd 0.010826f
C5471 vdd.n3378 gnd 0.010826f
C5472 vdd.n3379 gnd 0.008714f
C5473 vdd.n3380 gnd 0.010826f
C5474 vdd.n3381 gnd 0.77999f
C5475 vdd.n3382 gnd 0.010826f
C5476 vdd.n3383 gnd 0.008714f
C5477 vdd.n3384 gnd 0.010826f
C5478 vdd.n3385 gnd 0.010826f
C5479 vdd.n3386 gnd 0.010826f
C5480 vdd.n3387 gnd 0.010826f
C5481 vdd.n3388 gnd 0.010826f
C5482 vdd.n3389 gnd 0.008714f
C5483 vdd.n3390 gnd 0.008714f
C5484 vdd.n3391 gnd 0.010826f
C5485 vdd.t108 gnd 0.553185f
C5486 vdd.n3392 gnd 0.918287f
C5487 vdd.n3393 gnd 0.010826f
C5488 vdd.n3394 gnd 0.008714f
C5489 vdd.n3395 gnd 0.010826f
C5490 vdd.n3396 gnd 0.010826f
C5491 vdd.n3397 gnd 0.010826f
C5492 vdd.n3398 gnd 0.008714f
C5493 vdd.n3399 gnd 0.010826f
C5494 vdd.n3400 gnd 0.8685f
C5495 vdd.n3401 gnd 0.010826f
C5496 vdd.n3402 gnd 0.010826f
C5497 vdd.n3403 gnd 0.008714f
C5498 vdd.n3404 gnd 0.008714f
C5499 vdd.n3405 gnd 0.010826f
C5500 vdd.n3406 gnd 0.010826f
C5501 vdd.n3407 gnd 0.010826f
C5502 vdd.n3408 gnd 0.008714f
C5503 vdd.n3409 gnd 0.010826f
C5504 vdd.n3410 gnd 0.008714f
C5505 vdd.n3411 gnd 0.008714f
C5506 vdd.n3412 gnd 0.010826f
C5507 vdd.n3413 gnd 0.010826f
C5508 vdd.n3414 gnd 0.010826f
C5509 vdd.n3415 gnd 0.008714f
C5510 vdd.n3416 gnd 0.010826f
C5511 vdd.n3417 gnd 0.008714f
C5512 vdd.n3418 gnd 0.008714f
C5513 vdd.n3419 gnd 0.010826f
C5514 vdd.n3420 gnd 0.010826f
C5515 vdd.n3421 gnd 0.010826f
C5516 vdd.n3422 gnd 0.008714f
C5517 vdd.n3423 gnd 0.918287f
C5518 vdd.n3424 gnd 0.010826f
C5519 vdd.n3425 gnd 0.008714f
C5520 vdd.n3426 gnd 0.008714f
C5521 vdd.n3427 gnd 0.010826f
C5522 vdd.n3428 gnd 0.010826f
C5523 vdd.n3429 gnd 0.010826f
C5524 vdd.n3430 gnd 0.008714f
C5525 vdd.n3431 gnd 0.010826f
C5526 vdd.n3432 gnd 0.008714f
C5527 vdd.n3433 gnd 0.008714f
C5528 vdd.n3434 gnd 0.010826f
C5529 vdd.n3435 gnd 0.010826f
C5530 vdd.n3436 gnd 0.010826f
C5531 vdd.n3437 gnd 0.008714f
C5532 vdd.n3438 gnd 0.010826f
C5533 vdd.n3439 gnd 0.008714f
C5534 vdd.n3440 gnd 0.007232f
C5535 vdd.n3441 gnd 0.026189f
C5536 vdd.n3442 gnd 0.02675f
C5537 vdd.n3443 gnd 0.004139f
C5538 vdd.n3444 gnd 0.02675f
C5539 vdd.n3446 gnd 2.6221f
C5540 vdd.n3447 gnd 1.6319f
C5541 vdd.n3448 gnd 0.026189f
C5542 vdd.n3449 gnd 0.007232f
C5543 vdd.n3450 gnd 0.008714f
C5544 vdd.n3451 gnd 0.008714f
C5545 vdd.n3452 gnd 0.010826f
C5546 vdd.n3453 gnd 1.10637f
C5547 vdd.n3454 gnd 1.10637f
C5548 vdd.n3455 gnd 1.01233f
C5549 vdd.n3456 gnd 0.010826f
C5550 vdd.n3457 gnd 0.008714f
C5551 vdd.n3458 gnd 0.008714f
C5552 vdd.n3459 gnd 0.008714f
C5553 vdd.n3460 gnd 0.010826f
C5554 vdd.n3461 gnd 0.824245f
C5555 vdd.t136 gnd 0.553185f
C5556 vdd.n3462 gnd 0.835309f
C5557 vdd.n3463 gnd 0.636162f
C5558 vdd.n3464 gnd 0.010826f
C5559 vdd.n3465 gnd 0.008714f
C5560 vdd.n3466 gnd 0.008714f
C5561 vdd.n3467 gnd 0.008714f
C5562 vdd.n3468 gnd 0.010826f
C5563 vdd.n3469 gnd 0.65829f
C5564 vdd.n3470 gnd 0.813182f
C5565 vdd.t90 gnd 0.553185f
C5566 vdd.n3471 gnd 0.846373f
C5567 vdd.n3472 gnd 0.010826f
C5568 vdd.n3473 gnd 0.008714f
C5569 vdd.n3474 gnd 0.008714f
C5570 vdd.n3475 gnd 0.008714f
C5571 vdd.n3476 gnd 0.010826f
C5572 vdd.n3477 gnd 0.918287f
C5573 vdd.t35 gnd 0.553185f
C5574 vdd.n3478 gnd 0.669354f
C5575 vdd.n3479 gnd 0.802118f
C5576 vdd.n3480 gnd 0.010826f
C5577 vdd.n3481 gnd 0.008714f
C5578 vdd.n3482 gnd 0.008714f
C5579 vdd.n3483 gnd 0.008714f
C5580 vdd.n3484 gnd 0.010826f
C5581 vdd.n3485 gnd 0.614035f
C5582 vdd.t47 gnd 0.553185f
C5583 vdd.n3486 gnd 0.918287f
C5584 vdd.t39 gnd 0.553185f
C5585 vdd.n3487 gnd 0.680417f
C5586 vdd.n3488 gnd 0.010826f
C5587 vdd.n3489 gnd 0.008714f
C5588 vdd.n3490 gnd 0.00832f
C5589 vdd.n3491 gnd 0.63856f
C5590 vdd.n3492 gnd 2.89944f
C5591 a_n8300_8799.t31 gnd 0.112715f
C5592 a_n8300_8799.t21 gnd 0.112715f
C5593 a_n8300_8799.t20 gnd 0.112715f
C5594 a_n8300_8799.n0 gnd 0.998201f
C5595 a_n8300_8799.t26 gnd 0.112715f
C5596 a_n8300_8799.t25 gnd 0.112715f
C5597 a_n8300_8799.n1 gnd 0.995986f
C5598 a_n8300_8799.n2 gnd 0.793351f
C5599 a_n8300_8799.t0 gnd 0.144919f
C5600 a_n8300_8799.t4 gnd 0.144919f
C5601 a_n8300_8799.n3 gnd 1.143f
C5602 a_n8300_8799.t2 gnd 0.144919f
C5603 a_n8300_8799.t5 gnd 0.144919f
C5604 a_n8300_8799.n4 gnd 1.14111f
C5605 a_n8300_8799.n5 gnd 1.02572f
C5606 a_n8300_8799.t7 gnd 0.144919f
C5607 a_n8300_8799.t8 gnd 0.144919f
C5608 a_n8300_8799.n6 gnd 1.14111f
C5609 a_n8300_8799.n7 gnd 0.505597f
C5610 a_n8300_8799.t12 gnd 0.144919f
C5611 a_n8300_8799.t10 gnd 0.144919f
C5612 a_n8300_8799.n8 gnd 1.14111f
C5613 a_n8300_8799.n9 gnd 3.23842f
C5614 a_n8300_8799.t39 gnd 0.144919f
C5615 a_n8300_8799.t6 gnd 0.144919f
C5616 a_n8300_8799.n10 gnd 1.143f
C5617 a_n8300_8799.t9 gnd 0.144919f
C5618 a_n8300_8799.t11 gnd 0.144919f
C5619 a_n8300_8799.n11 gnd 1.14111f
C5620 a_n8300_8799.n12 gnd 1.02572f
C5621 a_n8300_8799.t1 gnd 0.144919f
C5622 a_n8300_8799.t13 gnd 0.144919f
C5623 a_n8300_8799.n13 gnd 1.14111f
C5624 a_n8300_8799.n14 gnd 0.505597f
C5625 a_n8300_8799.t38 gnd 0.144919f
C5626 a_n8300_8799.t3 gnd 0.144919f
C5627 a_n8300_8799.n15 gnd 1.14111f
C5628 a_n8300_8799.n16 gnd 2.02754f
C5629 a_n8300_8799.n17 gnd 6.373569f
C5630 a_n8300_8799.n18 gnd 0.052234f
C5631 a_n8300_8799.t92 gnd 0.600901f
C5632 a_n8300_8799.n19 gnd 0.268374f
C5633 a_n8300_8799.n20 gnd 0.052234f
C5634 a_n8300_8799.n21 gnd 0.011853f
C5635 a_n8300_8799.t40 gnd 0.600901f
C5636 a_n8300_8799.n22 gnd 0.052234f
C5637 a_n8300_8799.t71 gnd 0.600901f
C5638 a_n8300_8799.n23 gnd 0.265315f
C5639 a_n8300_8799.t72 gnd 0.600901f
C5640 a_n8300_8799.n24 gnd 0.052234f
C5641 a_n8300_8799.t86 gnd 0.600901f
C5642 a_n8300_8799.n25 gnd 0.265637f
C5643 a_n8300_8799.n26 gnd 0.052234f
C5644 a_n8300_8799.n27 gnd 0.011853f
C5645 a_n8300_8799.t138 gnd 0.600901f
C5646 a_n8300_8799.n28 gnd 0.052234f
C5647 a_n8300_8799.t141 gnd 0.600901f
C5648 a_n8300_8799.n29 gnd 0.268374f
C5649 a_n8300_8799.n30 gnd 0.052234f
C5650 a_n8300_8799.n31 gnd 0.011853f
C5651 a_n8300_8799.t102 gnd 0.600901f
C5652 a_n8300_8799.n32 gnd 0.16502f
C5653 a_n8300_8799.t146 gnd 0.600901f
C5654 a_n8300_8799.t107 gnd 0.612274f
C5655 a_n8300_8799.n33 gnd 0.251902f
C5656 a_n8300_8799.n34 gnd 0.264671f
C5657 a_n8300_8799.n35 gnd 0.011853f
C5658 a_n8300_8799.t69 gnd 0.600901f
C5659 a_n8300_8799.n36 gnd 0.268374f
C5660 a_n8300_8799.n37 gnd 0.052234f
C5661 a_n8300_8799.n38 gnd 0.052234f
C5662 a_n8300_8799.n39 gnd 0.052234f
C5663 a_n8300_8799.n40 gnd 0.266281f
C5664 a_n8300_8799.t139 gnd 0.600901f
C5665 a_n8300_8799.n41 gnd 0.264993f
C5666 a_n8300_8799.n42 gnd 0.011853f
C5667 a_n8300_8799.n43 gnd 0.052234f
C5668 a_n8300_8799.n44 gnd 0.052234f
C5669 a_n8300_8799.n45 gnd 0.052234f
C5670 a_n8300_8799.n46 gnd 0.011853f
C5671 a_n8300_8799.t87 gnd 0.600901f
C5672 a_n8300_8799.n47 gnd 0.265959f
C5673 a_n8300_8799.t118 gnd 0.600901f
C5674 a_n8300_8799.n48 gnd 0.265315f
C5675 a_n8300_8799.n49 gnd 0.052234f
C5676 a_n8300_8799.n50 gnd 0.052234f
C5677 a_n8300_8799.n51 gnd 0.052234f
C5678 a_n8300_8799.n52 gnd 0.268374f
C5679 a_n8300_8799.n53 gnd 0.011853f
C5680 a_n8300_8799.t85 gnd 0.600901f
C5681 a_n8300_8799.n54 gnd 0.265637f
C5682 a_n8300_8799.n55 gnd 0.052234f
C5683 a_n8300_8799.n56 gnd 0.052234f
C5684 a_n8300_8799.n57 gnd 0.052234f
C5685 a_n8300_8799.n58 gnd 0.011853f
C5686 a_n8300_8799.t115 gnd 0.600901f
C5687 a_n8300_8799.n59 gnd 0.268374f
C5688 a_n8300_8799.n60 gnd 0.011853f
C5689 a_n8300_8799.n61 gnd 0.052234f
C5690 a_n8300_8799.n62 gnd 0.052234f
C5691 a_n8300_8799.n63 gnd 0.052234f
C5692 a_n8300_8799.n64 gnd 0.265959f
C5693 a_n8300_8799.n65 gnd 0.011853f
C5694 a_n8300_8799.t112 gnd 0.600901f
C5695 a_n8300_8799.n66 gnd 0.268374f
C5696 a_n8300_8799.n67 gnd 0.052234f
C5697 a_n8300_8799.n68 gnd 0.052234f
C5698 a_n8300_8799.n69 gnd 0.052234f
C5699 a_n8300_8799.n70 gnd 0.264993f
C5700 a_n8300_8799.t70 gnd 0.600901f
C5701 a_n8300_8799.n71 gnd 0.266281f
C5702 a_n8300_8799.n72 gnd 0.011853f
C5703 a_n8300_8799.n73 gnd 0.052234f
C5704 a_n8300_8799.n74 gnd 0.052234f
C5705 a_n8300_8799.n75 gnd 0.052234f
C5706 a_n8300_8799.n76 gnd 0.011853f
C5707 a_n8300_8799.t140 gnd 0.600901f
C5708 a_n8300_8799.n77 gnd 0.264671f
C5709 a_n8300_8799.t51 gnd 0.600901f
C5710 a_n8300_8799.n78 gnd 0.262899f
C5711 a_n8300_8799.n79 gnd 0.29615f
C5712 a_n8300_8799.n80 gnd 0.052234f
C5713 a_n8300_8799.t104 gnd 0.600901f
C5714 a_n8300_8799.n81 gnd 0.268374f
C5715 a_n8300_8799.n82 gnd 0.052234f
C5716 a_n8300_8799.n83 gnd 0.011853f
C5717 a_n8300_8799.t50 gnd 0.600901f
C5718 a_n8300_8799.n84 gnd 0.052234f
C5719 a_n8300_8799.t83 gnd 0.600901f
C5720 a_n8300_8799.n85 gnd 0.265315f
C5721 a_n8300_8799.t84 gnd 0.600901f
C5722 a_n8300_8799.n86 gnd 0.052234f
C5723 a_n8300_8799.t94 gnd 0.600901f
C5724 a_n8300_8799.n87 gnd 0.265637f
C5725 a_n8300_8799.n88 gnd 0.052234f
C5726 a_n8300_8799.n89 gnd 0.011853f
C5727 a_n8300_8799.t152 gnd 0.600901f
C5728 a_n8300_8799.n90 gnd 0.052234f
C5729 a_n8300_8799.t157 gnd 0.600901f
C5730 a_n8300_8799.n91 gnd 0.268374f
C5731 a_n8300_8799.n92 gnd 0.052234f
C5732 a_n8300_8799.n93 gnd 0.011853f
C5733 a_n8300_8799.t116 gnd 0.600901f
C5734 a_n8300_8799.n94 gnd 0.16502f
C5735 a_n8300_8799.t159 gnd 0.600901f
C5736 a_n8300_8799.t123 gnd 0.612274f
C5737 a_n8300_8799.n95 gnd 0.251902f
C5738 a_n8300_8799.n96 gnd 0.264671f
C5739 a_n8300_8799.n97 gnd 0.011853f
C5740 a_n8300_8799.t79 gnd 0.600901f
C5741 a_n8300_8799.n98 gnd 0.268374f
C5742 a_n8300_8799.n99 gnd 0.052234f
C5743 a_n8300_8799.n100 gnd 0.052234f
C5744 a_n8300_8799.n101 gnd 0.052234f
C5745 a_n8300_8799.n102 gnd 0.266281f
C5746 a_n8300_8799.t154 gnd 0.600901f
C5747 a_n8300_8799.n103 gnd 0.264993f
C5748 a_n8300_8799.n104 gnd 0.011853f
C5749 a_n8300_8799.n105 gnd 0.052234f
C5750 a_n8300_8799.n106 gnd 0.052234f
C5751 a_n8300_8799.n107 gnd 0.052234f
C5752 a_n8300_8799.n108 gnd 0.011853f
C5753 a_n8300_8799.t97 gnd 0.600901f
C5754 a_n8300_8799.n109 gnd 0.265959f
C5755 a_n8300_8799.t135 gnd 0.600901f
C5756 a_n8300_8799.n110 gnd 0.265315f
C5757 a_n8300_8799.n111 gnd 0.052234f
C5758 a_n8300_8799.n112 gnd 0.052234f
C5759 a_n8300_8799.n113 gnd 0.052234f
C5760 a_n8300_8799.n114 gnd 0.268374f
C5761 a_n8300_8799.n115 gnd 0.011853f
C5762 a_n8300_8799.t93 gnd 0.600901f
C5763 a_n8300_8799.n116 gnd 0.265637f
C5764 a_n8300_8799.n117 gnd 0.052234f
C5765 a_n8300_8799.n118 gnd 0.052234f
C5766 a_n8300_8799.n119 gnd 0.052234f
C5767 a_n8300_8799.n120 gnd 0.011853f
C5768 a_n8300_8799.t133 gnd 0.600901f
C5769 a_n8300_8799.n121 gnd 0.268374f
C5770 a_n8300_8799.n122 gnd 0.011853f
C5771 a_n8300_8799.n123 gnd 0.052234f
C5772 a_n8300_8799.n124 gnd 0.052234f
C5773 a_n8300_8799.n125 gnd 0.052234f
C5774 a_n8300_8799.n126 gnd 0.265959f
C5775 a_n8300_8799.n127 gnd 0.011853f
C5776 a_n8300_8799.t129 gnd 0.600901f
C5777 a_n8300_8799.n128 gnd 0.268374f
C5778 a_n8300_8799.n129 gnd 0.052234f
C5779 a_n8300_8799.n130 gnd 0.052234f
C5780 a_n8300_8799.n131 gnd 0.052234f
C5781 a_n8300_8799.n132 gnd 0.264993f
C5782 a_n8300_8799.t80 gnd 0.600901f
C5783 a_n8300_8799.n133 gnd 0.266281f
C5784 a_n8300_8799.n134 gnd 0.011853f
C5785 a_n8300_8799.n135 gnd 0.052234f
C5786 a_n8300_8799.n136 gnd 0.052234f
C5787 a_n8300_8799.n137 gnd 0.052234f
C5788 a_n8300_8799.n138 gnd 0.011853f
C5789 a_n8300_8799.t155 gnd 0.600901f
C5790 a_n8300_8799.n139 gnd 0.264671f
C5791 a_n8300_8799.t63 gnd 0.600901f
C5792 a_n8300_8799.n140 gnd 0.262899f
C5793 a_n8300_8799.n141 gnd 0.130193f
C5794 a_n8300_8799.n142 gnd 0.903372f
C5795 a_n8300_8799.n143 gnd 0.052234f
C5796 a_n8300_8799.t108 gnd 0.600901f
C5797 a_n8300_8799.n144 gnd 0.268374f
C5798 a_n8300_8799.n145 gnd 0.052234f
C5799 a_n8300_8799.n146 gnd 0.011853f
C5800 a_n8300_8799.t91 gnd 0.600901f
C5801 a_n8300_8799.n147 gnd 0.052234f
C5802 a_n8300_8799.t145 gnd 0.600901f
C5803 a_n8300_8799.n148 gnd 0.265315f
C5804 a_n8300_8799.t117 gnd 0.600901f
C5805 a_n8300_8799.n149 gnd 0.052234f
C5806 a_n8300_8799.t41 gnd 0.600901f
C5807 a_n8300_8799.n150 gnd 0.265637f
C5808 a_n8300_8799.n151 gnd 0.052234f
C5809 a_n8300_8799.n152 gnd 0.011853f
C5810 a_n8300_8799.t142 gnd 0.600901f
C5811 a_n8300_8799.n153 gnd 0.052234f
C5812 a_n8300_8799.t90 gnd 0.600901f
C5813 a_n8300_8799.n154 gnd 0.268374f
C5814 a_n8300_8799.n155 gnd 0.052234f
C5815 a_n8300_8799.n156 gnd 0.011853f
C5816 a_n8300_8799.t52 gnd 0.600901f
C5817 a_n8300_8799.n157 gnd 0.16502f
C5818 a_n8300_8799.t74 gnd 0.600901f
C5819 a_n8300_8799.t125 gnd 0.612274f
C5820 a_n8300_8799.n158 gnd 0.251902f
C5821 a_n8300_8799.n159 gnd 0.264671f
C5822 a_n8300_8799.n160 gnd 0.011853f
C5823 a_n8300_8799.t95 gnd 0.600901f
C5824 a_n8300_8799.n161 gnd 0.268374f
C5825 a_n8300_8799.n162 gnd 0.052234f
C5826 a_n8300_8799.n163 gnd 0.052234f
C5827 a_n8300_8799.n164 gnd 0.052234f
C5828 a_n8300_8799.n165 gnd 0.266281f
C5829 a_n8300_8799.t113 gnd 0.600901f
C5830 a_n8300_8799.n166 gnd 0.264993f
C5831 a_n8300_8799.n167 gnd 0.011853f
C5832 a_n8300_8799.n168 gnd 0.052234f
C5833 a_n8300_8799.n169 gnd 0.052234f
C5834 a_n8300_8799.n170 gnd 0.052234f
C5835 a_n8300_8799.n171 gnd 0.011853f
C5836 a_n8300_8799.t134 gnd 0.600901f
C5837 a_n8300_8799.n172 gnd 0.265959f
C5838 a_n8300_8799.t81 gnd 0.600901f
C5839 a_n8300_8799.n173 gnd 0.265315f
C5840 a_n8300_8799.n174 gnd 0.052234f
C5841 a_n8300_8799.n175 gnd 0.052234f
C5842 a_n8300_8799.n176 gnd 0.052234f
C5843 a_n8300_8799.n177 gnd 0.268374f
C5844 a_n8300_8799.n178 gnd 0.011853f
C5845 a_n8300_8799.t57 gnd 0.600901f
C5846 a_n8300_8799.n179 gnd 0.265637f
C5847 a_n8300_8799.n180 gnd 0.052234f
C5848 a_n8300_8799.n181 gnd 0.052234f
C5849 a_n8300_8799.n182 gnd 0.052234f
C5850 a_n8300_8799.n183 gnd 0.011853f
C5851 a_n8300_8799.t98 gnd 0.600901f
C5852 a_n8300_8799.n184 gnd 0.268374f
C5853 a_n8300_8799.n185 gnd 0.011853f
C5854 a_n8300_8799.n186 gnd 0.052234f
C5855 a_n8300_8799.n187 gnd 0.052234f
C5856 a_n8300_8799.n188 gnd 0.052234f
C5857 a_n8300_8799.n189 gnd 0.265959f
C5858 a_n8300_8799.n190 gnd 0.011853f
C5859 a_n8300_8799.t151 gnd 0.600901f
C5860 a_n8300_8799.n191 gnd 0.268374f
C5861 a_n8300_8799.n192 gnd 0.052234f
C5862 a_n8300_8799.n193 gnd 0.052234f
C5863 a_n8300_8799.n194 gnd 0.052234f
C5864 a_n8300_8799.n195 gnd 0.264993f
C5865 a_n8300_8799.t46 gnd 0.600901f
C5866 a_n8300_8799.n196 gnd 0.266281f
C5867 a_n8300_8799.n197 gnd 0.011853f
C5868 a_n8300_8799.n198 gnd 0.052234f
C5869 a_n8300_8799.n199 gnd 0.052234f
C5870 a_n8300_8799.n200 gnd 0.052234f
C5871 a_n8300_8799.n201 gnd 0.011853f
C5872 a_n8300_8799.t61 gnd 0.600901f
C5873 a_n8300_8799.n202 gnd 0.264671f
C5874 a_n8300_8799.t130 gnd 0.600901f
C5875 a_n8300_8799.n203 gnd 0.262899f
C5876 a_n8300_8799.n204 gnd 0.130193f
C5877 a_n8300_8799.n205 gnd 1.62818f
C5878 a_n8300_8799.n206 gnd 0.052234f
C5879 a_n8300_8799.t89 gnd 0.600901f
C5880 a_n8300_8799.t65 gnd 0.600901f
C5881 a_n8300_8799.t144 gnd 0.600901f
C5882 a_n8300_8799.n207 gnd 0.268374f
C5883 a_n8300_8799.n208 gnd 0.052234f
C5884 a_n8300_8799.t106 gnd 0.600901f
C5885 a_n8300_8799.t103 gnd 0.600901f
C5886 a_n8300_8799.n209 gnd 0.052234f
C5887 a_n8300_8799.t43 gnd 0.600901f
C5888 a_n8300_8799.n210 gnd 0.268374f
C5889 a_n8300_8799.n211 gnd 0.052234f
C5890 a_n8300_8799.t111 gnd 0.600901f
C5891 a_n8300_8799.t110 gnd 0.600901f
C5892 a_n8300_8799.n212 gnd 0.052234f
C5893 a_n8300_8799.t45 gnd 0.600901f
C5894 a_n8300_8799.n213 gnd 0.268374f
C5895 a_n8300_8799.n214 gnd 0.052234f
C5896 a_n8300_8799.t44 gnd 0.600901f
C5897 a_n8300_8799.t132 gnd 0.600901f
C5898 a_n8300_8799.n215 gnd 0.052234f
C5899 a_n8300_8799.t60 gnd 0.600901f
C5900 a_n8300_8799.n216 gnd 0.268374f
C5901 a_n8300_8799.n217 gnd 0.052234f
C5902 a_n8300_8799.t49 gnd 0.600901f
C5903 a_n8300_8799.t136 gnd 0.600901f
C5904 a_n8300_8799.n218 gnd 0.052234f
C5905 a_n8300_8799.t88 gnd 0.600901f
C5906 a_n8300_8799.n219 gnd 0.268374f
C5907 a_n8300_8799.n220 gnd 0.052234f
C5908 a_n8300_8799.t64 gnd 0.600901f
C5909 a_n8300_8799.t156 gnd 0.600901f
C5910 a_n8300_8799.n221 gnd 0.052234f
C5911 a_n8300_8799.t105 gnd 0.600901f
C5912 a_n8300_8799.n222 gnd 0.268374f
C5913 a_n8300_8799.t149 gnd 0.612274f
C5914 a_n8300_8799.n223 gnd 0.251902f
C5915 a_n8300_8799.t67 gnd 0.600901f
C5916 a_n8300_8799.n224 gnd 0.264671f
C5917 a_n8300_8799.n225 gnd 0.011853f
C5918 a_n8300_8799.n226 gnd 0.16502f
C5919 a_n8300_8799.n227 gnd 0.052234f
C5920 a_n8300_8799.n228 gnd 0.052234f
C5921 a_n8300_8799.n229 gnd 0.011853f
C5922 a_n8300_8799.n230 gnd 0.266281f
C5923 a_n8300_8799.n231 gnd 0.264993f
C5924 a_n8300_8799.n232 gnd 0.011853f
C5925 a_n8300_8799.n233 gnd 0.052234f
C5926 a_n8300_8799.n234 gnd 0.052234f
C5927 a_n8300_8799.n235 gnd 0.052234f
C5928 a_n8300_8799.n236 gnd 0.011853f
C5929 a_n8300_8799.n237 gnd 0.265959f
C5930 a_n8300_8799.n238 gnd 0.265315f
C5931 a_n8300_8799.n239 gnd 0.011853f
C5932 a_n8300_8799.n240 gnd 0.052234f
C5933 a_n8300_8799.n241 gnd 0.052234f
C5934 a_n8300_8799.n242 gnd 0.052234f
C5935 a_n8300_8799.n243 gnd 0.011853f
C5936 a_n8300_8799.n244 gnd 0.265637f
C5937 a_n8300_8799.n245 gnd 0.265637f
C5938 a_n8300_8799.n246 gnd 0.011853f
C5939 a_n8300_8799.n247 gnd 0.052234f
C5940 a_n8300_8799.n248 gnd 0.052234f
C5941 a_n8300_8799.n249 gnd 0.052234f
C5942 a_n8300_8799.n250 gnd 0.011853f
C5943 a_n8300_8799.n251 gnd 0.265315f
C5944 a_n8300_8799.n252 gnd 0.265959f
C5945 a_n8300_8799.n253 gnd 0.011853f
C5946 a_n8300_8799.n254 gnd 0.052234f
C5947 a_n8300_8799.n255 gnd 0.052234f
C5948 a_n8300_8799.n256 gnd 0.052234f
C5949 a_n8300_8799.n257 gnd 0.011853f
C5950 a_n8300_8799.n258 gnd 0.264993f
C5951 a_n8300_8799.n259 gnd 0.266281f
C5952 a_n8300_8799.n260 gnd 0.011853f
C5953 a_n8300_8799.n261 gnd 0.052234f
C5954 a_n8300_8799.n262 gnd 0.052234f
C5955 a_n8300_8799.n263 gnd 0.052234f
C5956 a_n8300_8799.n264 gnd 0.011853f
C5957 a_n8300_8799.n265 gnd 0.264671f
C5958 a_n8300_8799.n266 gnd 0.262899f
C5959 a_n8300_8799.n267 gnd 0.29615f
C5960 a_n8300_8799.n268 gnd 0.052234f
C5961 a_n8300_8799.t100 gnd 0.600901f
C5962 a_n8300_8799.t76 gnd 0.600901f
C5963 a_n8300_8799.t158 gnd 0.600901f
C5964 a_n8300_8799.n269 gnd 0.268374f
C5965 a_n8300_8799.n270 gnd 0.052234f
C5966 a_n8300_8799.t121 gnd 0.600901f
C5967 a_n8300_8799.t120 gnd 0.600901f
C5968 a_n8300_8799.n271 gnd 0.052234f
C5969 a_n8300_8799.t54 gnd 0.600901f
C5970 a_n8300_8799.n272 gnd 0.268374f
C5971 a_n8300_8799.n273 gnd 0.052234f
C5972 a_n8300_8799.t128 gnd 0.600901f
C5973 a_n8300_8799.t127 gnd 0.600901f
C5974 a_n8300_8799.n274 gnd 0.052234f
C5975 a_n8300_8799.t56 gnd 0.600901f
C5976 a_n8300_8799.n275 gnd 0.268374f
C5977 a_n8300_8799.n276 gnd 0.052234f
C5978 a_n8300_8799.t55 gnd 0.600901f
C5979 a_n8300_8799.t148 gnd 0.600901f
C5980 a_n8300_8799.n277 gnd 0.052234f
C5981 a_n8300_8799.t73 gnd 0.600901f
C5982 a_n8300_8799.n278 gnd 0.268374f
C5983 a_n8300_8799.n279 gnd 0.052234f
C5984 a_n8300_8799.t59 gnd 0.600901f
C5985 a_n8300_8799.t150 gnd 0.600901f
C5986 a_n8300_8799.n280 gnd 0.052234f
C5987 a_n8300_8799.t101 gnd 0.600901f
C5988 a_n8300_8799.n281 gnd 0.268374f
C5989 a_n8300_8799.n282 gnd 0.052234f
C5990 a_n8300_8799.t77 gnd 0.600901f
C5991 a_n8300_8799.t47 gnd 0.600901f
C5992 a_n8300_8799.n283 gnd 0.052234f
C5993 a_n8300_8799.t122 gnd 0.600901f
C5994 a_n8300_8799.n284 gnd 0.268374f
C5995 a_n8300_8799.t42 gnd 0.612274f
C5996 a_n8300_8799.n285 gnd 0.251902f
C5997 a_n8300_8799.t78 gnd 0.600901f
C5998 a_n8300_8799.n286 gnd 0.264671f
C5999 a_n8300_8799.n287 gnd 0.011853f
C6000 a_n8300_8799.n288 gnd 0.16502f
C6001 a_n8300_8799.n289 gnd 0.052234f
C6002 a_n8300_8799.n290 gnd 0.052234f
C6003 a_n8300_8799.n291 gnd 0.011853f
C6004 a_n8300_8799.n292 gnd 0.266281f
C6005 a_n8300_8799.n293 gnd 0.264993f
C6006 a_n8300_8799.n294 gnd 0.011853f
C6007 a_n8300_8799.n295 gnd 0.052234f
C6008 a_n8300_8799.n296 gnd 0.052234f
C6009 a_n8300_8799.n297 gnd 0.052234f
C6010 a_n8300_8799.n298 gnd 0.011853f
C6011 a_n8300_8799.n299 gnd 0.265959f
C6012 a_n8300_8799.n300 gnd 0.265315f
C6013 a_n8300_8799.n301 gnd 0.011853f
C6014 a_n8300_8799.n302 gnd 0.052234f
C6015 a_n8300_8799.n303 gnd 0.052234f
C6016 a_n8300_8799.n304 gnd 0.052234f
C6017 a_n8300_8799.n305 gnd 0.011853f
C6018 a_n8300_8799.n306 gnd 0.265637f
C6019 a_n8300_8799.n307 gnd 0.265637f
C6020 a_n8300_8799.n308 gnd 0.011853f
C6021 a_n8300_8799.n309 gnd 0.052234f
C6022 a_n8300_8799.n310 gnd 0.052234f
C6023 a_n8300_8799.n311 gnd 0.052234f
C6024 a_n8300_8799.n312 gnd 0.011853f
C6025 a_n8300_8799.n313 gnd 0.265315f
C6026 a_n8300_8799.n314 gnd 0.265959f
C6027 a_n8300_8799.n315 gnd 0.011853f
C6028 a_n8300_8799.n316 gnd 0.052234f
C6029 a_n8300_8799.n317 gnd 0.052234f
C6030 a_n8300_8799.n318 gnd 0.052234f
C6031 a_n8300_8799.n319 gnd 0.011853f
C6032 a_n8300_8799.n320 gnd 0.264993f
C6033 a_n8300_8799.n321 gnd 0.266281f
C6034 a_n8300_8799.n322 gnd 0.011853f
C6035 a_n8300_8799.n323 gnd 0.052234f
C6036 a_n8300_8799.n324 gnd 0.052234f
C6037 a_n8300_8799.n325 gnd 0.052234f
C6038 a_n8300_8799.n326 gnd 0.011853f
C6039 a_n8300_8799.n327 gnd 0.264671f
C6040 a_n8300_8799.n328 gnd 0.262899f
C6041 a_n8300_8799.n329 gnd 0.130193f
C6042 a_n8300_8799.n330 gnd 0.903372f
C6043 a_n8300_8799.n331 gnd 0.052234f
C6044 a_n8300_8799.t131 gnd 0.600901f
C6045 a_n8300_8799.t62 gnd 0.600901f
C6046 a_n8300_8799.t109 gnd 0.600901f
C6047 a_n8300_8799.n332 gnd 0.268374f
C6048 a_n8300_8799.n333 gnd 0.052234f
C6049 a_n8300_8799.t48 gnd 0.600901f
C6050 a_n8300_8799.t68 gnd 0.600901f
C6051 a_n8300_8799.n334 gnd 0.052234f
C6052 a_n8300_8799.t153 gnd 0.600901f
C6053 a_n8300_8799.n335 gnd 0.268374f
C6054 a_n8300_8799.n336 gnd 0.052234f
C6055 a_n8300_8799.t119 gnd 0.600901f
C6056 a_n8300_8799.t147 gnd 0.600901f
C6057 a_n8300_8799.n337 gnd 0.052234f
C6058 a_n8300_8799.t99 gnd 0.600901f
C6059 a_n8300_8799.n338 gnd 0.268374f
C6060 a_n8300_8799.n339 gnd 0.052234f
C6061 a_n8300_8799.t126 gnd 0.600901f
C6062 a_n8300_8799.t58 gnd 0.600901f
C6063 a_n8300_8799.n340 gnd 0.052234f
C6064 a_n8300_8799.t143 gnd 0.600901f
C6065 a_n8300_8799.n341 gnd 0.268374f
C6066 a_n8300_8799.n342 gnd 0.052234f
C6067 a_n8300_8799.t82 gnd 0.600901f
C6068 a_n8300_8799.t137 gnd 0.600901f
C6069 a_n8300_8799.n343 gnd 0.052234f
C6070 a_n8300_8799.t66 gnd 0.600901f
C6071 a_n8300_8799.n344 gnd 0.268374f
C6072 a_n8300_8799.n345 gnd 0.052234f
C6073 a_n8300_8799.t114 gnd 0.600901f
C6074 a_n8300_8799.t53 gnd 0.600901f
C6075 a_n8300_8799.n346 gnd 0.052234f
C6076 a_n8300_8799.t96 gnd 0.600901f
C6077 a_n8300_8799.n347 gnd 0.268374f
C6078 a_n8300_8799.t124 gnd 0.612274f
C6079 a_n8300_8799.n348 gnd 0.251902f
C6080 a_n8300_8799.t75 gnd 0.600901f
C6081 a_n8300_8799.n349 gnd 0.264671f
C6082 a_n8300_8799.n350 gnd 0.011853f
C6083 a_n8300_8799.n351 gnd 0.16502f
C6084 a_n8300_8799.n352 gnd 0.052234f
C6085 a_n8300_8799.n353 gnd 0.052234f
C6086 a_n8300_8799.n354 gnd 0.011853f
C6087 a_n8300_8799.n355 gnd 0.266281f
C6088 a_n8300_8799.n356 gnd 0.264993f
C6089 a_n8300_8799.n357 gnd 0.011853f
C6090 a_n8300_8799.n358 gnd 0.052234f
C6091 a_n8300_8799.n359 gnd 0.052234f
C6092 a_n8300_8799.n360 gnd 0.052234f
C6093 a_n8300_8799.n361 gnd 0.011853f
C6094 a_n8300_8799.n362 gnd 0.265959f
C6095 a_n8300_8799.n363 gnd 0.265315f
C6096 a_n8300_8799.n364 gnd 0.011853f
C6097 a_n8300_8799.n365 gnd 0.052234f
C6098 a_n8300_8799.n366 gnd 0.052234f
C6099 a_n8300_8799.n367 gnd 0.052234f
C6100 a_n8300_8799.n368 gnd 0.011853f
C6101 a_n8300_8799.n369 gnd 0.265637f
C6102 a_n8300_8799.n370 gnd 0.265637f
C6103 a_n8300_8799.n371 gnd 0.011853f
C6104 a_n8300_8799.n372 gnd 0.052234f
C6105 a_n8300_8799.n373 gnd 0.052234f
C6106 a_n8300_8799.n374 gnd 0.052234f
C6107 a_n8300_8799.n375 gnd 0.011853f
C6108 a_n8300_8799.n376 gnd 0.265315f
C6109 a_n8300_8799.n377 gnd 0.265959f
C6110 a_n8300_8799.n378 gnd 0.011853f
C6111 a_n8300_8799.n379 gnd 0.052234f
C6112 a_n8300_8799.n380 gnd 0.052234f
C6113 a_n8300_8799.n381 gnd 0.052234f
C6114 a_n8300_8799.n382 gnd 0.011853f
C6115 a_n8300_8799.n383 gnd 0.264993f
C6116 a_n8300_8799.n384 gnd 0.266281f
C6117 a_n8300_8799.n385 gnd 0.011853f
C6118 a_n8300_8799.n386 gnd 0.052234f
C6119 a_n8300_8799.n387 gnd 0.052234f
C6120 a_n8300_8799.n388 gnd 0.052234f
C6121 a_n8300_8799.n389 gnd 0.011853f
C6122 a_n8300_8799.n390 gnd 0.264671f
C6123 a_n8300_8799.n391 gnd 0.262899f
C6124 a_n8300_8799.n392 gnd 0.130193f
C6125 a_n8300_8799.n393 gnd 1.19295f
C6126 a_n8300_8799.n394 gnd 14.034901f
C6127 a_n8300_8799.n395 gnd 4.39773f
C6128 a_n8300_8799.t22 gnd 0.112715f
C6129 a_n8300_8799.t23 gnd 0.112715f
C6130 a_n8300_8799.n396 gnd 0.998202f
C6131 a_n8300_8799.t16 gnd 0.112715f
C6132 a_n8300_8799.t17 gnd 0.112715f
C6133 a_n8300_8799.n397 gnd 0.995987f
C6134 a_n8300_8799.n398 gnd 0.793349f
C6135 a_n8300_8799.t15 gnd 0.112715f
C6136 a_n8300_8799.t33 gnd 0.112715f
C6137 a_n8300_8799.n399 gnd 0.995987f
C6138 a_n8300_8799.n400 gnd 0.331276f
C6139 a_n8300_8799.n401 gnd 0.472955f
C6140 a_n8300_8799.t35 gnd 0.112715f
C6141 a_n8300_8799.t28 gnd 0.112715f
C6142 a_n8300_8799.n402 gnd 0.995987f
C6143 a_n8300_8799.n403 gnd 0.331276f
C6144 a_n8300_8799.t30 gnd 0.112715f
C6145 a_n8300_8799.t14 gnd 0.112715f
C6146 a_n8300_8799.n404 gnd 0.995987f
C6147 a_n8300_8799.n405 gnd 0.389575f
C6148 a_n8300_8799.t32 gnd 0.112715f
C6149 a_n8300_8799.t34 gnd 0.112715f
C6150 a_n8300_8799.n406 gnd 0.995987f
C6151 a_n8300_8799.n407 gnd 2.8681f
C6152 a_n8300_8799.t29 gnd 0.112715f
C6153 a_n8300_8799.t27 gnd 0.112715f
C6154 a_n8300_8799.n408 gnd 0.998201f
C6155 a_n8300_8799.t18 gnd 0.112715f
C6156 a_n8300_8799.t24 gnd 0.112715f
C6157 a_n8300_8799.n409 gnd 0.995986f
C6158 a_n8300_8799.n410 gnd 0.793351f
C6159 a_n8300_8799.t36 gnd 0.112715f
C6160 a_n8300_8799.t19 gnd 0.112715f
C6161 a_n8300_8799.n411 gnd 0.995986f
C6162 a_n8300_8799.n412 gnd 0.331277f
C6163 a_n8300_8799.n413 gnd 2.41392f
C6164 a_n8300_8799.n414 gnd 0.331279f
C6165 a_n8300_8799.n415 gnd 0.995984f
C6166 a_n8300_8799.t37 gnd 0.112715f
C6167 a_n3827_n3924.n0 gnd 1.99733f
C6168 a_n3827_n3924.n1 gnd 2.17486f
C6169 a_n3827_n3924.n2 gnd 1.44807f
C6170 a_n3827_n3924.n3 gnd 1.31657f
C6171 a_n3827_n3924.n4 gnd 1.81285f
C6172 a_n3827_n3924.n5 gnd 0.914318f
C6173 a_n3827_n3924.n6 gnd 3.90473f
C6174 a_n3827_n3924.n7 gnd 0.886511f
C6175 a_n3827_n3924.n8 gnd 1.77302f
C6176 a_n3827_n3924.n9 gnd 2.49022f
C6177 a_n3827_n3924.n10 gnd 0.954549f
C6178 a_n3827_n3924.n11 gnd 0.724032f
C6179 a_n3827_n3924.n12 gnd 1.2733f
C6180 a_n3827_n3924.t1 gnd 1.26048f
C6181 a_n3827_n3924.t50 gnd 1.25868f
C6182 a_n3827_n3924.t5 gnd 1.25868f
C6183 a_n3827_n3924.t51 gnd 1.25868f
C6184 a_n3827_n3924.t21 gnd 1.25868f
C6185 a_n3827_n3924.t7 gnd 1.25868f
C6186 a_n3827_n3924.t49 gnd 1.25868f
C6187 a_n3827_n3924.t18 gnd 1.25868f
C6188 a_n3827_n3924.t57 gnd 1.25868f
C6189 a_n3827_n3924.t17 gnd 1.26084f
C6190 a_n3827_n3924.t36 gnd 1.01304f
C6191 a_n3827_n3924.t38 gnd 0.097472f
C6192 a_n3827_n3924.t33 gnd 0.097472f
C6193 a_n3827_n3924.n13 gnd 0.796068f
C6194 a_n3827_n3924.t26 gnd 0.097472f
C6195 a_n3827_n3924.t28 gnd 0.097472f
C6196 a_n3827_n3924.n14 gnd 0.796068f
C6197 a_n3827_n3924.t48 gnd 0.097472f
C6198 a_n3827_n3924.t42 gnd 0.097472f
C6199 a_n3827_n3924.n15 gnd 0.796068f
C6200 a_n3827_n3924.t44 gnd 0.097472f
C6201 a_n3827_n3924.t32 gnd 0.097472f
C6202 a_n3827_n3924.n16 gnd 0.796068f
C6203 a_n3827_n3924.t46 gnd 0.097472f
C6204 a_n3827_n3924.t31 gnd 0.097472f
C6205 a_n3827_n3924.n17 gnd 0.796068f
C6206 a_n3827_n3924.t29 gnd 1.01304f
C6207 a_n3827_n3924.t56 gnd 1.01304f
C6208 a_n3827_n3924.t15 gnd 0.097472f
C6209 a_n3827_n3924.t23 gnd 0.097472f
C6210 a_n3827_n3924.n18 gnd 0.796068f
C6211 a_n3827_n3924.t6 gnd 0.097472f
C6212 a_n3827_n3924.t12 gnd 0.097472f
C6213 a_n3827_n3924.n19 gnd 0.796068f
C6214 a_n3827_n3924.t20 gnd 0.097472f
C6215 a_n3827_n3924.t3 gnd 0.097472f
C6216 a_n3827_n3924.n20 gnd 0.796068f
C6217 a_n3827_n3924.t54 gnd 0.097472f
C6218 a_n3827_n3924.t53 gnd 0.097472f
C6219 a_n3827_n3924.n21 gnd 0.796068f
C6220 a_n3827_n3924.t16 gnd 0.097472f
C6221 a_n3827_n3924.t19 gnd 0.097472f
C6222 a_n3827_n3924.n22 gnd 0.796068f
C6223 a_n3827_n3924.t11 gnd 1.01304f
C6224 a_n3827_n3924.n23 gnd 0.914318f
C6225 a_n3827_n3924.t43 gnd 1.01304f
C6226 a_n3827_n3924.t35 gnd 0.097472f
C6227 a_n3827_n3924.t47 gnd 0.097472f
C6228 a_n3827_n3924.n24 gnd 0.796069f
C6229 a_n3827_n3924.t34 gnd 0.097472f
C6230 a_n3827_n3924.t25 gnd 0.097472f
C6231 a_n3827_n3924.n25 gnd 0.796069f
C6232 a_n3827_n3924.t45 gnd 0.097472f
C6233 a_n3827_n3924.t27 gnd 0.097472f
C6234 a_n3827_n3924.n26 gnd 0.796069f
C6235 a_n3827_n3924.t39 gnd 0.097472f
C6236 a_n3827_n3924.t41 gnd 0.097472f
C6237 a_n3827_n3924.n27 gnd 0.796069f
C6238 a_n3827_n3924.t37 gnd 0.097472f
C6239 a_n3827_n3924.t30 gnd 0.097472f
C6240 a_n3827_n3924.n28 gnd 0.796069f
C6241 a_n3827_n3924.t40 gnd 1.01304f
C6242 a_n3827_n3924.t2 gnd 1.01304f
C6243 a_n3827_n3924.t52 gnd 0.097472f
C6244 a_n3827_n3924.t55 gnd 0.097472f
C6245 a_n3827_n3924.n29 gnd 0.796069f
C6246 a_n3827_n3924.t8 gnd 0.097472f
C6247 a_n3827_n3924.t14 gnd 0.097472f
C6248 a_n3827_n3924.n30 gnd 0.796069f
C6249 a_n3827_n3924.t13 gnd 0.097472f
C6250 a_n3827_n3924.t24 gnd 0.097472f
C6251 a_n3827_n3924.n31 gnd 0.796069f
C6252 a_n3827_n3924.t22 gnd 0.097472f
C6253 a_n3827_n3924.t10 gnd 0.097472f
C6254 a_n3827_n3924.n32 gnd 0.796069f
C6255 a_n3827_n3924.t9 gnd 0.097472f
C6256 a_n3827_n3924.t4 gnd 0.097472f
C6257 a_n3827_n3924.n33 gnd 0.796069f
C6258 a_n3827_n3924.t0 gnd 1.01304f
C6259 plus.n0 gnd 0.0234f
C6260 plus.t21 gnd 0.330972f
C6261 plus.n1 gnd 0.0234f
C6262 plus.t22 gnd 0.330972f
C6263 plus.t16 gnd 0.330972f
C6264 plus.n2 gnd 0.147028f
C6265 plus.n3 gnd 0.0234f
C6266 plus.t17 gnd 0.330972f
C6267 plus.t11 gnd 0.330972f
C6268 plus.n4 gnd 0.147028f
C6269 plus.n5 gnd 0.0234f
C6270 plus.t5 gnd 0.330972f
C6271 plus.t6 gnd 0.330972f
C6272 plus.n6 gnd 0.147028f
C6273 plus.n7 gnd 0.0234f
C6274 plus.t23 gnd 0.330972f
C6275 plus.t24 gnd 0.330972f
C6276 plus.n8 gnd 0.147028f
C6277 plus.n9 gnd 0.0234f
C6278 plus.t18 gnd 0.330972f
C6279 plus.t13 gnd 0.330972f
C6280 plus.n10 gnd 0.151817f
C6281 plus.t15 gnd 0.342986f
C6282 plus.n11 gnd 0.13626f
C6283 plus.n12 gnd 0.100739f
C6284 plus.n13 gnd 0.00531f
C6285 plus.n14 gnd 0.147028f
C6286 plus.n15 gnd 0.00531f
C6287 plus.n16 gnd 0.0234f
C6288 plus.n17 gnd 0.0234f
C6289 plus.n18 gnd 0.0234f
C6290 plus.n19 gnd 0.00531f
C6291 plus.n20 gnd 0.147028f
C6292 plus.n21 gnd 0.00531f
C6293 plus.n22 gnd 0.0234f
C6294 plus.n23 gnd 0.0234f
C6295 plus.n24 gnd 0.0234f
C6296 plus.n25 gnd 0.00531f
C6297 plus.n26 gnd 0.147028f
C6298 plus.n27 gnd 0.00531f
C6299 plus.n28 gnd 0.0234f
C6300 plus.n29 gnd 0.0234f
C6301 plus.n30 gnd 0.0234f
C6302 plus.n31 gnd 0.00531f
C6303 plus.n32 gnd 0.147028f
C6304 plus.n33 gnd 0.00531f
C6305 plus.n34 gnd 0.0234f
C6306 plus.n35 gnd 0.0234f
C6307 plus.n36 gnd 0.0234f
C6308 plus.n37 gnd 0.00531f
C6309 plus.n38 gnd 0.147028f
C6310 plus.n39 gnd 0.00531f
C6311 plus.n40 gnd 0.147245f
C6312 plus.n41 gnd 0.264969f
C6313 plus.n42 gnd 0.0234f
C6314 plus.n43 gnd 0.00531f
C6315 plus.t10 gnd 0.330972f
C6316 plus.n44 gnd 0.0234f
C6317 plus.n45 gnd 0.00531f
C6318 plus.t12 gnd 0.330972f
C6319 plus.n46 gnd 0.0234f
C6320 plus.n47 gnd 0.00531f
C6321 plus.t7 gnd 0.330972f
C6322 plus.n48 gnd 0.0234f
C6323 plus.n49 gnd 0.00531f
C6324 plus.t27 gnd 0.330972f
C6325 plus.n50 gnd 0.0234f
C6326 plus.n51 gnd 0.00531f
C6327 plus.t26 gnd 0.330972f
C6328 plus.t20 gnd 0.342986f
C6329 plus.t19 gnd 0.330972f
C6330 plus.n52 gnd 0.151817f
C6331 plus.n53 gnd 0.13626f
C6332 plus.n54 gnd 0.100739f
C6333 plus.n55 gnd 0.0234f
C6334 plus.n56 gnd 0.147028f
C6335 plus.n57 gnd 0.00531f
C6336 plus.t25 gnd 0.330972f
C6337 plus.n58 gnd 0.147028f
C6338 plus.n59 gnd 0.0234f
C6339 plus.n60 gnd 0.0234f
C6340 plus.n61 gnd 0.0234f
C6341 plus.n62 gnd 0.147028f
C6342 plus.n63 gnd 0.00531f
C6343 plus.t9 gnd 0.330972f
C6344 plus.n64 gnd 0.147028f
C6345 plus.n65 gnd 0.0234f
C6346 plus.n66 gnd 0.0234f
C6347 plus.n67 gnd 0.0234f
C6348 plus.n68 gnd 0.147028f
C6349 plus.n69 gnd 0.00531f
C6350 plus.t14 gnd 0.330972f
C6351 plus.n70 gnd 0.147028f
C6352 plus.n71 gnd 0.0234f
C6353 plus.n72 gnd 0.0234f
C6354 plus.n73 gnd 0.0234f
C6355 plus.n74 gnd 0.147028f
C6356 plus.n75 gnd 0.00531f
C6357 plus.t28 gnd 0.330972f
C6358 plus.n76 gnd 0.147028f
C6359 plus.n77 gnd 0.0234f
C6360 plus.n78 gnd 0.0234f
C6361 plus.n79 gnd 0.0234f
C6362 plus.n80 gnd 0.147028f
C6363 plus.n81 gnd 0.00531f
C6364 plus.t8 gnd 0.330972f
C6365 plus.n82 gnd 0.147245f
C6366 plus.n83 gnd 0.774545f
C6367 plus.n84 gnd 1.15877f
C6368 plus.t1 gnd 0.040395f
C6369 plus.t2 gnd 0.007214f
C6370 plus.t3 gnd 0.007214f
C6371 plus.n85 gnd 0.023395f
C6372 plus.n86 gnd 0.181616f
C6373 plus.t0 gnd 0.007214f
C6374 plus.t4 gnd 0.007214f
C6375 plus.n87 gnd 0.023395f
C6376 plus.n88 gnd 0.136325f
C6377 plus.n89 gnd 2.94957f
.ends

