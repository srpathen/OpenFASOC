* NGSPICE file created from opamp72.ext - technology: sky130A

.subckt opamp72 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 a_n2472_13878.t27 a_n2650_13878.t28 a_n2650_13878.t29 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t101 a_n8300_8799.t40 vdd.t235 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878.t1 a_n2650_13878.t60 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t236 a_n8300_8799.t41 CSoutput.t100 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t153 gnd.t150 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X5 commonsourceibias.t47 commonsourceibias.t46 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X6 gnd.t221 commonsourceibias.t48 CSoutput.t118 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t149 gnd.t147 gnd.t148 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 a_n8300_8799.t39 plus.t5 a_n2903_n3924.t33 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 output.t19 outputibias.t8 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X10 output.t15 CSoutput.t144 vdd.t117 gnd.t37 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X11 CSoutput.t99 a_n8300_8799.t42 vdd.t209 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 CSoutput.t98 a_n8300_8799.t43 vdd.t211 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X13 gnd.t275 commonsourceibias.t49 CSoutput.t139 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 a_n2903_n3924.t32 plus.t6 a_n8300_8799.t33 gnd.t248 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X15 gnd.t4 commonsourceibias.t44 commonsourceibias.t45 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 a_n2650_8322.t25 a_n2650_13878.t61 a_n8300_8799.t23 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t235 commonsourceibias.t50 CSoutput.t120 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 outputibias.t7 outputibias.t6 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X19 output.t14 CSoutput.t145 vdd.t118 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t97 a_n8300_8799.t44 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t184 a_n8300_8799.t45 CSoutput.t96 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 a_n8300_8799.t20 a_n2650_13878.t62 a_n2650_8322.t24 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X23 a_n2650_13878.t41 minus.t5 a_n2903_n3924.t7 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n8300_8799.t35 plus.t7 a_n2903_n3924.t31 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 gnd.t234 commonsourceibias.t42 commonsourceibias.t43 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 vdd.t212 a_n8300_8799.t46 CSoutput.t95 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 a_n2650_13878.t42 minus.t6 a_n2903_n3924.t8 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 vdd.t214 a_n8300_8799.t47 CSoutput.t94 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 a_n8300_8799.t10 a_n2650_13878.t63 a_n2650_8322.t23 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X30 CSoutput.t110 commonsourceibias.t51 gnd.t187 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 CSoutput.t146 a_n2650_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 gnd.t185 commonsourceibias.t40 commonsourceibias.t41 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 CSoutput.t93 a_n8300_8799.t48 vdd.t249 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 a_n2903_n3924.t30 plus.t8 a_n8300_8799.t34 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X35 vdd.t23 CSoutput.t147 output.t13 gnd.t35 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X36 vdd.t24 CSoutput.t148 output.t12 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X37 CSoutput.t92 a_n8300_8799.t49 vdd.t250 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n2903_n3924.t46 minus.t7 a_n2650_13878.t59 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X39 CSoutput.t1 commonsourceibias.t52 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n2903_n3924.t3 diffpairibias.t16 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 vdd.t263 a_n8300_8799.t50 CSoutput.t91 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 CSoutput.t90 a_n8300_8799.t51 vdd.t264 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 CSoutput.t103 commonsourceibias.t53 gnd.t45 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 vdd.t100 vdd.t98 vdd.t99 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X45 a_n2472_13878.t26 a_n2650_13878.t10 a_n2650_13878.t11 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X46 a_n2650_13878.t35 a_n2650_13878.t34 a_n2472_13878.t25 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X47 CSoutput.t121 commonsourceibias.t54 gnd.t237 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X48 CSoutput.t89 a_n8300_8799.t52 vdd.t194 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 vdd.t97 vdd.t95 vdd.t96 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X50 vdd.t195 a_n8300_8799.t53 CSoutput.t88 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 plus.t4 gnd.t144 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X52 a_n2903_n3924.t29 plus.t9 a_n8300_8799.t8 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X53 gnd.t143 gnd.t141 gnd.t142 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X54 a_n2903_n3924.t28 plus.t10 a_n8300_8799.t3 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X55 diffpairibias.t15 diffpairibias.t14 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X56 a_n2650_13878.t27 a_n2650_13878.t26 a_n2472_13878.t24 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 gnd.t140 gnd.t138 gnd.t139 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X58 a_n8300_8799.t25 a_n2650_13878.t64 a_n2650_8322.t22 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X59 vdd.t247 a_n8300_8799.t54 CSoutput.t87 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 vdd.t248 a_n8300_8799.t55 CSoutput.t86 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 a_n2650_13878.t5 a_n2650_13878.t4 a_n2472_13878.t23 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X62 CSoutput.t85 a_n8300_8799.t56 vdd.t258 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 a_n8300_8799.t15 a_n2650_13878.t65 a_n2650_8322.t21 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X64 gnd.t17 commonsourceibias.t55 CSoutput.t0 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 gnd.t230 commonsourceibias.t56 CSoutput.t119 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 diffpairibias.t13 diffpairibias.t12 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X67 CSoutput.t84 a_n8300_8799.t57 vdd.t259 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 output.t11 CSoutput.t149 vdd.t228 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X69 gnd.t158 commonsourceibias.t57 CSoutput.t104 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 commonsourceibias.t39 commonsourceibias.t38 gnd.t184 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 vdd.t229 CSoutput.t150 output.t10 gnd.t32 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X72 a_n2650_8322.t20 a_n2650_13878.t66 a_n8300_8799.t22 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X73 vdd.t94 vdd.t92 vdd.t93 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X74 CSoutput.t83 a_n8300_8799.t58 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 a_n2903_n3924.t6 minus.t8 a_n2650_13878.t40 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X76 a_n2903_n3924.t27 plus.t11 a_n8300_8799.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X77 gnd.t137 gnd.t135 minus.t4 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X78 gnd.t284 commonsourceibias.t58 CSoutput.t140 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 a_n8300_8799.t38 plus.t12 a_n2903_n3924.t26 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X80 gnd.t134 gnd.t132 gnd.t133 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X81 commonsourceibias.t37 commonsourceibias.t36 gnd.t274 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 vdd.t126 a_n8300_8799.t59 CSoutput.t82 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 a_n2903_n3924.t4 diffpairibias.t17 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X84 gnd.t174 commonsourceibias.t34 commonsourceibias.t35 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 vdd.t196 a_n8300_8799.t60 CSoutput.t81 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t197 a_n8300_8799.t61 CSoutput.t80 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 vdd.t216 a_n8300_8799.t62 CSoutput.t79 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X88 a_n8300_8799.t9 a_n2650_13878.t67 a_n2650_8322.t19 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X89 a_n2650_13878.t9 a_n2650_13878.t8 a_n2472_13878.t22 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 a_n2903_n3924.t25 plus.t13 a_n8300_8799.t31 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X91 a_n2650_13878.t23 a_n2650_13878.t22 a_n2472_13878.t21 vdd.t133 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X92 gnd.t253 commonsourceibias.t32 commonsourceibias.t33 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X93 commonsourceibias.t31 commonsourceibias.t30 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 outputibias.t5 outputibias.t4 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X95 CSoutput.t78 a_n8300_8799.t63 vdd.t217 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 vdd.t243 a_n8300_8799.t64 CSoutput.t77 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 CSoutput.t126 commonsourceibias.t59 gnd.t245 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t230 CSoutput.t151 output.t9 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X99 CSoutput.t76 a_n8300_8799.t65 vdd.t244 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 vdd.t91 vdd.t89 vdd.t90 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X101 CSoutput.t111 commonsourceibias.t60 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 vdd.t88 vdd.t85 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X103 gnd.t162 commonsourceibias.t61 CSoutput.t106 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t131 gnd.t128 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X105 commonsourceibias.t29 commonsourceibias.t28 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t112 a_n8300_8799.t66 CSoutput.t75 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 CSoutput.t74 a_n8300_8799.t67 vdd.t113 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 CSoutput.t107 commonsourceibias.t62 gnd.t163 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X109 CSoutput.t152 a_n2650_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X110 outputibias.t3 outputibias.t2 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X111 vdd.t84 vdd.t82 vdd.t83 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X112 a_n2650_8322.t33 a_n2650_13878.t68 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X113 vdd.t174 a_n2650_13878.t69 a_n2650_8322.t32 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 vdd.t81 vdd.t79 vdd.t80 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X115 a_n2650_13878.t31 a_n2650_13878.t30 a_n2472_13878.t20 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 CSoutput.t73 a_n8300_8799.t68 vdd.t206 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 a_n2903_n3924.t5 diffpairibias.t18 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X118 commonsourceibias.t27 commonsourceibias.t26 gnd.t229 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 vdd.t172 a_n2650_13878.t70 a_n2472_13878.t0 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 vdd.t78 vdd.t75 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 vdd.t207 a_n8300_8799.t69 CSoutput.t72 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 vdd.t237 a_n8300_8799.t70 CSoutput.t71 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 plus.t3 gnd.t125 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X124 gnd.t9 commonsourceibias.t24 commonsourceibias.t25 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 gnd.t219 commonsourceibias.t63 CSoutput.t117 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 gnd.t124 gnd.t122 minus.t3 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X127 a_n8300_8799.t24 a_n2650_13878.t71 a_n2650_8322.t18 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n2650_8322.t31 a_n2650_13878.t72 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X129 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X130 gnd.t254 commonsourceibias.t64 CSoutput.t127 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n2650_13878.t45 minus.t9 a_n2903_n3924.t11 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X132 a_n8300_8799.t37 plus.t14 a_n2903_n3924.t24 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X133 gnd.t213 commonsourceibias.t65 CSoutput.t113 gnd.t212 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X134 vdd.t238 a_n8300_8799.t71 CSoutput.t70 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 vdd.t251 a_n8300_8799.t72 CSoutput.t69 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 a_n2650_13878.t19 a_n2650_13878.t18 a_n2472_13878.t19 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 CSoutput.t68 a_n8300_8799.t73 vdd.t252 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 a_n8300_8799.t4 plus.t15 a_n2903_n3924.t23 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X139 diffpairibias.t11 diffpairibias.t10 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X140 CSoutput.t67 a_n8300_8799.t74 vdd.t265 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 a_n8300_8799.t14 a_n2650_13878.t73 a_n2650_8322.t17 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 gnd.t165 commonsourceibias.t66 CSoutput.t108 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n2472_13878.t18 a_n2650_13878.t32 a_n2650_13878.t33 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 outputibias.t1 outputibias.t0 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X145 gnd.t238 commonsourceibias.t67 CSoutput.t122 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 CSoutput.t153 a_n2650_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X147 a_n2472_13878.t17 a_n2650_13878.t14 a_n2650_13878.t15 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 CSoutput.t66 a_n8300_8799.t75 vdd.t266 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X149 vdd.t165 a_n2650_13878.t74 a_n2650_8322.t30 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X150 gnd.t121 gnd.t119 minus.t2 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X151 CSoutput.t102 commonsourceibias.t68 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 CSoutput.t154 a_n2650_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X153 a_n2650_13878.t21 a_n2650_13878.t20 a_n2472_13878.t16 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 vdd.t1 a_n8300_8799.t76 CSoutput.t65 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 vdd.t70 vdd.t68 vdd.t69 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X156 a_n2903_n3924.t22 plus.t16 a_n8300_8799.t30 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X157 a_n2650_13878.t44 minus.t10 a_n2903_n3924.t10 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X158 vdd.t3 a_n8300_8799.t77 CSoutput.t64 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 gnd.t118 gnd.t115 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X160 a_n2903_n3924.t47 diffpairibias.t19 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X161 CSoutput.t125 commonsourceibias.t69 gnd.t244 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n8300_8799.t5 plus.t17 a_n2903_n3924.t21 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X163 CSoutput.t123 commonsourceibias.t70 gnd.t239 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 a_n2903_n3924.t0 diffpairibias.t20 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X165 vdd.t270 CSoutput.t155 output.t8 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 vdd.t198 a_n8300_8799.t78 CSoutput.t63 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 gnd.t214 commonsourceibias.t71 CSoutput.t114 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X168 CSoutput.t115 commonsourceibias.t72 gnd.t215 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2472_13878.t15 a_n2650_13878.t12 a_n2650_13878.t13 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X170 a_n8300_8799.t2 plus.t18 a_n2903_n3924.t20 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X171 vdd.t67 vdd.t65 vdd.t66 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X172 a_n2650_8322.t16 a_n2650_13878.t75 a_n8300_8799.t21 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 CSoutput.t62 a_n8300_8799.t79 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 CSoutput.t61 a_n8300_8799.t80 vdd.t239 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X175 a_n2472_13878.t3 a_n2650_13878.t76 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 gnd.t114 gnd.t112 gnd.t113 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X177 diffpairibias.t9 diffpairibias.t8 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X178 vdd.t160 a_n2650_13878.t77 a_n2472_13878.t2 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X179 a_n2650_13878.t47 minus.t11 a_n2903_n3924.t13 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X180 vdd.t240 a_n8300_8799.t81 CSoutput.t60 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 CSoutput.t59 a_n8300_8799.t82 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 a_n2903_n3924.t19 plus.t19 a_n8300_8799.t1 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X183 CSoutput.t58 a_n8300_8799.t83 vdd.t222 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 vdd.t13 a_n8300_8799.t84 CSoutput.t57 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 CSoutput.t128 commonsourceibias.t73 gnd.t255 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X186 gnd.t285 commonsourceibias.t74 CSoutput.t141 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 a_n2472_13878.t14 a_n2650_13878.t0 a_n2650_13878.t1 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X188 gnd.t197 commonsourceibias.t22 commonsourceibias.t23 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 gnd.t261 commonsourceibias.t75 CSoutput.t130 gnd.t212 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X190 vdd.t14 a_n8300_8799.t85 CSoutput.t56 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 a_n2650_8322.t15 a_n2650_13878.t78 a_n8300_8799.t28 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X192 gnd.t287 commonsourceibias.t76 CSoutput.t143 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 a_n2903_n3924.t9 minus.t12 a_n2650_13878.t43 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 a_n2472_13878.t13 a_n2650_13878.t38 a_n2650_13878.t39 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X195 vdd.t218 a_n8300_8799.t86 CSoutput.t55 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t54 a_n8300_8799.t87 vdd.t219 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 diffpairibias.t7 diffpairibias.t6 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X198 vdd.t64 vdd.t62 vdd.t63 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X199 vdd.t16 a_n8300_8799.t88 CSoutput.t53 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 vdd.t156 a_n2650_13878.t79 a_n2650_8322.t29 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X201 gnd.t273 commonsourceibias.t20 commonsourceibias.t21 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 CSoutput.t129 commonsourceibias.t77 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 gnd.t111 gnd.t108 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X204 a_n2903_n3924.t12 minus.t13 a_n2650_13878.t46 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X205 gnd.t107 gnd.t105 gnd.t106 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 gnd.t104 gnd.t102 gnd.t103 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X207 CSoutput.t52 a_n8300_8799.t89 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 minus.t1 gnd.t99 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X209 gnd.t98 gnd.t96 plus.t2 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X210 CSoutput.t142 commonsourceibias.t78 gnd.t286 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 a_n2903_n3924.t35 minus.t14 a_n2650_13878.t48 gnd.t248 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X212 a_n2472_13878.t6 a_n2650_13878.t80 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X213 vdd.t61 vdd.t59 vdd.t60 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X214 vdd.t58 vdd.t55 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X215 vdd.t267 a_n8300_8799.t90 CSoutput.t51 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X216 CSoutput.t50 a_n8300_8799.t91 vdd.t268 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t272 commonsourceibias.t18 commonsourceibias.t19 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t201 a_n8300_8799.t92 CSoutput.t49 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X219 gnd.t95 gnd.t92 gnd.t94 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X220 a_n2650_8322.t14 a_n2650_13878.t81 a_n8300_8799.t17 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X221 vdd.t151 a_n2650_13878.t82 a_n2650_8322.t28 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 CSoutput.t131 commonsourceibias.t79 gnd.t262 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 a_n2903_n3924.t2 diffpairibias.t21 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 output.t7 CSoutput.t156 vdd.t271 gnd.t29 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X225 CSoutput.t48 a_n8300_8799.t93 vdd.t202 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 vdd.t54 vdd.t51 vdd.t53 vdd.t52 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X227 a_n8300_8799.t32 plus.t20 a_n2903_n3924.t18 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X228 a_n2650_13878.t55 minus.t15 a_n2903_n3924.t42 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X229 CSoutput.t124 commonsourceibias.t80 gnd.t240 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 vdd.t253 a_n8300_8799.t94 CSoutput.t47 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 vdd.t254 a_n8300_8799.t95 CSoutput.t46 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 vdd.t50 vdd.t48 vdd.t49 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X233 a_n2903_n3924.t41 minus.t16 a_n2650_13878.t54 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X234 CSoutput.t157 a_n2650_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X235 CSoutput.t109 commonsourceibias.t81 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 gnd.t217 commonsourceibias.t82 CSoutput.t116 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 output.t18 outputibias.t9 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X238 output.t6 CSoutput.t158 vdd.t231 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X239 vdd.t47 vdd.t44 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X240 vdd.t260 a_n8300_8799.t96 CSoutput.t45 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 a_n2903_n3924.t40 minus.t17 a_n2650_13878.t53 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X242 gnd.t91 gnd.t89 gnd.t90 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X243 CSoutput.t44 a_n8300_8799.t97 vdd.t261 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 CSoutput.t43 a_n8300_8799.t98 vdd.t127 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 a_n2472_13878.t12 a_n2650_13878.t16 a_n2650_13878.t17 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 a_n2903_n3924.t39 minus.t18 a_n2650_13878.t52 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X247 vdd.t43 vdd.t41 vdd.t42 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 vdd.t40 vdd.t37 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X249 a_n2650_8322.t13 a_n2650_13878.t83 a_n8300_8799.t16 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 gnd.t88 gnd.t86 gnd.t87 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 output.t17 outputibias.t10 gnd.t178 gnd.t177 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X252 diffpairibias.t5 diffpairibias.t4 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X253 CSoutput.t42 a_n8300_8799.t99 vdd.t128 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 CSoutput.t41 a_n8300_8799.t100 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 CSoutput.t40 a_n8300_8799.t101 vdd.t187 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 vdd.t226 a_n8300_8799.t102 CSoutput.t39 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 gnd.t21 commonsourceibias.t83 CSoutput.t2 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t105 commonsourceibias.t84 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X259 vdd.t227 a_n8300_8799.t103 CSoutput.t38 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X260 CSoutput.t37 a_n8300_8799.t104 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 a_n2650_8322.t27 a_n2650_13878.t84 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X262 gnd.t85 gnd.t83 plus.t1 gnd.t84 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X263 gnd.t269 commonsourceibias.t85 CSoutput.t138 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 gnd.t236 commonsourceibias.t16 commonsourceibias.t17 gnd.t212 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X265 output.t5 CSoutput.t159 vdd.t232 gnd.t27 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X266 vdd.t22 a_n8300_8799.t105 CSoutput.t36 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X267 a_n2903_n3924.t38 minus.t19 a_n2650_13878.t51 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X268 gnd.t82 gnd.t79 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X269 vdd.t146 a_n2650_13878.t85 a_n2472_13878.t5 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X270 CSoutput.t35 a_n8300_8799.t106 vdd.t225 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X271 gnd.t72 gnd.t69 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X272 CSoutput.t34 a_n8300_8799.t107 vdd.t256 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t33 a_n8300_8799.t108 vdd.t269 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 vdd.t203 a_n8300_8799.t109 CSoutput.t32 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t224 a_n8300_8799.t110 CSoutput.t31 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t241 a_n8300_8799.t111 CSoutput.t30 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 gnd.t78 gnd.t76 gnd.t77 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X278 CSoutput.t137 commonsourceibias.t86 gnd.t268 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 CSoutput.t136 commonsourceibias.t87 gnd.t267 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t68 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X281 vdd.t233 CSoutput.t160 output.t4 gnd.t26 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 a_n8300_8799.t26 a_n2650_13878.t86 a_n2650_8322.t12 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X283 a_n2650_8322.t11 a_n2650_13878.t87 a_n8300_8799.t18 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 a_n2472_13878.t4 a_n2650_13878.t88 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X285 vdd.t36 vdd.t33 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X286 vdd.t120 a_n8300_8799.t112 CSoutput.t29 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 CSoutput.t28 a_n8300_8799.t113 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 vdd.t32 vdd.t29 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X289 vdd.t28 vdd.t25 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 minus.t0 gnd.t73 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X291 gnd.t64 gnd.t62 plus.t0 gnd.t63 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X292 a_n2903_n3924.t17 plus.t21 a_n8300_8799.t7 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X293 output.t16 outputibias.t11 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X294 a_n2650_8322.t10 a_n2650_13878.t89 a_n8300_8799.t12 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X295 a_n8300_8799.t19 a_n2650_13878.t90 a_n2650_8322.t9 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X296 a_n2650_13878.t50 minus.t20 a_n2903_n3924.t37 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X297 CSoutput.t132 commonsourceibias.t88 gnd.t263 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t27 a_n8300_8799.t114 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 vdd.t123 a_n8300_8799.t115 CSoutput.t26 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 a_n2650_13878.t49 minus.t21 a_n2903_n3924.t36 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X301 gnd.t61 gnd.t58 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X302 vdd.t191 CSoutput.t161 output.t3 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X303 CSoutput.t25 a_n8300_8799.t116 vdd.t116 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t24 a_n8300_8799.t117 vdd.t255 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 a_n2472_13878.t11 a_n2650_13878.t24 a_n2650_13878.t25 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X306 commonsourceibias.t15 commonsourceibias.t14 gnd.t257 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 output.t2 CSoutput.t162 vdd.t192 gnd.t24 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X308 vdd.t245 a_n8300_8799.t118 CSoutput.t23 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 gnd.t266 commonsourceibias.t89 CSoutput.t135 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 gnd.t265 commonsourceibias.t90 CSoutput.t134 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 output.t1 CSoutput.t163 vdd.t193 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X312 vdd.t115 a_n8300_8799.t119 CSoutput.t22 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 gnd.t57 gnd.t54 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X314 a_n2903_n3924.t43 minus.t22 a_n2650_13878.t56 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X315 a_n2903_n3924.t1 diffpairibias.t22 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X316 CSoutput.t21 a_n8300_8799.t120 vdd.t208 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 a_n8300_8799.t13 a_n2650_13878.t91 a_n2650_8322.t8 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X318 a_n2650_13878.t37 a_n2650_13878.t36 a_n2472_13878.t10 vdd.t137 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X319 gnd.t211 commonsourceibias.t91 CSoutput.t112 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 commonsourceibias.t13 commonsourceibias.t12 gnd.t241 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t20 a_n8300_8799.t121 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t205 a_n8300_8799.t122 CSoutput.t19 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 CSoutput.t18 a_n8300_8799.t123 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 CSoutput.t17 a_n8300_8799.t124 vdd.t108 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 vdd.t106 a_n8300_8799.t125 CSoutput.t16 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 diffpairibias.t3 diffpairibias.t2 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X327 a_n2650_8322.t7 a_n2650_13878.t92 a_n8300_8799.t27 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X328 a_n2650_13878.t58 minus.t23 a_n2903_n3924.t45 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X329 vdd.t257 a_n8300_8799.t126 CSoutput.t15 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 commonsourceibias.t11 commonsourceibias.t10 gnd.t203 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 gnd.t264 commonsourceibias.t92 CSoutput.t133 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 CSoutput.t14 a_n8300_8799.t127 vdd.t246 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X333 CSoutput.t164 a_n2650_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X334 diffpairibias.t1 diffpairibias.t0 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X335 CSoutput.t5 commonsourceibias.t93 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t190 CSoutput.t165 output.t0 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 CSoutput.t13 a_n8300_8799.t128 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 vdd.t135 a_n2650_13878.t93 a_n2472_13878.t7 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X339 vdd.t104 a_n8300_8799.t129 CSoutput.t12 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 gnd.t53 gnd.t50 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X341 CSoutput.t3 commonsourceibias.t94 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 vdd.t262 a_n8300_8799.t130 CSoutput.t11 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 CSoutput.t10 a_n8300_8799.t131 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 commonsourceibias.t9 commonsourceibias.t8 gnd.t258 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 a_n8300_8799.t6 plus.t22 a_n2903_n3924.t16 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 a_n2650_8322.t6 a_n2650_13878.t94 a_n8300_8799.t11 vdd.t133 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X347 CSoutput.t4 commonsourceibias.t95 gnd.t40 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 a_n8300_8799.t29 plus.t23 a_n2903_n3924.t15 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X349 a_n2650_13878.t57 minus.t24 a_n2903_n3924.t44 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X350 vdd.t102 a_n8300_8799.t132 CSoutput.t9 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 CSoutput.t8 a_n8300_8799.t133 vdd.t242 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 vdd.t188 a_n8300_8799.t134 CSoutput.t7 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 gnd.t256 commonsourceibias.t6 commonsourceibias.t7 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 commonsourceibias.t5 commonsourceibias.t4 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 a_n2650_8322.t26 a_n2650_13878.t95 vdd.t132 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X356 a_n2472_13878.t9 a_n2650_13878.t6 a_n2650_13878.t7 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X357 a_n2903_n3924.t14 plus.t24 a_n8300_8799.t36 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X358 commonsourceibias.t3 commonsourceibias.t2 gnd.t186 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X359 a_n2650_13878.t3 a_n2650_13878.t2 a_n2472_13878.t8 vdd.t129 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X360 CSoutput.t6 a_n8300_8799.t135 vdd.t189 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 gnd.t189 commonsourceibias.t0 commonsourceibias.t1 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 a_n2903_n3924.t34 diffpairibias.t23 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X363 gnd.t49 gnd.t46 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
R0 a_n2650_13878.n109 a_n2650_13878.t80 512.366
R1 a_n2650_13878.n99 a_n2650_13878.t70 512.366
R2 a_n2650_13878.n110 a_n2650_13878.t60 512.366
R3 a_n2650_13878.n107 a_n2650_13878.t88 512.366
R4 a_n2650_13878.n100 a_n2650_13878.t77 512.366
R5 a_n2650_13878.n108 a_n2650_13878.t76 512.366
R6 a_n2650_13878.n105 a_n2650_13878.t84 512.366
R7 a_n2650_13878.n101 a_n2650_13878.t69 512.366
R8 a_n2650_13878.n106 a_n2650_13878.t68 512.366
R9 a_n2650_13878.n103 a_n2650_13878.t72 512.366
R10 a_n2650_13878.n102 a_n2650_13878.t82 512.366
R11 a_n2650_13878.n104 a_n2650_13878.t95 512.366
R12 a_n2650_13878.n117 a_n2650_13878.t94 512.366
R13 a_n2650_13878.n116 a_n2650_13878.t73 512.366
R14 a_n2650_13878.n73 a_n2650_13878.t78 512.366
R15 a_n2650_13878.n115 a_n2650_13878.t67 512.366
R16 a_n2650_13878.n114 a_n2650_13878.t83 512.366
R17 a_n2650_13878.n74 a_n2650_13878.t91 512.366
R18 a_n2650_13878.n113 a_n2650_13878.t92 512.366
R19 a_n2650_13878.n112 a_n2650_13878.t62 512.366
R20 a_n2650_13878.n75 a_n2650_13878.t75 512.366
R21 a_n2650_13878.n40 a_n2650_13878.t6 533.335
R22 a_n2650_13878.n118 a_n2650_13878.t18 512.366
R23 a_n2650_13878.n129 a_n2650_13878.t24 512.366
R24 a_n2650_13878.n134 a_n2650_13878.t4 512.366
R25 a_n2650_13878.n133 a_n2650_13878.t12 512.366
R26 a_n2650_13878.n71 a_n2650_13878.t30 512.366
R27 a_n2650_13878.n132 a_n2650_13878.t0 512.366
R28 a_n2650_13878.n131 a_n2650_13878.t36 512.366
R29 a_n2650_13878.n72 a_n2650_13878.t16 512.366
R30 a_n2650_13878.n130 a_n2650_13878.t8 512.366
R31 a_n2650_13878.n91 a_n2650_13878.t22 512.366
R32 a_n2650_13878.n92 a_n2650_13878.t28 512.366
R33 a_n2650_13878.n81 a_n2650_13878.t2 512.366
R34 a_n2650_13878.n93 a_n2650_13878.t32 512.366
R35 a_n2650_13878.n94 a_n2650_13878.t34 512.366
R36 a_n2650_13878.n95 a_n2650_13878.t10 512.366
R37 a_n2650_13878.n96 a_n2650_13878.t20 512.366
R38 a_n2650_13878.n80 a_n2650_13878.t14 512.366
R39 a_n2650_13878.n97 a_n2650_13878.t26 512.366
R40 a_n2650_13878.n84 a_n2650_13878.t66 512.366
R41 a_n2650_13878.n85 a_n2650_13878.t90 512.366
R42 a_n2650_13878.n83 a_n2650_13878.t89 512.366
R43 a_n2650_13878.n86 a_n2650_13878.t64 512.366
R44 a_n2650_13878.n87 a_n2650_13878.t87 512.366
R45 a_n2650_13878.n88 a_n2650_13878.t86 512.366
R46 a_n2650_13878.n89 a_n2650_13878.t61 512.366
R47 a_n2650_13878.n82 a_n2650_13878.t71 512.366
R48 a_n2650_13878.n90 a_n2650_13878.t81 512.366
R49 a_n2650_13878.n4 a_n2650_13878.n69 70.1674
R50 a_n2650_13878.n6 a_n2650_13878.n67 70.1674
R51 a_n2650_13878.n8 a_n2650_13878.n65 70.1674
R52 a_n2650_13878.n11 a_n2650_13878.n63 70.1674
R53 a_n2650_13878.n22 a_n2650_13878.n47 70.1674
R54 a_n2650_13878.n39 a_n2650_13878.n26 80.4688
R55 a_n2650_13878.n39 a_n2650_13878.n130 0.365327
R56 a_n2650_13878.n26 a_n2650_13878.n38 75.0448
R57 a_n2650_13878.n37 a_n2650_13878.n25 70.1674
R58 a_n2650_13878.n132 a_n2650_13878.n37 20.9683
R59 a_n2650_13878.n25 a_n2650_13878.n36 70.3058
R60 a_n2650_13878.n36 a_n2650_13878.n71 20.6913
R61 a_n2650_13878.n35 a_n2650_13878.n27 75.3623
R62 a_n2650_13878.n133 a_n2650_13878.n35 10.5784
R63 a_n2650_13878.n27 a_n2650_13878.n134 161.3
R64 a_n2650_13878.n129 a_n2650_13878.n70 11.843
R65 a_n2650_13878.n40 a_n2650_13878.n34 70.1674
R66 a_n2650_13878.n40 a_n2650_13878.n118 20.9683
R67 a_n2650_13878.n26 a_n2650_13878.n70 74.73
R68 a_n2650_13878.n47 a_n2650_13878.n75 20.9683
R69 a_n2650_13878.n46 a_n2650_13878.n22 74.73
R70 a_n2650_13878.n112 a_n2650_13878.n46 11.843
R71 a_n2650_13878.n45 a_n2650_13878.n21 80.4688
R72 a_n2650_13878.n45 a_n2650_13878.n113 0.365327
R73 a_n2650_13878.n21 a_n2650_13878.n44 75.0448
R74 a_n2650_13878.n43 a_n2650_13878.n23 70.1674
R75 a_n2650_13878.n115 a_n2650_13878.n43 20.9683
R76 a_n2650_13878.n23 a_n2650_13878.n42 70.3058
R77 a_n2650_13878.n42 a_n2650_13878.n73 20.6913
R78 a_n2650_13878.n41 a_n2650_13878.n24 75.3623
R79 a_n2650_13878.n116 a_n2650_13878.n41 10.5784
R80 a_n2650_13878.n24 a_n2650_13878.n117 161.3
R81 a_n2650_13878.n14 a_n2650_13878.n61 70.1674
R82 a_n2650_13878.n18 a_n2650_13878.n54 70.1674
R83 a_n2650_13878.n90 a_n2650_13878.n54 20.9683
R84 a_n2650_13878.n53 a_n2650_13878.n18 74.73
R85 a_n2650_13878.n53 a_n2650_13878.n82 11.843
R86 a_n2650_13878.n17 a_n2650_13878.n52 80.4688
R87 a_n2650_13878.n89 a_n2650_13878.n52 0.365327
R88 a_n2650_13878.n51 a_n2650_13878.n17 75.0448
R89 a_n2650_13878.n19 a_n2650_13878.n50 70.1674
R90 a_n2650_13878.n86 a_n2650_13878.n50 20.9683
R91 a_n2650_13878.n49 a_n2650_13878.n19 70.3058
R92 a_n2650_13878.n49 a_n2650_13878.n83 20.6913
R93 a_n2650_13878.n20 a_n2650_13878.n48 75.3623
R94 a_n2650_13878.n85 a_n2650_13878.n48 10.5784
R95 a_n2650_13878.n84 a_n2650_13878.n20 161.3
R96 a_n2650_13878.n97 a_n2650_13878.n61 20.9683
R97 a_n2650_13878.n60 a_n2650_13878.n14 74.73
R98 a_n2650_13878.n60 a_n2650_13878.n80 11.843
R99 a_n2650_13878.n13 a_n2650_13878.n59 80.4688
R100 a_n2650_13878.n96 a_n2650_13878.n59 0.365327
R101 a_n2650_13878.n58 a_n2650_13878.n13 75.0448
R102 a_n2650_13878.n15 a_n2650_13878.n57 70.1674
R103 a_n2650_13878.n93 a_n2650_13878.n57 20.9683
R104 a_n2650_13878.n56 a_n2650_13878.n15 70.3058
R105 a_n2650_13878.n56 a_n2650_13878.n81 20.6913
R106 a_n2650_13878.n16 a_n2650_13878.n55 75.3623
R107 a_n2650_13878.n92 a_n2650_13878.n55 10.5784
R108 a_n2650_13878.n91 a_n2650_13878.n16 161.3
R109 a_n2650_13878.n104 a_n2650_13878.n63 20.9683
R110 a_n2650_13878.n62 a_n2650_13878.n12 75.0448
R111 a_n2650_13878.n62 a_n2650_13878.n102 11.2134
R112 a_n2650_13878.n12 a_n2650_13878.n103 161.3
R113 a_n2650_13878.n106 a_n2650_13878.n65 20.9683
R114 a_n2650_13878.n64 a_n2650_13878.n9 75.0448
R115 a_n2650_13878.n64 a_n2650_13878.n101 11.2134
R116 a_n2650_13878.n9 a_n2650_13878.n105 161.3
R117 a_n2650_13878.n108 a_n2650_13878.n67 20.9683
R118 a_n2650_13878.n66 a_n2650_13878.n7 75.0448
R119 a_n2650_13878.n66 a_n2650_13878.n100 11.2134
R120 a_n2650_13878.n7 a_n2650_13878.n107 161.3
R121 a_n2650_13878.n110 a_n2650_13878.n69 20.9683
R122 a_n2650_13878.n68 a_n2650_13878.n5 75.0448
R123 a_n2650_13878.n68 a_n2650_13878.n99 11.2134
R124 a_n2650_13878.n5 a_n2650_13878.n109 161.3
R125 a_n2650_13878.n3 a_n2650_13878.n127 81.4626
R126 a_n2650_13878.n1 a_n2650_13878.n122 81.4626
R127 a_n2650_13878.n0 a_n2650_13878.n119 81.4626
R128 a_n2650_13878.n3 a_n2650_13878.n128 80.9324
R129 a_n2650_13878.n3 a_n2650_13878.n126 80.9324
R130 a_n2650_13878.n2 a_n2650_13878.n125 80.9324
R131 a_n2650_13878.n2 a_n2650_13878.n124 80.9324
R132 a_n2650_13878.n1 a_n2650_13878.n123 80.9324
R133 a_n2650_13878.n1 a_n2650_13878.n121 80.9324
R134 a_n2650_13878.n0 a_n2650_13878.n120 80.9324
R135 a_n2650_13878.n31 a_n2650_13878.t7 74.6477
R136 a_n2650_13878.n28 a_n2650_13878.t23 74.6477
R137 a_n2650_13878.n32 a_n2650_13878.t5 74.2899
R138 a_n2650_13878.n30 a_n2650_13878.t39 74.2897
R139 a_n2650_13878.n31 a_n2650_13878.n137 70.6783
R140 a_n2650_13878.n31 a_n2650_13878.n138 70.6783
R141 a_n2650_13878.n33 a_n2650_13878.n136 70.6783
R142 a_n2650_13878.n30 a_n2650_13878.n79 70.6783
R143 a_n2650_13878.n29 a_n2650_13878.n78 70.6783
R144 a_n2650_13878.n29 a_n2650_13878.n77 70.6783
R145 a_n2650_13878.n28 a_n2650_13878.n76 70.6783
R146 a_n2650_13878.n139 a_n2650_13878.n33 70.6782
R147 a_n2650_13878.n109 a_n2650_13878.n99 48.2005
R148 a_n2650_13878.t85 a_n2650_13878.n69 533.335
R149 a_n2650_13878.n107 a_n2650_13878.n100 48.2005
R150 a_n2650_13878.t93 a_n2650_13878.n67 533.335
R151 a_n2650_13878.n105 a_n2650_13878.n101 48.2005
R152 a_n2650_13878.t79 a_n2650_13878.n65 533.335
R153 a_n2650_13878.n103 a_n2650_13878.n102 48.2005
R154 a_n2650_13878.t74 a_n2650_13878.n63 533.335
R155 a_n2650_13878.n117 a_n2650_13878.n116 48.2005
R156 a_n2650_13878.n43 a_n2650_13878.n114 20.9683
R157 a_n2650_13878.n113 a_n2650_13878.n74 48.2005
R158 a_n2650_13878.t65 a_n2650_13878.n47 533.335
R159 a_n2650_13878.n134 a_n2650_13878.n133 48.2005
R160 a_n2650_13878.n37 a_n2650_13878.n131 20.9683
R161 a_n2650_13878.n130 a_n2650_13878.n72 48.2005
R162 a_n2650_13878.n92 a_n2650_13878.n91 48.2005
R163 a_n2650_13878.n94 a_n2650_13878.n57 20.9683
R164 a_n2650_13878.n96 a_n2650_13878.n95 48.2005
R165 a_n2650_13878.t38 a_n2650_13878.n61 533.335
R166 a_n2650_13878.n85 a_n2650_13878.n84 48.2005
R167 a_n2650_13878.n87 a_n2650_13878.n50 20.9683
R168 a_n2650_13878.n89 a_n2650_13878.n88 48.2005
R169 a_n2650_13878.t63 a_n2650_13878.n54 533.335
R170 a_n2650_13878.n115 a_n2650_13878.n42 21.4216
R171 a_n2650_13878.n132 a_n2650_13878.n36 21.4216
R172 a_n2650_13878.n93 a_n2650_13878.n56 21.4216
R173 a_n2650_13878.n86 a_n2650_13878.n49 21.4216
R174 a_n2650_13878.n2 a_n2650_13878.n1 32.7898
R175 a_n2650_13878.n46 a_n2650_13878.n75 34.4824
R176 a_n2650_13878.n70 a_n2650_13878.n118 34.4824
R177 a_n2650_13878.n97 a_n2650_13878.n60 34.4824
R178 a_n2650_13878.n90 a_n2650_13878.n53 34.4824
R179 a_n2650_13878.n110 a_n2650_13878.n68 35.3134
R180 a_n2650_13878.n108 a_n2650_13878.n66 35.3134
R181 a_n2650_13878.n106 a_n2650_13878.n64 35.3134
R182 a_n2650_13878.n104 a_n2650_13878.n62 35.3134
R183 a_n2650_13878.n114 a_n2650_13878.n44 35.3134
R184 a_n2650_13878.n44 a_n2650_13878.n74 11.2134
R185 a_n2650_13878.n131 a_n2650_13878.n38 35.3134
R186 a_n2650_13878.n38 a_n2650_13878.n72 11.2134
R187 a_n2650_13878.n94 a_n2650_13878.n58 35.3134
R188 a_n2650_13878.n95 a_n2650_13878.n58 11.2134
R189 a_n2650_13878.n87 a_n2650_13878.n51 35.3134
R190 a_n2650_13878.n88 a_n2650_13878.n51 11.2134
R191 a_n2650_13878.n26 a_n2650_13878.n3 23.891
R192 a_n2650_13878.n41 a_n2650_13878.n73 36.139
R193 a_n2650_13878.n35 a_n2650_13878.n71 36.139
R194 a_n2650_13878.n81 a_n2650_13878.n55 36.139
R195 a_n2650_13878.n83 a_n2650_13878.n48 36.139
R196 a_n2650_13878.n20 a_n2650_13878.n10 13.3641
R197 a_n2650_13878.n22 a_n2650_13878.n111 13.1596
R198 a_n2650_13878.n135 a_n2650_13878.n27 11.8547
R199 a_n2650_13878.n98 a_n2650_13878.n30 10.2167
R200 a_n2650_13878.n111 a_n2650_13878.n4 9.99103
R201 a_n2650_13878.n12 a_n2650_13878.n10 9.99103
R202 a_n2650_13878.n98 a_n2650_13878.n14 8.01944
R203 a_n2650_13878.n32 a_n2650_13878.n135 6.37334
R204 a_n2650_13878.n111 a_n2650_13878.n98 5.3452
R205 a_n2650_13878.n34 a_n2650_13878.n24 4.07247
R206 a_n2650_13878.n16 a_n2650_13878.n18 4.07247
R207 a_n2650_13878.n137 a_n2650_13878.t25 3.61217
R208 a_n2650_13878.n137 a_n2650_13878.t19 3.61217
R209 a_n2650_13878.n138 a_n2650_13878.t17 3.61217
R210 a_n2650_13878.n138 a_n2650_13878.t9 3.61217
R211 a_n2650_13878.n136 a_n2650_13878.t13 3.61217
R212 a_n2650_13878.n136 a_n2650_13878.t31 3.61217
R213 a_n2650_13878.n79 a_n2650_13878.t15 3.61217
R214 a_n2650_13878.n79 a_n2650_13878.t27 3.61217
R215 a_n2650_13878.n78 a_n2650_13878.t11 3.61217
R216 a_n2650_13878.n78 a_n2650_13878.t21 3.61217
R217 a_n2650_13878.n77 a_n2650_13878.t33 3.61217
R218 a_n2650_13878.n77 a_n2650_13878.t35 3.61217
R219 a_n2650_13878.n76 a_n2650_13878.t29 3.61217
R220 a_n2650_13878.n76 a_n2650_13878.t3 3.61217
R221 a_n2650_13878.t1 a_n2650_13878.n139 3.61217
R222 a_n2650_13878.n139 a_n2650_13878.t37 3.61217
R223 a_n2650_13878.n127 a_n2650_13878.t51 2.82907
R224 a_n2650_13878.n127 a_n2650_13878.t57 2.82907
R225 a_n2650_13878.n128 a_n2650_13878.t43 2.82907
R226 a_n2650_13878.n128 a_n2650_13878.t47 2.82907
R227 a_n2650_13878.n126 a_n2650_13878.t59 2.82907
R228 a_n2650_13878.n126 a_n2650_13878.t42 2.82907
R229 a_n2650_13878.n125 a_n2650_13878.t52 2.82907
R230 a_n2650_13878.n125 a_n2650_13878.t55 2.82907
R231 a_n2650_13878.n124 a_n2650_13878.t48 2.82907
R232 a_n2650_13878.n124 a_n2650_13878.t49 2.82907
R233 a_n2650_13878.n122 a_n2650_13878.t46 2.82907
R234 a_n2650_13878.n122 a_n2650_13878.t45 2.82907
R235 a_n2650_13878.n123 a_n2650_13878.t53 2.82907
R236 a_n2650_13878.n123 a_n2650_13878.t50 2.82907
R237 a_n2650_13878.n121 a_n2650_13878.t56 2.82907
R238 a_n2650_13878.n121 a_n2650_13878.t58 2.82907
R239 a_n2650_13878.n120 a_n2650_13878.t40 2.82907
R240 a_n2650_13878.n120 a_n2650_13878.t41 2.82907
R241 a_n2650_13878.n119 a_n2650_13878.t54 2.82907
R242 a_n2650_13878.n119 a_n2650_13878.t44 2.82907
R243 a_n2650_13878.n135 a_n2650_13878.n10 1.30542
R244 a_n2650_13878.n7 a_n2650_13878.n8 1.04595
R245 a_n2650_13878.n45 a_n2650_13878.n112 47.835
R246 a_n2650_13878.n39 a_n2650_13878.n129 47.835
R247 a_n2650_13878.n80 a_n2650_13878.n59 47.835
R248 a_n2650_13878.n82 a_n2650_13878.n52 47.835
R249 a_n2650_13878.n3 a_n2650_13878.n2 1.59102
R250 a_n2650_13878.n22 a_n2650_13878.n21 1.13686
R251 a_n2650_13878.n18 a_n2650_13878.n17 1.13686
R252 a_n2650_13878.n14 a_n2650_13878.n13 1.13686
R253 a_n2650_13878.n26 a_n2650_13878.n34 1.09898
R254 a_n2650_13878.n1 a_n2650_13878.n0 1.06084
R255 a_n2650_13878.n27 a_n2650_13878.n25 0.758076
R256 a_n2650_13878.n26 a_n2650_13878.n25 0.758076
R257 a_n2650_13878.n24 a_n2650_13878.n23 0.758076
R258 a_n2650_13878.n21 a_n2650_13878.n23 0.758076
R259 a_n2650_13878.n19 a_n2650_13878.n20 0.758076
R260 a_n2650_13878.n17 a_n2650_13878.n19 0.758076
R261 a_n2650_13878.n15 a_n2650_13878.n16 0.758076
R262 a_n2650_13878.n13 a_n2650_13878.n15 0.758076
R263 a_n2650_13878.n12 a_n2650_13878.n11 0.758076
R264 a_n2650_13878.n9 a_n2650_13878.n8 0.758076
R265 a_n2650_13878.n7 a_n2650_13878.n6 0.758076
R266 a_n2650_13878.n5 a_n2650_13878.n4 0.758076
R267 a_n2650_13878.n33 a_n2650_13878.n31 0.716017
R268 a_n2650_13878.n33 a_n2650_13878.n32 0.716017
R269 a_n2650_13878.n30 a_n2650_13878.n29 0.716017
R270 a_n2650_13878.n29 a_n2650_13878.n28 0.716017
R271 a_n2650_13878.n9 a_n2650_13878.n11 0.67853
R272 a_n2650_13878.n5 a_n2650_13878.n6 0.67853
R273 a_n2472_13878.n2 a_n2472_13878.n0 98.9633
R274 a_n2472_13878.n5 a_n2472_13878.n3 98.7517
R275 a_n2472_13878.n23 a_n2472_13878.n22 98.6055
R276 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R277 a_n2472_13878.n11 a_n2472_13878.n10 98.6055
R278 a_n2472_13878.n9 a_n2472_13878.n8 98.6055
R279 a_n2472_13878.n7 a_n2472_13878.n6 98.6055
R280 a_n2472_13878.n5 a_n2472_13878.n4 98.6055
R281 a_n2472_13878.n25 a_n2472_13878.n24 98.6054
R282 a_n2472_13878.n21 a_n2472_13878.n20 98.6054
R283 a_n2472_13878.n13 a_n2472_13878.t4 74.6477
R284 a_n2472_13878.n18 a_n2472_13878.t5 74.2899
R285 a_n2472_13878.n15 a_n2472_13878.t6 74.2899
R286 a_n2472_13878.n14 a_n2472_13878.t7 74.2899
R287 a_n2472_13878.n17 a_n2472_13878.n16 70.6783
R288 a_n2472_13878.n13 a_n2472_13878.n12 70.6783
R289 a_n2472_13878.n19 a_n2472_13878.n11 15.0004
R290 a_n2472_13878.n21 a_n2472_13878.n19 12.2917
R291 a_n2472_13878.n19 a_n2472_13878.n18 7.67184
R292 a_n2472_13878.n20 a_n2472_13878.t24 3.61217
R293 a_n2472_13878.n20 a_n2472_13878.t13 3.61217
R294 a_n2472_13878.n22 a_n2472_13878.t16 3.61217
R295 a_n2472_13878.n22 a_n2472_13878.t17 3.61217
R296 a_n2472_13878.n1 a_n2472_13878.t8 3.61217
R297 a_n2472_13878.n1 a_n2472_13878.t18 3.61217
R298 a_n2472_13878.n0 a_n2472_13878.t21 3.61217
R299 a_n2472_13878.n0 a_n2472_13878.t27 3.61217
R300 a_n2472_13878.n16 a_n2472_13878.t0 3.61217
R301 a_n2472_13878.n16 a_n2472_13878.t1 3.61217
R302 a_n2472_13878.n12 a_n2472_13878.t2 3.61217
R303 a_n2472_13878.n12 a_n2472_13878.t3 3.61217
R304 a_n2472_13878.n10 a_n2472_13878.t19 3.61217
R305 a_n2472_13878.n10 a_n2472_13878.t9 3.61217
R306 a_n2472_13878.n8 a_n2472_13878.t22 3.61217
R307 a_n2472_13878.n8 a_n2472_13878.t11 3.61217
R308 a_n2472_13878.n6 a_n2472_13878.t10 3.61217
R309 a_n2472_13878.n6 a_n2472_13878.t12 3.61217
R310 a_n2472_13878.n4 a_n2472_13878.t20 3.61217
R311 a_n2472_13878.n4 a_n2472_13878.t14 3.61217
R312 a_n2472_13878.n3 a_n2472_13878.t23 3.61217
R313 a_n2472_13878.n3 a_n2472_13878.t15 3.61217
R314 a_n2472_13878.n25 a_n2472_13878.t25 3.61217
R315 a_n2472_13878.t26 a_n2472_13878.n25 3.61217
R316 a_n2472_13878.n14 a_n2472_13878.n13 0.358259
R317 a_n2472_13878.n17 a_n2472_13878.n15 0.358259
R318 a_n2472_13878.n18 a_n2472_13878.n17 0.358259
R319 a_n2472_13878.n24 a_n2472_13878.n2 0.358259
R320 a_n2472_13878.n24 a_n2472_13878.n23 0.358259
R321 a_n2472_13878.n23 a_n2472_13878.n21 0.358259
R322 a_n2472_13878.n7 a_n2472_13878.n5 0.146627
R323 a_n2472_13878.n9 a_n2472_13878.n7 0.146627
R324 a_n2472_13878.n11 a_n2472_13878.n9 0.146627
R325 a_n2472_13878.n15 a_n2472_13878.n14 0.101793
R326 vdd.n315 vdd.n279 756.745
R327 vdd.n260 vdd.n224 756.745
R328 vdd.n217 vdd.n181 756.745
R329 vdd.n162 vdd.n126 756.745
R330 vdd.n120 vdd.n84 756.745
R331 vdd.n65 vdd.n29 756.745
R332 vdd.n1764 vdd.n1728 756.745
R333 vdd.n1819 vdd.n1783 756.745
R334 vdd.n1666 vdd.n1630 756.745
R335 vdd.n1721 vdd.n1685 756.745
R336 vdd.n1569 vdd.n1533 756.745
R337 vdd.n1624 vdd.n1588 756.745
R338 vdd.n1107 vdd.t33 640.208
R339 vdd.n968 vdd.t71 640.208
R340 vdd.n1101 vdd.t98 640.208
R341 vdd.n959 vdd.t95 640.208
R342 vdd.n856 vdd.t44 640.208
R343 vdd.n2678 vdd.t89 640.208
R344 vdd.n804 vdd.t65 640.208
R345 vdd.n2747 vdd.t75 640.208
R346 vdd.n768 vdd.t29 640.208
R347 vdd.n1029 vdd.t85 640.208
R348 vdd.n1228 vdd.t55 592.009
R349 vdd.n1384 vdd.t79 592.009
R350 vdd.n1420 vdd.t92 592.009
R351 vdd.n2117 vdd.t51 592.009
R352 vdd.n1967 vdd.t68 592.009
R353 vdd.n1927 vdd.t82 592.009
R354 vdd.n405 vdd.t59 592.009
R355 vdd.n419 vdd.t37 592.009
R356 vdd.n431 vdd.t62 592.009
R357 vdd.n723 vdd.t25 592.009
R358 vdd.n686 vdd.t41 592.009
R359 vdd.n3195 vdd.t48 592.009
R360 vdd.n316 vdd.n315 585
R361 vdd.n314 vdd.n281 585
R362 vdd.n313 vdd.n312 585
R363 vdd.n284 vdd.n282 585
R364 vdd.n307 vdd.n306 585
R365 vdd.n305 vdd.n304 585
R366 vdd.n288 vdd.n287 585
R367 vdd.n299 vdd.n298 585
R368 vdd.n297 vdd.n296 585
R369 vdd.n292 vdd.n291 585
R370 vdd.n261 vdd.n260 585
R371 vdd.n259 vdd.n226 585
R372 vdd.n258 vdd.n257 585
R373 vdd.n229 vdd.n227 585
R374 vdd.n252 vdd.n251 585
R375 vdd.n250 vdd.n249 585
R376 vdd.n233 vdd.n232 585
R377 vdd.n244 vdd.n243 585
R378 vdd.n242 vdd.n241 585
R379 vdd.n237 vdd.n236 585
R380 vdd.n218 vdd.n217 585
R381 vdd.n216 vdd.n183 585
R382 vdd.n215 vdd.n214 585
R383 vdd.n186 vdd.n184 585
R384 vdd.n209 vdd.n208 585
R385 vdd.n207 vdd.n206 585
R386 vdd.n190 vdd.n189 585
R387 vdd.n201 vdd.n200 585
R388 vdd.n199 vdd.n198 585
R389 vdd.n194 vdd.n193 585
R390 vdd.n163 vdd.n162 585
R391 vdd.n161 vdd.n128 585
R392 vdd.n160 vdd.n159 585
R393 vdd.n131 vdd.n129 585
R394 vdd.n154 vdd.n153 585
R395 vdd.n152 vdd.n151 585
R396 vdd.n135 vdd.n134 585
R397 vdd.n146 vdd.n145 585
R398 vdd.n144 vdd.n143 585
R399 vdd.n139 vdd.n138 585
R400 vdd.n121 vdd.n120 585
R401 vdd.n119 vdd.n86 585
R402 vdd.n118 vdd.n117 585
R403 vdd.n89 vdd.n87 585
R404 vdd.n112 vdd.n111 585
R405 vdd.n110 vdd.n109 585
R406 vdd.n93 vdd.n92 585
R407 vdd.n104 vdd.n103 585
R408 vdd.n102 vdd.n101 585
R409 vdd.n97 vdd.n96 585
R410 vdd.n66 vdd.n65 585
R411 vdd.n64 vdd.n31 585
R412 vdd.n63 vdd.n62 585
R413 vdd.n34 vdd.n32 585
R414 vdd.n57 vdd.n56 585
R415 vdd.n55 vdd.n54 585
R416 vdd.n38 vdd.n37 585
R417 vdd.n49 vdd.n48 585
R418 vdd.n47 vdd.n46 585
R419 vdd.n42 vdd.n41 585
R420 vdd.n1765 vdd.n1764 585
R421 vdd.n1763 vdd.n1730 585
R422 vdd.n1762 vdd.n1761 585
R423 vdd.n1733 vdd.n1731 585
R424 vdd.n1756 vdd.n1755 585
R425 vdd.n1754 vdd.n1753 585
R426 vdd.n1737 vdd.n1736 585
R427 vdd.n1748 vdd.n1747 585
R428 vdd.n1746 vdd.n1745 585
R429 vdd.n1741 vdd.n1740 585
R430 vdd.n1820 vdd.n1819 585
R431 vdd.n1818 vdd.n1785 585
R432 vdd.n1817 vdd.n1816 585
R433 vdd.n1788 vdd.n1786 585
R434 vdd.n1811 vdd.n1810 585
R435 vdd.n1809 vdd.n1808 585
R436 vdd.n1792 vdd.n1791 585
R437 vdd.n1803 vdd.n1802 585
R438 vdd.n1801 vdd.n1800 585
R439 vdd.n1796 vdd.n1795 585
R440 vdd.n1667 vdd.n1666 585
R441 vdd.n1665 vdd.n1632 585
R442 vdd.n1664 vdd.n1663 585
R443 vdd.n1635 vdd.n1633 585
R444 vdd.n1658 vdd.n1657 585
R445 vdd.n1656 vdd.n1655 585
R446 vdd.n1639 vdd.n1638 585
R447 vdd.n1650 vdd.n1649 585
R448 vdd.n1648 vdd.n1647 585
R449 vdd.n1643 vdd.n1642 585
R450 vdd.n1722 vdd.n1721 585
R451 vdd.n1720 vdd.n1687 585
R452 vdd.n1719 vdd.n1718 585
R453 vdd.n1690 vdd.n1688 585
R454 vdd.n1713 vdd.n1712 585
R455 vdd.n1711 vdd.n1710 585
R456 vdd.n1694 vdd.n1693 585
R457 vdd.n1705 vdd.n1704 585
R458 vdd.n1703 vdd.n1702 585
R459 vdd.n1698 vdd.n1697 585
R460 vdd.n1570 vdd.n1569 585
R461 vdd.n1568 vdd.n1535 585
R462 vdd.n1567 vdd.n1566 585
R463 vdd.n1538 vdd.n1536 585
R464 vdd.n1561 vdd.n1560 585
R465 vdd.n1559 vdd.n1558 585
R466 vdd.n1542 vdd.n1541 585
R467 vdd.n1553 vdd.n1552 585
R468 vdd.n1551 vdd.n1550 585
R469 vdd.n1546 vdd.n1545 585
R470 vdd.n1625 vdd.n1624 585
R471 vdd.n1623 vdd.n1590 585
R472 vdd.n1622 vdd.n1621 585
R473 vdd.n1593 vdd.n1591 585
R474 vdd.n1616 vdd.n1615 585
R475 vdd.n1614 vdd.n1613 585
R476 vdd.n1597 vdd.n1596 585
R477 vdd.n1608 vdd.n1607 585
R478 vdd.n1606 vdd.n1605 585
R479 vdd.n1601 vdd.n1600 585
R480 vdd.n445 vdd.n370 462.44
R481 vdd.n3433 vdd.n372 462.44
R482 vdd.n3328 vdd.n657 462.44
R483 vdd.n3326 vdd.n660 462.44
R484 vdd.n2112 vdd.n1127 462.44
R485 vdd.n2115 vdd.n2114 462.44
R486 vdd.n1455 vdd.n1225 462.44
R487 vdd.n1452 vdd.n1223 462.44
R488 vdd.n293 vdd.t246 329.043
R489 vdd.n238 vdd.t267 329.043
R490 vdd.n195 vdd.t211 329.043
R491 vdd.n140 vdd.t227 329.043
R492 vdd.n98 vdd.t225 329.043
R493 vdd.n43 vdd.t216 329.043
R494 vdd.n1742 vdd.t235 329.043
R495 vdd.n1797 vdd.t201 329.043
R496 vdd.n1644 vdd.t249 329.043
R497 vdd.n1699 vdd.t22 329.043
R498 vdd.n1547 vdd.t239 329.043
R499 vdd.n1602 vdd.t203 329.043
R500 vdd.n1228 vdd.t58 319.788
R501 vdd.n1384 vdd.t81 319.788
R502 vdd.n1420 vdd.t94 319.788
R503 vdd.n2117 vdd.t53 319.788
R504 vdd.n1967 vdd.t69 319.788
R505 vdd.n1927 vdd.t83 319.788
R506 vdd.n405 vdd.t60 319.788
R507 vdd.n419 vdd.t39 319.788
R508 vdd.n431 vdd.t63 319.788
R509 vdd.n723 vdd.t28 319.788
R510 vdd.n686 vdd.t43 319.788
R511 vdd.n3195 vdd.t50 319.788
R512 vdd.n1229 vdd.t57 303.69
R513 vdd.n1385 vdd.t80 303.69
R514 vdd.n1421 vdd.t93 303.69
R515 vdd.n2118 vdd.t54 303.69
R516 vdd.n1968 vdd.t70 303.69
R517 vdd.n1928 vdd.t84 303.69
R518 vdd.n406 vdd.t61 303.69
R519 vdd.n420 vdd.t40 303.69
R520 vdd.n432 vdd.t64 303.69
R521 vdd.n724 vdd.t27 303.69
R522 vdd.n687 vdd.t42 303.69
R523 vdd.n3196 vdd.t49 303.69
R524 vdd.n2933 vdd.n918 285.366
R525 vdd.n3157 vdd.n778 285.366
R526 vdd.n3094 vdd.n775 285.366
R527 vdd.n2812 vdd.n915 285.366
R528 vdd.n2642 vdd.n956 285.366
R529 vdd.n2573 vdd.n2572 285.366
R530 vdd.n2313 vdd.n1082 285.366
R531 vdd.n2383 vdd.n1084 285.366
R532 vdd.n3073 vdd.n776 285.366
R533 vdd.n3160 vdd.n3159 285.366
R534 vdd.n2926 vdd.n916 285.366
R535 vdd.n2935 vdd.n914 285.366
R536 vdd.n2570 vdd.n966 285.366
R537 vdd.n964 vdd.n938 285.366
R538 vdd.n2199 vdd.n1083 285.366
R539 vdd.n2385 vdd.n1080 285.366
R540 vdd.n1125 vdd.n1081 216.982
R541 vdd.n756 vdd.n658 216.982
R542 vdd.n3075 vdd.n776 185
R543 vdd.n3158 vdd.n776 185
R544 vdd.n3077 vdd.n3076 185
R545 vdd.n3076 vdd.n774 185
R546 vdd.n3078 vdd.n810 185
R547 vdd.n3088 vdd.n810 185
R548 vdd.n3079 vdd.n819 185
R549 vdd.n819 vdd.n817 185
R550 vdd.n3081 vdd.n3080 185
R551 vdd.n3082 vdd.n3081 185
R552 vdd.n3034 vdd.n818 185
R553 vdd.n818 vdd.n814 185
R554 vdd.n3033 vdd.n3032 185
R555 vdd.n3032 vdd.n3031 185
R556 vdd.n821 vdd.n820 185
R557 vdd.n822 vdd.n821 185
R558 vdd.n3024 vdd.n3023 185
R559 vdd.n3025 vdd.n3024 185
R560 vdd.n3022 vdd.n830 185
R561 vdd.n835 vdd.n830 185
R562 vdd.n3021 vdd.n3020 185
R563 vdd.n3020 vdd.n3019 185
R564 vdd.n832 vdd.n831 185
R565 vdd.n841 vdd.n832 185
R566 vdd.n3012 vdd.n3011 185
R567 vdd.n3013 vdd.n3012 185
R568 vdd.n3010 vdd.n842 185
R569 vdd.n848 vdd.n842 185
R570 vdd.n3009 vdd.n3008 185
R571 vdd.n3008 vdd.n3007 185
R572 vdd.n844 vdd.n843 185
R573 vdd.n845 vdd.n844 185
R574 vdd.n3000 vdd.n2999 185
R575 vdd.n3001 vdd.n3000 185
R576 vdd.n2998 vdd.n855 185
R577 vdd.n855 vdd.n852 185
R578 vdd.n2996 vdd.n2995 185
R579 vdd.n2995 vdd.n2994 185
R580 vdd.n858 vdd.n857 185
R581 vdd.n859 vdd.n858 185
R582 vdd.n2987 vdd.n2986 185
R583 vdd.n2988 vdd.n2987 185
R584 vdd.n2985 vdd.n867 185
R585 vdd.n872 vdd.n867 185
R586 vdd.n2984 vdd.n2983 185
R587 vdd.n2983 vdd.n2982 185
R588 vdd.n869 vdd.n868 185
R589 vdd.n2894 vdd.n869 185
R590 vdd.n2975 vdd.n2974 185
R591 vdd.n2976 vdd.n2975 185
R592 vdd.n2973 vdd.n879 185
R593 vdd.n879 vdd.n876 185
R594 vdd.n2972 vdd.n2971 185
R595 vdd.n2971 vdd.n2970 185
R596 vdd.n881 vdd.n880 185
R597 vdd.n882 vdd.n881 185
R598 vdd.n2963 vdd.n2962 185
R599 vdd.n2964 vdd.n2963 185
R600 vdd.n2961 vdd.n890 185
R601 vdd.n2906 vdd.n890 185
R602 vdd.n2960 vdd.n2959 185
R603 vdd.n2959 vdd.n2958 185
R604 vdd.n892 vdd.n891 185
R605 vdd.n901 vdd.n892 185
R606 vdd.n2951 vdd.n2950 185
R607 vdd.n2952 vdd.n2951 185
R608 vdd.n2949 vdd.n902 185
R609 vdd.n902 vdd.n898 185
R610 vdd.n2948 vdd.n2947 185
R611 vdd.n2947 vdd.n2946 185
R612 vdd.n904 vdd.n903 185
R613 vdd.n2918 vdd.n904 185
R614 vdd.n2939 vdd.n2938 185
R615 vdd.n2940 vdd.n2939 185
R616 vdd.n2937 vdd.n912 185
R617 vdd.n917 vdd.n912 185
R618 vdd.n2936 vdd.n2935 185
R619 vdd.n2935 vdd.n2934 185
R620 vdd.n914 vdd.n913 185
R621 vdd.n2682 vdd.n2681 185
R622 vdd.n2684 vdd.n2683 185
R623 vdd.n2686 vdd.n2685 185
R624 vdd.n2688 vdd.n2687 185
R625 vdd.n2690 vdd.n2689 185
R626 vdd.n2692 vdd.n2691 185
R627 vdd.n2694 vdd.n2693 185
R628 vdd.n2696 vdd.n2695 185
R629 vdd.n2698 vdd.n2697 185
R630 vdd.n2700 vdd.n2699 185
R631 vdd.n2702 vdd.n2701 185
R632 vdd.n2704 vdd.n2703 185
R633 vdd.n2706 vdd.n2705 185
R634 vdd.n2708 vdd.n2707 185
R635 vdd.n2710 vdd.n2709 185
R636 vdd.n2712 vdd.n2711 185
R637 vdd.n2714 vdd.n2713 185
R638 vdd.n2716 vdd.n2715 185
R639 vdd.n2718 vdd.n2717 185
R640 vdd.n2720 vdd.n2719 185
R641 vdd.n2722 vdd.n2721 185
R642 vdd.n2724 vdd.n2723 185
R643 vdd.n2726 vdd.n2725 185
R644 vdd.n2728 vdd.n2727 185
R645 vdd.n2730 vdd.n2729 185
R646 vdd.n2732 vdd.n2731 185
R647 vdd.n2734 vdd.n2733 185
R648 vdd.n2736 vdd.n2735 185
R649 vdd.n2738 vdd.n2737 185
R650 vdd.n2740 vdd.n2739 185
R651 vdd.n2742 vdd.n2741 185
R652 vdd.n2744 vdd.n2743 185
R653 vdd.n2745 vdd.n2677 185
R654 vdd.n2926 vdd.n2925 185
R655 vdd.n2927 vdd.n2926 185
R656 vdd.n3161 vdd.n3160 185
R657 vdd.n3162 vdd.n767 185
R658 vdd.n3164 vdd.n3163 185
R659 vdd.n3166 vdd.n765 185
R660 vdd.n3168 vdd.n3167 185
R661 vdd.n3169 vdd.n764 185
R662 vdd.n3171 vdd.n3170 185
R663 vdd.n3173 vdd.n762 185
R664 vdd.n3175 vdd.n3174 185
R665 vdd.n3176 vdd.n761 185
R666 vdd.n3178 vdd.n3177 185
R667 vdd.n3180 vdd.n759 185
R668 vdd.n3182 vdd.n3181 185
R669 vdd.n3183 vdd.n758 185
R670 vdd.n3185 vdd.n3184 185
R671 vdd.n3187 vdd.n757 185
R672 vdd.n3188 vdd.n754 185
R673 vdd.n3191 vdd.n3190 185
R674 vdd.n755 vdd.n753 185
R675 vdd.n3047 vdd.n3046 185
R676 vdd.n3049 vdd.n3048 185
R677 vdd.n3051 vdd.n3043 185
R678 vdd.n3053 vdd.n3052 185
R679 vdd.n3054 vdd.n3042 185
R680 vdd.n3056 vdd.n3055 185
R681 vdd.n3058 vdd.n3040 185
R682 vdd.n3060 vdd.n3059 185
R683 vdd.n3061 vdd.n3039 185
R684 vdd.n3063 vdd.n3062 185
R685 vdd.n3065 vdd.n3037 185
R686 vdd.n3067 vdd.n3066 185
R687 vdd.n3068 vdd.n3036 185
R688 vdd.n3070 vdd.n3069 185
R689 vdd.n3072 vdd.n3035 185
R690 vdd.n3074 vdd.n3073 185
R691 vdd.n3073 vdd.n756 185
R692 vdd.n3159 vdd.n771 185
R693 vdd.n3159 vdd.n3158 185
R694 vdd.n2825 vdd.n773 185
R695 vdd.n774 vdd.n773 185
R696 vdd.n2826 vdd.n809 185
R697 vdd.n3088 vdd.n809 185
R698 vdd.n2828 vdd.n2827 185
R699 vdd.n2827 vdd.n817 185
R700 vdd.n2829 vdd.n816 185
R701 vdd.n3082 vdd.n816 185
R702 vdd.n2831 vdd.n2830 185
R703 vdd.n2830 vdd.n814 185
R704 vdd.n2832 vdd.n824 185
R705 vdd.n3031 vdd.n824 185
R706 vdd.n2834 vdd.n2833 185
R707 vdd.n2833 vdd.n822 185
R708 vdd.n2835 vdd.n829 185
R709 vdd.n3025 vdd.n829 185
R710 vdd.n2837 vdd.n2836 185
R711 vdd.n2836 vdd.n835 185
R712 vdd.n2838 vdd.n834 185
R713 vdd.n3019 vdd.n834 185
R714 vdd.n2840 vdd.n2839 185
R715 vdd.n2839 vdd.n841 185
R716 vdd.n2841 vdd.n840 185
R717 vdd.n3013 vdd.n840 185
R718 vdd.n2843 vdd.n2842 185
R719 vdd.n2842 vdd.n848 185
R720 vdd.n2844 vdd.n847 185
R721 vdd.n3007 vdd.n847 185
R722 vdd.n2846 vdd.n2845 185
R723 vdd.n2845 vdd.n845 185
R724 vdd.n2847 vdd.n854 185
R725 vdd.n3001 vdd.n854 185
R726 vdd.n2849 vdd.n2848 185
R727 vdd.n2848 vdd.n852 185
R728 vdd.n2850 vdd.n861 185
R729 vdd.n2994 vdd.n861 185
R730 vdd.n2852 vdd.n2851 185
R731 vdd.n2851 vdd.n859 185
R732 vdd.n2853 vdd.n866 185
R733 vdd.n2988 vdd.n866 185
R734 vdd.n2855 vdd.n2854 185
R735 vdd.n2854 vdd.n872 185
R736 vdd.n2856 vdd.n871 185
R737 vdd.n2982 vdd.n871 185
R738 vdd.n2896 vdd.n2895 185
R739 vdd.n2895 vdd.n2894 185
R740 vdd.n2897 vdd.n878 185
R741 vdd.n2976 vdd.n878 185
R742 vdd.n2899 vdd.n2898 185
R743 vdd.n2898 vdd.n876 185
R744 vdd.n2900 vdd.n884 185
R745 vdd.n2970 vdd.n884 185
R746 vdd.n2902 vdd.n2901 185
R747 vdd.n2901 vdd.n882 185
R748 vdd.n2903 vdd.n889 185
R749 vdd.n2964 vdd.n889 185
R750 vdd.n2905 vdd.n2904 185
R751 vdd.n2906 vdd.n2905 185
R752 vdd.n2824 vdd.n894 185
R753 vdd.n2958 vdd.n894 185
R754 vdd.n2823 vdd.n2822 185
R755 vdd.n2822 vdd.n901 185
R756 vdd.n2821 vdd.n900 185
R757 vdd.n2952 vdd.n900 185
R758 vdd.n2820 vdd.n2819 185
R759 vdd.n2819 vdd.n898 185
R760 vdd.n2746 vdd.n906 185
R761 vdd.n2946 vdd.n906 185
R762 vdd.n2920 vdd.n2919 185
R763 vdd.n2919 vdd.n2918 185
R764 vdd.n2921 vdd.n911 185
R765 vdd.n2940 vdd.n911 185
R766 vdd.n2923 vdd.n2922 185
R767 vdd.n2922 vdd.n917 185
R768 vdd.n2924 vdd.n916 185
R769 vdd.n2934 vdd.n916 185
R770 vdd.n2112 vdd.n2111 185
R771 vdd.n2113 vdd.n2112 185
R772 vdd.n1128 vdd.n1126 185
R773 vdd.n1126 vdd.n1124 185
R774 vdd.n1894 vdd.n1893 185
R775 vdd.n1893 vdd.n1892 185
R776 vdd.n1131 vdd.n1130 185
R777 vdd.n1132 vdd.n1131 185
R778 vdd.n1881 vdd.n1880 185
R779 vdd.n1882 vdd.n1881 185
R780 vdd.n1140 vdd.n1139 185
R781 vdd.n1873 vdd.n1139 185
R782 vdd.n1876 vdd.n1875 185
R783 vdd.n1875 vdd.n1874 185
R784 vdd.n1143 vdd.n1142 185
R785 vdd.n1149 vdd.n1143 185
R786 vdd.n1864 vdd.n1863 185
R787 vdd.n1865 vdd.n1864 185
R788 vdd.n1151 vdd.n1150 185
R789 vdd.n1856 vdd.n1150 185
R790 vdd.n1859 vdd.n1858 185
R791 vdd.n1858 vdd.n1857 185
R792 vdd.n1154 vdd.n1153 185
R793 vdd.n1155 vdd.n1154 185
R794 vdd.n1847 vdd.n1846 185
R795 vdd.n1848 vdd.n1847 185
R796 vdd.n1163 vdd.n1162 185
R797 vdd.n1162 vdd.n1161 185
R798 vdd.n1842 vdd.n1841 185
R799 vdd.n1841 vdd.n1840 185
R800 vdd.n1166 vdd.n1165 185
R801 vdd.n1172 vdd.n1166 185
R802 vdd.n1831 vdd.n1830 185
R803 vdd.n1832 vdd.n1831 185
R804 vdd.n1174 vdd.n1173 185
R805 vdd.n1528 vdd.n1173 185
R806 vdd.n1531 vdd.n1530 185
R807 vdd.n1530 vdd.n1529 185
R808 vdd.n1177 vdd.n1176 185
R809 vdd.n1184 vdd.n1177 185
R810 vdd.n1519 vdd.n1518 185
R811 vdd.n1520 vdd.n1519 185
R812 vdd.n1186 vdd.n1185 185
R813 vdd.n1185 vdd.n1183 185
R814 vdd.n1514 vdd.n1513 185
R815 vdd.n1513 vdd.n1512 185
R816 vdd.n1189 vdd.n1188 185
R817 vdd.n1190 vdd.n1189 185
R818 vdd.n1503 vdd.n1502 185
R819 vdd.n1504 vdd.n1503 185
R820 vdd.n1197 vdd.n1196 185
R821 vdd.n1495 vdd.n1196 185
R822 vdd.n1498 vdd.n1497 185
R823 vdd.n1497 vdd.n1496 185
R824 vdd.n1200 vdd.n1199 185
R825 vdd.n1206 vdd.n1200 185
R826 vdd.n1486 vdd.n1485 185
R827 vdd.n1487 vdd.n1486 185
R828 vdd.n1208 vdd.n1207 185
R829 vdd.n1478 vdd.n1207 185
R830 vdd.n1481 vdd.n1480 185
R831 vdd.n1480 vdd.n1479 185
R832 vdd.n1211 vdd.n1210 185
R833 vdd.n1212 vdd.n1211 185
R834 vdd.n1469 vdd.n1468 185
R835 vdd.n1470 vdd.n1469 185
R836 vdd.n1220 vdd.n1219 185
R837 vdd.n1219 vdd.n1218 185
R838 vdd.n1464 vdd.n1463 185
R839 vdd.n1463 vdd.n1462 185
R840 vdd.n1223 vdd.n1222 185
R841 vdd.n1224 vdd.n1223 185
R842 vdd.n1452 vdd.n1451 185
R843 vdd.n1450 vdd.n1263 185
R844 vdd.n1265 vdd.n1262 185
R845 vdd.n1454 vdd.n1262 185
R846 vdd.n1446 vdd.n1267 185
R847 vdd.n1445 vdd.n1268 185
R848 vdd.n1444 vdd.n1269 185
R849 vdd.n1272 vdd.n1270 185
R850 vdd.n1440 vdd.n1273 185
R851 vdd.n1439 vdd.n1274 185
R852 vdd.n1438 vdd.n1275 185
R853 vdd.n1278 vdd.n1276 185
R854 vdd.n1434 vdd.n1279 185
R855 vdd.n1433 vdd.n1280 185
R856 vdd.n1432 vdd.n1281 185
R857 vdd.n1284 vdd.n1282 185
R858 vdd.n1428 vdd.n1285 185
R859 vdd.n1427 vdd.n1286 185
R860 vdd.n1426 vdd.n1287 185
R861 vdd.n1418 vdd.n1288 185
R862 vdd.n1422 vdd.n1419 185
R863 vdd.n1417 vdd.n1290 185
R864 vdd.n1416 vdd.n1291 185
R865 vdd.n1294 vdd.n1292 185
R866 vdd.n1412 vdd.n1295 185
R867 vdd.n1411 vdd.n1296 185
R868 vdd.n1410 vdd.n1297 185
R869 vdd.n1300 vdd.n1298 185
R870 vdd.n1406 vdd.n1301 185
R871 vdd.n1405 vdd.n1302 185
R872 vdd.n1404 vdd.n1303 185
R873 vdd.n1306 vdd.n1304 185
R874 vdd.n1400 vdd.n1307 185
R875 vdd.n1399 vdd.n1308 185
R876 vdd.n1398 vdd.n1309 185
R877 vdd.n1312 vdd.n1310 185
R878 vdd.n1394 vdd.n1313 185
R879 vdd.n1393 vdd.n1314 185
R880 vdd.n1392 vdd.n1315 185
R881 vdd.n1318 vdd.n1316 185
R882 vdd.n1388 vdd.n1319 185
R883 vdd.n1387 vdd.n1320 185
R884 vdd.n1386 vdd.n1383 185
R885 vdd.n1323 vdd.n1321 185
R886 vdd.n1379 vdd.n1324 185
R887 vdd.n1378 vdd.n1325 185
R888 vdd.n1377 vdd.n1326 185
R889 vdd.n1329 vdd.n1327 185
R890 vdd.n1373 vdd.n1330 185
R891 vdd.n1372 vdd.n1331 185
R892 vdd.n1371 vdd.n1332 185
R893 vdd.n1335 vdd.n1333 185
R894 vdd.n1367 vdd.n1336 185
R895 vdd.n1366 vdd.n1337 185
R896 vdd.n1365 vdd.n1338 185
R897 vdd.n1341 vdd.n1339 185
R898 vdd.n1361 vdd.n1342 185
R899 vdd.n1360 vdd.n1343 185
R900 vdd.n1359 vdd.n1344 185
R901 vdd.n1347 vdd.n1345 185
R902 vdd.n1355 vdd.n1348 185
R903 vdd.n1354 vdd.n1349 185
R904 vdd.n1353 vdd.n1350 185
R905 vdd.n1351 vdd.n1231 185
R906 vdd.n1456 vdd.n1455 185
R907 vdd.n1455 vdd.n1454 185
R908 vdd.n2116 vdd.n2115 185
R909 vdd.n2120 vdd.n1120 185
R910 vdd.n1996 vdd.n1119 185
R911 vdd.n1999 vdd.n1998 185
R912 vdd.n2001 vdd.n2000 185
R913 vdd.n2004 vdd.n2003 185
R914 vdd.n2006 vdd.n2005 185
R915 vdd.n2008 vdd.n1994 185
R916 vdd.n2010 vdd.n2009 185
R917 vdd.n2011 vdd.n1988 185
R918 vdd.n2013 vdd.n2012 185
R919 vdd.n2015 vdd.n1986 185
R920 vdd.n2017 vdd.n2016 185
R921 vdd.n2018 vdd.n1981 185
R922 vdd.n2020 vdd.n2019 185
R923 vdd.n2022 vdd.n1979 185
R924 vdd.n2024 vdd.n2023 185
R925 vdd.n2025 vdd.n1975 185
R926 vdd.n2027 vdd.n2026 185
R927 vdd.n2029 vdd.n1972 185
R928 vdd.n2031 vdd.n2030 185
R929 vdd.n1973 vdd.n1966 185
R930 vdd.n2035 vdd.n1970 185
R931 vdd.n2036 vdd.n1962 185
R932 vdd.n2038 vdd.n2037 185
R933 vdd.n2040 vdd.n1960 185
R934 vdd.n2042 vdd.n2041 185
R935 vdd.n2043 vdd.n1955 185
R936 vdd.n2045 vdd.n2044 185
R937 vdd.n2047 vdd.n1953 185
R938 vdd.n2049 vdd.n2048 185
R939 vdd.n2050 vdd.n1948 185
R940 vdd.n2052 vdd.n2051 185
R941 vdd.n2054 vdd.n1946 185
R942 vdd.n2056 vdd.n2055 185
R943 vdd.n2057 vdd.n1941 185
R944 vdd.n2059 vdd.n2058 185
R945 vdd.n2061 vdd.n1939 185
R946 vdd.n2063 vdd.n2062 185
R947 vdd.n2064 vdd.n1935 185
R948 vdd.n2066 vdd.n2065 185
R949 vdd.n2068 vdd.n1932 185
R950 vdd.n2070 vdd.n2069 185
R951 vdd.n1933 vdd.n1926 185
R952 vdd.n2074 vdd.n1930 185
R953 vdd.n2075 vdd.n1922 185
R954 vdd.n2077 vdd.n2076 185
R955 vdd.n2079 vdd.n1920 185
R956 vdd.n2081 vdd.n2080 185
R957 vdd.n2082 vdd.n1915 185
R958 vdd.n2084 vdd.n2083 185
R959 vdd.n2086 vdd.n1913 185
R960 vdd.n2088 vdd.n2087 185
R961 vdd.n2089 vdd.n1908 185
R962 vdd.n2091 vdd.n2090 185
R963 vdd.n2093 vdd.n1907 185
R964 vdd.n2094 vdd.n1904 185
R965 vdd.n2097 vdd.n2096 185
R966 vdd.n1906 vdd.n1902 185
R967 vdd.n2101 vdd.n1900 185
R968 vdd.n2103 vdd.n2102 185
R969 vdd.n2105 vdd.n1898 185
R970 vdd.n2107 vdd.n2106 185
R971 vdd.n2108 vdd.n1127 185
R972 vdd.n2114 vdd.n1123 185
R973 vdd.n2114 vdd.n2113 185
R974 vdd.n1135 vdd.n1122 185
R975 vdd.n1124 vdd.n1122 185
R976 vdd.n1891 vdd.n1890 185
R977 vdd.n1892 vdd.n1891 185
R978 vdd.n1134 vdd.n1133 185
R979 vdd.n1133 vdd.n1132 185
R980 vdd.n1884 vdd.n1883 185
R981 vdd.n1883 vdd.n1882 185
R982 vdd.n1138 vdd.n1137 185
R983 vdd.n1873 vdd.n1138 185
R984 vdd.n1872 vdd.n1871 185
R985 vdd.n1874 vdd.n1872 185
R986 vdd.n1145 vdd.n1144 185
R987 vdd.n1149 vdd.n1144 185
R988 vdd.n1867 vdd.n1866 185
R989 vdd.n1866 vdd.n1865 185
R990 vdd.n1148 vdd.n1147 185
R991 vdd.n1856 vdd.n1148 185
R992 vdd.n1855 vdd.n1854 185
R993 vdd.n1857 vdd.n1855 185
R994 vdd.n1157 vdd.n1156 185
R995 vdd.n1156 vdd.n1155 185
R996 vdd.n1850 vdd.n1849 185
R997 vdd.n1849 vdd.n1848 185
R998 vdd.n1160 vdd.n1159 185
R999 vdd.n1161 vdd.n1160 185
R1000 vdd.n1839 vdd.n1838 185
R1001 vdd.n1840 vdd.n1839 185
R1002 vdd.n1168 vdd.n1167 185
R1003 vdd.n1172 vdd.n1167 185
R1004 vdd.n1834 vdd.n1833 185
R1005 vdd.n1833 vdd.n1832 185
R1006 vdd.n1171 vdd.n1170 185
R1007 vdd.n1528 vdd.n1171 185
R1008 vdd.n1527 vdd.n1526 185
R1009 vdd.n1529 vdd.n1527 185
R1010 vdd.n1179 vdd.n1178 185
R1011 vdd.n1184 vdd.n1178 185
R1012 vdd.n1522 vdd.n1521 185
R1013 vdd.n1521 vdd.n1520 185
R1014 vdd.n1182 vdd.n1181 185
R1015 vdd.n1183 vdd.n1182 185
R1016 vdd.n1511 vdd.n1510 185
R1017 vdd.n1512 vdd.n1511 185
R1018 vdd.n1192 vdd.n1191 185
R1019 vdd.n1191 vdd.n1190 185
R1020 vdd.n1506 vdd.n1505 185
R1021 vdd.n1505 vdd.n1504 185
R1022 vdd.n1195 vdd.n1194 185
R1023 vdd.n1495 vdd.n1195 185
R1024 vdd.n1494 vdd.n1493 185
R1025 vdd.n1496 vdd.n1494 185
R1026 vdd.n1202 vdd.n1201 185
R1027 vdd.n1206 vdd.n1201 185
R1028 vdd.n1489 vdd.n1488 185
R1029 vdd.n1488 vdd.n1487 185
R1030 vdd.n1205 vdd.n1204 185
R1031 vdd.n1478 vdd.n1205 185
R1032 vdd.n1477 vdd.n1476 185
R1033 vdd.n1479 vdd.n1477 185
R1034 vdd.n1214 vdd.n1213 185
R1035 vdd.n1213 vdd.n1212 185
R1036 vdd.n1472 vdd.n1471 185
R1037 vdd.n1471 vdd.n1470 185
R1038 vdd.n1217 vdd.n1216 185
R1039 vdd.n1218 vdd.n1217 185
R1040 vdd.n1461 vdd.n1460 185
R1041 vdd.n1462 vdd.n1461 185
R1042 vdd.n1226 vdd.n1225 185
R1043 vdd.n1225 vdd.n1224 185
R1044 vdd.n958 vdd.n956 185
R1045 vdd.n2571 vdd.n956 185
R1046 vdd.n2493 vdd.n976 185
R1047 vdd.n976 vdd.n963 185
R1048 vdd.n2495 vdd.n2494 185
R1049 vdd.n2496 vdd.n2495 185
R1050 vdd.n2492 vdd.n975 185
R1051 vdd.n2251 vdd.n975 185
R1052 vdd.n2491 vdd.n2490 185
R1053 vdd.n2490 vdd.n2489 185
R1054 vdd.n978 vdd.n977 185
R1055 vdd.n979 vdd.n978 185
R1056 vdd.n2480 vdd.n2479 185
R1057 vdd.n2481 vdd.n2480 185
R1058 vdd.n2478 vdd.n989 185
R1059 vdd.n989 vdd.n986 185
R1060 vdd.n2477 vdd.n2476 185
R1061 vdd.n2476 vdd.n2475 185
R1062 vdd.n991 vdd.n990 185
R1063 vdd.n2263 vdd.n991 185
R1064 vdd.n2468 vdd.n2467 185
R1065 vdd.n2469 vdd.n2468 185
R1066 vdd.n2466 vdd.n999 185
R1067 vdd.n1004 vdd.n999 185
R1068 vdd.n2465 vdd.n2464 185
R1069 vdd.n2464 vdd.n2463 185
R1070 vdd.n1001 vdd.n1000 185
R1071 vdd.n1010 vdd.n1001 185
R1072 vdd.n2456 vdd.n2455 185
R1073 vdd.n2457 vdd.n2456 185
R1074 vdd.n2454 vdd.n1011 185
R1075 vdd.n2275 vdd.n1011 185
R1076 vdd.n2453 vdd.n2452 185
R1077 vdd.n2452 vdd.n2451 185
R1078 vdd.n1013 vdd.n1012 185
R1079 vdd.n1014 vdd.n1013 185
R1080 vdd.n2444 vdd.n2443 185
R1081 vdd.n2445 vdd.n2444 185
R1082 vdd.n2442 vdd.n1023 185
R1083 vdd.n1023 vdd.n1020 185
R1084 vdd.n2441 vdd.n2440 185
R1085 vdd.n2440 vdd.n2439 185
R1086 vdd.n1025 vdd.n1024 185
R1087 vdd.n1034 vdd.n1025 185
R1088 vdd.n2431 vdd.n2430 185
R1089 vdd.n2432 vdd.n2431 185
R1090 vdd.n2429 vdd.n1035 185
R1091 vdd.n1041 vdd.n1035 185
R1092 vdd.n2428 vdd.n2427 185
R1093 vdd.n2427 vdd.n2426 185
R1094 vdd.n1037 vdd.n1036 185
R1095 vdd.n1038 vdd.n1037 185
R1096 vdd.n2419 vdd.n2418 185
R1097 vdd.n2420 vdd.n2419 185
R1098 vdd.n2417 vdd.n1048 185
R1099 vdd.n1048 vdd.n1045 185
R1100 vdd.n2416 vdd.n2415 185
R1101 vdd.n2415 vdd.n2414 185
R1102 vdd.n1050 vdd.n1049 185
R1103 vdd.n1051 vdd.n1050 185
R1104 vdd.n2407 vdd.n2406 185
R1105 vdd.n2408 vdd.n2407 185
R1106 vdd.n2405 vdd.n1060 185
R1107 vdd.n1060 vdd.n1057 185
R1108 vdd.n2404 vdd.n2403 185
R1109 vdd.n2403 vdd.n2402 185
R1110 vdd.n1062 vdd.n1061 185
R1111 vdd.n1063 vdd.n1062 185
R1112 vdd.n2395 vdd.n2394 185
R1113 vdd.n2396 vdd.n2395 185
R1114 vdd.n2393 vdd.n1072 185
R1115 vdd.n1072 vdd.n1069 185
R1116 vdd.n2392 vdd.n2391 185
R1117 vdd.n2391 vdd.n2390 185
R1118 vdd.n1074 vdd.n1073 185
R1119 vdd.n1075 vdd.n1074 185
R1120 vdd.n2383 vdd.n2382 185
R1121 vdd.n2384 vdd.n2383 185
R1122 vdd.n2381 vdd.n1084 185
R1123 vdd.n2380 vdd.n2379 185
R1124 vdd.n2377 vdd.n1085 185
R1125 vdd.n2377 vdd.n1081 185
R1126 vdd.n2376 vdd.n2375 185
R1127 vdd.n2374 vdd.n2373 185
R1128 vdd.n2372 vdd.n1087 185
R1129 vdd.n2370 vdd.n2369 185
R1130 vdd.n2368 vdd.n1088 185
R1131 vdd.n2367 vdd.n2366 185
R1132 vdd.n2364 vdd.n1089 185
R1133 vdd.n2362 vdd.n2361 185
R1134 vdd.n2360 vdd.n1090 185
R1135 vdd.n2359 vdd.n2358 185
R1136 vdd.n2356 vdd.n1091 185
R1137 vdd.n2354 vdd.n2353 185
R1138 vdd.n2352 vdd.n1092 185
R1139 vdd.n2351 vdd.n2350 185
R1140 vdd.n2348 vdd.n1093 185
R1141 vdd.n2346 vdd.n2345 185
R1142 vdd.n2344 vdd.n1094 185
R1143 vdd.n2343 vdd.n2342 185
R1144 vdd.n2340 vdd.n1095 185
R1145 vdd.n2338 vdd.n2337 185
R1146 vdd.n2336 vdd.n1096 185
R1147 vdd.n2335 vdd.n2334 185
R1148 vdd.n2332 vdd.n1097 185
R1149 vdd.n2330 vdd.n2329 185
R1150 vdd.n2328 vdd.n1098 185
R1151 vdd.n2327 vdd.n2326 185
R1152 vdd.n2324 vdd.n1099 185
R1153 vdd.n2322 vdd.n2321 185
R1154 vdd.n2320 vdd.n1100 185
R1155 vdd.n2318 vdd.n2317 185
R1156 vdd.n2315 vdd.n1103 185
R1157 vdd.n2313 vdd.n2312 185
R1158 vdd.n2574 vdd.n2573 185
R1159 vdd.n2576 vdd.n2575 185
R1160 vdd.n2578 vdd.n2577 185
R1161 vdd.n2581 vdd.n2580 185
R1162 vdd.n2583 vdd.n2582 185
R1163 vdd.n2585 vdd.n2584 185
R1164 vdd.n2587 vdd.n2586 185
R1165 vdd.n2589 vdd.n2588 185
R1166 vdd.n2591 vdd.n2590 185
R1167 vdd.n2593 vdd.n2592 185
R1168 vdd.n2595 vdd.n2594 185
R1169 vdd.n2597 vdd.n2596 185
R1170 vdd.n2599 vdd.n2598 185
R1171 vdd.n2601 vdd.n2600 185
R1172 vdd.n2603 vdd.n2602 185
R1173 vdd.n2605 vdd.n2604 185
R1174 vdd.n2607 vdd.n2606 185
R1175 vdd.n2609 vdd.n2608 185
R1176 vdd.n2611 vdd.n2610 185
R1177 vdd.n2613 vdd.n2612 185
R1178 vdd.n2615 vdd.n2614 185
R1179 vdd.n2617 vdd.n2616 185
R1180 vdd.n2619 vdd.n2618 185
R1181 vdd.n2621 vdd.n2620 185
R1182 vdd.n2623 vdd.n2622 185
R1183 vdd.n2625 vdd.n2624 185
R1184 vdd.n2627 vdd.n2626 185
R1185 vdd.n2629 vdd.n2628 185
R1186 vdd.n2631 vdd.n2630 185
R1187 vdd.n2633 vdd.n2632 185
R1188 vdd.n2635 vdd.n2634 185
R1189 vdd.n2637 vdd.n2636 185
R1190 vdd.n2639 vdd.n2638 185
R1191 vdd.n2640 vdd.n957 185
R1192 vdd.n2642 vdd.n2641 185
R1193 vdd.n2643 vdd.n2642 185
R1194 vdd.n2572 vdd.n961 185
R1195 vdd.n2572 vdd.n2571 185
R1196 vdd.n2249 vdd.n962 185
R1197 vdd.n963 vdd.n962 185
R1198 vdd.n2250 vdd.n973 185
R1199 vdd.n2496 vdd.n973 185
R1200 vdd.n2253 vdd.n2252 185
R1201 vdd.n2252 vdd.n2251 185
R1202 vdd.n2254 vdd.n980 185
R1203 vdd.n2489 vdd.n980 185
R1204 vdd.n2256 vdd.n2255 185
R1205 vdd.n2255 vdd.n979 185
R1206 vdd.n2257 vdd.n987 185
R1207 vdd.n2481 vdd.n987 185
R1208 vdd.n2259 vdd.n2258 185
R1209 vdd.n2258 vdd.n986 185
R1210 vdd.n2260 vdd.n992 185
R1211 vdd.n2475 vdd.n992 185
R1212 vdd.n2262 vdd.n2261 185
R1213 vdd.n2263 vdd.n2262 185
R1214 vdd.n2248 vdd.n997 185
R1215 vdd.n2469 vdd.n997 185
R1216 vdd.n2247 vdd.n2246 185
R1217 vdd.n2246 vdd.n1004 185
R1218 vdd.n2245 vdd.n1002 185
R1219 vdd.n2463 vdd.n1002 185
R1220 vdd.n2244 vdd.n2243 185
R1221 vdd.n2243 vdd.n1010 185
R1222 vdd.n1104 vdd.n1008 185
R1223 vdd.n2457 vdd.n1008 185
R1224 vdd.n2277 vdd.n2276 185
R1225 vdd.n2276 vdd.n2275 185
R1226 vdd.n2278 vdd.n1015 185
R1227 vdd.n2451 vdd.n1015 185
R1228 vdd.n2280 vdd.n2279 185
R1229 vdd.n2279 vdd.n1014 185
R1230 vdd.n2281 vdd.n1021 185
R1231 vdd.n2445 vdd.n1021 185
R1232 vdd.n2283 vdd.n2282 185
R1233 vdd.n2282 vdd.n1020 185
R1234 vdd.n2284 vdd.n1026 185
R1235 vdd.n2439 vdd.n1026 185
R1236 vdd.n2286 vdd.n2285 185
R1237 vdd.n2285 vdd.n1034 185
R1238 vdd.n2287 vdd.n1032 185
R1239 vdd.n2432 vdd.n1032 185
R1240 vdd.n2289 vdd.n2288 185
R1241 vdd.n2288 vdd.n1041 185
R1242 vdd.n2290 vdd.n1039 185
R1243 vdd.n2426 vdd.n1039 185
R1244 vdd.n2292 vdd.n2291 185
R1245 vdd.n2291 vdd.n1038 185
R1246 vdd.n2293 vdd.n1046 185
R1247 vdd.n2420 vdd.n1046 185
R1248 vdd.n2295 vdd.n2294 185
R1249 vdd.n2294 vdd.n1045 185
R1250 vdd.n2296 vdd.n1052 185
R1251 vdd.n2414 vdd.n1052 185
R1252 vdd.n2298 vdd.n2297 185
R1253 vdd.n2297 vdd.n1051 185
R1254 vdd.n2299 vdd.n1058 185
R1255 vdd.n2408 vdd.n1058 185
R1256 vdd.n2301 vdd.n2300 185
R1257 vdd.n2300 vdd.n1057 185
R1258 vdd.n2302 vdd.n1064 185
R1259 vdd.n2402 vdd.n1064 185
R1260 vdd.n2304 vdd.n2303 185
R1261 vdd.n2303 vdd.n1063 185
R1262 vdd.n2305 vdd.n1070 185
R1263 vdd.n2396 vdd.n1070 185
R1264 vdd.n2307 vdd.n2306 185
R1265 vdd.n2306 vdd.n1069 185
R1266 vdd.n2308 vdd.n1076 185
R1267 vdd.n2390 vdd.n1076 185
R1268 vdd.n2310 vdd.n2309 185
R1269 vdd.n2309 vdd.n1075 185
R1270 vdd.n2311 vdd.n1082 185
R1271 vdd.n2384 vdd.n1082 185
R1272 vdd.n370 vdd.n369 185
R1273 vdd.n3436 vdd.n370 185
R1274 vdd.n3439 vdd.n3438 185
R1275 vdd.n3438 vdd.n3437 185
R1276 vdd.n3440 vdd.n364 185
R1277 vdd.n364 vdd.n363 185
R1278 vdd.n3442 vdd.n3441 185
R1279 vdd.n3443 vdd.n3442 185
R1280 vdd.n359 vdd.n358 185
R1281 vdd.n3444 vdd.n359 185
R1282 vdd.n3447 vdd.n3446 185
R1283 vdd.n3446 vdd.n3445 185
R1284 vdd.n3448 vdd.n353 185
R1285 vdd.n3418 vdd.n353 185
R1286 vdd.n3450 vdd.n3449 185
R1287 vdd.n3451 vdd.n3450 185
R1288 vdd.n348 vdd.n347 185
R1289 vdd.n3452 vdd.n348 185
R1290 vdd.n3455 vdd.n3454 185
R1291 vdd.n3454 vdd.n3453 185
R1292 vdd.n3456 vdd.n342 185
R1293 vdd.n349 vdd.n342 185
R1294 vdd.n3458 vdd.n3457 185
R1295 vdd.n3459 vdd.n3458 185
R1296 vdd.n338 vdd.n337 185
R1297 vdd.n3460 vdd.n338 185
R1298 vdd.n3463 vdd.n3462 185
R1299 vdd.n3462 vdd.n3461 185
R1300 vdd.n3464 vdd.n333 185
R1301 vdd.n333 vdd.n332 185
R1302 vdd.n3466 vdd.n3465 185
R1303 vdd.n3467 vdd.n3466 185
R1304 vdd.n327 vdd.n325 185
R1305 vdd.n3468 vdd.n327 185
R1306 vdd.n3471 vdd.n3470 185
R1307 vdd.n3470 vdd.n3469 185
R1308 vdd.n326 vdd.n324 185
R1309 vdd.n328 vdd.n326 185
R1310 vdd.n3394 vdd.n3393 185
R1311 vdd.n3395 vdd.n3394 185
R1312 vdd.n615 vdd.n614 185
R1313 vdd.n614 vdd.n613 185
R1314 vdd.n3389 vdd.n3388 185
R1315 vdd.n3388 vdd.n3387 185
R1316 vdd.n618 vdd.n617 185
R1317 vdd.n624 vdd.n618 185
R1318 vdd.n3375 vdd.n3374 185
R1319 vdd.n3376 vdd.n3375 185
R1320 vdd.n626 vdd.n625 185
R1321 vdd.n3367 vdd.n625 185
R1322 vdd.n3370 vdd.n3369 185
R1323 vdd.n3369 vdd.n3368 185
R1324 vdd.n629 vdd.n628 185
R1325 vdd.n636 vdd.n629 185
R1326 vdd.n3358 vdd.n3357 185
R1327 vdd.n3359 vdd.n3358 185
R1328 vdd.n638 vdd.n637 185
R1329 vdd.n637 vdd.n635 185
R1330 vdd.n3353 vdd.n3352 185
R1331 vdd.n3352 vdd.n3351 185
R1332 vdd.n641 vdd.n640 185
R1333 vdd.n642 vdd.n641 185
R1334 vdd.n3342 vdd.n3341 185
R1335 vdd.n3343 vdd.n3342 185
R1336 vdd.n650 vdd.n649 185
R1337 vdd.n649 vdd.n648 185
R1338 vdd.n3337 vdd.n3336 185
R1339 vdd.n3336 vdd.n3335 185
R1340 vdd.n653 vdd.n652 185
R1341 vdd.n659 vdd.n653 185
R1342 vdd.n3326 vdd.n3325 185
R1343 vdd.n3327 vdd.n3326 185
R1344 vdd.n3322 vdd.n660 185
R1345 vdd.n3321 vdd.n3320 185
R1346 vdd.n3318 vdd.n662 185
R1347 vdd.n3318 vdd.n658 185
R1348 vdd.n3317 vdd.n3316 185
R1349 vdd.n3315 vdd.n3314 185
R1350 vdd.n3313 vdd.n3312 185
R1351 vdd.n3311 vdd.n3310 185
R1352 vdd.n3309 vdd.n668 185
R1353 vdd.n3307 vdd.n3306 185
R1354 vdd.n3305 vdd.n669 185
R1355 vdd.n3304 vdd.n3303 185
R1356 vdd.n3301 vdd.n674 185
R1357 vdd.n3299 vdd.n3298 185
R1358 vdd.n3297 vdd.n675 185
R1359 vdd.n3296 vdd.n3295 185
R1360 vdd.n3293 vdd.n680 185
R1361 vdd.n3291 vdd.n3290 185
R1362 vdd.n3289 vdd.n681 185
R1363 vdd.n3288 vdd.n3287 185
R1364 vdd.n3285 vdd.n688 185
R1365 vdd.n3283 vdd.n3282 185
R1366 vdd.n3281 vdd.n689 185
R1367 vdd.n3280 vdd.n3279 185
R1368 vdd.n3277 vdd.n694 185
R1369 vdd.n3275 vdd.n3274 185
R1370 vdd.n3273 vdd.n695 185
R1371 vdd.n3272 vdd.n3271 185
R1372 vdd.n3269 vdd.n700 185
R1373 vdd.n3267 vdd.n3266 185
R1374 vdd.n3265 vdd.n701 185
R1375 vdd.n3264 vdd.n3263 185
R1376 vdd.n3261 vdd.n706 185
R1377 vdd.n3259 vdd.n3258 185
R1378 vdd.n3257 vdd.n707 185
R1379 vdd.n3256 vdd.n3255 185
R1380 vdd.n3253 vdd.n712 185
R1381 vdd.n3251 vdd.n3250 185
R1382 vdd.n3249 vdd.n713 185
R1383 vdd.n3248 vdd.n3247 185
R1384 vdd.n3245 vdd.n718 185
R1385 vdd.n3243 vdd.n3242 185
R1386 vdd.n3241 vdd.n719 185
R1387 vdd.n728 vdd.n722 185
R1388 vdd.n3237 vdd.n3236 185
R1389 vdd.n3234 vdd.n726 185
R1390 vdd.n3233 vdd.n3232 185
R1391 vdd.n3231 vdd.n3230 185
R1392 vdd.n3229 vdd.n732 185
R1393 vdd.n3227 vdd.n3226 185
R1394 vdd.n3225 vdd.n733 185
R1395 vdd.n3224 vdd.n3223 185
R1396 vdd.n3221 vdd.n738 185
R1397 vdd.n3219 vdd.n3218 185
R1398 vdd.n3217 vdd.n739 185
R1399 vdd.n3216 vdd.n3215 185
R1400 vdd.n3213 vdd.n744 185
R1401 vdd.n3211 vdd.n3210 185
R1402 vdd.n3209 vdd.n745 185
R1403 vdd.n3208 vdd.n3207 185
R1404 vdd.n3205 vdd.n3204 185
R1405 vdd.n3203 vdd.n3202 185
R1406 vdd.n3201 vdd.n3200 185
R1407 vdd.n3199 vdd.n3198 185
R1408 vdd.n3194 vdd.n657 185
R1409 vdd.n658 vdd.n657 185
R1410 vdd.n3433 vdd.n3432 185
R1411 vdd.n599 vdd.n404 185
R1412 vdd.n598 vdd.n597 185
R1413 vdd.n596 vdd.n595 185
R1414 vdd.n594 vdd.n409 185
R1415 vdd.n590 vdd.n589 185
R1416 vdd.n588 vdd.n587 185
R1417 vdd.n586 vdd.n585 185
R1418 vdd.n584 vdd.n411 185
R1419 vdd.n580 vdd.n579 185
R1420 vdd.n578 vdd.n577 185
R1421 vdd.n576 vdd.n575 185
R1422 vdd.n574 vdd.n413 185
R1423 vdd.n570 vdd.n569 185
R1424 vdd.n568 vdd.n567 185
R1425 vdd.n566 vdd.n565 185
R1426 vdd.n564 vdd.n415 185
R1427 vdd.n560 vdd.n559 185
R1428 vdd.n558 vdd.n557 185
R1429 vdd.n556 vdd.n555 185
R1430 vdd.n554 vdd.n417 185
R1431 vdd.n550 vdd.n549 185
R1432 vdd.n548 vdd.n547 185
R1433 vdd.n546 vdd.n545 185
R1434 vdd.n544 vdd.n421 185
R1435 vdd.n540 vdd.n539 185
R1436 vdd.n538 vdd.n537 185
R1437 vdd.n536 vdd.n535 185
R1438 vdd.n534 vdd.n423 185
R1439 vdd.n530 vdd.n529 185
R1440 vdd.n528 vdd.n527 185
R1441 vdd.n526 vdd.n525 185
R1442 vdd.n524 vdd.n425 185
R1443 vdd.n520 vdd.n519 185
R1444 vdd.n518 vdd.n517 185
R1445 vdd.n516 vdd.n515 185
R1446 vdd.n514 vdd.n427 185
R1447 vdd.n510 vdd.n509 185
R1448 vdd.n508 vdd.n507 185
R1449 vdd.n506 vdd.n505 185
R1450 vdd.n504 vdd.n429 185
R1451 vdd.n500 vdd.n499 185
R1452 vdd.n498 vdd.n497 185
R1453 vdd.n496 vdd.n495 185
R1454 vdd.n494 vdd.n433 185
R1455 vdd.n490 vdd.n489 185
R1456 vdd.n488 vdd.n487 185
R1457 vdd.n486 vdd.n485 185
R1458 vdd.n484 vdd.n435 185
R1459 vdd.n480 vdd.n479 185
R1460 vdd.n478 vdd.n477 185
R1461 vdd.n476 vdd.n475 185
R1462 vdd.n474 vdd.n437 185
R1463 vdd.n470 vdd.n469 185
R1464 vdd.n468 vdd.n467 185
R1465 vdd.n466 vdd.n465 185
R1466 vdd.n464 vdd.n439 185
R1467 vdd.n460 vdd.n459 185
R1468 vdd.n458 vdd.n457 185
R1469 vdd.n456 vdd.n455 185
R1470 vdd.n454 vdd.n441 185
R1471 vdd.n450 vdd.n449 185
R1472 vdd.n448 vdd.n447 185
R1473 vdd.n446 vdd.n445 185
R1474 vdd.n3429 vdd.n372 185
R1475 vdd.n3436 vdd.n372 185
R1476 vdd.n3428 vdd.n371 185
R1477 vdd.n3437 vdd.n371 185
R1478 vdd.n3427 vdd.n3426 185
R1479 vdd.n3426 vdd.n363 185
R1480 vdd.n602 vdd.n362 185
R1481 vdd.n3443 vdd.n362 185
R1482 vdd.n3422 vdd.n361 185
R1483 vdd.n3444 vdd.n361 185
R1484 vdd.n3421 vdd.n360 185
R1485 vdd.n3445 vdd.n360 185
R1486 vdd.n3420 vdd.n3419 185
R1487 vdd.n3419 vdd.n3418 185
R1488 vdd.n604 vdd.n352 185
R1489 vdd.n3451 vdd.n352 185
R1490 vdd.n3414 vdd.n351 185
R1491 vdd.n3452 vdd.n351 185
R1492 vdd.n3413 vdd.n350 185
R1493 vdd.n3453 vdd.n350 185
R1494 vdd.n3412 vdd.n3411 185
R1495 vdd.n3411 vdd.n349 185
R1496 vdd.n606 vdd.n341 185
R1497 vdd.n3459 vdd.n341 185
R1498 vdd.n3407 vdd.n340 185
R1499 vdd.n3460 vdd.n340 185
R1500 vdd.n3406 vdd.n339 185
R1501 vdd.n3461 vdd.n339 185
R1502 vdd.n3405 vdd.n3404 185
R1503 vdd.n3404 vdd.n332 185
R1504 vdd.n608 vdd.n331 185
R1505 vdd.n3467 vdd.n331 185
R1506 vdd.n3400 vdd.n330 185
R1507 vdd.n3468 vdd.n330 185
R1508 vdd.n3399 vdd.n329 185
R1509 vdd.n3469 vdd.n329 185
R1510 vdd.n3398 vdd.n3397 185
R1511 vdd.n3397 vdd.n328 185
R1512 vdd.n3396 vdd.n610 185
R1513 vdd.n3396 vdd.n3395 185
R1514 vdd.n3384 vdd.n612 185
R1515 vdd.n613 vdd.n612 185
R1516 vdd.n3386 vdd.n3385 185
R1517 vdd.n3387 vdd.n3386 185
R1518 vdd.n620 vdd.n619 185
R1519 vdd.n624 vdd.n619 185
R1520 vdd.n3378 vdd.n3377 185
R1521 vdd.n3377 vdd.n3376 185
R1522 vdd.n623 vdd.n622 185
R1523 vdd.n3367 vdd.n623 185
R1524 vdd.n3366 vdd.n3365 185
R1525 vdd.n3368 vdd.n3366 185
R1526 vdd.n631 vdd.n630 185
R1527 vdd.n636 vdd.n630 185
R1528 vdd.n3361 vdd.n3360 185
R1529 vdd.n3360 vdd.n3359 185
R1530 vdd.n634 vdd.n633 185
R1531 vdd.n635 vdd.n634 185
R1532 vdd.n3350 vdd.n3349 185
R1533 vdd.n3351 vdd.n3350 185
R1534 vdd.n644 vdd.n643 185
R1535 vdd.n643 vdd.n642 185
R1536 vdd.n3345 vdd.n3344 185
R1537 vdd.n3344 vdd.n3343 185
R1538 vdd.n647 vdd.n646 185
R1539 vdd.n648 vdd.n647 185
R1540 vdd.n3334 vdd.n3333 185
R1541 vdd.n3335 vdd.n3334 185
R1542 vdd.n655 vdd.n654 185
R1543 vdd.n659 vdd.n654 185
R1544 vdd.n3329 vdd.n3328 185
R1545 vdd.n3328 vdd.n3327 185
R1546 vdd.n2931 vdd.n918 185
R1547 vdd.n2930 vdd.n2929 185
R1548 vdd.n920 vdd.n919 185
R1549 vdd.n2927 vdd.n920 185
R1550 vdd.n2750 vdd.n2749 185
R1551 vdd.n2752 vdd.n2751 185
R1552 vdd.n2754 vdd.n2753 185
R1553 vdd.n2756 vdd.n2755 185
R1554 vdd.n2758 vdd.n2757 185
R1555 vdd.n2760 vdd.n2759 185
R1556 vdd.n2762 vdd.n2761 185
R1557 vdd.n2764 vdd.n2763 185
R1558 vdd.n2766 vdd.n2765 185
R1559 vdd.n2768 vdd.n2767 185
R1560 vdd.n2770 vdd.n2769 185
R1561 vdd.n2772 vdd.n2771 185
R1562 vdd.n2774 vdd.n2773 185
R1563 vdd.n2776 vdd.n2775 185
R1564 vdd.n2778 vdd.n2777 185
R1565 vdd.n2780 vdd.n2779 185
R1566 vdd.n2782 vdd.n2781 185
R1567 vdd.n2784 vdd.n2783 185
R1568 vdd.n2786 vdd.n2785 185
R1569 vdd.n2788 vdd.n2787 185
R1570 vdd.n2790 vdd.n2789 185
R1571 vdd.n2792 vdd.n2791 185
R1572 vdd.n2794 vdd.n2793 185
R1573 vdd.n2796 vdd.n2795 185
R1574 vdd.n2798 vdd.n2797 185
R1575 vdd.n2800 vdd.n2799 185
R1576 vdd.n2802 vdd.n2801 185
R1577 vdd.n2804 vdd.n2803 185
R1578 vdd.n2806 vdd.n2805 185
R1579 vdd.n2809 vdd.n2808 185
R1580 vdd.n2811 vdd.n2810 185
R1581 vdd.n2813 vdd.n2812 185
R1582 vdd.n3095 vdd.n3094 185
R1583 vdd.n3096 vdd.n803 185
R1584 vdd.n3098 vdd.n3097 185
R1585 vdd.n3100 vdd.n801 185
R1586 vdd.n3102 vdd.n3101 185
R1587 vdd.n3103 vdd.n800 185
R1588 vdd.n3105 vdd.n3104 185
R1589 vdd.n3107 vdd.n798 185
R1590 vdd.n3109 vdd.n3108 185
R1591 vdd.n3110 vdd.n797 185
R1592 vdd.n3112 vdd.n3111 185
R1593 vdd.n3114 vdd.n795 185
R1594 vdd.n3116 vdd.n3115 185
R1595 vdd.n3117 vdd.n794 185
R1596 vdd.n3119 vdd.n3118 185
R1597 vdd.n3121 vdd.n792 185
R1598 vdd.n3123 vdd.n3122 185
R1599 vdd.n3125 vdd.n791 185
R1600 vdd.n3127 vdd.n3126 185
R1601 vdd.n3129 vdd.n789 185
R1602 vdd.n3131 vdd.n3130 185
R1603 vdd.n3132 vdd.n788 185
R1604 vdd.n3134 vdd.n3133 185
R1605 vdd.n3136 vdd.n786 185
R1606 vdd.n3138 vdd.n3137 185
R1607 vdd.n3139 vdd.n785 185
R1608 vdd.n3141 vdd.n3140 185
R1609 vdd.n3143 vdd.n783 185
R1610 vdd.n3145 vdd.n3144 185
R1611 vdd.n3146 vdd.n782 185
R1612 vdd.n3148 vdd.n3147 185
R1613 vdd.n3150 vdd.n781 185
R1614 vdd.n3151 vdd.n780 185
R1615 vdd.n3154 vdd.n3153 185
R1616 vdd.n3155 vdd.n778 185
R1617 vdd.n778 vdd.n756 185
R1618 vdd.n3092 vdd.n775 185
R1619 vdd.n3158 vdd.n775 185
R1620 vdd.n3091 vdd.n3090 185
R1621 vdd.n3090 vdd.n774 185
R1622 vdd.n3089 vdd.n807 185
R1623 vdd.n3089 vdd.n3088 185
R1624 vdd.n2863 vdd.n808 185
R1625 vdd.n817 vdd.n808 185
R1626 vdd.n2864 vdd.n815 185
R1627 vdd.n3082 vdd.n815 185
R1628 vdd.n2866 vdd.n2865 185
R1629 vdd.n2865 vdd.n814 185
R1630 vdd.n2867 vdd.n823 185
R1631 vdd.n3031 vdd.n823 185
R1632 vdd.n2869 vdd.n2868 185
R1633 vdd.n2868 vdd.n822 185
R1634 vdd.n2870 vdd.n828 185
R1635 vdd.n3025 vdd.n828 185
R1636 vdd.n2872 vdd.n2871 185
R1637 vdd.n2871 vdd.n835 185
R1638 vdd.n2873 vdd.n833 185
R1639 vdd.n3019 vdd.n833 185
R1640 vdd.n2875 vdd.n2874 185
R1641 vdd.n2874 vdd.n841 185
R1642 vdd.n2876 vdd.n839 185
R1643 vdd.n3013 vdd.n839 185
R1644 vdd.n2878 vdd.n2877 185
R1645 vdd.n2877 vdd.n848 185
R1646 vdd.n2879 vdd.n846 185
R1647 vdd.n3007 vdd.n846 185
R1648 vdd.n2881 vdd.n2880 185
R1649 vdd.n2880 vdd.n845 185
R1650 vdd.n2882 vdd.n853 185
R1651 vdd.n3001 vdd.n853 185
R1652 vdd.n2884 vdd.n2883 185
R1653 vdd.n2883 vdd.n852 185
R1654 vdd.n2885 vdd.n860 185
R1655 vdd.n2994 vdd.n860 185
R1656 vdd.n2887 vdd.n2886 185
R1657 vdd.n2886 vdd.n859 185
R1658 vdd.n2888 vdd.n865 185
R1659 vdd.n2988 vdd.n865 185
R1660 vdd.n2890 vdd.n2889 185
R1661 vdd.n2889 vdd.n872 185
R1662 vdd.n2891 vdd.n870 185
R1663 vdd.n2982 vdd.n870 185
R1664 vdd.n2893 vdd.n2892 185
R1665 vdd.n2894 vdd.n2893 185
R1666 vdd.n2862 vdd.n877 185
R1667 vdd.n2976 vdd.n877 185
R1668 vdd.n2861 vdd.n2860 185
R1669 vdd.n2860 vdd.n876 185
R1670 vdd.n2859 vdd.n883 185
R1671 vdd.n2970 vdd.n883 185
R1672 vdd.n2858 vdd.n2857 185
R1673 vdd.n2857 vdd.n882 185
R1674 vdd.n2818 vdd.n888 185
R1675 vdd.n2964 vdd.n888 185
R1676 vdd.n2908 vdd.n2907 185
R1677 vdd.n2907 vdd.n2906 185
R1678 vdd.n2909 vdd.n893 185
R1679 vdd.n2958 vdd.n893 185
R1680 vdd.n2911 vdd.n2910 185
R1681 vdd.n2910 vdd.n901 185
R1682 vdd.n2912 vdd.n899 185
R1683 vdd.n2952 vdd.n899 185
R1684 vdd.n2914 vdd.n2913 185
R1685 vdd.n2913 vdd.n898 185
R1686 vdd.n2915 vdd.n905 185
R1687 vdd.n2946 vdd.n905 185
R1688 vdd.n2917 vdd.n2916 185
R1689 vdd.n2918 vdd.n2917 185
R1690 vdd.n2817 vdd.n910 185
R1691 vdd.n2940 vdd.n910 185
R1692 vdd.n2816 vdd.n2815 185
R1693 vdd.n2815 vdd.n917 185
R1694 vdd.n2814 vdd.n915 185
R1695 vdd.n2934 vdd.n915 185
R1696 vdd.n2933 vdd.n2932 185
R1697 vdd.n2934 vdd.n2933 185
R1698 vdd.n909 vdd.n908 185
R1699 vdd.n917 vdd.n909 185
R1700 vdd.n2942 vdd.n2941 185
R1701 vdd.n2941 vdd.n2940 185
R1702 vdd.n2943 vdd.n907 185
R1703 vdd.n2918 vdd.n907 185
R1704 vdd.n2945 vdd.n2944 185
R1705 vdd.n2946 vdd.n2945 185
R1706 vdd.n897 vdd.n896 185
R1707 vdd.n898 vdd.n897 185
R1708 vdd.n2954 vdd.n2953 185
R1709 vdd.n2953 vdd.n2952 185
R1710 vdd.n2955 vdd.n895 185
R1711 vdd.n901 vdd.n895 185
R1712 vdd.n2957 vdd.n2956 185
R1713 vdd.n2958 vdd.n2957 185
R1714 vdd.n887 vdd.n886 185
R1715 vdd.n2906 vdd.n887 185
R1716 vdd.n2966 vdd.n2965 185
R1717 vdd.n2965 vdd.n2964 185
R1718 vdd.n2967 vdd.n885 185
R1719 vdd.n885 vdd.n882 185
R1720 vdd.n2969 vdd.n2968 185
R1721 vdd.n2970 vdd.n2969 185
R1722 vdd.n875 vdd.n874 185
R1723 vdd.n876 vdd.n875 185
R1724 vdd.n2978 vdd.n2977 185
R1725 vdd.n2977 vdd.n2976 185
R1726 vdd.n2979 vdd.n873 185
R1727 vdd.n2894 vdd.n873 185
R1728 vdd.n2981 vdd.n2980 185
R1729 vdd.n2982 vdd.n2981 185
R1730 vdd.n864 vdd.n863 185
R1731 vdd.n872 vdd.n864 185
R1732 vdd.n2990 vdd.n2989 185
R1733 vdd.n2989 vdd.n2988 185
R1734 vdd.n2991 vdd.n862 185
R1735 vdd.n862 vdd.n859 185
R1736 vdd.n2993 vdd.n2992 185
R1737 vdd.n2994 vdd.n2993 185
R1738 vdd.n851 vdd.n850 185
R1739 vdd.n852 vdd.n851 185
R1740 vdd.n3003 vdd.n3002 185
R1741 vdd.n3002 vdd.n3001 185
R1742 vdd.n3004 vdd.n849 185
R1743 vdd.n849 vdd.n845 185
R1744 vdd.n3006 vdd.n3005 185
R1745 vdd.n3007 vdd.n3006 185
R1746 vdd.n838 vdd.n837 185
R1747 vdd.n848 vdd.n838 185
R1748 vdd.n3015 vdd.n3014 185
R1749 vdd.n3014 vdd.n3013 185
R1750 vdd.n3016 vdd.n836 185
R1751 vdd.n841 vdd.n836 185
R1752 vdd.n3018 vdd.n3017 185
R1753 vdd.n3019 vdd.n3018 185
R1754 vdd.n827 vdd.n826 185
R1755 vdd.n835 vdd.n827 185
R1756 vdd.n3027 vdd.n3026 185
R1757 vdd.n3026 vdd.n3025 185
R1758 vdd.n3028 vdd.n825 185
R1759 vdd.n825 vdd.n822 185
R1760 vdd.n3030 vdd.n3029 185
R1761 vdd.n3031 vdd.n3030 185
R1762 vdd.n813 vdd.n812 185
R1763 vdd.n814 vdd.n813 185
R1764 vdd.n3084 vdd.n3083 185
R1765 vdd.n3083 vdd.n3082 185
R1766 vdd.n3085 vdd.n811 185
R1767 vdd.n817 vdd.n811 185
R1768 vdd.n3087 vdd.n3086 185
R1769 vdd.n3088 vdd.n3087 185
R1770 vdd.n779 vdd.n777 185
R1771 vdd.n777 vdd.n774 185
R1772 vdd.n3157 vdd.n3156 185
R1773 vdd.n3158 vdd.n3157 185
R1774 vdd.n2570 vdd.n2569 185
R1775 vdd.n2571 vdd.n2570 185
R1776 vdd.n967 vdd.n965 185
R1777 vdd.n965 vdd.n963 185
R1778 vdd.n2485 vdd.n974 185
R1779 vdd.n2496 vdd.n974 185
R1780 vdd.n2486 vdd.n983 185
R1781 vdd.n2251 vdd.n983 185
R1782 vdd.n2488 vdd.n2487 185
R1783 vdd.n2489 vdd.n2488 185
R1784 vdd.n2484 vdd.n982 185
R1785 vdd.n982 vdd.n979 185
R1786 vdd.n2483 vdd.n2482 185
R1787 vdd.n2482 vdd.n2481 185
R1788 vdd.n985 vdd.n984 185
R1789 vdd.n986 vdd.n985 185
R1790 vdd.n2474 vdd.n2473 185
R1791 vdd.n2475 vdd.n2474 185
R1792 vdd.n2472 vdd.n994 185
R1793 vdd.n2263 vdd.n994 185
R1794 vdd.n2471 vdd.n2470 185
R1795 vdd.n2470 vdd.n2469 185
R1796 vdd.n996 vdd.n995 185
R1797 vdd.n1004 vdd.n996 185
R1798 vdd.n2462 vdd.n2461 185
R1799 vdd.n2463 vdd.n2462 185
R1800 vdd.n2460 vdd.n1005 185
R1801 vdd.n1010 vdd.n1005 185
R1802 vdd.n2459 vdd.n2458 185
R1803 vdd.n2458 vdd.n2457 185
R1804 vdd.n1007 vdd.n1006 185
R1805 vdd.n2275 vdd.n1007 185
R1806 vdd.n2450 vdd.n2449 185
R1807 vdd.n2451 vdd.n2450 185
R1808 vdd.n2448 vdd.n1017 185
R1809 vdd.n1017 vdd.n1014 185
R1810 vdd.n2447 vdd.n2446 185
R1811 vdd.n2446 vdd.n2445 185
R1812 vdd.n1019 vdd.n1018 185
R1813 vdd.n1020 vdd.n1019 185
R1814 vdd.n2438 vdd.n2437 185
R1815 vdd.n2439 vdd.n2438 185
R1816 vdd.n2435 vdd.n1028 185
R1817 vdd.n1034 vdd.n1028 185
R1818 vdd.n2434 vdd.n2433 185
R1819 vdd.n2433 vdd.n2432 185
R1820 vdd.n1031 vdd.n1030 185
R1821 vdd.n1041 vdd.n1031 185
R1822 vdd.n2425 vdd.n2424 185
R1823 vdd.n2426 vdd.n2425 185
R1824 vdd.n2423 vdd.n1042 185
R1825 vdd.n1042 vdd.n1038 185
R1826 vdd.n2422 vdd.n2421 185
R1827 vdd.n2421 vdd.n2420 185
R1828 vdd.n1044 vdd.n1043 185
R1829 vdd.n1045 vdd.n1044 185
R1830 vdd.n2413 vdd.n2412 185
R1831 vdd.n2414 vdd.n2413 185
R1832 vdd.n2411 vdd.n1054 185
R1833 vdd.n1054 vdd.n1051 185
R1834 vdd.n2410 vdd.n2409 185
R1835 vdd.n2409 vdd.n2408 185
R1836 vdd.n1056 vdd.n1055 185
R1837 vdd.n1057 vdd.n1056 185
R1838 vdd.n2401 vdd.n2400 185
R1839 vdd.n2402 vdd.n2401 185
R1840 vdd.n2399 vdd.n1066 185
R1841 vdd.n1066 vdd.n1063 185
R1842 vdd.n2398 vdd.n2397 185
R1843 vdd.n2397 vdd.n2396 185
R1844 vdd.n1068 vdd.n1067 185
R1845 vdd.n1069 vdd.n1068 185
R1846 vdd.n2389 vdd.n2388 185
R1847 vdd.n2390 vdd.n2389 185
R1848 vdd.n2387 vdd.n1078 185
R1849 vdd.n1078 vdd.n1075 185
R1850 vdd.n2386 vdd.n2385 185
R1851 vdd.n2385 vdd.n2384 185
R1852 vdd.n2501 vdd.n938 185
R1853 vdd.n2643 vdd.n938 185
R1854 vdd.n2503 vdd.n2502 185
R1855 vdd.n2505 vdd.n2504 185
R1856 vdd.n2507 vdd.n2506 185
R1857 vdd.n2509 vdd.n2508 185
R1858 vdd.n2511 vdd.n2510 185
R1859 vdd.n2513 vdd.n2512 185
R1860 vdd.n2515 vdd.n2514 185
R1861 vdd.n2517 vdd.n2516 185
R1862 vdd.n2519 vdd.n2518 185
R1863 vdd.n2521 vdd.n2520 185
R1864 vdd.n2523 vdd.n2522 185
R1865 vdd.n2525 vdd.n2524 185
R1866 vdd.n2527 vdd.n2526 185
R1867 vdd.n2529 vdd.n2528 185
R1868 vdd.n2531 vdd.n2530 185
R1869 vdd.n2533 vdd.n2532 185
R1870 vdd.n2535 vdd.n2534 185
R1871 vdd.n2537 vdd.n2536 185
R1872 vdd.n2539 vdd.n2538 185
R1873 vdd.n2541 vdd.n2540 185
R1874 vdd.n2543 vdd.n2542 185
R1875 vdd.n2545 vdd.n2544 185
R1876 vdd.n2547 vdd.n2546 185
R1877 vdd.n2549 vdd.n2548 185
R1878 vdd.n2551 vdd.n2550 185
R1879 vdd.n2553 vdd.n2552 185
R1880 vdd.n2555 vdd.n2554 185
R1881 vdd.n2557 vdd.n2556 185
R1882 vdd.n2559 vdd.n2558 185
R1883 vdd.n2561 vdd.n2560 185
R1884 vdd.n2563 vdd.n2562 185
R1885 vdd.n2565 vdd.n2564 185
R1886 vdd.n2567 vdd.n2566 185
R1887 vdd.n2568 vdd.n966 185
R1888 vdd.n2500 vdd.n964 185
R1889 vdd.n2571 vdd.n964 185
R1890 vdd.n2499 vdd.n2498 185
R1891 vdd.n2498 vdd.n963 185
R1892 vdd.n2497 vdd.n971 185
R1893 vdd.n2497 vdd.n2496 185
R1894 vdd.n2235 vdd.n972 185
R1895 vdd.n2251 vdd.n972 185
R1896 vdd.n2236 vdd.n981 185
R1897 vdd.n2489 vdd.n981 185
R1898 vdd.n2238 vdd.n2237 185
R1899 vdd.n2237 vdd.n979 185
R1900 vdd.n2239 vdd.n988 185
R1901 vdd.n2481 vdd.n988 185
R1902 vdd.n2241 vdd.n2240 185
R1903 vdd.n2240 vdd.n986 185
R1904 vdd.n2242 vdd.n993 185
R1905 vdd.n2475 vdd.n993 185
R1906 vdd.n2265 vdd.n2264 185
R1907 vdd.n2264 vdd.n2263 185
R1908 vdd.n2266 vdd.n998 185
R1909 vdd.n2469 vdd.n998 185
R1910 vdd.n2268 vdd.n2267 185
R1911 vdd.n2267 vdd.n1004 185
R1912 vdd.n2269 vdd.n1003 185
R1913 vdd.n2463 vdd.n1003 185
R1914 vdd.n2271 vdd.n2270 185
R1915 vdd.n2270 vdd.n1010 185
R1916 vdd.n2272 vdd.n1009 185
R1917 vdd.n2457 vdd.n1009 185
R1918 vdd.n2274 vdd.n2273 185
R1919 vdd.n2275 vdd.n2274 185
R1920 vdd.n2234 vdd.n1016 185
R1921 vdd.n2451 vdd.n1016 185
R1922 vdd.n2233 vdd.n2232 185
R1923 vdd.n2232 vdd.n1014 185
R1924 vdd.n2231 vdd.n1022 185
R1925 vdd.n2445 vdd.n1022 185
R1926 vdd.n2230 vdd.n2229 185
R1927 vdd.n2229 vdd.n1020 185
R1928 vdd.n2228 vdd.n1027 185
R1929 vdd.n2439 vdd.n1027 185
R1930 vdd.n2227 vdd.n2226 185
R1931 vdd.n2226 vdd.n1034 185
R1932 vdd.n2225 vdd.n1033 185
R1933 vdd.n2432 vdd.n1033 185
R1934 vdd.n2224 vdd.n2223 185
R1935 vdd.n2223 vdd.n1041 185
R1936 vdd.n2222 vdd.n1040 185
R1937 vdd.n2426 vdd.n1040 185
R1938 vdd.n2221 vdd.n2220 185
R1939 vdd.n2220 vdd.n1038 185
R1940 vdd.n2219 vdd.n1047 185
R1941 vdd.n2420 vdd.n1047 185
R1942 vdd.n2218 vdd.n2217 185
R1943 vdd.n2217 vdd.n1045 185
R1944 vdd.n2216 vdd.n1053 185
R1945 vdd.n2414 vdd.n1053 185
R1946 vdd.n2215 vdd.n2214 185
R1947 vdd.n2214 vdd.n1051 185
R1948 vdd.n2213 vdd.n1059 185
R1949 vdd.n2408 vdd.n1059 185
R1950 vdd.n2212 vdd.n2211 185
R1951 vdd.n2211 vdd.n1057 185
R1952 vdd.n2210 vdd.n1065 185
R1953 vdd.n2402 vdd.n1065 185
R1954 vdd.n2209 vdd.n2208 185
R1955 vdd.n2208 vdd.n1063 185
R1956 vdd.n2207 vdd.n1071 185
R1957 vdd.n2396 vdd.n1071 185
R1958 vdd.n2206 vdd.n2205 185
R1959 vdd.n2205 vdd.n1069 185
R1960 vdd.n2204 vdd.n1077 185
R1961 vdd.n2390 vdd.n1077 185
R1962 vdd.n2203 vdd.n2202 185
R1963 vdd.n2202 vdd.n1075 185
R1964 vdd.n2201 vdd.n1083 185
R1965 vdd.n2384 vdd.n1083 185
R1966 vdd.n1080 vdd.n1079 185
R1967 vdd.n2133 vdd.n2131 185
R1968 vdd.n2136 vdd.n2135 185
R1969 vdd.n2137 vdd.n2130 185
R1970 vdd.n2139 vdd.n2138 185
R1971 vdd.n2141 vdd.n2129 185
R1972 vdd.n2144 vdd.n2143 185
R1973 vdd.n2145 vdd.n2128 185
R1974 vdd.n2147 vdd.n2146 185
R1975 vdd.n2149 vdd.n2127 185
R1976 vdd.n2152 vdd.n2151 185
R1977 vdd.n2153 vdd.n2126 185
R1978 vdd.n2155 vdd.n2154 185
R1979 vdd.n2157 vdd.n2125 185
R1980 vdd.n2160 vdd.n2159 185
R1981 vdd.n2161 vdd.n2124 185
R1982 vdd.n2163 vdd.n2162 185
R1983 vdd.n2165 vdd.n2123 185
R1984 vdd.n2168 vdd.n2167 185
R1985 vdd.n2169 vdd.n1114 185
R1986 vdd.n2171 vdd.n2170 185
R1987 vdd.n2173 vdd.n1113 185
R1988 vdd.n2176 vdd.n2175 185
R1989 vdd.n2177 vdd.n1112 185
R1990 vdd.n2179 vdd.n2178 185
R1991 vdd.n2181 vdd.n1111 185
R1992 vdd.n2184 vdd.n2183 185
R1993 vdd.n2185 vdd.n1110 185
R1994 vdd.n2187 vdd.n2186 185
R1995 vdd.n2189 vdd.n1109 185
R1996 vdd.n2192 vdd.n2191 185
R1997 vdd.n2193 vdd.n1106 185
R1998 vdd.n2196 vdd.n2195 185
R1999 vdd.n2198 vdd.n1105 185
R2000 vdd.n2200 vdd.n2199 185
R2001 vdd.n2199 vdd.n1081 185
R2002 vdd.n315 vdd.n314 171.744
R2003 vdd.n314 vdd.n313 171.744
R2004 vdd.n313 vdd.n282 171.744
R2005 vdd.n306 vdd.n282 171.744
R2006 vdd.n306 vdd.n305 171.744
R2007 vdd.n305 vdd.n287 171.744
R2008 vdd.n298 vdd.n287 171.744
R2009 vdd.n298 vdd.n297 171.744
R2010 vdd.n297 vdd.n291 171.744
R2011 vdd.n260 vdd.n259 171.744
R2012 vdd.n259 vdd.n258 171.744
R2013 vdd.n258 vdd.n227 171.744
R2014 vdd.n251 vdd.n227 171.744
R2015 vdd.n251 vdd.n250 171.744
R2016 vdd.n250 vdd.n232 171.744
R2017 vdd.n243 vdd.n232 171.744
R2018 vdd.n243 vdd.n242 171.744
R2019 vdd.n242 vdd.n236 171.744
R2020 vdd.n217 vdd.n216 171.744
R2021 vdd.n216 vdd.n215 171.744
R2022 vdd.n215 vdd.n184 171.744
R2023 vdd.n208 vdd.n184 171.744
R2024 vdd.n208 vdd.n207 171.744
R2025 vdd.n207 vdd.n189 171.744
R2026 vdd.n200 vdd.n189 171.744
R2027 vdd.n200 vdd.n199 171.744
R2028 vdd.n199 vdd.n193 171.744
R2029 vdd.n162 vdd.n161 171.744
R2030 vdd.n161 vdd.n160 171.744
R2031 vdd.n160 vdd.n129 171.744
R2032 vdd.n153 vdd.n129 171.744
R2033 vdd.n153 vdd.n152 171.744
R2034 vdd.n152 vdd.n134 171.744
R2035 vdd.n145 vdd.n134 171.744
R2036 vdd.n145 vdd.n144 171.744
R2037 vdd.n144 vdd.n138 171.744
R2038 vdd.n120 vdd.n119 171.744
R2039 vdd.n119 vdd.n118 171.744
R2040 vdd.n118 vdd.n87 171.744
R2041 vdd.n111 vdd.n87 171.744
R2042 vdd.n111 vdd.n110 171.744
R2043 vdd.n110 vdd.n92 171.744
R2044 vdd.n103 vdd.n92 171.744
R2045 vdd.n103 vdd.n102 171.744
R2046 vdd.n102 vdd.n96 171.744
R2047 vdd.n65 vdd.n64 171.744
R2048 vdd.n64 vdd.n63 171.744
R2049 vdd.n63 vdd.n32 171.744
R2050 vdd.n56 vdd.n32 171.744
R2051 vdd.n56 vdd.n55 171.744
R2052 vdd.n55 vdd.n37 171.744
R2053 vdd.n48 vdd.n37 171.744
R2054 vdd.n48 vdd.n47 171.744
R2055 vdd.n47 vdd.n41 171.744
R2056 vdd.n1764 vdd.n1763 171.744
R2057 vdd.n1763 vdd.n1762 171.744
R2058 vdd.n1762 vdd.n1731 171.744
R2059 vdd.n1755 vdd.n1731 171.744
R2060 vdd.n1755 vdd.n1754 171.744
R2061 vdd.n1754 vdd.n1736 171.744
R2062 vdd.n1747 vdd.n1736 171.744
R2063 vdd.n1747 vdd.n1746 171.744
R2064 vdd.n1746 vdd.n1740 171.744
R2065 vdd.n1819 vdd.n1818 171.744
R2066 vdd.n1818 vdd.n1817 171.744
R2067 vdd.n1817 vdd.n1786 171.744
R2068 vdd.n1810 vdd.n1786 171.744
R2069 vdd.n1810 vdd.n1809 171.744
R2070 vdd.n1809 vdd.n1791 171.744
R2071 vdd.n1802 vdd.n1791 171.744
R2072 vdd.n1802 vdd.n1801 171.744
R2073 vdd.n1801 vdd.n1795 171.744
R2074 vdd.n1666 vdd.n1665 171.744
R2075 vdd.n1665 vdd.n1664 171.744
R2076 vdd.n1664 vdd.n1633 171.744
R2077 vdd.n1657 vdd.n1633 171.744
R2078 vdd.n1657 vdd.n1656 171.744
R2079 vdd.n1656 vdd.n1638 171.744
R2080 vdd.n1649 vdd.n1638 171.744
R2081 vdd.n1649 vdd.n1648 171.744
R2082 vdd.n1648 vdd.n1642 171.744
R2083 vdd.n1721 vdd.n1720 171.744
R2084 vdd.n1720 vdd.n1719 171.744
R2085 vdd.n1719 vdd.n1688 171.744
R2086 vdd.n1712 vdd.n1688 171.744
R2087 vdd.n1712 vdd.n1711 171.744
R2088 vdd.n1711 vdd.n1693 171.744
R2089 vdd.n1704 vdd.n1693 171.744
R2090 vdd.n1704 vdd.n1703 171.744
R2091 vdd.n1703 vdd.n1697 171.744
R2092 vdd.n1569 vdd.n1568 171.744
R2093 vdd.n1568 vdd.n1567 171.744
R2094 vdd.n1567 vdd.n1536 171.744
R2095 vdd.n1560 vdd.n1536 171.744
R2096 vdd.n1560 vdd.n1559 171.744
R2097 vdd.n1559 vdd.n1541 171.744
R2098 vdd.n1552 vdd.n1541 171.744
R2099 vdd.n1552 vdd.n1551 171.744
R2100 vdd.n1551 vdd.n1545 171.744
R2101 vdd.n1624 vdd.n1623 171.744
R2102 vdd.n1623 vdd.n1622 171.744
R2103 vdd.n1622 vdd.n1591 171.744
R2104 vdd.n1615 vdd.n1591 171.744
R2105 vdd.n1615 vdd.n1614 171.744
R2106 vdd.n1614 vdd.n1596 171.744
R2107 vdd.n1607 vdd.n1596 171.744
R2108 vdd.n1607 vdd.n1606 171.744
R2109 vdd.n1606 vdd.n1600 171.744
R2110 vdd.n449 vdd.n448 146.341
R2111 vdd.n455 vdd.n454 146.341
R2112 vdd.n459 vdd.n458 146.341
R2113 vdd.n465 vdd.n464 146.341
R2114 vdd.n469 vdd.n468 146.341
R2115 vdd.n475 vdd.n474 146.341
R2116 vdd.n479 vdd.n478 146.341
R2117 vdd.n485 vdd.n484 146.341
R2118 vdd.n489 vdd.n488 146.341
R2119 vdd.n495 vdd.n494 146.341
R2120 vdd.n499 vdd.n498 146.341
R2121 vdd.n505 vdd.n504 146.341
R2122 vdd.n509 vdd.n508 146.341
R2123 vdd.n515 vdd.n514 146.341
R2124 vdd.n519 vdd.n518 146.341
R2125 vdd.n525 vdd.n524 146.341
R2126 vdd.n529 vdd.n528 146.341
R2127 vdd.n535 vdd.n534 146.341
R2128 vdd.n539 vdd.n538 146.341
R2129 vdd.n545 vdd.n544 146.341
R2130 vdd.n549 vdd.n548 146.341
R2131 vdd.n555 vdd.n554 146.341
R2132 vdd.n559 vdd.n558 146.341
R2133 vdd.n565 vdd.n564 146.341
R2134 vdd.n569 vdd.n568 146.341
R2135 vdd.n575 vdd.n574 146.341
R2136 vdd.n579 vdd.n578 146.341
R2137 vdd.n585 vdd.n584 146.341
R2138 vdd.n589 vdd.n588 146.341
R2139 vdd.n595 vdd.n594 146.341
R2140 vdd.n597 vdd.n404 146.341
R2141 vdd.n3328 vdd.n654 146.341
R2142 vdd.n3334 vdd.n654 146.341
R2143 vdd.n3334 vdd.n647 146.341
R2144 vdd.n3344 vdd.n647 146.341
R2145 vdd.n3344 vdd.n643 146.341
R2146 vdd.n3350 vdd.n643 146.341
R2147 vdd.n3350 vdd.n634 146.341
R2148 vdd.n3360 vdd.n634 146.341
R2149 vdd.n3360 vdd.n630 146.341
R2150 vdd.n3366 vdd.n630 146.341
R2151 vdd.n3366 vdd.n623 146.341
R2152 vdd.n3377 vdd.n623 146.341
R2153 vdd.n3377 vdd.n619 146.341
R2154 vdd.n3386 vdd.n619 146.341
R2155 vdd.n3386 vdd.n612 146.341
R2156 vdd.n3396 vdd.n612 146.341
R2157 vdd.n3397 vdd.n3396 146.341
R2158 vdd.n3397 vdd.n329 146.341
R2159 vdd.n330 vdd.n329 146.341
R2160 vdd.n331 vdd.n330 146.341
R2161 vdd.n3404 vdd.n331 146.341
R2162 vdd.n3404 vdd.n339 146.341
R2163 vdd.n340 vdd.n339 146.341
R2164 vdd.n341 vdd.n340 146.341
R2165 vdd.n3411 vdd.n341 146.341
R2166 vdd.n3411 vdd.n350 146.341
R2167 vdd.n351 vdd.n350 146.341
R2168 vdd.n352 vdd.n351 146.341
R2169 vdd.n3419 vdd.n352 146.341
R2170 vdd.n3419 vdd.n360 146.341
R2171 vdd.n361 vdd.n360 146.341
R2172 vdd.n362 vdd.n361 146.341
R2173 vdd.n3426 vdd.n362 146.341
R2174 vdd.n3426 vdd.n371 146.341
R2175 vdd.n372 vdd.n371 146.341
R2176 vdd.n3320 vdd.n3318 146.341
R2177 vdd.n3318 vdd.n3317 146.341
R2178 vdd.n3314 vdd.n3313 146.341
R2179 vdd.n3310 vdd.n3309 146.341
R2180 vdd.n3307 vdd.n669 146.341
R2181 vdd.n3303 vdd.n3301 146.341
R2182 vdd.n3299 vdd.n675 146.341
R2183 vdd.n3295 vdd.n3293 146.341
R2184 vdd.n3291 vdd.n681 146.341
R2185 vdd.n3287 vdd.n3285 146.341
R2186 vdd.n3283 vdd.n689 146.341
R2187 vdd.n3279 vdd.n3277 146.341
R2188 vdd.n3275 vdd.n695 146.341
R2189 vdd.n3271 vdd.n3269 146.341
R2190 vdd.n3267 vdd.n701 146.341
R2191 vdd.n3263 vdd.n3261 146.341
R2192 vdd.n3259 vdd.n707 146.341
R2193 vdd.n3255 vdd.n3253 146.341
R2194 vdd.n3251 vdd.n713 146.341
R2195 vdd.n3247 vdd.n3245 146.341
R2196 vdd.n3243 vdd.n719 146.341
R2197 vdd.n3236 vdd.n728 146.341
R2198 vdd.n3234 vdd.n3233 146.341
R2199 vdd.n3230 vdd.n3229 146.341
R2200 vdd.n3227 vdd.n733 146.341
R2201 vdd.n3223 vdd.n3221 146.341
R2202 vdd.n3219 vdd.n739 146.341
R2203 vdd.n3215 vdd.n3213 146.341
R2204 vdd.n3211 vdd.n745 146.341
R2205 vdd.n3207 vdd.n3205 146.341
R2206 vdd.n3202 vdd.n3201 146.341
R2207 vdd.n3198 vdd.n657 146.341
R2208 vdd.n3326 vdd.n653 146.341
R2209 vdd.n3336 vdd.n653 146.341
R2210 vdd.n3336 vdd.n649 146.341
R2211 vdd.n3342 vdd.n649 146.341
R2212 vdd.n3342 vdd.n641 146.341
R2213 vdd.n3352 vdd.n641 146.341
R2214 vdd.n3352 vdd.n637 146.341
R2215 vdd.n3358 vdd.n637 146.341
R2216 vdd.n3358 vdd.n629 146.341
R2217 vdd.n3369 vdd.n629 146.341
R2218 vdd.n3369 vdd.n625 146.341
R2219 vdd.n3375 vdd.n625 146.341
R2220 vdd.n3375 vdd.n618 146.341
R2221 vdd.n3388 vdd.n618 146.341
R2222 vdd.n3388 vdd.n614 146.341
R2223 vdd.n3394 vdd.n614 146.341
R2224 vdd.n3394 vdd.n326 146.341
R2225 vdd.n3470 vdd.n326 146.341
R2226 vdd.n3470 vdd.n327 146.341
R2227 vdd.n3466 vdd.n327 146.341
R2228 vdd.n3466 vdd.n333 146.341
R2229 vdd.n3462 vdd.n333 146.341
R2230 vdd.n3462 vdd.n338 146.341
R2231 vdd.n3458 vdd.n338 146.341
R2232 vdd.n3458 vdd.n342 146.341
R2233 vdd.n3454 vdd.n342 146.341
R2234 vdd.n3454 vdd.n348 146.341
R2235 vdd.n3450 vdd.n348 146.341
R2236 vdd.n3450 vdd.n353 146.341
R2237 vdd.n3446 vdd.n353 146.341
R2238 vdd.n3446 vdd.n359 146.341
R2239 vdd.n3442 vdd.n359 146.341
R2240 vdd.n3442 vdd.n364 146.341
R2241 vdd.n3438 vdd.n364 146.341
R2242 vdd.n3438 vdd.n370 146.341
R2243 vdd.n2106 vdd.n2105 146.341
R2244 vdd.n2103 vdd.n1900 146.341
R2245 vdd.n2096 vdd.n1906 146.341
R2246 vdd.n2094 vdd.n2093 146.341
R2247 vdd.n2091 vdd.n1908 146.341
R2248 vdd.n2087 vdd.n2086 146.341
R2249 vdd.n2084 vdd.n1915 146.341
R2250 vdd.n2080 vdd.n2079 146.341
R2251 vdd.n2077 vdd.n1922 146.341
R2252 vdd.n1933 vdd.n1930 146.341
R2253 vdd.n2069 vdd.n2068 146.341
R2254 vdd.n2066 vdd.n1935 146.341
R2255 vdd.n2062 vdd.n2061 146.341
R2256 vdd.n2059 vdd.n1941 146.341
R2257 vdd.n2055 vdd.n2054 146.341
R2258 vdd.n2052 vdd.n1948 146.341
R2259 vdd.n2048 vdd.n2047 146.341
R2260 vdd.n2045 vdd.n1955 146.341
R2261 vdd.n2041 vdd.n2040 146.341
R2262 vdd.n2038 vdd.n1962 146.341
R2263 vdd.n1973 vdd.n1970 146.341
R2264 vdd.n2030 vdd.n2029 146.341
R2265 vdd.n2027 vdd.n1975 146.341
R2266 vdd.n2023 vdd.n2022 146.341
R2267 vdd.n2020 vdd.n1981 146.341
R2268 vdd.n2016 vdd.n2015 146.341
R2269 vdd.n2013 vdd.n1988 146.341
R2270 vdd.n2009 vdd.n2008 146.341
R2271 vdd.n2006 vdd.n2003 146.341
R2272 vdd.n2001 vdd.n1998 146.341
R2273 vdd.n1996 vdd.n1120 146.341
R2274 vdd.n1461 vdd.n1225 146.341
R2275 vdd.n1461 vdd.n1217 146.341
R2276 vdd.n1471 vdd.n1217 146.341
R2277 vdd.n1471 vdd.n1213 146.341
R2278 vdd.n1477 vdd.n1213 146.341
R2279 vdd.n1477 vdd.n1205 146.341
R2280 vdd.n1488 vdd.n1205 146.341
R2281 vdd.n1488 vdd.n1201 146.341
R2282 vdd.n1494 vdd.n1201 146.341
R2283 vdd.n1494 vdd.n1195 146.341
R2284 vdd.n1505 vdd.n1195 146.341
R2285 vdd.n1505 vdd.n1191 146.341
R2286 vdd.n1511 vdd.n1191 146.341
R2287 vdd.n1511 vdd.n1182 146.341
R2288 vdd.n1521 vdd.n1182 146.341
R2289 vdd.n1521 vdd.n1178 146.341
R2290 vdd.n1527 vdd.n1178 146.341
R2291 vdd.n1527 vdd.n1171 146.341
R2292 vdd.n1833 vdd.n1171 146.341
R2293 vdd.n1833 vdd.n1167 146.341
R2294 vdd.n1839 vdd.n1167 146.341
R2295 vdd.n1839 vdd.n1160 146.341
R2296 vdd.n1849 vdd.n1160 146.341
R2297 vdd.n1849 vdd.n1156 146.341
R2298 vdd.n1855 vdd.n1156 146.341
R2299 vdd.n1855 vdd.n1148 146.341
R2300 vdd.n1866 vdd.n1148 146.341
R2301 vdd.n1866 vdd.n1144 146.341
R2302 vdd.n1872 vdd.n1144 146.341
R2303 vdd.n1872 vdd.n1138 146.341
R2304 vdd.n1883 vdd.n1138 146.341
R2305 vdd.n1883 vdd.n1133 146.341
R2306 vdd.n1891 vdd.n1133 146.341
R2307 vdd.n1891 vdd.n1122 146.341
R2308 vdd.n2114 vdd.n1122 146.341
R2309 vdd.n1263 vdd.n1262 146.341
R2310 vdd.n1267 vdd.n1262 146.341
R2311 vdd.n1269 vdd.n1268 146.341
R2312 vdd.n1273 vdd.n1272 146.341
R2313 vdd.n1275 vdd.n1274 146.341
R2314 vdd.n1279 vdd.n1278 146.341
R2315 vdd.n1281 vdd.n1280 146.341
R2316 vdd.n1285 vdd.n1284 146.341
R2317 vdd.n1287 vdd.n1286 146.341
R2318 vdd.n1419 vdd.n1418 146.341
R2319 vdd.n1291 vdd.n1290 146.341
R2320 vdd.n1295 vdd.n1294 146.341
R2321 vdd.n1297 vdd.n1296 146.341
R2322 vdd.n1301 vdd.n1300 146.341
R2323 vdd.n1303 vdd.n1302 146.341
R2324 vdd.n1307 vdd.n1306 146.341
R2325 vdd.n1309 vdd.n1308 146.341
R2326 vdd.n1313 vdd.n1312 146.341
R2327 vdd.n1315 vdd.n1314 146.341
R2328 vdd.n1319 vdd.n1318 146.341
R2329 vdd.n1383 vdd.n1320 146.341
R2330 vdd.n1324 vdd.n1323 146.341
R2331 vdd.n1326 vdd.n1325 146.341
R2332 vdd.n1330 vdd.n1329 146.341
R2333 vdd.n1332 vdd.n1331 146.341
R2334 vdd.n1336 vdd.n1335 146.341
R2335 vdd.n1338 vdd.n1337 146.341
R2336 vdd.n1342 vdd.n1341 146.341
R2337 vdd.n1344 vdd.n1343 146.341
R2338 vdd.n1348 vdd.n1347 146.341
R2339 vdd.n1350 vdd.n1349 146.341
R2340 vdd.n1455 vdd.n1231 146.341
R2341 vdd.n1463 vdd.n1223 146.341
R2342 vdd.n1463 vdd.n1219 146.341
R2343 vdd.n1469 vdd.n1219 146.341
R2344 vdd.n1469 vdd.n1211 146.341
R2345 vdd.n1480 vdd.n1211 146.341
R2346 vdd.n1480 vdd.n1207 146.341
R2347 vdd.n1486 vdd.n1207 146.341
R2348 vdd.n1486 vdd.n1200 146.341
R2349 vdd.n1497 vdd.n1200 146.341
R2350 vdd.n1497 vdd.n1196 146.341
R2351 vdd.n1503 vdd.n1196 146.341
R2352 vdd.n1503 vdd.n1189 146.341
R2353 vdd.n1513 vdd.n1189 146.341
R2354 vdd.n1513 vdd.n1185 146.341
R2355 vdd.n1519 vdd.n1185 146.341
R2356 vdd.n1519 vdd.n1177 146.341
R2357 vdd.n1530 vdd.n1177 146.341
R2358 vdd.n1530 vdd.n1173 146.341
R2359 vdd.n1831 vdd.n1173 146.341
R2360 vdd.n1831 vdd.n1166 146.341
R2361 vdd.n1841 vdd.n1166 146.341
R2362 vdd.n1841 vdd.n1162 146.341
R2363 vdd.n1847 vdd.n1162 146.341
R2364 vdd.n1847 vdd.n1154 146.341
R2365 vdd.n1858 vdd.n1154 146.341
R2366 vdd.n1858 vdd.n1150 146.341
R2367 vdd.n1864 vdd.n1150 146.341
R2368 vdd.n1864 vdd.n1143 146.341
R2369 vdd.n1875 vdd.n1143 146.341
R2370 vdd.n1875 vdd.n1139 146.341
R2371 vdd.n1881 vdd.n1139 146.341
R2372 vdd.n1881 vdd.n1131 146.341
R2373 vdd.n1893 vdd.n1131 146.341
R2374 vdd.n1893 vdd.n1126 146.341
R2375 vdd.n2112 vdd.n1126 146.341
R2376 vdd.n1107 vdd.t36 127.284
R2377 vdd.n968 vdd.t73 127.284
R2378 vdd.n1101 vdd.t100 127.284
R2379 vdd.n959 vdd.t96 127.284
R2380 vdd.n856 vdd.t46 127.284
R2381 vdd.n856 vdd.t47 127.284
R2382 vdd.n2678 vdd.t91 127.284
R2383 vdd.n804 vdd.t66 127.284
R2384 vdd.n2747 vdd.t78 127.284
R2385 vdd.n768 vdd.t31 127.284
R2386 vdd.n1029 vdd.t87 127.284
R2387 vdd.n1029 vdd.t88 127.284
R2388 vdd.n22 vdd.n20 117.314
R2389 vdd.n17 vdd.n15 117.314
R2390 vdd.n27 vdd.n26 116.927
R2391 vdd.n24 vdd.n23 116.927
R2392 vdd.n22 vdd.n21 116.927
R2393 vdd.n17 vdd.n16 116.927
R2394 vdd.n19 vdd.n18 116.927
R2395 vdd.n27 vdd.n25 116.927
R2396 vdd.n1108 vdd.t35 111.188
R2397 vdd.n969 vdd.t74 111.188
R2398 vdd.n1102 vdd.t99 111.188
R2399 vdd.n960 vdd.t97 111.188
R2400 vdd.n2679 vdd.t90 111.188
R2401 vdd.n805 vdd.t67 111.188
R2402 vdd.n2748 vdd.t77 111.188
R2403 vdd.n769 vdd.t32 111.188
R2404 vdd.n2933 vdd.n909 99.5127
R2405 vdd.n2941 vdd.n909 99.5127
R2406 vdd.n2941 vdd.n907 99.5127
R2407 vdd.n2945 vdd.n907 99.5127
R2408 vdd.n2945 vdd.n897 99.5127
R2409 vdd.n2953 vdd.n897 99.5127
R2410 vdd.n2953 vdd.n895 99.5127
R2411 vdd.n2957 vdd.n895 99.5127
R2412 vdd.n2957 vdd.n887 99.5127
R2413 vdd.n2965 vdd.n887 99.5127
R2414 vdd.n2965 vdd.n885 99.5127
R2415 vdd.n2969 vdd.n885 99.5127
R2416 vdd.n2969 vdd.n875 99.5127
R2417 vdd.n2977 vdd.n875 99.5127
R2418 vdd.n2977 vdd.n873 99.5127
R2419 vdd.n2981 vdd.n873 99.5127
R2420 vdd.n2981 vdd.n864 99.5127
R2421 vdd.n2989 vdd.n864 99.5127
R2422 vdd.n2989 vdd.n862 99.5127
R2423 vdd.n2993 vdd.n862 99.5127
R2424 vdd.n2993 vdd.n851 99.5127
R2425 vdd.n3002 vdd.n851 99.5127
R2426 vdd.n3002 vdd.n849 99.5127
R2427 vdd.n3006 vdd.n849 99.5127
R2428 vdd.n3006 vdd.n838 99.5127
R2429 vdd.n3014 vdd.n838 99.5127
R2430 vdd.n3014 vdd.n836 99.5127
R2431 vdd.n3018 vdd.n836 99.5127
R2432 vdd.n3018 vdd.n827 99.5127
R2433 vdd.n3026 vdd.n827 99.5127
R2434 vdd.n3026 vdd.n825 99.5127
R2435 vdd.n3030 vdd.n825 99.5127
R2436 vdd.n3030 vdd.n813 99.5127
R2437 vdd.n3083 vdd.n813 99.5127
R2438 vdd.n3083 vdd.n811 99.5127
R2439 vdd.n3087 vdd.n811 99.5127
R2440 vdd.n3087 vdd.n777 99.5127
R2441 vdd.n3157 vdd.n777 99.5127
R2442 vdd.n3153 vdd.n778 99.5127
R2443 vdd.n3151 vdd.n3150 99.5127
R2444 vdd.n3148 vdd.n782 99.5127
R2445 vdd.n3144 vdd.n3143 99.5127
R2446 vdd.n3141 vdd.n785 99.5127
R2447 vdd.n3137 vdd.n3136 99.5127
R2448 vdd.n3134 vdd.n788 99.5127
R2449 vdd.n3130 vdd.n3129 99.5127
R2450 vdd.n3127 vdd.n791 99.5127
R2451 vdd.n3122 vdd.n3121 99.5127
R2452 vdd.n3119 vdd.n794 99.5127
R2453 vdd.n3115 vdd.n3114 99.5127
R2454 vdd.n3112 vdd.n797 99.5127
R2455 vdd.n3108 vdd.n3107 99.5127
R2456 vdd.n3105 vdd.n800 99.5127
R2457 vdd.n3101 vdd.n3100 99.5127
R2458 vdd.n3098 vdd.n803 99.5127
R2459 vdd.n2815 vdd.n915 99.5127
R2460 vdd.n2815 vdd.n910 99.5127
R2461 vdd.n2917 vdd.n910 99.5127
R2462 vdd.n2917 vdd.n905 99.5127
R2463 vdd.n2913 vdd.n905 99.5127
R2464 vdd.n2913 vdd.n899 99.5127
R2465 vdd.n2910 vdd.n899 99.5127
R2466 vdd.n2910 vdd.n893 99.5127
R2467 vdd.n2907 vdd.n893 99.5127
R2468 vdd.n2907 vdd.n888 99.5127
R2469 vdd.n2857 vdd.n888 99.5127
R2470 vdd.n2857 vdd.n883 99.5127
R2471 vdd.n2860 vdd.n883 99.5127
R2472 vdd.n2860 vdd.n877 99.5127
R2473 vdd.n2893 vdd.n877 99.5127
R2474 vdd.n2893 vdd.n870 99.5127
R2475 vdd.n2889 vdd.n870 99.5127
R2476 vdd.n2889 vdd.n865 99.5127
R2477 vdd.n2886 vdd.n865 99.5127
R2478 vdd.n2886 vdd.n860 99.5127
R2479 vdd.n2883 vdd.n860 99.5127
R2480 vdd.n2883 vdd.n853 99.5127
R2481 vdd.n2880 vdd.n853 99.5127
R2482 vdd.n2880 vdd.n846 99.5127
R2483 vdd.n2877 vdd.n846 99.5127
R2484 vdd.n2877 vdd.n839 99.5127
R2485 vdd.n2874 vdd.n839 99.5127
R2486 vdd.n2874 vdd.n833 99.5127
R2487 vdd.n2871 vdd.n833 99.5127
R2488 vdd.n2871 vdd.n828 99.5127
R2489 vdd.n2868 vdd.n828 99.5127
R2490 vdd.n2868 vdd.n823 99.5127
R2491 vdd.n2865 vdd.n823 99.5127
R2492 vdd.n2865 vdd.n815 99.5127
R2493 vdd.n815 vdd.n808 99.5127
R2494 vdd.n3089 vdd.n808 99.5127
R2495 vdd.n3090 vdd.n3089 99.5127
R2496 vdd.n3090 vdd.n775 99.5127
R2497 vdd.n2929 vdd.n920 99.5127
R2498 vdd.n2749 vdd.n920 99.5127
R2499 vdd.n2753 vdd.n2752 99.5127
R2500 vdd.n2757 vdd.n2756 99.5127
R2501 vdd.n2761 vdd.n2760 99.5127
R2502 vdd.n2765 vdd.n2764 99.5127
R2503 vdd.n2769 vdd.n2768 99.5127
R2504 vdd.n2773 vdd.n2772 99.5127
R2505 vdd.n2777 vdd.n2776 99.5127
R2506 vdd.n2781 vdd.n2780 99.5127
R2507 vdd.n2785 vdd.n2784 99.5127
R2508 vdd.n2789 vdd.n2788 99.5127
R2509 vdd.n2793 vdd.n2792 99.5127
R2510 vdd.n2797 vdd.n2796 99.5127
R2511 vdd.n2801 vdd.n2800 99.5127
R2512 vdd.n2805 vdd.n2804 99.5127
R2513 vdd.n2810 vdd.n2809 99.5127
R2514 vdd.n2642 vdd.n957 99.5127
R2515 vdd.n2638 vdd.n2637 99.5127
R2516 vdd.n2634 vdd.n2633 99.5127
R2517 vdd.n2630 vdd.n2629 99.5127
R2518 vdd.n2626 vdd.n2625 99.5127
R2519 vdd.n2622 vdd.n2621 99.5127
R2520 vdd.n2618 vdd.n2617 99.5127
R2521 vdd.n2614 vdd.n2613 99.5127
R2522 vdd.n2610 vdd.n2609 99.5127
R2523 vdd.n2606 vdd.n2605 99.5127
R2524 vdd.n2602 vdd.n2601 99.5127
R2525 vdd.n2598 vdd.n2597 99.5127
R2526 vdd.n2594 vdd.n2593 99.5127
R2527 vdd.n2590 vdd.n2589 99.5127
R2528 vdd.n2586 vdd.n2585 99.5127
R2529 vdd.n2582 vdd.n2581 99.5127
R2530 vdd.n2577 vdd.n2576 99.5127
R2531 vdd.n2309 vdd.n1082 99.5127
R2532 vdd.n2309 vdd.n1076 99.5127
R2533 vdd.n2306 vdd.n1076 99.5127
R2534 vdd.n2306 vdd.n1070 99.5127
R2535 vdd.n2303 vdd.n1070 99.5127
R2536 vdd.n2303 vdd.n1064 99.5127
R2537 vdd.n2300 vdd.n1064 99.5127
R2538 vdd.n2300 vdd.n1058 99.5127
R2539 vdd.n2297 vdd.n1058 99.5127
R2540 vdd.n2297 vdd.n1052 99.5127
R2541 vdd.n2294 vdd.n1052 99.5127
R2542 vdd.n2294 vdd.n1046 99.5127
R2543 vdd.n2291 vdd.n1046 99.5127
R2544 vdd.n2291 vdd.n1039 99.5127
R2545 vdd.n2288 vdd.n1039 99.5127
R2546 vdd.n2288 vdd.n1032 99.5127
R2547 vdd.n2285 vdd.n1032 99.5127
R2548 vdd.n2285 vdd.n1026 99.5127
R2549 vdd.n2282 vdd.n1026 99.5127
R2550 vdd.n2282 vdd.n1021 99.5127
R2551 vdd.n2279 vdd.n1021 99.5127
R2552 vdd.n2279 vdd.n1015 99.5127
R2553 vdd.n2276 vdd.n1015 99.5127
R2554 vdd.n2276 vdd.n1008 99.5127
R2555 vdd.n2243 vdd.n1008 99.5127
R2556 vdd.n2243 vdd.n1002 99.5127
R2557 vdd.n2246 vdd.n1002 99.5127
R2558 vdd.n2246 vdd.n997 99.5127
R2559 vdd.n2262 vdd.n997 99.5127
R2560 vdd.n2262 vdd.n992 99.5127
R2561 vdd.n2258 vdd.n992 99.5127
R2562 vdd.n2258 vdd.n987 99.5127
R2563 vdd.n2255 vdd.n987 99.5127
R2564 vdd.n2255 vdd.n980 99.5127
R2565 vdd.n2252 vdd.n980 99.5127
R2566 vdd.n2252 vdd.n973 99.5127
R2567 vdd.n973 vdd.n962 99.5127
R2568 vdd.n2572 vdd.n962 99.5127
R2569 vdd.n2379 vdd.n2377 99.5127
R2570 vdd.n2377 vdd.n2376 99.5127
R2571 vdd.n2373 vdd.n2372 99.5127
R2572 vdd.n2370 vdd.n1088 99.5127
R2573 vdd.n2366 vdd.n2364 99.5127
R2574 vdd.n2362 vdd.n1090 99.5127
R2575 vdd.n2358 vdd.n2356 99.5127
R2576 vdd.n2354 vdd.n1092 99.5127
R2577 vdd.n2350 vdd.n2348 99.5127
R2578 vdd.n2346 vdd.n1094 99.5127
R2579 vdd.n2342 vdd.n2340 99.5127
R2580 vdd.n2338 vdd.n1096 99.5127
R2581 vdd.n2334 vdd.n2332 99.5127
R2582 vdd.n2330 vdd.n1098 99.5127
R2583 vdd.n2326 vdd.n2324 99.5127
R2584 vdd.n2322 vdd.n1100 99.5127
R2585 vdd.n2317 vdd.n2315 99.5127
R2586 vdd.n2383 vdd.n1074 99.5127
R2587 vdd.n2391 vdd.n1074 99.5127
R2588 vdd.n2391 vdd.n1072 99.5127
R2589 vdd.n2395 vdd.n1072 99.5127
R2590 vdd.n2395 vdd.n1062 99.5127
R2591 vdd.n2403 vdd.n1062 99.5127
R2592 vdd.n2403 vdd.n1060 99.5127
R2593 vdd.n2407 vdd.n1060 99.5127
R2594 vdd.n2407 vdd.n1050 99.5127
R2595 vdd.n2415 vdd.n1050 99.5127
R2596 vdd.n2415 vdd.n1048 99.5127
R2597 vdd.n2419 vdd.n1048 99.5127
R2598 vdd.n2419 vdd.n1037 99.5127
R2599 vdd.n2427 vdd.n1037 99.5127
R2600 vdd.n2427 vdd.n1035 99.5127
R2601 vdd.n2431 vdd.n1035 99.5127
R2602 vdd.n2431 vdd.n1025 99.5127
R2603 vdd.n2440 vdd.n1025 99.5127
R2604 vdd.n2440 vdd.n1023 99.5127
R2605 vdd.n2444 vdd.n1023 99.5127
R2606 vdd.n2444 vdd.n1013 99.5127
R2607 vdd.n2452 vdd.n1013 99.5127
R2608 vdd.n2452 vdd.n1011 99.5127
R2609 vdd.n2456 vdd.n1011 99.5127
R2610 vdd.n2456 vdd.n1001 99.5127
R2611 vdd.n2464 vdd.n1001 99.5127
R2612 vdd.n2464 vdd.n999 99.5127
R2613 vdd.n2468 vdd.n999 99.5127
R2614 vdd.n2468 vdd.n991 99.5127
R2615 vdd.n2476 vdd.n991 99.5127
R2616 vdd.n2476 vdd.n989 99.5127
R2617 vdd.n2480 vdd.n989 99.5127
R2618 vdd.n2480 vdd.n978 99.5127
R2619 vdd.n2490 vdd.n978 99.5127
R2620 vdd.n2490 vdd.n975 99.5127
R2621 vdd.n2495 vdd.n975 99.5127
R2622 vdd.n2495 vdd.n976 99.5127
R2623 vdd.n976 vdd.n956 99.5127
R2624 vdd.n3073 vdd.n3072 99.5127
R2625 vdd.n3070 vdd.n3036 99.5127
R2626 vdd.n3066 vdd.n3065 99.5127
R2627 vdd.n3063 vdd.n3039 99.5127
R2628 vdd.n3059 vdd.n3058 99.5127
R2629 vdd.n3056 vdd.n3042 99.5127
R2630 vdd.n3052 vdd.n3051 99.5127
R2631 vdd.n3049 vdd.n3046 99.5127
R2632 vdd.n3190 vdd.n755 99.5127
R2633 vdd.n3188 vdd.n3187 99.5127
R2634 vdd.n3185 vdd.n758 99.5127
R2635 vdd.n3181 vdd.n3180 99.5127
R2636 vdd.n3178 vdd.n761 99.5127
R2637 vdd.n3174 vdd.n3173 99.5127
R2638 vdd.n3171 vdd.n764 99.5127
R2639 vdd.n3167 vdd.n3166 99.5127
R2640 vdd.n3164 vdd.n767 99.5127
R2641 vdd.n2922 vdd.n916 99.5127
R2642 vdd.n2922 vdd.n911 99.5127
R2643 vdd.n2919 vdd.n911 99.5127
R2644 vdd.n2919 vdd.n906 99.5127
R2645 vdd.n2819 vdd.n906 99.5127
R2646 vdd.n2819 vdd.n900 99.5127
R2647 vdd.n2822 vdd.n900 99.5127
R2648 vdd.n2822 vdd.n894 99.5127
R2649 vdd.n2905 vdd.n894 99.5127
R2650 vdd.n2905 vdd.n889 99.5127
R2651 vdd.n2901 vdd.n889 99.5127
R2652 vdd.n2901 vdd.n884 99.5127
R2653 vdd.n2898 vdd.n884 99.5127
R2654 vdd.n2898 vdd.n878 99.5127
R2655 vdd.n2895 vdd.n878 99.5127
R2656 vdd.n2895 vdd.n871 99.5127
R2657 vdd.n2854 vdd.n871 99.5127
R2658 vdd.n2854 vdd.n866 99.5127
R2659 vdd.n2851 vdd.n866 99.5127
R2660 vdd.n2851 vdd.n861 99.5127
R2661 vdd.n2848 vdd.n861 99.5127
R2662 vdd.n2848 vdd.n854 99.5127
R2663 vdd.n2845 vdd.n854 99.5127
R2664 vdd.n2845 vdd.n847 99.5127
R2665 vdd.n2842 vdd.n847 99.5127
R2666 vdd.n2842 vdd.n840 99.5127
R2667 vdd.n2839 vdd.n840 99.5127
R2668 vdd.n2839 vdd.n834 99.5127
R2669 vdd.n2836 vdd.n834 99.5127
R2670 vdd.n2836 vdd.n829 99.5127
R2671 vdd.n2833 vdd.n829 99.5127
R2672 vdd.n2833 vdd.n824 99.5127
R2673 vdd.n2830 vdd.n824 99.5127
R2674 vdd.n2830 vdd.n816 99.5127
R2675 vdd.n2827 vdd.n816 99.5127
R2676 vdd.n2827 vdd.n809 99.5127
R2677 vdd.n809 vdd.n773 99.5127
R2678 vdd.n3159 vdd.n773 99.5127
R2679 vdd.n2683 vdd.n2682 99.5127
R2680 vdd.n2687 vdd.n2686 99.5127
R2681 vdd.n2691 vdd.n2690 99.5127
R2682 vdd.n2695 vdd.n2694 99.5127
R2683 vdd.n2699 vdd.n2698 99.5127
R2684 vdd.n2703 vdd.n2702 99.5127
R2685 vdd.n2707 vdd.n2706 99.5127
R2686 vdd.n2711 vdd.n2710 99.5127
R2687 vdd.n2715 vdd.n2714 99.5127
R2688 vdd.n2719 vdd.n2718 99.5127
R2689 vdd.n2723 vdd.n2722 99.5127
R2690 vdd.n2727 vdd.n2726 99.5127
R2691 vdd.n2731 vdd.n2730 99.5127
R2692 vdd.n2735 vdd.n2734 99.5127
R2693 vdd.n2739 vdd.n2738 99.5127
R2694 vdd.n2743 vdd.n2742 99.5127
R2695 vdd.n2926 vdd.n2677 99.5127
R2696 vdd.n2935 vdd.n912 99.5127
R2697 vdd.n2939 vdd.n912 99.5127
R2698 vdd.n2939 vdd.n904 99.5127
R2699 vdd.n2947 vdd.n904 99.5127
R2700 vdd.n2947 vdd.n902 99.5127
R2701 vdd.n2951 vdd.n902 99.5127
R2702 vdd.n2951 vdd.n892 99.5127
R2703 vdd.n2959 vdd.n892 99.5127
R2704 vdd.n2959 vdd.n890 99.5127
R2705 vdd.n2963 vdd.n890 99.5127
R2706 vdd.n2963 vdd.n881 99.5127
R2707 vdd.n2971 vdd.n881 99.5127
R2708 vdd.n2971 vdd.n879 99.5127
R2709 vdd.n2975 vdd.n879 99.5127
R2710 vdd.n2975 vdd.n869 99.5127
R2711 vdd.n2983 vdd.n869 99.5127
R2712 vdd.n2983 vdd.n867 99.5127
R2713 vdd.n2987 vdd.n867 99.5127
R2714 vdd.n2987 vdd.n858 99.5127
R2715 vdd.n2995 vdd.n858 99.5127
R2716 vdd.n2995 vdd.n855 99.5127
R2717 vdd.n3000 vdd.n855 99.5127
R2718 vdd.n3000 vdd.n844 99.5127
R2719 vdd.n3008 vdd.n844 99.5127
R2720 vdd.n3008 vdd.n842 99.5127
R2721 vdd.n3012 vdd.n842 99.5127
R2722 vdd.n3012 vdd.n832 99.5127
R2723 vdd.n3020 vdd.n832 99.5127
R2724 vdd.n3020 vdd.n830 99.5127
R2725 vdd.n3024 vdd.n830 99.5127
R2726 vdd.n3024 vdd.n821 99.5127
R2727 vdd.n3032 vdd.n821 99.5127
R2728 vdd.n3032 vdd.n818 99.5127
R2729 vdd.n3081 vdd.n818 99.5127
R2730 vdd.n3081 vdd.n819 99.5127
R2731 vdd.n819 vdd.n810 99.5127
R2732 vdd.n3076 vdd.n810 99.5127
R2733 vdd.n3076 vdd.n776 99.5127
R2734 vdd.n2566 vdd.n2565 99.5127
R2735 vdd.n2562 vdd.n2561 99.5127
R2736 vdd.n2558 vdd.n2557 99.5127
R2737 vdd.n2554 vdd.n2553 99.5127
R2738 vdd.n2550 vdd.n2549 99.5127
R2739 vdd.n2546 vdd.n2545 99.5127
R2740 vdd.n2542 vdd.n2541 99.5127
R2741 vdd.n2538 vdd.n2537 99.5127
R2742 vdd.n2534 vdd.n2533 99.5127
R2743 vdd.n2530 vdd.n2529 99.5127
R2744 vdd.n2526 vdd.n2525 99.5127
R2745 vdd.n2522 vdd.n2521 99.5127
R2746 vdd.n2518 vdd.n2517 99.5127
R2747 vdd.n2514 vdd.n2513 99.5127
R2748 vdd.n2510 vdd.n2509 99.5127
R2749 vdd.n2506 vdd.n2505 99.5127
R2750 vdd.n2502 vdd.n938 99.5127
R2751 vdd.n2202 vdd.n1083 99.5127
R2752 vdd.n2202 vdd.n1077 99.5127
R2753 vdd.n2205 vdd.n1077 99.5127
R2754 vdd.n2205 vdd.n1071 99.5127
R2755 vdd.n2208 vdd.n1071 99.5127
R2756 vdd.n2208 vdd.n1065 99.5127
R2757 vdd.n2211 vdd.n1065 99.5127
R2758 vdd.n2211 vdd.n1059 99.5127
R2759 vdd.n2214 vdd.n1059 99.5127
R2760 vdd.n2214 vdd.n1053 99.5127
R2761 vdd.n2217 vdd.n1053 99.5127
R2762 vdd.n2217 vdd.n1047 99.5127
R2763 vdd.n2220 vdd.n1047 99.5127
R2764 vdd.n2220 vdd.n1040 99.5127
R2765 vdd.n2223 vdd.n1040 99.5127
R2766 vdd.n2223 vdd.n1033 99.5127
R2767 vdd.n2226 vdd.n1033 99.5127
R2768 vdd.n2226 vdd.n1027 99.5127
R2769 vdd.n2229 vdd.n1027 99.5127
R2770 vdd.n2229 vdd.n1022 99.5127
R2771 vdd.n2232 vdd.n1022 99.5127
R2772 vdd.n2232 vdd.n1016 99.5127
R2773 vdd.n2274 vdd.n1016 99.5127
R2774 vdd.n2274 vdd.n1009 99.5127
R2775 vdd.n2270 vdd.n1009 99.5127
R2776 vdd.n2270 vdd.n1003 99.5127
R2777 vdd.n2267 vdd.n1003 99.5127
R2778 vdd.n2267 vdd.n998 99.5127
R2779 vdd.n2264 vdd.n998 99.5127
R2780 vdd.n2264 vdd.n993 99.5127
R2781 vdd.n2240 vdd.n993 99.5127
R2782 vdd.n2240 vdd.n988 99.5127
R2783 vdd.n2237 vdd.n988 99.5127
R2784 vdd.n2237 vdd.n981 99.5127
R2785 vdd.n981 vdd.n972 99.5127
R2786 vdd.n2497 vdd.n972 99.5127
R2787 vdd.n2498 vdd.n2497 99.5127
R2788 vdd.n2498 vdd.n964 99.5127
R2789 vdd.n2135 vdd.n2133 99.5127
R2790 vdd.n2139 vdd.n2130 99.5127
R2791 vdd.n2143 vdd.n2141 99.5127
R2792 vdd.n2147 vdd.n2128 99.5127
R2793 vdd.n2151 vdd.n2149 99.5127
R2794 vdd.n2155 vdd.n2126 99.5127
R2795 vdd.n2159 vdd.n2157 99.5127
R2796 vdd.n2163 vdd.n2124 99.5127
R2797 vdd.n2167 vdd.n2165 99.5127
R2798 vdd.n2171 vdd.n1114 99.5127
R2799 vdd.n2175 vdd.n2173 99.5127
R2800 vdd.n2179 vdd.n1112 99.5127
R2801 vdd.n2183 vdd.n2181 99.5127
R2802 vdd.n2187 vdd.n1110 99.5127
R2803 vdd.n2191 vdd.n2189 99.5127
R2804 vdd.n2196 vdd.n1106 99.5127
R2805 vdd.n2199 vdd.n2198 99.5127
R2806 vdd.n2385 vdd.n1078 99.5127
R2807 vdd.n2389 vdd.n1078 99.5127
R2808 vdd.n2389 vdd.n1068 99.5127
R2809 vdd.n2397 vdd.n1068 99.5127
R2810 vdd.n2397 vdd.n1066 99.5127
R2811 vdd.n2401 vdd.n1066 99.5127
R2812 vdd.n2401 vdd.n1056 99.5127
R2813 vdd.n2409 vdd.n1056 99.5127
R2814 vdd.n2409 vdd.n1054 99.5127
R2815 vdd.n2413 vdd.n1054 99.5127
R2816 vdd.n2413 vdd.n1044 99.5127
R2817 vdd.n2421 vdd.n1044 99.5127
R2818 vdd.n2421 vdd.n1042 99.5127
R2819 vdd.n2425 vdd.n1042 99.5127
R2820 vdd.n2425 vdd.n1031 99.5127
R2821 vdd.n2433 vdd.n1031 99.5127
R2822 vdd.n2433 vdd.n1028 99.5127
R2823 vdd.n2438 vdd.n1028 99.5127
R2824 vdd.n2438 vdd.n1019 99.5127
R2825 vdd.n2446 vdd.n1019 99.5127
R2826 vdd.n2446 vdd.n1017 99.5127
R2827 vdd.n2450 vdd.n1017 99.5127
R2828 vdd.n2450 vdd.n1007 99.5127
R2829 vdd.n2458 vdd.n1007 99.5127
R2830 vdd.n2458 vdd.n1005 99.5127
R2831 vdd.n2462 vdd.n1005 99.5127
R2832 vdd.n2462 vdd.n996 99.5127
R2833 vdd.n2470 vdd.n996 99.5127
R2834 vdd.n2470 vdd.n994 99.5127
R2835 vdd.n2474 vdd.n994 99.5127
R2836 vdd.n2474 vdd.n985 99.5127
R2837 vdd.n2482 vdd.n985 99.5127
R2838 vdd.n2482 vdd.n982 99.5127
R2839 vdd.n2488 vdd.n982 99.5127
R2840 vdd.n2488 vdd.n983 99.5127
R2841 vdd.n983 vdd.n974 99.5127
R2842 vdd.n974 vdd.n965 99.5127
R2843 vdd.n2570 vdd.n965 99.5127
R2844 vdd.n9 vdd.n7 98.9633
R2845 vdd.n2 vdd.n0 98.9633
R2846 vdd.n9 vdd.n8 98.6055
R2847 vdd.n11 vdd.n10 98.6055
R2848 vdd.n13 vdd.n12 98.6055
R2849 vdd.n6 vdd.n5 98.6055
R2850 vdd.n4 vdd.n3 98.6055
R2851 vdd.n2 vdd.n1 98.6055
R2852 vdd.t246 vdd.n291 85.8723
R2853 vdd.t267 vdd.n236 85.8723
R2854 vdd.t211 vdd.n193 85.8723
R2855 vdd.t227 vdd.n138 85.8723
R2856 vdd.t225 vdd.n96 85.8723
R2857 vdd.t216 vdd.n41 85.8723
R2858 vdd.t235 vdd.n1740 85.8723
R2859 vdd.t201 vdd.n1795 85.8723
R2860 vdd.t249 vdd.n1642 85.8723
R2861 vdd.t22 vdd.n1697 85.8723
R2862 vdd.t239 vdd.n1545 85.8723
R2863 vdd.t203 vdd.n1600 85.8723
R2864 vdd.n2997 vdd.n856 78.546
R2865 vdd.n2436 vdd.n1029 78.546
R2866 vdd.n278 vdd.n277 75.1835
R2867 vdd.n276 vdd.n275 75.1835
R2868 vdd.n274 vdd.n273 75.1835
R2869 vdd.n272 vdd.n271 75.1835
R2870 vdd.n270 vdd.n269 75.1835
R2871 vdd.n268 vdd.n267 75.1835
R2872 vdd.n266 vdd.n265 75.1835
R2873 vdd.n180 vdd.n179 75.1835
R2874 vdd.n178 vdd.n177 75.1835
R2875 vdd.n176 vdd.n175 75.1835
R2876 vdd.n174 vdd.n173 75.1835
R2877 vdd.n172 vdd.n171 75.1835
R2878 vdd.n170 vdd.n169 75.1835
R2879 vdd.n168 vdd.n167 75.1835
R2880 vdd.n83 vdd.n82 75.1835
R2881 vdd.n81 vdd.n80 75.1835
R2882 vdd.n79 vdd.n78 75.1835
R2883 vdd.n77 vdd.n76 75.1835
R2884 vdd.n75 vdd.n74 75.1835
R2885 vdd.n73 vdd.n72 75.1835
R2886 vdd.n71 vdd.n70 75.1835
R2887 vdd.n1770 vdd.n1769 75.1835
R2888 vdd.n1772 vdd.n1771 75.1835
R2889 vdd.n1774 vdd.n1773 75.1835
R2890 vdd.n1776 vdd.n1775 75.1835
R2891 vdd.n1778 vdd.n1777 75.1835
R2892 vdd.n1780 vdd.n1779 75.1835
R2893 vdd.n1782 vdd.n1781 75.1835
R2894 vdd.n1672 vdd.n1671 75.1835
R2895 vdd.n1674 vdd.n1673 75.1835
R2896 vdd.n1676 vdd.n1675 75.1835
R2897 vdd.n1678 vdd.n1677 75.1835
R2898 vdd.n1680 vdd.n1679 75.1835
R2899 vdd.n1682 vdd.n1681 75.1835
R2900 vdd.n1684 vdd.n1683 75.1835
R2901 vdd.n1575 vdd.n1574 75.1835
R2902 vdd.n1577 vdd.n1576 75.1835
R2903 vdd.n1579 vdd.n1578 75.1835
R2904 vdd.n1581 vdd.n1580 75.1835
R2905 vdd.n1583 vdd.n1582 75.1835
R2906 vdd.n1585 vdd.n1584 75.1835
R2907 vdd.n1587 vdd.n1586 75.1835
R2908 vdd.n2927 vdd.n2660 72.8958
R2909 vdd.n2927 vdd.n2661 72.8958
R2910 vdd.n2927 vdd.n2662 72.8958
R2911 vdd.n2927 vdd.n2663 72.8958
R2912 vdd.n2927 vdd.n2664 72.8958
R2913 vdd.n2927 vdd.n2665 72.8958
R2914 vdd.n2927 vdd.n2666 72.8958
R2915 vdd.n2927 vdd.n2667 72.8958
R2916 vdd.n2927 vdd.n2668 72.8958
R2917 vdd.n2927 vdd.n2669 72.8958
R2918 vdd.n2927 vdd.n2670 72.8958
R2919 vdd.n2927 vdd.n2671 72.8958
R2920 vdd.n2927 vdd.n2672 72.8958
R2921 vdd.n2927 vdd.n2673 72.8958
R2922 vdd.n2927 vdd.n2674 72.8958
R2923 vdd.n2927 vdd.n2675 72.8958
R2924 vdd.n2927 vdd.n2676 72.8958
R2925 vdd.n772 vdd.n756 72.8958
R2926 vdd.n3165 vdd.n756 72.8958
R2927 vdd.n766 vdd.n756 72.8958
R2928 vdd.n3172 vdd.n756 72.8958
R2929 vdd.n763 vdd.n756 72.8958
R2930 vdd.n3179 vdd.n756 72.8958
R2931 vdd.n760 vdd.n756 72.8958
R2932 vdd.n3186 vdd.n756 72.8958
R2933 vdd.n3189 vdd.n756 72.8958
R2934 vdd.n3045 vdd.n756 72.8958
R2935 vdd.n3050 vdd.n756 72.8958
R2936 vdd.n3044 vdd.n756 72.8958
R2937 vdd.n3057 vdd.n756 72.8958
R2938 vdd.n3041 vdd.n756 72.8958
R2939 vdd.n3064 vdd.n756 72.8958
R2940 vdd.n3038 vdd.n756 72.8958
R2941 vdd.n3071 vdd.n756 72.8958
R2942 vdd.n2378 vdd.n1081 72.8958
R2943 vdd.n1086 vdd.n1081 72.8958
R2944 vdd.n2371 vdd.n1081 72.8958
R2945 vdd.n2365 vdd.n1081 72.8958
R2946 vdd.n2363 vdd.n1081 72.8958
R2947 vdd.n2357 vdd.n1081 72.8958
R2948 vdd.n2355 vdd.n1081 72.8958
R2949 vdd.n2349 vdd.n1081 72.8958
R2950 vdd.n2347 vdd.n1081 72.8958
R2951 vdd.n2341 vdd.n1081 72.8958
R2952 vdd.n2339 vdd.n1081 72.8958
R2953 vdd.n2333 vdd.n1081 72.8958
R2954 vdd.n2331 vdd.n1081 72.8958
R2955 vdd.n2325 vdd.n1081 72.8958
R2956 vdd.n2323 vdd.n1081 72.8958
R2957 vdd.n2316 vdd.n1081 72.8958
R2958 vdd.n2314 vdd.n1081 72.8958
R2959 vdd.n2643 vdd.n939 72.8958
R2960 vdd.n2643 vdd.n940 72.8958
R2961 vdd.n2643 vdd.n941 72.8958
R2962 vdd.n2643 vdd.n942 72.8958
R2963 vdd.n2643 vdd.n943 72.8958
R2964 vdd.n2643 vdd.n944 72.8958
R2965 vdd.n2643 vdd.n945 72.8958
R2966 vdd.n2643 vdd.n946 72.8958
R2967 vdd.n2643 vdd.n947 72.8958
R2968 vdd.n2643 vdd.n948 72.8958
R2969 vdd.n2643 vdd.n949 72.8958
R2970 vdd.n2643 vdd.n950 72.8958
R2971 vdd.n2643 vdd.n951 72.8958
R2972 vdd.n2643 vdd.n952 72.8958
R2973 vdd.n2643 vdd.n953 72.8958
R2974 vdd.n2643 vdd.n954 72.8958
R2975 vdd.n2643 vdd.n955 72.8958
R2976 vdd.n2928 vdd.n2927 72.8958
R2977 vdd.n2927 vdd.n2644 72.8958
R2978 vdd.n2927 vdd.n2645 72.8958
R2979 vdd.n2927 vdd.n2646 72.8958
R2980 vdd.n2927 vdd.n2647 72.8958
R2981 vdd.n2927 vdd.n2648 72.8958
R2982 vdd.n2927 vdd.n2649 72.8958
R2983 vdd.n2927 vdd.n2650 72.8958
R2984 vdd.n2927 vdd.n2651 72.8958
R2985 vdd.n2927 vdd.n2652 72.8958
R2986 vdd.n2927 vdd.n2653 72.8958
R2987 vdd.n2927 vdd.n2654 72.8958
R2988 vdd.n2927 vdd.n2655 72.8958
R2989 vdd.n2927 vdd.n2656 72.8958
R2990 vdd.n2927 vdd.n2657 72.8958
R2991 vdd.n2927 vdd.n2658 72.8958
R2992 vdd.n2927 vdd.n2659 72.8958
R2993 vdd.n3093 vdd.n756 72.8958
R2994 vdd.n3099 vdd.n756 72.8958
R2995 vdd.n802 vdd.n756 72.8958
R2996 vdd.n3106 vdd.n756 72.8958
R2997 vdd.n799 vdd.n756 72.8958
R2998 vdd.n3113 vdd.n756 72.8958
R2999 vdd.n796 vdd.n756 72.8958
R3000 vdd.n3120 vdd.n756 72.8958
R3001 vdd.n793 vdd.n756 72.8958
R3002 vdd.n3128 vdd.n756 72.8958
R3003 vdd.n790 vdd.n756 72.8958
R3004 vdd.n3135 vdd.n756 72.8958
R3005 vdd.n787 vdd.n756 72.8958
R3006 vdd.n3142 vdd.n756 72.8958
R3007 vdd.n784 vdd.n756 72.8958
R3008 vdd.n3149 vdd.n756 72.8958
R3009 vdd.n3152 vdd.n756 72.8958
R3010 vdd.n2643 vdd.n937 72.8958
R3011 vdd.n2643 vdd.n936 72.8958
R3012 vdd.n2643 vdd.n935 72.8958
R3013 vdd.n2643 vdd.n934 72.8958
R3014 vdd.n2643 vdd.n933 72.8958
R3015 vdd.n2643 vdd.n932 72.8958
R3016 vdd.n2643 vdd.n931 72.8958
R3017 vdd.n2643 vdd.n930 72.8958
R3018 vdd.n2643 vdd.n929 72.8958
R3019 vdd.n2643 vdd.n928 72.8958
R3020 vdd.n2643 vdd.n927 72.8958
R3021 vdd.n2643 vdd.n926 72.8958
R3022 vdd.n2643 vdd.n925 72.8958
R3023 vdd.n2643 vdd.n924 72.8958
R3024 vdd.n2643 vdd.n923 72.8958
R3025 vdd.n2643 vdd.n922 72.8958
R3026 vdd.n2643 vdd.n921 72.8958
R3027 vdd.n2132 vdd.n1081 72.8958
R3028 vdd.n2134 vdd.n1081 72.8958
R3029 vdd.n2140 vdd.n1081 72.8958
R3030 vdd.n2142 vdd.n1081 72.8958
R3031 vdd.n2148 vdd.n1081 72.8958
R3032 vdd.n2150 vdd.n1081 72.8958
R3033 vdd.n2156 vdd.n1081 72.8958
R3034 vdd.n2158 vdd.n1081 72.8958
R3035 vdd.n2164 vdd.n1081 72.8958
R3036 vdd.n2166 vdd.n1081 72.8958
R3037 vdd.n2172 vdd.n1081 72.8958
R3038 vdd.n2174 vdd.n1081 72.8958
R3039 vdd.n2180 vdd.n1081 72.8958
R3040 vdd.n2182 vdd.n1081 72.8958
R3041 vdd.n2188 vdd.n1081 72.8958
R3042 vdd.n2190 vdd.n1081 72.8958
R3043 vdd.n2197 vdd.n1081 72.8958
R3044 vdd.n1454 vdd.n1453 66.2847
R3045 vdd.n1454 vdd.n1232 66.2847
R3046 vdd.n1454 vdd.n1233 66.2847
R3047 vdd.n1454 vdd.n1234 66.2847
R3048 vdd.n1454 vdd.n1235 66.2847
R3049 vdd.n1454 vdd.n1236 66.2847
R3050 vdd.n1454 vdd.n1237 66.2847
R3051 vdd.n1454 vdd.n1238 66.2847
R3052 vdd.n1454 vdd.n1239 66.2847
R3053 vdd.n1454 vdd.n1240 66.2847
R3054 vdd.n1454 vdd.n1241 66.2847
R3055 vdd.n1454 vdd.n1242 66.2847
R3056 vdd.n1454 vdd.n1243 66.2847
R3057 vdd.n1454 vdd.n1244 66.2847
R3058 vdd.n1454 vdd.n1245 66.2847
R3059 vdd.n1454 vdd.n1246 66.2847
R3060 vdd.n1454 vdd.n1247 66.2847
R3061 vdd.n1454 vdd.n1248 66.2847
R3062 vdd.n1454 vdd.n1249 66.2847
R3063 vdd.n1454 vdd.n1250 66.2847
R3064 vdd.n1454 vdd.n1251 66.2847
R3065 vdd.n1454 vdd.n1252 66.2847
R3066 vdd.n1454 vdd.n1253 66.2847
R3067 vdd.n1454 vdd.n1254 66.2847
R3068 vdd.n1454 vdd.n1255 66.2847
R3069 vdd.n1454 vdd.n1256 66.2847
R3070 vdd.n1454 vdd.n1257 66.2847
R3071 vdd.n1454 vdd.n1258 66.2847
R3072 vdd.n1454 vdd.n1259 66.2847
R3073 vdd.n1454 vdd.n1260 66.2847
R3074 vdd.n1454 vdd.n1261 66.2847
R3075 vdd.n1125 vdd.n1121 66.2847
R3076 vdd.n1997 vdd.n1125 66.2847
R3077 vdd.n2002 vdd.n1125 66.2847
R3078 vdd.n2007 vdd.n1125 66.2847
R3079 vdd.n1995 vdd.n1125 66.2847
R3080 vdd.n2014 vdd.n1125 66.2847
R3081 vdd.n1987 vdd.n1125 66.2847
R3082 vdd.n2021 vdd.n1125 66.2847
R3083 vdd.n1980 vdd.n1125 66.2847
R3084 vdd.n2028 vdd.n1125 66.2847
R3085 vdd.n1974 vdd.n1125 66.2847
R3086 vdd.n1969 vdd.n1125 66.2847
R3087 vdd.n2039 vdd.n1125 66.2847
R3088 vdd.n1961 vdd.n1125 66.2847
R3089 vdd.n2046 vdd.n1125 66.2847
R3090 vdd.n1954 vdd.n1125 66.2847
R3091 vdd.n2053 vdd.n1125 66.2847
R3092 vdd.n1947 vdd.n1125 66.2847
R3093 vdd.n2060 vdd.n1125 66.2847
R3094 vdd.n1940 vdd.n1125 66.2847
R3095 vdd.n2067 vdd.n1125 66.2847
R3096 vdd.n1934 vdd.n1125 66.2847
R3097 vdd.n1929 vdd.n1125 66.2847
R3098 vdd.n2078 vdd.n1125 66.2847
R3099 vdd.n1921 vdd.n1125 66.2847
R3100 vdd.n2085 vdd.n1125 66.2847
R3101 vdd.n1914 vdd.n1125 66.2847
R3102 vdd.n2092 vdd.n1125 66.2847
R3103 vdd.n2095 vdd.n1125 66.2847
R3104 vdd.n1905 vdd.n1125 66.2847
R3105 vdd.n2104 vdd.n1125 66.2847
R3106 vdd.n1899 vdd.n1125 66.2847
R3107 vdd.n3319 vdd.n658 66.2847
R3108 vdd.n663 vdd.n658 66.2847
R3109 vdd.n666 vdd.n658 66.2847
R3110 vdd.n3308 vdd.n658 66.2847
R3111 vdd.n3302 vdd.n658 66.2847
R3112 vdd.n3300 vdd.n658 66.2847
R3113 vdd.n3294 vdd.n658 66.2847
R3114 vdd.n3292 vdd.n658 66.2847
R3115 vdd.n3286 vdd.n658 66.2847
R3116 vdd.n3284 vdd.n658 66.2847
R3117 vdd.n3278 vdd.n658 66.2847
R3118 vdd.n3276 vdd.n658 66.2847
R3119 vdd.n3270 vdd.n658 66.2847
R3120 vdd.n3268 vdd.n658 66.2847
R3121 vdd.n3262 vdd.n658 66.2847
R3122 vdd.n3260 vdd.n658 66.2847
R3123 vdd.n3254 vdd.n658 66.2847
R3124 vdd.n3252 vdd.n658 66.2847
R3125 vdd.n3246 vdd.n658 66.2847
R3126 vdd.n3244 vdd.n658 66.2847
R3127 vdd.n727 vdd.n658 66.2847
R3128 vdd.n3235 vdd.n658 66.2847
R3129 vdd.n729 vdd.n658 66.2847
R3130 vdd.n3228 vdd.n658 66.2847
R3131 vdd.n3222 vdd.n658 66.2847
R3132 vdd.n3220 vdd.n658 66.2847
R3133 vdd.n3214 vdd.n658 66.2847
R3134 vdd.n3212 vdd.n658 66.2847
R3135 vdd.n3206 vdd.n658 66.2847
R3136 vdd.n750 vdd.n658 66.2847
R3137 vdd.n752 vdd.n658 66.2847
R3138 vdd.n3435 vdd.n3434 66.2847
R3139 vdd.n3435 vdd.n403 66.2847
R3140 vdd.n3435 vdd.n402 66.2847
R3141 vdd.n3435 vdd.n401 66.2847
R3142 vdd.n3435 vdd.n400 66.2847
R3143 vdd.n3435 vdd.n399 66.2847
R3144 vdd.n3435 vdd.n398 66.2847
R3145 vdd.n3435 vdd.n397 66.2847
R3146 vdd.n3435 vdd.n396 66.2847
R3147 vdd.n3435 vdd.n395 66.2847
R3148 vdd.n3435 vdd.n394 66.2847
R3149 vdd.n3435 vdd.n393 66.2847
R3150 vdd.n3435 vdd.n392 66.2847
R3151 vdd.n3435 vdd.n391 66.2847
R3152 vdd.n3435 vdd.n390 66.2847
R3153 vdd.n3435 vdd.n389 66.2847
R3154 vdd.n3435 vdd.n388 66.2847
R3155 vdd.n3435 vdd.n387 66.2847
R3156 vdd.n3435 vdd.n386 66.2847
R3157 vdd.n3435 vdd.n385 66.2847
R3158 vdd.n3435 vdd.n384 66.2847
R3159 vdd.n3435 vdd.n383 66.2847
R3160 vdd.n3435 vdd.n382 66.2847
R3161 vdd.n3435 vdd.n381 66.2847
R3162 vdd.n3435 vdd.n380 66.2847
R3163 vdd.n3435 vdd.n379 66.2847
R3164 vdd.n3435 vdd.n378 66.2847
R3165 vdd.n3435 vdd.n377 66.2847
R3166 vdd.n3435 vdd.n376 66.2847
R3167 vdd.n3435 vdd.n375 66.2847
R3168 vdd.n3435 vdd.n374 66.2847
R3169 vdd.n3435 vdd.n373 66.2847
R3170 vdd.n448 vdd.n373 52.4337
R3171 vdd.n454 vdd.n374 52.4337
R3172 vdd.n458 vdd.n375 52.4337
R3173 vdd.n464 vdd.n376 52.4337
R3174 vdd.n468 vdd.n377 52.4337
R3175 vdd.n474 vdd.n378 52.4337
R3176 vdd.n478 vdd.n379 52.4337
R3177 vdd.n484 vdd.n380 52.4337
R3178 vdd.n488 vdd.n381 52.4337
R3179 vdd.n494 vdd.n382 52.4337
R3180 vdd.n498 vdd.n383 52.4337
R3181 vdd.n504 vdd.n384 52.4337
R3182 vdd.n508 vdd.n385 52.4337
R3183 vdd.n514 vdd.n386 52.4337
R3184 vdd.n518 vdd.n387 52.4337
R3185 vdd.n524 vdd.n388 52.4337
R3186 vdd.n528 vdd.n389 52.4337
R3187 vdd.n534 vdd.n390 52.4337
R3188 vdd.n538 vdd.n391 52.4337
R3189 vdd.n544 vdd.n392 52.4337
R3190 vdd.n548 vdd.n393 52.4337
R3191 vdd.n554 vdd.n394 52.4337
R3192 vdd.n558 vdd.n395 52.4337
R3193 vdd.n564 vdd.n396 52.4337
R3194 vdd.n568 vdd.n397 52.4337
R3195 vdd.n574 vdd.n398 52.4337
R3196 vdd.n578 vdd.n399 52.4337
R3197 vdd.n584 vdd.n400 52.4337
R3198 vdd.n588 vdd.n401 52.4337
R3199 vdd.n594 vdd.n402 52.4337
R3200 vdd.n597 vdd.n403 52.4337
R3201 vdd.n3434 vdd.n3433 52.4337
R3202 vdd.n3319 vdd.n660 52.4337
R3203 vdd.n3317 vdd.n663 52.4337
R3204 vdd.n3313 vdd.n666 52.4337
R3205 vdd.n3309 vdd.n3308 52.4337
R3206 vdd.n3302 vdd.n669 52.4337
R3207 vdd.n3301 vdd.n3300 52.4337
R3208 vdd.n3294 vdd.n675 52.4337
R3209 vdd.n3293 vdd.n3292 52.4337
R3210 vdd.n3286 vdd.n681 52.4337
R3211 vdd.n3285 vdd.n3284 52.4337
R3212 vdd.n3278 vdd.n689 52.4337
R3213 vdd.n3277 vdd.n3276 52.4337
R3214 vdd.n3270 vdd.n695 52.4337
R3215 vdd.n3269 vdd.n3268 52.4337
R3216 vdd.n3262 vdd.n701 52.4337
R3217 vdd.n3261 vdd.n3260 52.4337
R3218 vdd.n3254 vdd.n707 52.4337
R3219 vdd.n3253 vdd.n3252 52.4337
R3220 vdd.n3246 vdd.n713 52.4337
R3221 vdd.n3245 vdd.n3244 52.4337
R3222 vdd.n727 vdd.n719 52.4337
R3223 vdd.n3236 vdd.n3235 52.4337
R3224 vdd.n3233 vdd.n729 52.4337
R3225 vdd.n3229 vdd.n3228 52.4337
R3226 vdd.n3222 vdd.n733 52.4337
R3227 vdd.n3221 vdd.n3220 52.4337
R3228 vdd.n3214 vdd.n739 52.4337
R3229 vdd.n3213 vdd.n3212 52.4337
R3230 vdd.n3206 vdd.n745 52.4337
R3231 vdd.n3205 vdd.n750 52.4337
R3232 vdd.n3201 vdd.n752 52.4337
R3233 vdd.n2106 vdd.n1899 52.4337
R3234 vdd.n2104 vdd.n2103 52.4337
R3235 vdd.n1906 vdd.n1905 52.4337
R3236 vdd.n2095 vdd.n2094 52.4337
R3237 vdd.n2092 vdd.n2091 52.4337
R3238 vdd.n2087 vdd.n1914 52.4337
R3239 vdd.n2085 vdd.n2084 52.4337
R3240 vdd.n2080 vdd.n1921 52.4337
R3241 vdd.n2078 vdd.n2077 52.4337
R3242 vdd.n1930 vdd.n1929 52.4337
R3243 vdd.n2069 vdd.n1934 52.4337
R3244 vdd.n2067 vdd.n2066 52.4337
R3245 vdd.n2062 vdd.n1940 52.4337
R3246 vdd.n2060 vdd.n2059 52.4337
R3247 vdd.n2055 vdd.n1947 52.4337
R3248 vdd.n2053 vdd.n2052 52.4337
R3249 vdd.n2048 vdd.n1954 52.4337
R3250 vdd.n2046 vdd.n2045 52.4337
R3251 vdd.n2041 vdd.n1961 52.4337
R3252 vdd.n2039 vdd.n2038 52.4337
R3253 vdd.n1970 vdd.n1969 52.4337
R3254 vdd.n2030 vdd.n1974 52.4337
R3255 vdd.n2028 vdd.n2027 52.4337
R3256 vdd.n2023 vdd.n1980 52.4337
R3257 vdd.n2021 vdd.n2020 52.4337
R3258 vdd.n2016 vdd.n1987 52.4337
R3259 vdd.n2014 vdd.n2013 52.4337
R3260 vdd.n2009 vdd.n1995 52.4337
R3261 vdd.n2007 vdd.n2006 52.4337
R3262 vdd.n2002 vdd.n2001 52.4337
R3263 vdd.n1997 vdd.n1996 52.4337
R3264 vdd.n2115 vdd.n1121 52.4337
R3265 vdd.n1453 vdd.n1452 52.4337
R3266 vdd.n1267 vdd.n1232 52.4337
R3267 vdd.n1269 vdd.n1233 52.4337
R3268 vdd.n1273 vdd.n1234 52.4337
R3269 vdd.n1275 vdd.n1235 52.4337
R3270 vdd.n1279 vdd.n1236 52.4337
R3271 vdd.n1281 vdd.n1237 52.4337
R3272 vdd.n1285 vdd.n1238 52.4337
R3273 vdd.n1287 vdd.n1239 52.4337
R3274 vdd.n1419 vdd.n1240 52.4337
R3275 vdd.n1291 vdd.n1241 52.4337
R3276 vdd.n1295 vdd.n1242 52.4337
R3277 vdd.n1297 vdd.n1243 52.4337
R3278 vdd.n1301 vdd.n1244 52.4337
R3279 vdd.n1303 vdd.n1245 52.4337
R3280 vdd.n1307 vdd.n1246 52.4337
R3281 vdd.n1309 vdd.n1247 52.4337
R3282 vdd.n1313 vdd.n1248 52.4337
R3283 vdd.n1315 vdd.n1249 52.4337
R3284 vdd.n1319 vdd.n1250 52.4337
R3285 vdd.n1383 vdd.n1251 52.4337
R3286 vdd.n1324 vdd.n1252 52.4337
R3287 vdd.n1326 vdd.n1253 52.4337
R3288 vdd.n1330 vdd.n1254 52.4337
R3289 vdd.n1332 vdd.n1255 52.4337
R3290 vdd.n1336 vdd.n1256 52.4337
R3291 vdd.n1338 vdd.n1257 52.4337
R3292 vdd.n1342 vdd.n1258 52.4337
R3293 vdd.n1344 vdd.n1259 52.4337
R3294 vdd.n1348 vdd.n1260 52.4337
R3295 vdd.n1350 vdd.n1261 52.4337
R3296 vdd.n1453 vdd.n1263 52.4337
R3297 vdd.n1268 vdd.n1232 52.4337
R3298 vdd.n1272 vdd.n1233 52.4337
R3299 vdd.n1274 vdd.n1234 52.4337
R3300 vdd.n1278 vdd.n1235 52.4337
R3301 vdd.n1280 vdd.n1236 52.4337
R3302 vdd.n1284 vdd.n1237 52.4337
R3303 vdd.n1286 vdd.n1238 52.4337
R3304 vdd.n1418 vdd.n1239 52.4337
R3305 vdd.n1290 vdd.n1240 52.4337
R3306 vdd.n1294 vdd.n1241 52.4337
R3307 vdd.n1296 vdd.n1242 52.4337
R3308 vdd.n1300 vdd.n1243 52.4337
R3309 vdd.n1302 vdd.n1244 52.4337
R3310 vdd.n1306 vdd.n1245 52.4337
R3311 vdd.n1308 vdd.n1246 52.4337
R3312 vdd.n1312 vdd.n1247 52.4337
R3313 vdd.n1314 vdd.n1248 52.4337
R3314 vdd.n1318 vdd.n1249 52.4337
R3315 vdd.n1320 vdd.n1250 52.4337
R3316 vdd.n1323 vdd.n1251 52.4337
R3317 vdd.n1325 vdd.n1252 52.4337
R3318 vdd.n1329 vdd.n1253 52.4337
R3319 vdd.n1331 vdd.n1254 52.4337
R3320 vdd.n1335 vdd.n1255 52.4337
R3321 vdd.n1337 vdd.n1256 52.4337
R3322 vdd.n1341 vdd.n1257 52.4337
R3323 vdd.n1343 vdd.n1258 52.4337
R3324 vdd.n1347 vdd.n1259 52.4337
R3325 vdd.n1349 vdd.n1260 52.4337
R3326 vdd.n1261 vdd.n1231 52.4337
R3327 vdd.n1121 vdd.n1120 52.4337
R3328 vdd.n1998 vdd.n1997 52.4337
R3329 vdd.n2003 vdd.n2002 52.4337
R3330 vdd.n2008 vdd.n2007 52.4337
R3331 vdd.n1995 vdd.n1988 52.4337
R3332 vdd.n2015 vdd.n2014 52.4337
R3333 vdd.n1987 vdd.n1981 52.4337
R3334 vdd.n2022 vdd.n2021 52.4337
R3335 vdd.n1980 vdd.n1975 52.4337
R3336 vdd.n2029 vdd.n2028 52.4337
R3337 vdd.n1974 vdd.n1973 52.4337
R3338 vdd.n1969 vdd.n1962 52.4337
R3339 vdd.n2040 vdd.n2039 52.4337
R3340 vdd.n1961 vdd.n1955 52.4337
R3341 vdd.n2047 vdd.n2046 52.4337
R3342 vdd.n1954 vdd.n1948 52.4337
R3343 vdd.n2054 vdd.n2053 52.4337
R3344 vdd.n1947 vdd.n1941 52.4337
R3345 vdd.n2061 vdd.n2060 52.4337
R3346 vdd.n1940 vdd.n1935 52.4337
R3347 vdd.n2068 vdd.n2067 52.4337
R3348 vdd.n1934 vdd.n1933 52.4337
R3349 vdd.n1929 vdd.n1922 52.4337
R3350 vdd.n2079 vdd.n2078 52.4337
R3351 vdd.n1921 vdd.n1915 52.4337
R3352 vdd.n2086 vdd.n2085 52.4337
R3353 vdd.n1914 vdd.n1908 52.4337
R3354 vdd.n2093 vdd.n2092 52.4337
R3355 vdd.n2096 vdd.n2095 52.4337
R3356 vdd.n1905 vdd.n1900 52.4337
R3357 vdd.n2105 vdd.n2104 52.4337
R3358 vdd.n1899 vdd.n1127 52.4337
R3359 vdd.n3320 vdd.n3319 52.4337
R3360 vdd.n3314 vdd.n663 52.4337
R3361 vdd.n3310 vdd.n666 52.4337
R3362 vdd.n3308 vdd.n3307 52.4337
R3363 vdd.n3303 vdd.n3302 52.4337
R3364 vdd.n3300 vdd.n3299 52.4337
R3365 vdd.n3295 vdd.n3294 52.4337
R3366 vdd.n3292 vdd.n3291 52.4337
R3367 vdd.n3287 vdd.n3286 52.4337
R3368 vdd.n3284 vdd.n3283 52.4337
R3369 vdd.n3279 vdd.n3278 52.4337
R3370 vdd.n3276 vdd.n3275 52.4337
R3371 vdd.n3271 vdd.n3270 52.4337
R3372 vdd.n3268 vdd.n3267 52.4337
R3373 vdd.n3263 vdd.n3262 52.4337
R3374 vdd.n3260 vdd.n3259 52.4337
R3375 vdd.n3255 vdd.n3254 52.4337
R3376 vdd.n3252 vdd.n3251 52.4337
R3377 vdd.n3247 vdd.n3246 52.4337
R3378 vdd.n3244 vdd.n3243 52.4337
R3379 vdd.n728 vdd.n727 52.4337
R3380 vdd.n3235 vdd.n3234 52.4337
R3381 vdd.n3230 vdd.n729 52.4337
R3382 vdd.n3228 vdd.n3227 52.4337
R3383 vdd.n3223 vdd.n3222 52.4337
R3384 vdd.n3220 vdd.n3219 52.4337
R3385 vdd.n3215 vdd.n3214 52.4337
R3386 vdd.n3212 vdd.n3211 52.4337
R3387 vdd.n3207 vdd.n3206 52.4337
R3388 vdd.n3202 vdd.n750 52.4337
R3389 vdd.n3198 vdd.n752 52.4337
R3390 vdd.n3434 vdd.n404 52.4337
R3391 vdd.n595 vdd.n403 52.4337
R3392 vdd.n589 vdd.n402 52.4337
R3393 vdd.n585 vdd.n401 52.4337
R3394 vdd.n579 vdd.n400 52.4337
R3395 vdd.n575 vdd.n399 52.4337
R3396 vdd.n569 vdd.n398 52.4337
R3397 vdd.n565 vdd.n397 52.4337
R3398 vdd.n559 vdd.n396 52.4337
R3399 vdd.n555 vdd.n395 52.4337
R3400 vdd.n549 vdd.n394 52.4337
R3401 vdd.n545 vdd.n393 52.4337
R3402 vdd.n539 vdd.n392 52.4337
R3403 vdd.n535 vdd.n391 52.4337
R3404 vdd.n529 vdd.n390 52.4337
R3405 vdd.n525 vdd.n389 52.4337
R3406 vdd.n519 vdd.n388 52.4337
R3407 vdd.n515 vdd.n387 52.4337
R3408 vdd.n509 vdd.n386 52.4337
R3409 vdd.n505 vdd.n385 52.4337
R3410 vdd.n499 vdd.n384 52.4337
R3411 vdd.n495 vdd.n383 52.4337
R3412 vdd.n489 vdd.n382 52.4337
R3413 vdd.n485 vdd.n381 52.4337
R3414 vdd.n479 vdd.n380 52.4337
R3415 vdd.n475 vdd.n379 52.4337
R3416 vdd.n469 vdd.n378 52.4337
R3417 vdd.n465 vdd.n377 52.4337
R3418 vdd.n459 vdd.n376 52.4337
R3419 vdd.n455 vdd.n375 52.4337
R3420 vdd.n449 vdd.n374 52.4337
R3421 vdd.n445 vdd.n373 52.4337
R3422 vdd.t142 vdd.t155 51.4683
R3423 vdd.n266 vdd.n264 42.0461
R3424 vdd.n168 vdd.n166 42.0461
R3425 vdd.n71 vdd.n69 42.0461
R3426 vdd.n1770 vdd.n1768 42.0461
R3427 vdd.n1672 vdd.n1670 42.0461
R3428 vdd.n1575 vdd.n1573 42.0461
R3429 vdd.n320 vdd.n319 41.6884
R3430 vdd.n222 vdd.n221 41.6884
R3431 vdd.n125 vdd.n124 41.6884
R3432 vdd.n1824 vdd.n1823 41.6884
R3433 vdd.n1726 vdd.n1725 41.6884
R3434 vdd.n1629 vdd.n1628 41.6884
R3435 vdd.n1230 vdd.n1229 41.1157
R3436 vdd.n1386 vdd.n1385 41.1157
R3437 vdd.n1422 vdd.n1421 41.1157
R3438 vdd.n407 vdd.n406 41.1157
R3439 vdd.n547 vdd.n420 41.1157
R3440 vdd.n433 vdd.n432 41.1157
R3441 vdd.n3152 vdd.n3151 39.2114
R3442 vdd.n3149 vdd.n3148 39.2114
R3443 vdd.n3144 vdd.n784 39.2114
R3444 vdd.n3142 vdd.n3141 39.2114
R3445 vdd.n3137 vdd.n787 39.2114
R3446 vdd.n3135 vdd.n3134 39.2114
R3447 vdd.n3130 vdd.n790 39.2114
R3448 vdd.n3128 vdd.n3127 39.2114
R3449 vdd.n3122 vdd.n793 39.2114
R3450 vdd.n3120 vdd.n3119 39.2114
R3451 vdd.n3115 vdd.n796 39.2114
R3452 vdd.n3113 vdd.n3112 39.2114
R3453 vdd.n3108 vdd.n799 39.2114
R3454 vdd.n3106 vdd.n3105 39.2114
R3455 vdd.n3101 vdd.n802 39.2114
R3456 vdd.n3099 vdd.n3098 39.2114
R3457 vdd.n3094 vdd.n3093 39.2114
R3458 vdd.n2928 vdd.n918 39.2114
R3459 vdd.n2749 vdd.n2644 39.2114
R3460 vdd.n2753 vdd.n2645 39.2114
R3461 vdd.n2757 vdd.n2646 39.2114
R3462 vdd.n2761 vdd.n2647 39.2114
R3463 vdd.n2765 vdd.n2648 39.2114
R3464 vdd.n2769 vdd.n2649 39.2114
R3465 vdd.n2773 vdd.n2650 39.2114
R3466 vdd.n2777 vdd.n2651 39.2114
R3467 vdd.n2781 vdd.n2652 39.2114
R3468 vdd.n2785 vdd.n2653 39.2114
R3469 vdd.n2789 vdd.n2654 39.2114
R3470 vdd.n2793 vdd.n2655 39.2114
R3471 vdd.n2797 vdd.n2656 39.2114
R3472 vdd.n2801 vdd.n2657 39.2114
R3473 vdd.n2805 vdd.n2658 39.2114
R3474 vdd.n2810 vdd.n2659 39.2114
R3475 vdd.n2638 vdd.n955 39.2114
R3476 vdd.n2634 vdd.n954 39.2114
R3477 vdd.n2630 vdd.n953 39.2114
R3478 vdd.n2626 vdd.n952 39.2114
R3479 vdd.n2622 vdd.n951 39.2114
R3480 vdd.n2618 vdd.n950 39.2114
R3481 vdd.n2614 vdd.n949 39.2114
R3482 vdd.n2610 vdd.n948 39.2114
R3483 vdd.n2606 vdd.n947 39.2114
R3484 vdd.n2602 vdd.n946 39.2114
R3485 vdd.n2598 vdd.n945 39.2114
R3486 vdd.n2594 vdd.n944 39.2114
R3487 vdd.n2590 vdd.n943 39.2114
R3488 vdd.n2586 vdd.n942 39.2114
R3489 vdd.n2582 vdd.n941 39.2114
R3490 vdd.n2577 vdd.n940 39.2114
R3491 vdd.n2573 vdd.n939 39.2114
R3492 vdd.n2378 vdd.n1084 39.2114
R3493 vdd.n2376 vdd.n1086 39.2114
R3494 vdd.n2372 vdd.n2371 39.2114
R3495 vdd.n2365 vdd.n1088 39.2114
R3496 vdd.n2364 vdd.n2363 39.2114
R3497 vdd.n2357 vdd.n1090 39.2114
R3498 vdd.n2356 vdd.n2355 39.2114
R3499 vdd.n2349 vdd.n1092 39.2114
R3500 vdd.n2348 vdd.n2347 39.2114
R3501 vdd.n2341 vdd.n1094 39.2114
R3502 vdd.n2340 vdd.n2339 39.2114
R3503 vdd.n2333 vdd.n1096 39.2114
R3504 vdd.n2332 vdd.n2331 39.2114
R3505 vdd.n2325 vdd.n1098 39.2114
R3506 vdd.n2324 vdd.n2323 39.2114
R3507 vdd.n2316 vdd.n1100 39.2114
R3508 vdd.n2315 vdd.n2314 39.2114
R3509 vdd.n3071 vdd.n3070 39.2114
R3510 vdd.n3066 vdd.n3038 39.2114
R3511 vdd.n3064 vdd.n3063 39.2114
R3512 vdd.n3059 vdd.n3041 39.2114
R3513 vdd.n3057 vdd.n3056 39.2114
R3514 vdd.n3052 vdd.n3044 39.2114
R3515 vdd.n3050 vdd.n3049 39.2114
R3516 vdd.n3045 vdd.n755 39.2114
R3517 vdd.n3189 vdd.n3188 39.2114
R3518 vdd.n3186 vdd.n3185 39.2114
R3519 vdd.n3181 vdd.n760 39.2114
R3520 vdd.n3179 vdd.n3178 39.2114
R3521 vdd.n3174 vdd.n763 39.2114
R3522 vdd.n3172 vdd.n3171 39.2114
R3523 vdd.n3167 vdd.n766 39.2114
R3524 vdd.n3165 vdd.n3164 39.2114
R3525 vdd.n3160 vdd.n772 39.2114
R3526 vdd.n2660 vdd.n914 39.2114
R3527 vdd.n2683 vdd.n2661 39.2114
R3528 vdd.n2687 vdd.n2662 39.2114
R3529 vdd.n2691 vdd.n2663 39.2114
R3530 vdd.n2695 vdd.n2664 39.2114
R3531 vdd.n2699 vdd.n2665 39.2114
R3532 vdd.n2703 vdd.n2666 39.2114
R3533 vdd.n2707 vdd.n2667 39.2114
R3534 vdd.n2711 vdd.n2668 39.2114
R3535 vdd.n2715 vdd.n2669 39.2114
R3536 vdd.n2719 vdd.n2670 39.2114
R3537 vdd.n2723 vdd.n2671 39.2114
R3538 vdd.n2727 vdd.n2672 39.2114
R3539 vdd.n2731 vdd.n2673 39.2114
R3540 vdd.n2735 vdd.n2674 39.2114
R3541 vdd.n2739 vdd.n2675 39.2114
R3542 vdd.n2743 vdd.n2676 39.2114
R3543 vdd.n2682 vdd.n2660 39.2114
R3544 vdd.n2686 vdd.n2661 39.2114
R3545 vdd.n2690 vdd.n2662 39.2114
R3546 vdd.n2694 vdd.n2663 39.2114
R3547 vdd.n2698 vdd.n2664 39.2114
R3548 vdd.n2702 vdd.n2665 39.2114
R3549 vdd.n2706 vdd.n2666 39.2114
R3550 vdd.n2710 vdd.n2667 39.2114
R3551 vdd.n2714 vdd.n2668 39.2114
R3552 vdd.n2718 vdd.n2669 39.2114
R3553 vdd.n2722 vdd.n2670 39.2114
R3554 vdd.n2726 vdd.n2671 39.2114
R3555 vdd.n2730 vdd.n2672 39.2114
R3556 vdd.n2734 vdd.n2673 39.2114
R3557 vdd.n2738 vdd.n2674 39.2114
R3558 vdd.n2742 vdd.n2675 39.2114
R3559 vdd.n2677 vdd.n2676 39.2114
R3560 vdd.n772 vdd.n767 39.2114
R3561 vdd.n3166 vdd.n3165 39.2114
R3562 vdd.n766 vdd.n764 39.2114
R3563 vdd.n3173 vdd.n3172 39.2114
R3564 vdd.n763 vdd.n761 39.2114
R3565 vdd.n3180 vdd.n3179 39.2114
R3566 vdd.n760 vdd.n758 39.2114
R3567 vdd.n3187 vdd.n3186 39.2114
R3568 vdd.n3190 vdd.n3189 39.2114
R3569 vdd.n3046 vdd.n3045 39.2114
R3570 vdd.n3051 vdd.n3050 39.2114
R3571 vdd.n3044 vdd.n3042 39.2114
R3572 vdd.n3058 vdd.n3057 39.2114
R3573 vdd.n3041 vdd.n3039 39.2114
R3574 vdd.n3065 vdd.n3064 39.2114
R3575 vdd.n3038 vdd.n3036 39.2114
R3576 vdd.n3072 vdd.n3071 39.2114
R3577 vdd.n2379 vdd.n2378 39.2114
R3578 vdd.n2373 vdd.n1086 39.2114
R3579 vdd.n2371 vdd.n2370 39.2114
R3580 vdd.n2366 vdd.n2365 39.2114
R3581 vdd.n2363 vdd.n2362 39.2114
R3582 vdd.n2358 vdd.n2357 39.2114
R3583 vdd.n2355 vdd.n2354 39.2114
R3584 vdd.n2350 vdd.n2349 39.2114
R3585 vdd.n2347 vdd.n2346 39.2114
R3586 vdd.n2342 vdd.n2341 39.2114
R3587 vdd.n2339 vdd.n2338 39.2114
R3588 vdd.n2334 vdd.n2333 39.2114
R3589 vdd.n2331 vdd.n2330 39.2114
R3590 vdd.n2326 vdd.n2325 39.2114
R3591 vdd.n2323 vdd.n2322 39.2114
R3592 vdd.n2317 vdd.n2316 39.2114
R3593 vdd.n2314 vdd.n2313 39.2114
R3594 vdd.n2576 vdd.n939 39.2114
R3595 vdd.n2581 vdd.n940 39.2114
R3596 vdd.n2585 vdd.n941 39.2114
R3597 vdd.n2589 vdd.n942 39.2114
R3598 vdd.n2593 vdd.n943 39.2114
R3599 vdd.n2597 vdd.n944 39.2114
R3600 vdd.n2601 vdd.n945 39.2114
R3601 vdd.n2605 vdd.n946 39.2114
R3602 vdd.n2609 vdd.n947 39.2114
R3603 vdd.n2613 vdd.n948 39.2114
R3604 vdd.n2617 vdd.n949 39.2114
R3605 vdd.n2621 vdd.n950 39.2114
R3606 vdd.n2625 vdd.n951 39.2114
R3607 vdd.n2629 vdd.n952 39.2114
R3608 vdd.n2633 vdd.n953 39.2114
R3609 vdd.n2637 vdd.n954 39.2114
R3610 vdd.n957 vdd.n955 39.2114
R3611 vdd.n2929 vdd.n2928 39.2114
R3612 vdd.n2752 vdd.n2644 39.2114
R3613 vdd.n2756 vdd.n2645 39.2114
R3614 vdd.n2760 vdd.n2646 39.2114
R3615 vdd.n2764 vdd.n2647 39.2114
R3616 vdd.n2768 vdd.n2648 39.2114
R3617 vdd.n2772 vdd.n2649 39.2114
R3618 vdd.n2776 vdd.n2650 39.2114
R3619 vdd.n2780 vdd.n2651 39.2114
R3620 vdd.n2784 vdd.n2652 39.2114
R3621 vdd.n2788 vdd.n2653 39.2114
R3622 vdd.n2792 vdd.n2654 39.2114
R3623 vdd.n2796 vdd.n2655 39.2114
R3624 vdd.n2800 vdd.n2656 39.2114
R3625 vdd.n2804 vdd.n2657 39.2114
R3626 vdd.n2809 vdd.n2658 39.2114
R3627 vdd.n2812 vdd.n2659 39.2114
R3628 vdd.n3093 vdd.n803 39.2114
R3629 vdd.n3100 vdd.n3099 39.2114
R3630 vdd.n802 vdd.n800 39.2114
R3631 vdd.n3107 vdd.n3106 39.2114
R3632 vdd.n799 vdd.n797 39.2114
R3633 vdd.n3114 vdd.n3113 39.2114
R3634 vdd.n796 vdd.n794 39.2114
R3635 vdd.n3121 vdd.n3120 39.2114
R3636 vdd.n793 vdd.n791 39.2114
R3637 vdd.n3129 vdd.n3128 39.2114
R3638 vdd.n790 vdd.n788 39.2114
R3639 vdd.n3136 vdd.n3135 39.2114
R3640 vdd.n787 vdd.n785 39.2114
R3641 vdd.n3143 vdd.n3142 39.2114
R3642 vdd.n784 vdd.n782 39.2114
R3643 vdd.n3150 vdd.n3149 39.2114
R3644 vdd.n3153 vdd.n3152 39.2114
R3645 vdd.n966 vdd.n921 39.2114
R3646 vdd.n2565 vdd.n922 39.2114
R3647 vdd.n2561 vdd.n923 39.2114
R3648 vdd.n2557 vdd.n924 39.2114
R3649 vdd.n2553 vdd.n925 39.2114
R3650 vdd.n2549 vdd.n926 39.2114
R3651 vdd.n2545 vdd.n927 39.2114
R3652 vdd.n2541 vdd.n928 39.2114
R3653 vdd.n2537 vdd.n929 39.2114
R3654 vdd.n2533 vdd.n930 39.2114
R3655 vdd.n2529 vdd.n931 39.2114
R3656 vdd.n2525 vdd.n932 39.2114
R3657 vdd.n2521 vdd.n933 39.2114
R3658 vdd.n2517 vdd.n934 39.2114
R3659 vdd.n2513 vdd.n935 39.2114
R3660 vdd.n2509 vdd.n936 39.2114
R3661 vdd.n2505 vdd.n937 39.2114
R3662 vdd.n2132 vdd.n1080 39.2114
R3663 vdd.n2135 vdd.n2134 39.2114
R3664 vdd.n2140 vdd.n2139 39.2114
R3665 vdd.n2143 vdd.n2142 39.2114
R3666 vdd.n2148 vdd.n2147 39.2114
R3667 vdd.n2151 vdd.n2150 39.2114
R3668 vdd.n2156 vdd.n2155 39.2114
R3669 vdd.n2159 vdd.n2158 39.2114
R3670 vdd.n2164 vdd.n2163 39.2114
R3671 vdd.n2167 vdd.n2166 39.2114
R3672 vdd.n2172 vdd.n2171 39.2114
R3673 vdd.n2175 vdd.n2174 39.2114
R3674 vdd.n2180 vdd.n2179 39.2114
R3675 vdd.n2183 vdd.n2182 39.2114
R3676 vdd.n2188 vdd.n2187 39.2114
R3677 vdd.n2191 vdd.n2190 39.2114
R3678 vdd.n2197 vdd.n2196 39.2114
R3679 vdd.n2502 vdd.n937 39.2114
R3680 vdd.n2506 vdd.n936 39.2114
R3681 vdd.n2510 vdd.n935 39.2114
R3682 vdd.n2514 vdd.n934 39.2114
R3683 vdd.n2518 vdd.n933 39.2114
R3684 vdd.n2522 vdd.n932 39.2114
R3685 vdd.n2526 vdd.n931 39.2114
R3686 vdd.n2530 vdd.n930 39.2114
R3687 vdd.n2534 vdd.n929 39.2114
R3688 vdd.n2538 vdd.n928 39.2114
R3689 vdd.n2542 vdd.n927 39.2114
R3690 vdd.n2546 vdd.n926 39.2114
R3691 vdd.n2550 vdd.n925 39.2114
R3692 vdd.n2554 vdd.n924 39.2114
R3693 vdd.n2558 vdd.n923 39.2114
R3694 vdd.n2562 vdd.n922 39.2114
R3695 vdd.n2566 vdd.n921 39.2114
R3696 vdd.n2133 vdd.n2132 39.2114
R3697 vdd.n2134 vdd.n2130 39.2114
R3698 vdd.n2141 vdd.n2140 39.2114
R3699 vdd.n2142 vdd.n2128 39.2114
R3700 vdd.n2149 vdd.n2148 39.2114
R3701 vdd.n2150 vdd.n2126 39.2114
R3702 vdd.n2157 vdd.n2156 39.2114
R3703 vdd.n2158 vdd.n2124 39.2114
R3704 vdd.n2165 vdd.n2164 39.2114
R3705 vdd.n2166 vdd.n1114 39.2114
R3706 vdd.n2173 vdd.n2172 39.2114
R3707 vdd.n2174 vdd.n1112 39.2114
R3708 vdd.n2181 vdd.n2180 39.2114
R3709 vdd.n2182 vdd.n1110 39.2114
R3710 vdd.n2189 vdd.n2188 39.2114
R3711 vdd.n2190 vdd.n1106 39.2114
R3712 vdd.n2198 vdd.n2197 39.2114
R3713 vdd.n2119 vdd.n2118 37.2369
R3714 vdd.n2035 vdd.n1968 37.2369
R3715 vdd.n2074 vdd.n1928 37.2369
R3716 vdd.n3241 vdd.n724 37.2369
R3717 vdd.n688 vdd.n687 37.2369
R3718 vdd.n3197 vdd.n3196 37.2369
R3719 vdd.n2194 vdd.n1108 30.449
R3720 vdd.n970 vdd.n969 30.449
R3721 vdd.n2319 vdd.n1102 30.449
R3722 vdd.n2579 vdd.n960 30.449
R3723 vdd.n2680 vdd.n2679 30.449
R3724 vdd.n806 vdd.n805 30.449
R3725 vdd.n2807 vdd.n2748 30.449
R3726 vdd.n770 vdd.n769 30.449
R3727 vdd.n2382 vdd.n2381 30.4395
R3728 vdd.n2641 vdd.n958 30.4395
R3729 vdd.n2574 vdd.n961 30.4395
R3730 vdd.n2312 vdd.n2311 30.4395
R3731 vdd.n2814 vdd.n2813 30.4395
R3732 vdd.n3095 vdd.n3092 30.4395
R3733 vdd.n2932 vdd.n2931 30.4395
R3734 vdd.n3156 vdd.n3155 30.4395
R3735 vdd.n3075 vdd.n3074 30.4395
R3736 vdd.n3161 vdd.n771 30.4395
R3737 vdd.n2925 vdd.n2924 30.4395
R3738 vdd.n2936 vdd.n913 30.4395
R3739 vdd.n2386 vdd.n1079 30.4395
R3740 vdd.n2569 vdd.n2568 30.4395
R3741 vdd.n2501 vdd.n2500 30.4395
R3742 vdd.n2201 vdd.n2200 30.4395
R3743 vdd.n1460 vdd.n1226 19.3944
R3744 vdd.n1460 vdd.n1216 19.3944
R3745 vdd.n1472 vdd.n1216 19.3944
R3746 vdd.n1472 vdd.n1214 19.3944
R3747 vdd.n1476 vdd.n1214 19.3944
R3748 vdd.n1476 vdd.n1204 19.3944
R3749 vdd.n1489 vdd.n1204 19.3944
R3750 vdd.n1489 vdd.n1202 19.3944
R3751 vdd.n1493 vdd.n1202 19.3944
R3752 vdd.n1493 vdd.n1194 19.3944
R3753 vdd.n1506 vdd.n1194 19.3944
R3754 vdd.n1506 vdd.n1192 19.3944
R3755 vdd.n1510 vdd.n1192 19.3944
R3756 vdd.n1510 vdd.n1181 19.3944
R3757 vdd.n1522 vdd.n1181 19.3944
R3758 vdd.n1522 vdd.n1179 19.3944
R3759 vdd.n1526 vdd.n1179 19.3944
R3760 vdd.n1526 vdd.n1170 19.3944
R3761 vdd.n1834 vdd.n1170 19.3944
R3762 vdd.n1834 vdd.n1168 19.3944
R3763 vdd.n1838 vdd.n1168 19.3944
R3764 vdd.n1838 vdd.n1159 19.3944
R3765 vdd.n1850 vdd.n1159 19.3944
R3766 vdd.n1850 vdd.n1157 19.3944
R3767 vdd.n1854 vdd.n1157 19.3944
R3768 vdd.n1854 vdd.n1147 19.3944
R3769 vdd.n1867 vdd.n1147 19.3944
R3770 vdd.n1867 vdd.n1145 19.3944
R3771 vdd.n1871 vdd.n1145 19.3944
R3772 vdd.n1871 vdd.n1137 19.3944
R3773 vdd.n1884 vdd.n1137 19.3944
R3774 vdd.n1884 vdd.n1134 19.3944
R3775 vdd.n1890 vdd.n1134 19.3944
R3776 vdd.n1890 vdd.n1135 19.3944
R3777 vdd.n1135 vdd.n1123 19.3944
R3778 vdd.n1379 vdd.n1321 19.3944
R3779 vdd.n1379 vdd.n1378 19.3944
R3780 vdd.n1378 vdd.n1377 19.3944
R3781 vdd.n1377 vdd.n1327 19.3944
R3782 vdd.n1373 vdd.n1327 19.3944
R3783 vdd.n1373 vdd.n1372 19.3944
R3784 vdd.n1372 vdd.n1371 19.3944
R3785 vdd.n1371 vdd.n1333 19.3944
R3786 vdd.n1367 vdd.n1333 19.3944
R3787 vdd.n1367 vdd.n1366 19.3944
R3788 vdd.n1366 vdd.n1365 19.3944
R3789 vdd.n1365 vdd.n1339 19.3944
R3790 vdd.n1361 vdd.n1339 19.3944
R3791 vdd.n1361 vdd.n1360 19.3944
R3792 vdd.n1360 vdd.n1359 19.3944
R3793 vdd.n1359 vdd.n1345 19.3944
R3794 vdd.n1355 vdd.n1345 19.3944
R3795 vdd.n1355 vdd.n1354 19.3944
R3796 vdd.n1354 vdd.n1353 19.3944
R3797 vdd.n1353 vdd.n1351 19.3944
R3798 vdd.n1417 vdd.n1416 19.3944
R3799 vdd.n1416 vdd.n1292 19.3944
R3800 vdd.n1412 vdd.n1292 19.3944
R3801 vdd.n1412 vdd.n1411 19.3944
R3802 vdd.n1411 vdd.n1410 19.3944
R3803 vdd.n1410 vdd.n1298 19.3944
R3804 vdd.n1406 vdd.n1298 19.3944
R3805 vdd.n1406 vdd.n1405 19.3944
R3806 vdd.n1405 vdd.n1404 19.3944
R3807 vdd.n1404 vdd.n1304 19.3944
R3808 vdd.n1400 vdd.n1304 19.3944
R3809 vdd.n1400 vdd.n1399 19.3944
R3810 vdd.n1399 vdd.n1398 19.3944
R3811 vdd.n1398 vdd.n1310 19.3944
R3812 vdd.n1394 vdd.n1310 19.3944
R3813 vdd.n1394 vdd.n1393 19.3944
R3814 vdd.n1393 vdd.n1392 19.3944
R3815 vdd.n1392 vdd.n1316 19.3944
R3816 vdd.n1388 vdd.n1316 19.3944
R3817 vdd.n1388 vdd.n1387 19.3944
R3818 vdd.n1451 vdd.n1450 19.3944
R3819 vdd.n1450 vdd.n1265 19.3944
R3820 vdd.n1446 vdd.n1265 19.3944
R3821 vdd.n1446 vdd.n1445 19.3944
R3822 vdd.n1445 vdd.n1444 19.3944
R3823 vdd.n1444 vdd.n1270 19.3944
R3824 vdd.n1440 vdd.n1270 19.3944
R3825 vdd.n1440 vdd.n1439 19.3944
R3826 vdd.n1439 vdd.n1438 19.3944
R3827 vdd.n1438 vdd.n1276 19.3944
R3828 vdd.n1434 vdd.n1276 19.3944
R3829 vdd.n1434 vdd.n1433 19.3944
R3830 vdd.n1433 vdd.n1432 19.3944
R3831 vdd.n1432 vdd.n1282 19.3944
R3832 vdd.n1428 vdd.n1282 19.3944
R3833 vdd.n1428 vdd.n1427 19.3944
R3834 vdd.n1427 vdd.n1426 19.3944
R3835 vdd.n1426 vdd.n1288 19.3944
R3836 vdd.n2031 vdd.n1966 19.3944
R3837 vdd.n2031 vdd.n1972 19.3944
R3838 vdd.n2026 vdd.n1972 19.3944
R3839 vdd.n2026 vdd.n2025 19.3944
R3840 vdd.n2025 vdd.n2024 19.3944
R3841 vdd.n2024 vdd.n1979 19.3944
R3842 vdd.n2019 vdd.n1979 19.3944
R3843 vdd.n2019 vdd.n2018 19.3944
R3844 vdd.n2018 vdd.n2017 19.3944
R3845 vdd.n2017 vdd.n1986 19.3944
R3846 vdd.n2012 vdd.n1986 19.3944
R3847 vdd.n2012 vdd.n2011 19.3944
R3848 vdd.n2011 vdd.n2010 19.3944
R3849 vdd.n2010 vdd.n1994 19.3944
R3850 vdd.n2005 vdd.n1994 19.3944
R3851 vdd.n2005 vdd.n2004 19.3944
R3852 vdd.n2000 vdd.n1999 19.3944
R3853 vdd.n2120 vdd.n1119 19.3944
R3854 vdd.n2070 vdd.n1926 19.3944
R3855 vdd.n2070 vdd.n1932 19.3944
R3856 vdd.n2065 vdd.n1932 19.3944
R3857 vdd.n2065 vdd.n2064 19.3944
R3858 vdd.n2064 vdd.n2063 19.3944
R3859 vdd.n2063 vdd.n1939 19.3944
R3860 vdd.n2058 vdd.n1939 19.3944
R3861 vdd.n2058 vdd.n2057 19.3944
R3862 vdd.n2057 vdd.n2056 19.3944
R3863 vdd.n2056 vdd.n1946 19.3944
R3864 vdd.n2051 vdd.n1946 19.3944
R3865 vdd.n2051 vdd.n2050 19.3944
R3866 vdd.n2050 vdd.n2049 19.3944
R3867 vdd.n2049 vdd.n1953 19.3944
R3868 vdd.n2044 vdd.n1953 19.3944
R3869 vdd.n2044 vdd.n2043 19.3944
R3870 vdd.n2043 vdd.n2042 19.3944
R3871 vdd.n2042 vdd.n1960 19.3944
R3872 vdd.n2037 vdd.n1960 19.3944
R3873 vdd.n2037 vdd.n2036 19.3944
R3874 vdd.n2108 vdd.n2107 19.3944
R3875 vdd.n2107 vdd.n1898 19.3944
R3876 vdd.n2102 vdd.n2101 19.3944
R3877 vdd.n2097 vdd.n1902 19.3944
R3878 vdd.n2097 vdd.n1904 19.3944
R3879 vdd.n1907 vdd.n1904 19.3944
R3880 vdd.n2090 vdd.n1907 19.3944
R3881 vdd.n2090 vdd.n2089 19.3944
R3882 vdd.n2089 vdd.n2088 19.3944
R3883 vdd.n2088 vdd.n1913 19.3944
R3884 vdd.n2083 vdd.n1913 19.3944
R3885 vdd.n2083 vdd.n2082 19.3944
R3886 vdd.n2082 vdd.n2081 19.3944
R3887 vdd.n2081 vdd.n1920 19.3944
R3888 vdd.n2076 vdd.n1920 19.3944
R3889 vdd.n2076 vdd.n2075 19.3944
R3890 vdd.n1464 vdd.n1222 19.3944
R3891 vdd.n1464 vdd.n1220 19.3944
R3892 vdd.n1468 vdd.n1220 19.3944
R3893 vdd.n1468 vdd.n1210 19.3944
R3894 vdd.n1481 vdd.n1210 19.3944
R3895 vdd.n1481 vdd.n1208 19.3944
R3896 vdd.n1485 vdd.n1208 19.3944
R3897 vdd.n1485 vdd.n1199 19.3944
R3898 vdd.n1498 vdd.n1199 19.3944
R3899 vdd.n1498 vdd.n1197 19.3944
R3900 vdd.n1502 vdd.n1197 19.3944
R3901 vdd.n1502 vdd.n1188 19.3944
R3902 vdd.n1514 vdd.n1188 19.3944
R3903 vdd.n1514 vdd.n1186 19.3944
R3904 vdd.n1518 vdd.n1186 19.3944
R3905 vdd.n1518 vdd.n1176 19.3944
R3906 vdd.n1531 vdd.n1176 19.3944
R3907 vdd.n1531 vdd.n1174 19.3944
R3908 vdd.n1830 vdd.n1174 19.3944
R3909 vdd.n1830 vdd.n1165 19.3944
R3910 vdd.n1842 vdd.n1165 19.3944
R3911 vdd.n1842 vdd.n1163 19.3944
R3912 vdd.n1846 vdd.n1163 19.3944
R3913 vdd.n1846 vdd.n1153 19.3944
R3914 vdd.n1859 vdd.n1153 19.3944
R3915 vdd.n1859 vdd.n1151 19.3944
R3916 vdd.n1863 vdd.n1151 19.3944
R3917 vdd.n1863 vdd.n1142 19.3944
R3918 vdd.n1876 vdd.n1142 19.3944
R3919 vdd.n1876 vdd.n1140 19.3944
R3920 vdd.n1880 vdd.n1140 19.3944
R3921 vdd.n1880 vdd.n1130 19.3944
R3922 vdd.n1894 vdd.n1130 19.3944
R3923 vdd.n1894 vdd.n1128 19.3944
R3924 vdd.n2111 vdd.n1128 19.3944
R3925 vdd.n3329 vdd.n655 19.3944
R3926 vdd.n3333 vdd.n655 19.3944
R3927 vdd.n3333 vdd.n646 19.3944
R3928 vdd.n3345 vdd.n646 19.3944
R3929 vdd.n3345 vdd.n644 19.3944
R3930 vdd.n3349 vdd.n644 19.3944
R3931 vdd.n3349 vdd.n633 19.3944
R3932 vdd.n3361 vdd.n633 19.3944
R3933 vdd.n3361 vdd.n631 19.3944
R3934 vdd.n3365 vdd.n631 19.3944
R3935 vdd.n3365 vdd.n622 19.3944
R3936 vdd.n3378 vdd.n622 19.3944
R3937 vdd.n3378 vdd.n620 19.3944
R3938 vdd.n3385 vdd.n620 19.3944
R3939 vdd.n3385 vdd.n3384 19.3944
R3940 vdd.n3384 vdd.n610 19.3944
R3941 vdd.n3398 vdd.n610 19.3944
R3942 vdd.n3399 vdd.n3398 19.3944
R3943 vdd.n3400 vdd.n3399 19.3944
R3944 vdd.n3400 vdd.n608 19.3944
R3945 vdd.n3405 vdd.n608 19.3944
R3946 vdd.n3406 vdd.n3405 19.3944
R3947 vdd.n3407 vdd.n3406 19.3944
R3948 vdd.n3407 vdd.n606 19.3944
R3949 vdd.n3412 vdd.n606 19.3944
R3950 vdd.n3413 vdd.n3412 19.3944
R3951 vdd.n3414 vdd.n3413 19.3944
R3952 vdd.n3414 vdd.n604 19.3944
R3953 vdd.n3420 vdd.n604 19.3944
R3954 vdd.n3421 vdd.n3420 19.3944
R3955 vdd.n3422 vdd.n3421 19.3944
R3956 vdd.n3422 vdd.n602 19.3944
R3957 vdd.n3427 vdd.n602 19.3944
R3958 vdd.n3428 vdd.n3427 19.3944
R3959 vdd.n3429 vdd.n3428 19.3944
R3960 vdd.n550 vdd.n417 19.3944
R3961 vdd.n556 vdd.n417 19.3944
R3962 vdd.n557 vdd.n556 19.3944
R3963 vdd.n560 vdd.n557 19.3944
R3964 vdd.n560 vdd.n415 19.3944
R3965 vdd.n566 vdd.n415 19.3944
R3966 vdd.n567 vdd.n566 19.3944
R3967 vdd.n570 vdd.n567 19.3944
R3968 vdd.n570 vdd.n413 19.3944
R3969 vdd.n576 vdd.n413 19.3944
R3970 vdd.n577 vdd.n576 19.3944
R3971 vdd.n580 vdd.n577 19.3944
R3972 vdd.n580 vdd.n411 19.3944
R3973 vdd.n586 vdd.n411 19.3944
R3974 vdd.n587 vdd.n586 19.3944
R3975 vdd.n590 vdd.n587 19.3944
R3976 vdd.n590 vdd.n409 19.3944
R3977 vdd.n596 vdd.n409 19.3944
R3978 vdd.n598 vdd.n596 19.3944
R3979 vdd.n599 vdd.n598 19.3944
R3980 vdd.n497 vdd.n496 19.3944
R3981 vdd.n500 vdd.n497 19.3944
R3982 vdd.n500 vdd.n429 19.3944
R3983 vdd.n506 vdd.n429 19.3944
R3984 vdd.n507 vdd.n506 19.3944
R3985 vdd.n510 vdd.n507 19.3944
R3986 vdd.n510 vdd.n427 19.3944
R3987 vdd.n516 vdd.n427 19.3944
R3988 vdd.n517 vdd.n516 19.3944
R3989 vdd.n520 vdd.n517 19.3944
R3990 vdd.n520 vdd.n425 19.3944
R3991 vdd.n526 vdd.n425 19.3944
R3992 vdd.n527 vdd.n526 19.3944
R3993 vdd.n530 vdd.n527 19.3944
R3994 vdd.n530 vdd.n423 19.3944
R3995 vdd.n536 vdd.n423 19.3944
R3996 vdd.n537 vdd.n536 19.3944
R3997 vdd.n540 vdd.n537 19.3944
R3998 vdd.n540 vdd.n421 19.3944
R3999 vdd.n546 vdd.n421 19.3944
R4000 vdd.n447 vdd.n446 19.3944
R4001 vdd.n450 vdd.n447 19.3944
R4002 vdd.n450 vdd.n441 19.3944
R4003 vdd.n456 vdd.n441 19.3944
R4004 vdd.n457 vdd.n456 19.3944
R4005 vdd.n460 vdd.n457 19.3944
R4006 vdd.n460 vdd.n439 19.3944
R4007 vdd.n466 vdd.n439 19.3944
R4008 vdd.n467 vdd.n466 19.3944
R4009 vdd.n470 vdd.n467 19.3944
R4010 vdd.n470 vdd.n437 19.3944
R4011 vdd.n476 vdd.n437 19.3944
R4012 vdd.n477 vdd.n476 19.3944
R4013 vdd.n480 vdd.n477 19.3944
R4014 vdd.n480 vdd.n435 19.3944
R4015 vdd.n486 vdd.n435 19.3944
R4016 vdd.n487 vdd.n486 19.3944
R4017 vdd.n490 vdd.n487 19.3944
R4018 vdd.n3325 vdd.n652 19.3944
R4019 vdd.n3337 vdd.n652 19.3944
R4020 vdd.n3337 vdd.n650 19.3944
R4021 vdd.n3341 vdd.n650 19.3944
R4022 vdd.n3341 vdd.n640 19.3944
R4023 vdd.n3353 vdd.n640 19.3944
R4024 vdd.n3353 vdd.n638 19.3944
R4025 vdd.n3357 vdd.n638 19.3944
R4026 vdd.n3357 vdd.n628 19.3944
R4027 vdd.n3370 vdd.n628 19.3944
R4028 vdd.n3370 vdd.n626 19.3944
R4029 vdd.n3374 vdd.n626 19.3944
R4030 vdd.n3374 vdd.n617 19.3944
R4031 vdd.n3389 vdd.n617 19.3944
R4032 vdd.n3389 vdd.n615 19.3944
R4033 vdd.n3393 vdd.n615 19.3944
R4034 vdd.n3393 vdd.n324 19.3944
R4035 vdd.n3471 vdd.n324 19.3944
R4036 vdd.n3471 vdd.n325 19.3944
R4037 vdd.n3465 vdd.n325 19.3944
R4038 vdd.n3465 vdd.n3464 19.3944
R4039 vdd.n3464 vdd.n3463 19.3944
R4040 vdd.n3463 vdd.n337 19.3944
R4041 vdd.n3457 vdd.n337 19.3944
R4042 vdd.n3457 vdd.n3456 19.3944
R4043 vdd.n3456 vdd.n3455 19.3944
R4044 vdd.n3455 vdd.n347 19.3944
R4045 vdd.n3449 vdd.n347 19.3944
R4046 vdd.n3449 vdd.n3448 19.3944
R4047 vdd.n3448 vdd.n3447 19.3944
R4048 vdd.n3447 vdd.n358 19.3944
R4049 vdd.n3441 vdd.n358 19.3944
R4050 vdd.n3441 vdd.n3440 19.3944
R4051 vdd.n3440 vdd.n3439 19.3944
R4052 vdd.n3439 vdd.n369 19.3944
R4053 vdd.n3282 vdd.n3281 19.3944
R4054 vdd.n3281 vdd.n3280 19.3944
R4055 vdd.n3280 vdd.n694 19.3944
R4056 vdd.n3274 vdd.n694 19.3944
R4057 vdd.n3274 vdd.n3273 19.3944
R4058 vdd.n3273 vdd.n3272 19.3944
R4059 vdd.n3272 vdd.n700 19.3944
R4060 vdd.n3266 vdd.n700 19.3944
R4061 vdd.n3266 vdd.n3265 19.3944
R4062 vdd.n3265 vdd.n3264 19.3944
R4063 vdd.n3264 vdd.n706 19.3944
R4064 vdd.n3258 vdd.n706 19.3944
R4065 vdd.n3258 vdd.n3257 19.3944
R4066 vdd.n3257 vdd.n3256 19.3944
R4067 vdd.n3256 vdd.n712 19.3944
R4068 vdd.n3250 vdd.n712 19.3944
R4069 vdd.n3250 vdd.n3249 19.3944
R4070 vdd.n3249 vdd.n3248 19.3944
R4071 vdd.n3248 vdd.n718 19.3944
R4072 vdd.n3242 vdd.n718 19.3944
R4073 vdd.n3322 vdd.n3321 19.3944
R4074 vdd.n3321 vdd.n662 19.3944
R4075 vdd.n3316 vdd.n3315 19.3944
R4076 vdd.n3312 vdd.n3311 19.3944
R4077 vdd.n3311 vdd.n668 19.3944
R4078 vdd.n3306 vdd.n668 19.3944
R4079 vdd.n3306 vdd.n3305 19.3944
R4080 vdd.n3305 vdd.n3304 19.3944
R4081 vdd.n3304 vdd.n674 19.3944
R4082 vdd.n3298 vdd.n674 19.3944
R4083 vdd.n3298 vdd.n3297 19.3944
R4084 vdd.n3297 vdd.n3296 19.3944
R4085 vdd.n3296 vdd.n680 19.3944
R4086 vdd.n3290 vdd.n680 19.3944
R4087 vdd.n3290 vdd.n3289 19.3944
R4088 vdd.n3289 vdd.n3288 19.3944
R4089 vdd.n3237 vdd.n722 19.3944
R4090 vdd.n3237 vdd.n726 19.3944
R4091 vdd.n3232 vdd.n726 19.3944
R4092 vdd.n3232 vdd.n3231 19.3944
R4093 vdd.n3231 vdd.n732 19.3944
R4094 vdd.n3226 vdd.n732 19.3944
R4095 vdd.n3226 vdd.n3225 19.3944
R4096 vdd.n3225 vdd.n3224 19.3944
R4097 vdd.n3224 vdd.n738 19.3944
R4098 vdd.n3218 vdd.n738 19.3944
R4099 vdd.n3218 vdd.n3217 19.3944
R4100 vdd.n3217 vdd.n3216 19.3944
R4101 vdd.n3216 vdd.n744 19.3944
R4102 vdd.n3210 vdd.n744 19.3944
R4103 vdd.n3210 vdd.n3209 19.3944
R4104 vdd.n3209 vdd.n3208 19.3944
R4105 vdd.n3204 vdd.n3203 19.3944
R4106 vdd.n3200 vdd.n3199 19.3944
R4107 vdd.n1386 vdd.n1321 19.0066
R4108 vdd.n2035 vdd.n1966 19.0066
R4109 vdd.n550 vdd.n547 19.0066
R4110 vdd.n3241 vdd.n722 19.0066
R4111 vdd.n1454 vdd.n1224 18.5924
R4112 vdd.n2113 vdd.n1125 18.5924
R4113 vdd.n3327 vdd.n658 18.5924
R4114 vdd.n3436 vdd.n3435 18.5924
R4115 vdd.n1108 vdd.n1107 16.0975
R4116 vdd.n969 vdd.n968 16.0975
R4117 vdd.n1229 vdd.n1228 16.0975
R4118 vdd.n1385 vdd.n1384 16.0975
R4119 vdd.n1421 vdd.n1420 16.0975
R4120 vdd.n2118 vdd.n2117 16.0975
R4121 vdd.n1968 vdd.n1967 16.0975
R4122 vdd.n1928 vdd.n1927 16.0975
R4123 vdd.n1102 vdd.n1101 16.0975
R4124 vdd.n960 vdd.n959 16.0975
R4125 vdd.n2679 vdd.n2678 16.0975
R4126 vdd.n406 vdd.n405 16.0975
R4127 vdd.n420 vdd.n419 16.0975
R4128 vdd.n432 vdd.n431 16.0975
R4129 vdd.n724 vdd.n723 16.0975
R4130 vdd.n687 vdd.n686 16.0975
R4131 vdd.n805 vdd.n804 16.0975
R4132 vdd.n2748 vdd.n2747 16.0975
R4133 vdd.n3196 vdd.n3195 16.0975
R4134 vdd.n769 vdd.n768 16.0975
R4135 vdd.t155 vdd.n2643 15.4182
R4136 vdd.n2927 vdd.t142 15.4182
R4137 vdd.n28 vdd.n27 14.5238
R4138 vdd.n2384 vdd.n1081 13.6043
R4139 vdd.n3158 vdd.n756 13.6043
R4140 vdd.n316 vdd.n281 13.1884
R4141 vdd.n261 vdd.n226 13.1884
R4142 vdd.n218 vdd.n183 13.1884
R4143 vdd.n163 vdd.n128 13.1884
R4144 vdd.n121 vdd.n86 13.1884
R4145 vdd.n66 vdd.n31 13.1884
R4146 vdd.n1765 vdd.n1730 13.1884
R4147 vdd.n1820 vdd.n1785 13.1884
R4148 vdd.n1667 vdd.n1632 13.1884
R4149 vdd.n1722 vdd.n1687 13.1884
R4150 vdd.n1570 vdd.n1535 13.1884
R4151 vdd.n1625 vdd.n1590 13.1884
R4152 vdd.n1422 vdd.n1417 12.9944
R4153 vdd.n1422 vdd.n1288 12.9944
R4154 vdd.n2074 vdd.n1926 12.9944
R4155 vdd.n2075 vdd.n2074 12.9944
R4156 vdd.n496 vdd.n433 12.9944
R4157 vdd.n490 vdd.n433 12.9944
R4158 vdd.n3282 vdd.n688 12.9944
R4159 vdd.n3288 vdd.n688 12.9944
R4160 vdd.n317 vdd.n279 12.8005
R4161 vdd.n312 vdd.n283 12.8005
R4162 vdd.n262 vdd.n224 12.8005
R4163 vdd.n257 vdd.n228 12.8005
R4164 vdd.n219 vdd.n181 12.8005
R4165 vdd.n214 vdd.n185 12.8005
R4166 vdd.n164 vdd.n126 12.8005
R4167 vdd.n159 vdd.n130 12.8005
R4168 vdd.n122 vdd.n84 12.8005
R4169 vdd.n117 vdd.n88 12.8005
R4170 vdd.n67 vdd.n29 12.8005
R4171 vdd.n62 vdd.n33 12.8005
R4172 vdd.n1766 vdd.n1728 12.8005
R4173 vdd.n1761 vdd.n1732 12.8005
R4174 vdd.n1821 vdd.n1783 12.8005
R4175 vdd.n1816 vdd.n1787 12.8005
R4176 vdd.n1668 vdd.n1630 12.8005
R4177 vdd.n1663 vdd.n1634 12.8005
R4178 vdd.n1723 vdd.n1685 12.8005
R4179 vdd.n1718 vdd.n1689 12.8005
R4180 vdd.n1571 vdd.n1533 12.8005
R4181 vdd.n1566 vdd.n1537 12.8005
R4182 vdd.n1626 vdd.n1588 12.8005
R4183 vdd.n1621 vdd.n1592 12.8005
R4184 vdd.n311 vdd.n284 12.0247
R4185 vdd.n256 vdd.n229 12.0247
R4186 vdd.n213 vdd.n186 12.0247
R4187 vdd.n158 vdd.n131 12.0247
R4188 vdd.n116 vdd.n89 12.0247
R4189 vdd.n61 vdd.n34 12.0247
R4190 vdd.n1760 vdd.n1733 12.0247
R4191 vdd.n1815 vdd.n1788 12.0247
R4192 vdd.n1662 vdd.n1635 12.0247
R4193 vdd.n1717 vdd.n1690 12.0247
R4194 vdd.n1565 vdd.n1538 12.0247
R4195 vdd.n1620 vdd.n1593 12.0247
R4196 vdd.n1462 vdd.n1224 11.337
R4197 vdd.n1470 vdd.n1218 11.337
R4198 vdd.n1470 vdd.n1212 11.337
R4199 vdd.n1479 vdd.n1212 11.337
R4200 vdd.n1487 vdd.n1206 11.337
R4201 vdd.n1496 vdd.n1495 11.337
R4202 vdd.n1512 vdd.n1190 11.337
R4203 vdd.n1520 vdd.n1183 11.337
R4204 vdd.n1529 vdd.n1528 11.337
R4205 vdd.n1832 vdd.n1172 11.337
R4206 vdd.n1848 vdd.n1161 11.337
R4207 vdd.n1857 vdd.n1155 11.337
R4208 vdd.n1865 vdd.n1149 11.337
R4209 vdd.n1874 vdd.n1873 11.337
R4210 vdd.n1882 vdd.n1132 11.337
R4211 vdd.n1892 vdd.n1132 11.337
R4212 vdd.n2113 vdd.n1124 11.337
R4213 vdd.n3327 vdd.n659 11.337
R4214 vdd.n3335 vdd.n648 11.337
R4215 vdd.n3343 vdd.n648 11.337
R4216 vdd.n3351 vdd.n642 11.337
R4217 vdd.n3359 vdd.n635 11.337
R4218 vdd.n3368 vdd.n3367 11.337
R4219 vdd.n3376 vdd.n624 11.337
R4220 vdd.n3395 vdd.n613 11.337
R4221 vdd.n3469 vdd.n328 11.337
R4222 vdd.n3467 vdd.n332 11.337
R4223 vdd.n3461 vdd.n3460 11.337
R4224 vdd.n3453 vdd.n349 11.337
R4225 vdd.n3452 vdd.n3451 11.337
R4226 vdd.n3445 vdd.n3444 11.337
R4227 vdd.n3444 vdd.n3443 11.337
R4228 vdd.n3443 vdd.n363 11.337
R4229 vdd.n3437 vdd.n3436 11.337
R4230 vdd.n308 vdd.n307 11.249
R4231 vdd.n253 vdd.n252 11.249
R4232 vdd.n210 vdd.n209 11.249
R4233 vdd.n155 vdd.n154 11.249
R4234 vdd.n113 vdd.n112 11.249
R4235 vdd.n58 vdd.n57 11.249
R4236 vdd.n1757 vdd.n1756 11.249
R4237 vdd.n1812 vdd.n1811 11.249
R4238 vdd.n1659 vdd.n1658 11.249
R4239 vdd.n1714 vdd.n1713 11.249
R4240 vdd.n1562 vdd.n1561 11.249
R4241 vdd.n1617 vdd.n1616 11.249
R4242 vdd.n1882 vdd.t234 10.7702
R4243 vdd.n3343 vdd.t215 10.7702
R4244 vdd.n293 vdd.n292 10.7238
R4245 vdd.n238 vdd.n237 10.7238
R4246 vdd.n195 vdd.n194 10.7238
R4247 vdd.n140 vdd.n139 10.7238
R4248 vdd.n98 vdd.n97 10.7238
R4249 vdd.n43 vdd.n42 10.7238
R4250 vdd.n1742 vdd.n1741 10.7238
R4251 vdd.n1797 vdd.n1796 10.7238
R4252 vdd.n1644 vdd.n1643 10.7238
R4253 vdd.n1699 vdd.n1698 10.7238
R4254 vdd.n1547 vdd.n1546 10.7238
R4255 vdd.n1602 vdd.n1601 10.7238
R4256 vdd.n2382 vdd.n1073 10.6151
R4257 vdd.n2392 vdd.n1073 10.6151
R4258 vdd.n2393 vdd.n2392 10.6151
R4259 vdd.n2394 vdd.n2393 10.6151
R4260 vdd.n2394 vdd.n1061 10.6151
R4261 vdd.n2404 vdd.n1061 10.6151
R4262 vdd.n2405 vdd.n2404 10.6151
R4263 vdd.n2406 vdd.n2405 10.6151
R4264 vdd.n2406 vdd.n1049 10.6151
R4265 vdd.n2416 vdd.n1049 10.6151
R4266 vdd.n2417 vdd.n2416 10.6151
R4267 vdd.n2418 vdd.n2417 10.6151
R4268 vdd.n2418 vdd.n1036 10.6151
R4269 vdd.n2428 vdd.n1036 10.6151
R4270 vdd.n2429 vdd.n2428 10.6151
R4271 vdd.n2430 vdd.n2429 10.6151
R4272 vdd.n2430 vdd.n1024 10.6151
R4273 vdd.n2441 vdd.n1024 10.6151
R4274 vdd.n2442 vdd.n2441 10.6151
R4275 vdd.n2443 vdd.n2442 10.6151
R4276 vdd.n2443 vdd.n1012 10.6151
R4277 vdd.n2453 vdd.n1012 10.6151
R4278 vdd.n2454 vdd.n2453 10.6151
R4279 vdd.n2455 vdd.n2454 10.6151
R4280 vdd.n2455 vdd.n1000 10.6151
R4281 vdd.n2465 vdd.n1000 10.6151
R4282 vdd.n2466 vdd.n2465 10.6151
R4283 vdd.n2467 vdd.n2466 10.6151
R4284 vdd.n2467 vdd.n990 10.6151
R4285 vdd.n2477 vdd.n990 10.6151
R4286 vdd.n2478 vdd.n2477 10.6151
R4287 vdd.n2479 vdd.n2478 10.6151
R4288 vdd.n2479 vdd.n977 10.6151
R4289 vdd.n2491 vdd.n977 10.6151
R4290 vdd.n2492 vdd.n2491 10.6151
R4291 vdd.n2494 vdd.n2492 10.6151
R4292 vdd.n2494 vdd.n2493 10.6151
R4293 vdd.n2493 vdd.n958 10.6151
R4294 vdd.n2641 vdd.n2640 10.6151
R4295 vdd.n2640 vdd.n2639 10.6151
R4296 vdd.n2639 vdd.n2636 10.6151
R4297 vdd.n2636 vdd.n2635 10.6151
R4298 vdd.n2635 vdd.n2632 10.6151
R4299 vdd.n2632 vdd.n2631 10.6151
R4300 vdd.n2631 vdd.n2628 10.6151
R4301 vdd.n2628 vdd.n2627 10.6151
R4302 vdd.n2627 vdd.n2624 10.6151
R4303 vdd.n2624 vdd.n2623 10.6151
R4304 vdd.n2623 vdd.n2620 10.6151
R4305 vdd.n2620 vdd.n2619 10.6151
R4306 vdd.n2619 vdd.n2616 10.6151
R4307 vdd.n2616 vdd.n2615 10.6151
R4308 vdd.n2615 vdd.n2612 10.6151
R4309 vdd.n2612 vdd.n2611 10.6151
R4310 vdd.n2611 vdd.n2608 10.6151
R4311 vdd.n2608 vdd.n2607 10.6151
R4312 vdd.n2607 vdd.n2604 10.6151
R4313 vdd.n2604 vdd.n2603 10.6151
R4314 vdd.n2603 vdd.n2600 10.6151
R4315 vdd.n2600 vdd.n2599 10.6151
R4316 vdd.n2599 vdd.n2596 10.6151
R4317 vdd.n2596 vdd.n2595 10.6151
R4318 vdd.n2595 vdd.n2592 10.6151
R4319 vdd.n2592 vdd.n2591 10.6151
R4320 vdd.n2591 vdd.n2588 10.6151
R4321 vdd.n2588 vdd.n2587 10.6151
R4322 vdd.n2587 vdd.n2584 10.6151
R4323 vdd.n2584 vdd.n2583 10.6151
R4324 vdd.n2583 vdd.n2580 10.6151
R4325 vdd.n2578 vdd.n2575 10.6151
R4326 vdd.n2575 vdd.n2574 10.6151
R4327 vdd.n2311 vdd.n2310 10.6151
R4328 vdd.n2310 vdd.n2308 10.6151
R4329 vdd.n2308 vdd.n2307 10.6151
R4330 vdd.n2307 vdd.n2305 10.6151
R4331 vdd.n2305 vdd.n2304 10.6151
R4332 vdd.n2304 vdd.n2302 10.6151
R4333 vdd.n2302 vdd.n2301 10.6151
R4334 vdd.n2301 vdd.n2299 10.6151
R4335 vdd.n2299 vdd.n2298 10.6151
R4336 vdd.n2298 vdd.n2296 10.6151
R4337 vdd.n2296 vdd.n2295 10.6151
R4338 vdd.n2295 vdd.n2293 10.6151
R4339 vdd.n2293 vdd.n2292 10.6151
R4340 vdd.n2292 vdd.n2290 10.6151
R4341 vdd.n2290 vdd.n2289 10.6151
R4342 vdd.n2289 vdd.n2287 10.6151
R4343 vdd.n2287 vdd.n2286 10.6151
R4344 vdd.n2286 vdd.n2284 10.6151
R4345 vdd.n2284 vdd.n2283 10.6151
R4346 vdd.n2283 vdd.n2281 10.6151
R4347 vdd.n2281 vdd.n2280 10.6151
R4348 vdd.n2280 vdd.n2278 10.6151
R4349 vdd.n2278 vdd.n2277 10.6151
R4350 vdd.n2277 vdd.n1104 10.6151
R4351 vdd.n2244 vdd.n1104 10.6151
R4352 vdd.n2245 vdd.n2244 10.6151
R4353 vdd.n2247 vdd.n2245 10.6151
R4354 vdd.n2248 vdd.n2247 10.6151
R4355 vdd.n2261 vdd.n2248 10.6151
R4356 vdd.n2261 vdd.n2260 10.6151
R4357 vdd.n2260 vdd.n2259 10.6151
R4358 vdd.n2259 vdd.n2257 10.6151
R4359 vdd.n2257 vdd.n2256 10.6151
R4360 vdd.n2256 vdd.n2254 10.6151
R4361 vdd.n2254 vdd.n2253 10.6151
R4362 vdd.n2253 vdd.n2250 10.6151
R4363 vdd.n2250 vdd.n2249 10.6151
R4364 vdd.n2249 vdd.n961 10.6151
R4365 vdd.n2381 vdd.n2380 10.6151
R4366 vdd.n2380 vdd.n1085 10.6151
R4367 vdd.n2375 vdd.n1085 10.6151
R4368 vdd.n2375 vdd.n2374 10.6151
R4369 vdd.n2374 vdd.n1087 10.6151
R4370 vdd.n2369 vdd.n1087 10.6151
R4371 vdd.n2369 vdd.n2368 10.6151
R4372 vdd.n2368 vdd.n2367 10.6151
R4373 vdd.n2367 vdd.n1089 10.6151
R4374 vdd.n2361 vdd.n1089 10.6151
R4375 vdd.n2361 vdd.n2360 10.6151
R4376 vdd.n2360 vdd.n2359 10.6151
R4377 vdd.n2359 vdd.n1091 10.6151
R4378 vdd.n2353 vdd.n1091 10.6151
R4379 vdd.n2353 vdd.n2352 10.6151
R4380 vdd.n2352 vdd.n2351 10.6151
R4381 vdd.n2351 vdd.n1093 10.6151
R4382 vdd.n2345 vdd.n1093 10.6151
R4383 vdd.n2345 vdd.n2344 10.6151
R4384 vdd.n2344 vdd.n2343 10.6151
R4385 vdd.n2343 vdd.n1095 10.6151
R4386 vdd.n2337 vdd.n1095 10.6151
R4387 vdd.n2337 vdd.n2336 10.6151
R4388 vdd.n2336 vdd.n2335 10.6151
R4389 vdd.n2335 vdd.n1097 10.6151
R4390 vdd.n2329 vdd.n1097 10.6151
R4391 vdd.n2329 vdd.n2328 10.6151
R4392 vdd.n2328 vdd.n2327 10.6151
R4393 vdd.n2327 vdd.n1099 10.6151
R4394 vdd.n2321 vdd.n1099 10.6151
R4395 vdd.n2321 vdd.n2320 10.6151
R4396 vdd.n2318 vdd.n1103 10.6151
R4397 vdd.n2312 vdd.n1103 10.6151
R4398 vdd.n2816 vdd.n2814 10.6151
R4399 vdd.n2817 vdd.n2816 10.6151
R4400 vdd.n2916 vdd.n2817 10.6151
R4401 vdd.n2916 vdd.n2915 10.6151
R4402 vdd.n2915 vdd.n2914 10.6151
R4403 vdd.n2914 vdd.n2912 10.6151
R4404 vdd.n2912 vdd.n2911 10.6151
R4405 vdd.n2911 vdd.n2909 10.6151
R4406 vdd.n2909 vdd.n2908 10.6151
R4407 vdd.n2908 vdd.n2818 10.6151
R4408 vdd.n2858 vdd.n2818 10.6151
R4409 vdd.n2859 vdd.n2858 10.6151
R4410 vdd.n2861 vdd.n2859 10.6151
R4411 vdd.n2862 vdd.n2861 10.6151
R4412 vdd.n2892 vdd.n2862 10.6151
R4413 vdd.n2892 vdd.n2891 10.6151
R4414 vdd.n2891 vdd.n2890 10.6151
R4415 vdd.n2890 vdd.n2888 10.6151
R4416 vdd.n2888 vdd.n2887 10.6151
R4417 vdd.n2887 vdd.n2885 10.6151
R4418 vdd.n2885 vdd.n2884 10.6151
R4419 vdd.n2884 vdd.n2882 10.6151
R4420 vdd.n2882 vdd.n2881 10.6151
R4421 vdd.n2881 vdd.n2879 10.6151
R4422 vdd.n2879 vdd.n2878 10.6151
R4423 vdd.n2878 vdd.n2876 10.6151
R4424 vdd.n2876 vdd.n2875 10.6151
R4425 vdd.n2875 vdd.n2873 10.6151
R4426 vdd.n2873 vdd.n2872 10.6151
R4427 vdd.n2872 vdd.n2870 10.6151
R4428 vdd.n2870 vdd.n2869 10.6151
R4429 vdd.n2869 vdd.n2867 10.6151
R4430 vdd.n2867 vdd.n2866 10.6151
R4431 vdd.n2866 vdd.n2864 10.6151
R4432 vdd.n2864 vdd.n2863 10.6151
R4433 vdd.n2863 vdd.n807 10.6151
R4434 vdd.n3091 vdd.n807 10.6151
R4435 vdd.n3092 vdd.n3091 10.6151
R4436 vdd.n2931 vdd.n2930 10.6151
R4437 vdd.n2930 vdd.n919 10.6151
R4438 vdd.n2750 vdd.n919 10.6151
R4439 vdd.n2751 vdd.n2750 10.6151
R4440 vdd.n2754 vdd.n2751 10.6151
R4441 vdd.n2755 vdd.n2754 10.6151
R4442 vdd.n2758 vdd.n2755 10.6151
R4443 vdd.n2759 vdd.n2758 10.6151
R4444 vdd.n2762 vdd.n2759 10.6151
R4445 vdd.n2763 vdd.n2762 10.6151
R4446 vdd.n2766 vdd.n2763 10.6151
R4447 vdd.n2767 vdd.n2766 10.6151
R4448 vdd.n2770 vdd.n2767 10.6151
R4449 vdd.n2771 vdd.n2770 10.6151
R4450 vdd.n2774 vdd.n2771 10.6151
R4451 vdd.n2775 vdd.n2774 10.6151
R4452 vdd.n2778 vdd.n2775 10.6151
R4453 vdd.n2779 vdd.n2778 10.6151
R4454 vdd.n2782 vdd.n2779 10.6151
R4455 vdd.n2783 vdd.n2782 10.6151
R4456 vdd.n2786 vdd.n2783 10.6151
R4457 vdd.n2787 vdd.n2786 10.6151
R4458 vdd.n2790 vdd.n2787 10.6151
R4459 vdd.n2791 vdd.n2790 10.6151
R4460 vdd.n2794 vdd.n2791 10.6151
R4461 vdd.n2795 vdd.n2794 10.6151
R4462 vdd.n2798 vdd.n2795 10.6151
R4463 vdd.n2799 vdd.n2798 10.6151
R4464 vdd.n2802 vdd.n2799 10.6151
R4465 vdd.n2803 vdd.n2802 10.6151
R4466 vdd.n2806 vdd.n2803 10.6151
R4467 vdd.n2811 vdd.n2808 10.6151
R4468 vdd.n2813 vdd.n2811 10.6151
R4469 vdd.n2932 vdd.n908 10.6151
R4470 vdd.n2942 vdd.n908 10.6151
R4471 vdd.n2943 vdd.n2942 10.6151
R4472 vdd.n2944 vdd.n2943 10.6151
R4473 vdd.n2944 vdd.n896 10.6151
R4474 vdd.n2954 vdd.n896 10.6151
R4475 vdd.n2955 vdd.n2954 10.6151
R4476 vdd.n2956 vdd.n2955 10.6151
R4477 vdd.n2956 vdd.n886 10.6151
R4478 vdd.n2966 vdd.n886 10.6151
R4479 vdd.n2967 vdd.n2966 10.6151
R4480 vdd.n2968 vdd.n2967 10.6151
R4481 vdd.n2968 vdd.n874 10.6151
R4482 vdd.n2978 vdd.n874 10.6151
R4483 vdd.n2979 vdd.n2978 10.6151
R4484 vdd.n2980 vdd.n2979 10.6151
R4485 vdd.n2980 vdd.n863 10.6151
R4486 vdd.n2990 vdd.n863 10.6151
R4487 vdd.n2991 vdd.n2990 10.6151
R4488 vdd.n2992 vdd.n2991 10.6151
R4489 vdd.n2992 vdd.n850 10.6151
R4490 vdd.n3003 vdd.n850 10.6151
R4491 vdd.n3004 vdd.n3003 10.6151
R4492 vdd.n3005 vdd.n3004 10.6151
R4493 vdd.n3005 vdd.n837 10.6151
R4494 vdd.n3015 vdd.n837 10.6151
R4495 vdd.n3016 vdd.n3015 10.6151
R4496 vdd.n3017 vdd.n3016 10.6151
R4497 vdd.n3017 vdd.n826 10.6151
R4498 vdd.n3027 vdd.n826 10.6151
R4499 vdd.n3028 vdd.n3027 10.6151
R4500 vdd.n3029 vdd.n3028 10.6151
R4501 vdd.n3029 vdd.n812 10.6151
R4502 vdd.n3084 vdd.n812 10.6151
R4503 vdd.n3085 vdd.n3084 10.6151
R4504 vdd.n3086 vdd.n3085 10.6151
R4505 vdd.n3086 vdd.n779 10.6151
R4506 vdd.n3156 vdd.n779 10.6151
R4507 vdd.n3155 vdd.n3154 10.6151
R4508 vdd.n3154 vdd.n780 10.6151
R4509 vdd.n781 vdd.n780 10.6151
R4510 vdd.n3147 vdd.n781 10.6151
R4511 vdd.n3147 vdd.n3146 10.6151
R4512 vdd.n3146 vdd.n3145 10.6151
R4513 vdd.n3145 vdd.n783 10.6151
R4514 vdd.n3140 vdd.n783 10.6151
R4515 vdd.n3140 vdd.n3139 10.6151
R4516 vdd.n3139 vdd.n3138 10.6151
R4517 vdd.n3138 vdd.n786 10.6151
R4518 vdd.n3133 vdd.n786 10.6151
R4519 vdd.n3133 vdd.n3132 10.6151
R4520 vdd.n3132 vdd.n3131 10.6151
R4521 vdd.n3131 vdd.n789 10.6151
R4522 vdd.n3126 vdd.n789 10.6151
R4523 vdd.n3126 vdd.n3125 10.6151
R4524 vdd.n3125 vdd.n3123 10.6151
R4525 vdd.n3123 vdd.n792 10.6151
R4526 vdd.n3118 vdd.n792 10.6151
R4527 vdd.n3118 vdd.n3117 10.6151
R4528 vdd.n3117 vdd.n3116 10.6151
R4529 vdd.n3116 vdd.n795 10.6151
R4530 vdd.n3111 vdd.n795 10.6151
R4531 vdd.n3111 vdd.n3110 10.6151
R4532 vdd.n3110 vdd.n3109 10.6151
R4533 vdd.n3109 vdd.n798 10.6151
R4534 vdd.n3104 vdd.n798 10.6151
R4535 vdd.n3104 vdd.n3103 10.6151
R4536 vdd.n3103 vdd.n3102 10.6151
R4537 vdd.n3102 vdd.n801 10.6151
R4538 vdd.n3097 vdd.n3096 10.6151
R4539 vdd.n3096 vdd.n3095 10.6151
R4540 vdd.n3074 vdd.n3035 10.6151
R4541 vdd.n3069 vdd.n3035 10.6151
R4542 vdd.n3069 vdd.n3068 10.6151
R4543 vdd.n3068 vdd.n3067 10.6151
R4544 vdd.n3067 vdd.n3037 10.6151
R4545 vdd.n3062 vdd.n3037 10.6151
R4546 vdd.n3062 vdd.n3061 10.6151
R4547 vdd.n3061 vdd.n3060 10.6151
R4548 vdd.n3060 vdd.n3040 10.6151
R4549 vdd.n3055 vdd.n3040 10.6151
R4550 vdd.n3055 vdd.n3054 10.6151
R4551 vdd.n3054 vdd.n3053 10.6151
R4552 vdd.n3053 vdd.n3043 10.6151
R4553 vdd.n3048 vdd.n3043 10.6151
R4554 vdd.n3048 vdd.n3047 10.6151
R4555 vdd.n3047 vdd.n753 10.6151
R4556 vdd.n3191 vdd.n753 10.6151
R4557 vdd.n3191 vdd.n754 10.6151
R4558 vdd.n757 vdd.n754 10.6151
R4559 vdd.n3184 vdd.n757 10.6151
R4560 vdd.n3184 vdd.n3183 10.6151
R4561 vdd.n3183 vdd.n3182 10.6151
R4562 vdd.n3182 vdd.n759 10.6151
R4563 vdd.n3177 vdd.n759 10.6151
R4564 vdd.n3177 vdd.n3176 10.6151
R4565 vdd.n3176 vdd.n3175 10.6151
R4566 vdd.n3175 vdd.n762 10.6151
R4567 vdd.n3170 vdd.n762 10.6151
R4568 vdd.n3170 vdd.n3169 10.6151
R4569 vdd.n3169 vdd.n3168 10.6151
R4570 vdd.n3168 vdd.n765 10.6151
R4571 vdd.n3163 vdd.n3162 10.6151
R4572 vdd.n3162 vdd.n3161 10.6151
R4573 vdd.n2924 vdd.n2923 10.6151
R4574 vdd.n2923 vdd.n2921 10.6151
R4575 vdd.n2921 vdd.n2920 10.6151
R4576 vdd.n2920 vdd.n2746 10.6151
R4577 vdd.n2820 vdd.n2746 10.6151
R4578 vdd.n2821 vdd.n2820 10.6151
R4579 vdd.n2823 vdd.n2821 10.6151
R4580 vdd.n2824 vdd.n2823 10.6151
R4581 vdd.n2904 vdd.n2824 10.6151
R4582 vdd.n2904 vdd.n2903 10.6151
R4583 vdd.n2903 vdd.n2902 10.6151
R4584 vdd.n2902 vdd.n2900 10.6151
R4585 vdd.n2900 vdd.n2899 10.6151
R4586 vdd.n2899 vdd.n2897 10.6151
R4587 vdd.n2897 vdd.n2896 10.6151
R4588 vdd.n2896 vdd.n2856 10.6151
R4589 vdd.n2856 vdd.n2855 10.6151
R4590 vdd.n2855 vdd.n2853 10.6151
R4591 vdd.n2853 vdd.n2852 10.6151
R4592 vdd.n2852 vdd.n2850 10.6151
R4593 vdd.n2850 vdd.n2849 10.6151
R4594 vdd.n2849 vdd.n2847 10.6151
R4595 vdd.n2847 vdd.n2846 10.6151
R4596 vdd.n2846 vdd.n2844 10.6151
R4597 vdd.n2844 vdd.n2843 10.6151
R4598 vdd.n2843 vdd.n2841 10.6151
R4599 vdd.n2841 vdd.n2840 10.6151
R4600 vdd.n2840 vdd.n2838 10.6151
R4601 vdd.n2838 vdd.n2837 10.6151
R4602 vdd.n2837 vdd.n2835 10.6151
R4603 vdd.n2835 vdd.n2834 10.6151
R4604 vdd.n2834 vdd.n2832 10.6151
R4605 vdd.n2832 vdd.n2831 10.6151
R4606 vdd.n2831 vdd.n2829 10.6151
R4607 vdd.n2829 vdd.n2828 10.6151
R4608 vdd.n2828 vdd.n2826 10.6151
R4609 vdd.n2826 vdd.n2825 10.6151
R4610 vdd.n2825 vdd.n771 10.6151
R4611 vdd.n2681 vdd.n913 10.6151
R4612 vdd.n2684 vdd.n2681 10.6151
R4613 vdd.n2685 vdd.n2684 10.6151
R4614 vdd.n2688 vdd.n2685 10.6151
R4615 vdd.n2689 vdd.n2688 10.6151
R4616 vdd.n2692 vdd.n2689 10.6151
R4617 vdd.n2693 vdd.n2692 10.6151
R4618 vdd.n2696 vdd.n2693 10.6151
R4619 vdd.n2697 vdd.n2696 10.6151
R4620 vdd.n2700 vdd.n2697 10.6151
R4621 vdd.n2701 vdd.n2700 10.6151
R4622 vdd.n2704 vdd.n2701 10.6151
R4623 vdd.n2705 vdd.n2704 10.6151
R4624 vdd.n2708 vdd.n2705 10.6151
R4625 vdd.n2709 vdd.n2708 10.6151
R4626 vdd.n2712 vdd.n2709 10.6151
R4627 vdd.n2713 vdd.n2712 10.6151
R4628 vdd.n2716 vdd.n2713 10.6151
R4629 vdd.n2717 vdd.n2716 10.6151
R4630 vdd.n2720 vdd.n2717 10.6151
R4631 vdd.n2721 vdd.n2720 10.6151
R4632 vdd.n2724 vdd.n2721 10.6151
R4633 vdd.n2725 vdd.n2724 10.6151
R4634 vdd.n2728 vdd.n2725 10.6151
R4635 vdd.n2729 vdd.n2728 10.6151
R4636 vdd.n2732 vdd.n2729 10.6151
R4637 vdd.n2733 vdd.n2732 10.6151
R4638 vdd.n2736 vdd.n2733 10.6151
R4639 vdd.n2737 vdd.n2736 10.6151
R4640 vdd.n2740 vdd.n2737 10.6151
R4641 vdd.n2741 vdd.n2740 10.6151
R4642 vdd.n2745 vdd.n2744 10.6151
R4643 vdd.n2925 vdd.n2745 10.6151
R4644 vdd.n2937 vdd.n2936 10.6151
R4645 vdd.n2938 vdd.n2937 10.6151
R4646 vdd.n2938 vdd.n903 10.6151
R4647 vdd.n2948 vdd.n903 10.6151
R4648 vdd.n2949 vdd.n2948 10.6151
R4649 vdd.n2950 vdd.n2949 10.6151
R4650 vdd.n2950 vdd.n891 10.6151
R4651 vdd.n2960 vdd.n891 10.6151
R4652 vdd.n2961 vdd.n2960 10.6151
R4653 vdd.n2962 vdd.n2961 10.6151
R4654 vdd.n2962 vdd.n880 10.6151
R4655 vdd.n2972 vdd.n880 10.6151
R4656 vdd.n2973 vdd.n2972 10.6151
R4657 vdd.n2974 vdd.n2973 10.6151
R4658 vdd.n2974 vdd.n868 10.6151
R4659 vdd.n2984 vdd.n868 10.6151
R4660 vdd.n2985 vdd.n2984 10.6151
R4661 vdd.n2986 vdd.n2985 10.6151
R4662 vdd.n2986 vdd.n857 10.6151
R4663 vdd.n2996 vdd.n857 10.6151
R4664 vdd.n2999 vdd.n2998 10.6151
R4665 vdd.n2999 vdd.n843 10.6151
R4666 vdd.n3009 vdd.n843 10.6151
R4667 vdd.n3010 vdd.n3009 10.6151
R4668 vdd.n3011 vdd.n3010 10.6151
R4669 vdd.n3011 vdd.n831 10.6151
R4670 vdd.n3021 vdd.n831 10.6151
R4671 vdd.n3022 vdd.n3021 10.6151
R4672 vdd.n3023 vdd.n3022 10.6151
R4673 vdd.n3023 vdd.n820 10.6151
R4674 vdd.n3033 vdd.n820 10.6151
R4675 vdd.n3034 vdd.n3033 10.6151
R4676 vdd.n3080 vdd.n3034 10.6151
R4677 vdd.n3080 vdd.n3079 10.6151
R4678 vdd.n3079 vdd.n3078 10.6151
R4679 vdd.n3078 vdd.n3077 10.6151
R4680 vdd.n3077 vdd.n3075 10.6151
R4681 vdd.n2387 vdd.n2386 10.6151
R4682 vdd.n2388 vdd.n2387 10.6151
R4683 vdd.n2388 vdd.n1067 10.6151
R4684 vdd.n2398 vdd.n1067 10.6151
R4685 vdd.n2399 vdd.n2398 10.6151
R4686 vdd.n2400 vdd.n2399 10.6151
R4687 vdd.n2400 vdd.n1055 10.6151
R4688 vdd.n2410 vdd.n1055 10.6151
R4689 vdd.n2411 vdd.n2410 10.6151
R4690 vdd.n2412 vdd.n2411 10.6151
R4691 vdd.n2412 vdd.n1043 10.6151
R4692 vdd.n2422 vdd.n1043 10.6151
R4693 vdd.n2423 vdd.n2422 10.6151
R4694 vdd.n2424 vdd.n2423 10.6151
R4695 vdd.n2424 vdd.n1030 10.6151
R4696 vdd.n2434 vdd.n1030 10.6151
R4697 vdd.n2435 vdd.n2434 10.6151
R4698 vdd.n2437 vdd.n1018 10.6151
R4699 vdd.n2447 vdd.n1018 10.6151
R4700 vdd.n2448 vdd.n2447 10.6151
R4701 vdd.n2449 vdd.n2448 10.6151
R4702 vdd.n2449 vdd.n1006 10.6151
R4703 vdd.n2459 vdd.n1006 10.6151
R4704 vdd.n2460 vdd.n2459 10.6151
R4705 vdd.n2461 vdd.n2460 10.6151
R4706 vdd.n2461 vdd.n995 10.6151
R4707 vdd.n2471 vdd.n995 10.6151
R4708 vdd.n2472 vdd.n2471 10.6151
R4709 vdd.n2473 vdd.n2472 10.6151
R4710 vdd.n2473 vdd.n984 10.6151
R4711 vdd.n2483 vdd.n984 10.6151
R4712 vdd.n2484 vdd.n2483 10.6151
R4713 vdd.n2487 vdd.n2484 10.6151
R4714 vdd.n2487 vdd.n2486 10.6151
R4715 vdd.n2486 vdd.n2485 10.6151
R4716 vdd.n2485 vdd.n967 10.6151
R4717 vdd.n2569 vdd.n967 10.6151
R4718 vdd.n2568 vdd.n2567 10.6151
R4719 vdd.n2567 vdd.n2564 10.6151
R4720 vdd.n2564 vdd.n2563 10.6151
R4721 vdd.n2563 vdd.n2560 10.6151
R4722 vdd.n2560 vdd.n2559 10.6151
R4723 vdd.n2559 vdd.n2556 10.6151
R4724 vdd.n2556 vdd.n2555 10.6151
R4725 vdd.n2555 vdd.n2552 10.6151
R4726 vdd.n2552 vdd.n2551 10.6151
R4727 vdd.n2551 vdd.n2548 10.6151
R4728 vdd.n2548 vdd.n2547 10.6151
R4729 vdd.n2547 vdd.n2544 10.6151
R4730 vdd.n2544 vdd.n2543 10.6151
R4731 vdd.n2543 vdd.n2540 10.6151
R4732 vdd.n2540 vdd.n2539 10.6151
R4733 vdd.n2539 vdd.n2536 10.6151
R4734 vdd.n2536 vdd.n2535 10.6151
R4735 vdd.n2535 vdd.n2532 10.6151
R4736 vdd.n2532 vdd.n2531 10.6151
R4737 vdd.n2531 vdd.n2528 10.6151
R4738 vdd.n2528 vdd.n2527 10.6151
R4739 vdd.n2527 vdd.n2524 10.6151
R4740 vdd.n2524 vdd.n2523 10.6151
R4741 vdd.n2523 vdd.n2520 10.6151
R4742 vdd.n2520 vdd.n2519 10.6151
R4743 vdd.n2519 vdd.n2516 10.6151
R4744 vdd.n2516 vdd.n2515 10.6151
R4745 vdd.n2515 vdd.n2512 10.6151
R4746 vdd.n2512 vdd.n2511 10.6151
R4747 vdd.n2511 vdd.n2508 10.6151
R4748 vdd.n2508 vdd.n2507 10.6151
R4749 vdd.n2504 vdd.n2503 10.6151
R4750 vdd.n2503 vdd.n2501 10.6151
R4751 vdd.n2203 vdd.n2201 10.6151
R4752 vdd.n2204 vdd.n2203 10.6151
R4753 vdd.n2206 vdd.n2204 10.6151
R4754 vdd.n2207 vdd.n2206 10.6151
R4755 vdd.n2209 vdd.n2207 10.6151
R4756 vdd.n2210 vdd.n2209 10.6151
R4757 vdd.n2212 vdd.n2210 10.6151
R4758 vdd.n2213 vdd.n2212 10.6151
R4759 vdd.n2215 vdd.n2213 10.6151
R4760 vdd.n2216 vdd.n2215 10.6151
R4761 vdd.n2218 vdd.n2216 10.6151
R4762 vdd.n2219 vdd.n2218 10.6151
R4763 vdd.n2221 vdd.n2219 10.6151
R4764 vdd.n2222 vdd.n2221 10.6151
R4765 vdd.n2224 vdd.n2222 10.6151
R4766 vdd.n2225 vdd.n2224 10.6151
R4767 vdd.n2227 vdd.n2225 10.6151
R4768 vdd.n2228 vdd.n2227 10.6151
R4769 vdd.n2230 vdd.n2228 10.6151
R4770 vdd.n2231 vdd.n2230 10.6151
R4771 vdd.n2233 vdd.n2231 10.6151
R4772 vdd.n2234 vdd.n2233 10.6151
R4773 vdd.n2273 vdd.n2234 10.6151
R4774 vdd.n2273 vdd.n2272 10.6151
R4775 vdd.n2272 vdd.n2271 10.6151
R4776 vdd.n2271 vdd.n2269 10.6151
R4777 vdd.n2269 vdd.n2268 10.6151
R4778 vdd.n2268 vdd.n2266 10.6151
R4779 vdd.n2266 vdd.n2265 10.6151
R4780 vdd.n2265 vdd.n2242 10.6151
R4781 vdd.n2242 vdd.n2241 10.6151
R4782 vdd.n2241 vdd.n2239 10.6151
R4783 vdd.n2239 vdd.n2238 10.6151
R4784 vdd.n2238 vdd.n2236 10.6151
R4785 vdd.n2236 vdd.n2235 10.6151
R4786 vdd.n2235 vdd.n971 10.6151
R4787 vdd.n2499 vdd.n971 10.6151
R4788 vdd.n2500 vdd.n2499 10.6151
R4789 vdd.n2131 vdd.n1079 10.6151
R4790 vdd.n2136 vdd.n2131 10.6151
R4791 vdd.n2137 vdd.n2136 10.6151
R4792 vdd.n2138 vdd.n2137 10.6151
R4793 vdd.n2138 vdd.n2129 10.6151
R4794 vdd.n2144 vdd.n2129 10.6151
R4795 vdd.n2145 vdd.n2144 10.6151
R4796 vdd.n2146 vdd.n2145 10.6151
R4797 vdd.n2146 vdd.n2127 10.6151
R4798 vdd.n2152 vdd.n2127 10.6151
R4799 vdd.n2153 vdd.n2152 10.6151
R4800 vdd.n2154 vdd.n2153 10.6151
R4801 vdd.n2154 vdd.n2125 10.6151
R4802 vdd.n2160 vdd.n2125 10.6151
R4803 vdd.n2161 vdd.n2160 10.6151
R4804 vdd.n2162 vdd.n2161 10.6151
R4805 vdd.n2162 vdd.n2123 10.6151
R4806 vdd.n2168 vdd.n2123 10.6151
R4807 vdd.n2169 vdd.n2168 10.6151
R4808 vdd.n2170 vdd.n2169 10.6151
R4809 vdd.n2170 vdd.n1113 10.6151
R4810 vdd.n2176 vdd.n1113 10.6151
R4811 vdd.n2177 vdd.n2176 10.6151
R4812 vdd.n2178 vdd.n2177 10.6151
R4813 vdd.n2178 vdd.n1111 10.6151
R4814 vdd.n2184 vdd.n1111 10.6151
R4815 vdd.n2185 vdd.n2184 10.6151
R4816 vdd.n2186 vdd.n2185 10.6151
R4817 vdd.n2186 vdd.n1109 10.6151
R4818 vdd.n2192 vdd.n1109 10.6151
R4819 vdd.n2193 vdd.n2192 10.6151
R4820 vdd.n2195 vdd.n1105 10.6151
R4821 vdd.n2200 vdd.n1105 10.6151
R4822 vdd.t105 vdd.n1856 10.5435
R4823 vdd.n636 vdd.t107 10.5435
R4824 vdd.n304 vdd.n286 10.4732
R4825 vdd.n249 vdd.n231 10.4732
R4826 vdd.n206 vdd.n188 10.4732
R4827 vdd.n151 vdd.n133 10.4732
R4828 vdd.n109 vdd.n91 10.4732
R4829 vdd.n54 vdd.n36 10.4732
R4830 vdd.n1753 vdd.n1735 10.4732
R4831 vdd.n1808 vdd.n1790 10.4732
R4832 vdd.n1655 vdd.n1637 10.4732
R4833 vdd.n1710 vdd.n1692 10.4732
R4834 vdd.n1558 vdd.n1540 10.4732
R4835 vdd.n1613 vdd.n1595 10.4732
R4836 vdd.n1840 vdd.t220 10.3167
R4837 vdd.n3387 vdd.t119 10.3167
R4838 vdd.n2571 vdd.t175 10.2034
R4839 vdd.n2934 vdd.t159 10.2034
R4840 vdd.t2 vdd.n1184 10.09
R4841 vdd.n1892 vdd.t52 10.09
R4842 vdd.n3335 vdd.t26 10.09
R4843 vdd.n3468 vdd.t8 10.09
R4844 vdd.n2099 vdd.n1093 9.88581
R4845 vdd.n3125 vdd.n3124 9.88581
R4846 vdd.n3192 vdd.n3191 9.88581
R4847 vdd.n2123 vdd.n2122 9.88581
R4848 vdd.n1504 vdd.t17 9.86327
R4849 vdd.n3459 vdd.t101 9.86327
R4850 vdd.n303 vdd.n288 9.69747
R4851 vdd.n248 vdd.n233 9.69747
R4852 vdd.n205 vdd.n190 9.69747
R4853 vdd.n150 vdd.n135 9.69747
R4854 vdd.n108 vdd.n93 9.69747
R4855 vdd.n53 vdd.n38 9.69747
R4856 vdd.n1752 vdd.n1737 9.69747
R4857 vdd.n1807 vdd.n1792 9.69747
R4858 vdd.n1654 vdd.n1639 9.69747
R4859 vdd.n1709 vdd.n1694 9.69747
R4860 vdd.n1557 vdd.n1542 9.69747
R4861 vdd.n1612 vdd.n1597 9.69747
R4862 vdd.t21 vdd.n1478 9.63654
R4863 vdd.n3418 vdd.t210 9.63654
R4864 vdd.n319 vdd.n318 9.45567
R4865 vdd.n264 vdd.n263 9.45567
R4866 vdd.n221 vdd.n220 9.45567
R4867 vdd.n166 vdd.n165 9.45567
R4868 vdd.n124 vdd.n123 9.45567
R4869 vdd.n69 vdd.n68 9.45567
R4870 vdd.n1768 vdd.n1767 9.45567
R4871 vdd.n1823 vdd.n1822 9.45567
R4872 vdd.n1670 vdd.n1669 9.45567
R4873 vdd.n1725 vdd.n1724 9.45567
R4874 vdd.n1573 vdd.n1572 9.45567
R4875 vdd.n1628 vdd.n1627 9.45567
R4876 vdd.n2072 vdd.n1926 9.3005
R4877 vdd.n2071 vdd.n2070 9.3005
R4878 vdd.n1932 vdd.n1931 9.3005
R4879 vdd.n2065 vdd.n1936 9.3005
R4880 vdd.n2064 vdd.n1937 9.3005
R4881 vdd.n2063 vdd.n1938 9.3005
R4882 vdd.n1942 vdd.n1939 9.3005
R4883 vdd.n2058 vdd.n1943 9.3005
R4884 vdd.n2057 vdd.n1944 9.3005
R4885 vdd.n2056 vdd.n1945 9.3005
R4886 vdd.n1949 vdd.n1946 9.3005
R4887 vdd.n2051 vdd.n1950 9.3005
R4888 vdd.n2050 vdd.n1951 9.3005
R4889 vdd.n2049 vdd.n1952 9.3005
R4890 vdd.n1956 vdd.n1953 9.3005
R4891 vdd.n2044 vdd.n1957 9.3005
R4892 vdd.n2043 vdd.n1958 9.3005
R4893 vdd.n2042 vdd.n1959 9.3005
R4894 vdd.n1963 vdd.n1960 9.3005
R4895 vdd.n2037 vdd.n1964 9.3005
R4896 vdd.n2036 vdd.n1965 9.3005
R4897 vdd.n2035 vdd.n2034 9.3005
R4898 vdd.n2033 vdd.n1966 9.3005
R4899 vdd.n2032 vdd.n2031 9.3005
R4900 vdd.n1972 vdd.n1971 9.3005
R4901 vdd.n2026 vdd.n1976 9.3005
R4902 vdd.n2025 vdd.n1977 9.3005
R4903 vdd.n2024 vdd.n1978 9.3005
R4904 vdd.n1982 vdd.n1979 9.3005
R4905 vdd.n2019 vdd.n1983 9.3005
R4906 vdd.n2018 vdd.n1984 9.3005
R4907 vdd.n2017 vdd.n1985 9.3005
R4908 vdd.n1989 vdd.n1986 9.3005
R4909 vdd.n2012 vdd.n1990 9.3005
R4910 vdd.n2011 vdd.n1991 9.3005
R4911 vdd.n2010 vdd.n1992 9.3005
R4912 vdd.n1994 vdd.n1993 9.3005
R4913 vdd.n2005 vdd.n1115 9.3005
R4914 vdd.n2074 vdd.n2073 9.3005
R4915 vdd.n2098 vdd.n2097 9.3005
R4916 vdd.n1904 vdd.n1903 9.3005
R4917 vdd.n1909 vdd.n1907 9.3005
R4918 vdd.n2090 vdd.n1910 9.3005
R4919 vdd.n2089 vdd.n1911 9.3005
R4920 vdd.n2088 vdd.n1912 9.3005
R4921 vdd.n1916 vdd.n1913 9.3005
R4922 vdd.n2083 vdd.n1917 9.3005
R4923 vdd.n2082 vdd.n1918 9.3005
R4924 vdd.n2081 vdd.n1919 9.3005
R4925 vdd.n1923 vdd.n1920 9.3005
R4926 vdd.n2076 vdd.n1924 9.3005
R4927 vdd.n2075 vdd.n1925 9.3005
R4928 vdd.n2107 vdd.n1897 9.3005
R4929 vdd.n2109 vdd.n2108 9.3005
R4930 vdd.n1828 vdd.n1174 9.3005
R4931 vdd.n1830 vdd.n1829 9.3005
R4932 vdd.n1165 vdd.n1164 9.3005
R4933 vdd.n1843 vdd.n1842 9.3005
R4934 vdd.n1844 vdd.n1163 9.3005
R4935 vdd.n1846 vdd.n1845 9.3005
R4936 vdd.n1153 vdd.n1152 9.3005
R4937 vdd.n1860 vdd.n1859 9.3005
R4938 vdd.n1861 vdd.n1151 9.3005
R4939 vdd.n1863 vdd.n1862 9.3005
R4940 vdd.n1142 vdd.n1141 9.3005
R4941 vdd.n1877 vdd.n1876 9.3005
R4942 vdd.n1878 vdd.n1140 9.3005
R4943 vdd.n1880 vdd.n1879 9.3005
R4944 vdd.n1130 vdd.n1129 9.3005
R4945 vdd.n1895 vdd.n1894 9.3005
R4946 vdd.n1896 vdd.n1128 9.3005
R4947 vdd.n2111 vdd.n2110 9.3005
R4948 vdd.n295 vdd.n294 9.3005
R4949 vdd.n290 vdd.n289 9.3005
R4950 vdd.n301 vdd.n300 9.3005
R4951 vdd.n303 vdd.n302 9.3005
R4952 vdd.n286 vdd.n285 9.3005
R4953 vdd.n309 vdd.n308 9.3005
R4954 vdd.n311 vdd.n310 9.3005
R4955 vdd.n283 vdd.n280 9.3005
R4956 vdd.n318 vdd.n317 9.3005
R4957 vdd.n240 vdd.n239 9.3005
R4958 vdd.n235 vdd.n234 9.3005
R4959 vdd.n246 vdd.n245 9.3005
R4960 vdd.n248 vdd.n247 9.3005
R4961 vdd.n231 vdd.n230 9.3005
R4962 vdd.n254 vdd.n253 9.3005
R4963 vdd.n256 vdd.n255 9.3005
R4964 vdd.n228 vdd.n225 9.3005
R4965 vdd.n263 vdd.n262 9.3005
R4966 vdd.n197 vdd.n196 9.3005
R4967 vdd.n192 vdd.n191 9.3005
R4968 vdd.n203 vdd.n202 9.3005
R4969 vdd.n205 vdd.n204 9.3005
R4970 vdd.n188 vdd.n187 9.3005
R4971 vdd.n211 vdd.n210 9.3005
R4972 vdd.n213 vdd.n212 9.3005
R4973 vdd.n185 vdd.n182 9.3005
R4974 vdd.n220 vdd.n219 9.3005
R4975 vdd.n142 vdd.n141 9.3005
R4976 vdd.n137 vdd.n136 9.3005
R4977 vdd.n148 vdd.n147 9.3005
R4978 vdd.n150 vdd.n149 9.3005
R4979 vdd.n133 vdd.n132 9.3005
R4980 vdd.n156 vdd.n155 9.3005
R4981 vdd.n158 vdd.n157 9.3005
R4982 vdd.n130 vdd.n127 9.3005
R4983 vdd.n165 vdd.n164 9.3005
R4984 vdd.n100 vdd.n99 9.3005
R4985 vdd.n95 vdd.n94 9.3005
R4986 vdd.n106 vdd.n105 9.3005
R4987 vdd.n108 vdd.n107 9.3005
R4988 vdd.n91 vdd.n90 9.3005
R4989 vdd.n114 vdd.n113 9.3005
R4990 vdd.n116 vdd.n115 9.3005
R4991 vdd.n88 vdd.n85 9.3005
R4992 vdd.n123 vdd.n122 9.3005
R4993 vdd.n45 vdd.n44 9.3005
R4994 vdd.n40 vdd.n39 9.3005
R4995 vdd.n51 vdd.n50 9.3005
R4996 vdd.n53 vdd.n52 9.3005
R4997 vdd.n36 vdd.n35 9.3005
R4998 vdd.n59 vdd.n58 9.3005
R4999 vdd.n61 vdd.n60 9.3005
R5000 vdd.n33 vdd.n30 9.3005
R5001 vdd.n68 vdd.n67 9.3005
R5002 vdd.n3241 vdd.n3240 9.3005
R5003 vdd.n3242 vdd.n721 9.3005
R5004 vdd.n720 vdd.n718 9.3005
R5005 vdd.n3248 vdd.n717 9.3005
R5006 vdd.n3249 vdd.n716 9.3005
R5007 vdd.n3250 vdd.n715 9.3005
R5008 vdd.n714 vdd.n712 9.3005
R5009 vdd.n3256 vdd.n711 9.3005
R5010 vdd.n3257 vdd.n710 9.3005
R5011 vdd.n3258 vdd.n709 9.3005
R5012 vdd.n708 vdd.n706 9.3005
R5013 vdd.n3264 vdd.n705 9.3005
R5014 vdd.n3265 vdd.n704 9.3005
R5015 vdd.n3266 vdd.n703 9.3005
R5016 vdd.n702 vdd.n700 9.3005
R5017 vdd.n3272 vdd.n699 9.3005
R5018 vdd.n3273 vdd.n698 9.3005
R5019 vdd.n3274 vdd.n697 9.3005
R5020 vdd.n696 vdd.n694 9.3005
R5021 vdd.n3280 vdd.n693 9.3005
R5022 vdd.n3281 vdd.n692 9.3005
R5023 vdd.n3282 vdd.n691 9.3005
R5024 vdd.n690 vdd.n688 9.3005
R5025 vdd.n3288 vdd.n685 9.3005
R5026 vdd.n3289 vdd.n684 9.3005
R5027 vdd.n3290 vdd.n683 9.3005
R5028 vdd.n682 vdd.n680 9.3005
R5029 vdd.n3296 vdd.n679 9.3005
R5030 vdd.n3297 vdd.n678 9.3005
R5031 vdd.n3298 vdd.n677 9.3005
R5032 vdd.n676 vdd.n674 9.3005
R5033 vdd.n3304 vdd.n673 9.3005
R5034 vdd.n3305 vdd.n672 9.3005
R5035 vdd.n3306 vdd.n671 9.3005
R5036 vdd.n670 vdd.n668 9.3005
R5037 vdd.n3311 vdd.n667 9.3005
R5038 vdd.n3321 vdd.n661 9.3005
R5039 vdd.n3323 vdd.n3322 9.3005
R5040 vdd.n652 vdd.n651 9.3005
R5041 vdd.n3338 vdd.n3337 9.3005
R5042 vdd.n3339 vdd.n650 9.3005
R5043 vdd.n3341 vdd.n3340 9.3005
R5044 vdd.n640 vdd.n639 9.3005
R5045 vdd.n3354 vdd.n3353 9.3005
R5046 vdd.n3355 vdd.n638 9.3005
R5047 vdd.n3357 vdd.n3356 9.3005
R5048 vdd.n628 vdd.n627 9.3005
R5049 vdd.n3371 vdd.n3370 9.3005
R5050 vdd.n3372 vdd.n626 9.3005
R5051 vdd.n3374 vdd.n3373 9.3005
R5052 vdd.n617 vdd.n616 9.3005
R5053 vdd.n3390 vdd.n3389 9.3005
R5054 vdd.n3391 vdd.n615 9.3005
R5055 vdd.n3393 vdd.n3392 9.3005
R5056 vdd.n324 vdd.n322 9.3005
R5057 vdd.n3325 vdd.n3324 9.3005
R5058 vdd.n3472 vdd.n3471 9.3005
R5059 vdd.n325 vdd.n323 9.3005
R5060 vdd.n3465 vdd.n334 9.3005
R5061 vdd.n3464 vdd.n335 9.3005
R5062 vdd.n3463 vdd.n336 9.3005
R5063 vdd.n343 vdd.n337 9.3005
R5064 vdd.n3457 vdd.n344 9.3005
R5065 vdd.n3456 vdd.n345 9.3005
R5066 vdd.n3455 vdd.n346 9.3005
R5067 vdd.n354 vdd.n347 9.3005
R5068 vdd.n3449 vdd.n355 9.3005
R5069 vdd.n3448 vdd.n356 9.3005
R5070 vdd.n3447 vdd.n357 9.3005
R5071 vdd.n365 vdd.n358 9.3005
R5072 vdd.n3441 vdd.n366 9.3005
R5073 vdd.n3440 vdd.n367 9.3005
R5074 vdd.n3439 vdd.n368 9.3005
R5075 vdd.n443 vdd.n369 9.3005
R5076 vdd.n447 vdd.n442 9.3005
R5077 vdd.n451 vdd.n450 9.3005
R5078 vdd.n452 vdd.n441 9.3005
R5079 vdd.n456 vdd.n453 9.3005
R5080 vdd.n457 vdd.n440 9.3005
R5081 vdd.n461 vdd.n460 9.3005
R5082 vdd.n462 vdd.n439 9.3005
R5083 vdd.n466 vdd.n463 9.3005
R5084 vdd.n467 vdd.n438 9.3005
R5085 vdd.n471 vdd.n470 9.3005
R5086 vdd.n472 vdd.n437 9.3005
R5087 vdd.n476 vdd.n473 9.3005
R5088 vdd.n477 vdd.n436 9.3005
R5089 vdd.n481 vdd.n480 9.3005
R5090 vdd.n482 vdd.n435 9.3005
R5091 vdd.n486 vdd.n483 9.3005
R5092 vdd.n487 vdd.n434 9.3005
R5093 vdd.n491 vdd.n490 9.3005
R5094 vdd.n492 vdd.n433 9.3005
R5095 vdd.n496 vdd.n493 9.3005
R5096 vdd.n497 vdd.n430 9.3005
R5097 vdd.n501 vdd.n500 9.3005
R5098 vdd.n502 vdd.n429 9.3005
R5099 vdd.n506 vdd.n503 9.3005
R5100 vdd.n507 vdd.n428 9.3005
R5101 vdd.n511 vdd.n510 9.3005
R5102 vdd.n512 vdd.n427 9.3005
R5103 vdd.n516 vdd.n513 9.3005
R5104 vdd.n517 vdd.n426 9.3005
R5105 vdd.n521 vdd.n520 9.3005
R5106 vdd.n522 vdd.n425 9.3005
R5107 vdd.n526 vdd.n523 9.3005
R5108 vdd.n527 vdd.n424 9.3005
R5109 vdd.n531 vdd.n530 9.3005
R5110 vdd.n532 vdd.n423 9.3005
R5111 vdd.n536 vdd.n533 9.3005
R5112 vdd.n537 vdd.n422 9.3005
R5113 vdd.n541 vdd.n540 9.3005
R5114 vdd.n542 vdd.n421 9.3005
R5115 vdd.n546 vdd.n543 9.3005
R5116 vdd.n547 vdd.n418 9.3005
R5117 vdd.n551 vdd.n550 9.3005
R5118 vdd.n552 vdd.n417 9.3005
R5119 vdd.n556 vdd.n553 9.3005
R5120 vdd.n557 vdd.n416 9.3005
R5121 vdd.n561 vdd.n560 9.3005
R5122 vdd.n562 vdd.n415 9.3005
R5123 vdd.n566 vdd.n563 9.3005
R5124 vdd.n567 vdd.n414 9.3005
R5125 vdd.n571 vdd.n570 9.3005
R5126 vdd.n572 vdd.n413 9.3005
R5127 vdd.n576 vdd.n573 9.3005
R5128 vdd.n577 vdd.n412 9.3005
R5129 vdd.n581 vdd.n580 9.3005
R5130 vdd.n582 vdd.n411 9.3005
R5131 vdd.n586 vdd.n583 9.3005
R5132 vdd.n587 vdd.n410 9.3005
R5133 vdd.n591 vdd.n590 9.3005
R5134 vdd.n592 vdd.n409 9.3005
R5135 vdd.n596 vdd.n593 9.3005
R5136 vdd.n598 vdd.n408 9.3005
R5137 vdd.n600 vdd.n599 9.3005
R5138 vdd.n3432 vdd.n3431 9.3005
R5139 vdd.n446 vdd.n444 9.3005
R5140 vdd.n3331 vdd.n655 9.3005
R5141 vdd.n3333 vdd.n3332 9.3005
R5142 vdd.n646 vdd.n645 9.3005
R5143 vdd.n3346 vdd.n3345 9.3005
R5144 vdd.n3347 vdd.n644 9.3005
R5145 vdd.n3349 vdd.n3348 9.3005
R5146 vdd.n633 vdd.n632 9.3005
R5147 vdd.n3362 vdd.n3361 9.3005
R5148 vdd.n3363 vdd.n631 9.3005
R5149 vdd.n3365 vdd.n3364 9.3005
R5150 vdd.n622 vdd.n621 9.3005
R5151 vdd.n3379 vdd.n3378 9.3005
R5152 vdd.n3380 vdd.n620 9.3005
R5153 vdd.n3385 vdd.n3381 9.3005
R5154 vdd.n3384 vdd.n3383 9.3005
R5155 vdd.n3382 vdd.n610 9.3005
R5156 vdd.n3398 vdd.n611 9.3005
R5157 vdd.n3399 vdd.n609 9.3005
R5158 vdd.n3401 vdd.n3400 9.3005
R5159 vdd.n3402 vdd.n608 9.3005
R5160 vdd.n3405 vdd.n3403 9.3005
R5161 vdd.n3406 vdd.n607 9.3005
R5162 vdd.n3408 vdd.n3407 9.3005
R5163 vdd.n3409 vdd.n606 9.3005
R5164 vdd.n3412 vdd.n3410 9.3005
R5165 vdd.n3413 vdd.n605 9.3005
R5166 vdd.n3415 vdd.n3414 9.3005
R5167 vdd.n3416 vdd.n604 9.3005
R5168 vdd.n3420 vdd.n3417 9.3005
R5169 vdd.n3421 vdd.n603 9.3005
R5170 vdd.n3423 vdd.n3422 9.3005
R5171 vdd.n3424 vdd.n602 9.3005
R5172 vdd.n3427 vdd.n3425 9.3005
R5173 vdd.n3428 vdd.n601 9.3005
R5174 vdd.n3430 vdd.n3429 9.3005
R5175 vdd.n3330 vdd.n3329 9.3005
R5176 vdd.n3194 vdd.n656 9.3005
R5177 vdd.n3199 vdd.n3193 9.3005
R5178 vdd.n3209 vdd.n748 9.3005
R5179 vdd.n3210 vdd.n747 9.3005
R5180 vdd.n746 vdd.n744 9.3005
R5181 vdd.n3216 vdd.n743 9.3005
R5182 vdd.n3217 vdd.n742 9.3005
R5183 vdd.n3218 vdd.n741 9.3005
R5184 vdd.n740 vdd.n738 9.3005
R5185 vdd.n3224 vdd.n737 9.3005
R5186 vdd.n3225 vdd.n736 9.3005
R5187 vdd.n3226 vdd.n735 9.3005
R5188 vdd.n734 vdd.n732 9.3005
R5189 vdd.n3231 vdd.n731 9.3005
R5190 vdd.n3232 vdd.n730 9.3005
R5191 vdd.n726 vdd.n725 9.3005
R5192 vdd.n3238 vdd.n3237 9.3005
R5193 vdd.n3239 vdd.n722 9.3005
R5194 vdd.n2121 vdd.n2120 9.3005
R5195 vdd.n2116 vdd.n1118 9.3005
R5196 vdd.n1460 vdd.n1459 9.3005
R5197 vdd.n1216 vdd.n1215 9.3005
R5198 vdd.n1473 vdd.n1472 9.3005
R5199 vdd.n1474 vdd.n1214 9.3005
R5200 vdd.n1476 vdd.n1475 9.3005
R5201 vdd.n1204 vdd.n1203 9.3005
R5202 vdd.n1490 vdd.n1489 9.3005
R5203 vdd.n1491 vdd.n1202 9.3005
R5204 vdd.n1493 vdd.n1492 9.3005
R5205 vdd.n1194 vdd.n1193 9.3005
R5206 vdd.n1507 vdd.n1506 9.3005
R5207 vdd.n1508 vdd.n1192 9.3005
R5208 vdd.n1510 vdd.n1509 9.3005
R5209 vdd.n1181 vdd.n1180 9.3005
R5210 vdd.n1523 vdd.n1522 9.3005
R5211 vdd.n1524 vdd.n1179 9.3005
R5212 vdd.n1526 vdd.n1525 9.3005
R5213 vdd.n1170 vdd.n1169 9.3005
R5214 vdd.n1835 vdd.n1834 9.3005
R5215 vdd.n1836 vdd.n1168 9.3005
R5216 vdd.n1838 vdd.n1837 9.3005
R5217 vdd.n1159 vdd.n1158 9.3005
R5218 vdd.n1851 vdd.n1850 9.3005
R5219 vdd.n1852 vdd.n1157 9.3005
R5220 vdd.n1854 vdd.n1853 9.3005
R5221 vdd.n1147 vdd.n1146 9.3005
R5222 vdd.n1868 vdd.n1867 9.3005
R5223 vdd.n1869 vdd.n1145 9.3005
R5224 vdd.n1871 vdd.n1870 9.3005
R5225 vdd.n1137 vdd.n1136 9.3005
R5226 vdd.n1885 vdd.n1884 9.3005
R5227 vdd.n1886 vdd.n1134 9.3005
R5228 vdd.n1890 vdd.n1889 9.3005
R5229 vdd.n1888 vdd.n1135 9.3005
R5230 vdd.n1887 vdd.n1123 9.3005
R5231 vdd.n1458 vdd.n1226 9.3005
R5232 vdd.n1351 vdd.n1227 9.3005
R5233 vdd.n1353 vdd.n1352 9.3005
R5234 vdd.n1354 vdd.n1346 9.3005
R5235 vdd.n1356 vdd.n1355 9.3005
R5236 vdd.n1357 vdd.n1345 9.3005
R5237 vdd.n1359 vdd.n1358 9.3005
R5238 vdd.n1360 vdd.n1340 9.3005
R5239 vdd.n1362 vdd.n1361 9.3005
R5240 vdd.n1363 vdd.n1339 9.3005
R5241 vdd.n1365 vdd.n1364 9.3005
R5242 vdd.n1366 vdd.n1334 9.3005
R5243 vdd.n1368 vdd.n1367 9.3005
R5244 vdd.n1369 vdd.n1333 9.3005
R5245 vdd.n1371 vdd.n1370 9.3005
R5246 vdd.n1372 vdd.n1328 9.3005
R5247 vdd.n1374 vdd.n1373 9.3005
R5248 vdd.n1375 vdd.n1327 9.3005
R5249 vdd.n1377 vdd.n1376 9.3005
R5250 vdd.n1378 vdd.n1322 9.3005
R5251 vdd.n1380 vdd.n1379 9.3005
R5252 vdd.n1381 vdd.n1321 9.3005
R5253 vdd.n1386 vdd.n1382 9.3005
R5254 vdd.n1387 vdd.n1317 9.3005
R5255 vdd.n1389 vdd.n1388 9.3005
R5256 vdd.n1390 vdd.n1316 9.3005
R5257 vdd.n1392 vdd.n1391 9.3005
R5258 vdd.n1393 vdd.n1311 9.3005
R5259 vdd.n1395 vdd.n1394 9.3005
R5260 vdd.n1396 vdd.n1310 9.3005
R5261 vdd.n1398 vdd.n1397 9.3005
R5262 vdd.n1399 vdd.n1305 9.3005
R5263 vdd.n1401 vdd.n1400 9.3005
R5264 vdd.n1402 vdd.n1304 9.3005
R5265 vdd.n1404 vdd.n1403 9.3005
R5266 vdd.n1405 vdd.n1299 9.3005
R5267 vdd.n1407 vdd.n1406 9.3005
R5268 vdd.n1408 vdd.n1298 9.3005
R5269 vdd.n1410 vdd.n1409 9.3005
R5270 vdd.n1411 vdd.n1293 9.3005
R5271 vdd.n1413 vdd.n1412 9.3005
R5272 vdd.n1414 vdd.n1292 9.3005
R5273 vdd.n1416 vdd.n1415 9.3005
R5274 vdd.n1417 vdd.n1289 9.3005
R5275 vdd.n1423 vdd.n1422 9.3005
R5276 vdd.n1424 vdd.n1288 9.3005
R5277 vdd.n1426 vdd.n1425 9.3005
R5278 vdd.n1427 vdd.n1283 9.3005
R5279 vdd.n1429 vdd.n1428 9.3005
R5280 vdd.n1430 vdd.n1282 9.3005
R5281 vdd.n1432 vdd.n1431 9.3005
R5282 vdd.n1433 vdd.n1277 9.3005
R5283 vdd.n1435 vdd.n1434 9.3005
R5284 vdd.n1436 vdd.n1276 9.3005
R5285 vdd.n1438 vdd.n1437 9.3005
R5286 vdd.n1439 vdd.n1271 9.3005
R5287 vdd.n1441 vdd.n1440 9.3005
R5288 vdd.n1442 vdd.n1270 9.3005
R5289 vdd.n1444 vdd.n1443 9.3005
R5290 vdd.n1445 vdd.n1266 9.3005
R5291 vdd.n1447 vdd.n1446 9.3005
R5292 vdd.n1448 vdd.n1265 9.3005
R5293 vdd.n1450 vdd.n1449 9.3005
R5294 vdd.n1451 vdd.n1264 9.3005
R5295 vdd.n1457 vdd.n1456 9.3005
R5296 vdd.n1465 vdd.n1464 9.3005
R5297 vdd.n1466 vdd.n1220 9.3005
R5298 vdd.n1468 vdd.n1467 9.3005
R5299 vdd.n1210 vdd.n1209 9.3005
R5300 vdd.n1482 vdd.n1481 9.3005
R5301 vdd.n1483 vdd.n1208 9.3005
R5302 vdd.n1485 vdd.n1484 9.3005
R5303 vdd.n1199 vdd.n1198 9.3005
R5304 vdd.n1499 vdd.n1498 9.3005
R5305 vdd.n1500 vdd.n1197 9.3005
R5306 vdd.n1502 vdd.n1501 9.3005
R5307 vdd.n1188 vdd.n1187 9.3005
R5308 vdd.n1515 vdd.n1514 9.3005
R5309 vdd.n1516 vdd.n1186 9.3005
R5310 vdd.n1518 vdd.n1517 9.3005
R5311 vdd.n1176 vdd.n1175 9.3005
R5312 vdd.n1532 vdd.n1531 9.3005
R5313 vdd.n1222 vdd.n1221 9.3005
R5314 vdd.n1744 vdd.n1743 9.3005
R5315 vdd.n1739 vdd.n1738 9.3005
R5316 vdd.n1750 vdd.n1749 9.3005
R5317 vdd.n1752 vdd.n1751 9.3005
R5318 vdd.n1735 vdd.n1734 9.3005
R5319 vdd.n1758 vdd.n1757 9.3005
R5320 vdd.n1760 vdd.n1759 9.3005
R5321 vdd.n1732 vdd.n1729 9.3005
R5322 vdd.n1767 vdd.n1766 9.3005
R5323 vdd.n1799 vdd.n1798 9.3005
R5324 vdd.n1794 vdd.n1793 9.3005
R5325 vdd.n1805 vdd.n1804 9.3005
R5326 vdd.n1807 vdd.n1806 9.3005
R5327 vdd.n1790 vdd.n1789 9.3005
R5328 vdd.n1813 vdd.n1812 9.3005
R5329 vdd.n1815 vdd.n1814 9.3005
R5330 vdd.n1787 vdd.n1784 9.3005
R5331 vdd.n1822 vdd.n1821 9.3005
R5332 vdd.n1646 vdd.n1645 9.3005
R5333 vdd.n1641 vdd.n1640 9.3005
R5334 vdd.n1652 vdd.n1651 9.3005
R5335 vdd.n1654 vdd.n1653 9.3005
R5336 vdd.n1637 vdd.n1636 9.3005
R5337 vdd.n1660 vdd.n1659 9.3005
R5338 vdd.n1662 vdd.n1661 9.3005
R5339 vdd.n1634 vdd.n1631 9.3005
R5340 vdd.n1669 vdd.n1668 9.3005
R5341 vdd.n1701 vdd.n1700 9.3005
R5342 vdd.n1696 vdd.n1695 9.3005
R5343 vdd.n1707 vdd.n1706 9.3005
R5344 vdd.n1709 vdd.n1708 9.3005
R5345 vdd.n1692 vdd.n1691 9.3005
R5346 vdd.n1715 vdd.n1714 9.3005
R5347 vdd.n1717 vdd.n1716 9.3005
R5348 vdd.n1689 vdd.n1686 9.3005
R5349 vdd.n1724 vdd.n1723 9.3005
R5350 vdd.n1549 vdd.n1548 9.3005
R5351 vdd.n1544 vdd.n1543 9.3005
R5352 vdd.n1555 vdd.n1554 9.3005
R5353 vdd.n1557 vdd.n1556 9.3005
R5354 vdd.n1540 vdd.n1539 9.3005
R5355 vdd.n1563 vdd.n1562 9.3005
R5356 vdd.n1565 vdd.n1564 9.3005
R5357 vdd.n1537 vdd.n1534 9.3005
R5358 vdd.n1572 vdd.n1571 9.3005
R5359 vdd.n1604 vdd.n1603 9.3005
R5360 vdd.n1599 vdd.n1598 9.3005
R5361 vdd.n1610 vdd.n1609 9.3005
R5362 vdd.n1612 vdd.n1611 9.3005
R5363 vdd.n1595 vdd.n1594 9.3005
R5364 vdd.n1618 vdd.n1617 9.3005
R5365 vdd.n1620 vdd.n1619 9.3005
R5366 vdd.n1592 vdd.n1589 9.3005
R5367 vdd.n1627 vdd.n1626 9.3005
R5368 vdd.n1478 vdd.t10 9.18308
R5369 vdd.n3418 vdd.t111 9.18308
R5370 vdd.n1504 vdd.t114 8.95635
R5371 vdd.t124 vdd.n3459 8.95635
R5372 vdd.n300 vdd.n299 8.92171
R5373 vdd.n245 vdd.n244 8.92171
R5374 vdd.n202 vdd.n201 8.92171
R5375 vdd.n147 vdd.n146 8.92171
R5376 vdd.n105 vdd.n104 8.92171
R5377 vdd.n50 vdd.n49 8.92171
R5378 vdd.n1749 vdd.n1748 8.92171
R5379 vdd.n1804 vdd.n1803 8.92171
R5380 vdd.n1651 vdd.n1650 8.92171
R5381 vdd.n1706 vdd.n1705 8.92171
R5382 vdd.n1554 vdd.n1553 8.92171
R5383 vdd.n1609 vdd.n1608 8.92171
R5384 vdd.n223 vdd.n125 8.81535
R5385 vdd.n1727 vdd.n1629 8.81535
R5386 vdd.n1184 vdd.t6 8.72962
R5387 vdd.t213 vdd.n3468 8.72962
R5388 vdd.n1840 vdd.t0 8.50289
R5389 vdd.n3387 vdd.t181 8.50289
R5390 vdd.n28 vdd.n14 8.42249
R5391 vdd.n1856 vdd.t185 8.27616
R5392 vdd.t223 vdd.n636 8.27616
R5393 vdd.n3474 vdd.n3473 8.16225
R5394 vdd.n1827 vdd.n1826 8.16225
R5395 vdd.n296 vdd.n290 8.14595
R5396 vdd.n241 vdd.n235 8.14595
R5397 vdd.n198 vdd.n192 8.14595
R5398 vdd.n143 vdd.n137 8.14595
R5399 vdd.n101 vdd.n95 8.14595
R5400 vdd.n46 vdd.n40 8.14595
R5401 vdd.n1745 vdd.n1739 8.14595
R5402 vdd.n1800 vdd.n1794 8.14595
R5403 vdd.n1647 vdd.n1641 8.14595
R5404 vdd.n1702 vdd.n1696 8.14595
R5405 vdd.n1550 vdd.n1544 8.14595
R5406 vdd.n1605 vdd.n1599 8.14595
R5407 vdd.t56 vdd.n1218 7.8227
R5408 vdd.t38 vdd.n363 7.8227
R5409 vdd.n2384 vdd.n1075 7.70933
R5410 vdd.n2390 vdd.n1075 7.70933
R5411 vdd.n2396 vdd.n1069 7.70933
R5412 vdd.n2396 vdd.n1063 7.70933
R5413 vdd.n2402 vdd.n1063 7.70933
R5414 vdd.n2402 vdd.n1057 7.70933
R5415 vdd.n2408 vdd.n1057 7.70933
R5416 vdd.n2414 vdd.n1051 7.70933
R5417 vdd.n2420 vdd.n1045 7.70933
R5418 vdd.n2426 vdd.n1038 7.70933
R5419 vdd.n2426 vdd.n1041 7.70933
R5420 vdd.n2432 vdd.n1034 7.70933
R5421 vdd.n2439 vdd.n1020 7.70933
R5422 vdd.n2445 vdd.n1020 7.70933
R5423 vdd.n2451 vdd.n1014 7.70933
R5424 vdd.n2457 vdd.n1010 7.70933
R5425 vdd.n2463 vdd.n1004 7.70933
R5426 vdd.n2481 vdd.n986 7.70933
R5427 vdd.n2481 vdd.n979 7.70933
R5428 vdd.n2489 vdd.n979 7.70933
R5429 vdd.n2571 vdd.n963 7.70933
R5430 vdd.n2934 vdd.n917 7.70933
R5431 vdd.n2946 vdd.n898 7.70933
R5432 vdd.n2952 vdd.n898 7.70933
R5433 vdd.n2952 vdd.n901 7.70933
R5434 vdd.n2970 vdd.n882 7.70933
R5435 vdd.n2976 vdd.n876 7.70933
R5436 vdd.n2982 vdd.n872 7.70933
R5437 vdd.n2988 vdd.n859 7.70933
R5438 vdd.n2994 vdd.n859 7.70933
R5439 vdd.n3001 vdd.n852 7.70933
R5440 vdd.n3007 vdd.n845 7.70933
R5441 vdd.n3007 vdd.n848 7.70933
R5442 vdd.n3013 vdd.n841 7.70933
R5443 vdd.n3019 vdd.n835 7.70933
R5444 vdd.n3025 vdd.n822 7.70933
R5445 vdd.n3031 vdd.n822 7.70933
R5446 vdd.n3031 vdd.n814 7.70933
R5447 vdd.n3082 vdd.n814 7.70933
R5448 vdd.n3082 vdd.n817 7.70933
R5449 vdd.n3088 vdd.n774 7.70933
R5450 vdd.n3158 vdd.n774 7.70933
R5451 vdd.t178 vdd.n1051 7.59597
R5452 vdd.n2263 vdd.t130 7.59597
R5453 vdd.n2906 vdd.t133 7.59597
R5454 vdd.n835 vdd.t157 7.59597
R5455 vdd.n295 vdd.n292 7.3702
R5456 vdd.n240 vdd.n237 7.3702
R5457 vdd.n197 vdd.n194 7.3702
R5458 vdd.n142 vdd.n139 7.3702
R5459 vdd.n100 vdd.n97 7.3702
R5460 vdd.n45 vdd.n42 7.3702
R5461 vdd.n1744 vdd.n1741 7.3702
R5462 vdd.n1799 vdd.n1796 7.3702
R5463 vdd.n1646 vdd.n1643 7.3702
R5464 vdd.n1701 vdd.n1698 7.3702
R5465 vdd.n1549 vdd.n1546 7.3702
R5466 vdd.n1604 vdd.n1601 7.3702
R5467 vdd.n1387 vdd.n1386 6.98232
R5468 vdd.n2036 vdd.n2035 6.98232
R5469 vdd.n547 vdd.n546 6.98232
R5470 vdd.n3242 vdd.n3241 6.98232
R5471 vdd.n1874 vdd.t103 6.91577
R5472 vdd.n2420 vdd.t141 6.91577
R5473 vdd.n3013 vdd.t166 6.91577
R5474 vdd.n3351 vdd.t121 6.91577
R5475 vdd.n2998 vdd.n2997 6.86879
R5476 vdd.n2436 vdd.n2435 6.86879
R5477 vdd.n2496 vdd.t173 6.80241
R5478 vdd.n2940 vdd.t161 6.80241
R5479 vdd.t4 vdd.n1155 6.68904
R5480 vdd.n3367 vdd.t183 6.68904
R5481 vdd.n1832 vdd.t204 6.46231
R5482 vdd.n3395 vdd.t109 6.46231
R5483 vdd.n2263 vdd.t131 6.34895
R5484 vdd.n2906 vdd.t171 6.34895
R5485 vdd.n3474 vdd.n321 6.32949
R5486 vdd.n1826 vdd.n1825 6.32949
R5487 vdd.t199 vdd.n1183 6.23558
R5488 vdd.t15 vdd.n332 6.23558
R5489 vdd.n1496 vdd.t12 6.00885
R5490 vdd.t144 vdd.n1014 6.00885
R5491 vdd.n872 vdd.t149 6.00885
R5492 vdd.n3453 vdd.t19 6.00885
R5493 vdd.n296 vdd.n295 5.81868
R5494 vdd.n241 vdd.n240 5.81868
R5495 vdd.n198 vdd.n197 5.81868
R5496 vdd.n143 vdd.n142 5.81868
R5497 vdd.n101 vdd.n100 5.81868
R5498 vdd.n46 vdd.n45 5.81868
R5499 vdd.n1745 vdd.n1744 5.81868
R5500 vdd.n1800 vdd.n1799 5.81868
R5501 vdd.n1647 vdd.n1646 5.81868
R5502 vdd.n1702 vdd.n1701 5.81868
R5503 vdd.n1550 vdd.n1549 5.81868
R5504 vdd.n1605 vdd.n1604 5.81868
R5505 vdd.n2579 vdd.n2578 5.77611
R5506 vdd.n2319 vdd.n2318 5.77611
R5507 vdd.n2808 vdd.n2807 5.77611
R5508 vdd.n3097 vdd.n806 5.77611
R5509 vdd.n3163 vdd.n770 5.77611
R5510 vdd.n2744 vdd.n2680 5.77611
R5511 vdd.n2504 vdd.n970 5.77611
R5512 vdd.n2195 vdd.n2194 5.77611
R5513 vdd.n1456 vdd.n1230 5.62474
R5514 vdd.n2119 vdd.n2116 5.62474
R5515 vdd.n3432 vdd.n407 5.62474
R5516 vdd.n3197 vdd.n3194 5.62474
R5517 vdd.n2457 vdd.t169 5.44203
R5518 vdd.n2976 vdd.t145 5.44203
R5519 vdd.n1206 vdd.t12 5.32866
R5520 vdd.t19 vdd.n3452 5.32866
R5521 vdd.n1512 vdd.t199 5.10193
R5522 vdd.n2432 vdd.t158 5.10193
R5523 vdd.n2451 vdd.t177 5.10193
R5524 vdd.n2982 vdd.t167 5.10193
R5525 vdd.n3001 vdd.t136 5.10193
R5526 vdd.n3461 vdd.t15 5.10193
R5527 vdd.n299 vdd.n290 5.04292
R5528 vdd.n244 vdd.n235 5.04292
R5529 vdd.n201 vdd.n192 5.04292
R5530 vdd.n146 vdd.n137 5.04292
R5531 vdd.n104 vdd.n95 5.04292
R5532 vdd.n49 vdd.n40 5.04292
R5533 vdd.n1748 vdd.n1739 5.04292
R5534 vdd.n1803 vdd.n1794 5.04292
R5535 vdd.n1650 vdd.n1641 5.04292
R5536 vdd.n1705 vdd.n1696 5.04292
R5537 vdd.n1553 vdd.n1544 5.04292
R5538 vdd.n1608 vdd.n1599 5.04292
R5539 vdd.n1034 vdd.t86 4.98857
R5540 vdd.t45 vdd.n852 4.98857
R5541 vdd.n1528 vdd.t204 4.8752
R5542 vdd.t34 vdd.n1069 4.8752
R5543 vdd.t139 vdd.t150 4.8752
R5544 vdd.n2251 vdd.t72 4.8752
R5545 vdd.n2918 vdd.t76 4.8752
R5546 vdd.t179 vdd.t129 4.8752
R5547 vdd.n817 vdd.t30 4.8752
R5548 vdd.t109 vdd.n328 4.8752
R5549 vdd.n2580 vdd.n2579 4.83952
R5550 vdd.n2320 vdd.n2319 4.83952
R5551 vdd.n2807 vdd.n2806 4.83952
R5552 vdd.n806 vdd.n801 4.83952
R5553 vdd.n770 vdd.n765 4.83952
R5554 vdd.n2741 vdd.n2680 4.83952
R5555 vdd.n2507 vdd.n970 4.83952
R5556 vdd.n2194 vdd.n2193 4.83952
R5557 vdd.n2475 vdd.t164 4.76184
R5558 vdd.n2958 vdd.t153 4.76184
R5559 vdd.n2004 vdd.n1116 4.74817
R5560 vdd.n1999 vdd.n1117 4.74817
R5561 vdd.n1901 vdd.n1898 4.74817
R5562 vdd.n2100 vdd.n1902 4.74817
R5563 vdd.n2102 vdd.n1901 4.74817
R5564 vdd.n2101 vdd.n2100 4.74817
R5565 vdd.n664 vdd.n662 4.74817
R5566 vdd.n3312 vdd.n665 4.74817
R5567 vdd.n3315 vdd.n665 4.74817
R5568 vdd.n3316 vdd.n664 4.74817
R5569 vdd.n3204 vdd.n749 4.74817
R5570 vdd.n3200 vdd.n751 4.74817
R5571 vdd.n3203 vdd.n751 4.74817
R5572 vdd.n3208 vdd.n749 4.74817
R5573 vdd.n2000 vdd.n1116 4.74817
R5574 vdd.n1119 vdd.n1117 4.74817
R5575 vdd.n321 vdd.n320 4.7074
R5576 vdd.n223 vdd.n222 4.7074
R5577 vdd.n1825 vdd.n1824 4.7074
R5578 vdd.n1727 vdd.n1726 4.7074
R5579 vdd.n1848 vdd.t4 4.64847
R5580 vdd.n3376 vdd.t183 4.64847
R5581 vdd.n1149 vdd.t103 4.42174
R5582 vdd.t121 vdd.n635 4.42174
R5583 vdd.n2251 vdd.t147 4.30838
R5584 vdd.n2918 vdd.t134 4.30838
R5585 vdd.n300 vdd.n288 4.26717
R5586 vdd.n245 vdd.n233 4.26717
R5587 vdd.n202 vdd.n190 4.26717
R5588 vdd.n147 vdd.n135 4.26717
R5589 vdd.n105 vdd.n93 4.26717
R5590 vdd.n50 vdd.n38 4.26717
R5591 vdd.n1749 vdd.n1737 4.26717
R5592 vdd.n1804 vdd.n1792 4.26717
R5593 vdd.n1651 vdd.n1639 4.26717
R5594 vdd.n1706 vdd.n1694 4.26717
R5595 vdd.n1554 vdd.n1542 4.26717
R5596 vdd.n1609 vdd.n1597 4.26717
R5597 vdd.t140 vdd.n1045 4.19501
R5598 vdd.n1004 vdd.t152 4.19501
R5599 vdd.t168 vdd.n882 4.19501
R5600 vdd.n841 vdd.t163 4.19501
R5601 vdd.n321 vdd.n223 4.10845
R5602 vdd.n1825 vdd.n1727 4.10845
R5603 vdd.n277 vdd.t268 4.06363
R5604 vdd.n277 vdd.t196 4.06363
R5605 vdd.n275 vdd.t125 4.06363
R5606 vdd.n275 vdd.t102 4.06363
R5607 vdd.n273 vdd.t116 4.06363
R5608 vdd.n273 vdd.t198 4.06363
R5609 vdd.n271 vdd.t259 4.06363
R5610 vdd.n271 vdd.t214 4.06363
R5611 vdd.n269 vdd.t182 4.06363
R5612 vdd.n269 vdd.t120 4.06363
R5613 vdd.n267 vdd.t202 4.06363
R5614 vdd.n267 vdd.t184 4.06363
R5615 vdd.n265 vdd.t209 4.06363
R5616 vdd.n265 vdd.t253 4.06363
R5617 vdd.n179 vdd.t20 4.06363
R5618 vdd.n179 vdd.t207 4.06363
R5619 vdd.n177 vdd.t206 4.06363
R5620 vdd.n177 vdd.t212 4.06363
R5621 vdd.n175 vdd.t9 4.06363
R5622 vdd.n175 vdd.t16 4.06363
R5623 vdd.n173 vdd.t244 4.06363
R5624 vdd.n173 vdd.t247 4.06363
R5625 vdd.n171 vdd.t194 4.06363
R5626 vdd.n171 vdd.t257 4.06363
R5627 vdd.n169 vdd.t256 4.06363
R5628 vdd.n169 vdd.t195 4.06363
R5629 vdd.n167 vdd.t264 4.06363
R5630 vdd.n167 vdd.t224 4.06363
R5631 vdd.n82 vdd.t222 4.06363
R5632 vdd.n82 vdd.t112 4.06363
R5633 vdd.n80 vdd.t127 4.06363
R5634 vdd.n80 vdd.t263 4.06363
R5635 vdd.n78 vdd.t255 4.06363
R5636 vdd.n78 vdd.t126 4.06363
R5637 vdd.n76 vdd.t110 4.06363
R5638 vdd.n76 vdd.t251 4.06363
R5639 vdd.n74 vdd.t269 4.06363
R5640 vdd.n74 vdd.t248 4.06363
R5641 vdd.n72 vdd.t108 4.06363
R5642 vdd.n72 vdd.t218 4.06363
R5643 vdd.n70 vdd.t122 4.06363
R5644 vdd.n70 vdd.t226 4.06363
R5645 vdd.n1769 vdd.t217 4.06363
R5646 vdd.n1769 vdd.t254 4.06363
R5647 vdd.n1771 vdd.t261 4.06363
R5648 vdd.n1771 vdd.t243 4.06363
R5649 vdd.n1773 vdd.t266 4.06363
R5650 vdd.n1773 vdd.t1 4.06363
R5651 vdd.n1775 vdd.t187 4.06363
R5652 vdd.n1775 vdd.t245 4.06363
R5653 vdd.n1777 vdd.t208 4.06363
R5654 vdd.n1777 vdd.t3 4.06363
R5655 vdd.n1779 vdd.t18 4.06363
R5656 vdd.n1779 vdd.t115 4.06363
R5657 vdd.n1781 vdd.t11 4.06363
R5658 vdd.n1781 vdd.t197 4.06363
R5659 vdd.n1671 vdd.t265 4.06363
R5660 vdd.n1671 vdd.t241 4.06363
R5661 vdd.n1673 vdd.t5 4.06363
R5662 vdd.n1673 vdd.t238 4.06363
R5663 vdd.n1675 vdd.t221 4.06363
R5664 vdd.n1675 vdd.t240 4.06363
R5665 vdd.n1677 vdd.t7 4.06363
R5666 vdd.n1677 vdd.t262 4.06363
R5667 vdd.n1679 vdd.t242 4.06363
R5668 vdd.n1679 vdd.t14 4.06363
R5669 vdd.n1681 vdd.t128 4.06363
R5670 vdd.n1681 vdd.t188 4.06363
R5671 vdd.n1683 vdd.t189 4.06363
R5672 vdd.n1683 vdd.t237 4.06363
R5673 vdd.n1574 vdd.t186 4.06363
R5674 vdd.n1574 vdd.t104 4.06363
R5675 vdd.n1576 vdd.t219 4.06363
R5676 vdd.n1576 vdd.t106 4.06363
R5677 vdd.n1578 vdd.t258 4.06363
R5678 vdd.n1578 vdd.t236 4.06363
R5679 vdd.n1580 vdd.t252 4.06363
R5680 vdd.n1580 vdd.t205 4.06363
R5681 vdd.n1582 vdd.t200 4.06363
R5682 vdd.n1582 vdd.t123 4.06363
R5683 vdd.n1584 vdd.t250 4.06363
R5684 vdd.n1584 vdd.t260 4.06363
R5685 vdd.n1586 vdd.t113 4.06363
R5686 vdd.n1586 vdd.t13 4.06363
R5687 vdd.n26 vdd.t193 3.9605
R5688 vdd.n26 vdd.t190 3.9605
R5689 vdd.n23 vdd.t228 3.9605
R5690 vdd.n23 vdd.t233 3.9605
R5691 vdd.n21 vdd.t231 3.9605
R5692 vdd.n21 vdd.t270 3.9605
R5693 vdd.n20 vdd.t118 3.9605
R5694 vdd.n20 vdd.t23 3.9605
R5695 vdd.n15 vdd.t271 3.9605
R5696 vdd.n15 vdd.t24 3.9605
R5697 vdd.n16 vdd.t117 3.9605
R5698 vdd.n16 vdd.t191 3.9605
R5699 vdd.n18 vdd.t232 3.9605
R5700 vdd.n18 vdd.t229 3.9605
R5701 vdd.n25 vdd.t192 3.9605
R5702 vdd.n25 vdd.t230 3.9605
R5703 vdd.n2997 vdd.n2996 3.74684
R5704 vdd.n2437 vdd.n2436 3.74684
R5705 vdd.n7 vdd.t180 3.61217
R5706 vdd.n7 vdd.t146 3.61217
R5707 vdd.n8 vdd.t154 3.61217
R5708 vdd.n8 vdd.t172 3.61217
R5709 vdd.n10 vdd.t162 3.61217
R5710 vdd.n10 vdd.t135 3.61217
R5711 vdd.n12 vdd.t143 3.61217
R5712 vdd.n12 vdd.t160 3.61217
R5713 vdd.n5 vdd.t176 3.61217
R5714 vdd.n5 vdd.t156 3.61217
R5715 vdd.n3 vdd.t148 3.61217
R5716 vdd.n3 vdd.t174 3.61217
R5717 vdd.n1 vdd.t132 3.61217
R5718 vdd.n1 vdd.t165 3.61217
R5719 vdd.n0 vdd.t170 3.61217
R5720 vdd.n0 vdd.t151 3.61217
R5721 vdd.n1462 vdd.t56 3.51482
R5722 vdd.n2414 vdd.t140 3.51482
R5723 vdd.n2469 vdd.t152 3.51482
R5724 vdd.n2964 vdd.t168 3.51482
R5725 vdd.n3019 vdd.t163 3.51482
R5726 vdd.n3437 vdd.t38 3.51482
R5727 vdd.n304 vdd.n303 3.49141
R5728 vdd.n249 vdd.n248 3.49141
R5729 vdd.n206 vdd.n205 3.49141
R5730 vdd.n151 vdd.n150 3.49141
R5731 vdd.n109 vdd.n108 3.49141
R5732 vdd.n54 vdd.n53 3.49141
R5733 vdd.n1753 vdd.n1752 3.49141
R5734 vdd.n1808 vdd.n1807 3.49141
R5735 vdd.n1655 vdd.n1654 3.49141
R5736 vdd.n1710 vdd.n1709 3.49141
R5737 vdd.n1558 vdd.n1557 3.49141
R5738 vdd.n1613 vdd.n1612 3.49141
R5739 vdd.n2489 vdd.t147 3.40145
R5740 vdd.n2643 vdd.t175 3.40145
R5741 vdd.n2927 vdd.t159 3.40145
R5742 vdd.n2946 vdd.t134 3.40145
R5743 vdd.n1865 vdd.t185 3.06136
R5744 vdd.n3359 vdd.t223 3.06136
R5745 vdd.t164 vdd.n986 2.94799
R5746 vdd.n901 vdd.t153 2.94799
R5747 vdd.t0 vdd.n1161 2.83463
R5748 vdd.n2390 vdd.t34 2.83463
R5749 vdd.n2496 vdd.t72 2.83463
R5750 vdd.n2940 vdd.t76 2.83463
R5751 vdd.n3088 vdd.t30 2.83463
R5752 vdd.n624 vdd.t181 2.83463
R5753 vdd.n307 vdd.n286 2.71565
R5754 vdd.n252 vdd.n231 2.71565
R5755 vdd.n209 vdd.n188 2.71565
R5756 vdd.n154 vdd.n133 2.71565
R5757 vdd.n112 vdd.n91 2.71565
R5758 vdd.n57 vdd.n36 2.71565
R5759 vdd.n1756 vdd.n1735 2.71565
R5760 vdd.n1811 vdd.n1790 2.71565
R5761 vdd.n1658 vdd.n1637 2.71565
R5762 vdd.n1713 vdd.n1692 2.71565
R5763 vdd.n1561 vdd.n1540 2.71565
R5764 vdd.n1616 vdd.n1595 2.71565
R5765 vdd.n1529 vdd.t6 2.6079
R5766 vdd.n1041 vdd.t158 2.6079
R5767 vdd.n2275 vdd.t177 2.6079
R5768 vdd.n2894 vdd.t167 2.6079
R5769 vdd.t136 vdd.n845 2.6079
R5770 vdd.n3469 vdd.t213 2.6079
R5771 vdd.n294 vdd.n293 2.4129
R5772 vdd.n239 vdd.n238 2.4129
R5773 vdd.n196 vdd.n195 2.4129
R5774 vdd.n141 vdd.n140 2.4129
R5775 vdd.n99 vdd.n98 2.4129
R5776 vdd.n44 vdd.n43 2.4129
R5777 vdd.n1743 vdd.n1742 2.4129
R5778 vdd.n1798 vdd.n1797 2.4129
R5779 vdd.n1645 vdd.n1644 2.4129
R5780 vdd.n1700 vdd.n1699 2.4129
R5781 vdd.n1548 vdd.n1547 2.4129
R5782 vdd.n1603 vdd.n1602 2.4129
R5783 vdd.t114 vdd.n1190 2.38117
R5784 vdd.n3460 vdd.t124 2.38117
R5785 vdd.n2099 vdd.n1901 2.27742
R5786 vdd.n2100 vdd.n2099 2.27742
R5787 vdd.n3124 vdd.n665 2.27742
R5788 vdd.n3124 vdd.n664 2.27742
R5789 vdd.n3192 vdd.n751 2.27742
R5790 vdd.n3192 vdd.n749 2.27742
R5791 vdd.n2122 vdd.n1116 2.27742
R5792 vdd.n2122 vdd.n1117 2.27742
R5793 vdd.n2275 vdd.t169 2.2678
R5794 vdd.n2894 vdd.t145 2.2678
R5795 vdd.n1487 vdd.t10 2.15444
R5796 vdd.n3451 vdd.t111 2.15444
R5797 vdd.n2463 vdd.t150 2.04107
R5798 vdd.n2970 vdd.t179 2.04107
R5799 vdd.n308 vdd.n284 1.93989
R5800 vdd.n253 vdd.n229 1.93989
R5801 vdd.n210 vdd.n186 1.93989
R5802 vdd.n155 vdd.n131 1.93989
R5803 vdd.n113 vdd.n89 1.93989
R5804 vdd.n58 vdd.n34 1.93989
R5805 vdd.n1757 vdd.n1733 1.93989
R5806 vdd.n1812 vdd.n1788 1.93989
R5807 vdd.n1659 vdd.n1635 1.93989
R5808 vdd.n1714 vdd.n1690 1.93989
R5809 vdd.n1562 vdd.n1538 1.93989
R5810 vdd.n1617 vdd.n1593 1.93989
R5811 vdd.n1479 vdd.t21 1.70098
R5812 vdd.n2439 vdd.t137 1.70098
R5813 vdd.n2445 vdd.t144 1.70098
R5814 vdd.n2988 vdd.t149 1.70098
R5815 vdd.n2994 vdd.t138 1.70098
R5816 vdd.n3445 vdd.t210 1.70098
R5817 vdd.n1495 vdd.t17 1.47425
R5818 vdd.n349 vdd.t101 1.47425
R5819 vdd.n2469 vdd.t131 1.36088
R5820 vdd.n2964 vdd.t171 1.36088
R5821 vdd.n1520 vdd.t2 1.24752
R5822 vdd.t52 vdd.n1124 1.24752
R5823 vdd.n659 vdd.t26 1.24752
R5824 vdd.t8 vdd.n3467 1.24752
R5825 vdd.n319 vdd.n279 1.16414
R5826 vdd.n312 vdd.n311 1.16414
R5827 vdd.n264 vdd.n224 1.16414
R5828 vdd.n257 vdd.n256 1.16414
R5829 vdd.n221 vdd.n181 1.16414
R5830 vdd.n214 vdd.n213 1.16414
R5831 vdd.n166 vdd.n126 1.16414
R5832 vdd.n159 vdd.n158 1.16414
R5833 vdd.n124 vdd.n84 1.16414
R5834 vdd.n117 vdd.n116 1.16414
R5835 vdd.n69 vdd.n29 1.16414
R5836 vdd.n62 vdd.n61 1.16414
R5837 vdd.n1768 vdd.n1728 1.16414
R5838 vdd.n1761 vdd.n1760 1.16414
R5839 vdd.n1823 vdd.n1783 1.16414
R5840 vdd.n1816 vdd.n1815 1.16414
R5841 vdd.n1670 vdd.n1630 1.16414
R5842 vdd.n1663 vdd.n1662 1.16414
R5843 vdd.n1725 vdd.n1685 1.16414
R5844 vdd.n1718 vdd.n1717 1.16414
R5845 vdd.n1573 vdd.n1533 1.16414
R5846 vdd.n1566 vdd.n1565 1.16414
R5847 vdd.n1628 vdd.n1588 1.16414
R5848 vdd.n1621 vdd.n1620 1.16414
R5849 vdd.n1826 vdd.n28 1.06035
R5850 vdd vdd.n3474 1.05252
R5851 vdd.n1172 vdd.t220 1.02079
R5852 vdd.t86 vdd.t137 1.02079
R5853 vdd.t138 vdd.t45 1.02079
R5854 vdd.t119 vdd.n613 1.02079
R5855 vdd.n1351 vdd.n1230 0.970197
R5856 vdd.n2120 vdd.n2119 0.970197
R5857 vdd.n599 vdd.n407 0.970197
R5858 vdd.n3199 vdd.n3197 0.970197
R5859 vdd.t173 vdd.n963 0.907421
R5860 vdd.n917 vdd.t161 0.907421
R5861 vdd.n1857 vdd.t105 0.794056
R5862 vdd.t141 vdd.n1038 0.794056
R5863 vdd.n1010 vdd.t139 0.794056
R5864 vdd.t129 vdd.n876 0.794056
R5865 vdd.n848 vdd.t166 0.794056
R5866 vdd.n3368 vdd.t107 0.794056
R5867 vdd.n1873 vdd.t234 0.567326
R5868 vdd.t215 vdd.n642 0.567326
R5869 vdd.n2110 vdd.n2109 0.482207
R5870 vdd.n3324 vdd.n3323 0.482207
R5871 vdd.n444 vdd.n443 0.482207
R5872 vdd.n3431 vdd.n3430 0.482207
R5873 vdd.n3330 vdd.n656 0.482207
R5874 vdd.n1887 vdd.n1118 0.482207
R5875 vdd.n1458 vdd.n1457 0.482207
R5876 vdd.n1264 vdd.n1221 0.482207
R5877 vdd.n4 vdd.n2 0.459552
R5878 vdd.n11 vdd.n9 0.459552
R5879 vdd.n317 vdd.n316 0.388379
R5880 vdd.n283 vdd.n281 0.388379
R5881 vdd.n262 vdd.n261 0.388379
R5882 vdd.n228 vdd.n226 0.388379
R5883 vdd.n219 vdd.n218 0.388379
R5884 vdd.n185 vdd.n183 0.388379
R5885 vdd.n164 vdd.n163 0.388379
R5886 vdd.n130 vdd.n128 0.388379
R5887 vdd.n122 vdd.n121 0.388379
R5888 vdd.n88 vdd.n86 0.388379
R5889 vdd.n67 vdd.n66 0.388379
R5890 vdd.n33 vdd.n31 0.388379
R5891 vdd.n1766 vdd.n1765 0.388379
R5892 vdd.n1732 vdd.n1730 0.388379
R5893 vdd.n1821 vdd.n1820 0.388379
R5894 vdd.n1787 vdd.n1785 0.388379
R5895 vdd.n1668 vdd.n1667 0.388379
R5896 vdd.n1634 vdd.n1632 0.388379
R5897 vdd.n1723 vdd.n1722 0.388379
R5898 vdd.n1689 vdd.n1687 0.388379
R5899 vdd.n1571 vdd.n1570 0.388379
R5900 vdd.n1537 vdd.n1535 0.388379
R5901 vdd.n1626 vdd.n1625 0.388379
R5902 vdd.n1592 vdd.n1590 0.388379
R5903 vdd.n19 vdd.n17 0.387128
R5904 vdd.n24 vdd.n22 0.387128
R5905 vdd.n6 vdd.n4 0.358259
R5906 vdd.n13 vdd.n11 0.358259
R5907 vdd.n268 vdd.n266 0.358259
R5908 vdd.n270 vdd.n268 0.358259
R5909 vdd.n272 vdd.n270 0.358259
R5910 vdd.n274 vdd.n272 0.358259
R5911 vdd.n276 vdd.n274 0.358259
R5912 vdd.n278 vdd.n276 0.358259
R5913 vdd.n320 vdd.n278 0.358259
R5914 vdd.n170 vdd.n168 0.358259
R5915 vdd.n172 vdd.n170 0.358259
R5916 vdd.n174 vdd.n172 0.358259
R5917 vdd.n176 vdd.n174 0.358259
R5918 vdd.n178 vdd.n176 0.358259
R5919 vdd.n180 vdd.n178 0.358259
R5920 vdd.n222 vdd.n180 0.358259
R5921 vdd.n73 vdd.n71 0.358259
R5922 vdd.n75 vdd.n73 0.358259
R5923 vdd.n77 vdd.n75 0.358259
R5924 vdd.n79 vdd.n77 0.358259
R5925 vdd.n81 vdd.n79 0.358259
R5926 vdd.n83 vdd.n81 0.358259
R5927 vdd.n125 vdd.n83 0.358259
R5928 vdd.n1824 vdd.n1782 0.358259
R5929 vdd.n1782 vdd.n1780 0.358259
R5930 vdd.n1780 vdd.n1778 0.358259
R5931 vdd.n1778 vdd.n1776 0.358259
R5932 vdd.n1776 vdd.n1774 0.358259
R5933 vdd.n1774 vdd.n1772 0.358259
R5934 vdd.n1772 vdd.n1770 0.358259
R5935 vdd.n1726 vdd.n1684 0.358259
R5936 vdd.n1684 vdd.n1682 0.358259
R5937 vdd.n1682 vdd.n1680 0.358259
R5938 vdd.n1680 vdd.n1678 0.358259
R5939 vdd.n1678 vdd.n1676 0.358259
R5940 vdd.n1676 vdd.n1674 0.358259
R5941 vdd.n1674 vdd.n1672 0.358259
R5942 vdd.n1629 vdd.n1587 0.358259
R5943 vdd.n1587 vdd.n1585 0.358259
R5944 vdd.n1585 vdd.n1583 0.358259
R5945 vdd.n1583 vdd.n1581 0.358259
R5946 vdd.n1581 vdd.n1579 0.358259
R5947 vdd.n1579 vdd.n1577 0.358259
R5948 vdd.n1577 vdd.n1575 0.358259
R5949 vdd.n14 vdd.n6 0.334552
R5950 vdd.n14 vdd.n13 0.334552
R5951 vdd.n27 vdd.n19 0.21707
R5952 vdd.n27 vdd.n24 0.21707
R5953 vdd.n318 vdd.n280 0.155672
R5954 vdd.n310 vdd.n280 0.155672
R5955 vdd.n310 vdd.n309 0.155672
R5956 vdd.n309 vdd.n285 0.155672
R5957 vdd.n302 vdd.n285 0.155672
R5958 vdd.n302 vdd.n301 0.155672
R5959 vdd.n301 vdd.n289 0.155672
R5960 vdd.n294 vdd.n289 0.155672
R5961 vdd.n263 vdd.n225 0.155672
R5962 vdd.n255 vdd.n225 0.155672
R5963 vdd.n255 vdd.n254 0.155672
R5964 vdd.n254 vdd.n230 0.155672
R5965 vdd.n247 vdd.n230 0.155672
R5966 vdd.n247 vdd.n246 0.155672
R5967 vdd.n246 vdd.n234 0.155672
R5968 vdd.n239 vdd.n234 0.155672
R5969 vdd.n220 vdd.n182 0.155672
R5970 vdd.n212 vdd.n182 0.155672
R5971 vdd.n212 vdd.n211 0.155672
R5972 vdd.n211 vdd.n187 0.155672
R5973 vdd.n204 vdd.n187 0.155672
R5974 vdd.n204 vdd.n203 0.155672
R5975 vdd.n203 vdd.n191 0.155672
R5976 vdd.n196 vdd.n191 0.155672
R5977 vdd.n165 vdd.n127 0.155672
R5978 vdd.n157 vdd.n127 0.155672
R5979 vdd.n157 vdd.n156 0.155672
R5980 vdd.n156 vdd.n132 0.155672
R5981 vdd.n149 vdd.n132 0.155672
R5982 vdd.n149 vdd.n148 0.155672
R5983 vdd.n148 vdd.n136 0.155672
R5984 vdd.n141 vdd.n136 0.155672
R5985 vdd.n123 vdd.n85 0.155672
R5986 vdd.n115 vdd.n85 0.155672
R5987 vdd.n115 vdd.n114 0.155672
R5988 vdd.n114 vdd.n90 0.155672
R5989 vdd.n107 vdd.n90 0.155672
R5990 vdd.n107 vdd.n106 0.155672
R5991 vdd.n106 vdd.n94 0.155672
R5992 vdd.n99 vdd.n94 0.155672
R5993 vdd.n68 vdd.n30 0.155672
R5994 vdd.n60 vdd.n30 0.155672
R5995 vdd.n60 vdd.n59 0.155672
R5996 vdd.n59 vdd.n35 0.155672
R5997 vdd.n52 vdd.n35 0.155672
R5998 vdd.n52 vdd.n51 0.155672
R5999 vdd.n51 vdd.n39 0.155672
R6000 vdd.n44 vdd.n39 0.155672
R6001 vdd.n1767 vdd.n1729 0.155672
R6002 vdd.n1759 vdd.n1729 0.155672
R6003 vdd.n1759 vdd.n1758 0.155672
R6004 vdd.n1758 vdd.n1734 0.155672
R6005 vdd.n1751 vdd.n1734 0.155672
R6006 vdd.n1751 vdd.n1750 0.155672
R6007 vdd.n1750 vdd.n1738 0.155672
R6008 vdd.n1743 vdd.n1738 0.155672
R6009 vdd.n1822 vdd.n1784 0.155672
R6010 vdd.n1814 vdd.n1784 0.155672
R6011 vdd.n1814 vdd.n1813 0.155672
R6012 vdd.n1813 vdd.n1789 0.155672
R6013 vdd.n1806 vdd.n1789 0.155672
R6014 vdd.n1806 vdd.n1805 0.155672
R6015 vdd.n1805 vdd.n1793 0.155672
R6016 vdd.n1798 vdd.n1793 0.155672
R6017 vdd.n1669 vdd.n1631 0.155672
R6018 vdd.n1661 vdd.n1631 0.155672
R6019 vdd.n1661 vdd.n1660 0.155672
R6020 vdd.n1660 vdd.n1636 0.155672
R6021 vdd.n1653 vdd.n1636 0.155672
R6022 vdd.n1653 vdd.n1652 0.155672
R6023 vdd.n1652 vdd.n1640 0.155672
R6024 vdd.n1645 vdd.n1640 0.155672
R6025 vdd.n1724 vdd.n1686 0.155672
R6026 vdd.n1716 vdd.n1686 0.155672
R6027 vdd.n1716 vdd.n1715 0.155672
R6028 vdd.n1715 vdd.n1691 0.155672
R6029 vdd.n1708 vdd.n1691 0.155672
R6030 vdd.n1708 vdd.n1707 0.155672
R6031 vdd.n1707 vdd.n1695 0.155672
R6032 vdd.n1700 vdd.n1695 0.155672
R6033 vdd.n1572 vdd.n1534 0.155672
R6034 vdd.n1564 vdd.n1534 0.155672
R6035 vdd.n1564 vdd.n1563 0.155672
R6036 vdd.n1563 vdd.n1539 0.155672
R6037 vdd.n1556 vdd.n1539 0.155672
R6038 vdd.n1556 vdd.n1555 0.155672
R6039 vdd.n1555 vdd.n1543 0.155672
R6040 vdd.n1548 vdd.n1543 0.155672
R6041 vdd.n1627 vdd.n1589 0.155672
R6042 vdd.n1619 vdd.n1589 0.155672
R6043 vdd.n1619 vdd.n1618 0.155672
R6044 vdd.n1618 vdd.n1594 0.155672
R6045 vdd.n1611 vdd.n1594 0.155672
R6046 vdd.n1611 vdd.n1610 0.155672
R6047 vdd.n1610 vdd.n1598 0.155672
R6048 vdd.n1603 vdd.n1598 0.155672
R6049 vdd.n2098 vdd.n1903 0.152939
R6050 vdd.n1909 vdd.n1903 0.152939
R6051 vdd.n1910 vdd.n1909 0.152939
R6052 vdd.n1911 vdd.n1910 0.152939
R6053 vdd.n1912 vdd.n1911 0.152939
R6054 vdd.n1916 vdd.n1912 0.152939
R6055 vdd.n1917 vdd.n1916 0.152939
R6056 vdd.n1918 vdd.n1917 0.152939
R6057 vdd.n1919 vdd.n1918 0.152939
R6058 vdd.n1923 vdd.n1919 0.152939
R6059 vdd.n1924 vdd.n1923 0.152939
R6060 vdd.n1925 vdd.n1924 0.152939
R6061 vdd.n2073 vdd.n1925 0.152939
R6062 vdd.n2073 vdd.n2072 0.152939
R6063 vdd.n2072 vdd.n2071 0.152939
R6064 vdd.n2071 vdd.n1931 0.152939
R6065 vdd.n1936 vdd.n1931 0.152939
R6066 vdd.n1937 vdd.n1936 0.152939
R6067 vdd.n1938 vdd.n1937 0.152939
R6068 vdd.n1942 vdd.n1938 0.152939
R6069 vdd.n1943 vdd.n1942 0.152939
R6070 vdd.n1944 vdd.n1943 0.152939
R6071 vdd.n1945 vdd.n1944 0.152939
R6072 vdd.n1949 vdd.n1945 0.152939
R6073 vdd.n1950 vdd.n1949 0.152939
R6074 vdd.n1951 vdd.n1950 0.152939
R6075 vdd.n1952 vdd.n1951 0.152939
R6076 vdd.n1956 vdd.n1952 0.152939
R6077 vdd.n1957 vdd.n1956 0.152939
R6078 vdd.n1958 vdd.n1957 0.152939
R6079 vdd.n1959 vdd.n1958 0.152939
R6080 vdd.n1963 vdd.n1959 0.152939
R6081 vdd.n1964 vdd.n1963 0.152939
R6082 vdd.n1965 vdd.n1964 0.152939
R6083 vdd.n2034 vdd.n1965 0.152939
R6084 vdd.n2034 vdd.n2033 0.152939
R6085 vdd.n2033 vdd.n2032 0.152939
R6086 vdd.n2032 vdd.n1971 0.152939
R6087 vdd.n1976 vdd.n1971 0.152939
R6088 vdd.n1977 vdd.n1976 0.152939
R6089 vdd.n1978 vdd.n1977 0.152939
R6090 vdd.n1982 vdd.n1978 0.152939
R6091 vdd.n1983 vdd.n1982 0.152939
R6092 vdd.n1984 vdd.n1983 0.152939
R6093 vdd.n1985 vdd.n1984 0.152939
R6094 vdd.n1989 vdd.n1985 0.152939
R6095 vdd.n1990 vdd.n1989 0.152939
R6096 vdd.n1991 vdd.n1990 0.152939
R6097 vdd.n1992 vdd.n1991 0.152939
R6098 vdd.n1993 vdd.n1992 0.152939
R6099 vdd.n1993 vdd.n1115 0.152939
R6100 vdd.n2109 vdd.n1897 0.152939
R6101 vdd.n1829 vdd.n1828 0.152939
R6102 vdd.n1829 vdd.n1164 0.152939
R6103 vdd.n1843 vdd.n1164 0.152939
R6104 vdd.n1844 vdd.n1843 0.152939
R6105 vdd.n1845 vdd.n1844 0.152939
R6106 vdd.n1845 vdd.n1152 0.152939
R6107 vdd.n1860 vdd.n1152 0.152939
R6108 vdd.n1861 vdd.n1860 0.152939
R6109 vdd.n1862 vdd.n1861 0.152939
R6110 vdd.n1862 vdd.n1141 0.152939
R6111 vdd.n1877 vdd.n1141 0.152939
R6112 vdd.n1878 vdd.n1877 0.152939
R6113 vdd.n1879 vdd.n1878 0.152939
R6114 vdd.n1879 vdd.n1129 0.152939
R6115 vdd.n1895 vdd.n1129 0.152939
R6116 vdd.n1896 vdd.n1895 0.152939
R6117 vdd.n2110 vdd.n1896 0.152939
R6118 vdd.n670 vdd.n667 0.152939
R6119 vdd.n671 vdd.n670 0.152939
R6120 vdd.n672 vdd.n671 0.152939
R6121 vdd.n673 vdd.n672 0.152939
R6122 vdd.n676 vdd.n673 0.152939
R6123 vdd.n677 vdd.n676 0.152939
R6124 vdd.n678 vdd.n677 0.152939
R6125 vdd.n679 vdd.n678 0.152939
R6126 vdd.n682 vdd.n679 0.152939
R6127 vdd.n683 vdd.n682 0.152939
R6128 vdd.n684 vdd.n683 0.152939
R6129 vdd.n685 vdd.n684 0.152939
R6130 vdd.n690 vdd.n685 0.152939
R6131 vdd.n691 vdd.n690 0.152939
R6132 vdd.n692 vdd.n691 0.152939
R6133 vdd.n693 vdd.n692 0.152939
R6134 vdd.n696 vdd.n693 0.152939
R6135 vdd.n697 vdd.n696 0.152939
R6136 vdd.n698 vdd.n697 0.152939
R6137 vdd.n699 vdd.n698 0.152939
R6138 vdd.n702 vdd.n699 0.152939
R6139 vdd.n703 vdd.n702 0.152939
R6140 vdd.n704 vdd.n703 0.152939
R6141 vdd.n705 vdd.n704 0.152939
R6142 vdd.n708 vdd.n705 0.152939
R6143 vdd.n709 vdd.n708 0.152939
R6144 vdd.n710 vdd.n709 0.152939
R6145 vdd.n711 vdd.n710 0.152939
R6146 vdd.n714 vdd.n711 0.152939
R6147 vdd.n715 vdd.n714 0.152939
R6148 vdd.n716 vdd.n715 0.152939
R6149 vdd.n717 vdd.n716 0.152939
R6150 vdd.n720 vdd.n717 0.152939
R6151 vdd.n721 vdd.n720 0.152939
R6152 vdd.n3240 vdd.n721 0.152939
R6153 vdd.n3240 vdd.n3239 0.152939
R6154 vdd.n3239 vdd.n3238 0.152939
R6155 vdd.n3238 vdd.n725 0.152939
R6156 vdd.n730 vdd.n725 0.152939
R6157 vdd.n731 vdd.n730 0.152939
R6158 vdd.n734 vdd.n731 0.152939
R6159 vdd.n735 vdd.n734 0.152939
R6160 vdd.n736 vdd.n735 0.152939
R6161 vdd.n737 vdd.n736 0.152939
R6162 vdd.n740 vdd.n737 0.152939
R6163 vdd.n741 vdd.n740 0.152939
R6164 vdd.n742 vdd.n741 0.152939
R6165 vdd.n743 vdd.n742 0.152939
R6166 vdd.n746 vdd.n743 0.152939
R6167 vdd.n747 vdd.n746 0.152939
R6168 vdd.n748 vdd.n747 0.152939
R6169 vdd.n3323 vdd.n661 0.152939
R6170 vdd.n3324 vdd.n651 0.152939
R6171 vdd.n3338 vdd.n651 0.152939
R6172 vdd.n3339 vdd.n3338 0.152939
R6173 vdd.n3340 vdd.n3339 0.152939
R6174 vdd.n3340 vdd.n639 0.152939
R6175 vdd.n3354 vdd.n639 0.152939
R6176 vdd.n3355 vdd.n3354 0.152939
R6177 vdd.n3356 vdd.n3355 0.152939
R6178 vdd.n3356 vdd.n627 0.152939
R6179 vdd.n3371 vdd.n627 0.152939
R6180 vdd.n3372 vdd.n3371 0.152939
R6181 vdd.n3373 vdd.n3372 0.152939
R6182 vdd.n3373 vdd.n616 0.152939
R6183 vdd.n3390 vdd.n616 0.152939
R6184 vdd.n3391 vdd.n3390 0.152939
R6185 vdd.n3392 vdd.n3391 0.152939
R6186 vdd.n3392 vdd.n322 0.152939
R6187 vdd.n3472 vdd.n323 0.152939
R6188 vdd.n334 vdd.n323 0.152939
R6189 vdd.n335 vdd.n334 0.152939
R6190 vdd.n336 vdd.n335 0.152939
R6191 vdd.n343 vdd.n336 0.152939
R6192 vdd.n344 vdd.n343 0.152939
R6193 vdd.n345 vdd.n344 0.152939
R6194 vdd.n346 vdd.n345 0.152939
R6195 vdd.n354 vdd.n346 0.152939
R6196 vdd.n355 vdd.n354 0.152939
R6197 vdd.n356 vdd.n355 0.152939
R6198 vdd.n357 vdd.n356 0.152939
R6199 vdd.n365 vdd.n357 0.152939
R6200 vdd.n366 vdd.n365 0.152939
R6201 vdd.n367 vdd.n366 0.152939
R6202 vdd.n368 vdd.n367 0.152939
R6203 vdd.n443 vdd.n368 0.152939
R6204 vdd.n444 vdd.n442 0.152939
R6205 vdd.n451 vdd.n442 0.152939
R6206 vdd.n452 vdd.n451 0.152939
R6207 vdd.n453 vdd.n452 0.152939
R6208 vdd.n453 vdd.n440 0.152939
R6209 vdd.n461 vdd.n440 0.152939
R6210 vdd.n462 vdd.n461 0.152939
R6211 vdd.n463 vdd.n462 0.152939
R6212 vdd.n463 vdd.n438 0.152939
R6213 vdd.n471 vdd.n438 0.152939
R6214 vdd.n472 vdd.n471 0.152939
R6215 vdd.n473 vdd.n472 0.152939
R6216 vdd.n473 vdd.n436 0.152939
R6217 vdd.n481 vdd.n436 0.152939
R6218 vdd.n482 vdd.n481 0.152939
R6219 vdd.n483 vdd.n482 0.152939
R6220 vdd.n483 vdd.n434 0.152939
R6221 vdd.n491 vdd.n434 0.152939
R6222 vdd.n492 vdd.n491 0.152939
R6223 vdd.n493 vdd.n492 0.152939
R6224 vdd.n493 vdd.n430 0.152939
R6225 vdd.n501 vdd.n430 0.152939
R6226 vdd.n502 vdd.n501 0.152939
R6227 vdd.n503 vdd.n502 0.152939
R6228 vdd.n503 vdd.n428 0.152939
R6229 vdd.n511 vdd.n428 0.152939
R6230 vdd.n512 vdd.n511 0.152939
R6231 vdd.n513 vdd.n512 0.152939
R6232 vdd.n513 vdd.n426 0.152939
R6233 vdd.n521 vdd.n426 0.152939
R6234 vdd.n522 vdd.n521 0.152939
R6235 vdd.n523 vdd.n522 0.152939
R6236 vdd.n523 vdd.n424 0.152939
R6237 vdd.n531 vdd.n424 0.152939
R6238 vdd.n532 vdd.n531 0.152939
R6239 vdd.n533 vdd.n532 0.152939
R6240 vdd.n533 vdd.n422 0.152939
R6241 vdd.n541 vdd.n422 0.152939
R6242 vdd.n542 vdd.n541 0.152939
R6243 vdd.n543 vdd.n542 0.152939
R6244 vdd.n543 vdd.n418 0.152939
R6245 vdd.n551 vdd.n418 0.152939
R6246 vdd.n552 vdd.n551 0.152939
R6247 vdd.n553 vdd.n552 0.152939
R6248 vdd.n553 vdd.n416 0.152939
R6249 vdd.n561 vdd.n416 0.152939
R6250 vdd.n562 vdd.n561 0.152939
R6251 vdd.n563 vdd.n562 0.152939
R6252 vdd.n563 vdd.n414 0.152939
R6253 vdd.n571 vdd.n414 0.152939
R6254 vdd.n572 vdd.n571 0.152939
R6255 vdd.n573 vdd.n572 0.152939
R6256 vdd.n573 vdd.n412 0.152939
R6257 vdd.n581 vdd.n412 0.152939
R6258 vdd.n582 vdd.n581 0.152939
R6259 vdd.n583 vdd.n582 0.152939
R6260 vdd.n583 vdd.n410 0.152939
R6261 vdd.n591 vdd.n410 0.152939
R6262 vdd.n592 vdd.n591 0.152939
R6263 vdd.n593 vdd.n592 0.152939
R6264 vdd.n593 vdd.n408 0.152939
R6265 vdd.n600 vdd.n408 0.152939
R6266 vdd.n3431 vdd.n600 0.152939
R6267 vdd.n3331 vdd.n3330 0.152939
R6268 vdd.n3332 vdd.n3331 0.152939
R6269 vdd.n3332 vdd.n645 0.152939
R6270 vdd.n3346 vdd.n645 0.152939
R6271 vdd.n3347 vdd.n3346 0.152939
R6272 vdd.n3348 vdd.n3347 0.152939
R6273 vdd.n3348 vdd.n632 0.152939
R6274 vdd.n3362 vdd.n632 0.152939
R6275 vdd.n3363 vdd.n3362 0.152939
R6276 vdd.n3364 vdd.n3363 0.152939
R6277 vdd.n3364 vdd.n621 0.152939
R6278 vdd.n3379 vdd.n621 0.152939
R6279 vdd.n3380 vdd.n3379 0.152939
R6280 vdd.n3381 vdd.n3380 0.152939
R6281 vdd.n3383 vdd.n3381 0.152939
R6282 vdd.n3383 vdd.n3382 0.152939
R6283 vdd.n3382 vdd.n611 0.152939
R6284 vdd.n611 vdd.n609 0.152939
R6285 vdd.n3401 vdd.n609 0.152939
R6286 vdd.n3402 vdd.n3401 0.152939
R6287 vdd.n3403 vdd.n3402 0.152939
R6288 vdd.n3403 vdd.n607 0.152939
R6289 vdd.n3408 vdd.n607 0.152939
R6290 vdd.n3409 vdd.n3408 0.152939
R6291 vdd.n3410 vdd.n3409 0.152939
R6292 vdd.n3410 vdd.n605 0.152939
R6293 vdd.n3415 vdd.n605 0.152939
R6294 vdd.n3416 vdd.n3415 0.152939
R6295 vdd.n3417 vdd.n3416 0.152939
R6296 vdd.n3417 vdd.n603 0.152939
R6297 vdd.n3423 vdd.n603 0.152939
R6298 vdd.n3424 vdd.n3423 0.152939
R6299 vdd.n3425 vdd.n3424 0.152939
R6300 vdd.n3425 vdd.n601 0.152939
R6301 vdd.n3430 vdd.n601 0.152939
R6302 vdd.n3193 vdd.n656 0.152939
R6303 vdd.n2121 vdd.n1118 0.152939
R6304 vdd.n1459 vdd.n1458 0.152939
R6305 vdd.n1459 vdd.n1215 0.152939
R6306 vdd.n1473 vdd.n1215 0.152939
R6307 vdd.n1474 vdd.n1473 0.152939
R6308 vdd.n1475 vdd.n1474 0.152939
R6309 vdd.n1475 vdd.n1203 0.152939
R6310 vdd.n1490 vdd.n1203 0.152939
R6311 vdd.n1491 vdd.n1490 0.152939
R6312 vdd.n1492 vdd.n1491 0.152939
R6313 vdd.n1492 vdd.n1193 0.152939
R6314 vdd.n1507 vdd.n1193 0.152939
R6315 vdd.n1508 vdd.n1507 0.152939
R6316 vdd.n1509 vdd.n1508 0.152939
R6317 vdd.n1509 vdd.n1180 0.152939
R6318 vdd.n1523 vdd.n1180 0.152939
R6319 vdd.n1524 vdd.n1523 0.152939
R6320 vdd.n1525 vdd.n1524 0.152939
R6321 vdd.n1525 vdd.n1169 0.152939
R6322 vdd.n1835 vdd.n1169 0.152939
R6323 vdd.n1836 vdd.n1835 0.152939
R6324 vdd.n1837 vdd.n1836 0.152939
R6325 vdd.n1837 vdd.n1158 0.152939
R6326 vdd.n1851 vdd.n1158 0.152939
R6327 vdd.n1852 vdd.n1851 0.152939
R6328 vdd.n1853 vdd.n1852 0.152939
R6329 vdd.n1853 vdd.n1146 0.152939
R6330 vdd.n1868 vdd.n1146 0.152939
R6331 vdd.n1869 vdd.n1868 0.152939
R6332 vdd.n1870 vdd.n1869 0.152939
R6333 vdd.n1870 vdd.n1136 0.152939
R6334 vdd.n1885 vdd.n1136 0.152939
R6335 vdd.n1886 vdd.n1885 0.152939
R6336 vdd.n1889 vdd.n1886 0.152939
R6337 vdd.n1889 vdd.n1888 0.152939
R6338 vdd.n1888 vdd.n1887 0.152939
R6339 vdd.n1449 vdd.n1264 0.152939
R6340 vdd.n1449 vdd.n1448 0.152939
R6341 vdd.n1448 vdd.n1447 0.152939
R6342 vdd.n1447 vdd.n1266 0.152939
R6343 vdd.n1443 vdd.n1266 0.152939
R6344 vdd.n1443 vdd.n1442 0.152939
R6345 vdd.n1442 vdd.n1441 0.152939
R6346 vdd.n1441 vdd.n1271 0.152939
R6347 vdd.n1437 vdd.n1271 0.152939
R6348 vdd.n1437 vdd.n1436 0.152939
R6349 vdd.n1436 vdd.n1435 0.152939
R6350 vdd.n1435 vdd.n1277 0.152939
R6351 vdd.n1431 vdd.n1277 0.152939
R6352 vdd.n1431 vdd.n1430 0.152939
R6353 vdd.n1430 vdd.n1429 0.152939
R6354 vdd.n1429 vdd.n1283 0.152939
R6355 vdd.n1425 vdd.n1283 0.152939
R6356 vdd.n1425 vdd.n1424 0.152939
R6357 vdd.n1424 vdd.n1423 0.152939
R6358 vdd.n1423 vdd.n1289 0.152939
R6359 vdd.n1415 vdd.n1289 0.152939
R6360 vdd.n1415 vdd.n1414 0.152939
R6361 vdd.n1414 vdd.n1413 0.152939
R6362 vdd.n1413 vdd.n1293 0.152939
R6363 vdd.n1409 vdd.n1293 0.152939
R6364 vdd.n1409 vdd.n1408 0.152939
R6365 vdd.n1408 vdd.n1407 0.152939
R6366 vdd.n1407 vdd.n1299 0.152939
R6367 vdd.n1403 vdd.n1299 0.152939
R6368 vdd.n1403 vdd.n1402 0.152939
R6369 vdd.n1402 vdd.n1401 0.152939
R6370 vdd.n1401 vdd.n1305 0.152939
R6371 vdd.n1397 vdd.n1305 0.152939
R6372 vdd.n1397 vdd.n1396 0.152939
R6373 vdd.n1396 vdd.n1395 0.152939
R6374 vdd.n1395 vdd.n1311 0.152939
R6375 vdd.n1391 vdd.n1311 0.152939
R6376 vdd.n1391 vdd.n1390 0.152939
R6377 vdd.n1390 vdd.n1389 0.152939
R6378 vdd.n1389 vdd.n1317 0.152939
R6379 vdd.n1382 vdd.n1317 0.152939
R6380 vdd.n1382 vdd.n1381 0.152939
R6381 vdd.n1381 vdd.n1380 0.152939
R6382 vdd.n1380 vdd.n1322 0.152939
R6383 vdd.n1376 vdd.n1322 0.152939
R6384 vdd.n1376 vdd.n1375 0.152939
R6385 vdd.n1375 vdd.n1374 0.152939
R6386 vdd.n1374 vdd.n1328 0.152939
R6387 vdd.n1370 vdd.n1328 0.152939
R6388 vdd.n1370 vdd.n1369 0.152939
R6389 vdd.n1369 vdd.n1368 0.152939
R6390 vdd.n1368 vdd.n1334 0.152939
R6391 vdd.n1364 vdd.n1334 0.152939
R6392 vdd.n1364 vdd.n1363 0.152939
R6393 vdd.n1363 vdd.n1362 0.152939
R6394 vdd.n1362 vdd.n1340 0.152939
R6395 vdd.n1358 vdd.n1340 0.152939
R6396 vdd.n1358 vdd.n1357 0.152939
R6397 vdd.n1357 vdd.n1356 0.152939
R6398 vdd.n1356 vdd.n1346 0.152939
R6399 vdd.n1352 vdd.n1346 0.152939
R6400 vdd.n1352 vdd.n1227 0.152939
R6401 vdd.n1457 vdd.n1227 0.152939
R6402 vdd.n1465 vdd.n1221 0.152939
R6403 vdd.n1466 vdd.n1465 0.152939
R6404 vdd.n1467 vdd.n1466 0.152939
R6405 vdd.n1467 vdd.n1209 0.152939
R6406 vdd.n1482 vdd.n1209 0.152939
R6407 vdd.n1483 vdd.n1482 0.152939
R6408 vdd.n1484 vdd.n1483 0.152939
R6409 vdd.n1484 vdd.n1198 0.152939
R6410 vdd.n1499 vdd.n1198 0.152939
R6411 vdd.n1500 vdd.n1499 0.152939
R6412 vdd.n1501 vdd.n1500 0.152939
R6413 vdd.n1501 vdd.n1187 0.152939
R6414 vdd.n1515 vdd.n1187 0.152939
R6415 vdd.n1516 vdd.n1515 0.152939
R6416 vdd.n1517 vdd.n1516 0.152939
R6417 vdd.n1517 vdd.n1175 0.152939
R6418 vdd.n1532 vdd.n1175 0.152939
R6419 vdd.n2408 vdd.t178 0.113865
R6420 vdd.n2475 vdd.t130 0.113865
R6421 vdd.n2958 vdd.t133 0.113865
R6422 vdd.n3025 vdd.t157 0.113865
R6423 vdd.n2099 vdd.n1897 0.110256
R6424 vdd.n3124 vdd.n661 0.110256
R6425 vdd.n3193 vdd.n3192 0.110256
R6426 vdd.n2122 vdd.n2121 0.110256
R6427 vdd.n1828 vdd.n1827 0.0695946
R6428 vdd.n3473 vdd.n322 0.0695946
R6429 vdd.n3473 vdd.n3472 0.0695946
R6430 vdd.n1827 vdd.n1532 0.0695946
R6431 vdd.n2099 vdd.n2098 0.0431829
R6432 vdd.n2122 vdd.n1115 0.0431829
R6433 vdd.n3124 vdd.n667 0.0431829
R6434 vdd.n3192 vdd.n748 0.0431829
R6435 vdd vdd.n28 0.00833333
R6436 a_n8300_8799.n181 a_n8300_8799.t127 485.149
R6437 a_n8300_8799.n197 a_n8300_8799.t43 485.149
R6438 a_n8300_8799.n214 a_n8300_8799.t106 485.149
R6439 a_n8300_8799.n130 a_n8300_8799.t92 485.149
R6440 a_n8300_8799.n146 a_n8300_8799.t105 485.149
R6441 a_n8300_8799.n163 a_n8300_8799.t109 485.149
R6442 a_n8300_8799.n191 a_n8300_8799.t90 464.166
R6443 a_n8300_8799.n190 a_n8300_8799.t42 464.166
R6444 a_n8300_8799.n176 a_n8300_8799.t94 464.166
R6445 a_n8300_8799.n189 a_n8300_8799.t93 464.166
R6446 a_n8300_8799.n188 a_n8300_8799.t45 464.166
R6447 a_n8300_8799.n177 a_n8300_8799.t44 464.166
R6448 a_n8300_8799.n187 a_n8300_8799.t112 464.166
R6449 a_n8300_8799.n186 a_n8300_8799.t57 464.166
R6450 a_n8300_8799.n178 a_n8300_8799.t47 464.166
R6451 a_n8300_8799.n185 a_n8300_8799.t116 464.166
R6452 a_n8300_8799.n184 a_n8300_8799.t78 464.166
R6453 a_n8300_8799.n179 a_n8300_8799.t58 464.166
R6454 a_n8300_8799.n183 a_n8300_8799.t132 464.166
R6455 a_n8300_8799.n182 a_n8300_8799.t91 464.166
R6456 a_n8300_8799.n180 a_n8300_8799.t60 464.166
R6457 a_n8300_8799.n207 a_n8300_8799.t103 464.166
R6458 a_n8300_8799.n206 a_n8300_8799.t51 464.166
R6459 a_n8300_8799.n192 a_n8300_8799.t110 464.166
R6460 a_n8300_8799.n205 a_n8300_8799.t107 464.166
R6461 a_n8300_8799.n204 a_n8300_8799.t53 464.166
R6462 a_n8300_8799.n193 a_n8300_8799.t52 464.166
R6463 a_n8300_8799.n203 a_n8300_8799.t126 464.166
R6464 a_n8300_8799.n202 a_n8300_8799.t65 464.166
R6465 a_n8300_8799.n194 a_n8300_8799.t54 464.166
R6466 a_n8300_8799.n201 a_n8300_8799.t128 464.166
R6467 a_n8300_8799.n200 a_n8300_8799.t88 464.166
R6468 a_n8300_8799.n195 a_n8300_8799.t68 464.166
R6469 a_n8300_8799.n199 a_n8300_8799.t46 464.166
R6470 a_n8300_8799.n198 a_n8300_8799.t104 464.166
R6471 a_n8300_8799.n196 a_n8300_8799.t69 464.166
R6472 a_n8300_8799.n224 a_n8300_8799.t62 464.166
R6473 a_n8300_8799.n223 a_n8300_8799.t131 464.166
R6474 a_n8300_8799.n209 a_n8300_8799.t102 464.166
R6475 a_n8300_8799.n222 a_n8300_8799.t124 464.166
R6476 a_n8300_8799.n221 a_n8300_8799.t86 464.166
R6477 a_n8300_8799.n210 a_n8300_8799.t108 464.166
R6478 a_n8300_8799.n220 a_n8300_8799.t55 464.166
R6479 a_n8300_8799.n219 a_n8300_8799.t121 464.166
R6480 a_n8300_8799.n211 a_n8300_8799.t72 464.166
R6481 a_n8300_8799.n218 a_n8300_8799.t117 464.166
R6482 a_n8300_8799.n217 a_n8300_8799.t59 464.166
R6483 a_n8300_8799.n212 a_n8300_8799.t98 464.166
R6484 a_n8300_8799.n216 a_n8300_8799.t50 464.166
R6485 a_n8300_8799.n215 a_n8300_8799.t83 464.166
R6486 a_n8300_8799.n213 a_n8300_8799.t66 464.166
R6487 a_n8300_8799.n129 a_n8300_8799.t123 464.166
R6488 a_n8300_8799.n132 a_n8300_8799.t61 464.166
R6489 a_n8300_8799.n128 a_n8300_8799.t89 464.166
R6490 a_n8300_8799.n133 a_n8300_8799.t119 464.166
R6491 a_n8300_8799.n134 a_n8300_8799.t120 464.166
R6492 a_n8300_8799.n135 a_n8300_8799.t77 464.166
R6493 a_n8300_8799.n136 a_n8300_8799.t101 464.166
R6494 a_n8300_8799.n127 a_n8300_8799.t118 464.166
R6495 a_n8300_8799.n137 a_n8300_8799.t75 464.166
R6496 a_n8300_8799.n138 a_n8300_8799.t76 464.166
R6497 a_n8300_8799.n139 a_n8300_8799.t97 464.166
R6498 a_n8300_8799.n140 a_n8300_8799.t64 464.166
R6499 a_n8300_8799.n126 a_n8300_8799.t63 464.166
R6500 a_n8300_8799.n141 a_n8300_8799.t95 464.166
R6501 a_n8300_8799.n145 a_n8300_8799.t135 464.166
R6502 a_n8300_8799.n148 a_n8300_8799.t70 464.166
R6503 a_n8300_8799.n144 a_n8300_8799.t99 464.166
R6504 a_n8300_8799.n149 a_n8300_8799.t134 464.166
R6505 a_n8300_8799.n150 a_n8300_8799.t133 464.166
R6506 a_n8300_8799.n151 a_n8300_8799.t85 464.166
R6507 a_n8300_8799.n152 a_n8300_8799.t114 464.166
R6508 a_n8300_8799.n143 a_n8300_8799.t130 464.166
R6509 a_n8300_8799.n153 a_n8300_8799.t82 464.166
R6510 a_n8300_8799.n154 a_n8300_8799.t81 464.166
R6511 a_n8300_8799.n155 a_n8300_8799.t113 464.166
R6512 a_n8300_8799.n156 a_n8300_8799.t71 464.166
R6513 a_n8300_8799.n142 a_n8300_8799.t74 464.166
R6514 a_n8300_8799.n157 a_n8300_8799.t111 464.166
R6515 a_n8300_8799.n162 a_n8300_8799.t67 464.166
R6516 a_n8300_8799.n165 a_n8300_8799.t84 464.166
R6517 a_n8300_8799.n161 a_n8300_8799.t49 464.166
R6518 a_n8300_8799.n166 a_n8300_8799.t96 464.166
R6519 a_n8300_8799.n167 a_n8300_8799.t79 464.166
R6520 a_n8300_8799.n168 a_n8300_8799.t115 464.166
R6521 a_n8300_8799.n169 a_n8300_8799.t73 464.166
R6522 a_n8300_8799.n160 a_n8300_8799.t122 464.166
R6523 a_n8300_8799.n170 a_n8300_8799.t56 464.166
R6524 a_n8300_8799.n171 a_n8300_8799.t41 464.166
R6525 a_n8300_8799.n172 a_n8300_8799.t87 464.166
R6526 a_n8300_8799.n173 a_n8300_8799.t125 464.166
R6527 a_n8300_8799.n159 a_n8300_8799.t100 464.166
R6528 a_n8300_8799.n174 a_n8300_8799.t129 464.166
R6529 a_n8300_8799.n54 a_n8300_8799.n34 74.4178
R6530 a_n8300_8799.n182 a_n8300_8799.n54 12.4674
R6531 a_n8300_8799.n53 a_n8300_8799.n34 80.107
R6532 a_n8300_8799.n53 a_n8300_8799.n183 1.08907
R6533 a_n8300_8799.n35 a_n8300_8799.n52 75.3623
R6534 a_n8300_8799.n51 a_n8300_8799.n35 70.3058
R6535 a_n8300_8799.n37 a_n8300_8799.n50 70.1674
R6536 a_n8300_8799.n50 a_n8300_8799.n178 20.9683
R6537 a_n8300_8799.n49 a_n8300_8799.n37 75.0448
R6538 a_n8300_8799.n186 a_n8300_8799.n49 11.2134
R6539 a_n8300_8799.n48 a_n8300_8799.n36 80.4688
R6540 a_n8300_8799.n36 a_n8300_8799.n47 74.73
R6541 a_n8300_8799.n46 a_n8300_8799.n38 70.1674
R6542 a_n8300_8799.n189 a_n8300_8799.n46 20.9683
R6543 a_n8300_8799.n38 a_n8300_8799.n45 70.5844
R6544 a_n8300_8799.n45 a_n8300_8799.n176 20.1342
R6545 a_n8300_8799.n44 a_n8300_8799.n39 75.6825
R6546 a_n8300_8799.n190 a_n8300_8799.n44 9.93802
R6547 a_n8300_8799.n39 a_n8300_8799.n191 161.3
R6548 a_n8300_8799.n65 a_n8300_8799.n28 74.4178
R6549 a_n8300_8799.n198 a_n8300_8799.n65 12.4674
R6550 a_n8300_8799.n64 a_n8300_8799.n28 80.107
R6551 a_n8300_8799.n64 a_n8300_8799.n199 1.08907
R6552 a_n8300_8799.n29 a_n8300_8799.n63 75.3623
R6553 a_n8300_8799.n62 a_n8300_8799.n29 70.3058
R6554 a_n8300_8799.n31 a_n8300_8799.n61 70.1674
R6555 a_n8300_8799.n61 a_n8300_8799.n194 20.9683
R6556 a_n8300_8799.n60 a_n8300_8799.n31 75.0448
R6557 a_n8300_8799.n202 a_n8300_8799.n60 11.2134
R6558 a_n8300_8799.n59 a_n8300_8799.n30 80.4688
R6559 a_n8300_8799.n30 a_n8300_8799.n58 74.73
R6560 a_n8300_8799.n57 a_n8300_8799.n32 70.1674
R6561 a_n8300_8799.n205 a_n8300_8799.n57 20.9683
R6562 a_n8300_8799.n32 a_n8300_8799.n56 70.5844
R6563 a_n8300_8799.n56 a_n8300_8799.n192 20.1342
R6564 a_n8300_8799.n55 a_n8300_8799.n33 75.6825
R6565 a_n8300_8799.n206 a_n8300_8799.n55 9.93802
R6566 a_n8300_8799.n33 a_n8300_8799.n207 161.3
R6567 a_n8300_8799.n76 a_n8300_8799.n22 74.4178
R6568 a_n8300_8799.n215 a_n8300_8799.n76 12.4674
R6569 a_n8300_8799.n75 a_n8300_8799.n22 80.107
R6570 a_n8300_8799.n75 a_n8300_8799.n216 1.08907
R6571 a_n8300_8799.n23 a_n8300_8799.n74 75.3623
R6572 a_n8300_8799.n73 a_n8300_8799.n23 70.3058
R6573 a_n8300_8799.n25 a_n8300_8799.n72 70.1674
R6574 a_n8300_8799.n72 a_n8300_8799.n211 20.9683
R6575 a_n8300_8799.n71 a_n8300_8799.n25 75.0448
R6576 a_n8300_8799.n219 a_n8300_8799.n71 11.2134
R6577 a_n8300_8799.n70 a_n8300_8799.n24 80.4688
R6578 a_n8300_8799.n24 a_n8300_8799.n69 74.73
R6579 a_n8300_8799.n68 a_n8300_8799.n26 70.1674
R6580 a_n8300_8799.n222 a_n8300_8799.n68 20.9683
R6581 a_n8300_8799.n26 a_n8300_8799.n67 70.5844
R6582 a_n8300_8799.n67 a_n8300_8799.n209 20.1342
R6583 a_n8300_8799.n66 a_n8300_8799.n27 75.6825
R6584 a_n8300_8799.n223 a_n8300_8799.n66 9.93802
R6585 a_n8300_8799.n27 a_n8300_8799.n224 161.3
R6586 a_n8300_8799.n17 a_n8300_8799.n87 70.1674
R6587 a_n8300_8799.n141 a_n8300_8799.n87 20.9683
R6588 a_n8300_8799.n86 a_n8300_8799.n17 74.4178
R6589 a_n8300_8799.n86 a_n8300_8799.n126 12.4674
R6590 a_n8300_8799.n16 a_n8300_8799.n85 80.107
R6591 a_n8300_8799.n140 a_n8300_8799.n85 1.08907
R6592 a_n8300_8799.n84 a_n8300_8799.n16 75.3623
R6593 a_n8300_8799.n18 a_n8300_8799.n83 70.3058
R6594 a_n8300_8799.n82 a_n8300_8799.n18 70.1674
R6595 a_n8300_8799.n82 a_n8300_8799.n127 20.9683
R6596 a_n8300_8799.n19 a_n8300_8799.n81 75.0448
R6597 a_n8300_8799.n136 a_n8300_8799.n81 11.2134
R6598 a_n8300_8799.n80 a_n8300_8799.n19 80.4688
R6599 a_n8300_8799.n20 a_n8300_8799.n79 74.73
R6600 a_n8300_8799.n78 a_n8300_8799.n20 70.1674
R6601 a_n8300_8799.n78 a_n8300_8799.n128 20.9683
R6602 a_n8300_8799.n21 a_n8300_8799.n77 70.5844
R6603 a_n8300_8799.n132 a_n8300_8799.n77 20.1342
R6604 a_n8300_8799.n131 a_n8300_8799.n21 161.3
R6605 a_n8300_8799.n11 a_n8300_8799.n98 70.1674
R6606 a_n8300_8799.n157 a_n8300_8799.n98 20.9683
R6607 a_n8300_8799.n97 a_n8300_8799.n11 74.4178
R6608 a_n8300_8799.n97 a_n8300_8799.n142 12.4674
R6609 a_n8300_8799.n10 a_n8300_8799.n96 80.107
R6610 a_n8300_8799.n156 a_n8300_8799.n96 1.08907
R6611 a_n8300_8799.n95 a_n8300_8799.n10 75.3623
R6612 a_n8300_8799.n12 a_n8300_8799.n94 70.3058
R6613 a_n8300_8799.n93 a_n8300_8799.n12 70.1674
R6614 a_n8300_8799.n93 a_n8300_8799.n143 20.9683
R6615 a_n8300_8799.n13 a_n8300_8799.n92 75.0448
R6616 a_n8300_8799.n152 a_n8300_8799.n92 11.2134
R6617 a_n8300_8799.n91 a_n8300_8799.n13 80.4688
R6618 a_n8300_8799.n14 a_n8300_8799.n90 74.73
R6619 a_n8300_8799.n89 a_n8300_8799.n14 70.1674
R6620 a_n8300_8799.n89 a_n8300_8799.n144 20.9683
R6621 a_n8300_8799.n15 a_n8300_8799.n88 70.5844
R6622 a_n8300_8799.n148 a_n8300_8799.n88 20.1342
R6623 a_n8300_8799.n147 a_n8300_8799.n15 161.3
R6624 a_n8300_8799.n5 a_n8300_8799.n109 70.1674
R6625 a_n8300_8799.n174 a_n8300_8799.n109 20.9683
R6626 a_n8300_8799.n108 a_n8300_8799.n5 74.4178
R6627 a_n8300_8799.n108 a_n8300_8799.n159 12.4674
R6628 a_n8300_8799.n4 a_n8300_8799.n107 80.107
R6629 a_n8300_8799.n173 a_n8300_8799.n107 1.08907
R6630 a_n8300_8799.n106 a_n8300_8799.n4 75.3623
R6631 a_n8300_8799.n6 a_n8300_8799.n105 70.3058
R6632 a_n8300_8799.n104 a_n8300_8799.n6 70.1674
R6633 a_n8300_8799.n104 a_n8300_8799.n160 20.9683
R6634 a_n8300_8799.n7 a_n8300_8799.n103 75.0448
R6635 a_n8300_8799.n169 a_n8300_8799.n103 11.2134
R6636 a_n8300_8799.n102 a_n8300_8799.n7 80.4688
R6637 a_n8300_8799.n8 a_n8300_8799.n101 74.73
R6638 a_n8300_8799.n100 a_n8300_8799.n8 70.1674
R6639 a_n8300_8799.n100 a_n8300_8799.n161 20.9683
R6640 a_n8300_8799.n9 a_n8300_8799.n99 70.5844
R6641 a_n8300_8799.n165 a_n8300_8799.n99 20.1342
R6642 a_n8300_8799.n164 a_n8300_8799.n9 161.3
R6643 a_n8300_8799.n43 a_n8300_8799.n110 98.9633
R6644 a_n8300_8799.n40 a_n8300_8799.n111 98.9631
R6645 a_n8300_8799.n42 a_n8300_8799.n229 98.6055
R6646 a_n8300_8799.n42 a_n8300_8799.n230 98.6055
R6647 a_n8300_8799.n43 a_n8300_8799.n231 98.6055
R6648 a_n8300_8799.n40 a_n8300_8799.n112 98.6055
R6649 a_n8300_8799.n40 a_n8300_8799.n113 98.6055
R6650 a_n8300_8799.n41 a_n8300_8799.n114 98.6055
R6651 a_n8300_8799.n41 a_n8300_8799.n115 98.6055
R6652 a_n8300_8799.n232 a_n8300_8799.n43 98.6054
R6653 a_n8300_8799.n3 a_n8300_8799.n116 81.4626
R6654 a_n8300_8799.n1 a_n8300_8799.n122 81.4626
R6655 a_n8300_8799.n0 a_n8300_8799.n119 81.4626
R6656 a_n8300_8799.n2 a_n8300_8799.n124 80.9324
R6657 a_n8300_8799.n2 a_n8300_8799.n125 80.9324
R6658 a_n8300_8799.n3 a_n8300_8799.n118 80.9324
R6659 a_n8300_8799.n3 a_n8300_8799.n117 80.9324
R6660 a_n8300_8799.n1 a_n8300_8799.n123 80.9324
R6661 a_n8300_8799.n1 a_n8300_8799.n121 80.9324
R6662 a_n8300_8799.n0 a_n8300_8799.n120 80.9324
R6663 a_n8300_8799.n34 a_n8300_8799.n181 70.4033
R6664 a_n8300_8799.n28 a_n8300_8799.n197 70.4033
R6665 a_n8300_8799.n22 a_n8300_8799.n214 70.4033
R6666 a_n8300_8799.n21 a_n8300_8799.n130 70.4033
R6667 a_n8300_8799.n15 a_n8300_8799.n146 70.4033
R6668 a_n8300_8799.n9 a_n8300_8799.n163 70.4033
R6669 a_n8300_8799.n191 a_n8300_8799.n190 48.2005
R6670 a_n8300_8799.n46 a_n8300_8799.n188 20.9683
R6671 a_n8300_8799.n187 a_n8300_8799.n186 48.2005
R6672 a_n8300_8799.n185 a_n8300_8799.n50 20.9683
R6673 a_n8300_8799.n183 a_n8300_8799.n179 48.2005
R6674 a_n8300_8799.n207 a_n8300_8799.n206 48.2005
R6675 a_n8300_8799.n57 a_n8300_8799.n204 20.9683
R6676 a_n8300_8799.n203 a_n8300_8799.n202 48.2005
R6677 a_n8300_8799.n201 a_n8300_8799.n61 20.9683
R6678 a_n8300_8799.n199 a_n8300_8799.n195 48.2005
R6679 a_n8300_8799.n224 a_n8300_8799.n223 48.2005
R6680 a_n8300_8799.n68 a_n8300_8799.n221 20.9683
R6681 a_n8300_8799.n220 a_n8300_8799.n219 48.2005
R6682 a_n8300_8799.n218 a_n8300_8799.n72 20.9683
R6683 a_n8300_8799.n216 a_n8300_8799.n212 48.2005
R6684 a_n8300_8799.n133 a_n8300_8799.n78 20.9683
R6685 a_n8300_8799.n136 a_n8300_8799.n135 48.2005
R6686 a_n8300_8799.n137 a_n8300_8799.n82 20.9683
R6687 a_n8300_8799.n140 a_n8300_8799.n139 48.2005
R6688 a_n8300_8799.t40 a_n8300_8799.n87 485.135
R6689 a_n8300_8799.n149 a_n8300_8799.n89 20.9683
R6690 a_n8300_8799.n152 a_n8300_8799.n151 48.2005
R6691 a_n8300_8799.n153 a_n8300_8799.n93 20.9683
R6692 a_n8300_8799.n156 a_n8300_8799.n155 48.2005
R6693 a_n8300_8799.t48 a_n8300_8799.n98 485.135
R6694 a_n8300_8799.n166 a_n8300_8799.n100 20.9683
R6695 a_n8300_8799.n169 a_n8300_8799.n168 48.2005
R6696 a_n8300_8799.n170 a_n8300_8799.n104 20.9683
R6697 a_n8300_8799.n173 a_n8300_8799.n172 48.2005
R6698 a_n8300_8799.t80 a_n8300_8799.n109 485.135
R6699 a_n8300_8799.n48 a_n8300_8799.n177 47.835
R6700 a_n8300_8799.n51 a_n8300_8799.n184 20.6913
R6701 a_n8300_8799.n59 a_n8300_8799.n193 47.835
R6702 a_n8300_8799.n62 a_n8300_8799.n200 20.6913
R6703 a_n8300_8799.n70 a_n8300_8799.n210 47.835
R6704 a_n8300_8799.n73 a_n8300_8799.n217 20.6913
R6705 a_n8300_8799.n134 a_n8300_8799.n80 47.835
R6706 a_n8300_8799.n138 a_n8300_8799.n83 20.6913
R6707 a_n8300_8799.n150 a_n8300_8799.n91 47.835
R6708 a_n8300_8799.n154 a_n8300_8799.n94 20.6913
R6709 a_n8300_8799.n167 a_n8300_8799.n102 47.835
R6710 a_n8300_8799.n171 a_n8300_8799.n105 20.6913
R6711 a_n8300_8799.n189 a_n8300_8799.n45 22.3251
R6712 a_n8300_8799.n205 a_n8300_8799.n56 22.3251
R6713 a_n8300_8799.n222 a_n8300_8799.n67 22.3251
R6714 a_n8300_8799.n128 a_n8300_8799.n77 22.3251
R6715 a_n8300_8799.n144 a_n8300_8799.n88 22.3251
R6716 a_n8300_8799.n161 a_n8300_8799.n99 22.3251
R6717 a_n8300_8799.n2 a_n8300_8799.n1 33.5285
R6718 a_n8300_8799.n228 a_n8300_8799.n41 33.0756
R6719 a_n8300_8799.n54 a_n8300_8799.n180 33.6462
R6720 a_n8300_8799.n65 a_n8300_8799.n196 33.6462
R6721 a_n8300_8799.n76 a_n8300_8799.n213 33.6462
R6722 a_n8300_8799.n132 a_n8300_8799.n131 27.0217
R6723 a_n8300_8799.n141 a_n8300_8799.n86 33.6462
R6724 a_n8300_8799.n148 a_n8300_8799.n147 27.0217
R6725 a_n8300_8799.n157 a_n8300_8799.n97 33.6462
R6726 a_n8300_8799.n165 a_n8300_8799.n164 27.0217
R6727 a_n8300_8799.n174 a_n8300_8799.n108 33.6462
R6728 a_n8300_8799.n47 a_n8300_8799.n177 11.843
R6729 a_n8300_8799.n184 a_n8300_8799.n52 36.139
R6730 a_n8300_8799.n58 a_n8300_8799.n193 11.843
R6731 a_n8300_8799.n200 a_n8300_8799.n63 36.139
R6732 a_n8300_8799.n69 a_n8300_8799.n210 11.843
R6733 a_n8300_8799.n217 a_n8300_8799.n74 36.139
R6734 a_n8300_8799.n134 a_n8300_8799.n79 11.843
R6735 a_n8300_8799.n138 a_n8300_8799.n84 36.139
R6736 a_n8300_8799.n150 a_n8300_8799.n90 11.843
R6737 a_n8300_8799.n154 a_n8300_8799.n95 36.139
R6738 a_n8300_8799.n167 a_n8300_8799.n101 11.843
R6739 a_n8300_8799.n171 a_n8300_8799.n106 36.139
R6740 a_n8300_8799.n49 a_n8300_8799.n178 35.3134
R6741 a_n8300_8799.n60 a_n8300_8799.n194 35.3134
R6742 a_n8300_8799.n71 a_n8300_8799.n211 35.3134
R6743 a_n8300_8799.n127 a_n8300_8799.n81 35.3134
R6744 a_n8300_8799.n143 a_n8300_8799.n92 35.3134
R6745 a_n8300_8799.n160 a_n8300_8799.n103 35.3134
R6746 a_n8300_8799.n188 a_n8300_8799.n47 34.4824
R6747 a_n8300_8799.n52 a_n8300_8799.n179 10.5784
R6748 a_n8300_8799.n204 a_n8300_8799.n58 34.4824
R6749 a_n8300_8799.n63 a_n8300_8799.n195 10.5784
R6750 a_n8300_8799.n221 a_n8300_8799.n69 34.4824
R6751 a_n8300_8799.n74 a_n8300_8799.n212 10.5784
R6752 a_n8300_8799.n79 a_n8300_8799.n133 34.4824
R6753 a_n8300_8799.n139 a_n8300_8799.n84 10.5784
R6754 a_n8300_8799.n90 a_n8300_8799.n149 34.4824
R6755 a_n8300_8799.n155 a_n8300_8799.n95 10.5784
R6756 a_n8300_8799.n101 a_n8300_8799.n166 34.4824
R6757 a_n8300_8799.n172 a_n8300_8799.n106 10.5784
R6758 a_n8300_8799.n44 a_n8300_8799.n176 36.9592
R6759 a_n8300_8799.n55 a_n8300_8799.n192 36.9592
R6760 a_n8300_8799.n66 a_n8300_8799.n209 36.9592
R6761 a_n8300_8799.n131 a_n8300_8799.n129 21.1793
R6762 a_n8300_8799.n147 a_n8300_8799.n145 21.1793
R6763 a_n8300_8799.n164 a_n8300_8799.n162 21.1793
R6764 a_n8300_8799.n181 a_n8300_8799.n180 20.9576
R6765 a_n8300_8799.n197 a_n8300_8799.n196 20.9576
R6766 a_n8300_8799.n214 a_n8300_8799.n213 20.9576
R6767 a_n8300_8799.n130 a_n8300_8799.n129 20.9576
R6768 a_n8300_8799.n146 a_n8300_8799.n145 20.9576
R6769 a_n8300_8799.n163 a_n8300_8799.n162 20.9576
R6770 a_n8300_8799.n42 a_n8300_8799.n228 19.6671
R6771 a_n8300_8799.n227 a_n8300_8799.n3 12.3339
R6772 a_n8300_8799.n228 a_n8300_8799.n227 11.4887
R6773 a_n8300_8799.n208 a_n8300_8799.n39 9.07815
R6774 a_n8300_8799.n158 a_n8300_8799.n17 9.07815
R6775 a_n8300_8799.n226 a_n8300_8799.n175 7.10923
R6776 a_n8300_8799.n226 a_n8300_8799.n225 6.68968
R6777 a_n8300_8799.n208 a_n8300_8799.n33 4.9702
R6778 a_n8300_8799.n225 a_n8300_8799.n27 4.9702
R6779 a_n8300_8799.n158 a_n8300_8799.n11 4.9702
R6780 a_n8300_8799.n175 a_n8300_8799.n5 4.9702
R6781 a_n8300_8799.n225 a_n8300_8799.n208 4.10845
R6782 a_n8300_8799.n175 a_n8300_8799.n158 4.10845
R6783 a_n8300_8799.n229 a_n8300_8799.t21 3.61217
R6784 a_n8300_8799.n229 a_n8300_8799.t15 3.61217
R6785 a_n8300_8799.n230 a_n8300_8799.t27 3.61217
R6786 a_n8300_8799.n230 a_n8300_8799.t20 3.61217
R6787 a_n8300_8799.n231 a_n8300_8799.t16 3.61217
R6788 a_n8300_8799.n231 a_n8300_8799.t13 3.61217
R6789 a_n8300_8799.n110 a_n8300_8799.t11 3.61217
R6790 a_n8300_8799.n110 a_n8300_8799.t14 3.61217
R6791 a_n8300_8799.n111 a_n8300_8799.t17 3.61217
R6792 a_n8300_8799.n111 a_n8300_8799.t10 3.61217
R6793 a_n8300_8799.n112 a_n8300_8799.t23 3.61217
R6794 a_n8300_8799.n112 a_n8300_8799.t24 3.61217
R6795 a_n8300_8799.n113 a_n8300_8799.t18 3.61217
R6796 a_n8300_8799.n113 a_n8300_8799.t26 3.61217
R6797 a_n8300_8799.n114 a_n8300_8799.t12 3.61217
R6798 a_n8300_8799.n114 a_n8300_8799.t25 3.61217
R6799 a_n8300_8799.n115 a_n8300_8799.t22 3.61217
R6800 a_n8300_8799.n115 a_n8300_8799.t19 3.61217
R6801 a_n8300_8799.n232 a_n8300_8799.t28 3.61217
R6802 a_n8300_8799.t9 a_n8300_8799.n232 3.61217
R6803 a_n8300_8799.n227 a_n8300_8799.n226 3.4105
R6804 a_n8300_8799.n124 a_n8300_8799.t3 2.82907
R6805 a_n8300_8799.n124 a_n8300_8799.t29 2.82907
R6806 a_n8300_8799.n125 a_n8300_8799.t31 2.82907
R6807 a_n8300_8799.n125 a_n8300_8799.t4 2.82907
R6808 a_n8300_8799.n118 a_n8300_8799.t30 2.82907
R6809 a_n8300_8799.n118 a_n8300_8799.t5 2.82907
R6810 a_n8300_8799.n117 a_n8300_8799.t7 2.82907
R6811 a_n8300_8799.n117 a_n8300_8799.t32 2.82907
R6812 a_n8300_8799.n116 a_n8300_8799.t0 2.82907
R6813 a_n8300_8799.n116 a_n8300_8799.t39 2.82907
R6814 a_n8300_8799.n122 a_n8300_8799.t8 2.82907
R6815 a_n8300_8799.n122 a_n8300_8799.t37 2.82907
R6816 a_n8300_8799.n123 a_n8300_8799.t36 2.82907
R6817 a_n8300_8799.n123 a_n8300_8799.t6 2.82907
R6818 a_n8300_8799.n121 a_n8300_8799.t1 2.82907
R6819 a_n8300_8799.n121 a_n8300_8799.t2 2.82907
R6820 a_n8300_8799.n120 a_n8300_8799.t34 2.82907
R6821 a_n8300_8799.n120 a_n8300_8799.t35 2.82907
R6822 a_n8300_8799.n119 a_n8300_8799.t33 2.82907
R6823 a_n8300_8799.n119 a_n8300_8799.t38 2.82907
R6824 a_n8300_8799.n53 a_n8300_8799.n182 47.0982
R6825 a_n8300_8799.n64 a_n8300_8799.n198 47.0982
R6826 a_n8300_8799.n75 a_n8300_8799.n215 47.0982
R6827 a_n8300_8799.n126 a_n8300_8799.n85 47.0982
R6828 a_n8300_8799.n142 a_n8300_8799.n96 47.0982
R6829 a_n8300_8799.n159 a_n8300_8799.n107 47.0982
R6830 a_n8300_8799.n48 a_n8300_8799.n187 0.365327
R6831 a_n8300_8799.n185 a_n8300_8799.n51 21.4216
R6832 a_n8300_8799.n59 a_n8300_8799.n203 0.365327
R6833 a_n8300_8799.n201 a_n8300_8799.n62 21.4216
R6834 a_n8300_8799.n70 a_n8300_8799.n220 0.365327
R6835 a_n8300_8799.n218 a_n8300_8799.n73 21.4216
R6836 a_n8300_8799.n135 a_n8300_8799.n80 0.365327
R6837 a_n8300_8799.n83 a_n8300_8799.n137 21.4216
R6838 a_n8300_8799.n151 a_n8300_8799.n91 0.365327
R6839 a_n8300_8799.n94 a_n8300_8799.n153 21.4216
R6840 a_n8300_8799.n168 a_n8300_8799.n102 0.365327
R6841 a_n8300_8799.n105 a_n8300_8799.n170 21.4216
R6842 a_n8300_8799.n3 a_n8300_8799.n2 1.59102
R6843 a_n8300_8799.n35 a_n8300_8799.n34 1.13686
R6844 a_n8300_8799.n29 a_n8300_8799.n28 1.13686
R6845 a_n8300_8799.n23 a_n8300_8799.n22 1.13686
R6846 a_n8300_8799.n17 a_n8300_8799.n16 1.13686
R6847 a_n8300_8799.n11 a_n8300_8799.n10 1.13686
R6848 a_n8300_8799.n5 a_n8300_8799.n4 1.13686
R6849 a_n8300_8799.n43 a_n8300_8799.n42 1.07378
R6850 a_n8300_8799.n41 a_n8300_8799.n40 1.07378
R6851 a_n8300_8799.n1 a_n8300_8799.n0 1.06084
R6852 a_n8300_8799.n39 a_n8300_8799.n38 0.758076
R6853 a_n8300_8799.n36 a_n8300_8799.n38 0.758076
R6854 a_n8300_8799.n37 a_n8300_8799.n36 0.758076
R6855 a_n8300_8799.n37 a_n8300_8799.n35 0.758076
R6856 a_n8300_8799.n33 a_n8300_8799.n32 0.758076
R6857 a_n8300_8799.n30 a_n8300_8799.n32 0.758076
R6858 a_n8300_8799.n31 a_n8300_8799.n30 0.758076
R6859 a_n8300_8799.n31 a_n8300_8799.n29 0.758076
R6860 a_n8300_8799.n27 a_n8300_8799.n26 0.758076
R6861 a_n8300_8799.n24 a_n8300_8799.n26 0.758076
R6862 a_n8300_8799.n25 a_n8300_8799.n24 0.758076
R6863 a_n8300_8799.n25 a_n8300_8799.n23 0.758076
R6864 a_n8300_8799.n20 a_n8300_8799.n21 0.758076
R6865 a_n8300_8799.n19 a_n8300_8799.n20 0.758076
R6866 a_n8300_8799.n18 a_n8300_8799.n19 0.758076
R6867 a_n8300_8799.n16 a_n8300_8799.n18 0.758076
R6868 a_n8300_8799.n14 a_n8300_8799.n15 0.758076
R6869 a_n8300_8799.n13 a_n8300_8799.n14 0.758076
R6870 a_n8300_8799.n12 a_n8300_8799.n13 0.758076
R6871 a_n8300_8799.n10 a_n8300_8799.n12 0.758076
R6872 a_n8300_8799.n8 a_n8300_8799.n9 0.758076
R6873 a_n8300_8799.n7 a_n8300_8799.n8 0.758076
R6874 a_n8300_8799.n6 a_n8300_8799.n7 0.758076
R6875 a_n8300_8799.n4 a_n8300_8799.n6 0.758076
R6876 CSoutput.n19 CSoutput.t145 184.661
R6877 CSoutput.n78 CSoutput.n77 165.8
R6878 CSoutput.n76 CSoutput.n0 165.8
R6879 CSoutput.n75 CSoutput.n74 165.8
R6880 CSoutput.n73 CSoutput.n72 165.8
R6881 CSoutput.n71 CSoutput.n2 165.8
R6882 CSoutput.n69 CSoutput.n68 165.8
R6883 CSoutput.n67 CSoutput.n3 165.8
R6884 CSoutput.n66 CSoutput.n65 165.8
R6885 CSoutput.n63 CSoutput.n4 165.8
R6886 CSoutput.n61 CSoutput.n60 165.8
R6887 CSoutput.n59 CSoutput.n5 165.8
R6888 CSoutput.n58 CSoutput.n57 165.8
R6889 CSoutput.n55 CSoutput.n6 165.8
R6890 CSoutput.n54 CSoutput.n53 165.8
R6891 CSoutput.n52 CSoutput.n51 165.8
R6892 CSoutput.n50 CSoutput.n8 165.8
R6893 CSoutput.n48 CSoutput.n47 165.8
R6894 CSoutput.n46 CSoutput.n9 165.8
R6895 CSoutput.n45 CSoutput.n44 165.8
R6896 CSoutput.n42 CSoutput.n10 165.8
R6897 CSoutput.n41 CSoutput.n40 165.8
R6898 CSoutput.n39 CSoutput.n38 165.8
R6899 CSoutput.n37 CSoutput.n12 165.8
R6900 CSoutput.n35 CSoutput.n34 165.8
R6901 CSoutput.n33 CSoutput.n13 165.8
R6902 CSoutput.n32 CSoutput.n31 165.8
R6903 CSoutput.n29 CSoutput.n14 165.8
R6904 CSoutput.n28 CSoutput.n27 165.8
R6905 CSoutput.n26 CSoutput.n25 165.8
R6906 CSoutput.n24 CSoutput.n16 165.8
R6907 CSoutput.n22 CSoutput.n21 165.8
R6908 CSoutput.n20 CSoutput.n17 165.8
R6909 CSoutput.n77 CSoutput.t148 162.194
R6910 CSoutput.n18 CSoutput.t147 120.501
R6911 CSoutput.n23 CSoutput.t158 120.501
R6912 CSoutput.n15 CSoutput.t155 120.501
R6913 CSoutput.n30 CSoutput.t149 120.501
R6914 CSoutput.n36 CSoutput.t160 120.501
R6915 CSoutput.n11 CSoutput.t162 120.501
R6916 CSoutput.n43 CSoutput.t151 120.501
R6917 CSoutput.n49 CSoutput.t163 120.501
R6918 CSoutput.n7 CSoutput.t165 120.501
R6919 CSoutput.n56 CSoutput.t159 120.501
R6920 CSoutput.n62 CSoutput.t150 120.501
R6921 CSoutput.n64 CSoutput.t144 120.501
R6922 CSoutput.n70 CSoutput.t161 120.501
R6923 CSoutput.n1 CSoutput.t156 120.501
R6924 CSoutput.n310 CSoutput.n308 103.469
R6925 CSoutput.n294 CSoutput.n292 103.469
R6926 CSoutput.n279 CSoutput.n277 103.469
R6927 CSoutput.n112 CSoutput.n110 103.469
R6928 CSoutput.n96 CSoutput.n94 103.469
R6929 CSoutput.n81 CSoutput.n79 103.469
R6930 CSoutput.n320 CSoutput.n319 103.111
R6931 CSoutput.n318 CSoutput.n317 103.111
R6932 CSoutput.n316 CSoutput.n315 103.111
R6933 CSoutput.n314 CSoutput.n313 103.111
R6934 CSoutput.n312 CSoutput.n311 103.111
R6935 CSoutput.n310 CSoutput.n309 103.111
R6936 CSoutput.n306 CSoutput.n305 103.111
R6937 CSoutput.n304 CSoutput.n303 103.111
R6938 CSoutput.n302 CSoutput.n301 103.111
R6939 CSoutput.n300 CSoutput.n299 103.111
R6940 CSoutput.n298 CSoutput.n297 103.111
R6941 CSoutput.n296 CSoutput.n295 103.111
R6942 CSoutput.n294 CSoutput.n293 103.111
R6943 CSoutput.n291 CSoutput.n290 103.111
R6944 CSoutput.n289 CSoutput.n288 103.111
R6945 CSoutput.n287 CSoutput.n286 103.111
R6946 CSoutput.n285 CSoutput.n284 103.111
R6947 CSoutput.n283 CSoutput.n282 103.111
R6948 CSoutput.n281 CSoutput.n280 103.111
R6949 CSoutput.n279 CSoutput.n278 103.111
R6950 CSoutput.n112 CSoutput.n111 103.111
R6951 CSoutput.n114 CSoutput.n113 103.111
R6952 CSoutput.n116 CSoutput.n115 103.111
R6953 CSoutput.n118 CSoutput.n117 103.111
R6954 CSoutput.n120 CSoutput.n119 103.111
R6955 CSoutput.n122 CSoutput.n121 103.111
R6956 CSoutput.n124 CSoutput.n123 103.111
R6957 CSoutput.n96 CSoutput.n95 103.111
R6958 CSoutput.n98 CSoutput.n97 103.111
R6959 CSoutput.n100 CSoutput.n99 103.111
R6960 CSoutput.n102 CSoutput.n101 103.111
R6961 CSoutput.n104 CSoutput.n103 103.111
R6962 CSoutput.n106 CSoutput.n105 103.111
R6963 CSoutput.n108 CSoutput.n107 103.111
R6964 CSoutput.n81 CSoutput.n80 103.111
R6965 CSoutput.n83 CSoutput.n82 103.111
R6966 CSoutput.n85 CSoutput.n84 103.111
R6967 CSoutput.n87 CSoutput.n86 103.111
R6968 CSoutput.n89 CSoutput.n88 103.111
R6969 CSoutput.n91 CSoutput.n90 103.111
R6970 CSoutput.n93 CSoutput.n92 103.111
R6971 CSoutput.n322 CSoutput.n321 103.111
R6972 CSoutput.n338 CSoutput.n336 81.5057
R6973 CSoutput.n327 CSoutput.n325 81.5057
R6974 CSoutput.n362 CSoutput.n360 81.5057
R6975 CSoutput.n351 CSoutput.n349 81.5057
R6976 CSoutput.n346 CSoutput.n345 80.9324
R6977 CSoutput.n344 CSoutput.n343 80.9324
R6978 CSoutput.n342 CSoutput.n341 80.9324
R6979 CSoutput.n340 CSoutput.n339 80.9324
R6980 CSoutput.n338 CSoutput.n337 80.9324
R6981 CSoutput.n335 CSoutput.n334 80.9324
R6982 CSoutput.n333 CSoutput.n332 80.9324
R6983 CSoutput.n331 CSoutput.n330 80.9324
R6984 CSoutput.n329 CSoutput.n328 80.9324
R6985 CSoutput.n327 CSoutput.n326 80.9324
R6986 CSoutput.n362 CSoutput.n361 80.9324
R6987 CSoutput.n364 CSoutput.n363 80.9324
R6988 CSoutput.n366 CSoutput.n365 80.9324
R6989 CSoutput.n368 CSoutput.n367 80.9324
R6990 CSoutput.n370 CSoutput.n369 80.9324
R6991 CSoutput.n351 CSoutput.n350 80.9324
R6992 CSoutput.n353 CSoutput.n352 80.9324
R6993 CSoutput.n355 CSoutput.n354 80.9324
R6994 CSoutput.n357 CSoutput.n356 80.9324
R6995 CSoutput.n359 CSoutput.n358 80.9324
R6996 CSoutput.n25 CSoutput.n24 48.1486
R6997 CSoutput.n69 CSoutput.n3 48.1486
R6998 CSoutput.n38 CSoutput.n37 48.1486
R6999 CSoutput.n42 CSoutput.n41 48.1486
R7000 CSoutput.n51 CSoutput.n50 48.1486
R7001 CSoutput.n55 CSoutput.n54 48.1486
R7002 CSoutput.n22 CSoutput.n17 46.462
R7003 CSoutput.n72 CSoutput.n71 46.462
R7004 CSoutput.n20 CSoutput.n19 44.9055
R7005 CSoutput.n29 CSoutput.n28 43.7635
R7006 CSoutput.n65 CSoutput.n63 43.7635
R7007 CSoutput.n35 CSoutput.n13 41.7396
R7008 CSoutput.n57 CSoutput.n5 41.7396
R7009 CSoutput.n44 CSoutput.n9 37.0171
R7010 CSoutput.n48 CSoutput.n9 37.0171
R7011 CSoutput.n76 CSoutput.n75 34.9932
R7012 CSoutput.n31 CSoutput.n13 32.2947
R7013 CSoutput.n61 CSoutput.n5 32.2947
R7014 CSoutput.n30 CSoutput.n29 29.6014
R7015 CSoutput.n63 CSoutput.n62 29.6014
R7016 CSoutput.n19 CSoutput.n18 28.4085
R7017 CSoutput.n18 CSoutput.n17 25.1176
R7018 CSoutput.n72 CSoutput.n1 25.1176
R7019 CSoutput.n43 CSoutput.n42 22.0922
R7020 CSoutput.n50 CSoutput.n49 22.0922
R7021 CSoutput.n77 CSoutput.n76 21.8586
R7022 CSoutput.n37 CSoutput.n36 18.9681
R7023 CSoutput.n56 CSoutput.n55 18.9681
R7024 CSoutput.n25 CSoutput.n15 17.6292
R7025 CSoutput.n64 CSoutput.n3 17.6292
R7026 CSoutput.n24 CSoutput.n23 15.844
R7027 CSoutput.n70 CSoutput.n69 15.844
R7028 CSoutput.n38 CSoutput.n11 14.5051
R7029 CSoutput.n54 CSoutput.n7 14.5051
R7030 CSoutput.n373 CSoutput.n78 11.6139
R7031 CSoutput.n41 CSoutput.n11 11.3811
R7032 CSoutput.n51 CSoutput.n7 11.3811
R7033 CSoutput.n23 CSoutput.n22 10.0422
R7034 CSoutput.n71 CSoutput.n70 10.0422
R7035 CSoutput.n307 CSoutput.n291 9.25285
R7036 CSoutput.n109 CSoutput.n93 9.25285
R7037 CSoutput.n347 CSoutput.n335 8.97993
R7038 CSoutput.n371 CSoutput.n359 8.97993
R7039 CSoutput.n348 CSoutput.n324 8.51219
R7040 CSoutput.n28 CSoutput.n15 8.25698
R7041 CSoutput.n65 CSoutput.n64 8.25698
R7042 CSoutput.n348 CSoutput.n347 7.89345
R7043 CSoutput.n372 CSoutput.n371 7.89345
R7044 CSoutput.n324 CSoutput.n323 7.12641
R7045 CSoutput.n126 CSoutput.n125 7.12641
R7046 CSoutput.n36 CSoutput.n35 6.91809
R7047 CSoutput.n57 CSoutput.n56 6.91809
R7048 CSoutput.n347 CSoutput.n346 5.25266
R7049 CSoutput.n371 CSoutput.n370 5.25266
R7050 CSoutput.n323 CSoutput.n322 5.1449
R7051 CSoutput.n307 CSoutput.n306 5.1449
R7052 CSoutput.n125 CSoutput.n124 5.1449
R7053 CSoutput.n109 CSoutput.n108 5.1449
R7054 CSoutput.n373 CSoutput.n126 4.91975
R7055 CSoutput.n217 CSoutput.n170 4.5005
R7056 CSoutput.n186 CSoutput.n170 4.5005
R7057 CSoutput.n181 CSoutput.n165 4.5005
R7058 CSoutput.n181 CSoutput.n167 4.5005
R7059 CSoutput.n181 CSoutput.n164 4.5005
R7060 CSoutput.n181 CSoutput.n168 4.5005
R7061 CSoutput.n181 CSoutput.n163 4.5005
R7062 CSoutput.n181 CSoutput.t152 4.5005
R7063 CSoutput.n181 CSoutput.n162 4.5005
R7064 CSoutput.n181 CSoutput.n169 4.5005
R7065 CSoutput.n181 CSoutput.n170 4.5005
R7066 CSoutput.n179 CSoutput.n165 4.5005
R7067 CSoutput.n179 CSoutput.n167 4.5005
R7068 CSoutput.n179 CSoutput.n164 4.5005
R7069 CSoutput.n179 CSoutput.n168 4.5005
R7070 CSoutput.n179 CSoutput.n163 4.5005
R7071 CSoutput.n179 CSoutput.t152 4.5005
R7072 CSoutput.n179 CSoutput.n162 4.5005
R7073 CSoutput.n179 CSoutput.n169 4.5005
R7074 CSoutput.n179 CSoutput.n170 4.5005
R7075 CSoutput.n178 CSoutput.n165 4.5005
R7076 CSoutput.n178 CSoutput.n167 4.5005
R7077 CSoutput.n178 CSoutput.n164 4.5005
R7078 CSoutput.n178 CSoutput.n168 4.5005
R7079 CSoutput.n178 CSoutput.n163 4.5005
R7080 CSoutput.n178 CSoutput.t152 4.5005
R7081 CSoutput.n178 CSoutput.n162 4.5005
R7082 CSoutput.n178 CSoutput.n169 4.5005
R7083 CSoutput.n178 CSoutput.n170 4.5005
R7084 CSoutput.n263 CSoutput.n165 4.5005
R7085 CSoutput.n263 CSoutput.n167 4.5005
R7086 CSoutput.n263 CSoutput.n164 4.5005
R7087 CSoutput.n263 CSoutput.n168 4.5005
R7088 CSoutput.n263 CSoutput.n163 4.5005
R7089 CSoutput.n263 CSoutput.t152 4.5005
R7090 CSoutput.n263 CSoutput.n162 4.5005
R7091 CSoutput.n263 CSoutput.n169 4.5005
R7092 CSoutput.n263 CSoutput.n170 4.5005
R7093 CSoutput.n261 CSoutput.n165 4.5005
R7094 CSoutput.n261 CSoutput.n167 4.5005
R7095 CSoutput.n261 CSoutput.n164 4.5005
R7096 CSoutput.n261 CSoutput.n168 4.5005
R7097 CSoutput.n261 CSoutput.n163 4.5005
R7098 CSoutput.n261 CSoutput.t152 4.5005
R7099 CSoutput.n261 CSoutput.n162 4.5005
R7100 CSoutput.n261 CSoutput.n169 4.5005
R7101 CSoutput.n259 CSoutput.n165 4.5005
R7102 CSoutput.n259 CSoutput.n167 4.5005
R7103 CSoutput.n259 CSoutput.n164 4.5005
R7104 CSoutput.n259 CSoutput.n168 4.5005
R7105 CSoutput.n259 CSoutput.n163 4.5005
R7106 CSoutput.n259 CSoutput.t152 4.5005
R7107 CSoutput.n259 CSoutput.n162 4.5005
R7108 CSoutput.n259 CSoutput.n169 4.5005
R7109 CSoutput.n189 CSoutput.n165 4.5005
R7110 CSoutput.n189 CSoutput.n167 4.5005
R7111 CSoutput.n189 CSoutput.n164 4.5005
R7112 CSoutput.n189 CSoutput.n168 4.5005
R7113 CSoutput.n189 CSoutput.n163 4.5005
R7114 CSoutput.n189 CSoutput.t152 4.5005
R7115 CSoutput.n189 CSoutput.n162 4.5005
R7116 CSoutput.n189 CSoutput.n169 4.5005
R7117 CSoutput.n189 CSoutput.n170 4.5005
R7118 CSoutput.n188 CSoutput.n165 4.5005
R7119 CSoutput.n188 CSoutput.n167 4.5005
R7120 CSoutput.n188 CSoutput.n164 4.5005
R7121 CSoutput.n188 CSoutput.n168 4.5005
R7122 CSoutput.n188 CSoutput.n163 4.5005
R7123 CSoutput.n188 CSoutput.t152 4.5005
R7124 CSoutput.n188 CSoutput.n162 4.5005
R7125 CSoutput.n188 CSoutput.n169 4.5005
R7126 CSoutput.n188 CSoutput.n170 4.5005
R7127 CSoutput.n192 CSoutput.n165 4.5005
R7128 CSoutput.n192 CSoutput.n167 4.5005
R7129 CSoutput.n192 CSoutput.n164 4.5005
R7130 CSoutput.n192 CSoutput.n168 4.5005
R7131 CSoutput.n192 CSoutput.n163 4.5005
R7132 CSoutput.n192 CSoutput.t152 4.5005
R7133 CSoutput.n192 CSoutput.n162 4.5005
R7134 CSoutput.n192 CSoutput.n169 4.5005
R7135 CSoutput.n192 CSoutput.n170 4.5005
R7136 CSoutput.n191 CSoutput.n165 4.5005
R7137 CSoutput.n191 CSoutput.n167 4.5005
R7138 CSoutput.n191 CSoutput.n164 4.5005
R7139 CSoutput.n191 CSoutput.n168 4.5005
R7140 CSoutput.n191 CSoutput.n163 4.5005
R7141 CSoutput.n191 CSoutput.t152 4.5005
R7142 CSoutput.n191 CSoutput.n162 4.5005
R7143 CSoutput.n191 CSoutput.n169 4.5005
R7144 CSoutput.n191 CSoutput.n170 4.5005
R7145 CSoutput.n174 CSoutput.n165 4.5005
R7146 CSoutput.n174 CSoutput.n167 4.5005
R7147 CSoutput.n174 CSoutput.n164 4.5005
R7148 CSoutput.n174 CSoutput.n168 4.5005
R7149 CSoutput.n174 CSoutput.n163 4.5005
R7150 CSoutput.n174 CSoutput.t152 4.5005
R7151 CSoutput.n174 CSoutput.n162 4.5005
R7152 CSoutput.n174 CSoutput.n169 4.5005
R7153 CSoutput.n174 CSoutput.n170 4.5005
R7154 CSoutput.n266 CSoutput.n165 4.5005
R7155 CSoutput.n266 CSoutput.n167 4.5005
R7156 CSoutput.n266 CSoutput.n164 4.5005
R7157 CSoutput.n266 CSoutput.n168 4.5005
R7158 CSoutput.n266 CSoutput.n163 4.5005
R7159 CSoutput.n266 CSoutput.t152 4.5005
R7160 CSoutput.n266 CSoutput.n162 4.5005
R7161 CSoutput.n266 CSoutput.n169 4.5005
R7162 CSoutput.n266 CSoutput.n170 4.5005
R7163 CSoutput.n253 CSoutput.n224 4.5005
R7164 CSoutput.n253 CSoutput.n230 4.5005
R7165 CSoutput.n211 CSoutput.n200 4.5005
R7166 CSoutput.n211 CSoutput.n202 4.5005
R7167 CSoutput.n211 CSoutput.n199 4.5005
R7168 CSoutput.n211 CSoutput.n203 4.5005
R7169 CSoutput.n211 CSoutput.n198 4.5005
R7170 CSoutput.n211 CSoutput.t146 4.5005
R7171 CSoutput.n211 CSoutput.n197 4.5005
R7172 CSoutput.n211 CSoutput.n204 4.5005
R7173 CSoutput.n253 CSoutput.n211 4.5005
R7174 CSoutput.n232 CSoutput.n200 4.5005
R7175 CSoutput.n232 CSoutput.n202 4.5005
R7176 CSoutput.n232 CSoutput.n199 4.5005
R7177 CSoutput.n232 CSoutput.n203 4.5005
R7178 CSoutput.n232 CSoutput.n198 4.5005
R7179 CSoutput.n232 CSoutput.t146 4.5005
R7180 CSoutput.n232 CSoutput.n197 4.5005
R7181 CSoutput.n232 CSoutput.n204 4.5005
R7182 CSoutput.n253 CSoutput.n232 4.5005
R7183 CSoutput.n210 CSoutput.n200 4.5005
R7184 CSoutput.n210 CSoutput.n202 4.5005
R7185 CSoutput.n210 CSoutput.n199 4.5005
R7186 CSoutput.n210 CSoutput.n203 4.5005
R7187 CSoutput.n210 CSoutput.n198 4.5005
R7188 CSoutput.n210 CSoutput.t146 4.5005
R7189 CSoutput.n210 CSoutput.n197 4.5005
R7190 CSoutput.n210 CSoutput.n204 4.5005
R7191 CSoutput.n253 CSoutput.n210 4.5005
R7192 CSoutput.n234 CSoutput.n200 4.5005
R7193 CSoutput.n234 CSoutput.n202 4.5005
R7194 CSoutput.n234 CSoutput.n199 4.5005
R7195 CSoutput.n234 CSoutput.n203 4.5005
R7196 CSoutput.n234 CSoutput.n198 4.5005
R7197 CSoutput.n234 CSoutput.t146 4.5005
R7198 CSoutput.n234 CSoutput.n197 4.5005
R7199 CSoutput.n234 CSoutput.n204 4.5005
R7200 CSoutput.n253 CSoutput.n234 4.5005
R7201 CSoutput.n200 CSoutput.n195 4.5005
R7202 CSoutput.n202 CSoutput.n195 4.5005
R7203 CSoutput.n199 CSoutput.n195 4.5005
R7204 CSoutput.n203 CSoutput.n195 4.5005
R7205 CSoutput.n198 CSoutput.n195 4.5005
R7206 CSoutput.t146 CSoutput.n195 4.5005
R7207 CSoutput.n197 CSoutput.n195 4.5005
R7208 CSoutput.n204 CSoutput.n195 4.5005
R7209 CSoutput.n256 CSoutput.n200 4.5005
R7210 CSoutput.n256 CSoutput.n202 4.5005
R7211 CSoutput.n256 CSoutput.n199 4.5005
R7212 CSoutput.n256 CSoutput.n203 4.5005
R7213 CSoutput.n256 CSoutput.n198 4.5005
R7214 CSoutput.n256 CSoutput.t146 4.5005
R7215 CSoutput.n256 CSoutput.n197 4.5005
R7216 CSoutput.n256 CSoutput.n204 4.5005
R7217 CSoutput.n254 CSoutput.n200 4.5005
R7218 CSoutput.n254 CSoutput.n202 4.5005
R7219 CSoutput.n254 CSoutput.n199 4.5005
R7220 CSoutput.n254 CSoutput.n203 4.5005
R7221 CSoutput.n254 CSoutput.n198 4.5005
R7222 CSoutput.n254 CSoutput.t146 4.5005
R7223 CSoutput.n254 CSoutput.n197 4.5005
R7224 CSoutput.n254 CSoutput.n204 4.5005
R7225 CSoutput.n254 CSoutput.n253 4.5005
R7226 CSoutput.n236 CSoutput.n200 4.5005
R7227 CSoutput.n236 CSoutput.n202 4.5005
R7228 CSoutput.n236 CSoutput.n199 4.5005
R7229 CSoutput.n236 CSoutput.n203 4.5005
R7230 CSoutput.n236 CSoutput.n198 4.5005
R7231 CSoutput.n236 CSoutput.t146 4.5005
R7232 CSoutput.n236 CSoutput.n197 4.5005
R7233 CSoutput.n236 CSoutput.n204 4.5005
R7234 CSoutput.n253 CSoutput.n236 4.5005
R7235 CSoutput.n208 CSoutput.n200 4.5005
R7236 CSoutput.n208 CSoutput.n202 4.5005
R7237 CSoutput.n208 CSoutput.n199 4.5005
R7238 CSoutput.n208 CSoutput.n203 4.5005
R7239 CSoutput.n208 CSoutput.n198 4.5005
R7240 CSoutput.n208 CSoutput.t146 4.5005
R7241 CSoutput.n208 CSoutput.n197 4.5005
R7242 CSoutput.n208 CSoutput.n204 4.5005
R7243 CSoutput.n253 CSoutput.n208 4.5005
R7244 CSoutput.n238 CSoutput.n200 4.5005
R7245 CSoutput.n238 CSoutput.n202 4.5005
R7246 CSoutput.n238 CSoutput.n199 4.5005
R7247 CSoutput.n238 CSoutput.n203 4.5005
R7248 CSoutput.n238 CSoutput.n198 4.5005
R7249 CSoutput.n238 CSoutput.t146 4.5005
R7250 CSoutput.n238 CSoutput.n197 4.5005
R7251 CSoutput.n238 CSoutput.n204 4.5005
R7252 CSoutput.n253 CSoutput.n238 4.5005
R7253 CSoutput.n207 CSoutput.n200 4.5005
R7254 CSoutput.n207 CSoutput.n202 4.5005
R7255 CSoutput.n207 CSoutput.n199 4.5005
R7256 CSoutput.n207 CSoutput.n203 4.5005
R7257 CSoutput.n207 CSoutput.n198 4.5005
R7258 CSoutput.n207 CSoutput.t146 4.5005
R7259 CSoutput.n207 CSoutput.n197 4.5005
R7260 CSoutput.n207 CSoutput.n204 4.5005
R7261 CSoutput.n253 CSoutput.n207 4.5005
R7262 CSoutput.n252 CSoutput.n200 4.5005
R7263 CSoutput.n252 CSoutput.n202 4.5005
R7264 CSoutput.n252 CSoutput.n199 4.5005
R7265 CSoutput.n252 CSoutput.n203 4.5005
R7266 CSoutput.n252 CSoutput.n198 4.5005
R7267 CSoutput.n252 CSoutput.t146 4.5005
R7268 CSoutput.n252 CSoutput.n197 4.5005
R7269 CSoutput.n252 CSoutput.n204 4.5005
R7270 CSoutput.n253 CSoutput.n252 4.5005
R7271 CSoutput.n251 CSoutput.n136 4.5005
R7272 CSoutput.n152 CSoutput.n136 4.5005
R7273 CSoutput.n147 CSoutput.n131 4.5005
R7274 CSoutput.n147 CSoutput.n133 4.5005
R7275 CSoutput.n147 CSoutput.n130 4.5005
R7276 CSoutput.n147 CSoutput.n134 4.5005
R7277 CSoutput.n147 CSoutput.n129 4.5005
R7278 CSoutput.n147 CSoutput.t164 4.5005
R7279 CSoutput.n147 CSoutput.n128 4.5005
R7280 CSoutput.n147 CSoutput.n135 4.5005
R7281 CSoutput.n147 CSoutput.n136 4.5005
R7282 CSoutput.n145 CSoutput.n131 4.5005
R7283 CSoutput.n145 CSoutput.n133 4.5005
R7284 CSoutput.n145 CSoutput.n130 4.5005
R7285 CSoutput.n145 CSoutput.n134 4.5005
R7286 CSoutput.n145 CSoutput.n129 4.5005
R7287 CSoutput.n145 CSoutput.t164 4.5005
R7288 CSoutput.n145 CSoutput.n128 4.5005
R7289 CSoutput.n145 CSoutput.n135 4.5005
R7290 CSoutput.n145 CSoutput.n136 4.5005
R7291 CSoutput.n144 CSoutput.n131 4.5005
R7292 CSoutput.n144 CSoutput.n133 4.5005
R7293 CSoutput.n144 CSoutput.n130 4.5005
R7294 CSoutput.n144 CSoutput.n134 4.5005
R7295 CSoutput.n144 CSoutput.n129 4.5005
R7296 CSoutput.n144 CSoutput.t164 4.5005
R7297 CSoutput.n144 CSoutput.n128 4.5005
R7298 CSoutput.n144 CSoutput.n135 4.5005
R7299 CSoutput.n144 CSoutput.n136 4.5005
R7300 CSoutput.n273 CSoutput.n131 4.5005
R7301 CSoutput.n273 CSoutput.n133 4.5005
R7302 CSoutput.n273 CSoutput.n130 4.5005
R7303 CSoutput.n273 CSoutput.n134 4.5005
R7304 CSoutput.n273 CSoutput.n129 4.5005
R7305 CSoutput.n273 CSoutput.t164 4.5005
R7306 CSoutput.n273 CSoutput.n128 4.5005
R7307 CSoutput.n273 CSoutput.n135 4.5005
R7308 CSoutput.n273 CSoutput.n136 4.5005
R7309 CSoutput.n271 CSoutput.n131 4.5005
R7310 CSoutput.n271 CSoutput.n133 4.5005
R7311 CSoutput.n271 CSoutput.n130 4.5005
R7312 CSoutput.n271 CSoutput.n134 4.5005
R7313 CSoutput.n271 CSoutput.n129 4.5005
R7314 CSoutput.n271 CSoutput.t164 4.5005
R7315 CSoutput.n271 CSoutput.n128 4.5005
R7316 CSoutput.n271 CSoutput.n135 4.5005
R7317 CSoutput.n269 CSoutput.n131 4.5005
R7318 CSoutput.n269 CSoutput.n133 4.5005
R7319 CSoutput.n269 CSoutput.n130 4.5005
R7320 CSoutput.n269 CSoutput.n134 4.5005
R7321 CSoutput.n269 CSoutput.n129 4.5005
R7322 CSoutput.n269 CSoutput.t164 4.5005
R7323 CSoutput.n269 CSoutput.n128 4.5005
R7324 CSoutput.n269 CSoutput.n135 4.5005
R7325 CSoutput.n155 CSoutput.n131 4.5005
R7326 CSoutput.n155 CSoutput.n133 4.5005
R7327 CSoutput.n155 CSoutput.n130 4.5005
R7328 CSoutput.n155 CSoutput.n134 4.5005
R7329 CSoutput.n155 CSoutput.n129 4.5005
R7330 CSoutput.n155 CSoutput.t164 4.5005
R7331 CSoutput.n155 CSoutput.n128 4.5005
R7332 CSoutput.n155 CSoutput.n135 4.5005
R7333 CSoutput.n155 CSoutput.n136 4.5005
R7334 CSoutput.n154 CSoutput.n131 4.5005
R7335 CSoutput.n154 CSoutput.n133 4.5005
R7336 CSoutput.n154 CSoutput.n130 4.5005
R7337 CSoutput.n154 CSoutput.n134 4.5005
R7338 CSoutput.n154 CSoutput.n129 4.5005
R7339 CSoutput.n154 CSoutput.t164 4.5005
R7340 CSoutput.n154 CSoutput.n128 4.5005
R7341 CSoutput.n154 CSoutput.n135 4.5005
R7342 CSoutput.n154 CSoutput.n136 4.5005
R7343 CSoutput.n158 CSoutput.n131 4.5005
R7344 CSoutput.n158 CSoutput.n133 4.5005
R7345 CSoutput.n158 CSoutput.n130 4.5005
R7346 CSoutput.n158 CSoutput.n134 4.5005
R7347 CSoutput.n158 CSoutput.n129 4.5005
R7348 CSoutput.n158 CSoutput.t164 4.5005
R7349 CSoutput.n158 CSoutput.n128 4.5005
R7350 CSoutput.n158 CSoutput.n135 4.5005
R7351 CSoutput.n158 CSoutput.n136 4.5005
R7352 CSoutput.n157 CSoutput.n131 4.5005
R7353 CSoutput.n157 CSoutput.n133 4.5005
R7354 CSoutput.n157 CSoutput.n130 4.5005
R7355 CSoutput.n157 CSoutput.n134 4.5005
R7356 CSoutput.n157 CSoutput.n129 4.5005
R7357 CSoutput.n157 CSoutput.t164 4.5005
R7358 CSoutput.n157 CSoutput.n128 4.5005
R7359 CSoutput.n157 CSoutput.n135 4.5005
R7360 CSoutput.n157 CSoutput.n136 4.5005
R7361 CSoutput.n140 CSoutput.n131 4.5005
R7362 CSoutput.n140 CSoutput.n133 4.5005
R7363 CSoutput.n140 CSoutput.n130 4.5005
R7364 CSoutput.n140 CSoutput.n134 4.5005
R7365 CSoutput.n140 CSoutput.n129 4.5005
R7366 CSoutput.n140 CSoutput.t164 4.5005
R7367 CSoutput.n140 CSoutput.n128 4.5005
R7368 CSoutput.n140 CSoutput.n135 4.5005
R7369 CSoutput.n140 CSoutput.n136 4.5005
R7370 CSoutput.n276 CSoutput.n131 4.5005
R7371 CSoutput.n276 CSoutput.n133 4.5005
R7372 CSoutput.n276 CSoutput.n130 4.5005
R7373 CSoutput.n276 CSoutput.n134 4.5005
R7374 CSoutput.n276 CSoutput.n129 4.5005
R7375 CSoutput.n276 CSoutput.t164 4.5005
R7376 CSoutput.n276 CSoutput.n128 4.5005
R7377 CSoutput.n276 CSoutput.n135 4.5005
R7378 CSoutput.n276 CSoutput.n136 4.5005
R7379 CSoutput.n323 CSoutput.n307 4.10845
R7380 CSoutput.n125 CSoutput.n109 4.10845
R7381 CSoutput.n321 CSoutput.t81 4.06363
R7382 CSoutput.n321 CSoutput.t14 4.06363
R7383 CSoutput.n319 CSoutput.t9 4.06363
R7384 CSoutput.n319 CSoutput.t50 4.06363
R7385 CSoutput.n317 CSoutput.t63 4.06363
R7386 CSoutput.n317 CSoutput.t83 4.06363
R7387 CSoutput.n315 CSoutput.t94 4.06363
R7388 CSoutput.n315 CSoutput.t25 4.06363
R7389 CSoutput.n313 CSoutput.t29 4.06363
R7390 CSoutput.n313 CSoutput.t84 4.06363
R7391 CSoutput.n311 CSoutput.t96 4.06363
R7392 CSoutput.n311 CSoutput.t97 4.06363
R7393 CSoutput.n309 CSoutput.t47 4.06363
R7394 CSoutput.n309 CSoutput.t48 4.06363
R7395 CSoutput.n308 CSoutput.t51 4.06363
R7396 CSoutput.n308 CSoutput.t99 4.06363
R7397 CSoutput.n305 CSoutput.t72 4.06363
R7398 CSoutput.n305 CSoutput.t98 4.06363
R7399 CSoutput.n303 CSoutput.t95 4.06363
R7400 CSoutput.n303 CSoutput.t37 4.06363
R7401 CSoutput.n301 CSoutput.t53 4.06363
R7402 CSoutput.n301 CSoutput.t73 4.06363
R7403 CSoutput.n299 CSoutput.t87 4.06363
R7404 CSoutput.n299 CSoutput.t13 4.06363
R7405 CSoutput.n297 CSoutput.t15 4.06363
R7406 CSoutput.n297 CSoutput.t76 4.06363
R7407 CSoutput.n295 CSoutput.t88 4.06363
R7408 CSoutput.n295 CSoutput.t89 4.06363
R7409 CSoutput.n293 CSoutput.t31 4.06363
R7410 CSoutput.n293 CSoutput.t34 4.06363
R7411 CSoutput.n292 CSoutput.t38 4.06363
R7412 CSoutput.n292 CSoutput.t90 4.06363
R7413 CSoutput.n290 CSoutput.t75 4.06363
R7414 CSoutput.n290 CSoutput.t35 4.06363
R7415 CSoutput.n288 CSoutput.t91 4.06363
R7416 CSoutput.n288 CSoutput.t58 4.06363
R7417 CSoutput.n286 CSoutput.t82 4.06363
R7418 CSoutput.n286 CSoutput.t43 4.06363
R7419 CSoutput.n284 CSoutput.t69 4.06363
R7420 CSoutput.n284 CSoutput.t24 4.06363
R7421 CSoutput.n282 CSoutput.t86 4.06363
R7422 CSoutput.n282 CSoutput.t20 4.06363
R7423 CSoutput.n280 CSoutput.t55 4.06363
R7424 CSoutput.n280 CSoutput.t33 4.06363
R7425 CSoutput.n278 CSoutput.t39 4.06363
R7426 CSoutput.n278 CSoutput.t17 4.06363
R7427 CSoutput.n277 CSoutput.t79 4.06363
R7428 CSoutput.n277 CSoutput.t10 4.06363
R7429 CSoutput.n110 CSoutput.t46 4.06363
R7430 CSoutput.n110 CSoutput.t101 4.06363
R7431 CSoutput.n111 CSoutput.t77 4.06363
R7432 CSoutput.n111 CSoutput.t78 4.06363
R7433 CSoutput.n113 CSoutput.t65 4.06363
R7434 CSoutput.n113 CSoutput.t44 4.06363
R7435 CSoutput.n115 CSoutput.t23 4.06363
R7436 CSoutput.n115 CSoutput.t66 4.06363
R7437 CSoutput.n117 CSoutput.t64 4.06363
R7438 CSoutput.n117 CSoutput.t40 4.06363
R7439 CSoutput.n119 CSoutput.t22 4.06363
R7440 CSoutput.n119 CSoutput.t21 4.06363
R7441 CSoutput.n121 CSoutput.t80 4.06363
R7442 CSoutput.n121 CSoutput.t52 4.06363
R7443 CSoutput.n123 CSoutput.t49 4.06363
R7444 CSoutput.n123 CSoutput.t18 4.06363
R7445 CSoutput.n94 CSoutput.t30 4.06363
R7446 CSoutput.n94 CSoutput.t93 4.06363
R7447 CSoutput.n95 CSoutput.t70 4.06363
R7448 CSoutput.n95 CSoutput.t67 4.06363
R7449 CSoutput.n97 CSoutput.t60 4.06363
R7450 CSoutput.n97 CSoutput.t28 4.06363
R7451 CSoutput.n99 CSoutput.t11 4.06363
R7452 CSoutput.n99 CSoutput.t59 4.06363
R7453 CSoutput.n101 CSoutput.t56 4.06363
R7454 CSoutput.n101 CSoutput.t27 4.06363
R7455 CSoutput.n103 CSoutput.t7 4.06363
R7456 CSoutput.n103 CSoutput.t8 4.06363
R7457 CSoutput.n105 CSoutput.t71 4.06363
R7458 CSoutput.n105 CSoutput.t42 4.06363
R7459 CSoutput.n107 CSoutput.t36 4.06363
R7460 CSoutput.n107 CSoutput.t6 4.06363
R7461 CSoutput.n79 CSoutput.t12 4.06363
R7462 CSoutput.n79 CSoutput.t61 4.06363
R7463 CSoutput.n80 CSoutput.t16 4.06363
R7464 CSoutput.n80 CSoutput.t41 4.06363
R7465 CSoutput.n82 CSoutput.t100 4.06363
R7466 CSoutput.n82 CSoutput.t54 4.06363
R7467 CSoutput.n84 CSoutput.t19 4.06363
R7468 CSoutput.n84 CSoutput.t85 4.06363
R7469 CSoutput.n86 CSoutput.t26 4.06363
R7470 CSoutput.n86 CSoutput.t68 4.06363
R7471 CSoutput.n88 CSoutput.t45 4.06363
R7472 CSoutput.n88 CSoutput.t62 4.06363
R7473 CSoutput.n90 CSoutput.t57 4.06363
R7474 CSoutput.n90 CSoutput.t92 4.06363
R7475 CSoutput.n92 CSoutput.t32 4.06363
R7476 CSoutput.n92 CSoutput.t74 4.06363
R7477 CSoutput.n44 CSoutput.n43 3.79402
R7478 CSoutput.n49 CSoutput.n48 3.79402
R7479 CSoutput.n373 CSoutput.n372 3.57343
R7480 CSoutput.n345 CSoutput.t104 2.82907
R7481 CSoutput.n345 CSoutput.t121 2.82907
R7482 CSoutput.n343 CSoutput.t140 2.82907
R7483 CSoutput.n343 CSoutput.t102 2.82907
R7484 CSoutput.n341 CSoutput.t112 2.82907
R7485 CSoutput.n341 CSoutput.t111 2.82907
R7486 CSoutput.n339 CSoutput.t108 2.82907
R7487 CSoutput.n339 CSoutput.t129 2.82907
R7488 CSoutput.n337 CSoutput.t139 2.82907
R7489 CSoutput.n337 CSoutput.t4 2.82907
R7490 CSoutput.n336 CSoutput.t106 2.82907
R7491 CSoutput.n336 CSoutput.t115 2.82907
R7492 CSoutput.n334 CSoutput.t127 2.82907
R7493 CSoutput.n334 CSoutput.t107 2.82907
R7494 CSoutput.n332 CSoutput.t122 2.82907
R7495 CSoutput.n332 CSoutput.t142 2.82907
R7496 CSoutput.n330 CSoutput.t120 2.82907
R7497 CSoutput.n330 CSoutput.t125 2.82907
R7498 CSoutput.n328 CSoutput.t143 2.82907
R7499 CSoutput.n328 CSoutput.t137 2.82907
R7500 CSoutput.n326 CSoutput.t0 2.82907
R7501 CSoutput.n326 CSoutput.t103 2.82907
R7502 CSoutput.n325 CSoutput.t114 2.82907
R7503 CSoutput.n325 CSoutput.t109 2.82907
R7504 CSoutput.n360 CSoutput.t138 2.82907
R7505 CSoutput.n360 CSoutput.t128 2.82907
R7506 CSoutput.n361 CSoutput.t119 2.82907
R7507 CSoutput.n361 CSoutput.t5 2.82907
R7508 CSoutput.n363 CSoutput.t135 2.82907
R7509 CSoutput.n363 CSoutput.t131 2.82907
R7510 CSoutput.n365 CSoutput.t141 2.82907
R7511 CSoutput.n365 CSoutput.t136 2.82907
R7512 CSoutput.n367 CSoutput.t116 2.82907
R7513 CSoutput.n367 CSoutput.t123 2.82907
R7514 CSoutput.n369 CSoutput.t113 2.82907
R7515 CSoutput.n369 CSoutput.t1 2.82907
R7516 CSoutput.n349 CSoutput.t133 2.82907
R7517 CSoutput.n349 CSoutput.t105 2.82907
R7518 CSoutput.n350 CSoutput.t117 2.82907
R7519 CSoutput.n350 CSoutput.t110 2.82907
R7520 CSoutput.n352 CSoutput.t118 2.82907
R7521 CSoutput.n352 CSoutput.t132 2.82907
R7522 CSoutput.n354 CSoutput.t2 2.82907
R7523 CSoutput.n354 CSoutput.t3 2.82907
R7524 CSoutput.n356 CSoutput.t134 2.82907
R7525 CSoutput.n356 CSoutput.t124 2.82907
R7526 CSoutput.n358 CSoutput.t130 2.82907
R7527 CSoutput.n358 CSoutput.t126 2.82907
R7528 CSoutput.n324 CSoutput.n126 2.78353
R7529 CSoutput.n372 CSoutput.n348 2.75627
R7530 CSoutput.n75 CSoutput.n1 2.45513
R7531 CSoutput.n217 CSoutput.n215 2.251
R7532 CSoutput.n217 CSoutput.n214 2.251
R7533 CSoutput.n217 CSoutput.n213 2.251
R7534 CSoutput.n217 CSoutput.n212 2.251
R7535 CSoutput.n186 CSoutput.n185 2.251
R7536 CSoutput.n186 CSoutput.n184 2.251
R7537 CSoutput.n186 CSoutput.n183 2.251
R7538 CSoutput.n186 CSoutput.n182 2.251
R7539 CSoutput.n259 CSoutput.n258 2.251
R7540 CSoutput.n224 CSoutput.n222 2.251
R7541 CSoutput.n224 CSoutput.n221 2.251
R7542 CSoutput.n224 CSoutput.n220 2.251
R7543 CSoutput.n242 CSoutput.n224 2.251
R7544 CSoutput.n230 CSoutput.n229 2.251
R7545 CSoutput.n230 CSoutput.n228 2.251
R7546 CSoutput.n230 CSoutput.n227 2.251
R7547 CSoutput.n230 CSoutput.n226 2.251
R7548 CSoutput.n256 CSoutput.n196 2.251
R7549 CSoutput.n251 CSoutput.n249 2.251
R7550 CSoutput.n251 CSoutput.n248 2.251
R7551 CSoutput.n251 CSoutput.n247 2.251
R7552 CSoutput.n251 CSoutput.n246 2.251
R7553 CSoutput.n152 CSoutput.n151 2.251
R7554 CSoutput.n152 CSoutput.n150 2.251
R7555 CSoutput.n152 CSoutput.n149 2.251
R7556 CSoutput.n152 CSoutput.n148 2.251
R7557 CSoutput.n269 CSoutput.n268 2.251
R7558 CSoutput.n186 CSoutput.n166 2.2505
R7559 CSoutput.n181 CSoutput.n166 2.2505
R7560 CSoutput.n179 CSoutput.n166 2.2505
R7561 CSoutput.n178 CSoutput.n166 2.2505
R7562 CSoutput.n263 CSoutput.n166 2.2505
R7563 CSoutput.n261 CSoutput.n166 2.2505
R7564 CSoutput.n259 CSoutput.n166 2.2505
R7565 CSoutput.n189 CSoutput.n166 2.2505
R7566 CSoutput.n188 CSoutput.n166 2.2505
R7567 CSoutput.n192 CSoutput.n166 2.2505
R7568 CSoutput.n191 CSoutput.n166 2.2505
R7569 CSoutput.n174 CSoutput.n166 2.2505
R7570 CSoutput.n266 CSoutput.n166 2.2505
R7571 CSoutput.n266 CSoutput.n265 2.2505
R7572 CSoutput.n230 CSoutput.n201 2.2505
R7573 CSoutput.n211 CSoutput.n201 2.2505
R7574 CSoutput.n232 CSoutput.n201 2.2505
R7575 CSoutput.n210 CSoutput.n201 2.2505
R7576 CSoutput.n234 CSoutput.n201 2.2505
R7577 CSoutput.n201 CSoutput.n195 2.2505
R7578 CSoutput.n256 CSoutput.n201 2.2505
R7579 CSoutput.n254 CSoutput.n201 2.2505
R7580 CSoutput.n236 CSoutput.n201 2.2505
R7581 CSoutput.n208 CSoutput.n201 2.2505
R7582 CSoutput.n238 CSoutput.n201 2.2505
R7583 CSoutput.n207 CSoutput.n201 2.2505
R7584 CSoutput.n252 CSoutput.n201 2.2505
R7585 CSoutput.n252 CSoutput.n205 2.2505
R7586 CSoutput.n152 CSoutput.n132 2.2505
R7587 CSoutput.n147 CSoutput.n132 2.2505
R7588 CSoutput.n145 CSoutput.n132 2.2505
R7589 CSoutput.n144 CSoutput.n132 2.2505
R7590 CSoutput.n273 CSoutput.n132 2.2505
R7591 CSoutput.n271 CSoutput.n132 2.2505
R7592 CSoutput.n269 CSoutput.n132 2.2505
R7593 CSoutput.n155 CSoutput.n132 2.2505
R7594 CSoutput.n154 CSoutput.n132 2.2505
R7595 CSoutput.n158 CSoutput.n132 2.2505
R7596 CSoutput.n157 CSoutput.n132 2.2505
R7597 CSoutput.n140 CSoutput.n132 2.2505
R7598 CSoutput.n276 CSoutput.n132 2.2505
R7599 CSoutput.n276 CSoutput.n275 2.2505
R7600 CSoutput.n194 CSoutput.n187 2.25024
R7601 CSoutput.n194 CSoutput.n180 2.25024
R7602 CSoutput.n262 CSoutput.n194 2.25024
R7603 CSoutput.n194 CSoutput.n190 2.25024
R7604 CSoutput.n194 CSoutput.n193 2.25024
R7605 CSoutput.n194 CSoutput.n161 2.25024
R7606 CSoutput.n244 CSoutput.n241 2.25024
R7607 CSoutput.n244 CSoutput.n240 2.25024
R7608 CSoutput.n244 CSoutput.n239 2.25024
R7609 CSoutput.n244 CSoutput.n206 2.25024
R7610 CSoutput.n244 CSoutput.n243 2.25024
R7611 CSoutput.n245 CSoutput.n244 2.25024
R7612 CSoutput.n160 CSoutput.n153 2.25024
R7613 CSoutput.n160 CSoutput.n146 2.25024
R7614 CSoutput.n272 CSoutput.n160 2.25024
R7615 CSoutput.n160 CSoutput.n156 2.25024
R7616 CSoutput.n160 CSoutput.n159 2.25024
R7617 CSoutput.n160 CSoutput.n127 2.25024
R7618 CSoutput.n261 CSoutput.n171 1.50111
R7619 CSoutput.n209 CSoutput.n195 1.50111
R7620 CSoutput.n271 CSoutput.n137 1.50111
R7621 CSoutput.n217 CSoutput.n216 1.501
R7622 CSoutput.n224 CSoutput.n223 1.501
R7623 CSoutput.n251 CSoutput.n250 1.501
R7624 CSoutput.n265 CSoutput.n176 1.12536
R7625 CSoutput.n265 CSoutput.n177 1.12536
R7626 CSoutput.n265 CSoutput.n264 1.12536
R7627 CSoutput.n225 CSoutput.n205 1.12536
R7628 CSoutput.n231 CSoutput.n205 1.12536
R7629 CSoutput.n233 CSoutput.n205 1.12536
R7630 CSoutput.n275 CSoutput.n142 1.12536
R7631 CSoutput.n275 CSoutput.n143 1.12536
R7632 CSoutput.n275 CSoutput.n274 1.12536
R7633 CSoutput.n265 CSoutput.n172 1.12536
R7634 CSoutput.n265 CSoutput.n173 1.12536
R7635 CSoutput.n265 CSoutput.n175 1.12536
R7636 CSoutput.n255 CSoutput.n205 1.12536
R7637 CSoutput.n235 CSoutput.n205 1.12536
R7638 CSoutput.n237 CSoutput.n205 1.12536
R7639 CSoutput.n275 CSoutput.n138 1.12536
R7640 CSoutput.n275 CSoutput.n139 1.12536
R7641 CSoutput.n275 CSoutput.n141 1.12536
R7642 CSoutput.n31 CSoutput.n30 0.669944
R7643 CSoutput.n62 CSoutput.n61 0.669944
R7644 CSoutput.n340 CSoutput.n338 0.573776
R7645 CSoutput.n342 CSoutput.n340 0.573776
R7646 CSoutput.n344 CSoutput.n342 0.573776
R7647 CSoutput.n346 CSoutput.n344 0.573776
R7648 CSoutput.n329 CSoutput.n327 0.573776
R7649 CSoutput.n331 CSoutput.n329 0.573776
R7650 CSoutput.n333 CSoutput.n331 0.573776
R7651 CSoutput.n335 CSoutput.n333 0.573776
R7652 CSoutput.n370 CSoutput.n368 0.573776
R7653 CSoutput.n368 CSoutput.n366 0.573776
R7654 CSoutput.n366 CSoutput.n364 0.573776
R7655 CSoutput.n364 CSoutput.n362 0.573776
R7656 CSoutput.n359 CSoutput.n357 0.573776
R7657 CSoutput.n357 CSoutput.n355 0.573776
R7658 CSoutput.n355 CSoutput.n353 0.573776
R7659 CSoutput.n353 CSoutput.n351 0.573776
R7660 CSoutput.n373 CSoutput.n276 0.53442
R7661 CSoutput.n312 CSoutput.n310 0.358259
R7662 CSoutput.n314 CSoutput.n312 0.358259
R7663 CSoutput.n316 CSoutput.n314 0.358259
R7664 CSoutput.n318 CSoutput.n316 0.358259
R7665 CSoutput.n320 CSoutput.n318 0.358259
R7666 CSoutput.n322 CSoutput.n320 0.358259
R7667 CSoutput.n296 CSoutput.n294 0.358259
R7668 CSoutput.n298 CSoutput.n296 0.358259
R7669 CSoutput.n300 CSoutput.n298 0.358259
R7670 CSoutput.n302 CSoutput.n300 0.358259
R7671 CSoutput.n304 CSoutput.n302 0.358259
R7672 CSoutput.n306 CSoutput.n304 0.358259
R7673 CSoutput.n281 CSoutput.n279 0.358259
R7674 CSoutput.n283 CSoutput.n281 0.358259
R7675 CSoutput.n285 CSoutput.n283 0.358259
R7676 CSoutput.n287 CSoutput.n285 0.358259
R7677 CSoutput.n289 CSoutput.n287 0.358259
R7678 CSoutput.n291 CSoutput.n289 0.358259
R7679 CSoutput.n124 CSoutput.n122 0.358259
R7680 CSoutput.n122 CSoutput.n120 0.358259
R7681 CSoutput.n120 CSoutput.n118 0.358259
R7682 CSoutput.n118 CSoutput.n116 0.358259
R7683 CSoutput.n116 CSoutput.n114 0.358259
R7684 CSoutput.n114 CSoutput.n112 0.358259
R7685 CSoutput.n108 CSoutput.n106 0.358259
R7686 CSoutput.n106 CSoutput.n104 0.358259
R7687 CSoutput.n104 CSoutput.n102 0.358259
R7688 CSoutput.n102 CSoutput.n100 0.358259
R7689 CSoutput.n100 CSoutput.n98 0.358259
R7690 CSoutput.n98 CSoutput.n96 0.358259
R7691 CSoutput.n93 CSoutput.n91 0.358259
R7692 CSoutput.n91 CSoutput.n89 0.358259
R7693 CSoutput.n89 CSoutput.n87 0.358259
R7694 CSoutput.n87 CSoutput.n85 0.358259
R7695 CSoutput.n85 CSoutput.n83 0.358259
R7696 CSoutput.n83 CSoutput.n81 0.358259
R7697 CSoutput.n21 CSoutput.n20 0.169105
R7698 CSoutput.n21 CSoutput.n16 0.169105
R7699 CSoutput.n26 CSoutput.n16 0.169105
R7700 CSoutput.n27 CSoutput.n26 0.169105
R7701 CSoutput.n27 CSoutput.n14 0.169105
R7702 CSoutput.n32 CSoutput.n14 0.169105
R7703 CSoutput.n33 CSoutput.n32 0.169105
R7704 CSoutput.n34 CSoutput.n33 0.169105
R7705 CSoutput.n34 CSoutput.n12 0.169105
R7706 CSoutput.n39 CSoutput.n12 0.169105
R7707 CSoutput.n40 CSoutput.n39 0.169105
R7708 CSoutput.n40 CSoutput.n10 0.169105
R7709 CSoutput.n45 CSoutput.n10 0.169105
R7710 CSoutput.n46 CSoutput.n45 0.169105
R7711 CSoutput.n47 CSoutput.n46 0.169105
R7712 CSoutput.n47 CSoutput.n8 0.169105
R7713 CSoutput.n52 CSoutput.n8 0.169105
R7714 CSoutput.n53 CSoutput.n52 0.169105
R7715 CSoutput.n53 CSoutput.n6 0.169105
R7716 CSoutput.n58 CSoutput.n6 0.169105
R7717 CSoutput.n59 CSoutput.n58 0.169105
R7718 CSoutput.n60 CSoutput.n59 0.169105
R7719 CSoutput.n60 CSoutput.n4 0.169105
R7720 CSoutput.n66 CSoutput.n4 0.169105
R7721 CSoutput.n67 CSoutput.n66 0.169105
R7722 CSoutput.n68 CSoutput.n67 0.169105
R7723 CSoutput.n68 CSoutput.n2 0.169105
R7724 CSoutput.n73 CSoutput.n2 0.169105
R7725 CSoutput.n74 CSoutput.n73 0.169105
R7726 CSoutput.n74 CSoutput.n0 0.169105
R7727 CSoutput.n78 CSoutput.n0 0.169105
R7728 CSoutput.n219 CSoutput.n218 0.0910737
R7729 CSoutput.n270 CSoutput.n267 0.0723685
R7730 CSoutput.n224 CSoutput.n219 0.0522944
R7731 CSoutput.n267 CSoutput.n266 0.0499135
R7732 CSoutput.n218 CSoutput.n217 0.0499135
R7733 CSoutput.n252 CSoutput.n251 0.0464294
R7734 CSoutput.n260 CSoutput.n257 0.0391444
R7735 CSoutput.n219 CSoutput.t154 0.023435
R7736 CSoutput.n267 CSoutput.t153 0.02262
R7737 CSoutput.n218 CSoutput.t157 0.02262
R7738 CSoutput CSoutput.n373 0.0052
R7739 CSoutput.n189 CSoutput.n172 0.00365111
R7740 CSoutput.n192 CSoutput.n173 0.00365111
R7741 CSoutput.n175 CSoutput.n174 0.00365111
R7742 CSoutput.n217 CSoutput.n176 0.00365111
R7743 CSoutput.n181 CSoutput.n177 0.00365111
R7744 CSoutput.n264 CSoutput.n178 0.00365111
R7745 CSoutput.n255 CSoutput.n254 0.00365111
R7746 CSoutput.n235 CSoutput.n208 0.00365111
R7747 CSoutput.n237 CSoutput.n207 0.00365111
R7748 CSoutput.n225 CSoutput.n224 0.00365111
R7749 CSoutput.n231 CSoutput.n211 0.00365111
R7750 CSoutput.n233 CSoutput.n210 0.00365111
R7751 CSoutput.n155 CSoutput.n138 0.00365111
R7752 CSoutput.n158 CSoutput.n139 0.00365111
R7753 CSoutput.n141 CSoutput.n140 0.00365111
R7754 CSoutput.n251 CSoutput.n142 0.00365111
R7755 CSoutput.n147 CSoutput.n143 0.00365111
R7756 CSoutput.n274 CSoutput.n144 0.00365111
R7757 CSoutput.n186 CSoutput.n176 0.00340054
R7758 CSoutput.n179 CSoutput.n177 0.00340054
R7759 CSoutput.n264 CSoutput.n263 0.00340054
R7760 CSoutput.n259 CSoutput.n172 0.00340054
R7761 CSoutput.n188 CSoutput.n173 0.00340054
R7762 CSoutput.n191 CSoutput.n175 0.00340054
R7763 CSoutput.n230 CSoutput.n225 0.00340054
R7764 CSoutput.n232 CSoutput.n231 0.00340054
R7765 CSoutput.n234 CSoutput.n233 0.00340054
R7766 CSoutput.n256 CSoutput.n255 0.00340054
R7767 CSoutput.n236 CSoutput.n235 0.00340054
R7768 CSoutput.n238 CSoutput.n237 0.00340054
R7769 CSoutput.n152 CSoutput.n142 0.00340054
R7770 CSoutput.n145 CSoutput.n143 0.00340054
R7771 CSoutput.n274 CSoutput.n273 0.00340054
R7772 CSoutput.n269 CSoutput.n138 0.00340054
R7773 CSoutput.n154 CSoutput.n139 0.00340054
R7774 CSoutput.n157 CSoutput.n141 0.00340054
R7775 CSoutput.n187 CSoutput.n181 0.00252698
R7776 CSoutput.n180 CSoutput.n178 0.00252698
R7777 CSoutput.n262 CSoutput.n261 0.00252698
R7778 CSoutput.n190 CSoutput.n188 0.00252698
R7779 CSoutput.n193 CSoutput.n191 0.00252698
R7780 CSoutput.n266 CSoutput.n161 0.00252698
R7781 CSoutput.n187 CSoutput.n186 0.00252698
R7782 CSoutput.n180 CSoutput.n179 0.00252698
R7783 CSoutput.n263 CSoutput.n262 0.00252698
R7784 CSoutput.n190 CSoutput.n189 0.00252698
R7785 CSoutput.n193 CSoutput.n192 0.00252698
R7786 CSoutput.n174 CSoutput.n161 0.00252698
R7787 CSoutput.n241 CSoutput.n211 0.00252698
R7788 CSoutput.n240 CSoutput.n210 0.00252698
R7789 CSoutput.n239 CSoutput.n195 0.00252698
R7790 CSoutput.n236 CSoutput.n206 0.00252698
R7791 CSoutput.n243 CSoutput.n238 0.00252698
R7792 CSoutput.n252 CSoutput.n245 0.00252698
R7793 CSoutput.n241 CSoutput.n230 0.00252698
R7794 CSoutput.n240 CSoutput.n232 0.00252698
R7795 CSoutput.n239 CSoutput.n234 0.00252698
R7796 CSoutput.n254 CSoutput.n206 0.00252698
R7797 CSoutput.n243 CSoutput.n208 0.00252698
R7798 CSoutput.n245 CSoutput.n207 0.00252698
R7799 CSoutput.n153 CSoutput.n147 0.00252698
R7800 CSoutput.n146 CSoutput.n144 0.00252698
R7801 CSoutput.n272 CSoutput.n271 0.00252698
R7802 CSoutput.n156 CSoutput.n154 0.00252698
R7803 CSoutput.n159 CSoutput.n157 0.00252698
R7804 CSoutput.n276 CSoutput.n127 0.00252698
R7805 CSoutput.n153 CSoutput.n152 0.00252698
R7806 CSoutput.n146 CSoutput.n145 0.00252698
R7807 CSoutput.n273 CSoutput.n272 0.00252698
R7808 CSoutput.n156 CSoutput.n155 0.00252698
R7809 CSoutput.n159 CSoutput.n158 0.00252698
R7810 CSoutput.n140 CSoutput.n127 0.00252698
R7811 CSoutput.n261 CSoutput.n260 0.0020275
R7812 CSoutput.n260 CSoutput.n259 0.0020275
R7813 CSoutput.n257 CSoutput.n195 0.0020275
R7814 CSoutput.n257 CSoutput.n256 0.0020275
R7815 CSoutput.n271 CSoutput.n270 0.0020275
R7816 CSoutput.n270 CSoutput.n269 0.0020275
R7817 CSoutput.n171 CSoutput.n170 0.00166668
R7818 CSoutput.n253 CSoutput.n209 0.00166668
R7819 CSoutput.n137 CSoutput.n136 0.00166668
R7820 CSoutput.n275 CSoutput.n137 0.00133328
R7821 CSoutput.n209 CSoutput.n205 0.00133328
R7822 CSoutput.n265 CSoutput.n171 0.00133328
R7823 CSoutput.n268 CSoutput.n160 0.001
R7824 CSoutput.n246 CSoutput.n160 0.001
R7825 CSoutput.n148 CSoutput.n128 0.001
R7826 CSoutput.n247 CSoutput.n128 0.001
R7827 CSoutput.n149 CSoutput.n129 0.001
R7828 CSoutput.n248 CSoutput.n129 0.001
R7829 CSoutput.n150 CSoutput.n130 0.001
R7830 CSoutput.n249 CSoutput.n130 0.001
R7831 CSoutput.n151 CSoutput.n131 0.001
R7832 CSoutput.n250 CSoutput.n131 0.001
R7833 CSoutput.n244 CSoutput.n196 0.001
R7834 CSoutput.n244 CSoutput.n242 0.001
R7835 CSoutput.n226 CSoutput.n197 0.001
R7836 CSoutput.n220 CSoutput.n197 0.001
R7837 CSoutput.n227 CSoutput.n198 0.001
R7838 CSoutput.n221 CSoutput.n198 0.001
R7839 CSoutput.n228 CSoutput.n199 0.001
R7840 CSoutput.n222 CSoutput.n199 0.001
R7841 CSoutput.n229 CSoutput.n200 0.001
R7842 CSoutput.n223 CSoutput.n200 0.001
R7843 CSoutput.n258 CSoutput.n194 0.001
R7844 CSoutput.n212 CSoutput.n194 0.001
R7845 CSoutput.n182 CSoutput.n162 0.001
R7846 CSoutput.n213 CSoutput.n162 0.001
R7847 CSoutput.n183 CSoutput.n163 0.001
R7848 CSoutput.n214 CSoutput.n163 0.001
R7849 CSoutput.n184 CSoutput.n164 0.001
R7850 CSoutput.n215 CSoutput.n164 0.001
R7851 CSoutput.n185 CSoutput.n165 0.001
R7852 CSoutput.n216 CSoutput.n165 0.001
R7853 CSoutput.n216 CSoutput.n166 0.001
R7854 CSoutput.n215 CSoutput.n167 0.001
R7855 CSoutput.n214 CSoutput.n168 0.001
R7856 CSoutput.n213 CSoutput.t152 0.001
R7857 CSoutput.n212 CSoutput.n169 0.001
R7858 CSoutput.n185 CSoutput.n167 0.001
R7859 CSoutput.n184 CSoutput.n168 0.001
R7860 CSoutput.n183 CSoutput.t152 0.001
R7861 CSoutput.n182 CSoutput.n169 0.001
R7862 CSoutput.n258 CSoutput.n170 0.001
R7863 CSoutput.n223 CSoutput.n201 0.001
R7864 CSoutput.n222 CSoutput.n202 0.001
R7865 CSoutput.n221 CSoutput.n203 0.001
R7866 CSoutput.n220 CSoutput.t146 0.001
R7867 CSoutput.n242 CSoutput.n204 0.001
R7868 CSoutput.n229 CSoutput.n202 0.001
R7869 CSoutput.n228 CSoutput.n203 0.001
R7870 CSoutput.n227 CSoutput.t146 0.001
R7871 CSoutput.n226 CSoutput.n204 0.001
R7872 CSoutput.n253 CSoutput.n196 0.001
R7873 CSoutput.n250 CSoutput.n132 0.001
R7874 CSoutput.n249 CSoutput.n133 0.001
R7875 CSoutput.n248 CSoutput.n134 0.001
R7876 CSoutput.n247 CSoutput.t164 0.001
R7877 CSoutput.n246 CSoutput.n135 0.001
R7878 CSoutput.n151 CSoutput.n133 0.001
R7879 CSoutput.n150 CSoutput.n134 0.001
R7880 CSoutput.n149 CSoutput.t164 0.001
R7881 CSoutput.n148 CSoutput.n135 0.001
R7882 CSoutput.n268 CSoutput.n136 0.001
R7883 gnd.n6687 gnd.n6686 1758.55
R7884 gnd.n2317 gnd.n2316 931.112
R7885 gnd.n7045 gnd.n84 838.452
R7886 gnd.n7194 gnd.n80 838.452
R7887 gnd.n2936 gnd.n2669 838.452
R7888 gnd.n2857 gnd.n2671 838.452
R7889 gnd.n5925 gnd.n2538 838.452
R7890 gnd.n3842 gnd.n2536 838.452
R7891 gnd.n4048 gnd.n2320 838.452
R7892 gnd.n4005 gnd.n2322 838.452
R7893 gnd.n7192 gnd.n86 819.232
R7894 gnd.n155 gnd.n82 819.232
R7895 gnd.n3103 gnd.n2668 819.232
R7896 gnd.n5778 gnd.n2672 819.232
R7897 gnd.n5927 gnd.n2533 819.232
R7898 gnd.n4548 gnd.n2535 819.232
R7899 gnd.n4194 gnd.n2319 819.232
R7900 gnd.n6054 gnd.n2323 819.232
R7901 gnd.n3888 gnd.n2543 771.183
R7902 gnd.n5796 gnd.n2646 771.183
R7903 gnd.n3771 gnd.n3738 771.183
R7904 gnd.n5542 gnd.n2648 771.183
R7905 gnd.n2224 gnd.n868 766.379
R7906 gnd.n2227 gnd.n2226 766.379
R7907 gnd.n1464 gnd.n1367 766.379
R7908 gnd.n1460 gnd.n1365 766.379
R7909 gnd.n2315 gnd.n890 756.769
R7910 gnd.n2218 gnd.n2217 756.769
R7911 gnd.n1557 gnd.n1274 756.769
R7912 gnd.n1555 gnd.n1277 756.769
R7913 gnd.n6233 gnd.n696 670.282
R7914 gnd.n6688 gnd.n424 670.282
R7915 gnd.n6902 gnd.n6901 670.282
R7916 gnd.n6057 gnd.n861 670.282
R7917 gnd.n6229 gnd.n696 585
R7918 gnd.n696 gnd.n695 585
R7919 gnd.n6228 gnd.n6227 585
R7920 gnd.n6227 gnd.n6226 585
R7921 gnd.n699 gnd.n698 585
R7922 gnd.n6225 gnd.n699 585
R7923 gnd.n6223 gnd.n6222 585
R7924 gnd.n6224 gnd.n6223 585
R7925 gnd.n6221 gnd.n701 585
R7926 gnd.n701 gnd.n700 585
R7927 gnd.n6220 gnd.n6219 585
R7928 gnd.n6219 gnd.n6218 585
R7929 gnd.n707 gnd.n706 585
R7930 gnd.n6217 gnd.n707 585
R7931 gnd.n6215 gnd.n6214 585
R7932 gnd.n6216 gnd.n6215 585
R7933 gnd.n6213 gnd.n709 585
R7934 gnd.n709 gnd.n708 585
R7935 gnd.n6212 gnd.n6211 585
R7936 gnd.n6211 gnd.n6210 585
R7937 gnd.n715 gnd.n714 585
R7938 gnd.n6209 gnd.n715 585
R7939 gnd.n6207 gnd.n6206 585
R7940 gnd.n6208 gnd.n6207 585
R7941 gnd.n6205 gnd.n717 585
R7942 gnd.n717 gnd.n716 585
R7943 gnd.n6204 gnd.n6203 585
R7944 gnd.n6203 gnd.n6202 585
R7945 gnd.n723 gnd.n722 585
R7946 gnd.n6201 gnd.n723 585
R7947 gnd.n6199 gnd.n6198 585
R7948 gnd.n6200 gnd.n6199 585
R7949 gnd.n6197 gnd.n725 585
R7950 gnd.n725 gnd.n724 585
R7951 gnd.n6196 gnd.n6195 585
R7952 gnd.n6195 gnd.n6194 585
R7953 gnd.n731 gnd.n730 585
R7954 gnd.n6193 gnd.n731 585
R7955 gnd.n6191 gnd.n6190 585
R7956 gnd.n6192 gnd.n6191 585
R7957 gnd.n6189 gnd.n733 585
R7958 gnd.n733 gnd.n732 585
R7959 gnd.n6188 gnd.n6187 585
R7960 gnd.n6187 gnd.n6186 585
R7961 gnd.n739 gnd.n738 585
R7962 gnd.n6185 gnd.n739 585
R7963 gnd.n6183 gnd.n6182 585
R7964 gnd.n6184 gnd.n6183 585
R7965 gnd.n6181 gnd.n741 585
R7966 gnd.n741 gnd.n740 585
R7967 gnd.n6180 gnd.n6179 585
R7968 gnd.n6179 gnd.n6178 585
R7969 gnd.n747 gnd.n746 585
R7970 gnd.n6177 gnd.n747 585
R7971 gnd.n6175 gnd.n6174 585
R7972 gnd.n6176 gnd.n6175 585
R7973 gnd.n6173 gnd.n749 585
R7974 gnd.n749 gnd.n748 585
R7975 gnd.n6172 gnd.n6171 585
R7976 gnd.n6171 gnd.n6170 585
R7977 gnd.n755 gnd.n754 585
R7978 gnd.n6169 gnd.n755 585
R7979 gnd.n6167 gnd.n6166 585
R7980 gnd.n6168 gnd.n6167 585
R7981 gnd.n6165 gnd.n757 585
R7982 gnd.n757 gnd.n756 585
R7983 gnd.n6164 gnd.n6163 585
R7984 gnd.n6163 gnd.n6162 585
R7985 gnd.n763 gnd.n762 585
R7986 gnd.n6161 gnd.n763 585
R7987 gnd.n6159 gnd.n6158 585
R7988 gnd.n6160 gnd.n6159 585
R7989 gnd.n6157 gnd.n765 585
R7990 gnd.n765 gnd.n764 585
R7991 gnd.n6156 gnd.n6155 585
R7992 gnd.n6155 gnd.n6154 585
R7993 gnd.n771 gnd.n770 585
R7994 gnd.n6153 gnd.n771 585
R7995 gnd.n6151 gnd.n6150 585
R7996 gnd.n6152 gnd.n6151 585
R7997 gnd.n6149 gnd.n773 585
R7998 gnd.n773 gnd.n772 585
R7999 gnd.n6148 gnd.n6147 585
R8000 gnd.n6147 gnd.n6146 585
R8001 gnd.n779 gnd.n778 585
R8002 gnd.n6145 gnd.n779 585
R8003 gnd.n6143 gnd.n6142 585
R8004 gnd.n6144 gnd.n6143 585
R8005 gnd.n6141 gnd.n781 585
R8006 gnd.n781 gnd.n780 585
R8007 gnd.n6140 gnd.n6139 585
R8008 gnd.n6139 gnd.n6138 585
R8009 gnd.n787 gnd.n786 585
R8010 gnd.n6137 gnd.n787 585
R8011 gnd.n6135 gnd.n6134 585
R8012 gnd.n6136 gnd.n6135 585
R8013 gnd.n6133 gnd.n789 585
R8014 gnd.n789 gnd.n788 585
R8015 gnd.n6132 gnd.n6131 585
R8016 gnd.n6131 gnd.n6130 585
R8017 gnd.n795 gnd.n794 585
R8018 gnd.n6129 gnd.n795 585
R8019 gnd.n6127 gnd.n6126 585
R8020 gnd.n6128 gnd.n6127 585
R8021 gnd.n6125 gnd.n797 585
R8022 gnd.n797 gnd.n796 585
R8023 gnd.n6124 gnd.n6123 585
R8024 gnd.n6123 gnd.n6122 585
R8025 gnd.n803 gnd.n802 585
R8026 gnd.n6121 gnd.n803 585
R8027 gnd.n6119 gnd.n6118 585
R8028 gnd.n6120 gnd.n6119 585
R8029 gnd.n6117 gnd.n805 585
R8030 gnd.n805 gnd.n804 585
R8031 gnd.n6116 gnd.n6115 585
R8032 gnd.n6115 gnd.n6114 585
R8033 gnd.n811 gnd.n810 585
R8034 gnd.n6113 gnd.n811 585
R8035 gnd.n6111 gnd.n6110 585
R8036 gnd.n6112 gnd.n6111 585
R8037 gnd.n6109 gnd.n813 585
R8038 gnd.n813 gnd.n812 585
R8039 gnd.n6108 gnd.n6107 585
R8040 gnd.n6107 gnd.n6106 585
R8041 gnd.n819 gnd.n818 585
R8042 gnd.n6105 gnd.n819 585
R8043 gnd.n6103 gnd.n6102 585
R8044 gnd.n6104 gnd.n6103 585
R8045 gnd.n6101 gnd.n821 585
R8046 gnd.n821 gnd.n820 585
R8047 gnd.n6100 gnd.n6099 585
R8048 gnd.n6099 gnd.n6098 585
R8049 gnd.n827 gnd.n826 585
R8050 gnd.n6097 gnd.n827 585
R8051 gnd.n6095 gnd.n6094 585
R8052 gnd.n6096 gnd.n6095 585
R8053 gnd.n6093 gnd.n829 585
R8054 gnd.n829 gnd.n828 585
R8055 gnd.n6092 gnd.n6091 585
R8056 gnd.n6091 gnd.n6090 585
R8057 gnd.n835 gnd.n834 585
R8058 gnd.n6089 gnd.n835 585
R8059 gnd.n6087 gnd.n6086 585
R8060 gnd.n6088 gnd.n6087 585
R8061 gnd.n6085 gnd.n837 585
R8062 gnd.n837 gnd.n836 585
R8063 gnd.n6084 gnd.n6083 585
R8064 gnd.n6083 gnd.n6082 585
R8065 gnd.n843 gnd.n842 585
R8066 gnd.n6081 gnd.n843 585
R8067 gnd.n6079 gnd.n6078 585
R8068 gnd.n6080 gnd.n6079 585
R8069 gnd.n6077 gnd.n845 585
R8070 gnd.n845 gnd.n844 585
R8071 gnd.n6076 gnd.n6075 585
R8072 gnd.n6075 gnd.n6074 585
R8073 gnd.n851 gnd.n850 585
R8074 gnd.n6073 gnd.n851 585
R8075 gnd.n6071 gnd.n6070 585
R8076 gnd.n6072 gnd.n6071 585
R8077 gnd.n6069 gnd.n853 585
R8078 gnd.n853 gnd.n852 585
R8079 gnd.n6068 gnd.n6067 585
R8080 gnd.n6067 gnd.n6066 585
R8081 gnd.n859 gnd.n858 585
R8082 gnd.n6065 gnd.n859 585
R8083 gnd.n6063 gnd.n6062 585
R8084 gnd.n6064 gnd.n6063 585
R8085 gnd.n6233 gnd.n6232 585
R8086 gnd.n6234 gnd.n6233 585
R8087 gnd.n694 gnd.n693 585
R8088 gnd.n6235 gnd.n694 585
R8089 gnd.n6238 gnd.n6237 585
R8090 gnd.n6237 gnd.n6236 585
R8091 gnd.n691 gnd.n690 585
R8092 gnd.n690 gnd.n689 585
R8093 gnd.n6243 gnd.n6242 585
R8094 gnd.n6244 gnd.n6243 585
R8095 gnd.n688 gnd.n687 585
R8096 gnd.n6245 gnd.n688 585
R8097 gnd.n6248 gnd.n6247 585
R8098 gnd.n6247 gnd.n6246 585
R8099 gnd.n685 gnd.n684 585
R8100 gnd.n684 gnd.n683 585
R8101 gnd.n6253 gnd.n6252 585
R8102 gnd.n6254 gnd.n6253 585
R8103 gnd.n682 gnd.n681 585
R8104 gnd.n6255 gnd.n682 585
R8105 gnd.n6258 gnd.n6257 585
R8106 gnd.n6257 gnd.n6256 585
R8107 gnd.n679 gnd.n678 585
R8108 gnd.n678 gnd.n677 585
R8109 gnd.n6263 gnd.n6262 585
R8110 gnd.n6264 gnd.n6263 585
R8111 gnd.n676 gnd.n675 585
R8112 gnd.n6265 gnd.n676 585
R8113 gnd.n6268 gnd.n6267 585
R8114 gnd.n6267 gnd.n6266 585
R8115 gnd.n673 gnd.n672 585
R8116 gnd.n672 gnd.n671 585
R8117 gnd.n6273 gnd.n6272 585
R8118 gnd.n6274 gnd.n6273 585
R8119 gnd.n670 gnd.n669 585
R8120 gnd.n6275 gnd.n670 585
R8121 gnd.n6278 gnd.n6277 585
R8122 gnd.n6277 gnd.n6276 585
R8123 gnd.n667 gnd.n666 585
R8124 gnd.n666 gnd.n665 585
R8125 gnd.n6283 gnd.n6282 585
R8126 gnd.n6284 gnd.n6283 585
R8127 gnd.n664 gnd.n663 585
R8128 gnd.n6285 gnd.n664 585
R8129 gnd.n6288 gnd.n6287 585
R8130 gnd.n6287 gnd.n6286 585
R8131 gnd.n661 gnd.n660 585
R8132 gnd.n660 gnd.n659 585
R8133 gnd.n6293 gnd.n6292 585
R8134 gnd.n6294 gnd.n6293 585
R8135 gnd.n658 gnd.n657 585
R8136 gnd.n6295 gnd.n658 585
R8137 gnd.n6298 gnd.n6297 585
R8138 gnd.n6297 gnd.n6296 585
R8139 gnd.n655 gnd.n654 585
R8140 gnd.n654 gnd.n653 585
R8141 gnd.n6303 gnd.n6302 585
R8142 gnd.n6304 gnd.n6303 585
R8143 gnd.n652 gnd.n651 585
R8144 gnd.n6305 gnd.n652 585
R8145 gnd.n6308 gnd.n6307 585
R8146 gnd.n6307 gnd.n6306 585
R8147 gnd.n649 gnd.n648 585
R8148 gnd.n648 gnd.n647 585
R8149 gnd.n6313 gnd.n6312 585
R8150 gnd.n6314 gnd.n6313 585
R8151 gnd.n646 gnd.n645 585
R8152 gnd.n6315 gnd.n646 585
R8153 gnd.n6318 gnd.n6317 585
R8154 gnd.n6317 gnd.n6316 585
R8155 gnd.n643 gnd.n642 585
R8156 gnd.n642 gnd.n641 585
R8157 gnd.n6323 gnd.n6322 585
R8158 gnd.n6324 gnd.n6323 585
R8159 gnd.n640 gnd.n639 585
R8160 gnd.n6325 gnd.n640 585
R8161 gnd.n6328 gnd.n6327 585
R8162 gnd.n6327 gnd.n6326 585
R8163 gnd.n637 gnd.n636 585
R8164 gnd.n636 gnd.n635 585
R8165 gnd.n6333 gnd.n6332 585
R8166 gnd.n6334 gnd.n6333 585
R8167 gnd.n634 gnd.n633 585
R8168 gnd.n6335 gnd.n634 585
R8169 gnd.n6338 gnd.n6337 585
R8170 gnd.n6337 gnd.n6336 585
R8171 gnd.n631 gnd.n630 585
R8172 gnd.n630 gnd.n629 585
R8173 gnd.n6343 gnd.n6342 585
R8174 gnd.n6344 gnd.n6343 585
R8175 gnd.n628 gnd.n627 585
R8176 gnd.n6345 gnd.n628 585
R8177 gnd.n6348 gnd.n6347 585
R8178 gnd.n6347 gnd.n6346 585
R8179 gnd.n625 gnd.n624 585
R8180 gnd.n624 gnd.n623 585
R8181 gnd.n6353 gnd.n6352 585
R8182 gnd.n6354 gnd.n6353 585
R8183 gnd.n622 gnd.n621 585
R8184 gnd.n6355 gnd.n622 585
R8185 gnd.n6358 gnd.n6357 585
R8186 gnd.n6357 gnd.n6356 585
R8187 gnd.n619 gnd.n618 585
R8188 gnd.n618 gnd.n617 585
R8189 gnd.n6363 gnd.n6362 585
R8190 gnd.n6364 gnd.n6363 585
R8191 gnd.n616 gnd.n615 585
R8192 gnd.n6365 gnd.n616 585
R8193 gnd.n6368 gnd.n6367 585
R8194 gnd.n6367 gnd.n6366 585
R8195 gnd.n613 gnd.n612 585
R8196 gnd.n612 gnd.n611 585
R8197 gnd.n6373 gnd.n6372 585
R8198 gnd.n6374 gnd.n6373 585
R8199 gnd.n610 gnd.n609 585
R8200 gnd.n6375 gnd.n610 585
R8201 gnd.n6378 gnd.n6377 585
R8202 gnd.n6377 gnd.n6376 585
R8203 gnd.n607 gnd.n606 585
R8204 gnd.n606 gnd.n605 585
R8205 gnd.n6383 gnd.n6382 585
R8206 gnd.n6384 gnd.n6383 585
R8207 gnd.n604 gnd.n603 585
R8208 gnd.n6385 gnd.n604 585
R8209 gnd.n6388 gnd.n6387 585
R8210 gnd.n6387 gnd.n6386 585
R8211 gnd.n601 gnd.n600 585
R8212 gnd.n600 gnd.n599 585
R8213 gnd.n6393 gnd.n6392 585
R8214 gnd.n6394 gnd.n6393 585
R8215 gnd.n598 gnd.n597 585
R8216 gnd.n6395 gnd.n598 585
R8217 gnd.n6398 gnd.n6397 585
R8218 gnd.n6397 gnd.n6396 585
R8219 gnd.n595 gnd.n594 585
R8220 gnd.n594 gnd.n593 585
R8221 gnd.n6403 gnd.n6402 585
R8222 gnd.n6404 gnd.n6403 585
R8223 gnd.n592 gnd.n591 585
R8224 gnd.n6405 gnd.n592 585
R8225 gnd.n6408 gnd.n6407 585
R8226 gnd.n6407 gnd.n6406 585
R8227 gnd.n589 gnd.n588 585
R8228 gnd.n588 gnd.n587 585
R8229 gnd.n6413 gnd.n6412 585
R8230 gnd.n6414 gnd.n6413 585
R8231 gnd.n586 gnd.n585 585
R8232 gnd.n6415 gnd.n586 585
R8233 gnd.n6418 gnd.n6417 585
R8234 gnd.n6417 gnd.n6416 585
R8235 gnd.n583 gnd.n582 585
R8236 gnd.n582 gnd.n581 585
R8237 gnd.n6423 gnd.n6422 585
R8238 gnd.n6424 gnd.n6423 585
R8239 gnd.n580 gnd.n579 585
R8240 gnd.n6425 gnd.n580 585
R8241 gnd.n6428 gnd.n6427 585
R8242 gnd.n6427 gnd.n6426 585
R8243 gnd.n577 gnd.n576 585
R8244 gnd.n576 gnd.n575 585
R8245 gnd.n6433 gnd.n6432 585
R8246 gnd.n6434 gnd.n6433 585
R8247 gnd.n574 gnd.n573 585
R8248 gnd.n6435 gnd.n574 585
R8249 gnd.n6438 gnd.n6437 585
R8250 gnd.n6437 gnd.n6436 585
R8251 gnd.n571 gnd.n570 585
R8252 gnd.n570 gnd.n569 585
R8253 gnd.n6443 gnd.n6442 585
R8254 gnd.n6444 gnd.n6443 585
R8255 gnd.n568 gnd.n567 585
R8256 gnd.n6445 gnd.n568 585
R8257 gnd.n6448 gnd.n6447 585
R8258 gnd.n6447 gnd.n6446 585
R8259 gnd.n565 gnd.n564 585
R8260 gnd.n564 gnd.n563 585
R8261 gnd.n6453 gnd.n6452 585
R8262 gnd.n6454 gnd.n6453 585
R8263 gnd.n562 gnd.n561 585
R8264 gnd.n6455 gnd.n562 585
R8265 gnd.n6458 gnd.n6457 585
R8266 gnd.n6457 gnd.n6456 585
R8267 gnd.n559 gnd.n558 585
R8268 gnd.n558 gnd.n557 585
R8269 gnd.n6463 gnd.n6462 585
R8270 gnd.n6464 gnd.n6463 585
R8271 gnd.n556 gnd.n555 585
R8272 gnd.n6465 gnd.n556 585
R8273 gnd.n6468 gnd.n6467 585
R8274 gnd.n6467 gnd.n6466 585
R8275 gnd.n553 gnd.n552 585
R8276 gnd.n552 gnd.n551 585
R8277 gnd.n6473 gnd.n6472 585
R8278 gnd.n6474 gnd.n6473 585
R8279 gnd.n550 gnd.n549 585
R8280 gnd.n6475 gnd.n550 585
R8281 gnd.n6478 gnd.n6477 585
R8282 gnd.n6477 gnd.n6476 585
R8283 gnd.n547 gnd.n546 585
R8284 gnd.n546 gnd.n545 585
R8285 gnd.n6483 gnd.n6482 585
R8286 gnd.n6484 gnd.n6483 585
R8287 gnd.n544 gnd.n543 585
R8288 gnd.n6485 gnd.n544 585
R8289 gnd.n6488 gnd.n6487 585
R8290 gnd.n6487 gnd.n6486 585
R8291 gnd.n541 gnd.n540 585
R8292 gnd.n540 gnd.n539 585
R8293 gnd.n6493 gnd.n6492 585
R8294 gnd.n6494 gnd.n6493 585
R8295 gnd.n538 gnd.n537 585
R8296 gnd.n6495 gnd.n538 585
R8297 gnd.n6498 gnd.n6497 585
R8298 gnd.n6497 gnd.n6496 585
R8299 gnd.n535 gnd.n534 585
R8300 gnd.n534 gnd.n533 585
R8301 gnd.n6503 gnd.n6502 585
R8302 gnd.n6504 gnd.n6503 585
R8303 gnd.n532 gnd.n531 585
R8304 gnd.n6505 gnd.n532 585
R8305 gnd.n6508 gnd.n6507 585
R8306 gnd.n6507 gnd.n6506 585
R8307 gnd.n529 gnd.n528 585
R8308 gnd.n528 gnd.n527 585
R8309 gnd.n6513 gnd.n6512 585
R8310 gnd.n6514 gnd.n6513 585
R8311 gnd.n526 gnd.n525 585
R8312 gnd.n6515 gnd.n526 585
R8313 gnd.n6518 gnd.n6517 585
R8314 gnd.n6517 gnd.n6516 585
R8315 gnd.n523 gnd.n522 585
R8316 gnd.n522 gnd.n521 585
R8317 gnd.n6523 gnd.n6522 585
R8318 gnd.n6524 gnd.n6523 585
R8319 gnd.n520 gnd.n519 585
R8320 gnd.n6525 gnd.n520 585
R8321 gnd.n6528 gnd.n6527 585
R8322 gnd.n6527 gnd.n6526 585
R8323 gnd.n517 gnd.n516 585
R8324 gnd.n516 gnd.n515 585
R8325 gnd.n6533 gnd.n6532 585
R8326 gnd.n6534 gnd.n6533 585
R8327 gnd.n514 gnd.n513 585
R8328 gnd.n6535 gnd.n514 585
R8329 gnd.n6538 gnd.n6537 585
R8330 gnd.n6537 gnd.n6536 585
R8331 gnd.n511 gnd.n510 585
R8332 gnd.n510 gnd.n509 585
R8333 gnd.n6543 gnd.n6542 585
R8334 gnd.n6544 gnd.n6543 585
R8335 gnd.n508 gnd.n507 585
R8336 gnd.n6545 gnd.n508 585
R8337 gnd.n6548 gnd.n6547 585
R8338 gnd.n6547 gnd.n6546 585
R8339 gnd.n505 gnd.n504 585
R8340 gnd.n504 gnd.n503 585
R8341 gnd.n6553 gnd.n6552 585
R8342 gnd.n6554 gnd.n6553 585
R8343 gnd.n502 gnd.n501 585
R8344 gnd.n6555 gnd.n502 585
R8345 gnd.n6558 gnd.n6557 585
R8346 gnd.n6557 gnd.n6556 585
R8347 gnd.n499 gnd.n498 585
R8348 gnd.n498 gnd.n497 585
R8349 gnd.n6563 gnd.n6562 585
R8350 gnd.n6564 gnd.n6563 585
R8351 gnd.n496 gnd.n495 585
R8352 gnd.n6565 gnd.n496 585
R8353 gnd.n6568 gnd.n6567 585
R8354 gnd.n6567 gnd.n6566 585
R8355 gnd.n493 gnd.n492 585
R8356 gnd.n492 gnd.n491 585
R8357 gnd.n6573 gnd.n6572 585
R8358 gnd.n6574 gnd.n6573 585
R8359 gnd.n490 gnd.n489 585
R8360 gnd.n6575 gnd.n490 585
R8361 gnd.n6578 gnd.n6577 585
R8362 gnd.n6577 gnd.n6576 585
R8363 gnd.n487 gnd.n486 585
R8364 gnd.n486 gnd.n485 585
R8365 gnd.n6583 gnd.n6582 585
R8366 gnd.n6584 gnd.n6583 585
R8367 gnd.n484 gnd.n483 585
R8368 gnd.n6585 gnd.n484 585
R8369 gnd.n6588 gnd.n6587 585
R8370 gnd.n6587 gnd.n6586 585
R8371 gnd.n481 gnd.n480 585
R8372 gnd.n480 gnd.n479 585
R8373 gnd.n6593 gnd.n6592 585
R8374 gnd.n6594 gnd.n6593 585
R8375 gnd.n478 gnd.n477 585
R8376 gnd.n6595 gnd.n478 585
R8377 gnd.n6598 gnd.n6597 585
R8378 gnd.n6597 gnd.n6596 585
R8379 gnd.n475 gnd.n474 585
R8380 gnd.n474 gnd.n473 585
R8381 gnd.n6603 gnd.n6602 585
R8382 gnd.n6604 gnd.n6603 585
R8383 gnd.n472 gnd.n471 585
R8384 gnd.n6605 gnd.n472 585
R8385 gnd.n6608 gnd.n6607 585
R8386 gnd.n6607 gnd.n6606 585
R8387 gnd.n469 gnd.n468 585
R8388 gnd.n468 gnd.n467 585
R8389 gnd.n6613 gnd.n6612 585
R8390 gnd.n6614 gnd.n6613 585
R8391 gnd.n466 gnd.n465 585
R8392 gnd.n6615 gnd.n466 585
R8393 gnd.n6618 gnd.n6617 585
R8394 gnd.n6617 gnd.n6616 585
R8395 gnd.n463 gnd.n462 585
R8396 gnd.n462 gnd.n461 585
R8397 gnd.n6623 gnd.n6622 585
R8398 gnd.n6624 gnd.n6623 585
R8399 gnd.n460 gnd.n459 585
R8400 gnd.n6625 gnd.n460 585
R8401 gnd.n6628 gnd.n6627 585
R8402 gnd.n6627 gnd.n6626 585
R8403 gnd.n457 gnd.n456 585
R8404 gnd.n456 gnd.n455 585
R8405 gnd.n6633 gnd.n6632 585
R8406 gnd.n6634 gnd.n6633 585
R8407 gnd.n454 gnd.n453 585
R8408 gnd.n6635 gnd.n454 585
R8409 gnd.n6638 gnd.n6637 585
R8410 gnd.n6637 gnd.n6636 585
R8411 gnd.n451 gnd.n450 585
R8412 gnd.n450 gnd.n449 585
R8413 gnd.n6643 gnd.n6642 585
R8414 gnd.n6644 gnd.n6643 585
R8415 gnd.n448 gnd.n447 585
R8416 gnd.n6645 gnd.n448 585
R8417 gnd.n6648 gnd.n6647 585
R8418 gnd.n6647 gnd.n6646 585
R8419 gnd.n445 gnd.n444 585
R8420 gnd.n444 gnd.n443 585
R8421 gnd.n6653 gnd.n6652 585
R8422 gnd.n6654 gnd.n6653 585
R8423 gnd.n442 gnd.n441 585
R8424 gnd.n6655 gnd.n442 585
R8425 gnd.n6658 gnd.n6657 585
R8426 gnd.n6657 gnd.n6656 585
R8427 gnd.n439 gnd.n438 585
R8428 gnd.n438 gnd.n437 585
R8429 gnd.n6663 gnd.n6662 585
R8430 gnd.n6664 gnd.n6663 585
R8431 gnd.n436 gnd.n435 585
R8432 gnd.n6665 gnd.n436 585
R8433 gnd.n6668 gnd.n6667 585
R8434 gnd.n6667 gnd.n6666 585
R8435 gnd.n433 gnd.n432 585
R8436 gnd.n432 gnd.n431 585
R8437 gnd.n6673 gnd.n6672 585
R8438 gnd.n6674 gnd.n6673 585
R8439 gnd.n430 gnd.n429 585
R8440 gnd.n6675 gnd.n430 585
R8441 gnd.n6678 gnd.n6677 585
R8442 gnd.n6677 gnd.n6676 585
R8443 gnd.n427 gnd.n426 585
R8444 gnd.n426 gnd.n425 585
R8445 gnd.n6684 gnd.n6683 585
R8446 gnd.n6685 gnd.n6684 585
R8447 gnd.n6682 gnd.n424 585
R8448 gnd.n6686 gnd.n424 585
R8449 gnd.n6895 gnd.n298 585
R8450 gnd.n6899 gnd.n298 585
R8451 gnd.n6897 gnd.n6896 585
R8452 gnd.n6898 gnd.n6897 585
R8453 gnd.n302 gnd.n301 585
R8454 gnd.n301 gnd.n300 585
R8455 gnd.n6889 gnd.n6888 585
R8456 gnd.n6888 gnd.n6887 585
R8457 gnd.n305 gnd.n304 585
R8458 gnd.n6886 gnd.n305 585
R8459 gnd.n6884 gnd.n6883 585
R8460 gnd.n6885 gnd.n6884 585
R8461 gnd.n308 gnd.n307 585
R8462 gnd.n307 gnd.n306 585
R8463 gnd.n6879 gnd.n6878 585
R8464 gnd.n6878 gnd.n6877 585
R8465 gnd.n311 gnd.n310 585
R8466 gnd.n6876 gnd.n311 585
R8467 gnd.n6874 gnd.n6873 585
R8468 gnd.n6875 gnd.n6874 585
R8469 gnd.n314 gnd.n313 585
R8470 gnd.n313 gnd.n312 585
R8471 gnd.n6869 gnd.n6868 585
R8472 gnd.n6868 gnd.n6867 585
R8473 gnd.n317 gnd.n316 585
R8474 gnd.n6866 gnd.n317 585
R8475 gnd.n6864 gnd.n6863 585
R8476 gnd.n6865 gnd.n6864 585
R8477 gnd.n320 gnd.n319 585
R8478 gnd.n319 gnd.n318 585
R8479 gnd.n6859 gnd.n6858 585
R8480 gnd.n6858 gnd.n6857 585
R8481 gnd.n323 gnd.n322 585
R8482 gnd.n6856 gnd.n323 585
R8483 gnd.n6854 gnd.n6853 585
R8484 gnd.n6855 gnd.n6854 585
R8485 gnd.n326 gnd.n325 585
R8486 gnd.n325 gnd.n324 585
R8487 gnd.n6849 gnd.n6848 585
R8488 gnd.n6848 gnd.n6847 585
R8489 gnd.n329 gnd.n328 585
R8490 gnd.n6846 gnd.n329 585
R8491 gnd.n6844 gnd.n6843 585
R8492 gnd.n6845 gnd.n6844 585
R8493 gnd.n332 gnd.n331 585
R8494 gnd.n331 gnd.n330 585
R8495 gnd.n6839 gnd.n6838 585
R8496 gnd.n6838 gnd.n6837 585
R8497 gnd.n335 gnd.n334 585
R8498 gnd.n6836 gnd.n335 585
R8499 gnd.n6834 gnd.n6833 585
R8500 gnd.n6835 gnd.n6834 585
R8501 gnd.n338 gnd.n337 585
R8502 gnd.n337 gnd.n336 585
R8503 gnd.n6829 gnd.n6828 585
R8504 gnd.n6828 gnd.n6827 585
R8505 gnd.n341 gnd.n340 585
R8506 gnd.n6826 gnd.n341 585
R8507 gnd.n6824 gnd.n6823 585
R8508 gnd.n6825 gnd.n6824 585
R8509 gnd.n344 gnd.n343 585
R8510 gnd.n343 gnd.n342 585
R8511 gnd.n6819 gnd.n6818 585
R8512 gnd.n6818 gnd.n6817 585
R8513 gnd.n347 gnd.n346 585
R8514 gnd.n6816 gnd.n347 585
R8515 gnd.n6814 gnd.n6813 585
R8516 gnd.n6815 gnd.n6814 585
R8517 gnd.n350 gnd.n349 585
R8518 gnd.n349 gnd.n348 585
R8519 gnd.n6809 gnd.n6808 585
R8520 gnd.n6808 gnd.n6807 585
R8521 gnd.n353 gnd.n352 585
R8522 gnd.n6806 gnd.n353 585
R8523 gnd.n6804 gnd.n6803 585
R8524 gnd.n6805 gnd.n6804 585
R8525 gnd.n356 gnd.n355 585
R8526 gnd.n355 gnd.n354 585
R8527 gnd.n6799 gnd.n6798 585
R8528 gnd.n6798 gnd.n6797 585
R8529 gnd.n359 gnd.n358 585
R8530 gnd.n6796 gnd.n359 585
R8531 gnd.n6794 gnd.n6793 585
R8532 gnd.n6795 gnd.n6794 585
R8533 gnd.n362 gnd.n361 585
R8534 gnd.n361 gnd.n360 585
R8535 gnd.n6789 gnd.n6788 585
R8536 gnd.n6788 gnd.n6787 585
R8537 gnd.n365 gnd.n364 585
R8538 gnd.n6786 gnd.n365 585
R8539 gnd.n6784 gnd.n6783 585
R8540 gnd.n6785 gnd.n6784 585
R8541 gnd.n368 gnd.n367 585
R8542 gnd.n367 gnd.n366 585
R8543 gnd.n6779 gnd.n6778 585
R8544 gnd.n6778 gnd.n6777 585
R8545 gnd.n371 gnd.n370 585
R8546 gnd.n6776 gnd.n371 585
R8547 gnd.n6774 gnd.n6773 585
R8548 gnd.n6775 gnd.n6774 585
R8549 gnd.n374 gnd.n373 585
R8550 gnd.n373 gnd.n372 585
R8551 gnd.n6769 gnd.n6768 585
R8552 gnd.n6768 gnd.n6767 585
R8553 gnd.n377 gnd.n376 585
R8554 gnd.n6766 gnd.n377 585
R8555 gnd.n6764 gnd.n6763 585
R8556 gnd.n6765 gnd.n6764 585
R8557 gnd.n380 gnd.n379 585
R8558 gnd.n379 gnd.n378 585
R8559 gnd.n6759 gnd.n6758 585
R8560 gnd.n6758 gnd.n6757 585
R8561 gnd.n383 gnd.n382 585
R8562 gnd.n6756 gnd.n383 585
R8563 gnd.n6754 gnd.n6753 585
R8564 gnd.n6755 gnd.n6754 585
R8565 gnd.n386 gnd.n385 585
R8566 gnd.n385 gnd.n384 585
R8567 gnd.n6749 gnd.n6748 585
R8568 gnd.n6748 gnd.n6747 585
R8569 gnd.n389 gnd.n388 585
R8570 gnd.n6746 gnd.n389 585
R8571 gnd.n6744 gnd.n6743 585
R8572 gnd.n6745 gnd.n6744 585
R8573 gnd.n392 gnd.n391 585
R8574 gnd.n391 gnd.n390 585
R8575 gnd.n6739 gnd.n6738 585
R8576 gnd.n6738 gnd.n6737 585
R8577 gnd.n395 gnd.n394 585
R8578 gnd.n6736 gnd.n395 585
R8579 gnd.n6734 gnd.n6733 585
R8580 gnd.n6735 gnd.n6734 585
R8581 gnd.n398 gnd.n397 585
R8582 gnd.n397 gnd.n396 585
R8583 gnd.n6729 gnd.n6728 585
R8584 gnd.n6728 gnd.n6727 585
R8585 gnd.n401 gnd.n400 585
R8586 gnd.n6726 gnd.n401 585
R8587 gnd.n6724 gnd.n6723 585
R8588 gnd.n6725 gnd.n6724 585
R8589 gnd.n404 gnd.n403 585
R8590 gnd.n403 gnd.n402 585
R8591 gnd.n6719 gnd.n6718 585
R8592 gnd.n6718 gnd.n6717 585
R8593 gnd.n407 gnd.n406 585
R8594 gnd.n6716 gnd.n407 585
R8595 gnd.n6714 gnd.n6713 585
R8596 gnd.n6715 gnd.n6714 585
R8597 gnd.n410 gnd.n409 585
R8598 gnd.n409 gnd.n408 585
R8599 gnd.n6709 gnd.n6708 585
R8600 gnd.n6708 gnd.n6707 585
R8601 gnd.n413 gnd.n412 585
R8602 gnd.n6706 gnd.n413 585
R8603 gnd.n6704 gnd.n6703 585
R8604 gnd.n6705 gnd.n6704 585
R8605 gnd.n416 gnd.n415 585
R8606 gnd.n415 gnd.n414 585
R8607 gnd.n6699 gnd.n6698 585
R8608 gnd.n6698 gnd.n6697 585
R8609 gnd.n419 gnd.n418 585
R8610 gnd.n6696 gnd.n419 585
R8611 gnd.n6694 gnd.n6693 585
R8612 gnd.n6695 gnd.n6694 585
R8613 gnd.n422 gnd.n421 585
R8614 gnd.n421 gnd.n420 585
R8615 gnd.n6689 gnd.n6688 585
R8616 gnd.n6688 gnd.n6687 585
R8617 gnd.n5925 gnd.n5924 585
R8618 gnd.n5926 gnd.n5925 585
R8619 gnd.n2523 gnd.n2522 585
R8620 gnd.n4541 gnd.n2523 585
R8621 gnd.n5934 gnd.n5933 585
R8622 gnd.n5933 gnd.n5932 585
R8623 gnd.n5935 gnd.n2517 585
R8624 gnd.n4430 gnd.n2517 585
R8625 gnd.n5937 gnd.n5936 585
R8626 gnd.n5938 gnd.n5937 585
R8627 gnd.n2502 gnd.n2501 585
R8628 gnd.n4421 gnd.n2502 585
R8629 gnd.n5946 gnd.n5945 585
R8630 gnd.n5945 gnd.n5944 585
R8631 gnd.n5947 gnd.n2496 585
R8632 gnd.n4441 gnd.n2496 585
R8633 gnd.n5949 gnd.n5948 585
R8634 gnd.n5950 gnd.n5949 585
R8635 gnd.n2480 gnd.n2479 585
R8636 gnd.n4413 gnd.n2480 585
R8637 gnd.n5958 gnd.n5957 585
R8638 gnd.n5957 gnd.n5956 585
R8639 gnd.n5959 gnd.n2474 585
R8640 gnd.n4405 gnd.n2474 585
R8641 gnd.n5961 gnd.n5960 585
R8642 gnd.n5962 gnd.n5961 585
R8643 gnd.n2460 gnd.n2459 585
R8644 gnd.n4397 gnd.n2460 585
R8645 gnd.n5970 gnd.n5969 585
R8646 gnd.n5969 gnd.n5968 585
R8647 gnd.n5971 gnd.n2454 585
R8648 gnd.n4389 gnd.n2454 585
R8649 gnd.n5973 gnd.n5972 585
R8650 gnd.n5974 gnd.n5973 585
R8651 gnd.n2441 gnd.n2440 585
R8652 gnd.n4339 gnd.n2441 585
R8653 gnd.n5983 gnd.n5982 585
R8654 gnd.n5982 gnd.n5981 585
R8655 gnd.n5984 gnd.n2436 585
R8656 gnd.n4327 gnd.n2436 585
R8657 gnd.n5986 gnd.n5985 585
R8658 gnd.n5987 gnd.n5986 585
R8659 gnd.n2425 gnd.n2424 585
R8660 gnd.n4312 gnd.n2425 585
R8661 gnd.n5996 gnd.n5995 585
R8662 gnd.n5995 gnd.n5994 585
R8663 gnd.n5997 gnd.n2419 585
R8664 gnd.n4352 gnd.n2419 585
R8665 gnd.n5999 gnd.n5998 585
R8666 gnd.n6000 gnd.n5999 585
R8667 gnd.n2405 gnd.n2404 585
R8668 gnd.n4304 gnd.n2405 585
R8669 gnd.n6009 gnd.n6008 585
R8670 gnd.n6008 gnd.n6007 585
R8671 gnd.n6010 gnd.n2399 585
R8672 gnd.n4295 gnd.n2399 585
R8673 gnd.n6012 gnd.n6011 585
R8674 gnd.n6013 gnd.n6012 585
R8675 gnd.n2384 gnd.n2383 585
R8676 gnd.n4286 gnd.n2384 585
R8677 gnd.n6021 gnd.n6020 585
R8678 gnd.n6020 gnd.n6019 585
R8679 gnd.n6022 gnd.n2378 585
R8680 gnd.n4278 gnd.n2378 585
R8681 gnd.n6024 gnd.n6023 585
R8682 gnd.n6025 gnd.n6024 585
R8683 gnd.n2362 gnd.n2361 585
R8684 gnd.n4223 gnd.n2362 585
R8685 gnd.n6033 gnd.n6032 585
R8686 gnd.n6032 gnd.n6031 585
R8687 gnd.n6034 gnd.n2356 585
R8688 gnd.n4229 gnd.n2356 585
R8689 gnd.n6036 gnd.n6035 585
R8690 gnd.n6037 gnd.n6036 585
R8691 gnd.n2340 gnd.n2339 585
R8692 gnd.n4235 gnd.n2340 585
R8693 gnd.n6045 gnd.n6044 585
R8694 gnd.n6044 gnd.n6043 585
R8695 gnd.n6046 gnd.n2334 585
R8696 gnd.n4241 gnd.n2334 585
R8697 gnd.n6048 gnd.n6047 585
R8698 gnd.n6049 gnd.n6048 585
R8699 gnd.n2335 gnd.n2333 585
R8700 gnd.n4247 gnd.n2333 585
R8701 gnd.n4001 gnd.n2322 585
R8702 gnd.n6055 gnd.n2322 585
R8703 gnd.n4005 gnd.n4004 585
R8704 gnd.n4007 gnd.n3999 585
R8705 gnd.n4010 gnd.n4009 585
R8706 gnd.n3997 gnd.n3996 585
R8707 gnd.n4015 gnd.n4014 585
R8708 gnd.n4017 gnd.n3995 585
R8709 gnd.n4020 gnd.n4019 585
R8710 gnd.n3993 gnd.n3992 585
R8711 gnd.n4025 gnd.n4024 585
R8712 gnd.n4027 gnd.n3991 585
R8713 gnd.n4030 gnd.n4029 585
R8714 gnd.n3989 gnd.n3988 585
R8715 gnd.n4035 gnd.n4034 585
R8716 gnd.n4037 gnd.n3987 585
R8717 gnd.n4040 gnd.n4039 585
R8718 gnd.n3985 gnd.n3984 585
R8719 gnd.n4045 gnd.n4044 585
R8720 gnd.n4047 gnd.n3983 585
R8721 gnd.n4049 gnd.n4048 585
R8722 gnd.n4048 gnd.n2318 585
R8723 gnd.n3843 gnd.n3842 585
R8724 gnd.n3840 gnd.n3834 585
R8725 gnd.n3850 gnd.n3831 585
R8726 gnd.n3851 gnd.n3829 585
R8727 gnd.n3828 gnd.n3821 585
R8728 gnd.n3858 gnd.n3820 585
R8729 gnd.n3859 gnd.n3819 585
R8730 gnd.n3817 gnd.n3809 585
R8731 gnd.n3866 gnd.n3808 585
R8732 gnd.n3867 gnd.n3806 585
R8733 gnd.n3805 gnd.n3798 585
R8734 gnd.n3874 gnd.n3797 585
R8735 gnd.n3875 gnd.n3796 585
R8736 gnd.n3794 gnd.n3787 585
R8737 gnd.n3882 gnd.n3786 585
R8738 gnd.n3883 gnd.n3784 585
R8739 gnd.n3783 gnd.n3779 585
R8740 gnd.n3781 gnd.n3780 585
R8741 gnd.n2540 gnd.n2538 585
R8742 gnd.n3680 gnd.n2538 585
R8743 gnd.n3716 gnd.n2536 585
R8744 gnd.n5926 gnd.n2536 585
R8745 gnd.n4540 gnd.n4539 585
R8746 gnd.n4541 gnd.n4540 585
R8747 gnd.n3715 gnd.n2526 585
R8748 gnd.n5932 gnd.n2526 585
R8749 gnd.n4433 gnd.n4431 585
R8750 gnd.n4431 gnd.n4430 585
R8751 gnd.n4434 gnd.n2515 585
R8752 gnd.n5938 gnd.n2515 585
R8753 gnd.n4435 gnd.n3910 585
R8754 gnd.n4421 gnd.n3910 585
R8755 gnd.n3907 gnd.n2504 585
R8756 gnd.n5944 gnd.n2504 585
R8757 gnd.n4440 gnd.n4439 585
R8758 gnd.n4441 gnd.n4440 585
R8759 gnd.n3906 gnd.n2494 585
R8760 gnd.n5950 gnd.n2494 585
R8761 gnd.n4412 gnd.n4411 585
R8762 gnd.n4413 gnd.n4412 585
R8763 gnd.n3916 gnd.n2483 585
R8764 gnd.n5956 gnd.n2483 585
R8765 gnd.n4407 gnd.n4406 585
R8766 gnd.n4406 gnd.n4405 585
R8767 gnd.n3918 gnd.n2473 585
R8768 gnd.n5962 gnd.n2473 585
R8769 gnd.n4396 gnd.n4395 585
R8770 gnd.n4397 gnd.n4396 585
R8771 gnd.n3923 gnd.n2462 585
R8772 gnd.n5968 gnd.n2462 585
R8773 gnd.n4391 gnd.n4390 585
R8774 gnd.n4390 gnd.n4389 585
R8775 gnd.n3925 gnd.n2452 585
R8776 gnd.n5974 gnd.n2452 585
R8777 gnd.n4342 gnd.n4340 585
R8778 gnd.n4340 gnd.n4339 585
R8779 gnd.n4343 gnd.n2444 585
R8780 gnd.n5981 gnd.n2444 585
R8781 gnd.n4344 gnd.n3949 585
R8782 gnd.n4327 gnd.n3949 585
R8783 gnd.n3947 gnd.n2435 585
R8784 gnd.n5987 gnd.n2435 585
R8785 gnd.n4348 gnd.n3946 585
R8786 gnd.n4312 gnd.n3946 585
R8787 gnd.n4349 gnd.n2427 585
R8788 gnd.n5994 gnd.n2427 585
R8789 gnd.n4351 gnd.n4350 585
R8790 gnd.n4352 gnd.n4351 585
R8791 gnd.n3943 gnd.n2417 585
R8792 gnd.n6000 gnd.n2417 585
R8793 gnd.n4303 gnd.n4302 585
R8794 gnd.n4304 gnd.n4303 585
R8795 gnd.n3957 gnd.n2408 585
R8796 gnd.n6007 gnd.n2408 585
R8797 gnd.n4297 gnd.n4296 585
R8798 gnd.n4296 gnd.n4295 585
R8799 gnd.n3959 gnd.n2397 585
R8800 gnd.n6013 gnd.n2397 585
R8801 gnd.n4285 gnd.n4284 585
R8802 gnd.n4286 gnd.n4285 585
R8803 gnd.n3963 gnd.n2386 585
R8804 gnd.n6019 gnd.n2386 585
R8805 gnd.n4280 gnd.n4279 585
R8806 gnd.n4279 gnd.n4278 585
R8807 gnd.n3965 gnd.n2376 585
R8808 gnd.n6025 gnd.n2376 585
R8809 gnd.n4222 gnd.n4221 585
R8810 gnd.n4223 gnd.n4222 585
R8811 gnd.n4210 gnd.n2365 585
R8812 gnd.n6031 gnd.n2365 585
R8813 gnd.n4231 gnd.n4230 585
R8814 gnd.n4230 gnd.n4229 585
R8815 gnd.n4232 gnd.n2354 585
R8816 gnd.n6037 gnd.n2354 585
R8817 gnd.n4234 gnd.n4233 585
R8818 gnd.n4235 gnd.n4234 585
R8819 gnd.n4055 gnd.n2343 585
R8820 gnd.n6043 gnd.n2343 585
R8821 gnd.n4243 gnd.n4242 585
R8822 gnd.n4242 gnd.n4241 585
R8823 gnd.n4244 gnd.n2331 585
R8824 gnd.n6049 gnd.n2331 585
R8825 gnd.n4246 gnd.n4245 585
R8826 gnd.n4247 gnd.n4246 585
R8827 gnd.n3979 gnd.n2320 585
R8828 gnd.n6055 gnd.n2320 585
R8829 gnd.n165 gnd.n84 585
R8830 gnd.n7193 gnd.n84 585
R8831 gnd.n7113 gnd.n7112 585
R8832 gnd.n7114 gnd.n7113 585
R8833 gnd.n164 gnd.n163 585
R8834 gnd.n173 gnd.n163 585
R8835 gnd.n7041 gnd.n7040 585
R8836 gnd.n7040 gnd.n7039 585
R8837 gnd.n168 gnd.n167 585
R8838 gnd.n6926 gnd.n168 585
R8839 gnd.n7028 gnd.n7027 585
R8840 gnd.n7029 gnd.n7028 585
R8841 gnd.n184 gnd.n183 585
R8842 gnd.n6932 gnd.n183 585
R8843 gnd.n7023 gnd.n7022 585
R8844 gnd.n7022 gnd.n7021 585
R8845 gnd.n187 gnd.n186 585
R8846 gnd.n6915 gnd.n187 585
R8847 gnd.n7012 gnd.n7011 585
R8848 gnd.n7013 gnd.n7012 585
R8849 gnd.n199 gnd.n198 585
R8850 gnd.n6941 gnd.n198 585
R8851 gnd.n7007 gnd.n7006 585
R8852 gnd.n7006 gnd.n7005 585
R8853 gnd.n202 gnd.n201 585
R8854 gnd.n6945 gnd.n202 585
R8855 gnd.n6996 gnd.n6995 585
R8856 gnd.n6997 gnd.n6996 585
R8857 gnd.n216 gnd.n215 585
R8858 gnd.n6951 gnd.n215 585
R8859 gnd.n6991 gnd.n6990 585
R8860 gnd.n6990 gnd.n6989 585
R8861 gnd.n219 gnd.n218 585
R8862 gnd.n5700 gnd.n219 585
R8863 gnd.n6967 gnd.n6966 585
R8864 gnd.n6966 gnd.n6965 585
R8865 gnd.n6968 gnd.n248 585
R8866 gnd.n6961 gnd.n248 585
R8867 gnd.n5707 gnd.n246 585
R8868 gnd.n5708 gnd.n5707 585
R8869 gnd.n6972 gnd.n245 585
R8870 gnd.n2726 gnd.n245 585
R8871 gnd.n6973 gnd.n244 585
R8872 gnd.n5727 gnd.n244 585
R8873 gnd.n6974 gnd.n243 585
R8874 gnd.n5732 gnd.n243 585
R8875 gnd.n240 gnd.n238 585
R8876 gnd.n5716 gnd.n238 585
R8877 gnd.n6979 gnd.n6978 585
R8878 gnd.n6980 gnd.n6979 585
R8879 gnd.n239 gnd.n237 585
R8880 gnd.n5686 gnd.n237 585
R8881 gnd.n5749 gnd.n5748 585
R8882 gnd.n5748 gnd.n5747 585
R8883 gnd.n2703 gnd.n2702 585
R8884 gnd.n5744 gnd.n2703 585
R8885 gnd.n5753 gnd.n2701 585
R8886 gnd.n2740 gnd.n2701 585
R8887 gnd.n5754 gnd.n2700 585
R8888 gnd.n5678 gnd.n2700 585
R8889 gnd.n5755 gnd.n2699 585
R8890 gnd.n5631 gnd.n2699 585
R8891 gnd.n5667 gnd.n2697 585
R8892 gnd.n5668 gnd.n5667 585
R8893 gnd.n5759 gnd.n2696 585
R8894 gnd.n5640 gnd.n2696 585
R8895 gnd.n5760 gnd.n2695 585
R8896 gnd.n5582 gnd.n2695 585
R8897 gnd.n5761 gnd.n2694 585
R8898 gnd.n5625 gnd.n2694 585
R8899 gnd.n2775 gnd.n2692 585
R8900 gnd.n2776 gnd.n2775 585
R8901 gnd.n5765 gnd.n2691 585
R8902 gnd.n5615 gnd.n2691 585
R8903 gnd.n5766 gnd.n2690 585
R8904 gnd.n5603 gnd.n2690 585
R8905 gnd.n5767 gnd.n2689 585
R8906 gnd.n2794 gnd.n2689 585
R8907 gnd.n2686 gnd.n2684 585
R8908 gnd.n5594 gnd.n2684 585
R8909 gnd.n5772 gnd.n5771 585
R8910 gnd.n5773 gnd.n5772 585
R8911 gnd.n2685 gnd.n2683 585
R8912 gnd.n5566 gnd.n2683 585
R8913 gnd.n2853 gnd.n2671 585
R8914 gnd.n5779 gnd.n2671 585
R8915 gnd.n2857 gnd.n2856 585
R8916 gnd.n2859 gnd.n2850 585
R8917 gnd.n2862 gnd.n2861 585
R8918 gnd.n2843 gnd.n2842 585
R8919 gnd.n2876 gnd.n2875 585
R8920 gnd.n2878 gnd.n2841 585
R8921 gnd.n2881 gnd.n2880 585
R8922 gnd.n2834 gnd.n2833 585
R8923 gnd.n2895 gnd.n2894 585
R8924 gnd.n2897 gnd.n2832 585
R8925 gnd.n2900 gnd.n2899 585
R8926 gnd.n2825 gnd.n2824 585
R8927 gnd.n2914 gnd.n2913 585
R8928 gnd.n2916 gnd.n2823 585
R8929 gnd.n2919 gnd.n2918 585
R8930 gnd.n2816 gnd.n2815 585
R8931 gnd.n2933 gnd.n2932 585
R8932 gnd.n2935 gnd.n2814 585
R8933 gnd.n2937 gnd.n2936 585
R8934 gnd.n2936 gnd.n2659 585
R8935 gnd.n7082 gnd.n80 585
R8936 gnd.n7083 gnd.n7081 585
R8937 gnd.n7084 gnd.n7077 585
R8938 gnd.n7075 gnd.n7073 585
R8939 gnd.n7088 gnd.n7072 585
R8940 gnd.n7089 gnd.n7070 585
R8941 gnd.n7090 gnd.n7069 585
R8942 gnd.n7067 gnd.n7065 585
R8943 gnd.n7094 gnd.n7064 585
R8944 gnd.n7095 gnd.n7062 585
R8945 gnd.n7096 gnd.n7061 585
R8946 gnd.n7059 gnd.n7057 585
R8947 gnd.n7100 gnd.n7056 585
R8948 gnd.n7101 gnd.n7054 585
R8949 gnd.n7102 gnd.n7053 585
R8950 gnd.n7051 gnd.n7049 585
R8951 gnd.n7106 gnd.n7048 585
R8952 gnd.n7107 gnd.n7046 585
R8953 gnd.n7108 gnd.n7045 585
R8954 gnd.n7045 gnd.n94 585
R8955 gnd.n7195 gnd.n7194 585
R8956 gnd.n7194 gnd.n7193 585
R8957 gnd.n79 gnd.n77 585
R8958 gnd.n7114 gnd.n79 585
R8959 gnd.n7199 gnd.n76 585
R8960 gnd.n173 gnd.n76 585
R8961 gnd.n7200 gnd.n75 585
R8962 gnd.n7039 gnd.n75 585
R8963 gnd.n7201 gnd.n74 585
R8964 gnd.n6926 gnd.n74 585
R8965 gnd.n181 gnd.n72 585
R8966 gnd.n7029 gnd.n181 585
R8967 gnd.n7205 gnd.n71 585
R8968 gnd.n6932 gnd.n71 585
R8969 gnd.n7206 gnd.n70 585
R8970 gnd.n7021 gnd.n70 585
R8971 gnd.n7207 gnd.n69 585
R8972 gnd.n6915 gnd.n69 585
R8973 gnd.n196 gnd.n67 585
R8974 gnd.n7013 gnd.n196 585
R8975 gnd.n7211 gnd.n66 585
R8976 gnd.n6941 gnd.n66 585
R8977 gnd.n7212 gnd.n65 585
R8978 gnd.n7005 gnd.n65 585
R8979 gnd.n7213 gnd.n64 585
R8980 gnd.n6945 gnd.n64 585
R8981 gnd.n213 gnd.n62 585
R8982 gnd.n6997 gnd.n213 585
R8983 gnd.n7217 gnd.n61 585
R8984 gnd.n6951 gnd.n61 585
R8985 gnd.n7218 gnd.n60 585
R8986 gnd.n6989 gnd.n60 585
R8987 gnd.n7219 gnd.n59 585
R8988 gnd.n5700 gnd.n59 585
R8989 gnd.n250 gnd.n57 585
R8990 gnd.n6965 gnd.n250 585
R8991 gnd.n7223 gnd.n56 585
R8992 gnd.n6961 gnd.n56 585
R8993 gnd.n7224 gnd.n55 585
R8994 gnd.n5708 gnd.n55 585
R8995 gnd.n7225 gnd.n54 585
R8996 gnd.n2726 gnd.n54 585
R8997 gnd.n2719 gnd.n52 585
R8998 gnd.n5727 gnd.n2719 585
R8999 gnd.n5734 gnd.n5733 585
R9000 gnd.n5733 gnd.n5732 585
R9001 gnd.n5736 gnd.n2718 585
R9002 gnd.n5716 gnd.n2718 585
R9003 gnd.n5737 gnd.n235 585
R9004 gnd.n6980 gnd.n235 585
R9005 gnd.n5738 gnd.n2717 585
R9006 gnd.n5686 gnd.n2717 585
R9007 gnd.n2714 gnd.n2706 585
R9008 gnd.n5747 gnd.n2706 585
R9009 gnd.n5743 gnd.n5742 585
R9010 gnd.n5744 gnd.n5743 585
R9011 gnd.n2713 gnd.n2712 585
R9012 gnd.n2740 gnd.n2712 585
R9013 gnd.n5633 gnd.n2739 585
R9014 gnd.n5678 gnd.n2739 585
R9015 gnd.n5634 gnd.n5632 585
R9016 gnd.n5632 gnd.n5631 585
R9017 gnd.n2759 gnd.n2749 585
R9018 gnd.n5668 gnd.n2749 585
R9019 gnd.n5639 gnd.n5638 585
R9020 gnd.n5640 gnd.n5639 585
R9021 gnd.n2758 gnd.n2757 585
R9022 gnd.n5582 gnd.n2757 585
R9023 gnd.n5627 gnd.n5626 585
R9024 gnd.n5626 gnd.n5625 585
R9025 gnd.n2762 gnd.n2761 585
R9026 gnd.n2776 gnd.n2762 585
R9027 gnd.n2798 gnd.n2774 585
R9028 gnd.n5615 gnd.n2774 585
R9029 gnd.n5602 gnd.n5601 585
R9030 gnd.n5603 gnd.n5602 585
R9031 gnd.n2797 gnd.n2796 585
R9032 gnd.n2796 gnd.n2794 585
R9033 gnd.n5596 gnd.n5595 585
R9034 gnd.n5595 gnd.n5594 585
R9035 gnd.n2800 gnd.n2681 585
R9036 gnd.n5773 gnd.n2681 585
R9037 gnd.n5565 gnd.n5564 585
R9038 gnd.n5566 gnd.n5565 585
R9039 gnd.n2805 gnd.n2669 585
R9040 gnd.n5779 gnd.n2669 585
R9041 gnd.n2224 gnd.n2223 585
R9042 gnd.n2225 gnd.n2224 585
R9043 gnd.n943 gnd.n942 585
R9044 gnd.n949 gnd.n942 585
R9045 gnd.n2199 gnd.n961 585
R9046 gnd.n961 gnd.n948 585
R9047 gnd.n2201 gnd.n2200 585
R9048 gnd.n2202 gnd.n2201 585
R9049 gnd.n962 gnd.n960 585
R9050 gnd.n960 gnd.n956 585
R9051 gnd.n1933 gnd.n1932 585
R9052 gnd.n1932 gnd.n1931 585
R9053 gnd.n967 gnd.n966 585
R9054 gnd.n1902 gnd.n967 585
R9055 gnd.n1922 gnd.n1921 585
R9056 gnd.n1921 gnd.n1920 585
R9057 gnd.n974 gnd.n973 585
R9058 gnd.n1908 gnd.n974 585
R9059 gnd.n1878 gnd.n994 585
R9060 gnd.n994 gnd.n993 585
R9061 gnd.n1880 gnd.n1879 585
R9062 gnd.n1881 gnd.n1880 585
R9063 gnd.n995 gnd.n992 585
R9064 gnd.n1003 gnd.n992 585
R9065 gnd.n1856 gnd.n1015 585
R9066 gnd.n1015 gnd.n1002 585
R9067 gnd.n1858 gnd.n1857 585
R9068 gnd.n1859 gnd.n1858 585
R9069 gnd.n1016 gnd.n1014 585
R9070 gnd.n1014 gnd.n1010 585
R9071 gnd.n1844 gnd.n1843 585
R9072 gnd.n1843 gnd.n1842 585
R9073 gnd.n1021 gnd.n1020 585
R9074 gnd.n1030 gnd.n1021 585
R9075 gnd.n1833 gnd.n1832 585
R9076 gnd.n1832 gnd.n1831 585
R9077 gnd.n1028 gnd.n1027 585
R9078 gnd.n1819 gnd.n1028 585
R9079 gnd.n1791 gnd.n1047 585
R9080 gnd.n1047 gnd.n1037 585
R9081 gnd.n1793 gnd.n1792 585
R9082 gnd.n1794 gnd.n1793 585
R9083 gnd.n1048 gnd.n1046 585
R9084 gnd.n1056 gnd.n1046 585
R9085 gnd.n1769 gnd.n1068 585
R9086 gnd.n1068 gnd.n1055 585
R9087 gnd.n1771 gnd.n1770 585
R9088 gnd.n1772 gnd.n1771 585
R9089 gnd.n1069 gnd.n1067 585
R9090 gnd.n1067 gnd.n1063 585
R9091 gnd.n1757 gnd.n1756 585
R9092 gnd.n1756 gnd.n1755 585
R9093 gnd.n1074 gnd.n1073 585
R9094 gnd.n1083 gnd.n1074 585
R9095 gnd.n1746 gnd.n1745 585
R9096 gnd.n1745 gnd.n1744 585
R9097 gnd.n1081 gnd.n1080 585
R9098 gnd.n1732 gnd.n1081 585
R9099 gnd.n1170 gnd.n1169 585
R9100 gnd.n1170 gnd.n1090 585
R9101 gnd.n1689 gnd.n1688 585
R9102 gnd.n1688 gnd.n1687 585
R9103 gnd.n1690 gnd.n1164 585
R9104 gnd.n1175 gnd.n1164 585
R9105 gnd.n1692 gnd.n1691 585
R9106 gnd.n1693 gnd.n1692 585
R9107 gnd.n1165 gnd.n1163 585
R9108 gnd.n1188 gnd.n1163 585
R9109 gnd.n1148 gnd.n1147 585
R9110 gnd.n1151 gnd.n1148 585
R9111 gnd.n1703 gnd.n1702 585
R9112 gnd.n1702 gnd.n1701 585
R9113 gnd.n1704 gnd.n1142 585
R9114 gnd.n1663 gnd.n1142 585
R9115 gnd.n1706 gnd.n1705 585
R9116 gnd.n1707 gnd.n1706 585
R9117 gnd.n1143 gnd.n1141 585
R9118 gnd.n1202 gnd.n1141 585
R9119 gnd.n1655 gnd.n1654 585
R9120 gnd.n1654 gnd.n1653 585
R9121 gnd.n1199 gnd.n1198 585
R9122 gnd.n1637 gnd.n1199 585
R9123 gnd.n1624 gnd.n1218 585
R9124 gnd.n1218 gnd.n1217 585
R9125 gnd.n1626 gnd.n1625 585
R9126 gnd.n1627 gnd.n1626 585
R9127 gnd.n1219 gnd.n1216 585
R9128 gnd.n1225 gnd.n1216 585
R9129 gnd.n1605 gnd.n1604 585
R9130 gnd.n1606 gnd.n1605 585
R9131 gnd.n1236 gnd.n1235 585
R9132 gnd.n1235 gnd.n1231 585
R9133 gnd.n1595 gnd.n1594 585
R9134 gnd.n1596 gnd.n1595 585
R9135 gnd.n1246 gnd.n1245 585
R9136 gnd.n1251 gnd.n1245 585
R9137 gnd.n1573 gnd.n1264 585
R9138 gnd.n1264 gnd.n1250 585
R9139 gnd.n1575 gnd.n1574 585
R9140 gnd.n1576 gnd.n1575 585
R9141 gnd.n1265 gnd.n1263 585
R9142 gnd.n1263 gnd.n1259 585
R9143 gnd.n1564 gnd.n1563 585
R9144 gnd.n1565 gnd.n1564 585
R9145 gnd.n1272 gnd.n1271 585
R9146 gnd.n1276 gnd.n1271 585
R9147 gnd.n1541 gnd.n1293 585
R9148 gnd.n1293 gnd.n1275 585
R9149 gnd.n1543 gnd.n1542 585
R9150 gnd.n1544 gnd.n1543 585
R9151 gnd.n1294 gnd.n1292 585
R9152 gnd.n1292 gnd.n1283 585
R9153 gnd.n1536 gnd.n1535 585
R9154 gnd.n1535 gnd.n1534 585
R9155 gnd.n1341 gnd.n1340 585
R9156 gnd.n1342 gnd.n1341 585
R9157 gnd.n1495 gnd.n1494 585
R9158 gnd.n1496 gnd.n1495 585
R9159 gnd.n1351 gnd.n1350 585
R9160 gnd.n1350 gnd.n1349 585
R9161 gnd.n1490 gnd.n1489 585
R9162 gnd.n1489 gnd.n1488 585
R9163 gnd.n1354 gnd.n1353 585
R9164 gnd.n1355 gnd.n1354 585
R9165 gnd.n1479 gnd.n1478 585
R9166 gnd.n1480 gnd.n1479 585
R9167 gnd.n1362 gnd.n1361 585
R9168 gnd.n1471 gnd.n1361 585
R9169 gnd.n1474 gnd.n1473 585
R9170 gnd.n1473 gnd.n1472 585
R9171 gnd.n1365 gnd.n1364 585
R9172 gnd.n1366 gnd.n1365 585
R9173 gnd.n1460 gnd.n1459 585
R9174 gnd.n1458 gnd.n1384 585
R9175 gnd.n1457 gnd.n1383 585
R9176 gnd.n1462 gnd.n1383 585
R9177 gnd.n1456 gnd.n1455 585
R9178 gnd.n1454 gnd.n1453 585
R9179 gnd.n1452 gnd.n1451 585
R9180 gnd.n1450 gnd.n1449 585
R9181 gnd.n1448 gnd.n1447 585
R9182 gnd.n1446 gnd.n1445 585
R9183 gnd.n1444 gnd.n1443 585
R9184 gnd.n1442 gnd.n1441 585
R9185 gnd.n1440 gnd.n1439 585
R9186 gnd.n1438 gnd.n1437 585
R9187 gnd.n1436 gnd.n1435 585
R9188 gnd.n1434 gnd.n1433 585
R9189 gnd.n1432 gnd.n1431 585
R9190 gnd.n1430 gnd.n1429 585
R9191 gnd.n1428 gnd.n1427 585
R9192 gnd.n1426 gnd.n1425 585
R9193 gnd.n1424 gnd.n1423 585
R9194 gnd.n1422 gnd.n1421 585
R9195 gnd.n1420 gnd.n1419 585
R9196 gnd.n1418 gnd.n1417 585
R9197 gnd.n1416 gnd.n1415 585
R9198 gnd.n1414 gnd.n1413 585
R9199 gnd.n1371 gnd.n1370 585
R9200 gnd.n1465 gnd.n1464 585
R9201 gnd.n2228 gnd.n2227 585
R9202 gnd.n2230 gnd.n2229 585
R9203 gnd.n2232 gnd.n2231 585
R9204 gnd.n2234 gnd.n2233 585
R9205 gnd.n2236 gnd.n2235 585
R9206 gnd.n2238 gnd.n2237 585
R9207 gnd.n2240 gnd.n2239 585
R9208 gnd.n2242 gnd.n2241 585
R9209 gnd.n2244 gnd.n2243 585
R9210 gnd.n2246 gnd.n2245 585
R9211 gnd.n2248 gnd.n2247 585
R9212 gnd.n2250 gnd.n2249 585
R9213 gnd.n2252 gnd.n2251 585
R9214 gnd.n2254 gnd.n2253 585
R9215 gnd.n2256 gnd.n2255 585
R9216 gnd.n2258 gnd.n2257 585
R9217 gnd.n2260 gnd.n2259 585
R9218 gnd.n2262 gnd.n2261 585
R9219 gnd.n2264 gnd.n2263 585
R9220 gnd.n2266 gnd.n2265 585
R9221 gnd.n2268 gnd.n2267 585
R9222 gnd.n2270 gnd.n2269 585
R9223 gnd.n2272 gnd.n2271 585
R9224 gnd.n2274 gnd.n2273 585
R9225 gnd.n2276 gnd.n2275 585
R9226 gnd.n2277 gnd.n910 585
R9227 gnd.n2278 gnd.n868 585
R9228 gnd.n2316 gnd.n868 585
R9229 gnd.n2226 gnd.n940 585
R9230 gnd.n2226 gnd.n2225 585
R9231 gnd.n1895 gnd.n939 585
R9232 gnd.n949 gnd.n939 585
R9233 gnd.n1897 gnd.n1896 585
R9234 gnd.n1896 gnd.n948 585
R9235 gnd.n1898 gnd.n958 585
R9236 gnd.n2202 gnd.n958 585
R9237 gnd.n1900 gnd.n1899 585
R9238 gnd.n1899 gnd.n956 585
R9239 gnd.n1901 gnd.n969 585
R9240 gnd.n1931 gnd.n969 585
R9241 gnd.n1904 gnd.n1903 585
R9242 gnd.n1903 gnd.n1902 585
R9243 gnd.n1905 gnd.n976 585
R9244 gnd.n1920 gnd.n976 585
R9245 gnd.n1907 gnd.n1906 585
R9246 gnd.n1908 gnd.n1907 585
R9247 gnd.n986 gnd.n985 585
R9248 gnd.n993 gnd.n985 585
R9249 gnd.n1883 gnd.n1882 585
R9250 gnd.n1882 gnd.n1881 585
R9251 gnd.n989 gnd.n988 585
R9252 gnd.n1003 gnd.n989 585
R9253 gnd.n1807 gnd.n1806 585
R9254 gnd.n1806 gnd.n1002 585
R9255 gnd.n1808 gnd.n1012 585
R9256 gnd.n1859 gnd.n1012 585
R9257 gnd.n1810 gnd.n1809 585
R9258 gnd.n1809 gnd.n1010 585
R9259 gnd.n1811 gnd.n1023 585
R9260 gnd.n1842 gnd.n1023 585
R9261 gnd.n1813 gnd.n1812 585
R9262 gnd.n1812 gnd.n1030 585
R9263 gnd.n1814 gnd.n1029 585
R9264 gnd.n1831 gnd.n1029 585
R9265 gnd.n1816 gnd.n1815 585
R9266 gnd.n1819 gnd.n1816 585
R9267 gnd.n1040 gnd.n1039 585
R9268 gnd.n1039 gnd.n1037 585
R9269 gnd.n1796 gnd.n1795 585
R9270 gnd.n1795 gnd.n1794 585
R9271 gnd.n1043 gnd.n1042 585
R9272 gnd.n1056 gnd.n1043 585
R9273 gnd.n1720 gnd.n1719 585
R9274 gnd.n1719 gnd.n1055 585
R9275 gnd.n1721 gnd.n1065 585
R9276 gnd.n1772 gnd.n1065 585
R9277 gnd.n1723 gnd.n1722 585
R9278 gnd.n1722 gnd.n1063 585
R9279 gnd.n1724 gnd.n1076 585
R9280 gnd.n1755 gnd.n1076 585
R9281 gnd.n1726 gnd.n1725 585
R9282 gnd.n1725 gnd.n1083 585
R9283 gnd.n1727 gnd.n1082 585
R9284 gnd.n1744 gnd.n1082 585
R9285 gnd.n1729 gnd.n1728 585
R9286 gnd.n1732 gnd.n1729 585
R9287 gnd.n1093 gnd.n1092 585
R9288 gnd.n1092 gnd.n1090 585
R9289 gnd.n1172 gnd.n1171 585
R9290 gnd.n1687 gnd.n1171 585
R9291 gnd.n1174 gnd.n1173 585
R9292 gnd.n1175 gnd.n1174 585
R9293 gnd.n1185 gnd.n1161 585
R9294 gnd.n1693 gnd.n1161 585
R9295 gnd.n1187 gnd.n1186 585
R9296 gnd.n1188 gnd.n1187 585
R9297 gnd.n1184 gnd.n1183 585
R9298 gnd.n1184 gnd.n1151 585
R9299 gnd.n1182 gnd.n1149 585
R9300 gnd.n1701 gnd.n1149 585
R9301 gnd.n1138 gnd.n1136 585
R9302 gnd.n1663 gnd.n1138 585
R9303 gnd.n1709 gnd.n1708 585
R9304 gnd.n1708 gnd.n1707 585
R9305 gnd.n1137 gnd.n1135 585
R9306 gnd.n1202 gnd.n1137 585
R9307 gnd.n1634 gnd.n1201 585
R9308 gnd.n1653 gnd.n1201 585
R9309 gnd.n1636 gnd.n1635 585
R9310 gnd.n1637 gnd.n1636 585
R9311 gnd.n1211 gnd.n1210 585
R9312 gnd.n1217 gnd.n1210 585
R9313 gnd.n1629 gnd.n1628 585
R9314 gnd.n1628 gnd.n1627 585
R9315 gnd.n1214 gnd.n1213 585
R9316 gnd.n1225 gnd.n1214 585
R9317 gnd.n1514 gnd.n1233 585
R9318 gnd.n1606 gnd.n1233 585
R9319 gnd.n1516 gnd.n1515 585
R9320 gnd.n1515 gnd.n1231 585
R9321 gnd.n1517 gnd.n1244 585
R9322 gnd.n1596 gnd.n1244 585
R9323 gnd.n1519 gnd.n1518 585
R9324 gnd.n1519 gnd.n1251 585
R9325 gnd.n1521 gnd.n1520 585
R9326 gnd.n1520 gnd.n1250 585
R9327 gnd.n1522 gnd.n1261 585
R9328 gnd.n1576 gnd.n1261 585
R9329 gnd.n1524 gnd.n1523 585
R9330 gnd.n1523 gnd.n1259 585
R9331 gnd.n1525 gnd.n1270 585
R9332 gnd.n1565 gnd.n1270 585
R9333 gnd.n1527 gnd.n1526 585
R9334 gnd.n1527 gnd.n1276 585
R9335 gnd.n1529 gnd.n1528 585
R9336 gnd.n1528 gnd.n1275 585
R9337 gnd.n1530 gnd.n1291 585
R9338 gnd.n1544 gnd.n1291 585
R9339 gnd.n1531 gnd.n1344 585
R9340 gnd.n1344 gnd.n1283 585
R9341 gnd.n1533 gnd.n1532 585
R9342 gnd.n1534 gnd.n1533 585
R9343 gnd.n1345 gnd.n1343 585
R9344 gnd.n1343 gnd.n1342 585
R9345 gnd.n1498 gnd.n1497 585
R9346 gnd.n1497 gnd.n1496 585
R9347 gnd.n1348 gnd.n1347 585
R9348 gnd.n1349 gnd.n1348 585
R9349 gnd.n1487 gnd.n1486 585
R9350 gnd.n1488 gnd.n1487 585
R9351 gnd.n1357 gnd.n1356 585
R9352 gnd.n1356 gnd.n1355 585
R9353 gnd.n1482 gnd.n1481 585
R9354 gnd.n1481 gnd.n1480 585
R9355 gnd.n1360 gnd.n1359 585
R9356 gnd.n1471 gnd.n1360 585
R9357 gnd.n1470 gnd.n1469 585
R9358 gnd.n1472 gnd.n1470 585
R9359 gnd.n1368 gnd.n1367 585
R9360 gnd.n1367 gnd.n1366 585
R9361 gnd.n2211 gnd.n890 585
R9362 gnd.n890 gnd.n867 585
R9363 gnd.n2212 gnd.n951 585
R9364 gnd.n951 gnd.n941 585
R9365 gnd.n2214 gnd.n2213 585
R9366 gnd.n2215 gnd.n2214 585
R9367 gnd.n952 gnd.n950 585
R9368 gnd.n959 gnd.n950 585
R9369 gnd.n2205 gnd.n2204 585
R9370 gnd.n2204 gnd.n2203 585
R9371 gnd.n955 gnd.n954 585
R9372 gnd.n1930 gnd.n955 585
R9373 gnd.n1916 gnd.n978 585
R9374 gnd.n978 gnd.n968 585
R9375 gnd.n1918 gnd.n1917 585
R9376 gnd.n1919 gnd.n1918 585
R9377 gnd.n979 gnd.n977 585
R9378 gnd.n977 gnd.n975 585
R9379 gnd.n1911 gnd.n1910 585
R9380 gnd.n1910 gnd.n1909 585
R9381 gnd.n982 gnd.n981 585
R9382 gnd.n991 gnd.n982 585
R9383 gnd.n1867 gnd.n1005 585
R9384 gnd.n1005 gnd.n990 585
R9385 gnd.n1869 gnd.n1868 585
R9386 gnd.n1870 gnd.n1869 585
R9387 gnd.n1006 gnd.n1004 585
R9388 gnd.n1013 gnd.n1004 585
R9389 gnd.n1862 gnd.n1861 585
R9390 gnd.n1861 gnd.n1860 585
R9391 gnd.n1009 gnd.n1008 585
R9392 gnd.n1841 gnd.n1009 585
R9393 gnd.n1827 gnd.n1032 585
R9394 gnd.n1032 gnd.n1022 585
R9395 gnd.n1829 gnd.n1828 585
R9396 gnd.n1830 gnd.n1829 585
R9397 gnd.n1033 gnd.n1031 585
R9398 gnd.n1818 gnd.n1031 585
R9399 gnd.n1822 gnd.n1821 585
R9400 gnd.n1821 gnd.n1820 585
R9401 gnd.n1036 gnd.n1035 585
R9402 gnd.n1045 gnd.n1036 585
R9403 gnd.n1780 gnd.n1058 585
R9404 gnd.n1058 gnd.n1044 585
R9405 gnd.n1782 gnd.n1781 585
R9406 gnd.n1783 gnd.n1782 585
R9407 gnd.n1059 gnd.n1057 585
R9408 gnd.n1066 gnd.n1057 585
R9409 gnd.n1775 gnd.n1774 585
R9410 gnd.n1774 gnd.n1773 585
R9411 gnd.n1062 gnd.n1061 585
R9412 gnd.n1754 gnd.n1062 585
R9413 gnd.n1740 gnd.n1085 585
R9414 gnd.n1085 gnd.n1075 585
R9415 gnd.n1742 gnd.n1741 585
R9416 gnd.n1743 gnd.n1742 585
R9417 gnd.n1086 gnd.n1084 585
R9418 gnd.n1731 gnd.n1084 585
R9419 gnd.n1735 gnd.n1734 585
R9420 gnd.n1734 gnd.n1733 585
R9421 gnd.n1089 gnd.n1088 585
R9422 gnd.n1686 gnd.n1089 585
R9423 gnd.n1179 gnd.n1178 585
R9424 gnd.n1180 gnd.n1179 585
R9425 gnd.n1159 gnd.n1158 585
R9426 gnd.n1162 gnd.n1159 585
R9427 gnd.n1696 gnd.n1695 585
R9428 gnd.n1695 gnd.n1694 585
R9429 gnd.n1697 gnd.n1153 585
R9430 gnd.n1189 gnd.n1153 585
R9431 gnd.n1699 gnd.n1698 585
R9432 gnd.n1700 gnd.n1699 585
R9433 gnd.n1154 gnd.n1152 585
R9434 gnd.n1664 gnd.n1152 585
R9435 gnd.n1648 gnd.n1647 585
R9436 gnd.n1647 gnd.n1140 585
R9437 gnd.n1649 gnd.n1204 585
R9438 gnd.n1204 gnd.n1139 585
R9439 gnd.n1651 gnd.n1650 585
R9440 gnd.n1652 gnd.n1651 585
R9441 gnd.n1205 gnd.n1203 585
R9442 gnd.n1203 gnd.n1200 585
R9443 gnd.n1640 gnd.n1639 585
R9444 gnd.n1639 gnd.n1638 585
R9445 gnd.n1208 gnd.n1207 585
R9446 gnd.n1215 gnd.n1208 585
R9447 gnd.n1614 gnd.n1613 585
R9448 gnd.n1615 gnd.n1614 585
R9449 gnd.n1227 gnd.n1226 585
R9450 gnd.n1234 gnd.n1226 585
R9451 gnd.n1609 gnd.n1608 585
R9452 gnd.n1608 gnd.n1607 585
R9453 gnd.n1230 gnd.n1229 585
R9454 gnd.n1597 gnd.n1230 585
R9455 gnd.n1584 gnd.n1254 585
R9456 gnd.n1254 gnd.n1253 585
R9457 gnd.n1586 gnd.n1585 585
R9458 gnd.n1587 gnd.n1586 585
R9459 gnd.n1255 gnd.n1252 585
R9460 gnd.n1262 gnd.n1252 585
R9461 gnd.n1579 gnd.n1578 585
R9462 gnd.n1578 gnd.n1577 585
R9463 gnd.n1258 gnd.n1257 585
R9464 gnd.n1566 gnd.n1258 585
R9465 gnd.n1553 gnd.n1279 585
R9466 gnd.n1279 gnd.n1278 585
R9467 gnd.n1555 gnd.n1554 585
R9468 gnd.n1556 gnd.n1555 585
R9469 gnd.n1549 gnd.n1277 585
R9470 gnd.n1548 gnd.n1547 585
R9471 gnd.n1282 gnd.n1281 585
R9472 gnd.n1545 gnd.n1282 585
R9473 gnd.n1304 gnd.n1303 585
R9474 gnd.n1307 gnd.n1306 585
R9475 gnd.n1305 gnd.n1300 585
R9476 gnd.n1312 gnd.n1311 585
R9477 gnd.n1314 gnd.n1313 585
R9478 gnd.n1317 gnd.n1316 585
R9479 gnd.n1315 gnd.n1298 585
R9480 gnd.n1322 gnd.n1321 585
R9481 gnd.n1324 gnd.n1323 585
R9482 gnd.n1327 gnd.n1326 585
R9483 gnd.n1325 gnd.n1296 585
R9484 gnd.n1332 gnd.n1331 585
R9485 gnd.n1336 gnd.n1333 585
R9486 gnd.n1337 gnd.n1274 585
R9487 gnd.n2217 gnd.n905 585
R9488 gnd.n2284 gnd.n2283 585
R9489 gnd.n2286 gnd.n2285 585
R9490 gnd.n2288 gnd.n2287 585
R9491 gnd.n2290 gnd.n2289 585
R9492 gnd.n2292 gnd.n2291 585
R9493 gnd.n2294 gnd.n2293 585
R9494 gnd.n2296 gnd.n2295 585
R9495 gnd.n2298 gnd.n2297 585
R9496 gnd.n2300 gnd.n2299 585
R9497 gnd.n2302 gnd.n2301 585
R9498 gnd.n2304 gnd.n2303 585
R9499 gnd.n2306 gnd.n2305 585
R9500 gnd.n2309 gnd.n2308 585
R9501 gnd.n2307 gnd.n893 585
R9502 gnd.n2313 gnd.n891 585
R9503 gnd.n2315 gnd.n2314 585
R9504 gnd.n2316 gnd.n2315 585
R9505 gnd.n2218 gnd.n946 585
R9506 gnd.n2218 gnd.n867 585
R9507 gnd.n2220 gnd.n2219 585
R9508 gnd.n2219 gnd.n941 585
R9509 gnd.n2216 gnd.n945 585
R9510 gnd.n2216 gnd.n2215 585
R9511 gnd.n2195 gnd.n947 585
R9512 gnd.n959 gnd.n947 585
R9513 gnd.n2194 gnd.n957 585
R9514 gnd.n2203 gnd.n957 585
R9515 gnd.n1929 gnd.n964 585
R9516 gnd.n1930 gnd.n1929 585
R9517 gnd.n1928 gnd.n1927 585
R9518 gnd.n1928 gnd.n968 585
R9519 gnd.n1926 gnd.n970 585
R9520 gnd.n1919 gnd.n970 585
R9521 gnd.n983 gnd.n971 585
R9522 gnd.n983 gnd.n975 585
R9523 gnd.n1875 gnd.n984 585
R9524 gnd.n1909 gnd.n984 585
R9525 gnd.n1874 gnd.n1873 585
R9526 gnd.n1873 gnd.n991 585
R9527 gnd.n1872 gnd.n999 585
R9528 gnd.n1872 gnd.n990 585
R9529 gnd.n1871 gnd.n1001 585
R9530 gnd.n1871 gnd.n1870 585
R9531 gnd.n1850 gnd.n1000 585
R9532 gnd.n1013 gnd.n1000 585
R9533 gnd.n1849 gnd.n1011 585
R9534 gnd.n1860 gnd.n1011 585
R9535 gnd.n1840 gnd.n1018 585
R9536 gnd.n1841 gnd.n1840 585
R9537 gnd.n1839 gnd.n1838 585
R9538 gnd.n1839 gnd.n1022 585
R9539 gnd.n1837 gnd.n1024 585
R9540 gnd.n1830 gnd.n1024 585
R9541 gnd.n1817 gnd.n1025 585
R9542 gnd.n1818 gnd.n1817 585
R9543 gnd.n1788 gnd.n1038 585
R9544 gnd.n1820 gnd.n1038 585
R9545 gnd.n1787 gnd.n1786 585
R9546 gnd.n1786 gnd.n1045 585
R9547 gnd.n1785 gnd.n1052 585
R9548 gnd.n1785 gnd.n1044 585
R9549 gnd.n1784 gnd.n1054 585
R9550 gnd.n1784 gnd.n1783 585
R9551 gnd.n1763 gnd.n1053 585
R9552 gnd.n1066 gnd.n1053 585
R9553 gnd.n1762 gnd.n1064 585
R9554 gnd.n1773 gnd.n1064 585
R9555 gnd.n1753 gnd.n1071 585
R9556 gnd.n1754 gnd.n1753 585
R9557 gnd.n1752 gnd.n1751 585
R9558 gnd.n1752 gnd.n1075 585
R9559 gnd.n1750 gnd.n1077 585
R9560 gnd.n1743 gnd.n1077 585
R9561 gnd.n1730 gnd.n1078 585
R9562 gnd.n1731 gnd.n1730 585
R9563 gnd.n1683 gnd.n1091 585
R9564 gnd.n1733 gnd.n1091 585
R9565 gnd.n1685 gnd.n1684 585
R9566 gnd.n1686 gnd.n1685 585
R9567 gnd.n1678 gnd.n1181 585
R9568 gnd.n1181 gnd.n1180 585
R9569 gnd.n1676 gnd.n1675 585
R9570 gnd.n1675 gnd.n1162 585
R9571 gnd.n1673 gnd.n1160 585
R9572 gnd.n1694 gnd.n1160 585
R9573 gnd.n1191 gnd.n1190 585
R9574 gnd.n1190 gnd.n1189 585
R9575 gnd.n1667 gnd.n1150 585
R9576 gnd.n1700 gnd.n1150 585
R9577 gnd.n1666 gnd.n1665 585
R9578 gnd.n1665 gnd.n1664 585
R9579 gnd.n1662 gnd.n1193 585
R9580 gnd.n1662 gnd.n1140 585
R9581 gnd.n1661 gnd.n1660 585
R9582 gnd.n1661 gnd.n1139 585
R9583 gnd.n1196 gnd.n1195 585
R9584 gnd.n1652 gnd.n1195 585
R9585 gnd.n1620 gnd.n1619 585
R9586 gnd.n1619 gnd.n1200 585
R9587 gnd.n1621 gnd.n1209 585
R9588 gnd.n1638 gnd.n1209 585
R9589 gnd.n1618 gnd.n1617 585
R9590 gnd.n1617 gnd.n1215 585
R9591 gnd.n1616 gnd.n1223 585
R9592 gnd.n1616 gnd.n1615 585
R9593 gnd.n1601 gnd.n1224 585
R9594 gnd.n1234 gnd.n1224 585
R9595 gnd.n1600 gnd.n1232 585
R9596 gnd.n1607 gnd.n1232 585
R9597 gnd.n1599 gnd.n1598 585
R9598 gnd.n1598 gnd.n1597 585
R9599 gnd.n1243 gnd.n1240 585
R9600 gnd.n1253 gnd.n1243 585
R9601 gnd.n1589 gnd.n1588 585
R9602 gnd.n1588 gnd.n1587 585
R9603 gnd.n1249 gnd.n1248 585
R9604 gnd.n1262 gnd.n1249 585
R9605 gnd.n1569 gnd.n1260 585
R9606 gnd.n1577 gnd.n1260 585
R9607 gnd.n1568 gnd.n1567 585
R9608 gnd.n1567 gnd.n1566 585
R9609 gnd.n1269 gnd.n1267 585
R9610 gnd.n1278 gnd.n1269 585
R9611 gnd.n1558 gnd.n1557 585
R9612 gnd.n1557 gnd.n1556 585
R9613 gnd.n5928 gnd.n5927 585
R9614 gnd.n5927 gnd.n5926 585
R9615 gnd.n5929 gnd.n2528 585
R9616 gnd.n4541 gnd.n2528 585
R9617 gnd.n5931 gnd.n5930 585
R9618 gnd.n5932 gnd.n5931 585
R9619 gnd.n2512 gnd.n2511 585
R9620 gnd.n4430 gnd.n2512 585
R9621 gnd.n5940 gnd.n5939 585
R9622 gnd.n5939 gnd.n5938 585
R9623 gnd.n5941 gnd.n2506 585
R9624 gnd.n4421 gnd.n2506 585
R9625 gnd.n5943 gnd.n5942 585
R9626 gnd.n5944 gnd.n5943 585
R9627 gnd.n2491 gnd.n2490 585
R9628 gnd.n4441 gnd.n2491 585
R9629 gnd.n5952 gnd.n5951 585
R9630 gnd.n5951 gnd.n5950 585
R9631 gnd.n5953 gnd.n2485 585
R9632 gnd.n4413 gnd.n2485 585
R9633 gnd.n5955 gnd.n5954 585
R9634 gnd.n5956 gnd.n5955 585
R9635 gnd.n2470 gnd.n2469 585
R9636 gnd.n4405 gnd.n2470 585
R9637 gnd.n5964 gnd.n5963 585
R9638 gnd.n5963 gnd.n5962 585
R9639 gnd.n5965 gnd.n2464 585
R9640 gnd.n4397 gnd.n2464 585
R9641 gnd.n5967 gnd.n5966 585
R9642 gnd.n5968 gnd.n5967 585
R9643 gnd.n2449 gnd.n2448 585
R9644 gnd.n4389 gnd.n2449 585
R9645 gnd.n5976 gnd.n5975 585
R9646 gnd.n5975 gnd.n5974 585
R9647 gnd.n5977 gnd.n2446 585
R9648 gnd.n4339 gnd.n2446 585
R9649 gnd.n5980 gnd.n5979 585
R9650 gnd.n5981 gnd.n5980 585
R9651 gnd.n2447 gnd.n2432 585
R9652 gnd.n4327 gnd.n2432 585
R9653 gnd.n5989 gnd.n5988 585
R9654 gnd.n5988 gnd.n5987 585
R9655 gnd.n5990 gnd.n2429 585
R9656 gnd.n4312 gnd.n2429 585
R9657 gnd.n5993 gnd.n5992 585
R9658 gnd.n5994 gnd.n5993 585
R9659 gnd.n2430 gnd.n2414 585
R9660 gnd.n4352 gnd.n2414 585
R9661 gnd.n6002 gnd.n6001 585
R9662 gnd.n6001 gnd.n6000 585
R9663 gnd.n6003 gnd.n2410 585
R9664 gnd.n4304 gnd.n2410 585
R9665 gnd.n6006 gnd.n6005 585
R9666 gnd.n6007 gnd.n6006 585
R9667 gnd.n2394 gnd.n2393 585
R9668 gnd.n4295 gnd.n2394 585
R9669 gnd.n6015 gnd.n6014 585
R9670 gnd.n6014 gnd.n6013 585
R9671 gnd.n6016 gnd.n2388 585
R9672 gnd.n4286 gnd.n2388 585
R9673 gnd.n6018 gnd.n6017 585
R9674 gnd.n6019 gnd.n6018 585
R9675 gnd.n2373 gnd.n2372 585
R9676 gnd.n4278 gnd.n2373 585
R9677 gnd.n6027 gnd.n6026 585
R9678 gnd.n6026 gnd.n6025 585
R9679 gnd.n6028 gnd.n2367 585
R9680 gnd.n4223 gnd.n2367 585
R9681 gnd.n6030 gnd.n6029 585
R9682 gnd.n6031 gnd.n6030 585
R9683 gnd.n2351 gnd.n2350 585
R9684 gnd.n4229 gnd.n2351 585
R9685 gnd.n6039 gnd.n6038 585
R9686 gnd.n6038 gnd.n6037 585
R9687 gnd.n6040 gnd.n2345 585
R9688 gnd.n4235 gnd.n2345 585
R9689 gnd.n6042 gnd.n6041 585
R9690 gnd.n6043 gnd.n6042 585
R9691 gnd.n2329 gnd.n2328 585
R9692 gnd.n4241 gnd.n2329 585
R9693 gnd.n6051 gnd.n6050 585
R9694 gnd.n6050 gnd.n6049 585
R9695 gnd.n6052 gnd.n2324 585
R9696 gnd.n4247 gnd.n2324 585
R9697 gnd.n6054 gnd.n6053 585
R9698 gnd.n6055 gnd.n6054 585
R9699 gnd.n4100 gnd.n2323 585
R9700 gnd.n4103 gnd.n4102 585
R9701 gnd.n4098 gnd.n4097 585
R9702 gnd.n4097 gnd.n2318 585
R9703 gnd.n4108 gnd.n4107 585
R9704 gnd.n4110 gnd.n4096 585
R9705 gnd.n4113 gnd.n4112 585
R9706 gnd.n4094 gnd.n4093 585
R9707 gnd.n4118 gnd.n4117 585
R9708 gnd.n4120 gnd.n4092 585
R9709 gnd.n4123 gnd.n4122 585
R9710 gnd.n4090 gnd.n4089 585
R9711 gnd.n4128 gnd.n4127 585
R9712 gnd.n4130 gnd.n4088 585
R9713 gnd.n4133 gnd.n4132 585
R9714 gnd.n4086 gnd.n4085 585
R9715 gnd.n4138 gnd.n4137 585
R9716 gnd.n4140 gnd.n4081 585
R9717 gnd.n4143 gnd.n4142 585
R9718 gnd.n4079 gnd.n4078 585
R9719 gnd.n4148 gnd.n4147 585
R9720 gnd.n4150 gnd.n4077 585
R9721 gnd.n4153 gnd.n4152 585
R9722 gnd.n4075 gnd.n4074 585
R9723 gnd.n4158 gnd.n4157 585
R9724 gnd.n4160 gnd.n4073 585
R9725 gnd.n4163 gnd.n4162 585
R9726 gnd.n4071 gnd.n4070 585
R9727 gnd.n4168 gnd.n4167 585
R9728 gnd.n4170 gnd.n4069 585
R9729 gnd.n4173 gnd.n4172 585
R9730 gnd.n4067 gnd.n4066 585
R9731 gnd.n4178 gnd.n4177 585
R9732 gnd.n4180 gnd.n4065 585
R9733 gnd.n4183 gnd.n4182 585
R9734 gnd.n4063 gnd.n4062 585
R9735 gnd.n4189 gnd.n4188 585
R9736 gnd.n4191 gnd.n4061 585
R9737 gnd.n4192 gnd.n4060 585
R9738 gnd.n4195 gnd.n4194 585
R9739 gnd.n4548 gnd.n4547 585
R9740 gnd.n4550 gnd.n3710 585
R9741 gnd.n4552 gnd.n4551 585
R9742 gnd.n4553 gnd.n3703 585
R9743 gnd.n4555 gnd.n4554 585
R9744 gnd.n4557 gnd.n3701 585
R9745 gnd.n4559 gnd.n4558 585
R9746 gnd.n4560 gnd.n3696 585
R9747 gnd.n4562 gnd.n4561 585
R9748 gnd.n4564 gnd.n3694 585
R9749 gnd.n4566 gnd.n4565 585
R9750 gnd.n4567 gnd.n3689 585
R9751 gnd.n4569 gnd.n4568 585
R9752 gnd.n4571 gnd.n3687 585
R9753 gnd.n4573 gnd.n4572 585
R9754 gnd.n4574 gnd.n3682 585
R9755 gnd.n4576 gnd.n4575 585
R9756 gnd.n4578 gnd.n3681 585
R9757 gnd.n4579 gnd.n3624 585
R9758 gnd.n4582 gnd.n4581 585
R9759 gnd.n3625 gnd.n3617 585
R9760 gnd.n3653 gnd.n3618 585
R9761 gnd.n3655 gnd.n3654 585
R9762 gnd.n3657 gnd.n3656 585
R9763 gnd.n3659 gnd.n3658 585
R9764 gnd.n3661 gnd.n3660 585
R9765 gnd.n3663 gnd.n3662 585
R9766 gnd.n3665 gnd.n3664 585
R9767 gnd.n3667 gnd.n3666 585
R9768 gnd.n3669 gnd.n3668 585
R9769 gnd.n3671 gnd.n3670 585
R9770 gnd.n3673 gnd.n3672 585
R9771 gnd.n3675 gnd.n3674 585
R9772 gnd.n3676 gnd.n3635 585
R9773 gnd.n3678 gnd.n3677 585
R9774 gnd.n3636 gnd.n3634 585
R9775 gnd.n3637 gnd.n2533 585
R9776 gnd.n3680 gnd.n2533 585
R9777 gnd.n4544 gnd.n2535 585
R9778 gnd.n5926 gnd.n2535 585
R9779 gnd.n4543 gnd.n4542 585
R9780 gnd.n4542 gnd.n4541 585
R9781 gnd.n3714 gnd.n2525 585
R9782 gnd.n5932 gnd.n2525 585
R9783 gnd.n4429 gnd.n4428 585
R9784 gnd.n4430 gnd.n4429 585
R9785 gnd.n3911 gnd.n2514 585
R9786 gnd.n5938 gnd.n2514 585
R9787 gnd.n4423 gnd.n4422 585
R9788 gnd.n4422 gnd.n4421 585
R9789 gnd.n4420 gnd.n2503 585
R9790 gnd.n5944 gnd.n2503 585
R9791 gnd.n4419 gnd.n3905 585
R9792 gnd.n4441 gnd.n3905 585
R9793 gnd.n3913 gnd.n2493 585
R9794 gnd.n5950 gnd.n2493 585
R9795 gnd.n4415 gnd.n4414 585
R9796 gnd.n4414 gnd.n4413 585
R9797 gnd.n3915 gnd.n2482 585
R9798 gnd.n5956 gnd.n2482 585
R9799 gnd.n4404 gnd.n4403 585
R9800 gnd.n4405 gnd.n4404 585
R9801 gnd.n3920 gnd.n2472 585
R9802 gnd.n5962 gnd.n2472 585
R9803 gnd.n4399 gnd.n4398 585
R9804 gnd.n4398 gnd.n4397 585
R9805 gnd.n3922 gnd.n2461 585
R9806 gnd.n5968 gnd.n2461 585
R9807 gnd.n4335 gnd.n3926 585
R9808 gnd.n4389 gnd.n3926 585
R9809 gnd.n4336 gnd.n2451 585
R9810 gnd.n5974 gnd.n2451 585
R9811 gnd.n4338 gnd.n4337 585
R9812 gnd.n4339 gnd.n4338 585
R9813 gnd.n3950 gnd.n2443 585
R9814 gnd.n5981 gnd.n2443 585
R9815 gnd.n4329 gnd.n4328 585
R9816 gnd.n4328 gnd.n4327 585
R9817 gnd.n4315 gnd.n2434 585
R9818 gnd.n5987 gnd.n2434 585
R9819 gnd.n4314 gnd.n4313 585
R9820 gnd.n4313 gnd.n4312 585
R9821 gnd.n3952 gnd.n2426 585
R9822 gnd.n5994 gnd.n2426 585
R9823 gnd.n4308 gnd.n3942 585
R9824 gnd.n4352 gnd.n3942 585
R9825 gnd.n4307 gnd.n2416 585
R9826 gnd.n6000 gnd.n2416 585
R9827 gnd.n4306 gnd.n4305 585
R9828 gnd.n4305 gnd.n4304 585
R9829 gnd.n3955 gnd.n2407 585
R9830 gnd.n6007 gnd.n2407 585
R9831 gnd.n4294 gnd.n4293 585
R9832 gnd.n4295 gnd.n4294 585
R9833 gnd.n3960 gnd.n2396 585
R9834 gnd.n6013 gnd.n2396 585
R9835 gnd.n4288 gnd.n4287 585
R9836 gnd.n4287 gnd.n4286 585
R9837 gnd.n3962 gnd.n2385 585
R9838 gnd.n6019 gnd.n2385 585
R9839 gnd.n4217 gnd.n3966 585
R9840 gnd.n4278 gnd.n3966 585
R9841 gnd.n4218 gnd.n2375 585
R9842 gnd.n6025 gnd.n2375 585
R9843 gnd.n4225 gnd.n4224 585
R9844 gnd.n4224 gnd.n4223 585
R9845 gnd.n4226 gnd.n2364 585
R9846 gnd.n6031 gnd.n2364 585
R9847 gnd.n4228 gnd.n4227 585
R9848 gnd.n4229 gnd.n4228 585
R9849 gnd.n4205 gnd.n2353 585
R9850 gnd.n6037 gnd.n2353 585
R9851 gnd.n4237 gnd.n4236 585
R9852 gnd.n4236 gnd.n4235 585
R9853 gnd.n4238 gnd.n2342 585
R9854 gnd.n6043 gnd.n2342 585
R9855 gnd.n4240 gnd.n4239 585
R9856 gnd.n4241 gnd.n4240 585
R9857 gnd.n4056 gnd.n2330 585
R9858 gnd.n6049 gnd.n2330 585
R9859 gnd.n4199 gnd.n3978 585
R9860 gnd.n4247 gnd.n3978 585
R9861 gnd.n4198 gnd.n2319 585
R9862 gnd.n6055 gnd.n2319 585
R9863 gnd.n7192 gnd.n7191 585
R9864 gnd.n7193 gnd.n7192 585
R9865 gnd.n87 gnd.n85 585
R9866 gnd.n7114 gnd.n85 585
R9867 gnd.n7036 gnd.n174 585
R9868 gnd.n174 gnd.n173 585
R9869 gnd.n7038 gnd.n7037 585
R9870 gnd.n7039 gnd.n7038 585
R9871 gnd.n175 gnd.n172 585
R9872 gnd.n6926 gnd.n172 585
R9873 gnd.n7031 gnd.n7030 585
R9874 gnd.n7030 gnd.n7029 585
R9875 gnd.n178 gnd.n177 585
R9876 gnd.n6932 gnd.n178 585
R9877 gnd.n7020 gnd.n7019 585
R9878 gnd.n7021 gnd.n7020 585
R9879 gnd.n191 gnd.n190 585
R9880 gnd.n6915 gnd.n190 585
R9881 gnd.n7015 gnd.n7014 585
R9882 gnd.n7014 gnd.n7013 585
R9883 gnd.n194 gnd.n193 585
R9884 gnd.n6941 gnd.n194 585
R9885 gnd.n7004 gnd.n7003 585
R9886 gnd.n7005 gnd.n7004 585
R9887 gnd.n207 gnd.n206 585
R9888 gnd.n6945 gnd.n206 585
R9889 gnd.n6999 gnd.n6998 585
R9890 gnd.n6998 gnd.n6997 585
R9891 gnd.n210 gnd.n209 585
R9892 gnd.n6951 gnd.n210 585
R9893 gnd.n6988 gnd.n6987 585
R9894 gnd.n6989 gnd.n6988 585
R9895 gnd.n223 gnd.n222 585
R9896 gnd.n5700 gnd.n222 585
R9897 gnd.n6964 gnd.n6963 585
R9898 gnd.n6965 gnd.n6964 585
R9899 gnd.n6962 gnd.n254 585
R9900 gnd.n6962 gnd.n6961 585
R9901 gnd.n253 gnd.n252 585
R9902 gnd.n5708 gnd.n252 585
R9903 gnd.n2723 gnd.n2722 585
R9904 gnd.n2726 gnd.n2722 585
R9905 gnd.n5728 gnd.n2724 585
R9906 gnd.n5728 gnd.n5727 585
R9907 gnd.n5731 gnd.n5730 585
R9908 gnd.n5732 gnd.n5731 585
R9909 gnd.n5729 gnd.n232 585
R9910 gnd.n5716 gnd.n232 585
R9911 gnd.n6982 gnd.n6981 585
R9912 gnd.n6981 gnd.n6980 585
R9913 gnd.n6983 gnd.n231 585
R9914 gnd.n5686 gnd.n231 585
R9915 gnd.n5746 gnd.n230 585
R9916 gnd.n5747 gnd.n5746 585
R9917 gnd.n5745 gnd.n2709 585
R9918 gnd.n5745 gnd.n5744 585
R9919 gnd.n5675 gnd.n2708 585
R9920 gnd.n2740 gnd.n2708 585
R9921 gnd.n5677 gnd.n5676 585
R9922 gnd.n5678 gnd.n5677 585
R9923 gnd.n2743 gnd.n2742 585
R9924 gnd.n5631 gnd.n2742 585
R9925 gnd.n5670 gnd.n5669 585
R9926 gnd.n5669 gnd.n5668 585
R9927 gnd.n2746 gnd.n2745 585
R9928 gnd.n5640 gnd.n2746 585
R9929 gnd.n5622 gnd.n2767 585
R9930 gnd.n5582 gnd.n2767 585
R9931 gnd.n5624 gnd.n5623 585
R9932 gnd.n5625 gnd.n5624 585
R9933 gnd.n2768 gnd.n2766 585
R9934 gnd.n2776 gnd.n2766 585
R9935 gnd.n5617 gnd.n5616 585
R9936 gnd.n5616 gnd.n5615 585
R9937 gnd.n2771 gnd.n2770 585
R9938 gnd.n5603 gnd.n2771 585
R9939 gnd.n2793 gnd.n2792 585
R9940 gnd.n2794 gnd.n2793 585
R9941 gnd.n2678 gnd.n2677 585
R9942 gnd.n5594 gnd.n2678 585
R9943 gnd.n5775 gnd.n5774 585
R9944 gnd.n5774 gnd.n5773 585
R9945 gnd.n5776 gnd.n2673 585
R9946 gnd.n5566 gnd.n2673 585
R9947 gnd.n5778 gnd.n5777 585
R9948 gnd.n5779 gnd.n5778 585
R9949 gnd.n3030 gnd.n2672 585
R9950 gnd.n3033 gnd.n3032 585
R9951 gnd.n3028 gnd.n3027 585
R9952 gnd.n3027 gnd.n2659 585
R9953 gnd.n3038 gnd.n3037 585
R9954 gnd.n3040 gnd.n3026 585
R9955 gnd.n3043 gnd.n3042 585
R9956 gnd.n3024 gnd.n3023 585
R9957 gnd.n3048 gnd.n3047 585
R9958 gnd.n3050 gnd.n3022 585
R9959 gnd.n3053 gnd.n3052 585
R9960 gnd.n3020 gnd.n3019 585
R9961 gnd.n3059 gnd.n3058 585
R9962 gnd.n3061 gnd.n3018 585
R9963 gnd.n3062 gnd.n3015 585
R9964 gnd.n3065 gnd.n3064 585
R9965 gnd.n3017 gnd.n3012 585
R9966 gnd.n3146 gnd.n3145 585
R9967 gnd.n3143 gnd.n3072 585
R9968 gnd.n3141 gnd.n3140 585
R9969 gnd.n3139 gnd.n3073 585
R9970 gnd.n3138 gnd.n3137 585
R9971 gnd.n3135 gnd.n3078 585
R9972 gnd.n3133 gnd.n3132 585
R9973 gnd.n3131 gnd.n3079 585
R9974 gnd.n3130 gnd.n3129 585
R9975 gnd.n3127 gnd.n3084 585
R9976 gnd.n3125 gnd.n3124 585
R9977 gnd.n3123 gnd.n3085 585
R9978 gnd.n3122 gnd.n3121 585
R9979 gnd.n3119 gnd.n3090 585
R9980 gnd.n3117 gnd.n3116 585
R9981 gnd.n3115 gnd.n3091 585
R9982 gnd.n3114 gnd.n3113 585
R9983 gnd.n3111 gnd.n3096 585
R9984 gnd.n3109 gnd.n3108 585
R9985 gnd.n3100 gnd.n3097 585
R9986 gnd.n3104 gnd.n3103 585
R9987 gnd.n156 gnd.n155 585
R9988 gnd.n7121 gnd.n151 585
R9989 gnd.n7123 gnd.n7122 585
R9990 gnd.n7125 gnd.n149 585
R9991 gnd.n7127 gnd.n7126 585
R9992 gnd.n7128 gnd.n144 585
R9993 gnd.n7130 gnd.n7129 585
R9994 gnd.n7132 gnd.n142 585
R9995 gnd.n7134 gnd.n7133 585
R9996 gnd.n7135 gnd.n137 585
R9997 gnd.n7137 gnd.n7136 585
R9998 gnd.n7139 gnd.n135 585
R9999 gnd.n7141 gnd.n7140 585
R10000 gnd.n7142 gnd.n130 585
R10001 gnd.n7144 gnd.n7143 585
R10002 gnd.n7146 gnd.n128 585
R10003 gnd.n7148 gnd.n7147 585
R10004 gnd.n7149 gnd.n123 585
R10005 gnd.n7151 gnd.n7150 585
R10006 gnd.n7153 gnd.n121 585
R10007 gnd.n7155 gnd.n7154 585
R10008 gnd.n7159 gnd.n116 585
R10009 gnd.n7161 gnd.n7160 585
R10010 gnd.n7163 gnd.n114 585
R10011 gnd.n7165 gnd.n7164 585
R10012 gnd.n7166 gnd.n109 585
R10013 gnd.n7168 gnd.n7167 585
R10014 gnd.n7170 gnd.n107 585
R10015 gnd.n7172 gnd.n7171 585
R10016 gnd.n7173 gnd.n102 585
R10017 gnd.n7175 gnd.n7174 585
R10018 gnd.n7177 gnd.n100 585
R10019 gnd.n7179 gnd.n7178 585
R10020 gnd.n7180 gnd.n95 585
R10021 gnd.n7182 gnd.n7181 585
R10022 gnd.n7184 gnd.n92 585
R10023 gnd.n7186 gnd.n7185 585
R10024 gnd.n7187 gnd.n90 585
R10025 gnd.n7188 gnd.n86 585
R10026 gnd.n94 gnd.n86 585
R10027 gnd.n7117 gnd.n82 585
R10028 gnd.n7193 gnd.n82 585
R10029 gnd.n7116 gnd.n7115 585
R10030 gnd.n7115 gnd.n7114 585
R10031 gnd.n161 gnd.n160 585
R10032 gnd.n173 gnd.n161 585
R10033 gnd.n6925 gnd.n170 585
R10034 gnd.n7039 gnd.n170 585
R10035 gnd.n6928 gnd.n6927 585
R10036 gnd.n6927 gnd.n6926 585
R10037 gnd.n6929 gnd.n180 585
R10038 gnd.n7029 gnd.n180 585
R10039 gnd.n6931 gnd.n6930 585
R10040 gnd.n6932 gnd.n6931 585
R10041 gnd.n6913 gnd.n189 585
R10042 gnd.n7021 gnd.n189 585
R10043 gnd.n6917 gnd.n6916 585
R10044 gnd.n6916 gnd.n6915 585
R10045 gnd.n269 gnd.n195 585
R10046 gnd.n7013 gnd.n195 585
R10047 gnd.n6943 gnd.n6942 585
R10048 gnd.n6942 gnd.n6941 585
R10049 gnd.n6944 gnd.n204 585
R10050 gnd.n7005 gnd.n204 585
R10051 gnd.n6947 gnd.n6946 585
R10052 gnd.n6946 gnd.n6945 585
R10053 gnd.n6948 gnd.n212 585
R10054 gnd.n6997 gnd.n212 585
R10055 gnd.n6950 gnd.n6949 585
R10056 gnd.n6951 gnd.n6950 585
R10057 gnd.n263 gnd.n221 585
R10058 gnd.n6989 gnd.n221 585
R10059 gnd.n5702 gnd.n5701 585
R10060 gnd.n5701 gnd.n5700 585
R10061 gnd.n5703 gnd.n249 585
R10062 gnd.n6965 gnd.n249 585
R10063 gnd.n5704 gnd.n256 585
R10064 gnd.n6961 gnd.n256 585
R10065 gnd.n5709 gnd.n5705 585
R10066 gnd.n5709 gnd.n5708 585
R10067 gnd.n5711 gnd.n5710 585
R10068 gnd.n5710 gnd.n2726 585
R10069 gnd.n5712 gnd.n2725 585
R10070 gnd.n5727 gnd.n2725 585
R10071 gnd.n5713 gnd.n2720 585
R10072 gnd.n5732 gnd.n2720 585
R10073 gnd.n5715 gnd.n5714 585
R10074 gnd.n5716 gnd.n5715 585
R10075 gnd.n2731 gnd.n234 585
R10076 gnd.n6980 gnd.n234 585
R10077 gnd.n5688 gnd.n5687 585
R10078 gnd.n5687 gnd.n5686 585
R10079 gnd.n5685 gnd.n2705 585
R10080 gnd.n5747 gnd.n2705 585
R10081 gnd.n5684 gnd.n2711 585
R10082 gnd.n5744 gnd.n2711 585
R10083 gnd.n2737 gnd.n2733 585
R10084 gnd.n2740 gnd.n2737 585
R10085 gnd.n5680 gnd.n5679 585
R10086 gnd.n5679 gnd.n5678 585
R10087 gnd.n2736 gnd.n2735 585
R10088 gnd.n5631 gnd.n2736 585
R10089 gnd.n5580 gnd.n2748 585
R10090 gnd.n5668 gnd.n2748 585
R10091 gnd.n5581 gnd.n2756 585
R10092 gnd.n5640 gnd.n2756 585
R10093 gnd.n5584 gnd.n5583 585
R10094 gnd.n5583 gnd.n5582 585
R10095 gnd.n5585 gnd.n2764 585
R10096 gnd.n5625 gnd.n2764 585
R10097 gnd.n5587 gnd.n5586 585
R10098 gnd.n5586 gnd.n2776 585
R10099 gnd.n5588 gnd.n2773 585
R10100 gnd.n5615 gnd.n2773 585
R10101 gnd.n5589 gnd.n2795 585
R10102 gnd.n5603 gnd.n2795 585
R10103 gnd.n5590 gnd.n2801 585
R10104 gnd.n2801 gnd.n2794 585
R10105 gnd.n5592 gnd.n5591 585
R10106 gnd.n5594 gnd.n5592 585
R10107 gnd.n2802 gnd.n2680 585
R10108 gnd.n5773 gnd.n2680 585
R10109 gnd.n5568 gnd.n5567 585
R10110 gnd.n5567 gnd.n5566 585
R10111 gnd.n2804 gnd.n2668 585
R10112 gnd.n5779 gnd.n2668 585
R10113 gnd.n5430 gnd.n5429 585
R10114 gnd.n5431 gnd.n5430 585
R10115 gnd.n5341 gnd.n3154 585
R10116 gnd.n3160 gnd.n3154 585
R10117 gnd.n5340 gnd.n5339 585
R10118 gnd.n5339 gnd.n5338 585
R10119 gnd.n3157 gnd.n3156 585
R10120 gnd.n5256 gnd.n3157 585
R10121 gnd.n5327 gnd.n5326 585
R10122 gnd.n5328 gnd.n5327 585
R10123 gnd.n5325 gnd.n3170 585
R10124 gnd.n3170 gnd.n3166 585
R10125 gnd.n5324 gnd.n5323 585
R10126 gnd.n5323 gnd.n5322 585
R10127 gnd.n3172 gnd.n3171 585
R10128 gnd.n5265 gnd.n3172 585
R10129 gnd.n5294 gnd.n5293 585
R10130 gnd.n5295 gnd.n5294 585
R10131 gnd.n5292 gnd.n3184 585
R10132 gnd.n3184 gnd.n3182 585
R10133 gnd.n5291 gnd.n5290 585
R10134 gnd.n5290 gnd.n5289 585
R10135 gnd.n3186 gnd.n3185 585
R10136 gnd.n5274 gnd.n3186 585
R10137 gnd.n5246 gnd.n3203 585
R10138 gnd.n3203 gnd.n3195 585
R10139 gnd.n5248 gnd.n5247 585
R10140 gnd.n5249 gnd.n5248 585
R10141 gnd.n5245 gnd.n3202 585
R10142 gnd.n3208 gnd.n3202 585
R10143 gnd.n5244 gnd.n5243 585
R10144 gnd.n5243 gnd.n5242 585
R10145 gnd.n3205 gnd.n3204 585
R10146 gnd.n5154 gnd.n3205 585
R10147 gnd.n5230 gnd.n5229 585
R10148 gnd.n5231 gnd.n5230 585
R10149 gnd.n5228 gnd.n3219 585
R10150 gnd.n3219 gnd.n3215 585
R10151 gnd.n5227 gnd.n5226 585
R10152 gnd.n5226 gnd.n5225 585
R10153 gnd.n3221 gnd.n3220 585
R10154 gnd.n5163 gnd.n3221 585
R10155 gnd.n5201 gnd.n5200 585
R10156 gnd.n5202 gnd.n5201 585
R10157 gnd.n5199 gnd.n3232 585
R10158 gnd.n3232 gnd.n3229 585
R10159 gnd.n5198 gnd.n5197 585
R10160 gnd.n5197 gnd.n5196 585
R10161 gnd.n3234 gnd.n3233 585
R10162 gnd.n5170 gnd.n3234 585
R10163 gnd.n5183 gnd.n5182 585
R10164 gnd.n5184 gnd.n5183 585
R10165 gnd.n5181 gnd.n3246 585
R10166 gnd.n5176 gnd.n3246 585
R10167 gnd.n5180 gnd.n5179 585
R10168 gnd.n5179 gnd.n5178 585
R10169 gnd.n3248 gnd.n3247 585
R10170 gnd.n5149 gnd.n3248 585
R10171 gnd.n5135 gnd.n5134 585
R10172 gnd.n5134 gnd.n5133 585
R10173 gnd.n5136 gnd.n3264 585
R10174 gnd.n5131 gnd.n3264 585
R10175 gnd.n5138 gnd.n5137 585
R10176 gnd.n5139 gnd.n5138 585
R10177 gnd.n3265 gnd.n3263 585
R10178 gnd.n5125 gnd.n3263 585
R10179 gnd.n5122 gnd.n5121 585
R10180 gnd.n5123 gnd.n5122 585
R10181 gnd.n5120 gnd.n3270 585
R10182 gnd.n3276 gnd.n3270 585
R10183 gnd.n5119 gnd.n5118 585
R10184 gnd.n5118 gnd.n5117 585
R10185 gnd.n3272 gnd.n3271 585
R10186 gnd.n5105 gnd.n3272 585
R10187 gnd.n5093 gnd.n3289 585
R10188 gnd.n3289 gnd.n3282 585
R10189 gnd.n5095 gnd.n5094 585
R10190 gnd.n5096 gnd.n5095 585
R10191 gnd.n5092 gnd.n3288 585
R10192 gnd.n3294 gnd.n3288 585
R10193 gnd.n5091 gnd.n5090 585
R10194 gnd.n5090 gnd.n5089 585
R10195 gnd.n3291 gnd.n3290 585
R10196 gnd.n4978 gnd.n3291 585
R10197 gnd.n5077 gnd.n5076 585
R10198 gnd.n5078 gnd.n5077 585
R10199 gnd.n5075 gnd.n3306 585
R10200 gnd.n3306 gnd.n3302 585
R10201 gnd.n5074 gnd.n5073 585
R10202 gnd.n5073 gnd.n5072 585
R10203 gnd.n3308 gnd.n3307 585
R10204 gnd.n4987 gnd.n3308 585
R10205 gnd.n5025 gnd.n5024 585
R10206 gnd.n5026 gnd.n5025 585
R10207 gnd.n5023 gnd.n3320 585
R10208 gnd.n3320 gnd.n3317 585
R10209 gnd.n5022 gnd.n5021 585
R10210 gnd.n5021 gnd.n5020 585
R10211 gnd.n3322 gnd.n3321 585
R10212 gnd.n4994 gnd.n3322 585
R10213 gnd.n5007 gnd.n5006 585
R10214 gnd.n5008 gnd.n5007 585
R10215 gnd.n5005 gnd.n3335 585
R10216 gnd.n5000 gnd.n3335 585
R10217 gnd.n5004 gnd.n5003 585
R10218 gnd.n5003 gnd.n5002 585
R10219 gnd.n3337 gnd.n3336 585
R10220 gnd.n4973 gnd.n3337 585
R10221 gnd.n4959 gnd.n4958 585
R10222 gnd.n4958 gnd.n4957 585
R10223 gnd.n4960 gnd.n3353 585
R10224 gnd.n4955 gnd.n3353 585
R10225 gnd.n4962 gnd.n4961 585
R10226 gnd.n4963 gnd.n4962 585
R10227 gnd.n3354 gnd.n3352 585
R10228 gnd.n4949 gnd.n3352 585
R10229 gnd.n4946 gnd.n4945 585
R10230 gnd.n4947 gnd.n4946 585
R10231 gnd.n4944 gnd.n3357 585
R10232 gnd.n3363 gnd.n3357 585
R10233 gnd.n4943 gnd.n4942 585
R10234 gnd.n4942 gnd.n4941 585
R10235 gnd.n3359 gnd.n3358 585
R10236 gnd.n4929 gnd.n3359 585
R10237 gnd.n4917 gnd.n3378 585
R10238 gnd.n3378 gnd.n3369 585
R10239 gnd.n4919 gnd.n4918 585
R10240 gnd.n4920 gnd.n4919 585
R10241 gnd.n4916 gnd.n3377 585
R10242 gnd.n3383 gnd.n3377 585
R10243 gnd.n4915 gnd.n4914 585
R10244 gnd.n4914 gnd.n4913 585
R10245 gnd.n3380 gnd.n3379 585
R10246 gnd.n4801 gnd.n3380 585
R10247 gnd.n4901 gnd.n4900 585
R10248 gnd.n4902 gnd.n4901 585
R10249 gnd.n4899 gnd.n3394 585
R10250 gnd.n3394 gnd.n3390 585
R10251 gnd.n4898 gnd.n4897 585
R10252 gnd.n4897 gnd.n4896 585
R10253 gnd.n3396 gnd.n3395 585
R10254 gnd.n4809 gnd.n3396 585
R10255 gnd.n4848 gnd.n4847 585
R10256 gnd.n4849 gnd.n4848 585
R10257 gnd.n4846 gnd.n3407 585
R10258 gnd.n3411 gnd.n3407 585
R10259 gnd.n4845 gnd.n4844 585
R10260 gnd.n4844 gnd.n4843 585
R10261 gnd.n3409 gnd.n3408 585
R10262 gnd.n4817 gnd.n3409 585
R10263 gnd.n4830 gnd.n4829 585
R10264 gnd.n4831 gnd.n4830 585
R10265 gnd.n4828 gnd.n3422 585
R10266 gnd.n4823 gnd.n3422 585
R10267 gnd.n4827 gnd.n4826 585
R10268 gnd.n4826 gnd.n4825 585
R10269 gnd.n3424 gnd.n3423 585
R10270 gnd.n4796 gnd.n3424 585
R10271 gnd.n4782 gnd.n4781 585
R10272 gnd.n4781 gnd.n4780 585
R10273 gnd.n4783 gnd.n3438 585
R10274 gnd.n4729 gnd.n3438 585
R10275 gnd.n4785 gnd.n4784 585
R10276 gnd.n4786 gnd.n4785 585
R10277 gnd.n3439 gnd.n3437 585
R10278 gnd.n4733 gnd.n3437 585
R10279 gnd.n4761 gnd.n4760 585
R10280 gnd.n4762 gnd.n4761 585
R10281 gnd.n4759 gnd.n3450 585
R10282 gnd.n3454 gnd.n3450 585
R10283 gnd.n4758 gnd.n4757 585
R10284 gnd.n4757 gnd.n4756 585
R10285 gnd.n3452 gnd.n3451 585
R10286 gnd.n4743 gnd.n3452 585
R10287 gnd.n4722 gnd.n3468 585
R10288 gnd.n3468 gnd.n3460 585
R10289 gnd.n4724 gnd.n4723 585
R10290 gnd.n4725 gnd.n4724 585
R10291 gnd.n4721 gnd.n3467 585
R10292 gnd.n3473 gnd.n3467 585
R10293 gnd.n4720 gnd.n4719 585
R10294 gnd.n4719 gnd.n4718 585
R10295 gnd.n3470 gnd.n3469 585
R10296 gnd.n4653 gnd.n3470 585
R10297 gnd.n4705 gnd.n4704 585
R10298 gnd.n4706 gnd.n4705 585
R10299 gnd.n4703 gnd.n3483 585
R10300 gnd.n3483 gnd.n3480 585
R10301 gnd.n4702 gnd.n4701 585
R10302 gnd.n4701 gnd.n4700 585
R10303 gnd.n3485 gnd.n3484 585
R10304 gnd.n4661 gnd.n3485 585
R10305 gnd.n4675 gnd.n4674 585
R10306 gnd.n4676 gnd.n4675 585
R10307 gnd.n4672 gnd.n3497 585
R10308 gnd.n4671 gnd.n4670 585
R10309 gnd.n3519 gnd.n3518 585
R10310 gnd.n4668 gnd.n3519 585
R10311 gnd.n3560 gnd.n3559 585
R10312 gnd.n3562 gnd.n3561 585
R10313 gnd.n3564 gnd.n3563 585
R10314 gnd.n3566 gnd.n3565 585
R10315 gnd.n3568 gnd.n3567 585
R10316 gnd.n3570 gnd.n3569 585
R10317 gnd.n3572 gnd.n3571 585
R10318 gnd.n3574 gnd.n3573 585
R10319 gnd.n3576 gnd.n3575 585
R10320 gnd.n3578 gnd.n3577 585
R10321 gnd.n3580 gnd.n3579 585
R10322 gnd.n3582 gnd.n3581 585
R10323 gnd.n3584 gnd.n3583 585
R10324 gnd.n3586 gnd.n3585 585
R10325 gnd.n3588 gnd.n3587 585
R10326 gnd.n3590 gnd.n3589 585
R10327 gnd.n3592 gnd.n3591 585
R10328 gnd.n3594 gnd.n3593 585
R10329 gnd.n3596 gnd.n3595 585
R10330 gnd.n3598 gnd.n3597 585
R10331 gnd.n3600 gnd.n3599 585
R10332 gnd.n3602 gnd.n3601 585
R10333 gnd.n3604 gnd.n3603 585
R10334 gnd.n3606 gnd.n3605 585
R10335 gnd.n3608 gnd.n3607 585
R10336 gnd.n3610 gnd.n3609 585
R10337 gnd.n3612 gnd.n3611 585
R10338 gnd.n3614 gnd.n3613 585
R10339 gnd.n3616 gnd.n3615 585
R10340 gnd.n4589 gnd.n4588 585
R10341 gnd.n4591 gnd.n4590 585
R10342 gnd.n4593 gnd.n4592 585
R10343 gnd.n4595 gnd.n4594 585
R10344 gnd.n4598 gnd.n4597 585
R10345 gnd.n4600 gnd.n4599 585
R10346 gnd.n4602 gnd.n4601 585
R10347 gnd.n4604 gnd.n4603 585
R10348 gnd.n4606 gnd.n4605 585
R10349 gnd.n4608 gnd.n4607 585
R10350 gnd.n4610 gnd.n4609 585
R10351 gnd.n4612 gnd.n4611 585
R10352 gnd.n4614 gnd.n4613 585
R10353 gnd.n4616 gnd.n4615 585
R10354 gnd.n4618 gnd.n4617 585
R10355 gnd.n4620 gnd.n4619 585
R10356 gnd.n4622 gnd.n4621 585
R10357 gnd.n4624 gnd.n4623 585
R10358 gnd.n4626 gnd.n4625 585
R10359 gnd.n4628 gnd.n4627 585
R10360 gnd.n4630 gnd.n4629 585
R10361 gnd.n4632 gnd.n4631 585
R10362 gnd.n4634 gnd.n4633 585
R10363 gnd.n4636 gnd.n4635 585
R10364 gnd.n4638 gnd.n4637 585
R10365 gnd.n4640 gnd.n4639 585
R10366 gnd.n4642 gnd.n4641 585
R10367 gnd.n4644 gnd.n4643 585
R10368 gnd.n4646 gnd.n4645 585
R10369 gnd.n4648 gnd.n4647 585
R10370 gnd.n4650 gnd.n4649 585
R10371 gnd.n4651 gnd.n3553 585
R10372 gnd.n4666 gnd.n4665 585
R10373 gnd.n5434 gnd.n5433 585
R10374 gnd.n5436 gnd.n5435 585
R10375 gnd.n5438 gnd.n5437 585
R10376 gnd.n5440 gnd.n5439 585
R10377 gnd.n5442 gnd.n5441 585
R10378 gnd.n5444 gnd.n5443 585
R10379 gnd.n5446 gnd.n5445 585
R10380 gnd.n5448 gnd.n5447 585
R10381 gnd.n5450 gnd.n5449 585
R10382 gnd.n5452 gnd.n5451 585
R10383 gnd.n5454 gnd.n5453 585
R10384 gnd.n5456 gnd.n5455 585
R10385 gnd.n5458 gnd.n5457 585
R10386 gnd.n5460 gnd.n5459 585
R10387 gnd.n5462 gnd.n5461 585
R10388 gnd.n5464 gnd.n5463 585
R10389 gnd.n5466 gnd.n5465 585
R10390 gnd.n5468 gnd.n5467 585
R10391 gnd.n5470 gnd.n5469 585
R10392 gnd.n5472 gnd.n5471 585
R10393 gnd.n5474 gnd.n5473 585
R10394 gnd.n5476 gnd.n5475 585
R10395 gnd.n5478 gnd.n5477 585
R10396 gnd.n5480 gnd.n5479 585
R10397 gnd.n5482 gnd.n5481 585
R10398 gnd.n5484 gnd.n5483 585
R10399 gnd.n5486 gnd.n5485 585
R10400 gnd.n5488 gnd.n5487 585
R10401 gnd.n5490 gnd.n5489 585
R10402 gnd.n5493 gnd.n5492 585
R10403 gnd.n5495 gnd.n5494 585
R10404 gnd.n5497 gnd.n5496 585
R10405 gnd.n5499 gnd.n5498 585
R10406 gnd.n5363 gnd.n3148 585
R10407 gnd.n5365 gnd.n5364 585
R10408 gnd.n5367 gnd.n5366 585
R10409 gnd.n5369 gnd.n5368 585
R10410 gnd.n5372 gnd.n5371 585
R10411 gnd.n5374 gnd.n5373 585
R10412 gnd.n5376 gnd.n5375 585
R10413 gnd.n5378 gnd.n5377 585
R10414 gnd.n5380 gnd.n5379 585
R10415 gnd.n5382 gnd.n5381 585
R10416 gnd.n5384 gnd.n5383 585
R10417 gnd.n5386 gnd.n5385 585
R10418 gnd.n5388 gnd.n5387 585
R10419 gnd.n5390 gnd.n5389 585
R10420 gnd.n5392 gnd.n5391 585
R10421 gnd.n5394 gnd.n5393 585
R10422 gnd.n5396 gnd.n5395 585
R10423 gnd.n5398 gnd.n5397 585
R10424 gnd.n5400 gnd.n5399 585
R10425 gnd.n5402 gnd.n5401 585
R10426 gnd.n5404 gnd.n5403 585
R10427 gnd.n5406 gnd.n5405 585
R10428 gnd.n5408 gnd.n5407 585
R10429 gnd.n5410 gnd.n5409 585
R10430 gnd.n5412 gnd.n5411 585
R10431 gnd.n5414 gnd.n5413 585
R10432 gnd.n5416 gnd.n5415 585
R10433 gnd.n5418 gnd.n5417 585
R10434 gnd.n5420 gnd.n5419 585
R10435 gnd.n5422 gnd.n5421 585
R10436 gnd.n5424 gnd.n5423 585
R10437 gnd.n5426 gnd.n5425 585
R10438 gnd.n5427 gnd.n3155 585
R10439 gnd.n5432 gnd.n3151 585
R10440 gnd.n5432 gnd.n5431 585
R10441 gnd.n5253 gnd.n3152 585
R10442 gnd.n3160 gnd.n3152 585
R10443 gnd.n5254 gnd.n3159 585
R10444 gnd.n5338 gnd.n3159 585
R10445 gnd.n5258 gnd.n5257 585
R10446 gnd.n5257 gnd.n5256 585
R10447 gnd.n5259 gnd.n3167 585
R10448 gnd.n5328 gnd.n3167 585
R10449 gnd.n5261 gnd.n5260 585
R10450 gnd.n5260 gnd.n3166 585
R10451 gnd.n5262 gnd.n3174 585
R10452 gnd.n5322 gnd.n3174 585
R10453 gnd.n5267 gnd.n5266 585
R10454 gnd.n5266 gnd.n5265 585
R10455 gnd.n5268 gnd.n3183 585
R10456 gnd.n5295 gnd.n3183 585
R10457 gnd.n5270 gnd.n5269 585
R10458 gnd.n5269 gnd.n3182 585
R10459 gnd.n5271 gnd.n3188 585
R10460 gnd.n5289 gnd.n3188 585
R10461 gnd.n5273 gnd.n5272 585
R10462 gnd.n5274 gnd.n5273 585
R10463 gnd.n5252 gnd.n3197 585
R10464 gnd.n3197 gnd.n3195 585
R10465 gnd.n5251 gnd.n5250 585
R10466 gnd.n5250 gnd.n5249 585
R10467 gnd.n3199 gnd.n3198 585
R10468 gnd.n3208 gnd.n3199 585
R10469 gnd.n5153 gnd.n3207 585
R10470 gnd.n5242 gnd.n3207 585
R10471 gnd.n5156 gnd.n5155 585
R10472 gnd.n5155 gnd.n5154 585
R10473 gnd.n5157 gnd.n3217 585
R10474 gnd.n5231 gnd.n3217 585
R10475 gnd.n5159 gnd.n5158 585
R10476 gnd.n5158 gnd.n3215 585
R10477 gnd.n5160 gnd.n3222 585
R10478 gnd.n5225 gnd.n3222 585
R10479 gnd.n5165 gnd.n5164 585
R10480 gnd.n5164 gnd.n5163 585
R10481 gnd.n5166 gnd.n3230 585
R10482 gnd.n5202 gnd.n3230 585
R10483 gnd.n5168 gnd.n5167 585
R10484 gnd.n5167 gnd.n3229 585
R10485 gnd.n5169 gnd.n3236 585
R10486 gnd.n5196 gnd.n3236 585
R10487 gnd.n5172 gnd.n5171 585
R10488 gnd.n5171 gnd.n5170 585
R10489 gnd.n5173 gnd.n3244 585
R10490 gnd.n5184 gnd.n3244 585
R10491 gnd.n5175 gnd.n5174 585
R10492 gnd.n5176 gnd.n5175 585
R10493 gnd.n5152 gnd.n3251 585
R10494 gnd.n5178 gnd.n3251 585
R10495 gnd.n5151 gnd.n5150 585
R10496 gnd.n5150 gnd.n5149 585
R10497 gnd.n3253 gnd.n3252 585
R10498 gnd.n5133 gnd.n3253 585
R10499 gnd.n5130 gnd.n5129 585
R10500 gnd.n5131 gnd.n5130 585
R10501 gnd.n5128 gnd.n3261 585
R10502 gnd.n5139 gnd.n3261 585
R10503 gnd.n5127 gnd.n5126 585
R10504 gnd.n5126 gnd.n5125 585
R10505 gnd.n3267 gnd.n3266 585
R10506 gnd.n5123 gnd.n3267 585
R10507 gnd.n5101 gnd.n5100 585
R10508 gnd.n5100 gnd.n3276 585
R10509 gnd.n5102 gnd.n3274 585
R10510 gnd.n5117 gnd.n3274 585
R10511 gnd.n5104 gnd.n5103 585
R10512 gnd.n5105 gnd.n5104 585
R10513 gnd.n5099 gnd.n3284 585
R10514 gnd.n3284 gnd.n3282 585
R10515 gnd.n5098 gnd.n5097 585
R10516 gnd.n5097 gnd.n5096 585
R10517 gnd.n3286 gnd.n3285 585
R10518 gnd.n3294 gnd.n3286 585
R10519 gnd.n4977 gnd.n3293 585
R10520 gnd.n5089 gnd.n3293 585
R10521 gnd.n4980 gnd.n4979 585
R10522 gnd.n4979 gnd.n4978 585
R10523 gnd.n4981 gnd.n3304 585
R10524 gnd.n5078 gnd.n3304 585
R10525 gnd.n4983 gnd.n4982 585
R10526 gnd.n4982 gnd.n3302 585
R10527 gnd.n4984 gnd.n3310 585
R10528 gnd.n5072 gnd.n3310 585
R10529 gnd.n4989 gnd.n4988 585
R10530 gnd.n4988 gnd.n4987 585
R10531 gnd.n4990 gnd.n3318 585
R10532 gnd.n5026 gnd.n3318 585
R10533 gnd.n4992 gnd.n4991 585
R10534 gnd.n4991 gnd.n3317 585
R10535 gnd.n4993 gnd.n3324 585
R10536 gnd.n5020 gnd.n3324 585
R10537 gnd.n4996 gnd.n4995 585
R10538 gnd.n4995 gnd.n4994 585
R10539 gnd.n4997 gnd.n3333 585
R10540 gnd.n5008 gnd.n3333 585
R10541 gnd.n4999 gnd.n4998 585
R10542 gnd.n5000 gnd.n4999 585
R10543 gnd.n4976 gnd.n3339 585
R10544 gnd.n5002 gnd.n3339 585
R10545 gnd.n4975 gnd.n4974 585
R10546 gnd.n4974 gnd.n4973 585
R10547 gnd.n3341 gnd.n3340 585
R10548 gnd.n4957 gnd.n3341 585
R10549 gnd.n4954 gnd.n4953 585
R10550 gnd.n4955 gnd.n4954 585
R10551 gnd.n4952 gnd.n3350 585
R10552 gnd.n4963 gnd.n3350 585
R10553 gnd.n4951 gnd.n4950 585
R10554 gnd.n4950 gnd.n4949 585
R10555 gnd.n3356 gnd.n3355 585
R10556 gnd.n4947 gnd.n3356 585
R10557 gnd.n4925 gnd.n4924 585
R10558 gnd.n4924 gnd.n3363 585
R10559 gnd.n4926 gnd.n3361 585
R10560 gnd.n4941 gnd.n3361 585
R10561 gnd.n4928 gnd.n4927 585
R10562 gnd.n4929 gnd.n4928 585
R10563 gnd.n4923 gnd.n3371 585
R10564 gnd.n3371 gnd.n3369 585
R10565 gnd.n4922 gnd.n4921 585
R10566 gnd.n4921 gnd.n4920 585
R10567 gnd.n3373 gnd.n3372 585
R10568 gnd.n3383 gnd.n3373 585
R10569 gnd.n4800 gnd.n3382 585
R10570 gnd.n4913 gnd.n3382 585
R10571 gnd.n4803 gnd.n4802 585
R10572 gnd.n4802 gnd.n4801 585
R10573 gnd.n4804 gnd.n3392 585
R10574 gnd.n4902 gnd.n3392 585
R10575 gnd.n4806 gnd.n4805 585
R10576 gnd.n4805 gnd.n3390 585
R10577 gnd.n4807 gnd.n3398 585
R10578 gnd.n4896 gnd.n3398 585
R10579 gnd.n4811 gnd.n4810 585
R10580 gnd.n4810 gnd.n4809 585
R10581 gnd.n4812 gnd.n3405 585
R10582 gnd.n4849 gnd.n3405 585
R10583 gnd.n4814 gnd.n4813 585
R10584 gnd.n4813 gnd.n3411 585
R10585 gnd.n4815 gnd.n3410 585
R10586 gnd.n4843 gnd.n3410 585
R10587 gnd.n4819 gnd.n4818 585
R10588 gnd.n4818 gnd.n4817 585
R10589 gnd.n4820 gnd.n3419 585
R10590 gnd.n4831 gnd.n3419 585
R10591 gnd.n4822 gnd.n4821 585
R10592 gnd.n4823 gnd.n4822 585
R10593 gnd.n4799 gnd.n3426 585
R10594 gnd.n4825 gnd.n3426 585
R10595 gnd.n4798 gnd.n4797 585
R10596 gnd.n4797 gnd.n4796 585
R10597 gnd.n3428 gnd.n3427 585
R10598 gnd.n4780 gnd.n3428 585
R10599 gnd.n4731 gnd.n4730 585
R10600 gnd.n4730 gnd.n4729 585
R10601 gnd.n4732 gnd.n3435 585
R10602 gnd.n4786 gnd.n3435 585
R10603 gnd.n4735 gnd.n4734 585
R10604 gnd.n4734 gnd.n4733 585
R10605 gnd.n4736 gnd.n3448 585
R10606 gnd.n4762 gnd.n3448 585
R10607 gnd.n4738 gnd.n4737 585
R10608 gnd.n4737 gnd.n3454 585
R10609 gnd.n4739 gnd.n3453 585
R10610 gnd.n4756 gnd.n3453 585
R10611 gnd.n4741 gnd.n4740 585
R10612 gnd.n4743 gnd.n4741 585
R10613 gnd.n4728 gnd.n3462 585
R10614 gnd.n3462 gnd.n3460 585
R10615 gnd.n4727 gnd.n4726 585
R10616 gnd.n4726 gnd.n4725 585
R10617 gnd.n3464 gnd.n3463 585
R10618 gnd.n3473 gnd.n3464 585
R10619 gnd.n4652 gnd.n3472 585
R10620 gnd.n4718 gnd.n3472 585
R10621 gnd.n4655 gnd.n4654 585
R10622 gnd.n4654 gnd.n4653 585
R10623 gnd.n4656 gnd.n3482 585
R10624 gnd.n4706 gnd.n3482 585
R10625 gnd.n4658 gnd.n4657 585
R10626 gnd.n4657 gnd.n3480 585
R10627 gnd.n4659 gnd.n3487 585
R10628 gnd.n4700 gnd.n3487 585
R10629 gnd.n4663 gnd.n4662 585
R10630 gnd.n4662 gnd.n4661 585
R10631 gnd.n4664 gnd.n3495 585
R10632 gnd.n4676 gnd.n3495 585
R10633 gnd.n6061 gnd.n861 585
R10634 gnd.n2317 gnd.n861 585
R10635 gnd.n6901 gnd.n299 585
R10636 gnd.n6901 gnd.n6900 585
R10637 gnd.n6903 gnd.n6902 585
R10638 gnd.n6902 gnd.n83 585
R10639 gnd.n6904 gnd.n293 585
R10640 gnd.n293 gnd.n81 585
R10641 gnd.n6906 gnd.n6905 585
R10642 gnd.n6906 gnd.n162 585
R10643 gnd.n6907 gnd.n292 585
R10644 gnd.n6907 gnd.n171 585
R10645 gnd.n6909 gnd.n6908 585
R10646 gnd.n6908 gnd.n169 585
R10647 gnd.n6910 gnd.n287 585
R10648 gnd.n287 gnd.n182 585
R10649 gnd.n6912 gnd.n6911 585
R10650 gnd.n6912 gnd.n179 585
R10651 gnd.n6934 gnd.n286 585
R10652 gnd.n6934 gnd.n6933 585
R10653 gnd.n6936 gnd.n6935 585
R10654 gnd.n6935 gnd.n188 585
R10655 gnd.n6937 gnd.n271 585
R10656 gnd.n271 gnd.n197 585
R10657 gnd.n6939 gnd.n6938 585
R10658 gnd.n6940 gnd.n6939 585
R10659 gnd.n272 gnd.n270 585
R10660 gnd.n270 gnd.n205 585
R10661 gnd.n280 gnd.n279 585
R10662 gnd.n279 gnd.n203 585
R10663 gnd.n278 gnd.n277 585
R10664 gnd.n278 gnd.n214 585
R10665 gnd.n276 gnd.n262 585
R10666 gnd.n262 gnd.n211 585
R10667 gnd.n6953 gnd.n261 585
R10668 gnd.n6953 gnd.n6952 585
R10669 gnd.n6955 gnd.n6954 585
R10670 gnd.n6954 gnd.n220 585
R10671 gnd.n6956 gnd.n258 585
R10672 gnd.n258 gnd.n251 585
R10673 gnd.n6959 gnd.n6958 585
R10674 gnd.n6960 gnd.n6959 585
R10675 gnd.n259 gnd.n257 585
R10676 gnd.n257 gnd.n255 585
R10677 gnd.n5723 gnd.n2728 585
R10678 gnd.n5706 gnd.n2728 585
R10679 gnd.n5725 gnd.n5724 585
R10680 gnd.n5726 gnd.n5725 585
R10681 gnd.n5720 gnd.n2727 585
R10682 gnd.n2727 gnd.n2721 585
R10683 gnd.n5719 gnd.n5718 585
R10684 gnd.n5718 gnd.n5717 585
R10685 gnd.n5653 gnd.n2730 585
R10686 gnd.n2730 gnd.n236 585
R10687 gnd.n5655 gnd.n5654 585
R10688 gnd.n5654 gnd.n233 585
R10689 gnd.n5657 gnd.n5650 585
R10690 gnd.n5650 gnd.n2707 585
R10691 gnd.n5659 gnd.n5658 585
R10692 gnd.n5659 gnd.n2704 585
R10693 gnd.n5660 gnd.n5649 585
R10694 gnd.n5660 gnd.n2710 585
R10695 gnd.n5662 gnd.n5661 585
R10696 gnd.n5661 gnd.n2741 585
R10697 gnd.n5663 gnd.n2751 585
R10698 gnd.n2751 gnd.n2738 585
R10699 gnd.n5665 gnd.n5664 585
R10700 gnd.n5666 gnd.n5665 585
R10701 gnd.n2752 gnd.n2750 585
R10702 gnd.n2750 gnd.n2747 585
R10703 gnd.n5643 gnd.n5642 585
R10704 gnd.n5642 gnd.n5641 585
R10705 gnd.n2755 gnd.n2754 585
R10706 gnd.n2765 gnd.n2755 585
R10707 gnd.n5611 gnd.n2778 585
R10708 gnd.n2778 gnd.n2763 585
R10709 gnd.n5613 gnd.n5612 585
R10710 gnd.n5614 gnd.n5613 585
R10711 gnd.n2779 gnd.n2777 585
R10712 gnd.n2777 gnd.n2772 585
R10713 gnd.n5606 gnd.n5605 585
R10714 gnd.n5605 gnd.n5604 585
R10715 gnd.n2789 gnd.n2781 585
R10716 gnd.n5593 gnd.n2789 585
R10717 gnd.n2788 gnd.n2787 585
R10718 gnd.n2788 gnd.n2682 585
R10719 gnd.n2783 gnd.n2782 585
R10720 gnd.n2782 gnd.n2679 585
R10721 gnd.n2666 gnd.n2665 585
R10722 gnd.n2670 gnd.n2666 585
R10723 gnd.n5782 gnd.n5781 585
R10724 gnd.n5781 gnd.n5780 585
R10725 gnd.n5783 gnd.n2660 585
R10726 gnd.n2667 gnd.n2660 585
R10727 gnd.n5785 gnd.n5784 585
R10728 gnd.n5786 gnd.n5785 585
R10729 gnd.n2657 gnd.n2656 585
R10730 gnd.n5787 gnd.n2657 585
R10731 gnd.n5790 gnd.n5789 585
R10732 gnd.n5789 gnd.n5788 585
R10733 gnd.n5791 gnd.n2651 585
R10734 gnd.n2651 gnd.n2649 585
R10735 gnd.n5793 gnd.n5792 585
R10736 gnd.n5794 gnd.n5793 585
R10737 gnd.n2652 gnd.n2650 585
R10738 gnd.n2650 gnd.n2647 585
R10739 gnd.n5531 gnd.n5530 585
R10740 gnd.n5532 gnd.n5531 585
R10741 gnd.n2961 gnd.n2960 585
R10742 gnd.n5520 gnd.n2960 585
R10743 gnd.n5525 gnd.n5524 585
R10744 gnd.n5524 gnd.n5523 585
R10745 gnd.n2964 gnd.n2963 585
R10746 gnd.n5509 gnd.n2964 585
R10747 gnd.n5507 gnd.n5506 585
R10748 gnd.n5508 gnd.n5507 585
R10749 gnd.n2973 gnd.n2972 585
R10750 gnd.n5306 gnd.n2972 585
R10751 gnd.n5502 gnd.n5501 585
R10752 gnd.n5501 gnd.n5500 585
R10753 gnd.n2976 gnd.n2975 585
R10754 gnd.n3153 gnd.n2976 585
R10755 gnd.n5336 gnd.n5335 585
R10756 gnd.n5337 gnd.n5336 585
R10757 gnd.n3162 gnd.n3161 585
R10758 gnd.n5255 gnd.n3161 585
R10759 gnd.n5331 gnd.n5330 585
R10760 gnd.n5330 gnd.n5329 585
R10761 gnd.n3165 gnd.n3164 585
R10762 gnd.n3173 gnd.n3165 585
R10763 gnd.n5283 gnd.n3190 585
R10764 gnd.n5263 gnd.n3190 585
R10765 gnd.n5285 gnd.n5284 585
R10766 gnd.n5286 gnd.n5285 585
R10767 gnd.n3191 gnd.n3189 585
R10768 gnd.n3189 gnd.n3187 585
R10769 gnd.n5278 gnd.n5277 585
R10770 gnd.n5277 gnd.n5276 585
R10771 gnd.n3194 gnd.n3193 585
R10772 gnd.n3200 gnd.n3194 585
R10773 gnd.n5240 gnd.n5239 585
R10774 gnd.n5241 gnd.n5240 585
R10775 gnd.n3211 gnd.n3210 585
R10776 gnd.n3218 gnd.n3210 585
R10777 gnd.n5235 gnd.n5234 585
R10778 gnd.n5234 gnd.n5233 585
R10779 gnd.n3214 gnd.n3213 585
R10780 gnd.n5162 gnd.n3214 585
R10781 gnd.n5192 gnd.n3238 585
R10782 gnd.n3238 gnd.n3231 585
R10783 gnd.n5194 gnd.n5193 585
R10784 gnd.n5195 gnd.n5194 585
R10785 gnd.n3239 gnd.n3237 585
R10786 gnd.n3237 gnd.n3235 585
R10787 gnd.n5187 gnd.n5186 585
R10788 gnd.n5186 gnd.n5185 585
R10789 gnd.n3242 gnd.n3241 585
R10790 gnd.n5177 gnd.n3242 585
R10791 gnd.n5147 gnd.n5146 585
R10792 gnd.n5148 gnd.n5147 585
R10793 gnd.n3256 gnd.n3255 585
R10794 gnd.n5132 gnd.n3255 585
R10795 gnd.n5142 gnd.n5141 585
R10796 gnd.n5141 gnd.n5140 585
R10797 gnd.n3259 gnd.n3258 585
R10798 gnd.n5124 gnd.n3259 585
R10799 gnd.n5114 gnd.n5113 585
R10800 gnd.n5115 gnd.n5114 585
R10801 gnd.n3278 gnd.n3277 585
R10802 gnd.n3277 gnd.n3273 585
R10803 gnd.n5109 gnd.n5108 585
R10804 gnd.n5108 gnd.n5107 585
R10805 gnd.n3281 gnd.n3280 585
R10806 gnd.n3287 gnd.n3281 585
R10807 gnd.n5087 gnd.n5086 585
R10808 gnd.n5088 gnd.n5087 585
R10809 gnd.n3298 gnd.n3297 585
R10810 gnd.n3305 gnd.n3297 585
R10811 gnd.n5082 gnd.n5081 585
R10812 gnd.n5081 gnd.n5080 585
R10813 gnd.n3301 gnd.n3300 585
R10814 gnd.n3309 gnd.n3301 585
R10815 gnd.n5016 gnd.n3326 585
R10816 gnd.n3326 gnd.n3319 585
R10817 gnd.n5018 gnd.n5017 585
R10818 gnd.n5019 gnd.n5018 585
R10819 gnd.n3327 gnd.n3325 585
R10820 gnd.n3325 gnd.n3323 585
R10821 gnd.n5011 gnd.n5010 585
R10822 gnd.n5010 gnd.n5009 585
R10823 gnd.n3330 gnd.n3329 585
R10824 gnd.n5001 gnd.n3330 585
R10825 gnd.n4971 gnd.n4970 585
R10826 gnd.n4972 gnd.n4971 585
R10827 gnd.n3344 gnd.n3343 585
R10828 gnd.n4956 gnd.n3343 585
R10829 gnd.n4966 gnd.n4965 585
R10830 gnd.n4965 gnd.n4964 585
R10831 gnd.n3347 gnd.n3346 585
R10832 gnd.n4948 gnd.n3347 585
R10833 gnd.n4938 gnd.n4937 585
R10834 gnd.n4939 gnd.n4938 585
R10835 gnd.n3365 gnd.n3364 585
R10836 gnd.n3364 gnd.n3360 585
R10837 gnd.n4933 gnd.n4932 585
R10838 gnd.n4932 gnd.n4931 585
R10839 gnd.n3368 gnd.n3367 585
R10840 gnd.n3374 gnd.n3368 585
R10841 gnd.n4911 gnd.n4910 585
R10842 gnd.n4912 gnd.n4911 585
R10843 gnd.n3386 gnd.n3385 585
R10844 gnd.n3393 gnd.n3385 585
R10845 gnd.n4906 gnd.n4905 585
R10846 gnd.n4905 gnd.n4904 585
R10847 gnd.n3389 gnd.n3388 585
R10848 gnd.n3397 gnd.n3389 585
R10849 gnd.n4839 gnd.n3413 585
R10850 gnd.n3413 gnd.n3406 585
R10851 gnd.n4841 gnd.n4840 585
R10852 gnd.n4842 gnd.n4841 585
R10853 gnd.n3414 gnd.n3412 585
R10854 gnd.n4816 gnd.n3412 585
R10855 gnd.n4834 gnd.n4833 585
R10856 gnd.n4833 gnd.n4832 585
R10857 gnd.n3417 gnd.n3416 585
R10858 gnd.n4824 gnd.n3417 585
R10859 gnd.n4794 gnd.n4793 585
R10860 gnd.n4795 gnd.n4794 585
R10861 gnd.n3430 gnd.n3429 585
R10862 gnd.n3440 gnd.n3429 585
R10863 gnd.n4789 gnd.n4788 585
R10864 gnd.n4788 gnd.n4787 585
R10865 gnd.n3433 gnd.n3432 585
R10866 gnd.n3449 gnd.n3433 585
R10867 gnd.n4753 gnd.n4752 585
R10868 gnd.n4754 gnd.n4753 585
R10869 gnd.n3456 gnd.n3455 585
R10870 gnd.n4742 gnd.n3455 585
R10871 gnd.n4748 gnd.n4747 585
R10872 gnd.n4747 gnd.n4746 585
R10873 gnd.n3459 gnd.n3458 585
R10874 gnd.n3465 gnd.n3459 585
R10875 gnd.n4716 gnd.n4715 585
R10876 gnd.n4717 gnd.n4716 585
R10877 gnd.n3476 gnd.n3475 585
R10878 gnd.t97 gnd.n3475 585
R10879 gnd.n4711 gnd.n4710 585
R10880 gnd.n4710 gnd.n4709 585
R10881 gnd.n3479 gnd.n3478 585
R10882 gnd.n3486 gnd.n3479 585
R10883 gnd.n4501 gnd.n4500 585
R10884 gnd.n4500 gnd.n3496 585
R10885 gnd.n4502 gnd.n3747 585
R10886 gnd.n3747 gnd.n3494 585
R10887 gnd.n4504 gnd.n4503 585
R10888 gnd.n4505 gnd.n4504 585
R10889 gnd.n3748 gnd.n3746 585
R10890 gnd.n3746 gnd.n3745 585
R10891 gnd.n4494 gnd.n4493 585
R10892 gnd.n4493 gnd.n4492 585
R10893 gnd.n3751 gnd.n3750 585
R10894 gnd.n4489 gnd.n3751 585
R10895 gnd.n4484 gnd.n4483 585
R10896 gnd.n4485 gnd.n4484 585
R10897 gnd.n3754 gnd.n3753 585
R10898 gnd.n4475 gnd.n3753 585
R10899 gnd.n4479 gnd.n4478 585
R10900 gnd.n4478 gnd.n4477 585
R10901 gnd.n3757 gnd.n3756 585
R10902 gnd.n4473 gnd.n3757 585
R10903 gnd.n4471 gnd.n4470 585
R10904 gnd.n4472 gnd.n4471 585
R10905 gnd.n3892 gnd.n3891 585
R10906 gnd.n4463 gnd.n3891 585
R10907 gnd.n4466 gnd.n4465 585
R10908 gnd.n4465 gnd.n4464 585
R10909 gnd.n4461 gnd.n3894 585
R10910 gnd.n4462 gnd.n4461 585
R10911 gnd.n4460 gnd.n4458 585
R10912 gnd.n4460 gnd.n4459 585
R10913 gnd.n3896 gnd.n3895 585
R10914 gnd.n3895 gnd.n2537 585
R10915 gnd.n4454 gnd.n4453 585
R10916 gnd.n4453 gnd.n2534 585
R10917 gnd.n4452 gnd.n3898 585
R10918 gnd.n4452 gnd.n2527 585
R10919 gnd.n4451 gnd.n4450 585
R10920 gnd.n4451 gnd.n2524 585
R10921 gnd.n3900 gnd.n3899 585
R10922 gnd.n3899 gnd.n2516 585
R10923 gnd.n4446 gnd.n4445 585
R10924 gnd.n4445 gnd.n2513 585
R10925 gnd.n4444 gnd.n3902 585
R10926 gnd.n4444 gnd.n2505 585
R10927 gnd.n4443 gnd.n3904 585
R10928 gnd.n4443 gnd.n4442 585
R10929 gnd.n4376 gnd.n3903 585
R10930 gnd.n3903 gnd.n2495 585
R10931 gnd.n4378 gnd.n4377 585
R10932 gnd.n4377 gnd.n2492 585
R10933 gnd.n4379 gnd.n4369 585
R10934 gnd.n4369 gnd.n2484 585
R10935 gnd.n4381 gnd.n4380 585
R10936 gnd.n4381 gnd.n2481 585
R10937 gnd.n4382 gnd.n4368 585
R10938 gnd.n4382 gnd.n3919 585
R10939 gnd.n4384 gnd.n4383 585
R10940 gnd.n4383 gnd.n2471 585
R10941 gnd.n4385 gnd.n3928 585
R10942 gnd.n3928 gnd.n2463 585
R10943 gnd.n4387 gnd.n4386 585
R10944 gnd.n4388 gnd.n4387 585
R10945 gnd.n3929 gnd.n3927 585
R10946 gnd.n3927 gnd.n2453 585
R10947 gnd.n4318 gnd.n4317 585
R10948 gnd.n4318 gnd.n2450 585
R10949 gnd.n4320 gnd.n4319 585
R10950 gnd.n4319 gnd.n2445 585
R10951 gnd.n4322 gnd.n4321 585
R10952 gnd.n4322 gnd.n2442 585
R10953 gnd.n4325 gnd.n4324 585
R10954 gnd.n4326 gnd.n4325 585
R10955 gnd.n4323 gnd.n4316 585
R10956 gnd.n4316 gnd.n2433 585
R10957 gnd.n3940 gnd.n3939 585
R10958 gnd.n3939 gnd.n2428 585
R10959 gnd.n4354 gnd.n3941 585
R10960 gnd.n4354 gnd.n4353 585
R10961 gnd.n4356 gnd.n4355 585
R10962 gnd.n4355 gnd.n2418 585
R10963 gnd.n4358 gnd.n4357 585
R10964 gnd.n4358 gnd.n2415 585
R10965 gnd.n4359 gnd.n3937 585
R10966 gnd.n4359 gnd.n2409 585
R10967 gnd.n4361 gnd.n4360 585
R10968 gnd.n4360 gnd.n2406 585
R10969 gnd.n3938 gnd.n3936 585
R10970 gnd.n3938 gnd.n2398 585
R10971 gnd.n4273 gnd.n4272 585
R10972 gnd.n4272 gnd.n2395 585
R10973 gnd.n4274 gnd.n3968 585
R10974 gnd.n3968 gnd.n2387 585
R10975 gnd.n4276 gnd.n4275 585
R10976 gnd.n4277 gnd.n4276 585
R10977 gnd.n3969 gnd.n3967 585
R10978 gnd.n3967 gnd.n2377 585
R10979 gnd.n4266 gnd.n4265 585
R10980 gnd.n4265 gnd.n2374 585
R10981 gnd.n4264 gnd.n3971 585
R10982 gnd.n4264 gnd.n2366 585
R10983 gnd.n4263 gnd.n4262 585
R10984 gnd.n4263 gnd.n2363 585
R10985 gnd.n3973 gnd.n3972 585
R10986 gnd.n3972 gnd.n2355 585
R10987 gnd.n4258 gnd.n4257 585
R10988 gnd.n4257 gnd.n2352 585
R10989 gnd.n4256 gnd.n3975 585
R10990 gnd.n4256 gnd.n2344 585
R10991 gnd.n4255 gnd.n4254 585
R10992 gnd.n4255 gnd.n2341 585
R10993 gnd.n3977 gnd.n3976 585
R10994 gnd.n3976 gnd.n2332 585
R10995 gnd.n4250 gnd.n4249 585
R10996 gnd.n4249 gnd.n4248 585
R10997 gnd.n866 gnd.n865 585
R10998 gnd.n2321 gnd.n866 585
R10999 gnd.n6058 gnd.n6057 585
R11000 gnd.n6057 gnd.n6056 585
R11001 gnd.n5797 gnd.n5796 585
R11002 gnd.n5796 gnd.n5795 585
R11003 gnd.n5798 gnd.n2644 585
R11004 gnd.n5533 gnd.n2644 585
R11005 gnd.n5799 gnd.n2643 585
R11006 gnd.n5519 gnd.n2643 585
R11007 gnd.n5521 gnd.n2641 585
R11008 gnd.n5522 gnd.n5521 585
R11009 gnd.n5803 gnd.n2640 585
R11010 gnd.n2965 gnd.n2640 585
R11011 gnd.n5804 gnd.n2639 585
R11012 gnd.n5510 gnd.n2639 585
R11013 gnd.n5805 gnd.n2638 585
R11014 gnd.n2971 gnd.n2638 585
R11015 gnd.n5307 gnd.n2636 585
R11016 gnd.n5308 gnd.n5307 585
R11017 gnd.n5809 gnd.n2635 585
R11018 gnd.n2977 gnd.n2635 585
R11019 gnd.n5810 gnd.n2634 585
R11020 gnd.n5303 gnd.n2634 585
R11021 gnd.n5811 gnd.n2633 585
R11022 gnd.n3158 gnd.n2633 585
R11023 gnd.n3168 gnd.n2631 585
R11024 gnd.n3169 gnd.n3168 585
R11025 gnd.n5815 gnd.n2630 585
R11026 gnd.n5321 gnd.n2630 585
R11027 gnd.n5816 gnd.n2629 585
R11028 gnd.n5264 gnd.n2629 585
R11029 gnd.n5817 gnd.n2628 585
R11030 gnd.n5296 gnd.n2628 585
R11031 gnd.n5287 gnd.n2626 585
R11032 gnd.n5288 gnd.n5287 585
R11033 gnd.n5821 gnd.n2625 585
R11034 gnd.n5275 gnd.n2625 585
R11035 gnd.n5822 gnd.n2624 585
R11036 gnd.n3201 gnd.n2624 585
R11037 gnd.n5823 gnd.n2623 585
R11038 gnd.n3209 gnd.n2623 585
R11039 gnd.n3206 gnd.n2621 585
R11040 gnd.t154 gnd.n3206 585
R11041 gnd.n5827 gnd.n2620 585
R11042 gnd.n5232 gnd.n2620 585
R11043 gnd.n5828 gnd.n2619 585
R11044 gnd.n5224 gnd.n2619 585
R11045 gnd.n5829 gnd.n2618 585
R11046 gnd.n5161 gnd.n2618 585
R11047 gnd.n5203 gnd.n2616 585
R11048 gnd.n5204 gnd.n5203 585
R11049 gnd.n5833 gnd.n2615 585
R11050 gnd.n5196 gnd.n2615 585
R11051 gnd.n5834 gnd.n2614 585
R11052 gnd.n3245 gnd.n2614 585
R11053 gnd.n5835 gnd.n2613 585
R11054 gnd.n3243 gnd.n2613 585
R11055 gnd.n3249 gnd.n2611 585
R11056 gnd.n3250 gnd.n3249 585
R11057 gnd.n5839 gnd.n2610 585
R11058 gnd.n3254 gnd.n2610 585
R11059 gnd.n5840 gnd.n2609 585
R11060 gnd.n3262 gnd.n2609 585
R11061 gnd.n5841 gnd.n2608 585
R11062 gnd.n3260 gnd.n2608 585
R11063 gnd.n3268 gnd.n2606 585
R11064 gnd.n3269 gnd.n3268 585
R11065 gnd.n5845 gnd.n2605 585
R11066 gnd.n5116 gnd.n2605 585
R11067 gnd.n5846 gnd.n2604 585
R11068 gnd.n5106 gnd.n2604 585
R11069 gnd.n5847 gnd.n2603 585
R11070 gnd.n5035 gnd.n2603 585
R11071 gnd.n3295 gnd.n2601 585
R11072 gnd.n3296 gnd.n3295 585
R11073 gnd.n5851 gnd.n2600 585
R11074 gnd.n3292 gnd.n2600 585
R11075 gnd.n5852 gnd.n2599 585
R11076 gnd.n5079 gnd.n2599 585
R11077 gnd.n5853 gnd.n2598 585
R11078 gnd.n5071 gnd.n2598 585
R11079 gnd.n4985 gnd.n2596 585
R11080 gnd.n4986 gnd.n4985 585
R11081 gnd.n5857 gnd.n2595 585
R11082 gnd.n5027 gnd.n2595 585
R11083 gnd.n5858 gnd.n2594 585
R11084 gnd.n5020 gnd.n2594 585
R11085 gnd.n5859 gnd.n2593 585
R11086 gnd.n3334 gnd.n2593 585
R11087 gnd.n3331 gnd.n2591 585
R11088 gnd.n3332 gnd.n3331 585
R11089 gnd.n5863 gnd.n2590 585
R11090 gnd.n3338 gnd.n2590 585
R11091 gnd.n5864 gnd.n2589 585
R11092 gnd.n3342 gnd.n2589 585
R11093 gnd.n5865 gnd.n2588 585
R11094 gnd.n3351 gnd.n2588 585
R11095 gnd.n3348 gnd.n2586 585
R11096 gnd.n3349 gnd.n3348 585
R11097 gnd.n5869 gnd.n2585 585
R11098 gnd.n4861 gnd.n2585 585
R11099 gnd.n5870 gnd.n2584 585
R11100 gnd.n4940 gnd.n2584 585
R11101 gnd.n5871 gnd.n2583 585
R11102 gnd.n4930 gnd.n2583 585
R11103 gnd.n3375 gnd.n2581 585
R11104 gnd.n3376 gnd.n3375 585
R11105 gnd.n5875 gnd.n2580 585
R11106 gnd.n3384 gnd.n2580 585
R11107 gnd.n5876 gnd.n2579 585
R11108 gnd.n3381 gnd.n2579 585
R11109 gnd.n5877 gnd.n2578 585
R11110 gnd.n4903 gnd.n2578 585
R11111 gnd.n4894 gnd.n2576 585
R11112 gnd.n4895 gnd.n4894 585
R11113 gnd.n5881 gnd.n2575 585
R11114 gnd.n4808 gnd.n2575 585
R11115 gnd.n5882 gnd.n2574 585
R11116 gnd.n4850 gnd.n2574 585
R11117 gnd.n5883 gnd.n2573 585
R11118 gnd.n4843 gnd.n2573 585
R11119 gnd.n3420 gnd.n2571 585
R11120 gnd.n3421 gnd.n3420 585
R11121 gnd.n5887 gnd.n2570 585
R11122 gnd.n3418 gnd.n2570 585
R11123 gnd.n5888 gnd.n2569 585
R11124 gnd.n3425 gnd.n2569 585
R11125 gnd.n5889 gnd.n2568 585
R11126 gnd.n4779 gnd.n2568 585
R11127 gnd.n3436 gnd.n2566 585
R11128 gnd.t249 gnd.n3436 585
R11129 gnd.n5893 gnd.n2565 585
R11130 gnd.n3434 gnd.n2565 585
R11131 gnd.n5894 gnd.n2564 585
R11132 gnd.n4763 gnd.n2564 585
R11133 gnd.n5895 gnd.n2563 585
R11134 gnd.n4755 gnd.n2563 585
R11135 gnd.n4744 gnd.n2561 585
R11136 gnd.n4745 gnd.n4744 585
R11137 gnd.n5899 gnd.n2560 585
R11138 gnd.n3466 gnd.n2560 585
R11139 gnd.n5900 gnd.n2559 585
R11140 gnd.n3474 gnd.n2559 585
R11141 gnd.n5901 gnd.n2558 585
R11142 gnd.n3471 gnd.n2558 585
R11143 gnd.n4707 gnd.n2556 585
R11144 gnd.n4708 gnd.n4707 585
R11145 gnd.n5905 gnd.n2555 585
R11146 gnd.n4699 gnd.n2555 585
R11147 gnd.n5906 gnd.n2554 585
R11148 gnd.n4660 gnd.n2554 585
R11149 gnd.n5907 gnd.n2553 585
R11150 gnd.n4677 gnd.n2553 585
R11151 gnd.n3520 gnd.n2551 585
R11152 gnd.n3521 gnd.n3520 585
R11153 gnd.n5911 gnd.n2550 585
R11154 gnd.n4506 gnd.n2550 585
R11155 gnd.n5912 gnd.n2549 585
R11156 gnd.n4491 gnd.n2549 585
R11157 gnd.n5913 gnd.n2548 585
R11158 gnd.n4490 gnd.n2548 585
R11159 gnd.n4487 gnd.n2546 585
R11160 gnd.n4488 gnd.n4487 585
R11161 gnd.n5917 gnd.n2545 585
R11162 gnd.n3752 gnd.n2545 585
R11163 gnd.n5918 gnd.n2544 585
R11164 gnd.n4476 gnd.n2544 585
R11165 gnd.n5919 gnd.n2543 585
R11166 gnd.n4474 gnd.n2543 585
R11167 gnd.n3888 gnd.n3887 585
R11168 gnd.n3886 gnd.n3774 585
R11169 gnd.n3776 gnd.n3773 585
R11170 gnd.n3890 gnd.n3773 585
R11171 gnd.n3879 gnd.n3789 585
R11172 gnd.n3878 gnd.n3790 585
R11173 gnd.n3792 gnd.n3791 585
R11174 gnd.n3871 gnd.n3800 585
R11175 gnd.n3870 gnd.n3801 585
R11176 gnd.n3811 gnd.n3802 585
R11177 gnd.n3863 gnd.n3812 585
R11178 gnd.n3862 gnd.n3813 585
R11179 gnd.n3815 gnd.n3814 585
R11180 gnd.n3855 gnd.n3823 585
R11181 gnd.n3854 gnd.n3824 585
R11182 gnd.n3836 gnd.n3825 585
R11183 gnd.n3847 gnd.n3837 585
R11184 gnd.n3846 gnd.n3839 585
R11185 gnd.n3838 gnd.n3720 585
R11186 gnd.n4534 gnd.n3721 585
R11187 gnd.n4533 gnd.n3722 585
R11188 gnd.n4532 gnd.n3723 585
R11189 gnd.n3767 gnd.n3724 585
R11190 gnd.n4528 gnd.n3726 585
R11191 gnd.n4527 gnd.n3727 585
R11192 gnd.n4526 gnd.n3728 585
R11193 gnd.n4523 gnd.n3733 585
R11194 gnd.n4522 gnd.n3734 585
R11195 gnd.n4521 gnd.n3735 585
R11196 gnd.n3771 gnd.n3736 585
R11197 gnd.n5536 gnd.n2648 585
R11198 gnd.n5795 gnd.n2648 585
R11199 gnd.n5535 gnd.n5534 585
R11200 gnd.n5534 gnd.n5533 585
R11201 gnd.n2959 gnd.n2958 585
R11202 gnd.n5519 gnd.n2959 585
R11203 gnd.n5518 gnd.n5517 585
R11204 gnd.n5522 gnd.n5518 585
R11205 gnd.n2967 gnd.n2966 585
R11206 gnd.n2966 gnd.n2965 585
R11207 gnd.n5512 gnd.n5511 585
R11208 gnd.n5511 gnd.n5510 585
R11209 gnd.n2970 gnd.n2969 585
R11210 gnd.n2971 gnd.n2970 585
R11211 gnd.n5310 gnd.n5309 585
R11212 gnd.n5309 gnd.n5308 585
R11213 gnd.n5313 gnd.n5305 585
R11214 gnd.n5305 gnd.n2977 585
R11215 gnd.n5314 gnd.n5304 585
R11216 gnd.n5304 gnd.n5303 585
R11217 gnd.n5315 gnd.n5302 585
R11218 gnd.n5302 gnd.n3158 585
R11219 gnd.n3178 gnd.n3176 585
R11220 gnd.n3176 gnd.n3169 585
R11221 gnd.n5320 gnd.n5319 585
R11222 gnd.n5321 gnd.n5320 585
R11223 gnd.n3177 gnd.n3175 585
R11224 gnd.n5264 gnd.n3175 585
R11225 gnd.n5298 gnd.n5297 585
R11226 gnd.n5297 gnd.n5296 585
R11227 gnd.n3181 gnd.n3180 585
R11228 gnd.n5288 gnd.n3181 585
R11229 gnd.n5213 gnd.n3196 585
R11230 gnd.n5275 gnd.n3196 585
R11231 gnd.n5216 gnd.n5212 585
R11232 gnd.n5212 gnd.n3201 585
R11233 gnd.n5217 gnd.n5211 585
R11234 gnd.n5211 gnd.n3209 585
R11235 gnd.n5218 gnd.n5210 585
R11236 gnd.n5210 gnd.t154 585
R11237 gnd.n3225 gnd.n3216 585
R11238 gnd.n5232 gnd.n3216 585
R11239 gnd.n5223 gnd.n5222 585
R11240 gnd.n5224 gnd.n5223 585
R11241 gnd.n3224 gnd.n3223 585
R11242 gnd.n5161 gnd.n3223 585
R11243 gnd.n5206 gnd.n5205 585
R11244 gnd.n5205 gnd.n5204 585
R11245 gnd.n3228 gnd.n3227 585
R11246 gnd.n5196 gnd.n3228 585
R11247 gnd.n5048 gnd.n5047 585
R11248 gnd.n5047 gnd.n3245 585
R11249 gnd.n5051 gnd.n5046 585
R11250 gnd.n5046 gnd.n3243 585
R11251 gnd.n5052 gnd.n5045 585
R11252 gnd.n5045 gnd.n3250 585
R11253 gnd.n5053 gnd.n5044 585
R11254 gnd.n5044 gnd.n3254 585
R11255 gnd.n5043 gnd.n5041 585
R11256 gnd.n5043 gnd.n3262 585
R11257 gnd.n5057 gnd.n5040 585
R11258 gnd.n5040 gnd.n3260 585
R11259 gnd.n5058 gnd.n5039 585
R11260 gnd.n5039 gnd.n3269 585
R11261 gnd.n5059 gnd.n3275 585
R11262 gnd.n5116 gnd.n3275 585
R11263 gnd.n5037 gnd.n3283 585
R11264 gnd.n5106 gnd.n3283 585
R11265 gnd.n5063 gnd.n5036 585
R11266 gnd.n5036 gnd.n5035 585
R11267 gnd.n5064 gnd.n5034 585
R11268 gnd.n5034 gnd.n3296 585
R11269 gnd.n5065 gnd.n5033 585
R11270 gnd.n5033 gnd.n3292 585
R11271 gnd.n3313 gnd.n3303 585
R11272 gnd.n5079 gnd.n3303 585
R11273 gnd.n5070 gnd.n5069 585
R11274 gnd.n5071 gnd.n5070 585
R11275 gnd.n3312 gnd.n3311 585
R11276 gnd.n4986 gnd.n3311 585
R11277 gnd.n5029 gnd.n5028 585
R11278 gnd.n5028 gnd.n5027 585
R11279 gnd.n3316 gnd.n3315 585
R11280 gnd.n5020 gnd.n3316 585
R11281 gnd.n4871 gnd.n4870 585
R11282 gnd.n4870 gnd.n3334 585
R11283 gnd.n4874 gnd.n4869 585
R11284 gnd.n4869 gnd.n3332 585
R11285 gnd.n4875 gnd.n4868 585
R11286 gnd.n4868 gnd.n3338 585
R11287 gnd.n4876 gnd.n4867 585
R11288 gnd.n4867 gnd.n3342 585
R11289 gnd.n4866 gnd.n4864 585
R11290 gnd.n4866 gnd.n3351 585
R11291 gnd.n4880 gnd.n4863 585
R11292 gnd.n4863 gnd.n3349 585
R11293 gnd.n4881 gnd.n4862 585
R11294 gnd.n4862 gnd.n4861 585
R11295 gnd.n4882 gnd.n3362 585
R11296 gnd.n4940 gnd.n3362 585
R11297 gnd.n4859 gnd.n3370 585
R11298 gnd.n4930 gnd.n3370 585
R11299 gnd.n4886 gnd.n4858 585
R11300 gnd.n4858 gnd.n3376 585
R11301 gnd.n4887 gnd.n4857 585
R11302 gnd.n4857 gnd.n3384 585
R11303 gnd.n4888 gnd.n4856 585
R11304 gnd.n4856 gnd.n3381 585
R11305 gnd.n3401 gnd.n3391 585
R11306 gnd.n4903 gnd.n3391 585
R11307 gnd.n4893 gnd.n4892 585
R11308 gnd.n4895 gnd.n4893 585
R11309 gnd.n3400 gnd.n3399 585
R11310 gnd.n4808 gnd.n3399 585
R11311 gnd.n4852 gnd.n4851 585
R11312 gnd.n4851 gnd.n4850 585
R11313 gnd.n3404 gnd.n3403 585
R11314 gnd.n4843 gnd.n3404 585
R11315 gnd.n4772 gnd.n4771 585
R11316 gnd.n4771 gnd.n3421 585
R11317 gnd.n4773 gnd.n4770 585
R11318 gnd.n4770 gnd.n3418 585
R11319 gnd.n3444 gnd.n3442 585
R11320 gnd.n3442 gnd.n3425 585
R11321 gnd.n4778 gnd.n4777 585
R11322 gnd.n4779 gnd.n4778 585
R11323 gnd.n3443 gnd.n3441 585
R11324 gnd.n3441 gnd.t249 585
R11325 gnd.n4766 gnd.n4765 585
R11326 gnd.n4765 gnd.n3434 585
R11327 gnd.n4764 gnd.n3446 585
R11328 gnd.n4764 gnd.n4763 585
R11329 gnd.n4687 gnd.n3447 585
R11330 gnd.n4755 gnd.n3447 585
R11331 gnd.n4686 gnd.n3461 585
R11332 gnd.n4745 gnd.n3461 585
R11333 gnd.n4691 gnd.n4685 585
R11334 gnd.n4685 gnd.n3466 585
R11335 gnd.n4692 gnd.n4684 585
R11336 gnd.n4684 gnd.n3474 585
R11337 gnd.n4693 gnd.n4683 585
R11338 gnd.n4683 gnd.n3471 585
R11339 gnd.n3490 gnd.n3481 585
R11340 gnd.n4708 gnd.n3481 585
R11341 gnd.n4698 gnd.n4697 585
R11342 gnd.n4699 gnd.n4698 585
R11343 gnd.n3489 gnd.n3488 585
R11344 gnd.n4660 gnd.n3488 585
R11345 gnd.n4679 gnd.n4678 585
R11346 gnd.n4678 gnd.n4677 585
R11347 gnd.n3493 gnd.n3492 585
R11348 gnd.n3521 gnd.n3493 585
R11349 gnd.n4509 gnd.n4507 585
R11350 gnd.n4507 gnd.n4506 585
R11351 gnd.n4510 gnd.n3744 585
R11352 gnd.n4491 gnd.n3744 585
R11353 gnd.n4511 gnd.n3743 585
R11354 gnd.n4490 gnd.n3743 585
R11355 gnd.n4486 gnd.n3741 585
R11356 gnd.n4488 gnd.n4486 585
R11357 gnd.n4515 gnd.n3740 585
R11358 gnd.n3752 gnd.n3740 585
R11359 gnd.n4516 gnd.n3739 585
R11360 gnd.n4476 gnd.n3739 585
R11361 gnd.n4517 gnd.n3738 585
R11362 gnd.n4474 gnd.n3738 585
R11363 gnd.n5543 gnd.n5542 585
R11364 gnd.n5542 gnd.n2658 585
R11365 gnd.n5544 gnd.n5541 585
R11366 gnd.n5539 gnd.n2956 585
R11367 gnd.n5548 gnd.n2955 585
R11368 gnd.n5552 gnd.n2953 585
R11369 gnd.n5553 gnd.n2952 585
R11370 gnd.n2950 gnd.n2948 585
R11371 gnd.n5557 gnd.n2947 585
R11372 gnd.n5558 gnd.n2945 585
R11373 gnd.n5559 gnd.n2944 585
R11374 gnd.n2942 gnd.n2808 585
R11375 gnd.n2941 gnd.n2940 585
R11376 gnd.n2927 gnd.n2810 585
R11377 gnd.n2929 gnd.n2928 585
R11378 gnd.n2925 gnd.n2819 585
R11379 gnd.n2924 gnd.n2923 585
R11380 gnd.n2908 gnd.n2821 585
R11381 gnd.n2910 gnd.n2909 585
R11382 gnd.n2906 gnd.n2828 585
R11383 gnd.n2905 gnd.n2904 585
R11384 gnd.n2889 gnd.n2830 585
R11385 gnd.n2891 gnd.n2890 585
R11386 gnd.n2887 gnd.n2837 585
R11387 gnd.n2886 gnd.n2885 585
R11388 gnd.n2870 gnd.n2839 585
R11389 gnd.n2872 gnd.n2871 585
R11390 gnd.n2868 gnd.n2846 585
R11391 gnd.n2867 gnd.n2866 585
R11392 gnd.n2848 gnd.n2646 585
R11393 gnd.n6234 gnd.n695 476.536
R11394 gnd.n5430 gnd.n3155 468.476
R11395 gnd.n5433 gnd.n5432 468.476
R11396 gnd.n4666 gnd.n3495 468.476
R11397 gnd.n4675 gnd.n3497 468.476
R11398 gnd.n3554 gnd.t132 389.64
R11399 gnd.n3149 gnd.t108 389.64
R11400 gnd.n3556 gnd.t58 389.64
R11401 gnd.n5361 gnd.t141 389.64
R11402 gnd.n3729 gnd.t115 371.625
R11403 gnd.n7078 gnd.t102 371.625
R11404 gnd.n2812 gnd.t89 371.625
R11405 gnd.n3832 gnd.t112 371.625
R11406 gnd.n3069 gnd.t86 371.625
R11407 gnd.n3098 gnd.t54 371.625
R11408 gnd.n157 gnd.t50 371.625
R11409 gnd.n7156 gnd.t76 371.625
R11410 gnd.n4082 gnd.t147 371.625
R11411 gnd.n4058 gnd.t138 371.625
R11412 gnd.n3981 gnd.t128 371.625
R11413 gnd.n3708 gnd.t65 371.625
R11414 gnd.n3619 gnd.t105 371.625
R11415 gnd.n5549 gnd.t92 371.625
R11416 gnd.n6900 gnd.n6899 368.923
R11417 gnd.n1334 gnd.t46 323.425
R11418 gnd.n906 gnd.t69 323.425
R11419 gnd.n6687 gnd.n420 299.933
R11420 gnd.n6695 gnd.n420 299.933
R11421 gnd.n6696 gnd.n6695 299.933
R11422 gnd.n6697 gnd.n6696 299.933
R11423 gnd.n6697 gnd.n414 299.933
R11424 gnd.n6705 gnd.n414 299.933
R11425 gnd.n6706 gnd.n6705 299.933
R11426 gnd.n6707 gnd.n6706 299.933
R11427 gnd.n6707 gnd.n408 299.933
R11428 gnd.n6715 gnd.n408 299.933
R11429 gnd.n6716 gnd.n6715 299.933
R11430 gnd.n6717 gnd.n6716 299.933
R11431 gnd.n6717 gnd.n402 299.933
R11432 gnd.n6725 gnd.n402 299.933
R11433 gnd.n6726 gnd.n6725 299.933
R11434 gnd.n6727 gnd.n6726 299.933
R11435 gnd.n6727 gnd.n396 299.933
R11436 gnd.n6735 gnd.n396 299.933
R11437 gnd.n6736 gnd.n6735 299.933
R11438 gnd.n6737 gnd.n6736 299.933
R11439 gnd.n6737 gnd.n390 299.933
R11440 gnd.n6745 gnd.n390 299.933
R11441 gnd.n6746 gnd.n6745 299.933
R11442 gnd.n6747 gnd.n6746 299.933
R11443 gnd.n6747 gnd.n384 299.933
R11444 gnd.n6755 gnd.n384 299.933
R11445 gnd.n6756 gnd.n6755 299.933
R11446 gnd.n6757 gnd.n6756 299.933
R11447 gnd.n6757 gnd.n378 299.933
R11448 gnd.n6765 gnd.n378 299.933
R11449 gnd.n6766 gnd.n6765 299.933
R11450 gnd.n6767 gnd.n6766 299.933
R11451 gnd.n6767 gnd.n372 299.933
R11452 gnd.n6775 gnd.n372 299.933
R11453 gnd.n6776 gnd.n6775 299.933
R11454 gnd.n6777 gnd.n6776 299.933
R11455 gnd.n6777 gnd.n366 299.933
R11456 gnd.n6785 gnd.n366 299.933
R11457 gnd.n6786 gnd.n6785 299.933
R11458 gnd.n6787 gnd.n6786 299.933
R11459 gnd.n6787 gnd.n360 299.933
R11460 gnd.n6795 gnd.n360 299.933
R11461 gnd.n6796 gnd.n6795 299.933
R11462 gnd.n6797 gnd.n6796 299.933
R11463 gnd.n6797 gnd.n354 299.933
R11464 gnd.n6805 gnd.n354 299.933
R11465 gnd.n6806 gnd.n6805 299.933
R11466 gnd.n6807 gnd.n6806 299.933
R11467 gnd.n6807 gnd.n348 299.933
R11468 gnd.n6815 gnd.n348 299.933
R11469 gnd.n6816 gnd.n6815 299.933
R11470 gnd.n6817 gnd.n6816 299.933
R11471 gnd.n6817 gnd.n342 299.933
R11472 gnd.n6825 gnd.n342 299.933
R11473 gnd.n6826 gnd.n6825 299.933
R11474 gnd.n6827 gnd.n6826 299.933
R11475 gnd.n6827 gnd.n336 299.933
R11476 gnd.n6835 gnd.n336 299.933
R11477 gnd.n6836 gnd.n6835 299.933
R11478 gnd.n6837 gnd.n6836 299.933
R11479 gnd.n6837 gnd.n330 299.933
R11480 gnd.n6845 gnd.n330 299.933
R11481 gnd.n6846 gnd.n6845 299.933
R11482 gnd.n6847 gnd.n6846 299.933
R11483 gnd.n6847 gnd.n324 299.933
R11484 gnd.n6855 gnd.n324 299.933
R11485 gnd.n6856 gnd.n6855 299.933
R11486 gnd.n6857 gnd.n6856 299.933
R11487 gnd.n6857 gnd.n318 299.933
R11488 gnd.n6865 gnd.n318 299.933
R11489 gnd.n6866 gnd.n6865 299.933
R11490 gnd.n6867 gnd.n6866 299.933
R11491 gnd.n6867 gnd.n312 299.933
R11492 gnd.n6875 gnd.n312 299.933
R11493 gnd.n6876 gnd.n6875 299.933
R11494 gnd.n6877 gnd.n6876 299.933
R11495 gnd.n6877 gnd.n306 299.933
R11496 gnd.n6885 gnd.n306 299.933
R11497 gnd.n6886 gnd.n6885 299.933
R11498 gnd.n6887 gnd.n6886 299.933
R11499 gnd.n6887 gnd.n300 299.933
R11500 gnd.n6898 gnd.n300 299.933
R11501 gnd.n6899 gnd.n6898 299.933
R11502 gnd.n2184 gnd.n2158 289.615
R11503 gnd.n2152 gnd.n2126 289.615
R11504 gnd.n2120 gnd.n2094 289.615
R11505 gnd.n2089 gnd.n2063 289.615
R11506 gnd.n2057 gnd.n2031 289.615
R11507 gnd.n2025 gnd.n1999 289.615
R11508 gnd.n1993 gnd.n1967 289.615
R11509 gnd.n1962 gnd.n1936 289.615
R11510 gnd.n1408 gnd.t150 279.217
R11511 gnd.n932 gnd.t79 279.217
R11512 gnd.n3504 gnd.t64 260.649
R11513 gnd.n5353 gnd.t121 260.649
R11514 gnd.n4669 gnd.n4668 256.663
R11515 gnd.n4668 gnd.n3522 256.663
R11516 gnd.n4668 gnd.n3523 256.663
R11517 gnd.n4668 gnd.n3524 256.663
R11518 gnd.n4668 gnd.n3525 256.663
R11519 gnd.n4668 gnd.n3526 256.663
R11520 gnd.n4668 gnd.n3527 256.663
R11521 gnd.n4668 gnd.n3528 256.663
R11522 gnd.n4668 gnd.n3529 256.663
R11523 gnd.n4668 gnd.n3530 256.663
R11524 gnd.n4668 gnd.n3531 256.663
R11525 gnd.n4668 gnd.n3532 256.663
R11526 gnd.n4668 gnd.n3533 256.663
R11527 gnd.n4668 gnd.n3534 256.663
R11528 gnd.n4668 gnd.n3535 256.663
R11529 gnd.n4668 gnd.n3536 256.663
R11530 gnd.n4588 gnd.n4587 256.663
R11531 gnd.n4668 gnd.n3537 256.663
R11532 gnd.n4668 gnd.n3538 256.663
R11533 gnd.n4668 gnd.n3539 256.663
R11534 gnd.n4668 gnd.n3540 256.663
R11535 gnd.n4668 gnd.n3541 256.663
R11536 gnd.n4668 gnd.n3542 256.663
R11537 gnd.n4668 gnd.n3543 256.663
R11538 gnd.n4668 gnd.n3544 256.663
R11539 gnd.n4668 gnd.n3545 256.663
R11540 gnd.n4668 gnd.n3546 256.663
R11541 gnd.n4668 gnd.n3547 256.663
R11542 gnd.n4668 gnd.n3548 256.663
R11543 gnd.n4668 gnd.n3549 256.663
R11544 gnd.n4668 gnd.n3550 256.663
R11545 gnd.n4668 gnd.n3551 256.663
R11546 gnd.n4668 gnd.n3552 256.663
R11547 gnd.n4668 gnd.n4667 256.663
R11548 gnd.n5499 gnd.n2995 256.663
R11549 gnd.n5499 gnd.n2996 256.663
R11550 gnd.n5499 gnd.n2997 256.663
R11551 gnd.n5499 gnd.n2998 256.663
R11552 gnd.n5499 gnd.n2999 256.663
R11553 gnd.n5499 gnd.n3000 256.663
R11554 gnd.n5499 gnd.n3001 256.663
R11555 gnd.n5499 gnd.n3002 256.663
R11556 gnd.n5499 gnd.n3003 256.663
R11557 gnd.n5499 gnd.n3004 256.663
R11558 gnd.n5499 gnd.n3005 256.663
R11559 gnd.n5499 gnd.n3006 256.663
R11560 gnd.n5499 gnd.n3007 256.663
R11561 gnd.n5499 gnd.n3008 256.663
R11562 gnd.n5499 gnd.n3009 256.663
R11563 gnd.n5499 gnd.n3010 256.663
R11564 gnd.n3148 gnd.n3011 256.663
R11565 gnd.n5499 gnd.n2994 256.663
R11566 gnd.n5499 gnd.n2993 256.663
R11567 gnd.n5499 gnd.n2992 256.663
R11568 gnd.n5499 gnd.n2991 256.663
R11569 gnd.n5499 gnd.n2990 256.663
R11570 gnd.n5499 gnd.n2989 256.663
R11571 gnd.n5499 gnd.n2988 256.663
R11572 gnd.n5499 gnd.n2987 256.663
R11573 gnd.n5499 gnd.n2986 256.663
R11574 gnd.n5499 gnd.n2985 256.663
R11575 gnd.n5499 gnd.n2984 256.663
R11576 gnd.n5499 gnd.n2983 256.663
R11577 gnd.n5499 gnd.n2982 256.663
R11578 gnd.n5499 gnd.n2981 256.663
R11579 gnd.n5499 gnd.n2980 256.663
R11580 gnd.n5499 gnd.n2979 256.663
R11581 gnd.n5499 gnd.n2978 256.663
R11582 gnd.n4006 gnd.n2318 242.672
R11583 gnd.n4008 gnd.n2318 242.672
R11584 gnd.n4016 gnd.n2318 242.672
R11585 gnd.n4018 gnd.n2318 242.672
R11586 gnd.n4026 gnd.n2318 242.672
R11587 gnd.n4028 gnd.n2318 242.672
R11588 gnd.n4036 gnd.n2318 242.672
R11589 gnd.n4038 gnd.n2318 242.672
R11590 gnd.n4046 gnd.n2318 242.672
R11591 gnd.n3841 gnd.n3680 242.672
R11592 gnd.n3830 gnd.n3680 242.672
R11593 gnd.n3827 gnd.n3680 242.672
R11594 gnd.n3818 gnd.n3680 242.672
R11595 gnd.n3807 gnd.n3680 242.672
R11596 gnd.n3804 gnd.n3680 242.672
R11597 gnd.n3795 gnd.n3680 242.672
R11598 gnd.n3785 gnd.n3680 242.672
R11599 gnd.n3782 gnd.n3680 242.672
R11600 gnd.n2858 gnd.n2659 242.672
R11601 gnd.n2860 gnd.n2659 242.672
R11602 gnd.n2877 gnd.n2659 242.672
R11603 gnd.n2879 gnd.n2659 242.672
R11604 gnd.n2896 gnd.n2659 242.672
R11605 gnd.n2898 gnd.n2659 242.672
R11606 gnd.n2915 gnd.n2659 242.672
R11607 gnd.n2917 gnd.n2659 242.672
R11608 gnd.n2934 gnd.n2659 242.672
R11609 gnd.n7080 gnd.n94 242.672
R11610 gnd.n7076 gnd.n94 242.672
R11611 gnd.n7071 gnd.n94 242.672
R11612 gnd.n7068 gnd.n94 242.672
R11613 gnd.n7063 gnd.n94 242.672
R11614 gnd.n7060 gnd.n94 242.672
R11615 gnd.n7055 gnd.n94 242.672
R11616 gnd.n7052 gnd.n94 242.672
R11617 gnd.n7047 gnd.n94 242.672
R11618 gnd.n1462 gnd.n1461 242.672
R11619 gnd.n1462 gnd.n1372 242.672
R11620 gnd.n1462 gnd.n1373 242.672
R11621 gnd.n1462 gnd.n1374 242.672
R11622 gnd.n1462 gnd.n1375 242.672
R11623 gnd.n1462 gnd.n1376 242.672
R11624 gnd.n1462 gnd.n1377 242.672
R11625 gnd.n1462 gnd.n1378 242.672
R11626 gnd.n1462 gnd.n1379 242.672
R11627 gnd.n1462 gnd.n1380 242.672
R11628 gnd.n1462 gnd.n1381 242.672
R11629 gnd.n1462 gnd.n1382 242.672
R11630 gnd.n1463 gnd.n1462 242.672
R11631 gnd.n2316 gnd.n881 242.672
R11632 gnd.n2316 gnd.n880 242.672
R11633 gnd.n2316 gnd.n879 242.672
R11634 gnd.n2316 gnd.n878 242.672
R11635 gnd.n2316 gnd.n877 242.672
R11636 gnd.n2316 gnd.n876 242.672
R11637 gnd.n2316 gnd.n875 242.672
R11638 gnd.n2316 gnd.n874 242.672
R11639 gnd.n2316 gnd.n873 242.672
R11640 gnd.n2316 gnd.n872 242.672
R11641 gnd.n2316 gnd.n871 242.672
R11642 gnd.n2316 gnd.n870 242.672
R11643 gnd.n2316 gnd.n869 242.672
R11644 gnd.n1546 gnd.n1545 242.672
R11645 gnd.n1545 gnd.n1284 242.672
R11646 gnd.n1545 gnd.n1285 242.672
R11647 gnd.n1545 gnd.n1286 242.672
R11648 gnd.n1545 gnd.n1287 242.672
R11649 gnd.n1545 gnd.n1288 242.672
R11650 gnd.n1545 gnd.n1289 242.672
R11651 gnd.n1545 gnd.n1290 242.672
R11652 gnd.n2316 gnd.n882 242.672
R11653 gnd.n2316 gnd.n883 242.672
R11654 gnd.n2316 gnd.n884 242.672
R11655 gnd.n2316 gnd.n885 242.672
R11656 gnd.n2316 gnd.n886 242.672
R11657 gnd.n2316 gnd.n887 242.672
R11658 gnd.n2316 gnd.n888 242.672
R11659 gnd.n2316 gnd.n889 242.672
R11660 gnd.n4101 gnd.n2318 242.672
R11661 gnd.n4109 gnd.n2318 242.672
R11662 gnd.n4111 gnd.n2318 242.672
R11663 gnd.n4119 gnd.n2318 242.672
R11664 gnd.n4121 gnd.n2318 242.672
R11665 gnd.n4129 gnd.n2318 242.672
R11666 gnd.n4131 gnd.n2318 242.672
R11667 gnd.n4139 gnd.n2318 242.672
R11668 gnd.n4141 gnd.n2318 242.672
R11669 gnd.n4149 gnd.n2318 242.672
R11670 gnd.n4151 gnd.n2318 242.672
R11671 gnd.n4159 gnd.n2318 242.672
R11672 gnd.n4161 gnd.n2318 242.672
R11673 gnd.n4169 gnd.n2318 242.672
R11674 gnd.n4171 gnd.n2318 242.672
R11675 gnd.n4179 gnd.n2318 242.672
R11676 gnd.n4181 gnd.n2318 242.672
R11677 gnd.n4190 gnd.n2318 242.672
R11678 gnd.n4193 gnd.n2318 242.672
R11679 gnd.n4549 gnd.n3680 242.672
R11680 gnd.n3711 gnd.n3680 242.672
R11681 gnd.n4556 gnd.n3680 242.672
R11682 gnd.n3702 gnd.n3680 242.672
R11683 gnd.n4563 gnd.n3680 242.672
R11684 gnd.n3695 gnd.n3680 242.672
R11685 gnd.n4570 gnd.n3680 242.672
R11686 gnd.n3688 gnd.n3680 242.672
R11687 gnd.n4577 gnd.n3680 242.672
R11688 gnd.n4580 gnd.n3680 242.672
R11689 gnd.n3680 gnd.n3626 242.672
R11690 gnd.n4586 gnd.n3621 242.672
R11691 gnd.n3680 gnd.n3627 242.672
R11692 gnd.n3680 gnd.n3628 242.672
R11693 gnd.n3680 gnd.n3629 242.672
R11694 gnd.n3680 gnd.n3630 242.672
R11695 gnd.n3680 gnd.n3631 242.672
R11696 gnd.n3680 gnd.n3632 242.672
R11697 gnd.n3680 gnd.n3633 242.672
R11698 gnd.n3680 gnd.n3679 242.672
R11699 gnd.n3031 gnd.n2659 242.672
R11700 gnd.n3039 gnd.n2659 242.672
R11701 gnd.n3041 gnd.n2659 242.672
R11702 gnd.n3049 gnd.n2659 242.672
R11703 gnd.n3051 gnd.n2659 242.672
R11704 gnd.n3060 gnd.n2659 242.672
R11705 gnd.n3063 gnd.n2659 242.672
R11706 gnd.n3016 gnd.n2659 242.672
R11707 gnd.n3147 gnd.n3013 242.672
R11708 gnd.n3144 gnd.n2659 242.672
R11709 gnd.n3142 gnd.n2659 242.672
R11710 gnd.n3136 gnd.n2659 242.672
R11711 gnd.n3134 gnd.n2659 242.672
R11712 gnd.n3128 gnd.n2659 242.672
R11713 gnd.n3126 gnd.n2659 242.672
R11714 gnd.n3120 gnd.n2659 242.672
R11715 gnd.n3118 gnd.n2659 242.672
R11716 gnd.n3112 gnd.n2659 242.672
R11717 gnd.n3110 gnd.n2659 242.672
R11718 gnd.n3102 gnd.n2659 242.672
R11719 gnd.n154 gnd.n94 242.672
R11720 gnd.n7124 gnd.n94 242.672
R11721 gnd.n150 gnd.n94 242.672
R11722 gnd.n7131 gnd.n94 242.672
R11723 gnd.n143 gnd.n94 242.672
R11724 gnd.n7138 gnd.n94 242.672
R11725 gnd.n136 gnd.n94 242.672
R11726 gnd.n7145 gnd.n94 242.672
R11727 gnd.n129 gnd.n94 242.672
R11728 gnd.n7152 gnd.n94 242.672
R11729 gnd.n122 gnd.n94 242.672
R11730 gnd.n7162 gnd.n94 242.672
R11731 gnd.n115 gnd.n94 242.672
R11732 gnd.n7169 gnd.n94 242.672
R11733 gnd.n108 gnd.n94 242.672
R11734 gnd.n7176 gnd.n94 242.672
R11735 gnd.n101 gnd.n94 242.672
R11736 gnd.n7183 gnd.n94 242.672
R11737 gnd.n94 gnd.n93 242.672
R11738 gnd.n3890 gnd.n3889 242.672
R11739 gnd.n3890 gnd.n3758 242.672
R11740 gnd.n3890 gnd.n3759 242.672
R11741 gnd.n3890 gnd.n3760 242.672
R11742 gnd.n3890 gnd.n3761 242.672
R11743 gnd.n3890 gnd.n3762 242.672
R11744 gnd.n3890 gnd.n3763 242.672
R11745 gnd.n3890 gnd.n3764 242.672
R11746 gnd.n3890 gnd.n3765 242.672
R11747 gnd.n3890 gnd.n3766 242.672
R11748 gnd.n3890 gnd.n3768 242.672
R11749 gnd.n3890 gnd.n3769 242.672
R11750 gnd.n3890 gnd.n3770 242.672
R11751 gnd.n3890 gnd.n3772 242.672
R11752 gnd.n5540 gnd.n2658 242.672
R11753 gnd.n2954 gnd.n2658 242.672
R11754 gnd.n2951 gnd.n2658 242.672
R11755 gnd.n2946 gnd.n2658 242.672
R11756 gnd.n2943 gnd.n2658 242.672
R11757 gnd.n2809 gnd.n2658 242.672
R11758 gnd.n2926 gnd.n2658 242.672
R11759 gnd.n2820 gnd.n2658 242.672
R11760 gnd.n2907 gnd.n2658 242.672
R11761 gnd.n2829 gnd.n2658 242.672
R11762 gnd.n2888 gnd.n2658 242.672
R11763 gnd.n2838 gnd.n2658 242.672
R11764 gnd.n2869 gnd.n2658 242.672
R11765 gnd.n2847 gnd.n2658 242.672
R11766 gnd.n90 gnd.n86 240.244
R11767 gnd.n7185 gnd.n7184 240.244
R11768 gnd.n7182 gnd.n95 240.244
R11769 gnd.n7178 gnd.n7177 240.244
R11770 gnd.n7175 gnd.n102 240.244
R11771 gnd.n7171 gnd.n7170 240.244
R11772 gnd.n7168 gnd.n109 240.244
R11773 gnd.n7164 gnd.n7163 240.244
R11774 gnd.n7161 gnd.n116 240.244
R11775 gnd.n7154 gnd.n7153 240.244
R11776 gnd.n7151 gnd.n123 240.244
R11777 gnd.n7147 gnd.n7146 240.244
R11778 gnd.n7144 gnd.n130 240.244
R11779 gnd.n7140 gnd.n7139 240.244
R11780 gnd.n7137 gnd.n137 240.244
R11781 gnd.n7133 gnd.n7132 240.244
R11782 gnd.n7130 gnd.n144 240.244
R11783 gnd.n7126 gnd.n7125 240.244
R11784 gnd.n7123 gnd.n151 240.244
R11785 gnd.n5567 gnd.n2668 240.244
R11786 gnd.n5567 gnd.n2680 240.244
R11787 gnd.n5592 gnd.n2680 240.244
R11788 gnd.n5592 gnd.n2801 240.244
R11789 gnd.n2801 gnd.n2795 240.244
R11790 gnd.n2795 gnd.n2773 240.244
R11791 gnd.n5586 gnd.n2773 240.244
R11792 gnd.n5586 gnd.n2764 240.244
R11793 gnd.n5583 gnd.n2764 240.244
R11794 gnd.n5583 gnd.n2756 240.244
R11795 gnd.n2756 gnd.n2748 240.244
R11796 gnd.n2748 gnd.n2736 240.244
R11797 gnd.n5679 gnd.n2736 240.244
R11798 gnd.n5679 gnd.n2737 240.244
R11799 gnd.n2737 gnd.n2711 240.244
R11800 gnd.n2711 gnd.n2705 240.244
R11801 gnd.n5687 gnd.n2705 240.244
R11802 gnd.n5687 gnd.n234 240.244
R11803 gnd.n5715 gnd.n234 240.244
R11804 gnd.n5715 gnd.n2720 240.244
R11805 gnd.n2725 gnd.n2720 240.244
R11806 gnd.n5710 gnd.n2725 240.244
R11807 gnd.n5710 gnd.n5709 240.244
R11808 gnd.n5709 gnd.n256 240.244
R11809 gnd.n256 gnd.n249 240.244
R11810 gnd.n5701 gnd.n249 240.244
R11811 gnd.n5701 gnd.n221 240.244
R11812 gnd.n6950 gnd.n221 240.244
R11813 gnd.n6950 gnd.n212 240.244
R11814 gnd.n6946 gnd.n212 240.244
R11815 gnd.n6946 gnd.n204 240.244
R11816 gnd.n6942 gnd.n204 240.244
R11817 gnd.n6942 gnd.n195 240.244
R11818 gnd.n6916 gnd.n195 240.244
R11819 gnd.n6916 gnd.n189 240.244
R11820 gnd.n6931 gnd.n189 240.244
R11821 gnd.n6931 gnd.n180 240.244
R11822 gnd.n6927 gnd.n180 240.244
R11823 gnd.n6927 gnd.n170 240.244
R11824 gnd.n170 gnd.n161 240.244
R11825 gnd.n7115 gnd.n161 240.244
R11826 gnd.n7115 gnd.n82 240.244
R11827 gnd.n3032 gnd.n3027 240.244
R11828 gnd.n3038 gnd.n3027 240.244
R11829 gnd.n3042 gnd.n3040 240.244
R11830 gnd.n3048 gnd.n3023 240.244
R11831 gnd.n3052 gnd.n3050 240.244
R11832 gnd.n3059 gnd.n3019 240.244
R11833 gnd.n3062 gnd.n3061 240.244
R11834 gnd.n3064 gnd.n3017 240.244
R11835 gnd.n3145 gnd.n3143 240.244
R11836 gnd.n3141 gnd.n3073 240.244
R11837 gnd.n3137 gnd.n3135 240.244
R11838 gnd.n3133 gnd.n3079 240.244
R11839 gnd.n3129 gnd.n3127 240.244
R11840 gnd.n3125 gnd.n3085 240.244
R11841 gnd.n3121 gnd.n3119 240.244
R11842 gnd.n3117 gnd.n3091 240.244
R11843 gnd.n3113 gnd.n3111 240.244
R11844 gnd.n3109 gnd.n3097 240.244
R11845 gnd.n5778 gnd.n2673 240.244
R11846 gnd.n5774 gnd.n2673 240.244
R11847 gnd.n5774 gnd.n2678 240.244
R11848 gnd.n2793 gnd.n2678 240.244
R11849 gnd.n2793 gnd.n2771 240.244
R11850 gnd.n5616 gnd.n2771 240.244
R11851 gnd.n5616 gnd.n2766 240.244
R11852 gnd.n5624 gnd.n2766 240.244
R11853 gnd.n5624 gnd.n2767 240.244
R11854 gnd.n2767 gnd.n2746 240.244
R11855 gnd.n5669 gnd.n2746 240.244
R11856 gnd.n5669 gnd.n2742 240.244
R11857 gnd.n5677 gnd.n2742 240.244
R11858 gnd.n5677 gnd.n2708 240.244
R11859 gnd.n5745 gnd.n2708 240.244
R11860 gnd.n5746 gnd.n5745 240.244
R11861 gnd.n5746 gnd.n231 240.244
R11862 gnd.n6981 gnd.n231 240.244
R11863 gnd.n6981 gnd.n232 240.244
R11864 gnd.n5731 gnd.n232 240.244
R11865 gnd.n5731 gnd.n5728 240.244
R11866 gnd.n5728 gnd.n2722 240.244
R11867 gnd.n2722 gnd.n252 240.244
R11868 gnd.n6962 gnd.n252 240.244
R11869 gnd.n6964 gnd.n6962 240.244
R11870 gnd.n6964 gnd.n222 240.244
R11871 gnd.n6988 gnd.n222 240.244
R11872 gnd.n6988 gnd.n210 240.244
R11873 gnd.n6998 gnd.n210 240.244
R11874 gnd.n6998 gnd.n206 240.244
R11875 gnd.n7004 gnd.n206 240.244
R11876 gnd.n7004 gnd.n194 240.244
R11877 gnd.n7014 gnd.n194 240.244
R11878 gnd.n7014 gnd.n190 240.244
R11879 gnd.n7020 gnd.n190 240.244
R11880 gnd.n7020 gnd.n178 240.244
R11881 gnd.n7030 gnd.n178 240.244
R11882 gnd.n7030 gnd.n172 240.244
R11883 gnd.n7038 gnd.n172 240.244
R11884 gnd.n7038 gnd.n174 240.244
R11885 gnd.n174 gnd.n85 240.244
R11886 gnd.n7192 gnd.n85 240.244
R11887 gnd.n3634 gnd.n2533 240.244
R11888 gnd.n3678 gnd.n3635 240.244
R11889 gnd.n3674 gnd.n3673 240.244
R11890 gnd.n3670 gnd.n3669 240.244
R11891 gnd.n3666 gnd.n3665 240.244
R11892 gnd.n3662 gnd.n3661 240.244
R11893 gnd.n3658 gnd.n3657 240.244
R11894 gnd.n3654 gnd.n3653 240.244
R11895 gnd.n4581 gnd.n3625 240.244
R11896 gnd.n4579 gnd.n4578 240.244
R11897 gnd.n4576 gnd.n3682 240.244
R11898 gnd.n4572 gnd.n4571 240.244
R11899 gnd.n4569 gnd.n3689 240.244
R11900 gnd.n4565 gnd.n4564 240.244
R11901 gnd.n4562 gnd.n3696 240.244
R11902 gnd.n4558 gnd.n4557 240.244
R11903 gnd.n4555 gnd.n3703 240.244
R11904 gnd.n4551 gnd.n4550 240.244
R11905 gnd.n3978 gnd.n2319 240.244
R11906 gnd.n3978 gnd.n2330 240.244
R11907 gnd.n4240 gnd.n2330 240.244
R11908 gnd.n4240 gnd.n2342 240.244
R11909 gnd.n4236 gnd.n2342 240.244
R11910 gnd.n4236 gnd.n2353 240.244
R11911 gnd.n4228 gnd.n2353 240.244
R11912 gnd.n4228 gnd.n2364 240.244
R11913 gnd.n4224 gnd.n2364 240.244
R11914 gnd.n4224 gnd.n2375 240.244
R11915 gnd.n3966 gnd.n2375 240.244
R11916 gnd.n3966 gnd.n2385 240.244
R11917 gnd.n4287 gnd.n2385 240.244
R11918 gnd.n4287 gnd.n2396 240.244
R11919 gnd.n4294 gnd.n2396 240.244
R11920 gnd.n4294 gnd.n2407 240.244
R11921 gnd.n4305 gnd.n2407 240.244
R11922 gnd.n4305 gnd.n2416 240.244
R11923 gnd.n3942 gnd.n2416 240.244
R11924 gnd.n3942 gnd.n2426 240.244
R11925 gnd.n4313 gnd.n2426 240.244
R11926 gnd.n4313 gnd.n2434 240.244
R11927 gnd.n4328 gnd.n2434 240.244
R11928 gnd.n4328 gnd.n2443 240.244
R11929 gnd.n4338 gnd.n2443 240.244
R11930 gnd.n4338 gnd.n2451 240.244
R11931 gnd.n3926 gnd.n2451 240.244
R11932 gnd.n3926 gnd.n2461 240.244
R11933 gnd.n4398 gnd.n2461 240.244
R11934 gnd.n4398 gnd.n2472 240.244
R11935 gnd.n4404 gnd.n2472 240.244
R11936 gnd.n4404 gnd.n2482 240.244
R11937 gnd.n4414 gnd.n2482 240.244
R11938 gnd.n4414 gnd.n2493 240.244
R11939 gnd.n3905 gnd.n2493 240.244
R11940 gnd.n3905 gnd.n2503 240.244
R11941 gnd.n4422 gnd.n2503 240.244
R11942 gnd.n4422 gnd.n2514 240.244
R11943 gnd.n4429 gnd.n2514 240.244
R11944 gnd.n4429 gnd.n2525 240.244
R11945 gnd.n4542 gnd.n2525 240.244
R11946 gnd.n4542 gnd.n2535 240.244
R11947 gnd.n4102 gnd.n4097 240.244
R11948 gnd.n4108 gnd.n4097 240.244
R11949 gnd.n4112 gnd.n4110 240.244
R11950 gnd.n4118 gnd.n4093 240.244
R11951 gnd.n4122 gnd.n4120 240.244
R11952 gnd.n4128 gnd.n4089 240.244
R11953 gnd.n4132 gnd.n4130 240.244
R11954 gnd.n4138 gnd.n4085 240.244
R11955 gnd.n4142 gnd.n4140 240.244
R11956 gnd.n4148 gnd.n4078 240.244
R11957 gnd.n4152 gnd.n4150 240.244
R11958 gnd.n4158 gnd.n4074 240.244
R11959 gnd.n4162 gnd.n4160 240.244
R11960 gnd.n4168 gnd.n4070 240.244
R11961 gnd.n4172 gnd.n4170 240.244
R11962 gnd.n4178 gnd.n4066 240.244
R11963 gnd.n4182 gnd.n4180 240.244
R11964 gnd.n4189 gnd.n4062 240.244
R11965 gnd.n4192 gnd.n4191 240.244
R11966 gnd.n6054 gnd.n2324 240.244
R11967 gnd.n6050 gnd.n2324 240.244
R11968 gnd.n6050 gnd.n2329 240.244
R11969 gnd.n6042 gnd.n2329 240.244
R11970 gnd.n6042 gnd.n2345 240.244
R11971 gnd.n6038 gnd.n2345 240.244
R11972 gnd.n6038 gnd.n2351 240.244
R11973 gnd.n6030 gnd.n2351 240.244
R11974 gnd.n6030 gnd.n2367 240.244
R11975 gnd.n6026 gnd.n2367 240.244
R11976 gnd.n6026 gnd.n2373 240.244
R11977 gnd.n6018 gnd.n2373 240.244
R11978 gnd.n6018 gnd.n2388 240.244
R11979 gnd.n6014 gnd.n2388 240.244
R11980 gnd.n6014 gnd.n2394 240.244
R11981 gnd.n6006 gnd.n2394 240.244
R11982 gnd.n6006 gnd.n2410 240.244
R11983 gnd.n6001 gnd.n2410 240.244
R11984 gnd.n6001 gnd.n2414 240.244
R11985 gnd.n5993 gnd.n2414 240.244
R11986 gnd.n5993 gnd.n2429 240.244
R11987 gnd.n5988 gnd.n2429 240.244
R11988 gnd.n5988 gnd.n2432 240.244
R11989 gnd.n5980 gnd.n2432 240.244
R11990 gnd.n5980 gnd.n2446 240.244
R11991 gnd.n5975 gnd.n2446 240.244
R11992 gnd.n5975 gnd.n2449 240.244
R11993 gnd.n5967 gnd.n2449 240.244
R11994 gnd.n5967 gnd.n2464 240.244
R11995 gnd.n5963 gnd.n2464 240.244
R11996 gnd.n5963 gnd.n2470 240.244
R11997 gnd.n5955 gnd.n2470 240.244
R11998 gnd.n5955 gnd.n2485 240.244
R11999 gnd.n5951 gnd.n2485 240.244
R12000 gnd.n5951 gnd.n2491 240.244
R12001 gnd.n5943 gnd.n2491 240.244
R12002 gnd.n5943 gnd.n2506 240.244
R12003 gnd.n5939 gnd.n2506 240.244
R12004 gnd.n5939 gnd.n2512 240.244
R12005 gnd.n5931 gnd.n2512 240.244
R12006 gnd.n5931 gnd.n2528 240.244
R12007 gnd.n5927 gnd.n2528 240.244
R12008 gnd.n2315 gnd.n891 240.244
R12009 gnd.n2308 gnd.n2307 240.244
R12010 gnd.n2305 gnd.n2304 240.244
R12011 gnd.n2301 gnd.n2300 240.244
R12012 gnd.n2297 gnd.n2296 240.244
R12013 gnd.n2293 gnd.n2292 240.244
R12014 gnd.n2289 gnd.n2288 240.244
R12015 gnd.n2285 gnd.n2284 240.244
R12016 gnd.n1557 gnd.n1269 240.244
R12017 gnd.n1567 gnd.n1269 240.244
R12018 gnd.n1567 gnd.n1260 240.244
R12019 gnd.n1260 gnd.n1249 240.244
R12020 gnd.n1588 gnd.n1249 240.244
R12021 gnd.n1588 gnd.n1243 240.244
R12022 gnd.n1598 gnd.n1243 240.244
R12023 gnd.n1598 gnd.n1232 240.244
R12024 gnd.n1232 gnd.n1224 240.244
R12025 gnd.n1616 gnd.n1224 240.244
R12026 gnd.n1617 gnd.n1616 240.244
R12027 gnd.n1617 gnd.n1209 240.244
R12028 gnd.n1619 gnd.n1209 240.244
R12029 gnd.n1619 gnd.n1195 240.244
R12030 gnd.n1661 gnd.n1195 240.244
R12031 gnd.n1662 gnd.n1661 240.244
R12032 gnd.n1665 gnd.n1662 240.244
R12033 gnd.n1665 gnd.n1150 240.244
R12034 gnd.n1190 gnd.n1150 240.244
R12035 gnd.n1190 gnd.n1160 240.244
R12036 gnd.n1675 gnd.n1160 240.244
R12037 gnd.n1675 gnd.n1181 240.244
R12038 gnd.n1685 gnd.n1181 240.244
R12039 gnd.n1685 gnd.n1091 240.244
R12040 gnd.n1730 gnd.n1091 240.244
R12041 gnd.n1730 gnd.n1077 240.244
R12042 gnd.n1752 gnd.n1077 240.244
R12043 gnd.n1753 gnd.n1752 240.244
R12044 gnd.n1753 gnd.n1064 240.244
R12045 gnd.n1064 gnd.n1053 240.244
R12046 gnd.n1784 gnd.n1053 240.244
R12047 gnd.n1785 gnd.n1784 240.244
R12048 gnd.n1786 gnd.n1785 240.244
R12049 gnd.n1786 gnd.n1038 240.244
R12050 gnd.n1817 gnd.n1038 240.244
R12051 gnd.n1817 gnd.n1024 240.244
R12052 gnd.n1839 gnd.n1024 240.244
R12053 gnd.n1840 gnd.n1839 240.244
R12054 gnd.n1840 gnd.n1011 240.244
R12055 gnd.n1011 gnd.n1000 240.244
R12056 gnd.n1871 gnd.n1000 240.244
R12057 gnd.n1872 gnd.n1871 240.244
R12058 gnd.n1873 gnd.n1872 240.244
R12059 gnd.n1873 gnd.n984 240.244
R12060 gnd.n984 gnd.n983 240.244
R12061 gnd.n983 gnd.n970 240.244
R12062 gnd.n1928 gnd.n970 240.244
R12063 gnd.n1929 gnd.n1928 240.244
R12064 gnd.n1929 gnd.n957 240.244
R12065 gnd.n957 gnd.n947 240.244
R12066 gnd.n2216 gnd.n947 240.244
R12067 gnd.n2219 gnd.n2216 240.244
R12068 gnd.n2219 gnd.n2218 240.244
R12069 gnd.n1547 gnd.n1282 240.244
R12070 gnd.n1303 gnd.n1282 240.244
R12071 gnd.n1306 gnd.n1305 240.244
R12072 gnd.n1313 gnd.n1312 240.244
R12073 gnd.n1316 gnd.n1315 240.244
R12074 gnd.n1323 gnd.n1322 240.244
R12075 gnd.n1326 gnd.n1325 240.244
R12076 gnd.n1333 gnd.n1332 240.244
R12077 gnd.n1555 gnd.n1279 240.244
R12078 gnd.n1279 gnd.n1258 240.244
R12079 gnd.n1578 gnd.n1258 240.244
R12080 gnd.n1578 gnd.n1252 240.244
R12081 gnd.n1586 gnd.n1252 240.244
R12082 gnd.n1586 gnd.n1254 240.244
R12083 gnd.n1254 gnd.n1230 240.244
R12084 gnd.n1608 gnd.n1230 240.244
R12085 gnd.n1608 gnd.n1226 240.244
R12086 gnd.n1614 gnd.n1226 240.244
R12087 gnd.n1614 gnd.n1208 240.244
R12088 gnd.n1639 gnd.n1208 240.244
R12089 gnd.n1639 gnd.n1203 240.244
R12090 gnd.n1651 gnd.n1203 240.244
R12091 gnd.n1651 gnd.n1204 240.244
R12092 gnd.n1647 gnd.n1204 240.244
R12093 gnd.n1647 gnd.n1152 240.244
R12094 gnd.n1699 gnd.n1152 240.244
R12095 gnd.n1699 gnd.n1153 240.244
R12096 gnd.n1695 gnd.n1153 240.244
R12097 gnd.n1695 gnd.n1159 240.244
R12098 gnd.n1179 gnd.n1159 240.244
R12099 gnd.n1179 gnd.n1089 240.244
R12100 gnd.n1734 gnd.n1089 240.244
R12101 gnd.n1734 gnd.n1084 240.244
R12102 gnd.n1742 gnd.n1084 240.244
R12103 gnd.n1742 gnd.n1085 240.244
R12104 gnd.n1085 gnd.n1062 240.244
R12105 gnd.n1774 gnd.n1062 240.244
R12106 gnd.n1774 gnd.n1057 240.244
R12107 gnd.n1782 gnd.n1057 240.244
R12108 gnd.n1782 gnd.n1058 240.244
R12109 gnd.n1058 gnd.n1036 240.244
R12110 gnd.n1821 gnd.n1036 240.244
R12111 gnd.n1821 gnd.n1031 240.244
R12112 gnd.n1829 gnd.n1031 240.244
R12113 gnd.n1829 gnd.n1032 240.244
R12114 gnd.n1032 gnd.n1009 240.244
R12115 gnd.n1861 gnd.n1009 240.244
R12116 gnd.n1861 gnd.n1004 240.244
R12117 gnd.n1869 gnd.n1004 240.244
R12118 gnd.n1869 gnd.n1005 240.244
R12119 gnd.n1005 gnd.n982 240.244
R12120 gnd.n1910 gnd.n982 240.244
R12121 gnd.n1910 gnd.n977 240.244
R12122 gnd.n1918 gnd.n977 240.244
R12123 gnd.n1918 gnd.n978 240.244
R12124 gnd.n978 gnd.n955 240.244
R12125 gnd.n2204 gnd.n955 240.244
R12126 gnd.n2204 gnd.n950 240.244
R12127 gnd.n2214 gnd.n950 240.244
R12128 gnd.n2214 gnd.n951 240.244
R12129 gnd.n951 gnd.n890 240.244
R12130 gnd.n910 gnd.n868 240.244
R12131 gnd.n2275 gnd.n2274 240.244
R12132 gnd.n2271 gnd.n2270 240.244
R12133 gnd.n2267 gnd.n2266 240.244
R12134 gnd.n2263 gnd.n2262 240.244
R12135 gnd.n2259 gnd.n2258 240.244
R12136 gnd.n2255 gnd.n2254 240.244
R12137 gnd.n2251 gnd.n2250 240.244
R12138 gnd.n2247 gnd.n2246 240.244
R12139 gnd.n2243 gnd.n2242 240.244
R12140 gnd.n2239 gnd.n2238 240.244
R12141 gnd.n2235 gnd.n2234 240.244
R12142 gnd.n2231 gnd.n2230 240.244
R12143 gnd.n1470 gnd.n1367 240.244
R12144 gnd.n1470 gnd.n1360 240.244
R12145 gnd.n1481 gnd.n1360 240.244
R12146 gnd.n1481 gnd.n1356 240.244
R12147 gnd.n1487 gnd.n1356 240.244
R12148 gnd.n1487 gnd.n1348 240.244
R12149 gnd.n1497 gnd.n1348 240.244
R12150 gnd.n1497 gnd.n1343 240.244
R12151 gnd.n1533 gnd.n1343 240.244
R12152 gnd.n1533 gnd.n1344 240.244
R12153 gnd.n1344 gnd.n1291 240.244
R12154 gnd.n1528 gnd.n1291 240.244
R12155 gnd.n1528 gnd.n1527 240.244
R12156 gnd.n1527 gnd.n1270 240.244
R12157 gnd.n1523 gnd.n1270 240.244
R12158 gnd.n1523 gnd.n1261 240.244
R12159 gnd.n1520 gnd.n1261 240.244
R12160 gnd.n1520 gnd.n1519 240.244
R12161 gnd.n1519 gnd.n1244 240.244
R12162 gnd.n1515 gnd.n1244 240.244
R12163 gnd.n1515 gnd.n1233 240.244
R12164 gnd.n1233 gnd.n1214 240.244
R12165 gnd.n1628 gnd.n1214 240.244
R12166 gnd.n1628 gnd.n1210 240.244
R12167 gnd.n1636 gnd.n1210 240.244
R12168 gnd.n1636 gnd.n1201 240.244
R12169 gnd.n1201 gnd.n1137 240.244
R12170 gnd.n1708 gnd.n1137 240.244
R12171 gnd.n1708 gnd.n1138 240.244
R12172 gnd.n1149 gnd.n1138 240.244
R12173 gnd.n1184 gnd.n1149 240.244
R12174 gnd.n1187 gnd.n1184 240.244
R12175 gnd.n1187 gnd.n1161 240.244
R12176 gnd.n1174 gnd.n1161 240.244
R12177 gnd.n1174 gnd.n1171 240.244
R12178 gnd.n1171 gnd.n1092 240.244
R12179 gnd.n1729 gnd.n1092 240.244
R12180 gnd.n1729 gnd.n1082 240.244
R12181 gnd.n1725 gnd.n1082 240.244
R12182 gnd.n1725 gnd.n1076 240.244
R12183 gnd.n1722 gnd.n1076 240.244
R12184 gnd.n1722 gnd.n1065 240.244
R12185 gnd.n1719 gnd.n1065 240.244
R12186 gnd.n1719 gnd.n1043 240.244
R12187 gnd.n1795 gnd.n1043 240.244
R12188 gnd.n1795 gnd.n1039 240.244
R12189 gnd.n1816 gnd.n1039 240.244
R12190 gnd.n1816 gnd.n1029 240.244
R12191 gnd.n1812 gnd.n1029 240.244
R12192 gnd.n1812 gnd.n1023 240.244
R12193 gnd.n1809 gnd.n1023 240.244
R12194 gnd.n1809 gnd.n1012 240.244
R12195 gnd.n1806 gnd.n1012 240.244
R12196 gnd.n1806 gnd.n989 240.244
R12197 gnd.n1882 gnd.n989 240.244
R12198 gnd.n1882 gnd.n985 240.244
R12199 gnd.n1907 gnd.n985 240.244
R12200 gnd.n1907 gnd.n976 240.244
R12201 gnd.n1903 gnd.n976 240.244
R12202 gnd.n1903 gnd.n969 240.244
R12203 gnd.n1899 gnd.n969 240.244
R12204 gnd.n1899 gnd.n958 240.244
R12205 gnd.n1896 gnd.n958 240.244
R12206 gnd.n1896 gnd.n939 240.244
R12207 gnd.n2226 gnd.n939 240.244
R12208 gnd.n1384 gnd.n1383 240.244
R12209 gnd.n1455 gnd.n1383 240.244
R12210 gnd.n1453 gnd.n1452 240.244
R12211 gnd.n1449 gnd.n1448 240.244
R12212 gnd.n1445 gnd.n1444 240.244
R12213 gnd.n1441 gnd.n1440 240.244
R12214 gnd.n1437 gnd.n1436 240.244
R12215 gnd.n1433 gnd.n1432 240.244
R12216 gnd.n1429 gnd.n1428 240.244
R12217 gnd.n1425 gnd.n1424 240.244
R12218 gnd.n1421 gnd.n1420 240.244
R12219 gnd.n1417 gnd.n1416 240.244
R12220 gnd.n1413 gnd.n1371 240.244
R12221 gnd.n1473 gnd.n1365 240.244
R12222 gnd.n1473 gnd.n1361 240.244
R12223 gnd.n1479 gnd.n1361 240.244
R12224 gnd.n1479 gnd.n1354 240.244
R12225 gnd.n1489 gnd.n1354 240.244
R12226 gnd.n1489 gnd.n1350 240.244
R12227 gnd.n1495 gnd.n1350 240.244
R12228 gnd.n1495 gnd.n1341 240.244
R12229 gnd.n1535 gnd.n1341 240.244
R12230 gnd.n1535 gnd.n1292 240.244
R12231 gnd.n1543 gnd.n1292 240.244
R12232 gnd.n1543 gnd.n1293 240.244
R12233 gnd.n1293 gnd.n1271 240.244
R12234 gnd.n1564 gnd.n1271 240.244
R12235 gnd.n1564 gnd.n1263 240.244
R12236 gnd.n1575 gnd.n1263 240.244
R12237 gnd.n1575 gnd.n1264 240.244
R12238 gnd.n1264 gnd.n1245 240.244
R12239 gnd.n1595 gnd.n1245 240.244
R12240 gnd.n1595 gnd.n1235 240.244
R12241 gnd.n1605 gnd.n1235 240.244
R12242 gnd.n1605 gnd.n1216 240.244
R12243 gnd.n1626 gnd.n1216 240.244
R12244 gnd.n1626 gnd.n1218 240.244
R12245 gnd.n1218 gnd.n1199 240.244
R12246 gnd.n1654 gnd.n1199 240.244
R12247 gnd.n1654 gnd.n1141 240.244
R12248 gnd.n1706 gnd.n1141 240.244
R12249 gnd.n1706 gnd.n1142 240.244
R12250 gnd.n1702 gnd.n1142 240.244
R12251 gnd.n1702 gnd.n1148 240.244
R12252 gnd.n1163 gnd.n1148 240.244
R12253 gnd.n1692 gnd.n1163 240.244
R12254 gnd.n1692 gnd.n1164 240.244
R12255 gnd.n1688 gnd.n1164 240.244
R12256 gnd.n1688 gnd.n1170 240.244
R12257 gnd.n1170 gnd.n1081 240.244
R12258 gnd.n1745 gnd.n1081 240.244
R12259 gnd.n1745 gnd.n1074 240.244
R12260 gnd.n1756 gnd.n1074 240.244
R12261 gnd.n1756 gnd.n1067 240.244
R12262 gnd.n1771 gnd.n1067 240.244
R12263 gnd.n1771 gnd.n1068 240.244
R12264 gnd.n1068 gnd.n1046 240.244
R12265 gnd.n1793 gnd.n1046 240.244
R12266 gnd.n1793 gnd.n1047 240.244
R12267 gnd.n1047 gnd.n1028 240.244
R12268 gnd.n1832 gnd.n1028 240.244
R12269 gnd.n1832 gnd.n1021 240.244
R12270 gnd.n1843 gnd.n1021 240.244
R12271 gnd.n1843 gnd.n1014 240.244
R12272 gnd.n1858 gnd.n1014 240.244
R12273 gnd.n1858 gnd.n1015 240.244
R12274 gnd.n1015 gnd.n992 240.244
R12275 gnd.n1880 gnd.n992 240.244
R12276 gnd.n1880 gnd.n994 240.244
R12277 gnd.n994 gnd.n974 240.244
R12278 gnd.n1921 gnd.n974 240.244
R12279 gnd.n1921 gnd.n967 240.244
R12280 gnd.n1932 gnd.n967 240.244
R12281 gnd.n1932 gnd.n960 240.244
R12282 gnd.n2201 gnd.n960 240.244
R12283 gnd.n2201 gnd.n961 240.244
R12284 gnd.n961 gnd.n942 240.244
R12285 gnd.n2224 gnd.n942 240.244
R12286 gnd.n7046 gnd.n7045 240.244
R12287 gnd.n7051 gnd.n7048 240.244
R12288 gnd.n7054 gnd.n7053 240.244
R12289 gnd.n7059 gnd.n7056 240.244
R12290 gnd.n7062 gnd.n7061 240.244
R12291 gnd.n7067 gnd.n7064 240.244
R12292 gnd.n7070 gnd.n7069 240.244
R12293 gnd.n7075 gnd.n7072 240.244
R12294 gnd.n7081 gnd.n7077 240.244
R12295 gnd.n5565 gnd.n2669 240.244
R12296 gnd.n5565 gnd.n2681 240.244
R12297 gnd.n5595 gnd.n2681 240.244
R12298 gnd.n5595 gnd.n2796 240.244
R12299 gnd.n5602 gnd.n2796 240.244
R12300 gnd.n5602 gnd.n2774 240.244
R12301 gnd.n2774 gnd.n2762 240.244
R12302 gnd.n5626 gnd.n2762 240.244
R12303 gnd.n5626 gnd.n2757 240.244
R12304 gnd.n5639 gnd.n2757 240.244
R12305 gnd.n5639 gnd.n2749 240.244
R12306 gnd.n5632 gnd.n2749 240.244
R12307 gnd.n5632 gnd.n2739 240.244
R12308 gnd.n2739 gnd.n2712 240.244
R12309 gnd.n5743 gnd.n2712 240.244
R12310 gnd.n5743 gnd.n2706 240.244
R12311 gnd.n2717 gnd.n2706 240.244
R12312 gnd.n2717 gnd.n235 240.244
R12313 gnd.n2718 gnd.n235 240.244
R12314 gnd.n5733 gnd.n2718 240.244
R12315 gnd.n5733 gnd.n2719 240.244
R12316 gnd.n2719 gnd.n54 240.244
R12317 gnd.n55 gnd.n54 240.244
R12318 gnd.n56 gnd.n55 240.244
R12319 gnd.n250 gnd.n56 240.244
R12320 gnd.n250 gnd.n59 240.244
R12321 gnd.n60 gnd.n59 240.244
R12322 gnd.n61 gnd.n60 240.244
R12323 gnd.n213 gnd.n61 240.244
R12324 gnd.n213 gnd.n64 240.244
R12325 gnd.n65 gnd.n64 240.244
R12326 gnd.n66 gnd.n65 240.244
R12327 gnd.n196 gnd.n66 240.244
R12328 gnd.n196 gnd.n69 240.244
R12329 gnd.n70 gnd.n69 240.244
R12330 gnd.n71 gnd.n70 240.244
R12331 gnd.n181 gnd.n71 240.244
R12332 gnd.n181 gnd.n74 240.244
R12333 gnd.n75 gnd.n74 240.244
R12334 gnd.n76 gnd.n75 240.244
R12335 gnd.n79 gnd.n76 240.244
R12336 gnd.n7194 gnd.n79 240.244
R12337 gnd.n2861 gnd.n2859 240.244
R12338 gnd.n2876 gnd.n2842 240.244
R12339 gnd.n2880 gnd.n2878 240.244
R12340 gnd.n2895 gnd.n2833 240.244
R12341 gnd.n2899 gnd.n2897 240.244
R12342 gnd.n2914 gnd.n2824 240.244
R12343 gnd.n2918 gnd.n2916 240.244
R12344 gnd.n2933 gnd.n2815 240.244
R12345 gnd.n2936 gnd.n2935 240.244
R12346 gnd.n2683 gnd.n2671 240.244
R12347 gnd.n5772 gnd.n2683 240.244
R12348 gnd.n5772 gnd.n2684 240.244
R12349 gnd.n2689 gnd.n2684 240.244
R12350 gnd.n2690 gnd.n2689 240.244
R12351 gnd.n2691 gnd.n2690 240.244
R12352 gnd.n2775 gnd.n2691 240.244
R12353 gnd.n2775 gnd.n2694 240.244
R12354 gnd.n2695 gnd.n2694 240.244
R12355 gnd.n2696 gnd.n2695 240.244
R12356 gnd.n5667 gnd.n2696 240.244
R12357 gnd.n5667 gnd.n2699 240.244
R12358 gnd.n2700 gnd.n2699 240.244
R12359 gnd.n2701 gnd.n2700 240.244
R12360 gnd.n2703 gnd.n2701 240.244
R12361 gnd.n5748 gnd.n2703 240.244
R12362 gnd.n5748 gnd.n237 240.244
R12363 gnd.n6979 gnd.n237 240.244
R12364 gnd.n6979 gnd.n238 240.244
R12365 gnd.n243 gnd.n238 240.244
R12366 gnd.n244 gnd.n243 240.244
R12367 gnd.n245 gnd.n244 240.244
R12368 gnd.n5707 gnd.n245 240.244
R12369 gnd.n5707 gnd.n248 240.244
R12370 gnd.n6966 gnd.n248 240.244
R12371 gnd.n6966 gnd.n219 240.244
R12372 gnd.n6990 gnd.n219 240.244
R12373 gnd.n6990 gnd.n215 240.244
R12374 gnd.n6996 gnd.n215 240.244
R12375 gnd.n6996 gnd.n202 240.244
R12376 gnd.n7006 gnd.n202 240.244
R12377 gnd.n7006 gnd.n198 240.244
R12378 gnd.n7012 gnd.n198 240.244
R12379 gnd.n7012 gnd.n187 240.244
R12380 gnd.n7022 gnd.n187 240.244
R12381 gnd.n7022 gnd.n183 240.244
R12382 gnd.n7028 gnd.n183 240.244
R12383 gnd.n7028 gnd.n168 240.244
R12384 gnd.n7040 gnd.n168 240.244
R12385 gnd.n7040 gnd.n163 240.244
R12386 gnd.n7113 gnd.n163 240.244
R12387 gnd.n7113 gnd.n84 240.244
R12388 gnd.n3781 gnd.n2538 240.244
R12389 gnd.n3784 gnd.n3783 240.244
R12390 gnd.n3794 gnd.n3786 240.244
R12391 gnd.n3797 gnd.n3796 240.244
R12392 gnd.n3806 gnd.n3805 240.244
R12393 gnd.n3817 gnd.n3808 240.244
R12394 gnd.n3820 gnd.n3819 240.244
R12395 gnd.n3829 gnd.n3828 240.244
R12396 gnd.n3840 gnd.n3831 240.244
R12397 gnd.n4246 gnd.n2320 240.244
R12398 gnd.n4246 gnd.n2331 240.244
R12399 gnd.n4242 gnd.n2331 240.244
R12400 gnd.n4242 gnd.n2343 240.244
R12401 gnd.n4234 gnd.n2343 240.244
R12402 gnd.n4234 gnd.n2354 240.244
R12403 gnd.n4230 gnd.n2354 240.244
R12404 gnd.n4230 gnd.n2365 240.244
R12405 gnd.n4222 gnd.n2365 240.244
R12406 gnd.n4222 gnd.n2376 240.244
R12407 gnd.n4279 gnd.n2376 240.244
R12408 gnd.n4279 gnd.n2386 240.244
R12409 gnd.n4285 gnd.n2386 240.244
R12410 gnd.n4285 gnd.n2397 240.244
R12411 gnd.n4296 gnd.n2397 240.244
R12412 gnd.n4296 gnd.n2408 240.244
R12413 gnd.n4303 gnd.n2408 240.244
R12414 gnd.n4303 gnd.n2417 240.244
R12415 gnd.n4351 gnd.n2417 240.244
R12416 gnd.n4351 gnd.n2427 240.244
R12417 gnd.n3946 gnd.n2427 240.244
R12418 gnd.n3946 gnd.n2435 240.244
R12419 gnd.n3949 gnd.n2435 240.244
R12420 gnd.n3949 gnd.n2444 240.244
R12421 gnd.n4340 gnd.n2444 240.244
R12422 gnd.n4340 gnd.n2452 240.244
R12423 gnd.n4390 gnd.n2452 240.244
R12424 gnd.n4390 gnd.n2462 240.244
R12425 gnd.n4396 gnd.n2462 240.244
R12426 gnd.n4396 gnd.n2473 240.244
R12427 gnd.n4406 gnd.n2473 240.244
R12428 gnd.n4406 gnd.n2483 240.244
R12429 gnd.n4412 gnd.n2483 240.244
R12430 gnd.n4412 gnd.n2494 240.244
R12431 gnd.n4440 gnd.n2494 240.244
R12432 gnd.n4440 gnd.n2504 240.244
R12433 gnd.n3910 gnd.n2504 240.244
R12434 gnd.n3910 gnd.n2515 240.244
R12435 gnd.n4431 gnd.n2515 240.244
R12436 gnd.n4431 gnd.n2526 240.244
R12437 gnd.n4540 gnd.n2526 240.244
R12438 gnd.n4540 gnd.n2536 240.244
R12439 gnd.n4009 gnd.n4007 240.244
R12440 gnd.n4015 gnd.n3996 240.244
R12441 gnd.n4019 gnd.n4017 240.244
R12442 gnd.n4025 gnd.n3992 240.244
R12443 gnd.n4029 gnd.n4027 240.244
R12444 gnd.n4035 gnd.n3988 240.244
R12445 gnd.n4039 gnd.n4037 240.244
R12446 gnd.n4045 gnd.n3984 240.244
R12447 gnd.n4048 gnd.n4047 240.244
R12448 gnd.n2333 gnd.n2322 240.244
R12449 gnd.n6048 gnd.n2333 240.244
R12450 gnd.n6048 gnd.n2334 240.244
R12451 gnd.n6044 gnd.n2334 240.244
R12452 gnd.n6044 gnd.n2340 240.244
R12453 gnd.n6036 gnd.n2340 240.244
R12454 gnd.n6036 gnd.n2356 240.244
R12455 gnd.n6032 gnd.n2356 240.244
R12456 gnd.n6032 gnd.n2362 240.244
R12457 gnd.n6024 gnd.n2362 240.244
R12458 gnd.n6024 gnd.n2378 240.244
R12459 gnd.n6020 gnd.n2378 240.244
R12460 gnd.n6020 gnd.n2384 240.244
R12461 gnd.n6012 gnd.n2384 240.244
R12462 gnd.n6012 gnd.n2399 240.244
R12463 gnd.n6008 gnd.n2399 240.244
R12464 gnd.n6008 gnd.n2405 240.244
R12465 gnd.n5999 gnd.n2405 240.244
R12466 gnd.n5999 gnd.n2419 240.244
R12467 gnd.n5995 gnd.n2419 240.244
R12468 gnd.n5995 gnd.n2425 240.244
R12469 gnd.n5986 gnd.n2425 240.244
R12470 gnd.n5986 gnd.n2436 240.244
R12471 gnd.n5982 gnd.n2436 240.244
R12472 gnd.n5982 gnd.n2441 240.244
R12473 gnd.n5973 gnd.n2441 240.244
R12474 gnd.n5973 gnd.n2454 240.244
R12475 gnd.n5969 gnd.n2454 240.244
R12476 gnd.n5969 gnd.n2460 240.244
R12477 gnd.n5961 gnd.n2460 240.244
R12478 gnd.n5961 gnd.n2474 240.244
R12479 gnd.n5957 gnd.n2474 240.244
R12480 gnd.n5957 gnd.n2480 240.244
R12481 gnd.n5949 gnd.n2480 240.244
R12482 gnd.n5949 gnd.n2496 240.244
R12483 gnd.n5945 gnd.n2496 240.244
R12484 gnd.n5945 gnd.n2502 240.244
R12485 gnd.n5937 gnd.n2502 240.244
R12486 gnd.n5937 gnd.n2517 240.244
R12487 gnd.n5933 gnd.n2517 240.244
R12488 gnd.n5933 gnd.n2523 240.244
R12489 gnd.n5925 gnd.n2523 240.244
R12490 gnd.n6233 gnd.n694 240.244
R12491 gnd.n6237 gnd.n694 240.244
R12492 gnd.n6237 gnd.n690 240.244
R12493 gnd.n6243 gnd.n690 240.244
R12494 gnd.n6243 gnd.n688 240.244
R12495 gnd.n6247 gnd.n688 240.244
R12496 gnd.n6247 gnd.n684 240.244
R12497 gnd.n6253 gnd.n684 240.244
R12498 gnd.n6253 gnd.n682 240.244
R12499 gnd.n6257 gnd.n682 240.244
R12500 gnd.n6257 gnd.n678 240.244
R12501 gnd.n6263 gnd.n678 240.244
R12502 gnd.n6263 gnd.n676 240.244
R12503 gnd.n6267 gnd.n676 240.244
R12504 gnd.n6267 gnd.n672 240.244
R12505 gnd.n6273 gnd.n672 240.244
R12506 gnd.n6273 gnd.n670 240.244
R12507 gnd.n6277 gnd.n670 240.244
R12508 gnd.n6277 gnd.n666 240.244
R12509 gnd.n6283 gnd.n666 240.244
R12510 gnd.n6283 gnd.n664 240.244
R12511 gnd.n6287 gnd.n664 240.244
R12512 gnd.n6287 gnd.n660 240.244
R12513 gnd.n6293 gnd.n660 240.244
R12514 gnd.n6293 gnd.n658 240.244
R12515 gnd.n6297 gnd.n658 240.244
R12516 gnd.n6297 gnd.n654 240.244
R12517 gnd.n6303 gnd.n654 240.244
R12518 gnd.n6303 gnd.n652 240.244
R12519 gnd.n6307 gnd.n652 240.244
R12520 gnd.n6307 gnd.n648 240.244
R12521 gnd.n6313 gnd.n648 240.244
R12522 gnd.n6313 gnd.n646 240.244
R12523 gnd.n6317 gnd.n646 240.244
R12524 gnd.n6317 gnd.n642 240.244
R12525 gnd.n6323 gnd.n642 240.244
R12526 gnd.n6323 gnd.n640 240.244
R12527 gnd.n6327 gnd.n640 240.244
R12528 gnd.n6327 gnd.n636 240.244
R12529 gnd.n6333 gnd.n636 240.244
R12530 gnd.n6333 gnd.n634 240.244
R12531 gnd.n6337 gnd.n634 240.244
R12532 gnd.n6337 gnd.n630 240.244
R12533 gnd.n6343 gnd.n630 240.244
R12534 gnd.n6343 gnd.n628 240.244
R12535 gnd.n6347 gnd.n628 240.244
R12536 gnd.n6347 gnd.n624 240.244
R12537 gnd.n6353 gnd.n624 240.244
R12538 gnd.n6353 gnd.n622 240.244
R12539 gnd.n6357 gnd.n622 240.244
R12540 gnd.n6357 gnd.n618 240.244
R12541 gnd.n6363 gnd.n618 240.244
R12542 gnd.n6363 gnd.n616 240.244
R12543 gnd.n6367 gnd.n616 240.244
R12544 gnd.n6367 gnd.n612 240.244
R12545 gnd.n6373 gnd.n612 240.244
R12546 gnd.n6373 gnd.n610 240.244
R12547 gnd.n6377 gnd.n610 240.244
R12548 gnd.n6377 gnd.n606 240.244
R12549 gnd.n6383 gnd.n606 240.244
R12550 gnd.n6383 gnd.n604 240.244
R12551 gnd.n6387 gnd.n604 240.244
R12552 gnd.n6387 gnd.n600 240.244
R12553 gnd.n6393 gnd.n600 240.244
R12554 gnd.n6393 gnd.n598 240.244
R12555 gnd.n6397 gnd.n598 240.244
R12556 gnd.n6397 gnd.n594 240.244
R12557 gnd.n6403 gnd.n594 240.244
R12558 gnd.n6403 gnd.n592 240.244
R12559 gnd.n6407 gnd.n592 240.244
R12560 gnd.n6407 gnd.n588 240.244
R12561 gnd.n6413 gnd.n588 240.244
R12562 gnd.n6413 gnd.n586 240.244
R12563 gnd.n6417 gnd.n586 240.244
R12564 gnd.n6417 gnd.n582 240.244
R12565 gnd.n6423 gnd.n582 240.244
R12566 gnd.n6423 gnd.n580 240.244
R12567 gnd.n6427 gnd.n580 240.244
R12568 gnd.n6427 gnd.n576 240.244
R12569 gnd.n6433 gnd.n576 240.244
R12570 gnd.n6433 gnd.n574 240.244
R12571 gnd.n6437 gnd.n574 240.244
R12572 gnd.n6437 gnd.n570 240.244
R12573 gnd.n6443 gnd.n570 240.244
R12574 gnd.n6443 gnd.n568 240.244
R12575 gnd.n6447 gnd.n568 240.244
R12576 gnd.n6447 gnd.n564 240.244
R12577 gnd.n6453 gnd.n564 240.244
R12578 gnd.n6453 gnd.n562 240.244
R12579 gnd.n6457 gnd.n562 240.244
R12580 gnd.n6457 gnd.n558 240.244
R12581 gnd.n6463 gnd.n558 240.244
R12582 gnd.n6463 gnd.n556 240.244
R12583 gnd.n6467 gnd.n556 240.244
R12584 gnd.n6467 gnd.n552 240.244
R12585 gnd.n6473 gnd.n552 240.244
R12586 gnd.n6473 gnd.n550 240.244
R12587 gnd.n6477 gnd.n550 240.244
R12588 gnd.n6477 gnd.n546 240.244
R12589 gnd.n6483 gnd.n546 240.244
R12590 gnd.n6483 gnd.n544 240.244
R12591 gnd.n6487 gnd.n544 240.244
R12592 gnd.n6487 gnd.n540 240.244
R12593 gnd.n6493 gnd.n540 240.244
R12594 gnd.n6493 gnd.n538 240.244
R12595 gnd.n6497 gnd.n538 240.244
R12596 gnd.n6497 gnd.n534 240.244
R12597 gnd.n6503 gnd.n534 240.244
R12598 gnd.n6503 gnd.n532 240.244
R12599 gnd.n6507 gnd.n532 240.244
R12600 gnd.n6507 gnd.n528 240.244
R12601 gnd.n6513 gnd.n528 240.244
R12602 gnd.n6513 gnd.n526 240.244
R12603 gnd.n6517 gnd.n526 240.244
R12604 gnd.n6517 gnd.n522 240.244
R12605 gnd.n6523 gnd.n522 240.244
R12606 gnd.n6523 gnd.n520 240.244
R12607 gnd.n6527 gnd.n520 240.244
R12608 gnd.n6527 gnd.n516 240.244
R12609 gnd.n6533 gnd.n516 240.244
R12610 gnd.n6533 gnd.n514 240.244
R12611 gnd.n6537 gnd.n514 240.244
R12612 gnd.n6537 gnd.n510 240.244
R12613 gnd.n6543 gnd.n510 240.244
R12614 gnd.n6543 gnd.n508 240.244
R12615 gnd.n6547 gnd.n508 240.244
R12616 gnd.n6547 gnd.n504 240.244
R12617 gnd.n6553 gnd.n504 240.244
R12618 gnd.n6553 gnd.n502 240.244
R12619 gnd.n6557 gnd.n502 240.244
R12620 gnd.n6557 gnd.n498 240.244
R12621 gnd.n6563 gnd.n498 240.244
R12622 gnd.n6563 gnd.n496 240.244
R12623 gnd.n6567 gnd.n496 240.244
R12624 gnd.n6567 gnd.n492 240.244
R12625 gnd.n6573 gnd.n492 240.244
R12626 gnd.n6573 gnd.n490 240.244
R12627 gnd.n6577 gnd.n490 240.244
R12628 gnd.n6577 gnd.n486 240.244
R12629 gnd.n6583 gnd.n486 240.244
R12630 gnd.n6583 gnd.n484 240.244
R12631 gnd.n6587 gnd.n484 240.244
R12632 gnd.n6587 gnd.n480 240.244
R12633 gnd.n6593 gnd.n480 240.244
R12634 gnd.n6593 gnd.n478 240.244
R12635 gnd.n6597 gnd.n478 240.244
R12636 gnd.n6597 gnd.n474 240.244
R12637 gnd.n6603 gnd.n474 240.244
R12638 gnd.n6603 gnd.n472 240.244
R12639 gnd.n6607 gnd.n472 240.244
R12640 gnd.n6607 gnd.n468 240.244
R12641 gnd.n6613 gnd.n468 240.244
R12642 gnd.n6613 gnd.n466 240.244
R12643 gnd.n6617 gnd.n466 240.244
R12644 gnd.n6617 gnd.n462 240.244
R12645 gnd.n6623 gnd.n462 240.244
R12646 gnd.n6623 gnd.n460 240.244
R12647 gnd.n6627 gnd.n460 240.244
R12648 gnd.n6627 gnd.n456 240.244
R12649 gnd.n6633 gnd.n456 240.244
R12650 gnd.n6633 gnd.n454 240.244
R12651 gnd.n6637 gnd.n454 240.244
R12652 gnd.n6637 gnd.n450 240.244
R12653 gnd.n6643 gnd.n450 240.244
R12654 gnd.n6643 gnd.n448 240.244
R12655 gnd.n6647 gnd.n448 240.244
R12656 gnd.n6647 gnd.n444 240.244
R12657 gnd.n6653 gnd.n444 240.244
R12658 gnd.n6653 gnd.n442 240.244
R12659 gnd.n6657 gnd.n442 240.244
R12660 gnd.n6657 gnd.n438 240.244
R12661 gnd.n6663 gnd.n438 240.244
R12662 gnd.n6663 gnd.n436 240.244
R12663 gnd.n6667 gnd.n436 240.244
R12664 gnd.n6667 gnd.n432 240.244
R12665 gnd.n6673 gnd.n432 240.244
R12666 gnd.n6673 gnd.n430 240.244
R12667 gnd.n6677 gnd.n430 240.244
R12668 gnd.n6677 gnd.n426 240.244
R12669 gnd.n6684 gnd.n426 240.244
R12670 gnd.n6684 gnd.n424 240.244
R12671 gnd.n6688 gnd.n421 240.244
R12672 gnd.n6694 gnd.n421 240.244
R12673 gnd.n6694 gnd.n419 240.244
R12674 gnd.n6698 gnd.n419 240.244
R12675 gnd.n6698 gnd.n415 240.244
R12676 gnd.n6704 gnd.n415 240.244
R12677 gnd.n6704 gnd.n413 240.244
R12678 gnd.n6708 gnd.n413 240.244
R12679 gnd.n6708 gnd.n409 240.244
R12680 gnd.n6714 gnd.n409 240.244
R12681 gnd.n6714 gnd.n407 240.244
R12682 gnd.n6718 gnd.n407 240.244
R12683 gnd.n6718 gnd.n403 240.244
R12684 gnd.n6724 gnd.n403 240.244
R12685 gnd.n6724 gnd.n401 240.244
R12686 gnd.n6728 gnd.n401 240.244
R12687 gnd.n6728 gnd.n397 240.244
R12688 gnd.n6734 gnd.n397 240.244
R12689 gnd.n6734 gnd.n395 240.244
R12690 gnd.n6738 gnd.n395 240.244
R12691 gnd.n6738 gnd.n391 240.244
R12692 gnd.n6744 gnd.n391 240.244
R12693 gnd.n6744 gnd.n389 240.244
R12694 gnd.n6748 gnd.n389 240.244
R12695 gnd.n6748 gnd.n385 240.244
R12696 gnd.n6754 gnd.n385 240.244
R12697 gnd.n6754 gnd.n383 240.244
R12698 gnd.n6758 gnd.n383 240.244
R12699 gnd.n6758 gnd.n379 240.244
R12700 gnd.n6764 gnd.n379 240.244
R12701 gnd.n6764 gnd.n377 240.244
R12702 gnd.n6768 gnd.n377 240.244
R12703 gnd.n6768 gnd.n373 240.244
R12704 gnd.n6774 gnd.n373 240.244
R12705 gnd.n6774 gnd.n371 240.244
R12706 gnd.n6778 gnd.n371 240.244
R12707 gnd.n6778 gnd.n367 240.244
R12708 gnd.n6784 gnd.n367 240.244
R12709 gnd.n6784 gnd.n365 240.244
R12710 gnd.n6788 gnd.n365 240.244
R12711 gnd.n6788 gnd.n361 240.244
R12712 gnd.n6794 gnd.n361 240.244
R12713 gnd.n6794 gnd.n359 240.244
R12714 gnd.n6798 gnd.n359 240.244
R12715 gnd.n6798 gnd.n355 240.244
R12716 gnd.n6804 gnd.n355 240.244
R12717 gnd.n6804 gnd.n353 240.244
R12718 gnd.n6808 gnd.n353 240.244
R12719 gnd.n6808 gnd.n349 240.244
R12720 gnd.n6814 gnd.n349 240.244
R12721 gnd.n6814 gnd.n347 240.244
R12722 gnd.n6818 gnd.n347 240.244
R12723 gnd.n6818 gnd.n343 240.244
R12724 gnd.n6824 gnd.n343 240.244
R12725 gnd.n6824 gnd.n341 240.244
R12726 gnd.n6828 gnd.n341 240.244
R12727 gnd.n6828 gnd.n337 240.244
R12728 gnd.n6834 gnd.n337 240.244
R12729 gnd.n6834 gnd.n335 240.244
R12730 gnd.n6838 gnd.n335 240.244
R12731 gnd.n6838 gnd.n331 240.244
R12732 gnd.n6844 gnd.n331 240.244
R12733 gnd.n6844 gnd.n329 240.244
R12734 gnd.n6848 gnd.n329 240.244
R12735 gnd.n6848 gnd.n325 240.244
R12736 gnd.n6854 gnd.n325 240.244
R12737 gnd.n6854 gnd.n323 240.244
R12738 gnd.n6858 gnd.n323 240.244
R12739 gnd.n6858 gnd.n319 240.244
R12740 gnd.n6864 gnd.n319 240.244
R12741 gnd.n6864 gnd.n317 240.244
R12742 gnd.n6868 gnd.n317 240.244
R12743 gnd.n6868 gnd.n313 240.244
R12744 gnd.n6874 gnd.n313 240.244
R12745 gnd.n6874 gnd.n311 240.244
R12746 gnd.n6878 gnd.n311 240.244
R12747 gnd.n6878 gnd.n307 240.244
R12748 gnd.n6884 gnd.n307 240.244
R12749 gnd.n6884 gnd.n305 240.244
R12750 gnd.n6888 gnd.n305 240.244
R12751 gnd.n6888 gnd.n301 240.244
R12752 gnd.n6897 gnd.n301 240.244
R12753 gnd.n6897 gnd.n298 240.244
R12754 gnd.n6901 gnd.n298 240.244
R12755 gnd.n6057 gnd.n866 240.244
R12756 gnd.n4249 gnd.n866 240.244
R12757 gnd.n4249 gnd.n3976 240.244
R12758 gnd.n4255 gnd.n3976 240.244
R12759 gnd.n4256 gnd.n4255 240.244
R12760 gnd.n4257 gnd.n4256 240.244
R12761 gnd.n4257 gnd.n3972 240.244
R12762 gnd.n4263 gnd.n3972 240.244
R12763 gnd.n4264 gnd.n4263 240.244
R12764 gnd.n4265 gnd.n4264 240.244
R12765 gnd.n4265 gnd.n3967 240.244
R12766 gnd.n4276 gnd.n3967 240.244
R12767 gnd.n4276 gnd.n3968 240.244
R12768 gnd.n4272 gnd.n3968 240.244
R12769 gnd.n4272 gnd.n3938 240.244
R12770 gnd.n4360 gnd.n3938 240.244
R12771 gnd.n4360 gnd.n4359 240.244
R12772 gnd.n4359 gnd.n4358 240.244
R12773 gnd.n4358 gnd.n4355 240.244
R12774 gnd.n4355 gnd.n4354 240.244
R12775 gnd.n4354 gnd.n3939 240.244
R12776 gnd.n4316 gnd.n3939 240.244
R12777 gnd.n4325 gnd.n4316 240.244
R12778 gnd.n4325 gnd.n4322 240.244
R12779 gnd.n4322 gnd.n4319 240.244
R12780 gnd.n4319 gnd.n4318 240.244
R12781 gnd.n4318 gnd.n3927 240.244
R12782 gnd.n4387 gnd.n3927 240.244
R12783 gnd.n4387 gnd.n3928 240.244
R12784 gnd.n4383 gnd.n3928 240.244
R12785 gnd.n4383 gnd.n4382 240.244
R12786 gnd.n4382 gnd.n4381 240.244
R12787 gnd.n4381 gnd.n4369 240.244
R12788 gnd.n4377 gnd.n4369 240.244
R12789 gnd.n4377 gnd.n3903 240.244
R12790 gnd.n4443 gnd.n3903 240.244
R12791 gnd.n4444 gnd.n4443 240.244
R12792 gnd.n4445 gnd.n4444 240.244
R12793 gnd.n4445 gnd.n3899 240.244
R12794 gnd.n4451 gnd.n3899 240.244
R12795 gnd.n4452 gnd.n4451 240.244
R12796 gnd.n4453 gnd.n4452 240.244
R12797 gnd.n4453 gnd.n3895 240.244
R12798 gnd.n4460 gnd.n3895 240.244
R12799 gnd.n4461 gnd.n4460 240.244
R12800 gnd.n4465 gnd.n4461 240.244
R12801 gnd.n4465 gnd.n3891 240.244
R12802 gnd.n4471 gnd.n3891 240.244
R12803 gnd.n4471 gnd.n3757 240.244
R12804 gnd.n4478 gnd.n3757 240.244
R12805 gnd.n4478 gnd.n3753 240.244
R12806 gnd.n4484 gnd.n3753 240.244
R12807 gnd.n4484 gnd.n3751 240.244
R12808 gnd.n4493 gnd.n3751 240.244
R12809 gnd.n4493 gnd.n3746 240.244
R12810 gnd.n4504 gnd.n3746 240.244
R12811 gnd.n4504 gnd.n3747 240.244
R12812 gnd.n4500 gnd.n3747 240.244
R12813 gnd.n4500 gnd.n3479 240.244
R12814 gnd.n4710 gnd.n3479 240.244
R12815 gnd.n4710 gnd.n3475 240.244
R12816 gnd.n4716 gnd.n3475 240.244
R12817 gnd.n4716 gnd.n3459 240.244
R12818 gnd.n4747 gnd.n3459 240.244
R12819 gnd.n4747 gnd.n3455 240.244
R12820 gnd.n4753 gnd.n3455 240.244
R12821 gnd.n4753 gnd.n3433 240.244
R12822 gnd.n4788 gnd.n3433 240.244
R12823 gnd.n4788 gnd.n3429 240.244
R12824 gnd.n4794 gnd.n3429 240.244
R12825 gnd.n4794 gnd.n3417 240.244
R12826 gnd.n4833 gnd.n3417 240.244
R12827 gnd.n4833 gnd.n3412 240.244
R12828 gnd.n4841 gnd.n3412 240.244
R12829 gnd.n4841 gnd.n3413 240.244
R12830 gnd.n3413 gnd.n3389 240.244
R12831 gnd.n4905 gnd.n3389 240.244
R12832 gnd.n4905 gnd.n3385 240.244
R12833 gnd.n4911 gnd.n3385 240.244
R12834 gnd.n4911 gnd.n3368 240.244
R12835 gnd.n4932 gnd.n3368 240.244
R12836 gnd.n4932 gnd.n3364 240.244
R12837 gnd.n4938 gnd.n3364 240.244
R12838 gnd.n4938 gnd.n3347 240.244
R12839 gnd.n4965 gnd.n3347 240.244
R12840 gnd.n4965 gnd.n3343 240.244
R12841 gnd.n4971 gnd.n3343 240.244
R12842 gnd.n4971 gnd.n3330 240.244
R12843 gnd.n5010 gnd.n3330 240.244
R12844 gnd.n5010 gnd.n3325 240.244
R12845 gnd.n5018 gnd.n3325 240.244
R12846 gnd.n5018 gnd.n3326 240.244
R12847 gnd.n3326 gnd.n3301 240.244
R12848 gnd.n5081 gnd.n3301 240.244
R12849 gnd.n5081 gnd.n3297 240.244
R12850 gnd.n5087 gnd.n3297 240.244
R12851 gnd.n5087 gnd.n3281 240.244
R12852 gnd.n5108 gnd.n3281 240.244
R12853 gnd.n5108 gnd.n3277 240.244
R12854 gnd.n5114 gnd.n3277 240.244
R12855 gnd.n5114 gnd.n3259 240.244
R12856 gnd.n5141 gnd.n3259 240.244
R12857 gnd.n5141 gnd.n3255 240.244
R12858 gnd.n5147 gnd.n3255 240.244
R12859 gnd.n5147 gnd.n3242 240.244
R12860 gnd.n5186 gnd.n3242 240.244
R12861 gnd.n5186 gnd.n3237 240.244
R12862 gnd.n5194 gnd.n3237 240.244
R12863 gnd.n5194 gnd.n3238 240.244
R12864 gnd.n3238 gnd.n3214 240.244
R12865 gnd.n5234 gnd.n3214 240.244
R12866 gnd.n5234 gnd.n3210 240.244
R12867 gnd.n5240 gnd.n3210 240.244
R12868 gnd.n5240 gnd.n3194 240.244
R12869 gnd.n5277 gnd.n3194 240.244
R12870 gnd.n5277 gnd.n3189 240.244
R12871 gnd.n5285 gnd.n3189 240.244
R12872 gnd.n5285 gnd.n3190 240.244
R12873 gnd.n3190 gnd.n3165 240.244
R12874 gnd.n5330 gnd.n3165 240.244
R12875 gnd.n5330 gnd.n3161 240.244
R12876 gnd.n5336 gnd.n3161 240.244
R12877 gnd.n5336 gnd.n2976 240.244
R12878 gnd.n5501 gnd.n2976 240.244
R12879 gnd.n5501 gnd.n2972 240.244
R12880 gnd.n5507 gnd.n2972 240.244
R12881 gnd.n5507 gnd.n2964 240.244
R12882 gnd.n5524 gnd.n2964 240.244
R12883 gnd.n5524 gnd.n2960 240.244
R12884 gnd.n5531 gnd.n2960 240.244
R12885 gnd.n5531 gnd.n2650 240.244
R12886 gnd.n5793 gnd.n2650 240.244
R12887 gnd.n5793 gnd.n2651 240.244
R12888 gnd.n5789 gnd.n2651 240.244
R12889 gnd.n5789 gnd.n2657 240.244
R12890 gnd.n5785 gnd.n2657 240.244
R12891 gnd.n5785 gnd.n2660 240.244
R12892 gnd.n5781 gnd.n2660 240.244
R12893 gnd.n5781 gnd.n2666 240.244
R12894 gnd.n2782 gnd.n2666 240.244
R12895 gnd.n2788 gnd.n2782 240.244
R12896 gnd.n2789 gnd.n2788 240.244
R12897 gnd.n5605 gnd.n2789 240.244
R12898 gnd.n5605 gnd.n2777 240.244
R12899 gnd.n5613 gnd.n2777 240.244
R12900 gnd.n5613 gnd.n2778 240.244
R12901 gnd.n2778 gnd.n2755 240.244
R12902 gnd.n5642 gnd.n2755 240.244
R12903 gnd.n5642 gnd.n2750 240.244
R12904 gnd.n5665 gnd.n2750 240.244
R12905 gnd.n5665 gnd.n2751 240.244
R12906 gnd.n5661 gnd.n2751 240.244
R12907 gnd.n5661 gnd.n5660 240.244
R12908 gnd.n5660 gnd.n5659 240.244
R12909 gnd.n5659 gnd.n5650 240.244
R12910 gnd.n5654 gnd.n5650 240.244
R12911 gnd.n5654 gnd.n2730 240.244
R12912 gnd.n5718 gnd.n2730 240.244
R12913 gnd.n5718 gnd.n2727 240.244
R12914 gnd.n5725 gnd.n2727 240.244
R12915 gnd.n5725 gnd.n2728 240.244
R12916 gnd.n2728 gnd.n257 240.244
R12917 gnd.n6959 gnd.n257 240.244
R12918 gnd.n6959 gnd.n258 240.244
R12919 gnd.n6954 gnd.n258 240.244
R12920 gnd.n6954 gnd.n6953 240.244
R12921 gnd.n6953 gnd.n262 240.244
R12922 gnd.n278 gnd.n262 240.244
R12923 gnd.n279 gnd.n278 240.244
R12924 gnd.n279 gnd.n270 240.244
R12925 gnd.n6939 gnd.n270 240.244
R12926 gnd.n6939 gnd.n271 240.244
R12927 gnd.n6935 gnd.n271 240.244
R12928 gnd.n6935 gnd.n6934 240.244
R12929 gnd.n6934 gnd.n6912 240.244
R12930 gnd.n6912 gnd.n287 240.244
R12931 gnd.n6908 gnd.n287 240.244
R12932 gnd.n6908 gnd.n6907 240.244
R12933 gnd.n6907 gnd.n6906 240.244
R12934 gnd.n6906 gnd.n293 240.244
R12935 gnd.n6902 gnd.n293 240.244
R12936 gnd.n6227 gnd.n696 240.244
R12937 gnd.n6227 gnd.n699 240.244
R12938 gnd.n6223 gnd.n699 240.244
R12939 gnd.n6223 gnd.n701 240.244
R12940 gnd.n6219 gnd.n701 240.244
R12941 gnd.n6219 gnd.n707 240.244
R12942 gnd.n6215 gnd.n707 240.244
R12943 gnd.n6215 gnd.n709 240.244
R12944 gnd.n6211 gnd.n709 240.244
R12945 gnd.n6211 gnd.n715 240.244
R12946 gnd.n6207 gnd.n715 240.244
R12947 gnd.n6207 gnd.n717 240.244
R12948 gnd.n6203 gnd.n717 240.244
R12949 gnd.n6203 gnd.n723 240.244
R12950 gnd.n6199 gnd.n723 240.244
R12951 gnd.n6199 gnd.n725 240.244
R12952 gnd.n6195 gnd.n725 240.244
R12953 gnd.n6195 gnd.n731 240.244
R12954 gnd.n6191 gnd.n731 240.244
R12955 gnd.n6191 gnd.n733 240.244
R12956 gnd.n6187 gnd.n733 240.244
R12957 gnd.n6187 gnd.n739 240.244
R12958 gnd.n6183 gnd.n739 240.244
R12959 gnd.n6183 gnd.n741 240.244
R12960 gnd.n6179 gnd.n741 240.244
R12961 gnd.n6179 gnd.n747 240.244
R12962 gnd.n6175 gnd.n747 240.244
R12963 gnd.n6175 gnd.n749 240.244
R12964 gnd.n6171 gnd.n749 240.244
R12965 gnd.n6171 gnd.n755 240.244
R12966 gnd.n6167 gnd.n755 240.244
R12967 gnd.n6167 gnd.n757 240.244
R12968 gnd.n6163 gnd.n757 240.244
R12969 gnd.n6163 gnd.n763 240.244
R12970 gnd.n6159 gnd.n763 240.244
R12971 gnd.n6159 gnd.n765 240.244
R12972 gnd.n6155 gnd.n765 240.244
R12973 gnd.n6155 gnd.n771 240.244
R12974 gnd.n6151 gnd.n771 240.244
R12975 gnd.n6151 gnd.n773 240.244
R12976 gnd.n6147 gnd.n773 240.244
R12977 gnd.n6147 gnd.n779 240.244
R12978 gnd.n6143 gnd.n779 240.244
R12979 gnd.n6143 gnd.n781 240.244
R12980 gnd.n6139 gnd.n781 240.244
R12981 gnd.n6139 gnd.n787 240.244
R12982 gnd.n6135 gnd.n787 240.244
R12983 gnd.n6135 gnd.n789 240.244
R12984 gnd.n6131 gnd.n789 240.244
R12985 gnd.n6131 gnd.n795 240.244
R12986 gnd.n6127 gnd.n795 240.244
R12987 gnd.n6127 gnd.n797 240.244
R12988 gnd.n6123 gnd.n797 240.244
R12989 gnd.n6123 gnd.n803 240.244
R12990 gnd.n6119 gnd.n803 240.244
R12991 gnd.n6119 gnd.n805 240.244
R12992 gnd.n6115 gnd.n805 240.244
R12993 gnd.n6115 gnd.n811 240.244
R12994 gnd.n6111 gnd.n811 240.244
R12995 gnd.n6111 gnd.n813 240.244
R12996 gnd.n6107 gnd.n813 240.244
R12997 gnd.n6107 gnd.n819 240.244
R12998 gnd.n6103 gnd.n819 240.244
R12999 gnd.n6103 gnd.n821 240.244
R13000 gnd.n6099 gnd.n821 240.244
R13001 gnd.n6099 gnd.n827 240.244
R13002 gnd.n6095 gnd.n827 240.244
R13003 gnd.n6095 gnd.n829 240.244
R13004 gnd.n6091 gnd.n829 240.244
R13005 gnd.n6091 gnd.n835 240.244
R13006 gnd.n6087 gnd.n835 240.244
R13007 gnd.n6087 gnd.n837 240.244
R13008 gnd.n6083 gnd.n837 240.244
R13009 gnd.n6083 gnd.n843 240.244
R13010 gnd.n6079 gnd.n843 240.244
R13011 gnd.n6079 gnd.n845 240.244
R13012 gnd.n6075 gnd.n845 240.244
R13013 gnd.n6075 gnd.n851 240.244
R13014 gnd.n6071 gnd.n851 240.244
R13015 gnd.n6071 gnd.n853 240.244
R13016 gnd.n6067 gnd.n853 240.244
R13017 gnd.n6067 gnd.n859 240.244
R13018 gnd.n6063 gnd.n859 240.244
R13019 gnd.n6063 gnd.n861 240.244
R13020 gnd.n2544 gnd.n2543 240.244
R13021 gnd.n2545 gnd.n2544 240.244
R13022 gnd.n4487 gnd.n2545 240.244
R13023 gnd.n4487 gnd.n2548 240.244
R13024 gnd.n2549 gnd.n2548 240.244
R13025 gnd.n2550 gnd.n2549 240.244
R13026 gnd.n3520 gnd.n2550 240.244
R13027 gnd.n3520 gnd.n2553 240.244
R13028 gnd.n2554 gnd.n2553 240.244
R13029 gnd.n2555 gnd.n2554 240.244
R13030 gnd.n4707 gnd.n2555 240.244
R13031 gnd.n4707 gnd.n2558 240.244
R13032 gnd.n2559 gnd.n2558 240.244
R13033 gnd.n2560 gnd.n2559 240.244
R13034 gnd.n4744 gnd.n2560 240.244
R13035 gnd.n4744 gnd.n2563 240.244
R13036 gnd.n2564 gnd.n2563 240.244
R13037 gnd.n2565 gnd.n2564 240.244
R13038 gnd.n3436 gnd.n2565 240.244
R13039 gnd.n3436 gnd.n2568 240.244
R13040 gnd.n2569 gnd.n2568 240.244
R13041 gnd.n2570 gnd.n2569 240.244
R13042 gnd.n3420 gnd.n2570 240.244
R13043 gnd.n3420 gnd.n2573 240.244
R13044 gnd.n2574 gnd.n2573 240.244
R13045 gnd.n2575 gnd.n2574 240.244
R13046 gnd.n4894 gnd.n2575 240.244
R13047 gnd.n4894 gnd.n2578 240.244
R13048 gnd.n2579 gnd.n2578 240.244
R13049 gnd.n2580 gnd.n2579 240.244
R13050 gnd.n3375 gnd.n2580 240.244
R13051 gnd.n3375 gnd.n2583 240.244
R13052 gnd.n2584 gnd.n2583 240.244
R13053 gnd.n2585 gnd.n2584 240.244
R13054 gnd.n3348 gnd.n2585 240.244
R13055 gnd.n3348 gnd.n2588 240.244
R13056 gnd.n2589 gnd.n2588 240.244
R13057 gnd.n2590 gnd.n2589 240.244
R13058 gnd.n3331 gnd.n2590 240.244
R13059 gnd.n3331 gnd.n2593 240.244
R13060 gnd.n2594 gnd.n2593 240.244
R13061 gnd.n2595 gnd.n2594 240.244
R13062 gnd.n4985 gnd.n2595 240.244
R13063 gnd.n4985 gnd.n2598 240.244
R13064 gnd.n2599 gnd.n2598 240.244
R13065 gnd.n2600 gnd.n2599 240.244
R13066 gnd.n3295 gnd.n2600 240.244
R13067 gnd.n3295 gnd.n2603 240.244
R13068 gnd.n2604 gnd.n2603 240.244
R13069 gnd.n2605 gnd.n2604 240.244
R13070 gnd.n3268 gnd.n2605 240.244
R13071 gnd.n3268 gnd.n2608 240.244
R13072 gnd.n2609 gnd.n2608 240.244
R13073 gnd.n2610 gnd.n2609 240.244
R13074 gnd.n3249 gnd.n2610 240.244
R13075 gnd.n3249 gnd.n2613 240.244
R13076 gnd.n2614 gnd.n2613 240.244
R13077 gnd.n2615 gnd.n2614 240.244
R13078 gnd.n5203 gnd.n2615 240.244
R13079 gnd.n5203 gnd.n2618 240.244
R13080 gnd.n2619 gnd.n2618 240.244
R13081 gnd.n2620 gnd.n2619 240.244
R13082 gnd.n3206 gnd.n2620 240.244
R13083 gnd.n3206 gnd.n2623 240.244
R13084 gnd.n2624 gnd.n2623 240.244
R13085 gnd.n2625 gnd.n2624 240.244
R13086 gnd.n5287 gnd.n2625 240.244
R13087 gnd.n5287 gnd.n2628 240.244
R13088 gnd.n2629 gnd.n2628 240.244
R13089 gnd.n2630 gnd.n2629 240.244
R13090 gnd.n3168 gnd.n2630 240.244
R13091 gnd.n3168 gnd.n2633 240.244
R13092 gnd.n2634 gnd.n2633 240.244
R13093 gnd.n2635 gnd.n2634 240.244
R13094 gnd.n5307 gnd.n2635 240.244
R13095 gnd.n5307 gnd.n2638 240.244
R13096 gnd.n2639 gnd.n2638 240.244
R13097 gnd.n2640 gnd.n2639 240.244
R13098 gnd.n5521 gnd.n2640 240.244
R13099 gnd.n5521 gnd.n2643 240.244
R13100 gnd.n2644 gnd.n2643 240.244
R13101 gnd.n5796 gnd.n2644 240.244
R13102 gnd.n3774 gnd.n3773 240.244
R13103 gnd.n3789 gnd.n3773 240.244
R13104 gnd.n3791 gnd.n3790 240.244
R13105 gnd.n3801 gnd.n3800 240.244
R13106 gnd.n3812 gnd.n3811 240.244
R13107 gnd.n3814 gnd.n3813 240.244
R13108 gnd.n3824 gnd.n3823 240.244
R13109 gnd.n3837 gnd.n3836 240.244
R13110 gnd.n3839 gnd.n3838 240.244
R13111 gnd.n3722 gnd.n3721 240.244
R13112 gnd.n3767 gnd.n3723 240.244
R13113 gnd.n3727 gnd.n3726 240.244
R13114 gnd.n3733 gnd.n3728 240.244
R13115 gnd.n3735 gnd.n3734 240.244
R13116 gnd.n3739 gnd.n3738 240.244
R13117 gnd.n3740 gnd.n3739 240.244
R13118 gnd.n4486 gnd.n3740 240.244
R13119 gnd.n4486 gnd.n3743 240.244
R13120 gnd.n3744 gnd.n3743 240.244
R13121 gnd.n4507 gnd.n3744 240.244
R13122 gnd.n4507 gnd.n3493 240.244
R13123 gnd.n4678 gnd.n3493 240.244
R13124 gnd.n4678 gnd.n3488 240.244
R13125 gnd.n4698 gnd.n3488 240.244
R13126 gnd.n4698 gnd.n3481 240.244
R13127 gnd.n4683 gnd.n3481 240.244
R13128 gnd.n4684 gnd.n4683 240.244
R13129 gnd.n4685 gnd.n4684 240.244
R13130 gnd.n4685 gnd.n3461 240.244
R13131 gnd.n3461 gnd.n3447 240.244
R13132 gnd.n4764 gnd.n3447 240.244
R13133 gnd.n4765 gnd.n4764 240.244
R13134 gnd.n4765 gnd.n3441 240.244
R13135 gnd.n4778 gnd.n3441 240.244
R13136 gnd.n4778 gnd.n3442 240.244
R13137 gnd.n4770 gnd.n3442 240.244
R13138 gnd.n4771 gnd.n4770 240.244
R13139 gnd.n4771 gnd.n3404 240.244
R13140 gnd.n4851 gnd.n3404 240.244
R13141 gnd.n4851 gnd.n3399 240.244
R13142 gnd.n4893 gnd.n3399 240.244
R13143 gnd.n4893 gnd.n3391 240.244
R13144 gnd.n4856 gnd.n3391 240.244
R13145 gnd.n4857 gnd.n4856 240.244
R13146 gnd.n4858 gnd.n4857 240.244
R13147 gnd.n4858 gnd.n3370 240.244
R13148 gnd.n3370 gnd.n3362 240.244
R13149 gnd.n4862 gnd.n3362 240.244
R13150 gnd.n4863 gnd.n4862 240.244
R13151 gnd.n4866 gnd.n4863 240.244
R13152 gnd.n4867 gnd.n4866 240.244
R13153 gnd.n4868 gnd.n4867 240.244
R13154 gnd.n4869 gnd.n4868 240.244
R13155 gnd.n4870 gnd.n4869 240.244
R13156 gnd.n4870 gnd.n3316 240.244
R13157 gnd.n5028 gnd.n3316 240.244
R13158 gnd.n5028 gnd.n3311 240.244
R13159 gnd.n5070 gnd.n3311 240.244
R13160 gnd.n5070 gnd.n3303 240.244
R13161 gnd.n5033 gnd.n3303 240.244
R13162 gnd.n5034 gnd.n5033 240.244
R13163 gnd.n5036 gnd.n5034 240.244
R13164 gnd.n5036 gnd.n3283 240.244
R13165 gnd.n3283 gnd.n3275 240.244
R13166 gnd.n5039 gnd.n3275 240.244
R13167 gnd.n5040 gnd.n5039 240.244
R13168 gnd.n5043 gnd.n5040 240.244
R13169 gnd.n5044 gnd.n5043 240.244
R13170 gnd.n5045 gnd.n5044 240.244
R13171 gnd.n5046 gnd.n5045 240.244
R13172 gnd.n5047 gnd.n5046 240.244
R13173 gnd.n5047 gnd.n3228 240.244
R13174 gnd.n5205 gnd.n3228 240.244
R13175 gnd.n5205 gnd.n3223 240.244
R13176 gnd.n5223 gnd.n3223 240.244
R13177 gnd.n5223 gnd.n3216 240.244
R13178 gnd.n5210 gnd.n3216 240.244
R13179 gnd.n5211 gnd.n5210 240.244
R13180 gnd.n5212 gnd.n5211 240.244
R13181 gnd.n5212 gnd.n3196 240.244
R13182 gnd.n3196 gnd.n3181 240.244
R13183 gnd.n5297 gnd.n3181 240.244
R13184 gnd.n5297 gnd.n3175 240.244
R13185 gnd.n5320 gnd.n3175 240.244
R13186 gnd.n5320 gnd.n3176 240.244
R13187 gnd.n5302 gnd.n3176 240.244
R13188 gnd.n5304 gnd.n5302 240.244
R13189 gnd.n5305 gnd.n5304 240.244
R13190 gnd.n5309 gnd.n5305 240.244
R13191 gnd.n5309 gnd.n2970 240.244
R13192 gnd.n5511 gnd.n2970 240.244
R13193 gnd.n5511 gnd.n2966 240.244
R13194 gnd.n5518 gnd.n2966 240.244
R13195 gnd.n5518 gnd.n2959 240.244
R13196 gnd.n5534 gnd.n2959 240.244
R13197 gnd.n5534 gnd.n2648 240.244
R13198 gnd.n2868 gnd.n2867 240.244
R13199 gnd.n2871 gnd.n2870 240.244
R13200 gnd.n2887 gnd.n2886 240.244
R13201 gnd.n2890 gnd.n2889 240.244
R13202 gnd.n2906 gnd.n2905 240.244
R13203 gnd.n2909 gnd.n2908 240.244
R13204 gnd.n2925 gnd.n2924 240.244
R13205 gnd.n2928 gnd.n2927 240.244
R13206 gnd.n2942 gnd.n2941 240.244
R13207 gnd.n2945 gnd.n2944 240.244
R13208 gnd.n2950 gnd.n2947 240.244
R13209 gnd.n2953 gnd.n2952 240.244
R13210 gnd.n5539 gnd.n2955 240.244
R13211 gnd.n5542 gnd.n5541 240.244
R13212 gnd.n3504 gnd.n3503 240.132
R13213 gnd.n5353 gnd.n5352 240.132
R13214 gnd.n6235 gnd.n6234 225.874
R13215 gnd.n6236 gnd.n6235 225.874
R13216 gnd.n6236 gnd.n689 225.874
R13217 gnd.n6244 gnd.n689 225.874
R13218 gnd.n6245 gnd.n6244 225.874
R13219 gnd.n6246 gnd.n6245 225.874
R13220 gnd.n6246 gnd.n683 225.874
R13221 gnd.n6254 gnd.n683 225.874
R13222 gnd.n6255 gnd.n6254 225.874
R13223 gnd.n6256 gnd.n6255 225.874
R13224 gnd.n6256 gnd.n677 225.874
R13225 gnd.n6264 gnd.n677 225.874
R13226 gnd.n6265 gnd.n6264 225.874
R13227 gnd.n6266 gnd.n6265 225.874
R13228 gnd.n6266 gnd.n671 225.874
R13229 gnd.n6274 gnd.n671 225.874
R13230 gnd.n6275 gnd.n6274 225.874
R13231 gnd.n6276 gnd.n6275 225.874
R13232 gnd.n6276 gnd.n665 225.874
R13233 gnd.n6284 gnd.n665 225.874
R13234 gnd.n6285 gnd.n6284 225.874
R13235 gnd.n6286 gnd.n6285 225.874
R13236 gnd.n6286 gnd.n659 225.874
R13237 gnd.n6294 gnd.n659 225.874
R13238 gnd.n6295 gnd.n6294 225.874
R13239 gnd.n6296 gnd.n6295 225.874
R13240 gnd.n6296 gnd.n653 225.874
R13241 gnd.n6304 gnd.n653 225.874
R13242 gnd.n6305 gnd.n6304 225.874
R13243 gnd.n6306 gnd.n6305 225.874
R13244 gnd.n6306 gnd.n647 225.874
R13245 gnd.n6314 gnd.n647 225.874
R13246 gnd.n6315 gnd.n6314 225.874
R13247 gnd.n6316 gnd.n6315 225.874
R13248 gnd.n6316 gnd.n641 225.874
R13249 gnd.n6324 gnd.n641 225.874
R13250 gnd.n6325 gnd.n6324 225.874
R13251 gnd.n6326 gnd.n6325 225.874
R13252 gnd.n6326 gnd.n635 225.874
R13253 gnd.n6334 gnd.n635 225.874
R13254 gnd.n6335 gnd.n6334 225.874
R13255 gnd.n6336 gnd.n6335 225.874
R13256 gnd.n6336 gnd.n629 225.874
R13257 gnd.n6344 gnd.n629 225.874
R13258 gnd.n6345 gnd.n6344 225.874
R13259 gnd.n6346 gnd.n6345 225.874
R13260 gnd.n6346 gnd.n623 225.874
R13261 gnd.n6354 gnd.n623 225.874
R13262 gnd.n6355 gnd.n6354 225.874
R13263 gnd.n6356 gnd.n6355 225.874
R13264 gnd.n6356 gnd.n617 225.874
R13265 gnd.n6364 gnd.n617 225.874
R13266 gnd.n6365 gnd.n6364 225.874
R13267 gnd.n6366 gnd.n6365 225.874
R13268 gnd.n6366 gnd.n611 225.874
R13269 gnd.n6374 gnd.n611 225.874
R13270 gnd.n6375 gnd.n6374 225.874
R13271 gnd.n6376 gnd.n6375 225.874
R13272 gnd.n6376 gnd.n605 225.874
R13273 gnd.n6384 gnd.n605 225.874
R13274 gnd.n6385 gnd.n6384 225.874
R13275 gnd.n6386 gnd.n6385 225.874
R13276 gnd.n6386 gnd.n599 225.874
R13277 gnd.n6394 gnd.n599 225.874
R13278 gnd.n6395 gnd.n6394 225.874
R13279 gnd.n6396 gnd.n6395 225.874
R13280 gnd.n6396 gnd.n593 225.874
R13281 gnd.n6404 gnd.n593 225.874
R13282 gnd.n6405 gnd.n6404 225.874
R13283 gnd.n6406 gnd.n6405 225.874
R13284 gnd.n6406 gnd.n587 225.874
R13285 gnd.n6414 gnd.n587 225.874
R13286 gnd.n6415 gnd.n6414 225.874
R13287 gnd.n6416 gnd.n6415 225.874
R13288 gnd.n6416 gnd.n581 225.874
R13289 gnd.n6424 gnd.n581 225.874
R13290 gnd.n6425 gnd.n6424 225.874
R13291 gnd.n6426 gnd.n6425 225.874
R13292 gnd.n6426 gnd.n575 225.874
R13293 gnd.n6434 gnd.n575 225.874
R13294 gnd.n6435 gnd.n6434 225.874
R13295 gnd.n6436 gnd.n6435 225.874
R13296 gnd.n6436 gnd.n569 225.874
R13297 gnd.n6444 gnd.n569 225.874
R13298 gnd.n6445 gnd.n6444 225.874
R13299 gnd.n6446 gnd.n6445 225.874
R13300 gnd.n6446 gnd.n563 225.874
R13301 gnd.n6454 gnd.n563 225.874
R13302 gnd.n6455 gnd.n6454 225.874
R13303 gnd.n6456 gnd.n6455 225.874
R13304 gnd.n6456 gnd.n557 225.874
R13305 gnd.n6464 gnd.n557 225.874
R13306 gnd.n6465 gnd.n6464 225.874
R13307 gnd.n6466 gnd.n6465 225.874
R13308 gnd.n6466 gnd.n551 225.874
R13309 gnd.n6474 gnd.n551 225.874
R13310 gnd.n6475 gnd.n6474 225.874
R13311 gnd.n6476 gnd.n6475 225.874
R13312 gnd.n6476 gnd.n545 225.874
R13313 gnd.n6484 gnd.n545 225.874
R13314 gnd.n6485 gnd.n6484 225.874
R13315 gnd.n6486 gnd.n6485 225.874
R13316 gnd.n6486 gnd.n539 225.874
R13317 gnd.n6494 gnd.n539 225.874
R13318 gnd.n6495 gnd.n6494 225.874
R13319 gnd.n6496 gnd.n6495 225.874
R13320 gnd.n6496 gnd.n533 225.874
R13321 gnd.n6504 gnd.n533 225.874
R13322 gnd.n6505 gnd.n6504 225.874
R13323 gnd.n6506 gnd.n6505 225.874
R13324 gnd.n6506 gnd.n527 225.874
R13325 gnd.n6514 gnd.n527 225.874
R13326 gnd.n6515 gnd.n6514 225.874
R13327 gnd.n6516 gnd.n6515 225.874
R13328 gnd.n6516 gnd.n521 225.874
R13329 gnd.n6524 gnd.n521 225.874
R13330 gnd.n6525 gnd.n6524 225.874
R13331 gnd.n6526 gnd.n6525 225.874
R13332 gnd.n6526 gnd.n515 225.874
R13333 gnd.n6534 gnd.n515 225.874
R13334 gnd.n6535 gnd.n6534 225.874
R13335 gnd.n6536 gnd.n6535 225.874
R13336 gnd.n6536 gnd.n509 225.874
R13337 gnd.n6544 gnd.n509 225.874
R13338 gnd.n6545 gnd.n6544 225.874
R13339 gnd.n6546 gnd.n6545 225.874
R13340 gnd.n6546 gnd.n503 225.874
R13341 gnd.n6554 gnd.n503 225.874
R13342 gnd.n6555 gnd.n6554 225.874
R13343 gnd.n6556 gnd.n6555 225.874
R13344 gnd.n6556 gnd.n497 225.874
R13345 gnd.n6564 gnd.n497 225.874
R13346 gnd.n6565 gnd.n6564 225.874
R13347 gnd.n6566 gnd.n6565 225.874
R13348 gnd.n6566 gnd.n491 225.874
R13349 gnd.n6574 gnd.n491 225.874
R13350 gnd.n6575 gnd.n6574 225.874
R13351 gnd.n6576 gnd.n6575 225.874
R13352 gnd.n6576 gnd.n485 225.874
R13353 gnd.n6584 gnd.n485 225.874
R13354 gnd.n6585 gnd.n6584 225.874
R13355 gnd.n6586 gnd.n6585 225.874
R13356 gnd.n6586 gnd.n479 225.874
R13357 gnd.n6594 gnd.n479 225.874
R13358 gnd.n6595 gnd.n6594 225.874
R13359 gnd.n6596 gnd.n6595 225.874
R13360 gnd.n6596 gnd.n473 225.874
R13361 gnd.n6604 gnd.n473 225.874
R13362 gnd.n6605 gnd.n6604 225.874
R13363 gnd.n6606 gnd.n6605 225.874
R13364 gnd.n6606 gnd.n467 225.874
R13365 gnd.n6614 gnd.n467 225.874
R13366 gnd.n6615 gnd.n6614 225.874
R13367 gnd.n6616 gnd.n6615 225.874
R13368 gnd.n6616 gnd.n461 225.874
R13369 gnd.n6624 gnd.n461 225.874
R13370 gnd.n6625 gnd.n6624 225.874
R13371 gnd.n6626 gnd.n6625 225.874
R13372 gnd.n6626 gnd.n455 225.874
R13373 gnd.n6634 gnd.n455 225.874
R13374 gnd.n6635 gnd.n6634 225.874
R13375 gnd.n6636 gnd.n6635 225.874
R13376 gnd.n6636 gnd.n449 225.874
R13377 gnd.n6644 gnd.n449 225.874
R13378 gnd.n6645 gnd.n6644 225.874
R13379 gnd.n6646 gnd.n6645 225.874
R13380 gnd.n6646 gnd.n443 225.874
R13381 gnd.n6654 gnd.n443 225.874
R13382 gnd.n6655 gnd.n6654 225.874
R13383 gnd.n6656 gnd.n6655 225.874
R13384 gnd.n6656 gnd.n437 225.874
R13385 gnd.n6664 gnd.n437 225.874
R13386 gnd.n6665 gnd.n6664 225.874
R13387 gnd.n6666 gnd.n6665 225.874
R13388 gnd.n6666 gnd.n431 225.874
R13389 gnd.n6674 gnd.n431 225.874
R13390 gnd.n6675 gnd.n6674 225.874
R13391 gnd.n6676 gnd.n6675 225.874
R13392 gnd.n6676 gnd.n425 225.874
R13393 gnd.n6685 gnd.n425 225.874
R13394 gnd.n6686 gnd.n6685 225.874
R13395 gnd.n1408 gnd.t153 224.174
R13396 gnd.n932 gnd.t81 224.174
R13397 gnd.n3016 gnd.n3013 199.319
R13398 gnd.n3144 gnd.n3013 199.319
R13399 gnd.n3627 gnd.n3621 199.319
R13400 gnd.n3626 gnd.n3621 199.319
R13401 gnd.n3505 gnd.n3502 186.49
R13402 gnd.n5354 gnd.n5351 186.49
R13403 gnd.n2185 gnd.n2184 185
R13404 gnd.n2183 gnd.n2182 185
R13405 gnd.n2162 gnd.n2161 185
R13406 gnd.n2177 gnd.n2176 185
R13407 gnd.n2175 gnd.n2174 185
R13408 gnd.n2166 gnd.n2165 185
R13409 gnd.n2169 gnd.n2168 185
R13410 gnd.n2153 gnd.n2152 185
R13411 gnd.n2151 gnd.n2150 185
R13412 gnd.n2130 gnd.n2129 185
R13413 gnd.n2145 gnd.n2144 185
R13414 gnd.n2143 gnd.n2142 185
R13415 gnd.n2134 gnd.n2133 185
R13416 gnd.n2137 gnd.n2136 185
R13417 gnd.n2121 gnd.n2120 185
R13418 gnd.n2119 gnd.n2118 185
R13419 gnd.n2098 gnd.n2097 185
R13420 gnd.n2113 gnd.n2112 185
R13421 gnd.n2111 gnd.n2110 185
R13422 gnd.n2102 gnd.n2101 185
R13423 gnd.n2105 gnd.n2104 185
R13424 gnd.n2090 gnd.n2089 185
R13425 gnd.n2088 gnd.n2087 185
R13426 gnd.n2067 gnd.n2066 185
R13427 gnd.n2082 gnd.n2081 185
R13428 gnd.n2080 gnd.n2079 185
R13429 gnd.n2071 gnd.n2070 185
R13430 gnd.n2074 gnd.n2073 185
R13431 gnd.n2058 gnd.n2057 185
R13432 gnd.n2056 gnd.n2055 185
R13433 gnd.n2035 gnd.n2034 185
R13434 gnd.n2050 gnd.n2049 185
R13435 gnd.n2048 gnd.n2047 185
R13436 gnd.n2039 gnd.n2038 185
R13437 gnd.n2042 gnd.n2041 185
R13438 gnd.n2026 gnd.n2025 185
R13439 gnd.n2024 gnd.n2023 185
R13440 gnd.n2003 gnd.n2002 185
R13441 gnd.n2018 gnd.n2017 185
R13442 gnd.n2016 gnd.n2015 185
R13443 gnd.n2007 gnd.n2006 185
R13444 gnd.n2010 gnd.n2009 185
R13445 gnd.n1994 gnd.n1993 185
R13446 gnd.n1992 gnd.n1991 185
R13447 gnd.n1971 gnd.n1970 185
R13448 gnd.n1986 gnd.n1985 185
R13449 gnd.n1984 gnd.n1983 185
R13450 gnd.n1975 gnd.n1974 185
R13451 gnd.n1978 gnd.n1977 185
R13452 gnd.n1963 gnd.n1962 185
R13453 gnd.n1961 gnd.n1960 185
R13454 gnd.n1940 gnd.n1939 185
R13455 gnd.n1955 gnd.n1954 185
R13456 gnd.n1953 gnd.n1952 185
R13457 gnd.n1944 gnd.n1943 185
R13458 gnd.n1947 gnd.n1946 185
R13459 gnd.n1409 gnd.t152 178.987
R13460 gnd.n933 gnd.t82 178.987
R13461 gnd.n1 gnd.t182 170.774
R13462 gnd.n7 gnd.t207 170.103
R13463 gnd.n6 gnd.t171 170.103
R13464 gnd.n5 gnd.t156 170.103
R13465 gnd.n4 gnd.t243 170.103
R13466 gnd.n3 gnd.t271 170.103
R13467 gnd.n2 gnd.t200 170.103
R13468 gnd.n1 gnd.t202 170.103
R13469 gnd.n5425 gnd.n5424 163.367
R13470 gnd.n5421 gnd.n5420 163.367
R13471 gnd.n5417 gnd.n5416 163.367
R13472 gnd.n5413 gnd.n5412 163.367
R13473 gnd.n5409 gnd.n5408 163.367
R13474 gnd.n5405 gnd.n5404 163.367
R13475 gnd.n5401 gnd.n5400 163.367
R13476 gnd.n5397 gnd.n5396 163.367
R13477 gnd.n5393 gnd.n5392 163.367
R13478 gnd.n5389 gnd.n5388 163.367
R13479 gnd.n5385 gnd.n5384 163.367
R13480 gnd.n5381 gnd.n5380 163.367
R13481 gnd.n5377 gnd.n5376 163.367
R13482 gnd.n5373 gnd.n5372 163.367
R13483 gnd.n5368 gnd.n5367 163.367
R13484 gnd.n5364 gnd.n5363 163.367
R13485 gnd.n5498 gnd.n5497 163.367
R13486 gnd.n5494 gnd.n5493 163.367
R13487 gnd.n5489 gnd.n5488 163.367
R13488 gnd.n5485 gnd.n5484 163.367
R13489 gnd.n5481 gnd.n5480 163.367
R13490 gnd.n5477 gnd.n5476 163.367
R13491 gnd.n5473 gnd.n5472 163.367
R13492 gnd.n5469 gnd.n5468 163.367
R13493 gnd.n5465 gnd.n5464 163.367
R13494 gnd.n5461 gnd.n5460 163.367
R13495 gnd.n5457 gnd.n5456 163.367
R13496 gnd.n5453 gnd.n5452 163.367
R13497 gnd.n5449 gnd.n5448 163.367
R13498 gnd.n5445 gnd.n5444 163.367
R13499 gnd.n5441 gnd.n5440 163.367
R13500 gnd.n5437 gnd.n5436 163.367
R13501 gnd.n4662 gnd.n3495 163.367
R13502 gnd.n4662 gnd.n3487 163.367
R13503 gnd.n4657 gnd.n3487 163.367
R13504 gnd.n4657 gnd.n3482 163.367
R13505 gnd.n4654 gnd.n3482 163.367
R13506 gnd.n4654 gnd.n3472 163.367
R13507 gnd.n3472 gnd.n3464 163.367
R13508 gnd.n4726 gnd.n3464 163.367
R13509 gnd.n4726 gnd.n3462 163.367
R13510 gnd.n4741 gnd.n3462 163.367
R13511 gnd.n4741 gnd.n3453 163.367
R13512 gnd.n4737 gnd.n3453 163.367
R13513 gnd.n4737 gnd.n3448 163.367
R13514 gnd.n4734 gnd.n3448 163.367
R13515 gnd.n4734 gnd.n3435 163.367
R13516 gnd.n4730 gnd.n3435 163.367
R13517 gnd.n4730 gnd.n3428 163.367
R13518 gnd.n4797 gnd.n3428 163.367
R13519 gnd.n4797 gnd.n3426 163.367
R13520 gnd.n4822 gnd.n3426 163.367
R13521 gnd.n4822 gnd.n3419 163.367
R13522 gnd.n4818 gnd.n3419 163.367
R13523 gnd.n4818 gnd.n3410 163.367
R13524 gnd.n4813 gnd.n3410 163.367
R13525 gnd.n4813 gnd.n3405 163.367
R13526 gnd.n4810 gnd.n3405 163.367
R13527 gnd.n4810 gnd.n3398 163.367
R13528 gnd.n4805 gnd.n3398 163.367
R13529 gnd.n4805 gnd.n3392 163.367
R13530 gnd.n4802 gnd.n3392 163.367
R13531 gnd.n4802 gnd.n3382 163.367
R13532 gnd.n3382 gnd.n3373 163.367
R13533 gnd.n4921 gnd.n3373 163.367
R13534 gnd.n4921 gnd.n3371 163.367
R13535 gnd.n4928 gnd.n3371 163.367
R13536 gnd.n4928 gnd.n3361 163.367
R13537 gnd.n4924 gnd.n3361 163.367
R13538 gnd.n4924 gnd.n3356 163.367
R13539 gnd.n4950 gnd.n3356 163.367
R13540 gnd.n4950 gnd.n3350 163.367
R13541 gnd.n4954 gnd.n3350 163.367
R13542 gnd.n4954 gnd.n3341 163.367
R13543 gnd.n4974 gnd.n3341 163.367
R13544 gnd.n4974 gnd.n3339 163.367
R13545 gnd.n4999 gnd.n3339 163.367
R13546 gnd.n4999 gnd.n3333 163.367
R13547 gnd.n4995 gnd.n3333 163.367
R13548 gnd.n4995 gnd.n3324 163.367
R13549 gnd.n4991 gnd.n3324 163.367
R13550 gnd.n4991 gnd.n3318 163.367
R13551 gnd.n4988 gnd.n3318 163.367
R13552 gnd.n4988 gnd.n3310 163.367
R13553 gnd.n4982 gnd.n3310 163.367
R13554 gnd.n4982 gnd.n3304 163.367
R13555 gnd.n4979 gnd.n3304 163.367
R13556 gnd.n4979 gnd.n3293 163.367
R13557 gnd.n3293 gnd.n3286 163.367
R13558 gnd.n5097 gnd.n3286 163.367
R13559 gnd.n5097 gnd.n3284 163.367
R13560 gnd.n5104 gnd.n3284 163.367
R13561 gnd.n5104 gnd.n3274 163.367
R13562 gnd.n5100 gnd.n3274 163.367
R13563 gnd.n5100 gnd.n3267 163.367
R13564 gnd.n5126 gnd.n3267 163.367
R13565 gnd.n5126 gnd.n3261 163.367
R13566 gnd.n5130 gnd.n3261 163.367
R13567 gnd.n5130 gnd.n3253 163.367
R13568 gnd.n5150 gnd.n3253 163.367
R13569 gnd.n5150 gnd.n3251 163.367
R13570 gnd.n5175 gnd.n3251 163.367
R13571 gnd.n5175 gnd.n3244 163.367
R13572 gnd.n5171 gnd.n3244 163.367
R13573 gnd.n5171 gnd.n3236 163.367
R13574 gnd.n5167 gnd.n3236 163.367
R13575 gnd.n5167 gnd.n3230 163.367
R13576 gnd.n5164 gnd.n3230 163.367
R13577 gnd.n5164 gnd.n3222 163.367
R13578 gnd.n5158 gnd.n3222 163.367
R13579 gnd.n5158 gnd.n3217 163.367
R13580 gnd.n5155 gnd.n3217 163.367
R13581 gnd.n5155 gnd.n3207 163.367
R13582 gnd.n3207 gnd.n3199 163.367
R13583 gnd.n5250 gnd.n3199 163.367
R13584 gnd.n5250 gnd.n3197 163.367
R13585 gnd.n5273 gnd.n3197 163.367
R13586 gnd.n5273 gnd.n3188 163.367
R13587 gnd.n5269 gnd.n3188 163.367
R13588 gnd.n5269 gnd.n3183 163.367
R13589 gnd.n5266 gnd.n3183 163.367
R13590 gnd.n5266 gnd.n3174 163.367
R13591 gnd.n5260 gnd.n3174 163.367
R13592 gnd.n5260 gnd.n3167 163.367
R13593 gnd.n5257 gnd.n3167 163.367
R13594 gnd.n5257 gnd.n3159 163.367
R13595 gnd.n3159 gnd.n3152 163.367
R13596 gnd.n5432 gnd.n3152 163.367
R13597 gnd.n4670 gnd.n3519 163.367
R13598 gnd.n3559 gnd.n3519 163.367
R13599 gnd.n3563 gnd.n3562 163.367
R13600 gnd.n3567 gnd.n3566 163.367
R13601 gnd.n3571 gnd.n3570 163.367
R13602 gnd.n3575 gnd.n3574 163.367
R13603 gnd.n3579 gnd.n3578 163.367
R13604 gnd.n3583 gnd.n3582 163.367
R13605 gnd.n3587 gnd.n3586 163.367
R13606 gnd.n3591 gnd.n3590 163.367
R13607 gnd.n3595 gnd.n3594 163.367
R13608 gnd.n3599 gnd.n3598 163.367
R13609 gnd.n3603 gnd.n3602 163.367
R13610 gnd.n3607 gnd.n3606 163.367
R13611 gnd.n3611 gnd.n3610 163.367
R13612 gnd.n3615 gnd.n3614 163.367
R13613 gnd.n4590 gnd.n4589 163.367
R13614 gnd.n4594 gnd.n4593 163.367
R13615 gnd.n4599 gnd.n4598 163.367
R13616 gnd.n4603 gnd.n4602 163.367
R13617 gnd.n4607 gnd.n4606 163.367
R13618 gnd.n4611 gnd.n4610 163.367
R13619 gnd.n4615 gnd.n4614 163.367
R13620 gnd.n4619 gnd.n4618 163.367
R13621 gnd.n4623 gnd.n4622 163.367
R13622 gnd.n4627 gnd.n4626 163.367
R13623 gnd.n4631 gnd.n4630 163.367
R13624 gnd.n4635 gnd.n4634 163.367
R13625 gnd.n4639 gnd.n4638 163.367
R13626 gnd.n4643 gnd.n4642 163.367
R13627 gnd.n4647 gnd.n4646 163.367
R13628 gnd.n4649 gnd.n3553 163.367
R13629 gnd.n4675 gnd.n3485 163.367
R13630 gnd.n4701 gnd.n3485 163.367
R13631 gnd.n4701 gnd.n3483 163.367
R13632 gnd.n4705 gnd.n3483 163.367
R13633 gnd.n4705 gnd.n3470 163.367
R13634 gnd.n4719 gnd.n3470 163.367
R13635 gnd.n4719 gnd.n3467 163.367
R13636 gnd.n4724 gnd.n3467 163.367
R13637 gnd.n4724 gnd.n3468 163.367
R13638 gnd.n3468 gnd.n3452 163.367
R13639 gnd.n4757 gnd.n3452 163.367
R13640 gnd.n4757 gnd.n3450 163.367
R13641 gnd.n4761 gnd.n3450 163.367
R13642 gnd.n4761 gnd.n3437 163.367
R13643 gnd.n4785 gnd.n3437 163.367
R13644 gnd.n4785 gnd.n3438 163.367
R13645 gnd.n4781 gnd.n3438 163.367
R13646 gnd.n4781 gnd.n3424 163.367
R13647 gnd.n4826 gnd.n3424 163.367
R13648 gnd.n4826 gnd.n3422 163.367
R13649 gnd.n4830 gnd.n3422 163.367
R13650 gnd.n4830 gnd.n3409 163.367
R13651 gnd.n4844 gnd.n3409 163.367
R13652 gnd.n4844 gnd.n3407 163.367
R13653 gnd.n4848 gnd.n3407 163.367
R13654 gnd.n4848 gnd.n3396 163.367
R13655 gnd.n4897 gnd.n3396 163.367
R13656 gnd.n4897 gnd.n3394 163.367
R13657 gnd.n4901 gnd.n3394 163.367
R13658 gnd.n4901 gnd.n3380 163.367
R13659 gnd.n4914 gnd.n3380 163.367
R13660 gnd.n4914 gnd.n3377 163.367
R13661 gnd.n4919 gnd.n3377 163.367
R13662 gnd.n4919 gnd.n3378 163.367
R13663 gnd.n3378 gnd.n3359 163.367
R13664 gnd.n4942 gnd.n3359 163.367
R13665 gnd.n4942 gnd.n3357 163.367
R13666 gnd.n4946 gnd.n3357 163.367
R13667 gnd.n4946 gnd.n3352 163.367
R13668 gnd.n4962 gnd.n3352 163.367
R13669 gnd.n4962 gnd.n3353 163.367
R13670 gnd.n4958 gnd.n3353 163.367
R13671 gnd.n4958 gnd.n3337 163.367
R13672 gnd.n5003 gnd.n3337 163.367
R13673 gnd.n5003 gnd.n3335 163.367
R13674 gnd.n5007 gnd.n3335 163.367
R13675 gnd.n5007 gnd.n3322 163.367
R13676 gnd.n5021 gnd.n3322 163.367
R13677 gnd.n5021 gnd.n3320 163.367
R13678 gnd.n5025 gnd.n3320 163.367
R13679 gnd.n5025 gnd.n3308 163.367
R13680 gnd.n5073 gnd.n3308 163.367
R13681 gnd.n5073 gnd.n3306 163.367
R13682 gnd.n5077 gnd.n3306 163.367
R13683 gnd.n5077 gnd.n3291 163.367
R13684 gnd.n5090 gnd.n3291 163.367
R13685 gnd.n5090 gnd.n3288 163.367
R13686 gnd.n5095 gnd.n3288 163.367
R13687 gnd.n5095 gnd.n3289 163.367
R13688 gnd.n3289 gnd.n3272 163.367
R13689 gnd.n5118 gnd.n3272 163.367
R13690 gnd.n5118 gnd.n3270 163.367
R13691 gnd.n5122 gnd.n3270 163.367
R13692 gnd.n5122 gnd.n3263 163.367
R13693 gnd.n5138 gnd.n3263 163.367
R13694 gnd.n5138 gnd.n3264 163.367
R13695 gnd.n5134 gnd.n3264 163.367
R13696 gnd.n5134 gnd.n3248 163.367
R13697 gnd.n5179 gnd.n3248 163.367
R13698 gnd.n5179 gnd.n3246 163.367
R13699 gnd.n5183 gnd.n3246 163.367
R13700 gnd.n5183 gnd.n3234 163.367
R13701 gnd.n5197 gnd.n3234 163.367
R13702 gnd.n5197 gnd.n3232 163.367
R13703 gnd.n5201 gnd.n3232 163.367
R13704 gnd.n5201 gnd.n3221 163.367
R13705 gnd.n5226 gnd.n3221 163.367
R13706 gnd.n5226 gnd.n3219 163.367
R13707 gnd.n5230 gnd.n3219 163.367
R13708 gnd.n5230 gnd.n3205 163.367
R13709 gnd.n5243 gnd.n3205 163.367
R13710 gnd.n5243 gnd.n3202 163.367
R13711 gnd.n5248 gnd.n3202 163.367
R13712 gnd.n5248 gnd.n3203 163.367
R13713 gnd.n3203 gnd.n3186 163.367
R13714 gnd.n5290 gnd.n3186 163.367
R13715 gnd.n5290 gnd.n3184 163.367
R13716 gnd.n5294 gnd.n3184 163.367
R13717 gnd.n5294 gnd.n3172 163.367
R13718 gnd.n5323 gnd.n3172 163.367
R13719 gnd.n5323 gnd.n3170 163.367
R13720 gnd.n5327 gnd.n3170 163.367
R13721 gnd.n5327 gnd.n3157 163.367
R13722 gnd.n5339 gnd.n3157 163.367
R13723 gnd.n5339 gnd.n3154 163.367
R13724 gnd.n5430 gnd.n3154 163.367
R13725 gnd.n5360 gnd.n5359 156.462
R13726 gnd.n2125 gnd.n2093 153.042
R13727 gnd.n2189 gnd.n2188 152.079
R13728 gnd.n2157 gnd.n2156 152.079
R13729 gnd.n2125 gnd.n2124 152.079
R13730 gnd.n3510 gnd.n3509 152
R13731 gnd.n3511 gnd.n3500 152
R13732 gnd.n3513 gnd.n3512 152
R13733 gnd.n3515 gnd.n3498 152
R13734 gnd.n3517 gnd.n3516 152
R13735 gnd.n5358 gnd.n5342 152
R13736 gnd.n5350 gnd.n5343 152
R13737 gnd.n5349 gnd.n5348 152
R13738 gnd.n5347 gnd.n5344 152
R13739 gnd.n5345 gnd.t119 150.546
R13740 gnd.t223 gnd.n2167 147.661
R13741 gnd.t180 gnd.n2135 147.661
R13742 gnd.t178 gnd.n2103 147.661
R13743 gnd.t279 gnd.n2072 147.661
R13744 gnd.t194 gnd.n2040 147.661
R13745 gnd.t205 gnd.n2008 147.661
R13746 gnd.t283 gnd.n1976 147.661
R13747 gnd.t281 gnd.n1945 147.661
R13748 gnd.n3011 gnd.n2994 143.351
R13749 gnd.n4587 gnd.n3536 143.351
R13750 gnd.n4587 gnd.n3537 143.351
R13751 gnd.n3507 gnd.t83 130.484
R13752 gnd.n3516 gnd.t62 126.766
R13753 gnd.n3514 gnd.t125 126.766
R13754 gnd.n3500 gnd.t96 126.766
R13755 gnd.n3508 gnd.t144 126.766
R13756 gnd.n5346 gnd.t99 126.766
R13757 gnd.n5348 gnd.t122 126.766
R13758 gnd.n5357 gnd.t73 126.766
R13759 gnd.n5359 gnd.t135 126.766
R13760 gnd.n2184 gnd.n2183 104.615
R13761 gnd.n2183 gnd.n2161 104.615
R13762 gnd.n2176 gnd.n2161 104.615
R13763 gnd.n2176 gnd.n2175 104.615
R13764 gnd.n2175 gnd.n2165 104.615
R13765 gnd.n2168 gnd.n2165 104.615
R13766 gnd.n2152 gnd.n2151 104.615
R13767 gnd.n2151 gnd.n2129 104.615
R13768 gnd.n2144 gnd.n2129 104.615
R13769 gnd.n2144 gnd.n2143 104.615
R13770 gnd.n2143 gnd.n2133 104.615
R13771 gnd.n2136 gnd.n2133 104.615
R13772 gnd.n2120 gnd.n2119 104.615
R13773 gnd.n2119 gnd.n2097 104.615
R13774 gnd.n2112 gnd.n2097 104.615
R13775 gnd.n2112 gnd.n2111 104.615
R13776 gnd.n2111 gnd.n2101 104.615
R13777 gnd.n2104 gnd.n2101 104.615
R13778 gnd.n2089 gnd.n2088 104.615
R13779 gnd.n2088 gnd.n2066 104.615
R13780 gnd.n2081 gnd.n2066 104.615
R13781 gnd.n2081 gnd.n2080 104.615
R13782 gnd.n2080 gnd.n2070 104.615
R13783 gnd.n2073 gnd.n2070 104.615
R13784 gnd.n2057 gnd.n2056 104.615
R13785 gnd.n2056 gnd.n2034 104.615
R13786 gnd.n2049 gnd.n2034 104.615
R13787 gnd.n2049 gnd.n2048 104.615
R13788 gnd.n2048 gnd.n2038 104.615
R13789 gnd.n2041 gnd.n2038 104.615
R13790 gnd.n2025 gnd.n2024 104.615
R13791 gnd.n2024 gnd.n2002 104.615
R13792 gnd.n2017 gnd.n2002 104.615
R13793 gnd.n2017 gnd.n2016 104.615
R13794 gnd.n2016 gnd.n2006 104.615
R13795 gnd.n2009 gnd.n2006 104.615
R13796 gnd.n1993 gnd.n1992 104.615
R13797 gnd.n1992 gnd.n1970 104.615
R13798 gnd.n1985 gnd.n1970 104.615
R13799 gnd.n1985 gnd.n1984 104.615
R13800 gnd.n1984 gnd.n1974 104.615
R13801 gnd.n1977 gnd.n1974 104.615
R13802 gnd.n1962 gnd.n1961 104.615
R13803 gnd.n1961 gnd.n1939 104.615
R13804 gnd.n1954 gnd.n1939 104.615
R13805 gnd.n1954 gnd.n1953 104.615
R13806 gnd.n1953 gnd.n1943 104.615
R13807 gnd.n1946 gnd.n1943 104.615
R13808 gnd.n1334 gnd.t49 100.632
R13809 gnd.n906 gnd.t71 100.632
R13810 gnd.n7185 gnd.n93 99.6594
R13811 gnd.n7183 gnd.n7182 99.6594
R13812 gnd.n7178 gnd.n101 99.6594
R13813 gnd.n7176 gnd.n7175 99.6594
R13814 gnd.n7171 gnd.n108 99.6594
R13815 gnd.n7169 gnd.n7168 99.6594
R13816 gnd.n7164 gnd.n115 99.6594
R13817 gnd.n7162 gnd.n7161 99.6594
R13818 gnd.n7154 gnd.n122 99.6594
R13819 gnd.n7152 gnd.n7151 99.6594
R13820 gnd.n7147 gnd.n129 99.6594
R13821 gnd.n7145 gnd.n7144 99.6594
R13822 gnd.n7140 gnd.n136 99.6594
R13823 gnd.n7138 gnd.n7137 99.6594
R13824 gnd.n7133 gnd.n143 99.6594
R13825 gnd.n7131 gnd.n7130 99.6594
R13826 gnd.n7126 gnd.n150 99.6594
R13827 gnd.n7124 gnd.n7123 99.6594
R13828 gnd.n155 gnd.n154 99.6594
R13829 gnd.n3031 gnd.n2672 99.6594
R13830 gnd.n3039 gnd.n3038 99.6594
R13831 gnd.n3042 gnd.n3041 99.6594
R13832 gnd.n3049 gnd.n3048 99.6594
R13833 gnd.n3052 gnd.n3051 99.6594
R13834 gnd.n3060 gnd.n3059 99.6594
R13835 gnd.n3063 gnd.n3062 99.6594
R13836 gnd.n3017 gnd.n3016 99.6594
R13837 gnd.n3143 gnd.n3142 99.6594
R13838 gnd.n3136 gnd.n3073 99.6594
R13839 gnd.n3135 gnd.n3134 99.6594
R13840 gnd.n3128 gnd.n3079 99.6594
R13841 gnd.n3127 gnd.n3126 99.6594
R13842 gnd.n3120 gnd.n3085 99.6594
R13843 gnd.n3119 gnd.n3118 99.6594
R13844 gnd.n3112 gnd.n3091 99.6594
R13845 gnd.n3111 gnd.n3110 99.6594
R13846 gnd.n3102 gnd.n3097 99.6594
R13847 gnd.n3679 gnd.n3678 99.6594
R13848 gnd.n3674 gnd.n3633 99.6594
R13849 gnd.n3670 gnd.n3632 99.6594
R13850 gnd.n3666 gnd.n3631 99.6594
R13851 gnd.n3662 gnd.n3630 99.6594
R13852 gnd.n3658 gnd.n3629 99.6594
R13853 gnd.n3654 gnd.n3628 99.6594
R13854 gnd.n3626 gnd.n3625 99.6594
R13855 gnd.n4580 gnd.n4579 99.6594
R13856 gnd.n4577 gnd.n4576 99.6594
R13857 gnd.n4572 gnd.n3688 99.6594
R13858 gnd.n4570 gnd.n4569 99.6594
R13859 gnd.n4565 gnd.n3695 99.6594
R13860 gnd.n4563 gnd.n4562 99.6594
R13861 gnd.n4558 gnd.n3702 99.6594
R13862 gnd.n4556 gnd.n4555 99.6594
R13863 gnd.n4551 gnd.n3711 99.6594
R13864 gnd.n4549 gnd.n4548 99.6594
R13865 gnd.n4101 gnd.n2323 99.6594
R13866 gnd.n4109 gnd.n4108 99.6594
R13867 gnd.n4112 gnd.n4111 99.6594
R13868 gnd.n4119 gnd.n4118 99.6594
R13869 gnd.n4122 gnd.n4121 99.6594
R13870 gnd.n4129 gnd.n4128 99.6594
R13871 gnd.n4132 gnd.n4131 99.6594
R13872 gnd.n4139 gnd.n4138 99.6594
R13873 gnd.n4142 gnd.n4141 99.6594
R13874 gnd.n4149 gnd.n4148 99.6594
R13875 gnd.n4152 gnd.n4151 99.6594
R13876 gnd.n4159 gnd.n4158 99.6594
R13877 gnd.n4162 gnd.n4161 99.6594
R13878 gnd.n4169 gnd.n4168 99.6594
R13879 gnd.n4172 gnd.n4171 99.6594
R13880 gnd.n4179 gnd.n4178 99.6594
R13881 gnd.n4182 gnd.n4181 99.6594
R13882 gnd.n4190 gnd.n4189 99.6594
R13883 gnd.n4193 gnd.n4192 99.6594
R13884 gnd.n2307 gnd.n889 99.6594
R13885 gnd.n2305 gnd.n888 99.6594
R13886 gnd.n2301 gnd.n887 99.6594
R13887 gnd.n2297 gnd.n886 99.6594
R13888 gnd.n2293 gnd.n885 99.6594
R13889 gnd.n2289 gnd.n884 99.6594
R13890 gnd.n2285 gnd.n883 99.6594
R13891 gnd.n2217 gnd.n882 99.6594
R13892 gnd.n1546 gnd.n1277 99.6594
R13893 gnd.n1303 gnd.n1284 99.6594
R13894 gnd.n1305 gnd.n1285 99.6594
R13895 gnd.n1313 gnd.n1286 99.6594
R13896 gnd.n1315 gnd.n1287 99.6594
R13897 gnd.n1323 gnd.n1288 99.6594
R13898 gnd.n1325 gnd.n1289 99.6594
R13899 gnd.n1333 gnd.n1290 99.6594
R13900 gnd.n2275 gnd.n869 99.6594
R13901 gnd.n2271 gnd.n870 99.6594
R13902 gnd.n2267 gnd.n871 99.6594
R13903 gnd.n2263 gnd.n872 99.6594
R13904 gnd.n2259 gnd.n873 99.6594
R13905 gnd.n2255 gnd.n874 99.6594
R13906 gnd.n2251 gnd.n875 99.6594
R13907 gnd.n2247 gnd.n876 99.6594
R13908 gnd.n2243 gnd.n877 99.6594
R13909 gnd.n2239 gnd.n878 99.6594
R13910 gnd.n2235 gnd.n879 99.6594
R13911 gnd.n2231 gnd.n880 99.6594
R13912 gnd.n2227 gnd.n881 99.6594
R13913 gnd.n1461 gnd.n1460 99.6594
R13914 gnd.n1455 gnd.n1372 99.6594
R13915 gnd.n1452 gnd.n1373 99.6594
R13916 gnd.n1448 gnd.n1374 99.6594
R13917 gnd.n1444 gnd.n1375 99.6594
R13918 gnd.n1440 gnd.n1376 99.6594
R13919 gnd.n1436 gnd.n1377 99.6594
R13920 gnd.n1432 gnd.n1378 99.6594
R13921 gnd.n1428 gnd.n1379 99.6594
R13922 gnd.n1424 gnd.n1380 99.6594
R13923 gnd.n1420 gnd.n1381 99.6594
R13924 gnd.n1416 gnd.n1382 99.6594
R13925 gnd.n1463 gnd.n1371 99.6594
R13926 gnd.n7048 gnd.n7047 99.6594
R13927 gnd.n7053 gnd.n7052 99.6594
R13928 gnd.n7056 gnd.n7055 99.6594
R13929 gnd.n7061 gnd.n7060 99.6594
R13930 gnd.n7064 gnd.n7063 99.6594
R13931 gnd.n7069 gnd.n7068 99.6594
R13932 gnd.n7072 gnd.n7071 99.6594
R13933 gnd.n7077 gnd.n7076 99.6594
R13934 gnd.n7080 gnd.n80 99.6594
R13935 gnd.n2858 gnd.n2857 99.6594
R13936 gnd.n2861 gnd.n2860 99.6594
R13937 gnd.n2877 gnd.n2876 99.6594
R13938 gnd.n2880 gnd.n2879 99.6594
R13939 gnd.n2896 gnd.n2895 99.6594
R13940 gnd.n2899 gnd.n2898 99.6594
R13941 gnd.n2915 gnd.n2914 99.6594
R13942 gnd.n2918 gnd.n2917 99.6594
R13943 gnd.n2934 gnd.n2933 99.6594
R13944 gnd.n3783 gnd.n3782 99.6594
R13945 gnd.n3786 gnd.n3785 99.6594
R13946 gnd.n3796 gnd.n3795 99.6594
R13947 gnd.n3805 gnd.n3804 99.6594
R13948 gnd.n3808 gnd.n3807 99.6594
R13949 gnd.n3819 gnd.n3818 99.6594
R13950 gnd.n3828 gnd.n3827 99.6594
R13951 gnd.n3831 gnd.n3830 99.6594
R13952 gnd.n3842 gnd.n3841 99.6594
R13953 gnd.n4006 gnd.n4005 99.6594
R13954 gnd.n4009 gnd.n4008 99.6594
R13955 gnd.n4016 gnd.n4015 99.6594
R13956 gnd.n4019 gnd.n4018 99.6594
R13957 gnd.n4026 gnd.n4025 99.6594
R13958 gnd.n4029 gnd.n4028 99.6594
R13959 gnd.n4036 gnd.n4035 99.6594
R13960 gnd.n4039 gnd.n4038 99.6594
R13961 gnd.n4046 gnd.n4045 99.6594
R13962 gnd.n4007 gnd.n4006 99.6594
R13963 gnd.n4008 gnd.n3996 99.6594
R13964 gnd.n4017 gnd.n4016 99.6594
R13965 gnd.n4018 gnd.n3992 99.6594
R13966 gnd.n4027 gnd.n4026 99.6594
R13967 gnd.n4028 gnd.n3988 99.6594
R13968 gnd.n4037 gnd.n4036 99.6594
R13969 gnd.n4038 gnd.n3984 99.6594
R13970 gnd.n4047 gnd.n4046 99.6594
R13971 gnd.n3841 gnd.n3840 99.6594
R13972 gnd.n3830 gnd.n3829 99.6594
R13973 gnd.n3827 gnd.n3820 99.6594
R13974 gnd.n3818 gnd.n3817 99.6594
R13975 gnd.n3807 gnd.n3806 99.6594
R13976 gnd.n3804 gnd.n3797 99.6594
R13977 gnd.n3795 gnd.n3794 99.6594
R13978 gnd.n3785 gnd.n3784 99.6594
R13979 gnd.n3782 gnd.n3781 99.6594
R13980 gnd.n2859 gnd.n2858 99.6594
R13981 gnd.n2860 gnd.n2842 99.6594
R13982 gnd.n2878 gnd.n2877 99.6594
R13983 gnd.n2879 gnd.n2833 99.6594
R13984 gnd.n2897 gnd.n2896 99.6594
R13985 gnd.n2898 gnd.n2824 99.6594
R13986 gnd.n2916 gnd.n2915 99.6594
R13987 gnd.n2917 gnd.n2815 99.6594
R13988 gnd.n2935 gnd.n2934 99.6594
R13989 gnd.n7081 gnd.n7080 99.6594
R13990 gnd.n7076 gnd.n7075 99.6594
R13991 gnd.n7071 gnd.n7070 99.6594
R13992 gnd.n7068 gnd.n7067 99.6594
R13993 gnd.n7063 gnd.n7062 99.6594
R13994 gnd.n7060 gnd.n7059 99.6594
R13995 gnd.n7055 gnd.n7054 99.6594
R13996 gnd.n7052 gnd.n7051 99.6594
R13997 gnd.n7047 gnd.n7046 99.6594
R13998 gnd.n1461 gnd.n1384 99.6594
R13999 gnd.n1453 gnd.n1372 99.6594
R14000 gnd.n1449 gnd.n1373 99.6594
R14001 gnd.n1445 gnd.n1374 99.6594
R14002 gnd.n1441 gnd.n1375 99.6594
R14003 gnd.n1437 gnd.n1376 99.6594
R14004 gnd.n1433 gnd.n1377 99.6594
R14005 gnd.n1429 gnd.n1378 99.6594
R14006 gnd.n1425 gnd.n1379 99.6594
R14007 gnd.n1421 gnd.n1380 99.6594
R14008 gnd.n1417 gnd.n1381 99.6594
R14009 gnd.n1413 gnd.n1382 99.6594
R14010 gnd.n1464 gnd.n1463 99.6594
R14011 gnd.n2230 gnd.n881 99.6594
R14012 gnd.n2234 gnd.n880 99.6594
R14013 gnd.n2238 gnd.n879 99.6594
R14014 gnd.n2242 gnd.n878 99.6594
R14015 gnd.n2246 gnd.n877 99.6594
R14016 gnd.n2250 gnd.n876 99.6594
R14017 gnd.n2254 gnd.n875 99.6594
R14018 gnd.n2258 gnd.n874 99.6594
R14019 gnd.n2262 gnd.n873 99.6594
R14020 gnd.n2266 gnd.n872 99.6594
R14021 gnd.n2270 gnd.n871 99.6594
R14022 gnd.n2274 gnd.n870 99.6594
R14023 gnd.n910 gnd.n869 99.6594
R14024 gnd.n1547 gnd.n1546 99.6594
R14025 gnd.n1306 gnd.n1284 99.6594
R14026 gnd.n1312 gnd.n1285 99.6594
R14027 gnd.n1316 gnd.n1286 99.6594
R14028 gnd.n1322 gnd.n1287 99.6594
R14029 gnd.n1326 gnd.n1288 99.6594
R14030 gnd.n1332 gnd.n1289 99.6594
R14031 gnd.n1290 gnd.n1274 99.6594
R14032 gnd.n2284 gnd.n882 99.6594
R14033 gnd.n2288 gnd.n883 99.6594
R14034 gnd.n2292 gnd.n884 99.6594
R14035 gnd.n2296 gnd.n885 99.6594
R14036 gnd.n2300 gnd.n886 99.6594
R14037 gnd.n2304 gnd.n887 99.6594
R14038 gnd.n2308 gnd.n888 99.6594
R14039 gnd.n891 gnd.n889 99.6594
R14040 gnd.n4102 gnd.n4101 99.6594
R14041 gnd.n4110 gnd.n4109 99.6594
R14042 gnd.n4111 gnd.n4093 99.6594
R14043 gnd.n4120 gnd.n4119 99.6594
R14044 gnd.n4121 gnd.n4089 99.6594
R14045 gnd.n4130 gnd.n4129 99.6594
R14046 gnd.n4131 gnd.n4085 99.6594
R14047 gnd.n4140 gnd.n4139 99.6594
R14048 gnd.n4141 gnd.n4078 99.6594
R14049 gnd.n4150 gnd.n4149 99.6594
R14050 gnd.n4151 gnd.n4074 99.6594
R14051 gnd.n4160 gnd.n4159 99.6594
R14052 gnd.n4161 gnd.n4070 99.6594
R14053 gnd.n4170 gnd.n4169 99.6594
R14054 gnd.n4171 gnd.n4066 99.6594
R14055 gnd.n4180 gnd.n4179 99.6594
R14056 gnd.n4181 gnd.n4062 99.6594
R14057 gnd.n4191 gnd.n4190 99.6594
R14058 gnd.n4194 gnd.n4193 99.6594
R14059 gnd.n4550 gnd.n4549 99.6594
R14060 gnd.n3711 gnd.n3703 99.6594
R14061 gnd.n4557 gnd.n4556 99.6594
R14062 gnd.n3702 gnd.n3696 99.6594
R14063 gnd.n4564 gnd.n4563 99.6594
R14064 gnd.n3695 gnd.n3689 99.6594
R14065 gnd.n4571 gnd.n4570 99.6594
R14066 gnd.n3688 gnd.n3682 99.6594
R14067 gnd.n4578 gnd.n4577 99.6594
R14068 gnd.n4581 gnd.n4580 99.6594
R14069 gnd.n3653 gnd.n3627 99.6594
R14070 gnd.n3657 gnd.n3628 99.6594
R14071 gnd.n3661 gnd.n3629 99.6594
R14072 gnd.n3665 gnd.n3630 99.6594
R14073 gnd.n3669 gnd.n3631 99.6594
R14074 gnd.n3673 gnd.n3632 99.6594
R14075 gnd.n3635 gnd.n3633 99.6594
R14076 gnd.n3679 gnd.n3634 99.6594
R14077 gnd.n3032 gnd.n3031 99.6594
R14078 gnd.n3040 gnd.n3039 99.6594
R14079 gnd.n3041 gnd.n3023 99.6594
R14080 gnd.n3050 gnd.n3049 99.6594
R14081 gnd.n3051 gnd.n3019 99.6594
R14082 gnd.n3061 gnd.n3060 99.6594
R14083 gnd.n3064 gnd.n3063 99.6594
R14084 gnd.n3145 gnd.n3144 99.6594
R14085 gnd.n3142 gnd.n3141 99.6594
R14086 gnd.n3137 gnd.n3136 99.6594
R14087 gnd.n3134 gnd.n3133 99.6594
R14088 gnd.n3129 gnd.n3128 99.6594
R14089 gnd.n3126 gnd.n3125 99.6594
R14090 gnd.n3121 gnd.n3120 99.6594
R14091 gnd.n3118 gnd.n3117 99.6594
R14092 gnd.n3113 gnd.n3112 99.6594
R14093 gnd.n3110 gnd.n3109 99.6594
R14094 gnd.n3103 gnd.n3102 99.6594
R14095 gnd.n154 gnd.n151 99.6594
R14096 gnd.n7125 gnd.n7124 99.6594
R14097 gnd.n150 gnd.n144 99.6594
R14098 gnd.n7132 gnd.n7131 99.6594
R14099 gnd.n143 gnd.n137 99.6594
R14100 gnd.n7139 gnd.n7138 99.6594
R14101 gnd.n136 gnd.n130 99.6594
R14102 gnd.n7146 gnd.n7145 99.6594
R14103 gnd.n129 gnd.n123 99.6594
R14104 gnd.n7153 gnd.n7152 99.6594
R14105 gnd.n122 gnd.n116 99.6594
R14106 gnd.n7163 gnd.n7162 99.6594
R14107 gnd.n115 gnd.n109 99.6594
R14108 gnd.n7170 gnd.n7169 99.6594
R14109 gnd.n108 gnd.n102 99.6594
R14110 gnd.n7177 gnd.n7176 99.6594
R14111 gnd.n101 gnd.n95 99.6594
R14112 gnd.n7184 gnd.n7183 99.6594
R14113 gnd.n93 gnd.n90 99.6594
R14114 gnd.n3889 gnd.n3888 99.6594
R14115 gnd.n3789 gnd.n3758 99.6594
R14116 gnd.n3791 gnd.n3759 99.6594
R14117 gnd.n3801 gnd.n3760 99.6594
R14118 gnd.n3812 gnd.n3761 99.6594
R14119 gnd.n3814 gnd.n3762 99.6594
R14120 gnd.n3824 gnd.n3763 99.6594
R14121 gnd.n3837 gnd.n3764 99.6594
R14122 gnd.n3838 gnd.n3765 99.6594
R14123 gnd.n3766 gnd.n3722 99.6594
R14124 gnd.n3768 gnd.n3767 99.6594
R14125 gnd.n3769 gnd.n3727 99.6594
R14126 gnd.n3770 gnd.n3733 99.6594
R14127 gnd.n3772 gnd.n3735 99.6594
R14128 gnd.n3889 gnd.n3774 99.6594
R14129 gnd.n3790 gnd.n3758 99.6594
R14130 gnd.n3800 gnd.n3759 99.6594
R14131 gnd.n3811 gnd.n3760 99.6594
R14132 gnd.n3813 gnd.n3761 99.6594
R14133 gnd.n3823 gnd.n3762 99.6594
R14134 gnd.n3836 gnd.n3763 99.6594
R14135 gnd.n3839 gnd.n3764 99.6594
R14136 gnd.n3765 gnd.n3721 99.6594
R14137 gnd.n3766 gnd.n3723 99.6594
R14138 gnd.n3768 gnd.n3726 99.6594
R14139 gnd.n3769 gnd.n3728 99.6594
R14140 gnd.n3770 gnd.n3734 99.6594
R14141 gnd.n3772 gnd.n3771 99.6594
R14142 gnd.n2867 gnd.n2847 99.6594
R14143 gnd.n2871 gnd.n2869 99.6594
R14144 gnd.n2886 gnd.n2838 99.6594
R14145 gnd.n2890 gnd.n2888 99.6594
R14146 gnd.n2905 gnd.n2829 99.6594
R14147 gnd.n2909 gnd.n2907 99.6594
R14148 gnd.n2924 gnd.n2820 99.6594
R14149 gnd.n2928 gnd.n2926 99.6594
R14150 gnd.n2941 gnd.n2809 99.6594
R14151 gnd.n2944 gnd.n2943 99.6594
R14152 gnd.n2947 gnd.n2946 99.6594
R14153 gnd.n2952 gnd.n2951 99.6594
R14154 gnd.n2955 gnd.n2954 99.6594
R14155 gnd.n5541 gnd.n5540 99.6594
R14156 gnd.n5540 gnd.n5539 99.6594
R14157 gnd.n2954 gnd.n2953 99.6594
R14158 gnd.n2951 gnd.n2950 99.6594
R14159 gnd.n2946 gnd.n2945 99.6594
R14160 gnd.n2943 gnd.n2942 99.6594
R14161 gnd.n2927 gnd.n2809 99.6594
R14162 gnd.n2926 gnd.n2925 99.6594
R14163 gnd.n2908 gnd.n2820 99.6594
R14164 gnd.n2907 gnd.n2906 99.6594
R14165 gnd.n2889 gnd.n2829 99.6594
R14166 gnd.n2888 gnd.n2887 99.6594
R14167 gnd.n2870 gnd.n2838 99.6594
R14168 gnd.n2869 gnd.n2868 99.6594
R14169 gnd.n2847 gnd.n2646 99.6594
R14170 gnd.n3729 gnd.t118 98.63
R14171 gnd.n7078 gnd.t103 98.63
R14172 gnd.n2812 gnd.t91 98.63
R14173 gnd.n3832 gnd.t113 98.63
R14174 gnd.n3069 gnd.t88 98.63
R14175 gnd.n3098 gnd.t57 98.63
R14176 gnd.n157 gnd.t52 98.63
R14177 gnd.n7156 gnd.t77 98.63
R14178 gnd.n4082 gnd.t149 98.63
R14179 gnd.n4058 gnd.t140 98.63
R14180 gnd.n3981 gnd.t131 98.63
R14181 gnd.n3708 gnd.t67 98.63
R14182 gnd.n3619 gnd.t106 98.63
R14183 gnd.n5549 gnd.t94 98.63
R14184 gnd.n3554 gnd.t134 96.6984
R14185 gnd.n3149 gnd.t110 96.6984
R14186 gnd.n3556 gnd.t61 96.6906
R14187 gnd.n5361 gnd.t142 96.6906
R14188 gnd.n3507 gnd.n3506 81.8399
R14189 gnd.n3148 gnd.n3147 77.1205
R14190 gnd.n4588 gnd.n4586 77.1205
R14191 gnd.n1335 gnd.t48 74.8376
R14192 gnd.n907 gnd.t72 74.8376
R14193 gnd.n3555 gnd.t133 72.8438
R14194 gnd.n3150 gnd.t111 72.8438
R14195 gnd.n3508 gnd.n3501 72.8411
R14196 gnd.n3514 gnd.n3499 72.8411
R14197 gnd.n5357 gnd.n5356 72.8411
R14198 gnd.n3730 gnd.t117 72.836
R14199 gnd.n3557 gnd.t60 72.836
R14200 gnd.n5362 gnd.t143 72.836
R14201 gnd.n7079 gnd.t104 72.836
R14202 gnd.n2813 gnd.t90 72.836
R14203 gnd.n3833 gnd.t114 72.836
R14204 gnd.n3070 gnd.t87 72.836
R14205 gnd.n3099 gnd.t56 72.836
R14206 gnd.n158 gnd.t53 72.836
R14207 gnd.n7157 gnd.t78 72.836
R14208 gnd.n4083 gnd.t148 72.836
R14209 gnd.n4059 gnd.t139 72.836
R14210 gnd.n3982 gnd.t130 72.836
R14211 gnd.n3709 gnd.t68 72.836
R14212 gnd.n3620 gnd.t107 72.836
R14213 gnd.n5550 gnd.t95 72.836
R14214 gnd.n5425 gnd.n2978 71.676
R14215 gnd.n5421 gnd.n2979 71.676
R14216 gnd.n5417 gnd.n2980 71.676
R14217 gnd.n5413 gnd.n2981 71.676
R14218 gnd.n5409 gnd.n2982 71.676
R14219 gnd.n5405 gnd.n2983 71.676
R14220 gnd.n5401 gnd.n2984 71.676
R14221 gnd.n5397 gnd.n2985 71.676
R14222 gnd.n5393 gnd.n2986 71.676
R14223 gnd.n5389 gnd.n2987 71.676
R14224 gnd.n5385 gnd.n2988 71.676
R14225 gnd.n5381 gnd.n2989 71.676
R14226 gnd.n5377 gnd.n2990 71.676
R14227 gnd.n5373 gnd.n2991 71.676
R14228 gnd.n5368 gnd.n2992 71.676
R14229 gnd.n5364 gnd.n2993 71.676
R14230 gnd.n5498 gnd.n3011 71.676
R14231 gnd.n5494 gnd.n3010 71.676
R14232 gnd.n5489 gnd.n3009 71.676
R14233 gnd.n5485 gnd.n3008 71.676
R14234 gnd.n5481 gnd.n3007 71.676
R14235 gnd.n5477 gnd.n3006 71.676
R14236 gnd.n5473 gnd.n3005 71.676
R14237 gnd.n5469 gnd.n3004 71.676
R14238 gnd.n5465 gnd.n3003 71.676
R14239 gnd.n5461 gnd.n3002 71.676
R14240 gnd.n5457 gnd.n3001 71.676
R14241 gnd.n5453 gnd.n3000 71.676
R14242 gnd.n5449 gnd.n2999 71.676
R14243 gnd.n5445 gnd.n2998 71.676
R14244 gnd.n5441 gnd.n2997 71.676
R14245 gnd.n5437 gnd.n2996 71.676
R14246 gnd.n5433 gnd.n2995 71.676
R14247 gnd.n4669 gnd.n3497 71.676
R14248 gnd.n3559 gnd.n3522 71.676
R14249 gnd.n3563 gnd.n3523 71.676
R14250 gnd.n3567 gnd.n3524 71.676
R14251 gnd.n3571 gnd.n3525 71.676
R14252 gnd.n3575 gnd.n3526 71.676
R14253 gnd.n3579 gnd.n3527 71.676
R14254 gnd.n3583 gnd.n3528 71.676
R14255 gnd.n3587 gnd.n3529 71.676
R14256 gnd.n3591 gnd.n3530 71.676
R14257 gnd.n3595 gnd.n3531 71.676
R14258 gnd.n3599 gnd.n3532 71.676
R14259 gnd.n3603 gnd.n3533 71.676
R14260 gnd.n3607 gnd.n3534 71.676
R14261 gnd.n3611 gnd.n3535 71.676
R14262 gnd.n3615 gnd.n3536 71.676
R14263 gnd.n4590 gnd.n3538 71.676
R14264 gnd.n4594 gnd.n3539 71.676
R14265 gnd.n4599 gnd.n3540 71.676
R14266 gnd.n4603 gnd.n3541 71.676
R14267 gnd.n4607 gnd.n3542 71.676
R14268 gnd.n4611 gnd.n3543 71.676
R14269 gnd.n4615 gnd.n3544 71.676
R14270 gnd.n4619 gnd.n3545 71.676
R14271 gnd.n4623 gnd.n3546 71.676
R14272 gnd.n4627 gnd.n3547 71.676
R14273 gnd.n4631 gnd.n3548 71.676
R14274 gnd.n4635 gnd.n3549 71.676
R14275 gnd.n4639 gnd.n3550 71.676
R14276 gnd.n4643 gnd.n3551 71.676
R14277 gnd.n4647 gnd.n3552 71.676
R14278 gnd.n4667 gnd.n3553 71.676
R14279 gnd.n4670 gnd.n4669 71.676
R14280 gnd.n3562 gnd.n3522 71.676
R14281 gnd.n3566 gnd.n3523 71.676
R14282 gnd.n3570 gnd.n3524 71.676
R14283 gnd.n3574 gnd.n3525 71.676
R14284 gnd.n3578 gnd.n3526 71.676
R14285 gnd.n3582 gnd.n3527 71.676
R14286 gnd.n3586 gnd.n3528 71.676
R14287 gnd.n3590 gnd.n3529 71.676
R14288 gnd.n3594 gnd.n3530 71.676
R14289 gnd.n3598 gnd.n3531 71.676
R14290 gnd.n3602 gnd.n3532 71.676
R14291 gnd.n3606 gnd.n3533 71.676
R14292 gnd.n3610 gnd.n3534 71.676
R14293 gnd.n3614 gnd.n3535 71.676
R14294 gnd.n4589 gnd.n3537 71.676
R14295 gnd.n4593 gnd.n3538 71.676
R14296 gnd.n4598 gnd.n3539 71.676
R14297 gnd.n4602 gnd.n3540 71.676
R14298 gnd.n4606 gnd.n3541 71.676
R14299 gnd.n4610 gnd.n3542 71.676
R14300 gnd.n4614 gnd.n3543 71.676
R14301 gnd.n4618 gnd.n3544 71.676
R14302 gnd.n4622 gnd.n3545 71.676
R14303 gnd.n4626 gnd.n3546 71.676
R14304 gnd.n4630 gnd.n3547 71.676
R14305 gnd.n4634 gnd.n3548 71.676
R14306 gnd.n4638 gnd.n3549 71.676
R14307 gnd.n4642 gnd.n3550 71.676
R14308 gnd.n4646 gnd.n3551 71.676
R14309 gnd.n4649 gnd.n3552 71.676
R14310 gnd.n4667 gnd.n4666 71.676
R14311 gnd.n5436 gnd.n2995 71.676
R14312 gnd.n5440 gnd.n2996 71.676
R14313 gnd.n5444 gnd.n2997 71.676
R14314 gnd.n5448 gnd.n2998 71.676
R14315 gnd.n5452 gnd.n2999 71.676
R14316 gnd.n5456 gnd.n3000 71.676
R14317 gnd.n5460 gnd.n3001 71.676
R14318 gnd.n5464 gnd.n3002 71.676
R14319 gnd.n5468 gnd.n3003 71.676
R14320 gnd.n5472 gnd.n3004 71.676
R14321 gnd.n5476 gnd.n3005 71.676
R14322 gnd.n5480 gnd.n3006 71.676
R14323 gnd.n5484 gnd.n3007 71.676
R14324 gnd.n5488 gnd.n3008 71.676
R14325 gnd.n5493 gnd.n3009 71.676
R14326 gnd.n5497 gnd.n3010 71.676
R14327 gnd.n5363 gnd.n2994 71.676
R14328 gnd.n5367 gnd.n2993 71.676
R14329 gnd.n5372 gnd.n2992 71.676
R14330 gnd.n5376 gnd.n2991 71.676
R14331 gnd.n5380 gnd.n2990 71.676
R14332 gnd.n5384 gnd.n2989 71.676
R14333 gnd.n5388 gnd.n2988 71.676
R14334 gnd.n5392 gnd.n2987 71.676
R14335 gnd.n5396 gnd.n2986 71.676
R14336 gnd.n5400 gnd.n2985 71.676
R14337 gnd.n5404 gnd.n2984 71.676
R14338 gnd.n5408 gnd.n2983 71.676
R14339 gnd.n5412 gnd.n2982 71.676
R14340 gnd.n5416 gnd.n2981 71.676
R14341 gnd.n5420 gnd.n2980 71.676
R14342 gnd.n5424 gnd.n2979 71.676
R14343 gnd.n3155 gnd.n2978 71.676
R14344 gnd.n8 gnd.t277 69.1507
R14345 gnd.n14 gnd.t1 68.4792
R14346 gnd.n13 gnd.t226 68.4792
R14347 gnd.n12 gnd.t191 68.4792
R14348 gnd.n11 gnd.t228 68.4792
R14349 gnd.n10 gnd.t167 68.4792
R14350 gnd.n9 gnd.t15 68.4792
R14351 gnd.n8 gnd.t169 68.4792
R14352 gnd.n1462 gnd.n1366 64.369
R14353 gnd.n4596 gnd.n3555 59.5399
R14354 gnd.n5491 gnd.n3150 59.5399
R14355 gnd.n3558 gnd.n3557 59.5399
R14356 gnd.n5370 gnd.n5362 59.5399
R14357 gnd.n4673 gnd.n3517 59.1804
R14358 gnd.n2316 gnd.n867 57.3586
R14359 gnd.n1121 gnd.t186 56.607
R14360 gnd.n40 gnd.t253 56.607
R14361 gnd.n1098 gnd.t255 56.407
R14362 gnd.n1109 gnd.t160 56.407
R14363 gnd.n17 gnd.t162 56.407
R14364 gnd.n28 gnd.t214 56.407
R14365 gnd.n1130 gnd.t236 55.8337
R14366 gnd.n1107 gnd.t213 55.8337
R14367 gnd.n1118 gnd.t261 55.8337
R14368 gnd.n49 gnd.t11 55.8337
R14369 gnd.n26 gnd.t237 55.8337
R14370 gnd.n37 gnd.t163 55.8337
R14371 gnd.n3505 gnd.n3504 54.358
R14372 gnd.n5354 gnd.n5353 54.358
R14373 gnd.n1121 gnd.n1120 53.0052
R14374 gnd.n1123 gnd.n1122 53.0052
R14375 gnd.n1125 gnd.n1124 53.0052
R14376 gnd.n1127 gnd.n1126 53.0052
R14377 gnd.n1129 gnd.n1128 53.0052
R14378 gnd.n1098 gnd.n1097 53.0052
R14379 gnd.n1100 gnd.n1099 53.0052
R14380 gnd.n1102 gnd.n1101 53.0052
R14381 gnd.n1104 gnd.n1103 53.0052
R14382 gnd.n1106 gnd.n1105 53.0052
R14383 gnd.n1109 gnd.n1108 53.0052
R14384 gnd.n1111 gnd.n1110 53.0052
R14385 gnd.n1113 gnd.n1112 53.0052
R14386 gnd.n1115 gnd.n1114 53.0052
R14387 gnd.n1117 gnd.n1116 53.0052
R14388 gnd.n48 gnd.n47 53.0052
R14389 gnd.n46 gnd.n45 53.0052
R14390 gnd.n44 gnd.n43 53.0052
R14391 gnd.n42 gnd.n41 53.0052
R14392 gnd.n40 gnd.n39 53.0052
R14393 gnd.n25 gnd.n24 53.0052
R14394 gnd.n23 gnd.n22 53.0052
R14395 gnd.n21 gnd.n20 53.0052
R14396 gnd.n19 gnd.n18 53.0052
R14397 gnd.n17 gnd.n16 53.0052
R14398 gnd.n36 gnd.n35 53.0052
R14399 gnd.n34 gnd.n33 53.0052
R14400 gnd.n32 gnd.n31 53.0052
R14401 gnd.n30 gnd.n29 53.0052
R14402 gnd.n28 gnd.n27 53.0052
R14403 gnd.n5345 gnd.n5344 52.4801
R14404 gnd.n2168 gnd.t223 52.3082
R14405 gnd.n2136 gnd.t180 52.3082
R14406 gnd.n2104 gnd.t178 52.3082
R14407 gnd.n2073 gnd.t279 52.3082
R14408 gnd.n2041 gnd.t194 52.3082
R14409 gnd.n2009 gnd.t205 52.3082
R14410 gnd.n1977 gnd.t283 52.3082
R14411 gnd.n1946 gnd.t281 52.3082
R14412 gnd.n1998 gnd.n1966 51.4173
R14413 gnd.n2062 gnd.n2061 50.455
R14414 gnd.n2030 gnd.n2029 50.455
R14415 gnd.n1998 gnd.n1997 50.455
R14416 gnd.n1409 gnd.n1408 45.1884
R14417 gnd.n933 gnd.n932 45.1884
R14418 gnd.n5428 gnd.n5360 44.3322
R14419 gnd.n3508 gnd.n3507 44.3189
R14420 gnd.n6226 gnd.n695 43.8514
R14421 gnd.n6226 gnd.n6225 43.8514
R14422 gnd.n6225 gnd.n6224 43.8514
R14423 gnd.n6224 gnd.n700 43.8514
R14424 gnd.n6218 gnd.n700 43.8514
R14425 gnd.n6218 gnd.n6217 43.8514
R14426 gnd.n6217 gnd.n6216 43.8514
R14427 gnd.n6216 gnd.n708 43.8514
R14428 gnd.n6210 gnd.n708 43.8514
R14429 gnd.n6210 gnd.n6209 43.8514
R14430 gnd.n6209 gnd.n6208 43.8514
R14431 gnd.n6208 gnd.n716 43.8514
R14432 gnd.n6202 gnd.n716 43.8514
R14433 gnd.n6202 gnd.n6201 43.8514
R14434 gnd.n6201 gnd.n6200 43.8514
R14435 gnd.n6200 gnd.n724 43.8514
R14436 gnd.n6194 gnd.n724 43.8514
R14437 gnd.n6194 gnd.n6193 43.8514
R14438 gnd.n6193 gnd.n6192 43.8514
R14439 gnd.n6192 gnd.n732 43.8514
R14440 gnd.n6186 gnd.n732 43.8514
R14441 gnd.n6186 gnd.n6185 43.8514
R14442 gnd.n6185 gnd.n6184 43.8514
R14443 gnd.n6184 gnd.n740 43.8514
R14444 gnd.n6178 gnd.n740 43.8514
R14445 gnd.n6178 gnd.n6177 43.8514
R14446 gnd.n6177 gnd.n6176 43.8514
R14447 gnd.n6176 gnd.n748 43.8514
R14448 gnd.n6170 gnd.n748 43.8514
R14449 gnd.n6170 gnd.n6169 43.8514
R14450 gnd.n6169 gnd.n6168 43.8514
R14451 gnd.n6168 gnd.n756 43.8514
R14452 gnd.n6162 gnd.n756 43.8514
R14453 gnd.n6162 gnd.n6161 43.8514
R14454 gnd.n6161 gnd.n6160 43.8514
R14455 gnd.n6160 gnd.n764 43.8514
R14456 gnd.n6154 gnd.n764 43.8514
R14457 gnd.n6154 gnd.n6153 43.8514
R14458 gnd.n6153 gnd.n6152 43.8514
R14459 gnd.n6152 gnd.n772 43.8514
R14460 gnd.n6146 gnd.n772 43.8514
R14461 gnd.n6146 gnd.n6145 43.8514
R14462 gnd.n6145 gnd.n6144 43.8514
R14463 gnd.n6144 gnd.n780 43.8514
R14464 gnd.n6138 gnd.n780 43.8514
R14465 gnd.n6138 gnd.n6137 43.8514
R14466 gnd.n6137 gnd.n6136 43.8514
R14467 gnd.n6136 gnd.n788 43.8514
R14468 gnd.n6130 gnd.n788 43.8514
R14469 gnd.n6130 gnd.n6129 43.8514
R14470 gnd.n6129 gnd.n6128 43.8514
R14471 gnd.n6128 gnd.n796 43.8514
R14472 gnd.n6122 gnd.n796 43.8514
R14473 gnd.n6122 gnd.n6121 43.8514
R14474 gnd.n6121 gnd.n6120 43.8514
R14475 gnd.n6120 gnd.n804 43.8514
R14476 gnd.n6114 gnd.n804 43.8514
R14477 gnd.n6114 gnd.n6113 43.8514
R14478 gnd.n6113 gnd.n6112 43.8514
R14479 gnd.n6112 gnd.n812 43.8514
R14480 gnd.n6106 gnd.n812 43.8514
R14481 gnd.n6106 gnd.n6105 43.8514
R14482 gnd.n6105 gnd.n6104 43.8514
R14483 gnd.n6104 gnd.n820 43.8514
R14484 gnd.n6098 gnd.n820 43.8514
R14485 gnd.n6098 gnd.n6097 43.8514
R14486 gnd.n6097 gnd.n6096 43.8514
R14487 gnd.n6096 gnd.n828 43.8514
R14488 gnd.n6090 gnd.n828 43.8514
R14489 gnd.n6090 gnd.n6089 43.8514
R14490 gnd.n6089 gnd.n6088 43.8514
R14491 gnd.n6088 gnd.n836 43.8514
R14492 gnd.n6082 gnd.n836 43.8514
R14493 gnd.n6082 gnd.n6081 43.8514
R14494 gnd.n6081 gnd.n6080 43.8514
R14495 gnd.n6080 gnd.n844 43.8514
R14496 gnd.n6074 gnd.n844 43.8514
R14497 gnd.n6074 gnd.n6073 43.8514
R14498 gnd.n6073 gnd.n6072 43.8514
R14499 gnd.n6072 gnd.n852 43.8514
R14500 gnd.n6066 gnd.n852 43.8514
R14501 gnd.n6066 gnd.n6065 43.8514
R14502 gnd.n6065 gnd.n6064 43.8514
R14503 gnd.n3731 gnd.n3730 42.2793
R14504 gnd.n1410 gnd.n1409 42.2793
R14505 gnd.n934 gnd.n933 42.2793
R14506 gnd.n1336 gnd.n1335 42.2793
R14507 gnd.n2283 gnd.n907 42.2793
R14508 gnd.n7083 gnd.n7079 42.2793
R14509 gnd.n2814 gnd.n2813 42.2793
R14510 gnd.n3834 gnd.n3833 42.2793
R14511 gnd.n3100 gnd.n3099 42.2793
R14512 gnd.n7121 gnd.n158 42.2793
R14513 gnd.n7158 gnd.n7157 42.2793
R14514 gnd.n4084 gnd.n4083 42.2793
R14515 gnd.n4060 gnd.n4059 42.2793
R14516 gnd.n3983 gnd.n3982 42.2793
R14517 gnd.n3710 gnd.n3709 42.2793
R14518 gnd.n5551 gnd.n5550 42.2793
R14519 gnd.n6056 gnd.n2318 42.0631
R14520 gnd.n94 gnd.n83 42.0631
R14521 gnd.n3506 gnd.n3505 41.6274
R14522 gnd.n5355 gnd.n5354 41.6274
R14523 gnd.n3515 gnd.n3514 40.8975
R14524 gnd.n5358 gnd.n5357 40.8975
R14525 gnd.n3147 gnd.n3070 36.9518
R14526 gnd.n4586 gnd.n3620 36.9518
R14527 gnd.n3514 gnd.n3513 35.055
R14528 gnd.n3509 gnd.n3508 35.055
R14529 gnd.n5347 gnd.n5346 35.055
R14530 gnd.n5357 gnd.n5343 35.055
R14531 gnd.n1472 gnd.n1366 31.8661
R14532 gnd.n1472 gnd.n1471 31.8661
R14533 gnd.n1480 gnd.n1355 31.8661
R14534 gnd.n1488 gnd.n1355 31.8661
R14535 gnd.n1488 gnd.n1349 31.8661
R14536 gnd.n1496 gnd.n1349 31.8661
R14537 gnd.n1496 gnd.n1342 31.8661
R14538 gnd.n1534 gnd.n1342 31.8661
R14539 gnd.n1544 gnd.n1275 31.8661
R14540 gnd.n4459 gnd.n2537 31.8661
R14541 gnd.n4464 gnd.n4462 31.8661
R14542 gnd.n4464 gnd.n4463 31.8661
R14543 gnd.n4473 gnd.n4472 31.8661
R14544 gnd.n5794 gnd.n2649 31.8661
R14545 gnd.n5788 gnd.n5787 31.8661
R14546 gnd.n5787 gnd.n5786 31.8661
R14547 gnd.n5780 gnd.n2667 31.8661
R14548 gnd.n5434 gnd.n3151 30.4395
R14549 gnd.n4665 gnd.n4664 30.4395
R14550 gnd.n6064 gnd.n860 26.311
R14551 gnd.n3730 gnd.n3729 25.7944
R14552 gnd.n1335 gnd.n1334 25.7944
R14553 gnd.n907 gnd.n906 25.7944
R14554 gnd.n7079 gnd.n7078 25.7944
R14555 gnd.n2813 gnd.n2812 25.7944
R14556 gnd.n3833 gnd.n3832 25.7944
R14557 gnd.n3070 gnd.n3069 25.7944
R14558 gnd.n3099 gnd.n3098 25.7944
R14559 gnd.n158 gnd.n157 25.7944
R14560 gnd.n7157 gnd.n7156 25.7944
R14561 gnd.n4083 gnd.n4082 25.7944
R14562 gnd.n4059 gnd.n4058 25.7944
R14563 gnd.n3982 gnd.n3981 25.7944
R14564 gnd.n3709 gnd.n3708 25.7944
R14565 gnd.n3620 gnd.n3619 25.7944
R14566 gnd.n5550 gnd.n5549 25.7944
R14567 gnd.n1556 gnd.n1276 24.8557
R14568 gnd.n1566 gnd.n1259 24.8557
R14569 gnd.n1262 gnd.n1250 24.8557
R14570 gnd.n1587 gnd.n1251 24.8557
R14571 gnd.n1597 gnd.n1231 24.8557
R14572 gnd.n1607 gnd.n1606 24.8557
R14573 gnd.n1217 gnd.n1215 24.8557
R14574 gnd.n1638 gnd.n1637 24.8557
R14575 gnd.n1653 gnd.n1200 24.8557
R14576 gnd.n1707 gnd.n1139 24.8557
R14577 gnd.n1663 gnd.n1140 24.8557
R14578 gnd.n1700 gnd.n1151 24.8557
R14579 gnd.n1189 gnd.n1188 24.8557
R14580 gnd.n1694 gnd.n1693 24.8557
R14581 gnd.n1175 gnd.n1162 24.8557
R14582 gnd.n1733 gnd.n1732 24.8557
R14583 gnd.n1743 gnd.n1083 24.8557
R14584 gnd.n1755 gnd.n1075 24.8557
R14585 gnd.n1754 gnd.n1063 24.8557
R14586 gnd.n1773 gnd.n1772 24.8557
R14587 gnd.n1783 gnd.n1056 24.8557
R14588 gnd.n1794 gnd.n1044 24.8557
R14589 gnd.n1820 gnd.n1819 24.8557
R14590 gnd.n1830 gnd.n1030 24.8557
R14591 gnd.n1842 gnd.n1022 24.8557
R14592 gnd.n1860 gnd.n1859 24.8557
R14593 gnd.n1013 gnd.n1002 24.8557
R14594 gnd.n1881 gnd.n990 24.8557
R14595 gnd.n1909 gnd.n1908 24.8557
R14596 gnd.n1920 gnd.n975 24.8557
R14597 gnd.n1931 gnd.n968 24.8557
R14598 gnd.n1930 gnd.n956 24.8557
R14599 gnd.n2203 gnd.n2202 24.8557
R14600 gnd.n2225 gnd.n941 24.8557
R14601 gnd.n3555 gnd.n3554 23.855
R14602 gnd.n3150 gnd.n3149 23.855
R14603 gnd.n3557 gnd.n3556 23.855
R14604 gnd.n5362 gnd.n5361 23.855
R14605 gnd.n1577 gnd.t280 23.2624
R14606 gnd.n1278 gnd.t47 22.6251
R14607 gnd.t278 gnd.n1283 21.3504
R14608 gnd.n6056 gnd.n6055 21.0318
R14609 gnd.n4247 gnd.n2321 21.0318
R14610 gnd.n4241 gnd.n2332 21.0318
R14611 gnd.n6043 gnd.n2341 21.0318
R14612 gnd.n4235 gnd.n2344 21.0318
R14613 gnd.n6037 gnd.n2352 21.0318
R14614 gnd.n6031 gnd.n2363 21.0318
R14615 gnd.n4223 gnd.n2366 21.0318
R14616 gnd.n6025 gnd.n2374 21.0318
R14617 gnd.n4278 gnd.n2377 21.0318
R14618 gnd.n4286 gnd.n2387 21.0318
R14619 gnd.n6013 gnd.n2395 21.0318
R14620 gnd.n6007 gnd.n2406 21.0318
R14621 gnd.n4304 gnd.n2409 21.0318
R14622 gnd.n6000 gnd.n2415 21.0318
R14623 gnd.n4352 gnd.n2418 21.0318
R14624 gnd.n4312 gnd.n2428 21.0318
R14625 gnd.n5987 gnd.n2433 21.0318
R14626 gnd.n4327 gnd.n4326 21.0318
R14627 gnd.n5981 gnd.n2442 21.0318
R14628 gnd.n5974 gnd.n2450 21.0318
R14629 gnd.n4389 gnd.n2453 21.0318
R14630 gnd.n4397 gnd.n2463 21.0318
R14631 gnd.n5962 gnd.n2471 21.0318
R14632 gnd.n4405 gnd.n3919 21.0318
R14633 gnd.n5956 gnd.n2481 21.0318
R14634 gnd.n5950 gnd.n2492 21.0318
R14635 gnd.n4441 gnd.n2495 21.0318
R14636 gnd.n4421 gnd.n2505 21.0318
R14637 gnd.n5938 gnd.n2513 21.0318
R14638 gnd.n4430 gnd.n2516 21.0318
R14639 gnd.n5932 gnd.n2524 21.0318
R14640 gnd.n5926 gnd.n2534 21.0318
R14641 gnd.n5779 gnd.n2670 21.0318
R14642 gnd.n5773 gnd.n2682 21.0318
R14643 gnd.n5594 gnd.n5593 21.0318
R14644 gnd.n5604 gnd.n2794 21.0318
R14645 gnd.n5603 gnd.n2772 21.0318
R14646 gnd.n2776 gnd.n2763 21.0318
R14647 gnd.n5625 gnd.n2765 21.0318
R14648 gnd.n5640 gnd.n2747 21.0318
R14649 gnd.n5668 gnd.n5666 21.0318
R14650 gnd.n5631 gnd.n2738 21.0318
R14651 gnd.n5678 gnd.n2741 21.0318
R14652 gnd.n5744 gnd.n2704 21.0318
R14653 gnd.n5747 gnd.n2707 21.0318
R14654 gnd.n6980 gnd.n236 21.0318
R14655 gnd.n5717 gnd.n5716 21.0318
R14656 gnd.n5732 gnd.n2721 21.0318
R14657 gnd.n5727 gnd.n5726 21.0318
R14658 gnd.n5708 gnd.n255 21.0318
R14659 gnd.n6961 gnd.n6960 21.0318
R14660 gnd.n6965 gnd.n251 21.0318
R14661 gnd.n5700 gnd.n220 21.0318
R14662 gnd.n6951 gnd.n211 21.0318
R14663 gnd.n6997 gnd.n214 21.0318
R14664 gnd.n7005 gnd.n205 21.0318
R14665 gnd.n6941 gnd.n6940 21.0318
R14666 gnd.n7013 gnd.n197 21.0318
R14667 gnd.n6915 gnd.n188 21.0318
R14668 gnd.n6932 gnd.n179 21.0318
R14669 gnd.n7029 gnd.n182 21.0318
R14670 gnd.n6926 gnd.n169 21.0318
R14671 gnd.n7039 gnd.n171 21.0318
R14672 gnd.n7114 gnd.n81 21.0318
R14673 gnd.n7193 gnd.n83 21.0318
R14674 gnd.t25 gnd.n1003 20.7131
R14675 gnd.n4295 gnd.t12 20.7131
R14676 gnd.t246 gnd.n2445 20.7131
R14677 gnd.t164 gnd.n233 20.7131
R14678 gnd.n6989 gnd.t173 20.7131
R14679 gnd.n4459 gnd.n3680 20.3945
R14680 gnd.n2667 gnd.n2659 20.3945
R14681 gnd.t27 gnd.n1037 20.0758
R14682 gnd.n4229 gnd.t212 20.0758
R14683 gnd.t196 gnd.n2484 20.0758
R14684 gnd.n5641 gnd.t175 20.0758
R14685 gnd.n7021 gnd.t10 20.0758
R14686 gnd.n3502 gnd.t146 19.8005
R14687 gnd.n3502 gnd.t85 19.8005
R14688 gnd.n3503 gnd.t127 19.8005
R14689 gnd.n3503 gnd.t98 19.8005
R14690 gnd.n5351 gnd.t75 19.8005
R14691 gnd.n5351 gnd.t137 19.8005
R14692 gnd.n5352 gnd.t101 19.8005
R14693 gnd.n5352 gnd.t124 19.8005
R14694 gnd.n3499 gnd.n3498 19.5087
R14695 gnd.n3512 gnd.n3499 19.5087
R14696 gnd.n3510 gnd.n3501 19.5087
R14697 gnd.n5356 gnd.n5350 19.5087
R14698 gnd.n1744 gnd.t31 19.4385
R14699 gnd.n4517 gnd.n4516 19.3944
R14700 gnd.n4516 gnd.n4515 19.3944
R14701 gnd.n4515 gnd.n3741 19.3944
R14702 gnd.n4511 gnd.n3741 19.3944
R14703 gnd.n4511 gnd.n4510 19.3944
R14704 gnd.n4510 gnd.n4509 19.3944
R14705 gnd.n4509 gnd.n3492 19.3944
R14706 gnd.n4679 gnd.n3492 19.3944
R14707 gnd.n4679 gnd.n3489 19.3944
R14708 gnd.n4697 gnd.n3489 19.3944
R14709 gnd.n4697 gnd.n3490 19.3944
R14710 gnd.n4693 gnd.n3490 19.3944
R14711 gnd.n4693 gnd.n4692 19.3944
R14712 gnd.n4692 gnd.n4691 19.3944
R14713 gnd.n4691 gnd.n4686 19.3944
R14714 gnd.n4687 gnd.n4686 19.3944
R14715 gnd.n4687 gnd.n3446 19.3944
R14716 gnd.n4766 gnd.n3446 19.3944
R14717 gnd.n4766 gnd.n3443 19.3944
R14718 gnd.n4777 gnd.n3443 19.3944
R14719 gnd.n4777 gnd.n3444 19.3944
R14720 gnd.n4773 gnd.n3444 19.3944
R14721 gnd.n4773 gnd.n4772 19.3944
R14722 gnd.n4772 gnd.n3403 19.3944
R14723 gnd.n4852 gnd.n3403 19.3944
R14724 gnd.n4852 gnd.n3400 19.3944
R14725 gnd.n4892 gnd.n3400 19.3944
R14726 gnd.n4892 gnd.n3401 19.3944
R14727 gnd.n4888 gnd.n3401 19.3944
R14728 gnd.n4888 gnd.n4887 19.3944
R14729 gnd.n4887 gnd.n4886 19.3944
R14730 gnd.n4886 gnd.n4859 19.3944
R14731 gnd.n4882 gnd.n4859 19.3944
R14732 gnd.n4882 gnd.n4881 19.3944
R14733 gnd.n4881 gnd.n4880 19.3944
R14734 gnd.n4880 gnd.n4864 19.3944
R14735 gnd.n4876 gnd.n4864 19.3944
R14736 gnd.n4876 gnd.n4875 19.3944
R14737 gnd.n4875 gnd.n4874 19.3944
R14738 gnd.n4874 gnd.n4871 19.3944
R14739 gnd.n4871 gnd.n3315 19.3944
R14740 gnd.n5029 gnd.n3315 19.3944
R14741 gnd.n5029 gnd.n3312 19.3944
R14742 gnd.n5069 gnd.n3312 19.3944
R14743 gnd.n5069 gnd.n3313 19.3944
R14744 gnd.n5065 gnd.n3313 19.3944
R14745 gnd.n5065 gnd.n5064 19.3944
R14746 gnd.n5064 gnd.n5063 19.3944
R14747 gnd.n5063 gnd.n5037 19.3944
R14748 gnd.n5059 gnd.n5037 19.3944
R14749 gnd.n5059 gnd.n5058 19.3944
R14750 gnd.n5058 gnd.n5057 19.3944
R14751 gnd.n5057 gnd.n5041 19.3944
R14752 gnd.n5053 gnd.n5041 19.3944
R14753 gnd.n5053 gnd.n5052 19.3944
R14754 gnd.n5052 gnd.n5051 19.3944
R14755 gnd.n5051 gnd.n5048 19.3944
R14756 gnd.n5048 gnd.n3227 19.3944
R14757 gnd.n5206 gnd.n3227 19.3944
R14758 gnd.n5206 gnd.n3224 19.3944
R14759 gnd.n5222 gnd.n3224 19.3944
R14760 gnd.n5222 gnd.n3225 19.3944
R14761 gnd.n5218 gnd.n3225 19.3944
R14762 gnd.n5218 gnd.n5217 19.3944
R14763 gnd.n5217 gnd.n5216 19.3944
R14764 gnd.n5216 gnd.n5213 19.3944
R14765 gnd.n5213 gnd.n3180 19.3944
R14766 gnd.n5298 gnd.n3180 19.3944
R14767 gnd.n5298 gnd.n3177 19.3944
R14768 gnd.n5319 gnd.n3177 19.3944
R14769 gnd.n5319 gnd.n3178 19.3944
R14770 gnd.n5315 gnd.n3178 19.3944
R14771 gnd.n5315 gnd.n5314 19.3944
R14772 gnd.n5314 gnd.n5313 19.3944
R14773 gnd.n5313 gnd.n5310 19.3944
R14774 gnd.n5310 gnd.n2969 19.3944
R14775 gnd.n5512 gnd.n2969 19.3944
R14776 gnd.n5512 gnd.n2967 19.3944
R14777 gnd.n5517 gnd.n2967 19.3944
R14778 gnd.n5517 gnd.n2958 19.3944
R14779 gnd.n5535 gnd.n2958 19.3944
R14780 gnd.n5536 gnd.n5535 19.3944
R14781 gnd.n4523 gnd.n4522 19.3944
R14782 gnd.n4522 gnd.n4521 19.3944
R14783 gnd.n4521 gnd.n3736 19.3944
R14784 gnd.n3887 gnd.n3886 19.3944
R14785 gnd.n3886 gnd.n3776 19.3944
R14786 gnd.n3879 gnd.n3776 19.3944
R14787 gnd.n3879 gnd.n3878 19.3944
R14788 gnd.n3878 gnd.n3792 19.3944
R14789 gnd.n3871 gnd.n3792 19.3944
R14790 gnd.n3871 gnd.n3870 19.3944
R14791 gnd.n3870 gnd.n3802 19.3944
R14792 gnd.n3863 gnd.n3802 19.3944
R14793 gnd.n3863 gnd.n3862 19.3944
R14794 gnd.n3862 gnd.n3815 19.3944
R14795 gnd.n3855 gnd.n3815 19.3944
R14796 gnd.n3855 gnd.n3854 19.3944
R14797 gnd.n3854 gnd.n3825 19.3944
R14798 gnd.n3847 gnd.n3825 19.3944
R14799 gnd.n3847 gnd.n3846 19.3944
R14800 gnd.n3846 gnd.n3720 19.3944
R14801 gnd.n4534 gnd.n3720 19.3944
R14802 gnd.n4534 gnd.n4533 19.3944
R14803 gnd.n4533 gnd.n4532 19.3944
R14804 gnd.n4532 gnd.n3724 19.3944
R14805 gnd.n4528 gnd.n3724 19.3944
R14806 gnd.n4528 gnd.n4527 19.3944
R14807 gnd.n4527 gnd.n4526 19.3944
R14808 gnd.n1459 gnd.n1458 19.3944
R14809 gnd.n1458 gnd.n1457 19.3944
R14810 gnd.n1457 gnd.n1456 19.3944
R14811 gnd.n1456 gnd.n1454 19.3944
R14812 gnd.n1454 gnd.n1451 19.3944
R14813 gnd.n1451 gnd.n1450 19.3944
R14814 gnd.n1450 gnd.n1447 19.3944
R14815 gnd.n1447 gnd.n1446 19.3944
R14816 gnd.n1446 gnd.n1443 19.3944
R14817 gnd.n1443 gnd.n1442 19.3944
R14818 gnd.n1442 gnd.n1439 19.3944
R14819 gnd.n1439 gnd.n1438 19.3944
R14820 gnd.n1438 gnd.n1435 19.3944
R14821 gnd.n1435 gnd.n1434 19.3944
R14822 gnd.n1434 gnd.n1431 19.3944
R14823 gnd.n1431 gnd.n1430 19.3944
R14824 gnd.n1430 gnd.n1427 19.3944
R14825 gnd.n1427 gnd.n1426 19.3944
R14826 gnd.n1426 gnd.n1423 19.3944
R14827 gnd.n1423 gnd.n1422 19.3944
R14828 gnd.n1422 gnd.n1419 19.3944
R14829 gnd.n1419 gnd.n1418 19.3944
R14830 gnd.n1415 gnd.n1414 19.3944
R14831 gnd.n1414 gnd.n1370 19.3944
R14832 gnd.n1465 gnd.n1370 19.3944
R14833 gnd.n2233 gnd.n2232 19.3944
R14834 gnd.n2232 gnd.n2229 19.3944
R14835 gnd.n2229 gnd.n2228 19.3944
R14836 gnd.n2278 gnd.n2277 19.3944
R14837 gnd.n2277 gnd.n2276 19.3944
R14838 gnd.n2276 gnd.n2273 19.3944
R14839 gnd.n2273 gnd.n2272 19.3944
R14840 gnd.n2272 gnd.n2269 19.3944
R14841 gnd.n2269 gnd.n2268 19.3944
R14842 gnd.n2268 gnd.n2265 19.3944
R14843 gnd.n2265 gnd.n2264 19.3944
R14844 gnd.n2264 gnd.n2261 19.3944
R14845 gnd.n2261 gnd.n2260 19.3944
R14846 gnd.n2260 gnd.n2257 19.3944
R14847 gnd.n2257 gnd.n2256 19.3944
R14848 gnd.n2256 gnd.n2253 19.3944
R14849 gnd.n2253 gnd.n2252 19.3944
R14850 gnd.n2252 gnd.n2249 19.3944
R14851 gnd.n2249 gnd.n2248 19.3944
R14852 gnd.n2248 gnd.n2245 19.3944
R14853 gnd.n2245 gnd.n2244 19.3944
R14854 gnd.n2244 gnd.n2241 19.3944
R14855 gnd.n2241 gnd.n2240 19.3944
R14856 gnd.n2240 gnd.n2237 19.3944
R14857 gnd.n2237 gnd.n2236 19.3944
R14858 gnd.n1558 gnd.n1267 19.3944
R14859 gnd.n1568 gnd.n1267 19.3944
R14860 gnd.n1569 gnd.n1568 19.3944
R14861 gnd.n1569 gnd.n1248 19.3944
R14862 gnd.n1589 gnd.n1248 19.3944
R14863 gnd.n1589 gnd.n1240 19.3944
R14864 gnd.n1599 gnd.n1240 19.3944
R14865 gnd.n1600 gnd.n1599 19.3944
R14866 gnd.n1601 gnd.n1600 19.3944
R14867 gnd.n1601 gnd.n1223 19.3944
R14868 gnd.n1618 gnd.n1223 19.3944
R14869 gnd.n1621 gnd.n1618 19.3944
R14870 gnd.n1621 gnd.n1620 19.3944
R14871 gnd.n1620 gnd.n1196 19.3944
R14872 gnd.n1660 gnd.n1196 19.3944
R14873 gnd.n1660 gnd.n1193 19.3944
R14874 gnd.n1666 gnd.n1193 19.3944
R14875 gnd.n1667 gnd.n1666 19.3944
R14876 gnd.n1667 gnd.n1191 19.3944
R14877 gnd.n1673 gnd.n1191 19.3944
R14878 gnd.n1676 gnd.n1673 19.3944
R14879 gnd.n1678 gnd.n1676 19.3944
R14880 gnd.n1684 gnd.n1678 19.3944
R14881 gnd.n1684 gnd.n1683 19.3944
R14882 gnd.n1683 gnd.n1078 19.3944
R14883 gnd.n1750 gnd.n1078 19.3944
R14884 gnd.n1751 gnd.n1750 19.3944
R14885 gnd.n1751 gnd.n1071 19.3944
R14886 gnd.n1762 gnd.n1071 19.3944
R14887 gnd.n1763 gnd.n1762 19.3944
R14888 gnd.n1763 gnd.n1054 19.3944
R14889 gnd.n1054 gnd.n1052 19.3944
R14890 gnd.n1787 gnd.n1052 19.3944
R14891 gnd.n1788 gnd.n1787 19.3944
R14892 gnd.n1788 gnd.n1025 19.3944
R14893 gnd.n1837 gnd.n1025 19.3944
R14894 gnd.n1838 gnd.n1837 19.3944
R14895 gnd.n1838 gnd.n1018 19.3944
R14896 gnd.n1849 gnd.n1018 19.3944
R14897 gnd.n1850 gnd.n1849 19.3944
R14898 gnd.n1850 gnd.n1001 19.3944
R14899 gnd.n1001 gnd.n999 19.3944
R14900 gnd.n1874 gnd.n999 19.3944
R14901 gnd.n1875 gnd.n1874 19.3944
R14902 gnd.n1875 gnd.n971 19.3944
R14903 gnd.n1926 gnd.n971 19.3944
R14904 gnd.n1927 gnd.n1926 19.3944
R14905 gnd.n1927 gnd.n964 19.3944
R14906 gnd.n2194 gnd.n964 19.3944
R14907 gnd.n2195 gnd.n2194 19.3944
R14908 gnd.n2195 gnd.n945 19.3944
R14909 gnd.n2220 gnd.n945 19.3944
R14910 gnd.n2220 gnd.n946 19.3944
R14911 gnd.n1549 gnd.n1548 19.3944
R14912 gnd.n1548 gnd.n1281 19.3944
R14913 gnd.n1304 gnd.n1281 19.3944
R14914 gnd.n1307 gnd.n1304 19.3944
R14915 gnd.n1307 gnd.n1300 19.3944
R14916 gnd.n1311 gnd.n1300 19.3944
R14917 gnd.n1314 gnd.n1311 19.3944
R14918 gnd.n1317 gnd.n1314 19.3944
R14919 gnd.n1317 gnd.n1298 19.3944
R14920 gnd.n1321 gnd.n1298 19.3944
R14921 gnd.n1324 gnd.n1321 19.3944
R14922 gnd.n1327 gnd.n1324 19.3944
R14923 gnd.n1327 gnd.n1296 19.3944
R14924 gnd.n1331 gnd.n1296 19.3944
R14925 gnd.n1554 gnd.n1553 19.3944
R14926 gnd.n1553 gnd.n1257 19.3944
R14927 gnd.n1579 gnd.n1257 19.3944
R14928 gnd.n1579 gnd.n1255 19.3944
R14929 gnd.n1585 gnd.n1255 19.3944
R14930 gnd.n1585 gnd.n1584 19.3944
R14931 gnd.n1584 gnd.n1229 19.3944
R14932 gnd.n1609 gnd.n1229 19.3944
R14933 gnd.n1609 gnd.n1227 19.3944
R14934 gnd.n1613 gnd.n1227 19.3944
R14935 gnd.n1613 gnd.n1207 19.3944
R14936 gnd.n1640 gnd.n1207 19.3944
R14937 gnd.n1640 gnd.n1205 19.3944
R14938 gnd.n1650 gnd.n1205 19.3944
R14939 gnd.n1650 gnd.n1649 19.3944
R14940 gnd.n1649 gnd.n1648 19.3944
R14941 gnd.n1648 gnd.n1154 19.3944
R14942 gnd.n1698 gnd.n1154 19.3944
R14943 gnd.n1698 gnd.n1697 19.3944
R14944 gnd.n1697 gnd.n1696 19.3944
R14945 gnd.n1696 gnd.n1158 19.3944
R14946 gnd.n1178 gnd.n1158 19.3944
R14947 gnd.n1178 gnd.n1088 19.3944
R14948 gnd.n1735 gnd.n1088 19.3944
R14949 gnd.n1735 gnd.n1086 19.3944
R14950 gnd.n1741 gnd.n1086 19.3944
R14951 gnd.n1741 gnd.n1740 19.3944
R14952 gnd.n1740 gnd.n1061 19.3944
R14953 gnd.n1775 gnd.n1061 19.3944
R14954 gnd.n1775 gnd.n1059 19.3944
R14955 gnd.n1781 gnd.n1059 19.3944
R14956 gnd.n1781 gnd.n1780 19.3944
R14957 gnd.n1780 gnd.n1035 19.3944
R14958 gnd.n1822 gnd.n1035 19.3944
R14959 gnd.n1822 gnd.n1033 19.3944
R14960 gnd.n1828 gnd.n1033 19.3944
R14961 gnd.n1828 gnd.n1827 19.3944
R14962 gnd.n1827 gnd.n1008 19.3944
R14963 gnd.n1862 gnd.n1008 19.3944
R14964 gnd.n1862 gnd.n1006 19.3944
R14965 gnd.n1868 gnd.n1006 19.3944
R14966 gnd.n1868 gnd.n1867 19.3944
R14967 gnd.n1867 gnd.n981 19.3944
R14968 gnd.n1911 gnd.n981 19.3944
R14969 gnd.n1911 gnd.n979 19.3944
R14970 gnd.n1917 gnd.n979 19.3944
R14971 gnd.n1917 gnd.n1916 19.3944
R14972 gnd.n1916 gnd.n954 19.3944
R14973 gnd.n2205 gnd.n954 19.3944
R14974 gnd.n2205 gnd.n952 19.3944
R14975 gnd.n2213 gnd.n952 19.3944
R14976 gnd.n2213 gnd.n2212 19.3944
R14977 gnd.n2212 gnd.n2211 19.3944
R14978 gnd.n2314 gnd.n2313 19.3944
R14979 gnd.n2313 gnd.n893 19.3944
R14980 gnd.n2309 gnd.n893 19.3944
R14981 gnd.n2309 gnd.n2306 19.3944
R14982 gnd.n2306 gnd.n2303 19.3944
R14983 gnd.n2303 gnd.n2302 19.3944
R14984 gnd.n2302 gnd.n2299 19.3944
R14985 gnd.n2299 gnd.n2298 19.3944
R14986 gnd.n2298 gnd.n2295 19.3944
R14987 gnd.n2295 gnd.n2294 19.3944
R14988 gnd.n2294 gnd.n2291 19.3944
R14989 gnd.n2291 gnd.n2290 19.3944
R14990 gnd.n2290 gnd.n2287 19.3944
R14991 gnd.n2287 gnd.n2286 19.3944
R14992 gnd.n1469 gnd.n1368 19.3944
R14993 gnd.n1469 gnd.n1359 19.3944
R14994 gnd.n1482 gnd.n1359 19.3944
R14995 gnd.n1482 gnd.n1357 19.3944
R14996 gnd.n1486 gnd.n1357 19.3944
R14997 gnd.n1486 gnd.n1347 19.3944
R14998 gnd.n1498 gnd.n1347 19.3944
R14999 gnd.n1498 gnd.n1345 19.3944
R15000 gnd.n1532 gnd.n1345 19.3944
R15001 gnd.n1532 gnd.n1531 19.3944
R15002 gnd.n1531 gnd.n1530 19.3944
R15003 gnd.n1530 gnd.n1529 19.3944
R15004 gnd.n1529 gnd.n1526 19.3944
R15005 gnd.n1526 gnd.n1525 19.3944
R15006 gnd.n1525 gnd.n1524 19.3944
R15007 gnd.n1524 gnd.n1522 19.3944
R15008 gnd.n1522 gnd.n1521 19.3944
R15009 gnd.n1521 gnd.n1518 19.3944
R15010 gnd.n1518 gnd.n1517 19.3944
R15011 gnd.n1517 gnd.n1516 19.3944
R15012 gnd.n1516 gnd.n1514 19.3944
R15013 gnd.n1514 gnd.n1213 19.3944
R15014 gnd.n1629 gnd.n1213 19.3944
R15015 gnd.n1629 gnd.n1211 19.3944
R15016 gnd.n1635 gnd.n1211 19.3944
R15017 gnd.n1635 gnd.n1634 19.3944
R15018 gnd.n1634 gnd.n1135 19.3944
R15019 gnd.n1709 gnd.n1135 19.3944
R15020 gnd.n1709 gnd.n1136 19.3944
R15021 gnd.n1183 gnd.n1182 19.3944
R15022 gnd.n1186 gnd.n1185 19.3944
R15023 gnd.n1173 gnd.n1172 19.3944
R15024 gnd.n1728 gnd.n1093 19.3944
R15025 gnd.n1728 gnd.n1727 19.3944
R15026 gnd.n1727 gnd.n1726 19.3944
R15027 gnd.n1726 gnd.n1724 19.3944
R15028 gnd.n1724 gnd.n1723 19.3944
R15029 gnd.n1723 gnd.n1721 19.3944
R15030 gnd.n1721 gnd.n1720 19.3944
R15031 gnd.n1720 gnd.n1042 19.3944
R15032 gnd.n1796 gnd.n1042 19.3944
R15033 gnd.n1796 gnd.n1040 19.3944
R15034 gnd.n1815 gnd.n1040 19.3944
R15035 gnd.n1815 gnd.n1814 19.3944
R15036 gnd.n1814 gnd.n1813 19.3944
R15037 gnd.n1813 gnd.n1811 19.3944
R15038 gnd.n1811 gnd.n1810 19.3944
R15039 gnd.n1810 gnd.n1808 19.3944
R15040 gnd.n1808 gnd.n1807 19.3944
R15041 gnd.n1807 gnd.n988 19.3944
R15042 gnd.n1883 gnd.n988 19.3944
R15043 gnd.n1883 gnd.n986 19.3944
R15044 gnd.n1906 gnd.n986 19.3944
R15045 gnd.n1906 gnd.n1905 19.3944
R15046 gnd.n1905 gnd.n1904 19.3944
R15047 gnd.n1904 gnd.n1901 19.3944
R15048 gnd.n1901 gnd.n1900 19.3944
R15049 gnd.n1900 gnd.n1898 19.3944
R15050 gnd.n1898 gnd.n1897 19.3944
R15051 gnd.n1897 gnd.n1895 19.3944
R15052 gnd.n1895 gnd.n940 19.3944
R15053 gnd.n1474 gnd.n1364 19.3944
R15054 gnd.n1474 gnd.n1362 19.3944
R15055 gnd.n1478 gnd.n1362 19.3944
R15056 gnd.n1478 gnd.n1353 19.3944
R15057 gnd.n1490 gnd.n1353 19.3944
R15058 gnd.n1490 gnd.n1351 19.3944
R15059 gnd.n1494 gnd.n1351 19.3944
R15060 gnd.n1494 gnd.n1340 19.3944
R15061 gnd.n1536 gnd.n1340 19.3944
R15062 gnd.n1536 gnd.n1294 19.3944
R15063 gnd.n1542 gnd.n1294 19.3944
R15064 gnd.n1542 gnd.n1541 19.3944
R15065 gnd.n1541 gnd.n1272 19.3944
R15066 gnd.n1563 gnd.n1272 19.3944
R15067 gnd.n1563 gnd.n1265 19.3944
R15068 gnd.n1574 gnd.n1265 19.3944
R15069 gnd.n1574 gnd.n1573 19.3944
R15070 gnd.n1573 gnd.n1246 19.3944
R15071 gnd.n1594 gnd.n1246 19.3944
R15072 gnd.n1594 gnd.n1236 19.3944
R15073 gnd.n1604 gnd.n1236 19.3944
R15074 gnd.n1604 gnd.n1219 19.3944
R15075 gnd.n1625 gnd.n1219 19.3944
R15076 gnd.n1625 gnd.n1624 19.3944
R15077 gnd.n1624 gnd.n1198 19.3944
R15078 gnd.n1655 gnd.n1198 19.3944
R15079 gnd.n1655 gnd.n1143 19.3944
R15080 gnd.n1705 gnd.n1143 19.3944
R15081 gnd.n1705 gnd.n1704 19.3944
R15082 gnd.n1704 gnd.n1703 19.3944
R15083 gnd.n1703 gnd.n1147 19.3944
R15084 gnd.n1165 gnd.n1147 19.3944
R15085 gnd.n1691 gnd.n1165 19.3944
R15086 gnd.n1691 gnd.n1690 19.3944
R15087 gnd.n1690 gnd.n1689 19.3944
R15088 gnd.n1689 gnd.n1169 19.3944
R15089 gnd.n1169 gnd.n1080 19.3944
R15090 gnd.n1746 gnd.n1080 19.3944
R15091 gnd.n1746 gnd.n1073 19.3944
R15092 gnd.n1757 gnd.n1073 19.3944
R15093 gnd.n1757 gnd.n1069 19.3944
R15094 gnd.n1770 gnd.n1069 19.3944
R15095 gnd.n1770 gnd.n1769 19.3944
R15096 gnd.n1769 gnd.n1048 19.3944
R15097 gnd.n1792 gnd.n1048 19.3944
R15098 gnd.n1792 gnd.n1791 19.3944
R15099 gnd.n1791 gnd.n1027 19.3944
R15100 gnd.n1833 gnd.n1027 19.3944
R15101 gnd.n1833 gnd.n1020 19.3944
R15102 gnd.n1844 gnd.n1020 19.3944
R15103 gnd.n1844 gnd.n1016 19.3944
R15104 gnd.n1857 gnd.n1016 19.3944
R15105 gnd.n1857 gnd.n1856 19.3944
R15106 gnd.n1856 gnd.n995 19.3944
R15107 gnd.n1879 gnd.n995 19.3944
R15108 gnd.n1879 gnd.n1878 19.3944
R15109 gnd.n1878 gnd.n973 19.3944
R15110 gnd.n1922 gnd.n973 19.3944
R15111 gnd.n1922 gnd.n966 19.3944
R15112 gnd.n1933 gnd.n966 19.3944
R15113 gnd.n1933 gnd.n962 19.3944
R15114 gnd.n2200 gnd.n962 19.3944
R15115 gnd.n2200 gnd.n2199 19.3944
R15116 gnd.n2199 gnd.n943 19.3944
R15117 gnd.n2223 gnd.n943 19.3944
R15118 gnd.n5564 gnd.n2805 19.3944
R15119 gnd.n5564 gnd.n2800 19.3944
R15120 gnd.n5596 gnd.n2800 19.3944
R15121 gnd.n5596 gnd.n2797 19.3944
R15122 gnd.n5601 gnd.n2797 19.3944
R15123 gnd.n5601 gnd.n2798 19.3944
R15124 gnd.n2798 gnd.n2761 19.3944
R15125 gnd.n5627 gnd.n2761 19.3944
R15126 gnd.n5627 gnd.n2758 19.3944
R15127 gnd.n5638 gnd.n2758 19.3944
R15128 gnd.n5638 gnd.n2759 19.3944
R15129 gnd.n5634 gnd.n2759 19.3944
R15130 gnd.n5634 gnd.n5633 19.3944
R15131 gnd.n5633 gnd.n2713 19.3944
R15132 gnd.n5742 gnd.n2713 19.3944
R15133 gnd.n5742 gnd.n2714 19.3944
R15134 gnd.n5738 gnd.n2714 19.3944
R15135 gnd.n5738 gnd.n5737 19.3944
R15136 gnd.n5737 gnd.n5736 19.3944
R15137 gnd.n5736 gnd.n5734 19.3944
R15138 gnd.n5734 gnd.n52 19.3944
R15139 gnd.n7225 gnd.n52 19.3944
R15140 gnd.n7225 gnd.n7224 19.3944
R15141 gnd.n7224 gnd.n7223 19.3944
R15142 gnd.n7223 gnd.n57 19.3944
R15143 gnd.n7219 gnd.n57 19.3944
R15144 gnd.n7219 gnd.n7218 19.3944
R15145 gnd.n7218 gnd.n7217 19.3944
R15146 gnd.n7217 gnd.n62 19.3944
R15147 gnd.n7213 gnd.n62 19.3944
R15148 gnd.n7213 gnd.n7212 19.3944
R15149 gnd.n7212 gnd.n7211 19.3944
R15150 gnd.n7211 gnd.n67 19.3944
R15151 gnd.n7207 gnd.n67 19.3944
R15152 gnd.n7207 gnd.n7206 19.3944
R15153 gnd.n7206 gnd.n7205 19.3944
R15154 gnd.n7205 gnd.n72 19.3944
R15155 gnd.n7201 gnd.n72 19.3944
R15156 gnd.n7201 gnd.n7200 19.3944
R15157 gnd.n7200 gnd.n7199 19.3944
R15158 gnd.n7199 gnd.n77 19.3944
R15159 gnd.n7195 gnd.n77 19.3944
R15160 gnd.n7108 gnd.n7107 19.3944
R15161 gnd.n7107 gnd.n7106 19.3944
R15162 gnd.n7106 gnd.n7049 19.3944
R15163 gnd.n7102 gnd.n7049 19.3944
R15164 gnd.n7102 gnd.n7101 19.3944
R15165 gnd.n7101 gnd.n7100 19.3944
R15166 gnd.n7100 gnd.n7057 19.3944
R15167 gnd.n7096 gnd.n7057 19.3944
R15168 gnd.n7096 gnd.n7095 19.3944
R15169 gnd.n7095 gnd.n7094 19.3944
R15170 gnd.n7094 gnd.n7065 19.3944
R15171 gnd.n7090 gnd.n7065 19.3944
R15172 gnd.n7090 gnd.n7089 19.3944
R15173 gnd.n7089 gnd.n7088 19.3944
R15174 gnd.n7088 gnd.n7073 19.3944
R15175 gnd.n7084 gnd.n7073 19.3944
R15176 gnd.n2856 gnd.n2850 19.3944
R15177 gnd.n2862 gnd.n2850 19.3944
R15178 gnd.n2862 gnd.n2843 19.3944
R15179 gnd.n2875 gnd.n2843 19.3944
R15180 gnd.n2875 gnd.n2841 19.3944
R15181 gnd.n2881 gnd.n2841 19.3944
R15182 gnd.n2881 gnd.n2834 19.3944
R15183 gnd.n2894 gnd.n2834 19.3944
R15184 gnd.n2894 gnd.n2832 19.3944
R15185 gnd.n2900 gnd.n2832 19.3944
R15186 gnd.n2900 gnd.n2825 19.3944
R15187 gnd.n2913 gnd.n2825 19.3944
R15188 gnd.n2913 gnd.n2823 19.3944
R15189 gnd.n2919 gnd.n2823 19.3944
R15190 gnd.n2919 gnd.n2816 19.3944
R15191 gnd.n2932 gnd.n2816 19.3944
R15192 gnd.n2853 gnd.n2685 19.3944
R15193 gnd.n5771 gnd.n2685 19.3944
R15194 gnd.n5771 gnd.n2686 19.3944
R15195 gnd.n5767 gnd.n2686 19.3944
R15196 gnd.n5767 gnd.n5766 19.3944
R15197 gnd.n5766 gnd.n5765 19.3944
R15198 gnd.n5765 gnd.n2692 19.3944
R15199 gnd.n5761 gnd.n2692 19.3944
R15200 gnd.n5761 gnd.n5760 19.3944
R15201 gnd.n5760 gnd.n5759 19.3944
R15202 gnd.n5759 gnd.n2697 19.3944
R15203 gnd.n5755 gnd.n2697 19.3944
R15204 gnd.n5755 gnd.n5754 19.3944
R15205 gnd.n5754 gnd.n5753 19.3944
R15206 gnd.n5753 gnd.n2702 19.3944
R15207 gnd.n5749 gnd.n2702 19.3944
R15208 gnd.n5749 gnd.n239 19.3944
R15209 gnd.n6978 gnd.n239 19.3944
R15210 gnd.n6978 gnd.n240 19.3944
R15211 gnd.n6974 gnd.n240 19.3944
R15212 gnd.n6974 gnd.n6973 19.3944
R15213 gnd.n6973 gnd.n6972 19.3944
R15214 gnd.n6972 gnd.n246 19.3944
R15215 gnd.n6968 gnd.n246 19.3944
R15216 gnd.n6968 gnd.n6967 19.3944
R15217 gnd.n6967 gnd.n218 19.3944
R15218 gnd.n6991 gnd.n218 19.3944
R15219 gnd.n6991 gnd.n216 19.3944
R15220 gnd.n6995 gnd.n216 19.3944
R15221 gnd.n6995 gnd.n201 19.3944
R15222 gnd.n7007 gnd.n201 19.3944
R15223 gnd.n7007 gnd.n199 19.3944
R15224 gnd.n7011 gnd.n199 19.3944
R15225 gnd.n7011 gnd.n186 19.3944
R15226 gnd.n7023 gnd.n186 19.3944
R15227 gnd.n7023 gnd.n184 19.3944
R15228 gnd.n7027 gnd.n184 19.3944
R15229 gnd.n7027 gnd.n167 19.3944
R15230 gnd.n7041 gnd.n167 19.3944
R15231 gnd.n7041 gnd.n164 19.3944
R15232 gnd.n7112 gnd.n164 19.3944
R15233 gnd.n7112 gnd.n165 19.3944
R15234 gnd.n3780 gnd.n2540 19.3944
R15235 gnd.n3780 gnd.n3779 19.3944
R15236 gnd.n3883 gnd.n3779 19.3944
R15237 gnd.n3883 gnd.n3882 19.3944
R15238 gnd.n3882 gnd.n3787 19.3944
R15239 gnd.n3875 gnd.n3787 19.3944
R15240 gnd.n3875 gnd.n3874 19.3944
R15241 gnd.n3874 gnd.n3798 19.3944
R15242 gnd.n3867 gnd.n3798 19.3944
R15243 gnd.n3867 gnd.n3866 19.3944
R15244 gnd.n3866 gnd.n3809 19.3944
R15245 gnd.n3859 gnd.n3809 19.3944
R15246 gnd.n3859 gnd.n3858 19.3944
R15247 gnd.n3858 gnd.n3821 19.3944
R15248 gnd.n3851 gnd.n3821 19.3944
R15249 gnd.n3851 gnd.n3850 19.3944
R15250 gnd.n6689 gnd.n422 19.3944
R15251 gnd.n6693 gnd.n422 19.3944
R15252 gnd.n6693 gnd.n418 19.3944
R15253 gnd.n6699 gnd.n418 19.3944
R15254 gnd.n6699 gnd.n416 19.3944
R15255 gnd.n6703 gnd.n416 19.3944
R15256 gnd.n6703 gnd.n412 19.3944
R15257 gnd.n6709 gnd.n412 19.3944
R15258 gnd.n6709 gnd.n410 19.3944
R15259 gnd.n6713 gnd.n410 19.3944
R15260 gnd.n6713 gnd.n406 19.3944
R15261 gnd.n6719 gnd.n406 19.3944
R15262 gnd.n6719 gnd.n404 19.3944
R15263 gnd.n6723 gnd.n404 19.3944
R15264 gnd.n6723 gnd.n400 19.3944
R15265 gnd.n6729 gnd.n400 19.3944
R15266 gnd.n6729 gnd.n398 19.3944
R15267 gnd.n6733 gnd.n398 19.3944
R15268 gnd.n6733 gnd.n394 19.3944
R15269 gnd.n6739 gnd.n394 19.3944
R15270 gnd.n6739 gnd.n392 19.3944
R15271 gnd.n6743 gnd.n392 19.3944
R15272 gnd.n6743 gnd.n388 19.3944
R15273 gnd.n6749 gnd.n388 19.3944
R15274 gnd.n6749 gnd.n386 19.3944
R15275 gnd.n6753 gnd.n386 19.3944
R15276 gnd.n6753 gnd.n382 19.3944
R15277 gnd.n6759 gnd.n382 19.3944
R15278 gnd.n6759 gnd.n380 19.3944
R15279 gnd.n6763 gnd.n380 19.3944
R15280 gnd.n6763 gnd.n376 19.3944
R15281 gnd.n6769 gnd.n376 19.3944
R15282 gnd.n6769 gnd.n374 19.3944
R15283 gnd.n6773 gnd.n374 19.3944
R15284 gnd.n6773 gnd.n370 19.3944
R15285 gnd.n6779 gnd.n370 19.3944
R15286 gnd.n6779 gnd.n368 19.3944
R15287 gnd.n6783 gnd.n368 19.3944
R15288 gnd.n6783 gnd.n364 19.3944
R15289 gnd.n6789 gnd.n364 19.3944
R15290 gnd.n6789 gnd.n362 19.3944
R15291 gnd.n6793 gnd.n362 19.3944
R15292 gnd.n6793 gnd.n358 19.3944
R15293 gnd.n6799 gnd.n358 19.3944
R15294 gnd.n6799 gnd.n356 19.3944
R15295 gnd.n6803 gnd.n356 19.3944
R15296 gnd.n6803 gnd.n352 19.3944
R15297 gnd.n6809 gnd.n352 19.3944
R15298 gnd.n6809 gnd.n350 19.3944
R15299 gnd.n6813 gnd.n350 19.3944
R15300 gnd.n6813 gnd.n346 19.3944
R15301 gnd.n6819 gnd.n346 19.3944
R15302 gnd.n6819 gnd.n344 19.3944
R15303 gnd.n6823 gnd.n344 19.3944
R15304 gnd.n6823 gnd.n340 19.3944
R15305 gnd.n6829 gnd.n340 19.3944
R15306 gnd.n6829 gnd.n338 19.3944
R15307 gnd.n6833 gnd.n338 19.3944
R15308 gnd.n6833 gnd.n334 19.3944
R15309 gnd.n6839 gnd.n334 19.3944
R15310 gnd.n6839 gnd.n332 19.3944
R15311 gnd.n6843 gnd.n332 19.3944
R15312 gnd.n6843 gnd.n328 19.3944
R15313 gnd.n6849 gnd.n328 19.3944
R15314 gnd.n6849 gnd.n326 19.3944
R15315 gnd.n6853 gnd.n326 19.3944
R15316 gnd.n6853 gnd.n322 19.3944
R15317 gnd.n6859 gnd.n322 19.3944
R15318 gnd.n6859 gnd.n320 19.3944
R15319 gnd.n6863 gnd.n320 19.3944
R15320 gnd.n6863 gnd.n316 19.3944
R15321 gnd.n6869 gnd.n316 19.3944
R15322 gnd.n6869 gnd.n314 19.3944
R15323 gnd.n6873 gnd.n314 19.3944
R15324 gnd.n6873 gnd.n310 19.3944
R15325 gnd.n6879 gnd.n310 19.3944
R15326 gnd.n6879 gnd.n308 19.3944
R15327 gnd.n6883 gnd.n308 19.3944
R15328 gnd.n6883 gnd.n304 19.3944
R15329 gnd.n6889 gnd.n304 19.3944
R15330 gnd.n6889 gnd.n302 19.3944
R15331 gnd.n6896 gnd.n302 19.3944
R15332 gnd.n6896 gnd.n6895 19.3944
R15333 gnd.n6895 gnd.n299 19.3944
R15334 gnd.n6232 gnd.n693 19.3944
R15335 gnd.n6238 gnd.n693 19.3944
R15336 gnd.n6238 gnd.n691 19.3944
R15337 gnd.n6242 gnd.n691 19.3944
R15338 gnd.n6242 gnd.n687 19.3944
R15339 gnd.n6248 gnd.n687 19.3944
R15340 gnd.n6248 gnd.n685 19.3944
R15341 gnd.n6252 gnd.n685 19.3944
R15342 gnd.n6252 gnd.n681 19.3944
R15343 gnd.n6258 gnd.n681 19.3944
R15344 gnd.n6258 gnd.n679 19.3944
R15345 gnd.n6262 gnd.n679 19.3944
R15346 gnd.n6262 gnd.n675 19.3944
R15347 gnd.n6268 gnd.n675 19.3944
R15348 gnd.n6268 gnd.n673 19.3944
R15349 gnd.n6272 gnd.n673 19.3944
R15350 gnd.n6272 gnd.n669 19.3944
R15351 gnd.n6278 gnd.n669 19.3944
R15352 gnd.n6278 gnd.n667 19.3944
R15353 gnd.n6282 gnd.n667 19.3944
R15354 gnd.n6282 gnd.n663 19.3944
R15355 gnd.n6288 gnd.n663 19.3944
R15356 gnd.n6288 gnd.n661 19.3944
R15357 gnd.n6292 gnd.n661 19.3944
R15358 gnd.n6292 gnd.n657 19.3944
R15359 gnd.n6298 gnd.n657 19.3944
R15360 gnd.n6298 gnd.n655 19.3944
R15361 gnd.n6302 gnd.n655 19.3944
R15362 gnd.n6302 gnd.n651 19.3944
R15363 gnd.n6308 gnd.n651 19.3944
R15364 gnd.n6308 gnd.n649 19.3944
R15365 gnd.n6312 gnd.n649 19.3944
R15366 gnd.n6312 gnd.n645 19.3944
R15367 gnd.n6318 gnd.n645 19.3944
R15368 gnd.n6318 gnd.n643 19.3944
R15369 gnd.n6322 gnd.n643 19.3944
R15370 gnd.n6322 gnd.n639 19.3944
R15371 gnd.n6328 gnd.n639 19.3944
R15372 gnd.n6328 gnd.n637 19.3944
R15373 gnd.n6332 gnd.n637 19.3944
R15374 gnd.n6332 gnd.n633 19.3944
R15375 gnd.n6338 gnd.n633 19.3944
R15376 gnd.n6338 gnd.n631 19.3944
R15377 gnd.n6342 gnd.n631 19.3944
R15378 gnd.n6342 gnd.n627 19.3944
R15379 gnd.n6348 gnd.n627 19.3944
R15380 gnd.n6348 gnd.n625 19.3944
R15381 gnd.n6352 gnd.n625 19.3944
R15382 gnd.n6352 gnd.n621 19.3944
R15383 gnd.n6358 gnd.n621 19.3944
R15384 gnd.n6358 gnd.n619 19.3944
R15385 gnd.n6362 gnd.n619 19.3944
R15386 gnd.n6362 gnd.n615 19.3944
R15387 gnd.n6368 gnd.n615 19.3944
R15388 gnd.n6368 gnd.n613 19.3944
R15389 gnd.n6372 gnd.n613 19.3944
R15390 gnd.n6372 gnd.n609 19.3944
R15391 gnd.n6378 gnd.n609 19.3944
R15392 gnd.n6378 gnd.n607 19.3944
R15393 gnd.n6382 gnd.n607 19.3944
R15394 gnd.n6382 gnd.n603 19.3944
R15395 gnd.n6388 gnd.n603 19.3944
R15396 gnd.n6388 gnd.n601 19.3944
R15397 gnd.n6392 gnd.n601 19.3944
R15398 gnd.n6392 gnd.n597 19.3944
R15399 gnd.n6398 gnd.n597 19.3944
R15400 gnd.n6398 gnd.n595 19.3944
R15401 gnd.n6402 gnd.n595 19.3944
R15402 gnd.n6402 gnd.n591 19.3944
R15403 gnd.n6408 gnd.n591 19.3944
R15404 gnd.n6408 gnd.n589 19.3944
R15405 gnd.n6412 gnd.n589 19.3944
R15406 gnd.n6412 gnd.n585 19.3944
R15407 gnd.n6418 gnd.n585 19.3944
R15408 gnd.n6418 gnd.n583 19.3944
R15409 gnd.n6422 gnd.n583 19.3944
R15410 gnd.n6422 gnd.n579 19.3944
R15411 gnd.n6428 gnd.n579 19.3944
R15412 gnd.n6428 gnd.n577 19.3944
R15413 gnd.n6432 gnd.n577 19.3944
R15414 gnd.n6432 gnd.n573 19.3944
R15415 gnd.n6438 gnd.n573 19.3944
R15416 gnd.n6438 gnd.n571 19.3944
R15417 gnd.n6442 gnd.n571 19.3944
R15418 gnd.n6442 gnd.n567 19.3944
R15419 gnd.n6448 gnd.n567 19.3944
R15420 gnd.n6448 gnd.n565 19.3944
R15421 gnd.n6452 gnd.n565 19.3944
R15422 gnd.n6452 gnd.n561 19.3944
R15423 gnd.n6458 gnd.n561 19.3944
R15424 gnd.n6458 gnd.n559 19.3944
R15425 gnd.n6462 gnd.n559 19.3944
R15426 gnd.n6462 gnd.n555 19.3944
R15427 gnd.n6468 gnd.n555 19.3944
R15428 gnd.n6468 gnd.n553 19.3944
R15429 gnd.n6472 gnd.n553 19.3944
R15430 gnd.n6472 gnd.n549 19.3944
R15431 gnd.n6478 gnd.n549 19.3944
R15432 gnd.n6478 gnd.n547 19.3944
R15433 gnd.n6482 gnd.n547 19.3944
R15434 gnd.n6482 gnd.n543 19.3944
R15435 gnd.n6488 gnd.n543 19.3944
R15436 gnd.n6488 gnd.n541 19.3944
R15437 gnd.n6492 gnd.n541 19.3944
R15438 gnd.n6492 gnd.n537 19.3944
R15439 gnd.n6498 gnd.n537 19.3944
R15440 gnd.n6498 gnd.n535 19.3944
R15441 gnd.n6502 gnd.n535 19.3944
R15442 gnd.n6502 gnd.n531 19.3944
R15443 gnd.n6508 gnd.n531 19.3944
R15444 gnd.n6508 gnd.n529 19.3944
R15445 gnd.n6512 gnd.n529 19.3944
R15446 gnd.n6512 gnd.n525 19.3944
R15447 gnd.n6518 gnd.n525 19.3944
R15448 gnd.n6518 gnd.n523 19.3944
R15449 gnd.n6522 gnd.n523 19.3944
R15450 gnd.n6522 gnd.n519 19.3944
R15451 gnd.n6528 gnd.n519 19.3944
R15452 gnd.n6528 gnd.n517 19.3944
R15453 gnd.n6532 gnd.n517 19.3944
R15454 gnd.n6532 gnd.n513 19.3944
R15455 gnd.n6538 gnd.n513 19.3944
R15456 gnd.n6538 gnd.n511 19.3944
R15457 gnd.n6542 gnd.n511 19.3944
R15458 gnd.n6542 gnd.n507 19.3944
R15459 gnd.n6548 gnd.n507 19.3944
R15460 gnd.n6548 gnd.n505 19.3944
R15461 gnd.n6552 gnd.n505 19.3944
R15462 gnd.n6552 gnd.n501 19.3944
R15463 gnd.n6558 gnd.n501 19.3944
R15464 gnd.n6558 gnd.n499 19.3944
R15465 gnd.n6562 gnd.n499 19.3944
R15466 gnd.n6562 gnd.n495 19.3944
R15467 gnd.n6568 gnd.n495 19.3944
R15468 gnd.n6568 gnd.n493 19.3944
R15469 gnd.n6572 gnd.n493 19.3944
R15470 gnd.n6572 gnd.n489 19.3944
R15471 gnd.n6578 gnd.n489 19.3944
R15472 gnd.n6578 gnd.n487 19.3944
R15473 gnd.n6582 gnd.n487 19.3944
R15474 gnd.n6582 gnd.n483 19.3944
R15475 gnd.n6588 gnd.n483 19.3944
R15476 gnd.n6588 gnd.n481 19.3944
R15477 gnd.n6592 gnd.n481 19.3944
R15478 gnd.n6592 gnd.n477 19.3944
R15479 gnd.n6598 gnd.n477 19.3944
R15480 gnd.n6598 gnd.n475 19.3944
R15481 gnd.n6602 gnd.n475 19.3944
R15482 gnd.n6602 gnd.n471 19.3944
R15483 gnd.n6608 gnd.n471 19.3944
R15484 gnd.n6608 gnd.n469 19.3944
R15485 gnd.n6612 gnd.n469 19.3944
R15486 gnd.n6612 gnd.n465 19.3944
R15487 gnd.n6618 gnd.n465 19.3944
R15488 gnd.n6618 gnd.n463 19.3944
R15489 gnd.n6622 gnd.n463 19.3944
R15490 gnd.n6622 gnd.n459 19.3944
R15491 gnd.n6628 gnd.n459 19.3944
R15492 gnd.n6628 gnd.n457 19.3944
R15493 gnd.n6632 gnd.n457 19.3944
R15494 gnd.n6632 gnd.n453 19.3944
R15495 gnd.n6638 gnd.n453 19.3944
R15496 gnd.n6638 gnd.n451 19.3944
R15497 gnd.n6642 gnd.n451 19.3944
R15498 gnd.n6642 gnd.n447 19.3944
R15499 gnd.n6648 gnd.n447 19.3944
R15500 gnd.n6648 gnd.n445 19.3944
R15501 gnd.n6652 gnd.n445 19.3944
R15502 gnd.n6652 gnd.n441 19.3944
R15503 gnd.n6658 gnd.n441 19.3944
R15504 gnd.n6658 gnd.n439 19.3944
R15505 gnd.n6662 gnd.n439 19.3944
R15506 gnd.n6662 gnd.n435 19.3944
R15507 gnd.n6668 gnd.n435 19.3944
R15508 gnd.n6668 gnd.n433 19.3944
R15509 gnd.n6672 gnd.n433 19.3944
R15510 gnd.n6672 gnd.n429 19.3944
R15511 gnd.n6678 gnd.n429 19.3944
R15512 gnd.n6678 gnd.n427 19.3944
R15513 gnd.n6683 gnd.n427 19.3944
R15514 gnd.n6683 gnd.n6682 19.3944
R15515 gnd.n3033 gnd.n3030 19.3944
R15516 gnd.n3033 gnd.n3028 19.3944
R15517 gnd.n3037 gnd.n3028 19.3944
R15518 gnd.n3037 gnd.n3026 19.3944
R15519 gnd.n3043 gnd.n3026 19.3944
R15520 gnd.n3043 gnd.n3024 19.3944
R15521 gnd.n3047 gnd.n3024 19.3944
R15522 gnd.n3047 gnd.n3022 19.3944
R15523 gnd.n3053 gnd.n3022 19.3944
R15524 gnd.n3053 gnd.n3020 19.3944
R15525 gnd.n3058 gnd.n3020 19.3944
R15526 gnd.n3058 gnd.n3018 19.3944
R15527 gnd.n3018 gnd.n3015 19.3944
R15528 gnd.n3065 gnd.n3015 19.3944
R15529 gnd.n3065 gnd.n3012 19.3944
R15530 gnd.n3146 gnd.n3072 19.3944
R15531 gnd.n3140 gnd.n3072 19.3944
R15532 gnd.n3140 gnd.n3139 19.3944
R15533 gnd.n3139 gnd.n3138 19.3944
R15534 gnd.n3138 gnd.n3078 19.3944
R15535 gnd.n3132 gnd.n3078 19.3944
R15536 gnd.n3132 gnd.n3131 19.3944
R15537 gnd.n3131 gnd.n3130 19.3944
R15538 gnd.n3130 gnd.n3084 19.3944
R15539 gnd.n3124 gnd.n3084 19.3944
R15540 gnd.n3124 gnd.n3123 19.3944
R15541 gnd.n3123 gnd.n3122 19.3944
R15542 gnd.n3122 gnd.n3090 19.3944
R15543 gnd.n3116 gnd.n3090 19.3944
R15544 gnd.n3116 gnd.n3115 19.3944
R15545 gnd.n3115 gnd.n3114 19.3944
R15546 gnd.n3114 gnd.n3096 19.3944
R15547 gnd.n3108 gnd.n3096 19.3944
R15548 gnd.n5568 gnd.n2804 19.3944
R15549 gnd.n5568 gnd.n2802 19.3944
R15550 gnd.n5591 gnd.n2802 19.3944
R15551 gnd.n5591 gnd.n5590 19.3944
R15552 gnd.n5590 gnd.n5589 19.3944
R15553 gnd.n5589 gnd.n5588 19.3944
R15554 gnd.n5588 gnd.n5587 19.3944
R15555 gnd.n5587 gnd.n5585 19.3944
R15556 gnd.n5585 gnd.n5584 19.3944
R15557 gnd.n5584 gnd.n5581 19.3944
R15558 gnd.n5581 gnd.n5580 19.3944
R15559 gnd.n5580 gnd.n2735 19.3944
R15560 gnd.n5680 gnd.n2735 19.3944
R15561 gnd.n5680 gnd.n2733 19.3944
R15562 gnd.n5684 gnd.n2733 19.3944
R15563 gnd.n5685 gnd.n5684 19.3944
R15564 gnd.n5688 gnd.n5685 19.3944
R15565 gnd.n5688 gnd.n2731 19.3944
R15566 gnd.n5714 gnd.n2731 19.3944
R15567 gnd.n5714 gnd.n5713 19.3944
R15568 gnd.n5713 gnd.n5712 19.3944
R15569 gnd.n5712 gnd.n5711 19.3944
R15570 gnd.n5711 gnd.n5705 19.3944
R15571 gnd.n5705 gnd.n5704 19.3944
R15572 gnd.n5704 gnd.n5703 19.3944
R15573 gnd.n5703 gnd.n5702 19.3944
R15574 gnd.n5702 gnd.n263 19.3944
R15575 gnd.n6949 gnd.n263 19.3944
R15576 gnd.n6949 gnd.n6948 19.3944
R15577 gnd.n6948 gnd.n6947 19.3944
R15578 gnd.n6947 gnd.n6944 19.3944
R15579 gnd.n6944 gnd.n6943 19.3944
R15580 gnd.n6943 gnd.n269 19.3944
R15581 gnd.n6917 gnd.n269 19.3944
R15582 gnd.n6917 gnd.n6913 19.3944
R15583 gnd.n6930 gnd.n6913 19.3944
R15584 gnd.n6930 gnd.n6929 19.3944
R15585 gnd.n6929 gnd.n6928 19.3944
R15586 gnd.n6928 gnd.n6925 19.3944
R15587 gnd.n6925 gnd.n160 19.3944
R15588 gnd.n7116 gnd.n160 19.3944
R15589 gnd.n7117 gnd.n7116 19.3944
R15590 gnd.n7155 gnd.n121 19.3944
R15591 gnd.n7150 gnd.n121 19.3944
R15592 gnd.n7150 gnd.n7149 19.3944
R15593 gnd.n7149 gnd.n7148 19.3944
R15594 gnd.n7148 gnd.n128 19.3944
R15595 gnd.n7143 gnd.n128 19.3944
R15596 gnd.n7143 gnd.n7142 19.3944
R15597 gnd.n7142 gnd.n7141 19.3944
R15598 gnd.n7141 gnd.n135 19.3944
R15599 gnd.n7136 gnd.n135 19.3944
R15600 gnd.n7136 gnd.n7135 19.3944
R15601 gnd.n7135 gnd.n7134 19.3944
R15602 gnd.n7134 gnd.n142 19.3944
R15603 gnd.n7129 gnd.n142 19.3944
R15604 gnd.n7129 gnd.n7128 19.3944
R15605 gnd.n7128 gnd.n7127 19.3944
R15606 gnd.n7127 gnd.n149 19.3944
R15607 gnd.n7122 gnd.n149 19.3944
R15608 gnd.n7188 gnd.n7187 19.3944
R15609 gnd.n7187 gnd.n7186 19.3944
R15610 gnd.n7186 gnd.n92 19.3944
R15611 gnd.n7181 gnd.n92 19.3944
R15612 gnd.n7181 gnd.n7180 19.3944
R15613 gnd.n7180 gnd.n7179 19.3944
R15614 gnd.n7179 gnd.n100 19.3944
R15615 gnd.n7174 gnd.n100 19.3944
R15616 gnd.n7174 gnd.n7173 19.3944
R15617 gnd.n7173 gnd.n7172 19.3944
R15618 gnd.n7172 gnd.n107 19.3944
R15619 gnd.n7167 gnd.n107 19.3944
R15620 gnd.n7167 gnd.n7166 19.3944
R15621 gnd.n7166 gnd.n7165 19.3944
R15622 gnd.n7165 gnd.n114 19.3944
R15623 gnd.n7160 gnd.n114 19.3944
R15624 gnd.n7160 gnd.n7159 19.3944
R15625 gnd.n5777 gnd.n5776 19.3944
R15626 gnd.n5776 gnd.n5775 19.3944
R15627 gnd.n5775 gnd.n2677 19.3944
R15628 gnd.n2792 gnd.n2677 19.3944
R15629 gnd.n2792 gnd.n2770 19.3944
R15630 gnd.n5617 gnd.n2770 19.3944
R15631 gnd.n5617 gnd.n2768 19.3944
R15632 gnd.n5623 gnd.n2768 19.3944
R15633 gnd.n5623 gnd.n5622 19.3944
R15634 gnd.n5622 gnd.n2745 19.3944
R15635 gnd.n5670 gnd.n2745 19.3944
R15636 gnd.n5670 gnd.n2743 19.3944
R15637 gnd.n5676 gnd.n2743 19.3944
R15638 gnd.n5676 gnd.n5675 19.3944
R15639 gnd.n5675 gnd.n2709 19.3944
R15640 gnd.n2709 gnd.n230 19.3944
R15641 gnd.n6983 gnd.n6982 19.3944
R15642 gnd.n5730 gnd.n5729 19.3944
R15643 gnd.n2724 gnd.n2723 19.3944
R15644 gnd.n254 gnd.n253 19.3944
R15645 gnd.n6963 gnd.n223 19.3944
R15646 gnd.n6987 gnd.n223 19.3944
R15647 gnd.n6987 gnd.n209 19.3944
R15648 gnd.n6999 gnd.n209 19.3944
R15649 gnd.n6999 gnd.n207 19.3944
R15650 gnd.n7003 gnd.n207 19.3944
R15651 gnd.n7003 gnd.n193 19.3944
R15652 gnd.n7015 gnd.n193 19.3944
R15653 gnd.n7015 gnd.n191 19.3944
R15654 gnd.n7019 gnd.n191 19.3944
R15655 gnd.n7019 gnd.n177 19.3944
R15656 gnd.n7031 gnd.n177 19.3944
R15657 gnd.n7031 gnd.n175 19.3944
R15658 gnd.n7037 gnd.n175 19.3944
R15659 gnd.n7037 gnd.n7036 19.3944
R15660 gnd.n7036 gnd.n87 19.3944
R15661 gnd.n7191 gnd.n87 19.3944
R15662 gnd.n6058 gnd.n865 19.3944
R15663 gnd.n4250 gnd.n865 19.3944
R15664 gnd.n4250 gnd.n3977 19.3944
R15665 gnd.n4254 gnd.n3977 19.3944
R15666 gnd.n4254 gnd.n3975 19.3944
R15667 gnd.n4258 gnd.n3975 19.3944
R15668 gnd.n4258 gnd.n3973 19.3944
R15669 gnd.n4262 gnd.n3973 19.3944
R15670 gnd.n4262 gnd.n3971 19.3944
R15671 gnd.n4266 gnd.n3971 19.3944
R15672 gnd.n4266 gnd.n3969 19.3944
R15673 gnd.n4275 gnd.n3969 19.3944
R15674 gnd.n4275 gnd.n4274 19.3944
R15675 gnd.n4274 gnd.n4273 19.3944
R15676 gnd.n4273 gnd.n3936 19.3944
R15677 gnd.n4361 gnd.n3936 19.3944
R15678 gnd.n4361 gnd.n3937 19.3944
R15679 gnd.n4357 gnd.n4356 19.3944
R15680 gnd.n3941 gnd.n3940 19.3944
R15681 gnd.n4324 gnd.n4323 19.3944
R15682 gnd.n4321 gnd.n4320 19.3944
R15683 gnd.n4317 gnd.n3929 19.3944
R15684 gnd.n4386 gnd.n3929 19.3944
R15685 gnd.n4386 gnd.n4385 19.3944
R15686 gnd.n4385 gnd.n4384 19.3944
R15687 gnd.n4384 gnd.n4368 19.3944
R15688 gnd.n4380 gnd.n4368 19.3944
R15689 gnd.n4380 gnd.n4379 19.3944
R15690 gnd.n4379 gnd.n4378 19.3944
R15691 gnd.n4378 gnd.n4376 19.3944
R15692 gnd.n4376 gnd.n3904 19.3944
R15693 gnd.n3904 gnd.n3902 19.3944
R15694 gnd.n4446 gnd.n3902 19.3944
R15695 gnd.n4446 gnd.n3900 19.3944
R15696 gnd.n4450 gnd.n3900 19.3944
R15697 gnd.n4450 gnd.n3898 19.3944
R15698 gnd.n4454 gnd.n3898 19.3944
R15699 gnd.n4454 gnd.n3896 19.3944
R15700 gnd.n4458 gnd.n3896 19.3944
R15701 gnd.n4458 gnd.n3894 19.3944
R15702 gnd.n4466 gnd.n3894 19.3944
R15703 gnd.n4466 gnd.n3892 19.3944
R15704 gnd.n4470 gnd.n3892 19.3944
R15705 gnd.n4470 gnd.n3756 19.3944
R15706 gnd.n4479 gnd.n3756 19.3944
R15707 gnd.n4479 gnd.n3754 19.3944
R15708 gnd.n4483 gnd.n3754 19.3944
R15709 gnd.n4483 gnd.n3750 19.3944
R15710 gnd.n4494 gnd.n3750 19.3944
R15711 gnd.n4494 gnd.n3748 19.3944
R15712 gnd.n4503 gnd.n3748 19.3944
R15713 gnd.n4503 gnd.n4502 19.3944
R15714 gnd.n4502 gnd.n4501 19.3944
R15715 gnd.n4501 gnd.n3478 19.3944
R15716 gnd.n4711 gnd.n3478 19.3944
R15717 gnd.n4711 gnd.n3476 19.3944
R15718 gnd.n4715 gnd.n3476 19.3944
R15719 gnd.n4715 gnd.n3458 19.3944
R15720 gnd.n4748 gnd.n3458 19.3944
R15721 gnd.n4748 gnd.n3456 19.3944
R15722 gnd.n4752 gnd.n3456 19.3944
R15723 gnd.n4752 gnd.n3432 19.3944
R15724 gnd.n4789 gnd.n3432 19.3944
R15725 gnd.n4789 gnd.n3430 19.3944
R15726 gnd.n4793 gnd.n3430 19.3944
R15727 gnd.n4793 gnd.n3416 19.3944
R15728 gnd.n4834 gnd.n3416 19.3944
R15729 gnd.n4834 gnd.n3414 19.3944
R15730 gnd.n4840 gnd.n3414 19.3944
R15731 gnd.n4840 gnd.n4839 19.3944
R15732 gnd.n4839 gnd.n3388 19.3944
R15733 gnd.n4906 gnd.n3388 19.3944
R15734 gnd.n4906 gnd.n3386 19.3944
R15735 gnd.n4910 gnd.n3386 19.3944
R15736 gnd.n4910 gnd.n3367 19.3944
R15737 gnd.n4933 gnd.n3367 19.3944
R15738 gnd.n4933 gnd.n3365 19.3944
R15739 gnd.n4937 gnd.n3365 19.3944
R15740 gnd.n4937 gnd.n3346 19.3944
R15741 gnd.n4966 gnd.n3346 19.3944
R15742 gnd.n4966 gnd.n3344 19.3944
R15743 gnd.n4970 gnd.n3344 19.3944
R15744 gnd.n4970 gnd.n3329 19.3944
R15745 gnd.n5011 gnd.n3329 19.3944
R15746 gnd.n5011 gnd.n3327 19.3944
R15747 gnd.n5017 gnd.n3327 19.3944
R15748 gnd.n5017 gnd.n5016 19.3944
R15749 gnd.n5016 gnd.n3300 19.3944
R15750 gnd.n5082 gnd.n3300 19.3944
R15751 gnd.n5082 gnd.n3298 19.3944
R15752 gnd.n5086 gnd.n3298 19.3944
R15753 gnd.n5086 gnd.n3280 19.3944
R15754 gnd.n5109 gnd.n3280 19.3944
R15755 gnd.n5109 gnd.n3278 19.3944
R15756 gnd.n5113 gnd.n3278 19.3944
R15757 gnd.n5113 gnd.n3258 19.3944
R15758 gnd.n5142 gnd.n3258 19.3944
R15759 gnd.n5142 gnd.n3256 19.3944
R15760 gnd.n5146 gnd.n3256 19.3944
R15761 gnd.n5146 gnd.n3241 19.3944
R15762 gnd.n5187 gnd.n3241 19.3944
R15763 gnd.n5187 gnd.n3239 19.3944
R15764 gnd.n5193 gnd.n3239 19.3944
R15765 gnd.n5193 gnd.n5192 19.3944
R15766 gnd.n5192 gnd.n3213 19.3944
R15767 gnd.n5235 gnd.n3213 19.3944
R15768 gnd.n5235 gnd.n3211 19.3944
R15769 gnd.n5239 gnd.n3211 19.3944
R15770 gnd.n5239 gnd.n3193 19.3944
R15771 gnd.n5278 gnd.n3193 19.3944
R15772 gnd.n5278 gnd.n3191 19.3944
R15773 gnd.n5284 gnd.n3191 19.3944
R15774 gnd.n5284 gnd.n5283 19.3944
R15775 gnd.n5283 gnd.n3164 19.3944
R15776 gnd.n5331 gnd.n3164 19.3944
R15777 gnd.n5331 gnd.n3162 19.3944
R15778 gnd.n5335 gnd.n3162 19.3944
R15779 gnd.n5335 gnd.n2975 19.3944
R15780 gnd.n5502 gnd.n2975 19.3944
R15781 gnd.n5502 gnd.n2973 19.3944
R15782 gnd.n5506 gnd.n2973 19.3944
R15783 gnd.n5506 gnd.n2963 19.3944
R15784 gnd.n5525 gnd.n2963 19.3944
R15785 gnd.n5525 gnd.n2961 19.3944
R15786 gnd.n5530 gnd.n2961 19.3944
R15787 gnd.n5530 gnd.n2652 19.3944
R15788 gnd.n5792 gnd.n2652 19.3944
R15789 gnd.n5792 gnd.n5791 19.3944
R15790 gnd.n5791 gnd.n5790 19.3944
R15791 gnd.n5790 gnd.n2656 19.3944
R15792 gnd.n5784 gnd.n2656 19.3944
R15793 gnd.n5784 gnd.n5783 19.3944
R15794 gnd.n5783 gnd.n5782 19.3944
R15795 gnd.n5782 gnd.n2665 19.3944
R15796 gnd.n2783 gnd.n2665 19.3944
R15797 gnd.n2787 gnd.n2783 19.3944
R15798 gnd.n2787 gnd.n2781 19.3944
R15799 gnd.n5606 gnd.n2781 19.3944
R15800 gnd.n5606 gnd.n2779 19.3944
R15801 gnd.n5612 gnd.n2779 19.3944
R15802 gnd.n5612 gnd.n5611 19.3944
R15803 gnd.n5611 gnd.n2754 19.3944
R15804 gnd.n5643 gnd.n2754 19.3944
R15805 gnd.n5643 gnd.n2752 19.3944
R15806 gnd.n5664 gnd.n2752 19.3944
R15807 gnd.n5664 gnd.n5663 19.3944
R15808 gnd.n5663 gnd.n5662 19.3944
R15809 gnd.n5662 gnd.n5649 19.3944
R15810 gnd.n5658 gnd.n5649 19.3944
R15811 gnd.n5658 gnd.n5657 19.3944
R15812 gnd.n5655 gnd.n5653 19.3944
R15813 gnd.n5720 gnd.n5719 19.3944
R15814 gnd.n5724 gnd.n5723 19.3944
R15815 gnd.n6958 gnd.n259 19.3944
R15816 gnd.n6956 gnd.n6955 19.3944
R15817 gnd.n6955 gnd.n261 19.3944
R15818 gnd.n276 gnd.n261 19.3944
R15819 gnd.n277 gnd.n276 19.3944
R15820 gnd.n280 gnd.n277 19.3944
R15821 gnd.n280 gnd.n272 19.3944
R15822 gnd.n6938 gnd.n272 19.3944
R15823 gnd.n6938 gnd.n6937 19.3944
R15824 gnd.n6937 gnd.n6936 19.3944
R15825 gnd.n6936 gnd.n286 19.3944
R15826 gnd.n6911 gnd.n286 19.3944
R15827 gnd.n6911 gnd.n6910 19.3944
R15828 gnd.n6910 gnd.n6909 19.3944
R15829 gnd.n6909 gnd.n292 19.3944
R15830 gnd.n6905 gnd.n292 19.3944
R15831 gnd.n6905 gnd.n6904 19.3944
R15832 gnd.n6904 gnd.n6903 19.3944
R15833 gnd.n4103 gnd.n4100 19.3944
R15834 gnd.n4103 gnd.n4098 19.3944
R15835 gnd.n4107 gnd.n4098 19.3944
R15836 gnd.n4107 gnd.n4096 19.3944
R15837 gnd.n4113 gnd.n4096 19.3944
R15838 gnd.n4113 gnd.n4094 19.3944
R15839 gnd.n4117 gnd.n4094 19.3944
R15840 gnd.n4117 gnd.n4092 19.3944
R15841 gnd.n4123 gnd.n4092 19.3944
R15842 gnd.n4123 gnd.n4090 19.3944
R15843 gnd.n4127 gnd.n4090 19.3944
R15844 gnd.n4127 gnd.n4088 19.3944
R15845 gnd.n4133 gnd.n4088 19.3944
R15846 gnd.n4133 gnd.n4086 19.3944
R15847 gnd.n4137 gnd.n4086 19.3944
R15848 gnd.n4137 gnd.n4081 19.3944
R15849 gnd.n4143 gnd.n4081 19.3944
R15850 gnd.n4147 gnd.n4079 19.3944
R15851 gnd.n4147 gnd.n4077 19.3944
R15852 gnd.n4153 gnd.n4077 19.3944
R15853 gnd.n4153 gnd.n4075 19.3944
R15854 gnd.n4157 gnd.n4075 19.3944
R15855 gnd.n4157 gnd.n4073 19.3944
R15856 gnd.n4163 gnd.n4073 19.3944
R15857 gnd.n4163 gnd.n4071 19.3944
R15858 gnd.n4167 gnd.n4071 19.3944
R15859 gnd.n4167 gnd.n4069 19.3944
R15860 gnd.n4173 gnd.n4069 19.3944
R15861 gnd.n4173 gnd.n4067 19.3944
R15862 gnd.n4177 gnd.n4067 19.3944
R15863 gnd.n4177 gnd.n4065 19.3944
R15864 gnd.n4183 gnd.n4065 19.3944
R15865 gnd.n4183 gnd.n4063 19.3944
R15866 gnd.n4188 gnd.n4063 19.3944
R15867 gnd.n4188 gnd.n4061 19.3944
R15868 gnd.n4001 gnd.n2335 19.3944
R15869 gnd.n6047 gnd.n2335 19.3944
R15870 gnd.n6047 gnd.n6046 19.3944
R15871 gnd.n6046 gnd.n6045 19.3944
R15872 gnd.n6045 gnd.n2339 19.3944
R15873 gnd.n6035 gnd.n2339 19.3944
R15874 gnd.n6035 gnd.n6034 19.3944
R15875 gnd.n6034 gnd.n6033 19.3944
R15876 gnd.n6033 gnd.n2361 19.3944
R15877 gnd.n6023 gnd.n2361 19.3944
R15878 gnd.n6023 gnd.n6022 19.3944
R15879 gnd.n6022 gnd.n6021 19.3944
R15880 gnd.n6021 gnd.n2383 19.3944
R15881 gnd.n6011 gnd.n2383 19.3944
R15882 gnd.n6011 gnd.n6010 19.3944
R15883 gnd.n6010 gnd.n6009 19.3944
R15884 gnd.n6009 gnd.n2404 19.3944
R15885 gnd.n5998 gnd.n2404 19.3944
R15886 gnd.n5998 gnd.n5997 19.3944
R15887 gnd.n5997 gnd.n5996 19.3944
R15888 gnd.n5996 gnd.n2424 19.3944
R15889 gnd.n5985 gnd.n2424 19.3944
R15890 gnd.n5985 gnd.n5984 19.3944
R15891 gnd.n5984 gnd.n5983 19.3944
R15892 gnd.n5983 gnd.n2440 19.3944
R15893 gnd.n5972 gnd.n2440 19.3944
R15894 gnd.n5972 gnd.n5971 19.3944
R15895 gnd.n5971 gnd.n5970 19.3944
R15896 gnd.n5970 gnd.n2459 19.3944
R15897 gnd.n5960 gnd.n2459 19.3944
R15898 gnd.n5960 gnd.n5959 19.3944
R15899 gnd.n5959 gnd.n5958 19.3944
R15900 gnd.n5958 gnd.n2479 19.3944
R15901 gnd.n5948 gnd.n2479 19.3944
R15902 gnd.n5948 gnd.n5947 19.3944
R15903 gnd.n5947 gnd.n5946 19.3944
R15904 gnd.n5946 gnd.n2501 19.3944
R15905 gnd.n5936 gnd.n2501 19.3944
R15906 gnd.n5936 gnd.n5935 19.3944
R15907 gnd.n5935 gnd.n5934 19.3944
R15908 gnd.n5934 gnd.n2522 19.3944
R15909 gnd.n5924 gnd.n2522 19.3944
R15910 gnd.n4004 gnd.n3999 19.3944
R15911 gnd.n4010 gnd.n3999 19.3944
R15912 gnd.n4010 gnd.n3997 19.3944
R15913 gnd.n4014 gnd.n3997 19.3944
R15914 gnd.n4014 gnd.n3995 19.3944
R15915 gnd.n4020 gnd.n3995 19.3944
R15916 gnd.n4020 gnd.n3993 19.3944
R15917 gnd.n4024 gnd.n3993 19.3944
R15918 gnd.n4024 gnd.n3991 19.3944
R15919 gnd.n4030 gnd.n3991 19.3944
R15920 gnd.n4030 gnd.n3989 19.3944
R15921 gnd.n4034 gnd.n3989 19.3944
R15922 gnd.n4034 gnd.n3987 19.3944
R15923 gnd.n4040 gnd.n3987 19.3944
R15924 gnd.n4040 gnd.n3985 19.3944
R15925 gnd.n4044 gnd.n3985 19.3944
R15926 gnd.n4245 gnd.n3979 19.3944
R15927 gnd.n4245 gnd.n4244 19.3944
R15928 gnd.n4244 gnd.n4243 19.3944
R15929 gnd.n4243 gnd.n4055 19.3944
R15930 gnd.n4233 gnd.n4055 19.3944
R15931 gnd.n4233 gnd.n4232 19.3944
R15932 gnd.n4232 gnd.n4231 19.3944
R15933 gnd.n4231 gnd.n4210 19.3944
R15934 gnd.n4221 gnd.n4210 19.3944
R15935 gnd.n4221 gnd.n3965 19.3944
R15936 gnd.n4280 gnd.n3965 19.3944
R15937 gnd.n4280 gnd.n3963 19.3944
R15938 gnd.n4284 gnd.n3963 19.3944
R15939 gnd.n4284 gnd.n3959 19.3944
R15940 gnd.n4297 gnd.n3959 19.3944
R15941 gnd.n4297 gnd.n3957 19.3944
R15942 gnd.n4302 gnd.n3957 19.3944
R15943 gnd.n4302 gnd.n3943 19.3944
R15944 gnd.n4350 gnd.n3943 19.3944
R15945 gnd.n4350 gnd.n4349 19.3944
R15946 gnd.n4349 gnd.n4348 19.3944
R15947 gnd.n4348 gnd.n3947 19.3944
R15948 gnd.n4344 gnd.n3947 19.3944
R15949 gnd.n4344 gnd.n4343 19.3944
R15950 gnd.n4343 gnd.n4342 19.3944
R15951 gnd.n4342 gnd.n3925 19.3944
R15952 gnd.n4391 gnd.n3925 19.3944
R15953 gnd.n4391 gnd.n3923 19.3944
R15954 gnd.n4395 gnd.n3923 19.3944
R15955 gnd.n4395 gnd.n3918 19.3944
R15956 gnd.n4407 gnd.n3918 19.3944
R15957 gnd.n4407 gnd.n3916 19.3944
R15958 gnd.n4411 gnd.n3916 19.3944
R15959 gnd.n4411 gnd.n3906 19.3944
R15960 gnd.n4439 gnd.n3906 19.3944
R15961 gnd.n4439 gnd.n3907 19.3944
R15962 gnd.n4435 gnd.n3907 19.3944
R15963 gnd.n4435 gnd.n4434 19.3944
R15964 gnd.n4434 gnd.n4433 19.3944
R15965 gnd.n4433 gnd.n3715 19.3944
R15966 gnd.n4539 gnd.n3715 19.3944
R15967 gnd.n4539 gnd.n3716 19.3944
R15968 gnd.n4199 gnd.n4198 19.3944
R15969 gnd.n4199 gnd.n4056 19.3944
R15970 gnd.n4239 gnd.n4056 19.3944
R15971 gnd.n4239 gnd.n4238 19.3944
R15972 gnd.n4238 gnd.n4237 19.3944
R15973 gnd.n4237 gnd.n4205 19.3944
R15974 gnd.n4227 gnd.n4205 19.3944
R15975 gnd.n4227 gnd.n4226 19.3944
R15976 gnd.n4226 gnd.n4225 19.3944
R15977 gnd.n4225 gnd.n4218 19.3944
R15978 gnd.n4218 gnd.n4217 19.3944
R15979 gnd.n4217 gnd.n3962 19.3944
R15980 gnd.n4288 gnd.n3962 19.3944
R15981 gnd.n4288 gnd.n3960 19.3944
R15982 gnd.n4293 gnd.n3960 19.3944
R15983 gnd.n4293 gnd.n3955 19.3944
R15984 gnd.n4306 gnd.n3955 19.3944
R15985 gnd.n4307 gnd.n4306 19.3944
R15986 gnd.n4308 gnd.n4307 19.3944
R15987 gnd.n4308 gnd.n3952 19.3944
R15988 gnd.n4314 gnd.n3952 19.3944
R15989 gnd.n4315 gnd.n4314 19.3944
R15990 gnd.n4329 gnd.n4315 19.3944
R15991 gnd.n4329 gnd.n3950 19.3944
R15992 gnd.n4337 gnd.n3950 19.3944
R15993 gnd.n4337 gnd.n4336 19.3944
R15994 gnd.n4336 gnd.n4335 19.3944
R15995 gnd.n4335 gnd.n3922 19.3944
R15996 gnd.n4399 gnd.n3922 19.3944
R15997 gnd.n4399 gnd.n3920 19.3944
R15998 gnd.n4403 gnd.n3920 19.3944
R15999 gnd.n4403 gnd.n3915 19.3944
R16000 gnd.n4415 gnd.n3915 19.3944
R16001 gnd.n4415 gnd.n3913 19.3944
R16002 gnd.n4419 gnd.n3913 19.3944
R16003 gnd.n4420 gnd.n4419 19.3944
R16004 gnd.n4423 gnd.n4420 19.3944
R16005 gnd.n4423 gnd.n3911 19.3944
R16006 gnd.n4428 gnd.n3911 19.3944
R16007 gnd.n4428 gnd.n3714 19.3944
R16008 gnd.n4543 gnd.n3714 19.3944
R16009 gnd.n4544 gnd.n4543 19.3944
R16010 gnd.n4582 gnd.n3617 19.3944
R16011 gnd.n4582 gnd.n3624 19.3944
R16012 gnd.n3681 gnd.n3624 19.3944
R16013 gnd.n4575 gnd.n3681 19.3944
R16014 gnd.n4575 gnd.n4574 19.3944
R16015 gnd.n4574 gnd.n4573 19.3944
R16016 gnd.n4573 gnd.n3687 19.3944
R16017 gnd.n4568 gnd.n3687 19.3944
R16018 gnd.n4568 gnd.n4567 19.3944
R16019 gnd.n4567 gnd.n4566 19.3944
R16020 gnd.n4566 gnd.n3694 19.3944
R16021 gnd.n4561 gnd.n3694 19.3944
R16022 gnd.n4561 gnd.n4560 19.3944
R16023 gnd.n4560 gnd.n4559 19.3944
R16024 gnd.n4559 gnd.n3701 19.3944
R16025 gnd.n4554 gnd.n3701 19.3944
R16026 gnd.n4554 gnd.n4553 19.3944
R16027 gnd.n4553 gnd.n4552 19.3944
R16028 gnd.n3637 gnd.n3636 19.3944
R16029 gnd.n3677 gnd.n3636 19.3944
R16030 gnd.n3677 gnd.n3676 19.3944
R16031 gnd.n3676 gnd.n3675 19.3944
R16032 gnd.n3675 gnd.n3672 19.3944
R16033 gnd.n3672 gnd.n3671 19.3944
R16034 gnd.n3671 gnd.n3668 19.3944
R16035 gnd.n3668 gnd.n3667 19.3944
R16036 gnd.n3667 gnd.n3664 19.3944
R16037 gnd.n3664 gnd.n3663 19.3944
R16038 gnd.n3663 gnd.n3660 19.3944
R16039 gnd.n3660 gnd.n3659 19.3944
R16040 gnd.n3659 gnd.n3656 19.3944
R16041 gnd.n3656 gnd.n3655 19.3944
R16042 gnd.n3655 gnd.n3618 19.3944
R16043 gnd.n6053 gnd.n6052 19.3944
R16044 gnd.n6052 gnd.n6051 19.3944
R16045 gnd.n6051 gnd.n2328 19.3944
R16046 gnd.n6041 gnd.n2328 19.3944
R16047 gnd.n6041 gnd.n6040 19.3944
R16048 gnd.n6040 gnd.n6039 19.3944
R16049 gnd.n6039 gnd.n2350 19.3944
R16050 gnd.n6029 gnd.n2350 19.3944
R16051 gnd.n6029 gnd.n6028 19.3944
R16052 gnd.n6028 gnd.n6027 19.3944
R16053 gnd.n6027 gnd.n2372 19.3944
R16054 gnd.n6017 gnd.n2372 19.3944
R16055 gnd.n6017 gnd.n6016 19.3944
R16056 gnd.n6016 gnd.n6015 19.3944
R16057 gnd.n6015 gnd.n2393 19.3944
R16058 gnd.n6005 gnd.n2393 19.3944
R16059 gnd.n6003 gnd.n6002 19.3944
R16060 gnd.n5992 gnd.n2430 19.3944
R16061 gnd.n5990 gnd.n5989 19.3944
R16062 gnd.n5979 gnd.n2447 19.3944
R16063 gnd.n5977 gnd.n5976 19.3944
R16064 gnd.n5976 gnd.n2448 19.3944
R16065 gnd.n5966 gnd.n2448 19.3944
R16066 gnd.n5966 gnd.n5965 19.3944
R16067 gnd.n5965 gnd.n5964 19.3944
R16068 gnd.n5964 gnd.n2469 19.3944
R16069 gnd.n5954 gnd.n2469 19.3944
R16070 gnd.n5954 gnd.n5953 19.3944
R16071 gnd.n5953 gnd.n5952 19.3944
R16072 gnd.n5952 gnd.n2490 19.3944
R16073 gnd.n5942 gnd.n2490 19.3944
R16074 gnd.n5942 gnd.n5941 19.3944
R16075 gnd.n5941 gnd.n5940 19.3944
R16076 gnd.n5940 gnd.n2511 19.3944
R16077 gnd.n5930 gnd.n2511 19.3944
R16078 gnd.n5930 gnd.n5929 19.3944
R16079 gnd.n5929 gnd.n5928 19.3944
R16080 gnd.n6229 gnd.n6228 19.3944
R16081 gnd.n6228 gnd.n698 19.3944
R16082 gnd.n6222 gnd.n698 19.3944
R16083 gnd.n6222 gnd.n6221 19.3944
R16084 gnd.n6221 gnd.n6220 19.3944
R16085 gnd.n6220 gnd.n706 19.3944
R16086 gnd.n6214 gnd.n706 19.3944
R16087 gnd.n6214 gnd.n6213 19.3944
R16088 gnd.n6213 gnd.n6212 19.3944
R16089 gnd.n6212 gnd.n714 19.3944
R16090 gnd.n6206 gnd.n714 19.3944
R16091 gnd.n6206 gnd.n6205 19.3944
R16092 gnd.n6205 gnd.n6204 19.3944
R16093 gnd.n6204 gnd.n722 19.3944
R16094 gnd.n6198 gnd.n722 19.3944
R16095 gnd.n6198 gnd.n6197 19.3944
R16096 gnd.n6197 gnd.n6196 19.3944
R16097 gnd.n6196 gnd.n730 19.3944
R16098 gnd.n6190 gnd.n730 19.3944
R16099 gnd.n6190 gnd.n6189 19.3944
R16100 gnd.n6189 gnd.n6188 19.3944
R16101 gnd.n6188 gnd.n738 19.3944
R16102 gnd.n6182 gnd.n738 19.3944
R16103 gnd.n6182 gnd.n6181 19.3944
R16104 gnd.n6181 gnd.n6180 19.3944
R16105 gnd.n6180 gnd.n746 19.3944
R16106 gnd.n6174 gnd.n746 19.3944
R16107 gnd.n6174 gnd.n6173 19.3944
R16108 gnd.n6173 gnd.n6172 19.3944
R16109 gnd.n6172 gnd.n754 19.3944
R16110 gnd.n6166 gnd.n754 19.3944
R16111 gnd.n6166 gnd.n6165 19.3944
R16112 gnd.n6165 gnd.n6164 19.3944
R16113 gnd.n6164 gnd.n762 19.3944
R16114 gnd.n6158 gnd.n762 19.3944
R16115 gnd.n6158 gnd.n6157 19.3944
R16116 gnd.n6157 gnd.n6156 19.3944
R16117 gnd.n6156 gnd.n770 19.3944
R16118 gnd.n6150 gnd.n770 19.3944
R16119 gnd.n6150 gnd.n6149 19.3944
R16120 gnd.n6149 gnd.n6148 19.3944
R16121 gnd.n6148 gnd.n778 19.3944
R16122 gnd.n6142 gnd.n778 19.3944
R16123 gnd.n6142 gnd.n6141 19.3944
R16124 gnd.n6141 gnd.n6140 19.3944
R16125 gnd.n6140 gnd.n786 19.3944
R16126 gnd.n6134 gnd.n786 19.3944
R16127 gnd.n6134 gnd.n6133 19.3944
R16128 gnd.n6133 gnd.n6132 19.3944
R16129 gnd.n6132 gnd.n794 19.3944
R16130 gnd.n6126 gnd.n794 19.3944
R16131 gnd.n6126 gnd.n6125 19.3944
R16132 gnd.n6125 gnd.n6124 19.3944
R16133 gnd.n6124 gnd.n802 19.3944
R16134 gnd.n6118 gnd.n802 19.3944
R16135 gnd.n6118 gnd.n6117 19.3944
R16136 gnd.n6117 gnd.n6116 19.3944
R16137 gnd.n6116 gnd.n810 19.3944
R16138 gnd.n6110 gnd.n810 19.3944
R16139 gnd.n6110 gnd.n6109 19.3944
R16140 gnd.n6109 gnd.n6108 19.3944
R16141 gnd.n6108 gnd.n818 19.3944
R16142 gnd.n6102 gnd.n818 19.3944
R16143 gnd.n6102 gnd.n6101 19.3944
R16144 gnd.n6101 gnd.n6100 19.3944
R16145 gnd.n6100 gnd.n826 19.3944
R16146 gnd.n6094 gnd.n826 19.3944
R16147 gnd.n6094 gnd.n6093 19.3944
R16148 gnd.n6093 gnd.n6092 19.3944
R16149 gnd.n6092 gnd.n834 19.3944
R16150 gnd.n6086 gnd.n834 19.3944
R16151 gnd.n6086 gnd.n6085 19.3944
R16152 gnd.n6085 gnd.n6084 19.3944
R16153 gnd.n6084 gnd.n842 19.3944
R16154 gnd.n6078 gnd.n842 19.3944
R16155 gnd.n6078 gnd.n6077 19.3944
R16156 gnd.n6077 gnd.n6076 19.3944
R16157 gnd.n6076 gnd.n850 19.3944
R16158 gnd.n6070 gnd.n850 19.3944
R16159 gnd.n6070 gnd.n6069 19.3944
R16160 gnd.n6069 gnd.n6068 19.3944
R16161 gnd.n6068 gnd.n858 19.3944
R16162 gnd.n6062 gnd.n858 19.3944
R16163 gnd.n6062 gnd.n6061 19.3944
R16164 gnd.n5919 gnd.n5918 19.3944
R16165 gnd.n5918 gnd.n5917 19.3944
R16166 gnd.n5917 gnd.n2546 19.3944
R16167 gnd.n5913 gnd.n2546 19.3944
R16168 gnd.n5913 gnd.n5912 19.3944
R16169 gnd.n5912 gnd.n5911 19.3944
R16170 gnd.n5911 gnd.n2551 19.3944
R16171 gnd.n5907 gnd.n2551 19.3944
R16172 gnd.n5907 gnd.n5906 19.3944
R16173 gnd.n5906 gnd.n5905 19.3944
R16174 gnd.n5905 gnd.n2556 19.3944
R16175 gnd.n5901 gnd.n2556 19.3944
R16176 gnd.n5901 gnd.n5900 19.3944
R16177 gnd.n5900 gnd.n5899 19.3944
R16178 gnd.n5899 gnd.n2561 19.3944
R16179 gnd.n5895 gnd.n2561 19.3944
R16180 gnd.n5895 gnd.n5894 19.3944
R16181 gnd.n5894 gnd.n5893 19.3944
R16182 gnd.n5893 gnd.n2566 19.3944
R16183 gnd.n5889 gnd.n2566 19.3944
R16184 gnd.n5889 gnd.n5888 19.3944
R16185 gnd.n5888 gnd.n5887 19.3944
R16186 gnd.n5887 gnd.n2571 19.3944
R16187 gnd.n5883 gnd.n2571 19.3944
R16188 gnd.n5883 gnd.n5882 19.3944
R16189 gnd.n5882 gnd.n5881 19.3944
R16190 gnd.n5881 gnd.n2576 19.3944
R16191 gnd.n5877 gnd.n2576 19.3944
R16192 gnd.n5877 gnd.n5876 19.3944
R16193 gnd.n5876 gnd.n5875 19.3944
R16194 gnd.n5875 gnd.n2581 19.3944
R16195 gnd.n5871 gnd.n2581 19.3944
R16196 gnd.n5871 gnd.n5870 19.3944
R16197 gnd.n5870 gnd.n5869 19.3944
R16198 gnd.n5869 gnd.n2586 19.3944
R16199 gnd.n5865 gnd.n2586 19.3944
R16200 gnd.n5865 gnd.n5864 19.3944
R16201 gnd.n5864 gnd.n5863 19.3944
R16202 gnd.n5863 gnd.n2591 19.3944
R16203 gnd.n5859 gnd.n2591 19.3944
R16204 gnd.n5859 gnd.n5858 19.3944
R16205 gnd.n5858 gnd.n5857 19.3944
R16206 gnd.n5857 gnd.n2596 19.3944
R16207 gnd.n5853 gnd.n2596 19.3944
R16208 gnd.n5853 gnd.n5852 19.3944
R16209 gnd.n5852 gnd.n5851 19.3944
R16210 gnd.n5851 gnd.n2601 19.3944
R16211 gnd.n5847 gnd.n2601 19.3944
R16212 gnd.n5847 gnd.n5846 19.3944
R16213 gnd.n5846 gnd.n5845 19.3944
R16214 gnd.n5845 gnd.n2606 19.3944
R16215 gnd.n5841 gnd.n2606 19.3944
R16216 gnd.n5841 gnd.n5840 19.3944
R16217 gnd.n5840 gnd.n5839 19.3944
R16218 gnd.n5839 gnd.n2611 19.3944
R16219 gnd.n5835 gnd.n2611 19.3944
R16220 gnd.n5835 gnd.n5834 19.3944
R16221 gnd.n5834 gnd.n5833 19.3944
R16222 gnd.n5833 gnd.n2616 19.3944
R16223 gnd.n5829 gnd.n2616 19.3944
R16224 gnd.n5829 gnd.n5828 19.3944
R16225 gnd.n5828 gnd.n5827 19.3944
R16226 gnd.n5827 gnd.n2621 19.3944
R16227 gnd.n5823 gnd.n2621 19.3944
R16228 gnd.n5823 gnd.n5822 19.3944
R16229 gnd.n5822 gnd.n5821 19.3944
R16230 gnd.n5821 gnd.n2626 19.3944
R16231 gnd.n5817 gnd.n2626 19.3944
R16232 gnd.n5817 gnd.n5816 19.3944
R16233 gnd.n5816 gnd.n5815 19.3944
R16234 gnd.n5815 gnd.n2631 19.3944
R16235 gnd.n5811 gnd.n2631 19.3944
R16236 gnd.n5811 gnd.n5810 19.3944
R16237 gnd.n5810 gnd.n5809 19.3944
R16238 gnd.n5809 gnd.n2636 19.3944
R16239 gnd.n5805 gnd.n2636 19.3944
R16240 gnd.n5805 gnd.n5804 19.3944
R16241 gnd.n5804 gnd.n5803 19.3944
R16242 gnd.n5803 gnd.n2641 19.3944
R16243 gnd.n5799 gnd.n2641 19.3944
R16244 gnd.n5799 gnd.n5798 19.3944
R16245 gnd.n5798 gnd.n5797 19.3944
R16246 gnd.n5548 gnd.n2956 19.3944
R16247 gnd.n5544 gnd.n2956 19.3944
R16248 gnd.n5544 gnd.n5543 19.3944
R16249 gnd.n2866 gnd.n2848 19.3944
R16250 gnd.n2866 gnd.n2846 19.3944
R16251 gnd.n2872 gnd.n2846 19.3944
R16252 gnd.n2872 gnd.n2839 19.3944
R16253 gnd.n2885 gnd.n2839 19.3944
R16254 gnd.n2885 gnd.n2837 19.3944
R16255 gnd.n2891 gnd.n2837 19.3944
R16256 gnd.n2891 gnd.n2830 19.3944
R16257 gnd.n2904 gnd.n2830 19.3944
R16258 gnd.n2904 gnd.n2828 19.3944
R16259 gnd.n2910 gnd.n2828 19.3944
R16260 gnd.n2910 gnd.n2821 19.3944
R16261 gnd.n2923 gnd.n2821 19.3944
R16262 gnd.n2923 gnd.n2819 19.3944
R16263 gnd.n2929 gnd.n2819 19.3944
R16264 gnd.n2929 gnd.n2810 19.3944
R16265 gnd.n2940 gnd.n2810 19.3944
R16266 gnd.n2940 gnd.n2808 19.3944
R16267 gnd.n5559 gnd.n2808 19.3944
R16268 gnd.n5559 gnd.n5558 19.3944
R16269 gnd.n5558 gnd.n5557 19.3944
R16270 gnd.n5557 gnd.n2948 19.3944
R16271 gnd.n5553 gnd.n2948 19.3944
R16272 gnd.n5553 gnd.n5552 19.3944
R16273 gnd.n1701 gnd.t33 18.8012
R16274 gnd.n1686 gnd.t179 18.8012
R16275 gnd.n1545 gnd.n1544 18.4825
R16276 gnd.n3147 gnd.n3012 18.4247
R16277 gnd.n4586 gnd.n3618 18.4247
R16278 gnd.n4674 gnd.n4673 18.2639
R16279 gnd.n5429 gnd.n5428 18.2639
R16280 gnd.n7084 gnd.n7083 18.2308
R16281 gnd.n2932 gnd.n2814 18.2308
R16282 gnd.n3850 gnd.n3834 18.2308
R16283 gnd.n4044 gnd.n3983 18.2308
R16284 gnd.t35 gnd.n1225 18.1639
R16285 gnd.n1253 gnd.t36 17.5266
R16286 gnd.n1652 gnd.t30 16.8893
R16287 gnd.n4541 gnd.t66 16.8893
R16288 gnd.n5566 gnd.t55 16.8893
R16289 gnd.n1831 gnd.n860 16.5706
R16290 gnd.n1480 gnd.t151 16.2519
R16291 gnd.n1180 gnd.t24 16.2519
R16292 gnd.n4463 gnd.n3890 15.9333
R16293 gnd.n4472 gnd.n3890 15.9333
R16294 gnd.n4474 gnd.n4473 15.9333
R16295 gnd.n4477 gnd.n4474 15.9333
R16296 gnd.n4477 gnd.n4476 15.9333
R16297 gnd.n4476 gnd.n4475 15.9333
R16298 gnd.n4485 gnd.n3752 15.9333
R16299 gnd.n4488 gnd.n4485 15.9333
R16300 gnd.n4489 gnd.n4488 15.9333
R16301 gnd.n4490 gnd.n4489 15.9333
R16302 gnd.n4492 gnd.n4490 15.9333
R16303 gnd.n4492 gnd.n4491 15.9333
R16304 gnd.n4491 gnd.n3745 15.9333
R16305 gnd.n4506 gnd.n3745 15.9333
R16306 gnd.n4505 gnd.n3521 15.9333
R16307 gnd.n4677 gnd.n3494 15.9333
R16308 gnd.n4660 gnd.n3496 15.9333
R16309 gnd.n4717 gnd.n3474 15.9333
R16310 gnd.n4755 gnd.n4754 15.9333
R16311 gnd.n4787 gnd.n3434 15.9333
R16312 gnd.n4832 gnd.n3418 15.9333
R16313 gnd.n4843 gnd.n4842 15.9333
R16314 gnd.n4808 gnd.n3406 15.9333
R16315 gnd.n4904 gnd.n4903 15.9333
R16316 gnd.n4912 gnd.n3384 15.9333
R16317 gnd.n4931 gnd.n4930 15.9333
R16318 gnd.n4940 gnd.n4939 15.9333
R16319 gnd.n4964 gnd.n3349 15.9333
R16320 gnd.n4972 gnd.n3342 15.9333
R16321 gnd.n5009 gnd.n3332 15.9333
R16322 gnd.n5020 gnd.n3323 15.9333
R16323 gnd.n5020 gnd.n5019 15.9333
R16324 gnd.n4986 gnd.n3319 15.9333
R16325 gnd.n5080 gnd.n5079 15.9333
R16326 gnd.n5088 gnd.n3296 15.9333
R16327 gnd.n5107 gnd.n5106 15.9333
R16328 gnd.n5116 gnd.n5115 15.9333
R16329 gnd.n5140 gnd.n3260 15.9333
R16330 gnd.n5148 gnd.n3254 15.9333
R16331 gnd.n5185 gnd.n3243 15.9333
R16332 gnd.n5196 gnd.n3235 15.9333
R16333 gnd.n5161 gnd.n3231 15.9333
R16334 gnd.n5241 gnd.n3209 15.9333
R16335 gnd.n5276 gnd.n5275 15.9333
R16336 gnd.n5288 gnd.n5286 15.9333
R16337 gnd.n5264 gnd.n3173 15.9333
R16338 gnd.n5500 gnd.n2977 15.9333
R16339 gnd.n5308 gnd.n5306 15.9333
R16340 gnd.n5508 gnd.n2971 15.9333
R16341 gnd.n5510 gnd.n5508 15.9333
R16342 gnd.n5510 gnd.n5509 15.9333
R16343 gnd.n5509 gnd.n2965 15.9333
R16344 gnd.n5523 gnd.n2965 15.9333
R16345 gnd.n5523 gnd.n5522 15.9333
R16346 gnd.n5522 gnd.n5520 15.9333
R16347 gnd.n5520 gnd.n5519 15.9333
R16348 gnd.n5533 gnd.n5532 15.9333
R16349 gnd.n5533 gnd.n2647 15.9333
R16350 gnd.n5795 gnd.n2647 15.9333
R16351 gnd.n5795 gnd.n5794 15.9333
R16352 gnd.n2658 gnd.n2649 15.9333
R16353 gnd.n5788 gnd.n2658 15.9333
R16354 gnd.n2169 gnd.n2167 15.6674
R16355 gnd.n2137 gnd.n2135 15.6674
R16356 gnd.n2105 gnd.n2103 15.6674
R16357 gnd.n2074 gnd.n2072 15.6674
R16358 gnd.n2042 gnd.n2040 15.6674
R16359 gnd.n2010 gnd.n2008 15.6674
R16360 gnd.n1978 gnd.n1976 15.6674
R16361 gnd.n1947 gnd.n1945 15.6674
R16362 gnd.n1471 gnd.t151 15.6146
R16363 gnd.t80 gnd.n948 15.6146
R16364 gnd.t70 gnd.n949 15.6146
R16365 gnd.t116 gnd.n3752 15.6146
R16366 gnd.n5519 gnd.t93 15.6146
R16367 gnd.n3466 gnd.n3460 15.296
R16368 gnd.n5296 gnd.n3182 15.296
R16369 gnd.n5346 gnd.n5345 15.0827
R16370 gnd.n3506 gnd.n3501 15.0481
R16371 gnd.n5356 gnd.n5355 15.0481
R16372 gnd.n1841 gnd.t37 14.9773
R16373 gnd.n6049 gnd.t129 14.9773
R16374 gnd.n4709 gnd.t276 14.9773
R16375 gnd.n5255 gnd.t206 14.9773
R16376 gnd.n173 gnd.t51 14.9773
R16377 gnd.n4661 gnd.n3486 14.6587
R16378 gnd.n4763 gnd.t248 14.6587
R16379 gnd.n4824 gnd.n4823 14.6587
R16380 gnd.n5163 gnd.n5162 14.6587
R16381 gnd.n3201 gnd.t208 14.6587
R16382 gnd.n5337 gnd.n3160 14.6587
R16383 gnd.t193 gnd.n991 14.34
R16384 gnd.n1919 gnd.t34 14.34
R16385 gnd.n4718 gnd.n3471 14.0214
R16386 gnd.n4786 gnd.t249 14.0214
R16387 gnd.n4913 gnd.n3381 14.0214
R16388 gnd.n4963 gnd.n3351 14.0214
R16389 gnd.n5089 gnd.n3292 14.0214
R16390 gnd.n5139 gnd.n3262 14.0214
R16391 gnd.n5242 gnd.t154 14.0214
R16392 gnd.n1627 gnd.t177 13.7027
R16393 gnd.n1337 gnd.n1336 13.5763
R16394 gnd.n2283 gnd.n905 13.5763
R16395 gnd.n3108 gnd.n3100 13.5763
R16396 gnd.n7122 gnd.n7121 13.5763
R16397 gnd.n4061 gnd.n4060 13.5763
R16398 gnd.n4552 gnd.n3710 13.5763
R16399 gnd.n1545 gnd.n1283 13.384
R16400 gnd.n4706 gnd.t97 13.384
R16401 gnd.n4780 gnd.n3440 13.384
R16402 gnd.n4816 gnd.t251 13.384
R16403 gnd.n4902 gnd.n3393 13.384
R16404 gnd.n4957 gnd.n4956 13.384
R16405 gnd.n5078 gnd.n3305 13.384
R16406 gnd.n5133 gnd.n5132 13.384
R16407 gnd.t224 gnd.n5195 13.384
R16408 gnd.n5231 gnd.n3218 13.384
R16409 gnd.n5322 gnd.t100 13.384
R16410 gnd.n5329 gnd.n5328 13.384
R16411 gnd.n3517 gnd.n3498 13.1884
R16412 gnd.n3512 gnd.n3511 13.1884
R16413 gnd.n3511 gnd.n3510 13.1884
R16414 gnd.n5349 gnd.n5344 13.1884
R16415 gnd.n5350 gnd.n5349 13.1884
R16416 gnd.n3513 gnd.n3500 13.146
R16417 gnd.n3509 gnd.n3500 13.146
R16418 gnd.n5348 gnd.n5347 13.146
R16419 gnd.n5348 gnd.n5343 13.146
R16420 gnd.n2170 gnd.n2166 12.8005
R16421 gnd.n2138 gnd.n2134 12.8005
R16422 gnd.n2106 gnd.n2102 12.8005
R16423 gnd.n2075 gnd.n2071 12.8005
R16424 gnd.n2043 gnd.n2039 12.8005
R16425 gnd.n2011 gnd.n2007 12.8005
R16426 gnd.n1979 gnd.n1975 12.8005
R16427 gnd.n1948 gnd.n1944 12.8005
R16428 gnd.n4699 gnd.n3480 12.7467
R16429 gnd.n4796 gnd.n3425 12.7467
R16430 gnd.n4895 gnd.n3390 12.7467
R16431 gnd.n4973 gnd.n3338 12.7467
R16432 gnd.n5071 gnd.n3302 12.7467
R16433 gnd.n5149 gnd.n3250 12.7467
R16434 gnd.n5224 gnd.n3215 12.7467
R16435 gnd.n1336 gnd.n1331 12.4126
R16436 gnd.n2286 gnd.n2283 12.4126
R16437 gnd.n3104 gnd.n3100 12.4126
R16438 gnd.n7121 gnd.n156 12.4126
R16439 gnd.n4195 gnd.n4060 12.4126
R16440 gnd.n4547 gnd.n3710 12.4126
R16441 gnd.n4673 gnd.n4672 12.1761
R16442 gnd.n5428 gnd.n5427 12.1761
R16443 gnd.n4733 gnd.n3449 12.1094
R16444 gnd.n3383 gnd.n3374 12.1094
R16445 gnd.n4949 gnd.n4948 12.1094
R16446 gnd.n3294 gnd.n3287 12.1094
R16447 gnd.n5125 gnd.n5124 12.1094
R16448 gnd.n3208 gnd.n3200 12.1094
R16449 gnd.n5265 gnd.n5263 12.1094
R16450 gnd.n2174 gnd.n2173 12.0247
R16451 gnd.n2142 gnd.n2141 12.0247
R16452 gnd.n2110 gnd.n2109 12.0247
R16453 gnd.n2079 gnd.n2078 12.0247
R16454 gnd.n2047 gnd.n2046 12.0247
R16455 gnd.n2015 gnd.n2014 12.0247
R16456 gnd.n1983 gnd.n1982 12.0247
R16457 gnd.n1952 gnd.n1951 12.0247
R16458 gnd.n5944 gnd.t159 11.7908
R16459 gnd.n5615 gnd.t161 11.7908
R16460 gnd.n4462 gnd.n3680 11.4721
R16461 gnd.n4831 gnd.n3421 11.4721
R16462 gnd.n4850 gnd.n4849 11.4721
R16463 gnd.n5008 gnd.n3334 11.4721
R16464 gnd.n5027 gnd.n5026 11.4721
R16465 gnd.n5184 gnd.n3245 11.4721
R16466 gnd.n5204 gnd.n5202 11.4721
R16467 gnd.t123 gnd.n3158 11.4721
R16468 gnd.n5431 gnd.n2977 11.4721
R16469 gnd.n5786 gnd.n2659 11.4721
R16470 gnd.n2177 gnd.n2164 11.249
R16471 gnd.n2145 gnd.n2132 11.249
R16472 gnd.n2113 gnd.n2100 11.249
R16473 gnd.n2082 gnd.n2069 11.249
R16474 gnd.n2050 gnd.n2037 11.249
R16475 gnd.n2018 gnd.n2005 11.249
R16476 gnd.n1986 gnd.n1973 11.249
R16477 gnd.n1955 gnd.n1942 11.249
R16478 gnd.n1615 gnd.t177 11.1535
R16479 gnd.n4277 gnd.t216 11.1535
R16480 gnd.n5968 gnd.t188 11.1535
R16481 gnd.n4506 gnd.t181 11.1535
R16482 gnd.t0 gnd.n2971 11.1535
R16483 gnd.n2740 gnd.t6 11.1535
R16484 gnd.t43 gnd.n203 11.1535
R16485 gnd.n6055 gnd.n2321 10.8348
R16486 gnd.n4248 gnd.n4247 10.8348
R16487 gnd.n6049 gnd.n2332 10.8348
R16488 gnd.n4241 gnd.n2341 10.8348
R16489 gnd.n6043 gnd.n2344 10.8348
R16490 gnd.n4235 gnd.n2352 10.8348
R16491 gnd.n6037 gnd.n2355 10.8348
R16492 gnd.n4229 gnd.n2363 10.8348
R16493 gnd.n6031 gnd.n2366 10.8348
R16494 gnd.n6025 gnd.n2377 10.8348
R16495 gnd.n4278 gnd.n4277 10.8348
R16496 gnd.n6019 gnd.n2387 10.8348
R16497 gnd.n4286 gnd.n2395 10.8348
R16498 gnd.n6013 gnd.n2398 10.8348
R16499 gnd.n4295 gnd.n2406 10.8348
R16500 gnd.n6007 gnd.n2409 10.8348
R16501 gnd.n6000 gnd.n2418 10.8348
R16502 gnd.n4353 gnd.n4352 10.8348
R16503 gnd.n5994 gnd.n2428 10.8348
R16504 gnd.n4312 gnd.n2433 10.8348
R16505 gnd.n4327 gnd.n2442 10.8348
R16506 gnd.n5981 gnd.n2445 10.8348
R16507 gnd.n4339 gnd.n2450 10.8348
R16508 gnd.n5974 gnd.n2453 10.8348
R16509 gnd.n4389 gnd.n4388 10.8348
R16510 gnd.n5968 gnd.n2463 10.8348
R16511 gnd.n4397 gnd.n2471 10.8348
R16512 gnd.n4405 gnd.n2481 10.8348
R16513 gnd.n5956 gnd.n2484 10.8348
R16514 gnd.n4413 gnd.n2492 10.8348
R16515 gnd.n5950 gnd.n2495 10.8348
R16516 gnd.n4442 gnd.n4441 10.8348
R16517 gnd.n5944 gnd.n2505 10.8348
R16518 gnd.n4421 gnd.n2513 10.8348
R16519 gnd.n5938 gnd.n2516 10.8348
R16520 gnd.n4430 gnd.n2524 10.8348
R16521 gnd.n5932 gnd.n2527 10.8348
R16522 gnd.n4541 gnd.n2534 10.8348
R16523 gnd.n5926 gnd.n2537 10.8348
R16524 gnd.t145 gnd.n3465 10.8348
R16525 gnd.n4743 gnd.n4742 10.8348
R16526 gnd.n4809 gnd.t5 10.8348
R16527 gnd.n4929 gnd.n3360 10.8348
R16528 gnd.n4941 gnd.n3360 10.8348
R16529 gnd.n5105 gnd.n3273 10.8348
R16530 gnd.n5117 gnd.n3273 10.8348
R16531 gnd.t183 gnd.n5176 10.8348
R16532 gnd.n5289 gnd.n3187 10.8348
R16533 gnd.n5780 gnd.n5779 10.8348
R16534 gnd.n5566 gnd.n2670 10.8348
R16535 gnd.n5773 gnd.n2679 10.8348
R16536 gnd.n5594 gnd.n2682 10.8348
R16537 gnd.n5593 gnd.n2794 10.8348
R16538 gnd.n5604 gnd.n5603 10.8348
R16539 gnd.n5615 gnd.n2772 10.8348
R16540 gnd.n5614 gnd.n2776 10.8348
R16541 gnd.n5625 gnd.n2763 10.8348
R16542 gnd.n5582 gnd.n2765 10.8348
R16543 gnd.n5641 gnd.n5640 10.8348
R16544 gnd.n5668 gnd.n2747 10.8348
R16545 gnd.n5678 gnd.n2738 10.8348
R16546 gnd.n2741 gnd.n2740 10.8348
R16547 gnd.n5744 gnd.n2710 10.8348
R16548 gnd.n5747 gnd.n2704 10.8348
R16549 gnd.n5686 gnd.n2707 10.8348
R16550 gnd.n6980 gnd.n233 10.8348
R16551 gnd.n5716 gnd.n236 10.8348
R16552 gnd.n5727 gnd.n2721 10.8348
R16553 gnd.n5726 gnd.n2726 10.8348
R16554 gnd.n5708 gnd.n5706 10.8348
R16555 gnd.n6961 gnd.n255 10.8348
R16556 gnd.n5700 gnd.n251 10.8348
R16557 gnd.n6989 gnd.n220 10.8348
R16558 gnd.n6952 gnd.n6951 10.8348
R16559 gnd.n6997 gnd.n211 10.8348
R16560 gnd.n6945 gnd.n214 10.8348
R16561 gnd.n7005 gnd.n203 10.8348
R16562 gnd.n6941 gnd.n205 10.8348
R16563 gnd.n6915 gnd.n197 10.8348
R16564 gnd.n7021 gnd.n188 10.8348
R16565 gnd.n6933 gnd.n6932 10.8348
R16566 gnd.n7029 gnd.n179 10.8348
R16567 gnd.n6926 gnd.n182 10.8348
R16568 gnd.n7039 gnd.n169 10.8348
R16569 gnd.n173 gnd.n171 10.8348
R16570 gnd.n7114 gnd.n162 10.8348
R16571 gnd.n7193 gnd.n81 10.8348
R16572 gnd.n5496 gnd.n5495 10.6151
R16573 gnd.n5495 gnd.n5492 10.6151
R16574 gnd.n5490 gnd.n5487 10.6151
R16575 gnd.n5487 gnd.n5486 10.6151
R16576 gnd.n5486 gnd.n5483 10.6151
R16577 gnd.n5483 gnd.n5482 10.6151
R16578 gnd.n5482 gnd.n5479 10.6151
R16579 gnd.n5479 gnd.n5478 10.6151
R16580 gnd.n5478 gnd.n5475 10.6151
R16581 gnd.n5475 gnd.n5474 10.6151
R16582 gnd.n5474 gnd.n5471 10.6151
R16583 gnd.n5471 gnd.n5470 10.6151
R16584 gnd.n5470 gnd.n5467 10.6151
R16585 gnd.n5467 gnd.n5466 10.6151
R16586 gnd.n5466 gnd.n5463 10.6151
R16587 gnd.n5463 gnd.n5462 10.6151
R16588 gnd.n5462 gnd.n5459 10.6151
R16589 gnd.n5459 gnd.n5458 10.6151
R16590 gnd.n5458 gnd.n5455 10.6151
R16591 gnd.n5455 gnd.n5454 10.6151
R16592 gnd.n5454 gnd.n5451 10.6151
R16593 gnd.n5451 gnd.n5450 10.6151
R16594 gnd.n5450 gnd.n5447 10.6151
R16595 gnd.n5447 gnd.n5446 10.6151
R16596 gnd.n5446 gnd.n5443 10.6151
R16597 gnd.n5443 gnd.n5442 10.6151
R16598 gnd.n5442 gnd.n5439 10.6151
R16599 gnd.n5439 gnd.n5438 10.6151
R16600 gnd.n5438 gnd.n5435 10.6151
R16601 gnd.n5435 gnd.n5434 10.6151
R16602 gnd.n4664 gnd.n4663 10.6151
R16603 gnd.n4663 gnd.n4659 10.6151
R16604 gnd.n4659 gnd.n4658 10.6151
R16605 gnd.n4658 gnd.n4656 10.6151
R16606 gnd.n4656 gnd.n4655 10.6151
R16607 gnd.n4655 gnd.n4652 10.6151
R16608 gnd.n4652 gnd.n3463 10.6151
R16609 gnd.n4727 gnd.n3463 10.6151
R16610 gnd.n4728 gnd.n4727 10.6151
R16611 gnd.n4740 gnd.n4728 10.6151
R16612 gnd.n4740 gnd.n4739 10.6151
R16613 gnd.n4739 gnd.n4738 10.6151
R16614 gnd.n4738 gnd.n4736 10.6151
R16615 gnd.n4736 gnd.n4735 10.6151
R16616 gnd.n4735 gnd.n4732 10.6151
R16617 gnd.n4732 gnd.n4731 10.6151
R16618 gnd.n4731 gnd.n3427 10.6151
R16619 gnd.n4798 gnd.n3427 10.6151
R16620 gnd.n4799 gnd.n4798 10.6151
R16621 gnd.n4821 gnd.n4799 10.6151
R16622 gnd.n4821 gnd.n4820 10.6151
R16623 gnd.n4820 gnd.n4819 10.6151
R16624 gnd.n4819 gnd.n4815 10.6151
R16625 gnd.n4815 gnd.n4814 10.6151
R16626 gnd.n4814 gnd.n4812 10.6151
R16627 gnd.n4812 gnd.n4811 10.6151
R16628 gnd.n4811 gnd.n4807 10.6151
R16629 gnd.n4807 gnd.n4806 10.6151
R16630 gnd.n4806 gnd.n4804 10.6151
R16631 gnd.n4804 gnd.n4803 10.6151
R16632 gnd.n4803 gnd.n4800 10.6151
R16633 gnd.n4800 gnd.n3372 10.6151
R16634 gnd.n4922 gnd.n3372 10.6151
R16635 gnd.n4923 gnd.n4922 10.6151
R16636 gnd.n4927 gnd.n4923 10.6151
R16637 gnd.n4927 gnd.n4926 10.6151
R16638 gnd.n4926 gnd.n4925 10.6151
R16639 gnd.n4925 gnd.n3355 10.6151
R16640 gnd.n4951 gnd.n3355 10.6151
R16641 gnd.n4952 gnd.n4951 10.6151
R16642 gnd.n4953 gnd.n4952 10.6151
R16643 gnd.n4953 gnd.n3340 10.6151
R16644 gnd.n4975 gnd.n3340 10.6151
R16645 gnd.n4976 gnd.n4975 10.6151
R16646 gnd.n4998 gnd.n4976 10.6151
R16647 gnd.n4998 gnd.n4997 10.6151
R16648 gnd.n4997 gnd.n4996 10.6151
R16649 gnd.n4996 gnd.n4993 10.6151
R16650 gnd.n4993 gnd.n4992 10.6151
R16651 gnd.n4992 gnd.n4990 10.6151
R16652 gnd.n4990 gnd.n4989 10.6151
R16653 gnd.n4989 gnd.n4984 10.6151
R16654 gnd.n4984 gnd.n4983 10.6151
R16655 gnd.n4983 gnd.n4981 10.6151
R16656 gnd.n4981 gnd.n4980 10.6151
R16657 gnd.n4980 gnd.n4977 10.6151
R16658 gnd.n4977 gnd.n3285 10.6151
R16659 gnd.n5098 gnd.n3285 10.6151
R16660 gnd.n5099 gnd.n5098 10.6151
R16661 gnd.n5103 gnd.n5099 10.6151
R16662 gnd.n5103 gnd.n5102 10.6151
R16663 gnd.n5102 gnd.n5101 10.6151
R16664 gnd.n5101 gnd.n3266 10.6151
R16665 gnd.n5127 gnd.n3266 10.6151
R16666 gnd.n5128 gnd.n5127 10.6151
R16667 gnd.n5129 gnd.n5128 10.6151
R16668 gnd.n5129 gnd.n3252 10.6151
R16669 gnd.n5151 gnd.n3252 10.6151
R16670 gnd.n5152 gnd.n5151 10.6151
R16671 gnd.n5174 gnd.n5152 10.6151
R16672 gnd.n5174 gnd.n5173 10.6151
R16673 gnd.n5173 gnd.n5172 10.6151
R16674 gnd.n5172 gnd.n5169 10.6151
R16675 gnd.n5169 gnd.n5168 10.6151
R16676 gnd.n5168 gnd.n5166 10.6151
R16677 gnd.n5166 gnd.n5165 10.6151
R16678 gnd.n5165 gnd.n5160 10.6151
R16679 gnd.n5160 gnd.n5159 10.6151
R16680 gnd.n5159 gnd.n5157 10.6151
R16681 gnd.n5157 gnd.n5156 10.6151
R16682 gnd.n5156 gnd.n5153 10.6151
R16683 gnd.n5153 gnd.n3198 10.6151
R16684 gnd.n5251 gnd.n3198 10.6151
R16685 gnd.n5252 gnd.n5251 10.6151
R16686 gnd.n5272 gnd.n5252 10.6151
R16687 gnd.n5272 gnd.n5271 10.6151
R16688 gnd.n5271 gnd.n5270 10.6151
R16689 gnd.n5270 gnd.n5268 10.6151
R16690 gnd.n5268 gnd.n5267 10.6151
R16691 gnd.n5267 gnd.n5262 10.6151
R16692 gnd.n5262 gnd.n5261 10.6151
R16693 gnd.n5261 gnd.n5259 10.6151
R16694 gnd.n5259 gnd.n5258 10.6151
R16695 gnd.n5258 gnd.n5254 10.6151
R16696 gnd.n5254 gnd.n5253 10.6151
R16697 gnd.n5253 gnd.n3151 10.6151
R16698 gnd.n4592 gnd.n4591 10.6151
R16699 gnd.n4595 gnd.n4592 10.6151
R16700 gnd.n4600 gnd.n4597 10.6151
R16701 gnd.n4601 gnd.n4600 10.6151
R16702 gnd.n4604 gnd.n4601 10.6151
R16703 gnd.n4605 gnd.n4604 10.6151
R16704 gnd.n4608 gnd.n4605 10.6151
R16705 gnd.n4609 gnd.n4608 10.6151
R16706 gnd.n4612 gnd.n4609 10.6151
R16707 gnd.n4613 gnd.n4612 10.6151
R16708 gnd.n4616 gnd.n4613 10.6151
R16709 gnd.n4617 gnd.n4616 10.6151
R16710 gnd.n4620 gnd.n4617 10.6151
R16711 gnd.n4621 gnd.n4620 10.6151
R16712 gnd.n4624 gnd.n4621 10.6151
R16713 gnd.n4625 gnd.n4624 10.6151
R16714 gnd.n4628 gnd.n4625 10.6151
R16715 gnd.n4629 gnd.n4628 10.6151
R16716 gnd.n4632 gnd.n4629 10.6151
R16717 gnd.n4633 gnd.n4632 10.6151
R16718 gnd.n4636 gnd.n4633 10.6151
R16719 gnd.n4637 gnd.n4636 10.6151
R16720 gnd.n4640 gnd.n4637 10.6151
R16721 gnd.n4641 gnd.n4640 10.6151
R16722 gnd.n4644 gnd.n4641 10.6151
R16723 gnd.n4645 gnd.n4644 10.6151
R16724 gnd.n4648 gnd.n4645 10.6151
R16725 gnd.n4650 gnd.n4648 10.6151
R16726 gnd.n4651 gnd.n4650 10.6151
R16727 gnd.n4665 gnd.n4651 10.6151
R16728 gnd.n4672 gnd.n4671 10.6151
R16729 gnd.n4671 gnd.n3518 10.6151
R16730 gnd.n3560 gnd.n3518 10.6151
R16731 gnd.n3561 gnd.n3560 10.6151
R16732 gnd.n3564 gnd.n3561 10.6151
R16733 gnd.n3565 gnd.n3564 10.6151
R16734 gnd.n3568 gnd.n3565 10.6151
R16735 gnd.n3569 gnd.n3568 10.6151
R16736 gnd.n3572 gnd.n3569 10.6151
R16737 gnd.n3573 gnd.n3572 10.6151
R16738 gnd.n3576 gnd.n3573 10.6151
R16739 gnd.n3577 gnd.n3576 10.6151
R16740 gnd.n3580 gnd.n3577 10.6151
R16741 gnd.n3581 gnd.n3580 10.6151
R16742 gnd.n3584 gnd.n3581 10.6151
R16743 gnd.n3585 gnd.n3584 10.6151
R16744 gnd.n3588 gnd.n3585 10.6151
R16745 gnd.n3589 gnd.n3588 10.6151
R16746 gnd.n3592 gnd.n3589 10.6151
R16747 gnd.n3593 gnd.n3592 10.6151
R16748 gnd.n3596 gnd.n3593 10.6151
R16749 gnd.n3597 gnd.n3596 10.6151
R16750 gnd.n3600 gnd.n3597 10.6151
R16751 gnd.n3601 gnd.n3600 10.6151
R16752 gnd.n3604 gnd.n3601 10.6151
R16753 gnd.n3605 gnd.n3604 10.6151
R16754 gnd.n3608 gnd.n3605 10.6151
R16755 gnd.n3609 gnd.n3608 10.6151
R16756 gnd.n3613 gnd.n3612 10.6151
R16757 gnd.n3616 gnd.n3613 10.6151
R16758 gnd.n5427 gnd.n5426 10.6151
R16759 gnd.n5426 gnd.n5423 10.6151
R16760 gnd.n5423 gnd.n5422 10.6151
R16761 gnd.n5422 gnd.n5419 10.6151
R16762 gnd.n5419 gnd.n5418 10.6151
R16763 gnd.n5418 gnd.n5415 10.6151
R16764 gnd.n5415 gnd.n5414 10.6151
R16765 gnd.n5414 gnd.n5411 10.6151
R16766 gnd.n5411 gnd.n5410 10.6151
R16767 gnd.n5410 gnd.n5407 10.6151
R16768 gnd.n5407 gnd.n5406 10.6151
R16769 gnd.n5406 gnd.n5403 10.6151
R16770 gnd.n5403 gnd.n5402 10.6151
R16771 gnd.n5402 gnd.n5399 10.6151
R16772 gnd.n5399 gnd.n5398 10.6151
R16773 gnd.n5398 gnd.n5395 10.6151
R16774 gnd.n5395 gnd.n5394 10.6151
R16775 gnd.n5394 gnd.n5391 10.6151
R16776 gnd.n5391 gnd.n5390 10.6151
R16777 gnd.n5390 gnd.n5387 10.6151
R16778 gnd.n5387 gnd.n5386 10.6151
R16779 gnd.n5386 gnd.n5383 10.6151
R16780 gnd.n5383 gnd.n5382 10.6151
R16781 gnd.n5382 gnd.n5379 10.6151
R16782 gnd.n5379 gnd.n5378 10.6151
R16783 gnd.n5378 gnd.n5375 10.6151
R16784 gnd.n5375 gnd.n5374 10.6151
R16785 gnd.n5374 gnd.n5371 10.6151
R16786 gnd.n5369 gnd.n5366 10.6151
R16787 gnd.n5366 gnd.n5365 10.6151
R16788 gnd.n4674 gnd.n3484 10.6151
R16789 gnd.n4702 gnd.n3484 10.6151
R16790 gnd.n4703 gnd.n4702 10.6151
R16791 gnd.n4704 gnd.n4703 10.6151
R16792 gnd.n4704 gnd.n3469 10.6151
R16793 gnd.n4720 gnd.n3469 10.6151
R16794 gnd.n4721 gnd.n4720 10.6151
R16795 gnd.n4723 gnd.n4721 10.6151
R16796 gnd.n4723 gnd.n4722 10.6151
R16797 gnd.n4722 gnd.n3451 10.6151
R16798 gnd.n4758 gnd.n3451 10.6151
R16799 gnd.n4759 gnd.n4758 10.6151
R16800 gnd.n4760 gnd.n4759 10.6151
R16801 gnd.n4760 gnd.n3439 10.6151
R16802 gnd.n4784 gnd.n3439 10.6151
R16803 gnd.n4784 gnd.n4783 10.6151
R16804 gnd.n4783 gnd.n4782 10.6151
R16805 gnd.n4782 gnd.n3423 10.6151
R16806 gnd.n4827 gnd.n3423 10.6151
R16807 gnd.n4828 gnd.n4827 10.6151
R16808 gnd.n4829 gnd.n4828 10.6151
R16809 gnd.n4829 gnd.n3408 10.6151
R16810 gnd.n4845 gnd.n3408 10.6151
R16811 gnd.n4846 gnd.n4845 10.6151
R16812 gnd.n4847 gnd.n4846 10.6151
R16813 gnd.n4847 gnd.n3395 10.6151
R16814 gnd.n4898 gnd.n3395 10.6151
R16815 gnd.n4899 gnd.n4898 10.6151
R16816 gnd.n4900 gnd.n4899 10.6151
R16817 gnd.n4900 gnd.n3379 10.6151
R16818 gnd.n4915 gnd.n3379 10.6151
R16819 gnd.n4916 gnd.n4915 10.6151
R16820 gnd.n4918 gnd.n4916 10.6151
R16821 gnd.n4918 gnd.n4917 10.6151
R16822 gnd.n4917 gnd.n3358 10.6151
R16823 gnd.n4943 gnd.n3358 10.6151
R16824 gnd.n4944 gnd.n4943 10.6151
R16825 gnd.n4945 gnd.n4944 10.6151
R16826 gnd.n4945 gnd.n3354 10.6151
R16827 gnd.n4961 gnd.n3354 10.6151
R16828 gnd.n4961 gnd.n4960 10.6151
R16829 gnd.n4960 gnd.n4959 10.6151
R16830 gnd.n4959 gnd.n3336 10.6151
R16831 gnd.n5004 gnd.n3336 10.6151
R16832 gnd.n5005 gnd.n5004 10.6151
R16833 gnd.n5006 gnd.n5005 10.6151
R16834 gnd.n5006 gnd.n3321 10.6151
R16835 gnd.n5022 gnd.n3321 10.6151
R16836 gnd.n5023 gnd.n5022 10.6151
R16837 gnd.n5024 gnd.n5023 10.6151
R16838 gnd.n5024 gnd.n3307 10.6151
R16839 gnd.n5074 gnd.n3307 10.6151
R16840 gnd.n5075 gnd.n5074 10.6151
R16841 gnd.n5076 gnd.n5075 10.6151
R16842 gnd.n5076 gnd.n3290 10.6151
R16843 gnd.n5091 gnd.n3290 10.6151
R16844 gnd.n5092 gnd.n5091 10.6151
R16845 gnd.n5094 gnd.n5092 10.6151
R16846 gnd.n5094 gnd.n5093 10.6151
R16847 gnd.n5093 gnd.n3271 10.6151
R16848 gnd.n5119 gnd.n3271 10.6151
R16849 gnd.n5120 gnd.n5119 10.6151
R16850 gnd.n5121 gnd.n5120 10.6151
R16851 gnd.n5121 gnd.n3265 10.6151
R16852 gnd.n5137 gnd.n3265 10.6151
R16853 gnd.n5137 gnd.n5136 10.6151
R16854 gnd.n5136 gnd.n5135 10.6151
R16855 gnd.n5135 gnd.n3247 10.6151
R16856 gnd.n5180 gnd.n3247 10.6151
R16857 gnd.n5181 gnd.n5180 10.6151
R16858 gnd.n5182 gnd.n5181 10.6151
R16859 gnd.n5182 gnd.n3233 10.6151
R16860 gnd.n5198 gnd.n3233 10.6151
R16861 gnd.n5199 gnd.n5198 10.6151
R16862 gnd.n5200 gnd.n5199 10.6151
R16863 gnd.n5200 gnd.n3220 10.6151
R16864 gnd.n5227 gnd.n3220 10.6151
R16865 gnd.n5228 gnd.n5227 10.6151
R16866 gnd.n5229 gnd.n5228 10.6151
R16867 gnd.n5229 gnd.n3204 10.6151
R16868 gnd.n5244 gnd.n3204 10.6151
R16869 gnd.n5245 gnd.n5244 10.6151
R16870 gnd.n5247 gnd.n5245 10.6151
R16871 gnd.n5247 gnd.n5246 10.6151
R16872 gnd.n5246 gnd.n3185 10.6151
R16873 gnd.n5291 gnd.n3185 10.6151
R16874 gnd.n5292 gnd.n5291 10.6151
R16875 gnd.n5293 gnd.n5292 10.6151
R16876 gnd.n5293 gnd.n3171 10.6151
R16877 gnd.n5324 gnd.n3171 10.6151
R16878 gnd.n5325 gnd.n5324 10.6151
R16879 gnd.n5326 gnd.n5325 10.6151
R16880 gnd.n5326 gnd.n3156 10.6151
R16881 gnd.n5340 gnd.n3156 10.6151
R16882 gnd.n5341 gnd.n5340 10.6151
R16883 gnd.n5429 gnd.n5341 10.6151
R16884 gnd.n1534 gnd.t278 10.5161
R16885 gnd.n993 gnd.t193 10.5161
R16886 gnd.n1902 gnd.t34 10.5161
R16887 gnd.t20 gnd.n2415 10.5161
R16888 gnd.n4353 gnd.t38 10.5161
R16889 gnd.n5994 gnd.t38 10.5161
R16890 gnd.n5987 gnd.t220 10.5161
R16891 gnd.n5732 gnd.t259 10.5161
R16892 gnd.t3 gnd.n2726 10.5161
R16893 gnd.n5706 gnd.t3 10.5161
R16894 gnd.n6960 gnd.t209 10.5161
R16895 gnd.n2178 gnd.n2162 10.4732
R16896 gnd.n2146 gnd.n2130 10.4732
R16897 gnd.n2114 gnd.n2098 10.4732
R16898 gnd.n2083 gnd.n2067 10.4732
R16899 gnd.n2051 gnd.n2035 10.4732
R16900 gnd.n2019 gnd.n2003 10.4732
R16901 gnd.n1987 gnd.n1971 10.4732
R16902 gnd.n1956 gnd.n1940 10.4732
R16903 gnd.n4746 gnd.t84 10.1975
R16904 gnd.n4817 gnd.n3421 10.1975
R16905 gnd.n4994 gnd.n3334 10.1975
R16906 gnd.n5027 gnd.n3317 10.1975
R16907 gnd.n5204 gnd.n3229 10.1975
R16908 gnd.t37 gnd.n1010 9.87883
R16909 gnd.t18 gnd.n2374 9.87883
R16910 gnd.n6019 gnd.t216 9.87883
R16911 gnd.n4388 gnd.t188 9.87883
R16912 gnd.n5962 gnd.t41 9.87883
R16913 gnd.n4668 gnd.n3494 9.87883
R16914 gnd.n5500 gnd.n5499 9.87883
R16915 gnd.n5631 gnd.t8 9.87883
R16916 gnd.t6 gnd.n2710 9.87883
R16917 gnd.n6945 gnd.t43 9.87883
R16918 gnd.n6940 gnd.t157 9.87883
R16919 gnd.n2182 gnd.n2181 9.69747
R16920 gnd.n2150 gnd.n2149 9.69747
R16921 gnd.n2118 gnd.n2117 9.69747
R16922 gnd.n2087 gnd.n2086 9.69747
R16923 gnd.n2055 gnd.n2054 9.69747
R16924 gnd.n2023 gnd.n2022 9.69747
R16925 gnd.n1991 gnd.n1990 9.69747
R16926 gnd.n1960 gnd.n1959 9.69747
R16927 gnd.n7228 gnd.n50 9.6512
R16928 gnd.n4725 gnd.n3465 9.56018
R16929 gnd.n4762 gnd.n3449 9.56018
R16930 gnd.n4920 gnd.n3374 9.56018
R16931 gnd.n3376 gnd.t232 9.56018
R16932 gnd.n4948 gnd.n4947 9.56018
R16933 gnd.n5096 gnd.n3287 9.56018
R16934 gnd.t231 gnd.n3269 9.56018
R16935 gnd.n5124 gnd.n5123 9.56018
R16936 gnd.n5249 gnd.n3200 9.56018
R16937 gnd.n5303 gnd.t74 9.56018
R16938 gnd.n5922 gnd.n2540 9.45599
R16939 gnd.n2856 gnd.n2855 9.45599
R16940 gnd.n2188 gnd.n2187 9.45567
R16941 gnd.n2156 gnd.n2155 9.45567
R16942 gnd.n2124 gnd.n2123 9.45567
R16943 gnd.n2093 gnd.n2092 9.45567
R16944 gnd.n2061 gnd.n2060 9.45567
R16945 gnd.n2029 gnd.n2028 9.45567
R16946 gnd.n1997 gnd.n1996 9.45567
R16947 gnd.n1966 gnd.n1965 9.45567
R16948 gnd.n1132 gnd.n1131 9.39724
R16949 gnd.n2187 gnd.n2186 9.3005
R16950 gnd.n2160 gnd.n2159 9.3005
R16951 gnd.n2181 gnd.n2180 9.3005
R16952 gnd.n2179 gnd.n2178 9.3005
R16953 gnd.n2164 gnd.n2163 9.3005
R16954 gnd.n2173 gnd.n2172 9.3005
R16955 gnd.n2171 gnd.n2170 9.3005
R16956 gnd.n2155 gnd.n2154 9.3005
R16957 gnd.n2128 gnd.n2127 9.3005
R16958 gnd.n2149 gnd.n2148 9.3005
R16959 gnd.n2147 gnd.n2146 9.3005
R16960 gnd.n2132 gnd.n2131 9.3005
R16961 gnd.n2141 gnd.n2140 9.3005
R16962 gnd.n2139 gnd.n2138 9.3005
R16963 gnd.n2123 gnd.n2122 9.3005
R16964 gnd.n2096 gnd.n2095 9.3005
R16965 gnd.n2117 gnd.n2116 9.3005
R16966 gnd.n2115 gnd.n2114 9.3005
R16967 gnd.n2100 gnd.n2099 9.3005
R16968 gnd.n2109 gnd.n2108 9.3005
R16969 gnd.n2107 gnd.n2106 9.3005
R16970 gnd.n2092 gnd.n2091 9.3005
R16971 gnd.n2065 gnd.n2064 9.3005
R16972 gnd.n2086 gnd.n2085 9.3005
R16973 gnd.n2084 gnd.n2083 9.3005
R16974 gnd.n2069 gnd.n2068 9.3005
R16975 gnd.n2078 gnd.n2077 9.3005
R16976 gnd.n2076 gnd.n2075 9.3005
R16977 gnd.n2060 gnd.n2059 9.3005
R16978 gnd.n2033 gnd.n2032 9.3005
R16979 gnd.n2054 gnd.n2053 9.3005
R16980 gnd.n2052 gnd.n2051 9.3005
R16981 gnd.n2037 gnd.n2036 9.3005
R16982 gnd.n2046 gnd.n2045 9.3005
R16983 gnd.n2044 gnd.n2043 9.3005
R16984 gnd.n2028 gnd.n2027 9.3005
R16985 gnd.n2001 gnd.n2000 9.3005
R16986 gnd.n2022 gnd.n2021 9.3005
R16987 gnd.n2020 gnd.n2019 9.3005
R16988 gnd.n2005 gnd.n2004 9.3005
R16989 gnd.n2014 gnd.n2013 9.3005
R16990 gnd.n2012 gnd.n2011 9.3005
R16991 gnd.n1996 gnd.n1995 9.3005
R16992 gnd.n1969 gnd.n1968 9.3005
R16993 gnd.n1990 gnd.n1989 9.3005
R16994 gnd.n1988 gnd.n1987 9.3005
R16995 gnd.n1973 gnd.n1972 9.3005
R16996 gnd.n1982 gnd.n1981 9.3005
R16997 gnd.n1980 gnd.n1979 9.3005
R16998 gnd.n1965 gnd.n1964 9.3005
R16999 gnd.n1938 gnd.n1937 9.3005
R17000 gnd.n1959 gnd.n1958 9.3005
R17001 gnd.n1957 gnd.n1956 9.3005
R17002 gnd.n1942 gnd.n1941 9.3005
R17003 gnd.n1951 gnd.n1950 9.3005
R17004 gnd.n1949 gnd.n1948 9.3005
R17005 gnd.n2313 gnd.n2312 9.3005
R17006 gnd.n2311 gnd.n893 9.3005
R17007 gnd.n2310 gnd.n2309 9.3005
R17008 gnd.n2306 gnd.n894 9.3005
R17009 gnd.n2303 gnd.n895 9.3005
R17010 gnd.n2302 gnd.n896 9.3005
R17011 gnd.n2299 gnd.n897 9.3005
R17012 gnd.n2298 gnd.n898 9.3005
R17013 gnd.n2295 gnd.n899 9.3005
R17014 gnd.n2294 gnd.n900 9.3005
R17015 gnd.n2291 gnd.n901 9.3005
R17016 gnd.n2290 gnd.n902 9.3005
R17017 gnd.n2287 gnd.n903 9.3005
R17018 gnd.n2286 gnd.n904 9.3005
R17019 gnd.n2283 gnd.n2282 9.3005
R17020 gnd.n2281 gnd.n905 9.3005
R17021 gnd.n2314 gnd.n892 9.3005
R17022 gnd.n1553 gnd.n1552 9.3005
R17023 gnd.n1257 gnd.n1256 9.3005
R17024 gnd.n1580 gnd.n1579 9.3005
R17025 gnd.n1581 gnd.n1255 9.3005
R17026 gnd.n1585 gnd.n1582 9.3005
R17027 gnd.n1584 gnd.n1583 9.3005
R17028 gnd.n1229 gnd.n1228 9.3005
R17029 gnd.n1610 gnd.n1609 9.3005
R17030 gnd.n1611 gnd.n1227 9.3005
R17031 gnd.n1613 gnd.n1612 9.3005
R17032 gnd.n1207 gnd.n1206 9.3005
R17033 gnd.n1641 gnd.n1640 9.3005
R17034 gnd.n1642 gnd.n1205 9.3005
R17035 gnd.n1650 gnd.n1643 9.3005
R17036 gnd.n1649 gnd.n1644 9.3005
R17037 gnd.n1648 gnd.n1646 9.3005
R17038 gnd.n1645 gnd.n1154 9.3005
R17039 gnd.n1698 gnd.n1155 9.3005
R17040 gnd.n1697 gnd.n1156 9.3005
R17041 gnd.n1696 gnd.n1157 9.3005
R17042 gnd.n1176 gnd.n1158 9.3005
R17043 gnd.n1178 gnd.n1177 9.3005
R17044 gnd.n1088 gnd.n1087 9.3005
R17045 gnd.n1736 gnd.n1735 9.3005
R17046 gnd.n1737 gnd.n1086 9.3005
R17047 gnd.n1741 gnd.n1738 9.3005
R17048 gnd.n1740 gnd.n1739 9.3005
R17049 gnd.n1061 gnd.n1060 9.3005
R17050 gnd.n1776 gnd.n1775 9.3005
R17051 gnd.n1777 gnd.n1059 9.3005
R17052 gnd.n1781 gnd.n1778 9.3005
R17053 gnd.n1780 gnd.n1779 9.3005
R17054 gnd.n1035 gnd.n1034 9.3005
R17055 gnd.n1823 gnd.n1822 9.3005
R17056 gnd.n1824 gnd.n1033 9.3005
R17057 gnd.n1828 gnd.n1825 9.3005
R17058 gnd.n1827 gnd.n1826 9.3005
R17059 gnd.n1008 gnd.n1007 9.3005
R17060 gnd.n1863 gnd.n1862 9.3005
R17061 gnd.n1864 gnd.n1006 9.3005
R17062 gnd.n1868 gnd.n1865 9.3005
R17063 gnd.n1867 gnd.n1866 9.3005
R17064 gnd.n981 gnd.n980 9.3005
R17065 gnd.n1912 gnd.n1911 9.3005
R17066 gnd.n1913 gnd.n979 9.3005
R17067 gnd.n1917 gnd.n1914 9.3005
R17068 gnd.n1916 gnd.n1915 9.3005
R17069 gnd.n954 gnd.n953 9.3005
R17070 gnd.n2206 gnd.n2205 9.3005
R17071 gnd.n2207 gnd.n952 9.3005
R17072 gnd.n2213 gnd.n2208 9.3005
R17073 gnd.n2212 gnd.n2209 9.3005
R17074 gnd.n2211 gnd.n2210 9.3005
R17075 gnd.n1554 gnd.n1551 9.3005
R17076 gnd.n1336 gnd.n1295 9.3005
R17077 gnd.n1331 gnd.n1330 9.3005
R17078 gnd.n1329 gnd.n1296 9.3005
R17079 gnd.n1328 gnd.n1327 9.3005
R17080 gnd.n1324 gnd.n1297 9.3005
R17081 gnd.n1321 gnd.n1320 9.3005
R17082 gnd.n1319 gnd.n1298 9.3005
R17083 gnd.n1318 gnd.n1317 9.3005
R17084 gnd.n1314 gnd.n1299 9.3005
R17085 gnd.n1311 gnd.n1310 9.3005
R17086 gnd.n1309 gnd.n1300 9.3005
R17087 gnd.n1308 gnd.n1307 9.3005
R17088 gnd.n1304 gnd.n1302 9.3005
R17089 gnd.n1301 gnd.n1281 9.3005
R17090 gnd.n1548 gnd.n1280 9.3005
R17091 gnd.n1550 gnd.n1549 9.3005
R17092 gnd.n1338 gnd.n1337 9.3005
R17093 gnd.n1561 gnd.n1267 9.3005
R17094 gnd.n1568 gnd.n1268 9.3005
R17095 gnd.n1570 gnd.n1569 9.3005
R17096 gnd.n1571 gnd.n1248 9.3005
R17097 gnd.n1590 gnd.n1589 9.3005
R17098 gnd.n1592 gnd.n1240 9.3005
R17099 gnd.n1599 gnd.n1242 9.3005
R17100 gnd.n1600 gnd.n1237 9.3005
R17101 gnd.n1602 gnd.n1601 9.3005
R17102 gnd.n1238 gnd.n1223 9.3005
R17103 gnd.n1618 gnd.n1221 9.3005
R17104 gnd.n1622 gnd.n1621 9.3005
R17105 gnd.n1620 gnd.n1197 9.3005
R17106 gnd.n1657 gnd.n1196 9.3005
R17107 gnd.n1660 gnd.n1659 9.3005
R17108 gnd.n1193 gnd.n1192 9.3005
R17109 gnd.n1666 gnd.n1194 9.3005
R17110 gnd.n1668 gnd.n1667 9.3005
R17111 gnd.n1670 gnd.n1191 9.3005
R17112 gnd.n1673 gnd.n1672 9.3005
R17113 gnd.n1676 gnd.n1674 9.3005
R17114 gnd.n1678 gnd.n1677 9.3005
R17115 gnd.n1684 gnd.n1679 9.3005
R17116 gnd.n1683 gnd.n1682 9.3005
R17117 gnd.n1079 gnd.n1078 9.3005
R17118 gnd.n1750 gnd.n1749 9.3005
R17119 gnd.n1751 gnd.n1072 9.3005
R17120 gnd.n1759 gnd.n1071 9.3005
R17121 gnd.n1762 gnd.n1761 9.3005
R17122 gnd.n1764 gnd.n1763 9.3005
R17123 gnd.n1767 gnd.n1054 9.3005
R17124 gnd.n1765 gnd.n1052 9.3005
R17125 gnd.n1787 gnd.n1050 9.3005
R17126 gnd.n1789 gnd.n1788 9.3005
R17127 gnd.n1026 gnd.n1025 9.3005
R17128 gnd.n1837 gnd.n1836 9.3005
R17129 gnd.n1838 gnd.n1019 9.3005
R17130 gnd.n1846 gnd.n1018 9.3005
R17131 gnd.n1849 gnd.n1848 9.3005
R17132 gnd.n1851 gnd.n1850 9.3005
R17133 gnd.n1854 gnd.n1001 9.3005
R17134 gnd.n1852 gnd.n999 9.3005
R17135 gnd.n1874 gnd.n997 9.3005
R17136 gnd.n1876 gnd.n1875 9.3005
R17137 gnd.n972 gnd.n971 9.3005
R17138 gnd.n1926 gnd.n1925 9.3005
R17139 gnd.n1927 gnd.n965 9.3005
R17140 gnd.n1935 gnd.n964 9.3005
R17141 gnd.n2194 gnd.n2193 9.3005
R17142 gnd.n2196 gnd.n2195 9.3005
R17143 gnd.n2197 gnd.n945 9.3005
R17144 gnd.n2221 gnd.n2220 9.3005
R17145 gnd.n946 gnd.n908 9.3005
R17146 gnd.n1559 gnd.n1558 9.3005
R17147 gnd.n2277 gnd.n909 9.3005
R17148 gnd.n2276 gnd.n911 9.3005
R17149 gnd.n2273 gnd.n912 9.3005
R17150 gnd.n2272 gnd.n913 9.3005
R17151 gnd.n2269 gnd.n914 9.3005
R17152 gnd.n2268 gnd.n915 9.3005
R17153 gnd.n2265 gnd.n916 9.3005
R17154 gnd.n2264 gnd.n917 9.3005
R17155 gnd.n2261 gnd.n918 9.3005
R17156 gnd.n2260 gnd.n919 9.3005
R17157 gnd.n2257 gnd.n920 9.3005
R17158 gnd.n2256 gnd.n921 9.3005
R17159 gnd.n2253 gnd.n922 9.3005
R17160 gnd.n2252 gnd.n923 9.3005
R17161 gnd.n2249 gnd.n924 9.3005
R17162 gnd.n2248 gnd.n925 9.3005
R17163 gnd.n2245 gnd.n926 9.3005
R17164 gnd.n2244 gnd.n927 9.3005
R17165 gnd.n2241 gnd.n928 9.3005
R17166 gnd.n2240 gnd.n929 9.3005
R17167 gnd.n2237 gnd.n930 9.3005
R17168 gnd.n2236 gnd.n931 9.3005
R17169 gnd.n2233 gnd.n935 9.3005
R17170 gnd.n2232 gnd.n936 9.3005
R17171 gnd.n2229 gnd.n937 9.3005
R17172 gnd.n2228 gnd.n938 9.3005
R17173 gnd.n2279 gnd.n2278 9.3005
R17174 gnd.n1728 gnd.n1712 9.3005
R17175 gnd.n1727 gnd.n1713 9.3005
R17176 gnd.n1726 gnd.n1714 9.3005
R17177 gnd.n1724 gnd.n1715 9.3005
R17178 gnd.n1723 gnd.n1716 9.3005
R17179 gnd.n1721 gnd.n1717 9.3005
R17180 gnd.n1720 gnd.n1718 9.3005
R17181 gnd.n1042 gnd.n1041 9.3005
R17182 gnd.n1797 gnd.n1796 9.3005
R17183 gnd.n1798 gnd.n1040 9.3005
R17184 gnd.n1815 gnd.n1799 9.3005
R17185 gnd.n1814 gnd.n1800 9.3005
R17186 gnd.n1813 gnd.n1801 9.3005
R17187 gnd.n1811 gnd.n1802 9.3005
R17188 gnd.n1810 gnd.n1803 9.3005
R17189 gnd.n1808 gnd.n1804 9.3005
R17190 gnd.n1807 gnd.n1805 9.3005
R17191 gnd.n988 gnd.n987 9.3005
R17192 gnd.n1884 gnd.n1883 9.3005
R17193 gnd.n1885 gnd.n986 9.3005
R17194 gnd.n1906 gnd.n1886 9.3005
R17195 gnd.n1905 gnd.n1887 9.3005
R17196 gnd.n1904 gnd.n1888 9.3005
R17197 gnd.n1901 gnd.n1889 9.3005
R17198 gnd.n1900 gnd.n1890 9.3005
R17199 gnd.n1898 gnd.n1891 9.3005
R17200 gnd.n1897 gnd.n1892 9.3005
R17201 gnd.n1895 gnd.n1894 9.3005
R17202 gnd.n1893 gnd.n940 9.3005
R17203 gnd.n1469 gnd.n1468 9.3005
R17204 gnd.n1359 gnd.n1358 9.3005
R17205 gnd.n1483 gnd.n1482 9.3005
R17206 gnd.n1484 gnd.n1357 9.3005
R17207 gnd.n1486 gnd.n1485 9.3005
R17208 gnd.n1347 gnd.n1346 9.3005
R17209 gnd.n1499 gnd.n1498 9.3005
R17210 gnd.n1500 gnd.n1345 9.3005
R17211 gnd.n1532 gnd.n1501 9.3005
R17212 gnd.n1531 gnd.n1502 9.3005
R17213 gnd.n1530 gnd.n1503 9.3005
R17214 gnd.n1529 gnd.n1504 9.3005
R17215 gnd.n1526 gnd.n1505 9.3005
R17216 gnd.n1525 gnd.n1506 9.3005
R17217 gnd.n1524 gnd.n1507 9.3005
R17218 gnd.n1522 gnd.n1508 9.3005
R17219 gnd.n1521 gnd.n1509 9.3005
R17220 gnd.n1518 gnd.n1510 9.3005
R17221 gnd.n1517 gnd.n1511 9.3005
R17222 gnd.n1516 gnd.n1512 9.3005
R17223 gnd.n1514 gnd.n1513 9.3005
R17224 gnd.n1213 gnd.n1212 9.3005
R17225 gnd.n1630 gnd.n1629 9.3005
R17226 gnd.n1631 gnd.n1211 9.3005
R17227 gnd.n1635 gnd.n1632 9.3005
R17228 gnd.n1634 gnd.n1633 9.3005
R17229 gnd.n1135 gnd.n1134 9.3005
R17230 gnd.n1710 gnd.n1709 9.3005
R17231 gnd.n1467 gnd.n1368 9.3005
R17232 gnd.n1370 gnd.n1369 9.3005
R17233 gnd.n1414 gnd.n1412 9.3005
R17234 gnd.n1415 gnd.n1411 9.3005
R17235 gnd.n1418 gnd.n1407 9.3005
R17236 gnd.n1419 gnd.n1406 9.3005
R17237 gnd.n1422 gnd.n1405 9.3005
R17238 gnd.n1423 gnd.n1404 9.3005
R17239 gnd.n1426 gnd.n1403 9.3005
R17240 gnd.n1427 gnd.n1402 9.3005
R17241 gnd.n1430 gnd.n1401 9.3005
R17242 gnd.n1431 gnd.n1400 9.3005
R17243 gnd.n1434 gnd.n1399 9.3005
R17244 gnd.n1435 gnd.n1398 9.3005
R17245 gnd.n1438 gnd.n1397 9.3005
R17246 gnd.n1439 gnd.n1396 9.3005
R17247 gnd.n1442 gnd.n1395 9.3005
R17248 gnd.n1443 gnd.n1394 9.3005
R17249 gnd.n1446 gnd.n1393 9.3005
R17250 gnd.n1447 gnd.n1392 9.3005
R17251 gnd.n1450 gnd.n1391 9.3005
R17252 gnd.n1451 gnd.n1390 9.3005
R17253 gnd.n1454 gnd.n1389 9.3005
R17254 gnd.n1456 gnd.n1388 9.3005
R17255 gnd.n1457 gnd.n1387 9.3005
R17256 gnd.n1458 gnd.n1386 9.3005
R17257 gnd.n1459 gnd.n1385 9.3005
R17258 gnd.n1466 gnd.n1465 9.3005
R17259 gnd.n1475 gnd.n1474 9.3005
R17260 gnd.n1476 gnd.n1362 9.3005
R17261 gnd.n1478 gnd.n1477 9.3005
R17262 gnd.n1353 gnd.n1352 9.3005
R17263 gnd.n1491 gnd.n1490 9.3005
R17264 gnd.n1492 gnd.n1351 9.3005
R17265 gnd.n1494 gnd.n1493 9.3005
R17266 gnd.n1340 gnd.n1339 9.3005
R17267 gnd.n1537 gnd.n1536 9.3005
R17268 gnd.n1538 gnd.n1294 9.3005
R17269 gnd.n1542 gnd.n1540 9.3005
R17270 gnd.n1541 gnd.n1273 9.3005
R17271 gnd.n1560 gnd.n1272 9.3005
R17272 gnd.n1563 gnd.n1562 9.3005
R17273 gnd.n1266 gnd.n1265 9.3005
R17274 gnd.n1574 gnd.n1572 9.3005
R17275 gnd.n1573 gnd.n1247 9.3005
R17276 gnd.n1591 gnd.n1246 9.3005
R17277 gnd.n1594 gnd.n1593 9.3005
R17278 gnd.n1241 gnd.n1236 9.3005
R17279 gnd.n1604 gnd.n1603 9.3005
R17280 gnd.n1239 gnd.n1219 9.3005
R17281 gnd.n1625 gnd.n1220 9.3005
R17282 gnd.n1624 gnd.n1623 9.3005
R17283 gnd.n1222 gnd.n1198 9.3005
R17284 gnd.n1656 gnd.n1655 9.3005
R17285 gnd.n1658 gnd.n1143 9.3005
R17286 gnd.n1705 gnd.n1144 9.3005
R17287 gnd.n1704 gnd.n1145 9.3005
R17288 gnd.n1703 gnd.n1146 9.3005
R17289 gnd.n1669 gnd.n1147 9.3005
R17290 gnd.n1671 gnd.n1165 9.3005
R17291 gnd.n1691 gnd.n1166 9.3005
R17292 gnd.n1690 gnd.n1167 9.3005
R17293 gnd.n1689 gnd.n1168 9.3005
R17294 gnd.n1680 gnd.n1169 9.3005
R17295 gnd.n1681 gnd.n1080 9.3005
R17296 gnd.n1747 gnd.n1746 9.3005
R17297 gnd.n1748 gnd.n1073 9.3005
R17298 gnd.n1758 gnd.n1757 9.3005
R17299 gnd.n1760 gnd.n1069 9.3005
R17300 gnd.n1770 gnd.n1070 9.3005
R17301 gnd.n1769 gnd.n1768 9.3005
R17302 gnd.n1766 gnd.n1048 9.3005
R17303 gnd.n1792 gnd.n1049 9.3005
R17304 gnd.n1791 gnd.n1790 9.3005
R17305 gnd.n1051 gnd.n1027 9.3005
R17306 gnd.n1834 gnd.n1833 9.3005
R17307 gnd.n1835 gnd.n1020 9.3005
R17308 gnd.n1845 gnd.n1844 9.3005
R17309 gnd.n1847 gnd.n1016 9.3005
R17310 gnd.n1857 gnd.n1017 9.3005
R17311 gnd.n1856 gnd.n1855 9.3005
R17312 gnd.n1853 gnd.n995 9.3005
R17313 gnd.n1879 gnd.n996 9.3005
R17314 gnd.n1878 gnd.n1877 9.3005
R17315 gnd.n998 gnd.n973 9.3005
R17316 gnd.n1923 gnd.n1922 9.3005
R17317 gnd.n1924 gnd.n966 9.3005
R17318 gnd.n1934 gnd.n1933 9.3005
R17319 gnd.n2192 gnd.n962 9.3005
R17320 gnd.n2200 gnd.n963 9.3005
R17321 gnd.n2199 gnd.n2198 9.3005
R17322 gnd.n944 gnd.n943 9.3005
R17323 gnd.n2223 gnd.n2222 9.3005
R17324 gnd.n1364 gnd.n1363 9.3005
R17325 gnd.n6232 gnd.n6231 9.3005
R17326 gnd.n693 gnd.n692 9.3005
R17327 gnd.n6239 gnd.n6238 9.3005
R17328 gnd.n6240 gnd.n691 9.3005
R17329 gnd.n6242 gnd.n6241 9.3005
R17330 gnd.n687 gnd.n686 9.3005
R17331 gnd.n6249 gnd.n6248 9.3005
R17332 gnd.n6250 gnd.n685 9.3005
R17333 gnd.n6252 gnd.n6251 9.3005
R17334 gnd.n681 gnd.n680 9.3005
R17335 gnd.n6259 gnd.n6258 9.3005
R17336 gnd.n6260 gnd.n679 9.3005
R17337 gnd.n6262 gnd.n6261 9.3005
R17338 gnd.n675 gnd.n674 9.3005
R17339 gnd.n6269 gnd.n6268 9.3005
R17340 gnd.n6270 gnd.n673 9.3005
R17341 gnd.n6272 gnd.n6271 9.3005
R17342 gnd.n669 gnd.n668 9.3005
R17343 gnd.n6279 gnd.n6278 9.3005
R17344 gnd.n6280 gnd.n667 9.3005
R17345 gnd.n6282 gnd.n6281 9.3005
R17346 gnd.n663 gnd.n662 9.3005
R17347 gnd.n6289 gnd.n6288 9.3005
R17348 gnd.n6290 gnd.n661 9.3005
R17349 gnd.n6292 gnd.n6291 9.3005
R17350 gnd.n657 gnd.n656 9.3005
R17351 gnd.n6299 gnd.n6298 9.3005
R17352 gnd.n6300 gnd.n655 9.3005
R17353 gnd.n6302 gnd.n6301 9.3005
R17354 gnd.n651 gnd.n650 9.3005
R17355 gnd.n6309 gnd.n6308 9.3005
R17356 gnd.n6310 gnd.n649 9.3005
R17357 gnd.n6312 gnd.n6311 9.3005
R17358 gnd.n645 gnd.n644 9.3005
R17359 gnd.n6319 gnd.n6318 9.3005
R17360 gnd.n6320 gnd.n643 9.3005
R17361 gnd.n6322 gnd.n6321 9.3005
R17362 gnd.n639 gnd.n638 9.3005
R17363 gnd.n6329 gnd.n6328 9.3005
R17364 gnd.n6330 gnd.n637 9.3005
R17365 gnd.n6332 gnd.n6331 9.3005
R17366 gnd.n633 gnd.n632 9.3005
R17367 gnd.n6339 gnd.n6338 9.3005
R17368 gnd.n6340 gnd.n631 9.3005
R17369 gnd.n6342 gnd.n6341 9.3005
R17370 gnd.n627 gnd.n626 9.3005
R17371 gnd.n6349 gnd.n6348 9.3005
R17372 gnd.n6350 gnd.n625 9.3005
R17373 gnd.n6352 gnd.n6351 9.3005
R17374 gnd.n621 gnd.n620 9.3005
R17375 gnd.n6359 gnd.n6358 9.3005
R17376 gnd.n6360 gnd.n619 9.3005
R17377 gnd.n6362 gnd.n6361 9.3005
R17378 gnd.n615 gnd.n614 9.3005
R17379 gnd.n6369 gnd.n6368 9.3005
R17380 gnd.n6370 gnd.n613 9.3005
R17381 gnd.n6372 gnd.n6371 9.3005
R17382 gnd.n609 gnd.n608 9.3005
R17383 gnd.n6379 gnd.n6378 9.3005
R17384 gnd.n6380 gnd.n607 9.3005
R17385 gnd.n6382 gnd.n6381 9.3005
R17386 gnd.n603 gnd.n602 9.3005
R17387 gnd.n6389 gnd.n6388 9.3005
R17388 gnd.n6390 gnd.n601 9.3005
R17389 gnd.n6392 gnd.n6391 9.3005
R17390 gnd.n597 gnd.n596 9.3005
R17391 gnd.n6399 gnd.n6398 9.3005
R17392 gnd.n6400 gnd.n595 9.3005
R17393 gnd.n6402 gnd.n6401 9.3005
R17394 gnd.n591 gnd.n590 9.3005
R17395 gnd.n6409 gnd.n6408 9.3005
R17396 gnd.n6410 gnd.n589 9.3005
R17397 gnd.n6412 gnd.n6411 9.3005
R17398 gnd.n585 gnd.n584 9.3005
R17399 gnd.n6419 gnd.n6418 9.3005
R17400 gnd.n6420 gnd.n583 9.3005
R17401 gnd.n6422 gnd.n6421 9.3005
R17402 gnd.n579 gnd.n578 9.3005
R17403 gnd.n6429 gnd.n6428 9.3005
R17404 gnd.n6430 gnd.n577 9.3005
R17405 gnd.n6432 gnd.n6431 9.3005
R17406 gnd.n573 gnd.n572 9.3005
R17407 gnd.n6439 gnd.n6438 9.3005
R17408 gnd.n6440 gnd.n571 9.3005
R17409 gnd.n6442 gnd.n6441 9.3005
R17410 gnd.n567 gnd.n566 9.3005
R17411 gnd.n6449 gnd.n6448 9.3005
R17412 gnd.n6450 gnd.n565 9.3005
R17413 gnd.n6452 gnd.n6451 9.3005
R17414 gnd.n561 gnd.n560 9.3005
R17415 gnd.n6459 gnd.n6458 9.3005
R17416 gnd.n6460 gnd.n559 9.3005
R17417 gnd.n6462 gnd.n6461 9.3005
R17418 gnd.n555 gnd.n554 9.3005
R17419 gnd.n6469 gnd.n6468 9.3005
R17420 gnd.n6470 gnd.n553 9.3005
R17421 gnd.n6472 gnd.n6471 9.3005
R17422 gnd.n549 gnd.n548 9.3005
R17423 gnd.n6479 gnd.n6478 9.3005
R17424 gnd.n6480 gnd.n547 9.3005
R17425 gnd.n6482 gnd.n6481 9.3005
R17426 gnd.n543 gnd.n542 9.3005
R17427 gnd.n6489 gnd.n6488 9.3005
R17428 gnd.n6490 gnd.n541 9.3005
R17429 gnd.n6492 gnd.n6491 9.3005
R17430 gnd.n537 gnd.n536 9.3005
R17431 gnd.n6499 gnd.n6498 9.3005
R17432 gnd.n6500 gnd.n535 9.3005
R17433 gnd.n6502 gnd.n6501 9.3005
R17434 gnd.n531 gnd.n530 9.3005
R17435 gnd.n6509 gnd.n6508 9.3005
R17436 gnd.n6510 gnd.n529 9.3005
R17437 gnd.n6512 gnd.n6511 9.3005
R17438 gnd.n525 gnd.n524 9.3005
R17439 gnd.n6519 gnd.n6518 9.3005
R17440 gnd.n6520 gnd.n523 9.3005
R17441 gnd.n6522 gnd.n6521 9.3005
R17442 gnd.n519 gnd.n518 9.3005
R17443 gnd.n6529 gnd.n6528 9.3005
R17444 gnd.n6530 gnd.n517 9.3005
R17445 gnd.n6532 gnd.n6531 9.3005
R17446 gnd.n513 gnd.n512 9.3005
R17447 gnd.n6539 gnd.n6538 9.3005
R17448 gnd.n6540 gnd.n511 9.3005
R17449 gnd.n6542 gnd.n6541 9.3005
R17450 gnd.n507 gnd.n506 9.3005
R17451 gnd.n6549 gnd.n6548 9.3005
R17452 gnd.n6550 gnd.n505 9.3005
R17453 gnd.n6552 gnd.n6551 9.3005
R17454 gnd.n501 gnd.n500 9.3005
R17455 gnd.n6559 gnd.n6558 9.3005
R17456 gnd.n6560 gnd.n499 9.3005
R17457 gnd.n6562 gnd.n6561 9.3005
R17458 gnd.n495 gnd.n494 9.3005
R17459 gnd.n6569 gnd.n6568 9.3005
R17460 gnd.n6570 gnd.n493 9.3005
R17461 gnd.n6572 gnd.n6571 9.3005
R17462 gnd.n489 gnd.n488 9.3005
R17463 gnd.n6579 gnd.n6578 9.3005
R17464 gnd.n6580 gnd.n487 9.3005
R17465 gnd.n6582 gnd.n6581 9.3005
R17466 gnd.n483 gnd.n482 9.3005
R17467 gnd.n6589 gnd.n6588 9.3005
R17468 gnd.n6590 gnd.n481 9.3005
R17469 gnd.n6592 gnd.n6591 9.3005
R17470 gnd.n477 gnd.n476 9.3005
R17471 gnd.n6599 gnd.n6598 9.3005
R17472 gnd.n6600 gnd.n475 9.3005
R17473 gnd.n6602 gnd.n6601 9.3005
R17474 gnd.n471 gnd.n470 9.3005
R17475 gnd.n6609 gnd.n6608 9.3005
R17476 gnd.n6610 gnd.n469 9.3005
R17477 gnd.n6612 gnd.n6611 9.3005
R17478 gnd.n465 gnd.n464 9.3005
R17479 gnd.n6619 gnd.n6618 9.3005
R17480 gnd.n6620 gnd.n463 9.3005
R17481 gnd.n6622 gnd.n6621 9.3005
R17482 gnd.n459 gnd.n458 9.3005
R17483 gnd.n6629 gnd.n6628 9.3005
R17484 gnd.n6630 gnd.n457 9.3005
R17485 gnd.n6632 gnd.n6631 9.3005
R17486 gnd.n453 gnd.n452 9.3005
R17487 gnd.n6639 gnd.n6638 9.3005
R17488 gnd.n6640 gnd.n451 9.3005
R17489 gnd.n6642 gnd.n6641 9.3005
R17490 gnd.n447 gnd.n446 9.3005
R17491 gnd.n6649 gnd.n6648 9.3005
R17492 gnd.n6650 gnd.n445 9.3005
R17493 gnd.n6652 gnd.n6651 9.3005
R17494 gnd.n441 gnd.n440 9.3005
R17495 gnd.n6659 gnd.n6658 9.3005
R17496 gnd.n6660 gnd.n439 9.3005
R17497 gnd.n6662 gnd.n6661 9.3005
R17498 gnd.n435 gnd.n434 9.3005
R17499 gnd.n6669 gnd.n6668 9.3005
R17500 gnd.n6670 gnd.n433 9.3005
R17501 gnd.n6672 gnd.n6671 9.3005
R17502 gnd.n429 gnd.n428 9.3005
R17503 gnd.n6679 gnd.n6678 9.3005
R17504 gnd.n6680 gnd.n427 9.3005
R17505 gnd.n6683 gnd.n6681 9.3005
R17506 gnd.n6682 gnd.n423 9.3005
R17507 gnd.n6691 gnd.n422 9.3005
R17508 gnd.n6693 gnd.n6692 9.3005
R17509 gnd.n418 gnd.n417 9.3005
R17510 gnd.n6700 gnd.n6699 9.3005
R17511 gnd.n6701 gnd.n416 9.3005
R17512 gnd.n6703 gnd.n6702 9.3005
R17513 gnd.n412 gnd.n411 9.3005
R17514 gnd.n6710 gnd.n6709 9.3005
R17515 gnd.n6711 gnd.n410 9.3005
R17516 gnd.n6713 gnd.n6712 9.3005
R17517 gnd.n406 gnd.n405 9.3005
R17518 gnd.n6720 gnd.n6719 9.3005
R17519 gnd.n6721 gnd.n404 9.3005
R17520 gnd.n6723 gnd.n6722 9.3005
R17521 gnd.n400 gnd.n399 9.3005
R17522 gnd.n6730 gnd.n6729 9.3005
R17523 gnd.n6731 gnd.n398 9.3005
R17524 gnd.n6733 gnd.n6732 9.3005
R17525 gnd.n394 gnd.n393 9.3005
R17526 gnd.n6740 gnd.n6739 9.3005
R17527 gnd.n6741 gnd.n392 9.3005
R17528 gnd.n6743 gnd.n6742 9.3005
R17529 gnd.n388 gnd.n387 9.3005
R17530 gnd.n6750 gnd.n6749 9.3005
R17531 gnd.n6751 gnd.n386 9.3005
R17532 gnd.n6753 gnd.n6752 9.3005
R17533 gnd.n382 gnd.n381 9.3005
R17534 gnd.n6760 gnd.n6759 9.3005
R17535 gnd.n6761 gnd.n380 9.3005
R17536 gnd.n6763 gnd.n6762 9.3005
R17537 gnd.n376 gnd.n375 9.3005
R17538 gnd.n6770 gnd.n6769 9.3005
R17539 gnd.n6771 gnd.n374 9.3005
R17540 gnd.n6773 gnd.n6772 9.3005
R17541 gnd.n370 gnd.n369 9.3005
R17542 gnd.n6780 gnd.n6779 9.3005
R17543 gnd.n6781 gnd.n368 9.3005
R17544 gnd.n6783 gnd.n6782 9.3005
R17545 gnd.n364 gnd.n363 9.3005
R17546 gnd.n6790 gnd.n6789 9.3005
R17547 gnd.n6791 gnd.n362 9.3005
R17548 gnd.n6793 gnd.n6792 9.3005
R17549 gnd.n358 gnd.n357 9.3005
R17550 gnd.n6800 gnd.n6799 9.3005
R17551 gnd.n6801 gnd.n356 9.3005
R17552 gnd.n6803 gnd.n6802 9.3005
R17553 gnd.n352 gnd.n351 9.3005
R17554 gnd.n6810 gnd.n6809 9.3005
R17555 gnd.n6811 gnd.n350 9.3005
R17556 gnd.n6813 gnd.n6812 9.3005
R17557 gnd.n346 gnd.n345 9.3005
R17558 gnd.n6820 gnd.n6819 9.3005
R17559 gnd.n6821 gnd.n344 9.3005
R17560 gnd.n6823 gnd.n6822 9.3005
R17561 gnd.n340 gnd.n339 9.3005
R17562 gnd.n6830 gnd.n6829 9.3005
R17563 gnd.n6831 gnd.n338 9.3005
R17564 gnd.n6833 gnd.n6832 9.3005
R17565 gnd.n334 gnd.n333 9.3005
R17566 gnd.n6840 gnd.n6839 9.3005
R17567 gnd.n6841 gnd.n332 9.3005
R17568 gnd.n6843 gnd.n6842 9.3005
R17569 gnd.n328 gnd.n327 9.3005
R17570 gnd.n6850 gnd.n6849 9.3005
R17571 gnd.n6851 gnd.n326 9.3005
R17572 gnd.n6853 gnd.n6852 9.3005
R17573 gnd.n322 gnd.n321 9.3005
R17574 gnd.n6860 gnd.n6859 9.3005
R17575 gnd.n6861 gnd.n320 9.3005
R17576 gnd.n6863 gnd.n6862 9.3005
R17577 gnd.n316 gnd.n315 9.3005
R17578 gnd.n6870 gnd.n6869 9.3005
R17579 gnd.n6871 gnd.n314 9.3005
R17580 gnd.n6873 gnd.n6872 9.3005
R17581 gnd.n310 gnd.n309 9.3005
R17582 gnd.n6880 gnd.n6879 9.3005
R17583 gnd.n6881 gnd.n308 9.3005
R17584 gnd.n6883 gnd.n6882 9.3005
R17585 gnd.n304 gnd.n303 9.3005
R17586 gnd.n6890 gnd.n6889 9.3005
R17587 gnd.n6891 gnd.n302 9.3005
R17588 gnd.n6896 gnd.n6892 9.3005
R17589 gnd.n6895 gnd.n6894 9.3005
R17590 gnd.n6893 gnd.n299 9.3005
R17591 gnd.n6690 gnd.n6689 9.3005
R17592 gnd.n7187 gnd.n89 9.3005
R17593 gnd.n7186 gnd.n91 9.3005
R17594 gnd.n96 gnd.n92 9.3005
R17595 gnd.n7181 gnd.n97 9.3005
R17596 gnd.n7180 gnd.n98 9.3005
R17597 gnd.n7179 gnd.n99 9.3005
R17598 gnd.n103 gnd.n100 9.3005
R17599 gnd.n7174 gnd.n104 9.3005
R17600 gnd.n7173 gnd.n105 9.3005
R17601 gnd.n7172 gnd.n106 9.3005
R17602 gnd.n110 gnd.n107 9.3005
R17603 gnd.n7167 gnd.n111 9.3005
R17604 gnd.n7166 gnd.n112 9.3005
R17605 gnd.n7165 gnd.n113 9.3005
R17606 gnd.n117 gnd.n114 9.3005
R17607 gnd.n7160 gnd.n118 9.3005
R17608 gnd.n7159 gnd.n119 9.3005
R17609 gnd.n7155 gnd.n120 9.3005
R17610 gnd.n124 gnd.n121 9.3005
R17611 gnd.n7150 gnd.n125 9.3005
R17612 gnd.n7149 gnd.n126 9.3005
R17613 gnd.n7148 gnd.n127 9.3005
R17614 gnd.n131 gnd.n128 9.3005
R17615 gnd.n7143 gnd.n132 9.3005
R17616 gnd.n7142 gnd.n133 9.3005
R17617 gnd.n7141 gnd.n134 9.3005
R17618 gnd.n138 gnd.n135 9.3005
R17619 gnd.n7136 gnd.n139 9.3005
R17620 gnd.n7135 gnd.n140 9.3005
R17621 gnd.n7134 gnd.n141 9.3005
R17622 gnd.n145 gnd.n142 9.3005
R17623 gnd.n7129 gnd.n146 9.3005
R17624 gnd.n7128 gnd.n147 9.3005
R17625 gnd.n7127 gnd.n148 9.3005
R17626 gnd.n152 gnd.n149 9.3005
R17627 gnd.n7122 gnd.n153 9.3005
R17628 gnd.n7121 gnd.n7120 9.3005
R17629 gnd.n7119 gnd.n156 9.3005
R17630 gnd.n7189 gnd.n7188 9.3005
R17631 gnd.n5569 gnd.n5568 9.3005
R17632 gnd.n5570 gnd.n2802 9.3005
R17633 gnd.n5591 gnd.n5571 9.3005
R17634 gnd.n5590 gnd.n5572 9.3005
R17635 gnd.n5589 gnd.n5573 9.3005
R17636 gnd.n5588 gnd.n5574 9.3005
R17637 gnd.n5587 gnd.n5575 9.3005
R17638 gnd.n5585 gnd.n5576 9.3005
R17639 gnd.n5584 gnd.n5577 9.3005
R17640 gnd.n5581 gnd.n5578 9.3005
R17641 gnd.n5580 gnd.n5579 9.3005
R17642 gnd.n2735 gnd.n2734 9.3005
R17643 gnd.n5681 gnd.n5680 9.3005
R17644 gnd.n5682 gnd.n2733 9.3005
R17645 gnd.n5684 gnd.n5683 9.3005
R17646 gnd.n5685 gnd.n2732 9.3005
R17647 gnd.n5689 gnd.n5688 9.3005
R17648 gnd.n5690 gnd.n2731 9.3005
R17649 gnd.n5714 gnd.n5691 9.3005
R17650 gnd.n5713 gnd.n5692 9.3005
R17651 gnd.n5712 gnd.n5693 9.3005
R17652 gnd.n5711 gnd.n5694 9.3005
R17653 gnd.n5705 gnd.n5695 9.3005
R17654 gnd.n5704 gnd.n5696 9.3005
R17655 gnd.n5703 gnd.n5697 9.3005
R17656 gnd.n5702 gnd.n5699 9.3005
R17657 gnd.n5698 gnd.n263 9.3005
R17658 gnd.n6949 gnd.n264 9.3005
R17659 gnd.n6948 gnd.n265 9.3005
R17660 gnd.n6947 gnd.n266 9.3005
R17661 gnd.n6944 gnd.n267 9.3005
R17662 gnd.n6943 gnd.n268 9.3005
R17663 gnd.n6914 gnd.n269 9.3005
R17664 gnd.n6918 gnd.n6917 9.3005
R17665 gnd.n6919 gnd.n6913 9.3005
R17666 gnd.n6930 gnd.n6920 9.3005
R17667 gnd.n6929 gnd.n6921 9.3005
R17668 gnd.n6928 gnd.n6922 9.3005
R17669 gnd.n6925 gnd.n6924 9.3005
R17670 gnd.n6923 gnd.n160 9.3005
R17671 gnd.n7116 gnd.n159 9.3005
R17672 gnd.n7118 gnd.n7117 9.3005
R17673 gnd.n2804 gnd.n2803 9.3005
R17674 gnd.n3108 gnd.n3107 9.3005
R17675 gnd.n3101 gnd.n3096 9.3005
R17676 gnd.n3114 gnd.n3095 9.3005
R17677 gnd.n3115 gnd.n3094 9.3005
R17678 gnd.n3116 gnd.n3093 9.3005
R17679 gnd.n3092 gnd.n3090 9.3005
R17680 gnd.n3122 gnd.n3089 9.3005
R17681 gnd.n3123 gnd.n3088 9.3005
R17682 gnd.n3124 gnd.n3087 9.3005
R17683 gnd.n3086 gnd.n3084 9.3005
R17684 gnd.n3130 gnd.n3083 9.3005
R17685 gnd.n3131 gnd.n3082 9.3005
R17686 gnd.n3132 gnd.n3081 9.3005
R17687 gnd.n3080 gnd.n3078 9.3005
R17688 gnd.n3138 gnd.n3077 9.3005
R17689 gnd.n3139 gnd.n3076 9.3005
R17690 gnd.n3140 gnd.n3075 9.3005
R17691 gnd.n3074 gnd.n3072 9.3005
R17692 gnd.n3146 gnd.n3071 9.3005
R17693 gnd.n3067 gnd.n3012 9.3005
R17694 gnd.n3066 gnd.n3065 9.3005
R17695 gnd.n3015 gnd.n3014 9.3005
R17696 gnd.n3056 gnd.n3018 9.3005
R17697 gnd.n3058 gnd.n3057 9.3005
R17698 gnd.n3055 gnd.n3020 9.3005
R17699 gnd.n3054 gnd.n3053 9.3005
R17700 gnd.n3022 gnd.n3021 9.3005
R17701 gnd.n3047 gnd.n3046 9.3005
R17702 gnd.n3045 gnd.n3024 9.3005
R17703 gnd.n3044 gnd.n3043 9.3005
R17704 gnd.n3026 gnd.n3025 9.3005
R17705 gnd.n3037 gnd.n3036 9.3005
R17706 gnd.n3035 gnd.n3028 9.3005
R17707 gnd.n3034 gnd.n3033 9.3005
R17708 gnd.n3030 gnd.n3029 9.3005
R17709 gnd.n3106 gnd.n3100 9.3005
R17710 gnd.n3105 gnd.n3104 9.3005
R17711 gnd.n5776 gnd.n2675 9.3005
R17712 gnd.n5775 gnd.n2676 9.3005
R17713 gnd.n2790 gnd.n2677 9.3005
R17714 gnd.n2792 gnd.n2791 9.3005
R17715 gnd.n2770 gnd.n2769 9.3005
R17716 gnd.n5618 gnd.n5617 9.3005
R17717 gnd.n5619 gnd.n2768 9.3005
R17718 gnd.n5623 gnd.n5620 9.3005
R17719 gnd.n5622 gnd.n5621 9.3005
R17720 gnd.n2745 gnd.n2744 9.3005
R17721 gnd.n5671 gnd.n5670 9.3005
R17722 gnd.n5672 gnd.n2743 9.3005
R17723 gnd.n5676 gnd.n5673 9.3005
R17724 gnd.n5675 gnd.n5674 9.3005
R17725 gnd.n2709 gnd.n224 9.3005
R17726 gnd.n6987 gnd.n6986 9.3005
R17727 gnd.n209 gnd.n208 9.3005
R17728 gnd.n7000 gnd.n6999 9.3005
R17729 gnd.n7001 gnd.n207 9.3005
R17730 gnd.n7003 gnd.n7002 9.3005
R17731 gnd.n193 gnd.n192 9.3005
R17732 gnd.n7016 gnd.n7015 9.3005
R17733 gnd.n7017 gnd.n191 9.3005
R17734 gnd.n7019 gnd.n7018 9.3005
R17735 gnd.n177 gnd.n176 9.3005
R17736 gnd.n7032 gnd.n7031 9.3005
R17737 gnd.n7033 gnd.n175 9.3005
R17738 gnd.n7037 gnd.n7034 9.3005
R17739 gnd.n7036 gnd.n7035 9.3005
R17740 gnd.n88 gnd.n87 9.3005
R17741 gnd.n7191 gnd.n7190 9.3005
R17742 gnd.n5777 gnd.n2674 9.3005
R17743 gnd.n6985 gnd.n223 9.3005
R17744 gnd.n4364 gnd.n3929 9.3005
R17745 gnd.n4386 gnd.n4365 9.3005
R17746 gnd.n4385 gnd.n4366 9.3005
R17747 gnd.n4384 gnd.n4367 9.3005
R17748 gnd.n4370 gnd.n4368 9.3005
R17749 gnd.n4380 gnd.n4371 9.3005
R17750 gnd.n4379 gnd.n4372 9.3005
R17751 gnd.n4378 gnd.n4373 9.3005
R17752 gnd.n4376 gnd.n4375 9.3005
R17753 gnd.n4374 gnd.n3904 9.3005
R17754 gnd.n3902 gnd.n3901 9.3005
R17755 gnd.n4447 gnd.n4446 9.3005
R17756 gnd.n4448 gnd.n3900 9.3005
R17757 gnd.n4450 gnd.n4449 9.3005
R17758 gnd.n3898 gnd.n3897 9.3005
R17759 gnd.n4455 gnd.n4454 9.3005
R17760 gnd.n4456 gnd.n3896 9.3005
R17761 gnd.n4458 gnd.n4457 9.3005
R17762 gnd.n3894 gnd.n3893 9.3005
R17763 gnd.n4467 gnd.n4466 9.3005
R17764 gnd.n4468 gnd.n3892 9.3005
R17765 gnd.n4470 gnd.n4469 9.3005
R17766 gnd.n3756 gnd.n3755 9.3005
R17767 gnd.n4480 gnd.n4479 9.3005
R17768 gnd.n4481 gnd.n3754 9.3005
R17769 gnd.n4483 gnd.n4482 9.3005
R17770 gnd.n3750 gnd.n3749 9.3005
R17771 gnd.n4495 gnd.n4494 9.3005
R17772 gnd.n4496 gnd.n3748 9.3005
R17773 gnd.n4503 gnd.n4497 9.3005
R17774 gnd.n4502 gnd.n4498 9.3005
R17775 gnd.n4501 gnd.n4499 9.3005
R17776 gnd.n3478 gnd.n3477 9.3005
R17777 gnd.n4712 gnd.n4711 9.3005
R17778 gnd.n4713 gnd.n3476 9.3005
R17779 gnd.n4715 gnd.n4714 9.3005
R17780 gnd.n3458 gnd.n3457 9.3005
R17781 gnd.n4749 gnd.n4748 9.3005
R17782 gnd.n4750 gnd.n3456 9.3005
R17783 gnd.n4752 gnd.n4751 9.3005
R17784 gnd.n3432 gnd.n3431 9.3005
R17785 gnd.n4790 gnd.n4789 9.3005
R17786 gnd.n4791 gnd.n3430 9.3005
R17787 gnd.n4793 gnd.n4792 9.3005
R17788 gnd.n3416 gnd.n3415 9.3005
R17789 gnd.n4835 gnd.n4834 9.3005
R17790 gnd.n4836 gnd.n3414 9.3005
R17791 gnd.n4840 gnd.n4837 9.3005
R17792 gnd.n4839 gnd.n4838 9.3005
R17793 gnd.n3388 gnd.n3387 9.3005
R17794 gnd.n4907 gnd.n4906 9.3005
R17795 gnd.n4908 gnd.n3386 9.3005
R17796 gnd.n4910 gnd.n4909 9.3005
R17797 gnd.n3367 gnd.n3366 9.3005
R17798 gnd.n4934 gnd.n4933 9.3005
R17799 gnd.n4935 gnd.n3365 9.3005
R17800 gnd.n4937 gnd.n4936 9.3005
R17801 gnd.n3346 gnd.n3345 9.3005
R17802 gnd.n4967 gnd.n4966 9.3005
R17803 gnd.n4968 gnd.n3344 9.3005
R17804 gnd.n4970 gnd.n4969 9.3005
R17805 gnd.n3329 gnd.n3328 9.3005
R17806 gnd.n5012 gnd.n5011 9.3005
R17807 gnd.n5013 gnd.n3327 9.3005
R17808 gnd.n5017 gnd.n5014 9.3005
R17809 gnd.n5016 gnd.n5015 9.3005
R17810 gnd.n3300 gnd.n3299 9.3005
R17811 gnd.n5083 gnd.n5082 9.3005
R17812 gnd.n5084 gnd.n3298 9.3005
R17813 gnd.n5086 gnd.n5085 9.3005
R17814 gnd.n3280 gnd.n3279 9.3005
R17815 gnd.n5110 gnd.n5109 9.3005
R17816 gnd.n5111 gnd.n3278 9.3005
R17817 gnd.n5113 gnd.n5112 9.3005
R17818 gnd.n3258 gnd.n3257 9.3005
R17819 gnd.n5143 gnd.n5142 9.3005
R17820 gnd.n5144 gnd.n3256 9.3005
R17821 gnd.n5146 gnd.n5145 9.3005
R17822 gnd.n3241 gnd.n3240 9.3005
R17823 gnd.n5188 gnd.n5187 9.3005
R17824 gnd.n5189 gnd.n3239 9.3005
R17825 gnd.n5193 gnd.n5190 9.3005
R17826 gnd.n5192 gnd.n5191 9.3005
R17827 gnd.n3213 gnd.n3212 9.3005
R17828 gnd.n5236 gnd.n5235 9.3005
R17829 gnd.n5237 gnd.n3211 9.3005
R17830 gnd.n5239 gnd.n5238 9.3005
R17831 gnd.n3193 gnd.n3192 9.3005
R17832 gnd.n5279 gnd.n5278 9.3005
R17833 gnd.n5280 gnd.n3191 9.3005
R17834 gnd.n5284 gnd.n5281 9.3005
R17835 gnd.n5283 gnd.n5282 9.3005
R17836 gnd.n3164 gnd.n3163 9.3005
R17837 gnd.n5332 gnd.n5331 9.3005
R17838 gnd.n5333 gnd.n3162 9.3005
R17839 gnd.n5335 gnd.n5334 9.3005
R17840 gnd.n2975 gnd.n2974 9.3005
R17841 gnd.n5503 gnd.n5502 9.3005
R17842 gnd.n5504 gnd.n2973 9.3005
R17843 gnd.n5506 gnd.n5505 9.3005
R17844 gnd.n2963 gnd.n2962 9.3005
R17845 gnd.n5526 gnd.n5525 9.3005
R17846 gnd.n5527 gnd.n2961 9.3005
R17847 gnd.n5530 gnd.n5529 9.3005
R17848 gnd.n5528 gnd.n2652 9.3005
R17849 gnd.n5792 gnd.n2653 9.3005
R17850 gnd.n5791 gnd.n2654 9.3005
R17851 gnd.n5790 gnd.n2655 9.3005
R17852 gnd.n2661 gnd.n2656 9.3005
R17853 gnd.n5784 gnd.n2662 9.3005
R17854 gnd.n5783 gnd.n2663 9.3005
R17855 gnd.n5782 gnd.n2664 9.3005
R17856 gnd.n2784 gnd.n2665 9.3005
R17857 gnd.n2785 gnd.n2783 9.3005
R17858 gnd.n2787 gnd.n2786 9.3005
R17859 gnd.n2781 gnd.n2780 9.3005
R17860 gnd.n5607 gnd.n5606 9.3005
R17861 gnd.n5608 gnd.n2779 9.3005
R17862 gnd.n5612 gnd.n5609 9.3005
R17863 gnd.n5611 gnd.n5610 9.3005
R17864 gnd.n2754 gnd.n2753 9.3005
R17865 gnd.n5644 gnd.n5643 9.3005
R17866 gnd.n5645 gnd.n2752 9.3005
R17867 gnd.n5664 gnd.n5646 9.3005
R17868 gnd.n5663 gnd.n5647 9.3005
R17869 gnd.n5662 gnd.n5648 9.3005
R17870 gnd.n5651 gnd.n5649 9.3005
R17871 gnd.n5658 gnd.n5652 9.3005
R17872 gnd.n6955 gnd.n260 9.3005
R17873 gnd.n274 gnd.n261 9.3005
R17874 gnd.n276 gnd.n275 9.3005
R17875 gnd.n277 gnd.n273 9.3005
R17876 gnd.n281 gnd.n280 9.3005
R17877 gnd.n282 gnd.n272 9.3005
R17878 gnd.n6938 gnd.n283 9.3005
R17879 gnd.n6937 gnd.n284 9.3005
R17880 gnd.n6936 gnd.n285 9.3005
R17881 gnd.n288 gnd.n286 9.3005
R17882 gnd.n6911 gnd.n289 9.3005
R17883 gnd.n6910 gnd.n290 9.3005
R17884 gnd.n6909 gnd.n291 9.3005
R17885 gnd.n294 gnd.n292 9.3005
R17886 gnd.n6905 gnd.n295 9.3005
R17887 gnd.n6904 gnd.n296 9.3005
R17888 gnd.n6903 gnd.n297 9.3005
R17889 gnd.n4348 gnd.n4347 9.3005
R17890 gnd.n4245 gnd.n4052 9.3005
R17891 gnd.n4244 gnd.n4053 9.3005
R17892 gnd.n4243 gnd.n4054 9.3005
R17893 gnd.n4206 gnd.n4055 9.3005
R17894 gnd.n4233 gnd.n4207 9.3005
R17895 gnd.n4232 gnd.n4208 9.3005
R17896 gnd.n4231 gnd.n4209 9.3005
R17897 gnd.n4219 gnd.n4210 9.3005
R17898 gnd.n4221 gnd.n4220 9.3005
R17899 gnd.n3965 gnd.n3964 9.3005
R17900 gnd.n4281 gnd.n4280 9.3005
R17901 gnd.n4282 gnd.n3963 9.3005
R17902 gnd.n4284 gnd.n4283 9.3005
R17903 gnd.n3959 gnd.n3958 9.3005
R17904 gnd.n4298 gnd.n4297 9.3005
R17905 gnd.n4299 gnd.n3957 9.3005
R17906 gnd.n4302 gnd.n4301 9.3005
R17907 gnd.n4300 gnd.n3943 9.3005
R17908 gnd.n4350 gnd.n3944 9.3005
R17909 gnd.n4349 gnd.n3945 9.3005
R17910 gnd.n4051 gnd.n3979 9.3005
R17911 gnd.n4044 gnd.n4043 9.3005
R17912 gnd.n4042 gnd.n3985 9.3005
R17913 gnd.n4041 gnd.n4040 9.3005
R17914 gnd.n3987 gnd.n3986 9.3005
R17915 gnd.n4034 gnd.n4033 9.3005
R17916 gnd.n4032 gnd.n3989 9.3005
R17917 gnd.n4031 gnd.n4030 9.3005
R17918 gnd.n3991 gnd.n3990 9.3005
R17919 gnd.n4024 gnd.n4023 9.3005
R17920 gnd.n4022 gnd.n3993 9.3005
R17921 gnd.n4021 gnd.n4020 9.3005
R17922 gnd.n3995 gnd.n3994 9.3005
R17923 gnd.n4014 gnd.n4013 9.3005
R17924 gnd.n4012 gnd.n3997 9.3005
R17925 gnd.n4011 gnd.n4010 9.3005
R17926 gnd.n3999 gnd.n3998 9.3005
R17927 gnd.n4004 gnd.n4003 9.3005
R17928 gnd.n3983 gnd.n3980 9.3005
R17929 gnd.n4050 gnd.n4049 9.3005
R17930 gnd.n4000 gnd.n2335 9.3005
R17931 gnd.n6047 gnd.n2336 9.3005
R17932 gnd.n6046 gnd.n2337 9.3005
R17933 gnd.n6045 gnd.n2338 9.3005
R17934 gnd.n2357 gnd.n2339 9.3005
R17935 gnd.n6035 gnd.n2358 9.3005
R17936 gnd.n6034 gnd.n2359 9.3005
R17937 gnd.n6033 gnd.n2360 9.3005
R17938 gnd.n2379 gnd.n2361 9.3005
R17939 gnd.n6023 gnd.n2380 9.3005
R17940 gnd.n6022 gnd.n2381 9.3005
R17941 gnd.n6021 gnd.n2382 9.3005
R17942 gnd.n2400 gnd.n2383 9.3005
R17943 gnd.n6011 gnd.n2401 9.3005
R17944 gnd.n6010 gnd.n2402 9.3005
R17945 gnd.n6009 gnd.n2403 9.3005
R17946 gnd.n2420 gnd.n2404 9.3005
R17947 gnd.n5998 gnd.n2421 9.3005
R17948 gnd.n5997 gnd.n2422 9.3005
R17949 gnd.n5996 gnd.n2423 9.3005
R17950 gnd.n3953 gnd.n2424 9.3005
R17951 gnd.n5985 gnd.n2437 9.3005
R17952 gnd.n5984 gnd.n2438 9.3005
R17953 gnd.n5983 gnd.n2439 9.3005
R17954 gnd.n2455 gnd.n2440 9.3005
R17955 gnd.n5972 gnd.n2456 9.3005
R17956 gnd.n5971 gnd.n2457 9.3005
R17957 gnd.n5970 gnd.n2458 9.3005
R17958 gnd.n2475 gnd.n2459 9.3005
R17959 gnd.n5960 gnd.n2476 9.3005
R17960 gnd.n5959 gnd.n2477 9.3005
R17961 gnd.n5958 gnd.n2478 9.3005
R17962 gnd.n2497 gnd.n2479 9.3005
R17963 gnd.n5948 gnd.n2498 9.3005
R17964 gnd.n5947 gnd.n2499 9.3005
R17965 gnd.n5946 gnd.n2500 9.3005
R17966 gnd.n2518 gnd.n2501 9.3005
R17967 gnd.n5936 gnd.n2519 9.3005
R17968 gnd.n5935 gnd.n2520 9.3005
R17969 gnd.n5934 gnd.n2521 9.3005
R17970 gnd.n2539 gnd.n2522 9.3005
R17971 gnd.n5924 gnd.n5923 9.3005
R17972 gnd.n4002 gnd.n4001 9.3005
R17973 gnd.n3622 gnd.n3618 9.3005
R17974 gnd.n3655 gnd.n3652 9.3005
R17975 gnd.n3656 gnd.n3651 9.3005
R17976 gnd.n3659 gnd.n3650 9.3005
R17977 gnd.n3660 gnd.n3649 9.3005
R17978 gnd.n3663 gnd.n3648 9.3005
R17979 gnd.n3664 gnd.n3647 9.3005
R17980 gnd.n3667 gnd.n3646 9.3005
R17981 gnd.n3668 gnd.n3645 9.3005
R17982 gnd.n3671 gnd.n3644 9.3005
R17983 gnd.n3672 gnd.n3643 9.3005
R17984 gnd.n3675 gnd.n3642 9.3005
R17985 gnd.n3676 gnd.n3641 9.3005
R17986 gnd.n3677 gnd.n3640 9.3005
R17987 gnd.n3639 gnd.n3636 9.3005
R17988 gnd.n3638 gnd.n3637 9.3005
R17989 gnd.n4583 gnd.n4582 9.3005
R17990 gnd.n3624 gnd.n3623 9.3005
R17991 gnd.n3683 gnd.n3681 9.3005
R17992 gnd.n4575 gnd.n3684 9.3005
R17993 gnd.n4574 gnd.n3685 9.3005
R17994 gnd.n4573 gnd.n3686 9.3005
R17995 gnd.n3690 gnd.n3687 9.3005
R17996 gnd.n4568 gnd.n3691 9.3005
R17997 gnd.n4567 gnd.n3692 9.3005
R17998 gnd.n4566 gnd.n3693 9.3005
R17999 gnd.n3697 gnd.n3694 9.3005
R18000 gnd.n4561 gnd.n3698 9.3005
R18001 gnd.n4560 gnd.n3699 9.3005
R18002 gnd.n4559 gnd.n3700 9.3005
R18003 gnd.n3704 gnd.n3701 9.3005
R18004 gnd.n4554 gnd.n3705 9.3005
R18005 gnd.n4553 gnd.n3706 9.3005
R18006 gnd.n4552 gnd.n3707 9.3005
R18007 gnd.n3712 gnd.n3710 9.3005
R18008 gnd.n4547 gnd.n4546 9.3005
R18009 gnd.n4584 gnd.n3617 9.3005
R18010 gnd.n4200 gnd.n4199 9.3005
R18011 gnd.n4201 gnd.n4056 9.3005
R18012 gnd.n4239 gnd.n4202 9.3005
R18013 gnd.n4238 gnd.n4203 9.3005
R18014 gnd.n4237 gnd.n4204 9.3005
R18015 gnd.n4211 gnd.n4205 9.3005
R18016 gnd.n4227 gnd.n4212 9.3005
R18017 gnd.n4226 gnd.n4213 9.3005
R18018 gnd.n4225 gnd.n4214 9.3005
R18019 gnd.n4218 gnd.n4215 9.3005
R18020 gnd.n4217 gnd.n4216 9.3005
R18021 gnd.n3962 gnd.n3961 9.3005
R18022 gnd.n4289 gnd.n4288 9.3005
R18023 gnd.n4290 gnd.n3960 9.3005
R18024 gnd.n4293 gnd.n4292 9.3005
R18025 gnd.n4291 gnd.n3955 9.3005
R18026 gnd.n4306 gnd.n3956 9.3005
R18027 gnd.n4307 gnd.n3954 9.3005
R18028 gnd.n4309 gnd.n4308 9.3005
R18029 gnd.n4310 gnd.n3952 9.3005
R18030 gnd.n4314 gnd.n4311 9.3005
R18031 gnd.n4315 gnd.n3951 9.3005
R18032 gnd.n4330 gnd.n4329 9.3005
R18033 gnd.n4331 gnd.n3950 9.3005
R18034 gnd.n4337 gnd.n4332 9.3005
R18035 gnd.n4336 gnd.n4333 9.3005
R18036 gnd.n4335 gnd.n4334 9.3005
R18037 gnd.n3922 gnd.n3921 9.3005
R18038 gnd.n4400 gnd.n4399 9.3005
R18039 gnd.n4401 gnd.n3920 9.3005
R18040 gnd.n4403 gnd.n4402 9.3005
R18041 gnd.n3915 gnd.n3914 9.3005
R18042 gnd.n4416 gnd.n4415 9.3005
R18043 gnd.n4417 gnd.n3913 9.3005
R18044 gnd.n4419 gnd.n4418 9.3005
R18045 gnd.n4420 gnd.n3912 9.3005
R18046 gnd.n4424 gnd.n4423 9.3005
R18047 gnd.n4425 gnd.n3911 9.3005
R18048 gnd.n4428 gnd.n4427 9.3005
R18049 gnd.n4426 gnd.n3714 9.3005
R18050 gnd.n4543 gnd.n3713 9.3005
R18051 gnd.n4545 gnd.n4544 9.3005
R18052 gnd.n4198 gnd.n4197 9.3005
R18053 gnd.n4186 gnd.n4061 9.3005
R18054 gnd.n4188 gnd.n4187 9.3005
R18055 gnd.n4185 gnd.n4063 9.3005
R18056 gnd.n4184 gnd.n4183 9.3005
R18057 gnd.n4065 gnd.n4064 9.3005
R18058 gnd.n4177 gnd.n4176 9.3005
R18059 gnd.n4175 gnd.n4067 9.3005
R18060 gnd.n4174 gnd.n4173 9.3005
R18061 gnd.n4069 gnd.n4068 9.3005
R18062 gnd.n4167 gnd.n4166 9.3005
R18063 gnd.n4165 gnd.n4071 9.3005
R18064 gnd.n4164 gnd.n4163 9.3005
R18065 gnd.n4073 gnd.n4072 9.3005
R18066 gnd.n4157 gnd.n4156 9.3005
R18067 gnd.n4155 gnd.n4075 9.3005
R18068 gnd.n4154 gnd.n4153 9.3005
R18069 gnd.n4077 gnd.n4076 9.3005
R18070 gnd.n4147 gnd.n4146 9.3005
R18071 gnd.n4145 gnd.n4079 9.3005
R18072 gnd.n4144 gnd.n4143 9.3005
R18073 gnd.n4081 gnd.n4080 9.3005
R18074 gnd.n4137 gnd.n4136 9.3005
R18075 gnd.n4135 gnd.n4086 9.3005
R18076 gnd.n4134 gnd.n4133 9.3005
R18077 gnd.n4088 gnd.n4087 9.3005
R18078 gnd.n4127 gnd.n4126 9.3005
R18079 gnd.n4125 gnd.n4090 9.3005
R18080 gnd.n4124 gnd.n4123 9.3005
R18081 gnd.n4092 gnd.n4091 9.3005
R18082 gnd.n4117 gnd.n4116 9.3005
R18083 gnd.n4115 gnd.n4094 9.3005
R18084 gnd.n4114 gnd.n4113 9.3005
R18085 gnd.n4096 gnd.n4095 9.3005
R18086 gnd.n4107 gnd.n4106 9.3005
R18087 gnd.n4105 gnd.n4098 9.3005
R18088 gnd.n4104 gnd.n4103 9.3005
R18089 gnd.n4100 gnd.n4099 9.3005
R18090 gnd.n4060 gnd.n4057 9.3005
R18091 gnd.n4196 gnd.n4195 9.3005
R18092 gnd.n6052 gnd.n2326 9.3005
R18093 gnd.n6051 gnd.n2327 9.3005
R18094 gnd.n2346 gnd.n2328 9.3005
R18095 gnd.n6041 gnd.n2347 9.3005
R18096 gnd.n6040 gnd.n2348 9.3005
R18097 gnd.n6039 gnd.n2349 9.3005
R18098 gnd.n2368 gnd.n2350 9.3005
R18099 gnd.n6029 gnd.n2369 9.3005
R18100 gnd.n6028 gnd.n2370 9.3005
R18101 gnd.n6027 gnd.n2371 9.3005
R18102 gnd.n2389 gnd.n2372 9.3005
R18103 gnd.n6017 gnd.n2390 9.3005
R18104 gnd.n6016 gnd.n2391 9.3005
R18105 gnd.n6015 gnd.n2392 9.3005
R18106 gnd.n2411 gnd.n2393 9.3005
R18107 gnd.n2465 gnd.n2448 9.3005
R18108 gnd.n5966 gnd.n2466 9.3005
R18109 gnd.n5965 gnd.n2467 9.3005
R18110 gnd.n5964 gnd.n2468 9.3005
R18111 gnd.n2486 gnd.n2469 9.3005
R18112 gnd.n5954 gnd.n2487 9.3005
R18113 gnd.n5953 gnd.n2488 9.3005
R18114 gnd.n5952 gnd.n2489 9.3005
R18115 gnd.n2507 gnd.n2490 9.3005
R18116 gnd.n5942 gnd.n2508 9.3005
R18117 gnd.n5941 gnd.n2509 9.3005
R18118 gnd.n5940 gnd.n2510 9.3005
R18119 gnd.n2529 gnd.n2511 9.3005
R18120 gnd.n5930 gnd.n2530 9.3005
R18121 gnd.n5929 gnd.n2531 9.3005
R18122 gnd.n5928 gnd.n2532 9.3005
R18123 gnd.n6053 gnd.n2325 9.3005
R18124 gnd.n5976 gnd.n2412 9.3005
R18125 gnd.n865 gnd.n864 9.3005
R18126 gnd.n4251 gnd.n4250 9.3005
R18127 gnd.n4252 gnd.n3977 9.3005
R18128 gnd.n4254 gnd.n4253 9.3005
R18129 gnd.n3975 gnd.n3974 9.3005
R18130 gnd.n4259 gnd.n4258 9.3005
R18131 gnd.n4260 gnd.n3973 9.3005
R18132 gnd.n4262 gnd.n4261 9.3005
R18133 gnd.n3971 gnd.n3970 9.3005
R18134 gnd.n4267 gnd.n4266 9.3005
R18135 gnd.n4268 gnd.n3969 9.3005
R18136 gnd.n4275 gnd.n4269 9.3005
R18137 gnd.n4274 gnd.n4270 9.3005
R18138 gnd.n4273 gnd.n4271 9.3005
R18139 gnd.n3936 gnd.n3935 9.3005
R18140 gnd.n4362 gnd.n4361 9.3005
R18141 gnd.n6059 gnd.n6058 9.3005
R18142 gnd.n6062 gnd.n863 9.3005
R18143 gnd.n862 gnd.n858 9.3005
R18144 gnd.n6068 gnd.n857 9.3005
R18145 gnd.n6069 gnd.n856 9.3005
R18146 gnd.n6070 gnd.n855 9.3005
R18147 gnd.n854 gnd.n850 9.3005
R18148 gnd.n6076 gnd.n849 9.3005
R18149 gnd.n6077 gnd.n848 9.3005
R18150 gnd.n6078 gnd.n847 9.3005
R18151 gnd.n846 gnd.n842 9.3005
R18152 gnd.n6084 gnd.n841 9.3005
R18153 gnd.n6085 gnd.n840 9.3005
R18154 gnd.n6086 gnd.n839 9.3005
R18155 gnd.n838 gnd.n834 9.3005
R18156 gnd.n6092 gnd.n833 9.3005
R18157 gnd.n6093 gnd.n832 9.3005
R18158 gnd.n6094 gnd.n831 9.3005
R18159 gnd.n830 gnd.n826 9.3005
R18160 gnd.n6100 gnd.n825 9.3005
R18161 gnd.n6101 gnd.n824 9.3005
R18162 gnd.n6102 gnd.n823 9.3005
R18163 gnd.n822 gnd.n818 9.3005
R18164 gnd.n6108 gnd.n817 9.3005
R18165 gnd.n6109 gnd.n816 9.3005
R18166 gnd.n6110 gnd.n815 9.3005
R18167 gnd.n814 gnd.n810 9.3005
R18168 gnd.n6116 gnd.n809 9.3005
R18169 gnd.n6117 gnd.n808 9.3005
R18170 gnd.n6118 gnd.n807 9.3005
R18171 gnd.n806 gnd.n802 9.3005
R18172 gnd.n6124 gnd.n801 9.3005
R18173 gnd.n6125 gnd.n800 9.3005
R18174 gnd.n6126 gnd.n799 9.3005
R18175 gnd.n798 gnd.n794 9.3005
R18176 gnd.n6132 gnd.n793 9.3005
R18177 gnd.n6133 gnd.n792 9.3005
R18178 gnd.n6134 gnd.n791 9.3005
R18179 gnd.n790 gnd.n786 9.3005
R18180 gnd.n6140 gnd.n785 9.3005
R18181 gnd.n6141 gnd.n784 9.3005
R18182 gnd.n6142 gnd.n783 9.3005
R18183 gnd.n782 gnd.n778 9.3005
R18184 gnd.n6148 gnd.n777 9.3005
R18185 gnd.n6149 gnd.n776 9.3005
R18186 gnd.n6150 gnd.n775 9.3005
R18187 gnd.n774 gnd.n770 9.3005
R18188 gnd.n6156 gnd.n769 9.3005
R18189 gnd.n6157 gnd.n768 9.3005
R18190 gnd.n6158 gnd.n767 9.3005
R18191 gnd.n766 gnd.n762 9.3005
R18192 gnd.n6164 gnd.n761 9.3005
R18193 gnd.n6165 gnd.n760 9.3005
R18194 gnd.n6166 gnd.n759 9.3005
R18195 gnd.n758 gnd.n754 9.3005
R18196 gnd.n6172 gnd.n753 9.3005
R18197 gnd.n6173 gnd.n752 9.3005
R18198 gnd.n6174 gnd.n751 9.3005
R18199 gnd.n750 gnd.n746 9.3005
R18200 gnd.n6180 gnd.n745 9.3005
R18201 gnd.n6181 gnd.n744 9.3005
R18202 gnd.n6182 gnd.n743 9.3005
R18203 gnd.n742 gnd.n738 9.3005
R18204 gnd.n6188 gnd.n737 9.3005
R18205 gnd.n6189 gnd.n736 9.3005
R18206 gnd.n6190 gnd.n735 9.3005
R18207 gnd.n734 gnd.n730 9.3005
R18208 gnd.n6196 gnd.n729 9.3005
R18209 gnd.n6197 gnd.n728 9.3005
R18210 gnd.n6198 gnd.n727 9.3005
R18211 gnd.n726 gnd.n722 9.3005
R18212 gnd.n6204 gnd.n721 9.3005
R18213 gnd.n6205 gnd.n720 9.3005
R18214 gnd.n6206 gnd.n719 9.3005
R18215 gnd.n718 gnd.n714 9.3005
R18216 gnd.n6212 gnd.n713 9.3005
R18217 gnd.n6213 gnd.n712 9.3005
R18218 gnd.n6214 gnd.n711 9.3005
R18219 gnd.n710 gnd.n706 9.3005
R18220 gnd.n6220 gnd.n705 9.3005
R18221 gnd.n6221 gnd.n704 9.3005
R18222 gnd.n6222 gnd.n703 9.3005
R18223 gnd.n702 gnd.n698 9.3005
R18224 gnd.n6228 gnd.n697 9.3005
R18225 gnd.n6230 gnd.n6229 9.3005
R18226 gnd.n6061 gnd.n6060 9.3005
R18227 gnd.n2866 gnd.n2865 9.3005
R18228 gnd.n2846 gnd.n2844 9.3005
R18229 gnd.n2873 gnd.n2872 9.3005
R18230 gnd.n2840 gnd.n2839 9.3005
R18231 gnd.n2885 gnd.n2884 9.3005
R18232 gnd.n2837 gnd.n2835 9.3005
R18233 gnd.n2892 gnd.n2891 9.3005
R18234 gnd.n2831 gnd.n2830 9.3005
R18235 gnd.n2904 gnd.n2903 9.3005
R18236 gnd.n2828 gnd.n2826 9.3005
R18237 gnd.n2911 gnd.n2910 9.3005
R18238 gnd.n2822 gnd.n2821 9.3005
R18239 gnd.n2923 gnd.n2922 9.3005
R18240 gnd.n2819 gnd.n2817 9.3005
R18241 gnd.n2930 gnd.n2929 9.3005
R18242 gnd.n2811 gnd.n2810 9.3005
R18243 gnd.n2940 gnd.n2939 9.3005
R18244 gnd.n2808 gnd.n2806 9.3005
R18245 gnd.n2849 gnd.n2848 9.3005
R18246 gnd.n2932 gnd.n2931 9.3005
R18247 gnd.n2921 gnd.n2816 9.3005
R18248 gnd.n2920 gnd.n2919 9.3005
R18249 gnd.n2827 gnd.n2823 9.3005
R18250 gnd.n2913 gnd.n2912 9.3005
R18251 gnd.n2902 gnd.n2825 9.3005
R18252 gnd.n2901 gnd.n2900 9.3005
R18253 gnd.n2836 gnd.n2832 9.3005
R18254 gnd.n2894 gnd.n2893 9.3005
R18255 gnd.n2883 gnd.n2834 9.3005
R18256 gnd.n2882 gnd.n2881 9.3005
R18257 gnd.n2845 gnd.n2841 9.3005
R18258 gnd.n2875 gnd.n2874 9.3005
R18259 gnd.n2864 gnd.n2843 9.3005
R18260 gnd.n2863 gnd.n2862 9.3005
R18261 gnd.n2851 gnd.n2850 9.3005
R18262 gnd.n2818 gnd.n2814 9.3005
R18263 gnd.n2938 gnd.n2937 9.3005
R18264 gnd.n5560 gnd.n5559 9.3005
R18265 gnd.n5558 gnd.n2807 9.3005
R18266 gnd.n5557 gnd.n5556 9.3005
R18267 gnd.n5555 gnd.n2948 9.3005
R18268 gnd.n5554 gnd.n5553 9.3005
R18269 gnd.n5552 gnd.n2949 9.3005
R18270 gnd.n5548 gnd.n5547 9.3005
R18271 gnd.n5546 gnd.n2956 9.3005
R18272 gnd.n5545 gnd.n5544 9.3005
R18273 gnd.n5543 gnd.n5538 9.3005
R18274 gnd.n4516 gnd.n3737 9.3005
R18275 gnd.n4515 gnd.n4514 9.3005
R18276 gnd.n4513 gnd.n3741 9.3005
R18277 gnd.n4512 gnd.n4511 9.3005
R18278 gnd.n4510 gnd.n3742 9.3005
R18279 gnd.n4509 gnd.n4508 9.3005
R18280 gnd.n3492 gnd.n3491 9.3005
R18281 gnd.n4680 gnd.n4679 9.3005
R18282 gnd.n4681 gnd.n3489 9.3005
R18283 gnd.n4697 gnd.n4696 9.3005
R18284 gnd.n4695 gnd.n3490 9.3005
R18285 gnd.n4694 gnd.n4693 9.3005
R18286 gnd.n4692 gnd.n4682 9.3005
R18287 gnd.n4691 gnd.n4690 9.3005
R18288 gnd.n4689 gnd.n4686 9.3005
R18289 gnd.n4688 gnd.n4687 9.3005
R18290 gnd.n3446 gnd.n3445 9.3005
R18291 gnd.n4767 gnd.n4766 9.3005
R18292 gnd.n4768 gnd.n3443 9.3005
R18293 gnd.n4777 gnd.n4776 9.3005
R18294 gnd.n4775 gnd.n3444 9.3005
R18295 gnd.n4774 gnd.n4773 9.3005
R18296 gnd.n4772 gnd.n4769 9.3005
R18297 gnd.n3403 gnd.n3402 9.3005
R18298 gnd.n4853 gnd.n4852 9.3005
R18299 gnd.n4854 gnd.n3400 9.3005
R18300 gnd.n4892 gnd.n4891 9.3005
R18301 gnd.n4890 gnd.n3401 9.3005
R18302 gnd.n4889 gnd.n4888 9.3005
R18303 gnd.n4887 gnd.n4855 9.3005
R18304 gnd.n4886 gnd.n4885 9.3005
R18305 gnd.n4884 gnd.n4859 9.3005
R18306 gnd.n4883 gnd.n4882 9.3005
R18307 gnd.n4881 gnd.n4860 9.3005
R18308 gnd.n4880 gnd.n4879 9.3005
R18309 gnd.n4878 gnd.n4864 9.3005
R18310 gnd.n4877 gnd.n4876 9.3005
R18311 gnd.n4875 gnd.n4865 9.3005
R18312 gnd.n4874 gnd.n4873 9.3005
R18313 gnd.n4872 gnd.n4871 9.3005
R18314 gnd.n3315 gnd.n3314 9.3005
R18315 gnd.n5030 gnd.n5029 9.3005
R18316 gnd.n5031 gnd.n3312 9.3005
R18317 gnd.n5069 gnd.n5068 9.3005
R18318 gnd.n5067 gnd.n3313 9.3005
R18319 gnd.n5066 gnd.n5065 9.3005
R18320 gnd.n5064 gnd.n5032 9.3005
R18321 gnd.n5063 gnd.n5062 9.3005
R18322 gnd.n5061 gnd.n5037 9.3005
R18323 gnd.n5060 gnd.n5059 9.3005
R18324 gnd.n5058 gnd.n5038 9.3005
R18325 gnd.n5057 gnd.n5056 9.3005
R18326 gnd.n5055 gnd.n5041 9.3005
R18327 gnd.n5054 gnd.n5053 9.3005
R18328 gnd.n5052 gnd.n5042 9.3005
R18329 gnd.n5051 gnd.n5050 9.3005
R18330 gnd.n5049 gnd.n5048 9.3005
R18331 gnd.n3227 gnd.n3226 9.3005
R18332 gnd.n5207 gnd.n5206 9.3005
R18333 gnd.n5208 gnd.n3224 9.3005
R18334 gnd.n5222 gnd.n5221 9.3005
R18335 gnd.n5220 gnd.n3225 9.3005
R18336 gnd.n5219 gnd.n5218 9.3005
R18337 gnd.n5217 gnd.n5209 9.3005
R18338 gnd.n5216 gnd.n5215 9.3005
R18339 gnd.n5214 gnd.n5213 9.3005
R18340 gnd.n3180 gnd.n3179 9.3005
R18341 gnd.n5299 gnd.n5298 9.3005
R18342 gnd.n5300 gnd.n3177 9.3005
R18343 gnd.n5319 gnd.n5318 9.3005
R18344 gnd.n5317 gnd.n3178 9.3005
R18345 gnd.n5316 gnd.n5315 9.3005
R18346 gnd.n5314 gnd.n5301 9.3005
R18347 gnd.n5313 gnd.n5312 9.3005
R18348 gnd.n5311 gnd.n5310 9.3005
R18349 gnd.n2969 gnd.n2968 9.3005
R18350 gnd.n5513 gnd.n5512 9.3005
R18351 gnd.n5514 gnd.n2967 9.3005
R18352 gnd.n5517 gnd.n5516 9.3005
R18353 gnd.n5515 gnd.n2958 9.3005
R18354 gnd.n5535 gnd.n2957 9.3005
R18355 gnd.n5537 gnd.n5536 9.3005
R18356 gnd.n4518 gnd.n4517 9.3005
R18357 gnd.n4521 gnd.n4520 9.3005
R18358 gnd.n4522 gnd.n3732 9.3005
R18359 gnd.n4524 gnd.n4523 9.3005
R18360 gnd.n4526 gnd.n4525 9.3005
R18361 gnd.n4527 gnd.n3725 9.3005
R18362 gnd.n4529 gnd.n4528 9.3005
R18363 gnd.n4530 gnd.n3724 9.3005
R18364 gnd.n4532 gnd.n4531 9.3005
R18365 gnd.n4533 gnd.n3718 9.3005
R18366 gnd.n4519 gnd.n3736 9.3005
R18367 gnd.n4346 gnd.n3947 9.3005
R18368 gnd.n4345 gnd.n4344 9.3005
R18369 gnd.n4343 gnd.n3948 9.3005
R18370 gnd.n4342 gnd.n4341 9.3005
R18371 gnd.n3925 gnd.n3924 9.3005
R18372 gnd.n4392 gnd.n4391 9.3005
R18373 gnd.n4393 gnd.n3923 9.3005
R18374 gnd.n4395 gnd.n4394 9.3005
R18375 gnd.n3918 gnd.n3917 9.3005
R18376 gnd.n4408 gnd.n4407 9.3005
R18377 gnd.n4409 gnd.n3916 9.3005
R18378 gnd.n4411 gnd.n4410 9.3005
R18379 gnd.n3908 gnd.n3906 9.3005
R18380 gnd.n4439 gnd.n4438 9.3005
R18381 gnd.n4437 gnd.n3907 9.3005
R18382 gnd.n4436 gnd.n4435 9.3005
R18383 gnd.n4434 gnd.n3909 9.3005
R18384 gnd.n4433 gnd.n4432 9.3005
R18385 gnd.n3717 gnd.n3715 9.3005
R18386 gnd.n4539 gnd.n4538 9.3005
R18387 gnd.n4537 gnd.n3716 9.3005
R18388 gnd.n4535 gnd.n4534 9.3005
R18389 gnd.n3720 gnd.n3719 9.3005
R18390 gnd.n3846 gnd.n3845 9.3005
R18391 gnd.n3848 gnd.n3847 9.3005
R18392 gnd.n3826 gnd.n3825 9.3005
R18393 gnd.n3854 gnd.n3853 9.3005
R18394 gnd.n3856 gnd.n3855 9.3005
R18395 gnd.n3816 gnd.n3815 9.3005
R18396 gnd.n3862 gnd.n3861 9.3005
R18397 gnd.n3864 gnd.n3863 9.3005
R18398 gnd.n3803 gnd.n3802 9.3005
R18399 gnd.n3870 gnd.n3869 9.3005
R18400 gnd.n3872 gnd.n3871 9.3005
R18401 gnd.n3793 gnd.n3792 9.3005
R18402 gnd.n3878 gnd.n3877 9.3005
R18403 gnd.n3880 gnd.n3879 9.3005
R18404 gnd.n3778 gnd.n3776 9.3005
R18405 gnd.n3886 gnd.n3885 9.3005
R18406 gnd.n3887 gnd.n3775 9.3005
R18407 gnd.n3780 gnd.n2541 9.3005
R18408 gnd.n3779 gnd.n3777 9.3005
R18409 gnd.n3884 gnd.n3883 9.3005
R18410 gnd.n3882 gnd.n3881 9.3005
R18411 gnd.n3788 gnd.n3787 9.3005
R18412 gnd.n3876 gnd.n3875 9.3005
R18413 gnd.n3874 gnd.n3873 9.3005
R18414 gnd.n3799 gnd.n3798 9.3005
R18415 gnd.n3868 gnd.n3867 9.3005
R18416 gnd.n3866 gnd.n3865 9.3005
R18417 gnd.n3810 gnd.n3809 9.3005
R18418 gnd.n3860 gnd.n3859 9.3005
R18419 gnd.n3858 gnd.n3857 9.3005
R18420 gnd.n3822 gnd.n3821 9.3005
R18421 gnd.n3852 gnd.n3851 9.3005
R18422 gnd.n3850 gnd.n3849 9.3005
R18423 gnd.n3835 gnd.n3834 9.3005
R18424 gnd.n3844 gnd.n3843 9.3005
R18425 gnd.n5918 gnd.n2542 9.3005
R18426 gnd.n5917 gnd.n5916 9.3005
R18427 gnd.n5915 gnd.n2546 9.3005
R18428 gnd.n5914 gnd.n5913 9.3005
R18429 gnd.n5912 gnd.n2547 9.3005
R18430 gnd.n5911 gnd.n5910 9.3005
R18431 gnd.n5909 gnd.n2551 9.3005
R18432 gnd.n5908 gnd.n5907 9.3005
R18433 gnd.n5906 gnd.n2552 9.3005
R18434 gnd.n5905 gnd.n5904 9.3005
R18435 gnd.n5903 gnd.n2556 9.3005
R18436 gnd.n5902 gnd.n5901 9.3005
R18437 gnd.n5900 gnd.n2557 9.3005
R18438 gnd.n5899 gnd.n5898 9.3005
R18439 gnd.n5897 gnd.n2561 9.3005
R18440 gnd.n5896 gnd.n5895 9.3005
R18441 gnd.n5894 gnd.n2562 9.3005
R18442 gnd.n5893 gnd.n5892 9.3005
R18443 gnd.n5891 gnd.n2566 9.3005
R18444 gnd.n5890 gnd.n5889 9.3005
R18445 gnd.n5888 gnd.n2567 9.3005
R18446 gnd.n5887 gnd.n5886 9.3005
R18447 gnd.n5885 gnd.n2571 9.3005
R18448 gnd.n5884 gnd.n5883 9.3005
R18449 gnd.n5882 gnd.n2572 9.3005
R18450 gnd.n5881 gnd.n5880 9.3005
R18451 gnd.n5879 gnd.n2576 9.3005
R18452 gnd.n5878 gnd.n5877 9.3005
R18453 gnd.n5876 gnd.n2577 9.3005
R18454 gnd.n5875 gnd.n5874 9.3005
R18455 gnd.n5873 gnd.n2581 9.3005
R18456 gnd.n5872 gnd.n5871 9.3005
R18457 gnd.n5870 gnd.n2582 9.3005
R18458 gnd.n5869 gnd.n5868 9.3005
R18459 gnd.n5867 gnd.n2586 9.3005
R18460 gnd.n5866 gnd.n5865 9.3005
R18461 gnd.n5864 gnd.n2587 9.3005
R18462 gnd.n5863 gnd.n5862 9.3005
R18463 gnd.n5861 gnd.n2591 9.3005
R18464 gnd.n5860 gnd.n5859 9.3005
R18465 gnd.n5858 gnd.n2592 9.3005
R18466 gnd.n5857 gnd.n5856 9.3005
R18467 gnd.n5855 gnd.n2596 9.3005
R18468 gnd.n5854 gnd.n5853 9.3005
R18469 gnd.n5852 gnd.n2597 9.3005
R18470 gnd.n5851 gnd.n5850 9.3005
R18471 gnd.n5849 gnd.n2601 9.3005
R18472 gnd.n5848 gnd.n5847 9.3005
R18473 gnd.n5846 gnd.n2602 9.3005
R18474 gnd.n5845 gnd.n5844 9.3005
R18475 gnd.n5843 gnd.n2606 9.3005
R18476 gnd.n5842 gnd.n5841 9.3005
R18477 gnd.n5840 gnd.n2607 9.3005
R18478 gnd.n5839 gnd.n5838 9.3005
R18479 gnd.n5837 gnd.n2611 9.3005
R18480 gnd.n5836 gnd.n5835 9.3005
R18481 gnd.n5834 gnd.n2612 9.3005
R18482 gnd.n5833 gnd.n5832 9.3005
R18483 gnd.n5831 gnd.n2616 9.3005
R18484 gnd.n5830 gnd.n5829 9.3005
R18485 gnd.n5828 gnd.n2617 9.3005
R18486 gnd.n5827 gnd.n5826 9.3005
R18487 gnd.n5825 gnd.n2621 9.3005
R18488 gnd.n5824 gnd.n5823 9.3005
R18489 gnd.n5822 gnd.n2622 9.3005
R18490 gnd.n5821 gnd.n5820 9.3005
R18491 gnd.n5819 gnd.n2626 9.3005
R18492 gnd.n5818 gnd.n5817 9.3005
R18493 gnd.n5816 gnd.n2627 9.3005
R18494 gnd.n5815 gnd.n5814 9.3005
R18495 gnd.n5813 gnd.n2631 9.3005
R18496 gnd.n5812 gnd.n5811 9.3005
R18497 gnd.n5810 gnd.n2632 9.3005
R18498 gnd.n5809 gnd.n5808 9.3005
R18499 gnd.n5807 gnd.n2636 9.3005
R18500 gnd.n5806 gnd.n5805 9.3005
R18501 gnd.n5804 gnd.n2637 9.3005
R18502 gnd.n5803 gnd.n5802 9.3005
R18503 gnd.n5801 gnd.n2641 9.3005
R18504 gnd.n5800 gnd.n5799 9.3005
R18505 gnd.n5798 gnd.n2642 9.3005
R18506 gnd.n5797 gnd.n2645 9.3005
R18507 gnd.n5920 gnd.n5919 9.3005
R18508 gnd.n2687 gnd.n2685 9.3005
R18509 gnd.n5771 gnd.n5770 9.3005
R18510 gnd.n5769 gnd.n2686 9.3005
R18511 gnd.n5768 gnd.n5767 9.3005
R18512 gnd.n5766 gnd.n2688 9.3005
R18513 gnd.n5765 gnd.n5764 9.3005
R18514 gnd.n5763 gnd.n2692 9.3005
R18515 gnd.n5762 gnd.n5761 9.3005
R18516 gnd.n5760 gnd.n2693 9.3005
R18517 gnd.n5759 gnd.n5758 9.3005
R18518 gnd.n5757 gnd.n2697 9.3005
R18519 gnd.n5756 gnd.n5755 9.3005
R18520 gnd.n5754 gnd.n2698 9.3005
R18521 gnd.n5753 gnd.n5752 9.3005
R18522 gnd.n5751 gnd.n2702 9.3005
R18523 gnd.n5750 gnd.n5749 9.3005
R18524 gnd.n241 gnd.n239 9.3005
R18525 gnd.n6978 gnd.n6977 9.3005
R18526 gnd.n6976 gnd.n240 9.3005
R18527 gnd.n6975 gnd.n6974 9.3005
R18528 gnd.n6973 gnd.n242 9.3005
R18529 gnd.n6972 gnd.n6971 9.3005
R18530 gnd.n6970 gnd.n246 9.3005
R18531 gnd.n6969 gnd.n6968 9.3005
R18532 gnd.n6967 gnd.n247 9.3005
R18533 gnd.n218 gnd.n217 9.3005
R18534 gnd.n6992 gnd.n6991 9.3005
R18535 gnd.n6993 gnd.n216 9.3005
R18536 gnd.n6995 gnd.n6994 9.3005
R18537 gnd.n201 gnd.n200 9.3005
R18538 gnd.n7008 gnd.n7007 9.3005
R18539 gnd.n7009 gnd.n199 9.3005
R18540 gnd.n7011 gnd.n7010 9.3005
R18541 gnd.n186 gnd.n185 9.3005
R18542 gnd.n7024 gnd.n7023 9.3005
R18543 gnd.n7025 gnd.n184 9.3005
R18544 gnd.n7027 gnd.n7026 9.3005
R18545 gnd.n167 gnd.n166 9.3005
R18546 gnd.n7042 gnd.n7041 9.3005
R18547 gnd.n7043 gnd.n164 9.3005
R18548 gnd.n7112 gnd.n7111 9.3005
R18549 gnd.n7110 gnd.n165 9.3005
R18550 gnd.n2854 gnd.n2853 9.3005
R18551 gnd.n7107 gnd.n7044 9.3005
R18552 gnd.n7106 gnd.n7105 9.3005
R18553 gnd.n7104 gnd.n7049 9.3005
R18554 gnd.n7103 gnd.n7102 9.3005
R18555 gnd.n7101 gnd.n7050 9.3005
R18556 gnd.n7100 gnd.n7099 9.3005
R18557 gnd.n7098 gnd.n7057 9.3005
R18558 gnd.n7097 gnd.n7096 9.3005
R18559 gnd.n7095 gnd.n7058 9.3005
R18560 gnd.n7094 gnd.n7093 9.3005
R18561 gnd.n7092 gnd.n7065 9.3005
R18562 gnd.n7091 gnd.n7090 9.3005
R18563 gnd.n7089 gnd.n7066 9.3005
R18564 gnd.n7088 gnd.n7087 9.3005
R18565 gnd.n7086 gnd.n7073 9.3005
R18566 gnd.n7085 gnd.n7084 9.3005
R18567 gnd.n7083 gnd.n7074 9.3005
R18568 gnd.n7082 gnd.n78 9.3005
R18569 gnd.n7109 gnd.n7108 9.3005
R18570 gnd.n5564 gnd.n5563 9.3005
R18571 gnd.n2800 gnd.n2799 9.3005
R18572 gnd.n5597 gnd.n5596 9.3005
R18573 gnd.n5598 gnd.n2797 9.3005
R18574 gnd.n5601 gnd.n5600 9.3005
R18575 gnd.n5599 gnd.n2798 9.3005
R18576 gnd.n2761 gnd.n2760 9.3005
R18577 gnd.n5628 gnd.n5627 9.3005
R18578 gnd.n5629 gnd.n2758 9.3005
R18579 gnd.n5638 gnd.n5637 9.3005
R18580 gnd.n5636 gnd.n2759 9.3005
R18581 gnd.n5635 gnd.n5634 9.3005
R18582 gnd.n5633 gnd.n5630 9.3005
R18583 gnd.n2715 gnd.n2713 9.3005
R18584 gnd.n5742 gnd.n5741 9.3005
R18585 gnd.n5740 gnd.n2714 9.3005
R18586 gnd.n5739 gnd.n5738 9.3005
R18587 gnd.n5737 gnd.n2716 9.3005
R18588 gnd.n5736 gnd.n5735 9.3005
R18589 gnd.n5734 gnd.n51 9.3005
R18590 gnd.n7227 gnd.n52 9.3005
R18591 gnd.n7226 gnd.n7225 9.3005
R18592 gnd.n7224 gnd.n53 9.3005
R18593 gnd.n7223 gnd.n7222 9.3005
R18594 gnd.n7221 gnd.n57 9.3005
R18595 gnd.n7220 gnd.n7219 9.3005
R18596 gnd.n7218 gnd.n58 9.3005
R18597 gnd.n7217 gnd.n7216 9.3005
R18598 gnd.n7215 gnd.n62 9.3005
R18599 gnd.n7214 gnd.n7213 9.3005
R18600 gnd.n7212 gnd.n63 9.3005
R18601 gnd.n7211 gnd.n7210 9.3005
R18602 gnd.n7209 gnd.n67 9.3005
R18603 gnd.n7208 gnd.n7207 9.3005
R18604 gnd.n7206 gnd.n68 9.3005
R18605 gnd.n7205 gnd.n7204 9.3005
R18606 gnd.n7203 gnd.n72 9.3005
R18607 gnd.n7202 gnd.n7201 9.3005
R18608 gnd.n7200 gnd.n73 9.3005
R18609 gnd.n7199 gnd.n7198 9.3005
R18610 gnd.n7197 gnd.n77 9.3005
R18611 gnd.n7196 gnd.n7195 9.3005
R18612 gnd.n5562 gnd.n2805 9.3005
R18613 gnd.t22 gnd.n1055 9.24152
R18614 gnd.n959 gnd.t80 9.24152
R18615 gnd.n2215 gnd.t70 9.24152
R18616 gnd.n4442 gnd.t159 9.24152
R18617 gnd.n4795 gnd.t168 9.24152
R18618 gnd.n5233 gnd.t170 9.24152
R18619 gnd.t161 gnd.n5614 9.24152
R18620 gnd.t204 gnd.t22 8.92286
R18621 gnd.n4825 gnd.n3425 8.92286
R18622 gnd.n4896 gnd.n4895 8.92286
R18623 gnd.n5002 gnd.n3338 8.92286
R18624 gnd.n5072 gnd.n5071 8.92286
R18625 gnd.n5178 gnd.n3250 8.92286
R18626 gnd.n5225 gnd.n5224 8.92286
R18627 gnd.n5338 gnd.n3158 8.92286
R18628 gnd.n2185 gnd.n2160 8.92171
R18629 gnd.n2153 gnd.n2128 8.92171
R18630 gnd.n2121 gnd.n2096 8.92171
R18631 gnd.n2090 gnd.n2065 8.92171
R18632 gnd.n2058 gnd.n2033 8.92171
R18633 gnd.n2026 gnd.n2001 8.92171
R18634 gnd.n1994 gnd.n1969 8.92171
R18635 gnd.n1963 gnd.n1938 8.92171
R18636 gnd.n5360 gnd.n5342 8.72777
R18637 gnd.n1687 gnd.t24 8.60421
R18638 gnd.n2318 gnd.n2317 8.60421
R18639 gnd.t166 gnd.n5000 8.60421
R18640 gnd.n4987 gnd.t242 8.60421
R18641 gnd.n6900 gnd.n94 8.60421
R18642 gnd.n1119 gnd.n1107 8.43467
R18643 gnd.n38 gnd.n26 8.43467
R18644 gnd.n4347 gnd.n0 8.41456
R18645 gnd.n7228 gnd.n7227 8.41456
R18646 gnd.n1818 gnd.n860 8.28555
R18647 gnd.n4653 gnd.t97 8.28555
R18648 gnd.n4729 gnd.n3440 8.28555
R18649 gnd.n4801 gnd.n3393 8.28555
R18650 gnd.n4956 gnd.n4955 8.28555
R18651 gnd.n4978 gnd.n3305 8.28555
R18652 gnd.n5132 gnd.n5131 8.28555
R18653 gnd.n5154 gnd.n3218 8.28555
R18654 gnd.n5329 gnd.n3166 8.28555
R18655 gnd.n2186 gnd.n2158 8.14595
R18656 gnd.n2154 gnd.n2126 8.14595
R18657 gnd.n2122 gnd.n2094 8.14595
R18658 gnd.n2091 gnd.n2063 8.14595
R18659 gnd.n2059 gnd.n2031 8.14595
R18660 gnd.n2027 gnd.n1999 8.14595
R18661 gnd.n1995 gnd.n1967 8.14595
R18662 gnd.n1964 gnd.n1936 8.14595
R18663 gnd.n2191 gnd.n2190 7.97301
R18664 gnd.t30 gnd.n1202 7.9669
R18665 gnd.n4756 gnd.t201 7.9669
R18666 gnd.n5274 gnd.t225 7.9669
R18667 gnd.n7083 gnd.n7082 7.75808
R18668 gnd.n2937 gnd.n2814 7.75808
R18669 gnd.n3843 gnd.n3834 7.75808
R18670 gnd.n4049 gnd.n3983 7.75808
R18671 gnd.n4729 gnd.t249 7.64824
R18672 gnd.t192 gnd.n3363 7.64824
R18673 gnd.n4861 gnd.t192 7.64824
R18674 gnd.n5035 gnd.t195 7.64824
R18675 gnd.t195 gnd.n3282 7.64824
R18676 gnd.n5154 gnd.t154 7.64824
R18677 gnd.n1596 gnd.t36 7.32958
R18678 gnd.n3516 gnd.n3515 7.30353
R18679 gnd.n5359 gnd.n5358 7.30353
R18680 gnd.n1556 gnd.n1275 7.01093
R18681 gnd.n1278 gnd.n1276 7.01093
R18682 gnd.n1566 gnd.n1565 7.01093
R18683 gnd.n1577 gnd.n1259 7.01093
R18684 gnd.n1576 gnd.n1262 7.01093
R18685 gnd.n1587 gnd.n1250 7.01093
R18686 gnd.n1253 gnd.n1251 7.01093
R18687 gnd.n1597 gnd.n1596 7.01093
R18688 gnd.n1607 gnd.n1231 7.01093
R18689 gnd.n1606 gnd.n1234 7.01093
R18690 gnd.n1615 gnd.n1225 7.01093
R18691 gnd.n1627 gnd.n1215 7.01093
R18692 gnd.n1637 gnd.n1200 7.01093
R18693 gnd.n1653 gnd.n1652 7.01093
R18694 gnd.n1202 gnd.n1139 7.01093
R18695 gnd.n1707 gnd.n1140 7.01093
R18696 gnd.n1701 gnd.n1700 7.01093
R18697 gnd.n1189 gnd.n1151 7.01093
R18698 gnd.n1693 gnd.n1162 7.01093
R18699 gnd.n1180 gnd.n1175 7.01093
R18700 gnd.n1687 gnd.n1686 7.01093
R18701 gnd.n1733 gnd.n1090 7.01093
R18702 gnd.n1732 gnd.n1731 7.01093
R18703 gnd.n1744 gnd.n1743 7.01093
R18704 gnd.n1083 gnd.n1075 7.01093
R18705 gnd.n1773 gnd.n1063 7.01093
R18706 gnd.n1772 gnd.n1066 7.01093
R18707 gnd.n1783 gnd.n1055 7.01093
R18708 gnd.n1056 gnd.n1044 7.01093
R18709 gnd.n1794 gnd.n1045 7.01093
R18710 gnd.n1820 gnd.n1037 7.01093
R18711 gnd.n1819 gnd.n1818 7.01093
R18712 gnd.n1842 gnd.n1841 7.01093
R18713 gnd.n1860 gnd.n1010 7.01093
R18714 gnd.n1859 gnd.n1013 7.01093
R18715 gnd.n1870 gnd.n1002 7.01093
R18716 gnd.n1003 gnd.n990 7.01093
R18717 gnd.n1881 gnd.n991 7.01093
R18718 gnd.n1908 gnd.n975 7.01093
R18719 gnd.n1920 gnd.n1919 7.01093
R18720 gnd.n1902 gnd.n968 7.01093
R18721 gnd.n1931 gnd.n1930 7.01093
R18722 gnd.n2203 gnd.n956 7.01093
R18723 gnd.n2202 gnd.n959 7.01093
R18724 gnd.n2215 gnd.n948 7.01093
R18725 gnd.n949 gnd.n941 7.01093
R18726 gnd.n2225 gnd.n867 7.01093
R18727 gnd.n4700 gnd.n3486 7.01093
R18728 gnd.n4896 gnd.n3397 7.01093
R18729 gnd.t198 gnd.n3351 7.01093
R18730 gnd.n5002 gnd.n5001 7.01093
R18731 gnd.n5072 gnd.n3309 7.01093
R18732 gnd.t233 gnd.n3292 7.01093
R18733 gnd.n5178 gnd.n5177 7.01093
R18734 gnd.n5338 gnd.n5337 7.01093
R18735 gnd.n1234 gnd.t35 6.69227
R18736 gnd.n1066 gnd.t204 6.69227
R18737 gnd.n1909 gnd.t29 6.69227
R18738 gnd.n4779 gnd.t168 6.69227
R18739 gnd.t170 gnd.n5232 6.69227
R18740 gnd.n5492 gnd.n5491 6.5566
R18741 gnd.n4596 gnd.n4595 6.5566
R18742 gnd.n3612 gnd.n3558 6.5566
R18743 gnd.n5370 gnd.n5369 6.5566
R18744 gnd.n4725 gnd.n3466 6.37362
R18745 gnd.n4763 gnd.n4762 6.37362
R18746 gnd.n4920 gnd.n3376 6.37362
R18747 gnd.n5123 gnd.n3269 6.37362
R18748 gnd.n5249 gnd.n3201 6.37362
R18749 gnd.n5296 gnd.n5295 6.37362
R18750 gnd.t74 gnd.n3153 6.37362
R18751 gnd.n4523 gnd.n3731 6.20656
R18752 gnd.n7158 gnd.n7155 6.20656
R18753 gnd.n4084 gnd.n4079 6.20656
R18754 gnd.n5551 gnd.n5548 6.20656
R18755 gnd.t282 gnd.n1663 6.05496
R18756 gnd.n1664 gnd.t33 6.05496
R18757 gnd.t179 gnd.n1090 6.05496
R18758 gnd.t32 gnd.n1830 6.05496
R18759 gnd.n4248 gnd.t129 6.05496
R18760 gnd.n4668 gnd.n3521 6.05496
R18761 gnd.t51 gnd.n162 6.05496
R18762 gnd.n2188 gnd.n2158 5.81868
R18763 gnd.n2156 gnd.n2126 5.81868
R18764 gnd.n2124 gnd.n2094 5.81868
R18765 gnd.n2093 gnd.n2063 5.81868
R18766 gnd.n2061 gnd.n2031 5.81868
R18767 gnd.n2029 gnd.n1999 5.81868
R18768 gnd.n1997 gnd.n1967 5.81868
R18769 gnd.n1966 gnd.n1936 5.81868
R18770 gnd.n4677 gnd.t63 5.73631
R18771 gnd.t63 gnd.n4676 5.73631
R18772 gnd.t84 gnd.n4745 5.73631
R18773 gnd.n4825 gnd.t250 5.73631
R18774 gnd.n4817 gnd.n4816 5.73631
R18775 gnd.n4842 gnd.n3411 5.73631
R18776 gnd.t232 gnd.n3369 5.73631
R18777 gnd.n5001 gnd.t252 5.73631
R18778 gnd.n4994 gnd.n3323 5.73631
R18779 gnd.n5019 gnd.n3317 5.73631
R18780 gnd.t2 gnd.n3309 5.73631
R18781 gnd.n3276 gnd.t231 5.73631
R18782 gnd.n5170 gnd.n3235 5.73631
R18783 gnd.n5195 gnd.n3229 5.73631
R18784 gnd.n5225 gnd.t172 5.73631
R18785 gnd.n5263 gnd.t120 5.73631
R18786 gnd.n5496 gnd.n3148 5.62001
R18787 gnd.n4591 gnd.n4588 5.62001
R18788 gnd.n4588 gnd.n3616 5.62001
R18789 gnd.n5365 gnd.n3148 5.62001
R18790 gnd.n1415 gnd.n1410 5.4308
R18791 gnd.n2233 gnd.n934 5.4308
R18792 gnd.n1731 gnd.t31 5.41765
R18793 gnd.t23 gnd.n1754 5.41765
R18794 gnd.t222 gnd.n1022 5.41765
R18795 gnd.n4850 gnd.t199 5.41765
R18796 gnd.t190 gnd.n3245 5.41765
R18797 gnd.t126 gnd.n4699 5.09899
R18798 gnd.n4745 gnd.n4743 5.09899
R18799 gnd.n4756 gnd.n4755 5.09899
R18800 gnd.t16 gnd.n3381 5.09899
R18801 gnd.n4930 gnd.n4929 5.09899
R18802 gnd.n4941 gnd.n4940 5.09899
R18803 gnd.n5106 gnd.n5105 5.09899
R18804 gnd.n5117 gnd.n5116 5.09899
R18805 gnd.t218 gnd.n3262 5.09899
R18806 gnd.n5275 gnd.n5274 5.09899
R18807 gnd.n5289 gnd.n5288 5.09899
R18808 gnd.n2186 gnd.n2185 5.04292
R18809 gnd.n2154 gnd.n2153 5.04292
R18810 gnd.n2122 gnd.n2121 5.04292
R18811 gnd.n2091 gnd.n2090 5.04292
R18812 gnd.n2059 gnd.n2058 5.04292
R18813 gnd.n2027 gnd.n2026 5.04292
R18814 gnd.n1995 gnd.n1994 5.04292
R18815 gnd.n1964 gnd.n1963 5.04292
R18816 gnd.n1131 gnd.n1130 4.82753
R18817 gnd.n50 gnd.n49 4.82753
R18818 gnd.n1694 gnd.t26 4.78034
R18819 gnd.n1045 gnd.t27 4.78034
R18820 gnd.t181 gnd.n4505 4.78034
R18821 gnd.n3411 gnd.t199 4.78034
R18822 gnd.n5170 gnd.t190 4.78034
R18823 gnd.n5499 gnd.t136 4.78034
R18824 gnd.n5306 gnd.t0 4.78034
R18825 gnd.n1136 gnd.n1133 4.74817
R18826 gnd.n1186 gnd.n1096 4.74817
R18827 gnd.n1173 gnd.n1095 4.74817
R18828 gnd.n1094 gnd.n1093 4.74817
R18829 gnd.n1182 gnd.n1133 4.74817
R18830 gnd.n1183 gnd.n1096 4.74817
R18831 gnd.n1185 gnd.n1095 4.74817
R18832 gnd.n1172 gnd.n1094 4.74817
R18833 gnd.n6984 gnd.n6983 4.74817
R18834 gnd.n5729 gnd.n229 4.74817
R18835 gnd.n2724 gnd.n228 4.74817
R18836 gnd.n253 gnd.n227 4.74817
R18837 gnd.n6963 gnd.n226 4.74817
R18838 gnd.n6984 gnd.n230 4.74817
R18839 gnd.n6982 gnd.n229 4.74817
R18840 gnd.n5730 gnd.n228 4.74817
R18841 gnd.n2723 gnd.n227 4.74817
R18842 gnd.n254 gnd.n226 4.74817
R18843 gnd.n3937 gnd.n3934 4.74817
R18844 gnd.n3941 gnd.n3933 4.74817
R18845 gnd.n4323 gnd.n3932 4.74817
R18846 gnd.n4321 gnd.n3931 4.74817
R18847 gnd.n4317 gnd.n3930 4.74817
R18848 gnd.n5656 gnd.n5655 4.74817
R18849 gnd.n5719 gnd.n2729 4.74817
R18850 gnd.n5724 gnd.n5721 4.74817
R18851 gnd.n5722 gnd.n259 4.74817
R18852 gnd.n6957 gnd.n6956 4.74817
R18853 gnd.n5657 gnd.n5656 4.74817
R18854 gnd.n5653 gnd.n2729 4.74817
R18855 gnd.n5721 gnd.n5720 4.74817
R18856 gnd.n5723 gnd.n5722 4.74817
R18857 gnd.n6958 gnd.n6957 4.74817
R18858 gnd.n6004 gnd.n6003 4.74817
R18859 gnd.n2430 gnd.n2413 4.74817
R18860 gnd.n5991 gnd.n5990 4.74817
R18861 gnd.n2447 gnd.n2431 4.74817
R18862 gnd.n5978 gnd.n5977 4.74817
R18863 gnd.n6005 gnd.n6004 4.74817
R18864 gnd.n6002 gnd.n2413 4.74817
R18865 gnd.n5992 gnd.n5991 4.74817
R18866 gnd.n5989 gnd.n2431 4.74817
R18867 gnd.n5979 gnd.n5978 4.74817
R18868 gnd.n4357 gnd.n3934 4.74817
R18869 gnd.n4356 gnd.n3933 4.74817
R18870 gnd.n3940 gnd.n3932 4.74817
R18871 gnd.n4324 gnd.n3931 4.74817
R18872 gnd.n4320 gnd.n3930 4.74817
R18873 gnd.n1119 gnd.n1118 4.7074
R18874 gnd.n38 gnd.n37 4.7074
R18875 gnd.n1131 gnd.n1119 4.65959
R18876 gnd.n50 gnd.n38 4.65959
R18877 gnd.n3147 gnd.n3068 4.6132
R18878 gnd.n4586 gnd.n4585 4.6132
R18879 gnd.n4676 gnd.n3496 4.46168
R18880 gnd.n4653 gnd.t59 4.46168
R18881 gnd.n4832 gnd.n4831 4.46168
R18882 gnd.n4849 gnd.n3406 4.46168
R18883 gnd.n5009 gnd.n5008 4.46168
R18884 gnd.n5026 gnd.n3319 4.46168
R18885 gnd.n5185 gnd.n5184 4.46168
R18886 gnd.n5202 gnd.n3231 4.46168
R18887 gnd.t109 gnd.n3166 4.46168
R18888 gnd.n5431 gnd.n3153 4.46168
R18889 gnd.n5355 gnd.n5342 4.46111
R18890 gnd.n2171 gnd.n2167 4.38594
R18891 gnd.n2139 gnd.n2135 4.38594
R18892 gnd.n2107 gnd.n2103 4.38594
R18893 gnd.n2076 gnd.n2072 4.38594
R18894 gnd.n2044 gnd.n2040 4.38594
R18895 gnd.n2012 gnd.n2008 4.38594
R18896 gnd.n1980 gnd.n1976 4.38594
R18897 gnd.n1949 gnd.n1945 4.38594
R18898 gnd.n2182 gnd.n2160 4.26717
R18899 gnd.n2150 gnd.n2128 4.26717
R18900 gnd.n2118 gnd.n2096 4.26717
R18901 gnd.n2087 gnd.n2065 4.26717
R18902 gnd.n2055 gnd.n2033 4.26717
R18903 gnd.n2023 gnd.n2001 4.26717
R18904 gnd.n1991 gnd.n1969 4.26717
R18905 gnd.n1960 gnd.n1938 4.26717
R18906 gnd.n1638 gnd.t28 4.14303
R18907 gnd.n1870 gnd.t25 4.14303
R18908 gnd.t66 gnd.n2527 4.14303
R18909 gnd.n4947 gnd.t270 4.14303
R18910 gnd.n5096 gnd.t227 4.14303
R18911 gnd.t55 gnd.n2679 4.14303
R18912 gnd.n2190 gnd.n2189 4.08274
R18913 gnd.n5491 gnd.n5490 4.05904
R18914 gnd.n4597 gnd.n4596 4.05904
R18915 gnd.n3609 gnd.n3558 4.05904
R18916 gnd.n5371 gnd.n5370 4.05904
R18917 gnd.n15 gnd.n7 3.99943
R18918 gnd.n4700 gnd.t126 3.82437
R18919 gnd.n3474 gnd.n3473 3.82437
R18920 gnd.n4733 gnd.n3434 3.82437
R18921 gnd.t5 gnd.n3397 3.82437
R18922 gnd.n3384 gnd.n3383 3.82437
R18923 gnd.n4949 gnd.n3349 3.82437
R18924 gnd.n3296 gnd.n3294 3.82437
R18925 gnd.n5125 gnd.n3260 3.82437
R18926 gnd.n5177 gnd.t183 3.82437
R18927 gnd.n3209 gnd.n3208 3.82437
R18928 gnd.n5295 gnd.t120 3.82437
R18929 gnd.n5265 gnd.n5264 3.82437
R18930 gnd.n2190 gnd.n2062 3.70378
R18931 gnd.n1711 gnd.n1132 3.65935
R18932 gnd.n15 gnd.n14 3.60163
R18933 gnd.n2181 gnd.n2162 3.49141
R18934 gnd.n2149 gnd.n2130 3.49141
R18935 gnd.n2117 gnd.n2098 3.49141
R18936 gnd.n2086 gnd.n2067 3.49141
R18937 gnd.n2054 gnd.n2035 3.49141
R18938 gnd.n2022 gnd.n2003 3.49141
R18939 gnd.n1990 gnd.n1971 3.49141
R18940 gnd.n1959 gnd.n1940 3.49141
R18941 gnd.n4709 gnd.n3480 3.18706
R18942 gnd.t59 gnd.n3471 3.18706
R18943 gnd.n4796 gnd.n4795 3.18706
R18944 gnd.n4904 gnd.n3390 3.18706
R18945 gnd.n4973 gnd.n4972 3.18706
R18946 gnd.n5080 gnd.n3302 3.18706
R18947 gnd.n5149 gnd.n5148 3.18706
R18948 gnd.n5233 gnd.n3215 3.18706
R18949 gnd.n5321 gnd.t109 3.18706
R18950 gnd.n5256 gnd.n5255 3.18706
R18951 gnd.n1217 gnd.t28 2.8684
R18952 gnd.n4742 gnd.t201 2.8684
R18953 gnd.t225 gnd.n3187 2.8684
R18954 gnd.n1120 gnd.t184 2.82907
R18955 gnd.n1120 gnd.t197 2.82907
R18956 gnd.n1122 gnd.t247 2.82907
R18957 gnd.n1122 gnd.t189 2.82907
R18958 gnd.n1124 gnd.t241 2.82907
R18959 gnd.n1124 gnd.t256 2.82907
R18960 gnd.n1126 gnd.t13 2.82907
R18961 gnd.n1126 gnd.t234 2.82907
R18962 gnd.n1128 gnd.t258 2.82907
R18963 gnd.n1128 gnd.t272 2.82907
R18964 gnd.n1097 gnd.t42 2.82907
R18965 gnd.n1097 gnd.t269 2.82907
R18966 gnd.n1099 gnd.t262 2.82907
R18967 gnd.n1099 gnd.t230 2.82907
R18968 gnd.n1101 gnd.t267 2.82907
R18969 gnd.n1101 gnd.t266 2.82907
R18970 gnd.n1103 gnd.t239 2.82907
R18971 gnd.n1103 gnd.t285 2.82907
R18972 gnd.n1105 gnd.t19 2.82907
R18973 gnd.n1105 gnd.t217 2.82907
R18974 gnd.n1108 gnd.t187 2.82907
R18975 gnd.n1108 gnd.t264 2.82907
R18976 gnd.n1110 gnd.t263 2.82907
R18977 gnd.n1110 gnd.t219 2.82907
R18978 gnd.n1112 gnd.t39 2.82907
R18979 gnd.n1112 gnd.t221 2.82907
R18980 gnd.n1114 gnd.t240 2.82907
R18981 gnd.n1114 gnd.t21 2.82907
R18982 gnd.n1116 gnd.t245 2.82907
R18983 gnd.n1116 gnd.t265 2.82907
R18984 gnd.n47 gnd.t203 2.82907
R18985 gnd.n47 gnd.t185 2.82907
R18986 gnd.n45 gnd.t229 2.82907
R18987 gnd.n45 gnd.t174 2.82907
R18988 gnd.n43 gnd.t274 2.82907
R18989 gnd.n43 gnd.t4 2.82907
R18990 gnd.n41 gnd.t7 2.82907
R18991 gnd.n41 gnd.t273 2.82907
R18992 gnd.n39 gnd.t257 2.82907
R18993 gnd.n39 gnd.t9 2.82907
R18994 gnd.n24 gnd.t44 2.82907
R18995 gnd.n24 gnd.t158 2.82907
R18996 gnd.n22 gnd.t210 2.82907
R18997 gnd.n22 gnd.t284 2.82907
R18998 gnd.n20 gnd.t260 2.82907
R18999 gnd.n20 gnd.t211 2.82907
R19000 gnd.n18 gnd.t40 2.82907
R19001 gnd.n18 gnd.t165 2.82907
R19002 gnd.n16 gnd.t215 2.82907
R19003 gnd.n16 gnd.t275 2.82907
R19004 gnd.n35 gnd.t286 2.82907
R19005 gnd.n35 gnd.t254 2.82907
R19006 gnd.n33 gnd.t244 2.82907
R19007 gnd.n33 gnd.t238 2.82907
R19008 gnd.n31 gnd.t268 2.82907
R19009 gnd.n31 gnd.t235 2.82907
R19010 gnd.n29 gnd.t45 2.82907
R19011 gnd.n29 gnd.t287 2.82907
R19012 gnd.n27 gnd.t176 2.82907
R19013 gnd.n27 gnd.t17 2.82907
R19014 gnd.n2178 gnd.n2177 2.71565
R19015 gnd.n2146 gnd.n2145 2.71565
R19016 gnd.n2114 gnd.n2113 2.71565
R19017 gnd.n2083 gnd.n2082 2.71565
R19018 gnd.n2051 gnd.n2050 2.71565
R19019 gnd.n2019 gnd.n2018 2.71565
R19020 gnd.n1987 gnd.n1986 2.71565
R19021 gnd.n1956 gnd.n1955 2.71565
R19022 gnd.n4708 gnd.n4706 2.54975
R19023 gnd.n4780 gnd.n4779 2.54975
R19024 gnd.n4843 gnd.t251 2.54975
R19025 gnd.n4903 gnd.n4902 2.54975
R19026 gnd.n4801 gnd.t16 2.54975
R19027 gnd.n4957 gnd.n3342 2.54975
R19028 gnd.n5079 gnd.n5078 2.54975
R19029 gnd.n5131 gnd.t218 2.54975
R19030 gnd.n5133 gnd.n3254 2.54975
R19031 gnd.n5196 gnd.t224 2.54975
R19032 gnd.n5232 gnd.n5231 2.54975
R19033 gnd.n5328 gnd.n3169 2.54975
R19034 gnd.n1711 gnd.n1133 2.27742
R19035 gnd.n1711 gnd.n1096 2.27742
R19036 gnd.n1711 gnd.n1095 2.27742
R19037 gnd.n1711 gnd.n1094 2.27742
R19038 gnd.n6985 gnd.n6984 2.27742
R19039 gnd.n6985 gnd.n229 2.27742
R19040 gnd.n6985 gnd.n228 2.27742
R19041 gnd.n6985 gnd.n227 2.27742
R19042 gnd.n6985 gnd.n226 2.27742
R19043 gnd.n5656 gnd.n225 2.27742
R19044 gnd.n2729 gnd.n225 2.27742
R19045 gnd.n5721 gnd.n225 2.27742
R19046 gnd.n5722 gnd.n225 2.27742
R19047 gnd.n6957 gnd.n225 2.27742
R19048 gnd.n6004 gnd.n2412 2.27742
R19049 gnd.n2413 gnd.n2412 2.27742
R19050 gnd.n5991 gnd.n2412 2.27742
R19051 gnd.n2431 gnd.n2412 2.27742
R19052 gnd.n5978 gnd.n2412 2.27742
R19053 gnd.n4363 gnd.n3934 2.27742
R19054 gnd.n4363 gnd.n3933 2.27742
R19055 gnd.n4363 gnd.n3932 2.27742
R19056 gnd.n4363 gnd.n3931 2.27742
R19057 gnd.n4363 gnd.n3930 2.27742
R19058 gnd.n1565 gnd.t47 2.23109
R19059 gnd.n1188 gnd.t26 2.23109
R19060 gnd.n4861 gnd.t270 2.23109
R19061 gnd.n5035 gnd.t227 2.23109
R19062 gnd.n2174 gnd.n2164 1.93989
R19063 gnd.n2142 gnd.n2132 1.93989
R19064 gnd.n2110 gnd.n2100 1.93989
R19065 gnd.n2079 gnd.n2069 1.93989
R19066 gnd.n2047 gnd.n2037 1.93989
R19067 gnd.n2015 gnd.n2005 1.93989
R19068 gnd.n1983 gnd.n1973 1.93989
R19069 gnd.n1952 gnd.n1942 1.93989
R19070 gnd.n4718 gnd.n4717 1.91244
R19071 gnd.n4787 gnd.n4786 1.91244
R19072 gnd.n4964 gnd.n4963 1.91244
R19073 gnd.n5089 gnd.n5088 1.91244
R19074 gnd.n5242 gnd.n5241 1.91244
R19075 gnd.n5322 gnd.n3173 1.91244
R19076 gnd.t280 gnd.n1576 1.59378
R19077 gnd.n1755 gnd.t23 1.59378
R19078 gnd.n1030 gnd.t222 1.59378
R19079 gnd.t14 gnd.n4912 1.59378
R19080 gnd.n5140 gnd.t155 1.59378
R19081 gnd.n4661 gnd.n4660 1.27512
R19082 gnd.n3473 gnd.t145 1.27512
R19083 gnd.t250 gnd.n4824 1.27512
R19084 gnd.n4823 gnd.n3418 1.27512
R19085 gnd.n4809 gnd.n4808 1.27512
R19086 gnd.n5000 gnd.n3332 1.27512
R19087 gnd.n4987 gnd.n4986 1.27512
R19088 gnd.n5176 gnd.n3243 1.27512
R19089 gnd.n5163 gnd.n5161 1.27512
R19090 gnd.n5162 gnd.t172 1.27512
R19091 gnd.n5256 gnd.t123 1.27512
R19092 gnd.n5303 gnd.n3160 1.27512
R19093 gnd.n5308 gnd.t136 1.27512
R19094 gnd.n1418 gnd.n1410 1.16414
R19095 gnd.n2236 gnd.n934 1.16414
R19096 gnd.n2173 gnd.n2166 1.16414
R19097 gnd.n2141 gnd.n2134 1.16414
R19098 gnd.n2109 gnd.n2102 1.16414
R19099 gnd.n2078 gnd.n2071 1.16414
R19100 gnd.n2046 gnd.n2039 1.16414
R19101 gnd.n2014 gnd.n2007 1.16414
R19102 gnd.n1982 gnd.n1975 1.16414
R19103 gnd.n1951 gnd.n1944 1.16414
R19104 gnd.n3147 gnd.n3146 0.970197
R19105 gnd.n4586 gnd.n3617 0.970197
R19106 gnd.n2157 gnd.n2125 0.962709
R19107 gnd.n2189 gnd.n2157 0.962709
R19108 gnd.n2030 gnd.n1998 0.962709
R19109 gnd.n2062 gnd.n2030 0.962709
R19110 gnd.n1664 gnd.t282 0.956468
R19111 gnd.n1831 gnd.t32 0.956468
R19112 gnd.t212 gnd.n2355 0.956468
R19113 gnd.n4223 gnd.t18 0.956468
R19114 gnd.n3919 gnd.t41 0.956468
R19115 gnd.n4413 gnd.t196 0.956468
R19116 gnd.t276 gnd.n4708 0.956468
R19117 gnd.t206 gnd.n3169 0.956468
R19118 gnd.n5582 gnd.t175 0.956468
R19119 gnd.n5666 gnd.t8 0.956468
R19120 gnd.n7013 gnd.t157 0.956468
R19121 gnd.n6933 gnd.t10 0.956468
R19122 gnd.n1127 gnd.n1125 0.773756
R19123 gnd.n46 gnd.n44 0.773756
R19124 gnd.n1130 gnd.n1129 0.773756
R19125 gnd.n1129 gnd.n1127 0.773756
R19126 gnd.n1125 gnd.n1123 0.773756
R19127 gnd.n1123 gnd.n1121 0.773756
R19128 gnd.n42 gnd.n40 0.773756
R19129 gnd.n44 gnd.n42 0.773756
R19130 gnd.n48 gnd.n46 0.773756
R19131 gnd.n49 gnd.n48 0.773756
R19132 gnd.n2 gnd.n1 0.672012
R19133 gnd.n3 gnd.n2 0.672012
R19134 gnd.n4 gnd.n3 0.672012
R19135 gnd.n5 gnd.n4 0.672012
R19136 gnd.n6 gnd.n5 0.672012
R19137 gnd.n7 gnd.n6 0.672012
R19138 gnd.n9 gnd.n8 0.672012
R19139 gnd.n10 gnd.n9 0.672012
R19140 gnd.n11 gnd.n10 0.672012
R19141 gnd.n12 gnd.n11 0.672012
R19142 gnd.n13 gnd.n12 0.672012
R19143 gnd.n14 gnd.n13 0.672012
R19144 gnd.n4746 gnd.n3460 0.637812
R19145 gnd.n4754 gnd.n3454 0.637812
R19146 gnd.n3454 gnd.t248 0.637812
R19147 gnd.n4931 gnd.n3369 0.637812
R19148 gnd.n4939 gnd.n3363 0.637812
R19149 gnd.n4955 gnd.t198 0.637812
R19150 gnd.n4978 gnd.t233 0.637812
R19151 gnd.n5107 gnd.n3282 0.637812
R19152 gnd.n5115 gnd.n3276 0.637812
R19153 gnd.t208 gnd.n3195 0.637812
R19154 gnd.n5276 gnd.n3195 0.637812
R19155 gnd.n5286 gnd.n3182 0.637812
R19156 gnd.t100 gnd.n5321 0.637812
R19157 gnd.n1107 gnd.n1106 0.573776
R19158 gnd.n1106 gnd.n1104 0.573776
R19159 gnd.n1104 gnd.n1102 0.573776
R19160 gnd.n1102 gnd.n1100 0.573776
R19161 gnd.n1100 gnd.n1098 0.573776
R19162 gnd.n1118 gnd.n1117 0.573776
R19163 gnd.n1117 gnd.n1115 0.573776
R19164 gnd.n1115 gnd.n1113 0.573776
R19165 gnd.n1113 gnd.n1111 0.573776
R19166 gnd.n1111 gnd.n1109 0.573776
R19167 gnd.n19 gnd.n17 0.573776
R19168 gnd.n21 gnd.n19 0.573776
R19169 gnd.n23 gnd.n21 0.573776
R19170 gnd.n25 gnd.n23 0.573776
R19171 gnd.n26 gnd.n25 0.573776
R19172 gnd.n30 gnd.n28 0.573776
R19173 gnd.n32 gnd.n30 0.573776
R19174 gnd.n34 gnd.n32 0.573776
R19175 gnd.n36 gnd.n34 0.573776
R19176 gnd.n37 gnd.n36 0.573776
R19177 gnd gnd.n0 0.551497
R19178 gnd.n6985 gnd.n225 0.548625
R19179 gnd.n4363 gnd.n2412 0.548625
R19180 gnd.n4051 gnd.n4050 0.532512
R19181 gnd.n4003 gnd.n4002 0.532512
R19182 gnd.n7110 gnd.n7109 0.532512
R19183 gnd.n7196 gnd.n78 0.532512
R19184 gnd.n5921 gnd.n5920 0.523366
R19185 gnd.n2852 gnd.n2645 0.523366
R19186 gnd.n7190 gnd.n7189 0.520317
R19187 gnd.n7119 gnd.n7118 0.520317
R19188 gnd.n3105 gnd.n2803 0.520317
R19189 gnd.n3029 gnd.n2674 0.520317
R19190 gnd.n3638 gnd.n2532 0.520317
R19191 gnd.n4546 gnd.n4545 0.520317
R19192 gnd.n4197 gnd.n4196 0.520317
R19193 gnd.n4099 gnd.n2325 0.520317
R19194 gnd.n5538 gnd.n5537 0.489829
R19195 gnd.n4519 gnd.n4518 0.489829
R19196 gnd.n1893 gnd.n938 0.486781
R19197 gnd.n1467 gnd.n1466 0.48678
R19198 gnd.n2210 gnd.n892 0.480683
R19199 gnd.n1551 gnd.n1550 0.480683
R19200 gnd.n7229 gnd.n7228 0.470187
R19201 gnd.n5923 gnd.n5922 0.432431
R19202 gnd.n2855 gnd.n2854 0.432431
R19203 gnd.n6231 gnd.n6230 0.425805
R19204 gnd.n6690 gnd.n423 0.425805
R19205 gnd.n6893 gnd.n297 0.425805
R19206 gnd.n6060 gnd.n6059 0.425805
R19207 gnd.n4526 gnd.n3731 0.388379
R19208 gnd.n2170 gnd.n2169 0.388379
R19209 gnd.n2138 gnd.n2137 0.388379
R19210 gnd.n2106 gnd.n2105 0.388379
R19211 gnd.n2075 gnd.n2074 0.388379
R19212 gnd.n2043 gnd.n2042 0.388379
R19213 gnd.n2011 gnd.n2010 0.388379
R19214 gnd.n1979 gnd.n1978 0.388379
R19215 gnd.n1948 gnd.n1947 0.388379
R19216 gnd.n7159 gnd.n7158 0.388379
R19217 gnd.n4143 gnd.n4084 0.388379
R19218 gnd.n5552 gnd.n5551 0.388379
R19219 gnd.n7229 gnd.n15 0.374463
R19220 gnd.n993 gnd.t29 0.319156
R19221 gnd.t12 gnd.n2398 0.319156
R19222 gnd.n4304 gnd.t20 0.319156
R19223 gnd.n4326 gnd.t220 0.319156
R19224 gnd.n4339 gnd.t246 0.319156
R19225 gnd.n4475 gnd.t116 0.319156
R19226 gnd.n4913 gnd.t14 0.319156
R19227 gnd.t252 gnd.t166 0.319156
R19228 gnd.t242 gnd.t2 0.319156
R19229 gnd.t155 gnd.n5139 0.319156
R19230 gnd.n5532 gnd.t93 0.319156
R19231 gnd.n5686 gnd.t164 0.319156
R19232 gnd.n5717 gnd.t259 0.319156
R19233 gnd.n6965 gnd.t209 0.319156
R19234 gnd.n6952 gnd.t173 0.319156
R19235 gnd.n1385 gnd.n1363 0.311721
R19236 gnd.n4537 gnd.n4536 0.302329
R19237 gnd.n5562 gnd.n5561 0.302329
R19238 gnd gnd.n7229 0.295112
R19239 gnd.n2281 gnd.n2280 0.268793
R19240 gnd.n2280 gnd.n2279 0.241354
R19241 gnd.n3068 gnd.n3067 0.229039
R19242 gnd.n3071 gnd.n3068 0.229039
R19243 gnd.n4585 gnd.n3622 0.229039
R19244 gnd.n4585 gnd.n4584 0.229039
R19245 gnd.n1539 gnd.n1338 0.206293
R19246 gnd.n2187 gnd.n2159 0.155672
R19247 gnd.n2180 gnd.n2159 0.155672
R19248 gnd.n2180 gnd.n2179 0.155672
R19249 gnd.n2179 gnd.n2163 0.155672
R19250 gnd.n2172 gnd.n2163 0.155672
R19251 gnd.n2172 gnd.n2171 0.155672
R19252 gnd.n2155 gnd.n2127 0.155672
R19253 gnd.n2148 gnd.n2127 0.155672
R19254 gnd.n2148 gnd.n2147 0.155672
R19255 gnd.n2147 gnd.n2131 0.155672
R19256 gnd.n2140 gnd.n2131 0.155672
R19257 gnd.n2140 gnd.n2139 0.155672
R19258 gnd.n2123 gnd.n2095 0.155672
R19259 gnd.n2116 gnd.n2095 0.155672
R19260 gnd.n2116 gnd.n2115 0.155672
R19261 gnd.n2115 gnd.n2099 0.155672
R19262 gnd.n2108 gnd.n2099 0.155672
R19263 gnd.n2108 gnd.n2107 0.155672
R19264 gnd.n2092 gnd.n2064 0.155672
R19265 gnd.n2085 gnd.n2064 0.155672
R19266 gnd.n2085 gnd.n2084 0.155672
R19267 gnd.n2084 gnd.n2068 0.155672
R19268 gnd.n2077 gnd.n2068 0.155672
R19269 gnd.n2077 gnd.n2076 0.155672
R19270 gnd.n2060 gnd.n2032 0.155672
R19271 gnd.n2053 gnd.n2032 0.155672
R19272 gnd.n2053 gnd.n2052 0.155672
R19273 gnd.n2052 gnd.n2036 0.155672
R19274 gnd.n2045 gnd.n2036 0.155672
R19275 gnd.n2045 gnd.n2044 0.155672
R19276 gnd.n2028 gnd.n2000 0.155672
R19277 gnd.n2021 gnd.n2000 0.155672
R19278 gnd.n2021 gnd.n2020 0.155672
R19279 gnd.n2020 gnd.n2004 0.155672
R19280 gnd.n2013 gnd.n2004 0.155672
R19281 gnd.n2013 gnd.n2012 0.155672
R19282 gnd.n1996 gnd.n1968 0.155672
R19283 gnd.n1989 gnd.n1968 0.155672
R19284 gnd.n1989 gnd.n1988 0.155672
R19285 gnd.n1988 gnd.n1972 0.155672
R19286 gnd.n1981 gnd.n1972 0.155672
R19287 gnd.n1981 gnd.n1980 0.155672
R19288 gnd.n1965 gnd.n1937 0.155672
R19289 gnd.n1958 gnd.n1937 0.155672
R19290 gnd.n1958 gnd.n1957 0.155672
R19291 gnd.n1957 gnd.n1941 0.155672
R19292 gnd.n1950 gnd.n1941 0.155672
R19293 gnd.n1950 gnd.n1949 0.155672
R19294 gnd.n2312 gnd.n892 0.152939
R19295 gnd.n2312 gnd.n2311 0.152939
R19296 gnd.n2311 gnd.n2310 0.152939
R19297 gnd.n2310 gnd.n894 0.152939
R19298 gnd.n895 gnd.n894 0.152939
R19299 gnd.n896 gnd.n895 0.152939
R19300 gnd.n897 gnd.n896 0.152939
R19301 gnd.n898 gnd.n897 0.152939
R19302 gnd.n899 gnd.n898 0.152939
R19303 gnd.n900 gnd.n899 0.152939
R19304 gnd.n901 gnd.n900 0.152939
R19305 gnd.n902 gnd.n901 0.152939
R19306 gnd.n903 gnd.n902 0.152939
R19307 gnd.n904 gnd.n903 0.152939
R19308 gnd.n2282 gnd.n904 0.152939
R19309 gnd.n2282 gnd.n2281 0.152939
R19310 gnd.n1552 gnd.n1551 0.152939
R19311 gnd.n1552 gnd.n1256 0.152939
R19312 gnd.n1580 gnd.n1256 0.152939
R19313 gnd.n1581 gnd.n1580 0.152939
R19314 gnd.n1582 gnd.n1581 0.152939
R19315 gnd.n1583 gnd.n1582 0.152939
R19316 gnd.n1583 gnd.n1228 0.152939
R19317 gnd.n1610 gnd.n1228 0.152939
R19318 gnd.n1611 gnd.n1610 0.152939
R19319 gnd.n1612 gnd.n1611 0.152939
R19320 gnd.n1612 gnd.n1206 0.152939
R19321 gnd.n1641 gnd.n1206 0.152939
R19322 gnd.n1642 gnd.n1641 0.152939
R19323 gnd.n1643 gnd.n1642 0.152939
R19324 gnd.n1644 gnd.n1643 0.152939
R19325 gnd.n1646 gnd.n1644 0.152939
R19326 gnd.n1646 gnd.n1645 0.152939
R19327 gnd.n1645 gnd.n1155 0.152939
R19328 gnd.n1156 gnd.n1155 0.152939
R19329 gnd.n1157 gnd.n1156 0.152939
R19330 gnd.n1176 gnd.n1157 0.152939
R19331 gnd.n1177 gnd.n1176 0.152939
R19332 gnd.n1177 gnd.n1087 0.152939
R19333 gnd.n1736 gnd.n1087 0.152939
R19334 gnd.n1737 gnd.n1736 0.152939
R19335 gnd.n1738 gnd.n1737 0.152939
R19336 gnd.n1739 gnd.n1738 0.152939
R19337 gnd.n1739 gnd.n1060 0.152939
R19338 gnd.n1776 gnd.n1060 0.152939
R19339 gnd.n1777 gnd.n1776 0.152939
R19340 gnd.n1778 gnd.n1777 0.152939
R19341 gnd.n1779 gnd.n1778 0.152939
R19342 gnd.n1779 gnd.n1034 0.152939
R19343 gnd.n1823 gnd.n1034 0.152939
R19344 gnd.n1824 gnd.n1823 0.152939
R19345 gnd.n1825 gnd.n1824 0.152939
R19346 gnd.n1826 gnd.n1825 0.152939
R19347 gnd.n1826 gnd.n1007 0.152939
R19348 gnd.n1863 gnd.n1007 0.152939
R19349 gnd.n1864 gnd.n1863 0.152939
R19350 gnd.n1865 gnd.n1864 0.152939
R19351 gnd.n1866 gnd.n1865 0.152939
R19352 gnd.n1866 gnd.n980 0.152939
R19353 gnd.n1912 gnd.n980 0.152939
R19354 gnd.n1913 gnd.n1912 0.152939
R19355 gnd.n1914 gnd.n1913 0.152939
R19356 gnd.n1915 gnd.n1914 0.152939
R19357 gnd.n1915 gnd.n953 0.152939
R19358 gnd.n2206 gnd.n953 0.152939
R19359 gnd.n2207 gnd.n2206 0.152939
R19360 gnd.n2208 gnd.n2207 0.152939
R19361 gnd.n2209 gnd.n2208 0.152939
R19362 gnd.n2210 gnd.n2209 0.152939
R19363 gnd.n1550 gnd.n1280 0.152939
R19364 gnd.n1301 gnd.n1280 0.152939
R19365 gnd.n1302 gnd.n1301 0.152939
R19366 gnd.n1308 gnd.n1302 0.152939
R19367 gnd.n1309 gnd.n1308 0.152939
R19368 gnd.n1310 gnd.n1309 0.152939
R19369 gnd.n1310 gnd.n1299 0.152939
R19370 gnd.n1318 gnd.n1299 0.152939
R19371 gnd.n1319 gnd.n1318 0.152939
R19372 gnd.n1320 gnd.n1319 0.152939
R19373 gnd.n1320 gnd.n1297 0.152939
R19374 gnd.n1328 gnd.n1297 0.152939
R19375 gnd.n1329 gnd.n1328 0.152939
R19376 gnd.n1330 gnd.n1329 0.152939
R19377 gnd.n1330 gnd.n1295 0.152939
R19378 gnd.n1338 gnd.n1295 0.152939
R19379 gnd.n2279 gnd.n909 0.152939
R19380 gnd.n911 gnd.n909 0.152939
R19381 gnd.n912 gnd.n911 0.152939
R19382 gnd.n913 gnd.n912 0.152939
R19383 gnd.n914 gnd.n913 0.152939
R19384 gnd.n915 gnd.n914 0.152939
R19385 gnd.n916 gnd.n915 0.152939
R19386 gnd.n917 gnd.n916 0.152939
R19387 gnd.n918 gnd.n917 0.152939
R19388 gnd.n919 gnd.n918 0.152939
R19389 gnd.n920 gnd.n919 0.152939
R19390 gnd.n921 gnd.n920 0.152939
R19391 gnd.n922 gnd.n921 0.152939
R19392 gnd.n923 gnd.n922 0.152939
R19393 gnd.n924 gnd.n923 0.152939
R19394 gnd.n925 gnd.n924 0.152939
R19395 gnd.n926 gnd.n925 0.152939
R19396 gnd.n927 gnd.n926 0.152939
R19397 gnd.n928 gnd.n927 0.152939
R19398 gnd.n929 gnd.n928 0.152939
R19399 gnd.n930 gnd.n929 0.152939
R19400 gnd.n931 gnd.n930 0.152939
R19401 gnd.n935 gnd.n931 0.152939
R19402 gnd.n936 gnd.n935 0.152939
R19403 gnd.n937 gnd.n936 0.152939
R19404 gnd.n938 gnd.n937 0.152939
R19405 gnd.n1713 gnd.n1712 0.152939
R19406 gnd.n1714 gnd.n1713 0.152939
R19407 gnd.n1715 gnd.n1714 0.152939
R19408 gnd.n1716 gnd.n1715 0.152939
R19409 gnd.n1717 gnd.n1716 0.152939
R19410 gnd.n1718 gnd.n1717 0.152939
R19411 gnd.n1718 gnd.n1041 0.152939
R19412 gnd.n1797 gnd.n1041 0.152939
R19413 gnd.n1798 gnd.n1797 0.152939
R19414 gnd.n1799 gnd.n1798 0.152939
R19415 gnd.n1800 gnd.n1799 0.152939
R19416 gnd.n1801 gnd.n1800 0.152939
R19417 gnd.n1802 gnd.n1801 0.152939
R19418 gnd.n1803 gnd.n1802 0.152939
R19419 gnd.n1804 gnd.n1803 0.152939
R19420 gnd.n1805 gnd.n1804 0.152939
R19421 gnd.n1805 gnd.n987 0.152939
R19422 gnd.n1884 gnd.n987 0.152939
R19423 gnd.n1885 gnd.n1884 0.152939
R19424 gnd.n1886 gnd.n1885 0.152939
R19425 gnd.n1887 gnd.n1886 0.152939
R19426 gnd.n1888 gnd.n1887 0.152939
R19427 gnd.n1889 gnd.n1888 0.152939
R19428 gnd.n1890 gnd.n1889 0.152939
R19429 gnd.n1891 gnd.n1890 0.152939
R19430 gnd.n1892 gnd.n1891 0.152939
R19431 gnd.n1894 gnd.n1892 0.152939
R19432 gnd.n1894 gnd.n1893 0.152939
R19433 gnd.n1468 gnd.n1467 0.152939
R19434 gnd.n1468 gnd.n1358 0.152939
R19435 gnd.n1483 gnd.n1358 0.152939
R19436 gnd.n1484 gnd.n1483 0.152939
R19437 gnd.n1485 gnd.n1484 0.152939
R19438 gnd.n1485 gnd.n1346 0.152939
R19439 gnd.n1499 gnd.n1346 0.152939
R19440 gnd.n1500 gnd.n1499 0.152939
R19441 gnd.n1501 gnd.n1500 0.152939
R19442 gnd.n1502 gnd.n1501 0.152939
R19443 gnd.n1503 gnd.n1502 0.152939
R19444 gnd.n1504 gnd.n1503 0.152939
R19445 gnd.n1505 gnd.n1504 0.152939
R19446 gnd.n1506 gnd.n1505 0.152939
R19447 gnd.n1507 gnd.n1506 0.152939
R19448 gnd.n1508 gnd.n1507 0.152939
R19449 gnd.n1509 gnd.n1508 0.152939
R19450 gnd.n1510 gnd.n1509 0.152939
R19451 gnd.n1511 gnd.n1510 0.152939
R19452 gnd.n1512 gnd.n1511 0.152939
R19453 gnd.n1513 gnd.n1512 0.152939
R19454 gnd.n1513 gnd.n1212 0.152939
R19455 gnd.n1630 gnd.n1212 0.152939
R19456 gnd.n1631 gnd.n1630 0.152939
R19457 gnd.n1632 gnd.n1631 0.152939
R19458 gnd.n1633 gnd.n1632 0.152939
R19459 gnd.n1633 gnd.n1134 0.152939
R19460 gnd.n1710 gnd.n1134 0.152939
R19461 gnd.n1386 gnd.n1385 0.152939
R19462 gnd.n1387 gnd.n1386 0.152939
R19463 gnd.n1388 gnd.n1387 0.152939
R19464 gnd.n1389 gnd.n1388 0.152939
R19465 gnd.n1390 gnd.n1389 0.152939
R19466 gnd.n1391 gnd.n1390 0.152939
R19467 gnd.n1392 gnd.n1391 0.152939
R19468 gnd.n1393 gnd.n1392 0.152939
R19469 gnd.n1394 gnd.n1393 0.152939
R19470 gnd.n1395 gnd.n1394 0.152939
R19471 gnd.n1396 gnd.n1395 0.152939
R19472 gnd.n1397 gnd.n1396 0.152939
R19473 gnd.n1398 gnd.n1397 0.152939
R19474 gnd.n1399 gnd.n1398 0.152939
R19475 gnd.n1400 gnd.n1399 0.152939
R19476 gnd.n1401 gnd.n1400 0.152939
R19477 gnd.n1402 gnd.n1401 0.152939
R19478 gnd.n1403 gnd.n1402 0.152939
R19479 gnd.n1404 gnd.n1403 0.152939
R19480 gnd.n1405 gnd.n1404 0.152939
R19481 gnd.n1406 gnd.n1405 0.152939
R19482 gnd.n1407 gnd.n1406 0.152939
R19483 gnd.n1411 gnd.n1407 0.152939
R19484 gnd.n1412 gnd.n1411 0.152939
R19485 gnd.n1412 gnd.n1369 0.152939
R19486 gnd.n1466 gnd.n1369 0.152939
R19487 gnd.n6231 gnd.n692 0.152939
R19488 gnd.n6239 gnd.n692 0.152939
R19489 gnd.n6240 gnd.n6239 0.152939
R19490 gnd.n6241 gnd.n6240 0.152939
R19491 gnd.n6241 gnd.n686 0.152939
R19492 gnd.n6249 gnd.n686 0.152939
R19493 gnd.n6250 gnd.n6249 0.152939
R19494 gnd.n6251 gnd.n6250 0.152939
R19495 gnd.n6251 gnd.n680 0.152939
R19496 gnd.n6259 gnd.n680 0.152939
R19497 gnd.n6260 gnd.n6259 0.152939
R19498 gnd.n6261 gnd.n6260 0.152939
R19499 gnd.n6261 gnd.n674 0.152939
R19500 gnd.n6269 gnd.n674 0.152939
R19501 gnd.n6270 gnd.n6269 0.152939
R19502 gnd.n6271 gnd.n6270 0.152939
R19503 gnd.n6271 gnd.n668 0.152939
R19504 gnd.n6279 gnd.n668 0.152939
R19505 gnd.n6280 gnd.n6279 0.152939
R19506 gnd.n6281 gnd.n6280 0.152939
R19507 gnd.n6281 gnd.n662 0.152939
R19508 gnd.n6289 gnd.n662 0.152939
R19509 gnd.n6290 gnd.n6289 0.152939
R19510 gnd.n6291 gnd.n6290 0.152939
R19511 gnd.n6291 gnd.n656 0.152939
R19512 gnd.n6299 gnd.n656 0.152939
R19513 gnd.n6300 gnd.n6299 0.152939
R19514 gnd.n6301 gnd.n6300 0.152939
R19515 gnd.n6301 gnd.n650 0.152939
R19516 gnd.n6309 gnd.n650 0.152939
R19517 gnd.n6310 gnd.n6309 0.152939
R19518 gnd.n6311 gnd.n6310 0.152939
R19519 gnd.n6311 gnd.n644 0.152939
R19520 gnd.n6319 gnd.n644 0.152939
R19521 gnd.n6320 gnd.n6319 0.152939
R19522 gnd.n6321 gnd.n6320 0.152939
R19523 gnd.n6321 gnd.n638 0.152939
R19524 gnd.n6329 gnd.n638 0.152939
R19525 gnd.n6330 gnd.n6329 0.152939
R19526 gnd.n6331 gnd.n6330 0.152939
R19527 gnd.n6331 gnd.n632 0.152939
R19528 gnd.n6339 gnd.n632 0.152939
R19529 gnd.n6340 gnd.n6339 0.152939
R19530 gnd.n6341 gnd.n6340 0.152939
R19531 gnd.n6341 gnd.n626 0.152939
R19532 gnd.n6349 gnd.n626 0.152939
R19533 gnd.n6350 gnd.n6349 0.152939
R19534 gnd.n6351 gnd.n6350 0.152939
R19535 gnd.n6351 gnd.n620 0.152939
R19536 gnd.n6359 gnd.n620 0.152939
R19537 gnd.n6360 gnd.n6359 0.152939
R19538 gnd.n6361 gnd.n6360 0.152939
R19539 gnd.n6361 gnd.n614 0.152939
R19540 gnd.n6369 gnd.n614 0.152939
R19541 gnd.n6370 gnd.n6369 0.152939
R19542 gnd.n6371 gnd.n6370 0.152939
R19543 gnd.n6371 gnd.n608 0.152939
R19544 gnd.n6379 gnd.n608 0.152939
R19545 gnd.n6380 gnd.n6379 0.152939
R19546 gnd.n6381 gnd.n6380 0.152939
R19547 gnd.n6381 gnd.n602 0.152939
R19548 gnd.n6389 gnd.n602 0.152939
R19549 gnd.n6390 gnd.n6389 0.152939
R19550 gnd.n6391 gnd.n6390 0.152939
R19551 gnd.n6391 gnd.n596 0.152939
R19552 gnd.n6399 gnd.n596 0.152939
R19553 gnd.n6400 gnd.n6399 0.152939
R19554 gnd.n6401 gnd.n6400 0.152939
R19555 gnd.n6401 gnd.n590 0.152939
R19556 gnd.n6409 gnd.n590 0.152939
R19557 gnd.n6410 gnd.n6409 0.152939
R19558 gnd.n6411 gnd.n6410 0.152939
R19559 gnd.n6411 gnd.n584 0.152939
R19560 gnd.n6419 gnd.n584 0.152939
R19561 gnd.n6420 gnd.n6419 0.152939
R19562 gnd.n6421 gnd.n6420 0.152939
R19563 gnd.n6421 gnd.n578 0.152939
R19564 gnd.n6429 gnd.n578 0.152939
R19565 gnd.n6430 gnd.n6429 0.152939
R19566 gnd.n6431 gnd.n6430 0.152939
R19567 gnd.n6431 gnd.n572 0.152939
R19568 gnd.n6439 gnd.n572 0.152939
R19569 gnd.n6440 gnd.n6439 0.152939
R19570 gnd.n6441 gnd.n6440 0.152939
R19571 gnd.n6441 gnd.n566 0.152939
R19572 gnd.n6449 gnd.n566 0.152939
R19573 gnd.n6450 gnd.n6449 0.152939
R19574 gnd.n6451 gnd.n6450 0.152939
R19575 gnd.n6451 gnd.n560 0.152939
R19576 gnd.n6459 gnd.n560 0.152939
R19577 gnd.n6460 gnd.n6459 0.152939
R19578 gnd.n6461 gnd.n6460 0.152939
R19579 gnd.n6461 gnd.n554 0.152939
R19580 gnd.n6469 gnd.n554 0.152939
R19581 gnd.n6470 gnd.n6469 0.152939
R19582 gnd.n6471 gnd.n6470 0.152939
R19583 gnd.n6471 gnd.n548 0.152939
R19584 gnd.n6479 gnd.n548 0.152939
R19585 gnd.n6480 gnd.n6479 0.152939
R19586 gnd.n6481 gnd.n6480 0.152939
R19587 gnd.n6481 gnd.n542 0.152939
R19588 gnd.n6489 gnd.n542 0.152939
R19589 gnd.n6490 gnd.n6489 0.152939
R19590 gnd.n6491 gnd.n6490 0.152939
R19591 gnd.n6491 gnd.n536 0.152939
R19592 gnd.n6499 gnd.n536 0.152939
R19593 gnd.n6500 gnd.n6499 0.152939
R19594 gnd.n6501 gnd.n6500 0.152939
R19595 gnd.n6501 gnd.n530 0.152939
R19596 gnd.n6509 gnd.n530 0.152939
R19597 gnd.n6510 gnd.n6509 0.152939
R19598 gnd.n6511 gnd.n6510 0.152939
R19599 gnd.n6511 gnd.n524 0.152939
R19600 gnd.n6519 gnd.n524 0.152939
R19601 gnd.n6520 gnd.n6519 0.152939
R19602 gnd.n6521 gnd.n6520 0.152939
R19603 gnd.n6521 gnd.n518 0.152939
R19604 gnd.n6529 gnd.n518 0.152939
R19605 gnd.n6530 gnd.n6529 0.152939
R19606 gnd.n6531 gnd.n6530 0.152939
R19607 gnd.n6531 gnd.n512 0.152939
R19608 gnd.n6539 gnd.n512 0.152939
R19609 gnd.n6540 gnd.n6539 0.152939
R19610 gnd.n6541 gnd.n6540 0.152939
R19611 gnd.n6541 gnd.n506 0.152939
R19612 gnd.n6549 gnd.n506 0.152939
R19613 gnd.n6550 gnd.n6549 0.152939
R19614 gnd.n6551 gnd.n6550 0.152939
R19615 gnd.n6551 gnd.n500 0.152939
R19616 gnd.n6559 gnd.n500 0.152939
R19617 gnd.n6560 gnd.n6559 0.152939
R19618 gnd.n6561 gnd.n6560 0.152939
R19619 gnd.n6561 gnd.n494 0.152939
R19620 gnd.n6569 gnd.n494 0.152939
R19621 gnd.n6570 gnd.n6569 0.152939
R19622 gnd.n6571 gnd.n6570 0.152939
R19623 gnd.n6571 gnd.n488 0.152939
R19624 gnd.n6579 gnd.n488 0.152939
R19625 gnd.n6580 gnd.n6579 0.152939
R19626 gnd.n6581 gnd.n6580 0.152939
R19627 gnd.n6581 gnd.n482 0.152939
R19628 gnd.n6589 gnd.n482 0.152939
R19629 gnd.n6590 gnd.n6589 0.152939
R19630 gnd.n6591 gnd.n6590 0.152939
R19631 gnd.n6591 gnd.n476 0.152939
R19632 gnd.n6599 gnd.n476 0.152939
R19633 gnd.n6600 gnd.n6599 0.152939
R19634 gnd.n6601 gnd.n6600 0.152939
R19635 gnd.n6601 gnd.n470 0.152939
R19636 gnd.n6609 gnd.n470 0.152939
R19637 gnd.n6610 gnd.n6609 0.152939
R19638 gnd.n6611 gnd.n6610 0.152939
R19639 gnd.n6611 gnd.n464 0.152939
R19640 gnd.n6619 gnd.n464 0.152939
R19641 gnd.n6620 gnd.n6619 0.152939
R19642 gnd.n6621 gnd.n6620 0.152939
R19643 gnd.n6621 gnd.n458 0.152939
R19644 gnd.n6629 gnd.n458 0.152939
R19645 gnd.n6630 gnd.n6629 0.152939
R19646 gnd.n6631 gnd.n6630 0.152939
R19647 gnd.n6631 gnd.n452 0.152939
R19648 gnd.n6639 gnd.n452 0.152939
R19649 gnd.n6640 gnd.n6639 0.152939
R19650 gnd.n6641 gnd.n6640 0.152939
R19651 gnd.n6641 gnd.n446 0.152939
R19652 gnd.n6649 gnd.n446 0.152939
R19653 gnd.n6650 gnd.n6649 0.152939
R19654 gnd.n6651 gnd.n6650 0.152939
R19655 gnd.n6651 gnd.n440 0.152939
R19656 gnd.n6659 gnd.n440 0.152939
R19657 gnd.n6660 gnd.n6659 0.152939
R19658 gnd.n6661 gnd.n6660 0.152939
R19659 gnd.n6661 gnd.n434 0.152939
R19660 gnd.n6669 gnd.n434 0.152939
R19661 gnd.n6670 gnd.n6669 0.152939
R19662 gnd.n6671 gnd.n6670 0.152939
R19663 gnd.n6671 gnd.n428 0.152939
R19664 gnd.n6679 gnd.n428 0.152939
R19665 gnd.n6680 gnd.n6679 0.152939
R19666 gnd.n6681 gnd.n6680 0.152939
R19667 gnd.n6681 gnd.n423 0.152939
R19668 gnd.n6691 gnd.n6690 0.152939
R19669 gnd.n6692 gnd.n6691 0.152939
R19670 gnd.n6692 gnd.n417 0.152939
R19671 gnd.n6700 gnd.n417 0.152939
R19672 gnd.n6701 gnd.n6700 0.152939
R19673 gnd.n6702 gnd.n6701 0.152939
R19674 gnd.n6702 gnd.n411 0.152939
R19675 gnd.n6710 gnd.n411 0.152939
R19676 gnd.n6711 gnd.n6710 0.152939
R19677 gnd.n6712 gnd.n6711 0.152939
R19678 gnd.n6712 gnd.n405 0.152939
R19679 gnd.n6720 gnd.n405 0.152939
R19680 gnd.n6721 gnd.n6720 0.152939
R19681 gnd.n6722 gnd.n6721 0.152939
R19682 gnd.n6722 gnd.n399 0.152939
R19683 gnd.n6730 gnd.n399 0.152939
R19684 gnd.n6731 gnd.n6730 0.152939
R19685 gnd.n6732 gnd.n6731 0.152939
R19686 gnd.n6732 gnd.n393 0.152939
R19687 gnd.n6740 gnd.n393 0.152939
R19688 gnd.n6741 gnd.n6740 0.152939
R19689 gnd.n6742 gnd.n6741 0.152939
R19690 gnd.n6742 gnd.n387 0.152939
R19691 gnd.n6750 gnd.n387 0.152939
R19692 gnd.n6751 gnd.n6750 0.152939
R19693 gnd.n6752 gnd.n6751 0.152939
R19694 gnd.n6752 gnd.n381 0.152939
R19695 gnd.n6760 gnd.n381 0.152939
R19696 gnd.n6761 gnd.n6760 0.152939
R19697 gnd.n6762 gnd.n6761 0.152939
R19698 gnd.n6762 gnd.n375 0.152939
R19699 gnd.n6770 gnd.n375 0.152939
R19700 gnd.n6771 gnd.n6770 0.152939
R19701 gnd.n6772 gnd.n6771 0.152939
R19702 gnd.n6772 gnd.n369 0.152939
R19703 gnd.n6780 gnd.n369 0.152939
R19704 gnd.n6781 gnd.n6780 0.152939
R19705 gnd.n6782 gnd.n6781 0.152939
R19706 gnd.n6782 gnd.n363 0.152939
R19707 gnd.n6790 gnd.n363 0.152939
R19708 gnd.n6791 gnd.n6790 0.152939
R19709 gnd.n6792 gnd.n6791 0.152939
R19710 gnd.n6792 gnd.n357 0.152939
R19711 gnd.n6800 gnd.n357 0.152939
R19712 gnd.n6801 gnd.n6800 0.152939
R19713 gnd.n6802 gnd.n6801 0.152939
R19714 gnd.n6802 gnd.n351 0.152939
R19715 gnd.n6810 gnd.n351 0.152939
R19716 gnd.n6811 gnd.n6810 0.152939
R19717 gnd.n6812 gnd.n6811 0.152939
R19718 gnd.n6812 gnd.n345 0.152939
R19719 gnd.n6820 gnd.n345 0.152939
R19720 gnd.n6821 gnd.n6820 0.152939
R19721 gnd.n6822 gnd.n6821 0.152939
R19722 gnd.n6822 gnd.n339 0.152939
R19723 gnd.n6830 gnd.n339 0.152939
R19724 gnd.n6831 gnd.n6830 0.152939
R19725 gnd.n6832 gnd.n6831 0.152939
R19726 gnd.n6832 gnd.n333 0.152939
R19727 gnd.n6840 gnd.n333 0.152939
R19728 gnd.n6841 gnd.n6840 0.152939
R19729 gnd.n6842 gnd.n6841 0.152939
R19730 gnd.n6842 gnd.n327 0.152939
R19731 gnd.n6850 gnd.n327 0.152939
R19732 gnd.n6851 gnd.n6850 0.152939
R19733 gnd.n6852 gnd.n6851 0.152939
R19734 gnd.n6852 gnd.n321 0.152939
R19735 gnd.n6860 gnd.n321 0.152939
R19736 gnd.n6861 gnd.n6860 0.152939
R19737 gnd.n6862 gnd.n6861 0.152939
R19738 gnd.n6862 gnd.n315 0.152939
R19739 gnd.n6870 gnd.n315 0.152939
R19740 gnd.n6871 gnd.n6870 0.152939
R19741 gnd.n6872 gnd.n6871 0.152939
R19742 gnd.n6872 gnd.n309 0.152939
R19743 gnd.n6880 gnd.n309 0.152939
R19744 gnd.n6881 gnd.n6880 0.152939
R19745 gnd.n6882 gnd.n6881 0.152939
R19746 gnd.n6882 gnd.n303 0.152939
R19747 gnd.n6890 gnd.n303 0.152939
R19748 gnd.n6891 gnd.n6890 0.152939
R19749 gnd.n6892 gnd.n6891 0.152939
R19750 gnd.n6894 gnd.n6892 0.152939
R19751 gnd.n6894 gnd.n6893 0.152939
R19752 gnd.n274 gnd.n260 0.152939
R19753 gnd.n275 gnd.n274 0.152939
R19754 gnd.n275 gnd.n273 0.152939
R19755 gnd.n281 gnd.n273 0.152939
R19756 gnd.n282 gnd.n281 0.152939
R19757 gnd.n283 gnd.n282 0.152939
R19758 gnd.n284 gnd.n283 0.152939
R19759 gnd.n285 gnd.n284 0.152939
R19760 gnd.n288 gnd.n285 0.152939
R19761 gnd.n289 gnd.n288 0.152939
R19762 gnd.n290 gnd.n289 0.152939
R19763 gnd.n291 gnd.n290 0.152939
R19764 gnd.n294 gnd.n291 0.152939
R19765 gnd.n295 gnd.n294 0.152939
R19766 gnd.n296 gnd.n295 0.152939
R19767 gnd.n297 gnd.n296 0.152939
R19768 gnd.n6986 gnd.n6985 0.152939
R19769 gnd.n6986 gnd.n208 0.152939
R19770 gnd.n7000 gnd.n208 0.152939
R19771 gnd.n7001 gnd.n7000 0.152939
R19772 gnd.n7002 gnd.n7001 0.152939
R19773 gnd.n7002 gnd.n192 0.152939
R19774 gnd.n7016 gnd.n192 0.152939
R19775 gnd.n7017 gnd.n7016 0.152939
R19776 gnd.n7018 gnd.n7017 0.152939
R19777 gnd.n7018 gnd.n176 0.152939
R19778 gnd.n7032 gnd.n176 0.152939
R19779 gnd.n7033 gnd.n7032 0.152939
R19780 gnd.n7034 gnd.n7033 0.152939
R19781 gnd.n7035 gnd.n7034 0.152939
R19782 gnd.n7035 gnd.n88 0.152939
R19783 gnd.n7190 gnd.n88 0.152939
R19784 gnd.n7189 gnd.n89 0.152939
R19785 gnd.n91 gnd.n89 0.152939
R19786 gnd.n96 gnd.n91 0.152939
R19787 gnd.n97 gnd.n96 0.152939
R19788 gnd.n98 gnd.n97 0.152939
R19789 gnd.n99 gnd.n98 0.152939
R19790 gnd.n103 gnd.n99 0.152939
R19791 gnd.n104 gnd.n103 0.152939
R19792 gnd.n105 gnd.n104 0.152939
R19793 gnd.n106 gnd.n105 0.152939
R19794 gnd.n110 gnd.n106 0.152939
R19795 gnd.n111 gnd.n110 0.152939
R19796 gnd.n112 gnd.n111 0.152939
R19797 gnd.n113 gnd.n112 0.152939
R19798 gnd.n117 gnd.n113 0.152939
R19799 gnd.n118 gnd.n117 0.152939
R19800 gnd.n119 gnd.n118 0.152939
R19801 gnd.n120 gnd.n119 0.152939
R19802 gnd.n124 gnd.n120 0.152939
R19803 gnd.n125 gnd.n124 0.152939
R19804 gnd.n126 gnd.n125 0.152939
R19805 gnd.n127 gnd.n126 0.152939
R19806 gnd.n131 gnd.n127 0.152939
R19807 gnd.n132 gnd.n131 0.152939
R19808 gnd.n133 gnd.n132 0.152939
R19809 gnd.n134 gnd.n133 0.152939
R19810 gnd.n138 gnd.n134 0.152939
R19811 gnd.n139 gnd.n138 0.152939
R19812 gnd.n140 gnd.n139 0.152939
R19813 gnd.n141 gnd.n140 0.152939
R19814 gnd.n145 gnd.n141 0.152939
R19815 gnd.n146 gnd.n145 0.152939
R19816 gnd.n147 gnd.n146 0.152939
R19817 gnd.n148 gnd.n147 0.152939
R19818 gnd.n152 gnd.n148 0.152939
R19819 gnd.n153 gnd.n152 0.152939
R19820 gnd.n7120 gnd.n153 0.152939
R19821 gnd.n7120 gnd.n7119 0.152939
R19822 gnd.n5569 gnd.n2803 0.152939
R19823 gnd.n5570 gnd.n5569 0.152939
R19824 gnd.n5571 gnd.n5570 0.152939
R19825 gnd.n5572 gnd.n5571 0.152939
R19826 gnd.n5573 gnd.n5572 0.152939
R19827 gnd.n5574 gnd.n5573 0.152939
R19828 gnd.n5575 gnd.n5574 0.152939
R19829 gnd.n5576 gnd.n5575 0.152939
R19830 gnd.n5577 gnd.n5576 0.152939
R19831 gnd.n5578 gnd.n5577 0.152939
R19832 gnd.n5579 gnd.n5578 0.152939
R19833 gnd.n5579 gnd.n2734 0.152939
R19834 gnd.n5681 gnd.n2734 0.152939
R19835 gnd.n5682 gnd.n5681 0.152939
R19836 gnd.n5683 gnd.n5682 0.152939
R19837 gnd.n5683 gnd.n2732 0.152939
R19838 gnd.n5689 gnd.n2732 0.152939
R19839 gnd.n5690 gnd.n5689 0.152939
R19840 gnd.n5691 gnd.n5690 0.152939
R19841 gnd.n5692 gnd.n5691 0.152939
R19842 gnd.n5693 gnd.n5692 0.152939
R19843 gnd.n5694 gnd.n5693 0.152939
R19844 gnd.n5695 gnd.n5694 0.152939
R19845 gnd.n5696 gnd.n5695 0.152939
R19846 gnd.n5697 gnd.n5696 0.152939
R19847 gnd.n5699 gnd.n5697 0.152939
R19848 gnd.n5699 gnd.n5698 0.152939
R19849 gnd.n5698 gnd.n264 0.152939
R19850 gnd.n265 gnd.n264 0.152939
R19851 gnd.n266 gnd.n265 0.152939
R19852 gnd.n267 gnd.n266 0.152939
R19853 gnd.n268 gnd.n267 0.152939
R19854 gnd.n6914 gnd.n268 0.152939
R19855 gnd.n6918 gnd.n6914 0.152939
R19856 gnd.n6919 gnd.n6918 0.152939
R19857 gnd.n6920 gnd.n6919 0.152939
R19858 gnd.n6921 gnd.n6920 0.152939
R19859 gnd.n6922 gnd.n6921 0.152939
R19860 gnd.n6924 gnd.n6922 0.152939
R19861 gnd.n6924 gnd.n6923 0.152939
R19862 gnd.n6923 gnd.n159 0.152939
R19863 gnd.n7118 gnd.n159 0.152939
R19864 gnd.n3034 gnd.n3029 0.152939
R19865 gnd.n3035 gnd.n3034 0.152939
R19866 gnd.n3036 gnd.n3035 0.152939
R19867 gnd.n3036 gnd.n3025 0.152939
R19868 gnd.n3044 gnd.n3025 0.152939
R19869 gnd.n3045 gnd.n3044 0.152939
R19870 gnd.n3046 gnd.n3045 0.152939
R19871 gnd.n3046 gnd.n3021 0.152939
R19872 gnd.n3054 gnd.n3021 0.152939
R19873 gnd.n3055 gnd.n3054 0.152939
R19874 gnd.n3057 gnd.n3055 0.152939
R19875 gnd.n3057 gnd.n3056 0.152939
R19876 gnd.n3056 gnd.n3014 0.152939
R19877 gnd.n3066 gnd.n3014 0.152939
R19878 gnd.n3067 gnd.n3066 0.152939
R19879 gnd.n3074 gnd.n3071 0.152939
R19880 gnd.n3075 gnd.n3074 0.152939
R19881 gnd.n3076 gnd.n3075 0.152939
R19882 gnd.n3077 gnd.n3076 0.152939
R19883 gnd.n3080 gnd.n3077 0.152939
R19884 gnd.n3081 gnd.n3080 0.152939
R19885 gnd.n3082 gnd.n3081 0.152939
R19886 gnd.n3083 gnd.n3082 0.152939
R19887 gnd.n3086 gnd.n3083 0.152939
R19888 gnd.n3087 gnd.n3086 0.152939
R19889 gnd.n3088 gnd.n3087 0.152939
R19890 gnd.n3089 gnd.n3088 0.152939
R19891 gnd.n3092 gnd.n3089 0.152939
R19892 gnd.n3093 gnd.n3092 0.152939
R19893 gnd.n3094 gnd.n3093 0.152939
R19894 gnd.n3095 gnd.n3094 0.152939
R19895 gnd.n3101 gnd.n3095 0.152939
R19896 gnd.n3107 gnd.n3101 0.152939
R19897 gnd.n3107 gnd.n3106 0.152939
R19898 gnd.n3106 gnd.n3105 0.152939
R19899 gnd.n2675 gnd.n2674 0.152939
R19900 gnd.n2676 gnd.n2675 0.152939
R19901 gnd.n2790 gnd.n2676 0.152939
R19902 gnd.n2791 gnd.n2790 0.152939
R19903 gnd.n2791 gnd.n2769 0.152939
R19904 gnd.n5618 gnd.n2769 0.152939
R19905 gnd.n5619 gnd.n5618 0.152939
R19906 gnd.n5620 gnd.n5619 0.152939
R19907 gnd.n5621 gnd.n5620 0.152939
R19908 gnd.n5621 gnd.n2744 0.152939
R19909 gnd.n5671 gnd.n2744 0.152939
R19910 gnd.n5672 gnd.n5671 0.152939
R19911 gnd.n5673 gnd.n5672 0.152939
R19912 gnd.n5674 gnd.n5673 0.152939
R19913 gnd.n5674 gnd.n224 0.152939
R19914 gnd.n6985 gnd.n224 0.152939
R19915 gnd.n4365 gnd.n4364 0.152939
R19916 gnd.n4366 gnd.n4365 0.152939
R19917 gnd.n4367 gnd.n4366 0.152939
R19918 gnd.n4370 gnd.n4367 0.152939
R19919 gnd.n4371 gnd.n4370 0.152939
R19920 gnd.n4372 gnd.n4371 0.152939
R19921 gnd.n4373 gnd.n4372 0.152939
R19922 gnd.n4375 gnd.n4373 0.152939
R19923 gnd.n4375 gnd.n4374 0.152939
R19924 gnd.n4374 gnd.n3901 0.152939
R19925 gnd.n4447 gnd.n3901 0.152939
R19926 gnd.n4448 gnd.n4447 0.152939
R19927 gnd.n4449 gnd.n4448 0.152939
R19928 gnd.n4449 gnd.n3897 0.152939
R19929 gnd.n4455 gnd.n3897 0.152939
R19930 gnd.n4456 gnd.n4455 0.152939
R19931 gnd.n4457 gnd.n4456 0.152939
R19932 gnd.n4457 gnd.n3893 0.152939
R19933 gnd.n4467 gnd.n3893 0.152939
R19934 gnd.n4468 gnd.n4467 0.152939
R19935 gnd.n4469 gnd.n4468 0.152939
R19936 gnd.n4469 gnd.n3755 0.152939
R19937 gnd.n4480 gnd.n3755 0.152939
R19938 gnd.n4481 gnd.n4480 0.152939
R19939 gnd.n4482 gnd.n4481 0.152939
R19940 gnd.n4482 gnd.n3749 0.152939
R19941 gnd.n4495 gnd.n3749 0.152939
R19942 gnd.n4496 gnd.n4495 0.152939
R19943 gnd.n4497 gnd.n4496 0.152939
R19944 gnd.n4498 gnd.n4497 0.152939
R19945 gnd.n4499 gnd.n4498 0.152939
R19946 gnd.n4499 gnd.n3477 0.152939
R19947 gnd.n4712 gnd.n3477 0.152939
R19948 gnd.n4713 gnd.n4712 0.152939
R19949 gnd.n4714 gnd.n4713 0.152939
R19950 gnd.n4714 gnd.n3457 0.152939
R19951 gnd.n4749 gnd.n3457 0.152939
R19952 gnd.n4750 gnd.n4749 0.152939
R19953 gnd.n4751 gnd.n4750 0.152939
R19954 gnd.n4751 gnd.n3431 0.152939
R19955 gnd.n4790 gnd.n3431 0.152939
R19956 gnd.n4791 gnd.n4790 0.152939
R19957 gnd.n4792 gnd.n4791 0.152939
R19958 gnd.n4792 gnd.n3415 0.152939
R19959 gnd.n4835 gnd.n3415 0.152939
R19960 gnd.n4836 gnd.n4835 0.152939
R19961 gnd.n4837 gnd.n4836 0.152939
R19962 gnd.n4838 gnd.n4837 0.152939
R19963 gnd.n4838 gnd.n3387 0.152939
R19964 gnd.n4907 gnd.n3387 0.152939
R19965 gnd.n4908 gnd.n4907 0.152939
R19966 gnd.n4909 gnd.n4908 0.152939
R19967 gnd.n4909 gnd.n3366 0.152939
R19968 gnd.n4934 gnd.n3366 0.152939
R19969 gnd.n4935 gnd.n4934 0.152939
R19970 gnd.n4936 gnd.n4935 0.152939
R19971 gnd.n4936 gnd.n3345 0.152939
R19972 gnd.n4967 gnd.n3345 0.152939
R19973 gnd.n4968 gnd.n4967 0.152939
R19974 gnd.n4969 gnd.n4968 0.152939
R19975 gnd.n4969 gnd.n3328 0.152939
R19976 gnd.n5012 gnd.n3328 0.152939
R19977 gnd.n5013 gnd.n5012 0.152939
R19978 gnd.n5014 gnd.n5013 0.152939
R19979 gnd.n5015 gnd.n5014 0.152939
R19980 gnd.n5015 gnd.n3299 0.152939
R19981 gnd.n5083 gnd.n3299 0.152939
R19982 gnd.n5084 gnd.n5083 0.152939
R19983 gnd.n5085 gnd.n5084 0.152939
R19984 gnd.n5085 gnd.n3279 0.152939
R19985 gnd.n5110 gnd.n3279 0.152939
R19986 gnd.n5111 gnd.n5110 0.152939
R19987 gnd.n5112 gnd.n5111 0.152939
R19988 gnd.n5112 gnd.n3257 0.152939
R19989 gnd.n5143 gnd.n3257 0.152939
R19990 gnd.n5144 gnd.n5143 0.152939
R19991 gnd.n5145 gnd.n5144 0.152939
R19992 gnd.n5145 gnd.n3240 0.152939
R19993 gnd.n5188 gnd.n3240 0.152939
R19994 gnd.n5189 gnd.n5188 0.152939
R19995 gnd.n5190 gnd.n5189 0.152939
R19996 gnd.n5191 gnd.n5190 0.152939
R19997 gnd.n5191 gnd.n3212 0.152939
R19998 gnd.n5236 gnd.n3212 0.152939
R19999 gnd.n5237 gnd.n5236 0.152939
R20000 gnd.n5238 gnd.n5237 0.152939
R20001 gnd.n5238 gnd.n3192 0.152939
R20002 gnd.n5279 gnd.n3192 0.152939
R20003 gnd.n5280 gnd.n5279 0.152939
R20004 gnd.n5281 gnd.n5280 0.152939
R20005 gnd.n5282 gnd.n5281 0.152939
R20006 gnd.n5282 gnd.n3163 0.152939
R20007 gnd.n5332 gnd.n3163 0.152939
R20008 gnd.n5333 gnd.n5332 0.152939
R20009 gnd.n5334 gnd.n5333 0.152939
R20010 gnd.n5334 gnd.n2974 0.152939
R20011 gnd.n5503 gnd.n2974 0.152939
R20012 gnd.n5504 gnd.n5503 0.152939
R20013 gnd.n5505 gnd.n5504 0.152939
R20014 gnd.n5505 gnd.n2962 0.152939
R20015 gnd.n5526 gnd.n2962 0.152939
R20016 gnd.n5527 gnd.n5526 0.152939
R20017 gnd.n5529 gnd.n5527 0.152939
R20018 gnd.n5529 gnd.n5528 0.152939
R20019 gnd.n5528 gnd.n2653 0.152939
R20020 gnd.n2654 gnd.n2653 0.152939
R20021 gnd.n2655 gnd.n2654 0.152939
R20022 gnd.n2661 gnd.n2655 0.152939
R20023 gnd.n2662 gnd.n2661 0.152939
R20024 gnd.n2663 gnd.n2662 0.152939
R20025 gnd.n2664 gnd.n2663 0.152939
R20026 gnd.n2784 gnd.n2664 0.152939
R20027 gnd.n2785 gnd.n2784 0.152939
R20028 gnd.n2786 gnd.n2785 0.152939
R20029 gnd.n2786 gnd.n2780 0.152939
R20030 gnd.n5607 gnd.n2780 0.152939
R20031 gnd.n5608 gnd.n5607 0.152939
R20032 gnd.n5609 gnd.n5608 0.152939
R20033 gnd.n5610 gnd.n5609 0.152939
R20034 gnd.n5610 gnd.n2753 0.152939
R20035 gnd.n5644 gnd.n2753 0.152939
R20036 gnd.n5645 gnd.n5644 0.152939
R20037 gnd.n5646 gnd.n5645 0.152939
R20038 gnd.n5647 gnd.n5646 0.152939
R20039 gnd.n5648 gnd.n5647 0.152939
R20040 gnd.n5651 gnd.n5648 0.152939
R20041 gnd.n5652 gnd.n5651 0.152939
R20042 gnd.n4052 gnd.n4051 0.152939
R20043 gnd.n4053 gnd.n4052 0.152939
R20044 gnd.n4054 gnd.n4053 0.152939
R20045 gnd.n4206 gnd.n4054 0.152939
R20046 gnd.n4207 gnd.n4206 0.152939
R20047 gnd.n4208 gnd.n4207 0.152939
R20048 gnd.n4209 gnd.n4208 0.152939
R20049 gnd.n4219 gnd.n4209 0.152939
R20050 gnd.n4220 gnd.n4219 0.152939
R20051 gnd.n4220 gnd.n3964 0.152939
R20052 gnd.n4281 gnd.n3964 0.152939
R20053 gnd.n4282 gnd.n4281 0.152939
R20054 gnd.n4283 gnd.n4282 0.152939
R20055 gnd.n4283 gnd.n3958 0.152939
R20056 gnd.n4298 gnd.n3958 0.152939
R20057 gnd.n4299 gnd.n4298 0.152939
R20058 gnd.n4301 gnd.n4299 0.152939
R20059 gnd.n4301 gnd.n4300 0.152939
R20060 gnd.n4300 gnd.n3944 0.152939
R20061 gnd.n3945 gnd.n3944 0.152939
R20062 gnd.n4003 gnd.n3998 0.152939
R20063 gnd.n4011 gnd.n3998 0.152939
R20064 gnd.n4012 gnd.n4011 0.152939
R20065 gnd.n4013 gnd.n4012 0.152939
R20066 gnd.n4013 gnd.n3994 0.152939
R20067 gnd.n4021 gnd.n3994 0.152939
R20068 gnd.n4022 gnd.n4021 0.152939
R20069 gnd.n4023 gnd.n4022 0.152939
R20070 gnd.n4023 gnd.n3990 0.152939
R20071 gnd.n4031 gnd.n3990 0.152939
R20072 gnd.n4032 gnd.n4031 0.152939
R20073 gnd.n4033 gnd.n4032 0.152939
R20074 gnd.n4033 gnd.n3986 0.152939
R20075 gnd.n4041 gnd.n3986 0.152939
R20076 gnd.n4042 gnd.n4041 0.152939
R20077 gnd.n4043 gnd.n4042 0.152939
R20078 gnd.n4043 gnd.n3980 0.152939
R20079 gnd.n4050 gnd.n3980 0.152939
R20080 gnd.n4002 gnd.n4000 0.152939
R20081 gnd.n4000 gnd.n2336 0.152939
R20082 gnd.n2337 gnd.n2336 0.152939
R20083 gnd.n2338 gnd.n2337 0.152939
R20084 gnd.n2357 gnd.n2338 0.152939
R20085 gnd.n2358 gnd.n2357 0.152939
R20086 gnd.n2359 gnd.n2358 0.152939
R20087 gnd.n2360 gnd.n2359 0.152939
R20088 gnd.n2379 gnd.n2360 0.152939
R20089 gnd.n2380 gnd.n2379 0.152939
R20090 gnd.n2381 gnd.n2380 0.152939
R20091 gnd.n2382 gnd.n2381 0.152939
R20092 gnd.n2400 gnd.n2382 0.152939
R20093 gnd.n2401 gnd.n2400 0.152939
R20094 gnd.n2402 gnd.n2401 0.152939
R20095 gnd.n2403 gnd.n2402 0.152939
R20096 gnd.n2420 gnd.n2403 0.152939
R20097 gnd.n2421 gnd.n2420 0.152939
R20098 gnd.n2422 gnd.n2421 0.152939
R20099 gnd.n2423 gnd.n2422 0.152939
R20100 gnd.n3953 gnd.n2423 0.152939
R20101 gnd.n3953 gnd.n2437 0.152939
R20102 gnd.n2438 gnd.n2437 0.152939
R20103 gnd.n2439 gnd.n2438 0.152939
R20104 gnd.n2455 gnd.n2439 0.152939
R20105 gnd.n2456 gnd.n2455 0.152939
R20106 gnd.n2457 gnd.n2456 0.152939
R20107 gnd.n2458 gnd.n2457 0.152939
R20108 gnd.n2475 gnd.n2458 0.152939
R20109 gnd.n2476 gnd.n2475 0.152939
R20110 gnd.n2477 gnd.n2476 0.152939
R20111 gnd.n2478 gnd.n2477 0.152939
R20112 gnd.n2497 gnd.n2478 0.152939
R20113 gnd.n2498 gnd.n2497 0.152939
R20114 gnd.n2499 gnd.n2498 0.152939
R20115 gnd.n2500 gnd.n2499 0.152939
R20116 gnd.n2518 gnd.n2500 0.152939
R20117 gnd.n2519 gnd.n2518 0.152939
R20118 gnd.n2520 gnd.n2519 0.152939
R20119 gnd.n2521 gnd.n2520 0.152939
R20120 gnd.n2539 gnd.n2521 0.152939
R20121 gnd.n5923 gnd.n2539 0.152939
R20122 gnd.n2465 gnd.n2412 0.152939
R20123 gnd.n2466 gnd.n2465 0.152939
R20124 gnd.n2467 gnd.n2466 0.152939
R20125 gnd.n2468 gnd.n2467 0.152939
R20126 gnd.n2486 gnd.n2468 0.152939
R20127 gnd.n2487 gnd.n2486 0.152939
R20128 gnd.n2488 gnd.n2487 0.152939
R20129 gnd.n2489 gnd.n2488 0.152939
R20130 gnd.n2507 gnd.n2489 0.152939
R20131 gnd.n2508 gnd.n2507 0.152939
R20132 gnd.n2509 gnd.n2508 0.152939
R20133 gnd.n2510 gnd.n2509 0.152939
R20134 gnd.n2529 gnd.n2510 0.152939
R20135 gnd.n2530 gnd.n2529 0.152939
R20136 gnd.n2531 gnd.n2530 0.152939
R20137 gnd.n2532 gnd.n2531 0.152939
R20138 gnd.n3639 gnd.n3638 0.152939
R20139 gnd.n3640 gnd.n3639 0.152939
R20140 gnd.n3641 gnd.n3640 0.152939
R20141 gnd.n3642 gnd.n3641 0.152939
R20142 gnd.n3643 gnd.n3642 0.152939
R20143 gnd.n3644 gnd.n3643 0.152939
R20144 gnd.n3645 gnd.n3644 0.152939
R20145 gnd.n3646 gnd.n3645 0.152939
R20146 gnd.n3647 gnd.n3646 0.152939
R20147 gnd.n3648 gnd.n3647 0.152939
R20148 gnd.n3649 gnd.n3648 0.152939
R20149 gnd.n3650 gnd.n3649 0.152939
R20150 gnd.n3651 gnd.n3650 0.152939
R20151 gnd.n3652 gnd.n3651 0.152939
R20152 gnd.n3652 gnd.n3622 0.152939
R20153 gnd.n4584 gnd.n4583 0.152939
R20154 gnd.n4583 gnd.n3623 0.152939
R20155 gnd.n3683 gnd.n3623 0.152939
R20156 gnd.n3684 gnd.n3683 0.152939
R20157 gnd.n3685 gnd.n3684 0.152939
R20158 gnd.n3686 gnd.n3685 0.152939
R20159 gnd.n3690 gnd.n3686 0.152939
R20160 gnd.n3691 gnd.n3690 0.152939
R20161 gnd.n3692 gnd.n3691 0.152939
R20162 gnd.n3693 gnd.n3692 0.152939
R20163 gnd.n3697 gnd.n3693 0.152939
R20164 gnd.n3698 gnd.n3697 0.152939
R20165 gnd.n3699 gnd.n3698 0.152939
R20166 gnd.n3700 gnd.n3699 0.152939
R20167 gnd.n3704 gnd.n3700 0.152939
R20168 gnd.n3705 gnd.n3704 0.152939
R20169 gnd.n3706 gnd.n3705 0.152939
R20170 gnd.n3707 gnd.n3706 0.152939
R20171 gnd.n3712 gnd.n3707 0.152939
R20172 gnd.n4546 gnd.n3712 0.152939
R20173 gnd.n4200 gnd.n4197 0.152939
R20174 gnd.n4201 gnd.n4200 0.152939
R20175 gnd.n4202 gnd.n4201 0.152939
R20176 gnd.n4203 gnd.n4202 0.152939
R20177 gnd.n4204 gnd.n4203 0.152939
R20178 gnd.n4211 gnd.n4204 0.152939
R20179 gnd.n4212 gnd.n4211 0.152939
R20180 gnd.n4213 gnd.n4212 0.152939
R20181 gnd.n4214 gnd.n4213 0.152939
R20182 gnd.n4215 gnd.n4214 0.152939
R20183 gnd.n4216 gnd.n4215 0.152939
R20184 gnd.n4216 gnd.n3961 0.152939
R20185 gnd.n4289 gnd.n3961 0.152939
R20186 gnd.n4290 gnd.n4289 0.152939
R20187 gnd.n4292 gnd.n4290 0.152939
R20188 gnd.n4292 gnd.n4291 0.152939
R20189 gnd.n4291 gnd.n3956 0.152939
R20190 gnd.n3956 gnd.n3954 0.152939
R20191 gnd.n4309 gnd.n3954 0.152939
R20192 gnd.n4310 gnd.n4309 0.152939
R20193 gnd.n4311 gnd.n4310 0.152939
R20194 gnd.n4311 gnd.n3951 0.152939
R20195 gnd.n4330 gnd.n3951 0.152939
R20196 gnd.n4331 gnd.n4330 0.152939
R20197 gnd.n4332 gnd.n4331 0.152939
R20198 gnd.n4333 gnd.n4332 0.152939
R20199 gnd.n4334 gnd.n4333 0.152939
R20200 gnd.n4334 gnd.n3921 0.152939
R20201 gnd.n4400 gnd.n3921 0.152939
R20202 gnd.n4401 gnd.n4400 0.152939
R20203 gnd.n4402 gnd.n4401 0.152939
R20204 gnd.n4402 gnd.n3914 0.152939
R20205 gnd.n4416 gnd.n3914 0.152939
R20206 gnd.n4417 gnd.n4416 0.152939
R20207 gnd.n4418 gnd.n4417 0.152939
R20208 gnd.n4418 gnd.n3912 0.152939
R20209 gnd.n4424 gnd.n3912 0.152939
R20210 gnd.n4425 gnd.n4424 0.152939
R20211 gnd.n4427 gnd.n4425 0.152939
R20212 gnd.n4427 gnd.n4426 0.152939
R20213 gnd.n4426 gnd.n3713 0.152939
R20214 gnd.n4545 gnd.n3713 0.152939
R20215 gnd.n4104 gnd.n4099 0.152939
R20216 gnd.n4105 gnd.n4104 0.152939
R20217 gnd.n4106 gnd.n4105 0.152939
R20218 gnd.n4106 gnd.n4095 0.152939
R20219 gnd.n4114 gnd.n4095 0.152939
R20220 gnd.n4115 gnd.n4114 0.152939
R20221 gnd.n4116 gnd.n4115 0.152939
R20222 gnd.n4116 gnd.n4091 0.152939
R20223 gnd.n4124 gnd.n4091 0.152939
R20224 gnd.n4125 gnd.n4124 0.152939
R20225 gnd.n4126 gnd.n4125 0.152939
R20226 gnd.n4126 gnd.n4087 0.152939
R20227 gnd.n4134 gnd.n4087 0.152939
R20228 gnd.n4135 gnd.n4134 0.152939
R20229 gnd.n4136 gnd.n4135 0.152939
R20230 gnd.n4136 gnd.n4080 0.152939
R20231 gnd.n4144 gnd.n4080 0.152939
R20232 gnd.n4145 gnd.n4144 0.152939
R20233 gnd.n4146 gnd.n4145 0.152939
R20234 gnd.n4146 gnd.n4076 0.152939
R20235 gnd.n4154 gnd.n4076 0.152939
R20236 gnd.n4155 gnd.n4154 0.152939
R20237 gnd.n4156 gnd.n4155 0.152939
R20238 gnd.n4156 gnd.n4072 0.152939
R20239 gnd.n4164 gnd.n4072 0.152939
R20240 gnd.n4165 gnd.n4164 0.152939
R20241 gnd.n4166 gnd.n4165 0.152939
R20242 gnd.n4166 gnd.n4068 0.152939
R20243 gnd.n4174 gnd.n4068 0.152939
R20244 gnd.n4175 gnd.n4174 0.152939
R20245 gnd.n4176 gnd.n4175 0.152939
R20246 gnd.n4176 gnd.n4064 0.152939
R20247 gnd.n4184 gnd.n4064 0.152939
R20248 gnd.n4185 gnd.n4184 0.152939
R20249 gnd.n4187 gnd.n4185 0.152939
R20250 gnd.n4187 gnd.n4186 0.152939
R20251 gnd.n4186 gnd.n4057 0.152939
R20252 gnd.n4196 gnd.n4057 0.152939
R20253 gnd.n2326 gnd.n2325 0.152939
R20254 gnd.n2327 gnd.n2326 0.152939
R20255 gnd.n2346 gnd.n2327 0.152939
R20256 gnd.n2347 gnd.n2346 0.152939
R20257 gnd.n2348 gnd.n2347 0.152939
R20258 gnd.n2349 gnd.n2348 0.152939
R20259 gnd.n2368 gnd.n2349 0.152939
R20260 gnd.n2369 gnd.n2368 0.152939
R20261 gnd.n2370 gnd.n2369 0.152939
R20262 gnd.n2371 gnd.n2370 0.152939
R20263 gnd.n2389 gnd.n2371 0.152939
R20264 gnd.n2390 gnd.n2389 0.152939
R20265 gnd.n2391 gnd.n2390 0.152939
R20266 gnd.n2392 gnd.n2391 0.152939
R20267 gnd.n2411 gnd.n2392 0.152939
R20268 gnd.n2412 gnd.n2411 0.152939
R20269 gnd.n6059 gnd.n864 0.152939
R20270 gnd.n4251 gnd.n864 0.152939
R20271 gnd.n4252 gnd.n4251 0.152939
R20272 gnd.n4253 gnd.n4252 0.152939
R20273 gnd.n4253 gnd.n3974 0.152939
R20274 gnd.n4259 gnd.n3974 0.152939
R20275 gnd.n4260 gnd.n4259 0.152939
R20276 gnd.n4261 gnd.n4260 0.152939
R20277 gnd.n4261 gnd.n3970 0.152939
R20278 gnd.n4267 gnd.n3970 0.152939
R20279 gnd.n4268 gnd.n4267 0.152939
R20280 gnd.n4269 gnd.n4268 0.152939
R20281 gnd.n4270 gnd.n4269 0.152939
R20282 gnd.n4271 gnd.n4270 0.152939
R20283 gnd.n4271 gnd.n3935 0.152939
R20284 gnd.n4362 gnd.n3935 0.152939
R20285 gnd.n6230 gnd.n697 0.152939
R20286 gnd.n702 gnd.n697 0.152939
R20287 gnd.n703 gnd.n702 0.152939
R20288 gnd.n704 gnd.n703 0.152939
R20289 gnd.n705 gnd.n704 0.152939
R20290 gnd.n710 gnd.n705 0.152939
R20291 gnd.n711 gnd.n710 0.152939
R20292 gnd.n712 gnd.n711 0.152939
R20293 gnd.n713 gnd.n712 0.152939
R20294 gnd.n718 gnd.n713 0.152939
R20295 gnd.n719 gnd.n718 0.152939
R20296 gnd.n720 gnd.n719 0.152939
R20297 gnd.n721 gnd.n720 0.152939
R20298 gnd.n726 gnd.n721 0.152939
R20299 gnd.n727 gnd.n726 0.152939
R20300 gnd.n728 gnd.n727 0.152939
R20301 gnd.n729 gnd.n728 0.152939
R20302 gnd.n734 gnd.n729 0.152939
R20303 gnd.n735 gnd.n734 0.152939
R20304 gnd.n736 gnd.n735 0.152939
R20305 gnd.n737 gnd.n736 0.152939
R20306 gnd.n742 gnd.n737 0.152939
R20307 gnd.n743 gnd.n742 0.152939
R20308 gnd.n744 gnd.n743 0.152939
R20309 gnd.n745 gnd.n744 0.152939
R20310 gnd.n750 gnd.n745 0.152939
R20311 gnd.n751 gnd.n750 0.152939
R20312 gnd.n752 gnd.n751 0.152939
R20313 gnd.n753 gnd.n752 0.152939
R20314 gnd.n758 gnd.n753 0.152939
R20315 gnd.n759 gnd.n758 0.152939
R20316 gnd.n760 gnd.n759 0.152939
R20317 gnd.n761 gnd.n760 0.152939
R20318 gnd.n766 gnd.n761 0.152939
R20319 gnd.n767 gnd.n766 0.152939
R20320 gnd.n768 gnd.n767 0.152939
R20321 gnd.n769 gnd.n768 0.152939
R20322 gnd.n774 gnd.n769 0.152939
R20323 gnd.n775 gnd.n774 0.152939
R20324 gnd.n776 gnd.n775 0.152939
R20325 gnd.n777 gnd.n776 0.152939
R20326 gnd.n782 gnd.n777 0.152939
R20327 gnd.n783 gnd.n782 0.152939
R20328 gnd.n784 gnd.n783 0.152939
R20329 gnd.n785 gnd.n784 0.152939
R20330 gnd.n790 gnd.n785 0.152939
R20331 gnd.n791 gnd.n790 0.152939
R20332 gnd.n792 gnd.n791 0.152939
R20333 gnd.n793 gnd.n792 0.152939
R20334 gnd.n798 gnd.n793 0.152939
R20335 gnd.n799 gnd.n798 0.152939
R20336 gnd.n800 gnd.n799 0.152939
R20337 gnd.n801 gnd.n800 0.152939
R20338 gnd.n806 gnd.n801 0.152939
R20339 gnd.n807 gnd.n806 0.152939
R20340 gnd.n808 gnd.n807 0.152939
R20341 gnd.n809 gnd.n808 0.152939
R20342 gnd.n814 gnd.n809 0.152939
R20343 gnd.n815 gnd.n814 0.152939
R20344 gnd.n816 gnd.n815 0.152939
R20345 gnd.n817 gnd.n816 0.152939
R20346 gnd.n822 gnd.n817 0.152939
R20347 gnd.n823 gnd.n822 0.152939
R20348 gnd.n824 gnd.n823 0.152939
R20349 gnd.n825 gnd.n824 0.152939
R20350 gnd.n830 gnd.n825 0.152939
R20351 gnd.n831 gnd.n830 0.152939
R20352 gnd.n832 gnd.n831 0.152939
R20353 gnd.n833 gnd.n832 0.152939
R20354 gnd.n838 gnd.n833 0.152939
R20355 gnd.n839 gnd.n838 0.152939
R20356 gnd.n840 gnd.n839 0.152939
R20357 gnd.n841 gnd.n840 0.152939
R20358 gnd.n846 gnd.n841 0.152939
R20359 gnd.n847 gnd.n846 0.152939
R20360 gnd.n848 gnd.n847 0.152939
R20361 gnd.n849 gnd.n848 0.152939
R20362 gnd.n854 gnd.n849 0.152939
R20363 gnd.n855 gnd.n854 0.152939
R20364 gnd.n856 gnd.n855 0.152939
R20365 gnd.n857 gnd.n856 0.152939
R20366 gnd.n862 gnd.n857 0.152939
R20367 gnd.n863 gnd.n862 0.152939
R20368 gnd.n6060 gnd.n863 0.152939
R20369 gnd.n5560 gnd.n2807 0.152939
R20370 gnd.n5556 gnd.n2807 0.152939
R20371 gnd.n5556 gnd.n5555 0.152939
R20372 gnd.n5555 gnd.n5554 0.152939
R20373 gnd.n5554 gnd.n2949 0.152939
R20374 gnd.n5547 gnd.n2949 0.152939
R20375 gnd.n5547 gnd.n5546 0.152939
R20376 gnd.n5546 gnd.n5545 0.152939
R20377 gnd.n5545 gnd.n5538 0.152939
R20378 gnd.n4518 gnd.n3737 0.152939
R20379 gnd.n4514 gnd.n3737 0.152939
R20380 gnd.n4514 gnd.n4513 0.152939
R20381 gnd.n4513 gnd.n4512 0.152939
R20382 gnd.n4512 gnd.n3742 0.152939
R20383 gnd.n4508 gnd.n3742 0.152939
R20384 gnd.n4508 gnd.n3491 0.152939
R20385 gnd.n4680 gnd.n3491 0.152939
R20386 gnd.n4681 gnd.n4680 0.152939
R20387 gnd.n4696 gnd.n4681 0.152939
R20388 gnd.n4696 gnd.n4695 0.152939
R20389 gnd.n4695 gnd.n4694 0.152939
R20390 gnd.n4694 gnd.n4682 0.152939
R20391 gnd.n4690 gnd.n4682 0.152939
R20392 gnd.n4690 gnd.n4689 0.152939
R20393 gnd.n4689 gnd.n4688 0.152939
R20394 gnd.n4688 gnd.n3445 0.152939
R20395 gnd.n4767 gnd.n3445 0.152939
R20396 gnd.n4768 gnd.n4767 0.152939
R20397 gnd.n4776 gnd.n4768 0.152939
R20398 gnd.n4776 gnd.n4775 0.152939
R20399 gnd.n4775 gnd.n4774 0.152939
R20400 gnd.n4774 gnd.n4769 0.152939
R20401 gnd.n4769 gnd.n3402 0.152939
R20402 gnd.n4853 gnd.n3402 0.152939
R20403 gnd.n4854 gnd.n4853 0.152939
R20404 gnd.n4891 gnd.n4854 0.152939
R20405 gnd.n4891 gnd.n4890 0.152939
R20406 gnd.n4890 gnd.n4889 0.152939
R20407 gnd.n4889 gnd.n4855 0.152939
R20408 gnd.n4885 gnd.n4855 0.152939
R20409 gnd.n4885 gnd.n4884 0.152939
R20410 gnd.n4884 gnd.n4883 0.152939
R20411 gnd.n4883 gnd.n4860 0.152939
R20412 gnd.n4879 gnd.n4860 0.152939
R20413 gnd.n4879 gnd.n4878 0.152939
R20414 gnd.n4878 gnd.n4877 0.152939
R20415 gnd.n4877 gnd.n4865 0.152939
R20416 gnd.n4873 gnd.n4865 0.152939
R20417 gnd.n4873 gnd.n4872 0.152939
R20418 gnd.n4872 gnd.n3314 0.152939
R20419 gnd.n5030 gnd.n3314 0.152939
R20420 gnd.n5031 gnd.n5030 0.152939
R20421 gnd.n5068 gnd.n5031 0.152939
R20422 gnd.n5068 gnd.n5067 0.152939
R20423 gnd.n5067 gnd.n5066 0.152939
R20424 gnd.n5066 gnd.n5032 0.152939
R20425 gnd.n5062 gnd.n5032 0.152939
R20426 gnd.n5062 gnd.n5061 0.152939
R20427 gnd.n5061 gnd.n5060 0.152939
R20428 gnd.n5060 gnd.n5038 0.152939
R20429 gnd.n5056 gnd.n5038 0.152939
R20430 gnd.n5056 gnd.n5055 0.152939
R20431 gnd.n5055 gnd.n5054 0.152939
R20432 gnd.n5054 gnd.n5042 0.152939
R20433 gnd.n5050 gnd.n5042 0.152939
R20434 gnd.n5050 gnd.n5049 0.152939
R20435 gnd.n5049 gnd.n3226 0.152939
R20436 gnd.n5207 gnd.n3226 0.152939
R20437 gnd.n5208 gnd.n5207 0.152939
R20438 gnd.n5221 gnd.n5208 0.152939
R20439 gnd.n5221 gnd.n5220 0.152939
R20440 gnd.n5220 gnd.n5219 0.152939
R20441 gnd.n5219 gnd.n5209 0.152939
R20442 gnd.n5215 gnd.n5209 0.152939
R20443 gnd.n5215 gnd.n5214 0.152939
R20444 gnd.n5214 gnd.n3179 0.152939
R20445 gnd.n5299 gnd.n3179 0.152939
R20446 gnd.n5300 gnd.n5299 0.152939
R20447 gnd.n5318 gnd.n5300 0.152939
R20448 gnd.n5318 gnd.n5317 0.152939
R20449 gnd.n5317 gnd.n5316 0.152939
R20450 gnd.n5316 gnd.n5301 0.152939
R20451 gnd.n5312 gnd.n5301 0.152939
R20452 gnd.n5312 gnd.n5311 0.152939
R20453 gnd.n5311 gnd.n2968 0.152939
R20454 gnd.n5513 gnd.n2968 0.152939
R20455 gnd.n5514 gnd.n5513 0.152939
R20456 gnd.n5516 gnd.n5514 0.152939
R20457 gnd.n5516 gnd.n5515 0.152939
R20458 gnd.n5515 gnd.n2957 0.152939
R20459 gnd.n5537 gnd.n2957 0.152939
R20460 gnd.n4531 gnd.n3718 0.152939
R20461 gnd.n4531 gnd.n4530 0.152939
R20462 gnd.n4530 gnd.n4529 0.152939
R20463 gnd.n4529 gnd.n3725 0.152939
R20464 gnd.n4525 gnd.n3725 0.152939
R20465 gnd.n4525 gnd.n4524 0.152939
R20466 gnd.n4524 gnd.n3732 0.152939
R20467 gnd.n4520 gnd.n3732 0.152939
R20468 gnd.n4520 gnd.n4519 0.152939
R20469 gnd.n4346 gnd.n4345 0.152939
R20470 gnd.n4345 gnd.n3948 0.152939
R20471 gnd.n4341 gnd.n3948 0.152939
R20472 gnd.n4341 gnd.n3924 0.152939
R20473 gnd.n4392 gnd.n3924 0.152939
R20474 gnd.n4393 gnd.n4392 0.152939
R20475 gnd.n4394 gnd.n4393 0.152939
R20476 gnd.n4394 gnd.n3917 0.152939
R20477 gnd.n4408 gnd.n3917 0.152939
R20478 gnd.n4409 gnd.n4408 0.152939
R20479 gnd.n4410 gnd.n4409 0.152939
R20480 gnd.n4410 gnd.n3908 0.152939
R20481 gnd.n4438 gnd.n3908 0.152939
R20482 gnd.n4438 gnd.n4437 0.152939
R20483 gnd.n4437 gnd.n4436 0.152939
R20484 gnd.n4436 gnd.n3909 0.152939
R20485 gnd.n4432 gnd.n3909 0.152939
R20486 gnd.n4432 gnd.n3717 0.152939
R20487 gnd.n4538 gnd.n3717 0.152939
R20488 gnd.n4538 gnd.n4537 0.152939
R20489 gnd.n5920 gnd.n2542 0.152939
R20490 gnd.n5916 gnd.n2542 0.152939
R20491 gnd.n5916 gnd.n5915 0.152939
R20492 gnd.n5915 gnd.n5914 0.152939
R20493 gnd.n5914 gnd.n2547 0.152939
R20494 gnd.n5910 gnd.n2547 0.152939
R20495 gnd.n5910 gnd.n5909 0.152939
R20496 gnd.n5909 gnd.n5908 0.152939
R20497 gnd.n5908 gnd.n2552 0.152939
R20498 gnd.n5904 gnd.n2552 0.152939
R20499 gnd.n5904 gnd.n5903 0.152939
R20500 gnd.n5903 gnd.n5902 0.152939
R20501 gnd.n5902 gnd.n2557 0.152939
R20502 gnd.n5898 gnd.n2557 0.152939
R20503 gnd.n5898 gnd.n5897 0.152939
R20504 gnd.n5897 gnd.n5896 0.152939
R20505 gnd.n5896 gnd.n2562 0.152939
R20506 gnd.n5892 gnd.n2562 0.152939
R20507 gnd.n5892 gnd.n5891 0.152939
R20508 gnd.n5891 gnd.n5890 0.152939
R20509 gnd.n5890 gnd.n2567 0.152939
R20510 gnd.n5886 gnd.n2567 0.152939
R20511 gnd.n5886 gnd.n5885 0.152939
R20512 gnd.n5885 gnd.n5884 0.152939
R20513 gnd.n5884 gnd.n2572 0.152939
R20514 gnd.n5880 gnd.n2572 0.152939
R20515 gnd.n5880 gnd.n5879 0.152939
R20516 gnd.n5879 gnd.n5878 0.152939
R20517 gnd.n5878 gnd.n2577 0.152939
R20518 gnd.n5874 gnd.n2577 0.152939
R20519 gnd.n5874 gnd.n5873 0.152939
R20520 gnd.n5873 gnd.n5872 0.152939
R20521 gnd.n5872 gnd.n2582 0.152939
R20522 gnd.n5868 gnd.n2582 0.152939
R20523 gnd.n5868 gnd.n5867 0.152939
R20524 gnd.n5867 gnd.n5866 0.152939
R20525 gnd.n5866 gnd.n2587 0.152939
R20526 gnd.n5862 gnd.n2587 0.152939
R20527 gnd.n5862 gnd.n5861 0.152939
R20528 gnd.n5861 gnd.n5860 0.152939
R20529 gnd.n5860 gnd.n2592 0.152939
R20530 gnd.n5856 gnd.n2592 0.152939
R20531 gnd.n5856 gnd.n5855 0.152939
R20532 gnd.n5855 gnd.n5854 0.152939
R20533 gnd.n5854 gnd.n2597 0.152939
R20534 gnd.n5850 gnd.n2597 0.152939
R20535 gnd.n5850 gnd.n5849 0.152939
R20536 gnd.n5849 gnd.n5848 0.152939
R20537 gnd.n5848 gnd.n2602 0.152939
R20538 gnd.n5844 gnd.n2602 0.152939
R20539 gnd.n5844 gnd.n5843 0.152939
R20540 gnd.n5843 gnd.n5842 0.152939
R20541 gnd.n5842 gnd.n2607 0.152939
R20542 gnd.n5838 gnd.n2607 0.152939
R20543 gnd.n5838 gnd.n5837 0.152939
R20544 gnd.n5837 gnd.n5836 0.152939
R20545 gnd.n5836 gnd.n2612 0.152939
R20546 gnd.n5832 gnd.n2612 0.152939
R20547 gnd.n5832 gnd.n5831 0.152939
R20548 gnd.n5831 gnd.n5830 0.152939
R20549 gnd.n5830 gnd.n2617 0.152939
R20550 gnd.n5826 gnd.n2617 0.152939
R20551 gnd.n5826 gnd.n5825 0.152939
R20552 gnd.n5825 gnd.n5824 0.152939
R20553 gnd.n5824 gnd.n2622 0.152939
R20554 gnd.n5820 gnd.n2622 0.152939
R20555 gnd.n5820 gnd.n5819 0.152939
R20556 gnd.n5819 gnd.n5818 0.152939
R20557 gnd.n5818 gnd.n2627 0.152939
R20558 gnd.n5814 gnd.n2627 0.152939
R20559 gnd.n5814 gnd.n5813 0.152939
R20560 gnd.n5813 gnd.n5812 0.152939
R20561 gnd.n5812 gnd.n2632 0.152939
R20562 gnd.n5808 gnd.n2632 0.152939
R20563 gnd.n5808 gnd.n5807 0.152939
R20564 gnd.n5807 gnd.n5806 0.152939
R20565 gnd.n5806 gnd.n2637 0.152939
R20566 gnd.n5802 gnd.n2637 0.152939
R20567 gnd.n5802 gnd.n5801 0.152939
R20568 gnd.n5801 gnd.n5800 0.152939
R20569 gnd.n5800 gnd.n2642 0.152939
R20570 gnd.n2645 gnd.n2642 0.152939
R20571 gnd.n2854 gnd.n2687 0.152939
R20572 gnd.n5770 gnd.n2687 0.152939
R20573 gnd.n5770 gnd.n5769 0.152939
R20574 gnd.n5769 gnd.n5768 0.152939
R20575 gnd.n5768 gnd.n2688 0.152939
R20576 gnd.n5764 gnd.n2688 0.152939
R20577 gnd.n5764 gnd.n5763 0.152939
R20578 gnd.n5763 gnd.n5762 0.152939
R20579 gnd.n5762 gnd.n2693 0.152939
R20580 gnd.n5758 gnd.n2693 0.152939
R20581 gnd.n5758 gnd.n5757 0.152939
R20582 gnd.n5757 gnd.n5756 0.152939
R20583 gnd.n5756 gnd.n2698 0.152939
R20584 gnd.n5752 gnd.n2698 0.152939
R20585 gnd.n5752 gnd.n5751 0.152939
R20586 gnd.n5751 gnd.n5750 0.152939
R20587 gnd.n5750 gnd.n241 0.152939
R20588 gnd.n6977 gnd.n241 0.152939
R20589 gnd.n6977 gnd.n6976 0.152939
R20590 gnd.n6976 gnd.n6975 0.152939
R20591 gnd.n6975 gnd.n242 0.152939
R20592 gnd.n6971 gnd.n242 0.152939
R20593 gnd.n6971 gnd.n6970 0.152939
R20594 gnd.n6970 gnd.n6969 0.152939
R20595 gnd.n6969 gnd.n247 0.152939
R20596 gnd.n247 gnd.n217 0.152939
R20597 gnd.n6992 gnd.n217 0.152939
R20598 gnd.n6993 gnd.n6992 0.152939
R20599 gnd.n6994 gnd.n6993 0.152939
R20600 gnd.n6994 gnd.n200 0.152939
R20601 gnd.n7008 gnd.n200 0.152939
R20602 gnd.n7009 gnd.n7008 0.152939
R20603 gnd.n7010 gnd.n7009 0.152939
R20604 gnd.n7010 gnd.n185 0.152939
R20605 gnd.n7024 gnd.n185 0.152939
R20606 gnd.n7025 gnd.n7024 0.152939
R20607 gnd.n7026 gnd.n7025 0.152939
R20608 gnd.n7026 gnd.n166 0.152939
R20609 gnd.n7042 gnd.n166 0.152939
R20610 gnd.n7043 gnd.n7042 0.152939
R20611 gnd.n7111 gnd.n7043 0.152939
R20612 gnd.n7111 gnd.n7110 0.152939
R20613 gnd.n7109 gnd.n7044 0.152939
R20614 gnd.n7105 gnd.n7044 0.152939
R20615 gnd.n7105 gnd.n7104 0.152939
R20616 gnd.n7104 gnd.n7103 0.152939
R20617 gnd.n7103 gnd.n7050 0.152939
R20618 gnd.n7099 gnd.n7050 0.152939
R20619 gnd.n7099 gnd.n7098 0.152939
R20620 gnd.n7098 gnd.n7097 0.152939
R20621 gnd.n7097 gnd.n7058 0.152939
R20622 gnd.n7093 gnd.n7058 0.152939
R20623 gnd.n7093 gnd.n7092 0.152939
R20624 gnd.n7092 gnd.n7091 0.152939
R20625 gnd.n7091 gnd.n7066 0.152939
R20626 gnd.n7087 gnd.n7066 0.152939
R20627 gnd.n7087 gnd.n7086 0.152939
R20628 gnd.n7086 gnd.n7085 0.152939
R20629 gnd.n7085 gnd.n7074 0.152939
R20630 gnd.n7074 gnd.n78 0.152939
R20631 gnd.n5563 gnd.n5562 0.152939
R20632 gnd.n5563 gnd.n2799 0.152939
R20633 gnd.n5597 gnd.n2799 0.152939
R20634 gnd.n5598 gnd.n5597 0.152939
R20635 gnd.n5600 gnd.n5598 0.152939
R20636 gnd.n5600 gnd.n5599 0.152939
R20637 gnd.n5599 gnd.n2760 0.152939
R20638 gnd.n5628 gnd.n2760 0.152939
R20639 gnd.n5629 gnd.n5628 0.152939
R20640 gnd.n5637 gnd.n5629 0.152939
R20641 gnd.n5637 gnd.n5636 0.152939
R20642 gnd.n5636 gnd.n5635 0.152939
R20643 gnd.n5635 gnd.n5630 0.152939
R20644 gnd.n5630 gnd.n2715 0.152939
R20645 gnd.n5741 gnd.n2715 0.152939
R20646 gnd.n5741 gnd.n5740 0.152939
R20647 gnd.n5740 gnd.n5739 0.152939
R20648 gnd.n5739 gnd.n2716 0.152939
R20649 gnd.n5735 gnd.n2716 0.152939
R20650 gnd.n5735 gnd.n51 0.152939
R20651 gnd.n7227 gnd.n51 0.152939
R20652 gnd.n7227 gnd.n7226 0.152939
R20653 gnd.n7226 gnd.n53 0.152939
R20654 gnd.n7222 gnd.n53 0.152939
R20655 gnd.n7222 gnd.n7221 0.152939
R20656 gnd.n7221 gnd.n7220 0.152939
R20657 gnd.n7220 gnd.n58 0.152939
R20658 gnd.n7216 gnd.n58 0.152939
R20659 gnd.n7216 gnd.n7215 0.152939
R20660 gnd.n7215 gnd.n7214 0.152939
R20661 gnd.n7214 gnd.n63 0.152939
R20662 gnd.n7210 gnd.n63 0.152939
R20663 gnd.n7210 gnd.n7209 0.152939
R20664 gnd.n7209 gnd.n7208 0.152939
R20665 gnd.n7208 gnd.n68 0.152939
R20666 gnd.n7204 gnd.n68 0.152939
R20667 gnd.n7204 gnd.n7203 0.152939
R20668 gnd.n7203 gnd.n7202 0.152939
R20669 gnd.n7202 gnd.n73 0.152939
R20670 gnd.n7198 gnd.n73 0.152939
R20671 gnd.n7198 gnd.n7197 0.152939
R20672 gnd.n7197 gnd.n7196 0.152939
R20673 gnd.n5561 gnd.n5560 0.151415
R20674 gnd.n4536 gnd.n3718 0.151415
R20675 gnd.n4347 gnd.n3945 0.145814
R20676 gnd.n4347 gnd.n4346 0.145814
R20677 gnd.n1132 gnd.n0 0.127478
R20678 gnd.n260 gnd.n225 0.10111
R20679 gnd.n4363 gnd.n4362 0.10111
R20680 gnd.n1712 gnd.n1711 0.0767195
R20681 gnd.n1711 gnd.n1710 0.0767195
R20682 gnd.n5922 gnd.n5921 0.063
R20683 gnd.n2855 gnd.n2852 0.063
R20684 gnd.n4364 gnd.n4363 0.0523293
R20685 gnd.n5652 gnd.n225 0.0523293
R20686 gnd.n2280 gnd.n908 0.0477147
R20687 gnd.n1475 gnd.n1363 0.0442063
R20688 gnd.n1476 gnd.n1475 0.0442063
R20689 gnd.n1477 gnd.n1476 0.0442063
R20690 gnd.n1477 gnd.n1352 0.0442063
R20691 gnd.n1491 gnd.n1352 0.0442063
R20692 gnd.n1492 gnd.n1491 0.0442063
R20693 gnd.n1493 gnd.n1492 0.0442063
R20694 gnd.n1493 gnd.n1339 0.0442063
R20695 gnd.n1537 gnd.n1339 0.0442063
R20696 gnd.n1538 gnd.n1537 0.0442063
R20697 gnd.n1540 gnd.n1273 0.0344674
R20698 gnd.n2939 gnd.n2806 0.0344674
R20699 gnd.n4535 gnd.n3719 0.0344674
R20700 gnd.n1560 gnd.n1559 0.0269946
R20701 gnd.n1562 gnd.n1561 0.0269946
R20702 gnd.n1268 gnd.n1266 0.0269946
R20703 gnd.n1572 gnd.n1570 0.0269946
R20704 gnd.n1571 gnd.n1247 0.0269946
R20705 gnd.n1591 gnd.n1590 0.0269946
R20706 gnd.n1593 gnd.n1592 0.0269946
R20707 gnd.n1242 gnd.n1241 0.0269946
R20708 gnd.n1603 gnd.n1237 0.0269946
R20709 gnd.n1602 gnd.n1239 0.0269946
R20710 gnd.n1238 gnd.n1220 0.0269946
R20711 gnd.n1623 gnd.n1221 0.0269946
R20712 gnd.n1622 gnd.n1222 0.0269946
R20713 gnd.n1656 gnd.n1197 0.0269946
R20714 gnd.n1658 gnd.n1657 0.0269946
R20715 gnd.n1659 gnd.n1144 0.0269946
R20716 gnd.n1192 gnd.n1145 0.0269946
R20717 gnd.n1194 gnd.n1146 0.0269946
R20718 gnd.n1669 gnd.n1668 0.0269946
R20719 gnd.n1671 gnd.n1670 0.0269946
R20720 gnd.n1672 gnd.n1166 0.0269946
R20721 gnd.n1674 gnd.n1167 0.0269946
R20722 gnd.n1677 gnd.n1168 0.0269946
R20723 gnd.n1680 gnd.n1679 0.0269946
R20724 gnd.n1682 gnd.n1681 0.0269946
R20725 gnd.n1747 gnd.n1079 0.0269946
R20726 gnd.n1749 gnd.n1748 0.0269946
R20727 gnd.n1758 gnd.n1072 0.0269946
R20728 gnd.n1760 gnd.n1759 0.0269946
R20729 gnd.n1761 gnd.n1070 0.0269946
R20730 gnd.n1768 gnd.n1764 0.0269946
R20731 gnd.n1767 gnd.n1766 0.0269946
R20732 gnd.n1765 gnd.n1049 0.0269946
R20733 gnd.n1790 gnd.n1050 0.0269946
R20734 gnd.n1789 gnd.n1051 0.0269946
R20735 gnd.n1834 gnd.n1026 0.0269946
R20736 gnd.n1836 gnd.n1835 0.0269946
R20737 gnd.n1845 gnd.n1019 0.0269946
R20738 gnd.n1847 gnd.n1846 0.0269946
R20739 gnd.n1848 gnd.n1017 0.0269946
R20740 gnd.n1855 gnd.n1851 0.0269946
R20741 gnd.n1854 gnd.n1853 0.0269946
R20742 gnd.n1852 gnd.n996 0.0269946
R20743 gnd.n1877 gnd.n997 0.0269946
R20744 gnd.n1876 gnd.n998 0.0269946
R20745 gnd.n1923 gnd.n972 0.0269946
R20746 gnd.n1925 gnd.n1924 0.0269946
R20747 gnd.n1934 gnd.n965 0.0269946
R20748 gnd.n2193 gnd.n963 0.0269946
R20749 gnd.n2198 gnd.n2196 0.0269946
R20750 gnd.n2197 gnd.n944 0.0269946
R20751 gnd.n2222 gnd.n2221 0.0269946
R20752 gnd.n2852 gnd.n2851 0.0246168
R20753 gnd.n5921 gnd.n2541 0.0246168
R20754 gnd.n1540 gnd.n1539 0.0202011
R20755 gnd.n2851 gnd.n2849 0.0174837
R20756 gnd.n2863 gnd.n2849 0.0174837
R20757 gnd.n2865 gnd.n2863 0.0174837
R20758 gnd.n2865 gnd.n2864 0.0174837
R20759 gnd.n2864 gnd.n2844 0.0174837
R20760 gnd.n2874 gnd.n2844 0.0174837
R20761 gnd.n2874 gnd.n2873 0.0174837
R20762 gnd.n2873 gnd.n2845 0.0174837
R20763 gnd.n2845 gnd.n2840 0.0174837
R20764 gnd.n2882 gnd.n2840 0.0174837
R20765 gnd.n2884 gnd.n2882 0.0174837
R20766 gnd.n2884 gnd.n2883 0.0174837
R20767 gnd.n2883 gnd.n2835 0.0174837
R20768 gnd.n2893 gnd.n2835 0.0174837
R20769 gnd.n2893 gnd.n2892 0.0174837
R20770 gnd.n2892 gnd.n2836 0.0174837
R20771 gnd.n2836 gnd.n2831 0.0174837
R20772 gnd.n2901 gnd.n2831 0.0174837
R20773 gnd.n2903 gnd.n2901 0.0174837
R20774 gnd.n2903 gnd.n2902 0.0174837
R20775 gnd.n2902 gnd.n2826 0.0174837
R20776 gnd.n2912 gnd.n2826 0.0174837
R20777 gnd.n2912 gnd.n2911 0.0174837
R20778 gnd.n2911 gnd.n2827 0.0174837
R20779 gnd.n2827 gnd.n2822 0.0174837
R20780 gnd.n2920 gnd.n2822 0.0174837
R20781 gnd.n2922 gnd.n2920 0.0174837
R20782 gnd.n2922 gnd.n2921 0.0174837
R20783 gnd.n2921 gnd.n2817 0.0174837
R20784 gnd.n2931 gnd.n2817 0.0174837
R20785 gnd.n2931 gnd.n2930 0.0174837
R20786 gnd.n2930 gnd.n2818 0.0174837
R20787 gnd.n2818 gnd.n2811 0.0174837
R20788 gnd.n2938 gnd.n2811 0.0174837
R20789 gnd.n2939 gnd.n2938 0.0174837
R20790 gnd.n3775 gnd.n2541 0.0174837
R20791 gnd.n3777 gnd.n3775 0.0174837
R20792 gnd.n3885 gnd.n3777 0.0174837
R20793 gnd.n3885 gnd.n3884 0.0174837
R20794 gnd.n3884 gnd.n3778 0.0174837
R20795 gnd.n3881 gnd.n3778 0.0174837
R20796 gnd.n3881 gnd.n3880 0.0174837
R20797 gnd.n3880 gnd.n3788 0.0174837
R20798 gnd.n3877 gnd.n3788 0.0174837
R20799 gnd.n3877 gnd.n3876 0.0174837
R20800 gnd.n3876 gnd.n3793 0.0174837
R20801 gnd.n3873 gnd.n3793 0.0174837
R20802 gnd.n3873 gnd.n3872 0.0174837
R20803 gnd.n3872 gnd.n3799 0.0174837
R20804 gnd.n3869 gnd.n3799 0.0174837
R20805 gnd.n3869 gnd.n3868 0.0174837
R20806 gnd.n3868 gnd.n3803 0.0174837
R20807 gnd.n3865 gnd.n3803 0.0174837
R20808 gnd.n3865 gnd.n3864 0.0174837
R20809 gnd.n3864 gnd.n3810 0.0174837
R20810 gnd.n3861 gnd.n3810 0.0174837
R20811 gnd.n3861 gnd.n3860 0.0174837
R20812 gnd.n3860 gnd.n3816 0.0174837
R20813 gnd.n3857 gnd.n3816 0.0174837
R20814 gnd.n3857 gnd.n3856 0.0174837
R20815 gnd.n3856 gnd.n3822 0.0174837
R20816 gnd.n3853 gnd.n3822 0.0174837
R20817 gnd.n3853 gnd.n3852 0.0174837
R20818 gnd.n3852 gnd.n3826 0.0174837
R20819 gnd.n3849 gnd.n3826 0.0174837
R20820 gnd.n3849 gnd.n3848 0.0174837
R20821 gnd.n3848 gnd.n3835 0.0174837
R20822 gnd.n3845 gnd.n3835 0.0174837
R20823 gnd.n3845 gnd.n3844 0.0174837
R20824 gnd.n3844 gnd.n3719 0.0174837
R20825 gnd.n1539 gnd.n1538 0.0148637
R20826 gnd.n2191 gnd.n1935 0.0144266
R20827 gnd.n2192 gnd.n2191 0.0130679
R20828 gnd.n1559 gnd.n1273 0.00797283
R20829 gnd.n1561 gnd.n1560 0.00797283
R20830 gnd.n1562 gnd.n1268 0.00797283
R20831 gnd.n1570 gnd.n1266 0.00797283
R20832 gnd.n1572 gnd.n1571 0.00797283
R20833 gnd.n1590 gnd.n1247 0.00797283
R20834 gnd.n1592 gnd.n1591 0.00797283
R20835 gnd.n1593 gnd.n1242 0.00797283
R20836 gnd.n1241 gnd.n1237 0.00797283
R20837 gnd.n1603 gnd.n1602 0.00797283
R20838 gnd.n1239 gnd.n1238 0.00797283
R20839 gnd.n1221 gnd.n1220 0.00797283
R20840 gnd.n1623 gnd.n1622 0.00797283
R20841 gnd.n1222 gnd.n1197 0.00797283
R20842 gnd.n1657 gnd.n1656 0.00797283
R20843 gnd.n1659 gnd.n1658 0.00797283
R20844 gnd.n1192 gnd.n1144 0.00797283
R20845 gnd.n1194 gnd.n1145 0.00797283
R20846 gnd.n1668 gnd.n1146 0.00797283
R20847 gnd.n1670 gnd.n1669 0.00797283
R20848 gnd.n1672 gnd.n1671 0.00797283
R20849 gnd.n1674 gnd.n1166 0.00797283
R20850 gnd.n1677 gnd.n1167 0.00797283
R20851 gnd.n1679 gnd.n1168 0.00797283
R20852 gnd.n1682 gnd.n1680 0.00797283
R20853 gnd.n1681 gnd.n1079 0.00797283
R20854 gnd.n1749 gnd.n1747 0.00797283
R20855 gnd.n1748 gnd.n1072 0.00797283
R20856 gnd.n1759 gnd.n1758 0.00797283
R20857 gnd.n1761 gnd.n1760 0.00797283
R20858 gnd.n1764 gnd.n1070 0.00797283
R20859 gnd.n1768 gnd.n1767 0.00797283
R20860 gnd.n1766 gnd.n1765 0.00797283
R20861 gnd.n1050 gnd.n1049 0.00797283
R20862 gnd.n1790 gnd.n1789 0.00797283
R20863 gnd.n1051 gnd.n1026 0.00797283
R20864 gnd.n1836 gnd.n1834 0.00797283
R20865 gnd.n1835 gnd.n1019 0.00797283
R20866 gnd.n1846 gnd.n1845 0.00797283
R20867 gnd.n1848 gnd.n1847 0.00797283
R20868 gnd.n1851 gnd.n1017 0.00797283
R20869 gnd.n1855 gnd.n1854 0.00797283
R20870 gnd.n1853 gnd.n1852 0.00797283
R20871 gnd.n997 gnd.n996 0.00797283
R20872 gnd.n1877 gnd.n1876 0.00797283
R20873 gnd.n998 gnd.n972 0.00797283
R20874 gnd.n1925 gnd.n1923 0.00797283
R20875 gnd.n1924 gnd.n965 0.00797283
R20876 gnd.n1935 gnd.n1934 0.00797283
R20877 gnd.n2193 gnd.n2192 0.00797283
R20878 gnd.n2196 gnd.n963 0.00797283
R20879 gnd.n2198 gnd.n2197 0.00797283
R20880 gnd.n2221 gnd.n944 0.00797283
R20881 gnd.n2222 gnd.n908 0.00797283
R20882 gnd.n5693 gnd.n242 0.00614909
R20883 gnd.n4311 gnd.n3953 0.00614909
R20884 gnd.n5561 gnd.n2806 0.000839674
R20885 gnd.n4536 gnd.n4535 0.000839674
R20886 commonsourceibias.n25 commonsourceibias.t46 230.006
R20887 commonsourceibias.n91 commonsourceibias.t62 230.006
R20888 commonsourceibias.n154 commonsourceibias.t54 230.006
R20889 commonsourceibias.n258 commonsourceibias.t16 230.006
R20890 commonsourceibias.n217 commonsourceibias.t75 230.006
R20891 commonsourceibias.n355 commonsourceibias.t65 230.006
R20892 commonsourceibias.n70 commonsourceibias.t32 207.983
R20893 commonsourceibias.n136 commonsourceibias.t71 207.983
R20894 commonsourceibias.n199 commonsourceibias.t61 207.983
R20895 commonsourceibias.n304 commonsourceibias.t2 207.983
R20896 commonsourceibias.n338 commonsourceibias.t84 207.983
R20897 commonsourceibias.n401 commonsourceibias.t73 207.983
R20898 commonsourceibias.n10 commonsourceibias.t14 168.701
R20899 commonsourceibias.n63 commonsourceibias.t24 168.701
R20900 commonsourceibias.n57 commonsourceibias.t30 168.701
R20901 commonsourceibias.n16 commonsourceibias.t20 168.701
R20902 commonsourceibias.n49 commonsourceibias.t36 168.701
R20903 commonsourceibias.n43 commonsourceibias.t44 168.701
R20904 commonsourceibias.n19 commonsourceibias.t26 168.701
R20905 commonsourceibias.n21 commonsourceibias.t34 168.701
R20906 commonsourceibias.n23 commonsourceibias.t10 168.701
R20907 commonsourceibias.n26 commonsourceibias.t40 168.701
R20908 commonsourceibias.n1 commonsourceibias.t81 168.701
R20909 commonsourceibias.n129 commonsourceibias.t55 168.701
R20910 commonsourceibias.n123 commonsourceibias.t53 168.701
R20911 commonsourceibias.n7 commonsourceibias.t76 168.701
R20912 commonsourceibias.n115 commonsourceibias.t86 168.701
R20913 commonsourceibias.n109 commonsourceibias.t50 168.701
R20914 commonsourceibias.n85 commonsourceibias.t69 168.701
R20915 commonsourceibias.n87 commonsourceibias.t67 168.701
R20916 commonsourceibias.n89 commonsourceibias.t78 168.701
R20917 commonsourceibias.n92 commonsourceibias.t64 168.701
R20918 commonsourceibias.n155 commonsourceibias.t57 168.701
R20919 commonsourceibias.n152 commonsourceibias.t68 168.701
R20920 commonsourceibias.n150 commonsourceibias.t58 168.701
R20921 commonsourceibias.n148 commonsourceibias.t60 168.701
R20922 commonsourceibias.n172 commonsourceibias.t91 168.701
R20923 commonsourceibias.n178 commonsourceibias.t77 168.701
R20924 commonsourceibias.n145 commonsourceibias.t66 168.701
R20925 commonsourceibias.n186 commonsourceibias.t95 168.701
R20926 commonsourceibias.n192 commonsourceibias.t49 168.701
R20927 commonsourceibias.n139 commonsourceibias.t72 168.701
R20928 commonsourceibias.n259 commonsourceibias.t8 168.701
R20929 commonsourceibias.n256 commonsourceibias.t18 168.701
R20930 commonsourceibias.n254 commonsourceibias.t4 168.701
R20931 commonsourceibias.n252 commonsourceibias.t42 168.701
R20932 commonsourceibias.n276 commonsourceibias.t12 168.701
R20933 commonsourceibias.n282 commonsourceibias.t6 168.701
R20934 commonsourceibias.n284 commonsourceibias.t28 168.701
R20935 commonsourceibias.n291 commonsourceibias.t0 168.701
R20936 commonsourceibias.n297 commonsourceibias.t38 168.701
R20937 commonsourceibias.n244 commonsourceibias.t22 168.701
R20938 commonsourceibias.n203 commonsourceibias.t92 168.701
R20939 commonsourceibias.n331 commonsourceibias.t51 168.701
R20940 commonsourceibias.n325 commonsourceibias.t63 168.701
R20941 commonsourceibias.n318 commonsourceibias.t88 168.701
R20942 commonsourceibias.n316 commonsourceibias.t48 168.701
R20943 commonsourceibias.n218 commonsourceibias.t59 168.701
R20944 commonsourceibias.n215 commonsourceibias.t90 168.701
R20945 commonsourceibias.n213 commonsourceibias.t80 168.701
R20946 commonsourceibias.n211 commonsourceibias.t83 168.701
R20947 commonsourceibias.n235 commonsourceibias.t94 168.701
R20948 commonsourceibias.n356 commonsourceibias.t52 168.701
R20949 commonsourceibias.n353 commonsourceibias.t82 168.701
R20950 commonsourceibias.n351 commonsourceibias.t70 168.701
R20951 commonsourceibias.n349 commonsourceibias.t74 168.701
R20952 commonsourceibias.n373 commonsourceibias.t87 168.701
R20953 commonsourceibias.n379 commonsourceibias.t89 168.701
R20954 commonsourceibias.n381 commonsourceibias.t79 168.701
R20955 commonsourceibias.n388 commonsourceibias.t56 168.701
R20956 commonsourceibias.n394 commonsourceibias.t93 168.701
R20957 commonsourceibias.n341 commonsourceibias.t85 168.701
R20958 commonsourceibias.n27 commonsourceibias.n24 161.3
R20959 commonsourceibias.n29 commonsourceibias.n28 161.3
R20960 commonsourceibias.n31 commonsourceibias.n30 161.3
R20961 commonsourceibias.n32 commonsourceibias.n22 161.3
R20962 commonsourceibias.n34 commonsourceibias.n33 161.3
R20963 commonsourceibias.n36 commonsourceibias.n35 161.3
R20964 commonsourceibias.n37 commonsourceibias.n20 161.3
R20965 commonsourceibias.n39 commonsourceibias.n38 161.3
R20966 commonsourceibias.n41 commonsourceibias.n40 161.3
R20967 commonsourceibias.n42 commonsourceibias.n18 161.3
R20968 commonsourceibias.n45 commonsourceibias.n44 161.3
R20969 commonsourceibias.n46 commonsourceibias.n17 161.3
R20970 commonsourceibias.n48 commonsourceibias.n47 161.3
R20971 commonsourceibias.n50 commonsourceibias.n15 161.3
R20972 commonsourceibias.n52 commonsourceibias.n51 161.3
R20973 commonsourceibias.n53 commonsourceibias.n14 161.3
R20974 commonsourceibias.n55 commonsourceibias.n54 161.3
R20975 commonsourceibias.n56 commonsourceibias.n13 161.3
R20976 commonsourceibias.n59 commonsourceibias.n58 161.3
R20977 commonsourceibias.n60 commonsourceibias.n12 161.3
R20978 commonsourceibias.n62 commonsourceibias.n61 161.3
R20979 commonsourceibias.n64 commonsourceibias.n11 161.3
R20980 commonsourceibias.n66 commonsourceibias.n65 161.3
R20981 commonsourceibias.n68 commonsourceibias.n67 161.3
R20982 commonsourceibias.n69 commonsourceibias.n9 161.3
R20983 commonsourceibias.n93 commonsourceibias.n90 161.3
R20984 commonsourceibias.n95 commonsourceibias.n94 161.3
R20985 commonsourceibias.n97 commonsourceibias.n96 161.3
R20986 commonsourceibias.n98 commonsourceibias.n88 161.3
R20987 commonsourceibias.n100 commonsourceibias.n99 161.3
R20988 commonsourceibias.n102 commonsourceibias.n101 161.3
R20989 commonsourceibias.n103 commonsourceibias.n86 161.3
R20990 commonsourceibias.n105 commonsourceibias.n104 161.3
R20991 commonsourceibias.n107 commonsourceibias.n106 161.3
R20992 commonsourceibias.n108 commonsourceibias.n84 161.3
R20993 commonsourceibias.n111 commonsourceibias.n110 161.3
R20994 commonsourceibias.n112 commonsourceibias.n8 161.3
R20995 commonsourceibias.n114 commonsourceibias.n113 161.3
R20996 commonsourceibias.n116 commonsourceibias.n6 161.3
R20997 commonsourceibias.n118 commonsourceibias.n117 161.3
R20998 commonsourceibias.n119 commonsourceibias.n5 161.3
R20999 commonsourceibias.n121 commonsourceibias.n120 161.3
R21000 commonsourceibias.n122 commonsourceibias.n4 161.3
R21001 commonsourceibias.n125 commonsourceibias.n124 161.3
R21002 commonsourceibias.n126 commonsourceibias.n3 161.3
R21003 commonsourceibias.n128 commonsourceibias.n127 161.3
R21004 commonsourceibias.n130 commonsourceibias.n2 161.3
R21005 commonsourceibias.n132 commonsourceibias.n131 161.3
R21006 commonsourceibias.n134 commonsourceibias.n133 161.3
R21007 commonsourceibias.n135 commonsourceibias.n0 161.3
R21008 commonsourceibias.n198 commonsourceibias.n138 161.3
R21009 commonsourceibias.n197 commonsourceibias.n196 161.3
R21010 commonsourceibias.n195 commonsourceibias.n194 161.3
R21011 commonsourceibias.n193 commonsourceibias.n140 161.3
R21012 commonsourceibias.n191 commonsourceibias.n190 161.3
R21013 commonsourceibias.n189 commonsourceibias.n141 161.3
R21014 commonsourceibias.n188 commonsourceibias.n187 161.3
R21015 commonsourceibias.n185 commonsourceibias.n142 161.3
R21016 commonsourceibias.n184 commonsourceibias.n183 161.3
R21017 commonsourceibias.n182 commonsourceibias.n143 161.3
R21018 commonsourceibias.n181 commonsourceibias.n180 161.3
R21019 commonsourceibias.n179 commonsourceibias.n144 161.3
R21020 commonsourceibias.n177 commonsourceibias.n176 161.3
R21021 commonsourceibias.n175 commonsourceibias.n146 161.3
R21022 commonsourceibias.n174 commonsourceibias.n173 161.3
R21023 commonsourceibias.n171 commonsourceibias.n147 161.3
R21024 commonsourceibias.n170 commonsourceibias.n169 161.3
R21025 commonsourceibias.n168 commonsourceibias.n167 161.3
R21026 commonsourceibias.n166 commonsourceibias.n149 161.3
R21027 commonsourceibias.n165 commonsourceibias.n164 161.3
R21028 commonsourceibias.n163 commonsourceibias.n162 161.3
R21029 commonsourceibias.n161 commonsourceibias.n151 161.3
R21030 commonsourceibias.n160 commonsourceibias.n159 161.3
R21031 commonsourceibias.n158 commonsourceibias.n157 161.3
R21032 commonsourceibias.n156 commonsourceibias.n153 161.3
R21033 commonsourceibias.n303 commonsourceibias.n243 161.3
R21034 commonsourceibias.n302 commonsourceibias.n301 161.3
R21035 commonsourceibias.n300 commonsourceibias.n299 161.3
R21036 commonsourceibias.n298 commonsourceibias.n245 161.3
R21037 commonsourceibias.n296 commonsourceibias.n295 161.3
R21038 commonsourceibias.n294 commonsourceibias.n246 161.3
R21039 commonsourceibias.n293 commonsourceibias.n292 161.3
R21040 commonsourceibias.n290 commonsourceibias.n247 161.3
R21041 commonsourceibias.n289 commonsourceibias.n288 161.3
R21042 commonsourceibias.n287 commonsourceibias.n248 161.3
R21043 commonsourceibias.n286 commonsourceibias.n285 161.3
R21044 commonsourceibias.n283 commonsourceibias.n249 161.3
R21045 commonsourceibias.n281 commonsourceibias.n280 161.3
R21046 commonsourceibias.n279 commonsourceibias.n250 161.3
R21047 commonsourceibias.n278 commonsourceibias.n277 161.3
R21048 commonsourceibias.n275 commonsourceibias.n251 161.3
R21049 commonsourceibias.n274 commonsourceibias.n273 161.3
R21050 commonsourceibias.n272 commonsourceibias.n271 161.3
R21051 commonsourceibias.n270 commonsourceibias.n253 161.3
R21052 commonsourceibias.n269 commonsourceibias.n268 161.3
R21053 commonsourceibias.n267 commonsourceibias.n266 161.3
R21054 commonsourceibias.n265 commonsourceibias.n255 161.3
R21055 commonsourceibias.n264 commonsourceibias.n263 161.3
R21056 commonsourceibias.n262 commonsourceibias.n261 161.3
R21057 commonsourceibias.n260 commonsourceibias.n257 161.3
R21058 commonsourceibias.n237 commonsourceibias.n236 161.3
R21059 commonsourceibias.n234 commonsourceibias.n210 161.3
R21060 commonsourceibias.n233 commonsourceibias.n232 161.3
R21061 commonsourceibias.n231 commonsourceibias.n230 161.3
R21062 commonsourceibias.n229 commonsourceibias.n212 161.3
R21063 commonsourceibias.n228 commonsourceibias.n227 161.3
R21064 commonsourceibias.n226 commonsourceibias.n225 161.3
R21065 commonsourceibias.n224 commonsourceibias.n214 161.3
R21066 commonsourceibias.n223 commonsourceibias.n222 161.3
R21067 commonsourceibias.n221 commonsourceibias.n220 161.3
R21068 commonsourceibias.n219 commonsourceibias.n216 161.3
R21069 commonsourceibias.n313 commonsourceibias.n209 161.3
R21070 commonsourceibias.n337 commonsourceibias.n202 161.3
R21071 commonsourceibias.n336 commonsourceibias.n335 161.3
R21072 commonsourceibias.n334 commonsourceibias.n333 161.3
R21073 commonsourceibias.n332 commonsourceibias.n204 161.3
R21074 commonsourceibias.n330 commonsourceibias.n329 161.3
R21075 commonsourceibias.n328 commonsourceibias.n205 161.3
R21076 commonsourceibias.n327 commonsourceibias.n326 161.3
R21077 commonsourceibias.n324 commonsourceibias.n206 161.3
R21078 commonsourceibias.n323 commonsourceibias.n322 161.3
R21079 commonsourceibias.n321 commonsourceibias.n207 161.3
R21080 commonsourceibias.n320 commonsourceibias.n319 161.3
R21081 commonsourceibias.n317 commonsourceibias.n208 161.3
R21082 commonsourceibias.n315 commonsourceibias.n314 161.3
R21083 commonsourceibias.n400 commonsourceibias.n340 161.3
R21084 commonsourceibias.n399 commonsourceibias.n398 161.3
R21085 commonsourceibias.n397 commonsourceibias.n396 161.3
R21086 commonsourceibias.n395 commonsourceibias.n342 161.3
R21087 commonsourceibias.n393 commonsourceibias.n392 161.3
R21088 commonsourceibias.n391 commonsourceibias.n343 161.3
R21089 commonsourceibias.n390 commonsourceibias.n389 161.3
R21090 commonsourceibias.n387 commonsourceibias.n344 161.3
R21091 commonsourceibias.n386 commonsourceibias.n385 161.3
R21092 commonsourceibias.n384 commonsourceibias.n345 161.3
R21093 commonsourceibias.n383 commonsourceibias.n382 161.3
R21094 commonsourceibias.n380 commonsourceibias.n346 161.3
R21095 commonsourceibias.n378 commonsourceibias.n377 161.3
R21096 commonsourceibias.n376 commonsourceibias.n347 161.3
R21097 commonsourceibias.n375 commonsourceibias.n374 161.3
R21098 commonsourceibias.n372 commonsourceibias.n348 161.3
R21099 commonsourceibias.n371 commonsourceibias.n370 161.3
R21100 commonsourceibias.n369 commonsourceibias.n368 161.3
R21101 commonsourceibias.n367 commonsourceibias.n350 161.3
R21102 commonsourceibias.n366 commonsourceibias.n365 161.3
R21103 commonsourceibias.n364 commonsourceibias.n363 161.3
R21104 commonsourceibias.n362 commonsourceibias.n352 161.3
R21105 commonsourceibias.n361 commonsourceibias.n360 161.3
R21106 commonsourceibias.n359 commonsourceibias.n358 161.3
R21107 commonsourceibias.n357 commonsourceibias.n354 161.3
R21108 commonsourceibias.n80 commonsourceibias.n78 81.5057
R21109 commonsourceibias.n240 commonsourceibias.n238 81.5057
R21110 commonsourceibias.n80 commonsourceibias.n79 80.9324
R21111 commonsourceibias.n82 commonsourceibias.n81 80.9324
R21112 commonsourceibias.n77 commonsourceibias.n76 80.9324
R21113 commonsourceibias.n75 commonsourceibias.n74 80.9324
R21114 commonsourceibias.n73 commonsourceibias.n72 80.9324
R21115 commonsourceibias.n307 commonsourceibias.n306 80.9324
R21116 commonsourceibias.n309 commonsourceibias.n308 80.9324
R21117 commonsourceibias.n311 commonsourceibias.n310 80.9324
R21118 commonsourceibias.n242 commonsourceibias.n241 80.9324
R21119 commonsourceibias.n240 commonsourceibias.n239 80.9324
R21120 commonsourceibias.n71 commonsourceibias.n70 80.6037
R21121 commonsourceibias.n137 commonsourceibias.n136 80.6037
R21122 commonsourceibias.n200 commonsourceibias.n199 80.6037
R21123 commonsourceibias.n305 commonsourceibias.n304 80.6037
R21124 commonsourceibias.n339 commonsourceibias.n338 80.6037
R21125 commonsourceibias.n402 commonsourceibias.n401 80.6037
R21126 commonsourceibias.n65 commonsourceibias.n64 56.5617
R21127 commonsourceibias.n51 commonsourceibias.n50 56.5617
R21128 commonsourceibias.n42 commonsourceibias.n41 56.5617
R21129 commonsourceibias.n28 commonsourceibias.n27 56.5617
R21130 commonsourceibias.n131 commonsourceibias.n130 56.5617
R21131 commonsourceibias.n117 commonsourceibias.n116 56.5617
R21132 commonsourceibias.n108 commonsourceibias.n107 56.5617
R21133 commonsourceibias.n94 commonsourceibias.n93 56.5617
R21134 commonsourceibias.n157 commonsourceibias.n156 56.5617
R21135 commonsourceibias.n171 commonsourceibias.n170 56.5617
R21136 commonsourceibias.n180 commonsourceibias.n179 56.5617
R21137 commonsourceibias.n194 commonsourceibias.n193 56.5617
R21138 commonsourceibias.n261 commonsourceibias.n260 56.5617
R21139 commonsourceibias.n275 commonsourceibias.n274 56.5617
R21140 commonsourceibias.n285 commonsourceibias.n283 56.5617
R21141 commonsourceibias.n299 commonsourceibias.n298 56.5617
R21142 commonsourceibias.n333 commonsourceibias.n332 56.5617
R21143 commonsourceibias.n319 commonsourceibias.n317 56.5617
R21144 commonsourceibias.n220 commonsourceibias.n219 56.5617
R21145 commonsourceibias.n234 commonsourceibias.n233 56.5617
R21146 commonsourceibias.n358 commonsourceibias.n357 56.5617
R21147 commonsourceibias.n372 commonsourceibias.n371 56.5617
R21148 commonsourceibias.n382 commonsourceibias.n380 56.5617
R21149 commonsourceibias.n396 commonsourceibias.n395 56.5617
R21150 commonsourceibias.n56 commonsourceibias.n55 56.0773
R21151 commonsourceibias.n37 commonsourceibias.n36 56.0773
R21152 commonsourceibias.n122 commonsourceibias.n121 56.0773
R21153 commonsourceibias.n103 commonsourceibias.n102 56.0773
R21154 commonsourceibias.n166 commonsourceibias.n165 56.0773
R21155 commonsourceibias.n185 commonsourceibias.n184 56.0773
R21156 commonsourceibias.n270 commonsourceibias.n269 56.0773
R21157 commonsourceibias.n290 commonsourceibias.n289 56.0773
R21158 commonsourceibias.n324 commonsourceibias.n323 56.0773
R21159 commonsourceibias.n229 commonsourceibias.n228 56.0773
R21160 commonsourceibias.n367 commonsourceibias.n366 56.0773
R21161 commonsourceibias.n387 commonsourceibias.n386 56.0773
R21162 commonsourceibias.n70 commonsourceibias.n69 46.0096
R21163 commonsourceibias.n136 commonsourceibias.n135 46.0096
R21164 commonsourceibias.n199 commonsourceibias.n198 46.0096
R21165 commonsourceibias.n304 commonsourceibias.n303 46.0096
R21166 commonsourceibias.n338 commonsourceibias.n337 46.0096
R21167 commonsourceibias.n401 commonsourceibias.n400 46.0096
R21168 commonsourceibias.n58 commonsourceibias.n12 41.5458
R21169 commonsourceibias.n33 commonsourceibias.n32 41.5458
R21170 commonsourceibias.n124 commonsourceibias.n3 41.5458
R21171 commonsourceibias.n99 commonsourceibias.n98 41.5458
R21172 commonsourceibias.n162 commonsourceibias.n161 41.5458
R21173 commonsourceibias.n187 commonsourceibias.n141 41.5458
R21174 commonsourceibias.n266 commonsourceibias.n265 41.5458
R21175 commonsourceibias.n292 commonsourceibias.n246 41.5458
R21176 commonsourceibias.n326 commonsourceibias.n205 41.5458
R21177 commonsourceibias.n225 commonsourceibias.n224 41.5458
R21178 commonsourceibias.n363 commonsourceibias.n362 41.5458
R21179 commonsourceibias.n389 commonsourceibias.n343 41.5458
R21180 commonsourceibias.n48 commonsourceibias.n17 40.577
R21181 commonsourceibias.n44 commonsourceibias.n17 40.577
R21182 commonsourceibias.n114 commonsourceibias.n8 40.577
R21183 commonsourceibias.n110 commonsourceibias.n8 40.577
R21184 commonsourceibias.n173 commonsourceibias.n146 40.577
R21185 commonsourceibias.n177 commonsourceibias.n146 40.577
R21186 commonsourceibias.n277 commonsourceibias.n250 40.577
R21187 commonsourceibias.n281 commonsourceibias.n250 40.577
R21188 commonsourceibias.n315 commonsourceibias.n209 40.577
R21189 commonsourceibias.n236 commonsourceibias.n209 40.577
R21190 commonsourceibias.n374 commonsourceibias.n347 40.577
R21191 commonsourceibias.n378 commonsourceibias.n347 40.577
R21192 commonsourceibias.n62 commonsourceibias.n12 39.6083
R21193 commonsourceibias.n32 commonsourceibias.n31 39.6083
R21194 commonsourceibias.n128 commonsourceibias.n3 39.6083
R21195 commonsourceibias.n98 commonsourceibias.n97 39.6083
R21196 commonsourceibias.n161 commonsourceibias.n160 39.6083
R21197 commonsourceibias.n191 commonsourceibias.n141 39.6083
R21198 commonsourceibias.n265 commonsourceibias.n264 39.6083
R21199 commonsourceibias.n296 commonsourceibias.n246 39.6083
R21200 commonsourceibias.n330 commonsourceibias.n205 39.6083
R21201 commonsourceibias.n224 commonsourceibias.n223 39.6083
R21202 commonsourceibias.n362 commonsourceibias.n361 39.6083
R21203 commonsourceibias.n393 commonsourceibias.n343 39.6083
R21204 commonsourceibias.n26 commonsourceibias.n25 33.0515
R21205 commonsourceibias.n92 commonsourceibias.n91 33.0515
R21206 commonsourceibias.n155 commonsourceibias.n154 33.0515
R21207 commonsourceibias.n259 commonsourceibias.n258 33.0515
R21208 commonsourceibias.n218 commonsourceibias.n217 33.0515
R21209 commonsourceibias.n356 commonsourceibias.n355 33.0515
R21210 commonsourceibias.n25 commonsourceibias.n24 28.5514
R21211 commonsourceibias.n91 commonsourceibias.n90 28.5514
R21212 commonsourceibias.n154 commonsourceibias.n153 28.5514
R21213 commonsourceibias.n258 commonsourceibias.n257 28.5514
R21214 commonsourceibias.n217 commonsourceibias.n216 28.5514
R21215 commonsourceibias.n355 commonsourceibias.n354 28.5514
R21216 commonsourceibias.n69 commonsourceibias.n68 26.0455
R21217 commonsourceibias.n135 commonsourceibias.n134 26.0455
R21218 commonsourceibias.n198 commonsourceibias.n197 26.0455
R21219 commonsourceibias.n303 commonsourceibias.n302 26.0455
R21220 commonsourceibias.n337 commonsourceibias.n336 26.0455
R21221 commonsourceibias.n400 commonsourceibias.n399 26.0455
R21222 commonsourceibias.n55 commonsourceibias.n14 25.0767
R21223 commonsourceibias.n38 commonsourceibias.n37 25.0767
R21224 commonsourceibias.n121 commonsourceibias.n5 25.0767
R21225 commonsourceibias.n104 commonsourceibias.n103 25.0767
R21226 commonsourceibias.n167 commonsourceibias.n166 25.0767
R21227 commonsourceibias.n184 commonsourceibias.n143 25.0767
R21228 commonsourceibias.n271 commonsourceibias.n270 25.0767
R21229 commonsourceibias.n289 commonsourceibias.n248 25.0767
R21230 commonsourceibias.n323 commonsourceibias.n207 25.0767
R21231 commonsourceibias.n230 commonsourceibias.n229 25.0767
R21232 commonsourceibias.n368 commonsourceibias.n367 25.0767
R21233 commonsourceibias.n386 commonsourceibias.n345 25.0767
R21234 commonsourceibias.n51 commonsourceibias.n16 24.3464
R21235 commonsourceibias.n41 commonsourceibias.n19 24.3464
R21236 commonsourceibias.n117 commonsourceibias.n7 24.3464
R21237 commonsourceibias.n107 commonsourceibias.n85 24.3464
R21238 commonsourceibias.n170 commonsourceibias.n148 24.3464
R21239 commonsourceibias.n180 commonsourceibias.n145 24.3464
R21240 commonsourceibias.n274 commonsourceibias.n252 24.3464
R21241 commonsourceibias.n285 commonsourceibias.n284 24.3464
R21242 commonsourceibias.n319 commonsourceibias.n318 24.3464
R21243 commonsourceibias.n233 commonsourceibias.n211 24.3464
R21244 commonsourceibias.n371 commonsourceibias.n349 24.3464
R21245 commonsourceibias.n382 commonsourceibias.n381 24.3464
R21246 commonsourceibias.n65 commonsourceibias.n10 23.8546
R21247 commonsourceibias.n27 commonsourceibias.n26 23.8546
R21248 commonsourceibias.n131 commonsourceibias.n1 23.8546
R21249 commonsourceibias.n93 commonsourceibias.n92 23.8546
R21250 commonsourceibias.n156 commonsourceibias.n155 23.8546
R21251 commonsourceibias.n194 commonsourceibias.n139 23.8546
R21252 commonsourceibias.n260 commonsourceibias.n259 23.8546
R21253 commonsourceibias.n299 commonsourceibias.n244 23.8546
R21254 commonsourceibias.n333 commonsourceibias.n203 23.8546
R21255 commonsourceibias.n219 commonsourceibias.n218 23.8546
R21256 commonsourceibias.n357 commonsourceibias.n356 23.8546
R21257 commonsourceibias.n396 commonsourceibias.n341 23.8546
R21258 commonsourceibias.n64 commonsourceibias.n63 16.9689
R21259 commonsourceibias.n28 commonsourceibias.n23 16.9689
R21260 commonsourceibias.n130 commonsourceibias.n129 16.9689
R21261 commonsourceibias.n94 commonsourceibias.n89 16.9689
R21262 commonsourceibias.n157 commonsourceibias.n152 16.9689
R21263 commonsourceibias.n193 commonsourceibias.n192 16.9689
R21264 commonsourceibias.n261 commonsourceibias.n256 16.9689
R21265 commonsourceibias.n298 commonsourceibias.n297 16.9689
R21266 commonsourceibias.n332 commonsourceibias.n331 16.9689
R21267 commonsourceibias.n220 commonsourceibias.n215 16.9689
R21268 commonsourceibias.n358 commonsourceibias.n353 16.9689
R21269 commonsourceibias.n395 commonsourceibias.n394 16.9689
R21270 commonsourceibias.n50 commonsourceibias.n49 16.477
R21271 commonsourceibias.n43 commonsourceibias.n42 16.477
R21272 commonsourceibias.n116 commonsourceibias.n115 16.477
R21273 commonsourceibias.n109 commonsourceibias.n108 16.477
R21274 commonsourceibias.n172 commonsourceibias.n171 16.477
R21275 commonsourceibias.n179 commonsourceibias.n178 16.477
R21276 commonsourceibias.n276 commonsourceibias.n275 16.477
R21277 commonsourceibias.n283 commonsourceibias.n282 16.477
R21278 commonsourceibias.n317 commonsourceibias.n316 16.477
R21279 commonsourceibias.n235 commonsourceibias.n234 16.477
R21280 commonsourceibias.n373 commonsourceibias.n372 16.477
R21281 commonsourceibias.n380 commonsourceibias.n379 16.477
R21282 commonsourceibias.n57 commonsourceibias.n56 15.9852
R21283 commonsourceibias.n36 commonsourceibias.n21 15.9852
R21284 commonsourceibias.n123 commonsourceibias.n122 15.9852
R21285 commonsourceibias.n102 commonsourceibias.n87 15.9852
R21286 commonsourceibias.n165 commonsourceibias.n150 15.9852
R21287 commonsourceibias.n186 commonsourceibias.n185 15.9852
R21288 commonsourceibias.n269 commonsourceibias.n254 15.9852
R21289 commonsourceibias.n291 commonsourceibias.n290 15.9852
R21290 commonsourceibias.n325 commonsourceibias.n324 15.9852
R21291 commonsourceibias.n228 commonsourceibias.n213 15.9852
R21292 commonsourceibias.n366 commonsourceibias.n351 15.9852
R21293 commonsourceibias.n388 commonsourceibias.n387 15.9852
R21294 commonsourceibias.n73 commonsourceibias.n71 13.2057
R21295 commonsourceibias.n307 commonsourceibias.n305 13.2057
R21296 commonsourceibias.n404 commonsourceibias.n201 11.9876
R21297 commonsourceibias.n404 commonsourceibias.n403 10.3347
R21298 commonsourceibias.n112 commonsourceibias.n83 9.50363
R21299 commonsourceibias.n313 commonsourceibias.n312 9.50363
R21300 commonsourceibias.n201 commonsourceibias.n137 8.732
R21301 commonsourceibias.n403 commonsourceibias.n339 8.732
R21302 commonsourceibias.n58 commonsourceibias.n57 8.60764
R21303 commonsourceibias.n33 commonsourceibias.n21 8.60764
R21304 commonsourceibias.n124 commonsourceibias.n123 8.60764
R21305 commonsourceibias.n99 commonsourceibias.n87 8.60764
R21306 commonsourceibias.n162 commonsourceibias.n150 8.60764
R21307 commonsourceibias.n187 commonsourceibias.n186 8.60764
R21308 commonsourceibias.n266 commonsourceibias.n254 8.60764
R21309 commonsourceibias.n292 commonsourceibias.n291 8.60764
R21310 commonsourceibias.n326 commonsourceibias.n325 8.60764
R21311 commonsourceibias.n225 commonsourceibias.n213 8.60764
R21312 commonsourceibias.n363 commonsourceibias.n351 8.60764
R21313 commonsourceibias.n389 commonsourceibias.n388 8.60764
R21314 commonsourceibias.n49 commonsourceibias.n48 8.11581
R21315 commonsourceibias.n44 commonsourceibias.n43 8.11581
R21316 commonsourceibias.n115 commonsourceibias.n114 8.11581
R21317 commonsourceibias.n110 commonsourceibias.n109 8.11581
R21318 commonsourceibias.n173 commonsourceibias.n172 8.11581
R21319 commonsourceibias.n178 commonsourceibias.n177 8.11581
R21320 commonsourceibias.n277 commonsourceibias.n276 8.11581
R21321 commonsourceibias.n282 commonsourceibias.n281 8.11581
R21322 commonsourceibias.n316 commonsourceibias.n315 8.11581
R21323 commonsourceibias.n236 commonsourceibias.n235 8.11581
R21324 commonsourceibias.n374 commonsourceibias.n373 8.11581
R21325 commonsourceibias.n379 commonsourceibias.n378 8.11581
R21326 commonsourceibias.n63 commonsourceibias.n62 7.62397
R21327 commonsourceibias.n31 commonsourceibias.n23 7.62397
R21328 commonsourceibias.n129 commonsourceibias.n128 7.62397
R21329 commonsourceibias.n97 commonsourceibias.n89 7.62397
R21330 commonsourceibias.n160 commonsourceibias.n152 7.62397
R21331 commonsourceibias.n192 commonsourceibias.n191 7.62397
R21332 commonsourceibias.n264 commonsourceibias.n256 7.62397
R21333 commonsourceibias.n297 commonsourceibias.n296 7.62397
R21334 commonsourceibias.n331 commonsourceibias.n330 7.62397
R21335 commonsourceibias.n223 commonsourceibias.n215 7.62397
R21336 commonsourceibias.n361 commonsourceibias.n353 7.62397
R21337 commonsourceibias.n394 commonsourceibias.n393 7.62397
R21338 commonsourceibias.n201 commonsourceibias.n200 5.00473
R21339 commonsourceibias.n403 commonsourceibias.n402 5.00473
R21340 commonsourceibias commonsourceibias.n404 3.87639
R21341 commonsourceibias.n78 commonsourceibias.t41 2.82907
R21342 commonsourceibias.n78 commonsourceibias.t47 2.82907
R21343 commonsourceibias.n79 commonsourceibias.t35 2.82907
R21344 commonsourceibias.n79 commonsourceibias.t11 2.82907
R21345 commonsourceibias.n81 commonsourceibias.t45 2.82907
R21346 commonsourceibias.n81 commonsourceibias.t27 2.82907
R21347 commonsourceibias.n76 commonsourceibias.t21 2.82907
R21348 commonsourceibias.n76 commonsourceibias.t37 2.82907
R21349 commonsourceibias.n74 commonsourceibias.t25 2.82907
R21350 commonsourceibias.n74 commonsourceibias.t31 2.82907
R21351 commonsourceibias.n72 commonsourceibias.t33 2.82907
R21352 commonsourceibias.n72 commonsourceibias.t15 2.82907
R21353 commonsourceibias.n306 commonsourceibias.t23 2.82907
R21354 commonsourceibias.n306 commonsourceibias.t3 2.82907
R21355 commonsourceibias.n308 commonsourceibias.t1 2.82907
R21356 commonsourceibias.n308 commonsourceibias.t39 2.82907
R21357 commonsourceibias.n310 commonsourceibias.t7 2.82907
R21358 commonsourceibias.n310 commonsourceibias.t29 2.82907
R21359 commonsourceibias.n241 commonsourceibias.t43 2.82907
R21360 commonsourceibias.n241 commonsourceibias.t13 2.82907
R21361 commonsourceibias.n239 commonsourceibias.t19 2.82907
R21362 commonsourceibias.n239 commonsourceibias.t5 2.82907
R21363 commonsourceibias.n238 commonsourceibias.t17 2.82907
R21364 commonsourceibias.n238 commonsourceibias.t9 2.82907
R21365 commonsourceibias.n68 commonsourceibias.n10 0.738255
R21366 commonsourceibias.n134 commonsourceibias.n1 0.738255
R21367 commonsourceibias.n197 commonsourceibias.n139 0.738255
R21368 commonsourceibias.n302 commonsourceibias.n244 0.738255
R21369 commonsourceibias.n336 commonsourceibias.n203 0.738255
R21370 commonsourceibias.n399 commonsourceibias.n341 0.738255
R21371 commonsourceibias.n75 commonsourceibias.n73 0.573776
R21372 commonsourceibias.n77 commonsourceibias.n75 0.573776
R21373 commonsourceibias.n82 commonsourceibias.n80 0.573776
R21374 commonsourceibias.n242 commonsourceibias.n240 0.573776
R21375 commonsourceibias.n311 commonsourceibias.n309 0.573776
R21376 commonsourceibias.n309 commonsourceibias.n307 0.573776
R21377 commonsourceibias.n83 commonsourceibias.n77 0.287138
R21378 commonsourceibias.n83 commonsourceibias.n82 0.287138
R21379 commonsourceibias.n312 commonsourceibias.n242 0.287138
R21380 commonsourceibias.n312 commonsourceibias.n311 0.287138
R21381 commonsourceibias.n71 commonsourceibias.n9 0.285035
R21382 commonsourceibias.n137 commonsourceibias.n0 0.285035
R21383 commonsourceibias.n200 commonsourceibias.n138 0.285035
R21384 commonsourceibias.n305 commonsourceibias.n243 0.285035
R21385 commonsourceibias.n339 commonsourceibias.n202 0.285035
R21386 commonsourceibias.n402 commonsourceibias.n340 0.285035
R21387 commonsourceibias.n16 commonsourceibias.n14 0.246418
R21388 commonsourceibias.n38 commonsourceibias.n19 0.246418
R21389 commonsourceibias.n7 commonsourceibias.n5 0.246418
R21390 commonsourceibias.n104 commonsourceibias.n85 0.246418
R21391 commonsourceibias.n167 commonsourceibias.n148 0.246418
R21392 commonsourceibias.n145 commonsourceibias.n143 0.246418
R21393 commonsourceibias.n271 commonsourceibias.n252 0.246418
R21394 commonsourceibias.n284 commonsourceibias.n248 0.246418
R21395 commonsourceibias.n318 commonsourceibias.n207 0.246418
R21396 commonsourceibias.n230 commonsourceibias.n211 0.246418
R21397 commonsourceibias.n368 commonsourceibias.n349 0.246418
R21398 commonsourceibias.n381 commonsourceibias.n345 0.246418
R21399 commonsourceibias.n67 commonsourceibias.n9 0.189894
R21400 commonsourceibias.n67 commonsourceibias.n66 0.189894
R21401 commonsourceibias.n66 commonsourceibias.n11 0.189894
R21402 commonsourceibias.n61 commonsourceibias.n11 0.189894
R21403 commonsourceibias.n61 commonsourceibias.n60 0.189894
R21404 commonsourceibias.n60 commonsourceibias.n59 0.189894
R21405 commonsourceibias.n59 commonsourceibias.n13 0.189894
R21406 commonsourceibias.n54 commonsourceibias.n13 0.189894
R21407 commonsourceibias.n54 commonsourceibias.n53 0.189894
R21408 commonsourceibias.n53 commonsourceibias.n52 0.189894
R21409 commonsourceibias.n52 commonsourceibias.n15 0.189894
R21410 commonsourceibias.n47 commonsourceibias.n15 0.189894
R21411 commonsourceibias.n47 commonsourceibias.n46 0.189894
R21412 commonsourceibias.n46 commonsourceibias.n45 0.189894
R21413 commonsourceibias.n45 commonsourceibias.n18 0.189894
R21414 commonsourceibias.n40 commonsourceibias.n18 0.189894
R21415 commonsourceibias.n40 commonsourceibias.n39 0.189894
R21416 commonsourceibias.n39 commonsourceibias.n20 0.189894
R21417 commonsourceibias.n35 commonsourceibias.n20 0.189894
R21418 commonsourceibias.n35 commonsourceibias.n34 0.189894
R21419 commonsourceibias.n34 commonsourceibias.n22 0.189894
R21420 commonsourceibias.n30 commonsourceibias.n22 0.189894
R21421 commonsourceibias.n30 commonsourceibias.n29 0.189894
R21422 commonsourceibias.n29 commonsourceibias.n24 0.189894
R21423 commonsourceibias.n111 commonsourceibias.n84 0.189894
R21424 commonsourceibias.n106 commonsourceibias.n84 0.189894
R21425 commonsourceibias.n106 commonsourceibias.n105 0.189894
R21426 commonsourceibias.n105 commonsourceibias.n86 0.189894
R21427 commonsourceibias.n101 commonsourceibias.n86 0.189894
R21428 commonsourceibias.n101 commonsourceibias.n100 0.189894
R21429 commonsourceibias.n100 commonsourceibias.n88 0.189894
R21430 commonsourceibias.n96 commonsourceibias.n88 0.189894
R21431 commonsourceibias.n96 commonsourceibias.n95 0.189894
R21432 commonsourceibias.n95 commonsourceibias.n90 0.189894
R21433 commonsourceibias.n133 commonsourceibias.n0 0.189894
R21434 commonsourceibias.n133 commonsourceibias.n132 0.189894
R21435 commonsourceibias.n132 commonsourceibias.n2 0.189894
R21436 commonsourceibias.n127 commonsourceibias.n2 0.189894
R21437 commonsourceibias.n127 commonsourceibias.n126 0.189894
R21438 commonsourceibias.n126 commonsourceibias.n125 0.189894
R21439 commonsourceibias.n125 commonsourceibias.n4 0.189894
R21440 commonsourceibias.n120 commonsourceibias.n4 0.189894
R21441 commonsourceibias.n120 commonsourceibias.n119 0.189894
R21442 commonsourceibias.n119 commonsourceibias.n118 0.189894
R21443 commonsourceibias.n118 commonsourceibias.n6 0.189894
R21444 commonsourceibias.n113 commonsourceibias.n6 0.189894
R21445 commonsourceibias.n196 commonsourceibias.n138 0.189894
R21446 commonsourceibias.n196 commonsourceibias.n195 0.189894
R21447 commonsourceibias.n195 commonsourceibias.n140 0.189894
R21448 commonsourceibias.n190 commonsourceibias.n140 0.189894
R21449 commonsourceibias.n190 commonsourceibias.n189 0.189894
R21450 commonsourceibias.n189 commonsourceibias.n188 0.189894
R21451 commonsourceibias.n188 commonsourceibias.n142 0.189894
R21452 commonsourceibias.n183 commonsourceibias.n142 0.189894
R21453 commonsourceibias.n183 commonsourceibias.n182 0.189894
R21454 commonsourceibias.n182 commonsourceibias.n181 0.189894
R21455 commonsourceibias.n181 commonsourceibias.n144 0.189894
R21456 commonsourceibias.n176 commonsourceibias.n144 0.189894
R21457 commonsourceibias.n176 commonsourceibias.n175 0.189894
R21458 commonsourceibias.n175 commonsourceibias.n174 0.189894
R21459 commonsourceibias.n174 commonsourceibias.n147 0.189894
R21460 commonsourceibias.n169 commonsourceibias.n147 0.189894
R21461 commonsourceibias.n169 commonsourceibias.n168 0.189894
R21462 commonsourceibias.n168 commonsourceibias.n149 0.189894
R21463 commonsourceibias.n164 commonsourceibias.n149 0.189894
R21464 commonsourceibias.n164 commonsourceibias.n163 0.189894
R21465 commonsourceibias.n163 commonsourceibias.n151 0.189894
R21466 commonsourceibias.n159 commonsourceibias.n151 0.189894
R21467 commonsourceibias.n159 commonsourceibias.n158 0.189894
R21468 commonsourceibias.n158 commonsourceibias.n153 0.189894
R21469 commonsourceibias.n262 commonsourceibias.n257 0.189894
R21470 commonsourceibias.n263 commonsourceibias.n262 0.189894
R21471 commonsourceibias.n263 commonsourceibias.n255 0.189894
R21472 commonsourceibias.n267 commonsourceibias.n255 0.189894
R21473 commonsourceibias.n268 commonsourceibias.n267 0.189894
R21474 commonsourceibias.n268 commonsourceibias.n253 0.189894
R21475 commonsourceibias.n272 commonsourceibias.n253 0.189894
R21476 commonsourceibias.n273 commonsourceibias.n272 0.189894
R21477 commonsourceibias.n273 commonsourceibias.n251 0.189894
R21478 commonsourceibias.n278 commonsourceibias.n251 0.189894
R21479 commonsourceibias.n279 commonsourceibias.n278 0.189894
R21480 commonsourceibias.n280 commonsourceibias.n279 0.189894
R21481 commonsourceibias.n280 commonsourceibias.n249 0.189894
R21482 commonsourceibias.n286 commonsourceibias.n249 0.189894
R21483 commonsourceibias.n287 commonsourceibias.n286 0.189894
R21484 commonsourceibias.n288 commonsourceibias.n287 0.189894
R21485 commonsourceibias.n288 commonsourceibias.n247 0.189894
R21486 commonsourceibias.n293 commonsourceibias.n247 0.189894
R21487 commonsourceibias.n294 commonsourceibias.n293 0.189894
R21488 commonsourceibias.n295 commonsourceibias.n294 0.189894
R21489 commonsourceibias.n295 commonsourceibias.n245 0.189894
R21490 commonsourceibias.n300 commonsourceibias.n245 0.189894
R21491 commonsourceibias.n301 commonsourceibias.n300 0.189894
R21492 commonsourceibias.n301 commonsourceibias.n243 0.189894
R21493 commonsourceibias.n221 commonsourceibias.n216 0.189894
R21494 commonsourceibias.n222 commonsourceibias.n221 0.189894
R21495 commonsourceibias.n222 commonsourceibias.n214 0.189894
R21496 commonsourceibias.n226 commonsourceibias.n214 0.189894
R21497 commonsourceibias.n227 commonsourceibias.n226 0.189894
R21498 commonsourceibias.n227 commonsourceibias.n212 0.189894
R21499 commonsourceibias.n231 commonsourceibias.n212 0.189894
R21500 commonsourceibias.n232 commonsourceibias.n231 0.189894
R21501 commonsourceibias.n232 commonsourceibias.n210 0.189894
R21502 commonsourceibias.n237 commonsourceibias.n210 0.189894
R21503 commonsourceibias.n314 commonsourceibias.n208 0.189894
R21504 commonsourceibias.n320 commonsourceibias.n208 0.189894
R21505 commonsourceibias.n321 commonsourceibias.n320 0.189894
R21506 commonsourceibias.n322 commonsourceibias.n321 0.189894
R21507 commonsourceibias.n322 commonsourceibias.n206 0.189894
R21508 commonsourceibias.n327 commonsourceibias.n206 0.189894
R21509 commonsourceibias.n328 commonsourceibias.n327 0.189894
R21510 commonsourceibias.n329 commonsourceibias.n328 0.189894
R21511 commonsourceibias.n329 commonsourceibias.n204 0.189894
R21512 commonsourceibias.n334 commonsourceibias.n204 0.189894
R21513 commonsourceibias.n335 commonsourceibias.n334 0.189894
R21514 commonsourceibias.n335 commonsourceibias.n202 0.189894
R21515 commonsourceibias.n359 commonsourceibias.n354 0.189894
R21516 commonsourceibias.n360 commonsourceibias.n359 0.189894
R21517 commonsourceibias.n360 commonsourceibias.n352 0.189894
R21518 commonsourceibias.n364 commonsourceibias.n352 0.189894
R21519 commonsourceibias.n365 commonsourceibias.n364 0.189894
R21520 commonsourceibias.n365 commonsourceibias.n350 0.189894
R21521 commonsourceibias.n369 commonsourceibias.n350 0.189894
R21522 commonsourceibias.n370 commonsourceibias.n369 0.189894
R21523 commonsourceibias.n370 commonsourceibias.n348 0.189894
R21524 commonsourceibias.n375 commonsourceibias.n348 0.189894
R21525 commonsourceibias.n376 commonsourceibias.n375 0.189894
R21526 commonsourceibias.n377 commonsourceibias.n376 0.189894
R21527 commonsourceibias.n377 commonsourceibias.n346 0.189894
R21528 commonsourceibias.n383 commonsourceibias.n346 0.189894
R21529 commonsourceibias.n384 commonsourceibias.n383 0.189894
R21530 commonsourceibias.n385 commonsourceibias.n384 0.189894
R21531 commonsourceibias.n385 commonsourceibias.n344 0.189894
R21532 commonsourceibias.n390 commonsourceibias.n344 0.189894
R21533 commonsourceibias.n391 commonsourceibias.n390 0.189894
R21534 commonsourceibias.n392 commonsourceibias.n391 0.189894
R21535 commonsourceibias.n392 commonsourceibias.n342 0.189894
R21536 commonsourceibias.n397 commonsourceibias.n342 0.189894
R21537 commonsourceibias.n398 commonsourceibias.n397 0.189894
R21538 commonsourceibias.n398 commonsourceibias.n340 0.189894
R21539 commonsourceibias.n112 commonsourceibias.n111 0.170955
R21540 commonsourceibias.n113 commonsourceibias.n112 0.170955
R21541 commonsourceibias.n313 commonsourceibias.n237 0.170955
R21542 commonsourceibias.n314 commonsourceibias.n313 0.170955
R21543 plus.n61 plus.t11 251.488
R21544 plus.n12 plus.t14 251.488
R21545 plus.n100 plus.t1 243.97
R21546 plus.n96 plus.t23 231.093
R21547 plus.n47 plus.t6 231.093
R21548 plus.n100 plus.n99 223.454
R21549 plus.n102 plus.n101 223.454
R21550 plus.n60 plus.t5 187.445
R21551 plus.n65 plus.t21 187.445
R21552 plus.n71 plus.t20 187.445
R21553 plus.n56 plus.t16 187.445
R21554 plus.n54 plus.t17 187.445
R21555 plus.n83 plus.t13 187.445
R21556 plus.n89 plus.t15 187.445
R21557 plus.n50 plus.t10 187.445
R21558 plus.n1 plus.t12 187.445
R21559 plus.n40 plus.t8 187.445
R21560 plus.n34 plus.t7 187.445
R21561 plus.n5 plus.t19 187.445
R21562 plus.n7 plus.t18 187.445
R21563 plus.n22 plus.t24 187.445
R21564 plus.n16 plus.t22 187.445
R21565 plus.n11 plus.t9 187.445
R21566 plus.n97 plus.n96 161.3
R21567 plus.n95 plus.n49 161.3
R21568 plus.n94 plus.n93 161.3
R21569 plus.n92 plus.n91 161.3
R21570 plus.n90 plus.n51 161.3
R21571 plus.n88 plus.n87 161.3
R21572 plus.n86 plus.n52 161.3
R21573 plus.n85 plus.n84 161.3
R21574 plus.n82 plus.n53 161.3
R21575 plus.n81 plus.n80 161.3
R21576 plus.n79 plus.n78 161.3
R21577 plus.n77 plus.n55 161.3
R21578 plus.n76 plus.n75 161.3
R21579 plus.n74 plus.n73 161.3
R21580 plus.n72 plus.n57 161.3
R21581 plus.n70 plus.n69 161.3
R21582 plus.n68 plus.n58 161.3
R21583 plus.n67 plus.n66 161.3
R21584 plus.n64 plus.n59 161.3
R21585 plus.n63 plus.n62 161.3
R21586 plus.n14 plus.n13 161.3
R21587 plus.n15 plus.n10 161.3
R21588 plus.n18 plus.n17 161.3
R21589 plus.n19 plus.n9 161.3
R21590 plus.n21 plus.n20 161.3
R21591 plus.n23 plus.n8 161.3
R21592 plus.n25 plus.n24 161.3
R21593 plus.n27 plus.n26 161.3
R21594 plus.n28 plus.n6 161.3
R21595 plus.n30 plus.n29 161.3
R21596 plus.n32 plus.n31 161.3
R21597 plus.n33 plus.n4 161.3
R21598 plus.n36 plus.n35 161.3
R21599 plus.n37 plus.n3 161.3
R21600 plus.n39 plus.n38 161.3
R21601 plus.n41 plus.n2 161.3
R21602 plus.n43 plus.n42 161.3
R21603 plus.n45 plus.n44 161.3
R21604 plus.n46 plus.n0 161.3
R21605 plus.n48 plus.n47 161.3
R21606 plus.n64 plus.n63 56.5617
R21607 plus.n91 plus.n90 56.5617
R21608 plus.n42 plus.n41 56.5617
R21609 plus.n15 plus.n14 56.5617
R21610 plus.n73 plus.n72 56.5617
R21611 plus.n82 plus.n81 56.5617
R21612 plus.n33 plus.n32 56.5617
R21613 plus.n24 plus.n23 56.5617
R21614 plus.n95 plus.n94 48.3272
R21615 plus.n46 plus.n45 48.3272
R21616 plus.n70 plus.n58 44.4521
R21617 plus.n84 plus.n52 44.4521
R21618 plus.n35 plus.n3 44.4521
R21619 plus.n21 plus.n9 44.4521
R21620 plus.n62 plus.n61 43.0014
R21621 plus.n13 plus.n12 43.0014
R21622 plus.n77 plus.n76 40.577
R21623 plus.n78 plus.n77 40.577
R21624 plus.n29 plus.n28 40.577
R21625 plus.n28 plus.n27 40.577
R21626 plus.n61 plus.n60 39.4345
R21627 plus.n12 plus.n11 39.4345
R21628 plus.n66 plus.n58 36.702
R21629 plus.n88 plus.n52 36.702
R21630 plus.n39 plus.n3 36.702
R21631 plus.n17 plus.n9 36.702
R21632 plus.n98 plus.n97 33.3471
R21633 plus.n65 plus.n64 20.9036
R21634 plus.n90 plus.n89 20.9036
R21635 plus.n41 plus.n40 20.9036
R21636 plus.n16 plus.n15 20.9036
R21637 plus.n99 plus.t2 19.8005
R21638 plus.n99 plus.t4 19.8005
R21639 plus.n101 plus.t0 19.8005
R21640 plus.n101 plus.t3 19.8005
R21641 plus.n73 plus.n56 18.9362
R21642 plus.n81 plus.n54 18.9362
R21643 plus.n32 plus.n5 18.9362
R21644 plus.n24 plus.n7 18.9362
R21645 plus.n72 plus.n71 16.9689
R21646 plus.n83 plus.n82 16.9689
R21647 plus.n34 plus.n33 16.9689
R21648 plus.n23 plus.n22 16.9689
R21649 plus.n63 plus.n60 15.0015
R21650 plus.n91 plus.n50 15.0015
R21651 plus.n42 plus.n1 15.0015
R21652 plus.n14 plus.n11 15.0015
R21653 plus plus.n103 14.2496
R21654 plus.n96 plus.n95 12.4157
R21655 plus.n47 plus.n46 12.4157
R21656 plus.n98 plus.n48 11.9418
R21657 plus.n94 plus.n50 9.59132
R21658 plus.n45 plus.n1 9.59132
R21659 plus.n71 plus.n70 7.62397
R21660 plus.n84 plus.n83 7.62397
R21661 plus.n35 plus.n34 7.62397
R21662 plus.n22 plus.n21 7.62397
R21663 plus.n76 plus.n56 5.65662
R21664 plus.n78 plus.n54 5.65662
R21665 plus.n29 plus.n5 5.65662
R21666 plus.n27 plus.n7 5.65662
R21667 plus.n103 plus.n102 5.40567
R21668 plus.n66 plus.n65 3.68928
R21669 plus.n89 plus.n88 3.68928
R21670 plus.n40 plus.n39 3.68928
R21671 plus.n17 plus.n16 3.68928
R21672 plus.n103 plus.n98 1.188
R21673 plus.n102 plus.n100 0.716017
R21674 plus.n62 plus.n59 0.189894
R21675 plus.n67 plus.n59 0.189894
R21676 plus.n68 plus.n67 0.189894
R21677 plus.n69 plus.n68 0.189894
R21678 plus.n69 plus.n57 0.189894
R21679 plus.n74 plus.n57 0.189894
R21680 plus.n75 plus.n74 0.189894
R21681 plus.n75 plus.n55 0.189894
R21682 plus.n79 plus.n55 0.189894
R21683 plus.n80 plus.n79 0.189894
R21684 plus.n80 plus.n53 0.189894
R21685 plus.n85 plus.n53 0.189894
R21686 plus.n86 plus.n85 0.189894
R21687 plus.n87 plus.n86 0.189894
R21688 plus.n87 plus.n51 0.189894
R21689 plus.n92 plus.n51 0.189894
R21690 plus.n93 plus.n92 0.189894
R21691 plus.n93 plus.n49 0.189894
R21692 plus.n97 plus.n49 0.189894
R21693 plus.n48 plus.n0 0.189894
R21694 plus.n44 plus.n0 0.189894
R21695 plus.n44 plus.n43 0.189894
R21696 plus.n43 plus.n2 0.189894
R21697 plus.n38 plus.n2 0.189894
R21698 plus.n38 plus.n37 0.189894
R21699 plus.n37 plus.n36 0.189894
R21700 plus.n36 plus.n4 0.189894
R21701 plus.n31 plus.n4 0.189894
R21702 plus.n31 plus.n30 0.189894
R21703 plus.n30 plus.n6 0.189894
R21704 plus.n26 plus.n6 0.189894
R21705 plus.n26 plus.n25 0.189894
R21706 plus.n25 plus.n8 0.189894
R21707 plus.n20 plus.n8 0.189894
R21708 plus.n20 plus.n19 0.189894
R21709 plus.n19 plus.n18 0.189894
R21710 plus.n18 plus.n10 0.189894
R21711 plus.n13 plus.n10 0.189894
R21712 a_n2903_n3924.n18 a_n2903_n3924.t2 214.624
R21713 a_n2903_n3924.n1 a_n2903_n3924.t5 214.321
R21714 a_n2903_n3924.n12 a_n2903_n3924.t1 214.321
R21715 a_n2903_n3924.n13 a_n2903_n3924.t0 214.321
R21716 a_n2903_n3924.n14 a_n2903_n3924.t34 214.321
R21717 a_n2903_n3924.n15 a_n2903_n3924.t47 214.321
R21718 a_n2903_n3924.n16 a_n2903_n3924.t3 214.321
R21719 a_n2903_n3924.n17 a_n2903_n3924.t4 214.321
R21720 a_n2903_n3924.n0 a_n2903_n3924.t27 55.8337
R21721 a_n2903_n3924.n2 a_n2903_n3924.t44 55.8337
R21722 a_n2903_n3924.n11 a_n2903_n3924.t35 55.8337
R21723 a_n2903_n3924.n41 a_n2903_n3924.t15 55.8335
R21724 a_n2903_n3924.n39 a_n2903_n3924.t11 55.8335
R21725 a_n2903_n3924.n30 a_n2903_n3924.t41 55.8335
R21726 a_n2903_n3924.n29 a_n2903_n3924.t24 55.8335
R21727 a_n2903_n3924.n20 a_n2903_n3924.t32 55.8335
R21728 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0052
R21729 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0052
R21730 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0052
R21731 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R21732 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R21733 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R21734 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R21735 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R21736 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R21737 a_n2903_n3924.n34 a_n2903_n3924.n33 53.0051
R21738 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R21739 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R21740 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R21741 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R21742 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0051
R21743 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R21744 a_n2903_n3924.n19 a_n2903_n3924.n11 12.2417
R21745 a_n2903_n3924.n41 a_n2903_n3924.n40 12.2417
R21746 a_n2903_n3924.n20 a_n2903_n3924.n19 5.16214
R21747 a_n2903_n3924.n40 a_n2903_n3924.n39 5.16214
R21748 a_n2903_n3924.n42 a_n2903_n3924.t23 2.82907
R21749 a_n2903_n3924.n42 a_n2903_n3924.t28 2.82907
R21750 a_n2903_n3924.n44 a_n2903_n3924.t21 2.82907
R21751 a_n2903_n3924.n44 a_n2903_n3924.t25 2.82907
R21752 a_n2903_n3924.n46 a_n2903_n3924.t18 2.82907
R21753 a_n2903_n3924.n46 a_n2903_n3924.t22 2.82907
R21754 a_n2903_n3924.n3 a_n2903_n3924.t13 2.82907
R21755 a_n2903_n3924.n3 a_n2903_n3924.t38 2.82907
R21756 a_n2903_n3924.n5 a_n2903_n3924.t8 2.82907
R21757 a_n2903_n3924.n5 a_n2903_n3924.t9 2.82907
R21758 a_n2903_n3924.n7 a_n2903_n3924.t42 2.82907
R21759 a_n2903_n3924.n7 a_n2903_n3924.t46 2.82907
R21760 a_n2903_n3924.n9 a_n2903_n3924.t36 2.82907
R21761 a_n2903_n3924.n9 a_n2903_n3924.t39 2.82907
R21762 a_n2903_n3924.n37 a_n2903_n3924.t37 2.82907
R21763 a_n2903_n3924.n37 a_n2903_n3924.t12 2.82907
R21764 a_n2903_n3924.n35 a_n2903_n3924.t45 2.82907
R21765 a_n2903_n3924.n35 a_n2903_n3924.t40 2.82907
R21766 a_n2903_n3924.n33 a_n2903_n3924.t7 2.82907
R21767 a_n2903_n3924.n33 a_n2903_n3924.t43 2.82907
R21768 a_n2903_n3924.n31 a_n2903_n3924.t10 2.82907
R21769 a_n2903_n3924.n31 a_n2903_n3924.t6 2.82907
R21770 a_n2903_n3924.n27 a_n2903_n3924.t16 2.82907
R21771 a_n2903_n3924.n27 a_n2903_n3924.t29 2.82907
R21772 a_n2903_n3924.n25 a_n2903_n3924.t20 2.82907
R21773 a_n2903_n3924.n25 a_n2903_n3924.t14 2.82907
R21774 a_n2903_n3924.n23 a_n2903_n3924.t31 2.82907
R21775 a_n2903_n3924.n23 a_n2903_n3924.t19 2.82907
R21776 a_n2903_n3924.n21 a_n2903_n3924.t26 2.82907
R21777 a_n2903_n3924.n21 a_n2903_n3924.t30 2.82907
R21778 a_n2903_n3924.t33 a_n2903_n3924.n49 2.82907
R21779 a_n2903_n3924.n49 a_n2903_n3924.t17 2.82907
R21780 a_n2903_n3924.n40 a_n2903_n3924.n1 2.18441
R21781 a_n2903_n3924.n19 a_n2903_n3924.n18 1.95694
R21782 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R21783 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R21784 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R21785 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R21786 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R21787 a_n2903_n3924.n12 a_n2903_n3924.n1 0.672012
R21788 a_n2903_n3924.n22 a_n2903_n3924.n20 0.530672
R21789 a_n2903_n3924.n24 a_n2903_n3924.n22 0.530672
R21790 a_n2903_n3924.n26 a_n2903_n3924.n24 0.530672
R21791 a_n2903_n3924.n28 a_n2903_n3924.n26 0.530672
R21792 a_n2903_n3924.n29 a_n2903_n3924.n28 0.530672
R21793 a_n2903_n3924.n32 a_n2903_n3924.n30 0.530672
R21794 a_n2903_n3924.n34 a_n2903_n3924.n32 0.530672
R21795 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R21796 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R21797 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R21798 a_n2903_n3924.n11 a_n2903_n3924.n10 0.530672
R21799 a_n2903_n3924.n10 a_n2903_n3924.n8 0.530672
R21800 a_n2903_n3924.n8 a_n2903_n3924.n6 0.530672
R21801 a_n2903_n3924.n6 a_n2903_n3924.n4 0.530672
R21802 a_n2903_n3924.n4 a_n2903_n3924.n2 0.530672
R21803 a_n2903_n3924.n48 a_n2903_n3924.n0 0.530672
R21804 a_n2903_n3924.n48 a_n2903_n3924.n47 0.530672
R21805 a_n2903_n3924.n47 a_n2903_n3924.n45 0.530672
R21806 a_n2903_n3924.n45 a_n2903_n3924.n43 0.530672
R21807 a_n2903_n3924.n43 a_n2903_n3924.n41 0.530672
R21808 a_n2903_n3924.n18 a_n2903_n3924.n17 0.370413
R21809 a_n2903_n3924.n30 a_n2903_n3924.n29 0.235414
R21810 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R21811 outputibias.n27 outputibias.n1 289.615
R21812 outputibias.n58 outputibias.n32 289.615
R21813 outputibias.n90 outputibias.n64 289.615
R21814 outputibias.n122 outputibias.n96 289.615
R21815 outputibias.n28 outputibias.n27 185
R21816 outputibias.n26 outputibias.n25 185
R21817 outputibias.n5 outputibias.n4 185
R21818 outputibias.n20 outputibias.n19 185
R21819 outputibias.n18 outputibias.n17 185
R21820 outputibias.n9 outputibias.n8 185
R21821 outputibias.n12 outputibias.n11 185
R21822 outputibias.n59 outputibias.n58 185
R21823 outputibias.n57 outputibias.n56 185
R21824 outputibias.n36 outputibias.n35 185
R21825 outputibias.n51 outputibias.n50 185
R21826 outputibias.n49 outputibias.n48 185
R21827 outputibias.n40 outputibias.n39 185
R21828 outputibias.n43 outputibias.n42 185
R21829 outputibias.n91 outputibias.n90 185
R21830 outputibias.n89 outputibias.n88 185
R21831 outputibias.n68 outputibias.n67 185
R21832 outputibias.n83 outputibias.n82 185
R21833 outputibias.n81 outputibias.n80 185
R21834 outputibias.n72 outputibias.n71 185
R21835 outputibias.n75 outputibias.n74 185
R21836 outputibias.n123 outputibias.n122 185
R21837 outputibias.n121 outputibias.n120 185
R21838 outputibias.n100 outputibias.n99 185
R21839 outputibias.n115 outputibias.n114 185
R21840 outputibias.n113 outputibias.n112 185
R21841 outputibias.n104 outputibias.n103 185
R21842 outputibias.n107 outputibias.n106 185
R21843 outputibias.n0 outputibias.t8 178.945
R21844 outputibias.n133 outputibias.t10 177.018
R21845 outputibias.n132 outputibias.t11 177.018
R21846 outputibias.n0 outputibias.t9 177.018
R21847 outputibias.t5 outputibias.n10 147.661
R21848 outputibias.t7 outputibias.n41 147.661
R21849 outputibias.t1 outputibias.n73 147.661
R21850 outputibias.t3 outputibias.n105 147.661
R21851 outputibias.n128 outputibias.t4 132.363
R21852 outputibias.n128 outputibias.t6 130.436
R21853 outputibias.n129 outputibias.t0 130.436
R21854 outputibias.n130 outputibias.t2 130.436
R21855 outputibias.n27 outputibias.n26 104.615
R21856 outputibias.n26 outputibias.n4 104.615
R21857 outputibias.n19 outputibias.n4 104.615
R21858 outputibias.n19 outputibias.n18 104.615
R21859 outputibias.n18 outputibias.n8 104.615
R21860 outputibias.n11 outputibias.n8 104.615
R21861 outputibias.n58 outputibias.n57 104.615
R21862 outputibias.n57 outputibias.n35 104.615
R21863 outputibias.n50 outputibias.n35 104.615
R21864 outputibias.n50 outputibias.n49 104.615
R21865 outputibias.n49 outputibias.n39 104.615
R21866 outputibias.n42 outputibias.n39 104.615
R21867 outputibias.n90 outputibias.n89 104.615
R21868 outputibias.n89 outputibias.n67 104.615
R21869 outputibias.n82 outputibias.n67 104.615
R21870 outputibias.n82 outputibias.n81 104.615
R21871 outputibias.n81 outputibias.n71 104.615
R21872 outputibias.n74 outputibias.n71 104.615
R21873 outputibias.n122 outputibias.n121 104.615
R21874 outputibias.n121 outputibias.n99 104.615
R21875 outputibias.n114 outputibias.n99 104.615
R21876 outputibias.n114 outputibias.n113 104.615
R21877 outputibias.n113 outputibias.n103 104.615
R21878 outputibias.n106 outputibias.n103 104.615
R21879 outputibias.n63 outputibias.n31 95.6354
R21880 outputibias.n63 outputibias.n62 94.6732
R21881 outputibias.n95 outputibias.n94 94.6732
R21882 outputibias.n127 outputibias.n126 94.6732
R21883 outputibias.n11 outputibias.t5 52.3082
R21884 outputibias.n42 outputibias.t7 52.3082
R21885 outputibias.n74 outputibias.t1 52.3082
R21886 outputibias.n106 outputibias.t3 52.3082
R21887 outputibias.n12 outputibias.n10 15.6674
R21888 outputibias.n43 outputibias.n41 15.6674
R21889 outputibias.n75 outputibias.n73 15.6674
R21890 outputibias.n107 outputibias.n105 15.6674
R21891 outputibias.n13 outputibias.n9 12.8005
R21892 outputibias.n44 outputibias.n40 12.8005
R21893 outputibias.n76 outputibias.n72 12.8005
R21894 outputibias.n108 outputibias.n104 12.8005
R21895 outputibias.n17 outputibias.n16 12.0247
R21896 outputibias.n48 outputibias.n47 12.0247
R21897 outputibias.n80 outputibias.n79 12.0247
R21898 outputibias.n112 outputibias.n111 12.0247
R21899 outputibias.n20 outputibias.n7 11.249
R21900 outputibias.n51 outputibias.n38 11.249
R21901 outputibias.n83 outputibias.n70 11.249
R21902 outputibias.n115 outputibias.n102 11.249
R21903 outputibias.n21 outputibias.n5 10.4732
R21904 outputibias.n52 outputibias.n36 10.4732
R21905 outputibias.n84 outputibias.n68 10.4732
R21906 outputibias.n116 outputibias.n100 10.4732
R21907 outputibias.n25 outputibias.n24 9.69747
R21908 outputibias.n56 outputibias.n55 9.69747
R21909 outputibias.n88 outputibias.n87 9.69747
R21910 outputibias.n120 outputibias.n119 9.69747
R21911 outputibias.n31 outputibias.n30 9.45567
R21912 outputibias.n62 outputibias.n61 9.45567
R21913 outputibias.n94 outputibias.n93 9.45567
R21914 outputibias.n126 outputibias.n125 9.45567
R21915 outputibias.n30 outputibias.n29 9.3005
R21916 outputibias.n3 outputibias.n2 9.3005
R21917 outputibias.n24 outputibias.n23 9.3005
R21918 outputibias.n22 outputibias.n21 9.3005
R21919 outputibias.n7 outputibias.n6 9.3005
R21920 outputibias.n16 outputibias.n15 9.3005
R21921 outputibias.n14 outputibias.n13 9.3005
R21922 outputibias.n61 outputibias.n60 9.3005
R21923 outputibias.n34 outputibias.n33 9.3005
R21924 outputibias.n55 outputibias.n54 9.3005
R21925 outputibias.n53 outputibias.n52 9.3005
R21926 outputibias.n38 outputibias.n37 9.3005
R21927 outputibias.n47 outputibias.n46 9.3005
R21928 outputibias.n45 outputibias.n44 9.3005
R21929 outputibias.n93 outputibias.n92 9.3005
R21930 outputibias.n66 outputibias.n65 9.3005
R21931 outputibias.n87 outputibias.n86 9.3005
R21932 outputibias.n85 outputibias.n84 9.3005
R21933 outputibias.n70 outputibias.n69 9.3005
R21934 outputibias.n79 outputibias.n78 9.3005
R21935 outputibias.n77 outputibias.n76 9.3005
R21936 outputibias.n125 outputibias.n124 9.3005
R21937 outputibias.n98 outputibias.n97 9.3005
R21938 outputibias.n119 outputibias.n118 9.3005
R21939 outputibias.n117 outputibias.n116 9.3005
R21940 outputibias.n102 outputibias.n101 9.3005
R21941 outputibias.n111 outputibias.n110 9.3005
R21942 outputibias.n109 outputibias.n108 9.3005
R21943 outputibias.n28 outputibias.n3 8.92171
R21944 outputibias.n59 outputibias.n34 8.92171
R21945 outputibias.n91 outputibias.n66 8.92171
R21946 outputibias.n123 outputibias.n98 8.92171
R21947 outputibias.n29 outputibias.n1 8.14595
R21948 outputibias.n60 outputibias.n32 8.14595
R21949 outputibias.n92 outputibias.n64 8.14595
R21950 outputibias.n124 outputibias.n96 8.14595
R21951 outputibias.n31 outputibias.n1 5.81868
R21952 outputibias.n62 outputibias.n32 5.81868
R21953 outputibias.n94 outputibias.n64 5.81868
R21954 outputibias.n126 outputibias.n96 5.81868
R21955 outputibias.n131 outputibias.n130 5.20947
R21956 outputibias.n29 outputibias.n28 5.04292
R21957 outputibias.n60 outputibias.n59 5.04292
R21958 outputibias.n92 outputibias.n91 5.04292
R21959 outputibias.n124 outputibias.n123 5.04292
R21960 outputibias.n131 outputibias.n127 4.42209
R21961 outputibias.n14 outputibias.n10 4.38594
R21962 outputibias.n45 outputibias.n41 4.38594
R21963 outputibias.n77 outputibias.n73 4.38594
R21964 outputibias.n109 outputibias.n105 4.38594
R21965 outputibias.n132 outputibias.n131 4.28454
R21966 outputibias.n25 outputibias.n3 4.26717
R21967 outputibias.n56 outputibias.n34 4.26717
R21968 outputibias.n88 outputibias.n66 4.26717
R21969 outputibias.n120 outputibias.n98 4.26717
R21970 outputibias.n24 outputibias.n5 3.49141
R21971 outputibias.n55 outputibias.n36 3.49141
R21972 outputibias.n87 outputibias.n68 3.49141
R21973 outputibias.n119 outputibias.n100 3.49141
R21974 outputibias.n21 outputibias.n20 2.71565
R21975 outputibias.n52 outputibias.n51 2.71565
R21976 outputibias.n84 outputibias.n83 2.71565
R21977 outputibias.n116 outputibias.n115 2.71565
R21978 outputibias.n17 outputibias.n7 1.93989
R21979 outputibias.n48 outputibias.n38 1.93989
R21980 outputibias.n80 outputibias.n70 1.93989
R21981 outputibias.n112 outputibias.n102 1.93989
R21982 outputibias.n130 outputibias.n129 1.9266
R21983 outputibias.n129 outputibias.n128 1.9266
R21984 outputibias.n133 outputibias.n132 1.92658
R21985 outputibias.n134 outputibias.n133 1.29913
R21986 outputibias.n16 outputibias.n9 1.16414
R21987 outputibias.n47 outputibias.n40 1.16414
R21988 outputibias.n79 outputibias.n72 1.16414
R21989 outputibias.n111 outputibias.n104 1.16414
R21990 outputibias.n127 outputibias.n95 0.962709
R21991 outputibias.n95 outputibias.n63 0.962709
R21992 outputibias.n13 outputibias.n12 0.388379
R21993 outputibias.n44 outputibias.n43 0.388379
R21994 outputibias.n76 outputibias.n75 0.388379
R21995 outputibias.n108 outputibias.n107 0.388379
R21996 outputibias.n134 outputibias.n0 0.337251
R21997 outputibias outputibias.n134 0.302375
R21998 outputibias.n30 outputibias.n2 0.155672
R21999 outputibias.n23 outputibias.n2 0.155672
R22000 outputibias.n23 outputibias.n22 0.155672
R22001 outputibias.n22 outputibias.n6 0.155672
R22002 outputibias.n15 outputibias.n6 0.155672
R22003 outputibias.n15 outputibias.n14 0.155672
R22004 outputibias.n61 outputibias.n33 0.155672
R22005 outputibias.n54 outputibias.n33 0.155672
R22006 outputibias.n54 outputibias.n53 0.155672
R22007 outputibias.n53 outputibias.n37 0.155672
R22008 outputibias.n46 outputibias.n37 0.155672
R22009 outputibias.n46 outputibias.n45 0.155672
R22010 outputibias.n93 outputibias.n65 0.155672
R22011 outputibias.n86 outputibias.n65 0.155672
R22012 outputibias.n86 outputibias.n85 0.155672
R22013 outputibias.n85 outputibias.n69 0.155672
R22014 outputibias.n78 outputibias.n69 0.155672
R22015 outputibias.n78 outputibias.n77 0.155672
R22016 outputibias.n125 outputibias.n97 0.155672
R22017 outputibias.n118 outputibias.n97 0.155672
R22018 outputibias.n118 outputibias.n117 0.155672
R22019 outputibias.n117 outputibias.n101 0.155672
R22020 outputibias.n110 outputibias.n101 0.155672
R22021 outputibias.n110 outputibias.n109 0.155672
R22022 output.n41 output.n15 289.615
R22023 output.n72 output.n46 289.615
R22024 output.n104 output.n78 289.615
R22025 output.n136 output.n110 289.615
R22026 output.n77 output.n45 197.26
R22027 output.n77 output.n76 196.298
R22028 output.n109 output.n108 196.298
R22029 output.n141 output.n140 196.298
R22030 output.n42 output.n41 185
R22031 output.n40 output.n39 185
R22032 output.n19 output.n18 185
R22033 output.n34 output.n33 185
R22034 output.n32 output.n31 185
R22035 output.n23 output.n22 185
R22036 output.n26 output.n25 185
R22037 output.n73 output.n72 185
R22038 output.n71 output.n70 185
R22039 output.n50 output.n49 185
R22040 output.n65 output.n64 185
R22041 output.n63 output.n62 185
R22042 output.n54 output.n53 185
R22043 output.n57 output.n56 185
R22044 output.n105 output.n104 185
R22045 output.n103 output.n102 185
R22046 output.n82 output.n81 185
R22047 output.n97 output.n96 185
R22048 output.n95 output.n94 185
R22049 output.n86 output.n85 185
R22050 output.n89 output.n88 185
R22051 output.n137 output.n136 185
R22052 output.n135 output.n134 185
R22053 output.n114 output.n113 185
R22054 output.n129 output.n128 185
R22055 output.n127 output.n126 185
R22056 output.n118 output.n117 185
R22057 output.n121 output.n120 185
R22058 output.t19 output.n24 147.661
R22059 output.t18 output.n55 147.661
R22060 output.t17 output.n87 147.661
R22061 output.t16 output.n119 147.661
R22062 output.n41 output.n40 104.615
R22063 output.n40 output.n18 104.615
R22064 output.n33 output.n18 104.615
R22065 output.n33 output.n32 104.615
R22066 output.n32 output.n22 104.615
R22067 output.n25 output.n22 104.615
R22068 output.n72 output.n71 104.615
R22069 output.n71 output.n49 104.615
R22070 output.n64 output.n49 104.615
R22071 output.n64 output.n63 104.615
R22072 output.n63 output.n53 104.615
R22073 output.n56 output.n53 104.615
R22074 output.n104 output.n103 104.615
R22075 output.n103 output.n81 104.615
R22076 output.n96 output.n81 104.615
R22077 output.n96 output.n95 104.615
R22078 output.n95 output.n85 104.615
R22079 output.n88 output.n85 104.615
R22080 output.n136 output.n135 104.615
R22081 output.n135 output.n113 104.615
R22082 output.n128 output.n113 104.615
R22083 output.n128 output.n127 104.615
R22084 output.n127 output.n117 104.615
R22085 output.n120 output.n117 104.615
R22086 output.n1 output.t12 77.056
R22087 output.n14 output.t14 76.6694
R22088 output.n1 output.n0 72.7095
R22089 output.n3 output.n2 72.7095
R22090 output.n5 output.n4 72.7095
R22091 output.n7 output.n6 72.7095
R22092 output.n9 output.n8 72.7095
R22093 output.n11 output.n10 72.7095
R22094 output.n13 output.n12 72.7095
R22095 output.n25 output.t19 52.3082
R22096 output.n56 output.t18 52.3082
R22097 output.n88 output.t17 52.3082
R22098 output.n120 output.t16 52.3082
R22099 output.n26 output.n24 15.6674
R22100 output.n57 output.n55 15.6674
R22101 output.n89 output.n87 15.6674
R22102 output.n121 output.n119 15.6674
R22103 output.n27 output.n23 12.8005
R22104 output.n58 output.n54 12.8005
R22105 output.n90 output.n86 12.8005
R22106 output.n122 output.n118 12.8005
R22107 output.n31 output.n30 12.0247
R22108 output.n62 output.n61 12.0247
R22109 output.n94 output.n93 12.0247
R22110 output.n126 output.n125 12.0247
R22111 output.n34 output.n21 11.249
R22112 output.n65 output.n52 11.249
R22113 output.n97 output.n84 11.249
R22114 output.n129 output.n116 11.249
R22115 output.n35 output.n19 10.4732
R22116 output.n66 output.n50 10.4732
R22117 output.n98 output.n82 10.4732
R22118 output.n130 output.n114 10.4732
R22119 output.n39 output.n38 9.69747
R22120 output.n70 output.n69 9.69747
R22121 output.n102 output.n101 9.69747
R22122 output.n134 output.n133 9.69747
R22123 output.n45 output.n44 9.45567
R22124 output.n76 output.n75 9.45567
R22125 output.n108 output.n107 9.45567
R22126 output.n140 output.n139 9.45567
R22127 output.n44 output.n43 9.3005
R22128 output.n17 output.n16 9.3005
R22129 output.n38 output.n37 9.3005
R22130 output.n36 output.n35 9.3005
R22131 output.n21 output.n20 9.3005
R22132 output.n30 output.n29 9.3005
R22133 output.n28 output.n27 9.3005
R22134 output.n75 output.n74 9.3005
R22135 output.n48 output.n47 9.3005
R22136 output.n69 output.n68 9.3005
R22137 output.n67 output.n66 9.3005
R22138 output.n52 output.n51 9.3005
R22139 output.n61 output.n60 9.3005
R22140 output.n59 output.n58 9.3005
R22141 output.n107 output.n106 9.3005
R22142 output.n80 output.n79 9.3005
R22143 output.n101 output.n100 9.3005
R22144 output.n99 output.n98 9.3005
R22145 output.n84 output.n83 9.3005
R22146 output.n93 output.n92 9.3005
R22147 output.n91 output.n90 9.3005
R22148 output.n139 output.n138 9.3005
R22149 output.n112 output.n111 9.3005
R22150 output.n133 output.n132 9.3005
R22151 output.n131 output.n130 9.3005
R22152 output.n116 output.n115 9.3005
R22153 output.n125 output.n124 9.3005
R22154 output.n123 output.n122 9.3005
R22155 output.n42 output.n17 8.92171
R22156 output.n73 output.n48 8.92171
R22157 output.n105 output.n80 8.92171
R22158 output.n137 output.n112 8.92171
R22159 output output.n141 8.15037
R22160 output.n43 output.n15 8.14595
R22161 output.n74 output.n46 8.14595
R22162 output.n106 output.n78 8.14595
R22163 output.n138 output.n110 8.14595
R22164 output.n45 output.n15 5.81868
R22165 output.n76 output.n46 5.81868
R22166 output.n108 output.n78 5.81868
R22167 output.n140 output.n110 5.81868
R22168 output.n43 output.n42 5.04292
R22169 output.n74 output.n73 5.04292
R22170 output.n106 output.n105 5.04292
R22171 output.n138 output.n137 5.04292
R22172 output.n28 output.n24 4.38594
R22173 output.n59 output.n55 4.38594
R22174 output.n91 output.n87 4.38594
R22175 output.n123 output.n119 4.38594
R22176 output.n39 output.n17 4.26717
R22177 output.n70 output.n48 4.26717
R22178 output.n102 output.n80 4.26717
R22179 output.n134 output.n112 4.26717
R22180 output.n0 output.t3 3.9605
R22181 output.n0 output.t7 3.9605
R22182 output.n2 output.t10 3.9605
R22183 output.n2 output.t15 3.9605
R22184 output.n4 output.t0 3.9605
R22185 output.n4 output.t5 3.9605
R22186 output.n6 output.t9 3.9605
R22187 output.n6 output.t1 3.9605
R22188 output.n8 output.t4 3.9605
R22189 output.n8 output.t2 3.9605
R22190 output.n10 output.t8 3.9605
R22191 output.n10 output.t11 3.9605
R22192 output.n12 output.t13 3.9605
R22193 output.n12 output.t6 3.9605
R22194 output.n38 output.n19 3.49141
R22195 output.n69 output.n50 3.49141
R22196 output.n101 output.n82 3.49141
R22197 output.n133 output.n114 3.49141
R22198 output.n35 output.n34 2.71565
R22199 output.n66 output.n65 2.71565
R22200 output.n98 output.n97 2.71565
R22201 output.n130 output.n129 2.71565
R22202 output.n31 output.n21 1.93989
R22203 output.n62 output.n52 1.93989
R22204 output.n94 output.n84 1.93989
R22205 output.n126 output.n116 1.93989
R22206 output.n30 output.n23 1.16414
R22207 output.n61 output.n54 1.16414
R22208 output.n93 output.n86 1.16414
R22209 output.n125 output.n118 1.16414
R22210 output.n141 output.n109 0.962709
R22211 output.n109 output.n77 0.962709
R22212 output.n27 output.n26 0.388379
R22213 output.n58 output.n57 0.388379
R22214 output.n90 output.n89 0.388379
R22215 output.n122 output.n121 0.388379
R22216 output.n14 output.n13 0.387128
R22217 output.n13 output.n11 0.387128
R22218 output.n11 output.n9 0.387128
R22219 output.n9 output.n7 0.387128
R22220 output.n7 output.n5 0.387128
R22221 output.n5 output.n3 0.387128
R22222 output.n3 output.n1 0.387128
R22223 output.n44 output.n16 0.155672
R22224 output.n37 output.n16 0.155672
R22225 output.n37 output.n36 0.155672
R22226 output.n36 output.n20 0.155672
R22227 output.n29 output.n20 0.155672
R22228 output.n29 output.n28 0.155672
R22229 output.n75 output.n47 0.155672
R22230 output.n68 output.n47 0.155672
R22231 output.n68 output.n67 0.155672
R22232 output.n67 output.n51 0.155672
R22233 output.n60 output.n51 0.155672
R22234 output.n60 output.n59 0.155672
R22235 output.n107 output.n79 0.155672
R22236 output.n100 output.n79 0.155672
R22237 output.n100 output.n99 0.155672
R22238 output.n99 output.n83 0.155672
R22239 output.n92 output.n83 0.155672
R22240 output.n92 output.n91 0.155672
R22241 output.n139 output.n111 0.155672
R22242 output.n132 output.n111 0.155672
R22243 output.n132 output.n131 0.155672
R22244 output.n131 output.n115 0.155672
R22245 output.n124 output.n115 0.155672
R22246 output.n124 output.n123 0.155672
R22247 output output.n14 0.126227
R22248 a_n2650_8322.n10 a_n2650_8322.t29 74.6477
R22249 a_n2650_8322.n1 a_n2650_8322.t21 74.6477
R22250 a_n2650_8322.n24 a_n2650_8322.t23 74.6474
R22251 a_n2650_8322.n18 a_n2650_8322.t20 74.2899
R22252 a_n2650_8322.n11 a_n2650_8322.t27 74.2899
R22253 a_n2650_8322.n12 a_n2650_8322.t30 74.2899
R22254 a_n2650_8322.n15 a_n2650_8322.t31 74.2899
R22255 a_n2650_8322.n8 a_n2650_8322.t6 74.2899
R22256 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R22257 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R22258 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R22259 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R22260 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R22261 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R22262 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R22263 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R22264 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R22265 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R22266 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R22267 a_n2650_8322.n17 a_n2650_8322.t2 9.58915
R22268 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R22269 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R22270 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R22271 a_n2650_8322.n23 a_n2650_8322.t18 3.61217
R22272 a_n2650_8322.n23 a_n2650_8322.t14 3.61217
R22273 a_n2650_8322.n21 a_n2650_8322.t22 3.61217
R22274 a_n2650_8322.n21 a_n2650_8322.t11 3.61217
R22275 a_n2650_8322.n19 a_n2650_8322.t9 3.61217
R22276 a_n2650_8322.n19 a_n2650_8322.t10 3.61217
R22277 a_n2650_8322.n9 a_n2650_8322.t32 3.61217
R22278 a_n2650_8322.n9 a_n2650_8322.t33 3.61217
R22279 a_n2650_8322.n13 a_n2650_8322.t28 3.61217
R22280 a_n2650_8322.n13 a_n2650_8322.t26 3.61217
R22281 a_n2650_8322.n0 a_n2650_8322.t24 3.61217
R22282 a_n2650_8322.n0 a_n2650_8322.t16 3.61217
R22283 a_n2650_8322.n2 a_n2650_8322.t8 3.61217
R22284 a_n2650_8322.n2 a_n2650_8322.t7 3.61217
R22285 a_n2650_8322.n4 a_n2650_8322.t19 3.61217
R22286 a_n2650_8322.n4 a_n2650_8322.t13 3.61217
R22287 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R22288 a_n2650_8322.n6 a_n2650_8322.t15 3.61217
R22289 a_n2650_8322.n26 a_n2650_8322.t12 3.61217
R22290 a_n2650_8322.t25 a_n2650_8322.n26 3.61217
R22291 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R22292 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R22293 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R22294 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R22295 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R22296 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R22297 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R22298 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R22299 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R22300 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R22301 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R22302 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R22303 a_n2650_8322.t3 a_n2650_8322.t0 0.0788333
R22304 a_n2650_8322.t4 a_n2650_8322.t5 0.0788333
R22305 a_n2650_8322.t2 a_n2650_8322.t1 0.0788333
R22306 a_n2650_8322.t4 a_n2650_8322.t3 0.0318333
R22307 a_n2650_8322.t2 a_n2650_8322.t5 0.0318333
R22308 a_n2650_8322.t0 a_n2650_8322.t5 0.0318333
R22309 a_n2650_8322.t1 a_n2650_8322.t4 0.0318333
R22310 minus.n61 minus.t24 251.488
R22311 minus.n12 minus.t16 251.488
R22312 minus.n102 minus.t4 243.255
R22313 minus.n96 minus.t14 231.093
R22314 minus.n47 minus.t9 231.093
R22315 minus.n101 minus.n99 224.169
R22316 minus.n101 minus.n100 223.454
R22317 minus.n50 minus.t21 187.445
R22318 minus.n89 minus.t18 187.445
R22319 minus.n83 minus.t15 187.445
R22320 minus.n54 minus.t7 187.445
R22321 minus.n56 minus.t6 187.445
R22322 minus.n71 minus.t12 187.445
R22323 minus.n65 minus.t11 187.445
R22324 minus.n60 minus.t19 187.445
R22325 minus.n11 minus.t10 187.445
R22326 minus.n16 minus.t8 187.445
R22327 minus.n22 minus.t5 187.445
R22328 minus.n7 minus.t22 187.445
R22329 minus.n5 minus.t23 187.445
R22330 minus.n34 minus.t17 187.445
R22331 minus.n40 minus.t20 187.445
R22332 minus.n1 minus.t13 187.445
R22333 minus.n63 minus.n62 161.3
R22334 minus.n64 minus.n59 161.3
R22335 minus.n67 minus.n66 161.3
R22336 minus.n68 minus.n58 161.3
R22337 minus.n70 minus.n69 161.3
R22338 minus.n72 minus.n57 161.3
R22339 minus.n74 minus.n73 161.3
R22340 minus.n76 minus.n75 161.3
R22341 minus.n77 minus.n55 161.3
R22342 minus.n79 minus.n78 161.3
R22343 minus.n81 minus.n80 161.3
R22344 minus.n82 minus.n53 161.3
R22345 minus.n85 minus.n84 161.3
R22346 minus.n86 minus.n52 161.3
R22347 minus.n88 minus.n87 161.3
R22348 minus.n90 minus.n51 161.3
R22349 minus.n92 minus.n91 161.3
R22350 minus.n94 minus.n93 161.3
R22351 minus.n95 minus.n49 161.3
R22352 minus.n97 minus.n96 161.3
R22353 minus.n48 minus.n47 161.3
R22354 minus.n46 minus.n0 161.3
R22355 minus.n45 minus.n44 161.3
R22356 minus.n43 minus.n42 161.3
R22357 minus.n41 minus.n2 161.3
R22358 minus.n39 minus.n38 161.3
R22359 minus.n37 minus.n3 161.3
R22360 minus.n36 minus.n35 161.3
R22361 minus.n33 minus.n4 161.3
R22362 minus.n32 minus.n31 161.3
R22363 minus.n30 minus.n29 161.3
R22364 minus.n28 minus.n6 161.3
R22365 minus.n27 minus.n26 161.3
R22366 minus.n25 minus.n24 161.3
R22367 minus.n23 minus.n8 161.3
R22368 minus.n21 minus.n20 161.3
R22369 minus.n19 minus.n9 161.3
R22370 minus.n18 minus.n17 161.3
R22371 minus.n15 minus.n10 161.3
R22372 minus.n14 minus.n13 161.3
R22373 minus.n91 minus.n90 56.5617
R22374 minus.n64 minus.n63 56.5617
R22375 minus.n15 minus.n14 56.5617
R22376 minus.n42 minus.n41 56.5617
R22377 minus.n82 minus.n81 56.5617
R22378 minus.n73 minus.n72 56.5617
R22379 minus.n24 minus.n23 56.5617
R22380 minus.n33 minus.n32 56.5617
R22381 minus.n95 minus.n94 48.3272
R22382 minus.n46 minus.n45 48.3272
R22383 minus.n84 minus.n52 44.4521
R22384 minus.n70 minus.n58 44.4521
R22385 minus.n21 minus.n9 44.4521
R22386 minus.n35 minus.n3 44.4521
R22387 minus.n13 minus.n12 43.0014
R22388 minus.n62 minus.n61 43.0014
R22389 minus.n78 minus.n77 40.577
R22390 minus.n77 minus.n76 40.577
R22391 minus.n28 minus.n27 40.577
R22392 minus.n29 minus.n28 40.577
R22393 minus.n61 minus.n60 39.4345
R22394 minus.n12 minus.n11 39.4345
R22395 minus.n88 minus.n52 36.702
R22396 minus.n66 minus.n58 36.702
R22397 minus.n17 minus.n9 36.702
R22398 minus.n39 minus.n3 36.702
R22399 minus.n98 minus.n97 33.563
R22400 minus.n90 minus.n89 20.9036
R22401 minus.n65 minus.n64 20.9036
R22402 minus.n16 minus.n15 20.9036
R22403 minus.n41 minus.n40 20.9036
R22404 minus.n100 minus.t3 19.8005
R22405 minus.n100 minus.t0 19.8005
R22406 minus.n99 minus.t2 19.8005
R22407 minus.n99 minus.t1 19.8005
R22408 minus.n81 minus.n54 18.9362
R22409 minus.n73 minus.n56 18.9362
R22410 minus.n24 minus.n7 18.9362
R22411 minus.n32 minus.n5 18.9362
R22412 minus.n83 minus.n82 16.9689
R22413 minus.n72 minus.n71 16.9689
R22414 minus.n23 minus.n22 16.9689
R22415 minus.n34 minus.n33 16.9689
R22416 minus.n91 minus.n50 15.0015
R22417 minus.n63 minus.n60 15.0015
R22418 minus.n14 minus.n11 15.0015
R22419 minus.n42 minus.n1 15.0015
R22420 minus.n96 minus.n95 12.4157
R22421 minus.n47 minus.n46 12.4157
R22422 minus.n98 minus.n48 12.1577
R22423 minus minus.n103 11.0699
R22424 minus.n94 minus.n50 9.59132
R22425 minus.n45 minus.n1 9.59132
R22426 minus.n84 minus.n83 7.62397
R22427 minus.n71 minus.n70 7.62397
R22428 minus.n22 minus.n21 7.62397
R22429 minus.n35 minus.n34 7.62397
R22430 minus.n78 minus.n54 5.65662
R22431 minus.n76 minus.n56 5.65662
R22432 minus.n27 minus.n7 5.65662
R22433 minus.n29 minus.n5 5.65662
R22434 minus.n103 minus.n102 4.80222
R22435 minus.n89 minus.n88 3.68928
R22436 minus.n66 minus.n65 3.68928
R22437 minus.n17 minus.n16 3.68928
R22438 minus.n40 minus.n39 3.68928
R22439 minus.n103 minus.n98 0.972091
R22440 minus.n102 minus.n101 0.716017
R22441 minus.n97 minus.n49 0.189894
R22442 minus.n93 minus.n49 0.189894
R22443 minus.n93 minus.n92 0.189894
R22444 minus.n92 minus.n51 0.189894
R22445 minus.n87 minus.n51 0.189894
R22446 minus.n87 minus.n86 0.189894
R22447 minus.n86 minus.n85 0.189894
R22448 minus.n85 minus.n53 0.189894
R22449 minus.n80 minus.n53 0.189894
R22450 minus.n80 minus.n79 0.189894
R22451 minus.n79 minus.n55 0.189894
R22452 minus.n75 minus.n55 0.189894
R22453 minus.n75 minus.n74 0.189894
R22454 minus.n74 minus.n57 0.189894
R22455 minus.n69 minus.n57 0.189894
R22456 minus.n69 minus.n68 0.189894
R22457 minus.n68 minus.n67 0.189894
R22458 minus.n67 minus.n59 0.189894
R22459 minus.n62 minus.n59 0.189894
R22460 minus.n13 minus.n10 0.189894
R22461 minus.n18 minus.n10 0.189894
R22462 minus.n19 minus.n18 0.189894
R22463 minus.n20 minus.n19 0.189894
R22464 minus.n20 minus.n8 0.189894
R22465 minus.n25 minus.n8 0.189894
R22466 minus.n26 minus.n25 0.189894
R22467 minus.n26 minus.n6 0.189894
R22468 minus.n30 minus.n6 0.189894
R22469 minus.n31 minus.n30 0.189894
R22470 minus.n31 minus.n4 0.189894
R22471 minus.n36 minus.n4 0.189894
R22472 minus.n37 minus.n36 0.189894
R22473 minus.n38 minus.n37 0.189894
R22474 minus.n38 minus.n2 0.189894
R22475 minus.n43 minus.n2 0.189894
R22476 minus.n44 minus.n43 0.189894
R22477 minus.n44 minus.n0 0.189894
R22478 minus.n48 minus.n0 0.189894
R22479 diffpairibias.n0 diffpairibias.t18 436.822
R22480 diffpairibias.n21 diffpairibias.t19 435.479
R22481 diffpairibias.n20 diffpairibias.t16 435.479
R22482 diffpairibias.n19 diffpairibias.t17 435.479
R22483 diffpairibias.n18 diffpairibias.t21 435.479
R22484 diffpairibias.n0 diffpairibias.t22 435.479
R22485 diffpairibias.n1 diffpairibias.t20 435.479
R22486 diffpairibias.n2 diffpairibias.t23 435.479
R22487 diffpairibias.n10 diffpairibias.t0 377.536
R22488 diffpairibias.n10 diffpairibias.t8 376.193
R22489 diffpairibias.n11 diffpairibias.t10 376.193
R22490 diffpairibias.n12 diffpairibias.t6 376.193
R22491 diffpairibias.n13 diffpairibias.t2 376.193
R22492 diffpairibias.n14 diffpairibias.t12 376.193
R22493 diffpairibias.n15 diffpairibias.t4 376.193
R22494 diffpairibias.n16 diffpairibias.t14 376.193
R22495 diffpairibias.n3 diffpairibias.t1 113.368
R22496 diffpairibias.n3 diffpairibias.t9 112.698
R22497 diffpairibias.n4 diffpairibias.t11 112.698
R22498 diffpairibias.n5 diffpairibias.t7 112.698
R22499 diffpairibias.n6 diffpairibias.t3 112.698
R22500 diffpairibias.n7 diffpairibias.t13 112.698
R22501 diffpairibias.n8 diffpairibias.t5 112.698
R22502 diffpairibias.n9 diffpairibias.t15 112.698
R22503 diffpairibias.n17 diffpairibias.n16 4.77242
R22504 diffpairibias.n17 diffpairibias.n9 4.30807
R22505 diffpairibias.n18 diffpairibias.n17 4.13945
R22506 diffpairibias.n16 diffpairibias.n15 1.34352
R22507 diffpairibias.n15 diffpairibias.n14 1.34352
R22508 diffpairibias.n14 diffpairibias.n13 1.34352
R22509 diffpairibias.n13 diffpairibias.n12 1.34352
R22510 diffpairibias.n12 diffpairibias.n11 1.34352
R22511 diffpairibias.n11 diffpairibias.n10 1.34352
R22512 diffpairibias.n2 diffpairibias.n1 1.34352
R22513 diffpairibias.n1 diffpairibias.n0 1.34352
R22514 diffpairibias.n19 diffpairibias.n18 1.34352
R22515 diffpairibias.n20 diffpairibias.n19 1.34352
R22516 diffpairibias.n21 diffpairibias.n20 1.34352
R22517 diffpairibias.n22 diffpairibias.n21 0.862419
R22518 diffpairibias diffpairibias.n22 0.684875
R22519 diffpairibias.n9 diffpairibias.n8 0.672012
R22520 diffpairibias.n8 diffpairibias.n7 0.672012
R22521 diffpairibias.n7 diffpairibias.n6 0.672012
R22522 diffpairibias.n6 diffpairibias.n5 0.672012
R22523 diffpairibias.n5 diffpairibias.n4 0.672012
R22524 diffpairibias.n4 diffpairibias.n3 0.672012
R22525 diffpairibias.n22 diffpairibias.n2 0.190907
C0 plus commonsourceibias 0.417817f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13571f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 0.117738p
C6 minus diffpairibias 5.12e-19
C7 commonsourceibias output 0.006808f
C8 vdd plus 0.091948f
C9 CSoutput minus 2.37773f
C10 plus diffpairibias 4.13e-19
C11 commonsourceibias outputibias 0.003832f
C12 CSoutput plus 0.85599f
C13 vdd commonsourceibias 0.004218f
C14 commonsourceibias diffpairibias 0.052851f
C15 minus plus 9.23291f
C16 CSoutput commonsourceibias 29.0223f
C17 minus commonsourceibias 0.462976f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118431p
C22 plus gnd 34.639297f
C23 minus gnd 27.083952f
C24 CSoutput gnd 87.43974f
C25 vdd gnd 0.47715p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031196f
C74 minus.t13 gnd 0.52455f
C75 minus.n1 gnd 0.212151f
C76 minus.n2 gnd 0.031196f
C77 minus.t20 gnd 0.52455f
C78 minus.n3 gnd 0.025838f
C79 minus.n4 gnd 0.031196f
C80 minus.t17 gnd 0.52455f
C81 minus.t23 gnd 0.52455f
C82 minus.n5 gnd 0.212151f
C83 minus.n6 gnd 0.031196f
C84 minus.t22 gnd 0.52455f
C85 minus.n7 gnd 0.212151f
C86 minus.n8 gnd 0.031196f
C87 minus.t5 gnd 0.52455f
C88 minus.n9 gnd 0.025838f
C89 minus.n10 gnd 0.031196f
C90 minus.t8 gnd 0.52455f
C91 minus.t10 gnd 0.52455f
C92 minus.n11 gnd 0.243966f
C93 minus.t16 gnd 0.587882f
C94 minus.n12 gnd 0.247088f
C95 minus.n13 gnd 0.133151f
C96 minus.n14 gnd 0.039389f
C97 minus.n15 gnd 0.035885f
C98 minus.n16 gnd 0.212151f
C99 minus.n17 gnd 0.038286f
C100 minus.n18 gnd 0.031196f
C101 minus.n19 gnd 0.031196f
C102 minus.n20 gnd 0.031196f
C103 minus.n21 gnd 0.040441f
C104 minus.n22 gnd 0.212151f
C105 minus.n23 gnd 0.038221f
C106 minus.n24 gnd 0.037053f
C107 minus.n25 gnd 0.031196f
C108 minus.n26 gnd 0.031196f
C109 minus.n27 gnd 0.039684f
C110 minus.n28 gnd 0.025196f
C111 minus.n29 gnd 0.039684f
C112 minus.n30 gnd 0.031196f
C113 minus.n31 gnd 0.031196f
C114 minus.n32 gnd 0.037053f
C115 minus.n33 gnd 0.038221f
C116 minus.n34 gnd 0.212151f
C117 minus.n35 gnd 0.040441f
C118 minus.n36 gnd 0.031196f
C119 minus.n37 gnd 0.031196f
C120 minus.n38 gnd 0.031196f
C121 minus.n39 gnd 0.038286f
C122 minus.n40 gnd 0.212151f
C123 minus.n41 gnd 0.035885f
C124 minus.n42 gnd 0.039389f
C125 minus.n43 gnd 0.031196f
C126 minus.n44 gnd 0.031196f
C127 minus.n45 gnd 0.040709f
C128 minus.n46 gnd 0.012082f
C129 minus.t9 gnd 0.567301f
C130 minus.n47 gnd 0.24602f
C131 minus.n48 gnd 0.366f
C132 minus.n49 gnd 0.031196f
C133 minus.t14 gnd 0.567301f
C134 minus.t21 gnd 0.52455f
C135 minus.n50 gnd 0.212151f
C136 minus.n51 gnd 0.031196f
C137 minus.t18 gnd 0.52455f
C138 minus.n52 gnd 0.025838f
C139 minus.n53 gnd 0.031196f
C140 minus.t15 gnd 0.52455f
C141 minus.t7 gnd 0.52455f
C142 minus.n54 gnd 0.212151f
C143 minus.n55 gnd 0.031196f
C144 minus.t6 gnd 0.52455f
C145 minus.n56 gnd 0.212151f
C146 minus.n57 gnd 0.031196f
C147 minus.t12 gnd 0.52455f
C148 minus.n58 gnd 0.025838f
C149 minus.n59 gnd 0.031196f
C150 minus.t11 gnd 0.52455f
C151 minus.t19 gnd 0.52455f
C152 minus.n60 gnd 0.243966f
C153 minus.t24 gnd 0.587882f
C154 minus.n61 gnd 0.247088f
C155 minus.n62 gnd 0.133151f
C156 minus.n63 gnd 0.039389f
C157 minus.n64 gnd 0.035885f
C158 minus.n65 gnd 0.212151f
C159 minus.n66 gnd 0.038286f
C160 minus.n67 gnd 0.031196f
C161 minus.n68 gnd 0.031196f
C162 minus.n69 gnd 0.031196f
C163 minus.n70 gnd 0.040441f
C164 minus.n71 gnd 0.212151f
C165 minus.n72 gnd 0.038221f
C166 minus.n73 gnd 0.037053f
C167 minus.n74 gnd 0.031196f
C168 minus.n75 gnd 0.031196f
C169 minus.n76 gnd 0.039684f
C170 minus.n77 gnd 0.025196f
C171 minus.n78 gnd 0.039684f
C172 minus.n79 gnd 0.031196f
C173 minus.n80 gnd 0.031196f
C174 minus.n81 gnd 0.037053f
C175 minus.n82 gnd 0.038221f
C176 minus.n83 gnd 0.212151f
C177 minus.n84 gnd 0.040441f
C178 minus.n85 gnd 0.031196f
C179 minus.n86 gnd 0.031196f
C180 minus.n87 gnd 0.031196f
C181 minus.n88 gnd 0.038286f
C182 minus.n89 gnd 0.212151f
C183 minus.n90 gnd 0.035885f
C184 minus.n91 gnd 0.039389f
C185 minus.n92 gnd 0.031196f
C186 minus.n93 gnd 0.031196f
C187 minus.n94 gnd 0.040709f
C188 minus.n95 gnd 0.012082f
C189 minus.n96 gnd 0.24602f
C190 minus.n97 gnd 1.0544f
C191 minus.n98 gnd 1.56697f
C192 minus.t2 gnd 0.009617f
C193 minus.t1 gnd 0.009617f
C194 minus.n99 gnd 0.031622f
C195 minus.t3 gnd 0.009617f
C196 minus.t0 gnd 0.009617f
C197 minus.n100 gnd 0.031189f
C198 minus.n101 gnd 0.266181f
C199 minus.t4 gnd 0.053525f
C200 minus.n102 gnd 0.145253f
C201 minus.n103 gnd 1.66979f
C202 a_n2650_8322.t12 gnd 0.098096f
C203 a_n2650_8322.t5 gnd 20.351f
C204 a_n2650_8322.t0 gnd 20.2083f
C205 a_n2650_8322.t3 gnd 20.2083f
C206 a_n2650_8322.t4 gnd 20.351f
C207 a_n2650_8322.t1 gnd 20.2083f
C208 a_n2650_8322.t2 gnd 27.901402f
C209 a_n2650_8322.t21 gnd 0.918523f
C210 a_n2650_8322.t24 gnd 0.098096f
C211 a_n2650_8322.t16 gnd 0.098096f
C212 a_n2650_8322.n0 gnd 0.69099f
C213 a_n2650_8322.n1 gnd 0.772079f
C214 a_n2650_8322.t8 gnd 0.098096f
C215 a_n2650_8322.t7 gnd 0.098096f
C216 a_n2650_8322.n2 gnd 0.69099f
C217 a_n2650_8322.n3 gnd 0.392283f
C218 a_n2650_8322.t19 gnd 0.098096f
C219 a_n2650_8322.t13 gnd 0.098096f
C220 a_n2650_8322.n4 gnd 0.69099f
C221 a_n2650_8322.n5 gnd 0.392283f
C222 a_n2650_8322.t17 gnd 0.098096f
C223 a_n2650_8322.t15 gnd 0.098096f
C224 a_n2650_8322.n6 gnd 0.69099f
C225 a_n2650_8322.n7 gnd 0.392283f
C226 a_n2650_8322.t6 gnd 0.916694f
C227 a_n2650_8322.n8 gnd 1.71065f
C228 a_n2650_8322.t29 gnd 0.918523f
C229 a_n2650_8322.t32 gnd 0.098096f
C230 a_n2650_8322.t33 gnd 0.098096f
C231 a_n2650_8322.n9 gnd 0.69099f
C232 a_n2650_8322.n10 gnd 0.772079f
C233 a_n2650_8322.t27 gnd 0.916694f
C234 a_n2650_8322.n11 gnd 0.388521f
C235 a_n2650_8322.t30 gnd 0.916694f
C236 a_n2650_8322.n12 gnd 0.388521f
C237 a_n2650_8322.t28 gnd 0.098096f
C238 a_n2650_8322.t26 gnd 0.098096f
C239 a_n2650_8322.n13 gnd 0.69099f
C240 a_n2650_8322.n14 gnd 0.392283f
C241 a_n2650_8322.t31 gnd 0.916694f
C242 a_n2650_8322.n15 gnd 1.27468f
C243 a_n2650_8322.n16 gnd 2.0827f
C244 a_n2650_8322.n17 gnd 3.05665f
C245 a_n2650_8322.t20 gnd 0.916694f
C246 a_n2650_8322.n18 gnd 0.997099f
C247 a_n2650_8322.t9 gnd 0.098096f
C248 a_n2650_8322.t10 gnd 0.098096f
C249 a_n2650_8322.n19 gnd 0.69099f
C250 a_n2650_8322.n20 gnd 0.392283f
C251 a_n2650_8322.t22 gnd 0.098096f
C252 a_n2650_8322.t11 gnd 0.098096f
C253 a_n2650_8322.n21 gnd 0.69099f
C254 a_n2650_8322.n22 gnd 0.392283f
C255 a_n2650_8322.t23 gnd 0.918521f
C256 a_n2650_8322.t18 gnd 0.098096f
C257 a_n2650_8322.t14 gnd 0.098096f
C258 a_n2650_8322.n23 gnd 0.69099f
C259 a_n2650_8322.n24 gnd 0.772081f
C260 a_n2650_8322.n25 gnd 0.392282f
C261 a_n2650_8322.n26 gnd 0.690992f
C262 a_n2650_8322.t25 gnd 0.098096f
C263 output.t12 gnd 0.464308f
C264 output.t3 gnd 0.044422f
C265 output.t7 gnd 0.044422f
C266 output.n0 gnd 0.364624f
C267 output.n1 gnd 0.614102f
C268 output.t10 gnd 0.044422f
C269 output.t15 gnd 0.044422f
C270 output.n2 gnd 0.364624f
C271 output.n3 gnd 0.350265f
C272 output.t0 gnd 0.044422f
C273 output.t5 gnd 0.044422f
C274 output.n4 gnd 0.364624f
C275 output.n5 gnd 0.350265f
C276 output.t9 gnd 0.044422f
C277 output.t1 gnd 0.044422f
C278 output.n6 gnd 0.364624f
C279 output.n7 gnd 0.350265f
C280 output.t4 gnd 0.044422f
C281 output.t2 gnd 0.044422f
C282 output.n8 gnd 0.364624f
C283 output.n9 gnd 0.350265f
C284 output.t8 gnd 0.044422f
C285 output.t11 gnd 0.044422f
C286 output.n10 gnd 0.364624f
C287 output.n11 gnd 0.350265f
C288 output.t13 gnd 0.044422f
C289 output.t6 gnd 0.044422f
C290 output.n12 gnd 0.364624f
C291 output.n13 gnd 0.350265f
C292 output.t14 gnd 0.462979f
C293 output.n14 gnd 0.28994f
C294 output.n15 gnd 0.015803f
C295 output.n16 gnd 0.011243f
C296 output.n17 gnd 0.006041f
C297 output.n18 gnd 0.01428f
C298 output.n19 gnd 0.006397f
C299 output.n20 gnd 0.011243f
C300 output.n21 gnd 0.006041f
C301 output.n22 gnd 0.01428f
C302 output.n23 gnd 0.006397f
C303 output.n24 gnd 0.048111f
C304 output.t19 gnd 0.023274f
C305 output.n25 gnd 0.01071f
C306 output.n26 gnd 0.008435f
C307 output.n27 gnd 0.006041f
C308 output.n28 gnd 0.267512f
C309 output.n29 gnd 0.011243f
C310 output.n30 gnd 0.006041f
C311 output.n31 gnd 0.006397f
C312 output.n32 gnd 0.01428f
C313 output.n33 gnd 0.01428f
C314 output.n34 gnd 0.006397f
C315 output.n35 gnd 0.006041f
C316 output.n36 gnd 0.011243f
C317 output.n37 gnd 0.011243f
C318 output.n38 gnd 0.006041f
C319 output.n39 gnd 0.006397f
C320 output.n40 gnd 0.01428f
C321 output.n41 gnd 0.030913f
C322 output.n42 gnd 0.006397f
C323 output.n43 gnd 0.006041f
C324 output.n44 gnd 0.025987f
C325 output.n45 gnd 0.097665f
C326 output.n46 gnd 0.015803f
C327 output.n47 gnd 0.011243f
C328 output.n48 gnd 0.006041f
C329 output.n49 gnd 0.01428f
C330 output.n50 gnd 0.006397f
C331 output.n51 gnd 0.011243f
C332 output.n52 gnd 0.006041f
C333 output.n53 gnd 0.01428f
C334 output.n54 gnd 0.006397f
C335 output.n55 gnd 0.048111f
C336 output.t18 gnd 0.023274f
C337 output.n56 gnd 0.01071f
C338 output.n57 gnd 0.008435f
C339 output.n58 gnd 0.006041f
C340 output.n59 gnd 0.267512f
C341 output.n60 gnd 0.011243f
C342 output.n61 gnd 0.006041f
C343 output.n62 gnd 0.006397f
C344 output.n63 gnd 0.01428f
C345 output.n64 gnd 0.01428f
C346 output.n65 gnd 0.006397f
C347 output.n66 gnd 0.006041f
C348 output.n67 gnd 0.011243f
C349 output.n68 gnd 0.011243f
C350 output.n69 gnd 0.006041f
C351 output.n70 gnd 0.006397f
C352 output.n71 gnd 0.01428f
C353 output.n72 gnd 0.030913f
C354 output.n73 gnd 0.006397f
C355 output.n74 gnd 0.006041f
C356 output.n75 gnd 0.025987f
C357 output.n76 gnd 0.09306f
C358 output.n77 gnd 1.65264f
C359 output.n78 gnd 0.015803f
C360 output.n79 gnd 0.011243f
C361 output.n80 gnd 0.006041f
C362 output.n81 gnd 0.01428f
C363 output.n82 gnd 0.006397f
C364 output.n83 gnd 0.011243f
C365 output.n84 gnd 0.006041f
C366 output.n85 gnd 0.01428f
C367 output.n86 gnd 0.006397f
C368 output.n87 gnd 0.048111f
C369 output.t17 gnd 0.023274f
C370 output.n88 gnd 0.01071f
C371 output.n89 gnd 0.008435f
C372 output.n90 gnd 0.006041f
C373 output.n91 gnd 0.267512f
C374 output.n92 gnd 0.011243f
C375 output.n93 gnd 0.006041f
C376 output.n94 gnd 0.006397f
C377 output.n95 gnd 0.01428f
C378 output.n96 gnd 0.01428f
C379 output.n97 gnd 0.006397f
C380 output.n98 gnd 0.006041f
C381 output.n99 gnd 0.011243f
C382 output.n100 gnd 0.011243f
C383 output.n101 gnd 0.006041f
C384 output.n102 gnd 0.006397f
C385 output.n103 gnd 0.01428f
C386 output.n104 gnd 0.030913f
C387 output.n105 gnd 0.006397f
C388 output.n106 gnd 0.006041f
C389 output.n107 gnd 0.025987f
C390 output.n108 gnd 0.09306f
C391 output.n109 gnd 0.713089f
C392 output.n110 gnd 0.015803f
C393 output.n111 gnd 0.011243f
C394 output.n112 gnd 0.006041f
C395 output.n113 gnd 0.01428f
C396 output.n114 gnd 0.006397f
C397 output.n115 gnd 0.011243f
C398 output.n116 gnd 0.006041f
C399 output.n117 gnd 0.01428f
C400 output.n118 gnd 0.006397f
C401 output.n119 gnd 0.048111f
C402 output.t16 gnd 0.023274f
C403 output.n120 gnd 0.01071f
C404 output.n121 gnd 0.008435f
C405 output.n122 gnd 0.006041f
C406 output.n123 gnd 0.267512f
C407 output.n124 gnd 0.011243f
C408 output.n125 gnd 0.006041f
C409 output.n126 gnd 0.006397f
C410 output.n127 gnd 0.01428f
C411 output.n128 gnd 0.01428f
C412 output.n129 gnd 0.006397f
C413 output.n130 gnd 0.006041f
C414 output.n131 gnd 0.011243f
C415 output.n132 gnd 0.011243f
C416 output.n133 gnd 0.006041f
C417 output.n134 gnd 0.006397f
C418 output.n135 gnd 0.01428f
C419 output.n136 gnd 0.030913f
C420 output.n137 gnd 0.006397f
C421 output.n138 gnd 0.006041f
C422 output.n139 gnd 0.025987f
C423 output.n140 gnd 0.09306f
C424 output.n141 gnd 1.67353f
C425 outputibias.t9 gnd 0.11477f
C426 outputibias.t8 gnd 0.115567f
C427 outputibias.n0 gnd 0.130108f
C428 outputibias.n1 gnd 0.001372f
C429 outputibias.n2 gnd 9.76e-19
C430 outputibias.n3 gnd 5.24e-19
C431 outputibias.n4 gnd 0.001239f
C432 outputibias.n5 gnd 5.55e-19
C433 outputibias.n6 gnd 9.76e-19
C434 outputibias.n7 gnd 5.24e-19
C435 outputibias.n8 gnd 0.001239f
C436 outputibias.n9 gnd 5.55e-19
C437 outputibias.n10 gnd 0.004176f
C438 outputibias.t5 gnd 0.00202f
C439 outputibias.n11 gnd 9.3e-19
C440 outputibias.n12 gnd 7.32e-19
C441 outputibias.n13 gnd 5.24e-19
C442 outputibias.n14 gnd 0.02322f
C443 outputibias.n15 gnd 9.76e-19
C444 outputibias.n16 gnd 5.24e-19
C445 outputibias.n17 gnd 5.55e-19
C446 outputibias.n18 gnd 0.001239f
C447 outputibias.n19 gnd 0.001239f
C448 outputibias.n20 gnd 5.55e-19
C449 outputibias.n21 gnd 5.24e-19
C450 outputibias.n22 gnd 9.76e-19
C451 outputibias.n23 gnd 9.76e-19
C452 outputibias.n24 gnd 5.24e-19
C453 outputibias.n25 gnd 5.55e-19
C454 outputibias.n26 gnd 0.001239f
C455 outputibias.n27 gnd 0.002683f
C456 outputibias.n28 gnd 5.55e-19
C457 outputibias.n29 gnd 5.24e-19
C458 outputibias.n30 gnd 0.002256f
C459 outputibias.n31 gnd 0.005781f
C460 outputibias.n32 gnd 0.001372f
C461 outputibias.n33 gnd 9.76e-19
C462 outputibias.n34 gnd 5.24e-19
C463 outputibias.n35 gnd 0.001239f
C464 outputibias.n36 gnd 5.55e-19
C465 outputibias.n37 gnd 9.76e-19
C466 outputibias.n38 gnd 5.24e-19
C467 outputibias.n39 gnd 0.001239f
C468 outputibias.n40 gnd 5.55e-19
C469 outputibias.n41 gnd 0.004176f
C470 outputibias.t7 gnd 0.00202f
C471 outputibias.n42 gnd 9.3e-19
C472 outputibias.n43 gnd 7.32e-19
C473 outputibias.n44 gnd 5.24e-19
C474 outputibias.n45 gnd 0.02322f
C475 outputibias.n46 gnd 9.76e-19
C476 outputibias.n47 gnd 5.24e-19
C477 outputibias.n48 gnd 5.55e-19
C478 outputibias.n49 gnd 0.001239f
C479 outputibias.n50 gnd 0.001239f
C480 outputibias.n51 gnd 5.55e-19
C481 outputibias.n52 gnd 5.24e-19
C482 outputibias.n53 gnd 9.76e-19
C483 outputibias.n54 gnd 9.76e-19
C484 outputibias.n55 gnd 5.24e-19
C485 outputibias.n56 gnd 5.55e-19
C486 outputibias.n57 gnd 0.001239f
C487 outputibias.n58 gnd 0.002683f
C488 outputibias.n59 gnd 5.55e-19
C489 outputibias.n60 gnd 5.24e-19
C490 outputibias.n61 gnd 0.002256f
C491 outputibias.n62 gnd 0.005197f
C492 outputibias.n63 gnd 0.121892f
C493 outputibias.n64 gnd 0.001372f
C494 outputibias.n65 gnd 9.76e-19
C495 outputibias.n66 gnd 5.24e-19
C496 outputibias.n67 gnd 0.001239f
C497 outputibias.n68 gnd 5.55e-19
C498 outputibias.n69 gnd 9.76e-19
C499 outputibias.n70 gnd 5.24e-19
C500 outputibias.n71 gnd 0.001239f
C501 outputibias.n72 gnd 5.55e-19
C502 outputibias.n73 gnd 0.004176f
C503 outputibias.t1 gnd 0.00202f
C504 outputibias.n74 gnd 9.3e-19
C505 outputibias.n75 gnd 7.32e-19
C506 outputibias.n76 gnd 5.24e-19
C507 outputibias.n77 gnd 0.02322f
C508 outputibias.n78 gnd 9.76e-19
C509 outputibias.n79 gnd 5.24e-19
C510 outputibias.n80 gnd 5.55e-19
C511 outputibias.n81 gnd 0.001239f
C512 outputibias.n82 gnd 0.001239f
C513 outputibias.n83 gnd 5.55e-19
C514 outputibias.n84 gnd 5.24e-19
C515 outputibias.n85 gnd 9.76e-19
C516 outputibias.n86 gnd 9.76e-19
C517 outputibias.n87 gnd 5.24e-19
C518 outputibias.n88 gnd 5.55e-19
C519 outputibias.n89 gnd 0.001239f
C520 outputibias.n90 gnd 0.002683f
C521 outputibias.n91 gnd 5.55e-19
C522 outputibias.n92 gnd 5.24e-19
C523 outputibias.n93 gnd 0.002256f
C524 outputibias.n94 gnd 0.005197f
C525 outputibias.n95 gnd 0.064513f
C526 outputibias.n96 gnd 0.001372f
C527 outputibias.n97 gnd 9.76e-19
C528 outputibias.n98 gnd 5.24e-19
C529 outputibias.n99 gnd 0.001239f
C530 outputibias.n100 gnd 5.55e-19
C531 outputibias.n101 gnd 9.76e-19
C532 outputibias.n102 gnd 5.24e-19
C533 outputibias.n103 gnd 0.001239f
C534 outputibias.n104 gnd 5.55e-19
C535 outputibias.n105 gnd 0.004176f
C536 outputibias.t3 gnd 0.00202f
C537 outputibias.n106 gnd 9.3e-19
C538 outputibias.n107 gnd 7.32e-19
C539 outputibias.n108 gnd 5.24e-19
C540 outputibias.n109 gnd 0.02322f
C541 outputibias.n110 gnd 9.76e-19
C542 outputibias.n111 gnd 5.24e-19
C543 outputibias.n112 gnd 5.55e-19
C544 outputibias.n113 gnd 0.001239f
C545 outputibias.n114 gnd 0.001239f
C546 outputibias.n115 gnd 5.55e-19
C547 outputibias.n116 gnd 5.24e-19
C548 outputibias.n117 gnd 9.76e-19
C549 outputibias.n118 gnd 9.76e-19
C550 outputibias.n119 gnd 5.24e-19
C551 outputibias.n120 gnd 5.55e-19
C552 outputibias.n121 gnd 0.001239f
C553 outputibias.n122 gnd 0.002683f
C554 outputibias.n123 gnd 5.55e-19
C555 outputibias.n124 gnd 5.24e-19
C556 outputibias.n125 gnd 0.002256f
C557 outputibias.n126 gnd 0.005197f
C558 outputibias.n127 gnd 0.084814f
C559 outputibias.t2 gnd 0.108319f
C560 outputibias.t0 gnd 0.108319f
C561 outputibias.t6 gnd 0.108319f
C562 outputibias.t4 gnd 0.109238f
C563 outputibias.n128 gnd 0.134674f
C564 outputibias.n129 gnd 0.07244f
C565 outputibias.n130 gnd 0.079818f
C566 outputibias.n131 gnd 0.164901f
C567 outputibias.t11 gnd 0.11477f
C568 outputibias.n132 gnd 0.067481f
C569 outputibias.t10 gnd 0.11477f
C570 outputibias.n133 gnd 0.065115f
C571 outputibias.n134 gnd 0.029159f
C572 a_n2903_n3924.t17 gnd 0.094851f
C573 a_n2903_n3924.t27 gnd 0.985803f
C574 a_n2903_n3924.n0 gnd 0.372677f
C575 a_n2903_n3924.t5 gnd 1.22484f
C576 a_n2903_n3924.n1 gnd 1.15477f
C577 a_n2903_n3924.t44 gnd 0.985803f
C578 a_n2903_n3924.n2 gnd 0.372677f
C579 a_n2903_n3924.t13 gnd 0.094851f
C580 a_n2903_n3924.t38 gnd 0.094851f
C581 a_n2903_n3924.n3 gnd 0.774663f
C582 a_n2903_n3924.n4 gnd 0.390386f
C583 a_n2903_n3924.t8 gnd 0.094851f
C584 a_n2903_n3924.t9 gnd 0.094851f
C585 a_n2903_n3924.n5 gnd 0.774663f
C586 a_n2903_n3924.n6 gnd 0.390386f
C587 a_n2903_n3924.t42 gnd 0.094851f
C588 a_n2903_n3924.t46 gnd 0.094851f
C589 a_n2903_n3924.n7 gnd 0.774663f
C590 a_n2903_n3924.n8 gnd 0.390386f
C591 a_n2903_n3924.t36 gnd 0.094851f
C592 a_n2903_n3924.t39 gnd 0.094851f
C593 a_n2903_n3924.n9 gnd 0.774663f
C594 a_n2903_n3924.n10 gnd 0.390386f
C595 a_n2903_n3924.t35 gnd 0.985803f
C596 a_n2903_n3924.n11 gnd 0.922787f
C597 a_n2903_n3924.t2 gnd 1.22537f
C598 a_n2903_n3924.t1 gnd 1.22484f
C599 a_n2903_n3924.n12 gnd 0.862674f
C600 a_n2903_n3924.t0 gnd 1.22484f
C601 a_n2903_n3924.n13 gnd 0.862674f
C602 a_n2903_n3924.t34 gnd 1.22484f
C603 a_n2903_n3924.n14 gnd 0.862674f
C604 a_n2903_n3924.t47 gnd 1.22484f
C605 a_n2903_n3924.n15 gnd 0.862674f
C606 a_n2903_n3924.t3 gnd 1.22484f
C607 a_n2903_n3924.n16 gnd 0.862674f
C608 a_n2903_n3924.t4 gnd 1.22484f
C609 a_n2903_n3924.n17 gnd 0.716127f
C610 a_n2903_n3924.n18 gnd 0.845678f
C611 a_n2903_n3924.n19 gnd 0.894202f
C612 a_n2903_n3924.t32 gnd 0.985799f
C613 a_n2903_n3924.n20 gnd 0.612329f
C614 a_n2903_n3924.t26 gnd 0.094851f
C615 a_n2903_n3924.t30 gnd 0.094851f
C616 a_n2903_n3924.n21 gnd 0.774662f
C617 a_n2903_n3924.n22 gnd 0.390388f
C618 a_n2903_n3924.t31 gnd 0.094851f
C619 a_n2903_n3924.t19 gnd 0.094851f
C620 a_n2903_n3924.n23 gnd 0.774662f
C621 a_n2903_n3924.n24 gnd 0.390388f
C622 a_n2903_n3924.t20 gnd 0.094851f
C623 a_n2903_n3924.t14 gnd 0.094851f
C624 a_n2903_n3924.n25 gnd 0.774662f
C625 a_n2903_n3924.n26 gnd 0.390388f
C626 a_n2903_n3924.t16 gnd 0.094851f
C627 a_n2903_n3924.t29 gnd 0.094851f
C628 a_n2903_n3924.n27 gnd 0.774662f
C629 a_n2903_n3924.n28 gnd 0.390388f
C630 a_n2903_n3924.t24 gnd 0.985799f
C631 a_n2903_n3924.n29 gnd 0.372681f
C632 a_n2903_n3924.t41 gnd 0.985799f
C633 a_n2903_n3924.n30 gnd 0.372681f
C634 a_n2903_n3924.t10 gnd 0.094851f
C635 a_n2903_n3924.t6 gnd 0.094851f
C636 a_n2903_n3924.n31 gnd 0.774662f
C637 a_n2903_n3924.n32 gnd 0.390388f
C638 a_n2903_n3924.t7 gnd 0.094851f
C639 a_n2903_n3924.t43 gnd 0.094851f
C640 a_n2903_n3924.n33 gnd 0.774662f
C641 a_n2903_n3924.n34 gnd 0.390388f
C642 a_n2903_n3924.t45 gnd 0.094851f
C643 a_n2903_n3924.t40 gnd 0.094851f
C644 a_n2903_n3924.n35 gnd 0.774662f
C645 a_n2903_n3924.n36 gnd 0.390388f
C646 a_n2903_n3924.t37 gnd 0.094851f
C647 a_n2903_n3924.t12 gnd 0.094851f
C648 a_n2903_n3924.n37 gnd 0.774662f
C649 a_n2903_n3924.n38 gnd 0.390388f
C650 a_n2903_n3924.t11 gnd 0.985799f
C651 a_n2903_n3924.n39 gnd 0.612329f
C652 a_n2903_n3924.n40 gnd 0.953249f
C653 a_n2903_n3924.t15 gnd 0.985799f
C654 a_n2903_n3924.n41 gnd 0.922791f
C655 a_n2903_n3924.t23 gnd 0.094851f
C656 a_n2903_n3924.t28 gnd 0.094851f
C657 a_n2903_n3924.n42 gnd 0.774663f
C658 a_n2903_n3924.n43 gnd 0.390386f
C659 a_n2903_n3924.t21 gnd 0.094851f
C660 a_n2903_n3924.t25 gnd 0.094851f
C661 a_n2903_n3924.n44 gnd 0.774663f
C662 a_n2903_n3924.n45 gnd 0.390386f
C663 a_n2903_n3924.t18 gnd 0.094851f
C664 a_n2903_n3924.t22 gnd 0.094851f
C665 a_n2903_n3924.n46 gnd 0.774663f
C666 a_n2903_n3924.n47 gnd 0.390386f
C667 a_n2903_n3924.n48 gnd 0.390385f
C668 a_n2903_n3924.n49 gnd 0.774665f
C669 a_n2903_n3924.t33 gnd 0.094851f
C670 plus.n0 gnd 0.023096f
C671 plus.t6 gnd 0.42001f
C672 plus.t12 gnd 0.388359f
C673 plus.n1 gnd 0.15707f
C674 plus.n2 gnd 0.023096f
C675 plus.t8 gnd 0.388359f
C676 plus.n3 gnd 0.019129f
C677 plus.n4 gnd 0.023096f
C678 plus.t7 gnd 0.388359f
C679 plus.t19 gnd 0.388359f
C680 plus.n5 gnd 0.15707f
C681 plus.n6 gnd 0.023096f
C682 plus.t18 gnd 0.388359f
C683 plus.n7 gnd 0.15707f
C684 plus.n8 gnd 0.023096f
C685 plus.t24 gnd 0.388359f
C686 plus.n9 gnd 0.019129f
C687 plus.n10 gnd 0.023096f
C688 plus.t22 gnd 0.388359f
C689 plus.t9 gnd 0.388359f
C690 plus.n11 gnd 0.180624f
C691 plus.t14 gnd 0.435248f
C692 plus.n12 gnd 0.182935f
C693 plus.n13 gnd 0.09858f
C694 plus.n14 gnd 0.029162f
C695 plus.n15 gnd 0.026568f
C696 plus.n16 gnd 0.15707f
C697 plus.n17 gnd 0.028346f
C698 plus.n18 gnd 0.023096f
C699 plus.n19 gnd 0.023096f
C700 plus.n20 gnd 0.023096f
C701 plus.n21 gnd 0.029941f
C702 plus.n22 gnd 0.15707f
C703 plus.n23 gnd 0.028297f
C704 plus.n24 gnd 0.027433f
C705 plus.n25 gnd 0.023096f
C706 plus.n26 gnd 0.023096f
C707 plus.n27 gnd 0.029381f
C708 plus.n28 gnd 0.018654f
C709 plus.n29 gnd 0.029381f
C710 plus.n30 gnd 0.023096f
C711 plus.n31 gnd 0.023096f
C712 plus.n32 gnd 0.027433f
C713 plus.n33 gnd 0.028297f
C714 plus.n34 gnd 0.15707f
C715 plus.n35 gnd 0.029941f
C716 plus.n36 gnd 0.023096f
C717 plus.n37 gnd 0.023096f
C718 plus.n38 gnd 0.023096f
C719 plus.n39 gnd 0.028346f
C720 plus.n40 gnd 0.15707f
C721 plus.n41 gnd 0.026568f
C722 plus.n42 gnd 0.029162f
C723 plus.n43 gnd 0.023096f
C724 plus.n44 gnd 0.023096f
C725 plus.n45 gnd 0.03014f
C726 plus.n46 gnd 0.008945f
C727 plus.n47 gnd 0.182145f
C728 plus.n48 gnd 0.265033f
C729 plus.n49 gnd 0.023096f
C730 plus.t10 gnd 0.388359f
C731 plus.n50 gnd 0.15707f
C732 plus.n51 gnd 0.023096f
C733 plus.t15 gnd 0.388359f
C734 plus.n52 gnd 0.019129f
C735 plus.n53 gnd 0.023096f
C736 plus.t13 gnd 0.388359f
C737 plus.t17 gnd 0.388359f
C738 plus.n54 gnd 0.15707f
C739 plus.n55 gnd 0.023096f
C740 plus.t16 gnd 0.388359f
C741 plus.n56 gnd 0.15707f
C742 plus.n57 gnd 0.023096f
C743 plus.t20 gnd 0.388359f
C744 plus.n58 gnd 0.019129f
C745 plus.n59 gnd 0.023096f
C746 plus.t21 gnd 0.388359f
C747 plus.t5 gnd 0.388359f
C748 plus.n60 gnd 0.180624f
C749 plus.t11 gnd 0.435248f
C750 plus.n61 gnd 0.182935f
C751 plus.n62 gnd 0.09858f
C752 plus.n63 gnd 0.029162f
C753 plus.n64 gnd 0.026568f
C754 plus.n65 gnd 0.15707f
C755 plus.n66 gnd 0.028346f
C756 plus.n67 gnd 0.023096f
C757 plus.n68 gnd 0.023096f
C758 plus.n69 gnd 0.023096f
C759 plus.n70 gnd 0.029941f
C760 plus.n71 gnd 0.15707f
C761 plus.n72 gnd 0.028297f
C762 plus.n73 gnd 0.027433f
C763 plus.n74 gnd 0.023096f
C764 plus.n75 gnd 0.023096f
C765 plus.n76 gnd 0.029381f
C766 plus.n77 gnd 0.018654f
C767 plus.n78 gnd 0.029381f
C768 plus.n79 gnd 0.023096f
C769 plus.n80 gnd 0.023096f
C770 plus.n81 gnd 0.027433f
C771 plus.n82 gnd 0.028297f
C772 plus.n83 gnd 0.15707f
C773 plus.n84 gnd 0.029941f
C774 plus.n85 gnd 0.023096f
C775 plus.n86 gnd 0.023096f
C776 plus.n87 gnd 0.023096f
C777 plus.n88 gnd 0.028346f
C778 plus.n89 gnd 0.15707f
C779 plus.n90 gnd 0.026568f
C780 plus.n91 gnd 0.029162f
C781 plus.n92 gnd 0.023096f
C782 plus.n93 gnd 0.023096f
C783 plus.n94 gnd 0.03014f
C784 plus.n95 gnd 0.008945f
C785 plus.t23 gnd 0.42001f
C786 plus.n96 gnd 0.182145f
C787 plus.n97 gnd 0.771394f
C788 plus.n98 gnd 1.15097f
C789 plus.t1 gnd 0.039871f
C790 plus.t2 gnd 0.00712f
C791 plus.t4 gnd 0.00712f
C792 plus.n99 gnd 0.023091f
C793 plus.n100 gnd 0.179258f
C794 plus.t0 gnd 0.00712f
C795 plus.t3 gnd 0.00712f
C796 plus.n101 gnd 0.023091f
C797 plus.n102 gnd 0.134555f
C798 plus.n103 gnd 2.47485f
C799 commonsourceibias.n0 gnd 0.010301f
C800 commonsourceibias.t71 gnd 0.155981f
C801 commonsourceibias.t81 gnd 0.144227f
C802 commonsourceibias.n1 gnd 0.057546f
C803 commonsourceibias.n2 gnd 0.00772f
C804 commonsourceibias.t55 gnd 0.144227f
C805 commonsourceibias.n3 gnd 0.006245f
C806 commonsourceibias.n4 gnd 0.00772f
C807 commonsourceibias.t53 gnd 0.144227f
C808 commonsourceibias.n5 gnd 0.007453f
C809 commonsourceibias.n6 gnd 0.00772f
C810 commonsourceibias.t76 gnd 0.144227f
C811 commonsourceibias.n7 gnd 0.057546f
C812 commonsourceibias.t86 gnd 0.144227f
C813 commonsourceibias.n8 gnd 0.006235f
C814 commonsourceibias.n9 gnd 0.010301f
C815 commonsourceibias.t32 gnd 0.155981f
C816 commonsourceibias.t14 gnd 0.144227f
C817 commonsourceibias.n10 gnd 0.057546f
C818 commonsourceibias.n11 gnd 0.00772f
C819 commonsourceibias.t24 gnd 0.144227f
C820 commonsourceibias.n12 gnd 0.006245f
C821 commonsourceibias.n13 gnd 0.00772f
C822 commonsourceibias.t30 gnd 0.144227f
C823 commonsourceibias.n14 gnd 0.007453f
C824 commonsourceibias.n15 gnd 0.00772f
C825 commonsourceibias.t20 gnd 0.144227f
C826 commonsourceibias.n16 gnd 0.057546f
C827 commonsourceibias.t36 gnd 0.144227f
C828 commonsourceibias.n17 gnd 0.006235f
C829 commonsourceibias.n18 gnd 0.00772f
C830 commonsourceibias.t44 gnd 0.144227f
C831 commonsourceibias.t26 gnd 0.144227f
C832 commonsourceibias.n19 gnd 0.057546f
C833 commonsourceibias.n20 gnd 0.00772f
C834 commonsourceibias.t34 gnd 0.144227f
C835 commonsourceibias.n21 gnd 0.057546f
C836 commonsourceibias.n22 gnd 0.00772f
C837 commonsourceibias.t10 gnd 0.144227f
C838 commonsourceibias.n23 gnd 0.057546f
C839 commonsourceibias.n24 gnd 0.038863f
C840 commonsourceibias.t40 gnd 0.144227f
C841 commonsourceibias.t46 gnd 0.162743f
C842 commonsourceibias.n25 gnd 0.066782f
C843 commonsourceibias.n26 gnd 0.069137f
C844 commonsourceibias.n27 gnd 0.009515f
C845 commonsourceibias.n28 gnd 0.010526f
C846 commonsourceibias.n29 gnd 0.00772f
C847 commonsourceibias.n30 gnd 0.00772f
C848 commonsourceibias.n31 gnd 0.010457f
C849 commonsourceibias.n32 gnd 0.006245f
C850 commonsourceibias.n33 gnd 0.010587f
C851 commonsourceibias.n34 gnd 0.00772f
C852 commonsourceibias.n35 gnd 0.00772f
C853 commonsourceibias.n36 gnd 0.010651f
C854 commonsourceibias.n37 gnd 0.009185f
C855 commonsourceibias.n38 gnd 0.007453f
C856 commonsourceibias.n39 gnd 0.00772f
C857 commonsourceibias.n40 gnd 0.00772f
C858 commonsourceibias.n41 gnd 0.009442f
C859 commonsourceibias.n42 gnd 0.010598f
C860 commonsourceibias.n43 gnd 0.057546f
C861 commonsourceibias.n44 gnd 0.010527f
C862 commonsourceibias.n45 gnd 0.00772f
C863 commonsourceibias.n46 gnd 0.00772f
C864 commonsourceibias.n47 gnd 0.00772f
C865 commonsourceibias.n48 gnd 0.010527f
C866 commonsourceibias.n49 gnd 0.057546f
C867 commonsourceibias.n50 gnd 0.010598f
C868 commonsourceibias.n51 gnd 0.009442f
C869 commonsourceibias.n52 gnd 0.00772f
C870 commonsourceibias.n53 gnd 0.00772f
C871 commonsourceibias.n54 gnd 0.00772f
C872 commonsourceibias.n55 gnd 0.009185f
C873 commonsourceibias.n56 gnd 0.010651f
C874 commonsourceibias.n57 gnd 0.057546f
C875 commonsourceibias.n58 gnd 0.010587f
C876 commonsourceibias.n59 gnd 0.00772f
C877 commonsourceibias.n60 gnd 0.00772f
C878 commonsourceibias.n61 gnd 0.00772f
C879 commonsourceibias.n62 gnd 0.010457f
C880 commonsourceibias.n63 gnd 0.057546f
C881 commonsourceibias.n64 gnd 0.010526f
C882 commonsourceibias.n65 gnd 0.009515f
C883 commonsourceibias.n66 gnd 0.00772f
C884 commonsourceibias.n67 gnd 0.00772f
C885 commonsourceibias.n68 gnd 0.007831f
C886 commonsourceibias.n69 gnd 0.008096f
C887 commonsourceibias.n70 gnd 0.068855f
C888 commonsourceibias.n71 gnd 0.076384f
C889 commonsourceibias.t33 gnd 0.016658f
C890 commonsourceibias.t15 gnd 0.016658f
C891 commonsourceibias.n72 gnd 0.147197f
C892 commonsourceibias.n73 gnd 0.12719f
C893 commonsourceibias.t25 gnd 0.016658f
C894 commonsourceibias.t31 gnd 0.016658f
C895 commonsourceibias.n74 gnd 0.147197f
C896 commonsourceibias.n75 gnd 0.067614f
C897 commonsourceibias.t21 gnd 0.016658f
C898 commonsourceibias.t37 gnd 0.016658f
C899 commonsourceibias.n76 gnd 0.147197f
C900 commonsourceibias.n77 gnd 0.056488f
C901 commonsourceibias.t41 gnd 0.016658f
C902 commonsourceibias.t47 gnd 0.016658f
C903 commonsourceibias.n78 gnd 0.14769f
C904 commonsourceibias.t35 gnd 0.016658f
C905 commonsourceibias.t11 gnd 0.016658f
C906 commonsourceibias.n79 gnd 0.147197f
C907 commonsourceibias.n80 gnd 0.13716f
C908 commonsourceibias.t45 gnd 0.016658f
C909 commonsourceibias.t27 gnd 0.016658f
C910 commonsourceibias.n81 gnd 0.147197f
C911 commonsourceibias.n82 gnd 0.056488f
C912 commonsourceibias.n83 gnd 0.068401f
C913 commonsourceibias.n84 gnd 0.00772f
C914 commonsourceibias.t50 gnd 0.144227f
C915 commonsourceibias.t69 gnd 0.144227f
C916 commonsourceibias.n85 gnd 0.057546f
C917 commonsourceibias.n86 gnd 0.00772f
C918 commonsourceibias.t67 gnd 0.144227f
C919 commonsourceibias.n87 gnd 0.057546f
C920 commonsourceibias.n88 gnd 0.00772f
C921 commonsourceibias.t78 gnd 0.144227f
C922 commonsourceibias.n89 gnd 0.057546f
C923 commonsourceibias.n90 gnd 0.038863f
C924 commonsourceibias.t64 gnd 0.144227f
C925 commonsourceibias.t62 gnd 0.162743f
C926 commonsourceibias.n91 gnd 0.066782f
C927 commonsourceibias.n92 gnd 0.069137f
C928 commonsourceibias.n93 gnd 0.009515f
C929 commonsourceibias.n94 gnd 0.010526f
C930 commonsourceibias.n95 gnd 0.00772f
C931 commonsourceibias.n96 gnd 0.00772f
C932 commonsourceibias.n97 gnd 0.010457f
C933 commonsourceibias.n98 gnd 0.006245f
C934 commonsourceibias.n99 gnd 0.010587f
C935 commonsourceibias.n100 gnd 0.00772f
C936 commonsourceibias.n101 gnd 0.00772f
C937 commonsourceibias.n102 gnd 0.010651f
C938 commonsourceibias.n103 gnd 0.009185f
C939 commonsourceibias.n104 gnd 0.007453f
C940 commonsourceibias.n105 gnd 0.00772f
C941 commonsourceibias.n106 gnd 0.00772f
C942 commonsourceibias.n107 gnd 0.009442f
C943 commonsourceibias.n108 gnd 0.010598f
C944 commonsourceibias.n109 gnd 0.057546f
C945 commonsourceibias.n110 gnd 0.010527f
C946 commonsourceibias.n111 gnd 0.007683f
C947 commonsourceibias.n112 gnd 0.055804f
C948 commonsourceibias.n113 gnd 0.007683f
C949 commonsourceibias.n114 gnd 0.010527f
C950 commonsourceibias.n115 gnd 0.057546f
C951 commonsourceibias.n116 gnd 0.010598f
C952 commonsourceibias.n117 gnd 0.009442f
C953 commonsourceibias.n118 gnd 0.00772f
C954 commonsourceibias.n119 gnd 0.00772f
C955 commonsourceibias.n120 gnd 0.00772f
C956 commonsourceibias.n121 gnd 0.009185f
C957 commonsourceibias.n122 gnd 0.010651f
C958 commonsourceibias.n123 gnd 0.057546f
C959 commonsourceibias.n124 gnd 0.010587f
C960 commonsourceibias.n125 gnd 0.00772f
C961 commonsourceibias.n126 gnd 0.00772f
C962 commonsourceibias.n127 gnd 0.00772f
C963 commonsourceibias.n128 gnd 0.010457f
C964 commonsourceibias.n129 gnd 0.057546f
C965 commonsourceibias.n130 gnd 0.010526f
C966 commonsourceibias.n131 gnd 0.009515f
C967 commonsourceibias.n132 gnd 0.00772f
C968 commonsourceibias.n133 gnd 0.00772f
C969 commonsourceibias.n134 gnd 0.007831f
C970 commonsourceibias.n135 gnd 0.008096f
C971 commonsourceibias.n136 gnd 0.068855f
C972 commonsourceibias.n137 gnd 0.04456f
C973 commonsourceibias.n138 gnd 0.010301f
C974 commonsourceibias.t72 gnd 0.144227f
C975 commonsourceibias.n139 gnd 0.057546f
C976 commonsourceibias.n140 gnd 0.00772f
C977 commonsourceibias.t49 gnd 0.144227f
C978 commonsourceibias.n141 gnd 0.006245f
C979 commonsourceibias.n142 gnd 0.00772f
C980 commonsourceibias.t95 gnd 0.144227f
C981 commonsourceibias.n143 gnd 0.007453f
C982 commonsourceibias.n144 gnd 0.00772f
C983 commonsourceibias.t66 gnd 0.144227f
C984 commonsourceibias.n145 gnd 0.057546f
C985 commonsourceibias.t77 gnd 0.144227f
C986 commonsourceibias.n146 gnd 0.006235f
C987 commonsourceibias.n147 gnd 0.00772f
C988 commonsourceibias.t91 gnd 0.144227f
C989 commonsourceibias.t60 gnd 0.144227f
C990 commonsourceibias.n148 gnd 0.057546f
C991 commonsourceibias.n149 gnd 0.00772f
C992 commonsourceibias.t58 gnd 0.144227f
C993 commonsourceibias.n150 gnd 0.057546f
C994 commonsourceibias.n151 gnd 0.00772f
C995 commonsourceibias.t68 gnd 0.144227f
C996 commonsourceibias.n152 gnd 0.057546f
C997 commonsourceibias.n153 gnd 0.038863f
C998 commonsourceibias.t57 gnd 0.144227f
C999 commonsourceibias.t54 gnd 0.162743f
C1000 commonsourceibias.n154 gnd 0.066782f
C1001 commonsourceibias.n155 gnd 0.069137f
C1002 commonsourceibias.n156 gnd 0.009515f
C1003 commonsourceibias.n157 gnd 0.010526f
C1004 commonsourceibias.n158 gnd 0.00772f
C1005 commonsourceibias.n159 gnd 0.00772f
C1006 commonsourceibias.n160 gnd 0.010457f
C1007 commonsourceibias.n161 gnd 0.006245f
C1008 commonsourceibias.n162 gnd 0.010587f
C1009 commonsourceibias.n163 gnd 0.00772f
C1010 commonsourceibias.n164 gnd 0.00772f
C1011 commonsourceibias.n165 gnd 0.010651f
C1012 commonsourceibias.n166 gnd 0.009185f
C1013 commonsourceibias.n167 gnd 0.007453f
C1014 commonsourceibias.n168 gnd 0.00772f
C1015 commonsourceibias.n169 gnd 0.00772f
C1016 commonsourceibias.n170 gnd 0.009442f
C1017 commonsourceibias.n171 gnd 0.010598f
C1018 commonsourceibias.n172 gnd 0.057546f
C1019 commonsourceibias.n173 gnd 0.010527f
C1020 commonsourceibias.n174 gnd 0.00772f
C1021 commonsourceibias.n175 gnd 0.00772f
C1022 commonsourceibias.n176 gnd 0.00772f
C1023 commonsourceibias.n177 gnd 0.010527f
C1024 commonsourceibias.n178 gnd 0.057546f
C1025 commonsourceibias.n179 gnd 0.010598f
C1026 commonsourceibias.n180 gnd 0.009442f
C1027 commonsourceibias.n181 gnd 0.00772f
C1028 commonsourceibias.n182 gnd 0.00772f
C1029 commonsourceibias.n183 gnd 0.00772f
C1030 commonsourceibias.n184 gnd 0.009185f
C1031 commonsourceibias.n185 gnd 0.010651f
C1032 commonsourceibias.n186 gnd 0.057546f
C1033 commonsourceibias.n187 gnd 0.010587f
C1034 commonsourceibias.n188 gnd 0.00772f
C1035 commonsourceibias.n189 gnd 0.00772f
C1036 commonsourceibias.n190 gnd 0.00772f
C1037 commonsourceibias.n191 gnd 0.010457f
C1038 commonsourceibias.n192 gnd 0.057546f
C1039 commonsourceibias.n193 gnd 0.010526f
C1040 commonsourceibias.n194 gnd 0.009515f
C1041 commonsourceibias.n195 gnd 0.00772f
C1042 commonsourceibias.n196 gnd 0.00772f
C1043 commonsourceibias.n197 gnd 0.007831f
C1044 commonsourceibias.n198 gnd 0.008096f
C1045 commonsourceibias.t61 gnd 0.155981f
C1046 commonsourceibias.n199 gnd 0.068855f
C1047 commonsourceibias.n200 gnd 0.023432f
C1048 commonsourceibias.n201 gnd 0.388694f
C1049 commonsourceibias.n202 gnd 0.010301f
C1050 commonsourceibias.t84 gnd 0.155981f
C1051 commonsourceibias.t92 gnd 0.144227f
C1052 commonsourceibias.n203 gnd 0.057546f
C1053 commonsourceibias.n204 gnd 0.00772f
C1054 commonsourceibias.t51 gnd 0.144227f
C1055 commonsourceibias.n205 gnd 0.006245f
C1056 commonsourceibias.n206 gnd 0.00772f
C1057 commonsourceibias.t63 gnd 0.144227f
C1058 commonsourceibias.n207 gnd 0.007453f
C1059 commonsourceibias.n208 gnd 0.00772f
C1060 commonsourceibias.t48 gnd 0.144227f
C1061 commonsourceibias.n209 gnd 0.006235f
C1062 commonsourceibias.n210 gnd 0.00772f
C1063 commonsourceibias.t94 gnd 0.144227f
C1064 commonsourceibias.t83 gnd 0.144227f
C1065 commonsourceibias.n211 gnd 0.057546f
C1066 commonsourceibias.n212 gnd 0.00772f
C1067 commonsourceibias.t80 gnd 0.144227f
C1068 commonsourceibias.n213 gnd 0.057546f
C1069 commonsourceibias.n214 gnd 0.00772f
C1070 commonsourceibias.t90 gnd 0.144227f
C1071 commonsourceibias.n215 gnd 0.057546f
C1072 commonsourceibias.n216 gnd 0.038863f
C1073 commonsourceibias.t59 gnd 0.144227f
C1074 commonsourceibias.t75 gnd 0.162743f
C1075 commonsourceibias.n217 gnd 0.066782f
C1076 commonsourceibias.n218 gnd 0.069137f
C1077 commonsourceibias.n219 gnd 0.009515f
C1078 commonsourceibias.n220 gnd 0.010526f
C1079 commonsourceibias.n221 gnd 0.00772f
C1080 commonsourceibias.n222 gnd 0.00772f
C1081 commonsourceibias.n223 gnd 0.010457f
C1082 commonsourceibias.n224 gnd 0.006245f
C1083 commonsourceibias.n225 gnd 0.010587f
C1084 commonsourceibias.n226 gnd 0.00772f
C1085 commonsourceibias.n227 gnd 0.00772f
C1086 commonsourceibias.n228 gnd 0.010651f
C1087 commonsourceibias.n229 gnd 0.009185f
C1088 commonsourceibias.n230 gnd 0.007453f
C1089 commonsourceibias.n231 gnd 0.00772f
C1090 commonsourceibias.n232 gnd 0.00772f
C1091 commonsourceibias.n233 gnd 0.009442f
C1092 commonsourceibias.n234 gnd 0.010598f
C1093 commonsourceibias.n235 gnd 0.057546f
C1094 commonsourceibias.n236 gnd 0.010527f
C1095 commonsourceibias.n237 gnd 0.007683f
C1096 commonsourceibias.t17 gnd 0.016658f
C1097 commonsourceibias.t9 gnd 0.016658f
C1098 commonsourceibias.n238 gnd 0.14769f
C1099 commonsourceibias.t19 gnd 0.016658f
C1100 commonsourceibias.t5 gnd 0.016658f
C1101 commonsourceibias.n239 gnd 0.147197f
C1102 commonsourceibias.n240 gnd 0.13716f
C1103 commonsourceibias.t43 gnd 0.016658f
C1104 commonsourceibias.t13 gnd 0.016658f
C1105 commonsourceibias.n241 gnd 0.147197f
C1106 commonsourceibias.n242 gnd 0.056488f
C1107 commonsourceibias.n243 gnd 0.010301f
C1108 commonsourceibias.t22 gnd 0.144227f
C1109 commonsourceibias.n244 gnd 0.057546f
C1110 commonsourceibias.n245 gnd 0.00772f
C1111 commonsourceibias.t38 gnd 0.144227f
C1112 commonsourceibias.n246 gnd 0.006245f
C1113 commonsourceibias.n247 gnd 0.00772f
C1114 commonsourceibias.t0 gnd 0.144227f
C1115 commonsourceibias.n248 gnd 0.007453f
C1116 commonsourceibias.n249 gnd 0.00772f
C1117 commonsourceibias.t6 gnd 0.144227f
C1118 commonsourceibias.n250 gnd 0.006235f
C1119 commonsourceibias.n251 gnd 0.00772f
C1120 commonsourceibias.t12 gnd 0.144227f
C1121 commonsourceibias.t42 gnd 0.144227f
C1122 commonsourceibias.n252 gnd 0.057546f
C1123 commonsourceibias.n253 gnd 0.00772f
C1124 commonsourceibias.t4 gnd 0.144227f
C1125 commonsourceibias.n254 gnd 0.057546f
C1126 commonsourceibias.n255 gnd 0.00772f
C1127 commonsourceibias.t18 gnd 0.144227f
C1128 commonsourceibias.n256 gnd 0.057546f
C1129 commonsourceibias.n257 gnd 0.038863f
C1130 commonsourceibias.t8 gnd 0.144227f
C1131 commonsourceibias.t16 gnd 0.162743f
C1132 commonsourceibias.n258 gnd 0.066782f
C1133 commonsourceibias.n259 gnd 0.069137f
C1134 commonsourceibias.n260 gnd 0.009515f
C1135 commonsourceibias.n261 gnd 0.010526f
C1136 commonsourceibias.n262 gnd 0.00772f
C1137 commonsourceibias.n263 gnd 0.00772f
C1138 commonsourceibias.n264 gnd 0.010457f
C1139 commonsourceibias.n265 gnd 0.006245f
C1140 commonsourceibias.n266 gnd 0.010587f
C1141 commonsourceibias.n267 gnd 0.00772f
C1142 commonsourceibias.n268 gnd 0.00772f
C1143 commonsourceibias.n269 gnd 0.010651f
C1144 commonsourceibias.n270 gnd 0.009185f
C1145 commonsourceibias.n271 gnd 0.007453f
C1146 commonsourceibias.n272 gnd 0.00772f
C1147 commonsourceibias.n273 gnd 0.00772f
C1148 commonsourceibias.n274 gnd 0.009442f
C1149 commonsourceibias.n275 gnd 0.010598f
C1150 commonsourceibias.n276 gnd 0.057546f
C1151 commonsourceibias.n277 gnd 0.010527f
C1152 commonsourceibias.n278 gnd 0.00772f
C1153 commonsourceibias.n279 gnd 0.00772f
C1154 commonsourceibias.n280 gnd 0.00772f
C1155 commonsourceibias.n281 gnd 0.010527f
C1156 commonsourceibias.n282 gnd 0.057546f
C1157 commonsourceibias.n283 gnd 0.010598f
C1158 commonsourceibias.t28 gnd 0.144227f
C1159 commonsourceibias.n284 gnd 0.057546f
C1160 commonsourceibias.n285 gnd 0.009442f
C1161 commonsourceibias.n286 gnd 0.00772f
C1162 commonsourceibias.n287 gnd 0.00772f
C1163 commonsourceibias.n288 gnd 0.00772f
C1164 commonsourceibias.n289 gnd 0.009185f
C1165 commonsourceibias.n290 gnd 0.010651f
C1166 commonsourceibias.n291 gnd 0.057546f
C1167 commonsourceibias.n292 gnd 0.010587f
C1168 commonsourceibias.n293 gnd 0.00772f
C1169 commonsourceibias.n294 gnd 0.00772f
C1170 commonsourceibias.n295 gnd 0.00772f
C1171 commonsourceibias.n296 gnd 0.010457f
C1172 commonsourceibias.n297 gnd 0.057546f
C1173 commonsourceibias.n298 gnd 0.010526f
C1174 commonsourceibias.n299 gnd 0.009515f
C1175 commonsourceibias.n300 gnd 0.00772f
C1176 commonsourceibias.n301 gnd 0.00772f
C1177 commonsourceibias.n302 gnd 0.007831f
C1178 commonsourceibias.n303 gnd 0.008096f
C1179 commonsourceibias.t2 gnd 0.155981f
C1180 commonsourceibias.n304 gnd 0.068855f
C1181 commonsourceibias.n305 gnd 0.076384f
C1182 commonsourceibias.t23 gnd 0.016658f
C1183 commonsourceibias.t3 gnd 0.016658f
C1184 commonsourceibias.n306 gnd 0.147197f
C1185 commonsourceibias.n307 gnd 0.12719f
C1186 commonsourceibias.t1 gnd 0.016658f
C1187 commonsourceibias.t39 gnd 0.016658f
C1188 commonsourceibias.n308 gnd 0.147197f
C1189 commonsourceibias.n309 gnd 0.067614f
C1190 commonsourceibias.t7 gnd 0.016658f
C1191 commonsourceibias.t29 gnd 0.016658f
C1192 commonsourceibias.n310 gnd 0.147197f
C1193 commonsourceibias.n311 gnd 0.056488f
C1194 commonsourceibias.n312 gnd 0.068401f
C1195 commonsourceibias.n313 gnd 0.055804f
C1196 commonsourceibias.n314 gnd 0.007683f
C1197 commonsourceibias.n315 gnd 0.010527f
C1198 commonsourceibias.n316 gnd 0.057546f
C1199 commonsourceibias.n317 gnd 0.010598f
C1200 commonsourceibias.t88 gnd 0.144227f
C1201 commonsourceibias.n318 gnd 0.057546f
C1202 commonsourceibias.n319 gnd 0.009442f
C1203 commonsourceibias.n320 gnd 0.00772f
C1204 commonsourceibias.n321 gnd 0.00772f
C1205 commonsourceibias.n322 gnd 0.00772f
C1206 commonsourceibias.n323 gnd 0.009185f
C1207 commonsourceibias.n324 gnd 0.010651f
C1208 commonsourceibias.n325 gnd 0.057546f
C1209 commonsourceibias.n326 gnd 0.010587f
C1210 commonsourceibias.n327 gnd 0.00772f
C1211 commonsourceibias.n328 gnd 0.00772f
C1212 commonsourceibias.n329 gnd 0.00772f
C1213 commonsourceibias.n330 gnd 0.010457f
C1214 commonsourceibias.n331 gnd 0.057546f
C1215 commonsourceibias.n332 gnd 0.010526f
C1216 commonsourceibias.n333 gnd 0.009515f
C1217 commonsourceibias.n334 gnd 0.00772f
C1218 commonsourceibias.n335 gnd 0.00772f
C1219 commonsourceibias.n336 gnd 0.007831f
C1220 commonsourceibias.n337 gnd 0.008096f
C1221 commonsourceibias.n338 gnd 0.068855f
C1222 commonsourceibias.n339 gnd 0.04456f
C1223 commonsourceibias.n340 gnd 0.010301f
C1224 commonsourceibias.t85 gnd 0.144227f
C1225 commonsourceibias.n341 gnd 0.057546f
C1226 commonsourceibias.n342 gnd 0.00772f
C1227 commonsourceibias.t93 gnd 0.144227f
C1228 commonsourceibias.n343 gnd 0.006245f
C1229 commonsourceibias.n344 gnd 0.00772f
C1230 commonsourceibias.t56 gnd 0.144227f
C1231 commonsourceibias.n345 gnd 0.007453f
C1232 commonsourceibias.n346 gnd 0.00772f
C1233 commonsourceibias.t89 gnd 0.144227f
C1234 commonsourceibias.n347 gnd 0.006235f
C1235 commonsourceibias.n348 gnd 0.00772f
C1236 commonsourceibias.t87 gnd 0.144227f
C1237 commonsourceibias.t74 gnd 0.144227f
C1238 commonsourceibias.n349 gnd 0.057546f
C1239 commonsourceibias.n350 gnd 0.00772f
C1240 commonsourceibias.t70 gnd 0.144227f
C1241 commonsourceibias.n351 gnd 0.057546f
C1242 commonsourceibias.n352 gnd 0.00772f
C1243 commonsourceibias.t82 gnd 0.144227f
C1244 commonsourceibias.n353 gnd 0.057546f
C1245 commonsourceibias.n354 gnd 0.038863f
C1246 commonsourceibias.t52 gnd 0.144227f
C1247 commonsourceibias.t65 gnd 0.162743f
C1248 commonsourceibias.n355 gnd 0.066782f
C1249 commonsourceibias.n356 gnd 0.069137f
C1250 commonsourceibias.n357 gnd 0.009515f
C1251 commonsourceibias.n358 gnd 0.010526f
C1252 commonsourceibias.n359 gnd 0.00772f
C1253 commonsourceibias.n360 gnd 0.00772f
C1254 commonsourceibias.n361 gnd 0.010457f
C1255 commonsourceibias.n362 gnd 0.006245f
C1256 commonsourceibias.n363 gnd 0.010587f
C1257 commonsourceibias.n364 gnd 0.00772f
C1258 commonsourceibias.n365 gnd 0.00772f
C1259 commonsourceibias.n366 gnd 0.010651f
C1260 commonsourceibias.n367 gnd 0.009185f
C1261 commonsourceibias.n368 gnd 0.007453f
C1262 commonsourceibias.n369 gnd 0.00772f
C1263 commonsourceibias.n370 gnd 0.00772f
C1264 commonsourceibias.n371 gnd 0.009442f
C1265 commonsourceibias.n372 gnd 0.010598f
C1266 commonsourceibias.n373 gnd 0.057546f
C1267 commonsourceibias.n374 gnd 0.010527f
C1268 commonsourceibias.n375 gnd 0.00772f
C1269 commonsourceibias.n376 gnd 0.00772f
C1270 commonsourceibias.n377 gnd 0.00772f
C1271 commonsourceibias.n378 gnd 0.010527f
C1272 commonsourceibias.n379 gnd 0.057546f
C1273 commonsourceibias.n380 gnd 0.010598f
C1274 commonsourceibias.t79 gnd 0.144227f
C1275 commonsourceibias.n381 gnd 0.057546f
C1276 commonsourceibias.n382 gnd 0.009442f
C1277 commonsourceibias.n383 gnd 0.00772f
C1278 commonsourceibias.n384 gnd 0.00772f
C1279 commonsourceibias.n385 gnd 0.00772f
C1280 commonsourceibias.n386 gnd 0.009185f
C1281 commonsourceibias.n387 gnd 0.010651f
C1282 commonsourceibias.n388 gnd 0.057546f
C1283 commonsourceibias.n389 gnd 0.010587f
C1284 commonsourceibias.n390 gnd 0.00772f
C1285 commonsourceibias.n391 gnd 0.00772f
C1286 commonsourceibias.n392 gnd 0.00772f
C1287 commonsourceibias.n393 gnd 0.010457f
C1288 commonsourceibias.n394 gnd 0.057546f
C1289 commonsourceibias.n395 gnd 0.010526f
C1290 commonsourceibias.n396 gnd 0.009515f
C1291 commonsourceibias.n397 gnd 0.00772f
C1292 commonsourceibias.n398 gnd 0.00772f
C1293 commonsourceibias.n399 gnd 0.007831f
C1294 commonsourceibias.n400 gnd 0.008096f
C1295 commonsourceibias.t73 gnd 0.155981f
C1296 commonsourceibias.n401 gnd 0.068855f
C1297 commonsourceibias.n402 gnd 0.023432f
C1298 commonsourceibias.n403 gnd 0.212991f
C1299 commonsourceibias.n404 gnd 4.01312f
C1300 CSoutput.n0 gnd 0.04487f
C1301 CSoutput.t156 gnd 0.296805f
C1302 CSoutput.n1 gnd 0.134022f
C1303 CSoutput.n2 gnd 0.04487f
C1304 CSoutput.t161 gnd 0.296805f
C1305 CSoutput.n3 gnd 0.035563f
C1306 CSoutput.n4 gnd 0.04487f
C1307 CSoutput.t150 gnd 0.296805f
C1308 CSoutput.n5 gnd 0.030666f
C1309 CSoutput.n6 gnd 0.04487f
C1310 CSoutput.t159 gnd 0.296805f
C1311 CSoutput.t165 gnd 0.296805f
C1312 CSoutput.n7 gnd 0.132562f
C1313 CSoutput.n8 gnd 0.04487f
C1314 CSoutput.t163 gnd 0.296805f
C1315 CSoutput.n9 gnd 0.029239f
C1316 CSoutput.n10 gnd 0.04487f
C1317 CSoutput.t151 gnd 0.296805f
C1318 CSoutput.t162 gnd 0.296805f
C1319 CSoutput.n11 gnd 0.132562f
C1320 CSoutput.n12 gnd 0.04487f
C1321 CSoutput.t160 gnd 0.296805f
C1322 CSoutput.n13 gnd 0.030666f
C1323 CSoutput.n14 gnd 0.04487f
C1324 CSoutput.t149 gnd 0.296805f
C1325 CSoutput.t155 gnd 0.296805f
C1326 CSoutput.n15 gnd 0.132562f
C1327 CSoutput.n16 gnd 0.04487f
C1328 CSoutput.t158 gnd 0.296805f
C1329 CSoutput.n17 gnd 0.032753f
C1330 CSoutput.t145 gnd 0.35469f
C1331 CSoutput.t147 gnd 0.296805f
C1332 CSoutput.n18 gnd 0.16923f
C1333 CSoutput.n19 gnd 0.164211f
C1334 CSoutput.n20 gnd 0.190505f
C1335 CSoutput.n21 gnd 0.04487f
C1336 CSoutput.n22 gnd 0.037449f
C1337 CSoutput.n23 gnd 0.132562f
C1338 CSoutput.n24 gnd 0.0361f
C1339 CSoutput.n25 gnd 0.035563f
C1340 CSoutput.n26 gnd 0.04487f
C1341 CSoutput.n27 gnd 0.04487f
C1342 CSoutput.n28 gnd 0.037161f
C1343 CSoutput.n29 gnd 0.031551f
C1344 CSoutput.n30 gnd 0.135513f
C1345 CSoutput.n31 gnd 0.031985f
C1346 CSoutput.n32 gnd 0.04487f
C1347 CSoutput.n33 gnd 0.04487f
C1348 CSoutput.n34 gnd 0.04487f
C1349 CSoutput.n35 gnd 0.036765f
C1350 CSoutput.n36 gnd 0.132562f
C1351 CSoutput.n37 gnd 0.035161f
C1352 CSoutput.n38 gnd 0.036502f
C1353 CSoutput.n39 gnd 0.04487f
C1354 CSoutput.n40 gnd 0.04487f
C1355 CSoutput.n41 gnd 0.037441f
C1356 CSoutput.n42 gnd 0.034222f
C1357 CSoutput.n43 gnd 0.132562f
C1358 CSoutput.n44 gnd 0.035089f
C1359 CSoutput.n45 gnd 0.04487f
C1360 CSoutput.n46 gnd 0.04487f
C1361 CSoutput.n47 gnd 0.04487f
C1362 CSoutput.n48 gnd 0.035089f
C1363 CSoutput.n49 gnd 0.132562f
C1364 CSoutput.n50 gnd 0.034222f
C1365 CSoutput.n51 gnd 0.037441f
C1366 CSoutput.n52 gnd 0.04487f
C1367 CSoutput.n53 gnd 0.04487f
C1368 CSoutput.n54 gnd 0.036502f
C1369 CSoutput.n55 gnd 0.035161f
C1370 CSoutput.n56 gnd 0.132562f
C1371 CSoutput.n57 gnd 0.036765f
C1372 CSoutput.n58 gnd 0.04487f
C1373 CSoutput.n59 gnd 0.04487f
C1374 CSoutput.n60 gnd 0.04487f
C1375 CSoutput.n61 gnd 0.031985f
C1376 CSoutput.n62 gnd 0.135513f
C1377 CSoutput.n63 gnd 0.031551f
C1378 CSoutput.t144 gnd 0.296805f
C1379 CSoutput.n64 gnd 0.132562f
C1380 CSoutput.n65 gnd 0.037161f
C1381 CSoutput.n66 gnd 0.04487f
C1382 CSoutput.n67 gnd 0.04487f
C1383 CSoutput.n68 gnd 0.04487f
C1384 CSoutput.n69 gnd 0.0361f
C1385 CSoutput.n70 gnd 0.132562f
C1386 CSoutput.n71 gnd 0.037449f
C1387 CSoutput.n72 gnd 0.032753f
C1388 CSoutput.n73 gnd 0.04487f
C1389 CSoutput.n74 gnd 0.04487f
C1390 CSoutput.n75 gnd 0.033967f
C1391 CSoutput.n76 gnd 0.020173f
C1392 CSoutput.t148 gnd 0.333482f
C1393 CSoutput.n77 gnd 0.16566f
C1394 CSoutput.n78 gnd 0.708845f
C1395 CSoutput.t12 gnd 0.055969f
C1396 CSoutput.t61 gnd 0.055969f
C1397 CSoutput.n79 gnd 0.43333f
C1398 CSoutput.t16 gnd 0.055969f
C1399 CSoutput.t41 gnd 0.055969f
C1400 CSoutput.n80 gnd 0.432557f
C1401 CSoutput.n81 gnd 0.439045f
C1402 CSoutput.t100 gnd 0.055969f
C1403 CSoutput.t54 gnd 0.055969f
C1404 CSoutput.n82 gnd 0.432557f
C1405 CSoutput.n83 gnd 0.216343f
C1406 CSoutput.t19 gnd 0.055969f
C1407 CSoutput.t85 gnd 0.055969f
C1408 CSoutput.n84 gnd 0.432557f
C1409 CSoutput.n85 gnd 0.216343f
C1410 CSoutput.t26 gnd 0.055969f
C1411 CSoutput.t68 gnd 0.055969f
C1412 CSoutput.n86 gnd 0.432557f
C1413 CSoutput.n87 gnd 0.216343f
C1414 CSoutput.t45 gnd 0.055969f
C1415 CSoutput.t62 gnd 0.055969f
C1416 CSoutput.n88 gnd 0.432557f
C1417 CSoutput.n89 gnd 0.216343f
C1418 CSoutput.t57 gnd 0.055969f
C1419 CSoutput.t92 gnd 0.055969f
C1420 CSoutput.n90 gnd 0.432557f
C1421 CSoutput.n91 gnd 0.216343f
C1422 CSoutput.t32 gnd 0.055969f
C1423 CSoutput.t74 gnd 0.055969f
C1424 CSoutput.n92 gnd 0.432557f
C1425 CSoutput.n93 gnd 0.396723f
C1426 CSoutput.t30 gnd 0.055969f
C1427 CSoutput.t93 gnd 0.055969f
C1428 CSoutput.n94 gnd 0.43333f
C1429 CSoutput.t70 gnd 0.055969f
C1430 CSoutput.t67 gnd 0.055969f
C1431 CSoutput.n95 gnd 0.432557f
C1432 CSoutput.n96 gnd 0.439045f
C1433 CSoutput.t60 gnd 0.055969f
C1434 CSoutput.t28 gnd 0.055969f
C1435 CSoutput.n97 gnd 0.432557f
C1436 CSoutput.n98 gnd 0.216343f
C1437 CSoutput.t11 gnd 0.055969f
C1438 CSoutput.t59 gnd 0.055969f
C1439 CSoutput.n99 gnd 0.432557f
C1440 CSoutput.n100 gnd 0.216343f
C1441 CSoutput.t56 gnd 0.055969f
C1442 CSoutput.t27 gnd 0.055969f
C1443 CSoutput.n101 gnd 0.432557f
C1444 CSoutput.n102 gnd 0.216343f
C1445 CSoutput.t7 gnd 0.055969f
C1446 CSoutput.t8 gnd 0.055969f
C1447 CSoutput.n103 gnd 0.432557f
C1448 CSoutput.n104 gnd 0.216343f
C1449 CSoutput.t71 gnd 0.055969f
C1450 CSoutput.t42 gnd 0.055969f
C1451 CSoutput.n105 gnd 0.432557f
C1452 CSoutput.n106 gnd 0.216343f
C1453 CSoutput.t36 gnd 0.055969f
C1454 CSoutput.t6 gnd 0.055969f
C1455 CSoutput.n107 gnd 0.432557f
C1456 CSoutput.n108 gnd 0.322622f
C1457 CSoutput.n109 gnd 0.406824f
C1458 CSoutput.t46 gnd 0.055969f
C1459 CSoutput.t101 gnd 0.055969f
C1460 CSoutput.n110 gnd 0.43333f
C1461 CSoutput.t77 gnd 0.055969f
C1462 CSoutput.t78 gnd 0.055969f
C1463 CSoutput.n111 gnd 0.432557f
C1464 CSoutput.n112 gnd 0.439045f
C1465 CSoutput.t65 gnd 0.055969f
C1466 CSoutput.t44 gnd 0.055969f
C1467 CSoutput.n113 gnd 0.432557f
C1468 CSoutput.n114 gnd 0.216343f
C1469 CSoutput.t23 gnd 0.055969f
C1470 CSoutput.t66 gnd 0.055969f
C1471 CSoutput.n115 gnd 0.432557f
C1472 CSoutput.n116 gnd 0.216343f
C1473 CSoutput.t64 gnd 0.055969f
C1474 CSoutput.t40 gnd 0.055969f
C1475 CSoutput.n117 gnd 0.432557f
C1476 CSoutput.n118 gnd 0.216343f
C1477 CSoutput.t22 gnd 0.055969f
C1478 CSoutput.t21 gnd 0.055969f
C1479 CSoutput.n119 gnd 0.432557f
C1480 CSoutput.n120 gnd 0.216343f
C1481 CSoutput.t80 gnd 0.055969f
C1482 CSoutput.t52 gnd 0.055969f
C1483 CSoutput.n121 gnd 0.432557f
C1484 CSoutput.n122 gnd 0.216343f
C1485 CSoutput.t49 gnd 0.055969f
C1486 CSoutput.t18 gnd 0.055969f
C1487 CSoutput.n123 gnd 0.432557f
C1488 CSoutput.n124 gnd 0.322622f
C1489 CSoutput.n125 gnd 0.454725f
C1490 CSoutput.n126 gnd 7.8714f
C1491 CSoutput.n128 gnd 0.793741f
C1492 CSoutput.n129 gnd 0.595306f
C1493 CSoutput.n130 gnd 0.793741f
C1494 CSoutput.n131 gnd 0.793741f
C1495 CSoutput.n132 gnd 2.137f
C1496 CSoutput.n133 gnd 0.793741f
C1497 CSoutput.n134 gnd 0.793741f
C1498 CSoutput.t164 gnd 0.992176f
C1499 CSoutput.n135 gnd 0.793741f
C1500 CSoutput.n136 gnd 0.793741f
C1501 CSoutput.n140 gnd 0.793741f
C1502 CSoutput.n144 gnd 0.793741f
C1503 CSoutput.n145 gnd 0.793741f
C1504 CSoutput.n147 gnd 0.793741f
C1505 CSoutput.n152 gnd 0.793741f
C1506 CSoutput.n154 gnd 0.793741f
C1507 CSoutput.n155 gnd 0.793741f
C1508 CSoutput.n157 gnd 0.793741f
C1509 CSoutput.n158 gnd 0.793741f
C1510 CSoutput.n160 gnd 0.793741f
C1511 CSoutput.t153 gnd 13.2633f
C1512 CSoutput.n162 gnd 0.793741f
C1513 CSoutput.n163 gnd 0.595306f
C1514 CSoutput.n164 gnd 0.793741f
C1515 CSoutput.n165 gnd 0.793741f
C1516 CSoutput.n166 gnd 2.137f
C1517 CSoutput.n167 gnd 0.793741f
C1518 CSoutput.n168 gnd 0.793741f
C1519 CSoutput.t152 gnd 0.992176f
C1520 CSoutput.n169 gnd 0.793741f
C1521 CSoutput.n170 gnd 0.793741f
C1522 CSoutput.n174 gnd 0.793741f
C1523 CSoutput.n178 gnd 0.793741f
C1524 CSoutput.n179 gnd 0.793741f
C1525 CSoutput.n181 gnd 0.793741f
C1526 CSoutput.n186 gnd 0.793741f
C1527 CSoutput.n188 gnd 0.793741f
C1528 CSoutput.n189 gnd 0.793741f
C1529 CSoutput.n191 gnd 0.793741f
C1530 CSoutput.n192 gnd 0.793741f
C1531 CSoutput.n194 gnd 0.793741f
C1532 CSoutput.n195 gnd 0.595306f
C1533 CSoutput.n197 gnd 0.793741f
C1534 CSoutput.n198 gnd 0.595306f
C1535 CSoutput.n199 gnd 0.793741f
C1536 CSoutput.n200 gnd 0.793741f
C1537 CSoutput.n201 gnd 2.137f
C1538 CSoutput.n202 gnd 0.793741f
C1539 CSoutput.n203 gnd 0.793741f
C1540 CSoutput.t146 gnd 0.992176f
C1541 CSoutput.n204 gnd 0.793741f
C1542 CSoutput.n205 gnd 2.137f
C1543 CSoutput.n207 gnd 0.793741f
C1544 CSoutput.n208 gnd 0.793741f
C1545 CSoutput.n210 gnd 0.793741f
C1546 CSoutput.n211 gnd 0.793741f
C1547 CSoutput.t154 gnd 13.0472f
C1548 CSoutput.t157 gnd 13.2633f
C1549 CSoutput.n217 gnd 2.49008f
C1550 CSoutput.n218 gnd 10.1437f
C1551 CSoutput.n219 gnd 10.5681f
C1552 CSoutput.n224 gnd 2.69743f
C1553 CSoutput.n230 gnd 0.793741f
C1554 CSoutput.n232 gnd 0.793741f
C1555 CSoutput.n234 gnd 0.793741f
C1556 CSoutput.n236 gnd 0.793741f
C1557 CSoutput.n238 gnd 0.793741f
C1558 CSoutput.n244 gnd 0.793741f
C1559 CSoutput.n251 gnd 1.45621f
C1560 CSoutput.n252 gnd 1.45621f
C1561 CSoutput.n253 gnd 0.793741f
C1562 CSoutput.n254 gnd 0.793741f
C1563 CSoutput.n256 gnd 0.595306f
C1564 CSoutput.n257 gnd 0.509826f
C1565 CSoutput.n259 gnd 0.595306f
C1566 CSoutput.n260 gnd 0.509826f
C1567 CSoutput.n261 gnd 0.595306f
C1568 CSoutput.n263 gnd 0.793741f
C1569 CSoutput.n265 gnd 2.137f
C1570 CSoutput.n266 gnd 2.49008f
C1571 CSoutput.n267 gnd 9.32958f
C1572 CSoutput.n269 gnd 0.595306f
C1573 CSoutput.n270 gnd 1.53176f
C1574 CSoutput.n271 gnd 0.595306f
C1575 CSoutput.n273 gnd 0.793741f
C1576 CSoutput.n275 gnd 2.137f
C1577 CSoutput.n276 gnd 4.65472f
C1578 CSoutput.t79 gnd 0.055969f
C1579 CSoutput.t10 gnd 0.055969f
C1580 CSoutput.n277 gnd 0.43333f
C1581 CSoutput.t39 gnd 0.055969f
C1582 CSoutput.t17 gnd 0.055969f
C1583 CSoutput.n278 gnd 0.432557f
C1584 CSoutput.n279 gnd 0.439045f
C1585 CSoutput.t55 gnd 0.055969f
C1586 CSoutput.t33 gnd 0.055969f
C1587 CSoutput.n280 gnd 0.432557f
C1588 CSoutput.n281 gnd 0.216343f
C1589 CSoutput.t86 gnd 0.055969f
C1590 CSoutput.t20 gnd 0.055969f
C1591 CSoutput.n282 gnd 0.432557f
C1592 CSoutput.n283 gnd 0.216343f
C1593 CSoutput.t69 gnd 0.055969f
C1594 CSoutput.t24 gnd 0.055969f
C1595 CSoutput.n284 gnd 0.432557f
C1596 CSoutput.n285 gnd 0.216343f
C1597 CSoutput.t82 gnd 0.055969f
C1598 CSoutput.t43 gnd 0.055969f
C1599 CSoutput.n286 gnd 0.432557f
C1600 CSoutput.n287 gnd 0.216343f
C1601 CSoutput.t91 gnd 0.055969f
C1602 CSoutput.t58 gnd 0.055969f
C1603 CSoutput.n288 gnd 0.432557f
C1604 CSoutput.n289 gnd 0.216343f
C1605 CSoutput.t75 gnd 0.055969f
C1606 CSoutput.t35 gnd 0.055969f
C1607 CSoutput.n290 gnd 0.432557f
C1608 CSoutput.n291 gnd 0.396723f
C1609 CSoutput.t38 gnd 0.055969f
C1610 CSoutput.t90 gnd 0.055969f
C1611 CSoutput.n292 gnd 0.43333f
C1612 CSoutput.t31 gnd 0.055969f
C1613 CSoutput.t34 gnd 0.055969f
C1614 CSoutput.n293 gnd 0.432557f
C1615 CSoutput.n294 gnd 0.439045f
C1616 CSoutput.t88 gnd 0.055969f
C1617 CSoutput.t89 gnd 0.055969f
C1618 CSoutput.n295 gnd 0.432557f
C1619 CSoutput.n296 gnd 0.216343f
C1620 CSoutput.t15 gnd 0.055969f
C1621 CSoutput.t76 gnd 0.055969f
C1622 CSoutput.n297 gnd 0.432557f
C1623 CSoutput.n298 gnd 0.216343f
C1624 CSoutput.t87 gnd 0.055969f
C1625 CSoutput.t13 gnd 0.055969f
C1626 CSoutput.n299 gnd 0.432557f
C1627 CSoutput.n300 gnd 0.216343f
C1628 CSoutput.t53 gnd 0.055969f
C1629 CSoutput.t73 gnd 0.055969f
C1630 CSoutput.n301 gnd 0.432557f
C1631 CSoutput.n302 gnd 0.216343f
C1632 CSoutput.t95 gnd 0.055969f
C1633 CSoutput.t37 gnd 0.055969f
C1634 CSoutput.n303 gnd 0.432557f
C1635 CSoutput.n304 gnd 0.216343f
C1636 CSoutput.t72 gnd 0.055969f
C1637 CSoutput.t98 gnd 0.055969f
C1638 CSoutput.n305 gnd 0.432557f
C1639 CSoutput.n306 gnd 0.322622f
C1640 CSoutput.n307 gnd 0.406824f
C1641 CSoutput.t51 gnd 0.055969f
C1642 CSoutput.t99 gnd 0.055969f
C1643 CSoutput.n308 gnd 0.43333f
C1644 CSoutput.t47 gnd 0.055969f
C1645 CSoutput.t48 gnd 0.055969f
C1646 CSoutput.n309 gnd 0.432557f
C1647 CSoutput.n310 gnd 0.439045f
C1648 CSoutput.t96 gnd 0.055969f
C1649 CSoutput.t97 gnd 0.055969f
C1650 CSoutput.n311 gnd 0.432557f
C1651 CSoutput.n312 gnd 0.216343f
C1652 CSoutput.t29 gnd 0.055969f
C1653 CSoutput.t84 gnd 0.055969f
C1654 CSoutput.n313 gnd 0.432557f
C1655 CSoutput.n314 gnd 0.216343f
C1656 CSoutput.t94 gnd 0.055969f
C1657 CSoutput.t25 gnd 0.055969f
C1658 CSoutput.n315 gnd 0.432557f
C1659 CSoutput.n316 gnd 0.216343f
C1660 CSoutput.t63 gnd 0.055969f
C1661 CSoutput.t83 gnd 0.055969f
C1662 CSoutput.n317 gnd 0.432557f
C1663 CSoutput.n318 gnd 0.216343f
C1664 CSoutput.t9 gnd 0.055969f
C1665 CSoutput.t50 gnd 0.055969f
C1666 CSoutput.n319 gnd 0.432557f
C1667 CSoutput.n320 gnd 0.216343f
C1668 CSoutput.t81 gnd 0.055969f
C1669 CSoutput.t14 gnd 0.055969f
C1670 CSoutput.n321 gnd 0.432556f
C1671 CSoutput.n322 gnd 0.322623f
C1672 CSoutput.n323 gnd 0.454725f
C1673 CSoutput.n324 gnd 11.534699f
C1674 CSoutput.t114 gnd 0.048973f
C1675 CSoutput.t109 gnd 0.048973f
C1676 CSoutput.n325 gnd 0.434189f
C1677 CSoutput.t0 gnd 0.048973f
C1678 CSoutput.t103 gnd 0.048973f
C1679 CSoutput.n326 gnd 0.432741f
C1680 CSoutput.n327 gnd 0.403234f
C1681 CSoutput.t143 gnd 0.048973f
C1682 CSoutput.t137 gnd 0.048973f
C1683 CSoutput.n328 gnd 0.432741f
C1684 CSoutput.n329 gnd 0.198775f
C1685 CSoutput.t120 gnd 0.048973f
C1686 CSoutput.t125 gnd 0.048973f
C1687 CSoutput.n330 gnd 0.432741f
C1688 CSoutput.n331 gnd 0.198775f
C1689 CSoutput.t122 gnd 0.048973f
C1690 CSoutput.t142 gnd 0.048973f
C1691 CSoutput.n332 gnd 0.432741f
C1692 CSoutput.n333 gnd 0.198775f
C1693 CSoutput.t127 gnd 0.048973f
C1694 CSoutput.t107 gnd 0.048973f
C1695 CSoutput.n334 gnd 0.432741f
C1696 CSoutput.n335 gnd 0.366582f
C1697 CSoutput.t106 gnd 0.048973f
C1698 CSoutput.t115 gnd 0.048973f
C1699 CSoutput.n336 gnd 0.434189f
C1700 CSoutput.t139 gnd 0.048973f
C1701 CSoutput.t4 gnd 0.048973f
C1702 CSoutput.n337 gnd 0.432741f
C1703 CSoutput.n338 gnd 0.403234f
C1704 CSoutput.t108 gnd 0.048973f
C1705 CSoutput.t129 gnd 0.048973f
C1706 CSoutput.n339 gnd 0.432741f
C1707 CSoutput.n340 gnd 0.198775f
C1708 CSoutput.t112 gnd 0.048973f
C1709 CSoutput.t111 gnd 0.048973f
C1710 CSoutput.n341 gnd 0.432741f
C1711 CSoutput.n342 gnd 0.198775f
C1712 CSoutput.t140 gnd 0.048973f
C1713 CSoutput.t102 gnd 0.048973f
C1714 CSoutput.n343 gnd 0.432741f
C1715 CSoutput.n344 gnd 0.198775f
C1716 CSoutput.t104 gnd 0.048973f
C1717 CSoutput.t121 gnd 0.048973f
C1718 CSoutput.n345 gnd 0.432741f
C1719 CSoutput.n346 gnd 0.301783f
C1720 CSoutput.n347 gnd 0.560736f
C1721 CSoutput.n348 gnd 11.547501f
C1722 CSoutput.t133 gnd 0.048973f
C1723 CSoutput.t105 gnd 0.048973f
C1724 CSoutput.n349 gnd 0.434189f
C1725 CSoutput.t117 gnd 0.048973f
C1726 CSoutput.t110 gnd 0.048973f
C1727 CSoutput.n350 gnd 0.432741f
C1728 CSoutput.n351 gnd 0.403234f
C1729 CSoutput.t118 gnd 0.048973f
C1730 CSoutput.t132 gnd 0.048973f
C1731 CSoutput.n352 gnd 0.432741f
C1732 CSoutput.n353 gnd 0.198775f
C1733 CSoutput.t2 gnd 0.048973f
C1734 CSoutput.t3 gnd 0.048973f
C1735 CSoutput.n354 gnd 0.432741f
C1736 CSoutput.n355 gnd 0.198775f
C1737 CSoutput.t134 gnd 0.048973f
C1738 CSoutput.t124 gnd 0.048973f
C1739 CSoutput.n356 gnd 0.432741f
C1740 CSoutput.n357 gnd 0.198775f
C1741 CSoutput.t130 gnd 0.048973f
C1742 CSoutput.t126 gnd 0.048973f
C1743 CSoutput.n358 gnd 0.432741f
C1744 CSoutput.n359 gnd 0.366582f
C1745 CSoutput.t138 gnd 0.048973f
C1746 CSoutput.t128 gnd 0.048973f
C1747 CSoutput.n360 gnd 0.434189f
C1748 CSoutput.t119 gnd 0.048973f
C1749 CSoutput.t5 gnd 0.048973f
C1750 CSoutput.n361 gnd 0.432741f
C1751 CSoutput.n362 gnd 0.403234f
C1752 CSoutput.t135 gnd 0.048973f
C1753 CSoutput.t131 gnd 0.048973f
C1754 CSoutput.n363 gnd 0.432741f
C1755 CSoutput.n364 gnd 0.198775f
C1756 CSoutput.t141 gnd 0.048973f
C1757 CSoutput.t136 gnd 0.048973f
C1758 CSoutput.n365 gnd 0.432741f
C1759 CSoutput.n366 gnd 0.198775f
C1760 CSoutput.t116 gnd 0.048973f
C1761 CSoutput.t123 gnd 0.048973f
C1762 CSoutput.n367 gnd 0.432741f
C1763 CSoutput.n368 gnd 0.198775f
C1764 CSoutput.t113 gnd 0.048973f
C1765 CSoutput.t1 gnd 0.048973f
C1766 CSoutput.n369 gnd 0.432741f
C1767 CSoutput.n370 gnd 0.301783f
C1768 CSoutput.n371 gnd 0.560736f
C1769 CSoutput.n372 gnd 6.53058f
C1770 CSoutput.n373 gnd 14.2841f
C1771 a_n8300_8799.n0 gnd 0.874504f
C1772 a_n8300_8799.n1 gnd 3.59374f
C1773 a_n8300_8799.n2 gnd 3.33612f
C1774 a_n8300_8799.n3 gnd 1.65793f
C1775 a_n8300_8799.n4 gnd 0.206879f
C1776 a_n8300_8799.n5 gnd 0.289153f
C1777 a_n8300_8799.n6 gnd 0.206879f
C1778 a_n8300_8799.n7 gnd 0.206879f
C1779 a_n8300_8799.n8 gnd 0.206879f
C1780 a_n8300_8799.n9 gnd 0.272554f
C1781 a_n8300_8799.n10 gnd 0.206879f
C1782 a_n8300_8799.n11 gnd 0.289153f
C1783 a_n8300_8799.n12 gnd 0.206879f
C1784 a_n8300_8799.n13 gnd 0.206879f
C1785 a_n8300_8799.n14 gnd 0.206879f
C1786 a_n8300_8799.n15 gnd 0.272554f
C1787 a_n8300_8799.n16 gnd 0.206879f
C1788 a_n8300_8799.n17 gnd 0.453159f
C1789 a_n8300_8799.n18 gnd 0.206879f
C1790 a_n8300_8799.n19 gnd 0.206879f
C1791 a_n8300_8799.n20 gnd 0.206879f
C1792 a_n8300_8799.n21 gnd 0.272554f
C1793 a_n8300_8799.n22 gnd 0.324274f
C1794 a_n8300_8799.n23 gnd 0.206879f
C1795 a_n8300_8799.n24 gnd 0.206879f
C1796 a_n8300_8799.n25 gnd 0.206879f
C1797 a_n8300_8799.n26 gnd 0.206879f
C1798 a_n8300_8799.n27 gnd 0.237433f
C1799 a_n8300_8799.n28 gnd 0.324274f
C1800 a_n8300_8799.n29 gnd 0.206879f
C1801 a_n8300_8799.n30 gnd 0.206879f
C1802 a_n8300_8799.n31 gnd 0.206879f
C1803 a_n8300_8799.n32 gnd 0.206879f
C1804 a_n8300_8799.n33 gnd 0.237433f
C1805 a_n8300_8799.n34 gnd 0.324274f
C1806 a_n8300_8799.n35 gnd 0.206879f
C1807 a_n8300_8799.n36 gnd 0.206879f
C1808 a_n8300_8799.n37 gnd 0.206879f
C1809 a_n8300_8799.n38 gnd 0.206879f
C1810 a_n8300_8799.n39 gnd 0.401439f
C1811 a_n8300_8799.n40 gnd 1.51626f
C1812 a_n8300_8799.n41 gnd 3.95f
C1813 a_n8300_8799.n42 gnd 2.73798f
C1814 a_n8300_8799.n43 gnd 1.51625f
C1815 a_n8300_8799.n44 gnd 0.008581f
C1816 a_n8300_8799.n45 gnd 0.001152f
C1817 a_n8300_8799.n47 gnd 0.007706f
C1818 a_n8300_8799.n48 gnd 0.011647f
C1819 a_n8300_8799.n49 gnd 0.00801f
C1820 a_n8300_8799.n51 gnd 4e-19
C1821 a_n8300_8799.n52 gnd 0.008301f
C1822 a_n8300_8799.n53 gnd 0.011465f
C1823 a_n8300_8799.n54 gnd 0.007388f
C1824 a_n8300_8799.n55 gnd 0.008581f
C1825 a_n8300_8799.n56 gnd 0.001152f
C1826 a_n8300_8799.n58 gnd 0.007706f
C1827 a_n8300_8799.n59 gnd 0.011647f
C1828 a_n8300_8799.n60 gnd 0.00801f
C1829 a_n8300_8799.n62 gnd 4e-19
C1830 a_n8300_8799.n63 gnd 0.008301f
C1831 a_n8300_8799.n64 gnd 0.011465f
C1832 a_n8300_8799.n65 gnd 0.007388f
C1833 a_n8300_8799.n66 gnd 0.008581f
C1834 a_n8300_8799.n67 gnd 0.001152f
C1835 a_n8300_8799.n69 gnd 0.007706f
C1836 a_n8300_8799.n70 gnd 0.011647f
C1837 a_n8300_8799.n71 gnd 0.00801f
C1838 a_n8300_8799.n73 gnd 4e-19
C1839 a_n8300_8799.n74 gnd 0.008301f
C1840 a_n8300_8799.n75 gnd 0.011465f
C1841 a_n8300_8799.n76 gnd 0.007388f
C1842 a_n8300_8799.n77 gnd 0.001152f
C1843 a_n8300_8799.n79 gnd 0.007706f
C1844 a_n8300_8799.n80 gnd 0.011647f
C1845 a_n8300_8799.n81 gnd 0.00801f
C1846 a_n8300_8799.n83 gnd 4e-19
C1847 a_n8300_8799.n84 gnd 0.008301f
C1848 a_n8300_8799.n85 gnd 0.011465f
C1849 a_n8300_8799.n86 gnd 0.007388f
C1850 a_n8300_8799.n87 gnd 0.249062f
C1851 a_n8300_8799.n88 gnd 0.001152f
C1852 a_n8300_8799.n90 gnd 0.007706f
C1853 a_n8300_8799.n91 gnd 0.011647f
C1854 a_n8300_8799.n92 gnd 0.00801f
C1855 a_n8300_8799.n94 gnd 4e-19
C1856 a_n8300_8799.n95 gnd 0.008301f
C1857 a_n8300_8799.n96 gnd 0.011465f
C1858 a_n8300_8799.n97 gnd 0.007388f
C1859 a_n8300_8799.n98 gnd 0.249062f
C1860 a_n8300_8799.n99 gnd 0.001152f
C1861 a_n8300_8799.n101 gnd 0.007706f
C1862 a_n8300_8799.n102 gnd 0.011647f
C1863 a_n8300_8799.n103 gnd 0.00801f
C1864 a_n8300_8799.n105 gnd 4e-19
C1865 a_n8300_8799.n106 gnd 0.008301f
C1866 a_n8300_8799.n107 gnd 0.011465f
C1867 a_n8300_8799.n108 gnd 0.007388f
C1868 a_n8300_8799.n109 gnd 0.249062f
C1869 a_n8300_8799.t28 gnd 0.143493f
C1870 a_n8300_8799.t11 gnd 0.143493f
C1871 a_n8300_8799.t14 gnd 0.143493f
C1872 a_n8300_8799.n110 gnd 1.13176f
C1873 a_n8300_8799.t17 gnd 0.143493f
C1874 a_n8300_8799.t10 gnd 0.143493f
C1875 a_n8300_8799.n111 gnd 1.13175f
C1876 a_n8300_8799.t23 gnd 0.143493f
C1877 a_n8300_8799.t24 gnd 0.143493f
C1878 a_n8300_8799.n112 gnd 1.12989f
C1879 a_n8300_8799.t18 gnd 0.143493f
C1880 a_n8300_8799.t26 gnd 0.143493f
C1881 a_n8300_8799.n113 gnd 1.12989f
C1882 a_n8300_8799.t12 gnd 0.143493f
C1883 a_n8300_8799.t25 gnd 0.143493f
C1884 a_n8300_8799.n114 gnd 1.12989f
C1885 a_n8300_8799.t22 gnd 0.143493f
C1886 a_n8300_8799.t19 gnd 0.143493f
C1887 a_n8300_8799.n115 gnd 1.12989f
C1888 a_n8300_8799.t0 gnd 0.111606f
C1889 a_n8300_8799.t39 gnd 0.111606f
C1890 a_n8300_8799.n116 gnd 0.989098f
C1891 a_n8300_8799.t7 gnd 0.111606f
C1892 a_n8300_8799.t32 gnd 0.111606f
C1893 a_n8300_8799.n117 gnd 0.98619f
C1894 a_n8300_8799.t30 gnd 0.111606f
C1895 a_n8300_8799.t5 gnd 0.111606f
C1896 a_n8300_8799.n118 gnd 0.98619f
C1897 a_n8300_8799.t33 gnd 0.111606f
C1898 a_n8300_8799.t38 gnd 0.111606f
C1899 a_n8300_8799.n119 gnd 0.989097f
C1900 a_n8300_8799.t34 gnd 0.111606f
C1901 a_n8300_8799.t35 gnd 0.111606f
C1902 a_n8300_8799.n120 gnd 0.986189f
C1903 a_n8300_8799.t1 gnd 0.111606f
C1904 a_n8300_8799.t2 gnd 0.111606f
C1905 a_n8300_8799.n121 gnd 0.986189f
C1906 a_n8300_8799.t8 gnd 0.111606f
C1907 a_n8300_8799.t37 gnd 0.111606f
C1908 a_n8300_8799.n122 gnd 0.989097f
C1909 a_n8300_8799.t36 gnd 0.111606f
C1910 a_n8300_8799.t6 gnd 0.111606f
C1911 a_n8300_8799.n123 gnd 0.986189f
C1912 a_n8300_8799.t3 gnd 0.111606f
C1913 a_n8300_8799.t29 gnd 0.111606f
C1914 a_n8300_8799.n124 gnd 0.98619f
C1915 a_n8300_8799.t31 gnd 0.111606f
C1916 a_n8300_8799.t4 gnd 0.111606f
C1917 a_n8300_8799.n125 gnd 0.98619f
C1918 a_n8300_8799.t63 gnd 0.594991f
C1919 a_n8300_8799.n126 gnd 0.266005f
C1920 a_n8300_8799.t97 gnd 0.594991f
C1921 a_n8300_8799.t118 gnd 0.594991f
C1922 a_n8300_8799.n127 gnd 0.269301f
C1923 a_n8300_8799.t75 gnd 0.594991f
C1924 a_n8300_8799.t77 gnd 0.594991f
C1925 a_n8300_8799.t89 gnd 0.594991f
C1926 a_n8300_8799.n128 gnd 0.271376f
C1927 a_n8300_8799.t119 gnd 0.594991f
C1928 a_n8300_8799.t123 gnd 0.594991f
C1929 a_n8300_8799.n129 gnd 0.264937f
C1930 a_n8300_8799.t92 gnd 0.606252f
C1931 a_n8300_8799.n130 gnd 0.249446f
C1932 a_n8300_8799.n131 gnd 0.011736f
C1933 a_n8300_8799.t61 gnd 0.594991f
C1934 a_n8300_8799.n132 gnd 0.265734f
C1935 a_n8300_8799.n133 gnd 0.269287f
C1936 a_n8300_8799.t120 gnd 0.594991f
C1937 a_n8300_8799.n134 gnd 0.265824f
C1938 a_n8300_8799.n135 gnd 0.260473f
C1939 a_n8300_8799.t101 gnd 0.594991f
C1940 a_n8300_8799.n136 gnd 0.265575f
C1941 a_n8300_8799.n137 gnd 0.271809f
C1942 a_n8300_8799.t76 gnd 0.594991f
C1943 a_n8300_8799.n138 gnd 0.269169f
C1944 a_n8300_8799.n139 gnd 0.265256f
C1945 a_n8300_8799.t64 gnd 0.594991f
C1946 a_n8300_8799.n140 gnd 0.260792f
C1947 a_n8300_8799.t95 gnd 0.594991f
C1948 a_n8300_8799.n141 gnd 0.269286f
C1949 a_n8300_8799.t40 gnd 0.606241f
C1950 a_n8300_8799.t74 gnd 0.594991f
C1951 a_n8300_8799.n142 gnd 0.266005f
C1952 a_n8300_8799.t113 gnd 0.594991f
C1953 a_n8300_8799.t130 gnd 0.594991f
C1954 a_n8300_8799.n143 gnd 0.269301f
C1955 a_n8300_8799.t82 gnd 0.594991f
C1956 a_n8300_8799.t85 gnd 0.594991f
C1957 a_n8300_8799.t99 gnd 0.594991f
C1958 a_n8300_8799.n144 gnd 0.271376f
C1959 a_n8300_8799.t134 gnd 0.594991f
C1960 a_n8300_8799.t135 gnd 0.594991f
C1961 a_n8300_8799.n145 gnd 0.264937f
C1962 a_n8300_8799.t105 gnd 0.606252f
C1963 a_n8300_8799.n146 gnd 0.249446f
C1964 a_n8300_8799.n147 gnd 0.011736f
C1965 a_n8300_8799.t70 gnd 0.594991f
C1966 a_n8300_8799.n148 gnd 0.265734f
C1967 a_n8300_8799.n149 gnd 0.269287f
C1968 a_n8300_8799.t133 gnd 0.594991f
C1969 a_n8300_8799.n150 gnd 0.265824f
C1970 a_n8300_8799.n151 gnd 0.260473f
C1971 a_n8300_8799.t114 gnd 0.594991f
C1972 a_n8300_8799.n152 gnd 0.265575f
C1973 a_n8300_8799.n153 gnd 0.271809f
C1974 a_n8300_8799.t81 gnd 0.594991f
C1975 a_n8300_8799.n154 gnd 0.269169f
C1976 a_n8300_8799.n155 gnd 0.265256f
C1977 a_n8300_8799.t71 gnd 0.594991f
C1978 a_n8300_8799.n156 gnd 0.260792f
C1979 a_n8300_8799.t111 gnd 0.594991f
C1980 a_n8300_8799.n157 gnd 0.269286f
C1981 a_n8300_8799.t48 gnd 0.606241f
C1982 a_n8300_8799.n158 gnd 0.896122f
C1983 a_n8300_8799.t100 gnd 0.594991f
C1984 a_n8300_8799.n159 gnd 0.266005f
C1985 a_n8300_8799.t87 gnd 0.594991f
C1986 a_n8300_8799.t122 gnd 0.594991f
C1987 a_n8300_8799.n160 gnd 0.269301f
C1988 a_n8300_8799.t56 gnd 0.594991f
C1989 a_n8300_8799.t115 gnd 0.594991f
C1990 a_n8300_8799.t49 gnd 0.594991f
C1991 a_n8300_8799.n161 gnd 0.271376f
C1992 a_n8300_8799.t96 gnd 0.594991f
C1993 a_n8300_8799.t67 gnd 0.594991f
C1994 a_n8300_8799.n162 gnd 0.264937f
C1995 a_n8300_8799.t109 gnd 0.606252f
C1996 a_n8300_8799.n163 gnd 0.249446f
C1997 a_n8300_8799.n164 gnd 0.011736f
C1998 a_n8300_8799.t84 gnd 0.594991f
C1999 a_n8300_8799.n165 gnd 0.265734f
C2000 a_n8300_8799.n166 gnd 0.269287f
C2001 a_n8300_8799.t79 gnd 0.594991f
C2002 a_n8300_8799.n167 gnd 0.265824f
C2003 a_n8300_8799.n168 gnd 0.260473f
C2004 a_n8300_8799.t73 gnd 0.594991f
C2005 a_n8300_8799.n169 gnd 0.265575f
C2006 a_n8300_8799.n170 gnd 0.271809f
C2007 a_n8300_8799.t41 gnd 0.594991f
C2008 a_n8300_8799.n171 gnd 0.269169f
C2009 a_n8300_8799.n172 gnd 0.265256f
C2010 a_n8300_8799.t125 gnd 0.594991f
C2011 a_n8300_8799.n173 gnd 0.260792f
C2012 a_n8300_8799.t129 gnd 0.594991f
C2013 a_n8300_8799.n174 gnd 0.269286f
C2014 a_n8300_8799.t80 gnd 0.606241f
C2015 a_n8300_8799.n175 gnd 1.74565f
C2016 a_n8300_8799.t90 gnd 0.594991f
C2017 a_n8300_8799.t42 gnd 0.594991f
C2018 a_n8300_8799.t94 gnd 0.594991f
C2019 a_n8300_8799.n176 gnd 0.26889f
C2020 a_n8300_8799.t93 gnd 0.594991f
C2021 a_n8300_8799.t45 gnd 0.594991f
C2022 a_n8300_8799.t44 gnd 0.594991f
C2023 a_n8300_8799.n177 gnd 0.265824f
C2024 a_n8300_8799.t112 gnd 0.594991f
C2025 a_n8300_8799.t57 gnd 0.594991f
C2026 a_n8300_8799.t47 gnd 0.594991f
C2027 a_n8300_8799.n178 gnd 0.269301f
C2028 a_n8300_8799.t116 gnd 0.594991f
C2029 a_n8300_8799.t78 gnd 0.594991f
C2030 a_n8300_8799.t58 gnd 0.594991f
C2031 a_n8300_8799.n179 gnd 0.265256f
C2032 a_n8300_8799.t132 gnd 0.594991f
C2033 a_n8300_8799.t91 gnd 0.594991f
C2034 a_n8300_8799.t60 gnd 0.594991f
C2035 a_n8300_8799.n180 gnd 0.269286f
C2036 a_n8300_8799.t127 gnd 0.606252f
C2037 a_n8300_8799.n181 gnd 0.249446f
C2038 a_n8300_8799.n182 gnd 0.266005f
C2039 a_n8300_8799.n183 gnd 0.260792f
C2040 a_n8300_8799.n184 gnd 0.269169f
C2041 a_n8300_8799.n185 gnd 0.271809f
C2042 a_n8300_8799.n186 gnd 0.265575f
C2043 a_n8300_8799.n187 gnd 0.260473f
C2044 a_n8300_8799.n188 gnd 0.269287f
C2045 a_n8300_8799.n189 gnd 0.271376f
C2046 a_n8300_8799.n190 gnd 0.264937f
C2047 a_n8300_8799.n191 gnd 0.260313f
C2048 a_n8300_8799.t103 gnd 0.594991f
C2049 a_n8300_8799.t51 gnd 0.594991f
C2050 a_n8300_8799.t110 gnd 0.594991f
C2051 a_n8300_8799.n192 gnd 0.26889f
C2052 a_n8300_8799.t107 gnd 0.594991f
C2053 a_n8300_8799.t53 gnd 0.594991f
C2054 a_n8300_8799.t52 gnd 0.594991f
C2055 a_n8300_8799.n193 gnd 0.265824f
C2056 a_n8300_8799.t126 gnd 0.594991f
C2057 a_n8300_8799.t65 gnd 0.594991f
C2058 a_n8300_8799.t54 gnd 0.594991f
C2059 a_n8300_8799.n194 gnd 0.269301f
C2060 a_n8300_8799.t128 gnd 0.594991f
C2061 a_n8300_8799.t88 gnd 0.594991f
C2062 a_n8300_8799.t68 gnd 0.594991f
C2063 a_n8300_8799.n195 gnd 0.265256f
C2064 a_n8300_8799.t46 gnd 0.594991f
C2065 a_n8300_8799.t104 gnd 0.594991f
C2066 a_n8300_8799.t69 gnd 0.594991f
C2067 a_n8300_8799.n196 gnd 0.269286f
C2068 a_n8300_8799.t43 gnd 0.606252f
C2069 a_n8300_8799.n197 gnd 0.249446f
C2070 a_n8300_8799.n198 gnd 0.266005f
C2071 a_n8300_8799.n199 gnd 0.260792f
C2072 a_n8300_8799.n200 gnd 0.269169f
C2073 a_n8300_8799.n201 gnd 0.271809f
C2074 a_n8300_8799.n202 gnd 0.265575f
C2075 a_n8300_8799.n203 gnd 0.260473f
C2076 a_n8300_8799.n204 gnd 0.269287f
C2077 a_n8300_8799.n205 gnd 0.271376f
C2078 a_n8300_8799.n206 gnd 0.264937f
C2079 a_n8300_8799.n207 gnd 0.260313f
C2080 a_n8300_8799.n208 gnd 0.896122f
C2081 a_n8300_8799.t62 gnd 0.594991f
C2082 a_n8300_8799.t131 gnd 0.594991f
C2083 a_n8300_8799.t102 gnd 0.594991f
C2084 a_n8300_8799.n209 gnd 0.26889f
C2085 a_n8300_8799.t124 gnd 0.594991f
C2086 a_n8300_8799.t86 gnd 0.594991f
C2087 a_n8300_8799.t108 gnd 0.594991f
C2088 a_n8300_8799.n210 gnd 0.265824f
C2089 a_n8300_8799.t55 gnd 0.594991f
C2090 a_n8300_8799.t121 gnd 0.594991f
C2091 a_n8300_8799.t72 gnd 0.594991f
C2092 a_n8300_8799.n211 gnd 0.269301f
C2093 a_n8300_8799.t117 gnd 0.594991f
C2094 a_n8300_8799.t59 gnd 0.594991f
C2095 a_n8300_8799.t98 gnd 0.594991f
C2096 a_n8300_8799.n212 gnd 0.265256f
C2097 a_n8300_8799.t50 gnd 0.594991f
C2098 a_n8300_8799.t83 gnd 0.594991f
C2099 a_n8300_8799.t66 gnd 0.594991f
C2100 a_n8300_8799.n213 gnd 0.269286f
C2101 a_n8300_8799.t106 gnd 0.606252f
C2102 a_n8300_8799.n214 gnd 0.249446f
C2103 a_n8300_8799.n215 gnd 0.266005f
C2104 a_n8300_8799.n216 gnd 0.260792f
C2105 a_n8300_8799.n217 gnd 0.269169f
C2106 a_n8300_8799.n218 gnd 0.271809f
C2107 a_n8300_8799.n219 gnd 0.265575f
C2108 a_n8300_8799.n220 gnd 0.260473f
C2109 a_n8300_8799.n221 gnd 0.269287f
C2110 a_n8300_8799.n222 gnd 0.271376f
C2111 a_n8300_8799.n223 gnd 0.264937f
C2112 a_n8300_8799.n224 gnd 0.260313f
C2113 a_n8300_8799.n225 gnd 1.27132f
C2114 a_n8300_8799.n226 gnd 15.599401f
C2115 a_n8300_8799.n227 gnd 4.35447f
C2116 a_n8300_8799.n228 gnd 6.95472f
C2117 a_n8300_8799.t21 gnd 0.143493f
C2118 a_n8300_8799.t15 gnd 0.143493f
C2119 a_n8300_8799.n229 gnd 1.12989f
C2120 a_n8300_8799.t27 gnd 0.143493f
C2121 a_n8300_8799.t20 gnd 0.143493f
C2122 a_n8300_8799.n230 gnd 1.12989f
C2123 a_n8300_8799.t16 gnd 0.143493f
C2124 a_n8300_8799.t13 gnd 0.143493f
C2125 a_n8300_8799.n231 gnd 1.12989f
C2126 a_n8300_8799.n232 gnd 1.12989f
C2127 a_n8300_8799.t9 gnd 0.143493f
C2128 vdd.t170 gnd 0.035882f
C2129 vdd.t151 gnd 0.035882f
C2130 vdd.n0 gnd 0.283008f
C2131 vdd.t132 gnd 0.035882f
C2132 vdd.t165 gnd 0.035882f
C2133 vdd.n1 gnd 0.28254f
C2134 vdd.n2 gnd 0.260556f
C2135 vdd.t148 gnd 0.035882f
C2136 vdd.t174 gnd 0.035882f
C2137 vdd.n3 gnd 0.28254f
C2138 vdd.n4 gnd 0.131773f
C2139 vdd.t176 gnd 0.035882f
C2140 vdd.t156 gnd 0.035882f
C2141 vdd.n5 gnd 0.28254f
C2142 vdd.n6 gnd 0.123645f
C2143 vdd.t180 gnd 0.035882f
C2144 vdd.t146 gnd 0.035882f
C2145 vdd.n7 gnd 0.283008f
C2146 vdd.t154 gnd 0.035882f
C2147 vdd.t172 gnd 0.035882f
C2148 vdd.n8 gnd 0.28254f
C2149 vdd.n9 gnd 0.260556f
C2150 vdd.t162 gnd 0.035882f
C2151 vdd.t135 gnd 0.035882f
C2152 vdd.n10 gnd 0.28254f
C2153 vdd.n11 gnd 0.131773f
C2154 vdd.t143 gnd 0.035882f
C2155 vdd.t160 gnd 0.035882f
C2156 vdd.n12 gnd 0.28254f
C2157 vdd.n13 gnd 0.123645f
C2158 vdd.n14 gnd 0.087414f
C2159 vdd.t271 gnd 0.019934f
C2160 vdd.t24 gnd 0.019934f
C2161 vdd.n15 gnd 0.183488f
C2162 vdd.t117 gnd 0.019934f
C2163 vdd.t191 gnd 0.019934f
C2164 vdd.n16 gnd 0.182952f
C2165 vdd.n17 gnd 0.318393f
C2166 vdd.t232 gnd 0.019934f
C2167 vdd.t229 gnd 0.019934f
C2168 vdd.n18 gnd 0.182952f
C2169 vdd.n19 gnd 0.131723f
C2170 vdd.t118 gnd 0.019934f
C2171 vdd.t23 gnd 0.019934f
C2172 vdd.n20 gnd 0.183488f
C2173 vdd.t231 gnd 0.019934f
C2174 vdd.t270 gnd 0.019934f
C2175 vdd.n21 gnd 0.182952f
C2176 vdd.n22 gnd 0.318393f
C2177 vdd.t228 gnd 0.019934f
C2178 vdd.t233 gnd 0.019934f
C2179 vdd.n23 gnd 0.182952f
C2180 vdd.n24 gnd 0.131723f
C2181 vdd.t192 gnd 0.019934f
C2182 vdd.t230 gnd 0.019934f
C2183 vdd.n25 gnd 0.182952f
C2184 vdd.t193 gnd 0.019934f
C2185 vdd.t190 gnd 0.019934f
C2186 vdd.n26 gnd 0.182952f
C2187 vdd.n27 gnd 20.858f
C2188 vdd.n28 gnd 7.85916f
C2189 vdd.n29 gnd 0.005437f
C2190 vdd.n30 gnd 0.005045f
C2191 vdd.n31 gnd 0.002791f
C2192 vdd.n32 gnd 0.006408f
C2193 vdd.n33 gnd 0.002711f
C2194 vdd.n34 gnd 0.002871f
C2195 vdd.n35 gnd 0.005045f
C2196 vdd.n36 gnd 0.002711f
C2197 vdd.n37 gnd 0.006408f
C2198 vdd.n38 gnd 0.002871f
C2199 vdd.n39 gnd 0.005045f
C2200 vdd.n40 gnd 0.002711f
C2201 vdd.n41 gnd 0.004806f
C2202 vdd.n42 gnd 0.00482f
C2203 vdd.t216 gnd 0.013767f
C2204 vdd.n43 gnd 0.030632f
C2205 vdd.n44 gnd 0.159414f
C2206 vdd.n45 gnd 0.002711f
C2207 vdd.n46 gnd 0.002871f
C2208 vdd.n47 gnd 0.006408f
C2209 vdd.n48 gnd 0.006408f
C2210 vdd.n49 gnd 0.002871f
C2211 vdd.n50 gnd 0.002711f
C2212 vdd.n51 gnd 0.005045f
C2213 vdd.n52 gnd 0.005045f
C2214 vdd.n53 gnd 0.002711f
C2215 vdd.n54 gnd 0.002871f
C2216 vdd.n55 gnd 0.006408f
C2217 vdd.n56 gnd 0.006408f
C2218 vdd.n57 gnd 0.002871f
C2219 vdd.n58 gnd 0.002711f
C2220 vdd.n59 gnd 0.005045f
C2221 vdd.n60 gnd 0.005045f
C2222 vdd.n61 gnd 0.002711f
C2223 vdd.n62 gnd 0.002871f
C2224 vdd.n63 gnd 0.006408f
C2225 vdd.n64 gnd 0.006408f
C2226 vdd.n65 gnd 0.01515f
C2227 vdd.n66 gnd 0.002791f
C2228 vdd.n67 gnd 0.002711f
C2229 vdd.n68 gnd 0.01304f
C2230 vdd.n69 gnd 0.009104f
C2231 vdd.t122 gnd 0.031895f
C2232 vdd.t226 gnd 0.031895f
C2233 vdd.n70 gnd 0.219206f
C2234 vdd.n71 gnd 0.172372f
C2235 vdd.t108 gnd 0.031895f
C2236 vdd.t218 gnd 0.031895f
C2237 vdd.n72 gnd 0.219206f
C2238 vdd.n73 gnd 0.139103f
C2239 vdd.t269 gnd 0.031895f
C2240 vdd.t248 gnd 0.031895f
C2241 vdd.n74 gnd 0.219206f
C2242 vdd.n75 gnd 0.139103f
C2243 vdd.t110 gnd 0.031895f
C2244 vdd.t251 gnd 0.031895f
C2245 vdd.n76 gnd 0.219206f
C2246 vdd.n77 gnd 0.139103f
C2247 vdd.t255 gnd 0.031895f
C2248 vdd.t126 gnd 0.031895f
C2249 vdd.n78 gnd 0.219206f
C2250 vdd.n79 gnd 0.139103f
C2251 vdd.t127 gnd 0.031895f
C2252 vdd.t263 gnd 0.031895f
C2253 vdd.n80 gnd 0.219206f
C2254 vdd.n81 gnd 0.139103f
C2255 vdd.t222 gnd 0.031895f
C2256 vdd.t112 gnd 0.031895f
C2257 vdd.n82 gnd 0.219206f
C2258 vdd.n83 gnd 0.139103f
C2259 vdd.n84 gnd 0.005437f
C2260 vdd.n85 gnd 0.005045f
C2261 vdd.n86 gnd 0.002791f
C2262 vdd.n87 gnd 0.006408f
C2263 vdd.n88 gnd 0.002711f
C2264 vdd.n89 gnd 0.002871f
C2265 vdd.n90 gnd 0.005045f
C2266 vdd.n91 gnd 0.002711f
C2267 vdd.n92 gnd 0.006408f
C2268 vdd.n93 gnd 0.002871f
C2269 vdd.n94 gnd 0.005045f
C2270 vdd.n95 gnd 0.002711f
C2271 vdd.n96 gnd 0.004806f
C2272 vdd.n97 gnd 0.00482f
C2273 vdd.t225 gnd 0.013767f
C2274 vdd.n98 gnd 0.030632f
C2275 vdd.n99 gnd 0.159414f
C2276 vdd.n100 gnd 0.002711f
C2277 vdd.n101 gnd 0.002871f
C2278 vdd.n102 gnd 0.006408f
C2279 vdd.n103 gnd 0.006408f
C2280 vdd.n104 gnd 0.002871f
C2281 vdd.n105 gnd 0.002711f
C2282 vdd.n106 gnd 0.005045f
C2283 vdd.n107 gnd 0.005045f
C2284 vdd.n108 gnd 0.002711f
C2285 vdd.n109 gnd 0.002871f
C2286 vdd.n110 gnd 0.006408f
C2287 vdd.n111 gnd 0.006408f
C2288 vdd.n112 gnd 0.002871f
C2289 vdd.n113 gnd 0.002711f
C2290 vdd.n114 gnd 0.005045f
C2291 vdd.n115 gnd 0.005045f
C2292 vdd.n116 gnd 0.002711f
C2293 vdd.n117 gnd 0.002871f
C2294 vdd.n118 gnd 0.006408f
C2295 vdd.n119 gnd 0.006408f
C2296 vdd.n120 gnd 0.01515f
C2297 vdd.n121 gnd 0.002791f
C2298 vdd.n122 gnd 0.002711f
C2299 vdd.n123 gnd 0.01304f
C2300 vdd.n124 gnd 0.008818f
C2301 vdd.n125 gnd 0.103493f
C2302 vdd.n126 gnd 0.005437f
C2303 vdd.n127 gnd 0.005045f
C2304 vdd.n128 gnd 0.002791f
C2305 vdd.n129 gnd 0.006408f
C2306 vdd.n130 gnd 0.002711f
C2307 vdd.n131 gnd 0.002871f
C2308 vdd.n132 gnd 0.005045f
C2309 vdd.n133 gnd 0.002711f
C2310 vdd.n134 gnd 0.006408f
C2311 vdd.n135 gnd 0.002871f
C2312 vdd.n136 gnd 0.005045f
C2313 vdd.n137 gnd 0.002711f
C2314 vdd.n138 gnd 0.004806f
C2315 vdd.n139 gnd 0.00482f
C2316 vdd.t227 gnd 0.013767f
C2317 vdd.n140 gnd 0.030632f
C2318 vdd.n141 gnd 0.159414f
C2319 vdd.n142 gnd 0.002711f
C2320 vdd.n143 gnd 0.002871f
C2321 vdd.n144 gnd 0.006408f
C2322 vdd.n145 gnd 0.006408f
C2323 vdd.n146 gnd 0.002871f
C2324 vdd.n147 gnd 0.002711f
C2325 vdd.n148 gnd 0.005045f
C2326 vdd.n149 gnd 0.005045f
C2327 vdd.n150 gnd 0.002711f
C2328 vdd.n151 gnd 0.002871f
C2329 vdd.n152 gnd 0.006408f
C2330 vdd.n153 gnd 0.006408f
C2331 vdd.n154 gnd 0.002871f
C2332 vdd.n155 gnd 0.002711f
C2333 vdd.n156 gnd 0.005045f
C2334 vdd.n157 gnd 0.005045f
C2335 vdd.n158 gnd 0.002711f
C2336 vdd.n159 gnd 0.002871f
C2337 vdd.n160 gnd 0.006408f
C2338 vdd.n161 gnd 0.006408f
C2339 vdd.n162 gnd 0.01515f
C2340 vdd.n163 gnd 0.002791f
C2341 vdd.n164 gnd 0.002711f
C2342 vdd.n165 gnd 0.01304f
C2343 vdd.n166 gnd 0.009104f
C2344 vdd.t264 gnd 0.031895f
C2345 vdd.t224 gnd 0.031895f
C2346 vdd.n167 gnd 0.219206f
C2347 vdd.n168 gnd 0.172372f
C2348 vdd.t256 gnd 0.031895f
C2349 vdd.t195 gnd 0.031895f
C2350 vdd.n169 gnd 0.219206f
C2351 vdd.n170 gnd 0.139103f
C2352 vdd.t194 gnd 0.031895f
C2353 vdd.t257 gnd 0.031895f
C2354 vdd.n171 gnd 0.219206f
C2355 vdd.n172 gnd 0.139103f
C2356 vdd.t244 gnd 0.031895f
C2357 vdd.t247 gnd 0.031895f
C2358 vdd.n173 gnd 0.219206f
C2359 vdd.n174 gnd 0.139103f
C2360 vdd.t9 gnd 0.031895f
C2361 vdd.t16 gnd 0.031895f
C2362 vdd.n175 gnd 0.219206f
C2363 vdd.n176 gnd 0.139103f
C2364 vdd.t206 gnd 0.031895f
C2365 vdd.t212 gnd 0.031895f
C2366 vdd.n177 gnd 0.219206f
C2367 vdd.n178 gnd 0.139103f
C2368 vdd.t20 gnd 0.031895f
C2369 vdd.t207 gnd 0.031895f
C2370 vdd.n179 gnd 0.219206f
C2371 vdd.n180 gnd 0.139103f
C2372 vdd.n181 gnd 0.005437f
C2373 vdd.n182 gnd 0.005045f
C2374 vdd.n183 gnd 0.002791f
C2375 vdd.n184 gnd 0.006408f
C2376 vdd.n185 gnd 0.002711f
C2377 vdd.n186 gnd 0.002871f
C2378 vdd.n187 gnd 0.005045f
C2379 vdd.n188 gnd 0.002711f
C2380 vdd.n189 gnd 0.006408f
C2381 vdd.n190 gnd 0.002871f
C2382 vdd.n191 gnd 0.005045f
C2383 vdd.n192 gnd 0.002711f
C2384 vdd.n193 gnd 0.004806f
C2385 vdd.n194 gnd 0.00482f
C2386 vdd.t211 gnd 0.013767f
C2387 vdd.n195 gnd 0.030632f
C2388 vdd.n196 gnd 0.159414f
C2389 vdd.n197 gnd 0.002711f
C2390 vdd.n198 gnd 0.002871f
C2391 vdd.n199 gnd 0.006408f
C2392 vdd.n200 gnd 0.006408f
C2393 vdd.n201 gnd 0.002871f
C2394 vdd.n202 gnd 0.002711f
C2395 vdd.n203 gnd 0.005045f
C2396 vdd.n204 gnd 0.005045f
C2397 vdd.n205 gnd 0.002711f
C2398 vdd.n206 gnd 0.002871f
C2399 vdd.n207 gnd 0.006408f
C2400 vdd.n208 gnd 0.006408f
C2401 vdd.n209 gnd 0.002871f
C2402 vdd.n210 gnd 0.002711f
C2403 vdd.n211 gnd 0.005045f
C2404 vdd.n212 gnd 0.005045f
C2405 vdd.n213 gnd 0.002711f
C2406 vdd.n214 gnd 0.002871f
C2407 vdd.n215 gnd 0.006408f
C2408 vdd.n216 gnd 0.006408f
C2409 vdd.n217 gnd 0.01515f
C2410 vdd.n218 gnd 0.002791f
C2411 vdd.n219 gnd 0.002711f
C2412 vdd.n220 gnd 0.01304f
C2413 vdd.n221 gnd 0.008818f
C2414 vdd.n222 gnd 0.061568f
C2415 vdd.n223 gnd 0.221846f
C2416 vdd.n224 gnd 0.005437f
C2417 vdd.n225 gnd 0.005045f
C2418 vdd.n226 gnd 0.002791f
C2419 vdd.n227 gnd 0.006408f
C2420 vdd.n228 gnd 0.002711f
C2421 vdd.n229 gnd 0.002871f
C2422 vdd.n230 gnd 0.005045f
C2423 vdd.n231 gnd 0.002711f
C2424 vdd.n232 gnd 0.006408f
C2425 vdd.n233 gnd 0.002871f
C2426 vdd.n234 gnd 0.005045f
C2427 vdd.n235 gnd 0.002711f
C2428 vdd.n236 gnd 0.004806f
C2429 vdd.n237 gnd 0.00482f
C2430 vdd.t267 gnd 0.013767f
C2431 vdd.n238 gnd 0.030632f
C2432 vdd.n239 gnd 0.159414f
C2433 vdd.n240 gnd 0.002711f
C2434 vdd.n241 gnd 0.002871f
C2435 vdd.n242 gnd 0.006408f
C2436 vdd.n243 gnd 0.006408f
C2437 vdd.n244 gnd 0.002871f
C2438 vdd.n245 gnd 0.002711f
C2439 vdd.n246 gnd 0.005045f
C2440 vdd.n247 gnd 0.005045f
C2441 vdd.n248 gnd 0.002711f
C2442 vdd.n249 gnd 0.002871f
C2443 vdd.n250 gnd 0.006408f
C2444 vdd.n251 gnd 0.006408f
C2445 vdd.n252 gnd 0.002871f
C2446 vdd.n253 gnd 0.002711f
C2447 vdd.n254 gnd 0.005045f
C2448 vdd.n255 gnd 0.005045f
C2449 vdd.n256 gnd 0.002711f
C2450 vdd.n257 gnd 0.002871f
C2451 vdd.n258 gnd 0.006408f
C2452 vdd.n259 gnd 0.006408f
C2453 vdd.n260 gnd 0.01515f
C2454 vdd.n261 gnd 0.002791f
C2455 vdd.n262 gnd 0.002711f
C2456 vdd.n263 gnd 0.01304f
C2457 vdd.n264 gnd 0.009104f
C2458 vdd.t209 gnd 0.031895f
C2459 vdd.t253 gnd 0.031895f
C2460 vdd.n265 gnd 0.219206f
C2461 vdd.n266 gnd 0.172372f
C2462 vdd.t202 gnd 0.031895f
C2463 vdd.t184 gnd 0.031895f
C2464 vdd.n267 gnd 0.219206f
C2465 vdd.n268 gnd 0.139103f
C2466 vdd.t182 gnd 0.031895f
C2467 vdd.t120 gnd 0.031895f
C2468 vdd.n269 gnd 0.219206f
C2469 vdd.n270 gnd 0.139103f
C2470 vdd.t259 gnd 0.031895f
C2471 vdd.t214 gnd 0.031895f
C2472 vdd.n271 gnd 0.219206f
C2473 vdd.n272 gnd 0.139103f
C2474 vdd.t116 gnd 0.031895f
C2475 vdd.t198 gnd 0.031895f
C2476 vdd.n273 gnd 0.219206f
C2477 vdd.n274 gnd 0.139103f
C2478 vdd.t125 gnd 0.031895f
C2479 vdd.t102 gnd 0.031895f
C2480 vdd.n275 gnd 0.219206f
C2481 vdd.n276 gnd 0.139103f
C2482 vdd.t268 gnd 0.031895f
C2483 vdd.t196 gnd 0.031895f
C2484 vdd.n277 gnd 0.219206f
C2485 vdd.n278 gnd 0.139103f
C2486 vdd.n279 gnd 0.005437f
C2487 vdd.n280 gnd 0.005045f
C2488 vdd.n281 gnd 0.002791f
C2489 vdd.n282 gnd 0.006408f
C2490 vdd.n283 gnd 0.002711f
C2491 vdd.n284 gnd 0.002871f
C2492 vdd.n285 gnd 0.005045f
C2493 vdd.n286 gnd 0.002711f
C2494 vdd.n287 gnd 0.006408f
C2495 vdd.n288 gnd 0.002871f
C2496 vdd.n289 gnd 0.005045f
C2497 vdd.n290 gnd 0.002711f
C2498 vdd.n291 gnd 0.004806f
C2499 vdd.n292 gnd 0.00482f
C2500 vdd.t246 gnd 0.013767f
C2501 vdd.n293 gnd 0.030632f
C2502 vdd.n294 gnd 0.159414f
C2503 vdd.n295 gnd 0.002711f
C2504 vdd.n296 gnd 0.002871f
C2505 vdd.n297 gnd 0.006408f
C2506 vdd.n298 gnd 0.006408f
C2507 vdd.n299 gnd 0.002871f
C2508 vdd.n300 gnd 0.002711f
C2509 vdd.n301 gnd 0.005045f
C2510 vdd.n302 gnd 0.005045f
C2511 vdd.n303 gnd 0.002711f
C2512 vdd.n304 gnd 0.002871f
C2513 vdd.n305 gnd 0.006408f
C2514 vdd.n306 gnd 0.006408f
C2515 vdd.n307 gnd 0.002871f
C2516 vdd.n308 gnd 0.002711f
C2517 vdd.n309 gnd 0.005045f
C2518 vdd.n310 gnd 0.005045f
C2519 vdd.n311 gnd 0.002711f
C2520 vdd.n312 gnd 0.002871f
C2521 vdd.n313 gnd 0.006408f
C2522 vdd.n314 gnd 0.006408f
C2523 vdd.n315 gnd 0.01515f
C2524 vdd.n316 gnd 0.002791f
C2525 vdd.n317 gnd 0.002711f
C2526 vdd.n318 gnd 0.01304f
C2527 vdd.n319 gnd 0.008818f
C2528 vdd.n320 gnd 0.061568f
C2529 vdd.n321 gnd 0.248438f
C2530 vdd.n322 gnd 0.007614f
C2531 vdd.n323 gnd 0.009907f
C2532 vdd.n324 gnd 0.007974f
C2533 vdd.n325 gnd 0.007974f
C2534 vdd.n326 gnd 0.009907f
C2535 vdd.n327 gnd 0.009907f
C2536 vdd.n328 gnd 0.723888f
C2537 vdd.n329 gnd 0.009907f
C2538 vdd.n330 gnd 0.009907f
C2539 vdd.n331 gnd 0.009907f
C2540 vdd.n332 gnd 0.784633f
C2541 vdd.n333 gnd 0.009907f
C2542 vdd.n334 gnd 0.009907f
C2543 vdd.n335 gnd 0.009907f
C2544 vdd.n336 gnd 0.009907f
C2545 vdd.n337 gnd 0.007974f
C2546 vdd.n338 gnd 0.009907f
C2547 vdd.t15 gnd 0.506215f
C2548 vdd.n339 gnd 0.009907f
C2549 vdd.n340 gnd 0.009907f
C2550 vdd.n341 gnd 0.009907f
C2551 vdd.t101 gnd 0.506215f
C2552 vdd.n342 gnd 0.009907f
C2553 vdd.n343 gnd 0.009907f
C2554 vdd.n344 gnd 0.009907f
C2555 vdd.n345 gnd 0.009907f
C2556 vdd.n346 gnd 0.009907f
C2557 vdd.n347 gnd 0.007974f
C2558 vdd.n348 gnd 0.009907f
C2559 vdd.n349 gnd 0.572023f
C2560 vdd.n350 gnd 0.009907f
C2561 vdd.n351 gnd 0.009907f
C2562 vdd.n352 gnd 0.009907f
C2563 vdd.t111 gnd 0.506215f
C2564 vdd.n353 gnd 0.009907f
C2565 vdd.n354 gnd 0.009907f
C2566 vdd.n355 gnd 0.009907f
C2567 vdd.n356 gnd 0.009907f
C2568 vdd.n357 gnd 0.009907f
C2569 vdd.n358 gnd 0.007974f
C2570 vdd.n359 gnd 0.009907f
C2571 vdd.t210 gnd 0.506215f
C2572 vdd.n360 gnd 0.009907f
C2573 vdd.n361 gnd 0.009907f
C2574 vdd.n362 gnd 0.009907f
C2575 vdd.n363 gnd 0.855503f
C2576 vdd.n364 gnd 0.009907f
C2577 vdd.n365 gnd 0.009907f
C2578 vdd.n366 gnd 0.009907f
C2579 vdd.n367 gnd 0.009907f
C2580 vdd.n368 gnd 0.009907f
C2581 vdd.n369 gnd 0.006618f
C2582 vdd.n370 gnd 0.02256f
C2583 vdd.t38 gnd 0.506215f
C2584 vdd.n371 gnd 0.009907f
C2585 vdd.n372 gnd 0.02256f
C2586 vdd.n404 gnd 0.009907f
C2587 vdd.t61 gnd 0.12188f
C2588 vdd.t60 gnd 0.130256f
C2589 vdd.t59 gnd 0.159174f
C2590 vdd.n405 gnd 0.204038f
C2591 vdd.n406 gnd 0.172226f
C2592 vdd.n407 gnd 0.013077f
C2593 vdd.n408 gnd 0.009907f
C2594 vdd.n409 gnd 0.007974f
C2595 vdd.n410 gnd 0.009907f
C2596 vdd.n411 gnd 0.007974f
C2597 vdd.n412 gnd 0.009907f
C2598 vdd.n413 gnd 0.007974f
C2599 vdd.n414 gnd 0.009907f
C2600 vdd.n415 gnd 0.007974f
C2601 vdd.n416 gnd 0.009907f
C2602 vdd.n417 gnd 0.007974f
C2603 vdd.n418 gnd 0.009907f
C2604 vdd.t40 gnd 0.12188f
C2605 vdd.t39 gnd 0.130256f
C2606 vdd.t37 gnd 0.159174f
C2607 vdd.n419 gnd 0.204038f
C2608 vdd.n420 gnd 0.172226f
C2609 vdd.n421 gnd 0.007974f
C2610 vdd.n422 gnd 0.009907f
C2611 vdd.n423 gnd 0.007974f
C2612 vdd.n424 gnd 0.009907f
C2613 vdd.n425 gnd 0.007974f
C2614 vdd.n426 gnd 0.009907f
C2615 vdd.n427 gnd 0.007974f
C2616 vdd.n428 gnd 0.009907f
C2617 vdd.n429 gnd 0.007974f
C2618 vdd.n430 gnd 0.009907f
C2619 vdd.t64 gnd 0.12188f
C2620 vdd.t63 gnd 0.130256f
C2621 vdd.t62 gnd 0.159174f
C2622 vdd.n431 gnd 0.204038f
C2623 vdd.n432 gnd 0.172226f
C2624 vdd.n433 gnd 0.017064f
C2625 vdd.n434 gnd 0.009907f
C2626 vdd.n435 gnd 0.007974f
C2627 vdd.n436 gnd 0.009907f
C2628 vdd.n437 gnd 0.007974f
C2629 vdd.n438 gnd 0.009907f
C2630 vdd.n439 gnd 0.007974f
C2631 vdd.n440 gnd 0.009907f
C2632 vdd.n441 gnd 0.007974f
C2633 vdd.n442 gnd 0.009907f
C2634 vdd.n443 gnd 0.02256f
C2635 vdd.n444 gnd 0.022714f
C2636 vdd.n445 gnd 0.022714f
C2637 vdd.n446 gnd 0.006618f
C2638 vdd.n447 gnd 0.007974f
C2639 vdd.n448 gnd 0.009907f
C2640 vdd.n449 gnd 0.009907f
C2641 vdd.n450 gnd 0.007974f
C2642 vdd.n451 gnd 0.009907f
C2643 vdd.n452 gnd 0.009907f
C2644 vdd.n453 gnd 0.009907f
C2645 vdd.n454 gnd 0.009907f
C2646 vdd.n455 gnd 0.009907f
C2647 vdd.n456 gnd 0.007974f
C2648 vdd.n457 gnd 0.007974f
C2649 vdd.n458 gnd 0.009907f
C2650 vdd.n459 gnd 0.009907f
C2651 vdd.n460 gnd 0.007974f
C2652 vdd.n461 gnd 0.009907f
C2653 vdd.n462 gnd 0.009907f
C2654 vdd.n463 gnd 0.009907f
C2655 vdd.n464 gnd 0.009907f
C2656 vdd.n465 gnd 0.009907f
C2657 vdd.n466 gnd 0.007974f
C2658 vdd.n467 gnd 0.007974f
C2659 vdd.n468 gnd 0.009907f
C2660 vdd.n469 gnd 0.009907f
C2661 vdd.n470 gnd 0.007974f
C2662 vdd.n471 gnd 0.009907f
C2663 vdd.n472 gnd 0.009907f
C2664 vdd.n473 gnd 0.009907f
C2665 vdd.n474 gnd 0.009907f
C2666 vdd.n475 gnd 0.009907f
C2667 vdd.n476 gnd 0.007974f
C2668 vdd.n477 gnd 0.007974f
C2669 vdd.n478 gnd 0.009907f
C2670 vdd.n479 gnd 0.009907f
C2671 vdd.n480 gnd 0.007974f
C2672 vdd.n481 gnd 0.009907f
C2673 vdd.n482 gnd 0.009907f
C2674 vdd.n483 gnd 0.009907f
C2675 vdd.n484 gnd 0.009907f
C2676 vdd.n485 gnd 0.009907f
C2677 vdd.n486 gnd 0.007974f
C2678 vdd.n487 gnd 0.007974f
C2679 vdd.n488 gnd 0.009907f
C2680 vdd.n489 gnd 0.009907f
C2681 vdd.n490 gnd 0.006658f
C2682 vdd.n491 gnd 0.009907f
C2683 vdd.n492 gnd 0.009907f
C2684 vdd.n493 gnd 0.009907f
C2685 vdd.n494 gnd 0.009907f
C2686 vdd.n495 gnd 0.009907f
C2687 vdd.n496 gnd 0.006658f
C2688 vdd.n497 gnd 0.007974f
C2689 vdd.n498 gnd 0.009907f
C2690 vdd.n499 gnd 0.009907f
C2691 vdd.n500 gnd 0.007974f
C2692 vdd.n501 gnd 0.009907f
C2693 vdd.n502 gnd 0.009907f
C2694 vdd.n503 gnd 0.009907f
C2695 vdd.n504 gnd 0.009907f
C2696 vdd.n505 gnd 0.009907f
C2697 vdd.n506 gnd 0.007974f
C2698 vdd.n507 gnd 0.007974f
C2699 vdd.n508 gnd 0.009907f
C2700 vdd.n509 gnd 0.009907f
C2701 vdd.n510 gnd 0.007974f
C2702 vdd.n511 gnd 0.009907f
C2703 vdd.n512 gnd 0.009907f
C2704 vdd.n513 gnd 0.009907f
C2705 vdd.n514 gnd 0.009907f
C2706 vdd.n515 gnd 0.009907f
C2707 vdd.n516 gnd 0.007974f
C2708 vdd.n517 gnd 0.007974f
C2709 vdd.n518 gnd 0.009907f
C2710 vdd.n519 gnd 0.009907f
C2711 vdd.n520 gnd 0.007974f
C2712 vdd.n521 gnd 0.009907f
C2713 vdd.n522 gnd 0.009907f
C2714 vdd.n523 gnd 0.009907f
C2715 vdd.n524 gnd 0.009907f
C2716 vdd.n525 gnd 0.009907f
C2717 vdd.n526 gnd 0.007974f
C2718 vdd.n527 gnd 0.007974f
C2719 vdd.n528 gnd 0.009907f
C2720 vdd.n529 gnd 0.009907f
C2721 vdd.n530 gnd 0.007974f
C2722 vdd.n531 gnd 0.009907f
C2723 vdd.n532 gnd 0.009907f
C2724 vdd.n533 gnd 0.009907f
C2725 vdd.n534 gnd 0.009907f
C2726 vdd.n535 gnd 0.009907f
C2727 vdd.n536 gnd 0.007974f
C2728 vdd.n537 gnd 0.007974f
C2729 vdd.n538 gnd 0.009907f
C2730 vdd.n539 gnd 0.009907f
C2731 vdd.n540 gnd 0.007974f
C2732 vdd.n541 gnd 0.009907f
C2733 vdd.n542 gnd 0.009907f
C2734 vdd.n543 gnd 0.009907f
C2735 vdd.n544 gnd 0.009907f
C2736 vdd.n545 gnd 0.009907f
C2737 vdd.n546 gnd 0.005422f
C2738 vdd.n547 gnd 0.017064f
C2739 vdd.n548 gnd 0.009907f
C2740 vdd.n549 gnd 0.009907f
C2741 vdd.n550 gnd 0.007894f
C2742 vdd.n551 gnd 0.009907f
C2743 vdd.n552 gnd 0.009907f
C2744 vdd.n553 gnd 0.009907f
C2745 vdd.n554 gnd 0.009907f
C2746 vdd.n555 gnd 0.009907f
C2747 vdd.n556 gnd 0.007974f
C2748 vdd.n557 gnd 0.007974f
C2749 vdd.n558 gnd 0.009907f
C2750 vdd.n559 gnd 0.009907f
C2751 vdd.n560 gnd 0.007974f
C2752 vdd.n561 gnd 0.009907f
C2753 vdd.n562 gnd 0.009907f
C2754 vdd.n563 gnd 0.009907f
C2755 vdd.n564 gnd 0.009907f
C2756 vdd.n565 gnd 0.009907f
C2757 vdd.n566 gnd 0.007974f
C2758 vdd.n567 gnd 0.007974f
C2759 vdd.n568 gnd 0.009907f
C2760 vdd.n569 gnd 0.009907f
C2761 vdd.n570 gnd 0.007974f
C2762 vdd.n571 gnd 0.009907f
C2763 vdd.n572 gnd 0.009907f
C2764 vdd.n573 gnd 0.009907f
C2765 vdd.n574 gnd 0.009907f
C2766 vdd.n575 gnd 0.009907f
C2767 vdd.n576 gnd 0.007974f
C2768 vdd.n577 gnd 0.007974f
C2769 vdd.n578 gnd 0.009907f
C2770 vdd.n579 gnd 0.009907f
C2771 vdd.n580 gnd 0.007974f
C2772 vdd.n581 gnd 0.009907f
C2773 vdd.n582 gnd 0.009907f
C2774 vdd.n583 gnd 0.009907f
C2775 vdd.n584 gnd 0.009907f
C2776 vdd.n585 gnd 0.009907f
C2777 vdd.n586 gnd 0.007974f
C2778 vdd.n587 gnd 0.007974f
C2779 vdd.n588 gnd 0.009907f
C2780 vdd.n589 gnd 0.009907f
C2781 vdd.n590 gnd 0.007974f
C2782 vdd.n591 gnd 0.009907f
C2783 vdd.n592 gnd 0.009907f
C2784 vdd.n593 gnd 0.009907f
C2785 vdd.n594 gnd 0.009907f
C2786 vdd.n595 gnd 0.009907f
C2787 vdd.n596 gnd 0.007974f
C2788 vdd.n597 gnd 0.009907f
C2789 vdd.n598 gnd 0.007974f
C2790 vdd.n599 gnd 0.004186f
C2791 vdd.n600 gnd 0.009907f
C2792 vdd.n601 gnd 0.009907f
C2793 vdd.n602 gnd 0.007974f
C2794 vdd.n603 gnd 0.009907f
C2795 vdd.n604 gnd 0.007974f
C2796 vdd.n605 gnd 0.009907f
C2797 vdd.n606 gnd 0.007974f
C2798 vdd.n607 gnd 0.009907f
C2799 vdd.n608 gnd 0.007974f
C2800 vdd.n609 gnd 0.009907f
C2801 vdd.n610 gnd 0.007974f
C2802 vdd.n611 gnd 0.009907f
C2803 vdd.n612 gnd 0.009907f
C2804 vdd.n613 gnd 0.551774f
C2805 vdd.t109 gnd 0.506215f
C2806 vdd.n614 gnd 0.009907f
C2807 vdd.n615 gnd 0.007974f
C2808 vdd.n616 gnd 0.009907f
C2809 vdd.n617 gnd 0.007974f
C2810 vdd.n618 gnd 0.009907f
C2811 vdd.t181 gnd 0.506215f
C2812 vdd.n619 gnd 0.009907f
C2813 vdd.n620 gnd 0.007974f
C2814 vdd.n621 gnd 0.009907f
C2815 vdd.n622 gnd 0.007974f
C2816 vdd.n623 gnd 0.009907f
C2817 vdd.t183 gnd 0.506215f
C2818 vdd.n624 gnd 0.632769f
C2819 vdd.n625 gnd 0.009907f
C2820 vdd.n626 gnd 0.007974f
C2821 vdd.n627 gnd 0.009907f
C2822 vdd.n628 gnd 0.007974f
C2823 vdd.n629 gnd 0.009907f
C2824 vdd.t107 gnd 0.506215f
C2825 vdd.n630 gnd 0.009907f
C2826 vdd.n631 gnd 0.007974f
C2827 vdd.n632 gnd 0.009907f
C2828 vdd.n633 gnd 0.007974f
C2829 vdd.n634 gnd 0.009907f
C2830 vdd.n635 gnd 0.703639f
C2831 vdd.n636 gnd 0.840317f
C2832 vdd.t223 gnd 0.506215f
C2833 vdd.n637 gnd 0.009907f
C2834 vdd.n638 gnd 0.007974f
C2835 vdd.n639 gnd 0.009907f
C2836 vdd.n640 gnd 0.007974f
C2837 vdd.n641 gnd 0.009907f
C2838 vdd.n642 gnd 0.531526f
C2839 vdd.n643 gnd 0.009907f
C2840 vdd.n644 gnd 0.007974f
C2841 vdd.n645 gnd 0.009907f
C2842 vdd.n646 gnd 0.007974f
C2843 vdd.n647 gnd 0.009907f
C2844 vdd.n648 gnd 1.01243f
C2845 vdd.t215 gnd 0.506215f
C2846 vdd.n649 gnd 0.009907f
C2847 vdd.n650 gnd 0.007974f
C2848 vdd.n651 gnd 0.009907f
C2849 vdd.n652 gnd 0.007974f
C2850 vdd.n653 gnd 0.009907f
C2851 vdd.t26 gnd 0.506215f
C2852 vdd.n654 gnd 0.009907f
C2853 vdd.n655 gnd 0.007974f
C2854 vdd.n656 gnd 0.022714f
C2855 vdd.n657 gnd 0.022714f
C2856 vdd.n658 gnd 10.5191f
C2857 vdd.n659 gnd 0.561899f
C2858 vdd.n660 gnd 0.022714f
C2859 vdd.n661 gnd 0.00852f
C2860 vdd.n662 gnd 0.007974f
C2861 vdd.n667 gnd 0.00634f
C2862 vdd.n668 gnd 0.007974f
C2863 vdd.n669 gnd 0.009907f
C2864 vdd.n670 gnd 0.009907f
C2865 vdd.n671 gnd 0.009907f
C2866 vdd.n672 gnd 0.009907f
C2867 vdd.n673 gnd 0.009907f
C2868 vdd.n674 gnd 0.007974f
C2869 vdd.n675 gnd 0.009907f
C2870 vdd.n676 gnd 0.009907f
C2871 vdd.n677 gnd 0.009907f
C2872 vdd.n678 gnd 0.009907f
C2873 vdd.n679 gnd 0.009907f
C2874 vdd.n680 gnd 0.007974f
C2875 vdd.n681 gnd 0.009907f
C2876 vdd.n682 gnd 0.009907f
C2877 vdd.n683 gnd 0.009907f
C2878 vdd.n684 gnd 0.009907f
C2879 vdd.n685 gnd 0.009907f
C2880 vdd.t42 gnd 0.12188f
C2881 vdd.t43 gnd 0.130256f
C2882 vdd.t41 gnd 0.159174f
C2883 vdd.n686 gnd 0.204038f
C2884 vdd.n687 gnd 0.171429f
C2885 vdd.n688 gnd 0.016267f
C2886 vdd.n689 gnd 0.009907f
C2887 vdd.n690 gnd 0.009907f
C2888 vdd.n691 gnd 0.009907f
C2889 vdd.n692 gnd 0.009907f
C2890 vdd.n693 gnd 0.009907f
C2891 vdd.n694 gnd 0.007974f
C2892 vdd.n695 gnd 0.009907f
C2893 vdd.n696 gnd 0.009907f
C2894 vdd.n697 gnd 0.009907f
C2895 vdd.n698 gnd 0.009907f
C2896 vdd.n699 gnd 0.009907f
C2897 vdd.n700 gnd 0.007974f
C2898 vdd.n701 gnd 0.009907f
C2899 vdd.n702 gnd 0.009907f
C2900 vdd.n703 gnd 0.009907f
C2901 vdd.n704 gnd 0.009907f
C2902 vdd.n705 gnd 0.009907f
C2903 vdd.n706 gnd 0.007974f
C2904 vdd.n707 gnd 0.009907f
C2905 vdd.n708 gnd 0.009907f
C2906 vdd.n709 gnd 0.009907f
C2907 vdd.n710 gnd 0.009907f
C2908 vdd.n711 gnd 0.009907f
C2909 vdd.n712 gnd 0.007974f
C2910 vdd.n713 gnd 0.009907f
C2911 vdd.n714 gnd 0.009907f
C2912 vdd.n715 gnd 0.009907f
C2913 vdd.n716 gnd 0.009907f
C2914 vdd.n717 gnd 0.009907f
C2915 vdd.n718 gnd 0.007974f
C2916 vdd.n719 gnd 0.009907f
C2917 vdd.n720 gnd 0.009907f
C2918 vdd.n721 gnd 0.009907f
C2919 vdd.n722 gnd 0.007894f
C2920 vdd.t27 gnd 0.12188f
C2921 vdd.t28 gnd 0.130256f
C2922 vdd.t25 gnd 0.159174f
C2923 vdd.n723 gnd 0.204038f
C2924 vdd.n724 gnd 0.171429f
C2925 vdd.n725 gnd 0.009907f
C2926 vdd.n726 gnd 0.007974f
C2927 vdd.n728 gnd 0.009907f
C2928 vdd.n730 gnd 0.009907f
C2929 vdd.n731 gnd 0.009907f
C2930 vdd.n732 gnd 0.007974f
C2931 vdd.n733 gnd 0.009907f
C2932 vdd.n734 gnd 0.009907f
C2933 vdd.n735 gnd 0.009907f
C2934 vdd.n736 gnd 0.009907f
C2935 vdd.n737 gnd 0.009907f
C2936 vdd.n738 gnd 0.007974f
C2937 vdd.n739 gnd 0.009907f
C2938 vdd.n740 gnd 0.009907f
C2939 vdd.n741 gnd 0.009907f
C2940 vdd.n742 gnd 0.009907f
C2941 vdd.n743 gnd 0.009907f
C2942 vdd.n744 gnd 0.007974f
C2943 vdd.n745 gnd 0.009907f
C2944 vdd.n746 gnd 0.009907f
C2945 vdd.n747 gnd 0.009907f
C2946 vdd.n748 gnd 0.00634f
C2947 vdd.n753 gnd 0.006737f
C2948 vdd.n754 gnd 0.006737f
C2949 vdd.n755 gnd 0.006737f
C2950 vdd.n756 gnd 10.2964f
C2951 vdd.n757 gnd 0.006737f
C2952 vdd.n758 gnd 0.006737f
C2953 vdd.n759 gnd 0.006737f
C2954 vdd.n761 gnd 0.006737f
C2955 vdd.n762 gnd 0.006737f
C2956 vdd.n764 gnd 0.006737f
C2957 vdd.n765 gnd 0.004904f
C2958 vdd.n767 gnd 0.006737f
C2959 vdd.t32 gnd 0.272227f
C2960 vdd.t31 gnd 0.278658f
C2961 vdd.t29 gnd 0.17772f
C2962 vdd.n768 gnd 0.096048f
C2963 vdd.n769 gnd 0.054481f
C2964 vdd.n770 gnd 0.009628f
C2965 vdd.n771 gnd 0.015444f
C2966 vdd.n773 gnd 0.006737f
C2967 vdd.n774 gnd 0.688453f
C2968 vdd.n775 gnd 0.01459f
C2969 vdd.n776 gnd 0.01459f
C2970 vdd.n777 gnd 0.006737f
C2971 vdd.n778 gnd 0.015527f
C2972 vdd.n779 gnd 0.006737f
C2973 vdd.n780 gnd 0.006737f
C2974 vdd.n781 gnd 0.006737f
C2975 vdd.n782 gnd 0.006737f
C2976 vdd.n783 gnd 0.006737f
C2977 vdd.n785 gnd 0.006737f
C2978 vdd.n786 gnd 0.006737f
C2979 vdd.n788 gnd 0.006737f
C2980 vdd.n789 gnd 0.006737f
C2981 vdd.n791 gnd 0.006737f
C2982 vdd.n792 gnd 0.006737f
C2983 vdd.n794 gnd 0.006737f
C2984 vdd.n795 gnd 0.006737f
C2985 vdd.n797 gnd 0.006737f
C2986 vdd.n798 gnd 0.006737f
C2987 vdd.n800 gnd 0.006737f
C2988 vdd.n801 gnd 0.004904f
C2989 vdd.n803 gnd 0.006737f
C2990 vdd.t67 gnd 0.272227f
C2991 vdd.t66 gnd 0.278658f
C2992 vdd.t65 gnd 0.17772f
C2993 vdd.n804 gnd 0.096048f
C2994 vdd.n805 gnd 0.054481f
C2995 vdd.n806 gnd 0.009628f
C2996 vdd.n807 gnd 0.006737f
C2997 vdd.n808 gnd 0.006737f
C2998 vdd.t30 gnd 0.344226f
C2999 vdd.n809 gnd 0.006737f
C3000 vdd.n810 gnd 0.006737f
C3001 vdd.n811 gnd 0.006737f
C3002 vdd.n812 gnd 0.006737f
C3003 vdd.n813 gnd 0.006737f
C3004 vdd.n814 gnd 0.688453f
C3005 vdd.n815 gnd 0.006737f
C3006 vdd.n816 gnd 0.006737f
C3007 vdd.n817 gnd 0.561899f
C3008 vdd.n818 gnd 0.006737f
C3009 vdd.n819 gnd 0.006737f
C3010 vdd.n820 gnd 0.006737f
C3011 vdd.n821 gnd 0.006737f
C3012 vdd.n822 gnd 0.688453f
C3013 vdd.n823 gnd 0.006737f
C3014 vdd.n824 gnd 0.006737f
C3015 vdd.n825 gnd 0.006737f
C3016 vdd.n826 gnd 0.006737f
C3017 vdd.n827 gnd 0.006737f
C3018 vdd.t157 gnd 0.344226f
C3019 vdd.n828 gnd 0.006737f
C3020 vdd.n829 gnd 0.006737f
C3021 vdd.n830 gnd 0.006737f
C3022 vdd.n831 gnd 0.006737f
C3023 vdd.n832 gnd 0.006737f
C3024 vdd.t163 gnd 0.344226f
C3025 vdd.n833 gnd 0.006737f
C3026 vdd.n834 gnd 0.006737f
C3027 vdd.n835 gnd 0.68339f
C3028 vdd.n836 gnd 0.006737f
C3029 vdd.n837 gnd 0.006737f
C3030 vdd.n838 gnd 0.006737f
C3031 vdd.t166 gnd 0.344226f
C3032 vdd.n839 gnd 0.006737f
C3033 vdd.n840 gnd 0.006737f
C3034 vdd.n841 gnd 0.531526f
C3035 vdd.n842 gnd 0.006737f
C3036 vdd.n843 gnd 0.006737f
C3037 vdd.n844 gnd 0.006737f
C3038 vdd.n845 gnd 0.460656f
C3039 vdd.n846 gnd 0.006737f
C3040 vdd.n847 gnd 0.006737f
C3041 vdd.n848 gnd 0.379661f
C3042 vdd.n849 gnd 0.006737f
C3043 vdd.n850 gnd 0.006737f
C3044 vdd.n851 gnd 0.006737f
C3045 vdd.n852 gnd 0.566961f
C3046 vdd.n853 gnd 0.006737f
C3047 vdd.n854 gnd 0.006737f
C3048 vdd.t136 gnd 0.344226f
C3049 vdd.n855 gnd 0.006737f
C3050 vdd.t46 gnd 0.278658f
C3051 vdd.t44 gnd 0.17772f
C3052 vdd.t47 gnd 0.278658f
C3053 vdd.n856 gnd 0.156617f
C3054 vdd.n857 gnd 0.006737f
C3055 vdd.n858 gnd 0.006737f
C3056 vdd.n859 gnd 0.688453f
C3057 vdd.n860 gnd 0.006737f
C3058 vdd.n861 gnd 0.006737f
C3059 vdd.t45 gnd 0.268294f
C3060 vdd.t138 gnd 0.121492f
C3061 vdd.n862 gnd 0.006737f
C3062 vdd.n863 gnd 0.006737f
C3063 vdd.n864 gnd 0.006737f
C3064 vdd.t149 gnd 0.344226f
C3065 vdd.n865 gnd 0.006737f
C3066 vdd.n866 gnd 0.006737f
C3067 vdd.n867 gnd 0.006737f
C3068 vdd.n868 gnd 0.006737f
C3069 vdd.n869 gnd 0.006737f
C3070 vdd.t167 gnd 0.344226f
C3071 vdd.n870 gnd 0.006737f
C3072 vdd.n871 gnd 0.006737f
C3073 vdd.n872 gnd 0.61252f
C3074 vdd.n873 gnd 0.006737f
C3075 vdd.n874 gnd 0.006737f
C3076 vdd.n875 gnd 0.006737f
C3077 vdd.n876 gnd 0.379661f
C3078 vdd.n877 gnd 0.006737f
C3079 vdd.n878 gnd 0.006737f
C3080 vdd.t145 gnd 0.344226f
C3081 vdd.n879 gnd 0.006737f
C3082 vdd.n880 gnd 0.006737f
C3083 vdd.n881 gnd 0.006737f
C3084 vdd.n882 gnd 0.531526f
C3085 vdd.n883 gnd 0.006737f
C3086 vdd.n884 gnd 0.006737f
C3087 vdd.t129 gnd 0.253108f
C3088 vdd.t179 gnd 0.308791f
C3089 vdd.n885 gnd 0.006737f
C3090 vdd.n886 gnd 0.006737f
C3091 vdd.n887 gnd 0.006737f
C3092 vdd.t171 gnd 0.344226f
C3093 vdd.n888 gnd 0.006737f
C3094 vdd.n889 gnd 0.006737f
C3095 vdd.t168 gnd 0.344226f
C3096 vdd.n890 gnd 0.006737f
C3097 vdd.n891 gnd 0.006737f
C3098 vdd.n892 gnd 0.006737f
C3099 vdd.t153 gnd 0.344226f
C3100 vdd.n893 gnd 0.006737f
C3101 vdd.n894 gnd 0.006737f
C3102 vdd.t133 gnd 0.344226f
C3103 vdd.n895 gnd 0.006737f
C3104 vdd.n896 gnd 0.006737f
C3105 vdd.n897 gnd 0.006737f
C3106 vdd.n898 gnd 0.688453f
C3107 vdd.n899 gnd 0.006737f
C3108 vdd.n900 gnd 0.006737f
C3109 vdd.n901 gnd 0.475842f
C3110 vdd.n902 gnd 0.006737f
C3111 vdd.n903 gnd 0.006737f
C3112 vdd.n904 gnd 0.006737f
C3113 vdd.t134 gnd 0.344226f
C3114 vdd.n905 gnd 0.006737f
C3115 vdd.n906 gnd 0.006737f
C3116 vdd.n907 gnd 0.006737f
C3117 vdd.n908 gnd 0.006737f
C3118 vdd.n909 gnd 0.006737f
C3119 vdd.t161 gnd 0.344226f
C3120 vdd.n910 gnd 0.006737f
C3121 vdd.n911 gnd 0.006737f
C3122 vdd.t76 gnd 0.344226f
C3123 vdd.n912 gnd 0.006737f
C3124 vdd.n913 gnd 0.015527f
C3125 vdd.n914 gnd 0.015527f
C3126 vdd.t159 gnd 0.607458f
C3127 vdd.n915 gnd 0.01459f
C3128 vdd.n916 gnd 0.01459f
C3129 vdd.n917 gnd 0.384723f
C3130 vdd.n918 gnd 0.015527f
C3131 vdd.n919 gnd 0.006737f
C3132 vdd.n920 gnd 0.006737f
C3133 vdd.t175 gnd 0.607458f
C3134 vdd.n938 gnd 0.015527f
C3135 vdd.n956 gnd 0.01459f
C3136 vdd.n957 gnd 0.006737f
C3137 vdd.n958 gnd 0.01459f
C3138 vdd.t97 gnd 0.272227f
C3139 vdd.t96 gnd 0.278658f
C3140 vdd.t95 gnd 0.17772f
C3141 vdd.n959 gnd 0.096048f
C3142 vdd.n960 gnd 0.054481f
C3143 vdd.n961 gnd 0.015444f
C3144 vdd.n962 gnd 0.006737f
C3145 vdd.n963 gnd 0.384723f
C3146 vdd.n964 gnd 0.01459f
C3147 vdd.n965 gnd 0.006737f
C3148 vdd.n966 gnd 0.015527f
C3149 vdd.n967 gnd 0.006737f
C3150 vdd.t74 gnd 0.272227f
C3151 vdd.t73 gnd 0.278658f
C3152 vdd.t71 gnd 0.17772f
C3153 vdd.n968 gnd 0.096048f
C3154 vdd.n969 gnd 0.054481f
C3155 vdd.n970 gnd 0.009628f
C3156 vdd.n971 gnd 0.006737f
C3157 vdd.n972 gnd 0.006737f
C3158 vdd.t72 gnd 0.344226f
C3159 vdd.n973 gnd 0.006737f
C3160 vdd.t173 gnd 0.344226f
C3161 vdd.n974 gnd 0.006737f
C3162 vdd.n975 gnd 0.006737f
C3163 vdd.n976 gnd 0.006737f
C3164 vdd.n977 gnd 0.006737f
C3165 vdd.n978 gnd 0.006737f
C3166 vdd.n979 gnd 0.688453f
C3167 vdd.n980 gnd 0.006737f
C3168 vdd.n981 gnd 0.006737f
C3169 vdd.t147 gnd 0.344226f
C3170 vdd.n982 gnd 0.006737f
C3171 vdd.n983 gnd 0.006737f
C3172 vdd.n984 gnd 0.006737f
C3173 vdd.n985 gnd 0.006737f
C3174 vdd.n986 gnd 0.475842f
C3175 vdd.n987 gnd 0.006737f
C3176 vdd.n988 gnd 0.006737f
C3177 vdd.n989 gnd 0.006737f
C3178 vdd.n990 gnd 0.006737f
C3179 vdd.n991 gnd 0.006737f
C3180 vdd.t130 gnd 0.344226f
C3181 vdd.n992 gnd 0.006737f
C3182 vdd.n993 gnd 0.006737f
C3183 vdd.t164 gnd 0.344226f
C3184 vdd.n994 gnd 0.006737f
C3185 vdd.n995 gnd 0.006737f
C3186 vdd.n996 gnd 0.006737f
C3187 vdd.t152 gnd 0.344226f
C3188 vdd.n997 gnd 0.006737f
C3189 vdd.n998 gnd 0.006737f
C3190 vdd.t131 gnd 0.344226f
C3191 vdd.n999 gnd 0.006737f
C3192 vdd.n1000 gnd 0.006737f
C3193 vdd.n1001 gnd 0.006737f
C3194 vdd.t150 gnd 0.308791f
C3195 vdd.n1002 gnd 0.006737f
C3196 vdd.n1003 gnd 0.006737f
C3197 vdd.n1004 gnd 0.531526f
C3198 vdd.n1005 gnd 0.006737f
C3199 vdd.n1006 gnd 0.006737f
C3200 vdd.n1007 gnd 0.006737f
C3201 vdd.t169 gnd 0.344226f
C3202 vdd.n1008 gnd 0.006737f
C3203 vdd.n1009 gnd 0.006737f
C3204 vdd.t139 gnd 0.253108f
C3205 vdd.n1010 gnd 0.379661f
C3206 vdd.n1011 gnd 0.006737f
C3207 vdd.n1012 gnd 0.006737f
C3208 vdd.n1013 gnd 0.006737f
C3209 vdd.n1014 gnd 0.61252f
C3210 vdd.n1015 gnd 0.006737f
C3211 vdd.n1016 gnd 0.006737f
C3212 vdd.t177 gnd 0.344226f
C3213 vdd.n1017 gnd 0.006737f
C3214 vdd.n1018 gnd 0.006737f
C3215 vdd.n1019 gnd 0.006737f
C3216 vdd.n1020 gnd 0.688453f
C3217 vdd.n1021 gnd 0.006737f
C3218 vdd.n1022 gnd 0.006737f
C3219 vdd.t144 gnd 0.344226f
C3220 vdd.n1023 gnd 0.006737f
C3221 vdd.n1024 gnd 0.006737f
C3222 vdd.n1025 gnd 0.006737f
C3223 vdd.t137 gnd 0.121492f
C3224 vdd.n1026 gnd 0.006737f
C3225 vdd.n1027 gnd 0.006737f
C3226 vdd.n1028 gnd 0.006737f
C3227 vdd.t87 gnd 0.278658f
C3228 vdd.t85 gnd 0.17772f
C3229 vdd.t88 gnd 0.278658f
C3230 vdd.n1029 gnd 0.156617f
C3231 vdd.n1030 gnd 0.006737f
C3232 vdd.n1031 gnd 0.006737f
C3233 vdd.t158 gnd 0.344226f
C3234 vdd.n1032 gnd 0.006737f
C3235 vdd.n1033 gnd 0.006737f
C3236 vdd.t86 gnd 0.268294f
C3237 vdd.n1034 gnd 0.566961f
C3238 vdd.n1035 gnd 0.006737f
C3239 vdd.n1036 gnd 0.006737f
C3240 vdd.n1037 gnd 0.006737f
C3241 vdd.n1038 gnd 0.379661f
C3242 vdd.n1039 gnd 0.006737f
C3243 vdd.n1040 gnd 0.006737f
C3244 vdd.n1041 gnd 0.460656f
C3245 vdd.n1042 gnd 0.006737f
C3246 vdd.n1043 gnd 0.006737f
C3247 vdd.n1044 gnd 0.006737f
C3248 vdd.n1045 gnd 0.531526f
C3249 vdd.n1046 gnd 0.006737f
C3250 vdd.n1047 gnd 0.006737f
C3251 vdd.t141 gnd 0.344226f
C3252 vdd.n1048 gnd 0.006737f
C3253 vdd.n1049 gnd 0.006737f
C3254 vdd.n1050 gnd 0.006737f
C3255 vdd.n1051 gnd 0.68339f
C3256 vdd.n1052 gnd 0.006737f
C3257 vdd.n1053 gnd 0.006737f
C3258 vdd.t140 gnd 0.344226f
C3259 vdd.n1054 gnd 0.006737f
C3260 vdd.n1055 gnd 0.006737f
C3261 vdd.n1056 gnd 0.006737f
C3262 vdd.n1057 gnd 0.688453f
C3263 vdd.n1058 gnd 0.006737f
C3264 vdd.n1059 gnd 0.006737f
C3265 vdd.t178 gnd 0.344226f
C3266 vdd.n1060 gnd 0.006737f
C3267 vdd.n1061 gnd 0.006737f
C3268 vdd.n1062 gnd 0.006737f
C3269 vdd.n1063 gnd 0.688453f
C3270 vdd.n1064 gnd 0.006737f
C3271 vdd.n1065 gnd 0.006737f
C3272 vdd.n1066 gnd 0.006737f
C3273 vdd.n1067 gnd 0.006737f
C3274 vdd.n1068 gnd 0.006737f
C3275 vdd.n1069 gnd 0.561899f
C3276 vdd.n1070 gnd 0.006737f
C3277 vdd.n1071 gnd 0.006737f
C3278 vdd.n1072 gnd 0.006737f
C3279 vdd.n1073 gnd 0.006737f
C3280 vdd.n1074 gnd 0.006737f
C3281 vdd.n1075 gnd 0.688453f
C3282 vdd.n1076 gnd 0.006737f
C3283 vdd.n1077 gnd 0.006737f
C3284 vdd.t34 gnd 0.344226f
C3285 vdd.n1078 gnd 0.006737f
C3286 vdd.n1079 gnd 0.015527f
C3287 vdd.n1080 gnd 0.015527f
C3288 vdd.n1081 gnd 10.2964f
C3289 vdd.n1082 gnd 0.01459f
C3290 vdd.n1083 gnd 0.01459f
C3291 vdd.n1084 gnd 0.015527f
C3292 vdd.n1085 gnd 0.006737f
C3293 vdd.n1087 gnd 0.006737f
C3294 vdd.n1088 gnd 0.006737f
C3295 vdd.n1089 gnd 0.006737f
C3296 vdd.n1090 gnd 0.006737f
C3297 vdd.n1091 gnd 0.006737f
C3298 vdd.n1092 gnd 0.006737f
C3299 vdd.n1093 gnd 0.035445f
C3300 vdd.n1094 gnd 0.006737f
C3301 vdd.n1095 gnd 0.006737f
C3302 vdd.n1096 gnd 0.006737f
C3303 vdd.n1097 gnd 0.006737f
C3304 vdd.n1098 gnd 0.006737f
C3305 vdd.n1099 gnd 0.006737f
C3306 vdd.n1100 gnd 0.006737f
C3307 vdd.t99 gnd 0.272227f
C3308 vdd.t100 gnd 0.278658f
C3309 vdd.t98 gnd 0.17772f
C3310 vdd.n1101 gnd 0.096048f
C3311 vdd.n1102 gnd 0.054481f
C3312 vdd.n1103 gnd 0.006737f
C3313 vdd.n1104 gnd 0.006737f
C3314 vdd.n1105 gnd 0.006737f
C3315 vdd.n1106 gnd 0.006737f
C3316 vdd.t35 gnd 0.272227f
C3317 vdd.t36 gnd 0.278658f
C3318 vdd.t33 gnd 0.17772f
C3319 vdd.n1107 gnd 0.096048f
C3320 vdd.n1108 gnd 0.054481f
C3321 vdd.n1109 gnd 0.006737f
C3322 vdd.n1110 gnd 0.006737f
C3323 vdd.n1111 gnd 0.006737f
C3324 vdd.n1112 gnd 0.006737f
C3325 vdd.n1113 gnd 0.006737f
C3326 vdd.n1114 gnd 0.006737f
C3327 vdd.n1115 gnd 0.00634f
C3328 vdd.n1118 gnd 0.022714f
C3329 vdd.n1119 gnd 0.007974f
C3330 vdd.n1120 gnd 0.009907f
C3331 vdd.n1122 gnd 0.009907f
C3332 vdd.n1123 gnd 0.006618f
C3333 vdd.n1124 gnd 0.561899f
C3334 vdd.n1125 gnd 10.5191f
C3335 vdd.n1126 gnd 0.009907f
C3336 vdd.n1127 gnd 0.022714f
C3337 vdd.n1128 gnd 0.007974f
C3338 vdd.n1129 gnd 0.009907f
C3339 vdd.n1130 gnd 0.007974f
C3340 vdd.n1131 gnd 0.009907f
C3341 vdd.n1132 gnd 1.01243f
C3342 vdd.n1133 gnd 0.009907f
C3343 vdd.n1134 gnd 0.007974f
C3344 vdd.n1135 gnd 0.007974f
C3345 vdd.n1136 gnd 0.009907f
C3346 vdd.n1137 gnd 0.007974f
C3347 vdd.n1138 gnd 0.009907f
C3348 vdd.t234 gnd 0.506215f
C3349 vdd.n1139 gnd 0.009907f
C3350 vdd.n1140 gnd 0.007974f
C3351 vdd.n1141 gnd 0.009907f
C3352 vdd.n1142 gnd 0.007974f
C3353 vdd.n1143 gnd 0.009907f
C3354 vdd.t103 gnd 0.506215f
C3355 vdd.n1144 gnd 0.009907f
C3356 vdd.n1145 gnd 0.007974f
C3357 vdd.n1146 gnd 0.009907f
C3358 vdd.n1147 gnd 0.007974f
C3359 vdd.n1148 gnd 0.009907f
C3360 vdd.t185 gnd 0.506215f
C3361 vdd.n1149 gnd 0.703639f
C3362 vdd.n1150 gnd 0.009907f
C3363 vdd.n1151 gnd 0.007974f
C3364 vdd.n1152 gnd 0.009907f
C3365 vdd.n1153 gnd 0.007974f
C3366 vdd.n1154 gnd 0.009907f
C3367 vdd.n1155 gnd 0.804882f
C3368 vdd.n1156 gnd 0.009907f
C3369 vdd.n1157 gnd 0.007974f
C3370 vdd.n1158 gnd 0.009907f
C3371 vdd.n1159 gnd 0.007974f
C3372 vdd.n1160 gnd 0.009907f
C3373 vdd.n1161 gnd 0.632769f
C3374 vdd.t4 gnd 0.506215f
C3375 vdd.n1162 gnd 0.009907f
C3376 vdd.n1163 gnd 0.007974f
C3377 vdd.n1164 gnd 0.009907f
C3378 vdd.n1165 gnd 0.007974f
C3379 vdd.n1166 gnd 0.009907f
C3380 vdd.t220 gnd 0.506215f
C3381 vdd.n1167 gnd 0.009907f
C3382 vdd.n1168 gnd 0.007974f
C3383 vdd.n1169 gnd 0.009907f
C3384 vdd.n1170 gnd 0.007974f
C3385 vdd.n1171 gnd 0.009907f
C3386 vdd.t204 gnd 0.506215f
C3387 vdd.n1172 gnd 0.551774f
C3388 vdd.n1173 gnd 0.009907f
C3389 vdd.n1174 gnd 0.007974f
C3390 vdd.n1175 gnd 0.009907f
C3391 vdd.n1176 gnd 0.007974f
C3392 vdd.n1177 gnd 0.009907f
C3393 vdd.t6 gnd 0.506215f
C3394 vdd.n1178 gnd 0.009907f
C3395 vdd.n1179 gnd 0.007974f
C3396 vdd.n1180 gnd 0.009907f
C3397 vdd.n1181 gnd 0.007974f
C3398 vdd.n1182 gnd 0.009907f
C3399 vdd.n1183 gnd 0.784633f
C3400 vdd.n1184 gnd 0.840317f
C3401 vdd.t2 gnd 0.506215f
C3402 vdd.n1185 gnd 0.009907f
C3403 vdd.n1186 gnd 0.007974f
C3404 vdd.n1187 gnd 0.009907f
C3405 vdd.n1188 gnd 0.007974f
C3406 vdd.n1189 gnd 0.009907f
C3407 vdd.n1190 gnd 0.61252f
C3408 vdd.n1191 gnd 0.009907f
C3409 vdd.n1192 gnd 0.007974f
C3410 vdd.n1193 gnd 0.009907f
C3411 vdd.n1194 gnd 0.007974f
C3412 vdd.n1195 gnd 0.009907f
C3413 vdd.t17 gnd 0.506215f
C3414 vdd.t114 gnd 0.506215f
C3415 vdd.n1196 gnd 0.009907f
C3416 vdd.n1197 gnd 0.007974f
C3417 vdd.n1198 gnd 0.009907f
C3418 vdd.n1199 gnd 0.007974f
C3419 vdd.n1200 gnd 0.009907f
C3420 vdd.t12 gnd 0.506215f
C3421 vdd.n1201 gnd 0.009907f
C3422 vdd.n1202 gnd 0.007974f
C3423 vdd.n1203 gnd 0.009907f
C3424 vdd.n1204 gnd 0.007974f
C3425 vdd.n1205 gnd 0.009907f
C3426 vdd.t10 gnd 0.506215f
C3427 vdd.n1206 gnd 0.744136f
C3428 vdd.n1207 gnd 0.009907f
C3429 vdd.n1208 gnd 0.007974f
C3430 vdd.n1209 gnd 0.009907f
C3431 vdd.n1210 gnd 0.007974f
C3432 vdd.n1211 gnd 0.009907f
C3433 vdd.n1212 gnd 1.01243f
C3434 vdd.n1213 gnd 0.009907f
C3435 vdd.n1214 gnd 0.007974f
C3436 vdd.n1215 gnd 0.009907f
C3437 vdd.n1216 gnd 0.007974f
C3438 vdd.n1217 gnd 0.009907f
C3439 vdd.n1218 gnd 0.855503f
C3440 vdd.n1219 gnd 0.009907f
C3441 vdd.n1220 gnd 0.007974f
C3442 vdd.n1221 gnd 0.02256f
C3443 vdd.n1222 gnd 0.006618f
C3444 vdd.n1223 gnd 0.02256f
C3445 vdd.n1224 gnd 1.33641f
C3446 vdd.n1225 gnd 0.02256f
C3447 vdd.n1226 gnd 0.006618f
C3448 vdd.n1227 gnd 0.009907f
C3449 vdd.t57 gnd 0.12188f
C3450 vdd.t58 gnd 0.130256f
C3451 vdd.t55 gnd 0.159174f
C3452 vdd.n1228 gnd 0.204038f
C3453 vdd.n1229 gnd 0.172226f
C3454 vdd.n1230 gnd 0.013077f
C3455 vdd.n1231 gnd 0.009907f
C3456 vdd.n1262 gnd 0.009907f
C3457 vdd.n1263 gnd 0.009907f
C3458 vdd.n1264 gnd 0.022714f
C3459 vdd.n1265 gnd 0.007974f
C3460 vdd.n1266 gnd 0.009907f
C3461 vdd.n1267 gnd 0.009907f
C3462 vdd.n1268 gnd 0.009907f
C3463 vdd.n1269 gnd 0.009907f
C3464 vdd.n1270 gnd 0.007974f
C3465 vdd.n1271 gnd 0.009907f
C3466 vdd.n1272 gnd 0.009907f
C3467 vdd.n1273 gnd 0.009907f
C3468 vdd.n1274 gnd 0.009907f
C3469 vdd.n1275 gnd 0.009907f
C3470 vdd.n1276 gnd 0.007974f
C3471 vdd.n1277 gnd 0.009907f
C3472 vdd.n1278 gnd 0.009907f
C3473 vdd.n1279 gnd 0.009907f
C3474 vdd.n1280 gnd 0.009907f
C3475 vdd.n1281 gnd 0.009907f
C3476 vdd.n1282 gnd 0.007974f
C3477 vdd.n1283 gnd 0.009907f
C3478 vdd.n1284 gnd 0.009907f
C3479 vdd.n1285 gnd 0.009907f
C3480 vdd.n1286 gnd 0.009907f
C3481 vdd.n1287 gnd 0.009907f
C3482 vdd.n1288 gnd 0.006658f
C3483 vdd.n1289 gnd 0.009907f
C3484 vdd.n1290 gnd 0.009907f
C3485 vdd.n1291 gnd 0.009907f
C3486 vdd.n1292 gnd 0.007974f
C3487 vdd.n1293 gnd 0.009907f
C3488 vdd.n1294 gnd 0.009907f
C3489 vdd.n1295 gnd 0.009907f
C3490 vdd.n1296 gnd 0.009907f
C3491 vdd.n1297 gnd 0.009907f
C3492 vdd.n1298 gnd 0.007974f
C3493 vdd.n1299 gnd 0.009907f
C3494 vdd.n1300 gnd 0.009907f
C3495 vdd.n1301 gnd 0.009907f
C3496 vdd.n1302 gnd 0.009907f
C3497 vdd.n1303 gnd 0.009907f
C3498 vdd.n1304 gnd 0.007974f
C3499 vdd.n1305 gnd 0.009907f
C3500 vdd.n1306 gnd 0.009907f
C3501 vdd.n1307 gnd 0.009907f
C3502 vdd.n1308 gnd 0.009907f
C3503 vdd.n1309 gnd 0.009907f
C3504 vdd.n1310 gnd 0.007974f
C3505 vdd.n1311 gnd 0.009907f
C3506 vdd.n1312 gnd 0.009907f
C3507 vdd.n1313 gnd 0.009907f
C3508 vdd.n1314 gnd 0.009907f
C3509 vdd.n1315 gnd 0.009907f
C3510 vdd.n1316 gnd 0.007974f
C3511 vdd.n1317 gnd 0.009907f
C3512 vdd.n1318 gnd 0.009907f
C3513 vdd.n1319 gnd 0.009907f
C3514 vdd.n1320 gnd 0.009907f
C3515 vdd.n1321 gnd 0.007894f
C3516 vdd.n1322 gnd 0.009907f
C3517 vdd.n1323 gnd 0.009907f
C3518 vdd.n1324 gnd 0.009907f
C3519 vdd.n1325 gnd 0.009907f
C3520 vdd.n1326 gnd 0.009907f
C3521 vdd.n1327 gnd 0.007974f
C3522 vdd.n1328 gnd 0.009907f
C3523 vdd.n1329 gnd 0.009907f
C3524 vdd.n1330 gnd 0.009907f
C3525 vdd.n1331 gnd 0.009907f
C3526 vdd.n1332 gnd 0.009907f
C3527 vdd.n1333 gnd 0.007974f
C3528 vdd.n1334 gnd 0.009907f
C3529 vdd.n1335 gnd 0.009907f
C3530 vdd.n1336 gnd 0.009907f
C3531 vdd.n1337 gnd 0.009907f
C3532 vdd.n1338 gnd 0.009907f
C3533 vdd.n1339 gnd 0.007974f
C3534 vdd.n1340 gnd 0.009907f
C3535 vdd.n1341 gnd 0.009907f
C3536 vdd.n1342 gnd 0.009907f
C3537 vdd.n1343 gnd 0.009907f
C3538 vdd.n1344 gnd 0.009907f
C3539 vdd.n1345 gnd 0.007974f
C3540 vdd.n1346 gnd 0.009907f
C3541 vdd.n1347 gnd 0.009907f
C3542 vdd.n1348 gnd 0.009907f
C3543 vdd.n1349 gnd 0.009907f
C3544 vdd.n1350 gnd 0.009907f
C3545 vdd.n1351 gnd 0.004186f
C3546 vdd.n1352 gnd 0.009907f
C3547 vdd.n1353 gnd 0.007974f
C3548 vdd.n1354 gnd 0.007974f
C3549 vdd.n1355 gnd 0.007974f
C3550 vdd.n1356 gnd 0.009907f
C3551 vdd.n1357 gnd 0.009907f
C3552 vdd.n1358 gnd 0.009907f
C3553 vdd.n1359 gnd 0.007974f
C3554 vdd.n1360 gnd 0.007974f
C3555 vdd.n1361 gnd 0.007974f
C3556 vdd.n1362 gnd 0.009907f
C3557 vdd.n1363 gnd 0.009907f
C3558 vdd.n1364 gnd 0.009907f
C3559 vdd.n1365 gnd 0.007974f
C3560 vdd.n1366 gnd 0.007974f
C3561 vdd.n1367 gnd 0.007974f
C3562 vdd.n1368 gnd 0.009907f
C3563 vdd.n1369 gnd 0.009907f
C3564 vdd.n1370 gnd 0.009907f
C3565 vdd.n1371 gnd 0.007974f
C3566 vdd.n1372 gnd 0.007974f
C3567 vdd.n1373 gnd 0.007974f
C3568 vdd.n1374 gnd 0.009907f
C3569 vdd.n1375 gnd 0.009907f
C3570 vdd.n1376 gnd 0.009907f
C3571 vdd.n1377 gnd 0.007974f
C3572 vdd.n1378 gnd 0.007974f
C3573 vdd.n1379 gnd 0.007974f
C3574 vdd.n1380 gnd 0.009907f
C3575 vdd.n1381 gnd 0.009907f
C3576 vdd.n1382 gnd 0.009907f
C3577 vdd.n1383 gnd 0.009907f
C3578 vdd.t80 gnd 0.12188f
C3579 vdd.t81 gnd 0.130256f
C3580 vdd.t79 gnd 0.159174f
C3581 vdd.n1384 gnd 0.204038f
C3582 vdd.n1385 gnd 0.172226f
C3583 vdd.n1386 gnd 0.017064f
C3584 vdd.n1387 gnd 0.005422f
C3585 vdd.n1388 gnd 0.007974f
C3586 vdd.n1389 gnd 0.009907f
C3587 vdd.n1390 gnd 0.009907f
C3588 vdd.n1391 gnd 0.009907f
C3589 vdd.n1392 gnd 0.007974f
C3590 vdd.n1393 gnd 0.007974f
C3591 vdd.n1394 gnd 0.007974f
C3592 vdd.n1395 gnd 0.009907f
C3593 vdd.n1396 gnd 0.009907f
C3594 vdd.n1397 gnd 0.009907f
C3595 vdd.n1398 gnd 0.007974f
C3596 vdd.n1399 gnd 0.007974f
C3597 vdd.n1400 gnd 0.007974f
C3598 vdd.n1401 gnd 0.009907f
C3599 vdd.n1402 gnd 0.009907f
C3600 vdd.n1403 gnd 0.009907f
C3601 vdd.n1404 gnd 0.007974f
C3602 vdd.n1405 gnd 0.007974f
C3603 vdd.n1406 gnd 0.007974f
C3604 vdd.n1407 gnd 0.009907f
C3605 vdd.n1408 gnd 0.009907f
C3606 vdd.n1409 gnd 0.009907f
C3607 vdd.n1410 gnd 0.007974f
C3608 vdd.n1411 gnd 0.007974f
C3609 vdd.n1412 gnd 0.007974f
C3610 vdd.n1413 gnd 0.009907f
C3611 vdd.n1414 gnd 0.009907f
C3612 vdd.n1415 gnd 0.009907f
C3613 vdd.n1416 gnd 0.007974f
C3614 vdd.n1417 gnd 0.006658f
C3615 vdd.n1418 gnd 0.009907f
C3616 vdd.n1419 gnd 0.009907f
C3617 vdd.t93 gnd 0.12188f
C3618 vdd.t94 gnd 0.130256f
C3619 vdd.t92 gnd 0.159174f
C3620 vdd.n1420 gnd 0.204038f
C3621 vdd.n1421 gnd 0.172226f
C3622 vdd.n1422 gnd 0.017064f
C3623 vdd.n1423 gnd 0.009907f
C3624 vdd.n1424 gnd 0.009907f
C3625 vdd.n1425 gnd 0.009907f
C3626 vdd.n1426 gnd 0.007974f
C3627 vdd.n1427 gnd 0.007974f
C3628 vdd.n1428 gnd 0.007974f
C3629 vdd.n1429 gnd 0.009907f
C3630 vdd.n1430 gnd 0.009907f
C3631 vdd.n1431 gnd 0.009907f
C3632 vdd.n1432 gnd 0.007974f
C3633 vdd.n1433 gnd 0.007974f
C3634 vdd.n1434 gnd 0.007974f
C3635 vdd.n1435 gnd 0.009907f
C3636 vdd.n1436 gnd 0.009907f
C3637 vdd.n1437 gnd 0.009907f
C3638 vdd.n1438 gnd 0.007974f
C3639 vdd.n1439 gnd 0.007974f
C3640 vdd.n1440 gnd 0.007974f
C3641 vdd.n1441 gnd 0.009907f
C3642 vdd.n1442 gnd 0.009907f
C3643 vdd.n1443 gnd 0.009907f
C3644 vdd.n1444 gnd 0.007974f
C3645 vdd.n1445 gnd 0.007974f
C3646 vdd.n1446 gnd 0.007974f
C3647 vdd.n1447 gnd 0.009907f
C3648 vdd.n1448 gnd 0.009907f
C3649 vdd.n1449 gnd 0.009907f
C3650 vdd.n1450 gnd 0.007974f
C3651 vdd.n1451 gnd 0.006618f
C3652 vdd.n1452 gnd 0.022714f
C3653 vdd.n1454 gnd 2.23747f
C3654 vdd.n1455 gnd 0.022714f
C3655 vdd.n1456 gnd 0.003788f
C3656 vdd.n1457 gnd 0.022714f
C3657 vdd.n1458 gnd 0.02256f
C3658 vdd.n1459 gnd 0.009907f
C3659 vdd.n1460 gnd 0.007974f
C3660 vdd.n1461 gnd 0.009907f
C3661 vdd.t56 gnd 0.506215f
C3662 vdd.n1462 gnd 0.663142f
C3663 vdd.n1463 gnd 0.009907f
C3664 vdd.n1464 gnd 0.007974f
C3665 vdd.n1465 gnd 0.009907f
C3666 vdd.n1466 gnd 0.009907f
C3667 vdd.n1467 gnd 0.009907f
C3668 vdd.n1468 gnd 0.007974f
C3669 vdd.n1469 gnd 0.009907f
C3670 vdd.n1470 gnd 1.01243f
C3671 vdd.n1471 gnd 0.009907f
C3672 vdd.n1472 gnd 0.007974f
C3673 vdd.n1473 gnd 0.009907f
C3674 vdd.n1474 gnd 0.009907f
C3675 vdd.n1475 gnd 0.009907f
C3676 vdd.n1476 gnd 0.007974f
C3677 vdd.n1477 gnd 0.009907f
C3678 vdd.n1478 gnd 0.840317f
C3679 vdd.t21 gnd 0.506215f
C3680 vdd.n1479 gnd 0.582147f
C3681 vdd.n1480 gnd 0.009907f
C3682 vdd.n1481 gnd 0.007974f
C3683 vdd.n1482 gnd 0.009907f
C3684 vdd.n1483 gnd 0.009907f
C3685 vdd.n1484 gnd 0.009907f
C3686 vdd.n1485 gnd 0.007974f
C3687 vdd.n1486 gnd 0.009907f
C3688 vdd.n1487 gnd 0.602396f
C3689 vdd.n1488 gnd 0.009907f
C3690 vdd.n1489 gnd 0.007974f
C3691 vdd.n1490 gnd 0.009907f
C3692 vdd.n1491 gnd 0.009907f
C3693 vdd.n1492 gnd 0.009907f
C3694 vdd.n1493 gnd 0.007974f
C3695 vdd.n1494 gnd 0.009907f
C3696 vdd.n1495 gnd 0.572023f
C3697 vdd.n1496 gnd 0.774509f
C3698 vdd.n1497 gnd 0.009907f
C3699 vdd.n1498 gnd 0.007974f
C3700 vdd.n1499 gnd 0.009907f
C3701 vdd.n1500 gnd 0.009907f
C3702 vdd.n1501 gnd 0.009907f
C3703 vdd.n1502 gnd 0.007974f
C3704 vdd.n1503 gnd 0.009907f
C3705 vdd.n1504 gnd 0.840317f
C3706 vdd.n1505 gnd 0.009907f
C3707 vdd.n1506 gnd 0.007974f
C3708 vdd.n1507 gnd 0.009907f
C3709 vdd.n1508 gnd 0.009907f
C3710 vdd.n1509 gnd 0.009907f
C3711 vdd.n1510 gnd 0.007974f
C3712 vdd.n1511 gnd 0.009907f
C3713 vdd.t199 gnd 0.506215f
C3714 vdd.n1512 gnd 0.734012f
C3715 vdd.n1513 gnd 0.009907f
C3716 vdd.n1514 gnd 0.007974f
C3717 vdd.n1515 gnd 0.009907f
C3718 vdd.n1516 gnd 0.009907f
C3719 vdd.n1517 gnd 0.009907f
C3720 vdd.n1518 gnd 0.007974f
C3721 vdd.n1519 gnd 0.009907f
C3722 vdd.n1520 gnd 0.561899f
C3723 vdd.n1521 gnd 0.009907f
C3724 vdd.n1522 gnd 0.007974f
C3725 vdd.n1523 gnd 0.009907f
C3726 vdd.n1524 gnd 0.009907f
C3727 vdd.n1525 gnd 0.009907f
C3728 vdd.n1526 gnd 0.007974f
C3729 vdd.n1527 gnd 0.009907f
C3730 vdd.n1528 gnd 0.723888f
C3731 vdd.n1529 gnd 0.622645f
C3732 vdd.n1530 gnd 0.009907f
C3733 vdd.n1531 gnd 0.007974f
C3734 vdd.n1532 gnd 0.007614f
C3735 vdd.n1533 gnd 0.005437f
C3736 vdd.n1534 gnd 0.005045f
C3737 vdd.n1535 gnd 0.002791f
C3738 vdd.n1536 gnd 0.006408f
C3739 vdd.n1537 gnd 0.002711f
C3740 vdd.n1538 gnd 0.002871f
C3741 vdd.n1539 gnd 0.005045f
C3742 vdd.n1540 gnd 0.002711f
C3743 vdd.n1541 gnd 0.006408f
C3744 vdd.n1542 gnd 0.002871f
C3745 vdd.n1543 gnd 0.005045f
C3746 vdd.n1544 gnd 0.002711f
C3747 vdd.n1545 gnd 0.004806f
C3748 vdd.n1546 gnd 0.00482f
C3749 vdd.t239 gnd 0.013767f
C3750 vdd.n1547 gnd 0.030632f
C3751 vdd.n1548 gnd 0.159414f
C3752 vdd.n1549 gnd 0.002711f
C3753 vdd.n1550 gnd 0.002871f
C3754 vdd.n1551 gnd 0.006408f
C3755 vdd.n1552 gnd 0.006408f
C3756 vdd.n1553 gnd 0.002871f
C3757 vdd.n1554 gnd 0.002711f
C3758 vdd.n1555 gnd 0.005045f
C3759 vdd.n1556 gnd 0.005045f
C3760 vdd.n1557 gnd 0.002711f
C3761 vdd.n1558 gnd 0.002871f
C3762 vdd.n1559 gnd 0.006408f
C3763 vdd.n1560 gnd 0.006408f
C3764 vdd.n1561 gnd 0.002871f
C3765 vdd.n1562 gnd 0.002711f
C3766 vdd.n1563 gnd 0.005045f
C3767 vdd.n1564 gnd 0.005045f
C3768 vdd.n1565 gnd 0.002711f
C3769 vdd.n1566 gnd 0.002871f
C3770 vdd.n1567 gnd 0.006408f
C3771 vdd.n1568 gnd 0.006408f
C3772 vdd.n1569 gnd 0.01515f
C3773 vdd.n1570 gnd 0.002791f
C3774 vdd.n1571 gnd 0.002711f
C3775 vdd.n1572 gnd 0.01304f
C3776 vdd.n1573 gnd 0.009104f
C3777 vdd.t186 gnd 0.031895f
C3778 vdd.t104 gnd 0.031895f
C3779 vdd.n1574 gnd 0.219206f
C3780 vdd.n1575 gnd 0.172372f
C3781 vdd.t219 gnd 0.031895f
C3782 vdd.t106 gnd 0.031895f
C3783 vdd.n1576 gnd 0.219206f
C3784 vdd.n1577 gnd 0.139103f
C3785 vdd.t258 gnd 0.031895f
C3786 vdd.t236 gnd 0.031895f
C3787 vdd.n1578 gnd 0.219206f
C3788 vdd.n1579 gnd 0.139103f
C3789 vdd.t252 gnd 0.031895f
C3790 vdd.t205 gnd 0.031895f
C3791 vdd.n1580 gnd 0.219206f
C3792 vdd.n1581 gnd 0.139103f
C3793 vdd.t200 gnd 0.031895f
C3794 vdd.t123 gnd 0.031895f
C3795 vdd.n1582 gnd 0.219206f
C3796 vdd.n1583 gnd 0.139103f
C3797 vdd.t250 gnd 0.031895f
C3798 vdd.t260 gnd 0.031895f
C3799 vdd.n1584 gnd 0.219206f
C3800 vdd.n1585 gnd 0.139103f
C3801 vdd.t113 gnd 0.031895f
C3802 vdd.t13 gnd 0.031895f
C3803 vdd.n1586 gnd 0.219206f
C3804 vdd.n1587 gnd 0.139103f
C3805 vdd.n1588 gnd 0.005437f
C3806 vdd.n1589 gnd 0.005045f
C3807 vdd.n1590 gnd 0.002791f
C3808 vdd.n1591 gnd 0.006408f
C3809 vdd.n1592 gnd 0.002711f
C3810 vdd.n1593 gnd 0.002871f
C3811 vdd.n1594 gnd 0.005045f
C3812 vdd.n1595 gnd 0.002711f
C3813 vdd.n1596 gnd 0.006408f
C3814 vdd.n1597 gnd 0.002871f
C3815 vdd.n1598 gnd 0.005045f
C3816 vdd.n1599 gnd 0.002711f
C3817 vdd.n1600 gnd 0.004806f
C3818 vdd.n1601 gnd 0.00482f
C3819 vdd.t203 gnd 0.013767f
C3820 vdd.n1602 gnd 0.030632f
C3821 vdd.n1603 gnd 0.159414f
C3822 vdd.n1604 gnd 0.002711f
C3823 vdd.n1605 gnd 0.002871f
C3824 vdd.n1606 gnd 0.006408f
C3825 vdd.n1607 gnd 0.006408f
C3826 vdd.n1608 gnd 0.002871f
C3827 vdd.n1609 gnd 0.002711f
C3828 vdd.n1610 gnd 0.005045f
C3829 vdd.n1611 gnd 0.005045f
C3830 vdd.n1612 gnd 0.002711f
C3831 vdd.n1613 gnd 0.002871f
C3832 vdd.n1614 gnd 0.006408f
C3833 vdd.n1615 gnd 0.006408f
C3834 vdd.n1616 gnd 0.002871f
C3835 vdd.n1617 gnd 0.002711f
C3836 vdd.n1618 gnd 0.005045f
C3837 vdd.n1619 gnd 0.005045f
C3838 vdd.n1620 gnd 0.002711f
C3839 vdd.n1621 gnd 0.002871f
C3840 vdd.n1622 gnd 0.006408f
C3841 vdd.n1623 gnd 0.006408f
C3842 vdd.n1624 gnd 0.01515f
C3843 vdd.n1625 gnd 0.002791f
C3844 vdd.n1626 gnd 0.002711f
C3845 vdd.n1627 gnd 0.01304f
C3846 vdd.n1628 gnd 0.008818f
C3847 vdd.n1629 gnd 0.103493f
C3848 vdd.n1630 gnd 0.005437f
C3849 vdd.n1631 gnd 0.005045f
C3850 vdd.n1632 gnd 0.002791f
C3851 vdd.n1633 gnd 0.006408f
C3852 vdd.n1634 gnd 0.002711f
C3853 vdd.n1635 gnd 0.002871f
C3854 vdd.n1636 gnd 0.005045f
C3855 vdd.n1637 gnd 0.002711f
C3856 vdd.n1638 gnd 0.006408f
C3857 vdd.n1639 gnd 0.002871f
C3858 vdd.n1640 gnd 0.005045f
C3859 vdd.n1641 gnd 0.002711f
C3860 vdd.n1642 gnd 0.004806f
C3861 vdd.n1643 gnd 0.00482f
C3862 vdd.t249 gnd 0.013767f
C3863 vdd.n1644 gnd 0.030632f
C3864 vdd.n1645 gnd 0.159414f
C3865 vdd.n1646 gnd 0.002711f
C3866 vdd.n1647 gnd 0.002871f
C3867 vdd.n1648 gnd 0.006408f
C3868 vdd.n1649 gnd 0.006408f
C3869 vdd.n1650 gnd 0.002871f
C3870 vdd.n1651 gnd 0.002711f
C3871 vdd.n1652 gnd 0.005045f
C3872 vdd.n1653 gnd 0.005045f
C3873 vdd.n1654 gnd 0.002711f
C3874 vdd.n1655 gnd 0.002871f
C3875 vdd.n1656 gnd 0.006408f
C3876 vdd.n1657 gnd 0.006408f
C3877 vdd.n1658 gnd 0.002871f
C3878 vdd.n1659 gnd 0.002711f
C3879 vdd.n1660 gnd 0.005045f
C3880 vdd.n1661 gnd 0.005045f
C3881 vdd.n1662 gnd 0.002711f
C3882 vdd.n1663 gnd 0.002871f
C3883 vdd.n1664 gnd 0.006408f
C3884 vdd.n1665 gnd 0.006408f
C3885 vdd.n1666 gnd 0.01515f
C3886 vdd.n1667 gnd 0.002791f
C3887 vdd.n1668 gnd 0.002711f
C3888 vdd.n1669 gnd 0.01304f
C3889 vdd.n1670 gnd 0.009104f
C3890 vdd.t265 gnd 0.031895f
C3891 vdd.t241 gnd 0.031895f
C3892 vdd.n1671 gnd 0.219206f
C3893 vdd.n1672 gnd 0.172372f
C3894 vdd.t5 gnd 0.031895f
C3895 vdd.t238 gnd 0.031895f
C3896 vdd.n1673 gnd 0.219206f
C3897 vdd.n1674 gnd 0.139103f
C3898 vdd.t221 gnd 0.031895f
C3899 vdd.t240 gnd 0.031895f
C3900 vdd.n1675 gnd 0.219206f
C3901 vdd.n1676 gnd 0.139103f
C3902 vdd.t7 gnd 0.031895f
C3903 vdd.t262 gnd 0.031895f
C3904 vdd.n1677 gnd 0.219206f
C3905 vdd.n1678 gnd 0.139103f
C3906 vdd.t242 gnd 0.031895f
C3907 vdd.t14 gnd 0.031895f
C3908 vdd.n1679 gnd 0.219206f
C3909 vdd.n1680 gnd 0.139103f
C3910 vdd.t128 gnd 0.031895f
C3911 vdd.t188 gnd 0.031895f
C3912 vdd.n1681 gnd 0.219206f
C3913 vdd.n1682 gnd 0.139103f
C3914 vdd.t189 gnd 0.031895f
C3915 vdd.t237 gnd 0.031895f
C3916 vdd.n1683 gnd 0.219206f
C3917 vdd.n1684 gnd 0.139103f
C3918 vdd.n1685 gnd 0.005437f
C3919 vdd.n1686 gnd 0.005045f
C3920 vdd.n1687 gnd 0.002791f
C3921 vdd.n1688 gnd 0.006408f
C3922 vdd.n1689 gnd 0.002711f
C3923 vdd.n1690 gnd 0.002871f
C3924 vdd.n1691 gnd 0.005045f
C3925 vdd.n1692 gnd 0.002711f
C3926 vdd.n1693 gnd 0.006408f
C3927 vdd.n1694 gnd 0.002871f
C3928 vdd.n1695 gnd 0.005045f
C3929 vdd.n1696 gnd 0.002711f
C3930 vdd.n1697 gnd 0.004806f
C3931 vdd.n1698 gnd 0.00482f
C3932 vdd.t22 gnd 0.013767f
C3933 vdd.n1699 gnd 0.030632f
C3934 vdd.n1700 gnd 0.159414f
C3935 vdd.n1701 gnd 0.002711f
C3936 vdd.n1702 gnd 0.002871f
C3937 vdd.n1703 gnd 0.006408f
C3938 vdd.n1704 gnd 0.006408f
C3939 vdd.n1705 gnd 0.002871f
C3940 vdd.n1706 gnd 0.002711f
C3941 vdd.n1707 gnd 0.005045f
C3942 vdd.n1708 gnd 0.005045f
C3943 vdd.n1709 gnd 0.002711f
C3944 vdd.n1710 gnd 0.002871f
C3945 vdd.n1711 gnd 0.006408f
C3946 vdd.n1712 gnd 0.006408f
C3947 vdd.n1713 gnd 0.002871f
C3948 vdd.n1714 gnd 0.002711f
C3949 vdd.n1715 gnd 0.005045f
C3950 vdd.n1716 gnd 0.005045f
C3951 vdd.n1717 gnd 0.002711f
C3952 vdd.n1718 gnd 0.002871f
C3953 vdd.n1719 gnd 0.006408f
C3954 vdd.n1720 gnd 0.006408f
C3955 vdd.n1721 gnd 0.01515f
C3956 vdd.n1722 gnd 0.002791f
C3957 vdd.n1723 gnd 0.002711f
C3958 vdd.n1724 gnd 0.01304f
C3959 vdd.n1725 gnd 0.008818f
C3960 vdd.n1726 gnd 0.061568f
C3961 vdd.n1727 gnd 0.221846f
C3962 vdd.n1728 gnd 0.005437f
C3963 vdd.n1729 gnd 0.005045f
C3964 vdd.n1730 gnd 0.002791f
C3965 vdd.n1731 gnd 0.006408f
C3966 vdd.n1732 gnd 0.002711f
C3967 vdd.n1733 gnd 0.002871f
C3968 vdd.n1734 gnd 0.005045f
C3969 vdd.n1735 gnd 0.002711f
C3970 vdd.n1736 gnd 0.006408f
C3971 vdd.n1737 gnd 0.002871f
C3972 vdd.n1738 gnd 0.005045f
C3973 vdd.n1739 gnd 0.002711f
C3974 vdd.n1740 gnd 0.004806f
C3975 vdd.n1741 gnd 0.00482f
C3976 vdd.t235 gnd 0.013767f
C3977 vdd.n1742 gnd 0.030632f
C3978 vdd.n1743 gnd 0.159414f
C3979 vdd.n1744 gnd 0.002711f
C3980 vdd.n1745 gnd 0.002871f
C3981 vdd.n1746 gnd 0.006408f
C3982 vdd.n1747 gnd 0.006408f
C3983 vdd.n1748 gnd 0.002871f
C3984 vdd.n1749 gnd 0.002711f
C3985 vdd.n1750 gnd 0.005045f
C3986 vdd.n1751 gnd 0.005045f
C3987 vdd.n1752 gnd 0.002711f
C3988 vdd.n1753 gnd 0.002871f
C3989 vdd.n1754 gnd 0.006408f
C3990 vdd.n1755 gnd 0.006408f
C3991 vdd.n1756 gnd 0.002871f
C3992 vdd.n1757 gnd 0.002711f
C3993 vdd.n1758 gnd 0.005045f
C3994 vdd.n1759 gnd 0.005045f
C3995 vdd.n1760 gnd 0.002711f
C3996 vdd.n1761 gnd 0.002871f
C3997 vdd.n1762 gnd 0.006408f
C3998 vdd.n1763 gnd 0.006408f
C3999 vdd.n1764 gnd 0.01515f
C4000 vdd.n1765 gnd 0.002791f
C4001 vdd.n1766 gnd 0.002711f
C4002 vdd.n1767 gnd 0.01304f
C4003 vdd.n1768 gnd 0.009104f
C4004 vdd.t217 gnd 0.031895f
C4005 vdd.t254 gnd 0.031895f
C4006 vdd.n1769 gnd 0.219206f
C4007 vdd.n1770 gnd 0.172372f
C4008 vdd.t261 gnd 0.031895f
C4009 vdd.t243 gnd 0.031895f
C4010 vdd.n1771 gnd 0.219206f
C4011 vdd.n1772 gnd 0.139103f
C4012 vdd.t266 gnd 0.031895f
C4013 vdd.t1 gnd 0.031895f
C4014 vdd.n1773 gnd 0.219206f
C4015 vdd.n1774 gnd 0.139103f
C4016 vdd.t187 gnd 0.031895f
C4017 vdd.t245 gnd 0.031895f
C4018 vdd.n1775 gnd 0.219206f
C4019 vdd.n1776 gnd 0.139103f
C4020 vdd.t208 gnd 0.031895f
C4021 vdd.t3 gnd 0.031895f
C4022 vdd.n1777 gnd 0.219206f
C4023 vdd.n1778 gnd 0.139103f
C4024 vdd.t18 gnd 0.031895f
C4025 vdd.t115 gnd 0.031895f
C4026 vdd.n1779 gnd 0.219206f
C4027 vdd.n1780 gnd 0.139103f
C4028 vdd.t11 gnd 0.031895f
C4029 vdd.t197 gnd 0.031895f
C4030 vdd.n1781 gnd 0.219206f
C4031 vdd.n1782 gnd 0.139103f
C4032 vdd.n1783 gnd 0.005437f
C4033 vdd.n1784 gnd 0.005045f
C4034 vdd.n1785 gnd 0.002791f
C4035 vdd.n1786 gnd 0.006408f
C4036 vdd.n1787 gnd 0.002711f
C4037 vdd.n1788 gnd 0.002871f
C4038 vdd.n1789 gnd 0.005045f
C4039 vdd.n1790 gnd 0.002711f
C4040 vdd.n1791 gnd 0.006408f
C4041 vdd.n1792 gnd 0.002871f
C4042 vdd.n1793 gnd 0.005045f
C4043 vdd.n1794 gnd 0.002711f
C4044 vdd.n1795 gnd 0.004806f
C4045 vdd.n1796 gnd 0.00482f
C4046 vdd.t201 gnd 0.013767f
C4047 vdd.n1797 gnd 0.030632f
C4048 vdd.n1798 gnd 0.159414f
C4049 vdd.n1799 gnd 0.002711f
C4050 vdd.n1800 gnd 0.002871f
C4051 vdd.n1801 gnd 0.006408f
C4052 vdd.n1802 gnd 0.006408f
C4053 vdd.n1803 gnd 0.002871f
C4054 vdd.n1804 gnd 0.002711f
C4055 vdd.n1805 gnd 0.005045f
C4056 vdd.n1806 gnd 0.005045f
C4057 vdd.n1807 gnd 0.002711f
C4058 vdd.n1808 gnd 0.002871f
C4059 vdd.n1809 gnd 0.006408f
C4060 vdd.n1810 gnd 0.006408f
C4061 vdd.n1811 gnd 0.002871f
C4062 vdd.n1812 gnd 0.002711f
C4063 vdd.n1813 gnd 0.005045f
C4064 vdd.n1814 gnd 0.005045f
C4065 vdd.n1815 gnd 0.002711f
C4066 vdd.n1816 gnd 0.002871f
C4067 vdd.n1817 gnd 0.006408f
C4068 vdd.n1818 gnd 0.006408f
C4069 vdd.n1819 gnd 0.01515f
C4070 vdd.n1820 gnd 0.002791f
C4071 vdd.n1821 gnd 0.002711f
C4072 vdd.n1822 gnd 0.01304f
C4073 vdd.n1823 gnd 0.008818f
C4074 vdd.n1824 gnd 0.061568f
C4075 vdd.n1825 gnd 0.248438f
C4076 vdd.n1826 gnd 2.60929f
C4077 vdd.n1827 gnd 0.584342f
C4078 vdd.n1828 gnd 0.007614f
C4079 vdd.n1829 gnd 0.009907f
C4080 vdd.n1830 gnd 0.007974f
C4081 vdd.n1831 gnd 0.009907f
C4082 vdd.n1832 gnd 0.794758f
C4083 vdd.n1833 gnd 0.009907f
C4084 vdd.n1834 gnd 0.007974f
C4085 vdd.n1835 gnd 0.009907f
C4086 vdd.n1836 gnd 0.009907f
C4087 vdd.n1837 gnd 0.009907f
C4088 vdd.n1838 gnd 0.007974f
C4089 vdd.n1839 gnd 0.009907f
C4090 vdd.t0 gnd 0.506215f
C4091 vdd.n1840 gnd 0.840317f
C4092 vdd.n1841 gnd 0.009907f
C4093 vdd.n1842 gnd 0.007974f
C4094 vdd.n1843 gnd 0.009907f
C4095 vdd.n1844 gnd 0.009907f
C4096 vdd.n1845 gnd 0.009907f
C4097 vdd.n1846 gnd 0.007974f
C4098 vdd.n1847 gnd 0.009907f
C4099 vdd.n1848 gnd 0.713763f
C4100 vdd.n1849 gnd 0.009907f
C4101 vdd.n1850 gnd 0.007974f
C4102 vdd.n1851 gnd 0.009907f
C4103 vdd.n1852 gnd 0.009907f
C4104 vdd.n1853 gnd 0.009907f
C4105 vdd.n1854 gnd 0.007974f
C4106 vdd.n1855 gnd 0.009907f
C4107 vdd.n1856 gnd 0.840317f
C4108 vdd.t105 gnd 0.506215f
C4109 vdd.n1857 gnd 0.54165f
C4110 vdd.n1858 gnd 0.009907f
C4111 vdd.n1859 gnd 0.007974f
C4112 vdd.n1860 gnd 0.009907f
C4113 vdd.n1861 gnd 0.009907f
C4114 vdd.n1862 gnd 0.009907f
C4115 vdd.n1863 gnd 0.007974f
C4116 vdd.n1864 gnd 0.009907f
C4117 vdd.n1865 gnd 0.642893f
C4118 vdd.n1866 gnd 0.009907f
C4119 vdd.n1867 gnd 0.007974f
C4120 vdd.n1868 gnd 0.009907f
C4121 vdd.n1869 gnd 0.009907f
C4122 vdd.n1870 gnd 0.009907f
C4123 vdd.n1871 gnd 0.007974f
C4124 vdd.n1872 gnd 0.009907f
C4125 vdd.n1873 gnd 0.531526f
C4126 vdd.n1874 gnd 0.815006f
C4127 vdd.n1875 gnd 0.009907f
C4128 vdd.n1876 gnd 0.007974f
C4129 vdd.n1877 gnd 0.009907f
C4130 vdd.n1878 gnd 0.009907f
C4131 vdd.n1879 gnd 0.009907f
C4132 vdd.n1880 gnd 0.007974f
C4133 vdd.n1881 gnd 0.009907f
C4134 vdd.n1882 gnd 0.987119f
C4135 vdd.n1883 gnd 0.009907f
C4136 vdd.n1884 gnd 0.007974f
C4137 vdd.n1885 gnd 0.009907f
C4138 vdd.n1886 gnd 0.009907f
C4139 vdd.n1887 gnd 0.02256f
C4140 vdd.n1888 gnd 0.009907f
C4141 vdd.n1889 gnd 0.009907f
C4142 vdd.n1890 gnd 0.007974f
C4143 vdd.n1891 gnd 0.009907f
C4144 vdd.t52 gnd 0.506215f
C4145 vdd.n1892 gnd 0.956746f
C4146 vdd.n1893 gnd 0.009907f
C4147 vdd.n1894 gnd 0.007974f
C4148 vdd.n1895 gnd 0.009907f
C4149 vdd.n1896 gnd 0.009907f
C4150 vdd.n1897 gnd 0.00852f
C4151 vdd.n1898 gnd 0.007974f
C4152 vdd.n1900 gnd 0.009907f
C4153 vdd.n1902 gnd 0.007974f
C4154 vdd.n1903 gnd 0.009907f
C4155 vdd.n1904 gnd 0.007974f
C4156 vdd.n1906 gnd 0.009907f
C4157 vdd.n1907 gnd 0.007974f
C4158 vdd.n1908 gnd 0.009907f
C4159 vdd.n1909 gnd 0.009907f
C4160 vdd.n1910 gnd 0.009907f
C4161 vdd.n1911 gnd 0.009907f
C4162 vdd.n1912 gnd 0.009907f
C4163 vdd.n1913 gnd 0.007974f
C4164 vdd.n1915 gnd 0.009907f
C4165 vdd.n1916 gnd 0.009907f
C4166 vdd.n1917 gnd 0.009907f
C4167 vdd.n1918 gnd 0.009907f
C4168 vdd.n1919 gnd 0.009907f
C4169 vdd.n1920 gnd 0.007974f
C4170 vdd.n1922 gnd 0.009907f
C4171 vdd.n1923 gnd 0.009907f
C4172 vdd.n1924 gnd 0.009907f
C4173 vdd.n1925 gnd 0.009907f
C4174 vdd.n1926 gnd 0.006658f
C4175 vdd.t84 gnd 0.12188f
C4176 vdd.t83 gnd 0.130256f
C4177 vdd.t82 gnd 0.159174f
C4178 vdd.n1927 gnd 0.204038f
C4179 vdd.n1928 gnd 0.171429f
C4180 vdd.n1930 gnd 0.009907f
C4181 vdd.n1931 gnd 0.009907f
C4182 vdd.n1932 gnd 0.007974f
C4183 vdd.n1933 gnd 0.009907f
C4184 vdd.n1935 gnd 0.009907f
C4185 vdd.n1936 gnd 0.009907f
C4186 vdd.n1937 gnd 0.009907f
C4187 vdd.n1938 gnd 0.009907f
C4188 vdd.n1939 gnd 0.007974f
C4189 vdd.n1941 gnd 0.009907f
C4190 vdd.n1942 gnd 0.009907f
C4191 vdd.n1943 gnd 0.009907f
C4192 vdd.n1944 gnd 0.009907f
C4193 vdd.n1945 gnd 0.009907f
C4194 vdd.n1946 gnd 0.007974f
C4195 vdd.n1948 gnd 0.009907f
C4196 vdd.n1949 gnd 0.009907f
C4197 vdd.n1950 gnd 0.009907f
C4198 vdd.n1951 gnd 0.009907f
C4199 vdd.n1952 gnd 0.009907f
C4200 vdd.n1953 gnd 0.007974f
C4201 vdd.n1955 gnd 0.009907f
C4202 vdd.n1956 gnd 0.009907f
C4203 vdd.n1957 gnd 0.009907f
C4204 vdd.n1958 gnd 0.009907f
C4205 vdd.n1959 gnd 0.009907f
C4206 vdd.n1960 gnd 0.007974f
C4207 vdd.n1962 gnd 0.009907f
C4208 vdd.n1963 gnd 0.009907f
C4209 vdd.n1964 gnd 0.009907f
C4210 vdd.n1965 gnd 0.009907f
C4211 vdd.n1966 gnd 0.007894f
C4212 vdd.t70 gnd 0.12188f
C4213 vdd.t69 gnd 0.130256f
C4214 vdd.t68 gnd 0.159174f
C4215 vdd.n1967 gnd 0.204038f
C4216 vdd.n1968 gnd 0.171429f
C4217 vdd.n1970 gnd 0.009907f
C4218 vdd.n1971 gnd 0.009907f
C4219 vdd.n1972 gnd 0.007974f
C4220 vdd.n1973 gnd 0.009907f
C4221 vdd.n1975 gnd 0.009907f
C4222 vdd.n1976 gnd 0.009907f
C4223 vdd.n1977 gnd 0.009907f
C4224 vdd.n1978 gnd 0.009907f
C4225 vdd.n1979 gnd 0.007974f
C4226 vdd.n1981 gnd 0.009907f
C4227 vdd.n1982 gnd 0.009907f
C4228 vdd.n1983 gnd 0.009907f
C4229 vdd.n1984 gnd 0.009907f
C4230 vdd.n1985 gnd 0.009907f
C4231 vdd.n1986 gnd 0.007974f
C4232 vdd.n1988 gnd 0.009907f
C4233 vdd.n1989 gnd 0.009907f
C4234 vdd.n1990 gnd 0.009907f
C4235 vdd.n1991 gnd 0.009907f
C4236 vdd.n1992 gnd 0.009907f
C4237 vdd.n1993 gnd 0.009907f
C4238 vdd.n1994 gnd 0.007974f
C4239 vdd.n1996 gnd 0.009907f
C4240 vdd.n1998 gnd 0.009907f
C4241 vdd.n1999 gnd 0.007974f
C4242 vdd.n2000 gnd 0.007974f
C4243 vdd.n2001 gnd 0.009907f
C4244 vdd.n2003 gnd 0.009907f
C4245 vdd.n2004 gnd 0.007974f
C4246 vdd.n2005 gnd 0.007974f
C4247 vdd.n2006 gnd 0.009907f
C4248 vdd.n2008 gnd 0.009907f
C4249 vdd.n2009 gnd 0.009907f
C4250 vdd.n2010 gnd 0.007974f
C4251 vdd.n2011 gnd 0.007974f
C4252 vdd.n2012 gnd 0.007974f
C4253 vdd.n2013 gnd 0.009907f
C4254 vdd.n2015 gnd 0.009907f
C4255 vdd.n2016 gnd 0.009907f
C4256 vdd.n2017 gnd 0.007974f
C4257 vdd.n2018 gnd 0.007974f
C4258 vdd.n2019 gnd 0.007974f
C4259 vdd.n2020 gnd 0.009907f
C4260 vdd.n2022 gnd 0.009907f
C4261 vdd.n2023 gnd 0.009907f
C4262 vdd.n2024 gnd 0.007974f
C4263 vdd.n2025 gnd 0.007974f
C4264 vdd.n2026 gnd 0.007974f
C4265 vdd.n2027 gnd 0.009907f
C4266 vdd.n2029 gnd 0.009907f
C4267 vdd.n2030 gnd 0.009907f
C4268 vdd.n2031 gnd 0.007974f
C4269 vdd.n2032 gnd 0.009907f
C4270 vdd.n2033 gnd 0.009907f
C4271 vdd.n2034 gnd 0.009907f
C4272 vdd.n2035 gnd 0.016267f
C4273 vdd.n2036 gnd 0.005422f
C4274 vdd.n2037 gnd 0.007974f
C4275 vdd.n2038 gnd 0.009907f
C4276 vdd.n2040 gnd 0.009907f
C4277 vdd.n2041 gnd 0.009907f
C4278 vdd.n2042 gnd 0.007974f
C4279 vdd.n2043 gnd 0.007974f
C4280 vdd.n2044 gnd 0.007974f
C4281 vdd.n2045 gnd 0.009907f
C4282 vdd.n2047 gnd 0.009907f
C4283 vdd.n2048 gnd 0.009907f
C4284 vdd.n2049 gnd 0.007974f
C4285 vdd.n2050 gnd 0.007974f
C4286 vdd.n2051 gnd 0.007974f
C4287 vdd.n2052 gnd 0.009907f
C4288 vdd.n2054 gnd 0.009907f
C4289 vdd.n2055 gnd 0.009907f
C4290 vdd.n2056 gnd 0.007974f
C4291 vdd.n2057 gnd 0.007974f
C4292 vdd.n2058 gnd 0.007974f
C4293 vdd.n2059 gnd 0.009907f
C4294 vdd.n2061 gnd 0.009907f
C4295 vdd.n2062 gnd 0.009907f
C4296 vdd.n2063 gnd 0.007974f
C4297 vdd.n2064 gnd 0.007974f
C4298 vdd.n2065 gnd 0.007974f
C4299 vdd.n2066 gnd 0.009907f
C4300 vdd.n2068 gnd 0.009907f
C4301 vdd.n2069 gnd 0.009907f
C4302 vdd.n2070 gnd 0.007974f
C4303 vdd.n2071 gnd 0.009907f
C4304 vdd.n2072 gnd 0.009907f
C4305 vdd.n2073 gnd 0.009907f
C4306 vdd.n2074 gnd 0.016267f
C4307 vdd.n2075 gnd 0.006658f
C4308 vdd.n2076 gnd 0.007974f
C4309 vdd.n2077 gnd 0.009907f
C4310 vdd.n2079 gnd 0.009907f
C4311 vdd.n2080 gnd 0.009907f
C4312 vdd.n2081 gnd 0.007974f
C4313 vdd.n2082 gnd 0.007974f
C4314 vdd.n2083 gnd 0.007974f
C4315 vdd.n2084 gnd 0.009907f
C4316 vdd.n2086 gnd 0.009907f
C4317 vdd.n2087 gnd 0.009907f
C4318 vdd.n2088 gnd 0.007974f
C4319 vdd.n2089 gnd 0.007974f
C4320 vdd.n2090 gnd 0.007974f
C4321 vdd.n2091 gnd 0.009907f
C4322 vdd.n2093 gnd 0.009907f
C4323 vdd.n2094 gnd 0.009907f
C4324 vdd.n2096 gnd 0.009907f
C4325 vdd.n2097 gnd 0.007974f
C4326 vdd.n2098 gnd 0.00634f
C4327 vdd.n2099 gnd 0.901205f
C4328 vdd.n2101 gnd 0.007974f
C4329 vdd.n2102 gnd 0.007974f
C4330 vdd.n2103 gnd 0.009907f
C4331 vdd.n2105 gnd 0.009907f
C4332 vdd.n2106 gnd 0.009907f
C4333 vdd.n2107 gnd 0.007974f
C4334 vdd.n2108 gnd 0.006618f
C4335 vdd.n2109 gnd 0.022714f
C4336 vdd.n2110 gnd 0.02256f
C4337 vdd.n2111 gnd 0.006618f
C4338 vdd.n2112 gnd 0.02256f
C4339 vdd.n2113 gnd 1.33641f
C4340 vdd.n2114 gnd 0.02256f
C4341 vdd.n2115 gnd 0.022714f
C4342 vdd.n2116 gnd 0.003788f
C4343 vdd.t54 gnd 0.12188f
C4344 vdd.t53 gnd 0.130256f
C4345 vdd.t51 gnd 0.159174f
C4346 vdd.n2117 gnd 0.204038f
C4347 vdd.n2118 gnd 0.171429f
C4348 vdd.n2119 gnd 0.01228f
C4349 vdd.n2120 gnd 0.004186f
C4350 vdd.n2121 gnd 0.00852f
C4351 vdd.n2122 gnd 0.901205f
C4352 vdd.n2123 gnd 0.035445f
C4353 vdd.n2124 gnd 0.006737f
C4354 vdd.n2125 gnd 0.006737f
C4355 vdd.n2126 gnd 0.006737f
C4356 vdd.n2127 gnd 0.006737f
C4357 vdd.n2128 gnd 0.006737f
C4358 vdd.n2129 gnd 0.006737f
C4359 vdd.n2130 gnd 0.006737f
C4360 vdd.n2131 gnd 0.006737f
C4361 vdd.n2133 gnd 0.006737f
C4362 vdd.n2135 gnd 0.006737f
C4363 vdd.n2136 gnd 0.006737f
C4364 vdd.n2137 gnd 0.006737f
C4365 vdd.n2138 gnd 0.006737f
C4366 vdd.n2139 gnd 0.006737f
C4367 vdd.n2141 gnd 0.006737f
C4368 vdd.n2143 gnd 0.006737f
C4369 vdd.n2144 gnd 0.006737f
C4370 vdd.n2145 gnd 0.006737f
C4371 vdd.n2146 gnd 0.006737f
C4372 vdd.n2147 gnd 0.006737f
C4373 vdd.n2149 gnd 0.006737f
C4374 vdd.n2151 gnd 0.006737f
C4375 vdd.n2152 gnd 0.006737f
C4376 vdd.n2153 gnd 0.006737f
C4377 vdd.n2154 gnd 0.006737f
C4378 vdd.n2155 gnd 0.006737f
C4379 vdd.n2157 gnd 0.006737f
C4380 vdd.n2159 gnd 0.006737f
C4381 vdd.n2160 gnd 0.006737f
C4382 vdd.n2161 gnd 0.006737f
C4383 vdd.n2162 gnd 0.006737f
C4384 vdd.n2163 gnd 0.006737f
C4385 vdd.n2165 gnd 0.006737f
C4386 vdd.n2167 gnd 0.006737f
C4387 vdd.n2168 gnd 0.006737f
C4388 vdd.n2169 gnd 0.006737f
C4389 vdd.n2170 gnd 0.006737f
C4390 vdd.n2171 gnd 0.006737f
C4391 vdd.n2173 gnd 0.006737f
C4392 vdd.n2175 gnd 0.006737f
C4393 vdd.n2176 gnd 0.006737f
C4394 vdd.n2177 gnd 0.006737f
C4395 vdd.n2178 gnd 0.006737f
C4396 vdd.n2179 gnd 0.006737f
C4397 vdd.n2181 gnd 0.006737f
C4398 vdd.n2183 gnd 0.006737f
C4399 vdd.n2184 gnd 0.006737f
C4400 vdd.n2185 gnd 0.006737f
C4401 vdd.n2186 gnd 0.006737f
C4402 vdd.n2187 gnd 0.006737f
C4403 vdd.n2189 gnd 0.006737f
C4404 vdd.n2191 gnd 0.006737f
C4405 vdd.n2192 gnd 0.006737f
C4406 vdd.n2193 gnd 0.004904f
C4407 vdd.n2194 gnd 0.009628f
C4408 vdd.n2195 gnd 0.005201f
C4409 vdd.n2196 gnd 0.006737f
C4410 vdd.n2198 gnd 0.006737f
C4411 vdd.n2199 gnd 0.015527f
C4412 vdd.n2200 gnd 0.015527f
C4413 vdd.n2201 gnd 0.01459f
C4414 vdd.n2202 gnd 0.006737f
C4415 vdd.n2203 gnd 0.006737f
C4416 vdd.n2204 gnd 0.006737f
C4417 vdd.n2205 gnd 0.006737f
C4418 vdd.n2206 gnd 0.006737f
C4419 vdd.n2207 gnd 0.006737f
C4420 vdd.n2208 gnd 0.006737f
C4421 vdd.n2209 gnd 0.006737f
C4422 vdd.n2210 gnd 0.006737f
C4423 vdd.n2211 gnd 0.006737f
C4424 vdd.n2212 gnd 0.006737f
C4425 vdd.n2213 gnd 0.006737f
C4426 vdd.n2214 gnd 0.006737f
C4427 vdd.n2215 gnd 0.006737f
C4428 vdd.n2216 gnd 0.006737f
C4429 vdd.n2217 gnd 0.006737f
C4430 vdd.n2218 gnd 0.006737f
C4431 vdd.n2219 gnd 0.006737f
C4432 vdd.n2220 gnd 0.006737f
C4433 vdd.n2221 gnd 0.006737f
C4434 vdd.n2222 gnd 0.006737f
C4435 vdd.n2223 gnd 0.006737f
C4436 vdd.n2224 gnd 0.006737f
C4437 vdd.n2225 gnd 0.006737f
C4438 vdd.n2226 gnd 0.006737f
C4439 vdd.n2227 gnd 0.006737f
C4440 vdd.n2228 gnd 0.006737f
C4441 vdd.n2229 gnd 0.006737f
C4442 vdd.n2230 gnd 0.006737f
C4443 vdd.n2231 gnd 0.006737f
C4444 vdd.n2232 gnd 0.006737f
C4445 vdd.n2233 gnd 0.006737f
C4446 vdd.n2234 gnd 0.006737f
C4447 vdd.n2235 gnd 0.006737f
C4448 vdd.n2236 gnd 0.006737f
C4449 vdd.n2237 gnd 0.006737f
C4450 vdd.n2238 gnd 0.006737f
C4451 vdd.n2239 gnd 0.006737f
C4452 vdd.n2240 gnd 0.006737f
C4453 vdd.n2241 gnd 0.006737f
C4454 vdd.n2242 gnd 0.006737f
C4455 vdd.n2243 gnd 0.006737f
C4456 vdd.n2244 gnd 0.006737f
C4457 vdd.n2245 gnd 0.006737f
C4458 vdd.n2246 gnd 0.006737f
C4459 vdd.n2247 gnd 0.006737f
C4460 vdd.n2248 gnd 0.006737f
C4461 vdd.n2249 gnd 0.006737f
C4462 vdd.n2250 gnd 0.006737f
C4463 vdd.n2251 gnd 0.410034f
C4464 vdd.n2252 gnd 0.006737f
C4465 vdd.n2253 gnd 0.006737f
C4466 vdd.n2254 gnd 0.006737f
C4467 vdd.n2255 gnd 0.006737f
C4468 vdd.n2256 gnd 0.006737f
C4469 vdd.n2257 gnd 0.006737f
C4470 vdd.n2258 gnd 0.006737f
C4471 vdd.n2259 gnd 0.006737f
C4472 vdd.n2260 gnd 0.006737f
C4473 vdd.n2261 gnd 0.006737f
C4474 vdd.n2262 gnd 0.006737f
C4475 vdd.n2263 gnd 0.622645f
C4476 vdd.n2264 gnd 0.006737f
C4477 vdd.n2265 gnd 0.006737f
C4478 vdd.n2266 gnd 0.006737f
C4479 vdd.n2267 gnd 0.006737f
C4480 vdd.n2268 gnd 0.006737f
C4481 vdd.n2269 gnd 0.006737f
C4482 vdd.n2270 gnd 0.006737f
C4483 vdd.n2271 gnd 0.006737f
C4484 vdd.n2272 gnd 0.006737f
C4485 vdd.n2273 gnd 0.006737f
C4486 vdd.n2274 gnd 0.006737f
C4487 vdd.n2275 gnd 0.217672f
C4488 vdd.n2276 gnd 0.006737f
C4489 vdd.n2277 gnd 0.006737f
C4490 vdd.n2278 gnd 0.006737f
C4491 vdd.n2279 gnd 0.006737f
C4492 vdd.n2280 gnd 0.006737f
C4493 vdd.n2281 gnd 0.006737f
C4494 vdd.n2282 gnd 0.006737f
C4495 vdd.n2283 gnd 0.006737f
C4496 vdd.n2284 gnd 0.006737f
C4497 vdd.n2285 gnd 0.006737f
C4498 vdd.n2286 gnd 0.006737f
C4499 vdd.n2287 gnd 0.006737f
C4500 vdd.n2288 gnd 0.006737f
C4501 vdd.n2289 gnd 0.006737f
C4502 vdd.n2290 gnd 0.006737f
C4503 vdd.n2291 gnd 0.006737f
C4504 vdd.n2292 gnd 0.006737f
C4505 vdd.n2293 gnd 0.006737f
C4506 vdd.n2294 gnd 0.006737f
C4507 vdd.n2295 gnd 0.006737f
C4508 vdd.n2296 gnd 0.006737f
C4509 vdd.n2297 gnd 0.006737f
C4510 vdd.n2298 gnd 0.006737f
C4511 vdd.n2299 gnd 0.006737f
C4512 vdd.n2300 gnd 0.006737f
C4513 vdd.n2301 gnd 0.006737f
C4514 vdd.n2302 gnd 0.006737f
C4515 vdd.n2303 gnd 0.006737f
C4516 vdd.n2304 gnd 0.006737f
C4517 vdd.n2305 gnd 0.006737f
C4518 vdd.n2306 gnd 0.006737f
C4519 vdd.n2307 gnd 0.006737f
C4520 vdd.n2308 gnd 0.006737f
C4521 vdd.n2309 gnd 0.006737f
C4522 vdd.n2310 gnd 0.006737f
C4523 vdd.n2311 gnd 0.01459f
C4524 vdd.n2312 gnd 0.015527f
C4525 vdd.n2313 gnd 0.015527f
C4526 vdd.n2315 gnd 0.006737f
C4527 vdd.n2317 gnd 0.006737f
C4528 vdd.n2318 gnd 0.005201f
C4529 vdd.n2319 gnd 0.009628f
C4530 vdd.n2320 gnd 0.004904f
C4531 vdd.n2321 gnd 0.006737f
C4532 vdd.n2322 gnd 0.006737f
C4533 vdd.n2324 gnd 0.006737f
C4534 vdd.n2326 gnd 0.006737f
C4535 vdd.n2327 gnd 0.006737f
C4536 vdd.n2328 gnd 0.006737f
C4537 vdd.n2329 gnd 0.006737f
C4538 vdd.n2330 gnd 0.006737f
C4539 vdd.n2332 gnd 0.006737f
C4540 vdd.n2334 gnd 0.006737f
C4541 vdd.n2335 gnd 0.006737f
C4542 vdd.n2336 gnd 0.006737f
C4543 vdd.n2337 gnd 0.006737f
C4544 vdd.n2338 gnd 0.006737f
C4545 vdd.n2340 gnd 0.006737f
C4546 vdd.n2342 gnd 0.006737f
C4547 vdd.n2343 gnd 0.006737f
C4548 vdd.n2344 gnd 0.006737f
C4549 vdd.n2345 gnd 0.006737f
C4550 vdd.n2346 gnd 0.006737f
C4551 vdd.n2348 gnd 0.006737f
C4552 vdd.n2350 gnd 0.006737f
C4553 vdd.n2351 gnd 0.006737f
C4554 vdd.n2352 gnd 0.006737f
C4555 vdd.n2353 gnd 0.006737f
C4556 vdd.n2354 gnd 0.006737f
C4557 vdd.n2356 gnd 0.006737f
C4558 vdd.n2358 gnd 0.006737f
C4559 vdd.n2359 gnd 0.006737f
C4560 vdd.n2360 gnd 0.006737f
C4561 vdd.n2361 gnd 0.006737f
C4562 vdd.n2362 gnd 0.006737f
C4563 vdd.n2364 gnd 0.006737f
C4564 vdd.n2366 gnd 0.006737f
C4565 vdd.n2367 gnd 0.006737f
C4566 vdd.n2368 gnd 0.006737f
C4567 vdd.n2369 gnd 0.006737f
C4568 vdd.n2370 gnd 0.006737f
C4569 vdd.n2372 gnd 0.006737f
C4570 vdd.n2373 gnd 0.006737f
C4571 vdd.n2374 gnd 0.006737f
C4572 vdd.n2375 gnd 0.006737f
C4573 vdd.n2376 gnd 0.006737f
C4574 vdd.n2377 gnd 0.006737f
C4575 vdd.n2379 gnd 0.006737f
C4576 vdd.n2380 gnd 0.006737f
C4577 vdd.n2381 gnd 0.015527f
C4578 vdd.n2382 gnd 0.01459f
C4579 vdd.n2383 gnd 0.01459f
C4580 vdd.n2384 gnd 0.951684f
C4581 vdd.n2385 gnd 0.01459f
C4582 vdd.n2386 gnd 0.01459f
C4583 vdd.n2387 gnd 0.006737f
C4584 vdd.n2388 gnd 0.006737f
C4585 vdd.n2389 gnd 0.006737f
C4586 vdd.n2390 gnd 0.47078f
C4587 vdd.n2391 gnd 0.006737f
C4588 vdd.n2392 gnd 0.006737f
C4589 vdd.n2393 gnd 0.006737f
C4590 vdd.n2394 gnd 0.006737f
C4591 vdd.n2395 gnd 0.006737f
C4592 vdd.n2396 gnd 0.688453f
C4593 vdd.n2397 gnd 0.006737f
C4594 vdd.n2398 gnd 0.006737f
C4595 vdd.n2399 gnd 0.006737f
C4596 vdd.n2400 gnd 0.006737f
C4597 vdd.n2401 gnd 0.006737f
C4598 vdd.n2402 gnd 0.688453f
C4599 vdd.n2403 gnd 0.006737f
C4600 vdd.n2404 gnd 0.006737f
C4601 vdd.n2405 gnd 0.006737f
C4602 vdd.n2406 gnd 0.006737f
C4603 vdd.n2407 gnd 0.006737f
C4604 vdd.n2408 gnd 0.349288f
C4605 vdd.n2409 gnd 0.006737f
C4606 vdd.n2410 gnd 0.006737f
C4607 vdd.n2411 gnd 0.006737f
C4608 vdd.n2412 gnd 0.006737f
C4609 vdd.n2413 gnd 0.006737f
C4610 vdd.n2414 gnd 0.501153f
C4611 vdd.n2415 gnd 0.006737f
C4612 vdd.n2416 gnd 0.006737f
C4613 vdd.n2417 gnd 0.006737f
C4614 vdd.n2418 gnd 0.006737f
C4615 vdd.n2419 gnd 0.006737f
C4616 vdd.n2420 gnd 0.653017f
C4617 vdd.n2421 gnd 0.006737f
C4618 vdd.n2422 gnd 0.006737f
C4619 vdd.n2423 gnd 0.006737f
C4620 vdd.n2424 gnd 0.006737f
C4621 vdd.n2425 gnd 0.006737f
C4622 vdd.n2426 gnd 0.688453f
C4623 vdd.n2427 gnd 0.006737f
C4624 vdd.n2428 gnd 0.006737f
C4625 vdd.n2429 gnd 0.006737f
C4626 vdd.n2430 gnd 0.006737f
C4627 vdd.n2431 gnd 0.006737f
C4628 vdd.n2432 gnd 0.572023f
C4629 vdd.n2433 gnd 0.006737f
C4630 vdd.n2434 gnd 0.006737f
C4631 vdd.n2435 gnd 0.005548f
C4632 vdd.n2436 gnd 0.019515f
C4633 vdd.n2437 gnd 0.004557f
C4634 vdd.n2438 gnd 0.006737f
C4635 vdd.n2439 gnd 0.420159f
C4636 vdd.n2440 gnd 0.006737f
C4637 vdd.n2441 gnd 0.006737f
C4638 vdd.n2442 gnd 0.006737f
C4639 vdd.n2443 gnd 0.006737f
C4640 vdd.n2444 gnd 0.006737f
C4641 vdd.n2445 gnd 0.420159f
C4642 vdd.n2446 gnd 0.006737f
C4643 vdd.n2447 gnd 0.006737f
C4644 vdd.n2448 gnd 0.006737f
C4645 vdd.n2449 gnd 0.006737f
C4646 vdd.n2450 gnd 0.006737f
C4647 vdd.n2451 gnd 0.572023f
C4648 vdd.n2452 gnd 0.006737f
C4649 vdd.n2453 gnd 0.006737f
C4650 vdd.n2454 gnd 0.006737f
C4651 vdd.n2455 gnd 0.006737f
C4652 vdd.n2456 gnd 0.006737f
C4653 vdd.n2457 gnd 0.587209f
C4654 vdd.n2458 gnd 0.006737f
C4655 vdd.n2459 gnd 0.006737f
C4656 vdd.n2460 gnd 0.006737f
C4657 vdd.n2461 gnd 0.006737f
C4658 vdd.n2462 gnd 0.006737f
C4659 vdd.n2463 gnd 0.435345f
C4660 vdd.n2464 gnd 0.006737f
C4661 vdd.n2465 gnd 0.006737f
C4662 vdd.n2466 gnd 0.006737f
C4663 vdd.n2467 gnd 0.006737f
C4664 vdd.n2468 gnd 0.006737f
C4665 vdd.n2469 gnd 0.217672f
C4666 vdd.n2470 gnd 0.006737f
C4667 vdd.n2471 gnd 0.006737f
C4668 vdd.n2472 gnd 0.006737f
C4669 vdd.n2473 gnd 0.006737f
C4670 vdd.n2474 gnd 0.006737f
C4671 vdd.n2475 gnd 0.217672f
C4672 vdd.n2476 gnd 0.006737f
C4673 vdd.n2477 gnd 0.006737f
C4674 vdd.n2478 gnd 0.006737f
C4675 vdd.n2479 gnd 0.006737f
C4676 vdd.n2480 gnd 0.006737f
C4677 vdd.n2481 gnd 0.688453f
C4678 vdd.n2482 gnd 0.006737f
C4679 vdd.n2483 gnd 0.006737f
C4680 vdd.n2484 gnd 0.006737f
C4681 vdd.n2485 gnd 0.006737f
C4682 vdd.n2486 gnd 0.006737f
C4683 vdd.n2487 gnd 0.006737f
C4684 vdd.n2488 gnd 0.006737f
C4685 vdd.n2489 gnd 0.496091f
C4686 vdd.n2490 gnd 0.006737f
C4687 vdd.n2491 gnd 0.006737f
C4688 vdd.n2492 gnd 0.006737f
C4689 vdd.n2493 gnd 0.006737f
C4690 vdd.n2494 gnd 0.006737f
C4691 vdd.n2495 gnd 0.006737f
C4692 vdd.n2496 gnd 0.430283f
C4693 vdd.n2497 gnd 0.006737f
C4694 vdd.n2498 gnd 0.006737f
C4695 vdd.n2499 gnd 0.006737f
C4696 vdd.n2500 gnd 0.015444f
C4697 vdd.n2501 gnd 0.014673f
C4698 vdd.n2502 gnd 0.006737f
C4699 vdd.n2503 gnd 0.006737f
C4700 vdd.n2504 gnd 0.005201f
C4701 vdd.n2505 gnd 0.006737f
C4702 vdd.n2506 gnd 0.006737f
C4703 vdd.n2507 gnd 0.004904f
C4704 vdd.n2508 gnd 0.006737f
C4705 vdd.n2509 gnd 0.006737f
C4706 vdd.n2510 gnd 0.006737f
C4707 vdd.n2511 gnd 0.006737f
C4708 vdd.n2512 gnd 0.006737f
C4709 vdd.n2513 gnd 0.006737f
C4710 vdd.n2514 gnd 0.006737f
C4711 vdd.n2515 gnd 0.006737f
C4712 vdd.n2516 gnd 0.006737f
C4713 vdd.n2517 gnd 0.006737f
C4714 vdd.n2518 gnd 0.006737f
C4715 vdd.n2519 gnd 0.006737f
C4716 vdd.n2520 gnd 0.006737f
C4717 vdd.n2521 gnd 0.006737f
C4718 vdd.n2522 gnd 0.006737f
C4719 vdd.n2523 gnd 0.006737f
C4720 vdd.n2524 gnd 0.006737f
C4721 vdd.n2525 gnd 0.006737f
C4722 vdd.n2526 gnd 0.006737f
C4723 vdd.n2527 gnd 0.006737f
C4724 vdd.n2528 gnd 0.006737f
C4725 vdd.n2529 gnd 0.006737f
C4726 vdd.n2530 gnd 0.006737f
C4727 vdd.n2531 gnd 0.006737f
C4728 vdd.n2532 gnd 0.006737f
C4729 vdd.n2533 gnd 0.006737f
C4730 vdd.n2534 gnd 0.006737f
C4731 vdd.n2535 gnd 0.006737f
C4732 vdd.n2536 gnd 0.006737f
C4733 vdd.n2537 gnd 0.006737f
C4734 vdd.n2538 gnd 0.006737f
C4735 vdd.n2539 gnd 0.006737f
C4736 vdd.n2540 gnd 0.006737f
C4737 vdd.n2541 gnd 0.006737f
C4738 vdd.n2542 gnd 0.006737f
C4739 vdd.n2543 gnd 0.006737f
C4740 vdd.n2544 gnd 0.006737f
C4741 vdd.n2545 gnd 0.006737f
C4742 vdd.n2546 gnd 0.006737f
C4743 vdd.n2547 gnd 0.006737f
C4744 vdd.n2548 gnd 0.006737f
C4745 vdd.n2549 gnd 0.006737f
C4746 vdd.n2550 gnd 0.006737f
C4747 vdd.n2551 gnd 0.006737f
C4748 vdd.n2552 gnd 0.006737f
C4749 vdd.n2553 gnd 0.006737f
C4750 vdd.n2554 gnd 0.006737f
C4751 vdd.n2555 gnd 0.006737f
C4752 vdd.n2556 gnd 0.006737f
C4753 vdd.n2557 gnd 0.006737f
C4754 vdd.n2558 gnd 0.006737f
C4755 vdd.n2559 gnd 0.006737f
C4756 vdd.n2560 gnd 0.006737f
C4757 vdd.n2561 gnd 0.006737f
C4758 vdd.n2562 gnd 0.006737f
C4759 vdd.n2563 gnd 0.006737f
C4760 vdd.n2564 gnd 0.006737f
C4761 vdd.n2565 gnd 0.006737f
C4762 vdd.n2566 gnd 0.006737f
C4763 vdd.n2567 gnd 0.006737f
C4764 vdd.n2568 gnd 0.015527f
C4765 vdd.n2569 gnd 0.01459f
C4766 vdd.n2570 gnd 0.01459f
C4767 vdd.n2571 gnd 0.79982f
C4768 vdd.n2572 gnd 0.01459f
C4769 vdd.n2573 gnd 0.015527f
C4770 vdd.n2574 gnd 0.014673f
C4771 vdd.n2575 gnd 0.006737f
C4772 vdd.n2576 gnd 0.006737f
C4773 vdd.n2577 gnd 0.006737f
C4774 vdd.n2578 gnd 0.005201f
C4775 vdd.n2579 gnd 0.009628f
C4776 vdd.n2580 gnd 0.004904f
C4777 vdd.n2581 gnd 0.006737f
C4778 vdd.n2582 gnd 0.006737f
C4779 vdd.n2583 gnd 0.006737f
C4780 vdd.n2584 gnd 0.006737f
C4781 vdd.n2585 gnd 0.006737f
C4782 vdd.n2586 gnd 0.006737f
C4783 vdd.n2587 gnd 0.006737f
C4784 vdd.n2588 gnd 0.006737f
C4785 vdd.n2589 gnd 0.006737f
C4786 vdd.n2590 gnd 0.006737f
C4787 vdd.n2591 gnd 0.006737f
C4788 vdd.n2592 gnd 0.006737f
C4789 vdd.n2593 gnd 0.006737f
C4790 vdd.n2594 gnd 0.006737f
C4791 vdd.n2595 gnd 0.006737f
C4792 vdd.n2596 gnd 0.006737f
C4793 vdd.n2597 gnd 0.006737f
C4794 vdd.n2598 gnd 0.006737f
C4795 vdd.n2599 gnd 0.006737f
C4796 vdd.n2600 gnd 0.006737f
C4797 vdd.n2601 gnd 0.006737f
C4798 vdd.n2602 gnd 0.006737f
C4799 vdd.n2603 gnd 0.006737f
C4800 vdd.n2604 gnd 0.006737f
C4801 vdd.n2605 gnd 0.006737f
C4802 vdd.n2606 gnd 0.006737f
C4803 vdd.n2607 gnd 0.006737f
C4804 vdd.n2608 gnd 0.006737f
C4805 vdd.n2609 gnd 0.006737f
C4806 vdd.n2610 gnd 0.006737f
C4807 vdd.n2611 gnd 0.006737f
C4808 vdd.n2612 gnd 0.006737f
C4809 vdd.n2613 gnd 0.006737f
C4810 vdd.n2614 gnd 0.006737f
C4811 vdd.n2615 gnd 0.006737f
C4812 vdd.n2616 gnd 0.006737f
C4813 vdd.n2617 gnd 0.006737f
C4814 vdd.n2618 gnd 0.006737f
C4815 vdd.n2619 gnd 0.006737f
C4816 vdd.n2620 gnd 0.006737f
C4817 vdd.n2621 gnd 0.006737f
C4818 vdd.n2622 gnd 0.006737f
C4819 vdd.n2623 gnd 0.006737f
C4820 vdd.n2624 gnd 0.006737f
C4821 vdd.n2625 gnd 0.006737f
C4822 vdd.n2626 gnd 0.006737f
C4823 vdd.n2627 gnd 0.006737f
C4824 vdd.n2628 gnd 0.006737f
C4825 vdd.n2629 gnd 0.006737f
C4826 vdd.n2630 gnd 0.006737f
C4827 vdd.n2631 gnd 0.006737f
C4828 vdd.n2632 gnd 0.006737f
C4829 vdd.n2633 gnd 0.006737f
C4830 vdd.n2634 gnd 0.006737f
C4831 vdd.n2635 gnd 0.006737f
C4832 vdd.n2636 gnd 0.006737f
C4833 vdd.n2637 gnd 0.006737f
C4834 vdd.n2638 gnd 0.006737f
C4835 vdd.n2639 gnd 0.006737f
C4836 vdd.n2640 gnd 0.006737f
C4837 vdd.n2641 gnd 0.015527f
C4838 vdd.n2642 gnd 0.015527f
C4839 vdd.n2643 gnd 0.840317f
C4840 vdd.t155 gnd 2.98667f
C4841 vdd.t142 gnd 2.98667f
C4842 vdd.n2677 gnd 0.006737f
C4843 vdd.t90 gnd 0.272227f
C4844 vdd.t91 gnd 0.278658f
C4845 vdd.t89 gnd 0.17772f
C4846 vdd.n2678 gnd 0.096048f
C4847 vdd.n2679 gnd 0.054481f
C4848 vdd.n2680 gnd 0.009628f
C4849 vdd.n2681 gnd 0.006737f
C4850 vdd.n2682 gnd 0.006737f
C4851 vdd.n2683 gnd 0.006737f
C4852 vdd.n2684 gnd 0.006737f
C4853 vdd.n2685 gnd 0.006737f
C4854 vdd.n2686 gnd 0.006737f
C4855 vdd.n2687 gnd 0.006737f
C4856 vdd.n2688 gnd 0.006737f
C4857 vdd.n2689 gnd 0.006737f
C4858 vdd.n2690 gnd 0.006737f
C4859 vdd.n2691 gnd 0.006737f
C4860 vdd.n2692 gnd 0.006737f
C4861 vdd.n2693 gnd 0.006737f
C4862 vdd.n2694 gnd 0.006737f
C4863 vdd.n2695 gnd 0.006737f
C4864 vdd.n2696 gnd 0.006737f
C4865 vdd.n2697 gnd 0.006737f
C4866 vdd.n2698 gnd 0.006737f
C4867 vdd.n2699 gnd 0.006737f
C4868 vdd.n2700 gnd 0.006737f
C4869 vdd.n2701 gnd 0.006737f
C4870 vdd.n2702 gnd 0.006737f
C4871 vdd.n2703 gnd 0.006737f
C4872 vdd.n2704 gnd 0.006737f
C4873 vdd.n2705 gnd 0.006737f
C4874 vdd.n2706 gnd 0.006737f
C4875 vdd.n2707 gnd 0.006737f
C4876 vdd.n2708 gnd 0.006737f
C4877 vdd.n2709 gnd 0.006737f
C4878 vdd.n2710 gnd 0.006737f
C4879 vdd.n2711 gnd 0.006737f
C4880 vdd.n2712 gnd 0.006737f
C4881 vdd.n2713 gnd 0.006737f
C4882 vdd.n2714 gnd 0.006737f
C4883 vdd.n2715 gnd 0.006737f
C4884 vdd.n2716 gnd 0.006737f
C4885 vdd.n2717 gnd 0.006737f
C4886 vdd.n2718 gnd 0.006737f
C4887 vdd.n2719 gnd 0.006737f
C4888 vdd.n2720 gnd 0.006737f
C4889 vdd.n2721 gnd 0.006737f
C4890 vdd.n2722 gnd 0.006737f
C4891 vdd.n2723 gnd 0.006737f
C4892 vdd.n2724 gnd 0.006737f
C4893 vdd.n2725 gnd 0.006737f
C4894 vdd.n2726 gnd 0.006737f
C4895 vdd.n2727 gnd 0.006737f
C4896 vdd.n2728 gnd 0.006737f
C4897 vdd.n2729 gnd 0.006737f
C4898 vdd.n2730 gnd 0.006737f
C4899 vdd.n2731 gnd 0.006737f
C4900 vdd.n2732 gnd 0.006737f
C4901 vdd.n2733 gnd 0.006737f
C4902 vdd.n2734 gnd 0.006737f
C4903 vdd.n2735 gnd 0.006737f
C4904 vdd.n2736 gnd 0.006737f
C4905 vdd.n2737 gnd 0.006737f
C4906 vdd.n2738 gnd 0.006737f
C4907 vdd.n2739 gnd 0.006737f
C4908 vdd.n2740 gnd 0.006737f
C4909 vdd.n2741 gnd 0.004904f
C4910 vdd.n2742 gnd 0.006737f
C4911 vdd.n2743 gnd 0.006737f
C4912 vdd.n2744 gnd 0.005201f
C4913 vdd.n2745 gnd 0.006737f
C4914 vdd.n2746 gnd 0.006737f
C4915 vdd.t77 gnd 0.272227f
C4916 vdd.t78 gnd 0.278658f
C4917 vdd.t75 gnd 0.17772f
C4918 vdd.n2747 gnd 0.096048f
C4919 vdd.n2748 gnd 0.054481f
C4920 vdd.n2749 gnd 0.006737f
C4921 vdd.n2750 gnd 0.006737f
C4922 vdd.n2751 gnd 0.006737f
C4923 vdd.n2752 gnd 0.006737f
C4924 vdd.n2753 gnd 0.006737f
C4925 vdd.n2754 gnd 0.006737f
C4926 vdd.n2755 gnd 0.006737f
C4927 vdd.n2756 gnd 0.006737f
C4928 vdd.n2757 gnd 0.006737f
C4929 vdd.n2758 gnd 0.006737f
C4930 vdd.n2759 gnd 0.006737f
C4931 vdd.n2760 gnd 0.006737f
C4932 vdd.n2761 gnd 0.006737f
C4933 vdd.n2762 gnd 0.006737f
C4934 vdd.n2763 gnd 0.006737f
C4935 vdd.n2764 gnd 0.006737f
C4936 vdd.n2765 gnd 0.006737f
C4937 vdd.n2766 gnd 0.006737f
C4938 vdd.n2767 gnd 0.006737f
C4939 vdd.n2768 gnd 0.006737f
C4940 vdd.n2769 gnd 0.006737f
C4941 vdd.n2770 gnd 0.006737f
C4942 vdd.n2771 gnd 0.006737f
C4943 vdd.n2772 gnd 0.006737f
C4944 vdd.n2773 gnd 0.006737f
C4945 vdd.n2774 gnd 0.006737f
C4946 vdd.n2775 gnd 0.006737f
C4947 vdd.n2776 gnd 0.006737f
C4948 vdd.n2777 gnd 0.006737f
C4949 vdd.n2778 gnd 0.006737f
C4950 vdd.n2779 gnd 0.006737f
C4951 vdd.n2780 gnd 0.006737f
C4952 vdd.n2781 gnd 0.006737f
C4953 vdd.n2782 gnd 0.006737f
C4954 vdd.n2783 gnd 0.006737f
C4955 vdd.n2784 gnd 0.006737f
C4956 vdd.n2785 gnd 0.006737f
C4957 vdd.n2786 gnd 0.006737f
C4958 vdd.n2787 gnd 0.006737f
C4959 vdd.n2788 gnd 0.006737f
C4960 vdd.n2789 gnd 0.006737f
C4961 vdd.n2790 gnd 0.006737f
C4962 vdd.n2791 gnd 0.006737f
C4963 vdd.n2792 gnd 0.006737f
C4964 vdd.n2793 gnd 0.006737f
C4965 vdd.n2794 gnd 0.006737f
C4966 vdd.n2795 gnd 0.006737f
C4967 vdd.n2796 gnd 0.006737f
C4968 vdd.n2797 gnd 0.006737f
C4969 vdd.n2798 gnd 0.006737f
C4970 vdd.n2799 gnd 0.006737f
C4971 vdd.n2800 gnd 0.006737f
C4972 vdd.n2801 gnd 0.006737f
C4973 vdd.n2802 gnd 0.006737f
C4974 vdd.n2803 gnd 0.006737f
C4975 vdd.n2804 gnd 0.006737f
C4976 vdd.n2805 gnd 0.006737f
C4977 vdd.n2806 gnd 0.004904f
C4978 vdd.n2807 gnd 0.009628f
C4979 vdd.n2808 gnd 0.005201f
C4980 vdd.n2809 gnd 0.006737f
C4981 vdd.n2810 gnd 0.006737f
C4982 vdd.n2811 gnd 0.006737f
C4983 vdd.n2812 gnd 0.015527f
C4984 vdd.n2813 gnd 0.015527f
C4985 vdd.n2814 gnd 0.01459f
C4986 vdd.n2815 gnd 0.006737f
C4987 vdd.n2816 gnd 0.006737f
C4988 vdd.n2817 gnd 0.006737f
C4989 vdd.n2818 gnd 0.006737f
C4990 vdd.n2819 gnd 0.006737f
C4991 vdd.n2820 gnd 0.006737f
C4992 vdd.n2821 gnd 0.006737f
C4993 vdd.n2822 gnd 0.006737f
C4994 vdd.n2823 gnd 0.006737f
C4995 vdd.n2824 gnd 0.006737f
C4996 vdd.n2825 gnd 0.006737f
C4997 vdd.n2826 gnd 0.006737f
C4998 vdd.n2827 gnd 0.006737f
C4999 vdd.n2828 gnd 0.006737f
C5000 vdd.n2829 gnd 0.006737f
C5001 vdd.n2830 gnd 0.006737f
C5002 vdd.n2831 gnd 0.006737f
C5003 vdd.n2832 gnd 0.006737f
C5004 vdd.n2833 gnd 0.006737f
C5005 vdd.n2834 gnd 0.006737f
C5006 vdd.n2835 gnd 0.006737f
C5007 vdd.n2836 gnd 0.006737f
C5008 vdd.n2837 gnd 0.006737f
C5009 vdd.n2838 gnd 0.006737f
C5010 vdd.n2839 gnd 0.006737f
C5011 vdd.n2840 gnd 0.006737f
C5012 vdd.n2841 gnd 0.006737f
C5013 vdd.n2842 gnd 0.006737f
C5014 vdd.n2843 gnd 0.006737f
C5015 vdd.n2844 gnd 0.006737f
C5016 vdd.n2845 gnd 0.006737f
C5017 vdd.n2846 gnd 0.006737f
C5018 vdd.n2847 gnd 0.006737f
C5019 vdd.n2848 gnd 0.006737f
C5020 vdd.n2849 gnd 0.006737f
C5021 vdd.n2850 gnd 0.006737f
C5022 vdd.n2851 gnd 0.006737f
C5023 vdd.n2852 gnd 0.006737f
C5024 vdd.n2853 gnd 0.006737f
C5025 vdd.n2854 gnd 0.006737f
C5026 vdd.n2855 gnd 0.006737f
C5027 vdd.n2856 gnd 0.006737f
C5028 vdd.n2857 gnd 0.006737f
C5029 vdd.n2858 gnd 0.006737f
C5030 vdd.n2859 gnd 0.006737f
C5031 vdd.n2860 gnd 0.006737f
C5032 vdd.n2861 gnd 0.006737f
C5033 vdd.n2862 gnd 0.006737f
C5034 vdd.n2863 gnd 0.006737f
C5035 vdd.n2864 gnd 0.006737f
C5036 vdd.n2865 gnd 0.006737f
C5037 vdd.n2866 gnd 0.006737f
C5038 vdd.n2867 gnd 0.006737f
C5039 vdd.n2868 gnd 0.006737f
C5040 vdd.n2869 gnd 0.006737f
C5041 vdd.n2870 gnd 0.006737f
C5042 vdd.n2871 gnd 0.006737f
C5043 vdd.n2872 gnd 0.006737f
C5044 vdd.n2873 gnd 0.006737f
C5045 vdd.n2874 gnd 0.006737f
C5046 vdd.n2875 gnd 0.006737f
C5047 vdd.n2876 gnd 0.006737f
C5048 vdd.n2877 gnd 0.006737f
C5049 vdd.n2878 gnd 0.006737f
C5050 vdd.n2879 gnd 0.006737f
C5051 vdd.n2880 gnd 0.006737f
C5052 vdd.n2881 gnd 0.006737f
C5053 vdd.n2882 gnd 0.006737f
C5054 vdd.n2883 gnd 0.006737f
C5055 vdd.n2884 gnd 0.006737f
C5056 vdd.n2885 gnd 0.006737f
C5057 vdd.n2886 gnd 0.006737f
C5058 vdd.n2887 gnd 0.006737f
C5059 vdd.n2888 gnd 0.006737f
C5060 vdd.n2889 gnd 0.006737f
C5061 vdd.n2890 gnd 0.006737f
C5062 vdd.n2891 gnd 0.006737f
C5063 vdd.n2892 gnd 0.006737f
C5064 vdd.n2893 gnd 0.006737f
C5065 vdd.n2894 gnd 0.217672f
C5066 vdd.n2895 gnd 0.006737f
C5067 vdd.n2896 gnd 0.006737f
C5068 vdd.n2897 gnd 0.006737f
C5069 vdd.n2898 gnd 0.006737f
C5070 vdd.n2899 gnd 0.006737f
C5071 vdd.n2900 gnd 0.006737f
C5072 vdd.n2901 gnd 0.006737f
C5073 vdd.n2902 gnd 0.006737f
C5074 vdd.n2903 gnd 0.006737f
C5075 vdd.n2904 gnd 0.006737f
C5076 vdd.n2905 gnd 0.006737f
C5077 vdd.n2906 gnd 0.622645f
C5078 vdd.n2907 gnd 0.006737f
C5079 vdd.n2908 gnd 0.006737f
C5080 vdd.n2909 gnd 0.006737f
C5081 vdd.n2910 gnd 0.006737f
C5082 vdd.n2911 gnd 0.006737f
C5083 vdd.n2912 gnd 0.006737f
C5084 vdd.n2913 gnd 0.006737f
C5085 vdd.n2914 gnd 0.006737f
C5086 vdd.n2915 gnd 0.006737f
C5087 vdd.n2916 gnd 0.006737f
C5088 vdd.n2917 gnd 0.006737f
C5089 vdd.n2918 gnd 0.410034f
C5090 vdd.n2919 gnd 0.006737f
C5091 vdd.n2920 gnd 0.006737f
C5092 vdd.n2921 gnd 0.006737f
C5093 vdd.n2922 gnd 0.006737f
C5094 vdd.n2923 gnd 0.006737f
C5095 vdd.n2924 gnd 0.01459f
C5096 vdd.n2925 gnd 0.015527f
C5097 vdd.n2926 gnd 0.015527f
C5098 vdd.n2927 gnd 0.840317f
C5099 vdd.n2929 gnd 0.006737f
C5100 vdd.n2930 gnd 0.006737f
C5101 vdd.n2931 gnd 0.015527f
C5102 vdd.n2932 gnd 0.01459f
C5103 vdd.n2933 gnd 0.01459f
C5104 vdd.n2934 gnd 0.79982f
C5105 vdd.n2935 gnd 0.01459f
C5106 vdd.n2936 gnd 0.01459f
C5107 vdd.n2937 gnd 0.006737f
C5108 vdd.n2938 gnd 0.006737f
C5109 vdd.n2939 gnd 0.006737f
C5110 vdd.n2940 gnd 0.430283f
C5111 vdd.n2941 gnd 0.006737f
C5112 vdd.n2942 gnd 0.006737f
C5113 vdd.n2943 gnd 0.006737f
C5114 vdd.n2944 gnd 0.006737f
C5115 vdd.n2945 gnd 0.006737f
C5116 vdd.n2946 gnd 0.496091f
C5117 vdd.n2947 gnd 0.006737f
C5118 vdd.n2948 gnd 0.006737f
C5119 vdd.n2949 gnd 0.006737f
C5120 vdd.n2950 gnd 0.006737f
C5121 vdd.n2951 gnd 0.006737f
C5122 vdd.n2952 gnd 0.688453f
C5123 vdd.n2953 gnd 0.006737f
C5124 vdd.n2954 gnd 0.006737f
C5125 vdd.n2955 gnd 0.006737f
C5126 vdd.n2956 gnd 0.006737f
C5127 vdd.n2957 gnd 0.006737f
C5128 vdd.n2958 gnd 0.217672f
C5129 vdd.n2959 gnd 0.006737f
C5130 vdd.n2960 gnd 0.006737f
C5131 vdd.n2961 gnd 0.006737f
C5132 vdd.n2962 gnd 0.006737f
C5133 vdd.n2963 gnd 0.006737f
C5134 vdd.n2964 gnd 0.217672f
C5135 vdd.n2965 gnd 0.006737f
C5136 vdd.n2966 gnd 0.006737f
C5137 vdd.n2967 gnd 0.006737f
C5138 vdd.n2968 gnd 0.006737f
C5139 vdd.n2969 gnd 0.006737f
C5140 vdd.n2970 gnd 0.435345f
C5141 vdd.n2971 gnd 0.006737f
C5142 vdd.n2972 gnd 0.006737f
C5143 vdd.n2973 gnd 0.006737f
C5144 vdd.n2974 gnd 0.006737f
C5145 vdd.n2975 gnd 0.006737f
C5146 vdd.n2976 gnd 0.587209f
C5147 vdd.n2977 gnd 0.006737f
C5148 vdd.n2978 gnd 0.006737f
C5149 vdd.n2979 gnd 0.006737f
C5150 vdd.n2980 gnd 0.006737f
C5151 vdd.n2981 gnd 0.006737f
C5152 vdd.n2982 gnd 0.572023f
C5153 vdd.n2983 gnd 0.006737f
C5154 vdd.n2984 gnd 0.006737f
C5155 vdd.n2985 gnd 0.006737f
C5156 vdd.n2986 gnd 0.006737f
C5157 vdd.n2987 gnd 0.006737f
C5158 vdd.n2988 gnd 0.420159f
C5159 vdd.n2989 gnd 0.006737f
C5160 vdd.n2990 gnd 0.006737f
C5161 vdd.n2991 gnd 0.006737f
C5162 vdd.n2992 gnd 0.006737f
C5163 vdd.n2993 gnd 0.006737f
C5164 vdd.n2994 gnd 0.420159f
C5165 vdd.n2995 gnd 0.006737f
C5166 vdd.n2996 gnd 0.004557f
C5167 vdd.n2997 gnd 0.019515f
C5168 vdd.n2998 gnd 0.005548f
C5169 vdd.n2999 gnd 0.006737f
C5170 vdd.n3000 gnd 0.006737f
C5171 vdd.n3001 gnd 0.572023f
C5172 vdd.n3002 gnd 0.006737f
C5173 vdd.n3003 gnd 0.006737f
C5174 vdd.n3004 gnd 0.006737f
C5175 vdd.n3005 gnd 0.006737f
C5176 vdd.n3006 gnd 0.006737f
C5177 vdd.n3007 gnd 0.688453f
C5178 vdd.n3008 gnd 0.006737f
C5179 vdd.n3009 gnd 0.006737f
C5180 vdd.n3010 gnd 0.006737f
C5181 vdd.n3011 gnd 0.006737f
C5182 vdd.n3012 gnd 0.006737f
C5183 vdd.n3013 gnd 0.653017f
C5184 vdd.n3014 gnd 0.006737f
C5185 vdd.n3015 gnd 0.006737f
C5186 vdd.n3016 gnd 0.006737f
C5187 vdd.n3017 gnd 0.006737f
C5188 vdd.n3018 gnd 0.006737f
C5189 vdd.n3019 gnd 0.501153f
C5190 vdd.n3020 gnd 0.006737f
C5191 vdd.n3021 gnd 0.006737f
C5192 vdd.n3022 gnd 0.006737f
C5193 vdd.n3023 gnd 0.006737f
C5194 vdd.n3024 gnd 0.006737f
C5195 vdd.n3025 gnd 0.349288f
C5196 vdd.n3026 gnd 0.006737f
C5197 vdd.n3027 gnd 0.006737f
C5198 vdd.n3028 gnd 0.006737f
C5199 vdd.n3029 gnd 0.006737f
C5200 vdd.n3030 gnd 0.006737f
C5201 vdd.n3031 gnd 0.688453f
C5202 vdd.n3032 gnd 0.006737f
C5203 vdd.n3033 gnd 0.006737f
C5204 vdd.n3034 gnd 0.006737f
C5205 vdd.n3035 gnd 0.006737f
C5206 vdd.n3036 gnd 0.006737f
C5207 vdd.n3037 gnd 0.006737f
C5208 vdd.n3039 gnd 0.006737f
C5209 vdd.n3040 gnd 0.006737f
C5210 vdd.n3042 gnd 0.006737f
C5211 vdd.n3043 gnd 0.006737f
C5212 vdd.n3046 gnd 0.006737f
C5213 vdd.n3047 gnd 0.006737f
C5214 vdd.n3048 gnd 0.006737f
C5215 vdd.n3049 gnd 0.006737f
C5216 vdd.n3051 gnd 0.006737f
C5217 vdd.n3052 gnd 0.006737f
C5218 vdd.n3053 gnd 0.006737f
C5219 vdd.n3054 gnd 0.006737f
C5220 vdd.n3055 gnd 0.006737f
C5221 vdd.n3056 gnd 0.006737f
C5222 vdd.n3058 gnd 0.006737f
C5223 vdd.n3059 gnd 0.006737f
C5224 vdd.n3060 gnd 0.006737f
C5225 vdd.n3061 gnd 0.006737f
C5226 vdd.n3062 gnd 0.006737f
C5227 vdd.n3063 gnd 0.006737f
C5228 vdd.n3065 gnd 0.006737f
C5229 vdd.n3066 gnd 0.006737f
C5230 vdd.n3067 gnd 0.006737f
C5231 vdd.n3068 gnd 0.006737f
C5232 vdd.n3069 gnd 0.006737f
C5233 vdd.n3070 gnd 0.006737f
C5234 vdd.n3072 gnd 0.006737f
C5235 vdd.n3073 gnd 0.015527f
C5236 vdd.n3074 gnd 0.015527f
C5237 vdd.n3075 gnd 0.01459f
C5238 vdd.n3076 gnd 0.006737f
C5239 vdd.n3077 gnd 0.006737f
C5240 vdd.n3078 gnd 0.006737f
C5241 vdd.n3079 gnd 0.006737f
C5242 vdd.n3080 gnd 0.006737f
C5243 vdd.n3081 gnd 0.006737f
C5244 vdd.n3082 gnd 0.688453f
C5245 vdd.n3083 gnd 0.006737f
C5246 vdd.n3084 gnd 0.006737f
C5247 vdd.n3085 gnd 0.006737f
C5248 vdd.n3086 gnd 0.006737f
C5249 vdd.n3087 gnd 0.006737f
C5250 vdd.n3088 gnd 0.47078f
C5251 vdd.n3089 gnd 0.006737f
C5252 vdd.n3090 gnd 0.006737f
C5253 vdd.n3091 gnd 0.006737f
C5254 vdd.n3092 gnd 0.015444f
C5255 vdd.n3094 gnd 0.015527f
C5256 vdd.n3095 gnd 0.014673f
C5257 vdd.n3096 gnd 0.006737f
C5258 vdd.n3097 gnd 0.005201f
C5259 vdd.n3098 gnd 0.006737f
C5260 vdd.n3100 gnd 0.006737f
C5261 vdd.n3101 gnd 0.006737f
C5262 vdd.n3102 gnd 0.006737f
C5263 vdd.n3103 gnd 0.006737f
C5264 vdd.n3104 gnd 0.006737f
C5265 vdd.n3105 gnd 0.006737f
C5266 vdd.n3107 gnd 0.006737f
C5267 vdd.n3108 gnd 0.006737f
C5268 vdd.n3109 gnd 0.006737f
C5269 vdd.n3110 gnd 0.006737f
C5270 vdd.n3111 gnd 0.006737f
C5271 vdd.n3112 gnd 0.006737f
C5272 vdd.n3114 gnd 0.006737f
C5273 vdd.n3115 gnd 0.006737f
C5274 vdd.n3116 gnd 0.006737f
C5275 vdd.n3117 gnd 0.006737f
C5276 vdd.n3118 gnd 0.006737f
C5277 vdd.n3119 gnd 0.006737f
C5278 vdd.n3121 gnd 0.006737f
C5279 vdd.n3122 gnd 0.006737f
C5280 vdd.n3123 gnd 0.006737f
C5281 vdd.n3124 gnd 0.905028f
C5282 vdd.n3125 gnd 0.031622f
C5283 vdd.n3126 gnd 0.006737f
C5284 vdd.n3127 gnd 0.006737f
C5285 vdd.n3129 gnd 0.006737f
C5286 vdd.n3130 gnd 0.006737f
C5287 vdd.n3131 gnd 0.006737f
C5288 vdd.n3132 gnd 0.006737f
C5289 vdd.n3133 gnd 0.006737f
C5290 vdd.n3134 gnd 0.006737f
C5291 vdd.n3136 gnd 0.006737f
C5292 vdd.n3137 gnd 0.006737f
C5293 vdd.n3138 gnd 0.006737f
C5294 vdd.n3139 gnd 0.006737f
C5295 vdd.n3140 gnd 0.006737f
C5296 vdd.n3141 gnd 0.006737f
C5297 vdd.n3143 gnd 0.006737f
C5298 vdd.n3144 gnd 0.006737f
C5299 vdd.n3145 gnd 0.006737f
C5300 vdd.n3146 gnd 0.006737f
C5301 vdd.n3147 gnd 0.006737f
C5302 vdd.n3148 gnd 0.006737f
C5303 vdd.n3150 gnd 0.006737f
C5304 vdd.n3151 gnd 0.006737f
C5305 vdd.n3153 gnd 0.006737f
C5306 vdd.n3154 gnd 0.006737f
C5307 vdd.n3155 gnd 0.015527f
C5308 vdd.n3156 gnd 0.01459f
C5309 vdd.n3157 gnd 0.01459f
C5310 vdd.n3158 gnd 0.951684f
C5311 vdd.n3159 gnd 0.01459f
C5312 vdd.n3160 gnd 0.015527f
C5313 vdd.n3161 gnd 0.014673f
C5314 vdd.n3162 gnd 0.006737f
C5315 vdd.n3163 gnd 0.005201f
C5316 vdd.n3164 gnd 0.006737f
C5317 vdd.n3166 gnd 0.006737f
C5318 vdd.n3167 gnd 0.006737f
C5319 vdd.n3168 gnd 0.006737f
C5320 vdd.n3169 gnd 0.006737f
C5321 vdd.n3170 gnd 0.006737f
C5322 vdd.n3171 gnd 0.006737f
C5323 vdd.n3173 gnd 0.006737f
C5324 vdd.n3174 gnd 0.006737f
C5325 vdd.n3175 gnd 0.006737f
C5326 vdd.n3176 gnd 0.006737f
C5327 vdd.n3177 gnd 0.006737f
C5328 vdd.n3178 gnd 0.006737f
C5329 vdd.n3180 gnd 0.006737f
C5330 vdd.n3181 gnd 0.006737f
C5331 vdd.n3182 gnd 0.006737f
C5332 vdd.n3183 gnd 0.006737f
C5333 vdd.n3184 gnd 0.006737f
C5334 vdd.n3185 gnd 0.006737f
C5335 vdd.n3187 gnd 0.006737f
C5336 vdd.n3188 gnd 0.006737f
C5337 vdd.n3190 gnd 0.006737f
C5338 vdd.n3191 gnd 0.031622f
C5339 vdd.n3192 gnd 0.905028f
C5340 vdd.n3193 gnd 0.00852f
C5341 vdd.n3194 gnd 0.003788f
C5342 vdd.t49 gnd 0.12188f
C5343 vdd.t50 gnd 0.130256f
C5344 vdd.t48 gnd 0.159174f
C5345 vdd.n3195 gnd 0.204038f
C5346 vdd.n3196 gnd 0.171429f
C5347 vdd.n3197 gnd 0.01228f
C5348 vdd.n3198 gnd 0.009907f
C5349 vdd.n3199 gnd 0.004186f
C5350 vdd.n3200 gnd 0.007974f
C5351 vdd.n3201 gnd 0.009907f
C5352 vdd.n3202 gnd 0.009907f
C5353 vdd.n3203 gnd 0.007974f
C5354 vdd.n3204 gnd 0.007974f
C5355 vdd.n3205 gnd 0.009907f
C5356 vdd.n3207 gnd 0.009907f
C5357 vdd.n3208 gnd 0.007974f
C5358 vdd.n3209 gnd 0.007974f
C5359 vdd.n3210 gnd 0.007974f
C5360 vdd.n3211 gnd 0.009907f
C5361 vdd.n3213 gnd 0.009907f
C5362 vdd.n3215 gnd 0.009907f
C5363 vdd.n3216 gnd 0.007974f
C5364 vdd.n3217 gnd 0.007974f
C5365 vdd.n3218 gnd 0.007974f
C5366 vdd.n3219 gnd 0.009907f
C5367 vdd.n3221 gnd 0.009907f
C5368 vdd.n3223 gnd 0.009907f
C5369 vdd.n3224 gnd 0.007974f
C5370 vdd.n3225 gnd 0.007974f
C5371 vdd.n3226 gnd 0.007974f
C5372 vdd.n3227 gnd 0.009907f
C5373 vdd.n3229 gnd 0.009907f
C5374 vdd.n3230 gnd 0.009907f
C5375 vdd.n3231 gnd 0.007974f
C5376 vdd.n3232 gnd 0.007974f
C5377 vdd.n3233 gnd 0.009907f
C5378 vdd.n3234 gnd 0.009907f
C5379 vdd.n3236 gnd 0.009907f
C5380 vdd.n3237 gnd 0.007974f
C5381 vdd.n3238 gnd 0.009907f
C5382 vdd.n3239 gnd 0.009907f
C5383 vdd.n3240 gnd 0.009907f
C5384 vdd.n3241 gnd 0.016267f
C5385 vdd.n3242 gnd 0.005422f
C5386 vdd.n3243 gnd 0.009907f
C5387 vdd.n3245 gnd 0.009907f
C5388 vdd.n3247 gnd 0.009907f
C5389 vdd.n3248 gnd 0.007974f
C5390 vdd.n3249 gnd 0.007974f
C5391 vdd.n3250 gnd 0.007974f
C5392 vdd.n3251 gnd 0.009907f
C5393 vdd.n3253 gnd 0.009907f
C5394 vdd.n3255 gnd 0.009907f
C5395 vdd.n3256 gnd 0.007974f
C5396 vdd.n3257 gnd 0.007974f
C5397 vdd.n3258 gnd 0.007974f
C5398 vdd.n3259 gnd 0.009907f
C5399 vdd.n3261 gnd 0.009907f
C5400 vdd.n3263 gnd 0.009907f
C5401 vdd.n3264 gnd 0.007974f
C5402 vdd.n3265 gnd 0.007974f
C5403 vdd.n3266 gnd 0.007974f
C5404 vdd.n3267 gnd 0.009907f
C5405 vdd.n3269 gnd 0.009907f
C5406 vdd.n3271 gnd 0.009907f
C5407 vdd.n3272 gnd 0.007974f
C5408 vdd.n3273 gnd 0.007974f
C5409 vdd.n3274 gnd 0.007974f
C5410 vdd.n3275 gnd 0.009907f
C5411 vdd.n3277 gnd 0.009907f
C5412 vdd.n3279 gnd 0.009907f
C5413 vdd.n3280 gnd 0.007974f
C5414 vdd.n3281 gnd 0.007974f
C5415 vdd.n3282 gnd 0.006658f
C5416 vdd.n3283 gnd 0.009907f
C5417 vdd.n3285 gnd 0.009907f
C5418 vdd.n3287 gnd 0.009907f
C5419 vdd.n3288 gnd 0.006658f
C5420 vdd.n3289 gnd 0.007974f
C5421 vdd.n3290 gnd 0.007974f
C5422 vdd.n3291 gnd 0.009907f
C5423 vdd.n3293 gnd 0.009907f
C5424 vdd.n3295 gnd 0.009907f
C5425 vdd.n3296 gnd 0.007974f
C5426 vdd.n3297 gnd 0.007974f
C5427 vdd.n3298 gnd 0.007974f
C5428 vdd.n3299 gnd 0.009907f
C5429 vdd.n3301 gnd 0.009907f
C5430 vdd.n3303 gnd 0.009907f
C5431 vdd.n3304 gnd 0.007974f
C5432 vdd.n3305 gnd 0.007974f
C5433 vdd.n3306 gnd 0.007974f
C5434 vdd.n3307 gnd 0.009907f
C5435 vdd.n3309 gnd 0.009907f
C5436 vdd.n3310 gnd 0.009907f
C5437 vdd.n3311 gnd 0.007974f
C5438 vdd.n3312 gnd 0.007974f
C5439 vdd.n3313 gnd 0.009907f
C5440 vdd.n3314 gnd 0.009907f
C5441 vdd.n3315 gnd 0.007974f
C5442 vdd.n3316 gnd 0.007974f
C5443 vdd.n3317 gnd 0.009907f
C5444 vdd.n3318 gnd 0.009907f
C5445 vdd.n3320 gnd 0.009907f
C5446 vdd.n3321 gnd 0.007974f
C5447 vdd.n3322 gnd 0.006618f
C5448 vdd.n3323 gnd 0.022714f
C5449 vdd.n3324 gnd 0.02256f
C5450 vdd.n3325 gnd 0.006618f
C5451 vdd.n3326 gnd 0.02256f
C5452 vdd.n3327 gnd 1.33641f
C5453 vdd.n3328 gnd 0.02256f
C5454 vdd.n3329 gnd 0.006618f
C5455 vdd.n3330 gnd 0.02256f
C5456 vdd.n3331 gnd 0.009907f
C5457 vdd.n3332 gnd 0.009907f
C5458 vdd.n3333 gnd 0.007974f
C5459 vdd.n3334 gnd 0.009907f
C5460 vdd.n3335 gnd 0.956746f
C5461 vdd.n3336 gnd 0.009907f
C5462 vdd.n3337 gnd 0.007974f
C5463 vdd.n3338 gnd 0.009907f
C5464 vdd.n3339 gnd 0.009907f
C5465 vdd.n3340 gnd 0.009907f
C5466 vdd.n3341 gnd 0.007974f
C5467 vdd.n3342 gnd 0.009907f
C5468 vdd.n3343 gnd 0.987119f
C5469 vdd.n3344 gnd 0.009907f
C5470 vdd.n3345 gnd 0.007974f
C5471 vdd.n3346 gnd 0.009907f
C5472 vdd.n3347 gnd 0.009907f
C5473 vdd.n3348 gnd 0.009907f
C5474 vdd.n3349 gnd 0.007974f
C5475 vdd.n3350 gnd 0.009907f
C5476 vdd.t121 gnd 0.506215f
C5477 vdd.n3351 gnd 0.815006f
C5478 vdd.n3352 gnd 0.009907f
C5479 vdd.n3353 gnd 0.007974f
C5480 vdd.n3354 gnd 0.009907f
C5481 vdd.n3355 gnd 0.009907f
C5482 vdd.n3356 gnd 0.009907f
C5483 vdd.n3357 gnd 0.007974f
C5484 vdd.n3358 gnd 0.009907f
C5485 vdd.n3359 gnd 0.642893f
C5486 vdd.n3360 gnd 0.009907f
C5487 vdd.n3361 gnd 0.007974f
C5488 vdd.n3362 gnd 0.009907f
C5489 vdd.n3363 gnd 0.009907f
C5490 vdd.n3364 gnd 0.009907f
C5491 vdd.n3365 gnd 0.007974f
C5492 vdd.n3366 gnd 0.009907f
C5493 vdd.n3367 gnd 0.804882f
C5494 vdd.n3368 gnd 0.54165f
C5495 vdd.n3369 gnd 0.009907f
C5496 vdd.n3370 gnd 0.007974f
C5497 vdd.n3371 gnd 0.009907f
C5498 vdd.n3372 gnd 0.009907f
C5499 vdd.n3373 gnd 0.009907f
C5500 vdd.n3374 gnd 0.007974f
C5501 vdd.n3375 gnd 0.009907f
C5502 vdd.n3376 gnd 0.713763f
C5503 vdd.n3377 gnd 0.009907f
C5504 vdd.n3378 gnd 0.007974f
C5505 vdd.n3379 gnd 0.009907f
C5506 vdd.n3380 gnd 0.009907f
C5507 vdd.n3381 gnd 0.009907f
C5508 vdd.n3382 gnd 0.009907f
C5509 vdd.n3383 gnd 0.009907f
C5510 vdd.n3384 gnd 0.007974f
C5511 vdd.n3385 gnd 0.007974f
C5512 vdd.n3386 gnd 0.009907f
C5513 vdd.t119 gnd 0.506215f
C5514 vdd.n3387 gnd 0.840317f
C5515 vdd.n3388 gnd 0.009907f
C5516 vdd.n3389 gnd 0.007974f
C5517 vdd.n3390 gnd 0.009907f
C5518 vdd.n3391 gnd 0.009907f
C5519 vdd.n3392 gnd 0.009907f
C5520 vdd.n3393 gnd 0.007974f
C5521 vdd.n3394 gnd 0.009907f
C5522 vdd.n3395 gnd 0.794758f
C5523 vdd.n3396 gnd 0.009907f
C5524 vdd.n3397 gnd 0.009907f
C5525 vdd.n3398 gnd 0.007974f
C5526 vdd.n3399 gnd 0.007974f
C5527 vdd.n3400 gnd 0.007974f
C5528 vdd.n3401 gnd 0.009907f
C5529 vdd.n3402 gnd 0.009907f
C5530 vdd.n3403 gnd 0.009907f
C5531 vdd.n3404 gnd 0.009907f
C5532 vdd.n3405 gnd 0.007974f
C5533 vdd.n3406 gnd 0.007974f
C5534 vdd.n3407 gnd 0.007974f
C5535 vdd.n3408 gnd 0.009907f
C5536 vdd.n3409 gnd 0.009907f
C5537 vdd.n3410 gnd 0.009907f
C5538 vdd.n3411 gnd 0.009907f
C5539 vdd.n3412 gnd 0.007974f
C5540 vdd.n3413 gnd 0.007974f
C5541 vdd.n3414 gnd 0.007974f
C5542 vdd.n3415 gnd 0.009907f
C5543 vdd.n3416 gnd 0.009907f
C5544 vdd.n3417 gnd 0.009907f
C5545 vdd.n3418 gnd 0.840317f
C5546 vdd.n3419 gnd 0.009907f
C5547 vdd.n3420 gnd 0.007974f
C5548 vdd.n3421 gnd 0.007974f
C5549 vdd.n3422 gnd 0.007974f
C5550 vdd.n3423 gnd 0.009907f
C5551 vdd.n3424 gnd 0.009907f
C5552 vdd.n3425 gnd 0.009907f
C5553 vdd.n3426 gnd 0.009907f
C5554 vdd.n3427 gnd 0.007974f
C5555 vdd.n3428 gnd 0.007974f
C5556 vdd.n3429 gnd 0.006618f
C5557 vdd.n3430 gnd 0.02256f
C5558 vdd.n3431 gnd 0.022714f
C5559 vdd.n3432 gnd 0.003788f
C5560 vdd.n3433 gnd 0.022714f
C5561 vdd.n3435 gnd 2.23747f
C5562 vdd.n3436 gnd 1.33641f
C5563 vdd.n3437 gnd 0.663142f
C5564 vdd.n3438 gnd 0.009907f
C5565 vdd.n3439 gnd 0.007974f
C5566 vdd.n3440 gnd 0.007974f
C5567 vdd.n3441 gnd 0.007974f
C5568 vdd.n3442 gnd 0.009907f
C5569 vdd.n3443 gnd 1.01243f
C5570 vdd.n3444 gnd 1.01243f
C5571 vdd.n3445 gnd 0.582147f
C5572 vdd.n3446 gnd 0.009907f
C5573 vdd.n3447 gnd 0.007974f
C5574 vdd.n3448 gnd 0.007974f
C5575 vdd.n3449 gnd 0.007974f
C5576 vdd.n3450 gnd 0.009907f
C5577 vdd.n3451 gnd 0.602396f
C5578 vdd.n3452 gnd 0.744136f
C5579 vdd.t19 gnd 0.506215f
C5580 vdd.n3453 gnd 0.774509f
C5581 vdd.n3454 gnd 0.009907f
C5582 vdd.n3455 gnd 0.007974f
C5583 vdd.n3456 gnd 0.007974f
C5584 vdd.n3457 gnd 0.007974f
C5585 vdd.n3458 gnd 0.009907f
C5586 vdd.n3459 gnd 0.840317f
C5587 vdd.t124 gnd 0.506215f
C5588 vdd.n3460 gnd 0.61252f
C5589 vdd.n3461 gnd 0.734012f
C5590 vdd.n3462 gnd 0.009907f
C5591 vdd.n3463 gnd 0.007974f
C5592 vdd.n3464 gnd 0.007974f
C5593 vdd.n3465 gnd 0.007974f
C5594 vdd.n3466 gnd 0.009907f
C5595 vdd.n3467 gnd 0.561899f
C5596 vdd.t8 gnd 0.506215f
C5597 vdd.n3468 gnd 0.840317f
C5598 vdd.t213 gnd 0.506215f
C5599 vdd.n3469 gnd 0.622645f
C5600 vdd.n3470 gnd 0.009907f
C5601 vdd.n3471 gnd 0.007974f
C5602 vdd.n3472 gnd 0.007614f
C5603 vdd.n3473 gnd 0.584342f
C5604 vdd.n3474 gnd 2.59845f
C5605 a_n2472_13878.t25 gnd 0.187389f
C5606 a_n2472_13878.t21 gnd 0.187389f
C5607 a_n2472_13878.t27 gnd 0.187389f
C5608 a_n2472_13878.n0 gnd 1.47796f
C5609 a_n2472_13878.t8 gnd 0.187389f
C5610 a_n2472_13878.t18 gnd 0.187389f
C5611 a_n2472_13878.n1 gnd 1.47552f
C5612 a_n2472_13878.n2 gnd 1.32632f
C5613 a_n2472_13878.t23 gnd 0.187389f
C5614 a_n2472_13878.t15 gnd 0.187389f
C5615 a_n2472_13878.n3 gnd 1.47709f
C5616 a_n2472_13878.t20 gnd 0.187389f
C5617 a_n2472_13878.t14 gnd 0.187389f
C5618 a_n2472_13878.n4 gnd 1.47552f
C5619 a_n2472_13878.n5 gnd 2.06176f
C5620 a_n2472_13878.t10 gnd 0.187389f
C5621 a_n2472_13878.t12 gnd 0.187389f
C5622 a_n2472_13878.n6 gnd 1.47552f
C5623 a_n2472_13878.n7 gnd 1.00568f
C5624 a_n2472_13878.t22 gnd 0.187389f
C5625 a_n2472_13878.t11 gnd 0.187389f
C5626 a_n2472_13878.n8 gnd 1.47552f
C5627 a_n2472_13878.n9 gnd 1.00568f
C5628 a_n2472_13878.t19 gnd 0.187389f
C5629 a_n2472_13878.t9 gnd 0.187389f
C5630 a_n2472_13878.n10 gnd 1.47552f
C5631 a_n2472_13878.n11 gnd 4.40118f
C5632 a_n2472_13878.t4 gnd 1.75461f
C5633 a_n2472_13878.t2 gnd 0.187389f
C5634 a_n2472_13878.t3 gnd 0.187389f
C5635 a_n2472_13878.n12 gnd 1.31997f
C5636 a_n2472_13878.n13 gnd 1.47487f
C5637 a_n2472_13878.t7 gnd 1.75112f
C5638 a_n2472_13878.n14 gnd 0.742173f
C5639 a_n2472_13878.t6 gnd 1.75112f
C5640 a_n2472_13878.n15 gnd 0.742173f
C5641 a_n2472_13878.t0 gnd 0.187389f
C5642 a_n2472_13878.t1 gnd 0.187389f
C5643 a_n2472_13878.n16 gnd 1.31997f
C5644 a_n2472_13878.n17 gnd 0.749361f
C5645 a_n2472_13878.t5 gnd 1.75112f
C5646 a_n2472_13878.n18 gnd 2.43496f
C5647 a_n2472_13878.n19 gnd 3.22551f
C5648 a_n2472_13878.t24 gnd 0.187389f
C5649 a_n2472_13878.t13 gnd 0.187389f
C5650 a_n2472_13878.n20 gnd 1.47552f
C5651 a_n2472_13878.n21 gnd 2.21835f
C5652 a_n2472_13878.t16 gnd 0.187389f
C5653 a_n2472_13878.t17 gnd 0.187389f
C5654 a_n2472_13878.n22 gnd 1.47552f
C5655 a_n2472_13878.n23 gnd 0.653766f
C5656 a_n2472_13878.n24 gnd 0.653763f
C5657 a_n2472_13878.n25 gnd 1.47553f
C5658 a_n2472_13878.t26 gnd 0.187389f
C5659 a_n2650_13878.n0 gnd 0.89022f
C5660 a_n2650_13878.n1 gnd 3.61027f
C5661 a_n2650_13878.n2 gnd 3.33797f
C5662 a_n2650_13878.n3 gnd 3.94237f
C5663 a_n2650_13878.n4 gnd 0.783099f
C5664 a_n2650_13878.n5 gnd 0.199822f
C5665 a_n2650_13878.n6 gnd 0.147172f
C5666 a_n2650_13878.n7 gnd 0.231308f
C5667 a_n2650_13878.n8 gnd 0.178659f
C5668 a_n2650_13878.n9 gnd 0.199822f
C5669 a_n2650_13878.n10 gnd 1.20992f
C5670 a_n2650_13878.n11 gnd 0.147172f
C5671 a_n2650_13878.n12 gnd 0.835748f
C5672 a_n2650_13878.n13 gnd 0.210597f
C5673 a_n2650_13878.n14 gnd 0.679581f
C5674 a_n2650_13878.n15 gnd 0.210597f
C5675 a_n2650_13878.n16 gnd 0.490668f
C5676 a_n2650_13878.n17 gnd 0.210597f
C5677 a_n2650_13878.n18 gnd 0.543317f
C5678 a_n2650_13878.n19 gnd 0.210597f
C5679 a_n2650_13878.n20 gnd 0.871815f
C5680 a_n2650_13878.n21 gnd 0.210597f
C5681 a_n2650_13878.n22 gnd 0.911906f
C5682 a_n2650_13878.n23 gnd 0.210597f
C5683 a_n2650_13878.n24 gnd 0.490668f
C5684 a_n2650_13878.n25 gnd 0.210597f
C5685 a_n2650_13878.n26 gnd 2.91769f
C5686 a_n2650_13878.n27 gnd 0.78318f
C5687 a_n2650_13878.n28 gnd 1.14968f
C5688 a_n2650_13878.n29 gnd 1.16828f
C5689 a_n2650_13878.n30 gnd 2.18252f
C5690 a_n2650_13878.n31 gnd 1.73382f
C5691 a_n2650_13878.n32 gnd 1.41042f
C5692 a_n2650_13878.n33 gnd 1.16827f
C5693 a_n2650_13878.n34 gnd 0.438019f
C5694 a_n2650_13878.n35 gnd 0.00845f
C5695 a_n2650_13878.n36 gnd 4.07e-19
C5696 a_n2650_13878.n38 gnd 0.008154f
C5697 a_n2650_13878.n39 gnd 0.011856f
C5698 a_n2650_13878.n40 gnd 0.278198f
C5699 a_n2650_13878.n41 gnd 0.00845f
C5700 a_n2650_13878.n42 gnd 4.07e-19
C5701 a_n2650_13878.n44 gnd 0.008154f
C5702 a_n2650_13878.n45 gnd 0.011856f
C5703 a_n2650_13878.n46 gnd 0.007844f
C5704 a_n2650_13878.n47 gnd 0.278198f
C5705 a_n2650_13878.n48 gnd 0.00845f
C5706 a_n2650_13878.n49 gnd 4.07e-19
C5707 a_n2650_13878.n51 gnd 0.008154f
C5708 a_n2650_13878.n52 gnd 0.011856f
C5709 a_n2650_13878.n53 gnd 0.007844f
C5710 a_n2650_13878.n54 gnd 0.278198f
C5711 a_n2650_13878.n55 gnd 0.00845f
C5712 a_n2650_13878.n56 gnd 4.07e-19
C5713 a_n2650_13878.n58 gnd 0.008154f
C5714 a_n2650_13878.n59 gnd 0.011856f
C5715 a_n2650_13878.n60 gnd 0.007844f
C5716 a_n2650_13878.n61 gnd 0.278198f
C5717 a_n2650_13878.n62 gnd 0.008154f
C5718 a_n2650_13878.n63 gnd 0.278198f
C5719 a_n2650_13878.n64 gnd 0.008154f
C5720 a_n2650_13878.n65 gnd 0.278198f
C5721 a_n2650_13878.n66 gnd 0.008154f
C5722 a_n2650_13878.n67 gnd 0.278198f
C5723 a_n2650_13878.n68 gnd 0.008154f
C5724 a_n2650_13878.n69 gnd 0.278198f
C5725 a_n2650_13878.n70 gnd 0.007844f
C5726 a_n2650_13878.t37 gnd 0.146072f
C5727 a_n2650_13878.t4 gnd 0.679457f
C5728 a_n2650_13878.t12 gnd 0.679457f
C5729 a_n2650_13878.t30 gnd 0.679457f
C5730 a_n2650_13878.n71 gnd 0.298598f
C5731 a_n2650_13878.t0 gnd 0.679457f
C5732 a_n2650_13878.t36 gnd 0.679457f
C5733 a_n2650_13878.t16 gnd 0.679457f
C5734 a_n2650_13878.n72 gnd 0.294939f
C5735 a_n2650_13878.t8 gnd 0.679457f
C5736 a_n2650_13878.t24 gnd 0.679457f
C5737 a_n2650_13878.t94 gnd 0.679457f
C5738 a_n2650_13878.t73 gnd 0.679457f
C5739 a_n2650_13878.t78 gnd 0.679457f
C5740 a_n2650_13878.n73 gnd 0.298598f
C5741 a_n2650_13878.t67 gnd 0.679457f
C5742 a_n2650_13878.t83 gnd 0.679457f
C5743 a_n2650_13878.t91 gnd 0.679457f
C5744 a_n2650_13878.n74 gnd 0.294939f
C5745 a_n2650_13878.t92 gnd 0.679457f
C5746 a_n2650_13878.t62 gnd 0.679457f
C5747 a_n2650_13878.t75 gnd 0.679457f
C5748 a_n2650_13878.n75 gnd 0.298717f
C5749 a_n2650_13878.t23 gnd 1.36775f
C5750 a_n2650_13878.t29 gnd 0.146072f
C5751 a_n2650_13878.t3 gnd 0.146072f
C5752 a_n2650_13878.n76 gnd 1.02893f
C5753 a_n2650_13878.t33 gnd 0.146072f
C5754 a_n2650_13878.t35 gnd 0.146072f
C5755 a_n2650_13878.n77 gnd 1.02893f
C5756 a_n2650_13878.t11 gnd 0.146072f
C5757 a_n2650_13878.t21 gnd 0.146072f
C5758 a_n2650_13878.n78 gnd 1.02893f
C5759 a_n2650_13878.t15 gnd 0.146072f
C5760 a_n2650_13878.t27 gnd 0.146072f
C5761 a_n2650_13878.n79 gnd 1.02893f
C5762 a_n2650_13878.t39 gnd 1.36502f
C5763 a_n2650_13878.t14 gnd 0.679457f
C5764 a_n2650_13878.n80 gnd 0.295192f
C5765 a_n2650_13878.t10 gnd 0.679457f
C5766 a_n2650_13878.t2 gnd 0.679457f
C5767 a_n2650_13878.n81 gnd 0.298598f
C5768 a_n2650_13878.t22 gnd 0.679457f
C5769 a_n2650_13878.t71 gnd 0.679457f
C5770 a_n2650_13878.n82 gnd 0.295192f
C5771 a_n2650_13878.t86 gnd 0.679457f
C5772 a_n2650_13878.t89 gnd 0.679457f
C5773 a_n2650_13878.n83 gnd 0.298598f
C5774 a_n2650_13878.t66 gnd 0.679457f
C5775 a_n2650_13878.n84 gnd 0.289583f
C5776 a_n2650_13878.t90 gnd 0.679457f
C5777 a_n2650_13878.n85 gnd 0.294614f
C5778 a_n2650_13878.t64 gnd 0.679457f
C5779 a_n2650_13878.n86 gnd 0.301285f
C5780 a_n2650_13878.t87 gnd 0.679457f
C5781 a_n2650_13878.n87 gnd 0.298732f
C5782 a_n2650_13878.n88 gnd 0.294939f
C5783 a_n2650_13878.t61 gnd 0.679457f
C5784 a_n2650_13878.n89 gnd 0.289745f
C5785 a_n2650_13878.t81 gnd 0.679457f
C5786 a_n2650_13878.n90 gnd 0.298717f
C5787 a_n2650_13878.t63 gnd 0.690842f
C5788 a_n2650_13878.n91 gnd 0.289583f
C5789 a_n2650_13878.t28 gnd 0.679457f
C5790 a_n2650_13878.n92 gnd 0.294614f
C5791 a_n2650_13878.t32 gnd 0.679457f
C5792 a_n2650_13878.n93 gnd 0.301285f
C5793 a_n2650_13878.t34 gnd 0.679457f
C5794 a_n2650_13878.n94 gnd 0.298732f
C5795 a_n2650_13878.n95 gnd 0.294939f
C5796 a_n2650_13878.t20 gnd 0.679457f
C5797 a_n2650_13878.n96 gnd 0.289745f
C5798 a_n2650_13878.t26 gnd 0.679457f
C5799 a_n2650_13878.n97 gnd 0.298717f
C5800 a_n2650_13878.t38 gnd 0.690842f
C5801 a_n2650_13878.n98 gnd 1.24181f
C5802 a_n2650_13878.t70 gnd 0.679457f
C5803 a_n2650_13878.n99 gnd 0.294939f
C5804 a_n2650_13878.t77 gnd 0.679457f
C5805 a_n2650_13878.n100 gnd 0.294939f
C5806 a_n2650_13878.t69 gnd 0.679457f
C5807 a_n2650_13878.n101 gnd 0.294939f
C5808 a_n2650_13878.t82 gnd 0.679457f
C5809 a_n2650_13878.n102 gnd 0.294939f
C5810 a_n2650_13878.t72 gnd 0.679457f
C5811 a_n2650_13878.n103 gnd 0.289583f
C5812 a_n2650_13878.t95 gnd 0.679457f
C5813 a_n2650_13878.n104 gnd 0.298732f
C5814 a_n2650_13878.t74 gnd 0.690842f
C5815 a_n2650_13878.t84 gnd 0.679457f
C5816 a_n2650_13878.n105 gnd 0.289583f
C5817 a_n2650_13878.t68 gnd 0.679457f
C5818 a_n2650_13878.n106 gnd 0.298732f
C5819 a_n2650_13878.t79 gnd 0.690842f
C5820 a_n2650_13878.t88 gnd 0.679457f
C5821 a_n2650_13878.n107 gnd 0.289583f
C5822 a_n2650_13878.t76 gnd 0.679457f
C5823 a_n2650_13878.n108 gnd 0.298732f
C5824 a_n2650_13878.t93 gnd 0.690842f
C5825 a_n2650_13878.t80 gnd 0.679457f
C5826 a_n2650_13878.n109 gnd 0.289583f
C5827 a_n2650_13878.t60 gnd 0.679457f
C5828 a_n2650_13878.n110 gnd 0.298732f
C5829 a_n2650_13878.t85 gnd 0.690842f
C5830 a_n2650_13878.n111 gnd 1.53361f
C5831 a_n2650_13878.t65 gnd 0.690842f
C5832 a_n2650_13878.n112 gnd 0.295192f
C5833 a_n2650_13878.n113 gnd 0.289745f
C5834 a_n2650_13878.n114 gnd 0.298732f
C5835 a_n2650_13878.n115 gnd 0.301285f
C5836 a_n2650_13878.n116 gnd 0.294614f
C5837 a_n2650_13878.n117 gnd 0.289583f
C5838 a_n2650_13878.t6 gnd 0.690842f
C5839 a_n2650_13878.t18 gnd 0.679457f
C5840 a_n2650_13878.n118 gnd 0.298717f
C5841 a_n2650_13878.t54 gnd 0.113612f
C5842 a_n2650_13878.t44 gnd 0.113612f
C5843 a_n2650_13878.n119 gnd 1.00687f
C5844 a_n2650_13878.t40 gnd 0.113612f
C5845 a_n2650_13878.t41 gnd 0.113612f
C5846 a_n2650_13878.n120 gnd 1.00391f
C5847 a_n2650_13878.t56 gnd 0.113612f
C5848 a_n2650_13878.t58 gnd 0.113612f
C5849 a_n2650_13878.n121 gnd 1.00391f
C5850 a_n2650_13878.t46 gnd 0.113612f
C5851 a_n2650_13878.t45 gnd 0.113612f
C5852 a_n2650_13878.n122 gnd 1.00687f
C5853 a_n2650_13878.t53 gnd 0.113612f
C5854 a_n2650_13878.t50 gnd 0.113612f
C5855 a_n2650_13878.n123 gnd 1.00391f
C5856 a_n2650_13878.t48 gnd 0.113612f
C5857 a_n2650_13878.t49 gnd 0.113612f
C5858 a_n2650_13878.n124 gnd 1.00391f
C5859 a_n2650_13878.t52 gnd 0.113612f
C5860 a_n2650_13878.t55 gnd 0.113612f
C5861 a_n2650_13878.n125 gnd 1.00391f
C5862 a_n2650_13878.t59 gnd 0.113612f
C5863 a_n2650_13878.t42 gnd 0.113612f
C5864 a_n2650_13878.n126 gnd 1.00391f
C5865 a_n2650_13878.t51 gnd 0.113612f
C5866 a_n2650_13878.t57 gnd 0.113612f
C5867 a_n2650_13878.n127 gnd 1.00687f
C5868 a_n2650_13878.t43 gnd 0.113612f
C5869 a_n2650_13878.t47 gnd 0.113612f
C5870 a_n2650_13878.n128 gnd 1.00391f
C5871 a_n2650_13878.n129 gnd 0.295192f
C5872 a_n2650_13878.n130 gnd 0.289745f
C5873 a_n2650_13878.n131 gnd 0.298732f
C5874 a_n2650_13878.n132 gnd 0.301285f
C5875 a_n2650_13878.n133 gnd 0.294614f
C5876 a_n2650_13878.n134 gnd 0.289583f
C5877 a_n2650_13878.n135 gnd 0.918226f
C5878 a_n2650_13878.t5 gnd 1.36502f
C5879 a_n2650_13878.t13 gnd 0.146072f
C5880 a_n2650_13878.t31 gnd 0.146072f
C5881 a_n2650_13878.n136 gnd 1.02893f
C5882 a_n2650_13878.t7 gnd 1.36775f
C5883 a_n2650_13878.t25 gnd 0.146072f
C5884 a_n2650_13878.t19 gnd 0.146072f
C5885 a_n2650_13878.n137 gnd 1.02893f
C5886 a_n2650_13878.t17 gnd 0.146072f
C5887 a_n2650_13878.t9 gnd 0.146072f
C5888 a_n2650_13878.n138 gnd 1.02893f
C5889 a_n2650_13878.n139 gnd 1.02894f
C5890 a_n2650_13878.t1 gnd 0.146072f
.ends

