* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 vdd.t102 vdd.t100 vdd.t101 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X1 CSoutput.t71 commonsourceibias.t32 gnd.t108 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X2 CSoutput.t34 a_n7677_7899.t20 vdd.t163 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X3 CSoutput.t35 a_n7677_7899.t21 vdd.t164 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X4 vdd.t212 a_n7677_7899.t22 CSoutput.t90 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 CSoutput.t70 commonsourceibias.t33 gnd.t107 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X6 vdd.t99 vdd.t97 vdd.t98 vdd.t68 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X7 a_n7677_7899.t14 plus.t5 a_n1455_n3628.t13 gnd.t217 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X8 vdd.t213 a_n7677_7899.t23 CSoutput.t91 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 a_n2511_10156.t19 a_n2686_12378.t25 a_n2686_12378.t26 vdd.t144 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X10 CSoutput.t72 a_n7677_7899.t24 vdd.t183 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 a_n2686_8022.t12 a_n2686_12378.t32 a_n7677_7899.t9 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X12 output.t15 CSoutput.t92 vdd.t198 gnd.t222 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X13 CSoutput.t73 a_n7677_7899.t25 vdd.t184 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 gnd.t106 commonsourceibias.t4 commonsourceibias.t5 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X15 vdd.t192 a_n7677_7899.t26 CSoutput.t80 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 CSoutput.t69 commonsourceibias.t34 gnd.t104 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X17 a_n2686_12378.t31 minus.t5 a_n1455_n3628.t19 gnd.t223 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X18 CSoutput.t81 a_n7677_7899.t27 vdd.t193 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t93 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X20 output.t14 CSoutput.t94 vdd.t12 gnd.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X21 a_n2686_12378.t18 a_n2686_12378.t17 a_n2511_10156.t18 vdd.t155 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X22 CSoutput.t86 a_n7677_7899.t28 vdd.t205 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t68 commonsourceibias.t35 gnd.t105 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X24 CSoutput.t67 commonsourceibias.t36 gnd.t103 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X25 a_n1455_n3628.t14 diffpairibias.t8 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X26 a_n1455_n3628.t5 minus.t6 a_n2686_12378.t2 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X27 CSoutput.t87 a_n7677_7899.t29 vdd.t206 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t102 commonsourceibias.t37 CSoutput.t66 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X29 diffpairibias.t7 diffpairibias.t6 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X30 plus.t4 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 gnd.t213 gnd.t210 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X32 vdd.t96 vdd.t94 vdd.t95 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X33 vdd.t93 vdd.t90 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X34 vdd.t152 a_n7677_7899.t30 CSoutput.t26 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t101 commonsourceibias.t38 CSoutput.t65 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X36 gnd.t209 gnd.t207 minus.t4 gnd.t208 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X37 gnd.t206 gnd.t203 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X38 gnd.t99 commonsourceibias.t30 commonsourceibias.t31 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X39 a_n2686_8022.t20 a_n2686_12378.t33 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X40 CSoutput.t64 commonsourceibias.t39 gnd.t100 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X41 gnd.t98 commonsourceibias.t40 CSoutput.t63 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X42 vdd.t153 a_n7677_7899.t31 CSoutput.t27 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t16 a_n7677_7899.t32 vdd.t119 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X44 commonsourceibias.t29 commonsourceibias.t28 gnd.t97 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X45 vdd.t13 CSoutput.t95 output.t13 gnd.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X46 diffpairibias.t5 diffpairibias.t4 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X47 commonsourceibias.t27 commonsourceibias.t26 gnd.t96 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X48 CSoutput.t17 a_n7677_7899.t33 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 gnd.t202 gnd.t200 gnd.t201 gnd.t110 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X50 a_n1455_n3628.t16 minus.t7 a_n2686_12378.t28 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X51 vdd.t18 a_n7677_7899.t34 CSoutput.t6 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 vdd.t20 a_n7677_7899.t35 CSoutput.t7 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 gnd.t199 gnd.t196 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X54 a_n2686_8022.t19 a_n2686_12378.t34 vdd.t143 vdd.t142 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X55 vdd.t89 vdd.t87 vdd.t88 vdd.t68 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X56 gnd.t195 gnd.t193 minus.t3 gnd.t194 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X57 output.t19 outputibias.t8 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X58 gnd.t95 commonsourceibias.t24 commonsourceibias.t25 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X59 CSoutput.t2 a_n7677_7899.t36 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 a_n1455_n3628.t1 diffpairibias.t9 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X61 CSoutput.t3 a_n7677_7899.t37 vdd.t11 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n7677_7899.t15 plus.t6 a_n1455_n3628.t12 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X63 gnd.t94 commonsourceibias.t22 commonsourceibias.t23 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X64 a_n2686_12378.t24 a_n2686_12378.t23 a_n2511_10156.t17 vdd.t172 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X65 a_n2686_12378.t10 a_n2686_12378.t9 a_n2511_10156.t16 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X66 commonsourceibias.t3 commonsourceibias.t2 gnd.t93 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X67 vdd.t86 vdd.t84 vdd.t85 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X68 plus.t3 gnd.t190 gnd.t192 gnd.t191 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X69 gnd.t90 commonsourceibias.t0 commonsourceibias.t1 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X70 output.t12 CSoutput.t96 vdd.t8 gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X71 gnd.t189 gnd.t187 gnd.t188 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X72 CSoutput.t62 commonsourceibias.t41 gnd.t92 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X73 a_n2686_8022.t11 a_n2686_12378.t35 a_n7677_7899.t12 vdd.t172 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X74 CSoutput.t12 a_n7677_7899.t38 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 vdd.t112 a_n7677_7899.t39 CSoutput.t13 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X76 CSoutput.t97 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X77 gnd.t91 commonsourceibias.t42 CSoutput.t61 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X78 a_n1455_n3628.t11 plus.t7 a_n7677_7899.t18 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X79 a_n2686_8022.t18 a_n2686_12378.t36 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X80 vdd.t104 a_n7677_7899.t40 CSoutput.t10 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X81 CSoutput.t98 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X82 gnd.t89 commonsourceibias.t43 CSoutput.t60 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X83 vdd.t83 vdd.t81 vdd.t82 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X84 a_n7677_7899.t19 a_n2686_12378.t37 a_n2686_8022.t10 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X85 vdd.t80 vdd.t78 vdd.t79 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X86 CSoutput.t59 commonsourceibias.t44 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X87 gnd.t86 commonsourceibias.t20 commonsourceibias.t21 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X88 a_n2511_10156.t15 a_n2686_12378.t7 a_n2686_12378.t8 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X89 vdd.t105 a_n7677_7899.t41 CSoutput.t11 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t99 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X91 vdd.t106 CSoutput.t100 output.t11 gnd.t16 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X92 CSoutput.t58 commonsourceibias.t45 gnd.t84 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X93 vdd.t24 a_n7677_7899.t42 CSoutput.t8 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 commonsourceibias.t19 commonsourceibias.t18 gnd.t83 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X95 gnd.t186 gnd.t184 gnd.t185 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X96 gnd.t82 commonsourceibias.t46 CSoutput.t57 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X97 vdd.t26 a_n7677_7899.t43 CSoutput.t9 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 CSoutput.t20 a_n7677_7899.t44 vdd.t132 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t183 gnd.t181 gnd.t182 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X100 vdd.t134 a_n7677_7899.t45 CSoutput.t21 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 CSoutput.t14 a_n7677_7899.t46 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 vdd.t77 vdd.t74 vdd.t76 vdd.t75 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X103 CSoutput.t56 commonsourceibias.t47 gnd.t81 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X104 vdd.t73 vdd.t71 vdd.t72 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X105 a_n7677_7899.t10 a_n2686_12378.t38 a_n2686_8022.t9 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X106 vdd.t146 a_n2686_12378.t39 a_n2511_10156.t7 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X107 vdd.t117 a_n7677_7899.t47 CSoutput.t15 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t180 gnd.t178 plus.t2 gnd.t179 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X109 a_n7677_7899.t1 plus.t8 a_n1455_n3628.t10 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X110 a_n2686_8022.t8 a_n2686_12378.t40 a_n7677_7899.t5 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X111 minus.t2 gnd.t175 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X112 commonsourceibias.t11 commonsourceibias.t10 gnd.t80 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X113 CSoutput.t78 a_n7677_7899.t48 vdd.t190 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X114 a_n2511_10156.t14 a_n2686_12378.t21 a_n2686_12378.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X115 vdd.t191 a_n7677_7899.t49 CSoutput.t79 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 a_n7677_7899.t0 a_n2686_12378.t41 a_n2686_8022.t7 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X117 outputibias.t7 outputibias.t6 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X118 vdd.t178 a_n2686_12378.t42 a_n2511_10156.t6 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X119 vdd.t166 a_n2686_12378.t43 a_n2686_8022.t17 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X120 gnd.t79 commonsourceibias.t48 CSoutput.t55 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X121 diffpairibias.t3 diffpairibias.t2 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X122 outputibias.t5 outputibias.t4 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X123 outputibias.t3 outputibias.t2 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X124 gnd.t174 gnd.t172 gnd.t173 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X125 CSoutput.t82 a_n7677_7899.t50 vdd.t199 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X126 a_n2686_8022.t6 a_n2686_12378.t44 a_n7677_7899.t7 vdd.t155 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X127 CSoutput.t54 commonsourceibias.t49 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X128 vdd.t107 CSoutput.t101 output.t10 gnd.t17 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X129 vdd.t202 a_n2686_12378.t45 a_n2686_8022.t16 vdd.t201 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X130 gnd.t76 commonsourceibias.t50 CSoutput.t53 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X131 gnd.t171 gnd.t169 gnd.t170 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X132 gnd.t75 commonsourceibias.t51 CSoutput.t52 gnd.t74 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X133 a_n1455_n3628.t4 minus.t8 a_n2686_12378.t1 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X134 CSoutput.t83 a_n7677_7899.t51 vdd.t200 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 a_n2686_8022.t5 a_n2686_12378.t46 a_n7677_7899.t4 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X136 vdd.t70 vdd.t67 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X137 vdd.t130 a_n7677_7899.t52 CSoutput.t18 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 vdd.t131 a_n7677_7899.t53 CSoutput.t19 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t168 gnd.t166 plus.t1 gnd.t167 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X140 vdd.t125 a_n2686_12378.t47 a_n2511_10156.t5 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X141 vdd.t66 vdd.t64 vdd.t65 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X142 a_n1455_n3628.t2 diffpairibias.t10 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X143 gnd.t165 gnd.t163 gnd.t164 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X144 a_n2511_10156.t4 a_n2686_12378.t48 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X145 CSoutput.t74 a_n7677_7899.t54 vdd.t185 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 CSoutput.t75 a_n7677_7899.t55 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 CSoutput.t51 commonsourceibias.t52 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X148 outputibias.t1 outputibias.t0 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X149 a_n2686_12378.t27 minus.t9 a_n1455_n3628.t15 gnd.t217 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X150 CSoutput.t0 a_n7677_7899.t56 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 a_n1455_n3628.t9 plus.t9 a_n7677_7899.t2 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X152 a_n7677_7899.t13 a_n2686_12378.t49 a_n2686_8022.t4 vdd.t176 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X153 output.t9 CSoutput.t102 vdd.t207 gnd.t225 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X154 gnd.t71 commonsourceibias.t53 CSoutput.t50 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X155 gnd.t70 commonsourceibias.t54 CSoutput.t49 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X156 gnd.t69 commonsourceibias.t55 CSoutput.t48 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X157 a_n7677_7899.t16 plus.t10 a_n1455_n3628.t8 gnd.t223 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X158 a_n2686_12378.t0 minus.t10 a_n1455_n3628.t3 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X159 CSoutput.t1 a_n7677_7899.t57 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 a_n1455_n3628.t7 plus.t11 a_n7677_7899.t17 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X161 vdd.t15 a_n7677_7899.t58 CSoutput.t4 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t63 vdd.t60 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X163 a_n2511_10156.t13 a_n2686_12378.t3 a_n2686_12378.t4 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X164 vdd.t17 a_n7677_7899.t59 CSoutput.t5 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n2686_12378.t16 a_n2686_12378.t15 a_n2511_10156.t12 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X166 vdd.t123 a_n2686_12378.t50 a_n2686_8022.t15 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X167 vdd.t208 CSoutput.t103 output.t8 gnd.t226 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X168 CSoutput.t24 a_n7677_7899.t60 vdd.t150 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 output.t7 CSoutput.t104 vdd.t209 gnd.t227 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X170 CSoutput.t25 a_n7677_7899.t61 vdd.t151 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n2686_12378.t20 a_n2686_12378.t19 a_n2511_10156.t11 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X172 gnd.t162 gnd.t159 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X173 gnd.t158 gnd.t155 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X174 a_n7677_7899.t6 a_n2686_12378.t51 a_n2686_8022.t3 vdd.t144 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X175 output.t6 CSoutput.t105 vdd.t196 gnd.t220 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 CSoutput.t38 a_n7677_7899.t62 vdd.t170 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n2686_8022.t2 a_n2686_12378.t52 a_n7677_7899.t11 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X178 vdd.t171 a_n7677_7899.t63 CSoutput.t39 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 commonsourceibias.t7 commonsourceibias.t6 gnd.t67 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X180 gnd.t66 commonsourceibias.t56 CSoutput.t47 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=2
X181 a_n1455_n3628.t18 minus.t11 a_n2686_12378.t30 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X182 gnd.t154 gnd.t152 gnd.t153 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X183 vdd.t59 vdd.t57 vdd.t58 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 a_n1455_n3628.t0 diffpairibias.t11 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X185 gnd.t151 gnd.t149 gnd.t150 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X186 vdd.t195 a_n2686_12378.t53 a_n2686_8022.t14 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X187 vdd.t161 a_n7677_7899.t64 CSoutput.t32 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 vdd.t56 vdd.t53 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X189 a_n2511_10156.t10 a_n2686_12378.t13 a_n2686_12378.t14 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X190 CSoutput.t106 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X191 gnd.t64 commonsourceibias.t14 commonsourceibias.t15 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X192 a_n2686_8022.t13 a_n2686_12378.t54 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X193 output.t5 CSoutput.t107 vdd.t197 gnd.t221 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X194 a_n2511_10156.t3 a_n2686_12378.t55 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X195 vdd.t162 a_n7677_7899.t65 CSoutput.t33 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X196 gnd.t148 gnd.t145 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X197 gnd.t144 gnd.t141 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X198 a_n2511_10156.t2 a_n2686_12378.t56 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X199 gnd.t63 commonsourceibias.t12 commonsourceibias.t13 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X200 vdd.t108 CSoutput.t108 output.t4 gnd.t19 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X201 a_n7677_7899.t8 a_n2686_12378.t57 a_n2686_8022.t1 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X202 minus.t1 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X203 CSoutput.t36 a_n7677_7899.t66 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 gnd.t61 commonsourceibias.t57 CSoutput.t46 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X205 gnd.t59 commonsourceibias.t58 CSoutput.t45 gnd.t58 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X206 CSoutput.t44 commonsourceibias.t59 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X207 vdd.t52 vdd.t50 vdd.t51 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X208 vdd.t169 a_n7677_7899.t67 CSoutput.t37 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 diffpairibias.t1 diffpairibias.t0 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X210 CSoutput.t30 a_n7677_7899.t68 vdd.t159 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 gnd.t137 gnd.t135 gnd.t136 gnd.t110 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X212 CSoutput.t43 commonsourceibias.t60 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=2
X213 vdd.t160 a_n7677_7899.t69 CSoutput.t31 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 vdd.t210 a_n7677_7899.t70 CSoutput.t88 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n2686_12378.t12 a_n2686_12378.t11 a_n2511_10156.t9 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X216 CSoutput.t109 a_n2686_8022.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X217 output.t18 outputibias.t9 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X218 commonsourceibias.t17 commonsourceibias.t16 gnd.t53 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X219 vdd.t211 a_n7677_7899.t71 CSoutput.t89 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X221 output.t17 outputibias.t10 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X222 gnd.t134 gnd.t131 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X223 vdd.t109 CSoutput.t110 output.t3 gnd.t20 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X224 vdd.t215 a_n2686_12378.t58 a_n2511_10156.t1 vdd.t214 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X225 vdd.t188 a_n7677_7899.t72 CSoutput.t76 vdd.t133 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X227 output.t16 outputibias.t11 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X228 vdd.t41 vdd.t39 vdd.t40 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X229 vdd.t126 CSoutput.t111 output.t2 gnd.t22 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X230 output.t1 CSoutput.t112 vdd.t127 gnd.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X231 CSoutput.t77 a_n7677_7899.t73 vdd.t189 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 vdd.t203 a_n7677_7899.t74 CSoutput.t84 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X233 CSoutput.t42 commonsourceibias.t61 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X234 CSoutput.t41 commonsourceibias.t62 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X235 a_n2511_10156.t0 a_n2686_12378.t59 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X236 gnd.t130 gnd.t127 gnd.t129 gnd.t128 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X237 vdd.t204 a_n7677_7899.t75 CSoutput.t85 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t126 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X239 CSoutput.t22 a_n7677_7899.t76 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X240 CSoutput.t23 a_n7677_7899.t77 vdd.t149 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 gnd.t122 gnd.t119 gnd.t121 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X242 gnd.t118 gnd.t116 plus.t0 gnd.t117 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X243 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X244 gnd.t48 commonsourceibias.t63 CSoutput.t40 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X245 vdd.t157 a_n7677_7899.t78 CSoutput.t28 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 vdd.t34 vdd.t31 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X247 vdd.t128 CSoutput.t113 output.t0 gnd.t24 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X248 a_n1455_n3628.t6 plus.t12 a_n7677_7899.t3 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X249 a_n2686_12378.t29 minus.t12 a_n1455_n3628.t17 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X250 commonsourceibias.t9 commonsourceibias.t8 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=2
X251 a_n2511_10156.t8 a_n2686_12378.t5 a_n2686_12378.t6 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X252 vdd.t30 vdd.t27 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X253 CSoutput.t29 a_n7677_7899.t79 vdd.t158 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t115 gnd.t113 minus.t0 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X255 gnd.t112 gnd.t109 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
R0 vdd.n2710 vdd.n112 452.195
R1 vdd.n2603 vdd.n110 452.195
R2 vdd.n316 vdd.n281 452.195
R3 vdd.n2496 vdd.n283 452.195
R4 vdd.n1411 vdd.n729 452.195
R5 vdd.n1414 vdd.n1413 452.195
R6 vdd.n900 vdd.n866 452.195
R7 vdd.n1077 vdd.n868 452.195
R8 vdd.n982 vdd.t42 371.625
R9 vdd.n1015 vdd.t57 371.625
R10 vdd.n1048 vdd.t84 371.625
R11 vdd.n718 vdd.t87 371.625
R12 vdd.n1290 vdd.t97 371.625
R13 vdd.n1255 vdd.t67 371.625
R14 vdd.n212 vdd.t27 371.625
R15 vdd.n179 vdd.t39 371.625
R16 vdd.n144 vdd.t71 371.625
R17 vdd.n354 vdd.t81 371.625
R18 vdd.n2463 vdd.t50 371.625
R19 vdd.n2380 vdd.t35 371.625
R20 vdd.n702 vdd.t64 347.526
R21 vdd.n553 vdd.t78 347.526
R22 vdd.n695 vdd.t31 347.526
R23 vdd.n563 vdd.t53 347.526
R24 vdd.n421 vdd.t74 347.526
R25 vdd.n1900 vdd.t100 347.526
R26 vdd.n404 vdd.t94 347.526
R27 vdd.n1906 vdd.t46 347.526
R28 vdd.n377 vdd.t60 347.526
R29 vdd.n663 vdd.t90 347.526
R30 vdd.n2140 vdd.n522 294.147
R31 vdd.n2344 vdd.n387 294.147
R32 vdd.n2296 vdd.n384 294.147
R33 vdd.n1967 vdd.n1884 294.147
R34 vdd.n1823 vdd.n561 294.147
R35 vdd.n1772 vdd.n1771 294.147
R36 vdd.n1597 vdd.n680 294.147
R37 vdd.n1648 vdd.n682 294.147
R38 vdd.n2275 vdd.n385 294.147
R39 vdd.n2347 vdd.n2346 294.147
R40 vdd.n2086 vdd.n1885 294.147
R41 vdd.n2138 vdd.n1887 294.147
R42 vdd.n1881 vdd.n550 294.147
R43 vdd.n1830 vdd.n549 294.147
R44 vdd.n1480 vdd.n681 294.147
R45 vdd.n1650 vdd.n678 294.147
R46 vdd.n702 vdd.t66 293.986
R47 vdd.n553 vdd.t79 293.986
R48 vdd.n695 vdd.t34 293.986
R49 vdd.n563 vdd.t55 293.986
R50 vdd.n421 vdd.t76 293.986
R51 vdd.n421 vdd.t77 293.986
R52 vdd.n1900 vdd.t102 293.986
R53 vdd.n404 vdd.t95 293.986
R54 vdd.n1906 vdd.t49 293.986
R55 vdd.n377 vdd.t62 293.986
R56 vdd.n663 vdd.t92 293.986
R57 vdd.n663 vdd.t93 293.986
R58 vdd.n703 vdd.t65 268.192
R59 vdd.n554 vdd.t80 268.192
R60 vdd.n696 vdd.t33 268.192
R61 vdd.n564 vdd.t56 268.192
R62 vdd.n1901 vdd.t101 268.192
R63 vdd.n405 vdd.t96 268.192
R64 vdd.n1907 vdd.t48 268.192
R65 vdd.n378 vdd.t63 268.192
R66 vdd.n2277 vdd.n385 185
R67 vdd.n2345 vdd.n385 185
R68 vdd.n2279 vdd.n2278 185
R69 vdd.n2278 vdd.n383 185
R70 vdd.n2280 vdd.n412 185
R71 vdd.n2290 vdd.n412 185
R72 vdd.n2281 vdd.n420 185
R73 vdd.n420 vdd.n410 185
R74 vdd.n2283 vdd.n2282 185
R75 vdd.n2284 vdd.n2283 185
R76 vdd.n2245 vdd.n419 185
R77 vdd.n419 vdd.n416 185
R78 vdd.n2243 vdd.n2242 185
R79 vdd.n2242 vdd.n2241 185
R80 vdd.n423 vdd.n422 185
R81 vdd.n424 vdd.n423 185
R82 vdd.n2234 vdd.n2233 185
R83 vdd.n2235 vdd.n2234 185
R84 vdd.n2232 vdd.n433 185
R85 vdd.n433 vdd.n430 185
R86 vdd.n2231 vdd.n2230 185
R87 vdd.n2230 vdd.n2229 185
R88 vdd.n435 vdd.n434 185
R89 vdd.n443 vdd.n435 185
R90 vdd.n2222 vdd.n2221 185
R91 vdd.n2223 vdd.n2222 185
R92 vdd.n2220 vdd.n444 185
R93 vdd.n449 vdd.n444 185
R94 vdd.n2219 vdd.n2218 185
R95 vdd.n2218 vdd.n2217 185
R96 vdd.n446 vdd.n445 185
R97 vdd.n455 vdd.n446 185
R98 vdd.n2210 vdd.n2209 185
R99 vdd.n2211 vdd.n2210 185
R100 vdd.n2208 vdd.n456 185
R101 vdd.n461 vdd.n456 185
R102 vdd.n2207 vdd.n2206 185
R103 vdd.n2206 vdd.n2205 185
R104 vdd.n458 vdd.n457 185
R105 vdd.n467 vdd.n458 185
R106 vdd.n2198 vdd.n2197 185
R107 vdd.n2199 vdd.n2198 185
R108 vdd.n2196 vdd.n468 185
R109 vdd.n2051 vdd.n468 185
R110 vdd.n2195 vdd.n2194 185
R111 vdd.n2194 vdd.n2193 185
R112 vdd.n470 vdd.n469 185
R113 vdd.n471 vdd.n470 185
R114 vdd.n2186 vdd.n2185 185
R115 vdd.n2187 vdd.n2186 185
R116 vdd.n2184 vdd.n479 185
R117 vdd.n2060 vdd.n479 185
R118 vdd.n2183 vdd.n2182 185
R119 vdd.n2182 vdd.n2181 185
R120 vdd.n481 vdd.n480 185
R121 vdd.n482 vdd.n481 185
R122 vdd.n2174 vdd.n2173 185
R123 vdd.n2175 vdd.n2174 185
R124 vdd.n2172 vdd.n491 185
R125 vdd.n491 vdd.n488 185
R126 vdd.n2171 vdd.n2170 185
R127 vdd.n2170 vdd.n2169 185
R128 vdd.n493 vdd.n492 185
R129 vdd.n502 vdd.n493 185
R130 vdd.n2162 vdd.n2161 185
R131 vdd.n2163 vdd.n2162 185
R132 vdd.n2160 vdd.n503 185
R133 vdd.n503 vdd.n499 185
R134 vdd.n2159 vdd.n2158 185
R135 vdd.n2158 vdd.n2157 185
R136 vdd.n505 vdd.n504 185
R137 vdd.n513 vdd.n505 185
R138 vdd.n2150 vdd.n2149 185
R139 vdd.n2151 vdd.n2150 185
R140 vdd.n2148 vdd.n514 185
R141 vdd.n519 vdd.n514 185
R142 vdd.n2147 vdd.n2146 185
R143 vdd.n2146 vdd.n2145 185
R144 vdd.n516 vdd.n515 185
R145 vdd.n1886 vdd.n516 185
R146 vdd.n2138 vdd.n2137 185
R147 vdd.n2139 vdd.n2138 185
R148 vdd.n2136 vdd.n1887 185
R149 vdd.n2135 vdd.n2134 185
R150 vdd.n2132 vdd.n1888 185
R151 vdd.n2130 vdd.n2129 185
R152 vdd.n2128 vdd.n1889 185
R153 vdd.n2127 vdd.n2126 185
R154 vdd.n2124 vdd.n1890 185
R155 vdd.n2122 vdd.n2121 185
R156 vdd.n2120 vdd.n1891 185
R157 vdd.n2119 vdd.n2118 185
R158 vdd.n2116 vdd.n1892 185
R159 vdd.n2114 vdd.n2113 185
R160 vdd.n2112 vdd.n1893 185
R161 vdd.n2111 vdd.n2110 185
R162 vdd.n2108 vdd.n1894 185
R163 vdd.n2106 vdd.n2105 185
R164 vdd.n2104 vdd.n1895 185
R165 vdd.n2103 vdd.n2102 185
R166 vdd.n2100 vdd.n1896 185
R167 vdd.n2098 vdd.n2097 185
R168 vdd.n2096 vdd.n1897 185
R169 vdd.n2095 vdd.n2094 185
R170 vdd.n2092 vdd.n1898 185
R171 vdd.n2090 vdd.n2089 185
R172 vdd.n2088 vdd.n1899 185
R173 vdd.n2087 vdd.n2086 185
R174 vdd.n2348 vdd.n2347 185
R175 vdd.n2349 vdd.n376 185
R176 vdd.n2351 vdd.n2350 185
R177 vdd.n2353 vdd.n374 185
R178 vdd.n2355 vdd.n2354 185
R179 vdd.n2356 vdd.n373 185
R180 vdd.n2358 vdd.n2357 185
R181 vdd.n2360 vdd.n371 185
R182 vdd.n2362 vdd.n2361 185
R183 vdd.n2363 vdd.n370 185
R184 vdd.n2365 vdd.n2364 185
R185 vdd.n2367 vdd.n368 185
R186 vdd.n2369 vdd.n2368 185
R187 vdd.n2254 vdd.n367 185
R188 vdd.n2256 vdd.n2255 185
R189 vdd.n2258 vdd.n2252 185
R190 vdd.n2260 vdd.n2259 185
R191 vdd.n2261 vdd.n2251 185
R192 vdd.n2263 vdd.n2262 185
R193 vdd.n2265 vdd.n2249 185
R194 vdd.n2267 vdd.n2266 185
R195 vdd.n2268 vdd.n2248 185
R196 vdd.n2270 vdd.n2269 185
R197 vdd.n2272 vdd.n2247 185
R198 vdd.n2273 vdd.n2246 185
R199 vdd.n2276 vdd.n2275 185
R200 vdd.n2346 vdd.n380 185
R201 vdd.n2346 vdd.n2345 185
R202 vdd.n2020 vdd.n382 185
R203 vdd.n383 vdd.n382 185
R204 vdd.n2021 vdd.n411 185
R205 vdd.n2290 vdd.n411 185
R206 vdd.n2023 vdd.n2022 185
R207 vdd.n2022 vdd.n410 185
R208 vdd.n2024 vdd.n418 185
R209 vdd.n2284 vdd.n418 185
R210 vdd.n2026 vdd.n2025 185
R211 vdd.n2025 vdd.n416 185
R212 vdd.n2027 vdd.n426 185
R213 vdd.n2241 vdd.n426 185
R214 vdd.n2029 vdd.n2028 185
R215 vdd.n2028 vdd.n424 185
R216 vdd.n2030 vdd.n432 185
R217 vdd.n2235 vdd.n432 185
R218 vdd.n2032 vdd.n2031 185
R219 vdd.n2031 vdd.n430 185
R220 vdd.n2033 vdd.n437 185
R221 vdd.n2229 vdd.n437 185
R222 vdd.n2035 vdd.n2034 185
R223 vdd.n2034 vdd.n443 185
R224 vdd.n2036 vdd.n442 185
R225 vdd.n2223 vdd.n442 185
R226 vdd.n2038 vdd.n2037 185
R227 vdd.n2037 vdd.n449 185
R228 vdd.n2039 vdd.n448 185
R229 vdd.n2217 vdd.n448 185
R230 vdd.n2041 vdd.n2040 185
R231 vdd.n2040 vdd.n455 185
R232 vdd.n2042 vdd.n454 185
R233 vdd.n2211 vdd.n454 185
R234 vdd.n2044 vdd.n2043 185
R235 vdd.n2043 vdd.n461 185
R236 vdd.n2045 vdd.n460 185
R237 vdd.n2205 vdd.n460 185
R238 vdd.n2047 vdd.n2046 185
R239 vdd.n2046 vdd.n467 185
R240 vdd.n2048 vdd.n466 185
R241 vdd.n2199 vdd.n466 185
R242 vdd.n2050 vdd.n2049 185
R243 vdd.n2051 vdd.n2050 185
R244 vdd.n2019 vdd.n473 185
R245 vdd.n2193 vdd.n473 185
R246 vdd.n2018 vdd.n2017 185
R247 vdd.n2017 vdd.n471 185
R248 vdd.n1903 vdd.n478 185
R249 vdd.n2187 vdd.n478 185
R250 vdd.n2062 vdd.n2061 185
R251 vdd.n2061 vdd.n2060 185
R252 vdd.n2063 vdd.n484 185
R253 vdd.n2181 vdd.n484 185
R254 vdd.n2065 vdd.n2064 185
R255 vdd.n2064 vdd.n482 185
R256 vdd.n2066 vdd.n490 185
R257 vdd.n2175 vdd.n490 185
R258 vdd.n2068 vdd.n2067 185
R259 vdd.n2067 vdd.n488 185
R260 vdd.n2069 vdd.n495 185
R261 vdd.n2169 vdd.n495 185
R262 vdd.n2071 vdd.n2070 185
R263 vdd.n2070 vdd.n502 185
R264 vdd.n2072 vdd.n501 185
R265 vdd.n2163 vdd.n501 185
R266 vdd.n2074 vdd.n2073 185
R267 vdd.n2073 vdd.n499 185
R268 vdd.n2075 vdd.n507 185
R269 vdd.n2157 vdd.n507 185
R270 vdd.n2077 vdd.n2076 185
R271 vdd.n2076 vdd.n513 185
R272 vdd.n2078 vdd.n512 185
R273 vdd.n2151 vdd.n512 185
R274 vdd.n2080 vdd.n2079 185
R275 vdd.n2079 vdd.n519 185
R276 vdd.n2081 vdd.n518 185
R277 vdd.n2145 vdd.n518 185
R278 vdd.n2083 vdd.n2082 185
R279 vdd.n2082 vdd.n1886 185
R280 vdd.n2084 vdd.n1885 185
R281 vdd.n2139 vdd.n1885 185
R282 vdd.n1411 vdd.n1410 185
R283 vdd.n1412 vdd.n1411 185
R284 vdd.n730 vdd.n728 185
R285 vdd.n728 vdd.n725 185
R286 vdd.n1224 vdd.n1223 185
R287 vdd.n1223 vdd.n1222 185
R288 vdd.n733 vdd.n732 185
R289 vdd.n734 vdd.n733 185
R290 vdd.n1212 vdd.n1211 185
R291 vdd.n1213 vdd.n1212 185
R292 vdd.n743 vdd.n742 185
R293 vdd.n742 vdd.n741 185
R294 vdd.n1207 vdd.n1206 185
R295 vdd.n1206 vdd.n1205 185
R296 vdd.n746 vdd.n745 185
R297 vdd.n753 vdd.n746 185
R298 vdd.n1196 vdd.n1195 185
R299 vdd.n1197 vdd.n1196 185
R300 vdd.n755 vdd.n754 185
R301 vdd.n754 vdd.n752 185
R302 vdd.n1191 vdd.n1190 185
R303 vdd.n1190 vdd.n1189 185
R304 vdd.n758 vdd.n757 185
R305 vdd.n759 vdd.n758 185
R306 vdd.n1180 vdd.n1179 185
R307 vdd.n1181 vdd.n1180 185
R308 vdd.n767 vdd.n766 185
R309 vdd.n766 vdd.n765 185
R310 vdd.n1175 vdd.n1174 185
R311 vdd.n1174 vdd.n1173 185
R312 vdd.n770 vdd.n769 185
R313 vdd.n777 vdd.n770 185
R314 vdd.n1164 vdd.n1163 185
R315 vdd.n1165 vdd.n1164 185
R316 vdd.n779 vdd.n778 185
R317 vdd.n778 vdd.n776 185
R318 vdd.n1159 vdd.n1158 185
R319 vdd.n1158 vdd.n1157 185
R320 vdd.n812 vdd.n811 185
R321 vdd.n813 vdd.n812 185
R322 vdd.n1148 vdd.n1147 185
R323 vdd.n1149 vdd.n1148 185
R324 vdd.n821 vdd.n820 185
R325 vdd.n820 vdd.n819 185
R326 vdd.n1142 vdd.n1141 185
R327 vdd.n1141 vdd.n1140 185
R328 vdd.n824 vdd.n823 185
R329 vdd.n831 vdd.n824 185
R330 vdd.n1131 vdd.n1130 185
R331 vdd.n1132 vdd.n1131 185
R332 vdd.n833 vdd.n832 185
R333 vdd.n832 vdd.n830 185
R334 vdd.n1126 vdd.n1125 185
R335 vdd.n1125 vdd.n1124 185
R336 vdd.n836 vdd.n835 185
R337 vdd.n837 vdd.n836 185
R338 vdd.n1115 vdd.n1114 185
R339 vdd.n1116 vdd.n1115 185
R340 vdd.n845 vdd.n844 185
R341 vdd.n844 vdd.n843 185
R342 vdd.n1110 vdd.n1109 185
R343 vdd.n1109 vdd.n1108 185
R344 vdd.n848 vdd.n847 185
R345 vdd.n855 vdd.n848 185
R346 vdd.n1099 vdd.n1098 185
R347 vdd.n1100 vdd.n1099 185
R348 vdd.n857 vdd.n856 185
R349 vdd.n856 vdd.n854 185
R350 vdd.n1094 vdd.n1093 185
R351 vdd.n1093 vdd.n1092 185
R352 vdd.n860 vdd.n859 185
R353 vdd.n861 vdd.n860 185
R354 vdd.n1083 vdd.n1082 185
R355 vdd.n1084 vdd.n1083 185
R356 vdd.n869 vdd.n868 185
R357 vdd.n868 vdd.n867 185
R358 vdd.n1078 vdd.n1077 185
R359 vdd.n872 vdd.n871 185
R360 vdd.n1074 vdd.n1073 185
R361 vdd.n1075 vdd.n1074 185
R362 vdd.n902 vdd.n901 185
R363 vdd.n1069 vdd.n904 185
R364 vdd.n1068 vdd.n905 185
R365 vdd.n1067 vdd.n906 185
R366 vdd.n908 vdd.n907 185
R367 vdd.n1063 vdd.n910 185
R368 vdd.n1062 vdd.n911 185
R369 vdd.n1061 vdd.n912 185
R370 vdd.n914 vdd.n913 185
R371 vdd.n1057 vdd.n916 185
R372 vdd.n1056 vdd.n917 185
R373 vdd.n1055 vdd.n918 185
R374 vdd.n920 vdd.n919 185
R375 vdd.n1051 vdd.n922 185
R376 vdd.n1050 vdd.n1047 185
R377 vdd.n1046 vdd.n923 185
R378 vdd.n925 vdd.n924 185
R379 vdd.n1042 vdd.n927 185
R380 vdd.n1041 vdd.n928 185
R381 vdd.n1040 vdd.n929 185
R382 vdd.n931 vdd.n930 185
R383 vdd.n1036 vdd.n933 185
R384 vdd.n1035 vdd.n934 185
R385 vdd.n1034 vdd.n935 185
R386 vdd.n937 vdd.n936 185
R387 vdd.n1030 vdd.n939 185
R388 vdd.n1029 vdd.n940 185
R389 vdd.n1028 vdd.n941 185
R390 vdd.n943 vdd.n942 185
R391 vdd.n1024 vdd.n945 185
R392 vdd.n1023 vdd.n946 185
R393 vdd.n1022 vdd.n947 185
R394 vdd.n949 vdd.n948 185
R395 vdd.n1018 vdd.n951 185
R396 vdd.n1017 vdd.n1014 185
R397 vdd.n1013 vdd.n952 185
R398 vdd.n954 vdd.n953 185
R399 vdd.n1009 vdd.n956 185
R400 vdd.n1008 vdd.n957 185
R401 vdd.n1007 vdd.n958 185
R402 vdd.n960 vdd.n959 185
R403 vdd.n1003 vdd.n962 185
R404 vdd.n1002 vdd.n963 185
R405 vdd.n1001 vdd.n964 185
R406 vdd.n966 vdd.n965 185
R407 vdd.n997 vdd.n968 185
R408 vdd.n996 vdd.n969 185
R409 vdd.n995 vdd.n970 185
R410 vdd.n972 vdd.n971 185
R411 vdd.n991 vdd.n974 185
R412 vdd.n990 vdd.n975 185
R413 vdd.n989 vdd.n976 185
R414 vdd.n978 vdd.n977 185
R415 vdd.n985 vdd.n980 185
R416 vdd.n981 vdd.n900 185
R417 vdd.n1075 vdd.n900 185
R418 vdd.n1415 vdd.n1414 185
R419 vdd.n721 vdd.n716 185
R420 vdd.n1419 vdd.n715 185
R421 vdd.n1420 vdd.n714 185
R422 vdd.n1421 vdd.n713 185
R423 vdd.n1311 vdd.n712 185
R424 vdd.n1313 vdd.n1312 185
R425 vdd.n1315 vdd.n1309 185
R426 vdd.n1317 vdd.n1316 185
R427 vdd.n1319 vdd.n1307 185
R428 vdd.n1321 vdd.n1320 185
R429 vdd.n1322 vdd.n1302 185
R430 vdd.n1324 vdd.n1323 185
R431 vdd.n1326 vdd.n1300 185
R432 vdd.n1328 vdd.n1327 185
R433 vdd.n1329 vdd.n1296 185
R434 vdd.n1331 vdd.n1330 185
R435 vdd.n1333 vdd.n1294 185
R436 vdd.n1335 vdd.n1334 185
R437 vdd.n1289 vdd.n1288 185
R438 vdd.n1340 vdd.n1339 185
R439 vdd.n1342 vdd.n1286 185
R440 vdd.n1344 vdd.n1343 185
R441 vdd.n1345 vdd.n1281 185
R442 vdd.n1347 vdd.n1346 185
R443 vdd.n1349 vdd.n1279 185
R444 vdd.n1351 vdd.n1350 185
R445 vdd.n1352 vdd.n1274 185
R446 vdd.n1354 vdd.n1353 185
R447 vdd.n1356 vdd.n1272 185
R448 vdd.n1358 vdd.n1357 185
R449 vdd.n1359 vdd.n1267 185
R450 vdd.n1361 vdd.n1360 185
R451 vdd.n1363 vdd.n1265 185
R452 vdd.n1365 vdd.n1364 185
R453 vdd.n1366 vdd.n1261 185
R454 vdd.n1368 vdd.n1367 185
R455 vdd.n1370 vdd.n1259 185
R456 vdd.n1372 vdd.n1371 185
R457 vdd.n1254 vdd.n1253 185
R458 vdd.n1377 vdd.n1376 185
R459 vdd.n1379 vdd.n1251 185
R460 vdd.n1381 vdd.n1380 185
R461 vdd.n1382 vdd.n1246 185
R462 vdd.n1384 vdd.n1383 185
R463 vdd.n1386 vdd.n1244 185
R464 vdd.n1388 vdd.n1387 185
R465 vdd.n1389 vdd.n1241 185
R466 vdd.n1391 vdd.n1390 185
R467 vdd.n1393 vdd.n1238 185
R468 vdd.n1395 vdd.n1394 185
R469 vdd.n1239 vdd.n1236 185
R470 vdd.n1399 vdd.n1235 185
R471 vdd.n1400 vdd.n1230 185
R472 vdd.n1402 vdd.n1401 185
R473 vdd.n1404 vdd.n1228 185
R474 vdd.n1406 vdd.n1405 185
R475 vdd.n1407 vdd.n729 185
R476 vdd.n1413 vdd.n724 185
R477 vdd.n1413 vdd.n1412 185
R478 vdd.n737 vdd.n723 185
R479 vdd.n725 vdd.n723 185
R480 vdd.n1221 vdd.n1220 185
R481 vdd.n1222 vdd.n1221 185
R482 vdd.n736 vdd.n735 185
R483 vdd.n735 vdd.n734 185
R484 vdd.n1215 vdd.n1214 185
R485 vdd.n1214 vdd.n1213 185
R486 vdd.n740 vdd.n739 185
R487 vdd.n741 vdd.n740 185
R488 vdd.n1204 vdd.n1203 185
R489 vdd.n1205 vdd.n1204 185
R490 vdd.n748 vdd.n747 185
R491 vdd.n753 vdd.n747 185
R492 vdd.n1199 vdd.n1198 185
R493 vdd.n1198 vdd.n1197 185
R494 vdd.n751 vdd.n750 185
R495 vdd.n752 vdd.n751 185
R496 vdd.n1188 vdd.n1187 185
R497 vdd.n1189 vdd.n1188 185
R498 vdd.n761 vdd.n760 185
R499 vdd.n760 vdd.n759 185
R500 vdd.n1183 vdd.n1182 185
R501 vdd.n1182 vdd.n1181 185
R502 vdd.n764 vdd.n763 185
R503 vdd.n765 vdd.n764 185
R504 vdd.n1172 vdd.n1171 185
R505 vdd.n1173 vdd.n1172 185
R506 vdd.n772 vdd.n771 185
R507 vdd.n777 vdd.n771 185
R508 vdd.n1167 vdd.n1166 185
R509 vdd.n1166 vdd.n1165 185
R510 vdd.n775 vdd.n774 185
R511 vdd.n776 vdd.n775 185
R512 vdd.n1156 vdd.n1155 185
R513 vdd.n1157 vdd.n1156 185
R514 vdd.n815 vdd.n814 185
R515 vdd.n814 vdd.n813 185
R516 vdd.n1151 vdd.n1150 185
R517 vdd.n1150 vdd.n1149 185
R518 vdd.n818 vdd.n817 185
R519 vdd.n819 vdd.n818 185
R520 vdd.n1139 vdd.n1138 185
R521 vdd.n1140 vdd.n1139 185
R522 vdd.n826 vdd.n825 185
R523 vdd.n831 vdd.n825 185
R524 vdd.n1134 vdd.n1133 185
R525 vdd.n1133 vdd.n1132 185
R526 vdd.n829 vdd.n828 185
R527 vdd.n830 vdd.n829 185
R528 vdd.n1123 vdd.n1122 185
R529 vdd.n1124 vdd.n1123 185
R530 vdd.n839 vdd.n838 185
R531 vdd.n838 vdd.n837 185
R532 vdd.n1118 vdd.n1117 185
R533 vdd.n1117 vdd.n1116 185
R534 vdd.n842 vdd.n841 185
R535 vdd.n843 vdd.n842 185
R536 vdd.n1107 vdd.n1106 185
R537 vdd.n1108 vdd.n1107 185
R538 vdd.n850 vdd.n849 185
R539 vdd.n855 vdd.n849 185
R540 vdd.n1102 vdd.n1101 185
R541 vdd.n1101 vdd.n1100 185
R542 vdd.n853 vdd.n852 185
R543 vdd.n854 vdd.n853 185
R544 vdd.n1091 vdd.n1090 185
R545 vdd.n1092 vdd.n1091 185
R546 vdd.n863 vdd.n862 185
R547 vdd.n862 vdd.n861 185
R548 vdd.n1086 vdd.n1085 185
R549 vdd.n1085 vdd.n1084 185
R550 vdd.n866 vdd.n865 185
R551 vdd.n867 vdd.n866 185
R552 vdd.n1825 vdd.n561 185
R553 vdd.n561 vdd.n523 185
R554 vdd.n1827 vdd.n1826 185
R555 vdd.n1828 vdd.n1827 185
R556 vdd.n562 vdd.n560 185
R557 vdd.n1766 vdd.n560 185
R558 vdd.n1756 vdd.n575 185
R559 vdd.n575 vdd.n567 185
R560 vdd.n1758 vdd.n1757 185
R561 vdd.n1759 vdd.n1758 185
R562 vdd.n1755 vdd.n574 185
R563 vdd.n574 vdd.n571 185
R564 vdd.n1754 vdd.n1753 185
R565 vdd.n1753 vdd.n1752 185
R566 vdd.n577 vdd.n576 185
R567 vdd.n578 vdd.n577 185
R568 vdd.n1745 vdd.n1744 185
R569 vdd.n1746 vdd.n1745 185
R570 vdd.n1743 vdd.n587 185
R571 vdd.n587 vdd.n584 185
R572 vdd.n1742 vdd.n1741 185
R573 vdd.n1741 vdd.n1740 185
R574 vdd.n589 vdd.n588 185
R575 vdd.n598 vdd.n589 185
R576 vdd.n1733 vdd.n1732 185
R577 vdd.n1734 vdd.n1733 185
R578 vdd.n1731 vdd.n599 185
R579 vdd.n599 vdd.n595 185
R580 vdd.n1730 vdd.n1729 185
R581 vdd.n1729 vdd.n1728 185
R582 vdd.n601 vdd.n600 185
R583 vdd.n1553 vdd.n601 185
R584 vdd.n1721 vdd.n1720 185
R585 vdd.n1722 vdd.n1721 185
R586 vdd.n1719 vdd.n610 185
R587 vdd.n610 vdd.n607 185
R588 vdd.n1718 vdd.n1717 185
R589 vdd.n1717 vdd.n1716 185
R590 vdd.n612 vdd.n611 185
R591 vdd.n1562 vdd.n612 185
R592 vdd.n1709 vdd.n1708 185
R593 vdd.n1710 vdd.n1709 185
R594 vdd.n1707 vdd.n621 185
R595 vdd.n621 vdd.n618 185
R596 vdd.n1706 vdd.n1705 185
R597 vdd.n1705 vdd.n1704 185
R598 vdd.n623 vdd.n622 185
R599 vdd.n624 vdd.n623 185
R600 vdd.n1697 vdd.n1696 185
R601 vdd.n1698 vdd.n1697 185
R602 vdd.n1695 vdd.n633 185
R603 vdd.n633 vdd.n630 185
R604 vdd.n1694 vdd.n1693 185
R605 vdd.n1693 vdd.n1692 185
R606 vdd.n635 vdd.n634 185
R607 vdd.n636 vdd.n635 185
R608 vdd.n1685 vdd.n1684 185
R609 vdd.n1686 vdd.n1685 185
R610 vdd.n1683 vdd.n645 185
R611 vdd.n645 vdd.n642 185
R612 vdd.n1682 vdd.n1681 185
R613 vdd.n1681 vdd.n1680 185
R614 vdd.n647 vdd.n646 185
R615 vdd.n648 vdd.n647 185
R616 vdd.n1673 vdd.n1672 185
R617 vdd.n1674 vdd.n1673 185
R618 vdd.n1671 vdd.n657 185
R619 vdd.n657 vdd.n654 185
R620 vdd.n1670 vdd.n1669 185
R621 vdd.n1669 vdd.n1668 185
R622 vdd.n659 vdd.n658 185
R623 vdd.n668 vdd.n659 185
R624 vdd.n1660 vdd.n1659 185
R625 vdd.n1661 vdd.n1660 185
R626 vdd.n1658 vdd.n669 185
R627 vdd.n675 vdd.n669 185
R628 vdd.n1657 vdd.n1656 185
R629 vdd.n1656 vdd.n1655 185
R630 vdd.n671 vdd.n670 185
R631 vdd.n672 vdd.n671 185
R632 vdd.n1648 vdd.n1647 185
R633 vdd.n1649 vdd.n1648 185
R634 vdd.n1646 vdd.n682 185
R635 vdd.n1645 vdd.n1644 185
R636 vdd.n1642 vdd.n683 185
R637 vdd.n1642 vdd.n679 185
R638 vdd.n1641 vdd.n1640 185
R639 vdd.n1639 vdd.n1638 185
R640 vdd.n1637 vdd.n685 185
R641 vdd.n1635 vdd.n1634 185
R642 vdd.n1633 vdd.n686 185
R643 vdd.n1632 vdd.n1631 185
R644 vdd.n1629 vdd.n687 185
R645 vdd.n1627 vdd.n1626 185
R646 vdd.n1625 vdd.n688 185
R647 vdd.n1624 vdd.n1623 185
R648 vdd.n1621 vdd.n1620 185
R649 vdd.n1619 vdd.n1618 185
R650 vdd.n1617 vdd.n691 185
R651 vdd.n1615 vdd.n1614 185
R652 vdd.n1613 vdd.n692 185
R653 vdd.n1612 vdd.n1611 185
R654 vdd.n1609 vdd.n693 185
R655 vdd.n1607 vdd.n1606 185
R656 vdd.n1605 vdd.n694 185
R657 vdd.n1604 vdd.n1603 185
R658 vdd.n1601 vdd.n1600 185
R659 vdd.n1599 vdd.n1598 185
R660 vdd.n1597 vdd.n1596 185
R661 vdd.n1597 vdd.n679 185
R662 vdd.n1773 vdd.n1772 185
R663 vdd.n1775 vdd.n1774 185
R664 vdd.n1777 vdd.n1776 185
R665 vdd.n1780 vdd.n1779 185
R666 vdd.n1782 vdd.n1781 185
R667 vdd.n1784 vdd.n1783 185
R668 vdd.n1786 vdd.n1785 185
R669 vdd.n1788 vdd.n1787 185
R670 vdd.n1790 vdd.n1789 185
R671 vdd.n1792 vdd.n1791 185
R672 vdd.n1794 vdd.n1793 185
R673 vdd.n1796 vdd.n1795 185
R674 vdd.n1798 vdd.n1797 185
R675 vdd.n1800 vdd.n1799 185
R676 vdd.n1802 vdd.n1801 185
R677 vdd.n1804 vdd.n1803 185
R678 vdd.n1806 vdd.n1805 185
R679 vdd.n1808 vdd.n1807 185
R680 vdd.n1810 vdd.n1809 185
R681 vdd.n1812 vdd.n1811 185
R682 vdd.n1814 vdd.n1813 185
R683 vdd.n1816 vdd.n1815 185
R684 vdd.n1818 vdd.n1817 185
R685 vdd.n1820 vdd.n1819 185
R686 vdd.n1822 vdd.n1821 185
R687 vdd.n1824 vdd.n1823 185
R688 vdd.n1771 vdd.n1770 185
R689 vdd.n1771 vdd.n523 185
R690 vdd.n1769 vdd.n558 185
R691 vdd.n1828 vdd.n558 185
R692 vdd.n1768 vdd.n1767 185
R693 vdd.n1767 vdd.n1766 185
R694 vdd.n566 vdd.n565 185
R695 vdd.n567 vdd.n566 185
R696 vdd.n1535 vdd.n572 185
R697 vdd.n1759 vdd.n572 185
R698 vdd.n1537 vdd.n1536 185
R699 vdd.n1536 vdd.n571 185
R700 vdd.n1538 vdd.n579 185
R701 vdd.n1752 vdd.n579 185
R702 vdd.n1540 vdd.n1539 185
R703 vdd.n1539 vdd.n578 185
R704 vdd.n1541 vdd.n585 185
R705 vdd.n1746 vdd.n585 185
R706 vdd.n1543 vdd.n1542 185
R707 vdd.n1542 vdd.n584 185
R708 vdd.n1544 vdd.n590 185
R709 vdd.n1740 vdd.n590 185
R710 vdd.n1546 vdd.n1545 185
R711 vdd.n1545 vdd.n598 185
R712 vdd.n1547 vdd.n596 185
R713 vdd.n1734 vdd.n596 185
R714 vdd.n1549 vdd.n1548 185
R715 vdd.n1548 vdd.n595 185
R716 vdd.n1550 vdd.n602 185
R717 vdd.n1728 vdd.n602 185
R718 vdd.n1552 vdd.n1551 185
R719 vdd.n1553 vdd.n1552 185
R720 vdd.n1534 vdd.n608 185
R721 vdd.n1722 vdd.n608 185
R722 vdd.n1533 vdd.n1532 185
R723 vdd.n1532 vdd.n607 185
R724 vdd.n699 vdd.n613 185
R725 vdd.n1716 vdd.n613 185
R726 vdd.n1564 vdd.n1563 185
R727 vdd.n1563 vdd.n1562 185
R728 vdd.n1565 vdd.n619 185
R729 vdd.n1710 vdd.n619 185
R730 vdd.n1567 vdd.n1566 185
R731 vdd.n1566 vdd.n618 185
R732 vdd.n1568 vdd.n625 185
R733 vdd.n1704 vdd.n625 185
R734 vdd.n1570 vdd.n1569 185
R735 vdd.n1569 vdd.n624 185
R736 vdd.n1571 vdd.n631 185
R737 vdd.n1698 vdd.n631 185
R738 vdd.n1573 vdd.n1572 185
R739 vdd.n1572 vdd.n630 185
R740 vdd.n1574 vdd.n637 185
R741 vdd.n1692 vdd.n637 185
R742 vdd.n1576 vdd.n1575 185
R743 vdd.n1575 vdd.n636 185
R744 vdd.n1577 vdd.n643 185
R745 vdd.n1686 vdd.n643 185
R746 vdd.n1579 vdd.n1578 185
R747 vdd.n1578 vdd.n642 185
R748 vdd.n1580 vdd.n649 185
R749 vdd.n1680 vdd.n649 185
R750 vdd.n1582 vdd.n1581 185
R751 vdd.n1581 vdd.n648 185
R752 vdd.n1583 vdd.n655 185
R753 vdd.n1674 vdd.n655 185
R754 vdd.n1585 vdd.n1584 185
R755 vdd.n1584 vdd.n654 185
R756 vdd.n1586 vdd.n660 185
R757 vdd.n1668 vdd.n660 185
R758 vdd.n1588 vdd.n1587 185
R759 vdd.n1587 vdd.n668 185
R760 vdd.n1589 vdd.n666 185
R761 vdd.n1661 vdd.n666 185
R762 vdd.n1591 vdd.n1590 185
R763 vdd.n1590 vdd.n675 185
R764 vdd.n1592 vdd.n673 185
R765 vdd.n1655 vdd.n673 185
R766 vdd.n1594 vdd.n1593 185
R767 vdd.n1593 vdd.n672 185
R768 vdd.n1595 vdd.n680 185
R769 vdd.n1649 vdd.n680 185
R770 vdd.n2710 vdd.n2709 185
R771 vdd.n2711 vdd.n2710 185
R772 vdd.n107 vdd.n106 185
R773 vdd.n2712 vdd.n107 185
R774 vdd.n2715 vdd.n2714 185
R775 vdd.n2714 vdd.n2713 185
R776 vdd.n2716 vdd.n101 185
R777 vdd.n101 vdd.n100 185
R778 vdd.n2718 vdd.n2717 185
R779 vdd.n2719 vdd.n2718 185
R780 vdd.n96 vdd.n95 185
R781 vdd.n2720 vdd.n96 185
R782 vdd.n2723 vdd.n2722 185
R783 vdd.n2722 vdd.n2721 185
R784 vdd.n2724 vdd.n90 185
R785 vdd.n90 vdd.n89 185
R786 vdd.n2726 vdd.n2725 185
R787 vdd.n2727 vdd.n2726 185
R788 vdd.n84 vdd.n83 185
R789 vdd.n2728 vdd.n84 185
R790 vdd.n2731 vdd.n2730 185
R791 vdd.n2730 vdd.n2729 185
R792 vdd.n2732 vdd.n78 185
R793 vdd.n85 vdd.n78 185
R794 vdd.n2734 vdd.n2733 185
R795 vdd.n2735 vdd.n2734 185
R796 vdd.n74 vdd.n73 185
R797 vdd.n2736 vdd.n74 185
R798 vdd.n2739 vdd.n2738 185
R799 vdd.n2738 vdd.n2737 185
R800 vdd.n2740 vdd.n69 185
R801 vdd.n69 vdd.n68 185
R802 vdd.n2742 vdd.n2741 185
R803 vdd.n2743 vdd.n2742 185
R804 vdd.n63 vdd.n61 185
R805 vdd.n2744 vdd.n63 185
R806 vdd.n2747 vdd.n2746 185
R807 vdd.n2746 vdd.n2745 185
R808 vdd.n62 vdd.n60 185
R809 vdd.n64 vdd.n62 185
R810 vdd.n2566 vdd.n2565 185
R811 vdd.n2567 vdd.n2566 185
R812 vdd.n236 vdd.n235 185
R813 vdd.n235 vdd.n234 185
R814 vdd.n2561 vdd.n2560 185
R815 vdd.n2560 vdd.n2559 185
R816 vdd.n239 vdd.n238 185
R817 vdd.n246 vdd.n239 185
R818 vdd.n2550 vdd.n2549 185
R819 vdd.n2551 vdd.n2550 185
R820 vdd.n248 vdd.n247 185
R821 vdd.n247 vdd.n245 185
R822 vdd.n2545 vdd.n2544 185
R823 vdd.n2544 vdd.n2543 185
R824 vdd.n251 vdd.n250 185
R825 vdd.n252 vdd.n251 185
R826 vdd.n2534 vdd.n2533 185
R827 vdd.n2535 vdd.n2534 185
R828 vdd.n260 vdd.n259 185
R829 vdd.n259 vdd.n258 185
R830 vdd.n2529 vdd.n2528 185
R831 vdd.n2528 vdd.n2527 185
R832 vdd.n263 vdd.n262 185
R833 vdd.n270 vdd.n263 185
R834 vdd.n2518 vdd.n2517 185
R835 vdd.n2519 vdd.n2518 185
R836 vdd.n272 vdd.n271 185
R837 vdd.n271 vdd.n269 185
R838 vdd.n2513 vdd.n2512 185
R839 vdd.n2512 vdd.n2511 185
R840 vdd.n275 vdd.n274 185
R841 vdd.n276 vdd.n275 185
R842 vdd.n2502 vdd.n2501 185
R843 vdd.n2503 vdd.n2502 185
R844 vdd.n284 vdd.n283 185
R845 vdd.n283 vdd.n282 185
R846 vdd.n2497 vdd.n2496 185
R847 vdd.n287 vdd.n286 185
R848 vdd.n2493 vdd.n2492 185
R849 vdd.n2494 vdd.n2493 185
R850 vdd.n2491 vdd.n317 185
R851 vdd.n2490 vdd.n2489 185
R852 vdd.n2488 vdd.n2487 185
R853 vdd.n324 vdd.n321 185
R854 vdd.n326 vdd.n325 185
R855 vdd.n2483 vdd.n327 185
R856 vdd.n2482 vdd.n2481 185
R857 vdd.n2480 vdd.n2479 185
R858 vdd.n2478 vdd.n2477 185
R859 vdd.n2476 vdd.n2475 185
R860 vdd.n2474 vdd.n2473 185
R861 vdd.n2472 vdd.n2471 185
R862 vdd.n2470 vdd.n2469 185
R863 vdd.n2468 vdd.n2467 185
R864 vdd.n2466 vdd.n2465 185
R865 vdd.n2457 vdd.n335 185
R866 vdd.n2459 vdd.n2458 185
R867 vdd.n2456 vdd.n2455 185
R868 vdd.n2454 vdd.n2453 185
R869 vdd.n2452 vdd.n2451 185
R870 vdd.n2450 vdd.n2449 185
R871 vdd.n2448 vdd.n2447 185
R872 vdd.n2446 vdd.n2445 185
R873 vdd.n2444 vdd.n2443 185
R874 vdd.n2442 vdd.n2441 185
R875 vdd.n2440 vdd.n2439 185
R876 vdd.n2438 vdd.n2437 185
R877 vdd.n2436 vdd.n2435 185
R878 vdd.n2434 vdd.n2433 185
R879 vdd.n2432 vdd.n2431 185
R880 vdd.n2430 vdd.n2429 185
R881 vdd.n2428 vdd.n2427 185
R882 vdd.n2426 vdd.n2425 185
R883 vdd.n2424 vdd.n2423 185
R884 vdd.n2422 vdd.n2421 185
R885 vdd.n2415 vdd.n353 185
R886 vdd.n2417 vdd.n2416 185
R887 vdd.n2414 vdd.n2413 185
R888 vdd.n2412 vdd.n2411 185
R889 vdd.n2410 vdd.n2409 185
R890 vdd.n2408 vdd.n2407 185
R891 vdd.n2406 vdd.n2405 185
R892 vdd.n2404 vdd.n2403 185
R893 vdd.n2402 vdd.n2401 185
R894 vdd.n2400 vdd.n2399 185
R895 vdd.n2398 vdd.n2397 185
R896 vdd.n2396 vdd.n2395 185
R897 vdd.n2371 vdd.n365 185
R898 vdd.n2373 vdd.n2372 185
R899 vdd.n2391 vdd.n2374 185
R900 vdd.n2390 vdd.n2389 185
R901 vdd.n2388 vdd.n2387 185
R902 vdd.n2386 vdd.n2385 185
R903 vdd.n2384 vdd.n2383 185
R904 vdd.n2379 vdd.n316 185
R905 vdd.n2494 vdd.n316 185
R906 vdd.n2603 vdd.n2602 185
R907 vdd.n2605 vdd.n210 185
R908 vdd.n2607 vdd.n2606 185
R909 vdd.n2608 vdd.n205 185
R910 vdd.n2610 vdd.n2609 185
R911 vdd.n2612 vdd.n203 185
R912 vdd.n2614 vdd.n2613 185
R913 vdd.n2615 vdd.n198 185
R914 vdd.n2617 vdd.n2616 185
R915 vdd.n2619 vdd.n196 185
R916 vdd.n2621 vdd.n2620 185
R917 vdd.n2622 vdd.n191 185
R918 vdd.n2624 vdd.n2623 185
R919 vdd.n2626 vdd.n189 185
R920 vdd.n2628 vdd.n2627 185
R921 vdd.n2629 vdd.n185 185
R922 vdd.n2631 vdd.n2630 185
R923 vdd.n2633 vdd.n183 185
R924 vdd.n2635 vdd.n2634 185
R925 vdd.n178 vdd.n177 185
R926 vdd.n2640 vdd.n2639 185
R927 vdd.n2642 vdd.n175 185
R928 vdd.n2644 vdd.n2643 185
R929 vdd.n2645 vdd.n170 185
R930 vdd.n2647 vdd.n2646 185
R931 vdd.n2649 vdd.n168 185
R932 vdd.n2651 vdd.n2650 185
R933 vdd.n2652 vdd.n163 185
R934 vdd.n2654 vdd.n2653 185
R935 vdd.n2656 vdd.n161 185
R936 vdd.n2658 vdd.n2657 185
R937 vdd.n2659 vdd.n156 185
R938 vdd.n2661 vdd.n2660 185
R939 vdd.n2663 vdd.n154 185
R940 vdd.n2665 vdd.n2664 185
R941 vdd.n2666 vdd.n150 185
R942 vdd.n2668 vdd.n2667 185
R943 vdd.n2670 vdd.n148 185
R944 vdd.n2672 vdd.n2671 185
R945 vdd.n143 vdd.n142 185
R946 vdd.n2677 vdd.n2676 185
R947 vdd.n2679 vdd.n140 185
R948 vdd.n2681 vdd.n2680 185
R949 vdd.n2682 vdd.n135 185
R950 vdd.n2684 vdd.n2683 185
R951 vdd.n2686 vdd.n133 185
R952 vdd.n2688 vdd.n2687 185
R953 vdd.n2689 vdd.n128 185
R954 vdd.n2691 vdd.n2690 185
R955 vdd.n2693 vdd.n126 185
R956 vdd.n2695 vdd.n2694 185
R957 vdd.n2696 vdd.n120 185
R958 vdd.n2698 vdd.n2697 185
R959 vdd.n2700 vdd.n119 185
R960 vdd.n2701 vdd.n118 185
R961 vdd.n2704 vdd.n2703 185
R962 vdd.n2705 vdd.n116 185
R963 vdd.n2706 vdd.n112 185
R964 vdd.n2599 vdd.n110 185
R965 vdd.n2711 vdd.n110 185
R966 vdd.n2598 vdd.n109 185
R967 vdd.n2712 vdd.n109 185
R968 vdd.n2597 vdd.n108 185
R969 vdd.n2713 vdd.n108 185
R970 vdd.n218 vdd.n217 185
R971 vdd.n217 vdd.n100 185
R972 vdd.n2593 vdd.n99 185
R973 vdd.n2719 vdd.n99 185
R974 vdd.n2592 vdd.n98 185
R975 vdd.n2720 vdd.n98 185
R976 vdd.n2591 vdd.n97 185
R977 vdd.n2721 vdd.n97 185
R978 vdd.n221 vdd.n220 185
R979 vdd.n220 vdd.n89 185
R980 vdd.n2587 vdd.n88 185
R981 vdd.n2727 vdd.n88 185
R982 vdd.n2586 vdd.n87 185
R983 vdd.n2728 vdd.n87 185
R984 vdd.n2585 vdd.n86 185
R985 vdd.n2729 vdd.n86 185
R986 vdd.n224 vdd.n223 185
R987 vdd.n223 vdd.n85 185
R988 vdd.n2581 vdd.n77 185
R989 vdd.n2735 vdd.n77 185
R990 vdd.n2580 vdd.n76 185
R991 vdd.n2736 vdd.n76 185
R992 vdd.n2579 vdd.n75 185
R993 vdd.n2737 vdd.n75 185
R994 vdd.n227 vdd.n226 185
R995 vdd.n226 vdd.n68 185
R996 vdd.n2575 vdd.n67 185
R997 vdd.n2743 vdd.n67 185
R998 vdd.n2574 vdd.n66 185
R999 vdd.n2744 vdd.n66 185
R1000 vdd.n2573 vdd.n65 185
R1001 vdd.n2745 vdd.n65 185
R1002 vdd.n233 vdd.n229 185
R1003 vdd.n233 vdd.n64 185
R1004 vdd.n2569 vdd.n2568 185
R1005 vdd.n2568 vdd.n2567 185
R1006 vdd.n232 vdd.n231 185
R1007 vdd.n234 vdd.n232 185
R1008 vdd.n2558 vdd.n2557 185
R1009 vdd.n2559 vdd.n2558 185
R1010 vdd.n241 vdd.n240 185
R1011 vdd.n246 vdd.n240 185
R1012 vdd.n2553 vdd.n2552 185
R1013 vdd.n2552 vdd.n2551 185
R1014 vdd.n244 vdd.n243 185
R1015 vdd.n245 vdd.n244 185
R1016 vdd.n2542 vdd.n2541 185
R1017 vdd.n2543 vdd.n2542 185
R1018 vdd.n254 vdd.n253 185
R1019 vdd.n253 vdd.n252 185
R1020 vdd.n2537 vdd.n2536 185
R1021 vdd.n2536 vdd.n2535 185
R1022 vdd.n257 vdd.n256 185
R1023 vdd.n258 vdd.n257 185
R1024 vdd.n2526 vdd.n2525 185
R1025 vdd.n2527 vdd.n2526 185
R1026 vdd.n265 vdd.n264 185
R1027 vdd.n270 vdd.n264 185
R1028 vdd.n2521 vdd.n2520 185
R1029 vdd.n2520 vdd.n2519 185
R1030 vdd.n268 vdd.n267 185
R1031 vdd.n269 vdd.n268 185
R1032 vdd.n2510 vdd.n2509 185
R1033 vdd.n2511 vdd.n2510 185
R1034 vdd.n278 vdd.n277 185
R1035 vdd.n277 vdd.n276 185
R1036 vdd.n2505 vdd.n2504 185
R1037 vdd.n2504 vdd.n2503 185
R1038 vdd.n281 vdd.n280 185
R1039 vdd.n282 vdd.n281 185
R1040 vdd.n522 vdd.n521 185
R1041 vdd.n1920 vdd.n1919 185
R1042 vdd.n1921 vdd.n1917 185
R1043 vdd.n1917 vdd.n1883 185
R1044 vdd.n1923 vdd.n1922 185
R1045 vdd.n1925 vdd.n1916 185
R1046 vdd.n1928 vdd.n1927 185
R1047 vdd.n1929 vdd.n1915 185
R1048 vdd.n1931 vdd.n1930 185
R1049 vdd.n1933 vdd.n1914 185
R1050 vdd.n1936 vdd.n1935 185
R1051 vdd.n1937 vdd.n1913 185
R1052 vdd.n1939 vdd.n1938 185
R1053 vdd.n1941 vdd.n1912 185
R1054 vdd.n1944 vdd.n1943 185
R1055 vdd.n1945 vdd.n1911 185
R1056 vdd.n1947 vdd.n1946 185
R1057 vdd.n1949 vdd.n1910 185
R1058 vdd.n1952 vdd.n1951 185
R1059 vdd.n1953 vdd.n1909 185
R1060 vdd.n1955 vdd.n1954 185
R1061 vdd.n1957 vdd.n1908 185
R1062 vdd.n1960 vdd.n1959 185
R1063 vdd.n1961 vdd.n1905 185
R1064 vdd.n1964 vdd.n1963 185
R1065 vdd.n1966 vdd.n1904 185
R1066 vdd.n1968 vdd.n1967 185
R1067 vdd.n1967 vdd.n1883 185
R1068 vdd.n2296 vdd.n2295 185
R1069 vdd.n2298 vdd.n406 185
R1070 vdd.n2300 vdd.n2299 185
R1071 vdd.n2302 vdd.n403 185
R1072 vdd.n2304 vdd.n2303 185
R1073 vdd.n2306 vdd.n401 185
R1074 vdd.n2308 vdd.n2307 185
R1075 vdd.n2309 vdd.n400 185
R1076 vdd.n2311 vdd.n2310 185
R1077 vdd.n2313 vdd.n398 185
R1078 vdd.n2315 vdd.n2314 185
R1079 vdd.n2316 vdd.n397 185
R1080 vdd.n2318 vdd.n2317 185
R1081 vdd.n2321 vdd.n2320 185
R1082 vdd.n2323 vdd.n2322 185
R1083 vdd.n2325 vdd.n395 185
R1084 vdd.n2327 vdd.n2326 185
R1085 vdd.n2328 vdd.n394 185
R1086 vdd.n2330 vdd.n2329 185
R1087 vdd.n2332 vdd.n392 185
R1088 vdd.n2334 vdd.n2333 185
R1089 vdd.n2335 vdd.n391 185
R1090 vdd.n2337 vdd.n2336 185
R1091 vdd.n2339 vdd.n389 185
R1092 vdd.n2341 vdd.n2340 185
R1093 vdd.n2342 vdd.n387 185
R1094 vdd.n2294 vdd.n384 185
R1095 vdd.n2345 vdd.n384 185
R1096 vdd.n2293 vdd.n2292 185
R1097 vdd.n2292 vdd.n383 185
R1098 vdd.n2291 vdd.n408 185
R1099 vdd.n2291 vdd.n2290 185
R1100 vdd.n1991 vdd.n409 185
R1101 vdd.n410 vdd.n409 185
R1102 vdd.n1992 vdd.n417 185
R1103 vdd.n2284 vdd.n417 185
R1104 vdd.n1994 vdd.n1993 185
R1105 vdd.n1993 vdd.n416 185
R1106 vdd.n1995 vdd.n425 185
R1107 vdd.n2241 vdd.n425 185
R1108 vdd.n1997 vdd.n1996 185
R1109 vdd.n1996 vdd.n424 185
R1110 vdd.n1998 vdd.n431 185
R1111 vdd.n2235 vdd.n431 185
R1112 vdd.n2000 vdd.n1999 185
R1113 vdd.n1999 vdd.n430 185
R1114 vdd.n2001 vdd.n436 185
R1115 vdd.n2229 vdd.n436 185
R1116 vdd.n2003 vdd.n2002 185
R1117 vdd.n2002 vdd.n443 185
R1118 vdd.n2004 vdd.n441 185
R1119 vdd.n2223 vdd.n441 185
R1120 vdd.n2006 vdd.n2005 185
R1121 vdd.n2005 vdd.n449 185
R1122 vdd.n2007 vdd.n447 185
R1123 vdd.n2217 vdd.n447 185
R1124 vdd.n2009 vdd.n2008 185
R1125 vdd.n2008 vdd.n455 185
R1126 vdd.n2010 vdd.n453 185
R1127 vdd.n2211 vdd.n453 185
R1128 vdd.n2012 vdd.n2011 185
R1129 vdd.n2011 vdd.n461 185
R1130 vdd.n2013 vdd.n459 185
R1131 vdd.n2205 vdd.n459 185
R1132 vdd.n2015 vdd.n2014 185
R1133 vdd.n2014 vdd.n467 185
R1134 vdd.n2016 vdd.n465 185
R1135 vdd.n2199 vdd.n465 185
R1136 vdd.n2053 vdd.n2052 185
R1137 vdd.n2052 vdd.n2051 185
R1138 vdd.n2054 vdd.n472 185
R1139 vdd.n2193 vdd.n472 185
R1140 vdd.n2056 vdd.n2055 185
R1141 vdd.n2055 vdd.n471 185
R1142 vdd.n2057 vdd.n477 185
R1143 vdd.n2187 vdd.n477 185
R1144 vdd.n2059 vdd.n2058 185
R1145 vdd.n2060 vdd.n2059 185
R1146 vdd.n1990 vdd.n483 185
R1147 vdd.n2181 vdd.n483 185
R1148 vdd.n1989 vdd.n1988 185
R1149 vdd.n1988 vdd.n482 185
R1150 vdd.n1987 vdd.n489 185
R1151 vdd.n2175 vdd.n489 185
R1152 vdd.n1986 vdd.n1985 185
R1153 vdd.n1985 vdd.n488 185
R1154 vdd.n1984 vdd.n494 185
R1155 vdd.n2169 vdd.n494 185
R1156 vdd.n1983 vdd.n1982 185
R1157 vdd.n1982 vdd.n502 185
R1158 vdd.n1981 vdd.n500 185
R1159 vdd.n2163 vdd.n500 185
R1160 vdd.n1980 vdd.n1979 185
R1161 vdd.n1979 vdd.n499 185
R1162 vdd.n1978 vdd.n506 185
R1163 vdd.n2157 vdd.n506 185
R1164 vdd.n1977 vdd.n1976 185
R1165 vdd.n1976 vdd.n513 185
R1166 vdd.n1975 vdd.n511 185
R1167 vdd.n2151 vdd.n511 185
R1168 vdd.n1974 vdd.n1973 185
R1169 vdd.n1973 vdd.n519 185
R1170 vdd.n1972 vdd.n517 185
R1171 vdd.n2145 vdd.n517 185
R1172 vdd.n1971 vdd.n1970 185
R1173 vdd.n1970 vdd.n1886 185
R1174 vdd.n1969 vdd.n1884 185
R1175 vdd.n2139 vdd.n1884 185
R1176 vdd.n2141 vdd.n2140 185
R1177 vdd.n2140 vdd.n2139 185
R1178 vdd.n2142 vdd.n520 185
R1179 vdd.n1886 vdd.n520 185
R1180 vdd.n2144 vdd.n2143 185
R1181 vdd.n2145 vdd.n2144 185
R1182 vdd.n510 vdd.n509 185
R1183 vdd.n519 vdd.n510 185
R1184 vdd.n2153 vdd.n2152 185
R1185 vdd.n2152 vdd.n2151 185
R1186 vdd.n2154 vdd.n508 185
R1187 vdd.n513 vdd.n508 185
R1188 vdd.n2156 vdd.n2155 185
R1189 vdd.n2157 vdd.n2156 185
R1190 vdd.n498 vdd.n497 185
R1191 vdd.n499 vdd.n498 185
R1192 vdd.n2165 vdd.n2164 185
R1193 vdd.n2164 vdd.n2163 185
R1194 vdd.n2166 vdd.n496 185
R1195 vdd.n502 vdd.n496 185
R1196 vdd.n2168 vdd.n2167 185
R1197 vdd.n2169 vdd.n2168 185
R1198 vdd.n487 vdd.n486 185
R1199 vdd.n488 vdd.n487 185
R1200 vdd.n2177 vdd.n2176 185
R1201 vdd.n2176 vdd.n2175 185
R1202 vdd.n2178 vdd.n485 185
R1203 vdd.n485 vdd.n482 185
R1204 vdd.n2180 vdd.n2179 185
R1205 vdd.n2181 vdd.n2180 185
R1206 vdd.n476 vdd.n475 185
R1207 vdd.n2060 vdd.n476 185
R1208 vdd.n2189 vdd.n2188 185
R1209 vdd.n2188 vdd.n2187 185
R1210 vdd.n2190 vdd.n474 185
R1211 vdd.n474 vdd.n471 185
R1212 vdd.n2192 vdd.n2191 185
R1213 vdd.n2193 vdd.n2192 185
R1214 vdd.n464 vdd.n463 185
R1215 vdd.n2051 vdd.n464 185
R1216 vdd.n2201 vdd.n2200 185
R1217 vdd.n2200 vdd.n2199 185
R1218 vdd.n2202 vdd.n462 185
R1219 vdd.n467 vdd.n462 185
R1220 vdd.n2204 vdd.n2203 185
R1221 vdd.n2205 vdd.n2204 185
R1222 vdd.n452 vdd.n451 185
R1223 vdd.n461 vdd.n452 185
R1224 vdd.n2213 vdd.n2212 185
R1225 vdd.n2212 vdd.n2211 185
R1226 vdd.n2214 vdd.n450 185
R1227 vdd.n455 vdd.n450 185
R1228 vdd.n2216 vdd.n2215 185
R1229 vdd.n2217 vdd.n2216 185
R1230 vdd.n440 vdd.n439 185
R1231 vdd.n449 vdd.n440 185
R1232 vdd.n2225 vdd.n2224 185
R1233 vdd.n2224 vdd.n2223 185
R1234 vdd.n2226 vdd.n438 185
R1235 vdd.n443 vdd.n438 185
R1236 vdd.n2228 vdd.n2227 185
R1237 vdd.n2229 vdd.n2228 185
R1238 vdd.n429 vdd.n428 185
R1239 vdd.n430 vdd.n429 185
R1240 vdd.n2237 vdd.n2236 185
R1241 vdd.n2236 vdd.n2235 185
R1242 vdd.n2238 vdd.n427 185
R1243 vdd.n427 vdd.n424 185
R1244 vdd.n2240 vdd.n2239 185
R1245 vdd.n2241 vdd.n2240 185
R1246 vdd.n415 vdd.n414 185
R1247 vdd.n416 vdd.n415 185
R1248 vdd.n2286 vdd.n2285 185
R1249 vdd.n2285 vdd.n2284 185
R1250 vdd.n2287 vdd.n413 185
R1251 vdd.n413 vdd.n410 185
R1252 vdd.n2289 vdd.n2288 185
R1253 vdd.n2290 vdd.n2289 185
R1254 vdd.n388 vdd.n386 185
R1255 vdd.n386 vdd.n383 185
R1256 vdd.n2344 vdd.n2343 185
R1257 vdd.n2345 vdd.n2344 185
R1258 vdd.n552 vdd.n550 185
R1259 vdd.n550 vdd.n523 185
R1260 vdd.n1763 vdd.n559 185
R1261 vdd.n1828 vdd.n559 185
R1262 vdd.n1765 vdd.n1764 185
R1263 vdd.n1766 vdd.n1765 185
R1264 vdd.n1762 vdd.n568 185
R1265 vdd.n568 vdd.n567 185
R1266 vdd.n1761 vdd.n1760 185
R1267 vdd.n1760 vdd.n1759 185
R1268 vdd.n570 vdd.n569 185
R1269 vdd.n571 vdd.n570 185
R1270 vdd.n1751 vdd.n1750 185
R1271 vdd.n1752 vdd.n1751 185
R1272 vdd.n1749 vdd.n581 185
R1273 vdd.n581 vdd.n578 185
R1274 vdd.n1748 vdd.n1747 185
R1275 vdd.n1747 vdd.n1746 185
R1276 vdd.n583 vdd.n582 185
R1277 vdd.n584 vdd.n583 185
R1278 vdd.n1739 vdd.n1738 185
R1279 vdd.n1740 vdd.n1739 185
R1280 vdd.n1737 vdd.n592 185
R1281 vdd.n598 vdd.n592 185
R1282 vdd.n1736 vdd.n1735 185
R1283 vdd.n1735 vdd.n1734 185
R1284 vdd.n594 vdd.n593 185
R1285 vdd.n595 vdd.n594 185
R1286 vdd.n1727 vdd.n1726 185
R1287 vdd.n1728 vdd.n1727 185
R1288 vdd.n1725 vdd.n604 185
R1289 vdd.n1553 vdd.n604 185
R1290 vdd.n1724 vdd.n1723 185
R1291 vdd.n1723 vdd.n1722 185
R1292 vdd.n606 vdd.n605 185
R1293 vdd.n607 vdd.n606 185
R1294 vdd.n1715 vdd.n1714 185
R1295 vdd.n1716 vdd.n1715 185
R1296 vdd.n1713 vdd.n615 185
R1297 vdd.n1562 vdd.n615 185
R1298 vdd.n1712 vdd.n1711 185
R1299 vdd.n1711 vdd.n1710 185
R1300 vdd.n617 vdd.n616 185
R1301 vdd.n618 vdd.n617 185
R1302 vdd.n1703 vdd.n1702 185
R1303 vdd.n1704 vdd.n1703 185
R1304 vdd.n1701 vdd.n627 185
R1305 vdd.n627 vdd.n624 185
R1306 vdd.n1700 vdd.n1699 185
R1307 vdd.n1699 vdd.n1698 185
R1308 vdd.n629 vdd.n628 185
R1309 vdd.n630 vdd.n629 185
R1310 vdd.n1691 vdd.n1690 185
R1311 vdd.n1692 vdd.n1691 185
R1312 vdd.n1689 vdd.n639 185
R1313 vdd.n639 vdd.n636 185
R1314 vdd.n1688 vdd.n1687 185
R1315 vdd.n1687 vdd.n1686 185
R1316 vdd.n641 vdd.n640 185
R1317 vdd.n642 vdd.n641 185
R1318 vdd.n1679 vdd.n1678 185
R1319 vdd.n1680 vdd.n1679 185
R1320 vdd.n1677 vdd.n651 185
R1321 vdd.n651 vdd.n648 185
R1322 vdd.n1676 vdd.n1675 185
R1323 vdd.n1675 vdd.n1674 185
R1324 vdd.n653 vdd.n652 185
R1325 vdd.n654 vdd.n653 185
R1326 vdd.n1667 vdd.n1666 185
R1327 vdd.n1668 vdd.n1667 185
R1328 vdd.n1664 vdd.n662 185
R1329 vdd.n668 vdd.n662 185
R1330 vdd.n1663 vdd.n1662 185
R1331 vdd.n1662 vdd.n1661 185
R1332 vdd.n665 vdd.n664 185
R1333 vdd.n675 vdd.n665 185
R1334 vdd.n1654 vdd.n1653 185
R1335 vdd.n1655 vdd.n1654 185
R1336 vdd.n1652 vdd.n676 185
R1337 vdd.n676 vdd.n672 185
R1338 vdd.n1651 vdd.n1650 185
R1339 vdd.n1650 vdd.n1649 185
R1340 vdd.n1832 vdd.n549 185
R1341 vdd.n1882 vdd.n549 185
R1342 vdd.n1834 vdd.n1833 185
R1343 vdd.n1836 vdd.n1835 185
R1344 vdd.n1838 vdd.n1837 185
R1345 vdd.n1840 vdd.n1839 185
R1346 vdd.n1842 vdd.n1841 185
R1347 vdd.n1844 vdd.n1843 185
R1348 vdd.n1846 vdd.n1845 185
R1349 vdd.n1848 vdd.n1847 185
R1350 vdd.n1850 vdd.n1849 185
R1351 vdd.n1852 vdd.n1851 185
R1352 vdd.n1854 vdd.n1853 185
R1353 vdd.n1856 vdd.n1855 185
R1354 vdd.n1858 vdd.n1857 185
R1355 vdd.n1860 vdd.n1859 185
R1356 vdd.n1862 vdd.n1861 185
R1357 vdd.n1864 vdd.n1863 185
R1358 vdd.n1866 vdd.n1865 185
R1359 vdd.n1868 vdd.n1867 185
R1360 vdd.n1870 vdd.n1869 185
R1361 vdd.n1872 vdd.n1871 185
R1362 vdd.n1874 vdd.n1873 185
R1363 vdd.n1876 vdd.n1875 185
R1364 vdd.n1878 vdd.n1877 185
R1365 vdd.n1879 vdd.n551 185
R1366 vdd.n1881 vdd.n1880 185
R1367 vdd.n1882 vdd.n1881 185
R1368 vdd.n1831 vdd.n1830 185
R1369 vdd.n1830 vdd.n523 185
R1370 vdd.n1829 vdd.n556 185
R1371 vdd.n1829 vdd.n1828 185
R1372 vdd.n1513 vdd.n557 185
R1373 vdd.n1766 vdd.n557 185
R1374 vdd.n1515 vdd.n1514 185
R1375 vdd.n1514 vdd.n567 185
R1376 vdd.n1516 vdd.n573 185
R1377 vdd.n1759 vdd.n573 185
R1378 vdd.n1518 vdd.n1517 185
R1379 vdd.n1517 vdd.n571 185
R1380 vdd.n1519 vdd.n580 185
R1381 vdd.n1752 vdd.n580 185
R1382 vdd.n1521 vdd.n1520 185
R1383 vdd.n1520 vdd.n578 185
R1384 vdd.n1522 vdd.n586 185
R1385 vdd.n1746 vdd.n586 185
R1386 vdd.n1524 vdd.n1523 185
R1387 vdd.n1523 vdd.n584 185
R1388 vdd.n1525 vdd.n591 185
R1389 vdd.n1740 vdd.n591 185
R1390 vdd.n1527 vdd.n1526 185
R1391 vdd.n1526 vdd.n598 185
R1392 vdd.n1528 vdd.n597 185
R1393 vdd.n1734 vdd.n597 185
R1394 vdd.n1530 vdd.n1529 185
R1395 vdd.n1529 vdd.n595 185
R1396 vdd.n1531 vdd.n603 185
R1397 vdd.n1728 vdd.n603 185
R1398 vdd.n1555 vdd.n1554 185
R1399 vdd.n1554 vdd.n1553 185
R1400 vdd.n1556 vdd.n609 185
R1401 vdd.n1722 vdd.n609 185
R1402 vdd.n1558 vdd.n1557 185
R1403 vdd.n1557 vdd.n607 185
R1404 vdd.n1559 vdd.n614 185
R1405 vdd.n1716 vdd.n614 185
R1406 vdd.n1561 vdd.n1560 185
R1407 vdd.n1562 vdd.n1561 185
R1408 vdd.n1512 vdd.n620 185
R1409 vdd.n1710 vdd.n620 185
R1410 vdd.n1511 vdd.n1510 185
R1411 vdd.n1510 vdd.n618 185
R1412 vdd.n1509 vdd.n626 185
R1413 vdd.n1704 vdd.n626 185
R1414 vdd.n1508 vdd.n1507 185
R1415 vdd.n1507 vdd.n624 185
R1416 vdd.n1506 vdd.n632 185
R1417 vdd.n1698 vdd.n632 185
R1418 vdd.n1505 vdd.n1504 185
R1419 vdd.n1504 vdd.n630 185
R1420 vdd.n1503 vdd.n638 185
R1421 vdd.n1692 vdd.n638 185
R1422 vdd.n1502 vdd.n1501 185
R1423 vdd.n1501 vdd.n636 185
R1424 vdd.n1500 vdd.n644 185
R1425 vdd.n1686 vdd.n644 185
R1426 vdd.n1499 vdd.n1498 185
R1427 vdd.n1498 vdd.n642 185
R1428 vdd.n1497 vdd.n650 185
R1429 vdd.n1680 vdd.n650 185
R1430 vdd.n1496 vdd.n1495 185
R1431 vdd.n1495 vdd.n648 185
R1432 vdd.n1494 vdd.n656 185
R1433 vdd.n1674 vdd.n656 185
R1434 vdd.n1493 vdd.n1492 185
R1435 vdd.n1492 vdd.n654 185
R1436 vdd.n1491 vdd.n661 185
R1437 vdd.n1668 vdd.n661 185
R1438 vdd.n1490 vdd.n1489 185
R1439 vdd.n1489 vdd.n668 185
R1440 vdd.n1488 vdd.n667 185
R1441 vdd.n1661 vdd.n667 185
R1442 vdd.n1487 vdd.n1486 185
R1443 vdd.n1486 vdd.n675 185
R1444 vdd.n1485 vdd.n674 185
R1445 vdd.n1655 vdd.n674 185
R1446 vdd.n1484 vdd.n1483 185
R1447 vdd.n1483 vdd.n672 185
R1448 vdd.n1482 vdd.n681 185
R1449 vdd.n1649 vdd.n681 185
R1450 vdd.n678 vdd.n677 185
R1451 vdd.n679 vdd.n678 185
R1452 vdd.n1433 vdd.n1432 185
R1453 vdd.n1434 vdd.n1430 185
R1454 vdd.n1436 vdd.n1435 185
R1455 vdd.n1438 vdd.n1429 185
R1456 vdd.n1441 vdd.n1440 185
R1457 vdd.n1442 vdd.n1428 185
R1458 vdd.n1444 vdd.n1443 185
R1459 vdd.n1446 vdd.n1427 185
R1460 vdd.n1449 vdd.n1448 185
R1461 vdd.n1450 vdd.n1426 185
R1462 vdd.n1452 vdd.n1451 185
R1463 vdd.n1454 vdd.n1425 185
R1464 vdd.n1457 vdd.n1456 185
R1465 vdd.n1458 vdd.n707 185
R1466 vdd.n1460 vdd.n1459 185
R1467 vdd.n1462 vdd.n706 185
R1468 vdd.n1465 vdd.n1464 185
R1469 vdd.n1466 vdd.n705 185
R1470 vdd.n1468 vdd.n1467 185
R1471 vdd.n1470 vdd.n704 185
R1472 vdd.n1473 vdd.n1472 185
R1473 vdd.n1474 vdd.n701 185
R1474 vdd.n1477 vdd.n1476 185
R1475 vdd.n1479 vdd.n700 185
R1476 vdd.n1481 vdd.n1480 185
R1477 vdd.n1480 vdd.n679 185
R1478 vdd.n727 vdd.n679 151.596
R1479 vdd.n2494 vdd.n288 151.596
R1480 vdd.n2703 vdd.n116 146.341
R1481 vdd.n2701 vdd.n2700 146.341
R1482 vdd.n2698 vdd.n120 146.341
R1483 vdd.n2694 vdd.n2693 146.341
R1484 vdd.n2691 vdd.n128 146.341
R1485 vdd.n2687 vdd.n2686 146.341
R1486 vdd.n2684 vdd.n135 146.341
R1487 vdd.n2680 vdd.n2679 146.341
R1488 vdd.n2677 vdd.n142 146.341
R1489 vdd.n2671 vdd.n2670 146.341
R1490 vdd.n2668 vdd.n150 146.341
R1491 vdd.n2664 vdd.n2663 146.341
R1492 vdd.n2661 vdd.n156 146.341
R1493 vdd.n2657 vdd.n2656 146.341
R1494 vdd.n2654 vdd.n163 146.341
R1495 vdd.n2650 vdd.n2649 146.341
R1496 vdd.n2647 vdd.n170 146.341
R1497 vdd.n2643 vdd.n2642 146.341
R1498 vdd.n2640 vdd.n177 146.341
R1499 vdd.n2634 vdd.n2633 146.341
R1500 vdd.n2631 vdd.n185 146.341
R1501 vdd.n2627 vdd.n2626 146.341
R1502 vdd.n2624 vdd.n191 146.341
R1503 vdd.n2620 vdd.n2619 146.341
R1504 vdd.n2617 vdd.n198 146.341
R1505 vdd.n2613 vdd.n2612 146.341
R1506 vdd.n2610 vdd.n205 146.341
R1507 vdd.n2606 vdd.n2605 146.341
R1508 vdd.n2504 vdd.n281 146.341
R1509 vdd.n2504 vdd.n277 146.341
R1510 vdd.n2510 vdd.n277 146.341
R1511 vdd.n2510 vdd.n268 146.341
R1512 vdd.n2520 vdd.n268 146.341
R1513 vdd.n2520 vdd.n264 146.341
R1514 vdd.n2526 vdd.n264 146.341
R1515 vdd.n2526 vdd.n257 146.341
R1516 vdd.n2536 vdd.n257 146.341
R1517 vdd.n2536 vdd.n253 146.341
R1518 vdd.n2542 vdd.n253 146.341
R1519 vdd.n2542 vdd.n244 146.341
R1520 vdd.n2552 vdd.n244 146.341
R1521 vdd.n2552 vdd.n240 146.341
R1522 vdd.n2558 vdd.n240 146.341
R1523 vdd.n2558 vdd.n232 146.341
R1524 vdd.n2568 vdd.n232 146.341
R1525 vdd.n2568 vdd.n233 146.341
R1526 vdd.n233 vdd.n65 146.341
R1527 vdd.n66 vdd.n65 146.341
R1528 vdd.n67 vdd.n66 146.341
R1529 vdd.n226 vdd.n67 146.341
R1530 vdd.n226 vdd.n75 146.341
R1531 vdd.n76 vdd.n75 146.341
R1532 vdd.n77 vdd.n76 146.341
R1533 vdd.n223 vdd.n77 146.341
R1534 vdd.n223 vdd.n86 146.341
R1535 vdd.n87 vdd.n86 146.341
R1536 vdd.n88 vdd.n87 146.341
R1537 vdd.n220 vdd.n88 146.341
R1538 vdd.n220 vdd.n97 146.341
R1539 vdd.n98 vdd.n97 146.341
R1540 vdd.n99 vdd.n98 146.341
R1541 vdd.n217 vdd.n99 146.341
R1542 vdd.n217 vdd.n108 146.341
R1543 vdd.n109 vdd.n108 146.341
R1544 vdd.n110 vdd.n109 146.341
R1545 vdd.n2493 vdd.n287 146.341
R1546 vdd.n2493 vdd.n317 146.341
R1547 vdd.n2489 vdd.n2488 146.341
R1548 vdd.n325 vdd.n324 146.341
R1549 vdd.n2481 vdd.n327 146.341
R1550 vdd.n2479 vdd.n2478 146.341
R1551 vdd.n2475 vdd.n2474 146.341
R1552 vdd.n2471 vdd.n2470 146.341
R1553 vdd.n2467 vdd.n2466 146.341
R1554 vdd.n2458 vdd.n2457 146.341
R1555 vdd.n2455 vdd.n2454 146.341
R1556 vdd.n2451 vdd.n2450 146.341
R1557 vdd.n2447 vdd.n2446 146.341
R1558 vdd.n2443 vdd.n2442 146.341
R1559 vdd.n2439 vdd.n2438 146.341
R1560 vdd.n2435 vdd.n2434 146.341
R1561 vdd.n2431 vdd.n2430 146.341
R1562 vdd.n2427 vdd.n2426 146.341
R1563 vdd.n2423 vdd.n2422 146.341
R1564 vdd.n2416 vdd.n2415 146.341
R1565 vdd.n2413 vdd.n2412 146.341
R1566 vdd.n2409 vdd.n2408 146.341
R1567 vdd.n2405 vdd.n2404 146.341
R1568 vdd.n2401 vdd.n2400 146.341
R1569 vdd.n2397 vdd.n2396 146.341
R1570 vdd.n2372 vdd.n2371 146.341
R1571 vdd.n2389 vdd.n2374 146.341
R1572 vdd.n2387 vdd.n2386 146.341
R1573 vdd.n2383 vdd.n316 146.341
R1574 vdd.n2502 vdd.n283 146.341
R1575 vdd.n2502 vdd.n275 146.341
R1576 vdd.n2512 vdd.n275 146.341
R1577 vdd.n2512 vdd.n271 146.341
R1578 vdd.n2518 vdd.n271 146.341
R1579 vdd.n2518 vdd.n263 146.341
R1580 vdd.n2528 vdd.n263 146.341
R1581 vdd.n2528 vdd.n259 146.341
R1582 vdd.n2534 vdd.n259 146.341
R1583 vdd.n2534 vdd.n251 146.341
R1584 vdd.n2544 vdd.n251 146.341
R1585 vdd.n2544 vdd.n247 146.341
R1586 vdd.n2550 vdd.n247 146.341
R1587 vdd.n2550 vdd.n239 146.341
R1588 vdd.n2560 vdd.n239 146.341
R1589 vdd.n2560 vdd.n235 146.341
R1590 vdd.n2566 vdd.n235 146.341
R1591 vdd.n2566 vdd.n62 146.341
R1592 vdd.n2746 vdd.n62 146.341
R1593 vdd.n2746 vdd.n63 146.341
R1594 vdd.n2742 vdd.n63 146.341
R1595 vdd.n2742 vdd.n69 146.341
R1596 vdd.n2738 vdd.n69 146.341
R1597 vdd.n2738 vdd.n74 146.341
R1598 vdd.n2734 vdd.n74 146.341
R1599 vdd.n2734 vdd.n78 146.341
R1600 vdd.n2730 vdd.n78 146.341
R1601 vdd.n2730 vdd.n84 146.341
R1602 vdd.n2726 vdd.n84 146.341
R1603 vdd.n2726 vdd.n90 146.341
R1604 vdd.n2722 vdd.n90 146.341
R1605 vdd.n2722 vdd.n96 146.341
R1606 vdd.n2718 vdd.n96 146.341
R1607 vdd.n2718 vdd.n101 146.341
R1608 vdd.n2714 vdd.n101 146.341
R1609 vdd.n2714 vdd.n107 146.341
R1610 vdd.n2710 vdd.n107 146.341
R1611 vdd.n1405 vdd.n1404 146.341
R1612 vdd.n1402 vdd.n1230 146.341
R1613 vdd.n1239 vdd.n1235 146.341
R1614 vdd.n1394 vdd.n1393 146.341
R1615 vdd.n1391 vdd.n1241 146.341
R1616 vdd.n1387 vdd.n1386 146.341
R1617 vdd.n1384 vdd.n1246 146.341
R1618 vdd.n1380 vdd.n1379 146.341
R1619 vdd.n1377 vdd.n1253 146.341
R1620 vdd.n1371 vdd.n1370 146.341
R1621 vdd.n1368 vdd.n1261 146.341
R1622 vdd.n1364 vdd.n1363 146.341
R1623 vdd.n1361 vdd.n1267 146.341
R1624 vdd.n1357 vdd.n1356 146.341
R1625 vdd.n1354 vdd.n1274 146.341
R1626 vdd.n1350 vdd.n1349 146.341
R1627 vdd.n1347 vdd.n1281 146.341
R1628 vdd.n1343 vdd.n1342 146.341
R1629 vdd.n1340 vdd.n1288 146.341
R1630 vdd.n1334 vdd.n1333 146.341
R1631 vdd.n1331 vdd.n1296 146.341
R1632 vdd.n1327 vdd.n1326 146.341
R1633 vdd.n1324 vdd.n1302 146.341
R1634 vdd.n1320 vdd.n1319 146.341
R1635 vdd.n1317 vdd.n1315 146.341
R1636 vdd.n1313 vdd.n1311 146.341
R1637 vdd.n714 vdd.n713 146.341
R1638 vdd.n721 vdd.n715 146.341
R1639 vdd.n1085 vdd.n866 146.341
R1640 vdd.n1085 vdd.n862 146.341
R1641 vdd.n1091 vdd.n862 146.341
R1642 vdd.n1091 vdd.n853 146.341
R1643 vdd.n1101 vdd.n853 146.341
R1644 vdd.n1101 vdd.n849 146.341
R1645 vdd.n1107 vdd.n849 146.341
R1646 vdd.n1107 vdd.n842 146.341
R1647 vdd.n1117 vdd.n842 146.341
R1648 vdd.n1117 vdd.n838 146.341
R1649 vdd.n1123 vdd.n838 146.341
R1650 vdd.n1123 vdd.n829 146.341
R1651 vdd.n1133 vdd.n829 146.341
R1652 vdd.n1133 vdd.n825 146.341
R1653 vdd.n1139 vdd.n825 146.341
R1654 vdd.n1139 vdd.n818 146.341
R1655 vdd.n1150 vdd.n818 146.341
R1656 vdd.n1150 vdd.n814 146.341
R1657 vdd.n1156 vdd.n814 146.341
R1658 vdd.n1156 vdd.n775 146.341
R1659 vdd.n1166 vdd.n775 146.341
R1660 vdd.n1166 vdd.n771 146.341
R1661 vdd.n1172 vdd.n771 146.341
R1662 vdd.n1172 vdd.n764 146.341
R1663 vdd.n1182 vdd.n764 146.341
R1664 vdd.n1182 vdd.n760 146.341
R1665 vdd.n1188 vdd.n760 146.341
R1666 vdd.n1188 vdd.n751 146.341
R1667 vdd.n1198 vdd.n751 146.341
R1668 vdd.n1198 vdd.n747 146.341
R1669 vdd.n1204 vdd.n747 146.341
R1670 vdd.n1204 vdd.n740 146.341
R1671 vdd.n1214 vdd.n740 146.341
R1672 vdd.n1214 vdd.n735 146.341
R1673 vdd.n1221 vdd.n735 146.341
R1674 vdd.n1221 vdd.n723 146.341
R1675 vdd.n1413 vdd.n723 146.341
R1676 vdd.n1074 vdd.n872 146.341
R1677 vdd.n1074 vdd.n901 146.341
R1678 vdd.n905 vdd.n904 146.341
R1679 vdd.n907 vdd.n906 146.341
R1680 vdd.n911 vdd.n910 146.341
R1681 vdd.n913 vdd.n912 146.341
R1682 vdd.n917 vdd.n916 146.341
R1683 vdd.n919 vdd.n918 146.341
R1684 vdd.n1047 vdd.n922 146.341
R1685 vdd.n924 vdd.n923 146.341
R1686 vdd.n928 vdd.n927 146.341
R1687 vdd.n930 vdd.n929 146.341
R1688 vdd.n934 vdd.n933 146.341
R1689 vdd.n936 vdd.n935 146.341
R1690 vdd.n940 vdd.n939 146.341
R1691 vdd.n942 vdd.n941 146.341
R1692 vdd.n946 vdd.n945 146.341
R1693 vdd.n948 vdd.n947 146.341
R1694 vdd.n1014 vdd.n951 146.341
R1695 vdd.n953 vdd.n952 146.341
R1696 vdd.n957 vdd.n956 146.341
R1697 vdd.n959 vdd.n958 146.341
R1698 vdd.n963 vdd.n962 146.341
R1699 vdd.n965 vdd.n964 146.341
R1700 vdd.n969 vdd.n968 146.341
R1701 vdd.n971 vdd.n970 146.341
R1702 vdd.n975 vdd.n974 146.341
R1703 vdd.n977 vdd.n976 146.341
R1704 vdd.n980 vdd.n900 146.341
R1705 vdd.n1083 vdd.n868 146.341
R1706 vdd.n1083 vdd.n860 146.341
R1707 vdd.n1093 vdd.n860 146.341
R1708 vdd.n1093 vdd.n856 146.341
R1709 vdd.n1099 vdd.n856 146.341
R1710 vdd.n1099 vdd.n848 146.341
R1711 vdd.n1109 vdd.n848 146.341
R1712 vdd.n1109 vdd.n844 146.341
R1713 vdd.n1115 vdd.n844 146.341
R1714 vdd.n1115 vdd.n836 146.341
R1715 vdd.n1125 vdd.n836 146.341
R1716 vdd.n1125 vdd.n832 146.341
R1717 vdd.n1131 vdd.n832 146.341
R1718 vdd.n1131 vdd.n824 146.341
R1719 vdd.n1141 vdd.n824 146.341
R1720 vdd.n1141 vdd.n820 146.341
R1721 vdd.n1148 vdd.n820 146.341
R1722 vdd.n1148 vdd.n812 146.341
R1723 vdd.n1158 vdd.n812 146.341
R1724 vdd.n1158 vdd.n778 146.341
R1725 vdd.n1164 vdd.n778 146.341
R1726 vdd.n1164 vdd.n770 146.341
R1727 vdd.n1174 vdd.n770 146.341
R1728 vdd.n1174 vdd.n766 146.341
R1729 vdd.n1180 vdd.n766 146.341
R1730 vdd.n1180 vdd.n758 146.341
R1731 vdd.n1190 vdd.n758 146.341
R1732 vdd.n1190 vdd.n754 146.341
R1733 vdd.n1196 vdd.n754 146.341
R1734 vdd.n1196 vdd.n746 146.341
R1735 vdd.n1206 vdd.n746 146.341
R1736 vdd.n1206 vdd.n742 146.341
R1737 vdd.n1212 vdd.n742 146.341
R1738 vdd.n1212 vdd.n733 146.341
R1739 vdd.n1223 vdd.n733 146.341
R1740 vdd.n1223 vdd.n728 146.341
R1741 vdd.n1411 vdd.n728 146.341
R1742 vdd.n982 vdd.t45 139.282
R1743 vdd.n1015 vdd.t59 139.282
R1744 vdd.n1048 vdd.t86 139.282
R1745 vdd.n718 vdd.t88 139.282
R1746 vdd.n1290 vdd.t98 139.282
R1747 vdd.n1255 vdd.t69 139.282
R1748 vdd.n212 vdd.t29 139.282
R1749 vdd.n179 vdd.t40 139.282
R1750 vdd.n144 vdd.t72 139.282
R1751 vdd.n354 vdd.t83 139.282
R1752 vdd.n2463 vdd.t52 139.282
R1753 vdd.n2380 vdd.t38 139.282
R1754 vdd.n22 vdd.n20 117.314
R1755 vdd.n17 vdd.n15 117.314
R1756 vdd.n27 vdd.n26 116.927
R1757 vdd.n24 vdd.n23 116.927
R1758 vdd.n22 vdd.n21 116.927
R1759 vdd.n17 vdd.n16 116.927
R1760 vdd.n19 vdd.n18 116.927
R1761 vdd.n27 vdd.n25 116.927
R1762 vdd.n983 vdd.t44 113.489
R1763 vdd.n1016 vdd.t58 113.489
R1764 vdd.n1049 vdd.t85 113.489
R1765 vdd.n719 vdd.t89 113.489
R1766 vdd.n1291 vdd.t99 113.489
R1767 vdd.n1256 vdd.t70 113.489
R1768 vdd.n213 vdd.t30 113.489
R1769 vdd.n180 vdd.t41 113.489
R1770 vdd.n145 vdd.t73 113.489
R1771 vdd.n355 vdd.t82 113.489
R1772 vdd.n2464 vdd.t51 113.489
R1773 vdd.n2381 vdd.t37 113.489
R1774 vdd.n9 vdd.n7 109.74
R1775 vdd.n2 vdd.n0 109.74
R1776 vdd.n9 vdd.n8 109.166
R1777 vdd.n11 vdd.n10 109.166
R1778 vdd.n13 vdd.n12 109.166
R1779 vdd.n6 vdd.n5 109.166
R1780 vdd.n4 vdd.n3 109.166
R1781 vdd.n2 vdd.n1 109.166
R1782 vdd.n2140 vdd.n520 99.5127
R1783 vdd.n2144 vdd.n520 99.5127
R1784 vdd.n2144 vdd.n510 99.5127
R1785 vdd.n2152 vdd.n510 99.5127
R1786 vdd.n2152 vdd.n508 99.5127
R1787 vdd.n2156 vdd.n508 99.5127
R1788 vdd.n2156 vdd.n498 99.5127
R1789 vdd.n2164 vdd.n498 99.5127
R1790 vdd.n2164 vdd.n496 99.5127
R1791 vdd.n2168 vdd.n496 99.5127
R1792 vdd.n2168 vdd.n487 99.5127
R1793 vdd.n2176 vdd.n487 99.5127
R1794 vdd.n2176 vdd.n485 99.5127
R1795 vdd.n2180 vdd.n485 99.5127
R1796 vdd.n2180 vdd.n476 99.5127
R1797 vdd.n2188 vdd.n476 99.5127
R1798 vdd.n2188 vdd.n474 99.5127
R1799 vdd.n2192 vdd.n474 99.5127
R1800 vdd.n2192 vdd.n464 99.5127
R1801 vdd.n2200 vdd.n464 99.5127
R1802 vdd.n2200 vdd.n462 99.5127
R1803 vdd.n2204 vdd.n462 99.5127
R1804 vdd.n2204 vdd.n452 99.5127
R1805 vdd.n2212 vdd.n452 99.5127
R1806 vdd.n2212 vdd.n450 99.5127
R1807 vdd.n2216 vdd.n450 99.5127
R1808 vdd.n2216 vdd.n440 99.5127
R1809 vdd.n2224 vdd.n440 99.5127
R1810 vdd.n2224 vdd.n438 99.5127
R1811 vdd.n2228 vdd.n438 99.5127
R1812 vdd.n2228 vdd.n429 99.5127
R1813 vdd.n2236 vdd.n429 99.5127
R1814 vdd.n2236 vdd.n427 99.5127
R1815 vdd.n2240 vdd.n427 99.5127
R1816 vdd.n2240 vdd.n415 99.5127
R1817 vdd.n2285 vdd.n415 99.5127
R1818 vdd.n2285 vdd.n413 99.5127
R1819 vdd.n2289 vdd.n413 99.5127
R1820 vdd.n2289 vdd.n386 99.5127
R1821 vdd.n2344 vdd.n386 99.5127
R1822 vdd.n2340 vdd.n2339 99.5127
R1823 vdd.n2337 vdd.n391 99.5127
R1824 vdd.n2333 vdd.n2332 99.5127
R1825 vdd.n2330 vdd.n394 99.5127
R1826 vdd.n2326 vdd.n2325 99.5127
R1827 vdd.n2323 vdd.n2320 99.5127
R1828 vdd.n2318 vdd.n397 99.5127
R1829 vdd.n2314 vdd.n2313 99.5127
R1830 vdd.n2311 vdd.n400 99.5127
R1831 vdd.n2307 vdd.n2306 99.5127
R1832 vdd.n2304 vdd.n403 99.5127
R1833 vdd.n2299 vdd.n2298 99.5127
R1834 vdd.n1970 vdd.n1884 99.5127
R1835 vdd.n1970 vdd.n517 99.5127
R1836 vdd.n1973 vdd.n517 99.5127
R1837 vdd.n1973 vdd.n511 99.5127
R1838 vdd.n1976 vdd.n511 99.5127
R1839 vdd.n1976 vdd.n506 99.5127
R1840 vdd.n1979 vdd.n506 99.5127
R1841 vdd.n1979 vdd.n500 99.5127
R1842 vdd.n1982 vdd.n500 99.5127
R1843 vdd.n1982 vdd.n494 99.5127
R1844 vdd.n1985 vdd.n494 99.5127
R1845 vdd.n1985 vdd.n489 99.5127
R1846 vdd.n1988 vdd.n489 99.5127
R1847 vdd.n1988 vdd.n483 99.5127
R1848 vdd.n2059 vdd.n483 99.5127
R1849 vdd.n2059 vdd.n477 99.5127
R1850 vdd.n2055 vdd.n477 99.5127
R1851 vdd.n2055 vdd.n472 99.5127
R1852 vdd.n2052 vdd.n472 99.5127
R1853 vdd.n2052 vdd.n465 99.5127
R1854 vdd.n2014 vdd.n465 99.5127
R1855 vdd.n2014 vdd.n459 99.5127
R1856 vdd.n2011 vdd.n459 99.5127
R1857 vdd.n2011 vdd.n453 99.5127
R1858 vdd.n2008 vdd.n453 99.5127
R1859 vdd.n2008 vdd.n447 99.5127
R1860 vdd.n2005 vdd.n447 99.5127
R1861 vdd.n2005 vdd.n441 99.5127
R1862 vdd.n2002 vdd.n441 99.5127
R1863 vdd.n2002 vdd.n436 99.5127
R1864 vdd.n1999 vdd.n436 99.5127
R1865 vdd.n1999 vdd.n431 99.5127
R1866 vdd.n1996 vdd.n431 99.5127
R1867 vdd.n1996 vdd.n425 99.5127
R1868 vdd.n1993 vdd.n425 99.5127
R1869 vdd.n1993 vdd.n417 99.5127
R1870 vdd.n417 vdd.n409 99.5127
R1871 vdd.n2291 vdd.n409 99.5127
R1872 vdd.n2292 vdd.n2291 99.5127
R1873 vdd.n2292 vdd.n384 99.5127
R1874 vdd.n1919 vdd.n1917 99.5127
R1875 vdd.n1923 vdd.n1917 99.5127
R1876 vdd.n1927 vdd.n1925 99.5127
R1877 vdd.n1931 vdd.n1915 99.5127
R1878 vdd.n1935 vdd.n1933 99.5127
R1879 vdd.n1939 vdd.n1913 99.5127
R1880 vdd.n1943 vdd.n1941 99.5127
R1881 vdd.n1947 vdd.n1911 99.5127
R1882 vdd.n1951 vdd.n1949 99.5127
R1883 vdd.n1955 vdd.n1909 99.5127
R1884 vdd.n1959 vdd.n1957 99.5127
R1885 vdd.n1964 vdd.n1905 99.5127
R1886 vdd.n1967 vdd.n1966 99.5127
R1887 vdd.n1821 vdd.n1820 99.5127
R1888 vdd.n1817 vdd.n1816 99.5127
R1889 vdd.n1813 vdd.n1812 99.5127
R1890 vdd.n1809 vdd.n1808 99.5127
R1891 vdd.n1805 vdd.n1804 99.5127
R1892 vdd.n1801 vdd.n1800 99.5127
R1893 vdd.n1797 vdd.n1796 99.5127
R1894 vdd.n1793 vdd.n1792 99.5127
R1895 vdd.n1789 vdd.n1788 99.5127
R1896 vdd.n1785 vdd.n1784 99.5127
R1897 vdd.n1781 vdd.n1780 99.5127
R1898 vdd.n1776 vdd.n1775 99.5127
R1899 vdd.n1593 vdd.n680 99.5127
R1900 vdd.n1593 vdd.n673 99.5127
R1901 vdd.n1590 vdd.n673 99.5127
R1902 vdd.n1590 vdd.n666 99.5127
R1903 vdd.n1587 vdd.n666 99.5127
R1904 vdd.n1587 vdd.n660 99.5127
R1905 vdd.n1584 vdd.n660 99.5127
R1906 vdd.n1584 vdd.n655 99.5127
R1907 vdd.n1581 vdd.n655 99.5127
R1908 vdd.n1581 vdd.n649 99.5127
R1909 vdd.n1578 vdd.n649 99.5127
R1910 vdd.n1578 vdd.n643 99.5127
R1911 vdd.n1575 vdd.n643 99.5127
R1912 vdd.n1575 vdd.n637 99.5127
R1913 vdd.n1572 vdd.n637 99.5127
R1914 vdd.n1572 vdd.n631 99.5127
R1915 vdd.n1569 vdd.n631 99.5127
R1916 vdd.n1569 vdd.n625 99.5127
R1917 vdd.n1566 vdd.n625 99.5127
R1918 vdd.n1566 vdd.n619 99.5127
R1919 vdd.n1563 vdd.n619 99.5127
R1920 vdd.n1563 vdd.n613 99.5127
R1921 vdd.n1532 vdd.n613 99.5127
R1922 vdd.n1532 vdd.n608 99.5127
R1923 vdd.n1552 vdd.n608 99.5127
R1924 vdd.n1552 vdd.n602 99.5127
R1925 vdd.n1548 vdd.n602 99.5127
R1926 vdd.n1548 vdd.n596 99.5127
R1927 vdd.n1545 vdd.n596 99.5127
R1928 vdd.n1545 vdd.n590 99.5127
R1929 vdd.n1542 vdd.n590 99.5127
R1930 vdd.n1542 vdd.n585 99.5127
R1931 vdd.n1539 vdd.n585 99.5127
R1932 vdd.n1539 vdd.n579 99.5127
R1933 vdd.n1536 vdd.n579 99.5127
R1934 vdd.n1536 vdd.n572 99.5127
R1935 vdd.n572 vdd.n566 99.5127
R1936 vdd.n1767 vdd.n566 99.5127
R1937 vdd.n1767 vdd.n558 99.5127
R1938 vdd.n1771 vdd.n558 99.5127
R1939 vdd.n1644 vdd.n1642 99.5127
R1940 vdd.n1642 vdd.n1641 99.5127
R1941 vdd.n1638 vdd.n1637 99.5127
R1942 vdd.n1635 vdd.n686 99.5127
R1943 vdd.n1631 vdd.n1629 99.5127
R1944 vdd.n1627 vdd.n688 99.5127
R1945 vdd.n1623 vdd.n1621 99.5127
R1946 vdd.n1618 vdd.n1617 99.5127
R1947 vdd.n1615 vdd.n692 99.5127
R1948 vdd.n1611 vdd.n1609 99.5127
R1949 vdd.n1607 vdd.n694 99.5127
R1950 vdd.n1603 vdd.n1601 99.5127
R1951 vdd.n1598 vdd.n1597 99.5127
R1952 vdd.n1648 vdd.n671 99.5127
R1953 vdd.n1656 vdd.n671 99.5127
R1954 vdd.n1656 vdd.n669 99.5127
R1955 vdd.n1660 vdd.n669 99.5127
R1956 vdd.n1660 vdd.n659 99.5127
R1957 vdd.n1669 vdd.n659 99.5127
R1958 vdd.n1669 vdd.n657 99.5127
R1959 vdd.n1673 vdd.n657 99.5127
R1960 vdd.n1673 vdd.n647 99.5127
R1961 vdd.n1681 vdd.n647 99.5127
R1962 vdd.n1681 vdd.n645 99.5127
R1963 vdd.n1685 vdd.n645 99.5127
R1964 vdd.n1685 vdd.n635 99.5127
R1965 vdd.n1693 vdd.n635 99.5127
R1966 vdd.n1693 vdd.n633 99.5127
R1967 vdd.n1697 vdd.n633 99.5127
R1968 vdd.n1697 vdd.n623 99.5127
R1969 vdd.n1705 vdd.n623 99.5127
R1970 vdd.n1705 vdd.n621 99.5127
R1971 vdd.n1709 vdd.n621 99.5127
R1972 vdd.n1709 vdd.n612 99.5127
R1973 vdd.n1717 vdd.n612 99.5127
R1974 vdd.n1717 vdd.n610 99.5127
R1975 vdd.n1721 vdd.n610 99.5127
R1976 vdd.n1721 vdd.n601 99.5127
R1977 vdd.n1729 vdd.n601 99.5127
R1978 vdd.n1729 vdd.n599 99.5127
R1979 vdd.n1733 vdd.n599 99.5127
R1980 vdd.n1733 vdd.n589 99.5127
R1981 vdd.n1741 vdd.n589 99.5127
R1982 vdd.n1741 vdd.n587 99.5127
R1983 vdd.n1745 vdd.n587 99.5127
R1984 vdd.n1745 vdd.n577 99.5127
R1985 vdd.n1753 vdd.n577 99.5127
R1986 vdd.n1753 vdd.n574 99.5127
R1987 vdd.n1758 vdd.n574 99.5127
R1988 vdd.n1758 vdd.n575 99.5127
R1989 vdd.n575 vdd.n560 99.5127
R1990 vdd.n1827 vdd.n560 99.5127
R1991 vdd.n1827 vdd.n561 99.5127
R1992 vdd.n2273 vdd.n2272 99.5127
R1993 vdd.n2270 vdd.n2248 99.5127
R1994 vdd.n2266 vdd.n2265 99.5127
R1995 vdd.n2263 vdd.n2251 99.5127
R1996 vdd.n2259 vdd.n2258 99.5127
R1997 vdd.n2256 vdd.n2254 99.5127
R1998 vdd.n2368 vdd.n2367 99.5127
R1999 vdd.n2365 vdd.n370 99.5127
R2000 vdd.n2361 vdd.n2360 99.5127
R2001 vdd.n2358 vdd.n373 99.5127
R2002 vdd.n2354 vdd.n2353 99.5127
R2003 vdd.n2351 vdd.n376 99.5127
R2004 vdd.n2082 vdd.n1885 99.5127
R2005 vdd.n2082 vdd.n518 99.5127
R2006 vdd.n2079 vdd.n518 99.5127
R2007 vdd.n2079 vdd.n512 99.5127
R2008 vdd.n2076 vdd.n512 99.5127
R2009 vdd.n2076 vdd.n507 99.5127
R2010 vdd.n2073 vdd.n507 99.5127
R2011 vdd.n2073 vdd.n501 99.5127
R2012 vdd.n2070 vdd.n501 99.5127
R2013 vdd.n2070 vdd.n495 99.5127
R2014 vdd.n2067 vdd.n495 99.5127
R2015 vdd.n2067 vdd.n490 99.5127
R2016 vdd.n2064 vdd.n490 99.5127
R2017 vdd.n2064 vdd.n484 99.5127
R2018 vdd.n2061 vdd.n484 99.5127
R2019 vdd.n2061 vdd.n478 99.5127
R2020 vdd.n2017 vdd.n478 99.5127
R2021 vdd.n2017 vdd.n473 99.5127
R2022 vdd.n2050 vdd.n473 99.5127
R2023 vdd.n2050 vdd.n466 99.5127
R2024 vdd.n2046 vdd.n466 99.5127
R2025 vdd.n2046 vdd.n460 99.5127
R2026 vdd.n2043 vdd.n460 99.5127
R2027 vdd.n2043 vdd.n454 99.5127
R2028 vdd.n2040 vdd.n454 99.5127
R2029 vdd.n2040 vdd.n448 99.5127
R2030 vdd.n2037 vdd.n448 99.5127
R2031 vdd.n2037 vdd.n442 99.5127
R2032 vdd.n2034 vdd.n442 99.5127
R2033 vdd.n2034 vdd.n437 99.5127
R2034 vdd.n2031 vdd.n437 99.5127
R2035 vdd.n2031 vdd.n432 99.5127
R2036 vdd.n2028 vdd.n432 99.5127
R2037 vdd.n2028 vdd.n426 99.5127
R2038 vdd.n2025 vdd.n426 99.5127
R2039 vdd.n2025 vdd.n418 99.5127
R2040 vdd.n2022 vdd.n418 99.5127
R2041 vdd.n2022 vdd.n411 99.5127
R2042 vdd.n411 vdd.n382 99.5127
R2043 vdd.n2346 vdd.n382 99.5127
R2044 vdd.n2134 vdd.n2132 99.5127
R2045 vdd.n2130 vdd.n1889 99.5127
R2046 vdd.n2126 vdd.n2124 99.5127
R2047 vdd.n2122 vdd.n1891 99.5127
R2048 vdd.n2118 vdd.n2116 99.5127
R2049 vdd.n2114 vdd.n1893 99.5127
R2050 vdd.n2110 vdd.n2108 99.5127
R2051 vdd.n2106 vdd.n1895 99.5127
R2052 vdd.n2102 vdd.n2100 99.5127
R2053 vdd.n2098 vdd.n1897 99.5127
R2054 vdd.n2094 vdd.n2092 99.5127
R2055 vdd.n2090 vdd.n1899 99.5127
R2056 vdd.n2138 vdd.n516 99.5127
R2057 vdd.n2146 vdd.n516 99.5127
R2058 vdd.n2146 vdd.n514 99.5127
R2059 vdd.n2150 vdd.n514 99.5127
R2060 vdd.n2150 vdd.n505 99.5127
R2061 vdd.n2158 vdd.n505 99.5127
R2062 vdd.n2158 vdd.n503 99.5127
R2063 vdd.n2162 vdd.n503 99.5127
R2064 vdd.n2162 vdd.n493 99.5127
R2065 vdd.n2170 vdd.n493 99.5127
R2066 vdd.n2170 vdd.n491 99.5127
R2067 vdd.n2174 vdd.n491 99.5127
R2068 vdd.n2174 vdd.n481 99.5127
R2069 vdd.n2182 vdd.n481 99.5127
R2070 vdd.n2182 vdd.n479 99.5127
R2071 vdd.n2186 vdd.n479 99.5127
R2072 vdd.n2186 vdd.n470 99.5127
R2073 vdd.n2194 vdd.n470 99.5127
R2074 vdd.n2194 vdd.n468 99.5127
R2075 vdd.n2198 vdd.n468 99.5127
R2076 vdd.n2198 vdd.n458 99.5127
R2077 vdd.n2206 vdd.n458 99.5127
R2078 vdd.n2206 vdd.n456 99.5127
R2079 vdd.n2210 vdd.n456 99.5127
R2080 vdd.n2210 vdd.n446 99.5127
R2081 vdd.n2218 vdd.n446 99.5127
R2082 vdd.n2218 vdd.n444 99.5127
R2083 vdd.n2222 vdd.n444 99.5127
R2084 vdd.n2222 vdd.n435 99.5127
R2085 vdd.n2230 vdd.n435 99.5127
R2086 vdd.n2230 vdd.n433 99.5127
R2087 vdd.n2234 vdd.n433 99.5127
R2088 vdd.n2234 vdd.n423 99.5127
R2089 vdd.n2242 vdd.n423 99.5127
R2090 vdd.n2242 vdd.n419 99.5127
R2091 vdd.n2283 vdd.n419 99.5127
R2092 vdd.n2283 vdd.n420 99.5127
R2093 vdd.n420 vdd.n412 99.5127
R2094 vdd.n2278 vdd.n412 99.5127
R2095 vdd.n2278 vdd.n385 99.5127
R2096 vdd.n1881 vdd.n551 99.5127
R2097 vdd.n1877 vdd.n1876 99.5127
R2098 vdd.n1873 vdd.n1872 99.5127
R2099 vdd.n1869 vdd.n1868 99.5127
R2100 vdd.n1865 vdd.n1864 99.5127
R2101 vdd.n1861 vdd.n1860 99.5127
R2102 vdd.n1857 vdd.n1856 99.5127
R2103 vdd.n1853 vdd.n1852 99.5127
R2104 vdd.n1849 vdd.n1848 99.5127
R2105 vdd.n1845 vdd.n1844 99.5127
R2106 vdd.n1841 vdd.n1840 99.5127
R2107 vdd.n1837 vdd.n1836 99.5127
R2108 vdd.n1833 vdd.n549 99.5127
R2109 vdd.n1483 vdd.n681 99.5127
R2110 vdd.n1483 vdd.n674 99.5127
R2111 vdd.n1486 vdd.n674 99.5127
R2112 vdd.n1486 vdd.n667 99.5127
R2113 vdd.n1489 vdd.n667 99.5127
R2114 vdd.n1489 vdd.n661 99.5127
R2115 vdd.n1492 vdd.n661 99.5127
R2116 vdd.n1492 vdd.n656 99.5127
R2117 vdd.n1495 vdd.n656 99.5127
R2118 vdd.n1495 vdd.n650 99.5127
R2119 vdd.n1498 vdd.n650 99.5127
R2120 vdd.n1498 vdd.n644 99.5127
R2121 vdd.n1501 vdd.n644 99.5127
R2122 vdd.n1501 vdd.n638 99.5127
R2123 vdd.n1504 vdd.n638 99.5127
R2124 vdd.n1504 vdd.n632 99.5127
R2125 vdd.n1507 vdd.n632 99.5127
R2126 vdd.n1507 vdd.n626 99.5127
R2127 vdd.n1510 vdd.n626 99.5127
R2128 vdd.n1510 vdd.n620 99.5127
R2129 vdd.n1561 vdd.n620 99.5127
R2130 vdd.n1561 vdd.n614 99.5127
R2131 vdd.n1557 vdd.n614 99.5127
R2132 vdd.n1557 vdd.n609 99.5127
R2133 vdd.n1554 vdd.n609 99.5127
R2134 vdd.n1554 vdd.n603 99.5127
R2135 vdd.n1529 vdd.n603 99.5127
R2136 vdd.n1529 vdd.n597 99.5127
R2137 vdd.n1526 vdd.n597 99.5127
R2138 vdd.n1526 vdd.n591 99.5127
R2139 vdd.n1523 vdd.n591 99.5127
R2140 vdd.n1523 vdd.n586 99.5127
R2141 vdd.n1520 vdd.n586 99.5127
R2142 vdd.n1520 vdd.n580 99.5127
R2143 vdd.n1517 vdd.n580 99.5127
R2144 vdd.n1517 vdd.n573 99.5127
R2145 vdd.n1514 vdd.n573 99.5127
R2146 vdd.n1514 vdd.n557 99.5127
R2147 vdd.n1829 vdd.n557 99.5127
R2148 vdd.n1830 vdd.n1829 99.5127
R2149 vdd.n1432 vdd.n678 99.5127
R2150 vdd.n1436 vdd.n1430 99.5127
R2151 vdd.n1440 vdd.n1438 99.5127
R2152 vdd.n1444 vdd.n1428 99.5127
R2153 vdd.n1448 vdd.n1446 99.5127
R2154 vdd.n1452 vdd.n1426 99.5127
R2155 vdd.n1456 vdd.n1454 99.5127
R2156 vdd.n1460 vdd.n707 99.5127
R2157 vdd.n1464 vdd.n1462 99.5127
R2158 vdd.n1468 vdd.n705 99.5127
R2159 vdd.n1472 vdd.n1470 99.5127
R2160 vdd.n1477 vdd.n701 99.5127
R2161 vdd.n1480 vdd.n1479 99.5127
R2162 vdd.n1650 vdd.n676 99.5127
R2163 vdd.n1654 vdd.n676 99.5127
R2164 vdd.n1654 vdd.n665 99.5127
R2165 vdd.n1662 vdd.n665 99.5127
R2166 vdd.n1662 vdd.n662 99.5127
R2167 vdd.n1667 vdd.n662 99.5127
R2168 vdd.n1667 vdd.n653 99.5127
R2169 vdd.n1675 vdd.n653 99.5127
R2170 vdd.n1675 vdd.n651 99.5127
R2171 vdd.n1679 vdd.n651 99.5127
R2172 vdd.n1679 vdd.n641 99.5127
R2173 vdd.n1687 vdd.n641 99.5127
R2174 vdd.n1687 vdd.n639 99.5127
R2175 vdd.n1691 vdd.n639 99.5127
R2176 vdd.n1691 vdd.n629 99.5127
R2177 vdd.n1699 vdd.n629 99.5127
R2178 vdd.n1699 vdd.n627 99.5127
R2179 vdd.n1703 vdd.n627 99.5127
R2180 vdd.n1703 vdd.n617 99.5127
R2181 vdd.n1711 vdd.n617 99.5127
R2182 vdd.n1711 vdd.n615 99.5127
R2183 vdd.n1715 vdd.n615 99.5127
R2184 vdd.n1715 vdd.n606 99.5127
R2185 vdd.n1723 vdd.n606 99.5127
R2186 vdd.n1723 vdd.n604 99.5127
R2187 vdd.n1727 vdd.n604 99.5127
R2188 vdd.n1727 vdd.n594 99.5127
R2189 vdd.n1735 vdd.n594 99.5127
R2190 vdd.n1735 vdd.n592 99.5127
R2191 vdd.n1739 vdd.n592 99.5127
R2192 vdd.n1739 vdd.n583 99.5127
R2193 vdd.n1747 vdd.n583 99.5127
R2194 vdd.n1747 vdd.n581 99.5127
R2195 vdd.n1751 vdd.n581 99.5127
R2196 vdd.n1751 vdd.n570 99.5127
R2197 vdd.n1760 vdd.n570 99.5127
R2198 vdd.n1760 vdd.n568 99.5127
R2199 vdd.n1765 vdd.n568 99.5127
R2200 vdd.n1765 vdd.n559 99.5127
R2201 vdd.n559 vdd.n550 99.5127
R2202 vdd.t174 vdd.t165 94.423
R2203 vdd.n49 vdd.t104 79.3769
R2204 vdd.n39 vdd.t162 79.3769
R2205 vdd.n30 vdd.t203 79.3769
R2206 vdd.n800 vdd.t163 79.3769
R2207 vdd.n790 vdd.t199 79.3769
R2208 vdd.n781 vdd.t119 79.3769
R2209 vdd.n56 vdd.t148 78.8036
R2210 vdd.n46 vdd.t190 78.8036
R2211 vdd.n37 vdd.t164 78.8036
R2212 vdd.n807 vdd.t15 78.8036
R2213 vdd.n797 vdd.t153 78.8036
R2214 vdd.n788 vdd.t112 78.8036
R2215 vdd.n2244 vdd.n421 78.546
R2216 vdd.n1665 vdd.n663 78.546
R2217 vdd.n55 vdd.n54 74.1601
R2218 vdd.n53 vdd.n52 74.1601
R2219 vdd.n51 vdd.n50 74.1601
R2220 vdd.n49 vdd.n48 74.1601
R2221 vdd.n45 vdd.n44 74.1601
R2222 vdd.n43 vdd.n42 74.1601
R2223 vdd.n41 vdd.n40 74.1601
R2224 vdd.n39 vdd.n38 74.1601
R2225 vdd.n36 vdd.n35 74.1601
R2226 vdd.n34 vdd.n33 74.1601
R2227 vdd.n32 vdd.n31 74.1601
R2228 vdd.n30 vdd.n29 74.1601
R2229 vdd.n800 vdd.n799 74.1601
R2230 vdd.n802 vdd.n801 74.1601
R2231 vdd.n804 vdd.n803 74.1601
R2232 vdd.n806 vdd.n805 74.1601
R2233 vdd.n790 vdd.n789 74.1601
R2234 vdd.n792 vdd.n791 74.1601
R2235 vdd.n794 vdd.n793 74.1601
R2236 vdd.n796 vdd.n795 74.1601
R2237 vdd.n781 vdd.n780 74.1601
R2238 vdd.n783 vdd.n782 74.1601
R2239 vdd.n785 vdd.n784 74.1601
R2240 vdd.n787 vdd.n786 74.1601
R2241 vdd.n2133 vdd.n1883 72.8958
R2242 vdd.n2131 vdd.n1883 72.8958
R2243 vdd.n2125 vdd.n1883 72.8958
R2244 vdd.n2123 vdd.n1883 72.8958
R2245 vdd.n2117 vdd.n1883 72.8958
R2246 vdd.n2115 vdd.n1883 72.8958
R2247 vdd.n2109 vdd.n1883 72.8958
R2248 vdd.n2107 vdd.n1883 72.8958
R2249 vdd.n2101 vdd.n1883 72.8958
R2250 vdd.n2099 vdd.n1883 72.8958
R2251 vdd.n2093 vdd.n1883 72.8958
R2252 vdd.n2091 vdd.n1883 72.8958
R2253 vdd.n2085 vdd.n1883 72.8958
R2254 vdd.n381 vdd.n288 72.8958
R2255 vdd.n2352 vdd.n288 72.8958
R2256 vdd.n375 vdd.n288 72.8958
R2257 vdd.n2359 vdd.n288 72.8958
R2258 vdd.n372 vdd.n288 72.8958
R2259 vdd.n2366 vdd.n288 72.8958
R2260 vdd.n369 vdd.n288 72.8958
R2261 vdd.n2257 vdd.n288 72.8958
R2262 vdd.n2253 vdd.n288 72.8958
R2263 vdd.n2264 vdd.n288 72.8958
R2264 vdd.n2250 vdd.n288 72.8958
R2265 vdd.n2271 vdd.n288 72.8958
R2266 vdd.n2274 vdd.n288 72.8958
R2267 vdd.n1643 vdd.n679 72.8958
R2268 vdd.n684 vdd.n679 72.8958
R2269 vdd.n1636 vdd.n679 72.8958
R2270 vdd.n1630 vdd.n679 72.8958
R2271 vdd.n1628 vdd.n679 72.8958
R2272 vdd.n1622 vdd.n679 72.8958
R2273 vdd.n690 vdd.n679 72.8958
R2274 vdd.n1616 vdd.n679 72.8958
R2275 vdd.n1610 vdd.n679 72.8958
R2276 vdd.n1608 vdd.n679 72.8958
R2277 vdd.n1602 vdd.n679 72.8958
R2278 vdd.n698 vdd.n679 72.8958
R2279 vdd.n1882 vdd.n536 72.8958
R2280 vdd.n1882 vdd.n535 72.8958
R2281 vdd.n1882 vdd.n534 72.8958
R2282 vdd.n1882 vdd.n533 72.8958
R2283 vdd.n1882 vdd.n532 72.8958
R2284 vdd.n1882 vdd.n531 72.8958
R2285 vdd.n1882 vdd.n530 72.8958
R2286 vdd.n1882 vdd.n529 72.8958
R2287 vdd.n1882 vdd.n528 72.8958
R2288 vdd.n1882 vdd.n527 72.8958
R2289 vdd.n1882 vdd.n526 72.8958
R2290 vdd.n1882 vdd.n525 72.8958
R2291 vdd.n1882 vdd.n524 72.8958
R2292 vdd.n1918 vdd.n1883 72.8958
R2293 vdd.n1924 vdd.n1883 72.8958
R2294 vdd.n1926 vdd.n1883 72.8958
R2295 vdd.n1932 vdd.n1883 72.8958
R2296 vdd.n1934 vdd.n1883 72.8958
R2297 vdd.n1940 vdd.n1883 72.8958
R2298 vdd.n1942 vdd.n1883 72.8958
R2299 vdd.n1948 vdd.n1883 72.8958
R2300 vdd.n1950 vdd.n1883 72.8958
R2301 vdd.n1956 vdd.n1883 72.8958
R2302 vdd.n1958 vdd.n1883 72.8958
R2303 vdd.n1965 vdd.n1883 72.8958
R2304 vdd.n2297 vdd.n288 72.8958
R2305 vdd.n407 vdd.n288 72.8958
R2306 vdd.n2305 vdd.n288 72.8958
R2307 vdd.n402 vdd.n288 72.8958
R2308 vdd.n2312 vdd.n288 72.8958
R2309 vdd.n399 vdd.n288 72.8958
R2310 vdd.n2319 vdd.n288 72.8958
R2311 vdd.n2324 vdd.n288 72.8958
R2312 vdd.n396 vdd.n288 72.8958
R2313 vdd.n2331 vdd.n288 72.8958
R2314 vdd.n393 vdd.n288 72.8958
R2315 vdd.n2338 vdd.n288 72.8958
R2316 vdd.n390 vdd.n288 72.8958
R2317 vdd.n1882 vdd.n548 72.8958
R2318 vdd.n1882 vdd.n547 72.8958
R2319 vdd.n1882 vdd.n546 72.8958
R2320 vdd.n1882 vdd.n545 72.8958
R2321 vdd.n1882 vdd.n544 72.8958
R2322 vdd.n1882 vdd.n543 72.8958
R2323 vdd.n1882 vdd.n542 72.8958
R2324 vdd.n1882 vdd.n541 72.8958
R2325 vdd.n1882 vdd.n540 72.8958
R2326 vdd.n1882 vdd.n539 72.8958
R2327 vdd.n1882 vdd.n538 72.8958
R2328 vdd.n1882 vdd.n537 72.8958
R2329 vdd.n1431 vdd.n679 72.8958
R2330 vdd.n1437 vdd.n679 72.8958
R2331 vdd.n1439 vdd.n679 72.8958
R2332 vdd.n1445 vdd.n679 72.8958
R2333 vdd.n1447 vdd.n679 72.8958
R2334 vdd.n1453 vdd.n679 72.8958
R2335 vdd.n1455 vdd.n679 72.8958
R2336 vdd.n1461 vdd.n679 72.8958
R2337 vdd.n1463 vdd.n679 72.8958
R2338 vdd.n1469 vdd.n679 72.8958
R2339 vdd.n1471 vdd.n679 72.8958
R2340 vdd.n1478 vdd.n679 72.8958
R2341 vdd.n1076 vdd.n1075 66.2847
R2342 vdd.n1075 vdd.n873 66.2847
R2343 vdd.n1075 vdd.n874 66.2847
R2344 vdd.n1075 vdd.n875 66.2847
R2345 vdd.n1075 vdd.n876 66.2847
R2346 vdd.n1075 vdd.n877 66.2847
R2347 vdd.n1075 vdd.n878 66.2847
R2348 vdd.n1075 vdd.n879 66.2847
R2349 vdd.n1075 vdd.n880 66.2847
R2350 vdd.n1075 vdd.n881 66.2847
R2351 vdd.n1075 vdd.n882 66.2847
R2352 vdd.n1075 vdd.n883 66.2847
R2353 vdd.n1075 vdd.n884 66.2847
R2354 vdd.n1075 vdd.n885 66.2847
R2355 vdd.n1075 vdd.n886 66.2847
R2356 vdd.n1075 vdd.n887 66.2847
R2357 vdd.n1075 vdd.n888 66.2847
R2358 vdd.n1075 vdd.n889 66.2847
R2359 vdd.n1075 vdd.n890 66.2847
R2360 vdd.n1075 vdd.n891 66.2847
R2361 vdd.n1075 vdd.n892 66.2847
R2362 vdd.n1075 vdd.n893 66.2847
R2363 vdd.n1075 vdd.n894 66.2847
R2364 vdd.n1075 vdd.n895 66.2847
R2365 vdd.n1075 vdd.n896 66.2847
R2366 vdd.n1075 vdd.n897 66.2847
R2367 vdd.n1075 vdd.n898 66.2847
R2368 vdd.n1075 vdd.n899 66.2847
R2369 vdd.n727 vdd.n722 66.2847
R2370 vdd.n727 vdd.n726 66.2847
R2371 vdd.n1310 vdd.n727 66.2847
R2372 vdd.n1314 vdd.n727 66.2847
R2373 vdd.n1318 vdd.n727 66.2847
R2374 vdd.n1308 vdd.n727 66.2847
R2375 vdd.n1325 vdd.n727 66.2847
R2376 vdd.n1301 vdd.n727 66.2847
R2377 vdd.n1332 vdd.n727 66.2847
R2378 vdd.n1295 vdd.n727 66.2847
R2379 vdd.n1341 vdd.n727 66.2847
R2380 vdd.n1287 vdd.n727 66.2847
R2381 vdd.n1348 vdd.n727 66.2847
R2382 vdd.n1280 vdd.n727 66.2847
R2383 vdd.n1355 vdd.n727 66.2847
R2384 vdd.n1273 vdd.n727 66.2847
R2385 vdd.n1362 vdd.n727 66.2847
R2386 vdd.n1266 vdd.n727 66.2847
R2387 vdd.n1369 vdd.n727 66.2847
R2388 vdd.n1260 vdd.n727 66.2847
R2389 vdd.n1378 vdd.n727 66.2847
R2390 vdd.n1252 vdd.n727 66.2847
R2391 vdd.n1385 vdd.n727 66.2847
R2392 vdd.n1245 vdd.n727 66.2847
R2393 vdd.n1392 vdd.n727 66.2847
R2394 vdd.n1240 vdd.n727 66.2847
R2395 vdd.n1234 vdd.n727 66.2847
R2396 vdd.n1403 vdd.n727 66.2847
R2397 vdd.n1229 vdd.n727 66.2847
R2398 vdd.n2495 vdd.n2494 66.2847
R2399 vdd.n2494 vdd.n289 66.2847
R2400 vdd.n2494 vdd.n290 66.2847
R2401 vdd.n2494 vdd.n291 66.2847
R2402 vdd.n2494 vdd.n292 66.2847
R2403 vdd.n2494 vdd.n293 66.2847
R2404 vdd.n2494 vdd.n294 66.2847
R2405 vdd.n2494 vdd.n295 66.2847
R2406 vdd.n2494 vdd.n296 66.2847
R2407 vdd.n2494 vdd.n297 66.2847
R2408 vdd.n2494 vdd.n298 66.2847
R2409 vdd.n2494 vdd.n299 66.2847
R2410 vdd.n2494 vdd.n300 66.2847
R2411 vdd.n2494 vdd.n301 66.2847
R2412 vdd.n2494 vdd.n302 66.2847
R2413 vdd.n2494 vdd.n303 66.2847
R2414 vdd.n2494 vdd.n304 66.2847
R2415 vdd.n2494 vdd.n305 66.2847
R2416 vdd.n2494 vdd.n306 66.2847
R2417 vdd.n2494 vdd.n307 66.2847
R2418 vdd.n2494 vdd.n308 66.2847
R2419 vdd.n2494 vdd.n309 66.2847
R2420 vdd.n2494 vdd.n310 66.2847
R2421 vdd.n2494 vdd.n311 66.2847
R2422 vdd.n2494 vdd.n312 66.2847
R2423 vdd.n2494 vdd.n313 66.2847
R2424 vdd.n2494 vdd.n314 66.2847
R2425 vdd.n2494 vdd.n315 66.2847
R2426 vdd.n2604 vdd.n111 66.2847
R2427 vdd.n211 vdd.n111 66.2847
R2428 vdd.n2611 vdd.n111 66.2847
R2429 vdd.n204 vdd.n111 66.2847
R2430 vdd.n2618 vdd.n111 66.2847
R2431 vdd.n197 vdd.n111 66.2847
R2432 vdd.n2625 vdd.n111 66.2847
R2433 vdd.n190 vdd.n111 66.2847
R2434 vdd.n2632 vdd.n111 66.2847
R2435 vdd.n184 vdd.n111 66.2847
R2436 vdd.n2641 vdd.n111 66.2847
R2437 vdd.n176 vdd.n111 66.2847
R2438 vdd.n2648 vdd.n111 66.2847
R2439 vdd.n169 vdd.n111 66.2847
R2440 vdd.n2655 vdd.n111 66.2847
R2441 vdd.n162 vdd.n111 66.2847
R2442 vdd.n2662 vdd.n111 66.2847
R2443 vdd.n155 vdd.n111 66.2847
R2444 vdd.n2669 vdd.n111 66.2847
R2445 vdd.n149 vdd.n111 66.2847
R2446 vdd.n2678 vdd.n111 66.2847
R2447 vdd.n141 vdd.n111 66.2847
R2448 vdd.n2685 vdd.n111 66.2847
R2449 vdd.n134 vdd.n111 66.2847
R2450 vdd.n2692 vdd.n111 66.2847
R2451 vdd.n127 vdd.n111 66.2847
R2452 vdd.n2699 vdd.n111 66.2847
R2453 vdd.n2702 vdd.n111 66.2847
R2454 vdd.n115 vdd.n111 66.2847
R2455 vdd.n116 vdd.n115 52.4337
R2456 vdd.n2702 vdd.n2701 52.4337
R2457 vdd.n2699 vdd.n2698 52.4337
R2458 vdd.n2694 vdd.n127 52.4337
R2459 vdd.n2692 vdd.n2691 52.4337
R2460 vdd.n2687 vdd.n134 52.4337
R2461 vdd.n2685 vdd.n2684 52.4337
R2462 vdd.n2680 vdd.n141 52.4337
R2463 vdd.n2678 vdd.n2677 52.4337
R2464 vdd.n2671 vdd.n149 52.4337
R2465 vdd.n2669 vdd.n2668 52.4337
R2466 vdd.n2664 vdd.n155 52.4337
R2467 vdd.n2662 vdd.n2661 52.4337
R2468 vdd.n2657 vdd.n162 52.4337
R2469 vdd.n2655 vdd.n2654 52.4337
R2470 vdd.n2650 vdd.n169 52.4337
R2471 vdd.n2648 vdd.n2647 52.4337
R2472 vdd.n2643 vdd.n176 52.4337
R2473 vdd.n2641 vdd.n2640 52.4337
R2474 vdd.n2634 vdd.n184 52.4337
R2475 vdd.n2632 vdd.n2631 52.4337
R2476 vdd.n2627 vdd.n190 52.4337
R2477 vdd.n2625 vdd.n2624 52.4337
R2478 vdd.n2620 vdd.n197 52.4337
R2479 vdd.n2618 vdd.n2617 52.4337
R2480 vdd.n2613 vdd.n204 52.4337
R2481 vdd.n2611 vdd.n2610 52.4337
R2482 vdd.n2606 vdd.n211 52.4337
R2483 vdd.n2604 vdd.n2603 52.4337
R2484 vdd.n2496 vdd.n2495 52.4337
R2485 vdd.n317 vdd.n289 52.4337
R2486 vdd.n2488 vdd.n290 52.4337
R2487 vdd.n325 vdd.n291 52.4337
R2488 vdd.n2481 vdd.n292 52.4337
R2489 vdd.n2478 vdd.n293 52.4337
R2490 vdd.n2474 vdd.n294 52.4337
R2491 vdd.n2470 vdd.n295 52.4337
R2492 vdd.n2466 vdd.n296 52.4337
R2493 vdd.n2458 vdd.n297 52.4337
R2494 vdd.n2454 vdd.n298 52.4337
R2495 vdd.n2450 vdd.n299 52.4337
R2496 vdd.n2446 vdd.n300 52.4337
R2497 vdd.n2442 vdd.n301 52.4337
R2498 vdd.n2438 vdd.n302 52.4337
R2499 vdd.n2434 vdd.n303 52.4337
R2500 vdd.n2430 vdd.n304 52.4337
R2501 vdd.n2426 vdd.n305 52.4337
R2502 vdd.n2422 vdd.n306 52.4337
R2503 vdd.n2416 vdd.n307 52.4337
R2504 vdd.n2412 vdd.n308 52.4337
R2505 vdd.n2408 vdd.n309 52.4337
R2506 vdd.n2404 vdd.n310 52.4337
R2507 vdd.n2400 vdd.n311 52.4337
R2508 vdd.n2396 vdd.n312 52.4337
R2509 vdd.n2372 vdd.n313 52.4337
R2510 vdd.n2389 vdd.n314 52.4337
R2511 vdd.n2386 vdd.n315 52.4337
R2512 vdd.n1405 vdd.n1229 52.4337
R2513 vdd.n1403 vdd.n1402 52.4337
R2514 vdd.n1235 vdd.n1234 52.4337
R2515 vdd.n1394 vdd.n1240 52.4337
R2516 vdd.n1392 vdd.n1391 52.4337
R2517 vdd.n1387 vdd.n1245 52.4337
R2518 vdd.n1385 vdd.n1384 52.4337
R2519 vdd.n1380 vdd.n1252 52.4337
R2520 vdd.n1378 vdd.n1377 52.4337
R2521 vdd.n1371 vdd.n1260 52.4337
R2522 vdd.n1369 vdd.n1368 52.4337
R2523 vdd.n1364 vdd.n1266 52.4337
R2524 vdd.n1362 vdd.n1361 52.4337
R2525 vdd.n1357 vdd.n1273 52.4337
R2526 vdd.n1355 vdd.n1354 52.4337
R2527 vdd.n1350 vdd.n1280 52.4337
R2528 vdd.n1348 vdd.n1347 52.4337
R2529 vdd.n1343 vdd.n1287 52.4337
R2530 vdd.n1341 vdd.n1340 52.4337
R2531 vdd.n1334 vdd.n1295 52.4337
R2532 vdd.n1332 vdd.n1331 52.4337
R2533 vdd.n1327 vdd.n1301 52.4337
R2534 vdd.n1325 vdd.n1324 52.4337
R2535 vdd.n1320 vdd.n1308 52.4337
R2536 vdd.n1318 vdd.n1317 52.4337
R2537 vdd.n1314 vdd.n1313 52.4337
R2538 vdd.n1310 vdd.n713 52.4337
R2539 vdd.n726 vdd.n715 52.4337
R2540 vdd.n1414 vdd.n722 52.4337
R2541 vdd.n1077 vdd.n1076 52.4337
R2542 vdd.n901 vdd.n873 52.4337
R2543 vdd.n905 vdd.n874 52.4337
R2544 vdd.n907 vdd.n875 52.4337
R2545 vdd.n911 vdd.n876 52.4337
R2546 vdd.n913 vdd.n877 52.4337
R2547 vdd.n917 vdd.n878 52.4337
R2548 vdd.n919 vdd.n879 52.4337
R2549 vdd.n1047 vdd.n880 52.4337
R2550 vdd.n924 vdd.n881 52.4337
R2551 vdd.n928 vdd.n882 52.4337
R2552 vdd.n930 vdd.n883 52.4337
R2553 vdd.n934 vdd.n884 52.4337
R2554 vdd.n936 vdd.n885 52.4337
R2555 vdd.n940 vdd.n886 52.4337
R2556 vdd.n942 vdd.n887 52.4337
R2557 vdd.n946 vdd.n888 52.4337
R2558 vdd.n948 vdd.n889 52.4337
R2559 vdd.n1014 vdd.n890 52.4337
R2560 vdd.n953 vdd.n891 52.4337
R2561 vdd.n957 vdd.n892 52.4337
R2562 vdd.n959 vdd.n893 52.4337
R2563 vdd.n963 vdd.n894 52.4337
R2564 vdd.n965 vdd.n895 52.4337
R2565 vdd.n969 vdd.n896 52.4337
R2566 vdd.n971 vdd.n897 52.4337
R2567 vdd.n975 vdd.n898 52.4337
R2568 vdd.n977 vdd.n899 52.4337
R2569 vdd.n1076 vdd.n872 52.4337
R2570 vdd.n904 vdd.n873 52.4337
R2571 vdd.n906 vdd.n874 52.4337
R2572 vdd.n910 vdd.n875 52.4337
R2573 vdd.n912 vdd.n876 52.4337
R2574 vdd.n916 vdd.n877 52.4337
R2575 vdd.n918 vdd.n878 52.4337
R2576 vdd.n922 vdd.n879 52.4337
R2577 vdd.n923 vdd.n880 52.4337
R2578 vdd.n927 vdd.n881 52.4337
R2579 vdd.n929 vdd.n882 52.4337
R2580 vdd.n933 vdd.n883 52.4337
R2581 vdd.n935 vdd.n884 52.4337
R2582 vdd.n939 vdd.n885 52.4337
R2583 vdd.n941 vdd.n886 52.4337
R2584 vdd.n945 vdd.n887 52.4337
R2585 vdd.n947 vdd.n888 52.4337
R2586 vdd.n951 vdd.n889 52.4337
R2587 vdd.n952 vdd.n890 52.4337
R2588 vdd.n956 vdd.n891 52.4337
R2589 vdd.n958 vdd.n892 52.4337
R2590 vdd.n962 vdd.n893 52.4337
R2591 vdd.n964 vdd.n894 52.4337
R2592 vdd.n968 vdd.n895 52.4337
R2593 vdd.n970 vdd.n896 52.4337
R2594 vdd.n974 vdd.n897 52.4337
R2595 vdd.n976 vdd.n898 52.4337
R2596 vdd.n980 vdd.n899 52.4337
R2597 vdd.n722 vdd.n721 52.4337
R2598 vdd.n726 vdd.n714 52.4337
R2599 vdd.n1311 vdd.n1310 52.4337
R2600 vdd.n1315 vdd.n1314 52.4337
R2601 vdd.n1319 vdd.n1318 52.4337
R2602 vdd.n1308 vdd.n1302 52.4337
R2603 vdd.n1326 vdd.n1325 52.4337
R2604 vdd.n1301 vdd.n1296 52.4337
R2605 vdd.n1333 vdd.n1332 52.4337
R2606 vdd.n1295 vdd.n1288 52.4337
R2607 vdd.n1342 vdd.n1341 52.4337
R2608 vdd.n1287 vdd.n1281 52.4337
R2609 vdd.n1349 vdd.n1348 52.4337
R2610 vdd.n1280 vdd.n1274 52.4337
R2611 vdd.n1356 vdd.n1355 52.4337
R2612 vdd.n1273 vdd.n1267 52.4337
R2613 vdd.n1363 vdd.n1362 52.4337
R2614 vdd.n1266 vdd.n1261 52.4337
R2615 vdd.n1370 vdd.n1369 52.4337
R2616 vdd.n1260 vdd.n1253 52.4337
R2617 vdd.n1379 vdd.n1378 52.4337
R2618 vdd.n1252 vdd.n1246 52.4337
R2619 vdd.n1386 vdd.n1385 52.4337
R2620 vdd.n1245 vdd.n1241 52.4337
R2621 vdd.n1393 vdd.n1392 52.4337
R2622 vdd.n1240 vdd.n1239 52.4337
R2623 vdd.n1234 vdd.n1230 52.4337
R2624 vdd.n1404 vdd.n1403 52.4337
R2625 vdd.n1229 vdd.n729 52.4337
R2626 vdd.n2495 vdd.n287 52.4337
R2627 vdd.n2489 vdd.n289 52.4337
R2628 vdd.n324 vdd.n290 52.4337
R2629 vdd.n327 vdd.n291 52.4337
R2630 vdd.n2479 vdd.n292 52.4337
R2631 vdd.n2475 vdd.n293 52.4337
R2632 vdd.n2471 vdd.n294 52.4337
R2633 vdd.n2467 vdd.n295 52.4337
R2634 vdd.n2457 vdd.n296 52.4337
R2635 vdd.n2455 vdd.n297 52.4337
R2636 vdd.n2451 vdd.n298 52.4337
R2637 vdd.n2447 vdd.n299 52.4337
R2638 vdd.n2443 vdd.n300 52.4337
R2639 vdd.n2439 vdd.n301 52.4337
R2640 vdd.n2435 vdd.n302 52.4337
R2641 vdd.n2431 vdd.n303 52.4337
R2642 vdd.n2427 vdd.n304 52.4337
R2643 vdd.n2423 vdd.n305 52.4337
R2644 vdd.n2415 vdd.n306 52.4337
R2645 vdd.n2413 vdd.n307 52.4337
R2646 vdd.n2409 vdd.n308 52.4337
R2647 vdd.n2405 vdd.n309 52.4337
R2648 vdd.n2401 vdd.n310 52.4337
R2649 vdd.n2397 vdd.n311 52.4337
R2650 vdd.n2371 vdd.n312 52.4337
R2651 vdd.n2374 vdd.n313 52.4337
R2652 vdd.n2387 vdd.n314 52.4337
R2653 vdd.n2383 vdd.n315 52.4337
R2654 vdd.n2605 vdd.n2604 52.4337
R2655 vdd.n211 vdd.n205 52.4337
R2656 vdd.n2612 vdd.n2611 52.4337
R2657 vdd.n204 vdd.n198 52.4337
R2658 vdd.n2619 vdd.n2618 52.4337
R2659 vdd.n197 vdd.n191 52.4337
R2660 vdd.n2626 vdd.n2625 52.4337
R2661 vdd.n190 vdd.n185 52.4337
R2662 vdd.n2633 vdd.n2632 52.4337
R2663 vdd.n184 vdd.n177 52.4337
R2664 vdd.n2642 vdd.n2641 52.4337
R2665 vdd.n176 vdd.n170 52.4337
R2666 vdd.n2649 vdd.n2648 52.4337
R2667 vdd.n169 vdd.n163 52.4337
R2668 vdd.n2656 vdd.n2655 52.4337
R2669 vdd.n162 vdd.n156 52.4337
R2670 vdd.n2663 vdd.n2662 52.4337
R2671 vdd.n155 vdd.n150 52.4337
R2672 vdd.n2670 vdd.n2669 52.4337
R2673 vdd.n149 vdd.n142 52.4337
R2674 vdd.n2679 vdd.n2678 52.4337
R2675 vdd.n141 vdd.n135 52.4337
R2676 vdd.n2686 vdd.n2685 52.4337
R2677 vdd.n134 vdd.n128 52.4337
R2678 vdd.n2693 vdd.n2692 52.4337
R2679 vdd.n127 vdd.n120 52.4337
R2680 vdd.n2700 vdd.n2699 52.4337
R2681 vdd.n2703 vdd.n2702 52.4337
R2682 vdd.n115 vdd.n112 52.4337
R2683 vdd.n2340 vdd.n390 39.2114
R2684 vdd.n2338 vdd.n2337 39.2114
R2685 vdd.n2333 vdd.n393 39.2114
R2686 vdd.n2331 vdd.n2330 39.2114
R2687 vdd.n2326 vdd.n396 39.2114
R2688 vdd.n2324 vdd.n2323 39.2114
R2689 vdd.n2319 vdd.n2318 39.2114
R2690 vdd.n2314 vdd.n399 39.2114
R2691 vdd.n2312 vdd.n2311 39.2114
R2692 vdd.n2307 vdd.n402 39.2114
R2693 vdd.n2305 vdd.n2304 39.2114
R2694 vdd.n2299 vdd.n407 39.2114
R2695 vdd.n2297 vdd.n2296 39.2114
R2696 vdd.n1918 vdd.n522 39.2114
R2697 vdd.n1924 vdd.n1923 39.2114
R2698 vdd.n1927 vdd.n1926 39.2114
R2699 vdd.n1932 vdd.n1931 39.2114
R2700 vdd.n1935 vdd.n1934 39.2114
R2701 vdd.n1940 vdd.n1939 39.2114
R2702 vdd.n1943 vdd.n1942 39.2114
R2703 vdd.n1948 vdd.n1947 39.2114
R2704 vdd.n1951 vdd.n1950 39.2114
R2705 vdd.n1956 vdd.n1955 39.2114
R2706 vdd.n1959 vdd.n1958 39.2114
R2707 vdd.n1965 vdd.n1964 39.2114
R2708 vdd.n1821 vdd.n524 39.2114
R2709 vdd.n1817 vdd.n525 39.2114
R2710 vdd.n1813 vdd.n526 39.2114
R2711 vdd.n1809 vdd.n527 39.2114
R2712 vdd.n1805 vdd.n528 39.2114
R2713 vdd.n1801 vdd.n529 39.2114
R2714 vdd.n1797 vdd.n530 39.2114
R2715 vdd.n1793 vdd.n531 39.2114
R2716 vdd.n1789 vdd.n532 39.2114
R2717 vdd.n1785 vdd.n533 39.2114
R2718 vdd.n1781 vdd.n534 39.2114
R2719 vdd.n1776 vdd.n535 39.2114
R2720 vdd.n1772 vdd.n536 39.2114
R2721 vdd.n1643 vdd.n682 39.2114
R2722 vdd.n1641 vdd.n684 39.2114
R2723 vdd.n1637 vdd.n1636 39.2114
R2724 vdd.n1630 vdd.n686 39.2114
R2725 vdd.n1629 vdd.n1628 39.2114
R2726 vdd.n1622 vdd.n688 39.2114
R2727 vdd.n1621 vdd.n690 39.2114
R2728 vdd.n1617 vdd.n1616 39.2114
R2729 vdd.n1610 vdd.n692 39.2114
R2730 vdd.n1609 vdd.n1608 39.2114
R2731 vdd.n1602 vdd.n694 39.2114
R2732 vdd.n1601 vdd.n698 39.2114
R2733 vdd.n2274 vdd.n2273 39.2114
R2734 vdd.n2271 vdd.n2270 39.2114
R2735 vdd.n2266 vdd.n2250 39.2114
R2736 vdd.n2264 vdd.n2263 39.2114
R2737 vdd.n2259 vdd.n2253 39.2114
R2738 vdd.n2257 vdd.n2256 39.2114
R2739 vdd.n2368 vdd.n369 39.2114
R2740 vdd.n2366 vdd.n2365 39.2114
R2741 vdd.n2361 vdd.n372 39.2114
R2742 vdd.n2359 vdd.n2358 39.2114
R2743 vdd.n2354 vdd.n375 39.2114
R2744 vdd.n2352 vdd.n2351 39.2114
R2745 vdd.n2347 vdd.n381 39.2114
R2746 vdd.n2133 vdd.n1887 39.2114
R2747 vdd.n2132 vdd.n2131 39.2114
R2748 vdd.n2125 vdd.n1889 39.2114
R2749 vdd.n2124 vdd.n2123 39.2114
R2750 vdd.n2117 vdd.n1891 39.2114
R2751 vdd.n2116 vdd.n2115 39.2114
R2752 vdd.n2109 vdd.n1893 39.2114
R2753 vdd.n2108 vdd.n2107 39.2114
R2754 vdd.n2101 vdd.n1895 39.2114
R2755 vdd.n2100 vdd.n2099 39.2114
R2756 vdd.n2093 vdd.n1897 39.2114
R2757 vdd.n2092 vdd.n2091 39.2114
R2758 vdd.n2085 vdd.n1899 39.2114
R2759 vdd.n2134 vdd.n2133 39.2114
R2760 vdd.n2131 vdd.n2130 39.2114
R2761 vdd.n2126 vdd.n2125 39.2114
R2762 vdd.n2123 vdd.n2122 39.2114
R2763 vdd.n2118 vdd.n2117 39.2114
R2764 vdd.n2115 vdd.n2114 39.2114
R2765 vdd.n2110 vdd.n2109 39.2114
R2766 vdd.n2107 vdd.n2106 39.2114
R2767 vdd.n2102 vdd.n2101 39.2114
R2768 vdd.n2099 vdd.n2098 39.2114
R2769 vdd.n2094 vdd.n2093 39.2114
R2770 vdd.n2091 vdd.n2090 39.2114
R2771 vdd.n2086 vdd.n2085 39.2114
R2772 vdd.n381 vdd.n376 39.2114
R2773 vdd.n2353 vdd.n2352 39.2114
R2774 vdd.n375 vdd.n373 39.2114
R2775 vdd.n2360 vdd.n2359 39.2114
R2776 vdd.n372 vdd.n370 39.2114
R2777 vdd.n2367 vdd.n2366 39.2114
R2778 vdd.n2254 vdd.n369 39.2114
R2779 vdd.n2258 vdd.n2257 39.2114
R2780 vdd.n2253 vdd.n2251 39.2114
R2781 vdd.n2265 vdd.n2264 39.2114
R2782 vdd.n2250 vdd.n2248 39.2114
R2783 vdd.n2272 vdd.n2271 39.2114
R2784 vdd.n2275 vdd.n2274 39.2114
R2785 vdd.n1644 vdd.n1643 39.2114
R2786 vdd.n1638 vdd.n684 39.2114
R2787 vdd.n1636 vdd.n1635 39.2114
R2788 vdd.n1631 vdd.n1630 39.2114
R2789 vdd.n1628 vdd.n1627 39.2114
R2790 vdd.n1623 vdd.n1622 39.2114
R2791 vdd.n1618 vdd.n690 39.2114
R2792 vdd.n1616 vdd.n1615 39.2114
R2793 vdd.n1611 vdd.n1610 39.2114
R2794 vdd.n1608 vdd.n1607 39.2114
R2795 vdd.n1603 vdd.n1602 39.2114
R2796 vdd.n1598 vdd.n698 39.2114
R2797 vdd.n1775 vdd.n536 39.2114
R2798 vdd.n1780 vdd.n535 39.2114
R2799 vdd.n1784 vdd.n534 39.2114
R2800 vdd.n1788 vdd.n533 39.2114
R2801 vdd.n1792 vdd.n532 39.2114
R2802 vdd.n1796 vdd.n531 39.2114
R2803 vdd.n1800 vdd.n530 39.2114
R2804 vdd.n1804 vdd.n529 39.2114
R2805 vdd.n1808 vdd.n528 39.2114
R2806 vdd.n1812 vdd.n527 39.2114
R2807 vdd.n1816 vdd.n526 39.2114
R2808 vdd.n1820 vdd.n525 39.2114
R2809 vdd.n1823 vdd.n524 39.2114
R2810 vdd.n1919 vdd.n1918 39.2114
R2811 vdd.n1925 vdd.n1924 39.2114
R2812 vdd.n1926 vdd.n1915 39.2114
R2813 vdd.n1933 vdd.n1932 39.2114
R2814 vdd.n1934 vdd.n1913 39.2114
R2815 vdd.n1941 vdd.n1940 39.2114
R2816 vdd.n1942 vdd.n1911 39.2114
R2817 vdd.n1949 vdd.n1948 39.2114
R2818 vdd.n1950 vdd.n1909 39.2114
R2819 vdd.n1957 vdd.n1956 39.2114
R2820 vdd.n1958 vdd.n1905 39.2114
R2821 vdd.n1966 vdd.n1965 39.2114
R2822 vdd.n2298 vdd.n2297 39.2114
R2823 vdd.n407 vdd.n403 39.2114
R2824 vdd.n2306 vdd.n2305 39.2114
R2825 vdd.n402 vdd.n400 39.2114
R2826 vdd.n2313 vdd.n2312 39.2114
R2827 vdd.n399 vdd.n397 39.2114
R2828 vdd.n2320 vdd.n2319 39.2114
R2829 vdd.n2325 vdd.n2324 39.2114
R2830 vdd.n396 vdd.n394 39.2114
R2831 vdd.n2332 vdd.n2331 39.2114
R2832 vdd.n393 vdd.n391 39.2114
R2833 vdd.n2339 vdd.n2338 39.2114
R2834 vdd.n390 vdd.n387 39.2114
R2835 vdd.n551 vdd.n537 39.2114
R2836 vdd.n1876 vdd.n538 39.2114
R2837 vdd.n1872 vdd.n539 39.2114
R2838 vdd.n1868 vdd.n540 39.2114
R2839 vdd.n1864 vdd.n541 39.2114
R2840 vdd.n1860 vdd.n542 39.2114
R2841 vdd.n1856 vdd.n543 39.2114
R2842 vdd.n1852 vdd.n544 39.2114
R2843 vdd.n1848 vdd.n545 39.2114
R2844 vdd.n1844 vdd.n546 39.2114
R2845 vdd.n1840 vdd.n547 39.2114
R2846 vdd.n1836 vdd.n548 39.2114
R2847 vdd.n1432 vdd.n1431 39.2114
R2848 vdd.n1437 vdd.n1436 39.2114
R2849 vdd.n1440 vdd.n1439 39.2114
R2850 vdd.n1445 vdd.n1444 39.2114
R2851 vdd.n1448 vdd.n1447 39.2114
R2852 vdd.n1453 vdd.n1452 39.2114
R2853 vdd.n1456 vdd.n1455 39.2114
R2854 vdd.n1461 vdd.n1460 39.2114
R2855 vdd.n1464 vdd.n1463 39.2114
R2856 vdd.n1469 vdd.n1468 39.2114
R2857 vdd.n1472 vdd.n1471 39.2114
R2858 vdd.n1478 vdd.n1477 39.2114
R2859 vdd.n1833 vdd.n548 39.2114
R2860 vdd.n1837 vdd.n547 39.2114
R2861 vdd.n1841 vdd.n546 39.2114
R2862 vdd.n1845 vdd.n545 39.2114
R2863 vdd.n1849 vdd.n544 39.2114
R2864 vdd.n1853 vdd.n543 39.2114
R2865 vdd.n1857 vdd.n542 39.2114
R2866 vdd.n1861 vdd.n541 39.2114
R2867 vdd.n1865 vdd.n540 39.2114
R2868 vdd.n1869 vdd.n539 39.2114
R2869 vdd.n1873 vdd.n538 39.2114
R2870 vdd.n1877 vdd.n537 39.2114
R2871 vdd.n1431 vdd.n1430 39.2114
R2872 vdd.n1438 vdd.n1437 39.2114
R2873 vdd.n1439 vdd.n1428 39.2114
R2874 vdd.n1446 vdd.n1445 39.2114
R2875 vdd.n1447 vdd.n1426 39.2114
R2876 vdd.n1454 vdd.n1453 39.2114
R2877 vdd.n1455 vdd.n707 39.2114
R2878 vdd.n1462 vdd.n1461 39.2114
R2879 vdd.n1463 vdd.n705 39.2114
R2880 vdd.n1470 vdd.n1469 39.2114
R2881 vdd.n1471 vdd.n701 39.2114
R2882 vdd.n1479 vdd.n1478 39.2114
R2883 vdd.n984 vdd.n983 37.4308
R2884 vdd.n1017 vdd.n1016 37.4308
R2885 vdd.n1050 vdd.n1049 37.4308
R2886 vdd.n720 vdd.n719 37.4308
R2887 vdd.n1339 vdd.n1291 37.4308
R2888 vdd.n1376 vdd.n1256 37.4308
R2889 vdd.n214 vdd.n213 37.4308
R2890 vdd.n2639 vdd.n180 37.4308
R2891 vdd.n2676 vdd.n145 37.4308
R2892 vdd.n2421 vdd.n355 37.4308
R2893 vdd.n2465 vdd.n2464 37.4308
R2894 vdd.n2382 vdd.n2381 37.4308
R2895 vdd.n1647 vdd.n1646 31.3761
R2896 vdd.n1825 vdd.n1824 31.3761
R2897 vdd.n1773 vdd.n1770 31.3761
R2898 vdd.n1596 vdd.n1595 31.3761
R2899 vdd.n1969 vdd.n1968 31.3761
R2900 vdd.n2295 vdd.n2294 31.3761
R2901 vdd.n2141 vdd.n521 31.3761
R2902 vdd.n2343 vdd.n2342 31.3761
R2903 vdd.n2277 vdd.n2276 31.3761
R2904 vdd.n2348 vdd.n380 31.3761
R2905 vdd.n2087 vdd.n2084 31.3761
R2906 vdd.n2137 vdd.n2136 31.3761
R2907 vdd.n1651 vdd.n677 31.3761
R2908 vdd.n1880 vdd.n552 31.3761
R2909 vdd.n1832 vdd.n1831 31.3761
R2910 vdd.n1482 vdd.n1481 31.3761
R2911 vdd.n1475 vdd.n703 30.449
R2912 vdd.n555 vdd.n554 30.449
R2913 vdd.n697 vdd.n696 30.449
R2914 vdd.n1778 vdd.n564 30.449
R2915 vdd.n1902 vdd.n1901 30.449
R2916 vdd.n2301 vdd.n405 30.449
R2917 vdd.n1962 vdd.n1907 30.449
R2918 vdd.n379 vdd.n378 30.449
R2919 vdd.n703 vdd.n702 25.7944
R2920 vdd.n554 vdd.n553 25.7944
R2921 vdd.n983 vdd.n982 25.7944
R2922 vdd.n1016 vdd.n1015 25.7944
R2923 vdd.n1049 vdd.n1048 25.7944
R2924 vdd.n719 vdd.n718 25.7944
R2925 vdd.n1291 vdd.n1290 25.7944
R2926 vdd.n1256 vdd.n1255 25.7944
R2927 vdd.n696 vdd.n695 25.7944
R2928 vdd.n564 vdd.n563 25.7944
R2929 vdd.n1901 vdd.n1900 25.7944
R2930 vdd.n213 vdd.n212 25.7944
R2931 vdd.n180 vdd.n179 25.7944
R2932 vdd.n145 vdd.n144 25.7944
R2933 vdd.n355 vdd.n354 25.7944
R2934 vdd.n2464 vdd.n2463 25.7944
R2935 vdd.n405 vdd.n404 25.7944
R2936 vdd.n1907 vdd.n1906 25.7944
R2937 vdd.n2381 vdd.n2380 25.7944
R2938 vdd.n378 vdd.n377 25.7944
R2939 vdd.n1075 vdd.n867 22.6677
R2940 vdd.n1412 vdd.n727 22.6677
R2941 vdd.n2494 vdd.n282 22.6677
R2942 vdd.n2711 vdd.n111 22.6677
R2943 vdd.n1086 vdd.n865 19.3944
R2944 vdd.n1086 vdd.n863 19.3944
R2945 vdd.n1090 vdd.n863 19.3944
R2946 vdd.n1090 vdd.n852 19.3944
R2947 vdd.n1102 vdd.n852 19.3944
R2948 vdd.n1102 vdd.n850 19.3944
R2949 vdd.n1106 vdd.n850 19.3944
R2950 vdd.n1106 vdd.n841 19.3944
R2951 vdd.n1118 vdd.n841 19.3944
R2952 vdd.n1118 vdd.n839 19.3944
R2953 vdd.n1122 vdd.n839 19.3944
R2954 vdd.n1122 vdd.n828 19.3944
R2955 vdd.n1134 vdd.n828 19.3944
R2956 vdd.n1134 vdd.n826 19.3944
R2957 vdd.n1138 vdd.n826 19.3944
R2958 vdd.n1138 vdd.n817 19.3944
R2959 vdd.n1151 vdd.n817 19.3944
R2960 vdd.n1151 vdd.n815 19.3944
R2961 vdd.n1155 vdd.n815 19.3944
R2962 vdd.n1155 vdd.n774 19.3944
R2963 vdd.n1167 vdd.n774 19.3944
R2964 vdd.n1167 vdd.n772 19.3944
R2965 vdd.n1171 vdd.n772 19.3944
R2966 vdd.n1171 vdd.n763 19.3944
R2967 vdd.n1183 vdd.n763 19.3944
R2968 vdd.n1183 vdd.n761 19.3944
R2969 vdd.n1187 vdd.n761 19.3944
R2970 vdd.n1187 vdd.n750 19.3944
R2971 vdd.n1199 vdd.n750 19.3944
R2972 vdd.n1199 vdd.n748 19.3944
R2973 vdd.n1203 vdd.n748 19.3944
R2974 vdd.n1203 vdd.n739 19.3944
R2975 vdd.n1215 vdd.n739 19.3944
R2976 vdd.n1215 vdd.n736 19.3944
R2977 vdd.n1220 vdd.n736 19.3944
R2978 vdd.n1220 vdd.n737 19.3944
R2979 vdd.n737 vdd.n724 19.3944
R2980 vdd.n1013 vdd.n954 19.3944
R2981 vdd.n1009 vdd.n954 19.3944
R2982 vdd.n1009 vdd.n1008 19.3944
R2983 vdd.n1008 vdd.n1007 19.3944
R2984 vdd.n1007 vdd.n960 19.3944
R2985 vdd.n1003 vdd.n960 19.3944
R2986 vdd.n1003 vdd.n1002 19.3944
R2987 vdd.n1002 vdd.n1001 19.3944
R2988 vdd.n1001 vdd.n966 19.3944
R2989 vdd.n997 vdd.n966 19.3944
R2990 vdd.n997 vdd.n996 19.3944
R2991 vdd.n996 vdd.n995 19.3944
R2992 vdd.n995 vdd.n972 19.3944
R2993 vdd.n991 vdd.n972 19.3944
R2994 vdd.n991 vdd.n990 19.3944
R2995 vdd.n990 vdd.n989 19.3944
R2996 vdd.n989 vdd.n978 19.3944
R2997 vdd.n985 vdd.n978 19.3944
R2998 vdd.n1046 vdd.n925 19.3944
R2999 vdd.n1042 vdd.n925 19.3944
R3000 vdd.n1042 vdd.n1041 19.3944
R3001 vdd.n1041 vdd.n1040 19.3944
R3002 vdd.n1040 vdd.n931 19.3944
R3003 vdd.n1036 vdd.n931 19.3944
R3004 vdd.n1036 vdd.n1035 19.3944
R3005 vdd.n1035 vdd.n1034 19.3944
R3006 vdd.n1034 vdd.n937 19.3944
R3007 vdd.n1030 vdd.n937 19.3944
R3008 vdd.n1030 vdd.n1029 19.3944
R3009 vdd.n1029 vdd.n1028 19.3944
R3010 vdd.n1028 vdd.n943 19.3944
R3011 vdd.n1024 vdd.n943 19.3944
R3012 vdd.n1024 vdd.n1023 19.3944
R3013 vdd.n1023 vdd.n1022 19.3944
R3014 vdd.n1022 vdd.n949 19.3944
R3015 vdd.n1018 vdd.n949 19.3944
R3016 vdd.n1078 vdd.n871 19.3944
R3017 vdd.n1073 vdd.n871 19.3944
R3018 vdd.n1073 vdd.n902 19.3944
R3019 vdd.n1069 vdd.n902 19.3944
R3020 vdd.n1069 vdd.n1068 19.3944
R3021 vdd.n1068 vdd.n1067 19.3944
R3022 vdd.n1067 vdd.n908 19.3944
R3023 vdd.n1063 vdd.n908 19.3944
R3024 vdd.n1063 vdd.n1062 19.3944
R3025 vdd.n1062 vdd.n1061 19.3944
R3026 vdd.n1061 vdd.n914 19.3944
R3027 vdd.n1057 vdd.n914 19.3944
R3028 vdd.n1057 vdd.n1056 19.3944
R3029 vdd.n1056 vdd.n1055 19.3944
R3030 vdd.n1055 vdd.n920 19.3944
R3031 vdd.n1051 vdd.n920 19.3944
R3032 vdd.n1335 vdd.n1289 19.3944
R3033 vdd.n1335 vdd.n1294 19.3944
R3034 vdd.n1330 vdd.n1294 19.3944
R3035 vdd.n1330 vdd.n1329 19.3944
R3036 vdd.n1329 vdd.n1328 19.3944
R3037 vdd.n1328 vdd.n1300 19.3944
R3038 vdd.n1323 vdd.n1300 19.3944
R3039 vdd.n1323 vdd.n1322 19.3944
R3040 vdd.n1322 vdd.n1321 19.3944
R3041 vdd.n1321 vdd.n1307 19.3944
R3042 vdd.n1316 vdd.n1307 19.3944
R3043 vdd.n1312 vdd.n1309 19.3944
R3044 vdd.n1421 vdd.n712 19.3944
R3045 vdd.n1421 vdd.n1420 19.3944
R3046 vdd.n1420 vdd.n1419 19.3944
R3047 vdd.n1419 vdd.n716 19.3944
R3048 vdd.n1372 vdd.n1254 19.3944
R3049 vdd.n1372 vdd.n1259 19.3944
R3050 vdd.n1367 vdd.n1259 19.3944
R3051 vdd.n1367 vdd.n1366 19.3944
R3052 vdd.n1366 vdd.n1365 19.3944
R3053 vdd.n1365 vdd.n1265 19.3944
R3054 vdd.n1360 vdd.n1265 19.3944
R3055 vdd.n1360 vdd.n1359 19.3944
R3056 vdd.n1359 vdd.n1358 19.3944
R3057 vdd.n1358 vdd.n1272 19.3944
R3058 vdd.n1353 vdd.n1272 19.3944
R3059 vdd.n1353 vdd.n1352 19.3944
R3060 vdd.n1352 vdd.n1351 19.3944
R3061 vdd.n1351 vdd.n1279 19.3944
R3062 vdd.n1346 vdd.n1279 19.3944
R3063 vdd.n1346 vdd.n1345 19.3944
R3064 vdd.n1345 vdd.n1344 19.3944
R3065 vdd.n1344 vdd.n1286 19.3944
R3066 vdd.n1407 vdd.n1406 19.3944
R3067 vdd.n1406 vdd.n1228 19.3944
R3068 vdd.n1401 vdd.n1228 19.3944
R3069 vdd.n1401 vdd.n1400 19.3944
R3070 vdd.n1400 vdd.n1399 19.3944
R3071 vdd.n1395 vdd.n1236 19.3944
R3072 vdd.n1390 vdd.n1238 19.3944
R3073 vdd.n1390 vdd.n1389 19.3944
R3074 vdd.n1389 vdd.n1388 19.3944
R3075 vdd.n1388 vdd.n1244 19.3944
R3076 vdd.n1383 vdd.n1244 19.3944
R3077 vdd.n1383 vdd.n1382 19.3944
R3078 vdd.n1382 vdd.n1381 19.3944
R3079 vdd.n1381 vdd.n1251 19.3944
R3080 vdd.n1082 vdd.n869 19.3944
R3081 vdd.n1082 vdd.n859 19.3944
R3082 vdd.n1094 vdd.n859 19.3944
R3083 vdd.n1094 vdd.n857 19.3944
R3084 vdd.n1098 vdd.n857 19.3944
R3085 vdd.n1098 vdd.n847 19.3944
R3086 vdd.n1110 vdd.n847 19.3944
R3087 vdd.n1110 vdd.n845 19.3944
R3088 vdd.n1114 vdd.n845 19.3944
R3089 vdd.n1114 vdd.n835 19.3944
R3090 vdd.n1126 vdd.n835 19.3944
R3091 vdd.n1126 vdd.n833 19.3944
R3092 vdd.n1130 vdd.n833 19.3944
R3093 vdd.n1130 vdd.n823 19.3944
R3094 vdd.n1142 vdd.n823 19.3944
R3095 vdd.n1142 vdd.n821 19.3944
R3096 vdd.n1147 vdd.n821 19.3944
R3097 vdd.n1147 vdd.n811 19.3944
R3098 vdd.n1159 vdd.n811 19.3944
R3099 vdd.n1159 vdd.n779 19.3944
R3100 vdd.n1163 vdd.n779 19.3944
R3101 vdd.n1163 vdd.n769 19.3944
R3102 vdd.n1175 vdd.n769 19.3944
R3103 vdd.n1175 vdd.n767 19.3944
R3104 vdd.n1179 vdd.n767 19.3944
R3105 vdd.n1179 vdd.n757 19.3944
R3106 vdd.n1191 vdd.n757 19.3944
R3107 vdd.n1191 vdd.n755 19.3944
R3108 vdd.n1195 vdd.n755 19.3944
R3109 vdd.n1195 vdd.n745 19.3944
R3110 vdd.n1207 vdd.n745 19.3944
R3111 vdd.n1207 vdd.n743 19.3944
R3112 vdd.n1211 vdd.n743 19.3944
R3113 vdd.n1211 vdd.n732 19.3944
R3114 vdd.n1224 vdd.n732 19.3944
R3115 vdd.n1224 vdd.n730 19.3944
R3116 vdd.n1410 vdd.n730 19.3944
R3117 vdd.n2505 vdd.n280 19.3944
R3118 vdd.n2505 vdd.n278 19.3944
R3119 vdd.n2509 vdd.n278 19.3944
R3120 vdd.n2509 vdd.n267 19.3944
R3121 vdd.n2521 vdd.n267 19.3944
R3122 vdd.n2521 vdd.n265 19.3944
R3123 vdd.n2525 vdd.n265 19.3944
R3124 vdd.n2525 vdd.n256 19.3944
R3125 vdd.n2537 vdd.n256 19.3944
R3126 vdd.n2537 vdd.n254 19.3944
R3127 vdd.n2541 vdd.n254 19.3944
R3128 vdd.n2541 vdd.n243 19.3944
R3129 vdd.n2553 vdd.n243 19.3944
R3130 vdd.n2553 vdd.n241 19.3944
R3131 vdd.n2557 vdd.n241 19.3944
R3132 vdd.n2557 vdd.n231 19.3944
R3133 vdd.n2569 vdd.n231 19.3944
R3134 vdd.n2569 vdd.n229 19.3944
R3135 vdd.n2573 vdd.n229 19.3944
R3136 vdd.n2574 vdd.n2573 19.3944
R3137 vdd.n2575 vdd.n2574 19.3944
R3138 vdd.n2575 vdd.n227 19.3944
R3139 vdd.n2579 vdd.n227 19.3944
R3140 vdd.n2580 vdd.n2579 19.3944
R3141 vdd.n2581 vdd.n2580 19.3944
R3142 vdd.n2581 vdd.n224 19.3944
R3143 vdd.n2585 vdd.n224 19.3944
R3144 vdd.n2586 vdd.n2585 19.3944
R3145 vdd.n2587 vdd.n2586 19.3944
R3146 vdd.n2587 vdd.n221 19.3944
R3147 vdd.n2591 vdd.n221 19.3944
R3148 vdd.n2592 vdd.n2591 19.3944
R3149 vdd.n2593 vdd.n2592 19.3944
R3150 vdd.n2593 vdd.n218 19.3944
R3151 vdd.n2597 vdd.n218 19.3944
R3152 vdd.n2598 vdd.n2597 19.3944
R3153 vdd.n2599 vdd.n2598 19.3944
R3154 vdd.n2635 vdd.n178 19.3944
R3155 vdd.n2635 vdd.n183 19.3944
R3156 vdd.n2630 vdd.n183 19.3944
R3157 vdd.n2630 vdd.n2629 19.3944
R3158 vdd.n2629 vdd.n2628 19.3944
R3159 vdd.n2628 vdd.n189 19.3944
R3160 vdd.n2623 vdd.n189 19.3944
R3161 vdd.n2623 vdd.n2622 19.3944
R3162 vdd.n2622 vdd.n2621 19.3944
R3163 vdd.n2621 vdd.n196 19.3944
R3164 vdd.n2616 vdd.n196 19.3944
R3165 vdd.n2616 vdd.n2615 19.3944
R3166 vdd.n2615 vdd.n2614 19.3944
R3167 vdd.n2614 vdd.n203 19.3944
R3168 vdd.n2609 vdd.n203 19.3944
R3169 vdd.n2609 vdd.n2608 19.3944
R3170 vdd.n2608 vdd.n2607 19.3944
R3171 vdd.n2607 vdd.n210 19.3944
R3172 vdd.n2672 vdd.n143 19.3944
R3173 vdd.n2672 vdd.n148 19.3944
R3174 vdd.n2667 vdd.n148 19.3944
R3175 vdd.n2667 vdd.n2666 19.3944
R3176 vdd.n2666 vdd.n2665 19.3944
R3177 vdd.n2665 vdd.n154 19.3944
R3178 vdd.n2660 vdd.n154 19.3944
R3179 vdd.n2660 vdd.n2659 19.3944
R3180 vdd.n2659 vdd.n2658 19.3944
R3181 vdd.n2658 vdd.n161 19.3944
R3182 vdd.n2653 vdd.n161 19.3944
R3183 vdd.n2653 vdd.n2652 19.3944
R3184 vdd.n2652 vdd.n2651 19.3944
R3185 vdd.n2651 vdd.n168 19.3944
R3186 vdd.n2646 vdd.n168 19.3944
R3187 vdd.n2646 vdd.n2645 19.3944
R3188 vdd.n2645 vdd.n2644 19.3944
R3189 vdd.n2644 vdd.n175 19.3944
R3190 vdd.n2706 vdd.n2705 19.3944
R3191 vdd.n2705 vdd.n2704 19.3944
R3192 vdd.n2704 vdd.n118 19.3944
R3193 vdd.n119 vdd.n118 19.3944
R3194 vdd.n2697 vdd.n119 19.3944
R3195 vdd.n2697 vdd.n2696 19.3944
R3196 vdd.n2696 vdd.n2695 19.3944
R3197 vdd.n2695 vdd.n126 19.3944
R3198 vdd.n2690 vdd.n126 19.3944
R3199 vdd.n2690 vdd.n2689 19.3944
R3200 vdd.n2689 vdd.n2688 19.3944
R3201 vdd.n2688 vdd.n133 19.3944
R3202 vdd.n2683 vdd.n133 19.3944
R3203 vdd.n2683 vdd.n2682 19.3944
R3204 vdd.n2682 vdd.n2681 19.3944
R3205 vdd.n2681 vdd.n140 19.3944
R3206 vdd.n2501 vdd.n284 19.3944
R3207 vdd.n2501 vdd.n274 19.3944
R3208 vdd.n2513 vdd.n274 19.3944
R3209 vdd.n2513 vdd.n272 19.3944
R3210 vdd.n2517 vdd.n272 19.3944
R3211 vdd.n2517 vdd.n262 19.3944
R3212 vdd.n2529 vdd.n262 19.3944
R3213 vdd.n2529 vdd.n260 19.3944
R3214 vdd.n2533 vdd.n260 19.3944
R3215 vdd.n2533 vdd.n250 19.3944
R3216 vdd.n2545 vdd.n250 19.3944
R3217 vdd.n2545 vdd.n248 19.3944
R3218 vdd.n2549 vdd.n248 19.3944
R3219 vdd.n2549 vdd.n238 19.3944
R3220 vdd.n2561 vdd.n238 19.3944
R3221 vdd.n2561 vdd.n236 19.3944
R3222 vdd.n2565 vdd.n236 19.3944
R3223 vdd.n2565 vdd.n60 19.3944
R3224 vdd.n2747 vdd.n60 19.3944
R3225 vdd.n2747 vdd.n61 19.3944
R3226 vdd.n2741 vdd.n61 19.3944
R3227 vdd.n2741 vdd.n2740 19.3944
R3228 vdd.n2740 vdd.n2739 19.3944
R3229 vdd.n2739 vdd.n73 19.3944
R3230 vdd.n2733 vdd.n73 19.3944
R3231 vdd.n2733 vdd.n2732 19.3944
R3232 vdd.n2732 vdd.n2731 19.3944
R3233 vdd.n2731 vdd.n83 19.3944
R3234 vdd.n2725 vdd.n83 19.3944
R3235 vdd.n2725 vdd.n2724 19.3944
R3236 vdd.n2724 vdd.n2723 19.3944
R3237 vdd.n2723 vdd.n95 19.3944
R3238 vdd.n2717 vdd.n95 19.3944
R3239 vdd.n2717 vdd.n2716 19.3944
R3240 vdd.n2716 vdd.n2715 19.3944
R3241 vdd.n2715 vdd.n106 19.3944
R3242 vdd.n2709 vdd.n106 19.3944
R3243 vdd.n2459 vdd.n335 19.3944
R3244 vdd.n2459 vdd.n2456 19.3944
R3245 vdd.n2456 vdd.n2453 19.3944
R3246 vdd.n2453 vdd.n2452 19.3944
R3247 vdd.n2452 vdd.n2449 19.3944
R3248 vdd.n2449 vdd.n2448 19.3944
R3249 vdd.n2448 vdd.n2445 19.3944
R3250 vdd.n2445 vdd.n2444 19.3944
R3251 vdd.n2444 vdd.n2441 19.3944
R3252 vdd.n2441 vdd.n2440 19.3944
R3253 vdd.n2440 vdd.n2437 19.3944
R3254 vdd.n2437 vdd.n2436 19.3944
R3255 vdd.n2436 vdd.n2433 19.3944
R3256 vdd.n2433 vdd.n2432 19.3944
R3257 vdd.n2432 vdd.n2429 19.3944
R3258 vdd.n2429 vdd.n2428 19.3944
R3259 vdd.n2428 vdd.n2425 19.3944
R3260 vdd.n2425 vdd.n2424 19.3944
R3261 vdd.n2497 vdd.n286 19.3944
R3262 vdd.n2492 vdd.n286 19.3944
R3263 vdd.n2492 vdd.n2491 19.3944
R3264 vdd.n2491 vdd.n2490 19.3944
R3265 vdd.n2490 vdd.n2487 19.3944
R3266 vdd.n326 vdd.n321 19.3944
R3267 vdd.n2483 vdd.n2482 19.3944
R3268 vdd.n2482 vdd.n2480 19.3944
R3269 vdd.n2480 vdd.n2477 19.3944
R3270 vdd.n2477 vdd.n2476 19.3944
R3271 vdd.n2476 vdd.n2473 19.3944
R3272 vdd.n2473 vdd.n2472 19.3944
R3273 vdd.n2472 vdd.n2469 19.3944
R3274 vdd.n2469 vdd.n2468 19.3944
R3275 vdd.n2417 vdd.n353 19.3944
R3276 vdd.n2417 vdd.n2414 19.3944
R3277 vdd.n2414 vdd.n2411 19.3944
R3278 vdd.n2411 vdd.n2410 19.3944
R3279 vdd.n2410 vdd.n2407 19.3944
R3280 vdd.n2407 vdd.n2406 19.3944
R3281 vdd.n2406 vdd.n2403 19.3944
R3282 vdd.n2403 vdd.n2402 19.3944
R3283 vdd.n2402 vdd.n2399 19.3944
R3284 vdd.n2399 vdd.n2398 19.3944
R3285 vdd.n2398 vdd.n2395 19.3944
R3286 vdd.n2373 vdd.n365 19.3944
R3287 vdd.n2391 vdd.n2390 19.3944
R3288 vdd.n2390 vdd.n2388 19.3944
R3289 vdd.n2388 vdd.n2385 19.3944
R3290 vdd.n2385 vdd.n2384 19.3944
R3291 vdd.n1017 vdd.n1013 19.0066
R3292 vdd.n1339 vdd.n1289 19.0066
R3293 vdd.n2639 vdd.n178 19.0066
R3294 vdd.n2421 vdd.n353 19.0066
R3295 vdd.n1649 vdd.n679 17.3257
R3296 vdd.n1882 vdd.n523 17.3257
R3297 vdd.n2139 vdd.n1883 17.3257
R3298 vdd.n2345 vdd.n288 17.3257
R3299 vdd.n1084 vdd.n867 14.4382
R3300 vdd.n1092 vdd.n861 14.4382
R3301 vdd.n1092 vdd.n854 14.4382
R3302 vdd.n1100 vdd.n854 14.4382
R3303 vdd.n1100 vdd.n855 14.4382
R3304 vdd.n1108 vdd.n843 14.4382
R3305 vdd.n1116 vdd.n843 14.4382
R3306 vdd.n1124 vdd.n837 14.4382
R3307 vdd.n1132 vdd.n830 14.4382
R3308 vdd.n1132 vdd.n831 14.4382
R3309 vdd.n1140 vdd.n819 14.4382
R3310 vdd.n1149 vdd.n819 14.4382
R3311 vdd.n1157 vdd.n813 14.4382
R3312 vdd.n1165 vdd.n776 14.4382
R3313 vdd.n1165 vdd.n777 14.4382
R3314 vdd.n1173 vdd.n765 14.4382
R3315 vdd.n1181 vdd.n765 14.4382
R3316 vdd.n1189 vdd.n759 14.4382
R3317 vdd.n1197 vdd.n752 14.4382
R3318 vdd.n1197 vdd.n753 14.4382
R3319 vdd.n1205 vdd.n741 14.4382
R3320 vdd.n1213 vdd.n741 14.4382
R3321 vdd.n1213 vdd.n734 14.4382
R3322 vdd.n1222 vdd.n734 14.4382
R3323 vdd.n1412 vdd.n725 14.4382
R3324 vdd.n2503 vdd.n282 14.4382
R3325 vdd.n2511 vdd.n276 14.4382
R3326 vdd.n2511 vdd.n269 14.4382
R3327 vdd.n2519 vdd.n269 14.4382
R3328 vdd.n2519 vdd.n270 14.4382
R3329 vdd.n2527 vdd.n258 14.4382
R3330 vdd.n2535 vdd.n258 14.4382
R3331 vdd.n2543 vdd.n252 14.4382
R3332 vdd.n2551 vdd.n245 14.4382
R3333 vdd.n2551 vdd.n246 14.4382
R3334 vdd.n2559 vdd.n234 14.4382
R3335 vdd.n2567 vdd.n234 14.4382
R3336 vdd.n2745 vdd.n64 14.4382
R3337 vdd.n2744 vdd.n2743 14.4382
R3338 vdd.n2743 vdd.n68 14.4382
R3339 vdd.n2737 vdd.n2736 14.4382
R3340 vdd.n2736 vdd.n2735 14.4382
R3341 vdd.n2729 vdd.n85 14.4382
R3342 vdd.n2728 vdd.n2727 14.4382
R3343 vdd.n2727 vdd.n89 14.4382
R3344 vdd.n2721 vdd.n2720 14.4382
R3345 vdd.n2720 vdd.n2719 14.4382
R3346 vdd.n2719 vdd.n100 14.4382
R3347 vdd.n2713 vdd.n100 14.4382
R3348 vdd.n2712 vdd.n2711 14.4382
R3349 vdd.n28 vdd.n27 14.3131
R3350 vdd.n1050 vdd.n1046 12.9944
R3351 vdd.n1051 vdd.n1050 12.9944
R3352 vdd.n1376 vdd.n1254 12.9944
R3353 vdd.n1376 vdd.n1251 12.9944
R3354 vdd.n2676 vdd.n143 12.9944
R3355 vdd.n2676 vdd.n140 12.9944
R3356 vdd.n2465 vdd.n335 12.9944
R3357 vdd.n2468 vdd.n2465 12.9944
R3358 vdd.n1124 vdd.t129 12.2725
R3359 vdd.t110 vdd.n759 12.2725
R3360 vdd.n2543 vdd.t23 12.2725
R3361 vdd.n85 vdd.t6 12.2725
R3362 vdd.t19 vdd.n813 11.9838
R3363 vdd.n1157 vdd.t120 11.9838
R3364 vdd.t156 vdd.n64 11.9838
R3365 vdd.n2745 vdd.t4 11.9838
R3366 vdd.t186 vdd.n837 11.695
R3367 vdd.n1189 vdd.t116 11.695
R3368 vdd.t9 vdd.n252 11.695
R3369 vdd.n2729 vdd.t25 11.695
R3370 vdd.n1647 vdd.n670 10.6151
R3371 vdd.n1657 vdd.n670 10.6151
R3372 vdd.n1658 vdd.n1657 10.6151
R3373 vdd.n1659 vdd.n1658 10.6151
R3374 vdd.n1659 vdd.n658 10.6151
R3375 vdd.n1670 vdd.n658 10.6151
R3376 vdd.n1671 vdd.n1670 10.6151
R3377 vdd.n1672 vdd.n1671 10.6151
R3378 vdd.n1672 vdd.n646 10.6151
R3379 vdd.n1682 vdd.n646 10.6151
R3380 vdd.n1683 vdd.n1682 10.6151
R3381 vdd.n1684 vdd.n1683 10.6151
R3382 vdd.n1684 vdd.n634 10.6151
R3383 vdd.n1694 vdd.n634 10.6151
R3384 vdd.n1695 vdd.n1694 10.6151
R3385 vdd.n1696 vdd.n1695 10.6151
R3386 vdd.n1696 vdd.n622 10.6151
R3387 vdd.n1706 vdd.n622 10.6151
R3388 vdd.n1707 vdd.n1706 10.6151
R3389 vdd.n1708 vdd.n1707 10.6151
R3390 vdd.n1708 vdd.n611 10.6151
R3391 vdd.n1718 vdd.n611 10.6151
R3392 vdd.n1719 vdd.n1718 10.6151
R3393 vdd.n1720 vdd.n1719 10.6151
R3394 vdd.n1720 vdd.n600 10.6151
R3395 vdd.n1730 vdd.n600 10.6151
R3396 vdd.n1731 vdd.n1730 10.6151
R3397 vdd.n1732 vdd.n1731 10.6151
R3398 vdd.n1732 vdd.n588 10.6151
R3399 vdd.n1742 vdd.n588 10.6151
R3400 vdd.n1743 vdd.n1742 10.6151
R3401 vdd.n1744 vdd.n1743 10.6151
R3402 vdd.n1744 vdd.n576 10.6151
R3403 vdd.n1754 vdd.n576 10.6151
R3404 vdd.n1755 vdd.n1754 10.6151
R3405 vdd.n1757 vdd.n1755 10.6151
R3406 vdd.n1757 vdd.n1756 10.6151
R3407 vdd.n1756 vdd.n562 10.6151
R3408 vdd.n1826 vdd.n562 10.6151
R3409 vdd.n1826 vdd.n1825 10.6151
R3410 vdd.n1824 vdd.n1822 10.6151
R3411 vdd.n1822 vdd.n1819 10.6151
R3412 vdd.n1819 vdd.n1818 10.6151
R3413 vdd.n1818 vdd.n1815 10.6151
R3414 vdd.n1815 vdd.n1814 10.6151
R3415 vdd.n1814 vdd.n1811 10.6151
R3416 vdd.n1811 vdd.n1810 10.6151
R3417 vdd.n1810 vdd.n1807 10.6151
R3418 vdd.n1807 vdd.n1806 10.6151
R3419 vdd.n1806 vdd.n1803 10.6151
R3420 vdd.n1803 vdd.n1802 10.6151
R3421 vdd.n1802 vdd.n1799 10.6151
R3422 vdd.n1799 vdd.n1798 10.6151
R3423 vdd.n1798 vdd.n1795 10.6151
R3424 vdd.n1795 vdd.n1794 10.6151
R3425 vdd.n1794 vdd.n1791 10.6151
R3426 vdd.n1791 vdd.n1790 10.6151
R3427 vdd.n1790 vdd.n1787 10.6151
R3428 vdd.n1787 vdd.n1786 10.6151
R3429 vdd.n1786 vdd.n1783 10.6151
R3430 vdd.n1783 vdd.n1782 10.6151
R3431 vdd.n1782 vdd.n1779 10.6151
R3432 vdd.n1777 vdd.n1774 10.6151
R3433 vdd.n1774 vdd.n1773 10.6151
R3434 vdd.n1595 vdd.n1594 10.6151
R3435 vdd.n1594 vdd.n1592 10.6151
R3436 vdd.n1592 vdd.n1591 10.6151
R3437 vdd.n1591 vdd.n1589 10.6151
R3438 vdd.n1589 vdd.n1588 10.6151
R3439 vdd.n1588 vdd.n1586 10.6151
R3440 vdd.n1586 vdd.n1585 10.6151
R3441 vdd.n1585 vdd.n1583 10.6151
R3442 vdd.n1583 vdd.n1582 10.6151
R3443 vdd.n1582 vdd.n1580 10.6151
R3444 vdd.n1580 vdd.n1579 10.6151
R3445 vdd.n1579 vdd.n1577 10.6151
R3446 vdd.n1577 vdd.n1576 10.6151
R3447 vdd.n1576 vdd.n1574 10.6151
R3448 vdd.n1574 vdd.n1573 10.6151
R3449 vdd.n1573 vdd.n1571 10.6151
R3450 vdd.n1571 vdd.n1570 10.6151
R3451 vdd.n1570 vdd.n1568 10.6151
R3452 vdd.n1568 vdd.n1567 10.6151
R3453 vdd.n1567 vdd.n1565 10.6151
R3454 vdd.n1565 vdd.n1564 10.6151
R3455 vdd.n1564 vdd.n699 10.6151
R3456 vdd.n1533 vdd.n699 10.6151
R3457 vdd.n1534 vdd.n1533 10.6151
R3458 vdd.n1551 vdd.n1534 10.6151
R3459 vdd.n1551 vdd.n1550 10.6151
R3460 vdd.n1550 vdd.n1549 10.6151
R3461 vdd.n1549 vdd.n1547 10.6151
R3462 vdd.n1547 vdd.n1546 10.6151
R3463 vdd.n1546 vdd.n1544 10.6151
R3464 vdd.n1544 vdd.n1543 10.6151
R3465 vdd.n1543 vdd.n1541 10.6151
R3466 vdd.n1541 vdd.n1540 10.6151
R3467 vdd.n1540 vdd.n1538 10.6151
R3468 vdd.n1538 vdd.n1537 10.6151
R3469 vdd.n1537 vdd.n1535 10.6151
R3470 vdd.n1535 vdd.n565 10.6151
R3471 vdd.n1768 vdd.n565 10.6151
R3472 vdd.n1769 vdd.n1768 10.6151
R3473 vdd.n1770 vdd.n1769 10.6151
R3474 vdd.n1646 vdd.n1645 10.6151
R3475 vdd.n1645 vdd.n683 10.6151
R3476 vdd.n1640 vdd.n683 10.6151
R3477 vdd.n1640 vdd.n1639 10.6151
R3478 vdd.n1639 vdd.n685 10.6151
R3479 vdd.n1634 vdd.n685 10.6151
R3480 vdd.n1634 vdd.n1633 10.6151
R3481 vdd.n1633 vdd.n1632 10.6151
R3482 vdd.n1632 vdd.n687 10.6151
R3483 vdd.n1626 vdd.n687 10.6151
R3484 vdd.n1626 vdd.n1625 10.6151
R3485 vdd.n1625 vdd.n1624 10.6151
R3486 vdd.n1620 vdd.n1619 10.6151
R3487 vdd.n1619 vdd.n691 10.6151
R3488 vdd.n1614 vdd.n691 10.6151
R3489 vdd.n1614 vdd.n1613 10.6151
R3490 vdd.n1613 vdd.n1612 10.6151
R3491 vdd.n1612 vdd.n693 10.6151
R3492 vdd.n1606 vdd.n693 10.6151
R3493 vdd.n1606 vdd.n1605 10.6151
R3494 vdd.n1605 vdd.n1604 10.6151
R3495 vdd.n1600 vdd.n1599 10.6151
R3496 vdd.n1599 vdd.n1596 10.6151
R3497 vdd.n1971 vdd.n1969 10.6151
R3498 vdd.n1972 vdd.n1971 10.6151
R3499 vdd.n1974 vdd.n1972 10.6151
R3500 vdd.n1975 vdd.n1974 10.6151
R3501 vdd.n1977 vdd.n1975 10.6151
R3502 vdd.n1978 vdd.n1977 10.6151
R3503 vdd.n1980 vdd.n1978 10.6151
R3504 vdd.n1981 vdd.n1980 10.6151
R3505 vdd.n1983 vdd.n1981 10.6151
R3506 vdd.n1984 vdd.n1983 10.6151
R3507 vdd.n1986 vdd.n1984 10.6151
R3508 vdd.n1987 vdd.n1986 10.6151
R3509 vdd.n1989 vdd.n1987 10.6151
R3510 vdd.n1990 vdd.n1989 10.6151
R3511 vdd.n2058 vdd.n1990 10.6151
R3512 vdd.n2058 vdd.n2057 10.6151
R3513 vdd.n2057 vdd.n2056 10.6151
R3514 vdd.n2056 vdd.n2054 10.6151
R3515 vdd.n2054 vdd.n2053 10.6151
R3516 vdd.n2053 vdd.n2016 10.6151
R3517 vdd.n2016 vdd.n2015 10.6151
R3518 vdd.n2015 vdd.n2013 10.6151
R3519 vdd.n2013 vdd.n2012 10.6151
R3520 vdd.n2012 vdd.n2010 10.6151
R3521 vdd.n2010 vdd.n2009 10.6151
R3522 vdd.n2009 vdd.n2007 10.6151
R3523 vdd.n2007 vdd.n2006 10.6151
R3524 vdd.n2006 vdd.n2004 10.6151
R3525 vdd.n2004 vdd.n2003 10.6151
R3526 vdd.n2003 vdd.n2001 10.6151
R3527 vdd.n2001 vdd.n2000 10.6151
R3528 vdd.n2000 vdd.n1998 10.6151
R3529 vdd.n1998 vdd.n1997 10.6151
R3530 vdd.n1997 vdd.n1995 10.6151
R3531 vdd.n1995 vdd.n1994 10.6151
R3532 vdd.n1994 vdd.n1992 10.6151
R3533 vdd.n1992 vdd.n1991 10.6151
R3534 vdd.n1991 vdd.n408 10.6151
R3535 vdd.n2293 vdd.n408 10.6151
R3536 vdd.n2294 vdd.n2293 10.6151
R3537 vdd.n1920 vdd.n521 10.6151
R3538 vdd.n1921 vdd.n1920 10.6151
R3539 vdd.n1922 vdd.n1921 10.6151
R3540 vdd.n1922 vdd.n1916 10.6151
R3541 vdd.n1928 vdd.n1916 10.6151
R3542 vdd.n1929 vdd.n1928 10.6151
R3543 vdd.n1930 vdd.n1929 10.6151
R3544 vdd.n1930 vdd.n1914 10.6151
R3545 vdd.n1936 vdd.n1914 10.6151
R3546 vdd.n1937 vdd.n1936 10.6151
R3547 vdd.n1938 vdd.n1937 10.6151
R3548 vdd.n1938 vdd.n1912 10.6151
R3549 vdd.n1944 vdd.n1912 10.6151
R3550 vdd.n1945 vdd.n1944 10.6151
R3551 vdd.n1946 vdd.n1945 10.6151
R3552 vdd.n1946 vdd.n1910 10.6151
R3553 vdd.n1952 vdd.n1910 10.6151
R3554 vdd.n1953 vdd.n1952 10.6151
R3555 vdd.n1954 vdd.n1953 10.6151
R3556 vdd.n1954 vdd.n1908 10.6151
R3557 vdd.n1960 vdd.n1908 10.6151
R3558 vdd.n1961 vdd.n1960 10.6151
R3559 vdd.n1963 vdd.n1904 10.6151
R3560 vdd.n1968 vdd.n1904 10.6151
R3561 vdd.n2142 vdd.n2141 10.6151
R3562 vdd.n2143 vdd.n2142 10.6151
R3563 vdd.n2143 vdd.n509 10.6151
R3564 vdd.n2153 vdd.n509 10.6151
R3565 vdd.n2154 vdd.n2153 10.6151
R3566 vdd.n2155 vdd.n2154 10.6151
R3567 vdd.n2155 vdd.n497 10.6151
R3568 vdd.n2165 vdd.n497 10.6151
R3569 vdd.n2166 vdd.n2165 10.6151
R3570 vdd.n2167 vdd.n2166 10.6151
R3571 vdd.n2167 vdd.n486 10.6151
R3572 vdd.n2177 vdd.n486 10.6151
R3573 vdd.n2178 vdd.n2177 10.6151
R3574 vdd.n2179 vdd.n2178 10.6151
R3575 vdd.n2179 vdd.n475 10.6151
R3576 vdd.n2189 vdd.n475 10.6151
R3577 vdd.n2190 vdd.n2189 10.6151
R3578 vdd.n2191 vdd.n2190 10.6151
R3579 vdd.n2191 vdd.n463 10.6151
R3580 vdd.n2201 vdd.n463 10.6151
R3581 vdd.n2202 vdd.n2201 10.6151
R3582 vdd.n2203 vdd.n2202 10.6151
R3583 vdd.n2203 vdd.n451 10.6151
R3584 vdd.n2213 vdd.n451 10.6151
R3585 vdd.n2214 vdd.n2213 10.6151
R3586 vdd.n2215 vdd.n2214 10.6151
R3587 vdd.n2215 vdd.n439 10.6151
R3588 vdd.n2225 vdd.n439 10.6151
R3589 vdd.n2226 vdd.n2225 10.6151
R3590 vdd.n2227 vdd.n2226 10.6151
R3591 vdd.n2227 vdd.n428 10.6151
R3592 vdd.n2237 vdd.n428 10.6151
R3593 vdd.n2238 vdd.n2237 10.6151
R3594 vdd.n2239 vdd.n2238 10.6151
R3595 vdd.n2239 vdd.n414 10.6151
R3596 vdd.n2286 vdd.n414 10.6151
R3597 vdd.n2287 vdd.n2286 10.6151
R3598 vdd.n2288 vdd.n2287 10.6151
R3599 vdd.n2288 vdd.n388 10.6151
R3600 vdd.n2343 vdd.n388 10.6151
R3601 vdd.n2342 vdd.n2341 10.6151
R3602 vdd.n2341 vdd.n389 10.6151
R3603 vdd.n2336 vdd.n389 10.6151
R3604 vdd.n2336 vdd.n2335 10.6151
R3605 vdd.n2335 vdd.n2334 10.6151
R3606 vdd.n2334 vdd.n392 10.6151
R3607 vdd.n2329 vdd.n392 10.6151
R3608 vdd.n2329 vdd.n2328 10.6151
R3609 vdd.n2328 vdd.n2327 10.6151
R3610 vdd.n2327 vdd.n395 10.6151
R3611 vdd.n2322 vdd.n395 10.6151
R3612 vdd.n2322 vdd.n2321 10.6151
R3613 vdd.n2317 vdd.n2316 10.6151
R3614 vdd.n2316 vdd.n2315 10.6151
R3615 vdd.n2315 vdd.n398 10.6151
R3616 vdd.n2310 vdd.n398 10.6151
R3617 vdd.n2310 vdd.n2309 10.6151
R3618 vdd.n2309 vdd.n2308 10.6151
R3619 vdd.n2308 vdd.n401 10.6151
R3620 vdd.n2303 vdd.n401 10.6151
R3621 vdd.n2303 vdd.n2302 10.6151
R3622 vdd.n2300 vdd.n406 10.6151
R3623 vdd.n2295 vdd.n406 10.6151
R3624 vdd.n2276 vdd.n2246 10.6151
R3625 vdd.n2247 vdd.n2246 10.6151
R3626 vdd.n2269 vdd.n2247 10.6151
R3627 vdd.n2269 vdd.n2268 10.6151
R3628 vdd.n2268 vdd.n2267 10.6151
R3629 vdd.n2267 vdd.n2249 10.6151
R3630 vdd.n2262 vdd.n2249 10.6151
R3631 vdd.n2262 vdd.n2261 10.6151
R3632 vdd.n2261 vdd.n2260 10.6151
R3633 vdd.n2260 vdd.n2252 10.6151
R3634 vdd.n2255 vdd.n2252 10.6151
R3635 vdd.n2255 vdd.n367 10.6151
R3636 vdd.n2369 vdd.n368 10.6151
R3637 vdd.n2364 vdd.n368 10.6151
R3638 vdd.n2364 vdd.n2363 10.6151
R3639 vdd.n2363 vdd.n2362 10.6151
R3640 vdd.n2362 vdd.n371 10.6151
R3641 vdd.n2357 vdd.n371 10.6151
R3642 vdd.n2357 vdd.n2356 10.6151
R3643 vdd.n2356 vdd.n2355 10.6151
R3644 vdd.n2355 vdd.n374 10.6151
R3645 vdd.n2350 vdd.n2349 10.6151
R3646 vdd.n2349 vdd.n2348 10.6151
R3647 vdd.n2084 vdd.n2083 10.6151
R3648 vdd.n2083 vdd.n2081 10.6151
R3649 vdd.n2081 vdd.n2080 10.6151
R3650 vdd.n2080 vdd.n2078 10.6151
R3651 vdd.n2078 vdd.n2077 10.6151
R3652 vdd.n2077 vdd.n2075 10.6151
R3653 vdd.n2075 vdd.n2074 10.6151
R3654 vdd.n2074 vdd.n2072 10.6151
R3655 vdd.n2072 vdd.n2071 10.6151
R3656 vdd.n2071 vdd.n2069 10.6151
R3657 vdd.n2069 vdd.n2068 10.6151
R3658 vdd.n2068 vdd.n2066 10.6151
R3659 vdd.n2066 vdd.n2065 10.6151
R3660 vdd.n2065 vdd.n2063 10.6151
R3661 vdd.n2063 vdd.n2062 10.6151
R3662 vdd.n2062 vdd.n1903 10.6151
R3663 vdd.n2018 vdd.n1903 10.6151
R3664 vdd.n2019 vdd.n2018 10.6151
R3665 vdd.n2049 vdd.n2019 10.6151
R3666 vdd.n2049 vdd.n2048 10.6151
R3667 vdd.n2048 vdd.n2047 10.6151
R3668 vdd.n2047 vdd.n2045 10.6151
R3669 vdd.n2045 vdd.n2044 10.6151
R3670 vdd.n2044 vdd.n2042 10.6151
R3671 vdd.n2042 vdd.n2041 10.6151
R3672 vdd.n2041 vdd.n2039 10.6151
R3673 vdd.n2039 vdd.n2038 10.6151
R3674 vdd.n2038 vdd.n2036 10.6151
R3675 vdd.n2036 vdd.n2035 10.6151
R3676 vdd.n2035 vdd.n2033 10.6151
R3677 vdd.n2033 vdd.n2032 10.6151
R3678 vdd.n2032 vdd.n2030 10.6151
R3679 vdd.n2030 vdd.n2029 10.6151
R3680 vdd.n2029 vdd.n2027 10.6151
R3681 vdd.n2027 vdd.n2026 10.6151
R3682 vdd.n2026 vdd.n2024 10.6151
R3683 vdd.n2024 vdd.n2023 10.6151
R3684 vdd.n2023 vdd.n2021 10.6151
R3685 vdd.n2021 vdd.n2020 10.6151
R3686 vdd.n2020 vdd.n380 10.6151
R3687 vdd.n2136 vdd.n2135 10.6151
R3688 vdd.n2135 vdd.n1888 10.6151
R3689 vdd.n2129 vdd.n1888 10.6151
R3690 vdd.n2129 vdd.n2128 10.6151
R3691 vdd.n2128 vdd.n2127 10.6151
R3692 vdd.n2127 vdd.n1890 10.6151
R3693 vdd.n2121 vdd.n1890 10.6151
R3694 vdd.n2121 vdd.n2120 10.6151
R3695 vdd.n2120 vdd.n2119 10.6151
R3696 vdd.n2119 vdd.n1892 10.6151
R3697 vdd.n2113 vdd.n1892 10.6151
R3698 vdd.n2113 vdd.n2112 10.6151
R3699 vdd.n2112 vdd.n2111 10.6151
R3700 vdd.n2111 vdd.n1894 10.6151
R3701 vdd.n2105 vdd.n1894 10.6151
R3702 vdd.n2105 vdd.n2104 10.6151
R3703 vdd.n2104 vdd.n2103 10.6151
R3704 vdd.n2103 vdd.n1896 10.6151
R3705 vdd.n2097 vdd.n1896 10.6151
R3706 vdd.n2097 vdd.n2096 10.6151
R3707 vdd.n2096 vdd.n2095 10.6151
R3708 vdd.n2095 vdd.n1898 10.6151
R3709 vdd.n2089 vdd.n2088 10.6151
R3710 vdd.n2088 vdd.n2087 10.6151
R3711 vdd.n2137 vdd.n515 10.6151
R3712 vdd.n2147 vdd.n515 10.6151
R3713 vdd.n2148 vdd.n2147 10.6151
R3714 vdd.n2149 vdd.n2148 10.6151
R3715 vdd.n2149 vdd.n504 10.6151
R3716 vdd.n2159 vdd.n504 10.6151
R3717 vdd.n2160 vdd.n2159 10.6151
R3718 vdd.n2161 vdd.n2160 10.6151
R3719 vdd.n2161 vdd.n492 10.6151
R3720 vdd.n2171 vdd.n492 10.6151
R3721 vdd.n2172 vdd.n2171 10.6151
R3722 vdd.n2173 vdd.n2172 10.6151
R3723 vdd.n2173 vdd.n480 10.6151
R3724 vdd.n2183 vdd.n480 10.6151
R3725 vdd.n2184 vdd.n2183 10.6151
R3726 vdd.n2185 vdd.n2184 10.6151
R3727 vdd.n2185 vdd.n469 10.6151
R3728 vdd.n2195 vdd.n469 10.6151
R3729 vdd.n2196 vdd.n2195 10.6151
R3730 vdd.n2197 vdd.n2196 10.6151
R3731 vdd.n2197 vdd.n457 10.6151
R3732 vdd.n2207 vdd.n457 10.6151
R3733 vdd.n2208 vdd.n2207 10.6151
R3734 vdd.n2209 vdd.n2208 10.6151
R3735 vdd.n2209 vdd.n445 10.6151
R3736 vdd.n2219 vdd.n445 10.6151
R3737 vdd.n2220 vdd.n2219 10.6151
R3738 vdd.n2221 vdd.n2220 10.6151
R3739 vdd.n2221 vdd.n434 10.6151
R3740 vdd.n2231 vdd.n434 10.6151
R3741 vdd.n2232 vdd.n2231 10.6151
R3742 vdd.n2233 vdd.n2232 10.6151
R3743 vdd.n2233 vdd.n422 10.6151
R3744 vdd.n2243 vdd.n422 10.6151
R3745 vdd.n2282 vdd.n2245 10.6151
R3746 vdd.n2282 vdd.n2281 10.6151
R3747 vdd.n2281 vdd.n2280 10.6151
R3748 vdd.n2280 vdd.n2279 10.6151
R3749 vdd.n2279 vdd.n2277 10.6151
R3750 vdd.n1652 vdd.n1651 10.6151
R3751 vdd.n1653 vdd.n1652 10.6151
R3752 vdd.n1653 vdd.n664 10.6151
R3753 vdd.n1663 vdd.n664 10.6151
R3754 vdd.n1664 vdd.n1663 10.6151
R3755 vdd.n1666 vdd.n652 10.6151
R3756 vdd.n1676 vdd.n652 10.6151
R3757 vdd.n1677 vdd.n1676 10.6151
R3758 vdd.n1678 vdd.n1677 10.6151
R3759 vdd.n1678 vdd.n640 10.6151
R3760 vdd.n1688 vdd.n640 10.6151
R3761 vdd.n1689 vdd.n1688 10.6151
R3762 vdd.n1690 vdd.n1689 10.6151
R3763 vdd.n1690 vdd.n628 10.6151
R3764 vdd.n1700 vdd.n628 10.6151
R3765 vdd.n1701 vdd.n1700 10.6151
R3766 vdd.n1702 vdd.n1701 10.6151
R3767 vdd.n1702 vdd.n616 10.6151
R3768 vdd.n1712 vdd.n616 10.6151
R3769 vdd.n1713 vdd.n1712 10.6151
R3770 vdd.n1714 vdd.n1713 10.6151
R3771 vdd.n1714 vdd.n605 10.6151
R3772 vdd.n1724 vdd.n605 10.6151
R3773 vdd.n1725 vdd.n1724 10.6151
R3774 vdd.n1726 vdd.n1725 10.6151
R3775 vdd.n1726 vdd.n593 10.6151
R3776 vdd.n1736 vdd.n593 10.6151
R3777 vdd.n1737 vdd.n1736 10.6151
R3778 vdd.n1738 vdd.n1737 10.6151
R3779 vdd.n1738 vdd.n582 10.6151
R3780 vdd.n1748 vdd.n582 10.6151
R3781 vdd.n1749 vdd.n1748 10.6151
R3782 vdd.n1750 vdd.n1749 10.6151
R3783 vdd.n1750 vdd.n569 10.6151
R3784 vdd.n1761 vdd.n569 10.6151
R3785 vdd.n1762 vdd.n1761 10.6151
R3786 vdd.n1764 vdd.n1762 10.6151
R3787 vdd.n1764 vdd.n1763 10.6151
R3788 vdd.n1763 vdd.n552 10.6151
R3789 vdd.n1880 vdd.n1879 10.6151
R3790 vdd.n1879 vdd.n1878 10.6151
R3791 vdd.n1878 vdd.n1875 10.6151
R3792 vdd.n1875 vdd.n1874 10.6151
R3793 vdd.n1874 vdd.n1871 10.6151
R3794 vdd.n1871 vdd.n1870 10.6151
R3795 vdd.n1870 vdd.n1867 10.6151
R3796 vdd.n1867 vdd.n1866 10.6151
R3797 vdd.n1866 vdd.n1863 10.6151
R3798 vdd.n1863 vdd.n1862 10.6151
R3799 vdd.n1862 vdd.n1859 10.6151
R3800 vdd.n1859 vdd.n1858 10.6151
R3801 vdd.n1858 vdd.n1855 10.6151
R3802 vdd.n1855 vdd.n1854 10.6151
R3803 vdd.n1854 vdd.n1851 10.6151
R3804 vdd.n1851 vdd.n1850 10.6151
R3805 vdd.n1850 vdd.n1847 10.6151
R3806 vdd.n1847 vdd.n1846 10.6151
R3807 vdd.n1846 vdd.n1843 10.6151
R3808 vdd.n1843 vdd.n1842 10.6151
R3809 vdd.n1842 vdd.n1839 10.6151
R3810 vdd.n1839 vdd.n1838 10.6151
R3811 vdd.n1835 vdd.n1834 10.6151
R3812 vdd.n1834 vdd.n1832 10.6151
R3813 vdd.n1484 vdd.n1482 10.6151
R3814 vdd.n1485 vdd.n1484 10.6151
R3815 vdd.n1487 vdd.n1485 10.6151
R3816 vdd.n1488 vdd.n1487 10.6151
R3817 vdd.n1490 vdd.n1488 10.6151
R3818 vdd.n1491 vdd.n1490 10.6151
R3819 vdd.n1493 vdd.n1491 10.6151
R3820 vdd.n1494 vdd.n1493 10.6151
R3821 vdd.n1496 vdd.n1494 10.6151
R3822 vdd.n1497 vdd.n1496 10.6151
R3823 vdd.n1499 vdd.n1497 10.6151
R3824 vdd.n1500 vdd.n1499 10.6151
R3825 vdd.n1502 vdd.n1500 10.6151
R3826 vdd.n1503 vdd.n1502 10.6151
R3827 vdd.n1505 vdd.n1503 10.6151
R3828 vdd.n1506 vdd.n1505 10.6151
R3829 vdd.n1508 vdd.n1506 10.6151
R3830 vdd.n1509 vdd.n1508 10.6151
R3831 vdd.n1511 vdd.n1509 10.6151
R3832 vdd.n1512 vdd.n1511 10.6151
R3833 vdd.n1560 vdd.n1512 10.6151
R3834 vdd.n1560 vdd.n1559 10.6151
R3835 vdd.n1559 vdd.n1558 10.6151
R3836 vdd.n1558 vdd.n1556 10.6151
R3837 vdd.n1556 vdd.n1555 10.6151
R3838 vdd.n1555 vdd.n1531 10.6151
R3839 vdd.n1531 vdd.n1530 10.6151
R3840 vdd.n1530 vdd.n1528 10.6151
R3841 vdd.n1528 vdd.n1527 10.6151
R3842 vdd.n1527 vdd.n1525 10.6151
R3843 vdd.n1525 vdd.n1524 10.6151
R3844 vdd.n1524 vdd.n1522 10.6151
R3845 vdd.n1522 vdd.n1521 10.6151
R3846 vdd.n1521 vdd.n1519 10.6151
R3847 vdd.n1519 vdd.n1518 10.6151
R3848 vdd.n1518 vdd.n1516 10.6151
R3849 vdd.n1516 vdd.n1515 10.6151
R3850 vdd.n1515 vdd.n1513 10.6151
R3851 vdd.n1513 vdd.n556 10.6151
R3852 vdd.n1831 vdd.n556 10.6151
R3853 vdd.n1433 vdd.n677 10.6151
R3854 vdd.n1434 vdd.n1433 10.6151
R3855 vdd.n1435 vdd.n1434 10.6151
R3856 vdd.n1435 vdd.n1429 10.6151
R3857 vdd.n1441 vdd.n1429 10.6151
R3858 vdd.n1442 vdd.n1441 10.6151
R3859 vdd.n1443 vdd.n1442 10.6151
R3860 vdd.n1443 vdd.n1427 10.6151
R3861 vdd.n1449 vdd.n1427 10.6151
R3862 vdd.n1450 vdd.n1449 10.6151
R3863 vdd.n1451 vdd.n1450 10.6151
R3864 vdd.n1451 vdd.n1425 10.6151
R3865 vdd.n1458 vdd.n1457 10.6151
R3866 vdd.n1459 vdd.n1458 10.6151
R3867 vdd.n1459 vdd.n706 10.6151
R3868 vdd.n1465 vdd.n706 10.6151
R3869 vdd.n1466 vdd.n1465 10.6151
R3870 vdd.n1467 vdd.n1466 10.6151
R3871 vdd.n1467 vdd.n704 10.6151
R3872 vdd.n1473 vdd.n704 10.6151
R3873 vdd.n1474 vdd.n1473 10.6151
R3874 vdd.n1476 vdd.n700 10.6151
R3875 vdd.n1481 vdd.n700 10.6151
R3876 vdd.n1084 vdd.t43 9.96251
R3877 vdd.t68 vdd.n725 9.96251
R3878 vdd.n2503 vdd.t36 9.96251
R3879 vdd.t28 vdd.n2712 9.96251
R3880 vdd.n1649 vdd.n672 9.81813
R3881 vdd.n1655 vdd.n672 9.81813
R3882 vdd.n1655 vdd.n675 9.81813
R3883 vdd.n1661 vdd.n668 9.81813
R3884 vdd.n1668 vdd.n654 9.81813
R3885 vdd.n1674 vdd.n654 9.81813
R3886 vdd.n1674 vdd.n648 9.81813
R3887 vdd.n1680 vdd.n648 9.81813
R3888 vdd.n1686 vdd.n642 9.81813
R3889 vdd.n1692 vdd.n636 9.81813
R3890 vdd.n1698 vdd.n630 9.81813
R3891 vdd.n1704 vdd.n624 9.81813
R3892 vdd.n1710 vdd.n618 9.81813
R3893 vdd.n1716 vdd.n607 9.81813
R3894 vdd.n1722 vdd.n607 9.81813
R3895 vdd.n1728 vdd.n595 9.81813
R3896 vdd.n1734 vdd.n595 9.81813
R3897 vdd.n1734 vdd.n598 9.81813
R3898 vdd.n1746 vdd.n584 9.81813
R3899 vdd.n1746 vdd.n578 9.81813
R3900 vdd.n1752 vdd.n578 9.81813
R3901 vdd.n1759 vdd.n571 9.81813
R3902 vdd.n1766 vdd.n567 9.81813
R3903 vdd.n1828 vdd.n523 9.81813
R3904 vdd.n2139 vdd.n1886 9.81813
R3905 vdd.n2145 vdd.n519 9.81813
R3906 vdd.n2151 vdd.n513 9.81813
R3907 vdd.n2157 vdd.n499 9.81813
R3908 vdd.n2163 vdd.n499 9.81813
R3909 vdd.n2163 vdd.n502 9.81813
R3910 vdd.n2175 vdd.n488 9.81813
R3911 vdd.n2175 vdd.n482 9.81813
R3912 vdd.n2181 vdd.n482 9.81813
R3913 vdd.n2187 vdd.n471 9.81813
R3914 vdd.n2193 vdd.n471 9.81813
R3915 vdd.n2199 vdd.n467 9.81813
R3916 vdd.n2205 vdd.n461 9.81813
R3917 vdd.n2211 vdd.n455 9.81813
R3918 vdd.n2217 vdd.n449 9.81813
R3919 vdd.n2223 vdd.n443 9.81813
R3920 vdd.n2229 vdd.n430 9.81813
R3921 vdd.n2235 vdd.n430 9.81813
R3922 vdd.n2235 vdd.n424 9.81813
R3923 vdd.n2241 vdd.n424 9.81813
R3924 vdd.n2284 vdd.n416 9.81813
R3925 vdd.n2290 vdd.n410 9.81813
R3926 vdd.n2290 vdd.n383 9.81813
R3927 vdd.n2345 vdd.n383 9.81813
R3928 vdd.n1397 vdd.n689 9.61581
R3929 vdd.n2485 vdd.n323 9.61581
R3930 vdd.n2393 vdd.n2370 9.61581
R3931 vdd.n1424 vdd.n1423 9.61581
R3932 vdd.t172 vdd.n618 9.385
R3933 vdd.n1562 vdd.t144 9.385
R3934 vdd.n2051 vdd.t137 9.385
R3935 vdd.n467 vdd.t21 9.385
R3936 vdd.n1374 vdd.n1254 9.3005
R3937 vdd.n1373 vdd.n1372 9.3005
R3938 vdd.n1259 vdd.n1258 9.3005
R3939 vdd.n1367 vdd.n1262 9.3005
R3940 vdd.n1366 vdd.n1263 9.3005
R3941 vdd.n1365 vdd.n1264 9.3005
R3942 vdd.n1268 vdd.n1265 9.3005
R3943 vdd.n1360 vdd.n1269 9.3005
R3944 vdd.n1359 vdd.n1270 9.3005
R3945 vdd.n1358 vdd.n1271 9.3005
R3946 vdd.n1275 vdd.n1272 9.3005
R3947 vdd.n1353 vdd.n1276 9.3005
R3948 vdd.n1352 vdd.n1277 9.3005
R3949 vdd.n1351 vdd.n1278 9.3005
R3950 vdd.n1282 vdd.n1279 9.3005
R3951 vdd.n1346 vdd.n1283 9.3005
R3952 vdd.n1345 vdd.n1284 9.3005
R3953 vdd.n1344 vdd.n1285 9.3005
R3954 vdd.n1292 vdd.n1286 9.3005
R3955 vdd.n1339 vdd.n1338 9.3005
R3956 vdd.n1337 vdd.n1289 9.3005
R3957 vdd.n1336 vdd.n1335 9.3005
R3958 vdd.n1294 vdd.n1293 9.3005
R3959 vdd.n1330 vdd.n1297 9.3005
R3960 vdd.n1329 vdd.n1298 9.3005
R3961 vdd.n1328 vdd.n1299 9.3005
R3962 vdd.n1303 vdd.n1300 9.3005
R3963 vdd.n1323 vdd.n1304 9.3005
R3964 vdd.n1322 vdd.n1305 9.3005
R3965 vdd.n1321 vdd.n1306 9.3005
R3966 vdd.n1307 vdd.n708 9.3005
R3967 vdd.n1376 vdd.n1375 9.3005
R3968 vdd.n1390 vdd.n1237 9.3005
R3969 vdd.n1389 vdd.n1242 9.3005
R3970 vdd.n1388 vdd.n1243 9.3005
R3971 vdd.n1247 vdd.n1244 9.3005
R3972 vdd.n1383 vdd.n1248 9.3005
R3973 vdd.n1382 vdd.n1249 9.3005
R3974 vdd.n1381 vdd.n1250 9.3005
R3975 vdd.n1257 vdd.n1251 9.3005
R3976 vdd.n1406 vdd.n1227 9.3005
R3977 vdd.n1231 vdd.n1228 9.3005
R3978 vdd.n1401 vdd.n1232 9.3005
R3979 vdd.n1400 vdd.n1233 9.3005
R3980 vdd.n1408 vdd.n1407 9.3005
R3981 vdd.n1160 vdd.n1159 9.3005
R3982 vdd.n1161 vdd.n779 9.3005
R3983 vdd.n1163 vdd.n1162 9.3005
R3984 vdd.n769 vdd.n768 9.3005
R3985 vdd.n1176 vdd.n1175 9.3005
R3986 vdd.n1177 vdd.n767 9.3005
R3987 vdd.n1179 vdd.n1178 9.3005
R3988 vdd.n757 vdd.n756 9.3005
R3989 vdd.n1192 vdd.n1191 9.3005
R3990 vdd.n1193 vdd.n755 9.3005
R3991 vdd.n1195 vdd.n1194 9.3005
R3992 vdd.n745 vdd.n744 9.3005
R3993 vdd.n1208 vdd.n1207 9.3005
R3994 vdd.n1209 vdd.n743 9.3005
R3995 vdd.n1211 vdd.n1210 9.3005
R3996 vdd.n732 vdd.n731 9.3005
R3997 vdd.n1225 vdd.n1224 9.3005
R3998 vdd.n1226 vdd.n730 9.3005
R3999 vdd.n1410 vdd.n1409 9.3005
R4000 vdd.n2421 vdd.n2420 9.3005
R4001 vdd.n2424 vdd.n352 9.3005
R4002 vdd.n2425 vdd.n351 9.3005
R4003 vdd.n2428 vdd.n350 9.3005
R4004 vdd.n2429 vdd.n349 9.3005
R4005 vdd.n2432 vdd.n348 9.3005
R4006 vdd.n2433 vdd.n347 9.3005
R4007 vdd.n2436 vdd.n346 9.3005
R4008 vdd.n2437 vdd.n345 9.3005
R4009 vdd.n2440 vdd.n344 9.3005
R4010 vdd.n2441 vdd.n343 9.3005
R4011 vdd.n2444 vdd.n342 9.3005
R4012 vdd.n2445 vdd.n341 9.3005
R4013 vdd.n2448 vdd.n340 9.3005
R4014 vdd.n2449 vdd.n339 9.3005
R4015 vdd.n2452 vdd.n338 9.3005
R4016 vdd.n2453 vdd.n337 9.3005
R4017 vdd.n2456 vdd.n336 9.3005
R4018 vdd.n2460 vdd.n2459 9.3005
R4019 vdd.n2461 vdd.n335 9.3005
R4020 vdd.n2465 vdd.n2462 9.3005
R4021 vdd.n2468 vdd.n334 9.3005
R4022 vdd.n2469 vdd.n333 9.3005
R4023 vdd.n2472 vdd.n332 9.3005
R4024 vdd.n2473 vdd.n331 9.3005
R4025 vdd.n2476 vdd.n330 9.3005
R4026 vdd.n2477 vdd.n329 9.3005
R4027 vdd.n2480 vdd.n328 9.3005
R4028 vdd.n2482 vdd.n322 9.3005
R4029 vdd.n2490 vdd.n320 9.3005
R4030 vdd.n2491 vdd.n319 9.3005
R4031 vdd.n2492 vdd.n318 9.3005
R4032 vdd.n286 vdd.n285 9.3005
R4033 vdd.n2498 vdd.n2497 9.3005
R4034 vdd.n2501 vdd.n2500 9.3005
R4035 vdd.n274 vdd.n273 9.3005
R4036 vdd.n2514 vdd.n2513 9.3005
R4037 vdd.n2515 vdd.n272 9.3005
R4038 vdd.n2517 vdd.n2516 9.3005
R4039 vdd.n262 vdd.n261 9.3005
R4040 vdd.n2530 vdd.n2529 9.3005
R4041 vdd.n2531 vdd.n260 9.3005
R4042 vdd.n2533 vdd.n2532 9.3005
R4043 vdd.n250 vdd.n249 9.3005
R4044 vdd.n2546 vdd.n2545 9.3005
R4045 vdd.n2547 vdd.n248 9.3005
R4046 vdd.n2549 vdd.n2548 9.3005
R4047 vdd.n238 vdd.n237 9.3005
R4048 vdd.n2562 vdd.n2561 9.3005
R4049 vdd.n2563 vdd.n236 9.3005
R4050 vdd.n2565 vdd.n2564 9.3005
R4051 vdd.n60 vdd.n58 9.3005
R4052 vdd.n2499 vdd.n284 9.3005
R4053 vdd.n2748 vdd.n2747 9.3005
R4054 vdd.n61 vdd.n59 9.3005
R4055 vdd.n2741 vdd.n70 9.3005
R4056 vdd.n2740 vdd.n71 9.3005
R4057 vdd.n2739 vdd.n72 9.3005
R4058 vdd.n79 vdd.n73 9.3005
R4059 vdd.n2733 vdd.n80 9.3005
R4060 vdd.n2732 vdd.n81 9.3005
R4061 vdd.n2731 vdd.n82 9.3005
R4062 vdd.n91 vdd.n83 9.3005
R4063 vdd.n2725 vdd.n92 9.3005
R4064 vdd.n2724 vdd.n93 9.3005
R4065 vdd.n2723 vdd.n94 9.3005
R4066 vdd.n102 vdd.n95 9.3005
R4067 vdd.n2717 vdd.n103 9.3005
R4068 vdd.n2716 vdd.n104 9.3005
R4069 vdd.n2715 vdd.n105 9.3005
R4070 vdd.n113 vdd.n106 9.3005
R4071 vdd.n2709 vdd.n2708 9.3005
R4072 vdd.n2705 vdd.n114 9.3005
R4073 vdd.n2704 vdd.n117 9.3005
R4074 vdd.n121 vdd.n118 9.3005
R4075 vdd.n122 vdd.n119 9.3005
R4076 vdd.n2697 vdd.n123 9.3005
R4077 vdd.n2696 vdd.n124 9.3005
R4078 vdd.n2695 vdd.n125 9.3005
R4079 vdd.n129 vdd.n126 9.3005
R4080 vdd.n2690 vdd.n130 9.3005
R4081 vdd.n2689 vdd.n131 9.3005
R4082 vdd.n2688 vdd.n132 9.3005
R4083 vdd.n136 vdd.n133 9.3005
R4084 vdd.n2683 vdd.n137 9.3005
R4085 vdd.n2682 vdd.n138 9.3005
R4086 vdd.n2681 vdd.n139 9.3005
R4087 vdd.n146 vdd.n140 9.3005
R4088 vdd.n2676 vdd.n2675 9.3005
R4089 vdd.n2674 vdd.n143 9.3005
R4090 vdd.n2673 vdd.n2672 9.3005
R4091 vdd.n148 vdd.n147 9.3005
R4092 vdd.n2667 vdd.n151 9.3005
R4093 vdd.n2666 vdd.n152 9.3005
R4094 vdd.n2665 vdd.n153 9.3005
R4095 vdd.n157 vdd.n154 9.3005
R4096 vdd.n2660 vdd.n158 9.3005
R4097 vdd.n2659 vdd.n159 9.3005
R4098 vdd.n2658 vdd.n160 9.3005
R4099 vdd.n164 vdd.n161 9.3005
R4100 vdd.n2653 vdd.n165 9.3005
R4101 vdd.n2652 vdd.n166 9.3005
R4102 vdd.n2651 vdd.n167 9.3005
R4103 vdd.n171 vdd.n168 9.3005
R4104 vdd.n2646 vdd.n172 9.3005
R4105 vdd.n2645 vdd.n173 9.3005
R4106 vdd.n2644 vdd.n174 9.3005
R4107 vdd.n181 vdd.n175 9.3005
R4108 vdd.n2639 vdd.n2638 9.3005
R4109 vdd.n2637 vdd.n178 9.3005
R4110 vdd.n2636 vdd.n2635 9.3005
R4111 vdd.n183 vdd.n182 9.3005
R4112 vdd.n2630 vdd.n186 9.3005
R4113 vdd.n2629 vdd.n187 9.3005
R4114 vdd.n2628 vdd.n188 9.3005
R4115 vdd.n192 vdd.n189 9.3005
R4116 vdd.n2623 vdd.n193 9.3005
R4117 vdd.n2622 vdd.n194 9.3005
R4118 vdd.n2621 vdd.n195 9.3005
R4119 vdd.n199 vdd.n196 9.3005
R4120 vdd.n2616 vdd.n200 9.3005
R4121 vdd.n2615 vdd.n201 9.3005
R4122 vdd.n2614 vdd.n202 9.3005
R4123 vdd.n206 vdd.n203 9.3005
R4124 vdd.n2609 vdd.n207 9.3005
R4125 vdd.n2608 vdd.n208 9.3005
R4126 vdd.n2607 vdd.n209 9.3005
R4127 vdd.n215 vdd.n210 9.3005
R4128 vdd.n2602 vdd.n2601 9.3005
R4129 vdd.n2707 vdd.n2706 9.3005
R4130 vdd.n2506 vdd.n2505 9.3005
R4131 vdd.n2507 vdd.n278 9.3005
R4132 vdd.n2509 vdd.n2508 9.3005
R4133 vdd.n267 vdd.n266 9.3005
R4134 vdd.n2522 vdd.n2521 9.3005
R4135 vdd.n2523 vdd.n265 9.3005
R4136 vdd.n2525 vdd.n2524 9.3005
R4137 vdd.n256 vdd.n255 9.3005
R4138 vdd.n2538 vdd.n2537 9.3005
R4139 vdd.n2539 vdd.n254 9.3005
R4140 vdd.n2541 vdd.n2540 9.3005
R4141 vdd.n243 vdd.n242 9.3005
R4142 vdd.n2554 vdd.n2553 9.3005
R4143 vdd.n2555 vdd.n241 9.3005
R4144 vdd.n2557 vdd.n2556 9.3005
R4145 vdd.n231 vdd.n230 9.3005
R4146 vdd.n2570 vdd.n2569 9.3005
R4147 vdd.n2571 vdd.n229 9.3005
R4148 vdd.n2573 vdd.n2572 9.3005
R4149 vdd.n2574 vdd.n228 9.3005
R4150 vdd.n2576 vdd.n2575 9.3005
R4151 vdd.n2577 vdd.n227 9.3005
R4152 vdd.n2579 vdd.n2578 9.3005
R4153 vdd.n2580 vdd.n225 9.3005
R4154 vdd.n2582 vdd.n2581 9.3005
R4155 vdd.n2583 vdd.n224 9.3005
R4156 vdd.n2585 vdd.n2584 9.3005
R4157 vdd.n2586 vdd.n222 9.3005
R4158 vdd.n2588 vdd.n2587 9.3005
R4159 vdd.n2589 vdd.n221 9.3005
R4160 vdd.n2591 vdd.n2590 9.3005
R4161 vdd.n2592 vdd.n219 9.3005
R4162 vdd.n2594 vdd.n2593 9.3005
R4163 vdd.n2595 vdd.n218 9.3005
R4164 vdd.n2597 vdd.n2596 9.3005
R4165 vdd.n2598 vdd.n216 9.3005
R4166 vdd.n2600 vdd.n2599 9.3005
R4167 vdd.n280 vdd.n279 9.3005
R4168 vdd.n2379 vdd.n2378 9.3005
R4169 vdd.n2384 vdd.n2377 9.3005
R4170 vdd.n2385 vdd.n2376 9.3005
R4171 vdd.n2388 vdd.n2375 9.3005
R4172 vdd.n2390 vdd.n366 9.3005
R4173 vdd.n2398 vdd.n364 9.3005
R4174 vdd.n2399 vdd.n363 9.3005
R4175 vdd.n2402 vdd.n362 9.3005
R4176 vdd.n2403 vdd.n361 9.3005
R4177 vdd.n2406 vdd.n360 9.3005
R4178 vdd.n2407 vdd.n359 9.3005
R4179 vdd.n2410 vdd.n358 9.3005
R4180 vdd.n2411 vdd.n357 9.3005
R4181 vdd.n2414 vdd.n356 9.3005
R4182 vdd.n2418 vdd.n2417 9.3005
R4183 vdd.n2419 vdd.n353 9.3005
R4184 vdd.n1422 vdd.n1421 9.3005
R4185 vdd.n1420 vdd.n711 9.3005
R4186 vdd.n1419 vdd.n1418 9.3005
R4187 vdd.n1417 vdd.n716 9.3005
R4188 vdd.n1416 vdd.n1415 9.3005
R4189 vdd.n1087 vdd.n1086 9.3005
R4190 vdd.n1088 vdd.n863 9.3005
R4191 vdd.n1090 vdd.n1089 9.3005
R4192 vdd.n852 vdd.n851 9.3005
R4193 vdd.n1103 vdd.n1102 9.3005
R4194 vdd.n1104 vdd.n850 9.3005
R4195 vdd.n1106 vdd.n1105 9.3005
R4196 vdd.n841 vdd.n840 9.3005
R4197 vdd.n1119 vdd.n1118 9.3005
R4198 vdd.n1120 vdd.n839 9.3005
R4199 vdd.n1122 vdd.n1121 9.3005
R4200 vdd.n828 vdd.n827 9.3005
R4201 vdd.n1135 vdd.n1134 9.3005
R4202 vdd.n1136 vdd.n826 9.3005
R4203 vdd.n1138 vdd.n1137 9.3005
R4204 vdd.n817 vdd.n816 9.3005
R4205 vdd.n1152 vdd.n1151 9.3005
R4206 vdd.n1153 vdd.n815 9.3005
R4207 vdd.n1155 vdd.n1154 9.3005
R4208 vdd.n774 vdd.n773 9.3005
R4209 vdd.n1168 vdd.n1167 9.3005
R4210 vdd.n1169 vdd.n772 9.3005
R4211 vdd.n1171 vdd.n1170 9.3005
R4212 vdd.n763 vdd.n762 9.3005
R4213 vdd.n1184 vdd.n1183 9.3005
R4214 vdd.n1185 vdd.n761 9.3005
R4215 vdd.n1187 vdd.n1186 9.3005
R4216 vdd.n750 vdd.n749 9.3005
R4217 vdd.n1200 vdd.n1199 9.3005
R4218 vdd.n1201 vdd.n748 9.3005
R4219 vdd.n1203 vdd.n1202 9.3005
R4220 vdd.n739 vdd.n738 9.3005
R4221 vdd.n1216 vdd.n1215 9.3005
R4222 vdd.n1217 vdd.n736 9.3005
R4223 vdd.n1220 vdd.n1219 9.3005
R4224 vdd.n1218 vdd.n737 9.3005
R4225 vdd.n724 vdd.n717 9.3005
R4226 vdd.n865 vdd.n864 9.3005
R4227 vdd.n986 vdd.n985 9.3005
R4228 vdd.n987 vdd.n978 9.3005
R4229 vdd.n989 vdd.n988 9.3005
R4230 vdd.n990 vdd.n973 9.3005
R4231 vdd.n992 vdd.n991 9.3005
R4232 vdd.n993 vdd.n972 9.3005
R4233 vdd.n995 vdd.n994 9.3005
R4234 vdd.n996 vdd.n967 9.3005
R4235 vdd.n998 vdd.n997 9.3005
R4236 vdd.n999 vdd.n966 9.3005
R4237 vdd.n1001 vdd.n1000 9.3005
R4238 vdd.n1002 vdd.n961 9.3005
R4239 vdd.n1004 vdd.n1003 9.3005
R4240 vdd.n1005 vdd.n960 9.3005
R4241 vdd.n1007 vdd.n1006 9.3005
R4242 vdd.n1008 vdd.n955 9.3005
R4243 vdd.n1010 vdd.n1009 9.3005
R4244 vdd.n1011 vdd.n954 9.3005
R4245 vdd.n1013 vdd.n1012 9.3005
R4246 vdd.n1017 vdd.n950 9.3005
R4247 vdd.n1019 vdd.n1018 9.3005
R4248 vdd.n1020 vdd.n949 9.3005
R4249 vdd.n1022 vdd.n1021 9.3005
R4250 vdd.n1023 vdd.n944 9.3005
R4251 vdd.n1025 vdd.n1024 9.3005
R4252 vdd.n1026 vdd.n943 9.3005
R4253 vdd.n1028 vdd.n1027 9.3005
R4254 vdd.n1029 vdd.n938 9.3005
R4255 vdd.n1031 vdd.n1030 9.3005
R4256 vdd.n1032 vdd.n937 9.3005
R4257 vdd.n1034 vdd.n1033 9.3005
R4258 vdd.n1035 vdd.n932 9.3005
R4259 vdd.n1037 vdd.n1036 9.3005
R4260 vdd.n1038 vdd.n931 9.3005
R4261 vdd.n1040 vdd.n1039 9.3005
R4262 vdd.n1041 vdd.n926 9.3005
R4263 vdd.n1043 vdd.n1042 9.3005
R4264 vdd.n1044 vdd.n925 9.3005
R4265 vdd.n1046 vdd.n1045 9.3005
R4266 vdd.n1050 vdd.n921 9.3005
R4267 vdd.n1052 vdd.n1051 9.3005
R4268 vdd.n1053 vdd.n920 9.3005
R4269 vdd.n1055 vdd.n1054 9.3005
R4270 vdd.n1056 vdd.n915 9.3005
R4271 vdd.n1058 vdd.n1057 9.3005
R4272 vdd.n1059 vdd.n914 9.3005
R4273 vdd.n1061 vdd.n1060 9.3005
R4274 vdd.n1062 vdd.n909 9.3005
R4275 vdd.n1064 vdd.n1063 9.3005
R4276 vdd.n1065 vdd.n908 9.3005
R4277 vdd.n1067 vdd.n1066 9.3005
R4278 vdd.n1068 vdd.n903 9.3005
R4279 vdd.n1070 vdd.n1069 9.3005
R4280 vdd.n1071 vdd.n902 9.3005
R4281 vdd.n1073 vdd.n1072 9.3005
R4282 vdd.n871 vdd.n870 9.3005
R4283 vdd.n1079 vdd.n1078 9.3005
R4284 vdd.n981 vdd.n979 9.3005
R4285 vdd.n1082 vdd.n1081 9.3005
R4286 vdd.n859 vdd.n858 9.3005
R4287 vdd.n1095 vdd.n1094 9.3005
R4288 vdd.n1096 vdd.n857 9.3005
R4289 vdd.n1098 vdd.n1097 9.3005
R4290 vdd.n847 vdd.n846 9.3005
R4291 vdd.n1111 vdd.n1110 9.3005
R4292 vdd.n1112 vdd.n845 9.3005
R4293 vdd.n1114 vdd.n1113 9.3005
R4294 vdd.n835 vdd.n834 9.3005
R4295 vdd.n1127 vdd.n1126 9.3005
R4296 vdd.n1128 vdd.n833 9.3005
R4297 vdd.n1130 vdd.n1129 9.3005
R4298 vdd.n823 vdd.n822 9.3005
R4299 vdd.n1143 vdd.n1142 9.3005
R4300 vdd.n1144 vdd.n821 9.3005
R4301 vdd.n1147 vdd.n1146 9.3005
R4302 vdd.n1145 vdd.n811 9.3005
R4303 vdd.n1080 vdd.n869 9.3005
R4304 vdd.n1661 vdd.t32 8.80749
R4305 vdd.n1759 vdd.t54 8.80749
R4306 vdd.n2151 vdd.t47 8.80749
R4307 vdd.n2284 vdd.t61 8.80749
R4308 vdd.t154 vdd.n630 8.51874
R4309 vdd.n1553 vdd.t22 8.51874
R4310 vdd.n2060 vdd.t176 8.51874
R4311 vdd.n455 vdd.t155 8.51874
R4312 vdd.n47 vdd.n37 8.43656
R4313 vdd.n798 vdd.n788 8.43656
R4314 vdd.n28 vdd.n14 8.32849
R4315 vdd.n2750 vdd.n2749 8.08725
R4316 vdd.n810 vdd.n809 8.08725
R4317 vdd.n1686 vdd.t135 7.79685
R4318 vdd.n2223 vdd.t124 7.79685
R4319 vdd.n855 vdd.t14 7.65248
R4320 vdd.n1205 vdd.t118 7.65248
R4321 vdd.t3 vdd.n642 7.65248
R4322 vdd.n598 vdd.t173 7.65248
R4323 vdd.t113 vdd.n488 7.65248
R4324 vdd.n443 vdd.t0 7.65248
R4325 vdd.n270 vdd.t103 7.65248
R4326 vdd.n2721 vdd.t147 7.65248
R4327 vdd.n831 vdd.t114 7.36372
R4328 vdd.n1173 vdd.t133 7.36372
R4329 vdd.n246 vdd.t167 7.36372
R4330 vdd.n2737 vdd.t16 7.36372
R4331 vdd.n2245 vdd.n2244 7.18099
R4332 vdd.n1665 vdd.n1664 7.18099
R4333 vdd.n1140 vdd.t114 7.07497
R4334 vdd.n777 vdd.t133 7.07497
R4335 vdd.n2559 vdd.t167 7.07497
R4336 vdd.t16 vdd.n68 7.07497
R4337 vdd.n1018 vdd.n1017 6.98232
R4338 vdd.n1339 vdd.n1286 6.98232
R4339 vdd.n2639 vdd.n175 6.98232
R4340 vdd.n2424 vdd.n2421 6.98232
R4341 vdd.n1698 vdd.t194 6.93059
R4342 vdd.n2211 vdd.t140 6.93059
R4343 vdd.n1108 vdd.t14 6.78621
R4344 vdd.n753 vdd.t118 6.78621
R4345 vdd.n2527 vdd.t103 6.78621
R4346 vdd.t147 vdd.n89 6.78621
R4347 vdd.n668 vdd.t91 6.64184
R4348 vdd.t75 vdd.n416 6.64184
R4349 vdd.n1710 vdd.t142 6.06433
R4350 vdd.n1828 vdd.t181 6.06433
R4351 vdd.n1886 vdd.t214 6.06433
R4352 vdd.n2199 vdd.t177 6.06433
R4353 vdd.n1779 vdd.n1778 5.77611
R4354 vdd.n1604 vdd.n697 5.77611
R4355 vdd.n1962 vdd.n1961 5.77611
R4356 vdd.n2302 vdd.n2301 5.77611
R4357 vdd.n379 vdd.n374 5.77611
R4358 vdd.n1902 vdd.n1898 5.77611
R4359 vdd.n1838 vdd.n555 5.77611
R4360 vdd.n1475 vdd.n1474 5.77611
R4361 vdd.n984 vdd.n981 5.62474
R4362 vdd.n1415 vdd.n720 5.62474
R4363 vdd.n2602 vdd.n214 5.62474
R4364 vdd.n2382 vdd.n2379 5.62474
R4365 vdd.n1740 vdd.t138 5.48682
R4366 vdd.n2169 vdd.t145 5.48682
R4367 vdd.n7 vdd.t141 5.418
R4368 vdd.n7 vdd.t125 5.418
R4369 vdd.n8 vdd.t180 5.418
R4370 vdd.n8 vdd.t178 5.418
R4371 vdd.n10 vdd.t2 5.418
R4372 vdd.n10 vdd.t146 5.418
R4373 vdd.n12 vdd.t175 5.418
R4374 vdd.n12 vdd.t215 5.418
R4375 vdd.n5 vdd.t182 5.418
R4376 vdd.n5 vdd.t166 5.418
R4377 vdd.n3 vdd.t139 5.418
R4378 vdd.n3 vdd.t123 5.418
R4379 vdd.n1 vdd.t143 5.418
R4380 vdd.n1 vdd.t202 5.418
R4381 vdd.n0 vdd.t136 5.418
R4382 vdd.n0 vdd.t195 5.418
R4383 vdd.n1624 vdd.n689 5.30782
R4384 vdd.n1620 vdd.n689 5.30782
R4385 vdd.n2321 vdd.n323 5.30782
R4386 vdd.n2317 vdd.n323 5.30782
R4387 vdd.n2370 vdd.n367 5.30782
R4388 vdd.n2370 vdd.n2369 5.30782
R4389 vdd.n1425 vdd.n1424 5.30782
R4390 vdd.n1457 vdd.n1424 5.30782
R4391 vdd.n1722 vdd.t201 5.19807
R4392 vdd.t122 vdd.n571 5.19807
R4393 vdd.t165 vdd.n1882 5.19807
R4394 vdd.n1883 vdd.t174 5.19807
R4395 vdd.n513 vdd.t1 5.19807
R4396 vdd.n2187 vdd.t179 5.19807
R4397 vdd.n2750 vdd.n57 5.19501
R4398 vdd.n809 vdd.n808 5.19501
R4399 vdd.n1778 vdd.n1777 4.83952
R4400 vdd.n1600 vdd.n697 4.83952
R4401 vdd.n1963 vdd.n1962 4.83952
R4402 vdd.n2301 vdd.n2300 4.83952
R4403 vdd.n2350 vdd.n379 4.83952
R4404 vdd.n2089 vdd.n1902 4.83952
R4405 vdd.n1835 vdd.n555 4.83952
R4406 vdd.n1476 vdd.n1475 4.83952
R4407 vdd.n1316 vdd.n709 4.74817
R4408 vdd.n1312 vdd.n710 4.74817
R4409 vdd.n1399 vdd.n1398 4.74817
R4410 vdd.n1396 vdd.n1238 4.74817
R4411 vdd.n1398 vdd.n1236 4.74817
R4412 vdd.n1396 vdd.n1395 4.74817
R4413 vdd.n2487 vdd.n2486 4.74817
R4414 vdd.n2484 vdd.n2483 4.74817
R4415 vdd.n2484 vdd.n326 4.74817
R4416 vdd.n2486 vdd.n321 4.74817
R4417 vdd.n2394 vdd.n365 4.74817
R4418 vdd.n2392 vdd.n2391 4.74817
R4419 vdd.n2392 vdd.n2373 4.74817
R4420 vdd.n2395 vdd.n2394 4.74817
R4421 vdd.n1309 vdd.n709 4.74817
R4422 vdd.n712 vdd.n710 4.74817
R4423 vdd.n57 vdd.n56 4.7074
R4424 vdd.n47 vdd.n46 4.7074
R4425 vdd.n808 vdd.n807 4.7074
R4426 vdd.n798 vdd.n797 4.7074
R4427 vdd.n54 vdd.t170 4.64407
R4428 vdd.n54 vdd.t26 4.64407
R4429 vdd.n52 vdd.t5 4.64407
R4430 vdd.n52 vdd.t18 4.64407
R4431 vdd.n50 vdd.t183 4.64407
R4432 vdd.n50 vdd.t157 4.64407
R4433 vdd.n48 vdd.t10 4.64407
R4434 vdd.n48 vdd.t160 4.64407
R4435 vdd.n44 vdd.t11 4.64407
R4436 vdd.n44 vdd.t211 4.64407
R4437 vdd.n42 vdd.t206 4.64407
R4438 vdd.n42 vdd.t17 4.64407
R4439 vdd.n40 vdd.t200 4.64407
R4440 vdd.n40 vdd.t191 4.64407
R4441 vdd.n38 vdd.t151 4.64407
R4442 vdd.n38 vdd.t24 4.64407
R4443 vdd.n35 vdd.t7 4.64407
R4444 vdd.n35 vdd.t210 4.64407
R4445 vdd.n33 vdd.t149 4.64407
R4446 vdd.n33 vdd.t152 4.64407
R4447 vdd.n31 vdd.t168 4.64407
R4448 vdd.n31 vdd.t161 4.64407
R4449 vdd.n29 vdd.t159 4.64407
R4450 vdd.n29 vdd.t212 4.64407
R4451 vdd.n799 vdd.t185 4.64407
R4452 vdd.n799 vdd.t204 4.64407
R4453 vdd.n801 vdd.t150 4.64407
R4454 vdd.n801 vdd.t188 4.64407
R4455 vdd.n803 vdd.t189 4.64407
R4456 vdd.n803 vdd.t105 4.64407
R4457 vdd.n805 vdd.t205 4.64407
R4458 vdd.n805 vdd.t130 4.64407
R4459 vdd.n789 vdd.t184 4.64407
R4460 vdd.n789 vdd.t117 4.64407
R4461 vdd.n791 vdd.t121 4.64407
R4462 vdd.n791 vdd.t134 4.64407
R4463 vdd.n793 vdd.t115 4.64407
R4464 vdd.n793 vdd.t169 4.64407
R4465 vdd.n795 vdd.t187 4.64407
R4466 vdd.n795 vdd.t213 4.64407
R4467 vdd.n780 vdd.t111 4.64407
R4468 vdd.n780 vdd.t192 4.64407
R4469 vdd.n782 vdd.t158 4.64407
R4470 vdd.n782 vdd.t171 4.64407
R4471 vdd.n784 vdd.t132 4.64407
R4472 vdd.n784 vdd.t20 4.64407
R4473 vdd.n786 vdd.t193 4.64407
R4474 vdd.n786 vdd.t131 4.64407
R4475 vdd.n1553 vdd.t201 4.62056
R4476 vdd.n1752 vdd.t122 4.62056
R4477 vdd.n2157 vdd.t1 4.62056
R4478 vdd.n2060 vdd.t179 4.62056
R4479 vdd.t43 vdd.n861 4.47618
R4480 vdd.n1222 vdd.t68 4.47618
R4481 vdd.t36 vdd.n276 4.47618
R4482 vdd.n2713 vdd.t28 4.47618
R4483 vdd.t138 vdd.n584 4.33181
R4484 vdd.n502 vdd.t145 4.33181
R4485 vdd.n26 vdd.t127 3.9605
R4486 vdd.n26 vdd.t128 3.9605
R4487 vdd.n23 vdd.t8 3.9605
R4488 vdd.n23 vdd.t108 3.9605
R4489 vdd.n21 vdd.t196 3.9605
R4490 vdd.n21 vdd.t107 3.9605
R4491 vdd.n20 vdd.t12 3.9605
R4492 vdd.n20 vdd.t126 3.9605
R4493 vdd.n15 vdd.t209 3.9605
R4494 vdd.n15 vdd.t13 3.9605
R4495 vdd.n16 vdd.t198 3.9605
R4496 vdd.n16 vdd.t109 3.9605
R4497 vdd.n18 vdd.t197 3.9605
R4498 vdd.n18 vdd.t106 3.9605
R4499 vdd.n25 vdd.t207 3.9605
R4500 vdd.n25 vdd.t208 3.9605
R4501 vdd.n1562 vdd.t142 3.7543
R4502 vdd.n1766 vdd.t181 3.7543
R4503 vdd.n2145 vdd.t214 3.7543
R4504 vdd.n2051 vdd.t177 3.7543
R4505 vdd.n57 vdd.n47 3.72967
R4506 vdd.n808 vdd.n798 3.72967
R4507 vdd.n2244 vdd.n2243 3.43465
R4508 vdd.n1666 vdd.n1665 3.43465
R4509 vdd.n1668 vdd.t91 3.17679
R4510 vdd.n2241 vdd.t75 3.17679
R4511 vdd.t194 vdd.n624 2.88804
R4512 vdd.n461 vdd.t140 2.88804
R4513 vdd.n1116 vdd.t186 2.74366
R4514 vdd.t116 vdd.n752 2.74366
R4515 vdd.n2535 vdd.t9 2.74366
R4516 vdd.t25 vdd.n2728 2.74366
R4517 vdd.n1149 vdd.t19 2.45491
R4518 vdd.t120 vdd.n776 2.45491
R4519 vdd.n2567 vdd.t156 2.45491
R4520 vdd.t4 vdd.n2744 2.45491
R4521 vdd.n1398 vdd.n1397 2.27742
R4522 vdd.n1397 vdd.n1396 2.27742
R4523 vdd.n2485 vdd.n2484 2.27742
R4524 vdd.n2486 vdd.n2485 2.27742
R4525 vdd.n2393 vdd.n2392 2.27742
R4526 vdd.n2394 vdd.n2393 2.27742
R4527 vdd.n1423 vdd.n709 2.27742
R4528 vdd.n1423 vdd.n710 2.27742
R4529 vdd.t129 vdd.n830 2.16615
R4530 vdd.n1181 vdd.t110 2.16615
R4531 vdd.n1680 vdd.t3 2.16615
R4532 vdd.n1740 vdd.t173 2.16615
R4533 vdd.n2169 vdd.t113 2.16615
R4534 vdd.n2229 vdd.t0 2.16615
R4535 vdd.t23 vdd.n245 2.16615
R4536 vdd.n2735 vdd.t6 2.16615
R4537 vdd.t135 vdd.n636 2.02178
R4538 vdd.n449 vdd.t124 2.02178
R4539 vdd.n1692 vdd.t154 1.29989
R4540 vdd.n1728 vdd.t22 1.29989
R4541 vdd.n2181 vdd.t176 1.29989
R4542 vdd.n2217 vdd.t155 1.29989
R4543 vdd.n675 vdd.t32 1.01114
R4544 vdd.t54 vdd.n567 1.01114
R4545 vdd.n519 vdd.t47 1.01114
R4546 vdd.t61 vdd.n410 1.01114
R4547 vdd.n985 vdd.n984 0.970197
R4548 vdd.n720 vdd.n716 0.970197
R4549 vdd.n214 vdd.n210 0.970197
R4550 vdd.n2384 vdd.n2382 0.970197
R4551 vdd.n809 vdd.n28 0.960867
R4552 vdd vdd.n2750 0.953033
R4553 vdd.n4 vdd.n2 0.728948
R4554 vdd.n11 vdd.n9 0.728948
R4555 vdd.n6 vdd.n4 0.573776
R4556 vdd.n13 vdd.n11 0.573776
R4557 vdd.n51 vdd.n49 0.573776
R4558 vdd.n53 vdd.n51 0.573776
R4559 vdd.n55 vdd.n53 0.573776
R4560 vdd.n56 vdd.n55 0.573776
R4561 vdd.n41 vdd.n39 0.573776
R4562 vdd.n43 vdd.n41 0.573776
R4563 vdd.n45 vdd.n43 0.573776
R4564 vdd.n46 vdd.n45 0.573776
R4565 vdd.n32 vdd.n30 0.573776
R4566 vdd.n34 vdd.n32 0.573776
R4567 vdd.n36 vdd.n34 0.573776
R4568 vdd.n37 vdd.n36 0.573776
R4569 vdd.n807 vdd.n806 0.573776
R4570 vdd.n806 vdd.n804 0.573776
R4571 vdd.n804 vdd.n802 0.573776
R4572 vdd.n802 vdd.n800 0.573776
R4573 vdd.n797 vdd.n796 0.573776
R4574 vdd.n796 vdd.n794 0.573776
R4575 vdd.n794 vdd.n792 0.573776
R4576 vdd.n792 vdd.n790 0.573776
R4577 vdd.n788 vdd.n787 0.573776
R4578 vdd.n787 vdd.n785 0.573776
R4579 vdd.n785 vdd.n783 0.573776
R4580 vdd.n783 vdd.n781 0.573776
R4581 vdd.n14 vdd.n6 0.49619
R4582 vdd.n14 vdd.n13 0.49619
R4583 vdd.n1409 vdd.n1408 0.471537
R4584 vdd.n2499 vdd.n2498 0.471537
R4585 vdd.n2708 vdd.n2707 0.471537
R4586 vdd.n2601 vdd.n2600 0.471537
R4587 vdd.n2378 vdd.n279 0.471537
R4588 vdd.n1416 vdd.n717 0.471537
R4589 vdd.n979 vdd.n864 0.471537
R4590 vdd.n1080 vdd.n1079 0.471537
R4591 vdd.n1704 vdd.t172 0.433631
R4592 vdd.n1716 vdd.t144 0.433631
R4593 vdd.n2193 vdd.t137 0.433631
R4594 vdd.n2205 vdd.t21 0.433631
R4595 vdd.n19 vdd.n17 0.387128
R4596 vdd.n24 vdd.n22 0.387128
R4597 vdd.n27 vdd.n19 0.21707
R4598 vdd.n27 vdd.n24 0.21707
R4599 vdd.n1242 vdd.n1237 0.152939
R4600 vdd.n1243 vdd.n1242 0.152939
R4601 vdd.n1247 vdd.n1243 0.152939
R4602 vdd.n1248 vdd.n1247 0.152939
R4603 vdd.n1249 vdd.n1248 0.152939
R4604 vdd.n1250 vdd.n1249 0.152939
R4605 vdd.n1257 vdd.n1250 0.152939
R4606 vdd.n1375 vdd.n1257 0.152939
R4607 vdd.n1375 vdd.n1374 0.152939
R4608 vdd.n1374 vdd.n1373 0.152939
R4609 vdd.n1373 vdd.n1258 0.152939
R4610 vdd.n1262 vdd.n1258 0.152939
R4611 vdd.n1263 vdd.n1262 0.152939
R4612 vdd.n1264 vdd.n1263 0.152939
R4613 vdd.n1268 vdd.n1264 0.152939
R4614 vdd.n1269 vdd.n1268 0.152939
R4615 vdd.n1270 vdd.n1269 0.152939
R4616 vdd.n1271 vdd.n1270 0.152939
R4617 vdd.n1275 vdd.n1271 0.152939
R4618 vdd.n1276 vdd.n1275 0.152939
R4619 vdd.n1277 vdd.n1276 0.152939
R4620 vdd.n1278 vdd.n1277 0.152939
R4621 vdd.n1282 vdd.n1278 0.152939
R4622 vdd.n1283 vdd.n1282 0.152939
R4623 vdd.n1284 vdd.n1283 0.152939
R4624 vdd.n1285 vdd.n1284 0.152939
R4625 vdd.n1292 vdd.n1285 0.152939
R4626 vdd.n1338 vdd.n1292 0.152939
R4627 vdd.n1338 vdd.n1337 0.152939
R4628 vdd.n1337 vdd.n1336 0.152939
R4629 vdd.n1336 vdd.n1293 0.152939
R4630 vdd.n1297 vdd.n1293 0.152939
R4631 vdd.n1298 vdd.n1297 0.152939
R4632 vdd.n1299 vdd.n1298 0.152939
R4633 vdd.n1303 vdd.n1299 0.152939
R4634 vdd.n1304 vdd.n1303 0.152939
R4635 vdd.n1305 vdd.n1304 0.152939
R4636 vdd.n1306 vdd.n1305 0.152939
R4637 vdd.n1306 vdd.n708 0.152939
R4638 vdd.n1408 vdd.n1227 0.152939
R4639 vdd.n1231 vdd.n1227 0.152939
R4640 vdd.n1232 vdd.n1231 0.152939
R4641 vdd.n1233 vdd.n1232 0.152939
R4642 vdd.n1161 vdd.n1160 0.152939
R4643 vdd.n1162 vdd.n1161 0.152939
R4644 vdd.n1162 vdd.n768 0.152939
R4645 vdd.n1176 vdd.n768 0.152939
R4646 vdd.n1177 vdd.n1176 0.152939
R4647 vdd.n1178 vdd.n1177 0.152939
R4648 vdd.n1178 vdd.n756 0.152939
R4649 vdd.n1192 vdd.n756 0.152939
R4650 vdd.n1193 vdd.n1192 0.152939
R4651 vdd.n1194 vdd.n1193 0.152939
R4652 vdd.n1194 vdd.n744 0.152939
R4653 vdd.n1208 vdd.n744 0.152939
R4654 vdd.n1209 vdd.n1208 0.152939
R4655 vdd.n1210 vdd.n1209 0.152939
R4656 vdd.n1210 vdd.n731 0.152939
R4657 vdd.n1225 vdd.n731 0.152939
R4658 vdd.n1226 vdd.n1225 0.152939
R4659 vdd.n1409 vdd.n1226 0.152939
R4660 vdd.n328 vdd.n322 0.152939
R4661 vdd.n329 vdd.n328 0.152939
R4662 vdd.n330 vdd.n329 0.152939
R4663 vdd.n331 vdd.n330 0.152939
R4664 vdd.n332 vdd.n331 0.152939
R4665 vdd.n333 vdd.n332 0.152939
R4666 vdd.n334 vdd.n333 0.152939
R4667 vdd.n2462 vdd.n334 0.152939
R4668 vdd.n2462 vdd.n2461 0.152939
R4669 vdd.n2461 vdd.n2460 0.152939
R4670 vdd.n2460 vdd.n336 0.152939
R4671 vdd.n337 vdd.n336 0.152939
R4672 vdd.n338 vdd.n337 0.152939
R4673 vdd.n339 vdd.n338 0.152939
R4674 vdd.n340 vdd.n339 0.152939
R4675 vdd.n341 vdd.n340 0.152939
R4676 vdd.n342 vdd.n341 0.152939
R4677 vdd.n343 vdd.n342 0.152939
R4678 vdd.n344 vdd.n343 0.152939
R4679 vdd.n345 vdd.n344 0.152939
R4680 vdd.n346 vdd.n345 0.152939
R4681 vdd.n347 vdd.n346 0.152939
R4682 vdd.n348 vdd.n347 0.152939
R4683 vdd.n349 vdd.n348 0.152939
R4684 vdd.n350 vdd.n349 0.152939
R4685 vdd.n351 vdd.n350 0.152939
R4686 vdd.n352 vdd.n351 0.152939
R4687 vdd.n2420 vdd.n352 0.152939
R4688 vdd.n2420 vdd.n2419 0.152939
R4689 vdd.n2419 vdd.n2418 0.152939
R4690 vdd.n2418 vdd.n356 0.152939
R4691 vdd.n357 vdd.n356 0.152939
R4692 vdd.n358 vdd.n357 0.152939
R4693 vdd.n359 vdd.n358 0.152939
R4694 vdd.n360 vdd.n359 0.152939
R4695 vdd.n361 vdd.n360 0.152939
R4696 vdd.n362 vdd.n361 0.152939
R4697 vdd.n363 vdd.n362 0.152939
R4698 vdd.n364 vdd.n363 0.152939
R4699 vdd.n2498 vdd.n285 0.152939
R4700 vdd.n318 vdd.n285 0.152939
R4701 vdd.n319 vdd.n318 0.152939
R4702 vdd.n320 vdd.n319 0.152939
R4703 vdd.n2500 vdd.n2499 0.152939
R4704 vdd.n2500 vdd.n273 0.152939
R4705 vdd.n2514 vdd.n273 0.152939
R4706 vdd.n2515 vdd.n2514 0.152939
R4707 vdd.n2516 vdd.n2515 0.152939
R4708 vdd.n2516 vdd.n261 0.152939
R4709 vdd.n2530 vdd.n261 0.152939
R4710 vdd.n2531 vdd.n2530 0.152939
R4711 vdd.n2532 vdd.n2531 0.152939
R4712 vdd.n2532 vdd.n249 0.152939
R4713 vdd.n2546 vdd.n249 0.152939
R4714 vdd.n2547 vdd.n2546 0.152939
R4715 vdd.n2548 vdd.n2547 0.152939
R4716 vdd.n2548 vdd.n237 0.152939
R4717 vdd.n2562 vdd.n237 0.152939
R4718 vdd.n2563 vdd.n2562 0.152939
R4719 vdd.n2564 vdd.n2563 0.152939
R4720 vdd.n2564 vdd.n58 0.152939
R4721 vdd.n2748 vdd.n59 0.152939
R4722 vdd.n70 vdd.n59 0.152939
R4723 vdd.n71 vdd.n70 0.152939
R4724 vdd.n72 vdd.n71 0.152939
R4725 vdd.n79 vdd.n72 0.152939
R4726 vdd.n80 vdd.n79 0.152939
R4727 vdd.n81 vdd.n80 0.152939
R4728 vdd.n82 vdd.n81 0.152939
R4729 vdd.n91 vdd.n82 0.152939
R4730 vdd.n92 vdd.n91 0.152939
R4731 vdd.n93 vdd.n92 0.152939
R4732 vdd.n94 vdd.n93 0.152939
R4733 vdd.n102 vdd.n94 0.152939
R4734 vdd.n103 vdd.n102 0.152939
R4735 vdd.n104 vdd.n103 0.152939
R4736 vdd.n105 vdd.n104 0.152939
R4737 vdd.n113 vdd.n105 0.152939
R4738 vdd.n2708 vdd.n113 0.152939
R4739 vdd.n2707 vdd.n114 0.152939
R4740 vdd.n117 vdd.n114 0.152939
R4741 vdd.n121 vdd.n117 0.152939
R4742 vdd.n122 vdd.n121 0.152939
R4743 vdd.n123 vdd.n122 0.152939
R4744 vdd.n124 vdd.n123 0.152939
R4745 vdd.n125 vdd.n124 0.152939
R4746 vdd.n129 vdd.n125 0.152939
R4747 vdd.n130 vdd.n129 0.152939
R4748 vdd.n131 vdd.n130 0.152939
R4749 vdd.n132 vdd.n131 0.152939
R4750 vdd.n136 vdd.n132 0.152939
R4751 vdd.n137 vdd.n136 0.152939
R4752 vdd.n138 vdd.n137 0.152939
R4753 vdd.n139 vdd.n138 0.152939
R4754 vdd.n146 vdd.n139 0.152939
R4755 vdd.n2675 vdd.n146 0.152939
R4756 vdd.n2675 vdd.n2674 0.152939
R4757 vdd.n2674 vdd.n2673 0.152939
R4758 vdd.n2673 vdd.n147 0.152939
R4759 vdd.n151 vdd.n147 0.152939
R4760 vdd.n152 vdd.n151 0.152939
R4761 vdd.n153 vdd.n152 0.152939
R4762 vdd.n157 vdd.n153 0.152939
R4763 vdd.n158 vdd.n157 0.152939
R4764 vdd.n159 vdd.n158 0.152939
R4765 vdd.n160 vdd.n159 0.152939
R4766 vdd.n164 vdd.n160 0.152939
R4767 vdd.n165 vdd.n164 0.152939
R4768 vdd.n166 vdd.n165 0.152939
R4769 vdd.n167 vdd.n166 0.152939
R4770 vdd.n171 vdd.n167 0.152939
R4771 vdd.n172 vdd.n171 0.152939
R4772 vdd.n173 vdd.n172 0.152939
R4773 vdd.n174 vdd.n173 0.152939
R4774 vdd.n181 vdd.n174 0.152939
R4775 vdd.n2638 vdd.n181 0.152939
R4776 vdd.n2638 vdd.n2637 0.152939
R4777 vdd.n2637 vdd.n2636 0.152939
R4778 vdd.n2636 vdd.n182 0.152939
R4779 vdd.n186 vdd.n182 0.152939
R4780 vdd.n187 vdd.n186 0.152939
R4781 vdd.n188 vdd.n187 0.152939
R4782 vdd.n192 vdd.n188 0.152939
R4783 vdd.n193 vdd.n192 0.152939
R4784 vdd.n194 vdd.n193 0.152939
R4785 vdd.n195 vdd.n194 0.152939
R4786 vdd.n199 vdd.n195 0.152939
R4787 vdd.n200 vdd.n199 0.152939
R4788 vdd.n201 vdd.n200 0.152939
R4789 vdd.n202 vdd.n201 0.152939
R4790 vdd.n206 vdd.n202 0.152939
R4791 vdd.n207 vdd.n206 0.152939
R4792 vdd.n208 vdd.n207 0.152939
R4793 vdd.n209 vdd.n208 0.152939
R4794 vdd.n215 vdd.n209 0.152939
R4795 vdd.n2601 vdd.n215 0.152939
R4796 vdd.n2506 vdd.n279 0.152939
R4797 vdd.n2507 vdd.n2506 0.152939
R4798 vdd.n2508 vdd.n2507 0.152939
R4799 vdd.n2508 vdd.n266 0.152939
R4800 vdd.n2522 vdd.n266 0.152939
R4801 vdd.n2523 vdd.n2522 0.152939
R4802 vdd.n2524 vdd.n2523 0.152939
R4803 vdd.n2524 vdd.n255 0.152939
R4804 vdd.n2538 vdd.n255 0.152939
R4805 vdd.n2539 vdd.n2538 0.152939
R4806 vdd.n2540 vdd.n2539 0.152939
R4807 vdd.n2540 vdd.n242 0.152939
R4808 vdd.n2554 vdd.n242 0.152939
R4809 vdd.n2555 vdd.n2554 0.152939
R4810 vdd.n2556 vdd.n2555 0.152939
R4811 vdd.n2556 vdd.n230 0.152939
R4812 vdd.n2570 vdd.n230 0.152939
R4813 vdd.n2571 vdd.n2570 0.152939
R4814 vdd.n2572 vdd.n2571 0.152939
R4815 vdd.n2572 vdd.n228 0.152939
R4816 vdd.n2576 vdd.n228 0.152939
R4817 vdd.n2577 vdd.n2576 0.152939
R4818 vdd.n2578 vdd.n2577 0.152939
R4819 vdd.n2578 vdd.n225 0.152939
R4820 vdd.n2582 vdd.n225 0.152939
R4821 vdd.n2583 vdd.n2582 0.152939
R4822 vdd.n2584 vdd.n2583 0.152939
R4823 vdd.n2584 vdd.n222 0.152939
R4824 vdd.n2588 vdd.n222 0.152939
R4825 vdd.n2589 vdd.n2588 0.152939
R4826 vdd.n2590 vdd.n2589 0.152939
R4827 vdd.n2590 vdd.n219 0.152939
R4828 vdd.n2594 vdd.n219 0.152939
R4829 vdd.n2595 vdd.n2594 0.152939
R4830 vdd.n2596 vdd.n2595 0.152939
R4831 vdd.n2596 vdd.n216 0.152939
R4832 vdd.n2600 vdd.n216 0.152939
R4833 vdd.n2375 vdd.n366 0.152939
R4834 vdd.n2376 vdd.n2375 0.152939
R4835 vdd.n2377 vdd.n2376 0.152939
R4836 vdd.n2378 vdd.n2377 0.152939
R4837 vdd.n1422 vdd.n711 0.152939
R4838 vdd.n1418 vdd.n711 0.152939
R4839 vdd.n1418 vdd.n1417 0.152939
R4840 vdd.n1417 vdd.n1416 0.152939
R4841 vdd.n1087 vdd.n864 0.152939
R4842 vdd.n1088 vdd.n1087 0.152939
R4843 vdd.n1089 vdd.n1088 0.152939
R4844 vdd.n1089 vdd.n851 0.152939
R4845 vdd.n1103 vdd.n851 0.152939
R4846 vdd.n1104 vdd.n1103 0.152939
R4847 vdd.n1105 vdd.n1104 0.152939
R4848 vdd.n1105 vdd.n840 0.152939
R4849 vdd.n1119 vdd.n840 0.152939
R4850 vdd.n1120 vdd.n1119 0.152939
R4851 vdd.n1121 vdd.n1120 0.152939
R4852 vdd.n1121 vdd.n827 0.152939
R4853 vdd.n1135 vdd.n827 0.152939
R4854 vdd.n1136 vdd.n1135 0.152939
R4855 vdd.n1137 vdd.n1136 0.152939
R4856 vdd.n1137 vdd.n816 0.152939
R4857 vdd.n1152 vdd.n816 0.152939
R4858 vdd.n1153 vdd.n1152 0.152939
R4859 vdd.n1154 vdd.n1153 0.152939
R4860 vdd.n1154 vdd.n773 0.152939
R4861 vdd.n1168 vdd.n773 0.152939
R4862 vdd.n1169 vdd.n1168 0.152939
R4863 vdd.n1170 vdd.n1169 0.152939
R4864 vdd.n1170 vdd.n762 0.152939
R4865 vdd.n1184 vdd.n762 0.152939
R4866 vdd.n1185 vdd.n1184 0.152939
R4867 vdd.n1186 vdd.n1185 0.152939
R4868 vdd.n1186 vdd.n749 0.152939
R4869 vdd.n1200 vdd.n749 0.152939
R4870 vdd.n1201 vdd.n1200 0.152939
R4871 vdd.n1202 vdd.n1201 0.152939
R4872 vdd.n1202 vdd.n738 0.152939
R4873 vdd.n1216 vdd.n738 0.152939
R4874 vdd.n1217 vdd.n1216 0.152939
R4875 vdd.n1219 vdd.n1217 0.152939
R4876 vdd.n1219 vdd.n1218 0.152939
R4877 vdd.n1218 vdd.n717 0.152939
R4878 vdd.n1079 vdd.n870 0.152939
R4879 vdd.n1072 vdd.n870 0.152939
R4880 vdd.n1072 vdd.n1071 0.152939
R4881 vdd.n1071 vdd.n1070 0.152939
R4882 vdd.n1070 vdd.n903 0.152939
R4883 vdd.n1066 vdd.n903 0.152939
R4884 vdd.n1066 vdd.n1065 0.152939
R4885 vdd.n1065 vdd.n1064 0.152939
R4886 vdd.n1064 vdd.n909 0.152939
R4887 vdd.n1060 vdd.n909 0.152939
R4888 vdd.n1060 vdd.n1059 0.152939
R4889 vdd.n1059 vdd.n1058 0.152939
R4890 vdd.n1058 vdd.n915 0.152939
R4891 vdd.n1054 vdd.n915 0.152939
R4892 vdd.n1054 vdd.n1053 0.152939
R4893 vdd.n1053 vdd.n1052 0.152939
R4894 vdd.n1052 vdd.n921 0.152939
R4895 vdd.n1045 vdd.n921 0.152939
R4896 vdd.n1045 vdd.n1044 0.152939
R4897 vdd.n1044 vdd.n1043 0.152939
R4898 vdd.n1043 vdd.n926 0.152939
R4899 vdd.n1039 vdd.n926 0.152939
R4900 vdd.n1039 vdd.n1038 0.152939
R4901 vdd.n1038 vdd.n1037 0.152939
R4902 vdd.n1037 vdd.n932 0.152939
R4903 vdd.n1033 vdd.n932 0.152939
R4904 vdd.n1033 vdd.n1032 0.152939
R4905 vdd.n1032 vdd.n1031 0.152939
R4906 vdd.n1031 vdd.n938 0.152939
R4907 vdd.n1027 vdd.n938 0.152939
R4908 vdd.n1027 vdd.n1026 0.152939
R4909 vdd.n1026 vdd.n1025 0.152939
R4910 vdd.n1025 vdd.n944 0.152939
R4911 vdd.n1021 vdd.n944 0.152939
R4912 vdd.n1021 vdd.n1020 0.152939
R4913 vdd.n1020 vdd.n1019 0.152939
R4914 vdd.n1019 vdd.n950 0.152939
R4915 vdd.n1012 vdd.n950 0.152939
R4916 vdd.n1012 vdd.n1011 0.152939
R4917 vdd.n1011 vdd.n1010 0.152939
R4918 vdd.n1010 vdd.n955 0.152939
R4919 vdd.n1006 vdd.n955 0.152939
R4920 vdd.n1006 vdd.n1005 0.152939
R4921 vdd.n1005 vdd.n1004 0.152939
R4922 vdd.n1004 vdd.n961 0.152939
R4923 vdd.n1000 vdd.n961 0.152939
R4924 vdd.n1000 vdd.n999 0.152939
R4925 vdd.n999 vdd.n998 0.152939
R4926 vdd.n998 vdd.n967 0.152939
R4927 vdd.n994 vdd.n967 0.152939
R4928 vdd.n994 vdd.n993 0.152939
R4929 vdd.n993 vdd.n992 0.152939
R4930 vdd.n992 vdd.n973 0.152939
R4931 vdd.n988 vdd.n973 0.152939
R4932 vdd.n988 vdd.n987 0.152939
R4933 vdd.n987 vdd.n986 0.152939
R4934 vdd.n986 vdd.n979 0.152939
R4935 vdd.n1081 vdd.n1080 0.152939
R4936 vdd.n1081 vdd.n858 0.152939
R4937 vdd.n1095 vdd.n858 0.152939
R4938 vdd.n1096 vdd.n1095 0.152939
R4939 vdd.n1097 vdd.n1096 0.152939
R4940 vdd.n1097 vdd.n846 0.152939
R4941 vdd.n1111 vdd.n846 0.152939
R4942 vdd.n1112 vdd.n1111 0.152939
R4943 vdd.n1113 vdd.n1112 0.152939
R4944 vdd.n1113 vdd.n834 0.152939
R4945 vdd.n1127 vdd.n834 0.152939
R4946 vdd.n1128 vdd.n1127 0.152939
R4947 vdd.n1129 vdd.n1128 0.152939
R4948 vdd.n1129 vdd.n822 0.152939
R4949 vdd.n1143 vdd.n822 0.152939
R4950 vdd.n1144 vdd.n1143 0.152939
R4951 vdd.n1146 vdd.n1144 0.152939
R4952 vdd.n1146 vdd.n1145 0.152939
R4953 vdd.n1397 vdd.n1233 0.110256
R4954 vdd.n2485 vdd.n320 0.110256
R4955 vdd.n2393 vdd.n366 0.110256
R4956 vdd.n1423 vdd.n1422 0.110256
R4957 vdd.n1160 vdd.n810 0.0695946
R4958 vdd.n2749 vdd.n58 0.0695946
R4959 vdd.n2749 vdd.n2748 0.0695946
R4960 vdd.n1145 vdd.n810 0.0695946
R4961 vdd.n1397 vdd.n1237 0.0431829
R4962 vdd.n1423 vdd.n708 0.0431829
R4963 vdd.n2485 vdd.n322 0.0431829
R4964 vdd.n2393 vdd.n364 0.0431829
R4965 vdd vdd.n28 0.00833333
R4966 commonsourceibias.n201 commonsourceibias.n139 161.3
R4967 commonsourceibias.n200 commonsourceibias.n199 161.3
R4968 commonsourceibias.n198 commonsourceibias.n140 161.3
R4969 commonsourceibias.n197 commonsourceibias.n196 161.3
R4970 commonsourceibias.n194 commonsourceibias.n141 161.3
R4971 commonsourceibias.n193 commonsourceibias.n192 161.3
R4972 commonsourceibias.n191 commonsourceibias.n142 161.3
R4973 commonsourceibias.n190 commonsourceibias.n189 161.3
R4974 commonsourceibias.n188 commonsourceibias.n143 161.3
R4975 commonsourceibias.n186 commonsourceibias.n185 161.3
R4976 commonsourceibias.n184 commonsourceibias.n144 161.3
R4977 commonsourceibias.n183 commonsourceibias.n182 161.3
R4978 commonsourceibias.n181 commonsourceibias.n145 161.3
R4979 commonsourceibias.n180 commonsourceibias.n179 161.3
R4980 commonsourceibias.n178 commonsourceibias.n177 161.3
R4981 commonsourceibias.n176 commonsourceibias.n147 161.3
R4982 commonsourceibias.n175 commonsourceibias.n174 161.3
R4983 commonsourceibias.n173 commonsourceibias.n148 161.3
R4984 commonsourceibias.n172 commonsourceibias.n171 161.3
R4985 commonsourceibias.n170 commonsourceibias.n149 161.3
R4986 commonsourceibias.n169 commonsourceibias.n168 161.3
R4987 commonsourceibias.n167 commonsourceibias.n151 161.3
R4988 commonsourceibias.n166 commonsourceibias.n165 161.3
R4989 commonsourceibias.n163 commonsourceibias.n152 161.3
R4990 commonsourceibias.n162 commonsourceibias.n161 161.3
R4991 commonsourceibias.n160 commonsourceibias.n153 161.3
R4992 commonsourceibias.n159 commonsourceibias.n158 161.3
R4993 commonsourceibias.n157 commonsourceibias.n154 161.3
R4994 commonsourceibias.n28 commonsourceibias.n25 161.3
R4995 commonsourceibias.n30 commonsourceibias.n29 161.3
R4996 commonsourceibias.n31 commonsourceibias.n24 161.3
R4997 commonsourceibias.n33 commonsourceibias.n32 161.3
R4998 commonsourceibias.n34 commonsourceibias.n23 161.3
R4999 commonsourceibias.n37 commonsourceibias.n36 161.3
R5000 commonsourceibias.n38 commonsourceibias.n22 161.3
R5001 commonsourceibias.n40 commonsourceibias.n39 161.3
R5002 commonsourceibias.n41 commonsourceibias.n20 161.3
R5003 commonsourceibias.n43 commonsourceibias.n42 161.3
R5004 commonsourceibias.n44 commonsourceibias.n19 161.3
R5005 commonsourceibias.n46 commonsourceibias.n45 161.3
R5006 commonsourceibias.n47 commonsourceibias.n18 161.3
R5007 commonsourceibias.n49 commonsourceibias.n48 161.3
R5008 commonsourceibias.n51 commonsourceibias.n50 161.3
R5009 commonsourceibias.n52 commonsourceibias.n16 161.3
R5010 commonsourceibias.n54 commonsourceibias.n53 161.3
R5011 commonsourceibias.n55 commonsourceibias.n15 161.3
R5012 commonsourceibias.n57 commonsourceibias.n56 161.3
R5013 commonsourceibias.n59 commonsourceibias.n14 161.3
R5014 commonsourceibias.n61 commonsourceibias.n60 161.3
R5015 commonsourceibias.n62 commonsourceibias.n13 161.3
R5016 commonsourceibias.n64 commonsourceibias.n63 161.3
R5017 commonsourceibias.n65 commonsourceibias.n12 161.3
R5018 commonsourceibias.n68 commonsourceibias.n67 161.3
R5019 commonsourceibias.n69 commonsourceibias.n11 161.3
R5020 commonsourceibias.n71 commonsourceibias.n70 161.3
R5021 commonsourceibias.n72 commonsourceibias.n10 161.3
R5022 commonsourceibias.n92 commonsourceibias.n89 161.3
R5023 commonsourceibias.n94 commonsourceibias.n93 161.3
R5024 commonsourceibias.n95 commonsourceibias.n88 161.3
R5025 commonsourceibias.n97 commonsourceibias.n96 161.3
R5026 commonsourceibias.n98 commonsourceibias.n87 161.3
R5027 commonsourceibias.n101 commonsourceibias.n100 161.3
R5028 commonsourceibias.n102 commonsourceibias.n86 161.3
R5029 commonsourceibias.n104 commonsourceibias.n103 161.3
R5030 commonsourceibias.n105 commonsourceibias.n84 161.3
R5031 commonsourceibias.n107 commonsourceibias.n106 161.3
R5032 commonsourceibias.n108 commonsourceibias.n9 161.3
R5033 commonsourceibias.n110 commonsourceibias.n109 161.3
R5034 commonsourceibias.n111 commonsourceibias.n8 161.3
R5035 commonsourceibias.n113 commonsourceibias.n112 161.3
R5036 commonsourceibias.n115 commonsourceibias.n114 161.3
R5037 commonsourceibias.n116 commonsourceibias.n6 161.3
R5038 commonsourceibias.n118 commonsourceibias.n117 161.3
R5039 commonsourceibias.n119 commonsourceibias.n5 161.3
R5040 commonsourceibias.n121 commonsourceibias.n120 161.3
R5041 commonsourceibias.n123 commonsourceibias.n4 161.3
R5042 commonsourceibias.n125 commonsourceibias.n124 161.3
R5043 commonsourceibias.n126 commonsourceibias.n3 161.3
R5044 commonsourceibias.n128 commonsourceibias.n127 161.3
R5045 commonsourceibias.n129 commonsourceibias.n2 161.3
R5046 commonsourceibias.n132 commonsourceibias.n131 161.3
R5047 commonsourceibias.n133 commonsourceibias.n1 161.3
R5048 commonsourceibias.n135 commonsourceibias.n134 161.3
R5049 commonsourceibias.n136 commonsourceibias.n0 161.3
R5050 commonsourceibias.n406 commonsourceibias.n344 161.3
R5051 commonsourceibias.n405 commonsourceibias.n404 161.3
R5052 commonsourceibias.n403 commonsourceibias.n345 161.3
R5053 commonsourceibias.n402 commonsourceibias.n401 161.3
R5054 commonsourceibias.n399 commonsourceibias.n346 161.3
R5055 commonsourceibias.n398 commonsourceibias.n397 161.3
R5056 commonsourceibias.n396 commonsourceibias.n347 161.3
R5057 commonsourceibias.n395 commonsourceibias.n394 161.3
R5058 commonsourceibias.n393 commonsourceibias.n348 161.3
R5059 commonsourceibias.n391 commonsourceibias.n390 161.3
R5060 commonsourceibias.n389 commonsourceibias.n349 161.3
R5061 commonsourceibias.n388 commonsourceibias.n387 161.3
R5062 commonsourceibias.n386 commonsourceibias.n350 161.3
R5063 commonsourceibias.n385 commonsourceibias.n384 161.3
R5064 commonsourceibias.n383 commonsourceibias.n382 161.3
R5065 commonsourceibias.n381 commonsourceibias.n352 161.3
R5066 commonsourceibias.n380 commonsourceibias.n379 161.3
R5067 commonsourceibias.n378 commonsourceibias.n353 161.3
R5068 commonsourceibias.n377 commonsourceibias.n376 161.3
R5069 commonsourceibias.n374 commonsourceibias.n354 161.3
R5070 commonsourceibias.n373 commonsourceibias.n372 161.3
R5071 commonsourceibias.n371 commonsourceibias.n355 161.3
R5072 commonsourceibias.n370 commonsourceibias.n369 161.3
R5073 commonsourceibias.n367 commonsourceibias.n356 161.3
R5074 commonsourceibias.n366 commonsourceibias.n365 161.3
R5075 commonsourceibias.n364 commonsourceibias.n357 161.3
R5076 commonsourceibias.n363 commonsourceibias.n362 161.3
R5077 commonsourceibias.n361 commonsourceibias.n358 161.3
R5078 commonsourceibias.n305 commonsourceibias.n243 161.3
R5079 commonsourceibias.n304 commonsourceibias.n303 161.3
R5080 commonsourceibias.n302 commonsourceibias.n244 161.3
R5081 commonsourceibias.n301 commonsourceibias.n300 161.3
R5082 commonsourceibias.n298 commonsourceibias.n245 161.3
R5083 commonsourceibias.n297 commonsourceibias.n296 161.3
R5084 commonsourceibias.n295 commonsourceibias.n246 161.3
R5085 commonsourceibias.n294 commonsourceibias.n293 161.3
R5086 commonsourceibias.n292 commonsourceibias.n247 161.3
R5087 commonsourceibias.n290 commonsourceibias.n289 161.3
R5088 commonsourceibias.n288 commonsourceibias.n248 161.3
R5089 commonsourceibias.n287 commonsourceibias.n286 161.3
R5090 commonsourceibias.n285 commonsourceibias.n249 161.3
R5091 commonsourceibias.n284 commonsourceibias.n283 161.3
R5092 commonsourceibias.n282 commonsourceibias.n281 161.3
R5093 commonsourceibias.n280 commonsourceibias.n251 161.3
R5094 commonsourceibias.n279 commonsourceibias.n278 161.3
R5095 commonsourceibias.n277 commonsourceibias.n252 161.3
R5096 commonsourceibias.n276 commonsourceibias.n275 161.3
R5097 commonsourceibias.n273 commonsourceibias.n253 161.3
R5098 commonsourceibias.n272 commonsourceibias.n271 161.3
R5099 commonsourceibias.n270 commonsourceibias.n254 161.3
R5100 commonsourceibias.n269 commonsourceibias.n268 161.3
R5101 commonsourceibias.n266 commonsourceibias.n255 161.3
R5102 commonsourceibias.n265 commonsourceibias.n264 161.3
R5103 commonsourceibias.n263 commonsourceibias.n256 161.3
R5104 commonsourceibias.n262 commonsourceibias.n261 161.3
R5105 commonsourceibias.n260 commonsourceibias.n257 161.3
R5106 commonsourceibias.n315 commonsourceibias.n314 161.3
R5107 commonsourceibias.n239 commonsourceibias.n214 161.3
R5108 commonsourceibias.n238 commonsourceibias.n237 161.3
R5109 commonsourceibias.n235 commonsourceibias.n215 161.3
R5110 commonsourceibias.n234 commonsourceibias.n233 161.3
R5111 commonsourceibias.n232 commonsourceibias.n216 161.3
R5112 commonsourceibias.n231 commonsourceibias.n230 161.3
R5113 commonsourceibias.n228 commonsourceibias.n217 161.3
R5114 commonsourceibias.n227 commonsourceibias.n226 161.3
R5115 commonsourceibias.n225 commonsourceibias.n218 161.3
R5116 commonsourceibias.n224 commonsourceibias.n223 161.3
R5117 commonsourceibias.n222 commonsourceibias.n219 161.3
R5118 commonsourceibias.n341 commonsourceibias.n205 161.3
R5119 commonsourceibias.n340 commonsourceibias.n339 161.3
R5120 commonsourceibias.n338 commonsourceibias.n206 161.3
R5121 commonsourceibias.n337 commonsourceibias.n336 161.3
R5122 commonsourceibias.n334 commonsourceibias.n207 161.3
R5123 commonsourceibias.n333 commonsourceibias.n332 161.3
R5124 commonsourceibias.n331 commonsourceibias.n208 161.3
R5125 commonsourceibias.n330 commonsourceibias.n329 161.3
R5126 commonsourceibias.n328 commonsourceibias.n209 161.3
R5127 commonsourceibias.n326 commonsourceibias.n325 161.3
R5128 commonsourceibias.n324 commonsourceibias.n210 161.3
R5129 commonsourceibias.n323 commonsourceibias.n322 161.3
R5130 commonsourceibias.n321 commonsourceibias.n211 161.3
R5131 commonsourceibias.n320 commonsourceibias.n319 161.3
R5132 commonsourceibias.n318 commonsourceibias.n317 161.3
R5133 commonsourceibias.n316 commonsourceibias.n213 161.3
R5134 commonsourceibias.n155 commonsourceibias.t39 102.697
R5135 commonsourceibias.n359 commonsourceibias.t50 102.697
R5136 commonsourceibias.n258 commonsourceibias.t24 102.697
R5137 commonsourceibias.n220 commonsourceibias.t56 102.697
R5138 commonsourceibias.n26 commonsourceibias.t26 102.697
R5139 commonsourceibias.n90 commonsourceibias.t44 102.697
R5140 commonsourceibias.n203 commonsourceibias.n202 90.9889
R5141 commonsourceibias.n74 commonsourceibias.n73 90.9889
R5142 commonsourceibias.n138 commonsourceibias.n137 90.9889
R5143 commonsourceibias.n408 commonsourceibias.n407 90.9889
R5144 commonsourceibias.n307 commonsourceibias.n306 90.9889
R5145 commonsourceibias.n343 commonsourceibias.n342 90.9889
R5146 commonsourceibias.n81 commonsourceibias.n79 85.0679
R5147 commonsourceibias.n242 commonsourceibias.n240 85.0679
R5148 commonsourceibias.n81 commonsourceibias.n80 84.0635
R5149 commonsourceibias.n78 commonsourceibias.n77 84.0635
R5150 commonsourceibias.n76 commonsourceibias.n75 84.0635
R5151 commonsourceibias.n309 commonsourceibias.n308 84.0635
R5152 commonsourceibias.n311 commonsourceibias.n310 84.0635
R5153 commonsourceibias.n242 commonsourceibias.n241 84.0635
R5154 commonsourceibias.n156 commonsourceibias.t37 72.3005
R5155 commonsourceibias.n164 commonsourceibias.t47 72.3005
R5156 commonsourceibias.n150 commonsourceibias.t46 72.3005
R5157 commonsourceibias.n146 commonsourceibias.t61 72.3005
R5158 commonsourceibias.n187 commonsourceibias.t63 72.3005
R5159 commonsourceibias.n195 commonsourceibias.t62 72.3005
R5160 commonsourceibias.n202 commonsourceibias.t48 72.3005
R5161 commonsourceibias.n73 commonsourceibias.t30 72.3005
R5162 commonsourceibias.n66 commonsourceibias.t16 72.3005
R5163 commonsourceibias.n58 commonsourceibias.t22 72.3005
R5164 commonsourceibias.n17 commonsourceibias.t18 72.3005
R5165 commonsourceibias.n21 commonsourceibias.t4 72.3005
R5166 commonsourceibias.n35 commonsourceibias.t10 72.3005
R5167 commonsourceibias.n27 commonsourceibias.t12 72.3005
R5168 commonsourceibias.n137 commonsourceibias.t55 72.3005
R5169 commonsourceibias.n130 commonsourceibias.t36 72.3005
R5170 commonsourceibias.n122 commonsourceibias.t40 72.3005
R5171 commonsourceibias.n7 commonsourceibias.t35 72.3005
R5172 commonsourceibias.n85 commonsourceibias.t51 72.3005
R5173 commonsourceibias.n99 commonsourceibias.t52 72.3005
R5174 commonsourceibias.n91 commonsourceibias.t42 72.3005
R5175 commonsourceibias.n360 commonsourceibias.t59 72.3005
R5176 commonsourceibias.n368 commonsourceibias.t38 72.3005
R5177 commonsourceibias.n375 commonsourceibias.t34 72.3005
R5178 commonsourceibias.n351 commonsourceibias.t53 72.3005
R5179 commonsourceibias.n392 commonsourceibias.t45 72.3005
R5180 commonsourceibias.n400 commonsourceibias.t54 72.3005
R5181 commonsourceibias.n407 commonsourceibias.t60 72.3005
R5182 commonsourceibias.n259 commonsourceibias.t6 72.3005
R5183 commonsourceibias.n267 commonsourceibias.t20 72.3005
R5184 commonsourceibias.n274 commonsourceibias.t8 72.3005
R5185 commonsourceibias.n250 commonsourceibias.t0 72.3005
R5186 commonsourceibias.n291 commonsourceibias.t2 72.3005
R5187 commonsourceibias.n299 commonsourceibias.t14 72.3005
R5188 commonsourceibias.n306 commonsourceibias.t28 72.3005
R5189 commonsourceibias.n342 commonsourceibias.t33 72.3005
R5190 commonsourceibias.n335 commonsourceibias.t58 72.3005
R5191 commonsourceibias.n327 commonsourceibias.t49 72.3005
R5192 commonsourceibias.n212 commonsourceibias.t57 72.3005
R5193 commonsourceibias.n221 commonsourceibias.t32 72.3005
R5194 commonsourceibias.n229 commonsourceibias.t43 72.3005
R5195 commonsourceibias.n236 commonsourceibias.t41 72.3005
R5196 commonsourceibias.n27 commonsourceibias.n26 66.3065
R5197 commonsourceibias.n91 commonsourceibias.n90 66.3065
R5198 commonsourceibias.n156 commonsourceibias.n155 66.3065
R5199 commonsourceibias.n360 commonsourceibias.n359 66.3065
R5200 commonsourceibias.n259 commonsourceibias.n258 66.3065
R5201 commonsourceibias.n221 commonsourceibias.n220 66.3065
R5202 commonsourceibias.n176 commonsourceibias.n175 56.5617
R5203 commonsourceibias.n200 commonsourceibias.n140 56.5617
R5204 commonsourceibias.n47 commonsourceibias.n46 56.5617
R5205 commonsourceibias.n111 commonsourceibias.n110 56.5617
R5206 commonsourceibias.n381 commonsourceibias.n380 56.5617
R5207 commonsourceibias.n405 commonsourceibias.n345 56.5617
R5208 commonsourceibias.n280 commonsourceibias.n279 56.5617
R5209 commonsourceibias.n304 commonsourceibias.n244 56.5617
R5210 commonsourceibias.n316 commonsourceibias.n315 56.5617
R5211 commonsourceibias.n71 commonsourceibias.n11 56.5617
R5212 commonsourceibias.n135 commonsourceibias.n1 56.5617
R5213 commonsourceibias.n340 commonsourceibias.n206 56.5617
R5214 commonsourceibias.n162 commonsourceibias.n153 49.296
R5215 commonsourceibias.n189 commonsourceibias.n142 49.296
R5216 commonsourceibias.n60 commonsourceibias.n13 49.296
R5217 commonsourceibias.n33 commonsourceibias.n24 49.296
R5218 commonsourceibias.n124 commonsourceibias.n3 49.296
R5219 commonsourceibias.n97 commonsourceibias.n88 49.296
R5220 commonsourceibias.n366 commonsourceibias.n357 49.296
R5221 commonsourceibias.n394 commonsourceibias.n347 49.296
R5222 commonsourceibias.n265 commonsourceibias.n256 49.296
R5223 commonsourceibias.n293 commonsourceibias.n246 49.296
R5224 commonsourceibias.n329 commonsourceibias.n208 49.296
R5225 commonsourceibias.n227 commonsourceibias.n218 49.296
R5226 commonsourceibias.n169 commonsourceibias.n151 48.3272
R5227 commonsourceibias.n182 commonsourceibias.n144 48.3272
R5228 commonsourceibias.n53 commonsourceibias.n15 48.3272
R5229 commonsourceibias.n40 commonsourceibias.n22 48.3272
R5230 commonsourceibias.n117 commonsourceibias.n5 48.3272
R5231 commonsourceibias.n104 commonsourceibias.n86 48.3272
R5232 commonsourceibias.n373 commonsourceibias.n355 48.3272
R5233 commonsourceibias.n387 commonsourceibias.n349 48.3272
R5234 commonsourceibias.n272 commonsourceibias.n254 48.3272
R5235 commonsourceibias.n286 commonsourceibias.n248 48.3272
R5236 commonsourceibias.n322 commonsourceibias.n210 48.3272
R5237 commonsourceibias.n234 commonsourceibias.n216 48.3272
R5238 commonsourceibias.n170 commonsourceibias.n169 32.8269
R5239 commonsourceibias.n182 commonsourceibias.n181 32.8269
R5240 commonsourceibias.n53 commonsourceibias.n52 32.8269
R5241 commonsourceibias.n41 commonsourceibias.n40 32.8269
R5242 commonsourceibias.n117 commonsourceibias.n116 32.8269
R5243 commonsourceibias.n105 commonsourceibias.n104 32.8269
R5244 commonsourceibias.n374 commonsourceibias.n373 32.8269
R5245 commonsourceibias.n387 commonsourceibias.n386 32.8269
R5246 commonsourceibias.n273 commonsourceibias.n272 32.8269
R5247 commonsourceibias.n286 commonsourceibias.n285 32.8269
R5248 commonsourceibias.n322 commonsourceibias.n321 32.8269
R5249 commonsourceibias.n235 commonsourceibias.n234 32.8269
R5250 commonsourceibias.n158 commonsourceibias.n153 31.8581
R5251 commonsourceibias.n193 commonsourceibias.n142 31.8581
R5252 commonsourceibias.n64 commonsourceibias.n13 31.8581
R5253 commonsourceibias.n29 commonsourceibias.n24 31.8581
R5254 commonsourceibias.n128 commonsourceibias.n3 31.8581
R5255 commonsourceibias.n93 commonsourceibias.n88 31.8581
R5256 commonsourceibias.n362 commonsourceibias.n357 31.8581
R5257 commonsourceibias.n398 commonsourceibias.n347 31.8581
R5258 commonsourceibias.n261 commonsourceibias.n256 31.8581
R5259 commonsourceibias.n297 commonsourceibias.n246 31.8581
R5260 commonsourceibias.n333 commonsourceibias.n208 31.8581
R5261 commonsourceibias.n223 commonsourceibias.n218 31.8581
R5262 commonsourceibias.n158 commonsourceibias.n157 24.5923
R5263 commonsourceibias.n165 commonsourceibias.n151 24.5923
R5264 commonsourceibias.n163 commonsourceibias.n162 24.5923
R5265 commonsourceibias.n175 commonsourceibias.n148 24.5923
R5266 commonsourceibias.n171 commonsourceibias.n170 24.5923
R5267 commonsourceibias.n181 commonsourceibias.n180 24.5923
R5268 commonsourceibias.n177 commonsourceibias.n176 24.5923
R5269 commonsourceibias.n189 commonsourceibias.n188 24.5923
R5270 commonsourceibias.n186 commonsourceibias.n144 24.5923
R5271 commonsourceibias.n196 commonsourceibias.n140 24.5923
R5272 commonsourceibias.n194 commonsourceibias.n193 24.5923
R5273 commonsourceibias.n201 commonsourceibias.n200 24.5923
R5274 commonsourceibias.n72 commonsourceibias.n71 24.5923
R5275 commonsourceibias.n67 commonsourceibias.n11 24.5923
R5276 commonsourceibias.n65 commonsourceibias.n64 24.5923
R5277 commonsourceibias.n60 commonsourceibias.n59 24.5923
R5278 commonsourceibias.n57 commonsourceibias.n15 24.5923
R5279 commonsourceibias.n52 commonsourceibias.n51 24.5923
R5280 commonsourceibias.n48 commonsourceibias.n47 24.5923
R5281 commonsourceibias.n46 commonsourceibias.n19 24.5923
R5282 commonsourceibias.n42 commonsourceibias.n41 24.5923
R5283 commonsourceibias.n36 commonsourceibias.n22 24.5923
R5284 commonsourceibias.n34 commonsourceibias.n33 24.5923
R5285 commonsourceibias.n29 commonsourceibias.n28 24.5923
R5286 commonsourceibias.n136 commonsourceibias.n135 24.5923
R5287 commonsourceibias.n131 commonsourceibias.n1 24.5923
R5288 commonsourceibias.n129 commonsourceibias.n128 24.5923
R5289 commonsourceibias.n124 commonsourceibias.n123 24.5923
R5290 commonsourceibias.n121 commonsourceibias.n5 24.5923
R5291 commonsourceibias.n116 commonsourceibias.n115 24.5923
R5292 commonsourceibias.n112 commonsourceibias.n111 24.5923
R5293 commonsourceibias.n110 commonsourceibias.n9 24.5923
R5294 commonsourceibias.n106 commonsourceibias.n105 24.5923
R5295 commonsourceibias.n100 commonsourceibias.n86 24.5923
R5296 commonsourceibias.n98 commonsourceibias.n97 24.5923
R5297 commonsourceibias.n93 commonsourceibias.n92 24.5923
R5298 commonsourceibias.n362 commonsourceibias.n361 24.5923
R5299 commonsourceibias.n367 commonsourceibias.n366 24.5923
R5300 commonsourceibias.n369 commonsourceibias.n355 24.5923
R5301 commonsourceibias.n376 commonsourceibias.n374 24.5923
R5302 commonsourceibias.n380 commonsourceibias.n353 24.5923
R5303 commonsourceibias.n382 commonsourceibias.n381 24.5923
R5304 commonsourceibias.n386 commonsourceibias.n385 24.5923
R5305 commonsourceibias.n391 commonsourceibias.n349 24.5923
R5306 commonsourceibias.n394 commonsourceibias.n393 24.5923
R5307 commonsourceibias.n399 commonsourceibias.n398 24.5923
R5308 commonsourceibias.n401 commonsourceibias.n345 24.5923
R5309 commonsourceibias.n406 commonsourceibias.n405 24.5923
R5310 commonsourceibias.n261 commonsourceibias.n260 24.5923
R5311 commonsourceibias.n266 commonsourceibias.n265 24.5923
R5312 commonsourceibias.n268 commonsourceibias.n254 24.5923
R5313 commonsourceibias.n275 commonsourceibias.n273 24.5923
R5314 commonsourceibias.n279 commonsourceibias.n252 24.5923
R5315 commonsourceibias.n281 commonsourceibias.n280 24.5923
R5316 commonsourceibias.n285 commonsourceibias.n284 24.5923
R5317 commonsourceibias.n290 commonsourceibias.n248 24.5923
R5318 commonsourceibias.n293 commonsourceibias.n292 24.5923
R5319 commonsourceibias.n298 commonsourceibias.n297 24.5923
R5320 commonsourceibias.n300 commonsourceibias.n244 24.5923
R5321 commonsourceibias.n305 commonsourceibias.n304 24.5923
R5322 commonsourceibias.n341 commonsourceibias.n340 24.5923
R5323 commonsourceibias.n334 commonsourceibias.n333 24.5923
R5324 commonsourceibias.n336 commonsourceibias.n206 24.5923
R5325 commonsourceibias.n326 commonsourceibias.n210 24.5923
R5326 commonsourceibias.n329 commonsourceibias.n328 24.5923
R5327 commonsourceibias.n317 commonsourceibias.n316 24.5923
R5328 commonsourceibias.n321 commonsourceibias.n320 24.5923
R5329 commonsourceibias.n223 commonsourceibias.n222 24.5923
R5330 commonsourceibias.n228 commonsourceibias.n227 24.5923
R5331 commonsourceibias.n230 commonsourceibias.n216 24.5923
R5332 commonsourceibias.n237 commonsourceibias.n235 24.5923
R5333 commonsourceibias.n315 commonsourceibias.n214 24.5923
R5334 commonsourceibias.n196 commonsourceibias.n195 20.9036
R5335 commonsourceibias.n67 commonsourceibias.n66 20.9036
R5336 commonsourceibias.n131 commonsourceibias.n130 20.9036
R5337 commonsourceibias.n401 commonsourceibias.n400 20.9036
R5338 commonsourceibias.n300 commonsourceibias.n299 20.9036
R5339 commonsourceibias.n336 commonsourceibias.n335 20.9036
R5340 commonsourceibias.n150 commonsourceibias.n148 20.4117
R5341 commonsourceibias.n177 commonsourceibias.n146 20.4117
R5342 commonsourceibias.n48 commonsourceibias.n17 20.4117
R5343 commonsourceibias.n21 commonsourceibias.n19 20.4117
R5344 commonsourceibias.n112 commonsourceibias.n7 20.4117
R5345 commonsourceibias.n85 commonsourceibias.n9 20.4117
R5346 commonsourceibias.n375 commonsourceibias.n353 20.4117
R5347 commonsourceibias.n382 commonsourceibias.n351 20.4117
R5348 commonsourceibias.n274 commonsourceibias.n252 20.4117
R5349 commonsourceibias.n281 commonsourceibias.n250 20.4117
R5350 commonsourceibias.n317 commonsourceibias.n212 20.4117
R5351 commonsourceibias.n236 commonsourceibias.n214 20.4117
R5352 commonsourceibias.n202 commonsourceibias.n201 19.9199
R5353 commonsourceibias.n73 commonsourceibias.n72 19.9199
R5354 commonsourceibias.n137 commonsourceibias.n136 19.9199
R5355 commonsourceibias.n407 commonsourceibias.n406 19.9199
R5356 commonsourceibias.n306 commonsourceibias.n305 19.9199
R5357 commonsourceibias.n342 commonsourceibias.n341 19.9199
R5358 commonsourceibias.n155 commonsourceibias.n154 13.3071
R5359 commonsourceibias.n359 commonsourceibias.n358 13.3071
R5360 commonsourceibias.n258 commonsourceibias.n257 13.3071
R5361 commonsourceibias.n220 commonsourceibias.n219 13.3071
R5362 commonsourceibias.n26 commonsourceibias.n25 13.3071
R5363 commonsourceibias.n90 commonsourceibias.n89 13.3071
R5364 commonsourceibias.n76 commonsourceibias.n74 13.0832
R5365 commonsourceibias.n309 commonsourceibias.n307 13.0832
R5366 commonsourceibias.n164 commonsourceibias.n163 12.5423
R5367 commonsourceibias.n188 commonsourceibias.n187 12.5423
R5368 commonsourceibias.n59 commonsourceibias.n58 12.5423
R5369 commonsourceibias.n35 commonsourceibias.n34 12.5423
R5370 commonsourceibias.n123 commonsourceibias.n122 12.5423
R5371 commonsourceibias.n99 commonsourceibias.n98 12.5423
R5372 commonsourceibias.n368 commonsourceibias.n367 12.5423
R5373 commonsourceibias.n393 commonsourceibias.n392 12.5423
R5374 commonsourceibias.n267 commonsourceibias.n266 12.5423
R5375 commonsourceibias.n292 commonsourceibias.n291 12.5423
R5376 commonsourceibias.n328 commonsourceibias.n327 12.5423
R5377 commonsourceibias.n229 commonsourceibias.n228 12.5423
R5378 commonsourceibias.n165 commonsourceibias.n164 12.0505
R5379 commonsourceibias.n187 commonsourceibias.n186 12.0505
R5380 commonsourceibias.n58 commonsourceibias.n57 12.0505
R5381 commonsourceibias.n36 commonsourceibias.n35 12.0505
R5382 commonsourceibias.n122 commonsourceibias.n121 12.0505
R5383 commonsourceibias.n100 commonsourceibias.n99 12.0505
R5384 commonsourceibias.n369 commonsourceibias.n368 12.0505
R5385 commonsourceibias.n392 commonsourceibias.n391 12.0505
R5386 commonsourceibias.n268 commonsourceibias.n267 12.0505
R5387 commonsourceibias.n291 commonsourceibias.n290 12.0505
R5388 commonsourceibias.n327 commonsourceibias.n326 12.0505
R5389 commonsourceibias.n230 commonsourceibias.n229 12.0505
R5390 commonsourceibias.n410 commonsourceibias.n204 11.4057
R5391 commonsourceibias.n410 commonsourceibias.n409 9.95595
R5392 commonsourceibias.n83 commonsourceibias.n82 9.50363
R5393 commonsourceibias.n313 commonsourceibias.n312 9.50363
R5394 commonsourceibias.n204 commonsourceibias.n138 8.39402
R5395 commonsourceibias.n409 commonsourceibias.n343 8.39402
R5396 commonsourceibias.n204 commonsourceibias.n203 5.04553
R5397 commonsourceibias.n409 commonsourceibias.n408 5.04553
R5398 commonsourceibias.n171 commonsourceibias.n150 4.18111
R5399 commonsourceibias.n180 commonsourceibias.n146 4.18111
R5400 commonsourceibias.n51 commonsourceibias.n17 4.18111
R5401 commonsourceibias.n42 commonsourceibias.n21 4.18111
R5402 commonsourceibias.n115 commonsourceibias.n7 4.18111
R5403 commonsourceibias.n106 commonsourceibias.n85 4.18111
R5404 commonsourceibias.n376 commonsourceibias.n375 4.18111
R5405 commonsourceibias.n385 commonsourceibias.n351 4.18111
R5406 commonsourceibias.n275 commonsourceibias.n274 4.18111
R5407 commonsourceibias.n284 commonsourceibias.n250 4.18111
R5408 commonsourceibias.n320 commonsourceibias.n212 4.18111
R5409 commonsourceibias.n237 commonsourceibias.n236 4.18111
R5410 commonsourceibias commonsourceibias.n410 3.92026
R5411 commonsourceibias.n157 commonsourceibias.n156 3.68928
R5412 commonsourceibias.n195 commonsourceibias.n194 3.68928
R5413 commonsourceibias.n66 commonsourceibias.n65 3.68928
R5414 commonsourceibias.n28 commonsourceibias.n27 3.68928
R5415 commonsourceibias.n130 commonsourceibias.n129 3.68928
R5416 commonsourceibias.n92 commonsourceibias.n91 3.68928
R5417 commonsourceibias.n361 commonsourceibias.n360 3.68928
R5418 commonsourceibias.n400 commonsourceibias.n399 3.68928
R5419 commonsourceibias.n260 commonsourceibias.n259 3.68928
R5420 commonsourceibias.n299 commonsourceibias.n298 3.68928
R5421 commonsourceibias.n335 commonsourceibias.n334 3.68928
R5422 commonsourceibias.n222 commonsourceibias.n221 3.68928
R5423 commonsourceibias.n79 commonsourceibias.t13 3.3005
R5424 commonsourceibias.n79 commonsourceibias.t27 3.3005
R5425 commonsourceibias.n80 commonsourceibias.t5 3.3005
R5426 commonsourceibias.n80 commonsourceibias.t11 3.3005
R5427 commonsourceibias.n77 commonsourceibias.t23 3.3005
R5428 commonsourceibias.n77 commonsourceibias.t19 3.3005
R5429 commonsourceibias.n75 commonsourceibias.t31 3.3005
R5430 commonsourceibias.n75 commonsourceibias.t17 3.3005
R5431 commonsourceibias.n308 commonsourceibias.t15 3.3005
R5432 commonsourceibias.n308 commonsourceibias.t29 3.3005
R5433 commonsourceibias.n310 commonsourceibias.t1 3.3005
R5434 commonsourceibias.n310 commonsourceibias.t3 3.3005
R5435 commonsourceibias.n241 commonsourceibias.t21 3.3005
R5436 commonsourceibias.n241 commonsourceibias.t9 3.3005
R5437 commonsourceibias.n240 commonsourceibias.t25 3.3005
R5438 commonsourceibias.n240 commonsourceibias.t7 3.3005
R5439 commonsourceibias.n78 commonsourceibias.n76 1.00481
R5440 commonsourceibias.n311 commonsourceibias.n309 1.00481
R5441 commonsourceibias.n82 commonsourceibias.n78 0.502655
R5442 commonsourceibias.n82 commonsourceibias.n81 0.502655
R5443 commonsourceibias.n312 commonsourceibias.n242 0.502655
R5444 commonsourceibias.n312 commonsourceibias.n311 0.502655
R5445 commonsourceibias.n203 commonsourceibias.n139 0.278335
R5446 commonsourceibias.n74 commonsourceibias.n10 0.278335
R5447 commonsourceibias.n138 commonsourceibias.n0 0.278335
R5448 commonsourceibias.n408 commonsourceibias.n344 0.278335
R5449 commonsourceibias.n307 commonsourceibias.n243 0.278335
R5450 commonsourceibias.n343 commonsourceibias.n205 0.278335
R5451 commonsourceibias.n199 commonsourceibias.n139 0.189894
R5452 commonsourceibias.n199 commonsourceibias.n198 0.189894
R5453 commonsourceibias.n198 commonsourceibias.n197 0.189894
R5454 commonsourceibias.n197 commonsourceibias.n141 0.189894
R5455 commonsourceibias.n192 commonsourceibias.n141 0.189894
R5456 commonsourceibias.n192 commonsourceibias.n191 0.189894
R5457 commonsourceibias.n191 commonsourceibias.n190 0.189894
R5458 commonsourceibias.n190 commonsourceibias.n143 0.189894
R5459 commonsourceibias.n185 commonsourceibias.n143 0.189894
R5460 commonsourceibias.n185 commonsourceibias.n184 0.189894
R5461 commonsourceibias.n184 commonsourceibias.n183 0.189894
R5462 commonsourceibias.n183 commonsourceibias.n145 0.189894
R5463 commonsourceibias.n179 commonsourceibias.n145 0.189894
R5464 commonsourceibias.n179 commonsourceibias.n178 0.189894
R5465 commonsourceibias.n178 commonsourceibias.n147 0.189894
R5466 commonsourceibias.n174 commonsourceibias.n147 0.189894
R5467 commonsourceibias.n174 commonsourceibias.n173 0.189894
R5468 commonsourceibias.n173 commonsourceibias.n172 0.189894
R5469 commonsourceibias.n172 commonsourceibias.n149 0.189894
R5470 commonsourceibias.n168 commonsourceibias.n149 0.189894
R5471 commonsourceibias.n168 commonsourceibias.n167 0.189894
R5472 commonsourceibias.n167 commonsourceibias.n166 0.189894
R5473 commonsourceibias.n166 commonsourceibias.n152 0.189894
R5474 commonsourceibias.n161 commonsourceibias.n152 0.189894
R5475 commonsourceibias.n161 commonsourceibias.n160 0.189894
R5476 commonsourceibias.n160 commonsourceibias.n159 0.189894
R5477 commonsourceibias.n159 commonsourceibias.n154 0.189894
R5478 commonsourceibias.n70 commonsourceibias.n10 0.189894
R5479 commonsourceibias.n70 commonsourceibias.n69 0.189894
R5480 commonsourceibias.n69 commonsourceibias.n68 0.189894
R5481 commonsourceibias.n68 commonsourceibias.n12 0.189894
R5482 commonsourceibias.n63 commonsourceibias.n12 0.189894
R5483 commonsourceibias.n63 commonsourceibias.n62 0.189894
R5484 commonsourceibias.n62 commonsourceibias.n61 0.189894
R5485 commonsourceibias.n61 commonsourceibias.n14 0.189894
R5486 commonsourceibias.n56 commonsourceibias.n14 0.189894
R5487 commonsourceibias.n56 commonsourceibias.n55 0.189894
R5488 commonsourceibias.n55 commonsourceibias.n54 0.189894
R5489 commonsourceibias.n54 commonsourceibias.n16 0.189894
R5490 commonsourceibias.n50 commonsourceibias.n16 0.189894
R5491 commonsourceibias.n50 commonsourceibias.n49 0.189894
R5492 commonsourceibias.n49 commonsourceibias.n18 0.189894
R5493 commonsourceibias.n45 commonsourceibias.n18 0.189894
R5494 commonsourceibias.n45 commonsourceibias.n44 0.189894
R5495 commonsourceibias.n44 commonsourceibias.n43 0.189894
R5496 commonsourceibias.n43 commonsourceibias.n20 0.189894
R5497 commonsourceibias.n39 commonsourceibias.n20 0.189894
R5498 commonsourceibias.n39 commonsourceibias.n38 0.189894
R5499 commonsourceibias.n38 commonsourceibias.n37 0.189894
R5500 commonsourceibias.n37 commonsourceibias.n23 0.189894
R5501 commonsourceibias.n32 commonsourceibias.n23 0.189894
R5502 commonsourceibias.n32 commonsourceibias.n31 0.189894
R5503 commonsourceibias.n31 commonsourceibias.n30 0.189894
R5504 commonsourceibias.n30 commonsourceibias.n25 0.189894
R5505 commonsourceibias.n109 commonsourceibias.n108 0.189894
R5506 commonsourceibias.n108 commonsourceibias.n107 0.189894
R5507 commonsourceibias.n107 commonsourceibias.n84 0.189894
R5508 commonsourceibias.n103 commonsourceibias.n84 0.189894
R5509 commonsourceibias.n103 commonsourceibias.n102 0.189894
R5510 commonsourceibias.n102 commonsourceibias.n101 0.189894
R5511 commonsourceibias.n101 commonsourceibias.n87 0.189894
R5512 commonsourceibias.n96 commonsourceibias.n87 0.189894
R5513 commonsourceibias.n96 commonsourceibias.n95 0.189894
R5514 commonsourceibias.n95 commonsourceibias.n94 0.189894
R5515 commonsourceibias.n94 commonsourceibias.n89 0.189894
R5516 commonsourceibias.n134 commonsourceibias.n0 0.189894
R5517 commonsourceibias.n134 commonsourceibias.n133 0.189894
R5518 commonsourceibias.n133 commonsourceibias.n132 0.189894
R5519 commonsourceibias.n132 commonsourceibias.n2 0.189894
R5520 commonsourceibias.n127 commonsourceibias.n2 0.189894
R5521 commonsourceibias.n127 commonsourceibias.n126 0.189894
R5522 commonsourceibias.n126 commonsourceibias.n125 0.189894
R5523 commonsourceibias.n125 commonsourceibias.n4 0.189894
R5524 commonsourceibias.n120 commonsourceibias.n4 0.189894
R5525 commonsourceibias.n120 commonsourceibias.n119 0.189894
R5526 commonsourceibias.n119 commonsourceibias.n118 0.189894
R5527 commonsourceibias.n118 commonsourceibias.n6 0.189894
R5528 commonsourceibias.n114 commonsourceibias.n6 0.189894
R5529 commonsourceibias.n114 commonsourceibias.n113 0.189894
R5530 commonsourceibias.n113 commonsourceibias.n8 0.189894
R5531 commonsourceibias.n363 commonsourceibias.n358 0.189894
R5532 commonsourceibias.n364 commonsourceibias.n363 0.189894
R5533 commonsourceibias.n365 commonsourceibias.n364 0.189894
R5534 commonsourceibias.n365 commonsourceibias.n356 0.189894
R5535 commonsourceibias.n370 commonsourceibias.n356 0.189894
R5536 commonsourceibias.n371 commonsourceibias.n370 0.189894
R5537 commonsourceibias.n372 commonsourceibias.n371 0.189894
R5538 commonsourceibias.n372 commonsourceibias.n354 0.189894
R5539 commonsourceibias.n377 commonsourceibias.n354 0.189894
R5540 commonsourceibias.n378 commonsourceibias.n377 0.189894
R5541 commonsourceibias.n379 commonsourceibias.n378 0.189894
R5542 commonsourceibias.n379 commonsourceibias.n352 0.189894
R5543 commonsourceibias.n383 commonsourceibias.n352 0.189894
R5544 commonsourceibias.n384 commonsourceibias.n383 0.189894
R5545 commonsourceibias.n384 commonsourceibias.n350 0.189894
R5546 commonsourceibias.n388 commonsourceibias.n350 0.189894
R5547 commonsourceibias.n389 commonsourceibias.n388 0.189894
R5548 commonsourceibias.n390 commonsourceibias.n389 0.189894
R5549 commonsourceibias.n390 commonsourceibias.n348 0.189894
R5550 commonsourceibias.n395 commonsourceibias.n348 0.189894
R5551 commonsourceibias.n396 commonsourceibias.n395 0.189894
R5552 commonsourceibias.n397 commonsourceibias.n396 0.189894
R5553 commonsourceibias.n397 commonsourceibias.n346 0.189894
R5554 commonsourceibias.n402 commonsourceibias.n346 0.189894
R5555 commonsourceibias.n403 commonsourceibias.n402 0.189894
R5556 commonsourceibias.n404 commonsourceibias.n403 0.189894
R5557 commonsourceibias.n404 commonsourceibias.n344 0.189894
R5558 commonsourceibias.n262 commonsourceibias.n257 0.189894
R5559 commonsourceibias.n263 commonsourceibias.n262 0.189894
R5560 commonsourceibias.n264 commonsourceibias.n263 0.189894
R5561 commonsourceibias.n264 commonsourceibias.n255 0.189894
R5562 commonsourceibias.n269 commonsourceibias.n255 0.189894
R5563 commonsourceibias.n270 commonsourceibias.n269 0.189894
R5564 commonsourceibias.n271 commonsourceibias.n270 0.189894
R5565 commonsourceibias.n271 commonsourceibias.n253 0.189894
R5566 commonsourceibias.n276 commonsourceibias.n253 0.189894
R5567 commonsourceibias.n277 commonsourceibias.n276 0.189894
R5568 commonsourceibias.n278 commonsourceibias.n277 0.189894
R5569 commonsourceibias.n278 commonsourceibias.n251 0.189894
R5570 commonsourceibias.n282 commonsourceibias.n251 0.189894
R5571 commonsourceibias.n283 commonsourceibias.n282 0.189894
R5572 commonsourceibias.n283 commonsourceibias.n249 0.189894
R5573 commonsourceibias.n287 commonsourceibias.n249 0.189894
R5574 commonsourceibias.n288 commonsourceibias.n287 0.189894
R5575 commonsourceibias.n289 commonsourceibias.n288 0.189894
R5576 commonsourceibias.n289 commonsourceibias.n247 0.189894
R5577 commonsourceibias.n294 commonsourceibias.n247 0.189894
R5578 commonsourceibias.n295 commonsourceibias.n294 0.189894
R5579 commonsourceibias.n296 commonsourceibias.n295 0.189894
R5580 commonsourceibias.n296 commonsourceibias.n245 0.189894
R5581 commonsourceibias.n301 commonsourceibias.n245 0.189894
R5582 commonsourceibias.n302 commonsourceibias.n301 0.189894
R5583 commonsourceibias.n303 commonsourceibias.n302 0.189894
R5584 commonsourceibias.n303 commonsourceibias.n243 0.189894
R5585 commonsourceibias.n224 commonsourceibias.n219 0.189894
R5586 commonsourceibias.n225 commonsourceibias.n224 0.189894
R5587 commonsourceibias.n226 commonsourceibias.n225 0.189894
R5588 commonsourceibias.n226 commonsourceibias.n217 0.189894
R5589 commonsourceibias.n231 commonsourceibias.n217 0.189894
R5590 commonsourceibias.n232 commonsourceibias.n231 0.189894
R5591 commonsourceibias.n233 commonsourceibias.n232 0.189894
R5592 commonsourceibias.n233 commonsourceibias.n215 0.189894
R5593 commonsourceibias.n238 commonsourceibias.n215 0.189894
R5594 commonsourceibias.n239 commonsourceibias.n238 0.189894
R5595 commonsourceibias.n314 commonsourceibias.n239 0.189894
R5596 commonsourceibias.n318 commonsourceibias.n213 0.189894
R5597 commonsourceibias.n319 commonsourceibias.n318 0.189894
R5598 commonsourceibias.n319 commonsourceibias.n211 0.189894
R5599 commonsourceibias.n323 commonsourceibias.n211 0.189894
R5600 commonsourceibias.n324 commonsourceibias.n323 0.189894
R5601 commonsourceibias.n325 commonsourceibias.n324 0.189894
R5602 commonsourceibias.n325 commonsourceibias.n209 0.189894
R5603 commonsourceibias.n330 commonsourceibias.n209 0.189894
R5604 commonsourceibias.n331 commonsourceibias.n330 0.189894
R5605 commonsourceibias.n332 commonsourceibias.n331 0.189894
R5606 commonsourceibias.n332 commonsourceibias.n207 0.189894
R5607 commonsourceibias.n337 commonsourceibias.n207 0.189894
R5608 commonsourceibias.n338 commonsourceibias.n337 0.189894
R5609 commonsourceibias.n339 commonsourceibias.n338 0.189894
R5610 commonsourceibias.n339 commonsourceibias.n205 0.189894
R5611 commonsourceibias.n109 commonsourceibias.n83 0.0762576
R5612 commonsourceibias.n83 commonsourceibias.n8 0.0762576
R5613 commonsourceibias.n314 commonsourceibias.n313 0.0762576
R5614 commonsourceibias.n313 commonsourceibias.n213 0.0762576
R5615 gnd.n3029 gnd.n2659 2144.37
R5616 gnd.n5116 gnd.n2012 982.702
R5617 gnd.n5010 gnd.n3606 766.379
R5618 gnd.n5032 gnd.n5031 766.379
R5619 gnd.n4035 gnd.n3934 766.379
R5620 gnd.n4033 gnd.n3936 766.379
R5621 gnd.n5807 gnd.n1622 766.379
R5622 gnd.n1043 gnd.n795 766.379
R5623 gnd.n5820 gnd.n1667 766.379
R5624 gnd.n6710 gnd.n993 766.379
R5625 gnd.n7207 gnd.n503 761.573
R5626 gnd.n7354 gnd.n499 761.573
R5627 gnd.n832 gnd.n788 761.573
R5628 gnd.n7014 gnd.n790 761.573
R5629 gnd.n1695 gnd.n1604 761.573
R5630 gnd.n5768 gnd.n1602 761.573
R5631 gnd.n2036 gnd.n2014 761.573
R5632 gnd.n5280 gnd.n2015 761.573
R5633 gnd.n5118 gnd.n3603 756.769
R5634 gnd.n3646 gnd.n3605 756.769
R5635 gnd.n4442 gnd.n3896 756.769
R5636 gnd.n4428 gnd.n3886 756.769
R5637 gnd.n7352 gnd.n505 742.355
R5638 gnd.n569 gnd.n501 742.355
R5639 gnd.n6899 gnd.n787 742.355
R5640 gnd.n7016 gnd.n785 742.355
R5641 gnd.n5957 gnd.n1606 742.355
R5642 gnd.n5959 gnd.n1600 742.355
R5643 gnd.n2172 gnd.n2013 742.355
R5644 gnd.n5282 gnd.n2011 742.355
R5645 gnd.n3376 gnd.n2322 689.5
R5646 gnd.n3030 gnd.n2660 689.5
R5647 gnd.n2898 gnd.n2792 689.5
R5648 gnd.n5169 gnd.n5168 689.5
R5649 gnd.n3377 gnd.n3376 585
R5650 gnd.n3376 gnd.n3375 585
R5651 gnd.n2320 gnd.n2319 585
R5652 gnd.n2319 gnd.n2318 585
R5653 gnd.n3382 gnd.n3381 585
R5654 gnd.n3383 gnd.n3382 585
R5655 gnd.n2317 gnd.n2316 585
R5656 gnd.n3384 gnd.n2317 585
R5657 gnd.n3387 gnd.n3386 585
R5658 gnd.n3386 gnd.n3385 585
R5659 gnd.n2314 gnd.n2313 585
R5660 gnd.n2313 gnd.n2312 585
R5661 gnd.n3392 gnd.n3391 585
R5662 gnd.n3393 gnd.n3392 585
R5663 gnd.n2311 gnd.n2310 585
R5664 gnd.n3394 gnd.n2311 585
R5665 gnd.n3397 gnd.n3396 585
R5666 gnd.n3396 gnd.n3395 585
R5667 gnd.n2308 gnd.n2307 585
R5668 gnd.n2307 gnd.n2306 585
R5669 gnd.n3402 gnd.n3401 585
R5670 gnd.n3403 gnd.n3402 585
R5671 gnd.n2305 gnd.n2304 585
R5672 gnd.n3404 gnd.n2305 585
R5673 gnd.n3407 gnd.n3406 585
R5674 gnd.n3406 gnd.n3405 585
R5675 gnd.n2302 gnd.n2301 585
R5676 gnd.n2301 gnd.n2300 585
R5677 gnd.n3412 gnd.n3411 585
R5678 gnd.n3413 gnd.n3412 585
R5679 gnd.n2299 gnd.n2298 585
R5680 gnd.n3414 gnd.n2299 585
R5681 gnd.n3417 gnd.n3416 585
R5682 gnd.n3416 gnd.n3415 585
R5683 gnd.n2296 gnd.n2295 585
R5684 gnd.n2295 gnd.n2294 585
R5685 gnd.n3422 gnd.n3421 585
R5686 gnd.n3423 gnd.n3422 585
R5687 gnd.n2293 gnd.n2292 585
R5688 gnd.n3424 gnd.n2293 585
R5689 gnd.n3427 gnd.n3426 585
R5690 gnd.n3426 gnd.n3425 585
R5691 gnd.n2290 gnd.n2289 585
R5692 gnd.n2289 gnd.n2288 585
R5693 gnd.n3432 gnd.n3431 585
R5694 gnd.n3433 gnd.n3432 585
R5695 gnd.n2287 gnd.n2286 585
R5696 gnd.n3434 gnd.n2287 585
R5697 gnd.n3437 gnd.n3436 585
R5698 gnd.n3436 gnd.n3435 585
R5699 gnd.n2284 gnd.n2283 585
R5700 gnd.n2283 gnd.n2282 585
R5701 gnd.n3442 gnd.n3441 585
R5702 gnd.n3443 gnd.n3442 585
R5703 gnd.n2281 gnd.n2280 585
R5704 gnd.n3444 gnd.n2281 585
R5705 gnd.n3447 gnd.n3446 585
R5706 gnd.n3446 gnd.n3445 585
R5707 gnd.n2278 gnd.n2277 585
R5708 gnd.n2277 gnd.n2276 585
R5709 gnd.n3452 gnd.n3451 585
R5710 gnd.n3453 gnd.n3452 585
R5711 gnd.n2275 gnd.n2274 585
R5712 gnd.n3454 gnd.n2275 585
R5713 gnd.n3457 gnd.n3456 585
R5714 gnd.n3456 gnd.n3455 585
R5715 gnd.n2272 gnd.n2271 585
R5716 gnd.n2271 gnd.n2270 585
R5717 gnd.n3462 gnd.n3461 585
R5718 gnd.n3463 gnd.n3462 585
R5719 gnd.n2269 gnd.n2268 585
R5720 gnd.n3464 gnd.n2269 585
R5721 gnd.n3467 gnd.n3466 585
R5722 gnd.n3466 gnd.n3465 585
R5723 gnd.n2266 gnd.n2265 585
R5724 gnd.n2265 gnd.n2264 585
R5725 gnd.n3472 gnd.n3471 585
R5726 gnd.n3473 gnd.n3472 585
R5727 gnd.n2263 gnd.n2262 585
R5728 gnd.n3474 gnd.n2263 585
R5729 gnd.n3477 gnd.n3476 585
R5730 gnd.n3476 gnd.n3475 585
R5731 gnd.n2260 gnd.n2259 585
R5732 gnd.n2259 gnd.n2258 585
R5733 gnd.n3482 gnd.n3481 585
R5734 gnd.n3483 gnd.n3482 585
R5735 gnd.n2257 gnd.n2256 585
R5736 gnd.n3484 gnd.n2257 585
R5737 gnd.n3487 gnd.n3486 585
R5738 gnd.n3486 gnd.n3485 585
R5739 gnd.n2254 gnd.n2253 585
R5740 gnd.n2253 gnd.n2252 585
R5741 gnd.n3492 gnd.n3491 585
R5742 gnd.n3493 gnd.n3492 585
R5743 gnd.n2251 gnd.n2250 585
R5744 gnd.n3494 gnd.n2251 585
R5745 gnd.n3497 gnd.n3496 585
R5746 gnd.n3496 gnd.n3495 585
R5747 gnd.n2248 gnd.n2247 585
R5748 gnd.n2247 gnd.n2246 585
R5749 gnd.n3502 gnd.n3501 585
R5750 gnd.n3503 gnd.n3502 585
R5751 gnd.n2245 gnd.n2244 585
R5752 gnd.n3504 gnd.n2245 585
R5753 gnd.n3507 gnd.n3506 585
R5754 gnd.n3506 gnd.n3505 585
R5755 gnd.n2242 gnd.n2241 585
R5756 gnd.n2241 gnd.n2240 585
R5757 gnd.n3512 gnd.n3511 585
R5758 gnd.n3513 gnd.n3512 585
R5759 gnd.n2239 gnd.n2238 585
R5760 gnd.n3514 gnd.n2239 585
R5761 gnd.n3517 gnd.n3516 585
R5762 gnd.n3516 gnd.n3515 585
R5763 gnd.n2236 gnd.n2235 585
R5764 gnd.n2235 gnd.n2234 585
R5765 gnd.n3522 gnd.n3521 585
R5766 gnd.n3523 gnd.n3522 585
R5767 gnd.n2233 gnd.n2232 585
R5768 gnd.n3524 gnd.n2233 585
R5769 gnd.n3527 gnd.n3526 585
R5770 gnd.n3526 gnd.n3525 585
R5771 gnd.n2230 gnd.n2229 585
R5772 gnd.n2229 gnd.n2228 585
R5773 gnd.n3532 gnd.n3531 585
R5774 gnd.n3533 gnd.n3532 585
R5775 gnd.n2227 gnd.n2226 585
R5776 gnd.n3534 gnd.n2227 585
R5777 gnd.n5163 gnd.n5162 585
R5778 gnd.n5162 gnd.n5161 585
R5779 gnd.n2224 gnd.n2223 585
R5780 gnd.n5160 gnd.n2223 585
R5781 gnd.n2325 gnd.n2322 585
R5782 gnd.n3374 gnd.n2322 585
R5783 gnd.n3372 gnd.n3371 585
R5784 gnd.n3373 gnd.n3372 585
R5785 gnd.n3370 gnd.n2324 585
R5786 gnd.n2324 gnd.n2323 585
R5787 gnd.n3369 gnd.n3368 585
R5788 gnd.n3368 gnd.n3367 585
R5789 gnd.n2330 gnd.n2329 585
R5790 gnd.n3366 gnd.n2330 585
R5791 gnd.n3364 gnd.n3363 585
R5792 gnd.n3365 gnd.n3364 585
R5793 gnd.n3362 gnd.n2332 585
R5794 gnd.n2332 gnd.n2331 585
R5795 gnd.n3361 gnd.n3360 585
R5796 gnd.n3360 gnd.n3359 585
R5797 gnd.n2338 gnd.n2337 585
R5798 gnd.n3358 gnd.n2338 585
R5799 gnd.n3356 gnd.n3355 585
R5800 gnd.n3357 gnd.n3356 585
R5801 gnd.n3354 gnd.n2340 585
R5802 gnd.n2340 gnd.n2339 585
R5803 gnd.n3353 gnd.n3352 585
R5804 gnd.n3352 gnd.n3351 585
R5805 gnd.n2346 gnd.n2345 585
R5806 gnd.n3350 gnd.n2346 585
R5807 gnd.n3348 gnd.n3347 585
R5808 gnd.n3349 gnd.n3348 585
R5809 gnd.n3346 gnd.n2348 585
R5810 gnd.n2348 gnd.n2347 585
R5811 gnd.n3345 gnd.n3344 585
R5812 gnd.n3344 gnd.n3343 585
R5813 gnd.n2354 gnd.n2353 585
R5814 gnd.n3342 gnd.n2354 585
R5815 gnd.n3340 gnd.n3339 585
R5816 gnd.n3341 gnd.n3340 585
R5817 gnd.n3338 gnd.n2356 585
R5818 gnd.n2356 gnd.n2355 585
R5819 gnd.n3337 gnd.n3336 585
R5820 gnd.n3336 gnd.n3335 585
R5821 gnd.n2362 gnd.n2361 585
R5822 gnd.n3334 gnd.n2362 585
R5823 gnd.n3332 gnd.n3331 585
R5824 gnd.n3333 gnd.n3332 585
R5825 gnd.n3330 gnd.n2364 585
R5826 gnd.n2364 gnd.n2363 585
R5827 gnd.n3329 gnd.n3328 585
R5828 gnd.n3328 gnd.n3327 585
R5829 gnd.n2370 gnd.n2369 585
R5830 gnd.n3326 gnd.n2370 585
R5831 gnd.n3324 gnd.n3323 585
R5832 gnd.n3325 gnd.n3324 585
R5833 gnd.n3322 gnd.n2372 585
R5834 gnd.n2372 gnd.n2371 585
R5835 gnd.n3321 gnd.n3320 585
R5836 gnd.n3320 gnd.n3319 585
R5837 gnd.n2378 gnd.n2377 585
R5838 gnd.n3318 gnd.n2378 585
R5839 gnd.n3316 gnd.n3315 585
R5840 gnd.n3317 gnd.n3316 585
R5841 gnd.n3314 gnd.n2380 585
R5842 gnd.n2380 gnd.n2379 585
R5843 gnd.n3313 gnd.n3312 585
R5844 gnd.n3312 gnd.n3311 585
R5845 gnd.n2386 gnd.n2385 585
R5846 gnd.n3310 gnd.n2386 585
R5847 gnd.n3308 gnd.n3307 585
R5848 gnd.n3309 gnd.n3308 585
R5849 gnd.n3306 gnd.n2388 585
R5850 gnd.n2388 gnd.n2387 585
R5851 gnd.n3305 gnd.n3304 585
R5852 gnd.n3304 gnd.n3303 585
R5853 gnd.n2394 gnd.n2393 585
R5854 gnd.n3302 gnd.n2394 585
R5855 gnd.n3300 gnd.n3299 585
R5856 gnd.n3301 gnd.n3300 585
R5857 gnd.n3298 gnd.n2396 585
R5858 gnd.n2396 gnd.n2395 585
R5859 gnd.n3297 gnd.n3296 585
R5860 gnd.n3296 gnd.n3295 585
R5861 gnd.n2402 gnd.n2401 585
R5862 gnd.n3294 gnd.n2402 585
R5863 gnd.n3292 gnd.n3291 585
R5864 gnd.n3293 gnd.n3292 585
R5865 gnd.n3290 gnd.n2404 585
R5866 gnd.n2404 gnd.n2403 585
R5867 gnd.n3289 gnd.n3288 585
R5868 gnd.n3288 gnd.n3287 585
R5869 gnd.n2410 gnd.n2409 585
R5870 gnd.n3286 gnd.n2410 585
R5871 gnd.n3284 gnd.n3283 585
R5872 gnd.n3285 gnd.n3284 585
R5873 gnd.n3282 gnd.n2412 585
R5874 gnd.n2412 gnd.n2411 585
R5875 gnd.n3281 gnd.n3280 585
R5876 gnd.n3280 gnd.n3279 585
R5877 gnd.n2418 gnd.n2417 585
R5878 gnd.n3278 gnd.n2418 585
R5879 gnd.n3276 gnd.n3275 585
R5880 gnd.n3277 gnd.n3276 585
R5881 gnd.n3274 gnd.n2420 585
R5882 gnd.n2420 gnd.n2419 585
R5883 gnd.n3273 gnd.n3272 585
R5884 gnd.n3272 gnd.n3271 585
R5885 gnd.n2426 gnd.n2425 585
R5886 gnd.n3270 gnd.n2426 585
R5887 gnd.n3268 gnd.n3267 585
R5888 gnd.n3269 gnd.n3268 585
R5889 gnd.n3266 gnd.n2428 585
R5890 gnd.n2428 gnd.n2427 585
R5891 gnd.n3265 gnd.n3264 585
R5892 gnd.n3264 gnd.n3263 585
R5893 gnd.n2434 gnd.n2433 585
R5894 gnd.n3262 gnd.n2434 585
R5895 gnd.n3260 gnd.n3259 585
R5896 gnd.n3261 gnd.n3260 585
R5897 gnd.n3258 gnd.n2436 585
R5898 gnd.n2436 gnd.n2435 585
R5899 gnd.n3257 gnd.n3256 585
R5900 gnd.n3256 gnd.n3255 585
R5901 gnd.n2442 gnd.n2441 585
R5902 gnd.n3254 gnd.n2442 585
R5903 gnd.n3252 gnd.n3251 585
R5904 gnd.n3253 gnd.n3252 585
R5905 gnd.n3250 gnd.n2444 585
R5906 gnd.n2444 gnd.n2443 585
R5907 gnd.n3249 gnd.n3248 585
R5908 gnd.n3248 gnd.n3247 585
R5909 gnd.n2450 gnd.n2449 585
R5910 gnd.n3246 gnd.n2450 585
R5911 gnd.n3244 gnd.n3243 585
R5912 gnd.n3245 gnd.n3244 585
R5913 gnd.n3242 gnd.n2452 585
R5914 gnd.n2452 gnd.n2451 585
R5915 gnd.n3241 gnd.n3240 585
R5916 gnd.n3240 gnd.n3239 585
R5917 gnd.n2458 gnd.n2457 585
R5918 gnd.n3238 gnd.n2458 585
R5919 gnd.n3236 gnd.n3235 585
R5920 gnd.n3237 gnd.n3236 585
R5921 gnd.n3234 gnd.n2460 585
R5922 gnd.n2460 gnd.n2459 585
R5923 gnd.n3233 gnd.n3232 585
R5924 gnd.n3232 gnd.n3231 585
R5925 gnd.n2466 gnd.n2465 585
R5926 gnd.n3230 gnd.n2466 585
R5927 gnd.n3228 gnd.n3227 585
R5928 gnd.n3229 gnd.n3228 585
R5929 gnd.n3226 gnd.n2468 585
R5930 gnd.n2468 gnd.n2467 585
R5931 gnd.n3225 gnd.n3224 585
R5932 gnd.n3224 gnd.n3223 585
R5933 gnd.n2474 gnd.n2473 585
R5934 gnd.n3222 gnd.n2474 585
R5935 gnd.n3220 gnd.n3219 585
R5936 gnd.n3221 gnd.n3220 585
R5937 gnd.n3218 gnd.n2476 585
R5938 gnd.n2476 gnd.n2475 585
R5939 gnd.n3217 gnd.n3216 585
R5940 gnd.n3216 gnd.n3215 585
R5941 gnd.n2482 gnd.n2481 585
R5942 gnd.n3214 gnd.n2482 585
R5943 gnd.n3212 gnd.n3211 585
R5944 gnd.n3213 gnd.n3212 585
R5945 gnd.n3210 gnd.n2484 585
R5946 gnd.n2484 gnd.n2483 585
R5947 gnd.n3209 gnd.n3208 585
R5948 gnd.n3208 gnd.n3207 585
R5949 gnd.n2490 gnd.n2489 585
R5950 gnd.n3206 gnd.n2490 585
R5951 gnd.n3204 gnd.n3203 585
R5952 gnd.n3205 gnd.n3204 585
R5953 gnd.n3202 gnd.n2492 585
R5954 gnd.n2492 gnd.n2491 585
R5955 gnd.n3201 gnd.n3200 585
R5956 gnd.n3200 gnd.n3199 585
R5957 gnd.n2498 gnd.n2497 585
R5958 gnd.n3198 gnd.n2498 585
R5959 gnd.n3196 gnd.n3195 585
R5960 gnd.n3197 gnd.n3196 585
R5961 gnd.n3194 gnd.n2500 585
R5962 gnd.n2500 gnd.n2499 585
R5963 gnd.n3193 gnd.n3192 585
R5964 gnd.n3192 gnd.n3191 585
R5965 gnd.n2506 gnd.n2505 585
R5966 gnd.n3190 gnd.n2506 585
R5967 gnd.n3188 gnd.n3187 585
R5968 gnd.n3189 gnd.n3188 585
R5969 gnd.n3186 gnd.n2508 585
R5970 gnd.n2508 gnd.n2507 585
R5971 gnd.n3185 gnd.n3184 585
R5972 gnd.n3184 gnd.n3183 585
R5973 gnd.n2514 gnd.n2513 585
R5974 gnd.n3182 gnd.n2514 585
R5975 gnd.n3180 gnd.n3179 585
R5976 gnd.n3181 gnd.n3180 585
R5977 gnd.n3178 gnd.n2516 585
R5978 gnd.n2516 gnd.n2515 585
R5979 gnd.n3177 gnd.n3176 585
R5980 gnd.n3176 gnd.n3175 585
R5981 gnd.n2522 gnd.n2521 585
R5982 gnd.n3174 gnd.n2522 585
R5983 gnd.n3172 gnd.n3171 585
R5984 gnd.n3173 gnd.n3172 585
R5985 gnd.n3170 gnd.n2524 585
R5986 gnd.n2524 gnd.n2523 585
R5987 gnd.n3169 gnd.n3168 585
R5988 gnd.n3168 gnd.n3167 585
R5989 gnd.n2530 gnd.n2529 585
R5990 gnd.n3166 gnd.n2530 585
R5991 gnd.n3164 gnd.n3163 585
R5992 gnd.n3165 gnd.n3164 585
R5993 gnd.n3162 gnd.n2532 585
R5994 gnd.n2532 gnd.n2531 585
R5995 gnd.n3161 gnd.n3160 585
R5996 gnd.n3160 gnd.n3159 585
R5997 gnd.n2538 gnd.n2537 585
R5998 gnd.n3158 gnd.n2538 585
R5999 gnd.n3156 gnd.n3155 585
R6000 gnd.n3157 gnd.n3156 585
R6001 gnd.n3154 gnd.n2540 585
R6002 gnd.n2540 gnd.n2539 585
R6003 gnd.n3153 gnd.n3152 585
R6004 gnd.n3152 gnd.n3151 585
R6005 gnd.n2546 gnd.n2545 585
R6006 gnd.n3150 gnd.n2546 585
R6007 gnd.n3148 gnd.n3147 585
R6008 gnd.n3149 gnd.n3148 585
R6009 gnd.n3146 gnd.n2548 585
R6010 gnd.n2548 gnd.n2547 585
R6011 gnd.n3145 gnd.n3144 585
R6012 gnd.n3144 gnd.n3143 585
R6013 gnd.n2554 gnd.n2553 585
R6014 gnd.n3142 gnd.n2554 585
R6015 gnd.n3140 gnd.n3139 585
R6016 gnd.n3141 gnd.n3140 585
R6017 gnd.n3138 gnd.n2556 585
R6018 gnd.n2556 gnd.n2555 585
R6019 gnd.n3137 gnd.n3136 585
R6020 gnd.n3136 gnd.n3135 585
R6021 gnd.n2562 gnd.n2561 585
R6022 gnd.n3134 gnd.n2562 585
R6023 gnd.n3132 gnd.n3131 585
R6024 gnd.n3133 gnd.n3132 585
R6025 gnd.n3130 gnd.n2564 585
R6026 gnd.n2564 gnd.n2563 585
R6027 gnd.n3129 gnd.n3128 585
R6028 gnd.n3128 gnd.n3127 585
R6029 gnd.n2570 gnd.n2569 585
R6030 gnd.n3126 gnd.n2570 585
R6031 gnd.n3124 gnd.n3123 585
R6032 gnd.n3125 gnd.n3124 585
R6033 gnd.n3122 gnd.n2572 585
R6034 gnd.n2572 gnd.n2571 585
R6035 gnd.n3121 gnd.n3120 585
R6036 gnd.n3120 gnd.n3119 585
R6037 gnd.n2578 gnd.n2577 585
R6038 gnd.n3118 gnd.n2578 585
R6039 gnd.n3116 gnd.n3115 585
R6040 gnd.n3117 gnd.n3116 585
R6041 gnd.n3114 gnd.n2580 585
R6042 gnd.n2580 gnd.n2579 585
R6043 gnd.n3113 gnd.n3112 585
R6044 gnd.n3112 gnd.n3111 585
R6045 gnd.n2586 gnd.n2585 585
R6046 gnd.n3110 gnd.n2586 585
R6047 gnd.n3108 gnd.n3107 585
R6048 gnd.n3109 gnd.n3108 585
R6049 gnd.n3106 gnd.n2588 585
R6050 gnd.n2588 gnd.n2587 585
R6051 gnd.n3105 gnd.n3104 585
R6052 gnd.n3104 gnd.n3103 585
R6053 gnd.n2594 gnd.n2593 585
R6054 gnd.n3102 gnd.n2594 585
R6055 gnd.n3100 gnd.n3099 585
R6056 gnd.n3101 gnd.n3100 585
R6057 gnd.n3098 gnd.n2596 585
R6058 gnd.n2596 gnd.n2595 585
R6059 gnd.n3097 gnd.n3096 585
R6060 gnd.n3096 gnd.n3095 585
R6061 gnd.n2602 gnd.n2601 585
R6062 gnd.n3094 gnd.n2602 585
R6063 gnd.n3092 gnd.n3091 585
R6064 gnd.n3093 gnd.n3092 585
R6065 gnd.n3090 gnd.n2604 585
R6066 gnd.n2604 gnd.n2603 585
R6067 gnd.n3089 gnd.n3088 585
R6068 gnd.n3088 gnd.n3087 585
R6069 gnd.n2610 gnd.n2609 585
R6070 gnd.n3086 gnd.n2610 585
R6071 gnd.n3084 gnd.n3083 585
R6072 gnd.n3085 gnd.n3084 585
R6073 gnd.n3082 gnd.n2612 585
R6074 gnd.n2612 gnd.n2611 585
R6075 gnd.n3081 gnd.n3080 585
R6076 gnd.n3080 gnd.n3079 585
R6077 gnd.n2618 gnd.n2617 585
R6078 gnd.n3078 gnd.n2618 585
R6079 gnd.n3076 gnd.n3075 585
R6080 gnd.n3077 gnd.n3076 585
R6081 gnd.n3074 gnd.n2620 585
R6082 gnd.n2620 gnd.n2619 585
R6083 gnd.n3073 gnd.n3072 585
R6084 gnd.n3072 gnd.n3071 585
R6085 gnd.n2626 gnd.n2625 585
R6086 gnd.n3070 gnd.n2626 585
R6087 gnd.n3068 gnd.n3067 585
R6088 gnd.n3069 gnd.n3068 585
R6089 gnd.n3066 gnd.n2628 585
R6090 gnd.n2628 gnd.n2627 585
R6091 gnd.n3065 gnd.n3064 585
R6092 gnd.n3064 gnd.n3063 585
R6093 gnd.n2634 gnd.n2633 585
R6094 gnd.n3062 gnd.n2634 585
R6095 gnd.n3060 gnd.n3059 585
R6096 gnd.n3061 gnd.n3060 585
R6097 gnd.n3058 gnd.n2636 585
R6098 gnd.n2636 gnd.n2635 585
R6099 gnd.n3057 gnd.n3056 585
R6100 gnd.n3056 gnd.n3055 585
R6101 gnd.n2642 gnd.n2641 585
R6102 gnd.n3054 gnd.n2642 585
R6103 gnd.n3052 gnd.n3051 585
R6104 gnd.n3053 gnd.n3052 585
R6105 gnd.n3050 gnd.n2644 585
R6106 gnd.n2644 gnd.n2643 585
R6107 gnd.n3049 gnd.n3048 585
R6108 gnd.n3048 gnd.n3047 585
R6109 gnd.n2650 gnd.n2649 585
R6110 gnd.n3046 gnd.n2650 585
R6111 gnd.n3044 gnd.n3043 585
R6112 gnd.n3045 gnd.n3044 585
R6113 gnd.n3042 gnd.n2652 585
R6114 gnd.n2652 gnd.n2651 585
R6115 gnd.n3041 gnd.n3040 585
R6116 gnd.n3040 gnd.n3039 585
R6117 gnd.n2658 gnd.n2657 585
R6118 gnd.n3038 gnd.n2658 585
R6119 gnd.n3036 gnd.n3035 585
R6120 gnd.n3037 gnd.n3036 585
R6121 gnd.n3034 gnd.n2660 585
R6122 gnd.n2660 gnd.n2659 585
R6123 gnd.n2899 gnd.n2791 585
R6124 gnd.n2900 gnd.n2899 585
R6125 gnd.n2903 gnd.n2902 585
R6126 gnd.n2902 gnd.n2901 585
R6127 gnd.n2904 gnd.n2786 585
R6128 gnd.n2786 gnd.n2785 585
R6129 gnd.n2906 gnd.n2905 585
R6130 gnd.n2907 gnd.n2906 585
R6131 gnd.n2784 gnd.n2783 585
R6132 gnd.n2908 gnd.n2784 585
R6133 gnd.n2911 gnd.n2910 585
R6134 gnd.n2910 gnd.n2909 585
R6135 gnd.n2912 gnd.n2778 585
R6136 gnd.n2778 gnd.n2777 585
R6137 gnd.n2914 gnd.n2913 585
R6138 gnd.n2915 gnd.n2914 585
R6139 gnd.n2776 gnd.n2775 585
R6140 gnd.n2916 gnd.n2776 585
R6141 gnd.n2919 gnd.n2918 585
R6142 gnd.n2918 gnd.n2917 585
R6143 gnd.n2920 gnd.n2770 585
R6144 gnd.n2770 gnd.n2769 585
R6145 gnd.n2922 gnd.n2921 585
R6146 gnd.n2923 gnd.n2922 585
R6147 gnd.n2768 gnd.n2767 585
R6148 gnd.n2924 gnd.n2768 585
R6149 gnd.n2927 gnd.n2926 585
R6150 gnd.n2926 gnd.n2925 585
R6151 gnd.n2928 gnd.n2762 585
R6152 gnd.n2762 gnd.n2761 585
R6153 gnd.n2930 gnd.n2929 585
R6154 gnd.n2931 gnd.n2930 585
R6155 gnd.n2760 gnd.n2759 585
R6156 gnd.n2932 gnd.n2760 585
R6157 gnd.n2935 gnd.n2934 585
R6158 gnd.n2934 gnd.n2933 585
R6159 gnd.n2936 gnd.n2754 585
R6160 gnd.n2754 gnd.n2753 585
R6161 gnd.n2938 gnd.n2937 585
R6162 gnd.n2939 gnd.n2938 585
R6163 gnd.n2752 gnd.n2751 585
R6164 gnd.n2940 gnd.n2752 585
R6165 gnd.n2943 gnd.n2942 585
R6166 gnd.n2942 gnd.n2941 585
R6167 gnd.n2944 gnd.n2746 585
R6168 gnd.n2746 gnd.n2745 585
R6169 gnd.n2946 gnd.n2945 585
R6170 gnd.n2947 gnd.n2946 585
R6171 gnd.n2744 gnd.n2743 585
R6172 gnd.n2948 gnd.n2744 585
R6173 gnd.n2951 gnd.n2950 585
R6174 gnd.n2950 gnd.n2949 585
R6175 gnd.n2952 gnd.n2738 585
R6176 gnd.n2738 gnd.n2737 585
R6177 gnd.n2954 gnd.n2953 585
R6178 gnd.n2955 gnd.n2954 585
R6179 gnd.n2736 gnd.n2735 585
R6180 gnd.n2956 gnd.n2736 585
R6181 gnd.n2959 gnd.n2958 585
R6182 gnd.n2958 gnd.n2957 585
R6183 gnd.n2960 gnd.n2730 585
R6184 gnd.n2730 gnd.n2729 585
R6185 gnd.n2962 gnd.n2961 585
R6186 gnd.n2963 gnd.n2962 585
R6187 gnd.n2728 gnd.n2727 585
R6188 gnd.n2964 gnd.n2728 585
R6189 gnd.n2967 gnd.n2966 585
R6190 gnd.n2966 gnd.n2965 585
R6191 gnd.n2968 gnd.n2722 585
R6192 gnd.n2722 gnd.n2721 585
R6193 gnd.n2970 gnd.n2969 585
R6194 gnd.n2971 gnd.n2970 585
R6195 gnd.n2720 gnd.n2719 585
R6196 gnd.n2972 gnd.n2720 585
R6197 gnd.n2975 gnd.n2974 585
R6198 gnd.n2974 gnd.n2973 585
R6199 gnd.n2976 gnd.n2714 585
R6200 gnd.n2714 gnd.n2713 585
R6201 gnd.n2978 gnd.n2977 585
R6202 gnd.n2979 gnd.n2978 585
R6203 gnd.n2712 gnd.n2711 585
R6204 gnd.n2980 gnd.n2712 585
R6205 gnd.n2983 gnd.n2982 585
R6206 gnd.n2982 gnd.n2981 585
R6207 gnd.n2984 gnd.n2706 585
R6208 gnd.n2706 gnd.n2705 585
R6209 gnd.n2986 gnd.n2985 585
R6210 gnd.n2987 gnd.n2986 585
R6211 gnd.n2704 gnd.n2703 585
R6212 gnd.n2988 gnd.n2704 585
R6213 gnd.n2991 gnd.n2990 585
R6214 gnd.n2990 gnd.n2989 585
R6215 gnd.n2992 gnd.n2698 585
R6216 gnd.n2698 gnd.n2697 585
R6217 gnd.n2994 gnd.n2993 585
R6218 gnd.n2995 gnd.n2994 585
R6219 gnd.n2696 gnd.n2695 585
R6220 gnd.n2996 gnd.n2696 585
R6221 gnd.n2999 gnd.n2998 585
R6222 gnd.n2998 gnd.n2997 585
R6223 gnd.n3000 gnd.n2690 585
R6224 gnd.n2690 gnd.n2689 585
R6225 gnd.n3002 gnd.n3001 585
R6226 gnd.n3003 gnd.n3002 585
R6227 gnd.n2688 gnd.n2687 585
R6228 gnd.n3004 gnd.n2688 585
R6229 gnd.n3007 gnd.n3006 585
R6230 gnd.n3006 gnd.n3005 585
R6231 gnd.n3008 gnd.n2682 585
R6232 gnd.n2682 gnd.n2681 585
R6233 gnd.n3010 gnd.n3009 585
R6234 gnd.n3011 gnd.n3010 585
R6235 gnd.n2680 gnd.n2679 585
R6236 gnd.n3012 gnd.n2680 585
R6237 gnd.n3015 gnd.n3014 585
R6238 gnd.n3014 gnd.n3013 585
R6239 gnd.n3016 gnd.n2674 585
R6240 gnd.n2674 gnd.n2673 585
R6241 gnd.n3018 gnd.n3017 585
R6242 gnd.n3019 gnd.n3018 585
R6243 gnd.n2672 gnd.n2671 585
R6244 gnd.n3020 gnd.n2672 585
R6245 gnd.n3023 gnd.n3022 585
R6246 gnd.n3022 gnd.n3021 585
R6247 gnd.n3024 gnd.n2667 585
R6248 gnd.n2667 gnd.n2666 585
R6249 gnd.n3026 gnd.n3025 585
R6250 gnd.n3027 gnd.n3026 585
R6251 gnd.n2665 gnd.n2664 585
R6252 gnd.n3028 gnd.n2665 585
R6253 gnd.n3031 gnd.n3030 585
R6254 gnd.n3030 gnd.n3029 585
R6255 gnd.n5900 gnd.n1604 585
R6256 gnd.n5958 gnd.n1604 585
R6257 gnd.n5901 gnd.n1615 585
R6258 gnd.n5728 gnd.n1615 585
R6259 gnd.n5903 gnd.n5902 585
R6260 gnd.n5904 gnd.n5903 585
R6261 gnd.n1616 gnd.n1614 585
R6262 gnd.n5559 gnd.n1614 585
R6263 gnd.n5709 gnd.n1763 585
R6264 gnd.n5721 gnd.n1763 585
R6265 gnd.n5710 gnd.n1774 585
R6266 gnd.n5563 gnd.n1774 585
R6267 gnd.n5712 gnd.n5711 585
R6268 gnd.n5713 gnd.n5712 585
R6269 gnd.n1775 gnd.n1773 585
R6270 gnd.n5569 gnd.n1773 585
R6271 gnd.n5702 gnd.n5701 585
R6272 gnd.n5701 gnd.n5700 585
R6273 gnd.n1778 gnd.n1777 585
R6274 gnd.n5497 gnd.n1778 585
R6275 gnd.n5691 gnd.n5690 585
R6276 gnd.n5692 gnd.n5691 585
R6277 gnd.n1793 gnd.n1792 585
R6278 gnd.n5501 gnd.n1792 585
R6279 gnd.n5686 gnd.n5685 585
R6280 gnd.n5685 gnd.n5684 585
R6281 gnd.n1796 gnd.n1795 585
R6282 gnd.n5505 gnd.n1796 585
R6283 gnd.n5675 gnd.n5674 585
R6284 gnd.n5676 gnd.n5675 585
R6285 gnd.n1810 gnd.n1809 585
R6286 gnd.n5511 gnd.n1809 585
R6287 gnd.n5670 gnd.n5669 585
R6288 gnd.n5669 gnd.n5668 585
R6289 gnd.n1813 gnd.n1812 585
R6290 gnd.n5484 gnd.n1813 585
R6291 gnd.n5659 gnd.n5658 585
R6292 gnd.n5660 gnd.n5659 585
R6293 gnd.n1828 gnd.n1827 585
R6294 gnd.n5480 gnd.n1827 585
R6295 gnd.n5654 gnd.n5653 585
R6296 gnd.n5653 gnd.n5652 585
R6297 gnd.n1831 gnd.n1830 585
R6298 gnd.n5596 gnd.n1831 585
R6299 gnd.n5617 gnd.n5616 585
R6300 gnd.n5618 gnd.n5617 585
R6301 gnd.n1885 gnd.n1879 585
R6302 gnd.n5623 gnd.n1879 585
R6303 gnd.n5612 gnd.n5611 585
R6304 gnd.n5611 gnd.n1875 585
R6305 gnd.n5610 gnd.n5609 585
R6306 gnd.n5610 gnd.n1868 585
R6307 gnd.n1858 gnd.n1857 585
R6308 gnd.n5632 gnd.n1858 585
R6309 gnd.n5639 gnd.n5638 585
R6310 gnd.n5638 gnd.n5637 585
R6311 gnd.n5640 gnd.n1852 585
R6312 gnd.n5405 gnd.n1852 585
R6313 gnd.n5642 gnd.n5641 585
R6314 gnd.n5643 gnd.n5642 585
R6315 gnd.n1853 gnd.n1851 585
R6316 gnd.n5397 gnd.n1851 585
R6317 gnd.n1936 gnd.n1935 585
R6318 gnd.n1935 gnd.n1934 585
R6319 gnd.n1937 gnd.n1913 585
R6320 gnd.n5388 gnd.n1913 585
R6321 gnd.n5375 gnd.n5374 585
R6322 gnd.n5374 gnd.n5373 585
R6323 gnd.n5376 gnd.n1926 585
R6324 gnd.n5356 gnd.n1926 585
R6325 gnd.n5378 gnd.n5377 585
R6326 gnd.n5379 gnd.n5378 585
R6327 gnd.n1927 gnd.n1925 585
R6328 gnd.n5362 gnd.n1925 585
R6329 gnd.n5333 gnd.n5332 585
R6330 gnd.n5332 gnd.n5331 585
R6331 gnd.n5334 gnd.n1953 585
R6332 gnd.n5348 gnd.n1953 585
R6333 gnd.n5335 gnd.n1965 585
R6334 gnd.n2206 gnd.n1965 585
R6335 gnd.n5337 gnd.n5336 585
R6336 gnd.n5338 gnd.n5337 585
R6337 gnd.n1966 gnd.n1964 585
R6338 gnd.n2212 gnd.n1964 585
R6339 gnd.n5323 gnd.n5322 585
R6340 gnd.n5322 gnd.n5321 585
R6341 gnd.n1969 gnd.n1968 585
R6342 gnd.n5221 gnd.n1969 585
R6343 gnd.n5312 gnd.n5311 585
R6344 gnd.n5313 gnd.n5312 585
R6345 gnd.n1983 gnd.n1982 585
R6346 gnd.n5227 gnd.n1982 585
R6347 gnd.n5307 gnd.n5306 585
R6348 gnd.n5306 gnd.n5305 585
R6349 gnd.n1986 gnd.n1985 585
R6350 gnd.n1987 gnd.n1986 585
R6351 gnd.n5296 gnd.n5295 585
R6352 gnd.n5297 gnd.n5296 585
R6353 gnd.n2001 gnd.n2000 585
R6354 gnd.n2000 gnd.n1996 585
R6355 gnd.n5291 gnd.n5290 585
R6356 gnd.n5290 gnd.n5289 585
R6357 gnd.n2004 gnd.n2003 585
R6358 gnd.n2005 gnd.n2004 585
R6359 gnd.n5280 gnd.n5279 585
R6360 gnd.n5281 gnd.n5280 585
R6361 gnd.n5276 gnd.n2015 585
R6362 gnd.n5275 gnd.n5274 585
R6363 gnd.n5272 gnd.n2017 585
R6364 gnd.n5270 gnd.n5269 585
R6365 gnd.n5268 gnd.n2018 585
R6366 gnd.n5267 gnd.n5266 585
R6367 gnd.n5264 gnd.n2023 585
R6368 gnd.n5262 gnd.n5261 585
R6369 gnd.n5260 gnd.n2024 585
R6370 gnd.n5259 gnd.n5258 585
R6371 gnd.n5256 gnd.n2029 585
R6372 gnd.n5254 gnd.n5253 585
R6373 gnd.n5252 gnd.n2030 585
R6374 gnd.n5251 gnd.n5250 585
R6375 gnd.n5248 gnd.n2035 585
R6376 gnd.n5246 gnd.n5245 585
R6377 gnd.n2037 gnd.n2036 585
R6378 gnd.n2036 gnd.n2012 585
R6379 gnd.n5769 gnd.n5768 585
R6380 gnd.n5770 gnd.n1747 585
R6381 gnd.n1746 gnd.n1737 585
R6382 gnd.n5777 gnd.n1736 585
R6383 gnd.n5778 gnd.n1735 585
R6384 gnd.n1733 gnd.n1725 585
R6385 gnd.n5785 gnd.n1724 585
R6386 gnd.n5786 gnd.n1722 585
R6387 gnd.n1721 gnd.n1714 585
R6388 gnd.n5793 gnd.n1713 585
R6389 gnd.n5794 gnd.n1712 585
R6390 gnd.n1710 gnd.n1703 585
R6391 gnd.n5801 gnd.n1702 585
R6392 gnd.n5802 gnd.n1700 585
R6393 gnd.n1699 gnd.n1694 585
R6394 gnd.n1697 gnd.n1696 585
R6395 gnd.n1695 gnd.n1619 585
R6396 gnd.n1695 gnd.n1567 585
R6397 gnd.n5731 gnd.n1602 585
R6398 gnd.n5958 gnd.n1602 585
R6399 gnd.n5730 gnd.n5729 585
R6400 gnd.n5729 gnd.n5728 585
R6401 gnd.n5727 gnd.n1612 585
R6402 gnd.n5904 gnd.n1612 585
R6403 gnd.n1759 gnd.n1755 585
R6404 gnd.n5559 gnd.n1759 585
R6405 gnd.n5723 gnd.n5722 585
R6406 gnd.n5722 gnd.n5721 585
R6407 gnd.n1758 gnd.n1757 585
R6408 gnd.n5563 gnd.n1758 585
R6409 gnd.n5571 gnd.n1771 585
R6410 gnd.n5713 gnd.n1771 585
R6411 gnd.n5572 gnd.n5570 585
R6412 gnd.n5570 gnd.n5569 585
R6413 gnd.n5430 gnd.n1781 585
R6414 gnd.n5700 gnd.n1781 585
R6415 gnd.n5576 gnd.n5429 585
R6416 gnd.n5497 gnd.n5429 585
R6417 gnd.n5577 gnd.n1790 585
R6418 gnd.n5692 gnd.n1790 585
R6419 gnd.n5578 gnd.n5428 585
R6420 gnd.n5501 gnd.n5428 585
R6421 gnd.n5426 gnd.n1799 585
R6422 gnd.n5684 gnd.n1799 585
R6423 gnd.n5582 gnd.n5425 585
R6424 gnd.n5505 gnd.n5425 585
R6425 gnd.n5583 gnd.n1807 585
R6426 gnd.n5676 gnd.n1807 585
R6427 gnd.n5584 gnd.n5424 585
R6428 gnd.n5511 gnd.n5424 585
R6429 gnd.n5422 gnd.n1816 585
R6430 gnd.n5668 gnd.n1816 585
R6431 gnd.n5588 gnd.n5421 585
R6432 gnd.n5484 gnd.n5421 585
R6433 gnd.n5589 gnd.n1825 585
R6434 gnd.n5660 gnd.n1825 585
R6435 gnd.n5590 gnd.n5420 585
R6436 gnd.n5480 gnd.n5420 585
R6437 gnd.n1895 gnd.n1834 585
R6438 gnd.n5652 gnd.n1834 585
R6439 gnd.n5595 gnd.n5594 585
R6440 gnd.n5596 gnd.n5595 585
R6441 gnd.n1894 gnd.n1883 585
R6442 gnd.n5618 gnd.n1883 585
R6443 gnd.n5416 gnd.n1877 585
R6444 gnd.n5623 gnd.n1877 585
R6445 gnd.n5415 gnd.n5414 585
R6446 gnd.n5414 gnd.n1875 585
R6447 gnd.n5413 gnd.n5412 585
R6448 gnd.n5413 gnd.n1868 585
R6449 gnd.n1897 gnd.n1867 585
R6450 gnd.n5632 gnd.n1867 585
R6451 gnd.n5408 gnd.n1861 585
R6452 gnd.n5637 gnd.n1861 585
R6453 gnd.n5407 gnd.n5406 585
R6454 gnd.n5406 gnd.n5405 585
R6455 gnd.n1899 gnd.n1849 585
R6456 gnd.n5643 gnd.n1849 585
R6457 gnd.n5396 gnd.n5395 585
R6458 gnd.n5397 gnd.n5396 585
R6459 gnd.n1906 gnd.n1905 585
R6460 gnd.n1934 gnd.n1905 585
R6461 gnd.n5390 gnd.n5389 585
R6462 gnd.n5389 gnd.n5388 585
R6463 gnd.n1909 gnd.n1908 585
R6464 gnd.n5373 gnd.n1909 585
R6465 gnd.n5358 gnd.n5357 585
R6466 gnd.n5357 gnd.n5356 585
R6467 gnd.n5359 gnd.n1923 585
R6468 gnd.n5379 gnd.n1923 585
R6469 gnd.n5361 gnd.n5360 585
R6470 gnd.n5362 gnd.n5361 585
R6471 gnd.n1946 gnd.n1945 585
R6472 gnd.n5331 gnd.n1945 585
R6473 gnd.n5350 gnd.n5349 585
R6474 gnd.n5349 gnd.n5348 585
R6475 gnd.n1949 gnd.n1948 585
R6476 gnd.n2206 gnd.n1949 585
R6477 gnd.n2198 gnd.n1962 585
R6478 gnd.n5338 gnd.n1962 585
R6479 gnd.n2214 gnd.n2213 585
R6480 gnd.n2213 gnd.n2212 585
R6481 gnd.n2215 gnd.n1971 585
R6482 gnd.n5321 gnd.n1971 585
R6483 gnd.n2217 gnd.n2216 585
R6484 gnd.n5221 gnd.n2217 585
R6485 gnd.n2046 gnd.n1980 585
R6486 gnd.n5313 gnd.n1980 585
R6487 gnd.n5229 gnd.n5228 585
R6488 gnd.n5228 gnd.n5227 585
R6489 gnd.n5230 gnd.n1989 585
R6490 gnd.n5305 gnd.n1989 585
R6491 gnd.n5232 gnd.n5231 585
R6492 gnd.n5231 gnd.n1987 585
R6493 gnd.n5233 gnd.n1998 585
R6494 gnd.n5297 gnd.n1998 585
R6495 gnd.n5235 gnd.n5234 585
R6496 gnd.n5234 gnd.n1996 585
R6497 gnd.n5236 gnd.n2007 585
R6498 gnd.n5289 gnd.n2007 585
R6499 gnd.n5238 gnd.n5237 585
R6500 gnd.n5237 gnd.n2005 585
R6501 gnd.n5239 gnd.n2014 585
R6502 gnd.n5281 gnd.n2014 585
R6503 gnd.n7267 gnd.n503 585
R6504 gnd.n7353 gnd.n503 585
R6505 gnd.n7268 gnd.n7205 585
R6506 gnd.n7205 gnd.n500 585
R6507 gnd.n7269 gnd.n577 585
R6508 gnd.n7283 gnd.n577 585
R6509 gnd.n589 gnd.n587 585
R6510 gnd.n587 gnd.n585 585
R6511 gnd.n7274 gnd.n7273 585
R6512 gnd.n7275 gnd.n7274 585
R6513 gnd.n588 gnd.n586 585
R6514 gnd.n596 gnd.n586 585
R6515 gnd.n7201 gnd.n7200 585
R6516 gnd.n7200 gnd.n7199 585
R6517 gnd.n592 gnd.n591 585
R6518 gnd.n2882 gnd.n592 585
R6519 gnd.n7190 gnd.n7189 585
R6520 gnd.n7191 gnd.n7190 585
R6521 gnd.n606 gnd.n605 585
R6522 gnd.n2888 gnd.n605 585
R6523 gnd.n7185 gnd.n7184 585
R6524 gnd.n7184 gnd.n7183 585
R6525 gnd.n609 gnd.n608 585
R6526 gnd.n2864 gnd.n609 585
R6527 gnd.n7174 gnd.n7173 585
R6528 gnd.n7175 gnd.n7174 585
R6529 gnd.n622 gnd.n621 585
R6530 gnd.n2860 gnd.n621 585
R6531 gnd.n7169 gnd.n7168 585
R6532 gnd.n7168 gnd.n7167 585
R6533 gnd.n625 gnd.n624 585
R6534 gnd.n2854 gnd.n625 585
R6535 gnd.n7158 gnd.n7157 585
R6536 gnd.n7159 gnd.n7158 585
R6537 gnd.n639 gnd.n638 585
R6538 gnd.n2850 gnd.n638 585
R6539 gnd.n7153 gnd.n7152 585
R6540 gnd.n7152 gnd.n7151 585
R6541 gnd.n642 gnd.n641 585
R6542 gnd.n2844 gnd.n642 585
R6543 gnd.n7142 gnd.n7141 585
R6544 gnd.n7143 gnd.n7142 585
R6545 gnd.n656 gnd.n655 585
R6546 gnd.n2840 gnd.n655 585
R6547 gnd.n7137 gnd.n7136 585
R6548 gnd.n7136 gnd.n7135 585
R6549 gnd.n659 gnd.n658 585
R6550 gnd.n6844 gnd.n659 585
R6551 gnd.n7127 gnd.n7126 585
R6552 gnd.n7128 gnd.n7127 585
R6553 gnd.n670 gnd.n669 585
R6554 gnd.n6848 gnd.n669 585
R6555 gnd.n7122 gnd.n7121 585
R6556 gnd.n7121 gnd.n7120 585
R6557 gnd.n674 gnd.n673 585
R6558 gnd.n6854 gnd.n674 585
R6559 gnd.n7111 gnd.n7110 585
R6560 gnd.n7112 gnd.n7111 585
R6561 gnd.n687 gnd.n686 585
R6562 gnd.n6793 gnd.n686 585
R6563 gnd.n7106 gnd.n7105 585
R6564 gnd.n7105 gnd.n7104 585
R6565 gnd.n690 gnd.n689 585
R6566 gnd.n6797 gnd.n690 585
R6567 gnd.n7095 gnd.n7094 585
R6568 gnd.n7096 gnd.n7095 585
R6569 gnd.n704 gnd.n703 585
R6570 gnd.n6801 gnd.n703 585
R6571 gnd.n7090 gnd.n7089 585
R6572 gnd.n7089 gnd.n7088 585
R6573 gnd.n707 gnd.n706 585
R6574 gnd.n6805 gnd.n707 585
R6575 gnd.n7078 gnd.n7077 585
R6576 gnd.n7079 gnd.n7078 585
R6577 gnd.n722 gnd.n721 585
R6578 gnd.n6811 gnd.n721 585
R6579 gnd.n7073 gnd.n7072 585
R6580 gnd.n7072 gnd.n7071 585
R6581 gnd.n725 gnd.n724 585
R6582 gnd.n6778 gnd.n725 585
R6583 gnd.n7062 gnd.n7061 585
R6584 gnd.n7063 gnd.n7062 585
R6585 gnd.n739 gnd.n738 585
R6586 gnd.n6774 gnd.n738 585
R6587 gnd.n7057 gnd.n7056 585
R6588 gnd.n7056 gnd.n7055 585
R6589 gnd.n742 gnd.n741 585
R6590 gnd.n6768 gnd.n742 585
R6591 gnd.n7046 gnd.n7045 585
R6592 gnd.n7047 gnd.n7046 585
R6593 gnd.n757 gnd.n756 585
R6594 gnd.n6764 gnd.n756 585
R6595 gnd.n7041 gnd.n7040 585
R6596 gnd.n7040 gnd.n7039 585
R6597 gnd.n760 gnd.n759 585
R6598 gnd.n6758 gnd.n760 585
R6599 gnd.n7030 gnd.n7029 585
R6600 gnd.n7031 gnd.n7030 585
R6601 gnd.n775 gnd.n774 585
R6602 gnd.n6892 gnd.n774 585
R6603 gnd.n7025 gnd.n7024 585
R6604 gnd.n7024 gnd.n7023 585
R6605 gnd.n778 gnd.n777 585
R6606 gnd.n1013 gnd.n778 585
R6607 gnd.n7014 gnd.n7013 585
R6608 gnd.n7015 gnd.n7014 585
R6609 gnd.n7010 gnd.n790 585
R6610 gnd.n7009 gnd.n792 585
R6611 gnd.n851 gnd.n793 585
R6612 gnd.n7002 gnd.n799 585
R6613 gnd.n7001 gnd.n800 585
R6614 gnd.n853 gnd.n801 585
R6615 gnd.n6994 gnd.n807 585
R6616 gnd.n6993 gnd.n808 585
R6617 gnd.n856 gnd.n809 585
R6618 gnd.n6986 gnd.n815 585
R6619 gnd.n6985 gnd.n816 585
R6620 gnd.n858 gnd.n817 585
R6621 gnd.n6978 gnd.n823 585
R6622 gnd.n6977 gnd.n824 585
R6623 gnd.n6965 gnd.n825 585
R6624 gnd.n6970 gnd.n6967 585
R6625 gnd.n832 gnd.n831 585
R6626 gnd.n6964 gnd.n832 585
R6627 gnd.n7240 gnd.n499 585
R6628 gnd.n7239 gnd.n7238 585
R6629 gnd.n7244 gnd.n7234 585
R6630 gnd.n7245 gnd.n7232 585
R6631 gnd.n7246 gnd.n7231 585
R6632 gnd.n7229 gnd.n7227 585
R6633 gnd.n7250 gnd.n7226 585
R6634 gnd.n7251 gnd.n7224 585
R6635 gnd.n7252 gnd.n7223 585
R6636 gnd.n7221 gnd.n7219 585
R6637 gnd.n7256 gnd.n7218 585
R6638 gnd.n7257 gnd.n7216 585
R6639 gnd.n7258 gnd.n7215 585
R6640 gnd.n7213 gnd.n7211 585
R6641 gnd.n7262 gnd.n7210 585
R6642 gnd.n7263 gnd.n7208 585
R6643 gnd.n7264 gnd.n7207 585
R6644 gnd.n7207 gnd.n502 585
R6645 gnd.n7355 gnd.n7354 585
R6646 gnd.n7354 gnd.n7353 585
R6647 gnd.n7356 gnd.n498 585
R6648 gnd.n500 gnd.n498 585
R6649 gnd.n576 gnd.n496 585
R6650 gnd.n7283 gnd.n576 585
R6651 gnd.n7360 gnd.n495 585
R6652 gnd.n585 gnd.n495 585
R6653 gnd.n7361 gnd.n494 585
R6654 gnd.n7275 gnd.n494 585
R6655 gnd.n7362 gnd.n493 585
R6656 gnd.n596 gnd.n493 585
R6657 gnd.n595 gnd.n491 585
R6658 gnd.n7199 gnd.n595 585
R6659 gnd.n7366 gnd.n490 585
R6660 gnd.n2882 gnd.n490 585
R6661 gnd.n7367 gnd.n489 585
R6662 gnd.n7191 gnd.n489 585
R6663 gnd.n7368 gnd.n488 585
R6664 gnd.n2888 gnd.n488 585
R6665 gnd.n612 gnd.n486 585
R6666 gnd.n7183 gnd.n612 585
R6667 gnd.n7372 gnd.n485 585
R6668 gnd.n2864 gnd.n485 585
R6669 gnd.n7373 gnd.n484 585
R6670 gnd.n7175 gnd.n484 585
R6671 gnd.n7374 gnd.n483 585
R6672 gnd.n2860 gnd.n483 585
R6673 gnd.n628 gnd.n481 585
R6674 gnd.n7167 gnd.n628 585
R6675 gnd.n7378 gnd.n480 585
R6676 gnd.n2854 gnd.n480 585
R6677 gnd.n7379 gnd.n479 585
R6678 gnd.n7159 gnd.n479 585
R6679 gnd.n7380 gnd.n478 585
R6680 gnd.n2850 gnd.n478 585
R6681 gnd.n645 gnd.n476 585
R6682 gnd.n7151 gnd.n645 585
R6683 gnd.n7384 gnd.n475 585
R6684 gnd.n2844 gnd.n475 585
R6685 gnd.n7385 gnd.n474 585
R6686 gnd.n7143 gnd.n474 585
R6687 gnd.n7386 gnd.n473 585
R6688 gnd.n2840 gnd.n473 585
R6689 gnd.n662 gnd.n471 585
R6690 gnd.n7135 gnd.n662 585
R6691 gnd.n7390 gnd.n470 585
R6692 gnd.n6844 gnd.n470 585
R6693 gnd.n7391 gnd.n469 585
R6694 gnd.n7128 gnd.n469 585
R6695 gnd.n7392 gnd.n468 585
R6696 gnd.n6848 gnd.n468 585
R6697 gnd.n677 gnd.n466 585
R6698 gnd.n7120 gnd.n677 585
R6699 gnd.n6856 gnd.n6855 585
R6700 gnd.n6855 gnd.n6854 585
R6701 gnd.n6857 gnd.n684 585
R6702 gnd.n7112 gnd.n684 585
R6703 gnd.n6860 gnd.n930 585
R6704 gnd.n6793 gnd.n930 585
R6705 gnd.n6861 gnd.n693 585
R6706 gnd.n7104 gnd.n693 585
R6707 gnd.n6862 gnd.n929 585
R6708 gnd.n6797 gnd.n929 585
R6709 gnd.n927 gnd.n701 585
R6710 gnd.n7096 gnd.n701 585
R6711 gnd.n6866 gnd.n926 585
R6712 gnd.n6801 gnd.n926 585
R6713 gnd.n6867 gnd.n710 585
R6714 gnd.n7088 gnd.n710 585
R6715 gnd.n6868 gnd.n925 585
R6716 gnd.n6805 gnd.n925 585
R6717 gnd.n923 gnd.n719 585
R6718 gnd.n7079 gnd.n719 585
R6719 gnd.n6872 gnd.n922 585
R6720 gnd.n6811 gnd.n922 585
R6721 gnd.n6873 gnd.n728 585
R6722 gnd.n7071 gnd.n728 585
R6723 gnd.n6874 gnd.n921 585
R6724 gnd.n6778 gnd.n921 585
R6725 gnd.n919 gnd.n736 585
R6726 gnd.n7063 gnd.n736 585
R6727 gnd.n6878 gnd.n918 585
R6728 gnd.n6774 gnd.n918 585
R6729 gnd.n6879 gnd.n745 585
R6730 gnd.n7055 gnd.n745 585
R6731 gnd.n6880 gnd.n917 585
R6732 gnd.n6768 gnd.n917 585
R6733 gnd.n915 gnd.n754 585
R6734 gnd.n7047 gnd.n754 585
R6735 gnd.n6884 gnd.n914 585
R6736 gnd.n6764 gnd.n914 585
R6737 gnd.n6885 gnd.n763 585
R6738 gnd.n7039 gnd.n763 585
R6739 gnd.n6886 gnd.n913 585
R6740 gnd.n6758 gnd.n913 585
R6741 gnd.n910 gnd.n772 585
R6742 gnd.n7031 gnd.n772 585
R6743 gnd.n6891 gnd.n6890 585
R6744 gnd.n6892 gnd.n6891 585
R6745 gnd.n909 gnd.n781 585
R6746 gnd.n7023 gnd.n781 585
R6747 gnd.n1015 gnd.n1014 585
R6748 gnd.n1014 gnd.n1013 585
R6749 gnd.n1016 gnd.n788 585
R6750 gnd.n7015 gnd.n788 585
R6751 gnd.n5011 gnd.n5010 585
R6752 gnd.n5010 gnd.n3604 585
R6753 gnd.n3592 gnd.n3591 585
R6754 gnd.n5015 gnd.n3592 585
R6755 gnd.n5126 gnd.n5125 585
R6756 gnd.n5125 gnd.n5124 585
R6757 gnd.n5127 gnd.n3586 585
R6758 gnd.n5023 gnd.n3586 585
R6759 gnd.n5129 gnd.n5128 585
R6760 gnd.n5130 gnd.n5129 585
R6761 gnd.n3587 gnd.n3585 585
R6762 gnd.n3585 gnd.n3581 585
R6763 gnd.n3567 gnd.n3566 585
R6764 gnd.n4731 gnd.n3567 585
R6765 gnd.n5140 gnd.n5139 585
R6766 gnd.n5139 gnd.n5138 585
R6767 gnd.n5141 gnd.n3561 585
R6768 gnd.n4737 gnd.n3561 585
R6769 gnd.n5143 gnd.n5142 585
R6770 gnd.n5144 gnd.n5143 585
R6771 gnd.n3562 gnd.n3560 585
R6772 gnd.n3560 gnd.n3557 585
R6773 gnd.n3545 gnd.n3544 585
R6774 gnd.n4716 gnd.n3545 585
R6775 gnd.n5154 gnd.n5153 585
R6776 gnd.n5153 gnd.n5152 585
R6777 gnd.n5155 gnd.n3539 585
R6778 gnd.n4669 gnd.n3539 585
R6779 gnd.n5157 gnd.n5156 585
R6780 gnd.n5158 gnd.n5157 585
R6781 gnd.n3540 gnd.n3538 585
R6782 gnd.n3703 gnd.n3538 585
R6783 gnd.n4696 gnd.n4695 585
R6784 gnd.n4695 gnd.n4694 585
R6785 gnd.n3700 gnd.n3699 585
R6786 gnd.n4678 gnd.n3700 585
R6787 gnd.n4654 gnd.n3719 585
R6788 gnd.n3719 gnd.n3710 585
R6789 gnd.n4656 gnd.n4655 585
R6790 gnd.n4657 gnd.n4656 585
R6791 gnd.n3720 gnd.n3718 585
R6792 gnd.n3726 gnd.n3718 585
R6793 gnd.n4635 gnd.n4634 585
R6794 gnd.n4636 gnd.n4635 585
R6795 gnd.n3737 gnd.n3736 585
R6796 gnd.n3736 gnd.n3732 585
R6797 gnd.n4625 gnd.n4624 585
R6798 gnd.n4626 gnd.n4625 585
R6799 gnd.n3748 gnd.n3747 585
R6800 gnd.n3752 gnd.n3747 585
R6801 gnd.n4603 gnd.n3764 585
R6802 gnd.n4106 gnd.n3764 585
R6803 gnd.n4605 gnd.n4604 585
R6804 gnd.n4606 gnd.n4605 585
R6805 gnd.n3765 gnd.n3763 585
R6806 gnd.n3763 gnd.n3759 585
R6807 gnd.n4594 gnd.n4593 585
R6808 gnd.n4595 gnd.n4594 585
R6809 gnd.n3773 gnd.n3772 585
R6810 gnd.n4114 gnd.n3772 585
R6811 gnd.n4572 gnd.n3789 585
R6812 gnd.n3789 gnd.n3777 585
R6813 gnd.n4574 gnd.n4573 585
R6814 gnd.n4575 gnd.n4574 585
R6815 gnd.n3790 gnd.n3788 585
R6816 gnd.n3788 gnd.n3784 585
R6817 gnd.n4563 gnd.n4562 585
R6818 gnd.n4564 gnd.n4563 585
R6819 gnd.n3798 gnd.n3797 585
R6820 gnd.n3803 gnd.n3797 585
R6821 gnd.n4541 gnd.n3815 585
R6822 gnd.n3815 gnd.n3802 585
R6823 gnd.n4543 gnd.n4542 585
R6824 gnd.n4544 gnd.n4543 585
R6825 gnd.n3816 gnd.n3814 585
R6826 gnd.n3814 gnd.n3810 585
R6827 gnd.n4532 gnd.n4531 585
R6828 gnd.n4533 gnd.n4532 585
R6829 gnd.n3823 gnd.n3822 585
R6830 gnd.n3828 gnd.n3822 585
R6831 gnd.n4510 gnd.n3841 585
R6832 gnd.n3841 gnd.n3827 585
R6833 gnd.n4512 gnd.n4511 585
R6834 gnd.n4513 gnd.n4512 585
R6835 gnd.n3842 gnd.n3840 585
R6836 gnd.n3840 gnd.n3836 585
R6837 gnd.n4501 gnd.n4500 585
R6838 gnd.n4502 gnd.n4501 585
R6839 gnd.n3849 gnd.n3848 585
R6840 gnd.n3854 gnd.n3848 585
R6841 gnd.n4479 gnd.n3867 585
R6842 gnd.n3867 gnd.n3853 585
R6843 gnd.n4481 gnd.n4480 585
R6844 gnd.n4482 gnd.n4481 585
R6845 gnd.n3868 gnd.n3866 585
R6846 gnd.n3866 gnd.n3862 585
R6847 gnd.n4470 gnd.n4469 585
R6848 gnd.n4471 gnd.n4470 585
R6849 gnd.n3876 gnd.n3875 585
R6850 gnd.n4360 gnd.n3875 585
R6851 gnd.n4448 gnd.n3892 585
R6852 gnd.n3892 gnd.n3880 585
R6853 gnd.n4450 gnd.n4449 585
R6854 gnd.n4451 gnd.n4450 585
R6855 gnd.n3893 gnd.n3891 585
R6856 gnd.n3891 gnd.n3887 585
R6857 gnd.n4439 gnd.n4438 585
R6858 gnd.n4440 gnd.n4439 585
R6859 gnd.n3900 gnd.n3899 585
R6860 gnd.n3899 gnd.n3897 585
R6861 gnd.n4433 gnd.n4432 585
R6862 gnd.n4432 gnd.n4431 585
R6863 gnd.n3904 gnd.n3903 585
R6864 gnd.n3912 gnd.n3904 585
R6865 gnd.n4065 gnd.n4064 585
R6866 gnd.n4066 gnd.n4065 585
R6867 gnd.n3914 gnd.n3913 585
R6868 gnd.n3913 gnd.n3911 585
R6869 gnd.n4060 gnd.n4059 585
R6870 gnd.n4059 gnd.n4058 585
R6871 gnd.n3917 gnd.n3916 585
R6872 gnd.n3918 gnd.n3917 585
R6873 gnd.n4049 gnd.n4048 585
R6874 gnd.n4050 gnd.n4049 585
R6875 gnd.n3926 gnd.n3925 585
R6876 gnd.n3925 gnd.n3924 585
R6877 gnd.n4044 gnd.n4043 585
R6878 gnd.n4043 gnd.n4042 585
R6879 gnd.n3929 gnd.n3928 585
R6880 gnd.n3930 gnd.n3929 585
R6881 gnd.n4033 gnd.n4032 585
R6882 gnd.n4034 gnd.n4033 585
R6883 gnd.n4029 gnd.n3936 585
R6884 gnd.n4028 gnd.n4027 585
R6885 gnd.n4025 gnd.n3938 585
R6886 gnd.n4025 gnd.n3935 585
R6887 gnd.n4024 gnd.n4023 585
R6888 gnd.n4022 gnd.n4021 585
R6889 gnd.n4020 gnd.n3943 585
R6890 gnd.n4018 gnd.n4017 585
R6891 gnd.n4016 gnd.n3944 585
R6892 gnd.n4015 gnd.n4014 585
R6893 gnd.n4012 gnd.n3949 585
R6894 gnd.n4010 gnd.n4009 585
R6895 gnd.n4008 gnd.n3950 585
R6896 gnd.n4007 gnd.n4006 585
R6897 gnd.n4004 gnd.n3955 585
R6898 gnd.n4002 gnd.n4001 585
R6899 gnd.n4000 gnd.n3956 585
R6900 gnd.n3999 gnd.n3998 585
R6901 gnd.n3996 gnd.n3961 585
R6902 gnd.n3994 gnd.n3993 585
R6903 gnd.n3992 gnd.n3962 585
R6904 gnd.n3991 gnd.n3990 585
R6905 gnd.n3988 gnd.n3967 585
R6906 gnd.n3986 gnd.n3985 585
R6907 gnd.n3983 gnd.n3968 585
R6908 gnd.n3982 gnd.n3981 585
R6909 gnd.n3979 gnd.n3977 585
R6910 gnd.n3975 gnd.n3934 585
R6911 gnd.n5033 gnd.n5032 585
R6912 gnd.n5035 gnd.n5034 585
R6913 gnd.n5037 gnd.n5036 585
R6914 gnd.n5039 gnd.n5038 585
R6915 gnd.n5041 gnd.n5040 585
R6916 gnd.n5043 gnd.n5042 585
R6917 gnd.n5045 gnd.n5044 585
R6918 gnd.n5047 gnd.n5046 585
R6919 gnd.n5049 gnd.n5048 585
R6920 gnd.n5051 gnd.n5050 585
R6921 gnd.n5053 gnd.n5052 585
R6922 gnd.n5055 gnd.n5054 585
R6923 gnd.n5057 gnd.n5056 585
R6924 gnd.n5059 gnd.n5058 585
R6925 gnd.n5061 gnd.n5060 585
R6926 gnd.n5063 gnd.n5062 585
R6927 gnd.n5065 gnd.n5064 585
R6928 gnd.n5067 gnd.n5066 585
R6929 gnd.n5069 gnd.n5068 585
R6930 gnd.n5071 gnd.n5070 585
R6931 gnd.n5073 gnd.n5072 585
R6932 gnd.n5075 gnd.n5074 585
R6933 gnd.n5077 gnd.n5076 585
R6934 gnd.n5079 gnd.n5078 585
R6935 gnd.n5081 gnd.n5080 585
R6936 gnd.n5082 gnd.n3652 585
R6937 gnd.n5083 gnd.n3606 585
R6938 gnd.n5116 gnd.n3606 585
R6939 gnd.n5031 gnd.n5030 585
R6940 gnd.n5031 gnd.n3604 585
R6941 gnd.n3682 gnd.n3681 585
R6942 gnd.n5015 gnd.n3681 585
R6943 gnd.n5026 gnd.n3593 585
R6944 gnd.n5124 gnd.n3593 585
R6945 gnd.n5025 gnd.n5024 585
R6946 gnd.n5024 gnd.n5023 585
R6947 gnd.n3684 gnd.n3583 585
R6948 gnd.n5130 gnd.n3583 585
R6949 gnd.n4728 gnd.n4727 585
R6950 gnd.n4728 gnd.n3581 585
R6951 gnd.n4733 gnd.n4732 585
R6952 gnd.n4732 gnd.n4731 585
R6953 gnd.n4734 gnd.n3569 585
R6954 gnd.n5138 gnd.n3569 585
R6955 gnd.n4736 gnd.n4735 585
R6956 gnd.n4737 gnd.n4736 585
R6957 gnd.n3690 gnd.n3559 585
R6958 gnd.n5144 gnd.n3559 585
R6959 gnd.n4719 gnd.n4718 585
R6960 gnd.n4718 gnd.n3557 585
R6961 gnd.n4717 gnd.n3692 585
R6962 gnd.n4717 gnd.n4716 585
R6963 gnd.n4668 gnd.n3547 585
R6964 gnd.n5152 gnd.n3547 585
R6965 gnd.n4671 gnd.n4670 585
R6966 gnd.n4670 gnd.n4669 585
R6967 gnd.n4672 gnd.n3536 585
R6968 gnd.n5158 gnd.n3536 585
R6969 gnd.n4674 gnd.n4673 585
R6970 gnd.n4673 gnd.n3703 585
R6971 gnd.n4675 gnd.n3702 585
R6972 gnd.n4694 gnd.n3702 585
R6973 gnd.n4677 gnd.n4676 585
R6974 gnd.n4678 gnd.n4677 585
R6975 gnd.n3713 gnd.n3712 585
R6976 gnd.n3712 gnd.n3710 585
R6977 gnd.n4659 gnd.n4658 585
R6978 gnd.n4658 gnd.n4657 585
R6979 gnd.n3716 gnd.n3715 585
R6980 gnd.n3726 gnd.n3716 585
R6981 gnd.n4100 gnd.n3734 585
R6982 gnd.n4636 gnd.n3734 585
R6983 gnd.n4102 gnd.n4101 585
R6984 gnd.n4101 gnd.n3732 585
R6985 gnd.n4103 gnd.n3746 585
R6986 gnd.n4626 gnd.n3746 585
R6987 gnd.n4105 gnd.n4104 585
R6988 gnd.n4105 gnd.n3752 585
R6989 gnd.n4108 gnd.n4107 585
R6990 gnd.n4107 gnd.n4106 585
R6991 gnd.n4109 gnd.n3761 585
R6992 gnd.n4606 gnd.n3761 585
R6993 gnd.n4111 gnd.n4110 585
R6994 gnd.n4110 gnd.n3759 585
R6995 gnd.n4112 gnd.n3771 585
R6996 gnd.n4595 gnd.n3771 585
R6997 gnd.n4115 gnd.n4113 585
R6998 gnd.n4115 gnd.n4114 585
R6999 gnd.n4117 gnd.n4116 585
R7000 gnd.n4116 gnd.n3777 585
R7001 gnd.n4118 gnd.n3786 585
R7002 gnd.n4575 gnd.n3786 585
R7003 gnd.n4121 gnd.n4120 585
R7004 gnd.n4120 gnd.n3784 585
R7005 gnd.n4122 gnd.n3796 585
R7006 gnd.n4564 gnd.n3796 585
R7007 gnd.n4125 gnd.n4124 585
R7008 gnd.n4124 gnd.n3803 585
R7009 gnd.n4123 gnd.n4090 585
R7010 gnd.n4123 gnd.n3802 585
R7011 gnd.n4339 gnd.n3812 585
R7012 gnd.n4544 gnd.n3812 585
R7013 gnd.n4341 gnd.n4340 585
R7014 gnd.n4340 gnd.n3810 585
R7015 gnd.n4342 gnd.n3821 585
R7016 gnd.n4533 gnd.n3821 585
R7017 gnd.n4344 gnd.n4343 585
R7018 gnd.n4344 gnd.n3828 585
R7019 gnd.n4346 gnd.n4345 585
R7020 gnd.n4345 gnd.n3827 585
R7021 gnd.n4347 gnd.n3838 585
R7022 gnd.n4513 gnd.n3838 585
R7023 gnd.n4349 gnd.n4348 585
R7024 gnd.n4348 gnd.n3836 585
R7025 gnd.n4350 gnd.n3847 585
R7026 gnd.n4502 gnd.n3847 585
R7027 gnd.n4352 gnd.n4351 585
R7028 gnd.n4352 gnd.n3854 585
R7029 gnd.n4354 gnd.n4353 585
R7030 gnd.n4353 gnd.n3853 585
R7031 gnd.n4355 gnd.n3864 585
R7032 gnd.n4482 gnd.n3864 585
R7033 gnd.n4357 gnd.n4356 585
R7034 gnd.n4356 gnd.n3862 585
R7035 gnd.n4358 gnd.n3874 585
R7036 gnd.n4471 gnd.n3874 585
R7037 gnd.n4361 gnd.n4359 585
R7038 gnd.n4361 gnd.n4360 585
R7039 gnd.n4363 gnd.n4362 585
R7040 gnd.n4362 gnd.n3880 585
R7041 gnd.n4364 gnd.n3889 585
R7042 gnd.n4451 gnd.n3889 585
R7043 gnd.n4366 gnd.n4365 585
R7044 gnd.n4365 gnd.n3887 585
R7045 gnd.n4367 gnd.n3898 585
R7046 gnd.n4440 gnd.n3898 585
R7047 gnd.n4368 gnd.n3906 585
R7048 gnd.n3906 gnd.n3897 585
R7049 gnd.n4370 gnd.n4369 585
R7050 gnd.n4431 gnd.n4370 585
R7051 gnd.n3907 gnd.n3905 585
R7052 gnd.n3912 gnd.n3905 585
R7053 gnd.n4068 gnd.n4067 585
R7054 gnd.n4067 gnd.n4066 585
R7055 gnd.n3910 gnd.n3909 585
R7056 gnd.n3911 gnd.n3910 585
R7057 gnd.n4057 gnd.n4056 585
R7058 gnd.n4058 gnd.n4057 585
R7059 gnd.n3920 gnd.n3919 585
R7060 gnd.n3919 gnd.n3918 585
R7061 gnd.n4052 gnd.n4051 585
R7062 gnd.n4051 gnd.n4050 585
R7063 gnd.n3923 gnd.n3922 585
R7064 gnd.n3924 gnd.n3923 585
R7065 gnd.n4041 gnd.n4040 585
R7066 gnd.n4042 gnd.n4041 585
R7067 gnd.n3932 gnd.n3931 585
R7068 gnd.n3931 gnd.n3930 585
R7069 gnd.n4036 gnd.n4035 585
R7070 gnd.n4035 gnd.n4034 585
R7071 gnd.n5119 gnd.n5118 585
R7072 gnd.n5118 gnd.n5117 585
R7073 gnd.n5120 gnd.n3596 585
R7074 gnd.n5016 gnd.n3596 585
R7075 gnd.n5122 gnd.n5121 585
R7076 gnd.n5123 gnd.n5122 585
R7077 gnd.n3597 gnd.n3595 585
R7078 gnd.n5022 gnd.n3595 585
R7079 gnd.n3580 gnd.n3579 585
R7080 gnd.n3584 gnd.n3580 585
R7081 gnd.n5133 gnd.n5132 585
R7082 gnd.n5132 gnd.n5131 585
R7083 gnd.n5134 gnd.n3572 585
R7084 gnd.n4730 gnd.n3572 585
R7085 gnd.n5136 gnd.n5135 585
R7086 gnd.n5137 gnd.n5136 585
R7087 gnd.n3573 gnd.n3571 585
R7088 gnd.n3571 gnd.n3568 585
R7089 gnd.n3556 gnd.n3555 585
R7090 gnd.n4738 gnd.n3556 585
R7091 gnd.n5147 gnd.n5146 585
R7092 gnd.n5146 gnd.n5145 585
R7093 gnd.n5148 gnd.n3550 585
R7094 gnd.n4715 gnd.n3550 585
R7095 gnd.n5150 gnd.n5149 585
R7096 gnd.n5151 gnd.n5150 585
R7097 gnd.n3551 gnd.n3549 585
R7098 gnd.n3549 gnd.n3546 585
R7099 gnd.n4689 gnd.n4688 585
R7100 gnd.n4688 gnd.n3537 585
R7101 gnd.n4690 gnd.n3705 585
R7102 gnd.n3705 gnd.n3535 585
R7103 gnd.n4692 gnd.n4691 585
R7104 gnd.n4693 gnd.n4692 585
R7105 gnd.n3706 gnd.n3704 585
R7106 gnd.n3704 gnd.n3701 585
R7107 gnd.n4681 gnd.n4680 585
R7108 gnd.n4680 gnd.n4679 585
R7109 gnd.n3709 gnd.n3708 585
R7110 gnd.n3717 gnd.n3709 585
R7111 gnd.n4644 gnd.n4643 585
R7112 gnd.n4645 gnd.n4644 585
R7113 gnd.n3728 gnd.n3727 585
R7114 gnd.n3735 gnd.n3727 585
R7115 gnd.n4639 gnd.n4638 585
R7116 gnd.n4638 gnd.n4637 585
R7117 gnd.n3731 gnd.n3730 585
R7118 gnd.n4627 gnd.n3731 585
R7119 gnd.n4614 gnd.n3754 585
R7120 gnd.n3754 gnd.n3745 585
R7121 gnd.n4616 gnd.n4615 585
R7122 gnd.n4617 gnd.n4616 585
R7123 gnd.n3755 gnd.n3753 585
R7124 gnd.n3762 gnd.n3753 585
R7125 gnd.n4609 gnd.n4608 585
R7126 gnd.n4608 gnd.n4607 585
R7127 gnd.n3758 gnd.n3757 585
R7128 gnd.n4596 gnd.n3758 585
R7129 gnd.n4583 gnd.n3779 585
R7130 gnd.n3779 gnd.n3770 585
R7131 gnd.n4585 gnd.n4584 585
R7132 gnd.n4586 gnd.n4585 585
R7133 gnd.n3780 gnd.n3778 585
R7134 gnd.n3787 gnd.n3778 585
R7135 gnd.n4578 gnd.n4577 585
R7136 gnd.n4577 gnd.n4576 585
R7137 gnd.n3783 gnd.n3782 585
R7138 gnd.n4565 gnd.n3783 585
R7139 gnd.n4552 gnd.n3805 585
R7140 gnd.n3805 gnd.n3795 585
R7141 gnd.n4554 gnd.n4553 585
R7142 gnd.n4555 gnd.n4554 585
R7143 gnd.n3806 gnd.n3804 585
R7144 gnd.n3813 gnd.n3804 585
R7145 gnd.n4547 gnd.n4546 585
R7146 gnd.n4546 gnd.n4545 585
R7147 gnd.n3809 gnd.n3808 585
R7148 gnd.n4534 gnd.n3809 585
R7149 gnd.n4521 gnd.n3831 585
R7150 gnd.n3831 gnd.n3830 585
R7151 gnd.n4523 gnd.n4522 585
R7152 gnd.n4524 gnd.n4523 585
R7153 gnd.n3832 gnd.n3829 585
R7154 gnd.n3839 gnd.n3829 585
R7155 gnd.n4516 gnd.n4515 585
R7156 gnd.n4515 gnd.n4514 585
R7157 gnd.n3835 gnd.n3834 585
R7158 gnd.n4503 gnd.n3835 585
R7159 gnd.n4490 gnd.n3857 585
R7160 gnd.n3857 gnd.n3856 585
R7161 gnd.n4492 gnd.n4491 585
R7162 gnd.n4493 gnd.n4492 585
R7163 gnd.n3858 gnd.n3855 585
R7164 gnd.n3865 gnd.n3855 585
R7165 gnd.n4485 gnd.n4484 585
R7166 gnd.n4484 gnd.n4483 585
R7167 gnd.n3861 gnd.n3860 585
R7168 gnd.n4472 gnd.n3861 585
R7169 gnd.n4459 gnd.n3882 585
R7170 gnd.n3882 gnd.n3873 585
R7171 gnd.n4461 gnd.n4460 585
R7172 gnd.n4462 gnd.n4461 585
R7173 gnd.n3883 gnd.n3881 585
R7174 gnd.n3890 gnd.n3881 585
R7175 gnd.n4454 gnd.n4453 585
R7176 gnd.n4453 gnd.n4452 585
R7177 gnd.n3886 gnd.n3885 585
R7178 gnd.n4441 gnd.n3886 585
R7179 gnd.n4428 gnd.n4427 585
R7180 gnd.n4426 gnd.n4379 585
R7181 gnd.n4425 gnd.n4378 585
R7182 gnd.n4430 gnd.n4378 585
R7183 gnd.n4424 gnd.n4423 585
R7184 gnd.n4422 gnd.n4421 585
R7185 gnd.n4420 gnd.n4419 585
R7186 gnd.n4418 gnd.n4417 585
R7187 gnd.n4416 gnd.n4415 585
R7188 gnd.n4414 gnd.n4413 585
R7189 gnd.n4412 gnd.n4411 585
R7190 gnd.n4410 gnd.n4409 585
R7191 gnd.n4408 gnd.n4407 585
R7192 gnd.n4406 gnd.n4405 585
R7193 gnd.n4404 gnd.n4403 585
R7194 gnd.n4402 gnd.n4401 585
R7195 gnd.n4400 gnd.n4399 585
R7196 gnd.n4395 gnd.n3896 585
R7197 gnd.n3647 gnd.n3646 585
R7198 gnd.n5089 gnd.n5088 585
R7199 gnd.n5091 gnd.n5090 585
R7200 gnd.n5093 gnd.n5092 585
R7201 gnd.n5095 gnd.n5094 585
R7202 gnd.n5097 gnd.n5096 585
R7203 gnd.n5099 gnd.n5098 585
R7204 gnd.n5101 gnd.n5100 585
R7205 gnd.n5103 gnd.n5102 585
R7206 gnd.n5105 gnd.n5104 585
R7207 gnd.n5107 gnd.n5106 585
R7208 gnd.n5109 gnd.n5108 585
R7209 gnd.n5111 gnd.n5110 585
R7210 gnd.n5112 gnd.n3628 585
R7211 gnd.n5114 gnd.n5113 585
R7212 gnd.n3629 gnd.n3627 585
R7213 gnd.n3630 gnd.n3603 585
R7214 gnd.n5116 gnd.n3603 585
R7215 gnd.n5014 gnd.n3605 585
R7216 gnd.n5117 gnd.n3605 585
R7217 gnd.n5018 gnd.n5017 585
R7218 gnd.n5017 gnd.n5016 585
R7219 gnd.n5019 gnd.n3594 585
R7220 gnd.n5123 gnd.n3594 585
R7221 gnd.n5021 gnd.n5020 585
R7222 gnd.n5022 gnd.n5021 585
R7223 gnd.n5006 gnd.n3685 585
R7224 gnd.n3685 gnd.n3584 585
R7225 gnd.n5004 gnd.n3582 585
R7226 gnd.n5131 gnd.n3582 585
R7227 gnd.n4729 gnd.n3686 585
R7228 gnd.n4730 gnd.n4729 585
R7229 gnd.n4742 gnd.n3570 585
R7230 gnd.n5137 gnd.n3570 585
R7231 gnd.n4741 gnd.n4740 585
R7232 gnd.n4740 gnd.n3568 585
R7233 gnd.n4739 gnd.n3688 585
R7234 gnd.n4739 gnd.n4738 585
R7235 gnd.n4712 gnd.n3558 585
R7236 gnd.n5145 gnd.n3558 585
R7237 gnd.n4714 gnd.n4713 585
R7238 gnd.n4715 gnd.n4714 585
R7239 gnd.n4706 gnd.n3548 585
R7240 gnd.n5151 gnd.n3548 585
R7241 gnd.n4705 gnd.n4704 585
R7242 gnd.n4704 gnd.n3546 585
R7243 gnd.n4703 gnd.n3694 585
R7244 gnd.n4703 gnd.n3537 585
R7245 gnd.n4702 gnd.n4701 585
R7246 gnd.n4702 gnd.n3535 585
R7247 gnd.n3697 gnd.n3696 585
R7248 gnd.n4693 gnd.n3696 585
R7249 gnd.n4650 gnd.n4649 585
R7250 gnd.n4649 gnd.n3701 585
R7251 gnd.n4651 gnd.n3711 585
R7252 gnd.n4679 gnd.n3711 585
R7253 gnd.n4648 gnd.n4647 585
R7254 gnd.n4647 gnd.n3717 585
R7255 gnd.n4646 gnd.n3724 585
R7256 gnd.n4646 gnd.n4645 585
R7257 gnd.n4631 gnd.n3725 585
R7258 gnd.n3735 gnd.n3725 585
R7259 gnd.n4630 gnd.n3733 585
R7260 gnd.n4637 gnd.n3733 585
R7261 gnd.n4629 gnd.n4628 585
R7262 gnd.n4628 gnd.n4627 585
R7263 gnd.n3744 gnd.n3741 585
R7264 gnd.n3745 gnd.n3744 585
R7265 gnd.n4619 gnd.n4618 585
R7266 gnd.n4618 gnd.n4617 585
R7267 gnd.n3751 gnd.n3750 585
R7268 gnd.n3762 gnd.n3751 585
R7269 gnd.n4599 gnd.n3760 585
R7270 gnd.n4607 gnd.n3760 585
R7271 gnd.n4598 gnd.n4597 585
R7272 gnd.n4597 gnd.n4596 585
R7273 gnd.n3769 gnd.n3767 585
R7274 gnd.n3770 gnd.n3769 585
R7275 gnd.n4588 gnd.n4587 585
R7276 gnd.n4587 gnd.n4586 585
R7277 gnd.n3776 gnd.n3775 585
R7278 gnd.n3787 gnd.n3776 585
R7279 gnd.n4568 gnd.n3785 585
R7280 gnd.n4576 gnd.n3785 585
R7281 gnd.n4567 gnd.n4566 585
R7282 gnd.n4566 gnd.n4565 585
R7283 gnd.n3794 gnd.n3792 585
R7284 gnd.n3795 gnd.n3794 585
R7285 gnd.n4557 gnd.n4556 585
R7286 gnd.n4556 gnd.n4555 585
R7287 gnd.n3801 gnd.n3800 585
R7288 gnd.n3813 gnd.n3801 585
R7289 gnd.n4537 gnd.n3811 585
R7290 gnd.n4545 gnd.n3811 585
R7291 gnd.n4536 gnd.n4535 585
R7292 gnd.n4535 gnd.n4534 585
R7293 gnd.n3820 gnd.n3818 585
R7294 gnd.n3830 gnd.n3820 585
R7295 gnd.n4526 gnd.n4525 585
R7296 gnd.n4525 gnd.n4524 585
R7297 gnd.n3826 gnd.n3825 585
R7298 gnd.n3839 gnd.n3826 585
R7299 gnd.n4506 gnd.n3837 585
R7300 gnd.n4514 gnd.n3837 585
R7301 gnd.n4505 gnd.n4504 585
R7302 gnd.n4504 gnd.n4503 585
R7303 gnd.n3846 gnd.n3844 585
R7304 gnd.n3856 gnd.n3846 585
R7305 gnd.n4495 gnd.n4494 585
R7306 gnd.n4494 gnd.n4493 585
R7307 gnd.n3852 gnd.n3851 585
R7308 gnd.n3865 gnd.n3852 585
R7309 gnd.n4475 gnd.n3863 585
R7310 gnd.n4483 gnd.n3863 585
R7311 gnd.n4474 gnd.n4473 585
R7312 gnd.n4473 gnd.n4472 585
R7313 gnd.n3872 gnd.n3870 585
R7314 gnd.n3873 gnd.n3872 585
R7315 gnd.n4464 gnd.n4463 585
R7316 gnd.n4463 gnd.n4462 585
R7317 gnd.n3879 gnd.n3878 585
R7318 gnd.n3890 gnd.n3879 585
R7319 gnd.n4444 gnd.n3888 585
R7320 gnd.n4452 gnd.n3888 585
R7321 gnd.n4443 gnd.n4442 585
R7322 gnd.n4442 gnd.n4441 585
R7323 gnd.n5957 gnd.n5956 585
R7324 gnd.n5958 gnd.n5957 585
R7325 gnd.n1607 gnd.n1605 585
R7326 gnd.n5728 gnd.n1605 585
R7327 gnd.n5906 gnd.n5905 585
R7328 gnd.n5905 gnd.n5904 585
R7329 gnd.n1610 gnd.n1609 585
R7330 gnd.n5559 gnd.n1610 585
R7331 gnd.n5720 gnd.n5719 585
R7332 gnd.n5721 gnd.n5720 585
R7333 gnd.n1765 gnd.n1764 585
R7334 gnd.n5563 gnd.n1764 585
R7335 gnd.n5715 gnd.n5714 585
R7336 gnd.n5714 gnd.n5713 585
R7337 gnd.n1768 gnd.n1767 585
R7338 gnd.n5569 gnd.n1768 585
R7339 gnd.n5699 gnd.n5698 585
R7340 gnd.n5700 gnd.n5699 585
R7341 gnd.n1784 gnd.n1783 585
R7342 gnd.n5497 gnd.n1783 585
R7343 gnd.n5694 gnd.n5693 585
R7344 gnd.n5693 gnd.n5692 585
R7345 gnd.n1787 gnd.n1786 585
R7346 gnd.n5501 gnd.n1787 585
R7347 gnd.n5683 gnd.n5682 585
R7348 gnd.n5684 gnd.n5683 585
R7349 gnd.n1802 gnd.n1801 585
R7350 gnd.n5505 gnd.n1801 585
R7351 gnd.n5678 gnd.n5677 585
R7352 gnd.n5677 gnd.n5676 585
R7353 gnd.n1805 gnd.n1804 585
R7354 gnd.n5511 gnd.n1805 585
R7355 gnd.n5667 gnd.n5666 585
R7356 gnd.n5668 gnd.n5667 585
R7357 gnd.n1819 gnd.n1818 585
R7358 gnd.n5484 gnd.n1818 585
R7359 gnd.n5662 gnd.n5661 585
R7360 gnd.n5661 gnd.n5660 585
R7361 gnd.n1822 gnd.n1821 585
R7362 gnd.n5480 gnd.n1822 585
R7363 gnd.n5651 gnd.n5650 585
R7364 gnd.n5652 gnd.n5651 585
R7365 gnd.n1837 gnd.n1836 585
R7366 gnd.n5596 gnd.n1836 585
R7367 gnd.n5619 gnd.n1881 585
R7368 gnd.n5619 gnd.n5618 585
R7369 gnd.n5622 gnd.n5621 585
R7370 gnd.n5623 gnd.n5622 585
R7371 gnd.n5620 gnd.n1880 585
R7372 gnd.n1880 gnd.n1875 585
R7373 gnd.n1864 gnd.n1863 585
R7374 gnd.n1868 gnd.n1863 585
R7375 gnd.n5633 gnd.n1865 585
R7376 gnd.n5633 gnd.n5632 585
R7377 gnd.n5636 gnd.n5635 585
R7378 gnd.n5637 gnd.n5636 585
R7379 gnd.n5634 gnd.n1846 585
R7380 gnd.n5405 gnd.n1846 585
R7381 gnd.n5645 gnd.n5644 585
R7382 gnd.n5644 gnd.n5643 585
R7383 gnd.n5646 gnd.n1845 585
R7384 gnd.n5397 gnd.n1845 585
R7385 gnd.n1915 gnd.n1844 585
R7386 gnd.n1934 gnd.n1915 585
R7387 gnd.n5387 gnd.n5386 585
R7388 gnd.n5388 gnd.n5387 585
R7389 gnd.n5385 gnd.n1914 585
R7390 gnd.n5373 gnd.n1914 585
R7391 gnd.n1920 gnd.n1916 585
R7392 gnd.n5356 gnd.n1920 585
R7393 gnd.n5381 gnd.n5380 585
R7394 gnd.n5380 gnd.n5379 585
R7395 gnd.n1919 gnd.n1918 585
R7396 gnd.n5362 gnd.n1919 585
R7397 gnd.n5345 gnd.n1955 585
R7398 gnd.n5331 gnd.n1955 585
R7399 gnd.n5347 gnd.n5346 585
R7400 gnd.n5348 gnd.n5347 585
R7401 gnd.n1956 gnd.n1954 585
R7402 gnd.n2206 gnd.n1954 585
R7403 gnd.n5340 gnd.n5339 585
R7404 gnd.n5339 gnd.n5338 585
R7405 gnd.n1959 gnd.n1958 585
R7406 gnd.n2212 gnd.n1959 585
R7407 gnd.n5320 gnd.n5319 585
R7408 gnd.n5321 gnd.n5320 585
R7409 gnd.n1974 gnd.n1973 585
R7410 gnd.n5221 gnd.n1973 585
R7411 gnd.n5315 gnd.n5314 585
R7412 gnd.n5314 gnd.n5313 585
R7413 gnd.n1977 gnd.n1976 585
R7414 gnd.n5227 gnd.n1977 585
R7415 gnd.n5304 gnd.n5303 585
R7416 gnd.n5305 gnd.n5304 585
R7417 gnd.n1992 gnd.n1991 585
R7418 gnd.n1991 gnd.n1987 585
R7419 gnd.n5299 gnd.n5298 585
R7420 gnd.n5298 gnd.n5297 585
R7421 gnd.n1995 gnd.n1994 585
R7422 gnd.n1996 gnd.n1995 585
R7423 gnd.n5288 gnd.n5287 585
R7424 gnd.n5289 gnd.n5288 585
R7425 gnd.n2009 gnd.n2008 585
R7426 gnd.n2008 gnd.n2005 585
R7427 gnd.n5283 gnd.n5282 585
R7428 gnd.n5282 gnd.n5281 585
R7429 gnd.n2085 gnd.n2011 585
R7430 gnd.n2088 gnd.n2087 585
R7431 gnd.n2084 gnd.n2083 585
R7432 gnd.n2083 gnd.n2012 585
R7433 gnd.n2093 gnd.n2092 585
R7434 gnd.n2095 gnd.n2082 585
R7435 gnd.n2098 gnd.n2097 585
R7436 gnd.n2080 gnd.n2079 585
R7437 gnd.n2103 gnd.n2102 585
R7438 gnd.n2105 gnd.n2078 585
R7439 gnd.n2108 gnd.n2107 585
R7440 gnd.n2076 gnd.n2075 585
R7441 gnd.n2113 gnd.n2112 585
R7442 gnd.n2115 gnd.n2074 585
R7443 gnd.n2118 gnd.n2117 585
R7444 gnd.n2072 gnd.n2071 585
R7445 gnd.n2126 gnd.n2125 585
R7446 gnd.n2128 gnd.n2070 585
R7447 gnd.n2131 gnd.n2130 585
R7448 gnd.n2068 gnd.n2067 585
R7449 gnd.n2136 gnd.n2135 585
R7450 gnd.n2138 gnd.n2066 585
R7451 gnd.n2141 gnd.n2140 585
R7452 gnd.n2064 gnd.n2063 585
R7453 gnd.n2146 gnd.n2145 585
R7454 gnd.n2148 gnd.n2062 585
R7455 gnd.n2151 gnd.n2150 585
R7456 gnd.n2060 gnd.n2059 585
R7457 gnd.n2156 gnd.n2155 585
R7458 gnd.n2158 gnd.n2058 585
R7459 gnd.n2161 gnd.n2160 585
R7460 gnd.n2056 gnd.n2055 585
R7461 gnd.n2167 gnd.n2166 585
R7462 gnd.n2169 gnd.n2054 585
R7463 gnd.n2170 gnd.n2053 585
R7464 gnd.n2173 gnd.n2172 585
R7465 gnd.n1600 gnd.n1593 585
R7466 gnd.n5964 gnd.n1590 585
R7467 gnd.n5966 gnd.n5965 585
R7468 gnd.n5968 gnd.n1588 585
R7469 gnd.n5970 gnd.n5969 585
R7470 gnd.n5971 gnd.n1583 585
R7471 gnd.n5973 gnd.n5972 585
R7472 gnd.n5975 gnd.n1581 585
R7473 gnd.n5977 gnd.n5976 585
R7474 gnd.n5978 gnd.n1576 585
R7475 gnd.n5980 gnd.n5979 585
R7476 gnd.n5982 gnd.n1574 585
R7477 gnd.n5984 gnd.n5983 585
R7478 gnd.n5985 gnd.n1569 585
R7479 gnd.n5987 gnd.n5986 585
R7480 gnd.n5989 gnd.n1568 585
R7481 gnd.n5990 gnd.n1564 585
R7482 gnd.n5993 gnd.n5992 585
R7483 gnd.n1565 gnd.n1557 585
R7484 gnd.n5928 gnd.n1558 585
R7485 gnd.n5932 gnd.n5931 585
R7486 gnd.n5934 gnd.n5925 585
R7487 gnd.n5936 gnd.n5935 585
R7488 gnd.n5937 gnd.n5920 585
R7489 gnd.n5939 gnd.n5938 585
R7490 gnd.n5941 gnd.n5918 585
R7491 gnd.n5943 gnd.n5942 585
R7492 gnd.n5944 gnd.n5912 585
R7493 gnd.n5946 gnd.n5945 585
R7494 gnd.n5948 gnd.n5911 585
R7495 gnd.n5949 gnd.n5910 585
R7496 gnd.n5952 gnd.n5951 585
R7497 gnd.n5953 gnd.n1606 585
R7498 gnd.n1606 gnd.n1567 585
R7499 gnd.n5960 gnd.n5959 585
R7500 gnd.n5959 gnd.n5958 585
R7501 gnd.n1598 gnd.n1597 585
R7502 gnd.n5728 gnd.n1598 585
R7503 gnd.n5439 gnd.n1611 585
R7504 gnd.n5904 gnd.n1611 585
R7505 gnd.n5561 gnd.n5560 585
R7506 gnd.n5560 gnd.n5559 585
R7507 gnd.n5562 gnd.n1761 585
R7508 gnd.n5721 gnd.n1761 585
R7509 gnd.n5565 gnd.n5564 585
R7510 gnd.n5564 gnd.n5563 585
R7511 gnd.n5566 gnd.n1770 585
R7512 gnd.n5713 gnd.n1770 585
R7513 gnd.n5568 gnd.n5567 585
R7514 gnd.n5569 gnd.n5568 585
R7515 gnd.n5432 gnd.n1780 585
R7516 gnd.n5700 gnd.n1780 585
R7517 gnd.n5499 gnd.n5498 585
R7518 gnd.n5498 gnd.n5497 585
R7519 gnd.n5500 gnd.n1789 585
R7520 gnd.n5692 gnd.n1789 585
R7521 gnd.n5503 gnd.n5502 585
R7522 gnd.n5502 gnd.n5501 585
R7523 gnd.n5504 gnd.n1798 585
R7524 gnd.n5684 gnd.n1798 585
R7525 gnd.n5507 gnd.n5506 585
R7526 gnd.n5506 gnd.n5505 585
R7527 gnd.n5508 gnd.n1806 585
R7528 gnd.n5676 gnd.n1806 585
R7529 gnd.n5510 gnd.n5509 585
R7530 gnd.n5511 gnd.n5510 585
R7531 gnd.n5476 gnd.n1815 585
R7532 gnd.n5668 gnd.n1815 585
R7533 gnd.n5486 gnd.n5485 585
R7534 gnd.n5485 gnd.n5484 585
R7535 gnd.n5483 gnd.n1824 585
R7536 gnd.n5660 gnd.n1824 585
R7537 gnd.n5482 gnd.n5481 585
R7538 gnd.n5481 gnd.n5480 585
R7539 gnd.n1893 gnd.n1833 585
R7540 gnd.n5652 gnd.n1833 585
R7541 gnd.n5598 gnd.n5597 585
R7542 gnd.n5597 gnd.n5596 585
R7543 gnd.n5599 gnd.n1882 585
R7544 gnd.n5618 gnd.n1882 585
R7545 gnd.n5600 gnd.n1876 585
R7546 gnd.n5623 gnd.n1876 585
R7547 gnd.n5602 gnd.n5601 585
R7548 gnd.n5602 gnd.n1875 585
R7549 gnd.n5604 gnd.n5603 585
R7550 gnd.n5603 gnd.n1868 585
R7551 gnd.n5605 gnd.n1866 585
R7552 gnd.n5632 gnd.n1866 585
R7553 gnd.n1888 gnd.n1860 585
R7554 gnd.n5637 gnd.n1860 585
R7555 gnd.n5404 gnd.n5403 585
R7556 gnd.n5405 gnd.n5404 585
R7557 gnd.n1900 gnd.n1848 585
R7558 gnd.n5643 gnd.n1848 585
R7559 gnd.n5399 gnd.n5398 585
R7560 gnd.n5398 gnd.n5397 585
R7561 gnd.n1903 gnd.n1902 585
R7562 gnd.n1934 gnd.n1903 585
R7563 gnd.n5370 gnd.n1911 585
R7564 gnd.n5388 gnd.n1911 585
R7565 gnd.n5372 gnd.n5371 585
R7566 gnd.n5373 gnd.n5372 585
R7567 gnd.n1940 gnd.n1939 585
R7568 gnd.n5356 gnd.n1939 585
R7569 gnd.n5365 gnd.n1922 585
R7570 gnd.n5379 gnd.n1922 585
R7571 gnd.n5364 gnd.n5363 585
R7572 gnd.n5363 gnd.n5362 585
R7573 gnd.n1943 gnd.n1942 585
R7574 gnd.n5331 gnd.n1943 585
R7575 gnd.n2205 gnd.n1951 585
R7576 gnd.n5348 gnd.n1951 585
R7577 gnd.n2208 gnd.n2207 585
R7578 gnd.n2207 gnd.n2206 585
R7579 gnd.n2209 gnd.n1961 585
R7580 gnd.n5338 gnd.n1961 585
R7581 gnd.n2211 gnd.n2210 585
R7582 gnd.n2212 gnd.n2211 585
R7583 gnd.n2192 gnd.n1970 585
R7584 gnd.n5321 gnd.n1970 585
R7585 gnd.n5223 gnd.n5222 585
R7586 gnd.n5222 gnd.n5221 585
R7587 gnd.n5224 gnd.n1979 585
R7588 gnd.n5313 gnd.n1979 585
R7589 gnd.n5226 gnd.n5225 585
R7590 gnd.n5227 gnd.n5226 585
R7591 gnd.n2047 gnd.n1988 585
R7592 gnd.n5305 gnd.n1988 585
R7593 gnd.n2186 gnd.n2185 585
R7594 gnd.n2185 gnd.n1987 585
R7595 gnd.n2184 gnd.n1997 585
R7596 gnd.n5297 gnd.n1997 585
R7597 gnd.n2183 gnd.n2182 585
R7598 gnd.n2182 gnd.n1996 585
R7599 gnd.n2049 gnd.n2006 585
R7600 gnd.n5289 gnd.n2006 585
R7601 gnd.n2178 gnd.n2177 585
R7602 gnd.n2177 gnd.n2005 585
R7603 gnd.n2176 gnd.n2013 585
R7604 gnd.n5281 gnd.n2013 585
R7605 gnd.n7352 gnd.n7351 585
R7606 gnd.n7353 gnd.n7352 585
R7607 gnd.n506 gnd.n504 585
R7608 gnd.n504 gnd.n500 585
R7609 gnd.n7282 gnd.n7281 585
R7610 gnd.n7283 gnd.n7282 585
R7611 gnd.n579 gnd.n578 585
R7612 gnd.n585 gnd.n578 585
R7613 gnd.n7277 gnd.n7276 585
R7614 gnd.n7276 gnd.n7275 585
R7615 gnd.n582 gnd.n581 585
R7616 gnd.n596 gnd.n582 585
R7617 gnd.n7198 gnd.n7197 585
R7618 gnd.n7199 gnd.n7198 585
R7619 gnd.n598 gnd.n597 585
R7620 gnd.n2882 gnd.n597 585
R7621 gnd.n7193 gnd.n7192 585
R7622 gnd.n7192 gnd.n7191 585
R7623 gnd.n601 gnd.n600 585
R7624 gnd.n2888 gnd.n601 585
R7625 gnd.n7182 gnd.n7181 585
R7626 gnd.n7183 gnd.n7182 585
R7627 gnd.n614 gnd.n613 585
R7628 gnd.n2864 gnd.n613 585
R7629 gnd.n7177 gnd.n7176 585
R7630 gnd.n7176 gnd.n7175 585
R7631 gnd.n617 gnd.n616 585
R7632 gnd.n2860 gnd.n617 585
R7633 gnd.n7166 gnd.n7165 585
R7634 gnd.n7167 gnd.n7166 585
R7635 gnd.n631 gnd.n630 585
R7636 gnd.n2854 gnd.n630 585
R7637 gnd.n7161 gnd.n7160 585
R7638 gnd.n7160 gnd.n7159 585
R7639 gnd.n634 gnd.n633 585
R7640 gnd.n2850 gnd.n634 585
R7641 gnd.n7150 gnd.n7149 585
R7642 gnd.n7151 gnd.n7150 585
R7643 gnd.n648 gnd.n647 585
R7644 gnd.n2844 gnd.n647 585
R7645 gnd.n7145 gnd.n7144 585
R7646 gnd.n7144 gnd.n7143 585
R7647 gnd.n651 gnd.n650 585
R7648 gnd.n2840 gnd.n651 585
R7649 gnd.n7134 gnd.n7133 585
R7650 gnd.n7135 gnd.n7134 585
R7651 gnd.n7131 gnd.n664 585
R7652 gnd.n6844 gnd.n664 585
R7653 gnd.n7130 gnd.n7129 585
R7654 gnd.n7129 gnd.n7128 585
R7655 gnd.n7117 gnd.n666 585
R7656 gnd.n6848 gnd.n666 585
R7657 gnd.n7119 gnd.n7118 585
R7658 gnd.n7120 gnd.n7119 585
R7659 gnd.n7115 gnd.n679 585
R7660 gnd.n6854 gnd.n679 585
R7661 gnd.n7114 gnd.n7113 585
R7662 gnd.n7113 gnd.n7112 585
R7663 gnd.n7101 gnd.n681 585
R7664 gnd.n6793 gnd.n681 585
R7665 gnd.n7103 gnd.n7102 585
R7666 gnd.n7104 gnd.n7103 585
R7667 gnd.n7099 gnd.n695 585
R7668 gnd.n6797 gnd.n695 585
R7669 gnd.n7098 gnd.n7097 585
R7670 gnd.n7097 gnd.n7096 585
R7671 gnd.n698 gnd.n696 585
R7672 gnd.n6801 gnd.n698 585
R7673 gnd.n7087 gnd.n7086 585
R7674 gnd.n7088 gnd.n7087 585
R7675 gnd.n713 gnd.n712 585
R7676 gnd.n6805 gnd.n712 585
R7677 gnd.n7081 gnd.n7080 585
R7678 gnd.n7080 gnd.n7079 585
R7679 gnd.n716 gnd.n715 585
R7680 gnd.n6811 gnd.n716 585
R7681 gnd.n7070 gnd.n7069 585
R7682 gnd.n7071 gnd.n7070 585
R7683 gnd.n730 gnd.n729 585
R7684 gnd.n6778 gnd.n729 585
R7685 gnd.n7065 gnd.n7064 585
R7686 gnd.n7064 gnd.n7063 585
R7687 gnd.n733 gnd.n732 585
R7688 gnd.n6774 gnd.n733 585
R7689 gnd.n7054 gnd.n7053 585
R7690 gnd.n7055 gnd.n7054 585
R7691 gnd.n748 gnd.n747 585
R7692 gnd.n6768 gnd.n747 585
R7693 gnd.n7049 gnd.n7048 585
R7694 gnd.n7048 gnd.n7047 585
R7695 gnd.n751 gnd.n750 585
R7696 gnd.n6764 gnd.n751 585
R7697 gnd.n7038 gnd.n7037 585
R7698 gnd.n7039 gnd.n7038 585
R7699 gnd.n766 gnd.n765 585
R7700 gnd.n6758 gnd.n765 585
R7701 gnd.n7033 gnd.n7032 585
R7702 gnd.n7032 gnd.n7031 585
R7703 gnd.n769 gnd.n768 585
R7704 gnd.n6892 gnd.n769 585
R7705 gnd.n7022 gnd.n7021 585
R7706 gnd.n7023 gnd.n7022 585
R7707 gnd.n783 gnd.n782 585
R7708 gnd.n1013 gnd.n782 585
R7709 gnd.n7017 gnd.n7016 585
R7710 gnd.n7016 gnd.n7015 585
R7711 gnd.n863 gnd.n785 585
R7712 gnd.n6962 gnd.n6961 585
R7713 gnd.n6960 gnd.n862 585
R7714 gnd.n6964 gnd.n862 585
R7715 gnd.n6959 gnd.n6958 585
R7716 gnd.n6957 gnd.n6956 585
R7717 gnd.n6955 gnd.n6954 585
R7718 gnd.n6953 gnd.n6952 585
R7719 gnd.n6951 gnd.n6950 585
R7720 gnd.n6949 gnd.n6948 585
R7721 gnd.n6947 gnd.n6946 585
R7722 gnd.n6945 gnd.n6944 585
R7723 gnd.n6943 gnd.n6942 585
R7724 gnd.n6941 gnd.n6940 585
R7725 gnd.n6939 gnd.n6938 585
R7726 gnd.n6936 gnd.n6935 585
R7727 gnd.n6934 gnd.n6933 585
R7728 gnd.n6932 gnd.n6931 585
R7729 gnd.n6930 gnd.n6929 585
R7730 gnd.n6928 gnd.n6927 585
R7731 gnd.n6926 gnd.n6925 585
R7732 gnd.n6924 gnd.n6923 585
R7733 gnd.n6922 gnd.n6921 585
R7734 gnd.n6920 gnd.n6919 585
R7735 gnd.n6918 gnd.n6917 585
R7736 gnd.n6916 gnd.n6915 585
R7737 gnd.n6914 gnd.n6913 585
R7738 gnd.n6912 gnd.n6911 585
R7739 gnd.n6910 gnd.n6909 585
R7740 gnd.n6908 gnd.n6907 585
R7741 gnd.n6906 gnd.n6905 585
R7742 gnd.n6904 gnd.n898 585
R7743 gnd.n902 gnd.n899 585
R7744 gnd.n6900 gnd.n6899 585
R7745 gnd.n570 gnd.n569 585
R7746 gnd.n7291 gnd.n565 585
R7747 gnd.n7293 gnd.n7292 585
R7748 gnd.n7295 gnd.n563 585
R7749 gnd.n7297 gnd.n7296 585
R7750 gnd.n7298 gnd.n558 585
R7751 gnd.n7300 gnd.n7299 585
R7752 gnd.n7302 gnd.n556 585
R7753 gnd.n7304 gnd.n7303 585
R7754 gnd.n7305 gnd.n551 585
R7755 gnd.n7307 gnd.n7306 585
R7756 gnd.n7309 gnd.n549 585
R7757 gnd.n7311 gnd.n7310 585
R7758 gnd.n7312 gnd.n544 585
R7759 gnd.n7314 gnd.n7313 585
R7760 gnd.n7316 gnd.n542 585
R7761 gnd.n7318 gnd.n7317 585
R7762 gnd.n7319 gnd.n534 585
R7763 gnd.n7321 gnd.n7320 585
R7764 gnd.n7323 gnd.n532 585
R7765 gnd.n7325 gnd.n7324 585
R7766 gnd.n7326 gnd.n527 585
R7767 gnd.n7328 gnd.n7327 585
R7768 gnd.n7330 gnd.n525 585
R7769 gnd.n7332 gnd.n7331 585
R7770 gnd.n7333 gnd.n520 585
R7771 gnd.n7335 gnd.n7334 585
R7772 gnd.n7337 gnd.n518 585
R7773 gnd.n7339 gnd.n7338 585
R7774 gnd.n7340 gnd.n513 585
R7775 gnd.n7342 gnd.n7341 585
R7776 gnd.n7344 gnd.n511 585
R7777 gnd.n7346 gnd.n7345 585
R7778 gnd.n7347 gnd.n509 585
R7779 gnd.n7348 gnd.n505 585
R7780 gnd.n505 gnd.n502 585
R7781 gnd.n7287 gnd.n501 585
R7782 gnd.n7353 gnd.n501 585
R7783 gnd.n7286 gnd.n7285 585
R7784 gnd.n7285 gnd.n500 585
R7785 gnd.n7284 gnd.n574 585
R7786 gnd.n7284 gnd.n7283 585
R7787 gnd.n2877 gnd.n575 585
R7788 gnd.n585 gnd.n575 585
R7789 gnd.n2878 gnd.n584 585
R7790 gnd.n7275 gnd.n584 585
R7791 gnd.n2880 gnd.n2879 585
R7792 gnd.n2879 gnd.n596 585
R7793 gnd.n2881 gnd.n594 585
R7794 gnd.n7199 gnd.n594 585
R7795 gnd.n2884 gnd.n2883 585
R7796 gnd.n2883 gnd.n2882 585
R7797 gnd.n2885 gnd.n603 585
R7798 gnd.n7191 gnd.n603 585
R7799 gnd.n2887 gnd.n2886 585
R7800 gnd.n2888 gnd.n2887 585
R7801 gnd.n2832 gnd.n611 585
R7802 gnd.n7183 gnd.n611 585
R7803 gnd.n2866 gnd.n2865 585
R7804 gnd.n2865 gnd.n2864 585
R7805 gnd.n2863 gnd.n619 585
R7806 gnd.n7175 gnd.n619 585
R7807 gnd.n2862 gnd.n2861 585
R7808 gnd.n2861 gnd.n2860 585
R7809 gnd.n2834 gnd.n627 585
R7810 gnd.n7167 gnd.n627 585
R7811 gnd.n2856 gnd.n2855 585
R7812 gnd.n2855 gnd.n2854 585
R7813 gnd.n2853 gnd.n636 585
R7814 gnd.n7159 gnd.n636 585
R7815 gnd.n2852 gnd.n2851 585
R7816 gnd.n2851 gnd.n2850 585
R7817 gnd.n2836 gnd.n644 585
R7818 gnd.n7151 gnd.n644 585
R7819 gnd.n2846 gnd.n2845 585
R7820 gnd.n2845 gnd.n2844 585
R7821 gnd.n2843 gnd.n653 585
R7822 gnd.n7143 gnd.n653 585
R7823 gnd.n2842 gnd.n2841 585
R7824 gnd.n2841 gnd.n2840 585
R7825 gnd.n936 gnd.n661 585
R7826 gnd.n7135 gnd.n661 585
R7827 gnd.n6846 gnd.n6845 585
R7828 gnd.n6845 gnd.n6844 585
R7829 gnd.n6847 gnd.n668 585
R7830 gnd.n7128 gnd.n668 585
R7831 gnd.n6850 gnd.n6849 585
R7832 gnd.n6849 gnd.n6848 585
R7833 gnd.n6851 gnd.n676 585
R7834 gnd.n7120 gnd.n676 585
R7835 gnd.n6853 gnd.n6852 585
R7836 gnd.n6854 gnd.n6853 585
R7837 gnd.n931 gnd.n683 585
R7838 gnd.n7112 gnd.n683 585
R7839 gnd.n6795 gnd.n6794 585
R7840 gnd.n6794 gnd.n6793 585
R7841 gnd.n6796 gnd.n692 585
R7842 gnd.n7104 gnd.n692 585
R7843 gnd.n6799 gnd.n6798 585
R7844 gnd.n6798 gnd.n6797 585
R7845 gnd.n6800 gnd.n700 585
R7846 gnd.n7096 gnd.n700 585
R7847 gnd.n6803 gnd.n6802 585
R7848 gnd.n6802 gnd.n6801 585
R7849 gnd.n6804 gnd.n709 585
R7850 gnd.n7088 gnd.n709 585
R7851 gnd.n6807 gnd.n6806 585
R7852 gnd.n6806 gnd.n6805 585
R7853 gnd.n6808 gnd.n718 585
R7854 gnd.n7079 gnd.n718 585
R7855 gnd.n6810 gnd.n6809 585
R7856 gnd.n6811 gnd.n6810 585
R7857 gnd.n6752 gnd.n727 585
R7858 gnd.n7071 gnd.n727 585
R7859 gnd.n6780 gnd.n6779 585
R7860 gnd.n6779 gnd.n6778 585
R7861 gnd.n6777 gnd.n735 585
R7862 gnd.n7063 gnd.n735 585
R7863 gnd.n6776 gnd.n6775 585
R7864 gnd.n6775 gnd.n6774 585
R7865 gnd.n6754 gnd.n744 585
R7866 gnd.n7055 gnd.n744 585
R7867 gnd.n6770 gnd.n6769 585
R7868 gnd.n6769 gnd.n6768 585
R7869 gnd.n6767 gnd.n753 585
R7870 gnd.n7047 gnd.n753 585
R7871 gnd.n6766 gnd.n6765 585
R7872 gnd.n6765 gnd.n6764 585
R7873 gnd.n6756 gnd.n762 585
R7874 gnd.n7039 gnd.n762 585
R7875 gnd.n6760 gnd.n6759 585
R7876 gnd.n6759 gnd.n6758 585
R7877 gnd.n907 gnd.n771 585
R7878 gnd.n7031 gnd.n771 585
R7879 gnd.n6894 gnd.n6893 585
R7880 gnd.n6893 gnd.n6892 585
R7881 gnd.n6895 gnd.n780 585
R7882 gnd.n7023 gnd.n780 585
R7883 gnd.n6896 gnd.n904 585
R7884 gnd.n1013 gnd.n904 585
R7885 gnd.n6897 gnd.n787 585
R7886 gnd.n7015 gnd.n787 585
R7887 gnd.n6607 gnd.n1113 585
R7888 gnd.n1182 gnd.n1113 585
R7889 gnd.n6609 gnd.n6608 585
R7890 gnd.n6610 gnd.n6609 585
R7891 gnd.n1114 gnd.n1112 585
R7892 gnd.n6495 gnd.n1112 585
R7893 gnd.n6492 gnd.n6491 585
R7894 gnd.n6493 gnd.n6492 585
R7895 gnd.n6490 gnd.n1186 585
R7896 gnd.n1191 gnd.n1186 585
R7897 gnd.n6489 gnd.n6488 585
R7898 gnd.n6488 gnd.n6487 585
R7899 gnd.n1188 gnd.n1187 585
R7900 gnd.n6459 gnd.n1188 585
R7901 gnd.n6472 gnd.n6471 585
R7902 gnd.n6473 gnd.n6472 585
R7903 gnd.n6470 gnd.n1203 585
R7904 gnd.n1203 gnd.n1199 585
R7905 gnd.n6469 gnd.n6468 585
R7906 gnd.n6468 gnd.n6467 585
R7907 gnd.n1205 gnd.n1204 585
R7908 gnd.n6447 gnd.n1205 585
R7909 gnd.n6432 gnd.n6431 585
R7910 gnd.n6431 gnd.n1220 585
R7911 gnd.n6433 gnd.n1231 585
R7912 gnd.n6419 gnd.n1231 585
R7913 gnd.n6435 gnd.n6434 585
R7914 gnd.n6436 gnd.n6435 585
R7915 gnd.n6430 gnd.n1230 585
R7916 gnd.n1230 gnd.n1227 585
R7917 gnd.n6429 gnd.n6428 585
R7918 gnd.n6428 gnd.n6427 585
R7919 gnd.n1233 gnd.n1232 585
R7920 gnd.n6410 gnd.n1233 585
R7921 gnd.n6396 gnd.n6395 585
R7922 gnd.n6395 gnd.n1248 585
R7923 gnd.n6397 gnd.n1260 585
R7924 gnd.n1273 gnd.n1260 585
R7925 gnd.n6399 gnd.n6398 585
R7926 gnd.n6400 gnd.n6399 585
R7927 gnd.n6394 gnd.n1259 585
R7928 gnd.n1259 gnd.n1255 585
R7929 gnd.n6393 gnd.n6392 585
R7930 gnd.n6392 gnd.n6391 585
R7931 gnd.n1262 gnd.n1261 585
R7932 gnd.n1279 gnd.n1262 585
R7933 gnd.n6327 gnd.n6326 585
R7934 gnd.n6326 gnd.n6325 585
R7935 gnd.n6328 gnd.n1290 585
R7936 gnd.n1294 gnd.n1290 585
R7937 gnd.n6330 gnd.n6329 585
R7938 gnd.n6331 gnd.n6330 585
R7939 gnd.n1291 gnd.n1289 585
R7940 gnd.n1289 gnd.n1285 585
R7941 gnd.n6309 gnd.n6308 585
R7942 gnd.n6310 gnd.n6309 585
R7943 gnd.n6307 gnd.n1301 585
R7944 gnd.n1306 gnd.n1301 585
R7945 gnd.n6306 gnd.n6305 585
R7946 gnd.n6305 gnd.n6304 585
R7947 gnd.n1303 gnd.n1302 585
R7948 gnd.n6259 gnd.n1303 585
R7949 gnd.n6262 gnd.n1330 585
R7950 gnd.n6262 gnd.n6261 585
R7951 gnd.n6264 gnd.n6263 585
R7952 gnd.n6263 gnd.n1314 585
R7953 gnd.n6265 gnd.n1328 585
R7954 gnd.n6250 gnd.n1328 585
R7955 gnd.n6267 gnd.n6266 585
R7956 gnd.n6268 gnd.n6267 585
R7957 gnd.n1329 gnd.n1327 585
R7958 gnd.n6227 gnd.n1327 585
R7959 gnd.n6217 gnd.n1345 585
R7960 gnd.n1345 gnd.n1338 585
R7961 gnd.n6219 gnd.n6218 585
R7962 gnd.n6220 gnd.n6219 585
R7963 gnd.n6216 gnd.n1344 585
R7964 gnd.n1351 gnd.n1344 585
R7965 gnd.n6215 gnd.n6214 585
R7966 gnd.n6214 gnd.n6213 585
R7967 gnd.n1347 gnd.n1346 585
R7968 gnd.n6106 gnd.n1347 585
R7969 gnd.n6201 gnd.n6200 585
R7970 gnd.n6202 gnd.n6201 585
R7971 gnd.n6199 gnd.n1363 585
R7972 gnd.n1363 gnd.n1359 585
R7973 gnd.n6198 gnd.n6197 585
R7974 gnd.n6197 gnd.n6196 585
R7975 gnd.n1365 gnd.n1364 585
R7976 gnd.n6096 gnd.n1365 585
R7977 gnd.n6169 gnd.n6168 585
R7978 gnd.n6170 gnd.n6169 585
R7979 gnd.n6167 gnd.n1377 585
R7980 gnd.n6162 gnd.n1377 585
R7981 gnd.n6166 gnd.n6165 585
R7982 gnd.n6165 gnd.n6164 585
R7983 gnd.n1379 gnd.n1378 585
R7984 gnd.n1393 gnd.n1379 585
R7985 gnd.n6138 gnd.n6137 585
R7986 gnd.n6137 gnd.n1391 585
R7987 gnd.n6139 gnd.n1402 585
R7988 gnd.n6125 gnd.n1402 585
R7989 gnd.n6141 gnd.n6140 585
R7990 gnd.n6142 gnd.n6141 585
R7991 gnd.n6136 gnd.n1401 585
R7992 gnd.n6131 gnd.n1401 585
R7993 gnd.n6135 gnd.n6134 585
R7994 gnd.n6134 gnd.n6133 585
R7995 gnd.n1404 gnd.n1403 585
R7996 gnd.n1496 gnd.n1404 585
R7997 gnd.n1486 gnd.n1465 585
R7998 gnd.n1465 gnd.n1425 585
R7999 gnd.n6057 gnd.n6056 585
R8000 gnd.n6055 gnd.n1464 585
R8001 gnd.n6054 gnd.n1463 585
R8002 gnd.n6059 gnd.n1463 585
R8003 gnd.n6053 gnd.n6052 585
R8004 gnd.n6051 gnd.n6050 585
R8005 gnd.n6049 gnd.n6048 585
R8006 gnd.n6047 gnd.n6046 585
R8007 gnd.n6045 gnd.n6044 585
R8008 gnd.n6043 gnd.n6042 585
R8009 gnd.n6041 gnd.n6040 585
R8010 gnd.n6039 gnd.n6038 585
R8011 gnd.n6037 gnd.n6036 585
R8012 gnd.n6035 gnd.n6034 585
R8013 gnd.n6033 gnd.n6032 585
R8014 gnd.n6031 gnd.n6030 585
R8015 gnd.n6029 gnd.n6028 585
R8016 gnd.n6027 gnd.n6026 585
R8017 gnd.n6025 gnd.n6024 585
R8018 gnd.n6023 gnd.n6022 585
R8019 gnd.n6021 gnd.n6020 585
R8020 gnd.n6019 gnd.n6018 585
R8021 gnd.n6017 gnd.n6016 585
R8022 gnd.n6015 gnd.n6014 585
R8023 gnd.n6013 gnd.n6012 585
R8024 gnd.n6011 gnd.n6010 585
R8025 gnd.n6009 gnd.n6008 585
R8026 gnd.n6006 gnd.n6005 585
R8027 gnd.n6004 gnd.n6003 585
R8028 gnd.n6002 gnd.n6001 585
R8029 gnd.n6000 gnd.n5999 585
R8030 gnd.n1556 gnd.n1555 585
R8031 gnd.n1554 gnd.n1553 585
R8032 gnd.n1552 gnd.n1551 585
R8033 gnd.n1550 gnd.n1549 585
R8034 gnd.n1548 gnd.n1547 585
R8035 gnd.n1546 gnd.n1545 585
R8036 gnd.n1544 gnd.n1543 585
R8037 gnd.n1542 gnd.n1541 585
R8038 gnd.n1540 gnd.n1539 585
R8039 gnd.n1538 gnd.n1537 585
R8040 gnd.n1536 gnd.n1535 585
R8041 gnd.n1534 gnd.n1533 585
R8042 gnd.n1532 gnd.n1531 585
R8043 gnd.n1530 gnd.n1529 585
R8044 gnd.n1528 gnd.n1527 585
R8045 gnd.n1526 gnd.n1525 585
R8046 gnd.n1524 gnd.n1523 585
R8047 gnd.n1522 gnd.n1521 585
R8048 gnd.n1520 gnd.n1519 585
R8049 gnd.n1518 gnd.n1517 585
R8050 gnd.n1516 gnd.n1515 585
R8051 gnd.n1514 gnd.n1513 585
R8052 gnd.n1512 gnd.n1511 585
R8053 gnd.n1510 gnd.n1509 585
R8054 gnd.n1508 gnd.n1507 585
R8055 gnd.n1506 gnd.n1505 585
R8056 gnd.n1504 gnd.n1503 585
R8057 gnd.n1502 gnd.n1501 585
R8058 gnd.n1500 gnd.n1499 585
R8059 gnd.n6501 gnd.n6500 585
R8060 gnd.n6503 gnd.n1180 585
R8061 gnd.n6505 gnd.n6504 585
R8062 gnd.n6506 gnd.n1179 585
R8063 gnd.n6508 gnd.n6507 585
R8064 gnd.n6510 gnd.n1177 585
R8065 gnd.n6512 gnd.n6511 585
R8066 gnd.n6513 gnd.n1176 585
R8067 gnd.n6515 gnd.n6514 585
R8068 gnd.n6517 gnd.n1174 585
R8069 gnd.n6519 gnd.n6518 585
R8070 gnd.n6520 gnd.n1173 585
R8071 gnd.n6522 gnd.n6521 585
R8072 gnd.n6524 gnd.n1171 585
R8073 gnd.n6526 gnd.n6525 585
R8074 gnd.n6527 gnd.n1170 585
R8075 gnd.n6529 gnd.n6528 585
R8076 gnd.n6531 gnd.n1168 585
R8077 gnd.n6533 gnd.n6532 585
R8078 gnd.n6534 gnd.n1167 585
R8079 gnd.n6536 gnd.n6535 585
R8080 gnd.n6538 gnd.n1165 585
R8081 gnd.n6540 gnd.n6539 585
R8082 gnd.n6541 gnd.n1164 585
R8083 gnd.n6543 gnd.n6542 585
R8084 gnd.n6545 gnd.n1163 585
R8085 gnd.n6547 gnd.n6546 585
R8086 gnd.n6548 gnd.n1158 585
R8087 gnd.n6550 gnd.n6549 585
R8088 gnd.n6554 gnd.n877 585
R8089 gnd.n6556 gnd.n6555 585
R8090 gnd.n6557 gnd.n1153 585
R8091 gnd.n6559 gnd.n6558 585
R8092 gnd.n6561 gnd.n1151 585
R8093 gnd.n6563 gnd.n6562 585
R8094 gnd.n6564 gnd.n1150 585
R8095 gnd.n6566 gnd.n6565 585
R8096 gnd.n6568 gnd.n1148 585
R8097 gnd.n6570 gnd.n6569 585
R8098 gnd.n6571 gnd.n1147 585
R8099 gnd.n6573 gnd.n6572 585
R8100 gnd.n6575 gnd.n1145 585
R8101 gnd.n6577 gnd.n6576 585
R8102 gnd.n6578 gnd.n1144 585
R8103 gnd.n6580 gnd.n6579 585
R8104 gnd.n6582 gnd.n1142 585
R8105 gnd.n6584 gnd.n6583 585
R8106 gnd.n6585 gnd.n1141 585
R8107 gnd.n6587 gnd.n6586 585
R8108 gnd.n6589 gnd.n1139 585
R8109 gnd.n6591 gnd.n6590 585
R8110 gnd.n6592 gnd.n1138 585
R8111 gnd.n6594 gnd.n6593 585
R8112 gnd.n6596 gnd.n1136 585
R8113 gnd.n6598 gnd.n6597 585
R8114 gnd.n6599 gnd.n1135 585
R8115 gnd.n6601 gnd.n6600 585
R8116 gnd.n6603 gnd.n1134 585
R8117 gnd.n6605 gnd.n6604 585
R8118 gnd.n6604 gnd.n1102 585
R8119 gnd.n6499 gnd.n1183 585
R8120 gnd.n1183 gnd.n1182 585
R8121 gnd.n6498 gnd.n1110 585
R8122 gnd.n6610 gnd.n1110 585
R8123 gnd.n6497 gnd.n6496 585
R8124 gnd.n6496 gnd.n6495 585
R8125 gnd.n1185 gnd.n1184 585
R8126 gnd.n6493 gnd.n1185 585
R8127 gnd.n6455 gnd.n6454 585
R8128 gnd.n6454 gnd.n1191 585
R8129 gnd.n6456 gnd.n1189 585
R8130 gnd.n6487 gnd.n1189 585
R8131 gnd.n6458 gnd.n6457 585
R8132 gnd.n6459 gnd.n6458 585
R8133 gnd.n6453 gnd.n1201 585
R8134 gnd.n6473 gnd.n1201 585
R8135 gnd.n6452 gnd.n6451 585
R8136 gnd.n6451 gnd.n1199 585
R8137 gnd.n6450 gnd.n1207 585
R8138 gnd.n6467 gnd.n1207 585
R8139 gnd.n6449 gnd.n6448 585
R8140 gnd.n6448 gnd.n6447 585
R8141 gnd.n1219 gnd.n1218 585
R8142 gnd.n1220 gnd.n1219 585
R8143 gnd.n6418 gnd.n6417 585
R8144 gnd.n6419 gnd.n6418 585
R8145 gnd.n6416 gnd.n1229 585
R8146 gnd.n6436 gnd.n1229 585
R8147 gnd.n6415 gnd.n6414 585
R8148 gnd.n6414 gnd.n1227 585
R8149 gnd.n6413 gnd.n1235 585
R8150 gnd.n6427 gnd.n1235 585
R8151 gnd.n6412 gnd.n6411 585
R8152 gnd.n6411 gnd.n6410 585
R8153 gnd.n1247 gnd.n1246 585
R8154 gnd.n1248 gnd.n1247 585
R8155 gnd.n6317 gnd.n6316 585
R8156 gnd.n6316 gnd.n1273 585
R8157 gnd.n6318 gnd.n1257 585
R8158 gnd.n6400 gnd.n1257 585
R8159 gnd.n6320 gnd.n6319 585
R8160 gnd.n6319 gnd.n1255 585
R8161 gnd.n6321 gnd.n1264 585
R8162 gnd.n6391 gnd.n1264 585
R8163 gnd.n6322 gnd.n1296 585
R8164 gnd.n1296 gnd.n1279 585
R8165 gnd.n6324 gnd.n6323 585
R8166 gnd.n6325 gnd.n6324 585
R8167 gnd.n6315 gnd.n1295 585
R8168 gnd.n1295 gnd.n1294 585
R8169 gnd.n6314 gnd.n1287 585
R8170 gnd.n6331 gnd.n1287 585
R8171 gnd.n6313 gnd.n6312 585
R8172 gnd.n6312 gnd.n1285 585
R8173 gnd.n6311 gnd.n1297 585
R8174 gnd.n6311 gnd.n6310 585
R8175 gnd.n6255 gnd.n1298 585
R8176 gnd.n1306 gnd.n1298 585
R8177 gnd.n6256 gnd.n1305 585
R8178 gnd.n6304 gnd.n1305 585
R8179 gnd.n6258 gnd.n6257 585
R8180 gnd.n6259 gnd.n6258 585
R8181 gnd.n6254 gnd.n1331 585
R8182 gnd.n6261 gnd.n1331 585
R8183 gnd.n6253 gnd.n6252 585
R8184 gnd.n6252 gnd.n1314 585
R8185 gnd.n6251 gnd.n1332 585
R8186 gnd.n6251 gnd.n6250 585
R8187 gnd.n6224 gnd.n1325 585
R8188 gnd.n6268 gnd.n1325 585
R8189 gnd.n6226 gnd.n6225 585
R8190 gnd.n6227 gnd.n6226 585
R8191 gnd.n6223 gnd.n1339 585
R8192 gnd.n1339 gnd.n1338 585
R8193 gnd.n6222 gnd.n6221 585
R8194 gnd.n6221 gnd.n6220 585
R8195 gnd.n1341 gnd.n1340 585
R8196 gnd.n1351 gnd.n1341 585
R8197 gnd.n6103 gnd.n1349 585
R8198 gnd.n6213 gnd.n1349 585
R8199 gnd.n6105 gnd.n6104 585
R8200 gnd.n6106 gnd.n6105 585
R8201 gnd.n6102 gnd.n1361 585
R8202 gnd.n6202 gnd.n1361 585
R8203 gnd.n6101 gnd.n6100 585
R8204 gnd.n6100 gnd.n1359 585
R8205 gnd.n6099 gnd.n1367 585
R8206 gnd.n6196 gnd.n1367 585
R8207 gnd.n6098 gnd.n6097 585
R8208 gnd.n6097 gnd.n6096 585
R8209 gnd.n6095 gnd.n1375 585
R8210 gnd.n6170 gnd.n1375 585
R8211 gnd.n6094 gnd.n1382 585
R8212 gnd.n6162 gnd.n1382 585
R8213 gnd.n6093 gnd.n1381 585
R8214 gnd.n6164 gnd.n1381 585
R8215 gnd.n6092 gnd.n6091 585
R8216 gnd.n6091 gnd.n1393 585
R8217 gnd.n1408 gnd.n1407 585
R8218 gnd.n1408 gnd.n1391 585
R8219 gnd.n6127 gnd.n6126 585
R8220 gnd.n6126 gnd.n6125 585
R8221 gnd.n6128 gnd.n1400 585
R8222 gnd.n6142 gnd.n1400 585
R8223 gnd.n6130 gnd.n6129 585
R8224 gnd.n6131 gnd.n6130 585
R8225 gnd.n1406 gnd.n1405 585
R8226 gnd.n6133 gnd.n1405 585
R8227 gnd.n1497 gnd.n1494 585
R8228 gnd.n1497 gnd.n1496 585
R8229 gnd.n1498 gnd.n1493 585
R8230 gnd.n1498 gnd.n1425 585
R8231 gnd.n5168 gnd.n5167 585
R8232 gnd.n5168 gnd.n1999 585
R8233 gnd.n2898 gnd.n2897 585
R8234 gnd.n2898 gnd.n583 585
R8235 gnd.n2894 gnd.n2792 585
R8236 gnd.n2792 gnd.n593 585
R8237 gnd.n2893 gnd.n2892 585
R8238 gnd.n2892 gnd.n604 585
R8239 gnd.n2891 gnd.n2795 585
R8240 gnd.n2891 gnd.n602 585
R8241 gnd.n2890 gnd.n2831 585
R8242 gnd.n2890 gnd.n2889 585
R8243 gnd.n2797 gnd.n2796 585
R8244 gnd.n2796 gnd.n610 585
R8245 gnd.n2826 gnd.n2825 585
R8246 gnd.n2825 gnd.n620 585
R8247 gnd.n2824 gnd.n2799 585
R8248 gnd.n2824 gnd.n618 585
R8249 gnd.n2823 gnd.n2822 585
R8250 gnd.n2823 gnd.n629 585
R8251 gnd.n2801 gnd.n2800 585
R8252 gnd.n2800 gnd.n626 585
R8253 gnd.n2818 gnd.n2817 585
R8254 gnd.n2817 gnd.n637 585
R8255 gnd.n2816 gnd.n2803 585
R8256 gnd.n2816 gnd.n635 585
R8257 gnd.n2815 gnd.n2814 585
R8258 gnd.n2815 gnd.n646 585
R8259 gnd.n2805 gnd.n2804 585
R8260 gnd.n2804 gnd.n643 585
R8261 gnd.n2810 gnd.n2809 585
R8262 gnd.n2809 gnd.n654 585
R8263 gnd.n2808 gnd.n2806 585
R8264 gnd.n2808 gnd.n652 585
R8265 gnd.n2807 gnd.n940 585
R8266 gnd.n2807 gnd.n663 585
R8267 gnd.n6840 gnd.n938 585
R8268 gnd.n938 gnd.n660 585
R8269 gnd.n6842 gnd.n6841 585
R8270 gnd.n6843 gnd.n6842 585
R8271 gnd.n6823 gnd.n937 585
R8272 gnd.n937 gnd.n667 585
R8273 gnd.n6825 gnd.n6824 585
R8274 gnd.n6825 gnd.n678 585
R8275 gnd.n6827 gnd.n6826 585
R8276 gnd.n6826 gnd.n675 585
R8277 gnd.n6829 gnd.n6828 585
R8278 gnd.n6829 gnd.n685 585
R8279 gnd.n6831 gnd.n6830 585
R8280 gnd.n6830 gnd.n682 585
R8281 gnd.n6833 gnd.n6832 585
R8282 gnd.n6833 gnd.n694 585
R8283 gnd.n6834 gnd.n947 585
R8284 gnd.n6834 gnd.n691 585
R8285 gnd.n6836 gnd.n6835 585
R8286 gnd.n6835 gnd.n702 585
R8287 gnd.n6822 gnd.n946 585
R8288 gnd.n6822 gnd.n699 585
R8289 gnd.n6821 gnd.n6820 585
R8290 gnd.n6821 gnd.n711 585
R8291 gnd.n949 gnd.n948 585
R8292 gnd.n948 gnd.n708 585
R8293 gnd.n6816 gnd.n6815 585
R8294 gnd.n6815 gnd.n720 585
R8295 gnd.n6814 gnd.n951 585
R8296 gnd.n6814 gnd.n717 585
R8297 gnd.n6813 gnd.n6751 585
R8298 gnd.n6813 gnd.n6812 585
R8299 gnd.n953 gnd.n952 585
R8300 gnd.n952 gnd.n726 585
R8301 gnd.n6747 gnd.n6746 585
R8302 gnd.n6746 gnd.n737 585
R8303 gnd.n6745 gnd.n955 585
R8304 gnd.n6745 gnd.n734 585
R8305 gnd.n6744 gnd.n6743 585
R8306 gnd.n6744 gnd.n746 585
R8307 gnd.n957 gnd.n956 585
R8308 gnd.n956 gnd.n743 585
R8309 gnd.n6739 gnd.n6738 585
R8310 gnd.n6738 gnd.n755 585
R8311 gnd.n6737 gnd.n959 585
R8312 gnd.n6737 gnd.n752 585
R8313 gnd.n6736 gnd.n6735 585
R8314 gnd.n6736 gnd.n764 585
R8315 gnd.n961 gnd.n960 585
R8316 gnd.n960 gnd.n761 585
R8317 gnd.n6731 gnd.n6730 585
R8318 gnd.n6730 gnd.n773 585
R8319 gnd.n6729 gnd.n963 585
R8320 gnd.n6729 gnd.n770 585
R8321 gnd.n6728 gnd.n6727 585
R8322 gnd.n6728 gnd.n908 585
R8323 gnd.n965 gnd.n964 585
R8324 gnd.n964 gnd.n779 585
R8325 gnd.n6723 gnd.n6722 585
R8326 gnd.n6722 gnd.n789 585
R8327 gnd.n6721 gnd.n967 585
R8328 gnd.n6721 gnd.n786 585
R8329 gnd.n6720 gnd.n6719 585
R8330 gnd.n6720 gnd.n861 585
R8331 gnd.n969 gnd.n968 585
R8332 gnd.n968 gnd.n833 585
R8333 gnd.n6715 gnd.n6714 585
R8334 gnd.n6714 gnd.n6713 585
R8335 gnd.n972 gnd.n971 585
R8336 gnd.n6712 gnd.n972 585
R8337 gnd.n6684 gnd.n6683 585
R8338 gnd.n6684 gnd.n973 585
R8339 gnd.n6687 gnd.n6680 585
R8340 gnd.n6687 gnd.n6686 585
R8341 gnd.n6689 gnd.n6688 585
R8342 gnd.n6688 gnd.n1041 585
R8343 gnd.n6690 gnd.n1053 585
R8344 gnd.n1053 gnd.n1040 585
R8345 gnd.n6692 gnd.n6691 585
R8346 gnd.n6693 gnd.n6692 585
R8347 gnd.n1054 gnd.n1052 585
R8348 gnd.n1052 gnd.n1049 585
R8349 gnd.n6674 gnd.n6673 585
R8350 gnd.n6673 gnd.n6672 585
R8351 gnd.n1057 gnd.n1056 585
R8352 gnd.n1066 gnd.n1057 585
R8353 gnd.n6648 gnd.n1078 585
R8354 gnd.n1078 gnd.n1065 585
R8355 gnd.n6650 gnd.n6649 585
R8356 gnd.n6651 gnd.n6650 585
R8357 gnd.n1079 gnd.n1077 585
R8358 gnd.n1077 gnd.n1074 585
R8359 gnd.n6643 gnd.n6642 585
R8360 gnd.n6642 gnd.n6641 585
R8361 gnd.n1082 gnd.n1081 585
R8362 gnd.n1091 gnd.n1082 585
R8363 gnd.n6618 gnd.n1104 585
R8364 gnd.n1104 gnd.n1090 585
R8365 gnd.n6620 gnd.n6619 585
R8366 gnd.n6621 gnd.n6620 585
R8367 gnd.n1105 gnd.n1103 585
R8368 gnd.n1103 gnd.n1099 585
R8369 gnd.n6613 gnd.n6612 585
R8370 gnd.n6612 gnd.n6611 585
R8371 gnd.n1108 gnd.n1107 585
R8372 gnd.n6494 gnd.n1108 585
R8373 gnd.n1216 gnd.n1215 585
R8374 gnd.n6354 gnd.n1216 585
R8375 gnd.n6462 gnd.n6461 585
R8376 gnd.n6461 gnd.n6460 585
R8377 gnd.n6463 gnd.n1209 585
R8378 gnd.n1209 gnd.n1202 585
R8379 gnd.n6465 gnd.n6464 585
R8380 gnd.n6466 gnd.n6465 585
R8381 gnd.n1210 gnd.n1208 585
R8382 gnd.n6446 gnd.n1208 585
R8383 gnd.n6422 gnd.n6421 585
R8384 gnd.n6421 gnd.n6420 585
R8385 gnd.n6423 gnd.n1238 585
R8386 gnd.n1244 gnd.n1238 585
R8387 gnd.n6425 gnd.n6424 585
R8388 gnd.n6426 gnd.n6425 585
R8389 gnd.n1239 gnd.n1237 585
R8390 gnd.n1237 gnd.n1234 585
R8391 gnd.n6385 gnd.n6384 585
R8392 gnd.n6384 gnd.n6383 585
R8393 gnd.n6386 gnd.n1267 585
R8394 gnd.n1267 gnd.n1258 585
R8395 gnd.n6388 gnd.n6387 585
R8396 gnd.n6389 gnd.n6388 585
R8397 gnd.n1268 gnd.n1266 585
R8398 gnd.n1266 gnd.n1263 585
R8399 gnd.n6295 gnd.n6294 585
R8400 gnd.n6295 gnd.n1292 585
R8401 gnd.n6296 gnd.n6290 585
R8402 gnd.n6296 gnd.n1288 585
R8403 gnd.n6299 gnd.n6298 585
R8404 gnd.n6298 gnd.n6297 585
R8405 gnd.n6300 gnd.n1309 585
R8406 gnd.n1309 gnd.n1299 585
R8407 gnd.n6302 gnd.n6301 585
R8408 gnd.n6303 gnd.n6302 585
R8409 gnd.n1310 gnd.n1308 585
R8410 gnd.n6260 gnd.n1308 585
R8411 gnd.n6284 gnd.n6283 585
R8412 gnd.n6283 gnd.n6282 585
R8413 gnd.n1313 gnd.n1312 585
R8414 gnd.n1326 gnd.n1313 585
R8415 gnd.n6184 gnd.n6180 585
R8416 gnd.n6180 gnd.n1323 585
R8417 gnd.n6186 gnd.n6185 585
R8418 gnd.n6186 gnd.n1343 585
R8419 gnd.n6188 gnd.n6179 585
R8420 gnd.n6188 gnd.n6187 585
R8421 gnd.n6190 gnd.n6189 585
R8422 gnd.n6189 gnd.n1348 585
R8423 gnd.n6191 gnd.n1370 585
R8424 gnd.n1370 gnd.n1362 585
R8425 gnd.n6193 gnd.n6192 585
R8426 gnd.n6194 gnd.n6193 585
R8427 gnd.n1371 gnd.n1369 585
R8428 gnd.n1369 gnd.n1366 585
R8429 gnd.n6173 gnd.n6172 585
R8430 gnd.n6172 gnd.n6171 585
R8431 gnd.n1374 gnd.n1373 585
R8432 gnd.n6163 gnd.n1374 585
R8433 gnd.n6150 gnd.n6149 585
R8434 gnd.n6151 gnd.n6150 585
R8435 gnd.n1395 gnd.n1394 585
R8436 gnd.n6124 gnd.n1394 585
R8437 gnd.n6145 gnd.n6144 585
R8438 gnd.n6144 gnd.n6143 585
R8439 gnd.n1398 gnd.n1397 585
R8440 gnd.n6132 gnd.n1398 585
R8441 gnd.n6068 gnd.n1427 585
R8442 gnd.n1427 gnd.n1415 585
R8443 gnd.n6070 gnd.n6069 585
R8444 gnd.n6071 gnd.n6070 585
R8445 gnd.n1428 gnd.n1426 585
R8446 gnd.n1426 gnd.n1423 585
R8447 gnd.n6063 gnd.n6062 585
R8448 gnd.n6062 gnd.n6061 585
R8449 gnd.n1431 gnd.n1430 585
R8450 gnd.n5874 gnd.n1431 585
R8451 gnd.n5857 gnd.n1645 585
R8452 gnd.n1645 gnd.n1634 585
R8453 gnd.n5859 gnd.n5858 585
R8454 gnd.n5860 gnd.n5859 585
R8455 gnd.n1646 gnd.n1644 585
R8456 gnd.n1644 gnd.n1642 585
R8457 gnd.n5852 gnd.n5851 585
R8458 gnd.n5851 gnd.n5850 585
R8459 gnd.n1649 gnd.n1648 585
R8460 gnd.n1650 gnd.n1649 585
R8461 gnd.n5837 gnd.n5836 585
R8462 gnd.n5838 gnd.n5837 585
R8463 gnd.n1659 gnd.n1658 585
R8464 gnd.n1658 gnd.n1656 585
R8465 gnd.n5832 gnd.n5831 585
R8466 gnd.n5831 gnd.n5830 585
R8467 gnd.n1662 gnd.n1661 585
R8468 gnd.n1663 gnd.n1662 585
R8469 gnd.n5817 gnd.n5816 585
R8470 gnd.n5818 gnd.n5817 585
R8471 gnd.n1671 gnd.n1670 585
R8472 gnd.n1670 gnd.n1668 585
R8473 gnd.n5812 gnd.n5811 585
R8474 gnd.n5811 gnd.n5810 585
R8475 gnd.n1674 gnd.n1673 585
R8476 gnd.n1675 gnd.n1674 585
R8477 gnd.n5547 gnd.n5546 585
R8478 gnd.n5546 gnd.n5545 585
R8479 gnd.n5548 gnd.n5539 585
R8480 gnd.n5544 gnd.n5539 585
R8481 gnd.n5551 gnd.n5549 585
R8482 gnd.n5551 gnd.n5550 585
R8483 gnd.n5552 gnd.n5538 585
R8484 gnd.n5552 gnd.n1603 585
R8485 gnd.n5554 gnd.n5553 585
R8486 gnd.n5553 gnd.n1601 585
R8487 gnd.n5555 gnd.n5441 585
R8488 gnd.n5441 gnd.n1613 585
R8489 gnd.n5557 gnd.n5556 585
R8490 gnd.n5558 gnd.n5557 585
R8491 gnd.n5442 gnd.n5440 585
R8492 gnd.n5440 gnd.n1762 585
R8493 gnd.n5532 gnd.n5531 585
R8494 gnd.n5531 gnd.n1760 585
R8495 gnd.n5530 gnd.n5444 585
R8496 gnd.n5530 gnd.n1772 585
R8497 gnd.n5529 gnd.n5528 585
R8498 gnd.n5529 gnd.n1769 585
R8499 gnd.n5446 gnd.n5445 585
R8500 gnd.n5445 gnd.n1782 585
R8501 gnd.n5524 gnd.n5523 585
R8502 gnd.n5523 gnd.n1779 585
R8503 gnd.n5522 gnd.n5448 585
R8504 gnd.n5522 gnd.n1791 585
R8505 gnd.n5521 gnd.n5520 585
R8506 gnd.n5521 gnd.n1788 585
R8507 gnd.n5450 gnd.n5449 585
R8508 gnd.n5449 gnd.n1800 585
R8509 gnd.n5516 gnd.n5515 585
R8510 gnd.n5515 gnd.n1797 585
R8511 gnd.n5514 gnd.n5452 585
R8512 gnd.n5514 gnd.n1808 585
R8513 gnd.n5513 gnd.n5475 585
R8514 gnd.n5513 gnd.n5512 585
R8515 gnd.n5454 gnd.n5453 585
R8516 gnd.n5453 gnd.n1817 585
R8517 gnd.n5471 gnd.n5470 585
R8518 gnd.n5470 gnd.n1814 585
R8519 gnd.n5469 gnd.n5456 585
R8520 gnd.n5469 gnd.n1826 585
R8521 gnd.n5468 gnd.n5467 585
R8522 gnd.n5468 gnd.n1823 585
R8523 gnd.n5458 gnd.n5457 585
R8524 gnd.n5457 gnd.n1835 585
R8525 gnd.n5463 gnd.n5462 585
R8526 gnd.n5462 gnd.n1832 585
R8527 gnd.n5461 gnd.n5460 585
R8528 gnd.n5461 gnd.n1884 585
R8529 gnd.n1873 gnd.n1872 585
R8530 gnd.n1878 gnd.n1873 585
R8531 gnd.n5626 gnd.n5625 585
R8532 gnd.n5625 gnd.n5624 585
R8533 gnd.n5628 gnd.n1870 585
R8534 gnd.n1874 gnd.n1870 585
R8535 gnd.n5630 gnd.n5629 585
R8536 gnd.n5631 gnd.n5630 585
R8537 gnd.n5193 gnd.n1869 585
R8538 gnd.n1869 gnd.n1862 585
R8539 gnd.n5195 gnd.n5194 585
R8540 gnd.n5195 gnd.n1859 585
R8541 gnd.n5197 gnd.n5196 585
R8542 gnd.n5196 gnd.n1850 585
R8543 gnd.n5198 gnd.n5191 585
R8544 gnd.n5191 gnd.n1847 585
R8545 gnd.n5201 gnd.n5200 585
R8546 gnd.n5201 gnd.n1904 585
R8547 gnd.n5202 gnd.n5190 585
R8548 gnd.n5202 gnd.n1912 585
R8549 gnd.n5204 gnd.n5203 585
R8550 gnd.n5203 gnd.n1910 585
R8551 gnd.n5205 gnd.n5184 585
R8552 gnd.n5184 gnd.n1938 585
R8553 gnd.n5207 gnd.n5206 585
R8554 gnd.n5207 gnd.n1924 585
R8555 gnd.n5208 gnd.n5183 585
R8556 gnd.n5208 gnd.n1921 585
R8557 gnd.n5210 gnd.n5209 585
R8558 gnd.n5209 gnd.n1944 585
R8559 gnd.n5211 gnd.n5178 585
R8560 gnd.n5178 gnd.n1952 585
R8561 gnd.n5213 gnd.n5212 585
R8562 gnd.n5213 gnd.n1950 585
R8563 gnd.n5214 gnd.n5177 585
R8564 gnd.n5214 gnd.n1963 585
R8565 gnd.n5216 gnd.n5215 585
R8566 gnd.n5215 gnd.n1960 585
R8567 gnd.n5217 gnd.n2219 585
R8568 gnd.n2219 gnd.n1972 585
R8569 gnd.n5219 gnd.n5218 585
R8570 gnd.n5220 gnd.n5219 585
R8571 gnd.n2220 gnd.n2218 585
R8572 gnd.n2218 gnd.n1981 585
R8573 gnd.n5171 gnd.n5170 585
R8574 gnd.n5170 gnd.n1978 585
R8575 gnd.n5169 gnd.n2222 585
R8576 gnd.n5169 gnd.n1990 585
R8577 gnd.n1045 gnd.n1043 585
R8578 gnd.n6685 gnd.n1043 585
R8579 gnd.n6702 gnd.n6701 585
R8580 gnd.n6703 gnd.n6702 585
R8581 gnd.n1044 gnd.n1042 585
R8582 gnd.n1051 gnd.n1042 585
R8583 gnd.n6696 gnd.n6695 585
R8584 gnd.n6695 gnd.n6694 585
R8585 gnd.n1048 gnd.n1047 585
R8586 gnd.n6671 gnd.n1048 585
R8587 gnd.n1070 gnd.n1068 585
R8588 gnd.n1068 gnd.n1058 585
R8589 gnd.n6660 gnd.n6659 585
R8590 gnd.n6661 gnd.n6660 585
R8591 gnd.n1069 gnd.n1067 585
R8592 gnd.n1076 gnd.n1067 585
R8593 gnd.n6654 gnd.n6653 585
R8594 gnd.n6653 gnd.n6652 585
R8595 gnd.n1073 gnd.n1072 585
R8596 gnd.n6640 gnd.n1073 585
R8597 gnd.n1095 gnd.n1093 585
R8598 gnd.n1093 gnd.n1083 585
R8599 gnd.n6630 gnd.n6629 585
R8600 gnd.n6631 gnd.n6630 585
R8601 gnd.n1094 gnd.n1092 585
R8602 gnd.n1101 gnd.n1092 585
R8603 gnd.n6624 gnd.n6623 585
R8604 gnd.n6623 gnd.n6622 585
R8605 gnd.n1098 gnd.n1097 585
R8606 gnd.n1111 gnd.n1098 585
R8607 gnd.n6480 gnd.n6479 585
R8608 gnd.n6479 gnd.n1109 585
R8609 gnd.n1195 gnd.n1193 585
R8610 gnd.n6355 gnd.n1193 585
R8611 gnd.n6485 gnd.n6484 585
R8612 gnd.n6486 gnd.n6485 585
R8613 gnd.n1194 gnd.n1192 585
R8614 gnd.n1217 gnd.n1192 585
R8615 gnd.n6476 gnd.n6475 585
R8616 gnd.n6475 gnd.n6474 585
R8617 gnd.n1198 gnd.n1197 585
R8618 gnd.n1206 gnd.n1198 585
R8619 gnd.n6444 gnd.n6443 585
R8620 gnd.n6445 gnd.n6444 585
R8621 gnd.n1223 gnd.n1222 585
R8622 gnd.n1245 gnd.n1222 585
R8623 gnd.n6439 gnd.n6438 585
R8624 gnd.n6438 gnd.n6437 585
R8625 gnd.n1226 gnd.n1225 585
R8626 gnd.n6427 gnd.n1226 585
R8627 gnd.n6408 gnd.n6407 585
R8628 gnd.n6409 gnd.n6408 585
R8629 gnd.n1251 gnd.n1250 585
R8630 gnd.n6382 gnd.n1250 585
R8631 gnd.n6403 gnd.n6402 585
R8632 gnd.n6402 gnd.n6401 585
R8633 gnd.n1254 gnd.n1253 585
R8634 gnd.n6390 gnd.n1254 585
R8635 gnd.n6339 gnd.n6338 585
R8636 gnd.n6340 gnd.n6339 585
R8637 gnd.n1281 gnd.n1280 585
R8638 gnd.n1293 gnd.n1280 585
R8639 gnd.n6334 gnd.n6333 585
R8640 gnd.n6333 gnd.n6332 585
R8641 gnd.n1284 gnd.n1283 585
R8642 gnd.n1300 gnd.n1284 585
R8643 gnd.n6275 gnd.n6274 585
R8644 gnd.n6274 gnd.n1307 585
R8645 gnd.n1319 gnd.n1317 585
R8646 gnd.n1317 gnd.n1304 585
R8647 gnd.n6280 gnd.n6279 585
R8648 gnd.n6281 gnd.n6280 585
R8649 gnd.n1318 gnd.n1316 585
R8650 gnd.n6249 gnd.n1316 585
R8651 gnd.n6271 gnd.n6270 585
R8652 gnd.n6270 gnd.n6269 585
R8653 gnd.n1322 gnd.n1321 585
R8654 gnd.n6228 gnd.n1322 585
R8655 gnd.n1355 gnd.n1353 585
R8656 gnd.n1353 gnd.n1342 585
R8657 gnd.n6211 gnd.n6210 585
R8658 gnd.n6212 gnd.n6211 585
R8659 gnd.n1354 gnd.n1352 585
R8660 gnd.n6106 gnd.n1352 585
R8661 gnd.n6205 gnd.n6204 585
R8662 gnd.n6204 gnd.n6203 585
R8663 gnd.n1358 gnd.n1357 585
R8664 gnd.n6195 gnd.n1358 585
R8665 gnd.n1387 gnd.n1385 585
R8666 gnd.n1385 gnd.n1376 585
R8667 gnd.n6160 gnd.n6159 585
R8668 gnd.n6161 gnd.n6160 585
R8669 gnd.n1386 gnd.n1384 585
R8670 gnd.n1384 gnd.n1380 585
R8671 gnd.n6154 gnd.n6153 585
R8672 gnd.n6153 gnd.n6152 585
R8673 gnd.n1390 gnd.n1389 585
R8674 gnd.n6123 gnd.n1390 585
R8675 gnd.n1419 gnd.n1417 585
R8676 gnd.n1417 gnd.n1399 585
R8677 gnd.n6080 gnd.n6079 585
R8678 gnd.n6081 gnd.n6080 585
R8679 gnd.n1418 gnd.n1416 585
R8680 gnd.n1495 gnd.n1416 585
R8681 gnd.n6074 gnd.n6073 585
R8682 gnd.n6073 gnd.n6072 585
R8683 gnd.n1422 gnd.n1421 585
R8684 gnd.n6060 gnd.n1422 585
R8685 gnd.n5878 gnd.n5877 585
R8686 gnd.n5877 gnd.n1432 585
R8687 gnd.n5881 gnd.n5876 585
R8688 gnd.n5876 gnd.n5875 585
R8689 gnd.n5882 gnd.n1633 585
R8690 gnd.n1643 gnd.n1633 585
R8691 gnd.n5883 gnd.n1632 585
R8692 gnd.n5861 gnd.n1632 585
R8693 gnd.n5848 gnd.n1630 585
R8694 gnd.n5849 gnd.n5848 585
R8695 gnd.n5887 gnd.n1629 585
R8696 gnd.n5847 gnd.n1629 585
R8697 gnd.n5888 gnd.n1628 585
R8698 gnd.n1657 gnd.n1628 585
R8699 gnd.n5889 gnd.n1627 585
R8700 gnd.n5839 gnd.n1627 585
R8701 gnd.n5828 gnd.n1625 585
R8702 gnd.n5829 gnd.n5828 585
R8703 gnd.n5893 gnd.n1624 585
R8704 gnd.n5827 gnd.n1624 585
R8705 gnd.n5894 gnd.n1623 585
R8706 gnd.n1669 gnd.n1623 585
R8707 gnd.n5895 gnd.n1622 585
R8708 gnd.n5819 gnd.n1622 585
R8709 gnd.n5807 gnd.n5806 585
R8710 gnd.n5805 gnd.n1689 585
R8711 gnd.n1691 gnd.n1688 585
R8712 gnd.n5809 gnd.n1688 585
R8713 gnd.n5798 gnd.n1705 585
R8714 gnd.n5797 gnd.n1706 585
R8715 gnd.n1708 gnd.n1707 585
R8716 gnd.n5790 gnd.n1716 585
R8717 gnd.n5789 gnd.n1717 585
R8718 gnd.n1727 gnd.n1718 585
R8719 gnd.n5782 gnd.n1728 585
R8720 gnd.n5781 gnd.n1729 585
R8721 gnd.n1731 gnd.n1730 585
R8722 gnd.n5774 gnd.n1739 585
R8723 gnd.n5773 gnd.n1740 585
R8724 gnd.n1749 gnd.n1741 585
R8725 gnd.n5764 gnd.n1750 585
R8726 gnd.n5763 gnd.n1751 585
R8727 gnd.n5762 gnd.n1752 585
R8728 gnd.n5735 gnd.n1753 585
R8729 gnd.n5758 gnd.n5736 585
R8730 gnd.n5757 gnd.n5737 585
R8731 gnd.n5756 gnd.n5738 585
R8732 gnd.n5744 gnd.n5739 585
R8733 gnd.n5752 gnd.n5745 585
R8734 gnd.n5751 gnd.n5746 585
R8735 gnd.n5750 gnd.n5747 585
R8736 gnd.n5748 gnd.n1667 585
R8737 gnd.n6706 gnd.n993 585
R8738 gnd.n6685 gnd.n993 585
R8739 gnd.n6705 gnd.n6704 585
R8740 gnd.n6704 gnd.n6703 585
R8741 gnd.n1039 gnd.n1038 585
R8742 gnd.n1051 gnd.n1039 585
R8743 gnd.n1061 gnd.n1050 585
R8744 gnd.n6694 gnd.n1050 585
R8745 gnd.n6670 gnd.n6669 585
R8746 gnd.n6671 gnd.n6670 585
R8747 gnd.n1060 gnd.n1059 585
R8748 gnd.n1059 gnd.n1058 585
R8749 gnd.n6663 gnd.n6662 585
R8750 gnd.n6662 gnd.n6661 585
R8751 gnd.n1064 gnd.n1063 585
R8752 gnd.n1076 gnd.n1064 585
R8753 gnd.n1086 gnd.n1075 585
R8754 gnd.n6652 gnd.n1075 585
R8755 gnd.n6639 gnd.n6638 585
R8756 gnd.n6640 gnd.n6639 585
R8757 gnd.n1085 gnd.n1084 585
R8758 gnd.n1084 gnd.n1083 585
R8759 gnd.n6633 gnd.n6632 585
R8760 gnd.n6632 gnd.n6631 585
R8761 gnd.n1089 gnd.n1088 585
R8762 gnd.n1101 gnd.n1089 585
R8763 gnd.n6359 gnd.n1100 585
R8764 gnd.n6622 gnd.n1100 585
R8765 gnd.n6362 gnd.n6358 585
R8766 gnd.n6358 gnd.n1111 585
R8767 gnd.n6363 gnd.n6357 585
R8768 gnd.n6357 gnd.n1109 585
R8769 gnd.n6364 gnd.n6356 585
R8770 gnd.n6356 gnd.n6355 585
R8771 gnd.n6352 gnd.n1190 585
R8772 gnd.n6486 gnd.n1190 585
R8773 gnd.n6368 gnd.n6351 585
R8774 gnd.n6351 gnd.n1217 585
R8775 gnd.n6369 gnd.n1200 585
R8776 gnd.n6474 gnd.n1200 585
R8777 gnd.n6370 gnd.n6350 585
R8778 gnd.n6350 gnd.n1206 585
R8779 gnd.n6348 gnd.n1221 585
R8780 gnd.n6445 gnd.n1221 585
R8781 gnd.n6374 gnd.n6347 585
R8782 gnd.n6347 gnd.n1245 585
R8783 gnd.n6375 gnd.n1228 585
R8784 gnd.n6437 gnd.n1228 585
R8785 gnd.n6376 gnd.n1236 585
R8786 gnd.n6427 gnd.n1236 585
R8787 gnd.n1275 gnd.n1249 585
R8788 gnd.n6409 gnd.n1249 585
R8789 gnd.n6381 gnd.n6380 585
R8790 gnd.n6382 gnd.n6381 585
R8791 gnd.n1274 gnd.n1256 585
R8792 gnd.n6401 gnd.n1256 585
R8793 gnd.n6343 gnd.n1265 585
R8794 gnd.n6390 gnd.n1265 585
R8795 gnd.n6342 gnd.n6341 585
R8796 gnd.n6341 gnd.n6340 585
R8797 gnd.n1278 gnd.n1277 585
R8798 gnd.n1293 gnd.n1278 585
R8799 gnd.n6237 gnd.n1286 585
R8800 gnd.n6332 gnd.n1286 585
R8801 gnd.n6241 gnd.n6236 585
R8802 gnd.n6236 gnd.n1300 585
R8803 gnd.n6242 gnd.n6235 585
R8804 gnd.n6235 gnd.n1307 585
R8805 gnd.n6243 gnd.n6234 585
R8806 gnd.n6234 gnd.n1304 585
R8807 gnd.n1334 gnd.n1315 585
R8808 gnd.n6281 gnd.n1315 585
R8809 gnd.n6248 gnd.n6247 585
R8810 gnd.n6249 gnd.n6248 585
R8811 gnd.n1333 gnd.n1324 585
R8812 gnd.n6269 gnd.n1324 585
R8813 gnd.n6230 gnd.n6229 585
R8814 gnd.n6229 gnd.n6228 585
R8815 gnd.n1337 gnd.n1336 585
R8816 gnd.n1342 gnd.n1337 585
R8817 gnd.n6109 gnd.n1350 585
R8818 gnd.n6212 gnd.n1350 585
R8819 gnd.n6110 gnd.n6107 585
R8820 gnd.n6107 gnd.n6106 585
R8821 gnd.n6111 gnd.n1360 585
R8822 gnd.n6203 gnd.n1360 585
R8823 gnd.n6089 gnd.n1368 585
R8824 gnd.n6195 gnd.n1368 585
R8825 gnd.n6115 gnd.n6088 585
R8826 gnd.n6088 gnd.n1376 585
R8827 gnd.n6116 gnd.n1383 585
R8828 gnd.n6161 gnd.n1383 585
R8829 gnd.n6117 gnd.n6087 585
R8830 gnd.n6087 gnd.n1380 585
R8831 gnd.n1411 gnd.n1392 585
R8832 gnd.n6152 gnd.n1392 585
R8833 gnd.n6122 gnd.n6121 585
R8834 gnd.n6123 gnd.n6122 585
R8835 gnd.n1410 gnd.n1409 585
R8836 gnd.n1409 gnd.n1399 585
R8837 gnd.n6083 gnd.n6082 585
R8838 gnd.n6082 gnd.n6081 585
R8839 gnd.n1414 gnd.n1413 585
R8840 gnd.n1495 gnd.n1414 585
R8841 gnd.n5867 gnd.n1424 585
R8842 gnd.n6072 gnd.n1424 585
R8843 gnd.n5868 gnd.n1433 585
R8844 gnd.n6060 gnd.n1433 585
R8845 gnd.n1638 gnd.n1636 585
R8846 gnd.n1636 gnd.n1432 585
R8847 gnd.n5873 gnd.n5872 585
R8848 gnd.n5875 gnd.n5873 585
R8849 gnd.n1637 gnd.n1635 585
R8850 gnd.n1643 gnd.n1635 585
R8851 gnd.n5863 gnd.n5862 585
R8852 gnd.n5862 gnd.n5861 585
R8853 gnd.n1641 gnd.n1640 585
R8854 gnd.n5849 gnd.n1641 585
R8855 gnd.n5846 gnd.n5845 585
R8856 gnd.n5847 gnd.n5846 585
R8857 gnd.n1652 gnd.n1651 585
R8858 gnd.n1657 gnd.n1651 585
R8859 gnd.n5841 gnd.n5840 585
R8860 gnd.n5840 gnd.n5839 585
R8861 gnd.n1655 gnd.n1654 585
R8862 gnd.n5829 gnd.n1655 585
R8863 gnd.n5826 gnd.n5825 585
R8864 gnd.n5827 gnd.n5826 585
R8865 gnd.n1665 gnd.n1664 585
R8866 gnd.n1669 gnd.n1664 585
R8867 gnd.n5821 gnd.n5820 585
R8868 gnd.n5820 gnd.n5819 585
R8869 gnd.n6710 gnd.n6709 585
R8870 gnd.n6711 gnd.n6710 585
R8871 gnd.n994 gnd.n992 585
R8872 gnd.n1034 gnd.n1033 585
R8873 gnd.n1032 gnd.n1031 585
R8874 gnd.n1029 gnd.n1000 585
R8875 gnd.n999 gnd.n998 585
R8876 gnd.n1025 gnd.n1024 585
R8877 gnd.n1023 gnd.n1022 585
R8878 gnd.n1021 gnd.n1004 585
R8879 gnd.n1003 gnd.n1002 585
R8880 gnd.n1010 gnd.n1009 585
R8881 gnd.n1008 gnd.n1007 585
R8882 gnd.n985 gnd.n829 585
R8883 gnd.n6973 gnd.n828 585
R8884 gnd.n6974 gnd.n827 585
R8885 gnd.n982 gnd.n821 585
R8886 gnd.n6981 gnd.n820 585
R8887 gnd.n6982 gnd.n819 585
R8888 gnd.n980 gnd.n813 585
R8889 gnd.n6989 gnd.n812 585
R8890 gnd.n6990 gnd.n811 585
R8891 gnd.n977 gnd.n805 585
R8892 gnd.n6997 gnd.n804 585
R8893 gnd.n6998 gnd.n803 585
R8894 gnd.n975 gnd.n797 585
R8895 gnd.n7005 gnd.n796 585
R8896 gnd.n7006 gnd.n795 585
R8897 gnd.n6604 gnd.n1113 521.33
R8898 gnd.n6501 gnd.n1183 521.33
R8899 gnd.n1499 gnd.n1498 521.33
R8900 gnd.n6057 gnd.n1465 521.33
R8901 gnd.n3375 gnd.n3374 468.854
R8902 gnd.n1490 gnd.t119 347.526
R8903 gnd.n1159 gnd.t155 347.526
R8904 gnd.n1488 gnd.t172 347.526
R8905 gnd.n1154 gnd.t187 347.526
R8906 gnd.n4396 gnd.t145 323.425
R8907 gnd.n3648 gnd.t141 323.425
R8908 gnd.n4292 gnd.n4266 289.615
R8909 gnd.n4329 gnd.n4303 289.615
R8910 gnd.n4153 gnd.n4127 289.615
R8911 gnd.n4190 gnd.n4164 289.615
R8912 gnd.n4222 gnd.n4196 289.615
R8913 gnd.n4259 gnd.n4233 289.615
R8914 gnd.n458 gnd.n432 289.615
R8915 gnd.n421 gnd.n395 289.615
R8916 gnd.n319 gnd.n293 289.615
R8917 gnd.n282 gnd.n256 289.615
R8918 gnd.n388 gnd.n362 289.615
R8919 gnd.n351 gnd.n325 289.615
R8920 gnd.n4995 gnd.n4969 289.615
R8921 gnd.n4963 gnd.n4937 289.615
R8922 gnd.n4931 gnd.n4905 289.615
R8923 gnd.n4900 gnd.n4874 289.615
R8924 gnd.n4868 gnd.n4842 289.615
R8925 gnd.n4836 gnd.n4810 289.615
R8926 gnd.n4804 gnd.n4778 289.615
R8927 gnd.n4773 gnd.n4747 289.615
R8928 gnd.n122 gnd.n96 289.615
R8929 gnd.n90 gnd.n64 289.615
R8930 gnd.n58 gnd.n32 289.615
R8931 gnd.n27 gnd.n1 289.615
R8932 gnd.n249 gnd.n223 289.615
R8933 gnd.n217 gnd.n191 289.615
R8934 gnd.n185 gnd.n159 289.615
R8935 gnd.n154 gnd.n128 289.615
R8936 gnd.n5741 gnd.t203 279.217
R8937 gnd.n3971 gnd.t196 279.217
R8938 gnd.n3674 gnd.t127 279.217
R8939 gnd.n7235 gnd.t159 279.217
R8940 gnd.n6968 gnd.t135 279.217
R8941 gnd.n1743 gnd.t131 279.217
R8942 gnd.n880 gnd.t109 279.217
R8943 gnd.n900 gnd.t200 279.217
R8944 gnd.n571 gnd.t169 279.217
R8945 gnd.n535 gnd.t184 279.217
R8946 gnd.n2122 gnd.t149 279.217
R8947 gnd.n2051 gnd.t123 279.217
R8948 gnd.n5243 gnd.t152 279.217
R8949 gnd.n1594 gnd.t163 279.217
R8950 gnd.n1559 gnd.t181 279.217
R8951 gnd.n996 gnd.t210 279.217
R8952 gnd.n1472 gnd.t180 260.649
R8953 gnd.n1126 gnd.t209 260.649
R8954 gnd.n6059 gnd.n6058 256.663
R8955 gnd.n6059 gnd.n1434 256.663
R8956 gnd.n6059 gnd.n1435 256.663
R8957 gnd.n6059 gnd.n1436 256.663
R8958 gnd.n6059 gnd.n1437 256.663
R8959 gnd.n6059 gnd.n1438 256.663
R8960 gnd.n6059 gnd.n1439 256.663
R8961 gnd.n6059 gnd.n1440 256.663
R8962 gnd.n6059 gnd.n1441 256.663
R8963 gnd.n6059 gnd.n1442 256.663
R8964 gnd.n6059 gnd.n1443 256.663
R8965 gnd.n6059 gnd.n1444 256.663
R8966 gnd.n6059 gnd.n1445 256.663
R8967 gnd.n6059 gnd.n1446 256.663
R8968 gnd.n6059 gnd.n1447 256.663
R8969 gnd.n5999 gnd.n5998 256.663
R8970 gnd.n6059 gnd.n1448 256.663
R8971 gnd.n6059 gnd.n1449 256.663
R8972 gnd.n6059 gnd.n1450 256.663
R8973 gnd.n6059 gnd.n1451 256.663
R8974 gnd.n6059 gnd.n1452 256.663
R8975 gnd.n6059 gnd.n1453 256.663
R8976 gnd.n6059 gnd.n1454 256.663
R8977 gnd.n6059 gnd.n1455 256.663
R8978 gnd.n6059 gnd.n1456 256.663
R8979 gnd.n6059 gnd.n1457 256.663
R8980 gnd.n6059 gnd.n1458 256.663
R8981 gnd.n6059 gnd.n1459 256.663
R8982 gnd.n6059 gnd.n1460 256.663
R8983 gnd.n6059 gnd.n1461 256.663
R8984 gnd.n6059 gnd.n1462 256.663
R8985 gnd.n6502 gnd.n1102 256.663
R8986 gnd.n1181 gnd.n1102 256.663
R8987 gnd.n6509 gnd.n1102 256.663
R8988 gnd.n1178 gnd.n1102 256.663
R8989 gnd.n6516 gnd.n1102 256.663
R8990 gnd.n1175 gnd.n1102 256.663
R8991 gnd.n6523 gnd.n1102 256.663
R8992 gnd.n1172 gnd.n1102 256.663
R8993 gnd.n6530 gnd.n1102 256.663
R8994 gnd.n1169 gnd.n1102 256.663
R8995 gnd.n6537 gnd.n1102 256.663
R8996 gnd.n1166 gnd.n1102 256.663
R8997 gnd.n6544 gnd.n1102 256.663
R8998 gnd.n1162 gnd.n1102 256.663
R8999 gnd.n6551 gnd.n1102 256.663
R9000 gnd.n6552 gnd.n877 256.663
R9001 gnd.n6553 gnd.n1102 256.663
R9002 gnd.n1157 gnd.n1102 256.663
R9003 gnd.n6560 gnd.n1102 256.663
R9004 gnd.n1152 gnd.n1102 256.663
R9005 gnd.n6567 gnd.n1102 256.663
R9006 gnd.n1149 gnd.n1102 256.663
R9007 gnd.n6574 gnd.n1102 256.663
R9008 gnd.n1146 gnd.n1102 256.663
R9009 gnd.n6581 gnd.n1102 256.663
R9010 gnd.n1143 gnd.n1102 256.663
R9011 gnd.n6588 gnd.n1102 256.663
R9012 gnd.n1140 gnd.n1102 256.663
R9013 gnd.n6595 gnd.n1102 256.663
R9014 gnd.n1137 gnd.n1102 256.663
R9015 gnd.n6602 gnd.n1102 256.663
R9016 gnd.n5273 gnd.n2012 242.672
R9017 gnd.n5271 gnd.n2012 242.672
R9018 gnd.n5265 gnd.n2012 242.672
R9019 gnd.n5263 gnd.n2012 242.672
R9020 gnd.n5257 gnd.n2012 242.672
R9021 gnd.n5255 gnd.n2012 242.672
R9022 gnd.n5249 gnd.n2012 242.672
R9023 gnd.n5247 gnd.n2012 242.672
R9024 gnd.n5767 gnd.n1567 242.672
R9025 gnd.n1745 gnd.n1567 242.672
R9026 gnd.n1734 gnd.n1567 242.672
R9027 gnd.n1723 gnd.n1567 242.672
R9028 gnd.n1720 gnd.n1567 242.672
R9029 gnd.n1711 gnd.n1567 242.672
R9030 gnd.n1701 gnd.n1567 242.672
R9031 gnd.n1698 gnd.n1567 242.672
R9032 gnd.n6964 gnd.n850 242.672
R9033 gnd.n6964 gnd.n852 242.672
R9034 gnd.n6964 gnd.n854 242.672
R9035 gnd.n6964 gnd.n855 242.672
R9036 gnd.n6964 gnd.n857 242.672
R9037 gnd.n6964 gnd.n859 242.672
R9038 gnd.n6964 gnd.n860 242.672
R9039 gnd.n6966 gnd.n6964 242.672
R9040 gnd.n7237 gnd.n502 242.672
R9041 gnd.n7233 gnd.n502 242.672
R9042 gnd.n7230 gnd.n502 242.672
R9043 gnd.n7225 gnd.n502 242.672
R9044 gnd.n7222 gnd.n502 242.672
R9045 gnd.n7217 gnd.n502 242.672
R9046 gnd.n7214 gnd.n502 242.672
R9047 gnd.n7209 gnd.n502 242.672
R9048 gnd.n4026 gnd.n3935 242.672
R9049 gnd.n3939 gnd.n3935 242.672
R9050 gnd.n4019 gnd.n3935 242.672
R9051 gnd.n4013 gnd.n3935 242.672
R9052 gnd.n4011 gnd.n3935 242.672
R9053 gnd.n4005 gnd.n3935 242.672
R9054 gnd.n4003 gnd.n3935 242.672
R9055 gnd.n3997 gnd.n3935 242.672
R9056 gnd.n3995 gnd.n3935 242.672
R9057 gnd.n3989 gnd.n3935 242.672
R9058 gnd.n3987 gnd.n3935 242.672
R9059 gnd.n3980 gnd.n3935 242.672
R9060 gnd.n3978 gnd.n3935 242.672
R9061 gnd.n5116 gnd.n3619 242.672
R9062 gnd.n5116 gnd.n3618 242.672
R9063 gnd.n5116 gnd.n3617 242.672
R9064 gnd.n5116 gnd.n3616 242.672
R9065 gnd.n5116 gnd.n3615 242.672
R9066 gnd.n5116 gnd.n3614 242.672
R9067 gnd.n5116 gnd.n3613 242.672
R9068 gnd.n5116 gnd.n3612 242.672
R9069 gnd.n5116 gnd.n3611 242.672
R9070 gnd.n5116 gnd.n3610 242.672
R9071 gnd.n5116 gnd.n3609 242.672
R9072 gnd.n5116 gnd.n3608 242.672
R9073 gnd.n5116 gnd.n3607 242.672
R9074 gnd.n4430 gnd.n4429 242.672
R9075 gnd.n4430 gnd.n4371 242.672
R9076 gnd.n4430 gnd.n4372 242.672
R9077 gnd.n4430 gnd.n4373 242.672
R9078 gnd.n4430 gnd.n4374 242.672
R9079 gnd.n4430 gnd.n4375 242.672
R9080 gnd.n4430 gnd.n4376 242.672
R9081 gnd.n4430 gnd.n4377 242.672
R9082 gnd.n5116 gnd.n3620 242.672
R9083 gnd.n5116 gnd.n3621 242.672
R9084 gnd.n5116 gnd.n3622 242.672
R9085 gnd.n5116 gnd.n3623 242.672
R9086 gnd.n5116 gnd.n3624 242.672
R9087 gnd.n5116 gnd.n3625 242.672
R9088 gnd.n5116 gnd.n3626 242.672
R9089 gnd.n5116 gnd.n5115 242.672
R9090 gnd.n2086 gnd.n2012 242.672
R9091 gnd.n2094 gnd.n2012 242.672
R9092 gnd.n2096 gnd.n2012 242.672
R9093 gnd.n2104 gnd.n2012 242.672
R9094 gnd.n2106 gnd.n2012 242.672
R9095 gnd.n2114 gnd.n2012 242.672
R9096 gnd.n2116 gnd.n2012 242.672
R9097 gnd.n2127 gnd.n2012 242.672
R9098 gnd.n2129 gnd.n2012 242.672
R9099 gnd.n2137 gnd.n2012 242.672
R9100 gnd.n2139 gnd.n2012 242.672
R9101 gnd.n2147 gnd.n2012 242.672
R9102 gnd.n2149 gnd.n2012 242.672
R9103 gnd.n2157 gnd.n2012 242.672
R9104 gnd.n2159 gnd.n2012 242.672
R9105 gnd.n2168 gnd.n2012 242.672
R9106 gnd.n2171 gnd.n2012 242.672
R9107 gnd.n1599 gnd.n1567 242.672
R9108 gnd.n5967 gnd.n1567 242.672
R9109 gnd.n1589 gnd.n1567 242.672
R9110 gnd.n5974 gnd.n1567 242.672
R9111 gnd.n1582 gnd.n1567 242.672
R9112 gnd.n5981 gnd.n1567 242.672
R9113 gnd.n1575 gnd.n1567 242.672
R9114 gnd.n5988 gnd.n1567 242.672
R9115 gnd.n5991 gnd.n1567 242.672
R9116 gnd.n1567 gnd.n1566 242.672
R9117 gnd.n5997 gnd.n1561 242.672
R9118 gnd.n5927 gnd.n1567 242.672
R9119 gnd.n5933 gnd.n1567 242.672
R9120 gnd.n5926 gnd.n1567 242.672
R9121 gnd.n5940 gnd.n1567 242.672
R9122 gnd.n5919 gnd.n1567 242.672
R9123 gnd.n5947 gnd.n1567 242.672
R9124 gnd.n5950 gnd.n1567 242.672
R9125 gnd.n6964 gnd.n6963 242.672
R9126 gnd.n6964 gnd.n834 242.672
R9127 gnd.n6964 gnd.n835 242.672
R9128 gnd.n6964 gnd.n836 242.672
R9129 gnd.n6964 gnd.n837 242.672
R9130 gnd.n6964 gnd.n838 242.672
R9131 gnd.n6964 gnd.n839 242.672
R9132 gnd.n6937 gnd.n878 242.672
R9133 gnd.n6964 gnd.n840 242.672
R9134 gnd.n6964 gnd.n841 242.672
R9135 gnd.n6964 gnd.n842 242.672
R9136 gnd.n6964 gnd.n843 242.672
R9137 gnd.n6964 gnd.n844 242.672
R9138 gnd.n6964 gnd.n845 242.672
R9139 gnd.n6964 gnd.n846 242.672
R9140 gnd.n6964 gnd.n847 242.672
R9141 gnd.n6964 gnd.n848 242.672
R9142 gnd.n6964 gnd.n849 242.672
R9143 gnd.n568 gnd.n502 242.672
R9144 gnd.n7294 gnd.n502 242.672
R9145 gnd.n564 gnd.n502 242.672
R9146 gnd.n7301 gnd.n502 242.672
R9147 gnd.n557 gnd.n502 242.672
R9148 gnd.n7308 gnd.n502 242.672
R9149 gnd.n550 gnd.n502 242.672
R9150 gnd.n7315 gnd.n502 242.672
R9151 gnd.n543 gnd.n502 242.672
R9152 gnd.n7322 gnd.n502 242.672
R9153 gnd.n533 gnd.n502 242.672
R9154 gnd.n7329 gnd.n502 242.672
R9155 gnd.n526 gnd.n502 242.672
R9156 gnd.n7336 gnd.n502 242.672
R9157 gnd.n519 gnd.n502 242.672
R9158 gnd.n7343 gnd.n502 242.672
R9159 gnd.n512 gnd.n502 242.672
R9160 gnd.n5809 gnd.n5808 242.672
R9161 gnd.n5809 gnd.n1676 242.672
R9162 gnd.n5809 gnd.n1677 242.672
R9163 gnd.n5809 gnd.n1678 242.672
R9164 gnd.n5809 gnd.n1679 242.672
R9165 gnd.n5809 gnd.n1680 242.672
R9166 gnd.n5809 gnd.n1681 242.672
R9167 gnd.n5809 gnd.n1682 242.672
R9168 gnd.n5809 gnd.n1683 242.672
R9169 gnd.n5809 gnd.n1684 242.672
R9170 gnd.n5809 gnd.n1685 242.672
R9171 gnd.n5809 gnd.n1686 242.672
R9172 gnd.n5809 gnd.n1687 242.672
R9173 gnd.n6711 gnd.n991 242.672
R9174 gnd.n6711 gnd.n990 242.672
R9175 gnd.n6711 gnd.n989 242.672
R9176 gnd.n6711 gnd.n988 242.672
R9177 gnd.n6711 gnd.n987 242.672
R9178 gnd.n6711 gnd.n986 242.672
R9179 gnd.n6711 gnd.n984 242.672
R9180 gnd.n6711 gnd.n983 242.672
R9181 gnd.n6711 gnd.n981 242.672
R9182 gnd.n6711 gnd.n979 242.672
R9183 gnd.n6711 gnd.n978 242.672
R9184 gnd.n6711 gnd.n976 242.672
R9185 gnd.n6711 gnd.n974 242.672
R9186 gnd.n509 gnd.n505 240.244
R9187 gnd.n7345 gnd.n7344 240.244
R9188 gnd.n7342 gnd.n513 240.244
R9189 gnd.n7338 gnd.n7337 240.244
R9190 gnd.n7335 gnd.n520 240.244
R9191 gnd.n7331 gnd.n7330 240.244
R9192 gnd.n7328 gnd.n527 240.244
R9193 gnd.n7324 gnd.n7323 240.244
R9194 gnd.n7321 gnd.n534 240.244
R9195 gnd.n7317 gnd.n7316 240.244
R9196 gnd.n7314 gnd.n544 240.244
R9197 gnd.n7310 gnd.n7309 240.244
R9198 gnd.n7307 gnd.n551 240.244
R9199 gnd.n7303 gnd.n7302 240.244
R9200 gnd.n7300 gnd.n558 240.244
R9201 gnd.n7296 gnd.n7295 240.244
R9202 gnd.n7293 gnd.n565 240.244
R9203 gnd.n904 gnd.n787 240.244
R9204 gnd.n904 gnd.n780 240.244
R9205 gnd.n6893 gnd.n780 240.244
R9206 gnd.n6893 gnd.n771 240.244
R9207 gnd.n6759 gnd.n771 240.244
R9208 gnd.n6759 gnd.n762 240.244
R9209 gnd.n6765 gnd.n762 240.244
R9210 gnd.n6765 gnd.n753 240.244
R9211 gnd.n6769 gnd.n753 240.244
R9212 gnd.n6769 gnd.n744 240.244
R9213 gnd.n6775 gnd.n744 240.244
R9214 gnd.n6775 gnd.n735 240.244
R9215 gnd.n6779 gnd.n735 240.244
R9216 gnd.n6779 gnd.n727 240.244
R9217 gnd.n6810 gnd.n727 240.244
R9218 gnd.n6810 gnd.n718 240.244
R9219 gnd.n6806 gnd.n718 240.244
R9220 gnd.n6806 gnd.n709 240.244
R9221 gnd.n6802 gnd.n709 240.244
R9222 gnd.n6802 gnd.n700 240.244
R9223 gnd.n6798 gnd.n700 240.244
R9224 gnd.n6798 gnd.n692 240.244
R9225 gnd.n6794 gnd.n692 240.244
R9226 gnd.n6794 gnd.n683 240.244
R9227 gnd.n6853 gnd.n683 240.244
R9228 gnd.n6853 gnd.n676 240.244
R9229 gnd.n6849 gnd.n676 240.244
R9230 gnd.n6849 gnd.n668 240.244
R9231 gnd.n6845 gnd.n668 240.244
R9232 gnd.n6845 gnd.n661 240.244
R9233 gnd.n2841 gnd.n661 240.244
R9234 gnd.n2841 gnd.n653 240.244
R9235 gnd.n2845 gnd.n653 240.244
R9236 gnd.n2845 gnd.n644 240.244
R9237 gnd.n2851 gnd.n644 240.244
R9238 gnd.n2851 gnd.n636 240.244
R9239 gnd.n2855 gnd.n636 240.244
R9240 gnd.n2855 gnd.n627 240.244
R9241 gnd.n2861 gnd.n627 240.244
R9242 gnd.n2861 gnd.n619 240.244
R9243 gnd.n2865 gnd.n619 240.244
R9244 gnd.n2865 gnd.n611 240.244
R9245 gnd.n2887 gnd.n611 240.244
R9246 gnd.n2887 gnd.n603 240.244
R9247 gnd.n2883 gnd.n603 240.244
R9248 gnd.n2883 gnd.n594 240.244
R9249 gnd.n2879 gnd.n594 240.244
R9250 gnd.n2879 gnd.n584 240.244
R9251 gnd.n584 gnd.n575 240.244
R9252 gnd.n7284 gnd.n575 240.244
R9253 gnd.n7285 gnd.n7284 240.244
R9254 gnd.n7285 gnd.n501 240.244
R9255 gnd.n6962 gnd.n862 240.244
R9256 gnd.n6958 gnd.n862 240.244
R9257 gnd.n6956 gnd.n6955 240.244
R9258 gnd.n6952 gnd.n6951 240.244
R9259 gnd.n6948 gnd.n6947 240.244
R9260 gnd.n6944 gnd.n6943 240.244
R9261 gnd.n6940 gnd.n6939 240.244
R9262 gnd.n6935 gnd.n6934 240.244
R9263 gnd.n6931 gnd.n6930 240.244
R9264 gnd.n6927 gnd.n6926 240.244
R9265 gnd.n6923 gnd.n6922 240.244
R9266 gnd.n6919 gnd.n6918 240.244
R9267 gnd.n6915 gnd.n6914 240.244
R9268 gnd.n6911 gnd.n6910 240.244
R9269 gnd.n6907 gnd.n6906 240.244
R9270 gnd.n899 gnd.n898 240.244
R9271 gnd.n7016 gnd.n782 240.244
R9272 gnd.n7022 gnd.n782 240.244
R9273 gnd.n7022 gnd.n769 240.244
R9274 gnd.n7032 gnd.n769 240.244
R9275 gnd.n7032 gnd.n765 240.244
R9276 gnd.n7038 gnd.n765 240.244
R9277 gnd.n7038 gnd.n751 240.244
R9278 gnd.n7048 gnd.n751 240.244
R9279 gnd.n7048 gnd.n747 240.244
R9280 gnd.n7054 gnd.n747 240.244
R9281 gnd.n7054 gnd.n733 240.244
R9282 gnd.n7064 gnd.n733 240.244
R9283 gnd.n7064 gnd.n729 240.244
R9284 gnd.n7070 gnd.n729 240.244
R9285 gnd.n7070 gnd.n716 240.244
R9286 gnd.n7080 gnd.n716 240.244
R9287 gnd.n7080 gnd.n712 240.244
R9288 gnd.n7087 gnd.n712 240.244
R9289 gnd.n7087 gnd.n698 240.244
R9290 gnd.n7097 gnd.n698 240.244
R9291 gnd.n7097 gnd.n695 240.244
R9292 gnd.n7103 gnd.n695 240.244
R9293 gnd.n7103 gnd.n681 240.244
R9294 gnd.n7113 gnd.n681 240.244
R9295 gnd.n7113 gnd.n679 240.244
R9296 gnd.n7119 gnd.n679 240.244
R9297 gnd.n7119 gnd.n666 240.244
R9298 gnd.n7129 gnd.n666 240.244
R9299 gnd.n7129 gnd.n664 240.244
R9300 gnd.n7134 gnd.n664 240.244
R9301 gnd.n7134 gnd.n651 240.244
R9302 gnd.n7144 gnd.n651 240.244
R9303 gnd.n7144 gnd.n647 240.244
R9304 gnd.n7150 gnd.n647 240.244
R9305 gnd.n7150 gnd.n634 240.244
R9306 gnd.n7160 gnd.n634 240.244
R9307 gnd.n7160 gnd.n630 240.244
R9308 gnd.n7166 gnd.n630 240.244
R9309 gnd.n7166 gnd.n617 240.244
R9310 gnd.n7176 gnd.n617 240.244
R9311 gnd.n7176 gnd.n613 240.244
R9312 gnd.n7182 gnd.n613 240.244
R9313 gnd.n7182 gnd.n601 240.244
R9314 gnd.n7192 gnd.n601 240.244
R9315 gnd.n7192 gnd.n597 240.244
R9316 gnd.n7198 gnd.n597 240.244
R9317 gnd.n7198 gnd.n582 240.244
R9318 gnd.n7276 gnd.n582 240.244
R9319 gnd.n7276 gnd.n578 240.244
R9320 gnd.n7282 gnd.n578 240.244
R9321 gnd.n7282 gnd.n504 240.244
R9322 gnd.n7352 gnd.n504 240.244
R9323 gnd.n5951 gnd.n1606 240.244
R9324 gnd.n5949 gnd.n5948 240.244
R9325 gnd.n5946 gnd.n5912 240.244
R9326 gnd.n5942 gnd.n5941 240.244
R9327 gnd.n5939 gnd.n5920 240.244
R9328 gnd.n5935 gnd.n5934 240.244
R9329 gnd.n5932 gnd.n5928 240.244
R9330 gnd.n5992 gnd.n1565 240.244
R9331 gnd.n5990 gnd.n5989 240.244
R9332 gnd.n5987 gnd.n1569 240.244
R9333 gnd.n5983 gnd.n5982 240.244
R9334 gnd.n5980 gnd.n1576 240.244
R9335 gnd.n5976 gnd.n5975 240.244
R9336 gnd.n5973 gnd.n1583 240.244
R9337 gnd.n5969 gnd.n5968 240.244
R9338 gnd.n5966 gnd.n1590 240.244
R9339 gnd.n2177 gnd.n2013 240.244
R9340 gnd.n2177 gnd.n2006 240.244
R9341 gnd.n2182 gnd.n2006 240.244
R9342 gnd.n2182 gnd.n1997 240.244
R9343 gnd.n2185 gnd.n1997 240.244
R9344 gnd.n2185 gnd.n1988 240.244
R9345 gnd.n5226 gnd.n1988 240.244
R9346 gnd.n5226 gnd.n1979 240.244
R9347 gnd.n5222 gnd.n1979 240.244
R9348 gnd.n5222 gnd.n1970 240.244
R9349 gnd.n2211 gnd.n1970 240.244
R9350 gnd.n2211 gnd.n1961 240.244
R9351 gnd.n2207 gnd.n1961 240.244
R9352 gnd.n2207 gnd.n1951 240.244
R9353 gnd.n1951 gnd.n1943 240.244
R9354 gnd.n5363 gnd.n1943 240.244
R9355 gnd.n5363 gnd.n1922 240.244
R9356 gnd.n1939 gnd.n1922 240.244
R9357 gnd.n5372 gnd.n1939 240.244
R9358 gnd.n5372 gnd.n1911 240.244
R9359 gnd.n1911 gnd.n1903 240.244
R9360 gnd.n5398 gnd.n1903 240.244
R9361 gnd.n5398 gnd.n1848 240.244
R9362 gnd.n5404 gnd.n1848 240.244
R9363 gnd.n5404 gnd.n1860 240.244
R9364 gnd.n1866 gnd.n1860 240.244
R9365 gnd.n5603 gnd.n1866 240.244
R9366 gnd.n5603 gnd.n5602 240.244
R9367 gnd.n5602 gnd.n1876 240.244
R9368 gnd.n1882 gnd.n1876 240.244
R9369 gnd.n5597 gnd.n1882 240.244
R9370 gnd.n5597 gnd.n1833 240.244
R9371 gnd.n5481 gnd.n1833 240.244
R9372 gnd.n5481 gnd.n1824 240.244
R9373 gnd.n5485 gnd.n1824 240.244
R9374 gnd.n5485 gnd.n1815 240.244
R9375 gnd.n5510 gnd.n1815 240.244
R9376 gnd.n5510 gnd.n1806 240.244
R9377 gnd.n5506 gnd.n1806 240.244
R9378 gnd.n5506 gnd.n1798 240.244
R9379 gnd.n5502 gnd.n1798 240.244
R9380 gnd.n5502 gnd.n1789 240.244
R9381 gnd.n5498 gnd.n1789 240.244
R9382 gnd.n5498 gnd.n1780 240.244
R9383 gnd.n5568 gnd.n1780 240.244
R9384 gnd.n5568 gnd.n1770 240.244
R9385 gnd.n5564 gnd.n1770 240.244
R9386 gnd.n5564 gnd.n1761 240.244
R9387 gnd.n5560 gnd.n1761 240.244
R9388 gnd.n5560 gnd.n1611 240.244
R9389 gnd.n1611 gnd.n1598 240.244
R9390 gnd.n5959 gnd.n1598 240.244
R9391 gnd.n2087 gnd.n2083 240.244
R9392 gnd.n2093 gnd.n2083 240.244
R9393 gnd.n2097 gnd.n2095 240.244
R9394 gnd.n2103 gnd.n2079 240.244
R9395 gnd.n2107 gnd.n2105 240.244
R9396 gnd.n2113 gnd.n2075 240.244
R9397 gnd.n2117 gnd.n2115 240.244
R9398 gnd.n2126 gnd.n2071 240.244
R9399 gnd.n2130 gnd.n2128 240.244
R9400 gnd.n2136 gnd.n2067 240.244
R9401 gnd.n2140 gnd.n2138 240.244
R9402 gnd.n2146 gnd.n2063 240.244
R9403 gnd.n2150 gnd.n2148 240.244
R9404 gnd.n2156 gnd.n2059 240.244
R9405 gnd.n2160 gnd.n2158 240.244
R9406 gnd.n2167 gnd.n2055 240.244
R9407 gnd.n2170 gnd.n2169 240.244
R9408 gnd.n5282 gnd.n2008 240.244
R9409 gnd.n5288 gnd.n2008 240.244
R9410 gnd.n5288 gnd.n1995 240.244
R9411 gnd.n5298 gnd.n1995 240.244
R9412 gnd.n5298 gnd.n1991 240.244
R9413 gnd.n5304 gnd.n1991 240.244
R9414 gnd.n5304 gnd.n1977 240.244
R9415 gnd.n5314 gnd.n1977 240.244
R9416 gnd.n5314 gnd.n1973 240.244
R9417 gnd.n5320 gnd.n1973 240.244
R9418 gnd.n5320 gnd.n1959 240.244
R9419 gnd.n5339 gnd.n1959 240.244
R9420 gnd.n5339 gnd.n1954 240.244
R9421 gnd.n5347 gnd.n1954 240.244
R9422 gnd.n5347 gnd.n1955 240.244
R9423 gnd.n1955 gnd.n1919 240.244
R9424 gnd.n5380 gnd.n1919 240.244
R9425 gnd.n5380 gnd.n1920 240.244
R9426 gnd.n1920 gnd.n1914 240.244
R9427 gnd.n5387 gnd.n1914 240.244
R9428 gnd.n5387 gnd.n1915 240.244
R9429 gnd.n1915 gnd.n1845 240.244
R9430 gnd.n5644 gnd.n1845 240.244
R9431 gnd.n5644 gnd.n1846 240.244
R9432 gnd.n5636 gnd.n1846 240.244
R9433 gnd.n5636 gnd.n5633 240.244
R9434 gnd.n5633 gnd.n1863 240.244
R9435 gnd.n1880 gnd.n1863 240.244
R9436 gnd.n5622 gnd.n1880 240.244
R9437 gnd.n5622 gnd.n5619 240.244
R9438 gnd.n5619 gnd.n1836 240.244
R9439 gnd.n5651 gnd.n1836 240.244
R9440 gnd.n5651 gnd.n1822 240.244
R9441 gnd.n5661 gnd.n1822 240.244
R9442 gnd.n5661 gnd.n1818 240.244
R9443 gnd.n5667 gnd.n1818 240.244
R9444 gnd.n5667 gnd.n1805 240.244
R9445 gnd.n5677 gnd.n1805 240.244
R9446 gnd.n5677 gnd.n1801 240.244
R9447 gnd.n5683 gnd.n1801 240.244
R9448 gnd.n5683 gnd.n1787 240.244
R9449 gnd.n5693 gnd.n1787 240.244
R9450 gnd.n5693 gnd.n1783 240.244
R9451 gnd.n5699 gnd.n1783 240.244
R9452 gnd.n5699 gnd.n1768 240.244
R9453 gnd.n5714 gnd.n1768 240.244
R9454 gnd.n5714 gnd.n1764 240.244
R9455 gnd.n5720 gnd.n1764 240.244
R9456 gnd.n5720 gnd.n1610 240.244
R9457 gnd.n5905 gnd.n1610 240.244
R9458 gnd.n5905 gnd.n1605 240.244
R9459 gnd.n5957 gnd.n1605 240.244
R9460 gnd.n3627 gnd.n3603 240.244
R9461 gnd.n5114 gnd.n3628 240.244
R9462 gnd.n5110 gnd.n5109 240.244
R9463 gnd.n5106 gnd.n5105 240.244
R9464 gnd.n5102 gnd.n5101 240.244
R9465 gnd.n5098 gnd.n5097 240.244
R9466 gnd.n5094 gnd.n5093 240.244
R9467 gnd.n5090 gnd.n5089 240.244
R9468 gnd.n4442 gnd.n3888 240.244
R9469 gnd.n3888 gnd.n3879 240.244
R9470 gnd.n4463 gnd.n3879 240.244
R9471 gnd.n4463 gnd.n3872 240.244
R9472 gnd.n4473 gnd.n3872 240.244
R9473 gnd.n4473 gnd.n3863 240.244
R9474 gnd.n3863 gnd.n3852 240.244
R9475 gnd.n4494 gnd.n3852 240.244
R9476 gnd.n4494 gnd.n3846 240.244
R9477 gnd.n4504 gnd.n3846 240.244
R9478 gnd.n4504 gnd.n3837 240.244
R9479 gnd.n3837 gnd.n3826 240.244
R9480 gnd.n4525 gnd.n3826 240.244
R9481 gnd.n4525 gnd.n3820 240.244
R9482 gnd.n4535 gnd.n3820 240.244
R9483 gnd.n4535 gnd.n3811 240.244
R9484 gnd.n3811 gnd.n3801 240.244
R9485 gnd.n4556 gnd.n3801 240.244
R9486 gnd.n4556 gnd.n3794 240.244
R9487 gnd.n4566 gnd.n3794 240.244
R9488 gnd.n4566 gnd.n3785 240.244
R9489 gnd.n3785 gnd.n3776 240.244
R9490 gnd.n4587 gnd.n3776 240.244
R9491 gnd.n4587 gnd.n3769 240.244
R9492 gnd.n4597 gnd.n3769 240.244
R9493 gnd.n4597 gnd.n3760 240.244
R9494 gnd.n3760 gnd.n3751 240.244
R9495 gnd.n4618 gnd.n3751 240.244
R9496 gnd.n4618 gnd.n3744 240.244
R9497 gnd.n4628 gnd.n3744 240.244
R9498 gnd.n4628 gnd.n3733 240.244
R9499 gnd.n3733 gnd.n3725 240.244
R9500 gnd.n4646 gnd.n3725 240.244
R9501 gnd.n4647 gnd.n4646 240.244
R9502 gnd.n4647 gnd.n3711 240.244
R9503 gnd.n4649 gnd.n3711 240.244
R9504 gnd.n4649 gnd.n3696 240.244
R9505 gnd.n4702 gnd.n3696 240.244
R9506 gnd.n4703 gnd.n4702 240.244
R9507 gnd.n4704 gnd.n4703 240.244
R9508 gnd.n4704 gnd.n3548 240.244
R9509 gnd.n4714 gnd.n3548 240.244
R9510 gnd.n4714 gnd.n3558 240.244
R9511 gnd.n4739 gnd.n3558 240.244
R9512 gnd.n4740 gnd.n4739 240.244
R9513 gnd.n4740 gnd.n3570 240.244
R9514 gnd.n4729 gnd.n3570 240.244
R9515 gnd.n4729 gnd.n3582 240.244
R9516 gnd.n3685 gnd.n3582 240.244
R9517 gnd.n5021 gnd.n3685 240.244
R9518 gnd.n5021 gnd.n3594 240.244
R9519 gnd.n5017 gnd.n3594 240.244
R9520 gnd.n5017 gnd.n3605 240.244
R9521 gnd.n4379 gnd.n4378 240.244
R9522 gnd.n4423 gnd.n4378 240.244
R9523 gnd.n4421 gnd.n4420 240.244
R9524 gnd.n4417 gnd.n4416 240.244
R9525 gnd.n4413 gnd.n4412 240.244
R9526 gnd.n4409 gnd.n4408 240.244
R9527 gnd.n4405 gnd.n4404 240.244
R9528 gnd.n4401 gnd.n4400 240.244
R9529 gnd.n4453 gnd.n3886 240.244
R9530 gnd.n4453 gnd.n3881 240.244
R9531 gnd.n4461 gnd.n3881 240.244
R9532 gnd.n4461 gnd.n3882 240.244
R9533 gnd.n3882 gnd.n3861 240.244
R9534 gnd.n4484 gnd.n3861 240.244
R9535 gnd.n4484 gnd.n3855 240.244
R9536 gnd.n4492 gnd.n3855 240.244
R9537 gnd.n4492 gnd.n3857 240.244
R9538 gnd.n3857 gnd.n3835 240.244
R9539 gnd.n4515 gnd.n3835 240.244
R9540 gnd.n4515 gnd.n3829 240.244
R9541 gnd.n4523 gnd.n3829 240.244
R9542 gnd.n4523 gnd.n3831 240.244
R9543 gnd.n3831 gnd.n3809 240.244
R9544 gnd.n4546 gnd.n3809 240.244
R9545 gnd.n4546 gnd.n3804 240.244
R9546 gnd.n4554 gnd.n3804 240.244
R9547 gnd.n4554 gnd.n3805 240.244
R9548 gnd.n3805 gnd.n3783 240.244
R9549 gnd.n4577 gnd.n3783 240.244
R9550 gnd.n4577 gnd.n3778 240.244
R9551 gnd.n4585 gnd.n3778 240.244
R9552 gnd.n4585 gnd.n3779 240.244
R9553 gnd.n3779 gnd.n3758 240.244
R9554 gnd.n4608 gnd.n3758 240.244
R9555 gnd.n4608 gnd.n3753 240.244
R9556 gnd.n4616 gnd.n3753 240.244
R9557 gnd.n4616 gnd.n3754 240.244
R9558 gnd.n3754 gnd.n3731 240.244
R9559 gnd.n4638 gnd.n3731 240.244
R9560 gnd.n4638 gnd.n3727 240.244
R9561 gnd.n4644 gnd.n3727 240.244
R9562 gnd.n4644 gnd.n3709 240.244
R9563 gnd.n4680 gnd.n3709 240.244
R9564 gnd.n4680 gnd.n3704 240.244
R9565 gnd.n4692 gnd.n3704 240.244
R9566 gnd.n4692 gnd.n3705 240.244
R9567 gnd.n4688 gnd.n3705 240.244
R9568 gnd.n4688 gnd.n3549 240.244
R9569 gnd.n5150 gnd.n3549 240.244
R9570 gnd.n5150 gnd.n3550 240.244
R9571 gnd.n5146 gnd.n3550 240.244
R9572 gnd.n5146 gnd.n3556 240.244
R9573 gnd.n3571 gnd.n3556 240.244
R9574 gnd.n5136 gnd.n3571 240.244
R9575 gnd.n5136 gnd.n3572 240.244
R9576 gnd.n5132 gnd.n3572 240.244
R9577 gnd.n5132 gnd.n3580 240.244
R9578 gnd.n3595 gnd.n3580 240.244
R9579 gnd.n5122 gnd.n3595 240.244
R9580 gnd.n5122 gnd.n3596 240.244
R9581 gnd.n5118 gnd.n3596 240.244
R9582 gnd.n3652 gnd.n3606 240.244
R9583 gnd.n5080 gnd.n5079 240.244
R9584 gnd.n5076 gnd.n5075 240.244
R9585 gnd.n5072 gnd.n5071 240.244
R9586 gnd.n5068 gnd.n5067 240.244
R9587 gnd.n5064 gnd.n5063 240.244
R9588 gnd.n5060 gnd.n5059 240.244
R9589 gnd.n5056 gnd.n5055 240.244
R9590 gnd.n5052 gnd.n5051 240.244
R9591 gnd.n5048 gnd.n5047 240.244
R9592 gnd.n5044 gnd.n5043 240.244
R9593 gnd.n5040 gnd.n5039 240.244
R9594 gnd.n5036 gnd.n5035 240.244
R9595 gnd.n4035 gnd.n3931 240.244
R9596 gnd.n4041 gnd.n3931 240.244
R9597 gnd.n4041 gnd.n3923 240.244
R9598 gnd.n4051 gnd.n3923 240.244
R9599 gnd.n4051 gnd.n3919 240.244
R9600 gnd.n4057 gnd.n3919 240.244
R9601 gnd.n4057 gnd.n3910 240.244
R9602 gnd.n4067 gnd.n3910 240.244
R9603 gnd.n4067 gnd.n3905 240.244
R9604 gnd.n4370 gnd.n3905 240.244
R9605 gnd.n4370 gnd.n3906 240.244
R9606 gnd.n3906 gnd.n3898 240.244
R9607 gnd.n4365 gnd.n3898 240.244
R9608 gnd.n4365 gnd.n3889 240.244
R9609 gnd.n4362 gnd.n3889 240.244
R9610 gnd.n4362 gnd.n4361 240.244
R9611 gnd.n4361 gnd.n3874 240.244
R9612 gnd.n4356 gnd.n3874 240.244
R9613 gnd.n4356 gnd.n3864 240.244
R9614 gnd.n4353 gnd.n3864 240.244
R9615 gnd.n4353 gnd.n4352 240.244
R9616 gnd.n4352 gnd.n3847 240.244
R9617 gnd.n4348 gnd.n3847 240.244
R9618 gnd.n4348 gnd.n3838 240.244
R9619 gnd.n4345 gnd.n3838 240.244
R9620 gnd.n4345 gnd.n4344 240.244
R9621 gnd.n4344 gnd.n3821 240.244
R9622 gnd.n4340 gnd.n3821 240.244
R9623 gnd.n4340 gnd.n3812 240.244
R9624 gnd.n4123 gnd.n3812 240.244
R9625 gnd.n4124 gnd.n4123 240.244
R9626 gnd.n4124 gnd.n3796 240.244
R9627 gnd.n4120 gnd.n3796 240.244
R9628 gnd.n4120 gnd.n3786 240.244
R9629 gnd.n4116 gnd.n3786 240.244
R9630 gnd.n4116 gnd.n4115 240.244
R9631 gnd.n4115 gnd.n3771 240.244
R9632 gnd.n4110 gnd.n3771 240.244
R9633 gnd.n4110 gnd.n3761 240.244
R9634 gnd.n4107 gnd.n3761 240.244
R9635 gnd.n4107 gnd.n4105 240.244
R9636 gnd.n4105 gnd.n3746 240.244
R9637 gnd.n4101 gnd.n3746 240.244
R9638 gnd.n4101 gnd.n3734 240.244
R9639 gnd.n3734 gnd.n3716 240.244
R9640 gnd.n4658 gnd.n3716 240.244
R9641 gnd.n4658 gnd.n3712 240.244
R9642 gnd.n4677 gnd.n3712 240.244
R9643 gnd.n4677 gnd.n3702 240.244
R9644 gnd.n4673 gnd.n3702 240.244
R9645 gnd.n4673 gnd.n3536 240.244
R9646 gnd.n4670 gnd.n3536 240.244
R9647 gnd.n4670 gnd.n3547 240.244
R9648 gnd.n4717 gnd.n3547 240.244
R9649 gnd.n4718 gnd.n4717 240.244
R9650 gnd.n4718 gnd.n3559 240.244
R9651 gnd.n4736 gnd.n3559 240.244
R9652 gnd.n4736 gnd.n3569 240.244
R9653 gnd.n4732 gnd.n3569 240.244
R9654 gnd.n4732 gnd.n4728 240.244
R9655 gnd.n4728 gnd.n3583 240.244
R9656 gnd.n5024 gnd.n3583 240.244
R9657 gnd.n5024 gnd.n3593 240.244
R9658 gnd.n3681 gnd.n3593 240.244
R9659 gnd.n5031 gnd.n3681 240.244
R9660 gnd.n4027 gnd.n4025 240.244
R9661 gnd.n4025 gnd.n4024 240.244
R9662 gnd.n4021 gnd.n4020 240.244
R9663 gnd.n4018 gnd.n3944 240.244
R9664 gnd.n4014 gnd.n4012 240.244
R9665 gnd.n4010 gnd.n3950 240.244
R9666 gnd.n4006 gnd.n4004 240.244
R9667 gnd.n4002 gnd.n3956 240.244
R9668 gnd.n3998 gnd.n3996 240.244
R9669 gnd.n3994 gnd.n3962 240.244
R9670 gnd.n3990 gnd.n3988 240.244
R9671 gnd.n3986 gnd.n3968 240.244
R9672 gnd.n3981 gnd.n3979 240.244
R9673 gnd.n4033 gnd.n3929 240.244
R9674 gnd.n4043 gnd.n3929 240.244
R9675 gnd.n4043 gnd.n3925 240.244
R9676 gnd.n4049 gnd.n3925 240.244
R9677 gnd.n4049 gnd.n3917 240.244
R9678 gnd.n4059 gnd.n3917 240.244
R9679 gnd.n4059 gnd.n3913 240.244
R9680 gnd.n4065 gnd.n3913 240.244
R9681 gnd.n4065 gnd.n3904 240.244
R9682 gnd.n4432 gnd.n3904 240.244
R9683 gnd.n4432 gnd.n3899 240.244
R9684 gnd.n4439 gnd.n3899 240.244
R9685 gnd.n4439 gnd.n3891 240.244
R9686 gnd.n4450 gnd.n3891 240.244
R9687 gnd.n4450 gnd.n3892 240.244
R9688 gnd.n3892 gnd.n3875 240.244
R9689 gnd.n4470 gnd.n3875 240.244
R9690 gnd.n4470 gnd.n3866 240.244
R9691 gnd.n4481 gnd.n3866 240.244
R9692 gnd.n4481 gnd.n3867 240.244
R9693 gnd.n3867 gnd.n3848 240.244
R9694 gnd.n4501 gnd.n3848 240.244
R9695 gnd.n4501 gnd.n3840 240.244
R9696 gnd.n4512 gnd.n3840 240.244
R9697 gnd.n4512 gnd.n3841 240.244
R9698 gnd.n3841 gnd.n3822 240.244
R9699 gnd.n4532 gnd.n3822 240.244
R9700 gnd.n4532 gnd.n3814 240.244
R9701 gnd.n4543 gnd.n3814 240.244
R9702 gnd.n4543 gnd.n3815 240.244
R9703 gnd.n3815 gnd.n3797 240.244
R9704 gnd.n4563 gnd.n3797 240.244
R9705 gnd.n4563 gnd.n3788 240.244
R9706 gnd.n4574 gnd.n3788 240.244
R9707 gnd.n4574 gnd.n3789 240.244
R9708 gnd.n3789 gnd.n3772 240.244
R9709 gnd.n4594 gnd.n3772 240.244
R9710 gnd.n4594 gnd.n3763 240.244
R9711 gnd.n4605 gnd.n3763 240.244
R9712 gnd.n4605 gnd.n3764 240.244
R9713 gnd.n3764 gnd.n3747 240.244
R9714 gnd.n4625 gnd.n3747 240.244
R9715 gnd.n4625 gnd.n3736 240.244
R9716 gnd.n4635 gnd.n3736 240.244
R9717 gnd.n4635 gnd.n3718 240.244
R9718 gnd.n4656 gnd.n3718 240.244
R9719 gnd.n4656 gnd.n3719 240.244
R9720 gnd.n3719 gnd.n3700 240.244
R9721 gnd.n4695 gnd.n3700 240.244
R9722 gnd.n4695 gnd.n3538 240.244
R9723 gnd.n5157 gnd.n3538 240.244
R9724 gnd.n5157 gnd.n3539 240.244
R9725 gnd.n5153 gnd.n3539 240.244
R9726 gnd.n5153 gnd.n3545 240.244
R9727 gnd.n3560 gnd.n3545 240.244
R9728 gnd.n5143 gnd.n3560 240.244
R9729 gnd.n5143 gnd.n3561 240.244
R9730 gnd.n5139 gnd.n3561 240.244
R9731 gnd.n5139 gnd.n3567 240.244
R9732 gnd.n3585 gnd.n3567 240.244
R9733 gnd.n5129 gnd.n3585 240.244
R9734 gnd.n5129 gnd.n3586 240.244
R9735 gnd.n5125 gnd.n3586 240.244
R9736 gnd.n5125 gnd.n3592 240.244
R9737 gnd.n5010 gnd.n3592 240.244
R9738 gnd.n7208 gnd.n7207 240.244
R9739 gnd.n7213 gnd.n7210 240.244
R9740 gnd.n7216 gnd.n7215 240.244
R9741 gnd.n7221 gnd.n7218 240.244
R9742 gnd.n7224 gnd.n7223 240.244
R9743 gnd.n7229 gnd.n7226 240.244
R9744 gnd.n7232 gnd.n7231 240.244
R9745 gnd.n7238 gnd.n7234 240.244
R9746 gnd.n1014 gnd.n788 240.244
R9747 gnd.n1014 gnd.n781 240.244
R9748 gnd.n6891 gnd.n781 240.244
R9749 gnd.n6891 gnd.n772 240.244
R9750 gnd.n913 gnd.n772 240.244
R9751 gnd.n913 gnd.n763 240.244
R9752 gnd.n914 gnd.n763 240.244
R9753 gnd.n914 gnd.n754 240.244
R9754 gnd.n917 gnd.n754 240.244
R9755 gnd.n917 gnd.n745 240.244
R9756 gnd.n918 gnd.n745 240.244
R9757 gnd.n918 gnd.n736 240.244
R9758 gnd.n921 gnd.n736 240.244
R9759 gnd.n921 gnd.n728 240.244
R9760 gnd.n922 gnd.n728 240.244
R9761 gnd.n922 gnd.n719 240.244
R9762 gnd.n925 gnd.n719 240.244
R9763 gnd.n925 gnd.n710 240.244
R9764 gnd.n926 gnd.n710 240.244
R9765 gnd.n926 gnd.n701 240.244
R9766 gnd.n929 gnd.n701 240.244
R9767 gnd.n929 gnd.n693 240.244
R9768 gnd.n930 gnd.n693 240.244
R9769 gnd.n930 gnd.n684 240.244
R9770 gnd.n6855 gnd.n684 240.244
R9771 gnd.n6855 gnd.n677 240.244
R9772 gnd.n677 gnd.n468 240.244
R9773 gnd.n469 gnd.n468 240.244
R9774 gnd.n470 gnd.n469 240.244
R9775 gnd.n662 gnd.n470 240.244
R9776 gnd.n662 gnd.n473 240.244
R9777 gnd.n474 gnd.n473 240.244
R9778 gnd.n475 gnd.n474 240.244
R9779 gnd.n645 gnd.n475 240.244
R9780 gnd.n645 gnd.n478 240.244
R9781 gnd.n479 gnd.n478 240.244
R9782 gnd.n480 gnd.n479 240.244
R9783 gnd.n628 gnd.n480 240.244
R9784 gnd.n628 gnd.n483 240.244
R9785 gnd.n484 gnd.n483 240.244
R9786 gnd.n485 gnd.n484 240.244
R9787 gnd.n612 gnd.n485 240.244
R9788 gnd.n612 gnd.n488 240.244
R9789 gnd.n489 gnd.n488 240.244
R9790 gnd.n490 gnd.n489 240.244
R9791 gnd.n595 gnd.n490 240.244
R9792 gnd.n595 gnd.n493 240.244
R9793 gnd.n494 gnd.n493 240.244
R9794 gnd.n495 gnd.n494 240.244
R9795 gnd.n576 gnd.n495 240.244
R9796 gnd.n576 gnd.n498 240.244
R9797 gnd.n7354 gnd.n498 240.244
R9798 gnd.n851 gnd.n792 240.244
R9799 gnd.n800 gnd.n799 240.244
R9800 gnd.n853 gnd.n807 240.244
R9801 gnd.n856 gnd.n808 240.244
R9802 gnd.n816 gnd.n815 240.244
R9803 gnd.n858 gnd.n823 240.244
R9804 gnd.n6965 gnd.n824 240.244
R9805 gnd.n6967 gnd.n832 240.244
R9806 gnd.n7014 gnd.n778 240.244
R9807 gnd.n7024 gnd.n778 240.244
R9808 gnd.n7024 gnd.n774 240.244
R9809 gnd.n7030 gnd.n774 240.244
R9810 gnd.n7030 gnd.n760 240.244
R9811 gnd.n7040 gnd.n760 240.244
R9812 gnd.n7040 gnd.n756 240.244
R9813 gnd.n7046 gnd.n756 240.244
R9814 gnd.n7046 gnd.n742 240.244
R9815 gnd.n7056 gnd.n742 240.244
R9816 gnd.n7056 gnd.n738 240.244
R9817 gnd.n7062 gnd.n738 240.244
R9818 gnd.n7062 gnd.n725 240.244
R9819 gnd.n7072 gnd.n725 240.244
R9820 gnd.n7072 gnd.n721 240.244
R9821 gnd.n7078 gnd.n721 240.244
R9822 gnd.n7078 gnd.n707 240.244
R9823 gnd.n7089 gnd.n707 240.244
R9824 gnd.n7089 gnd.n703 240.244
R9825 gnd.n7095 gnd.n703 240.244
R9826 gnd.n7095 gnd.n690 240.244
R9827 gnd.n7105 gnd.n690 240.244
R9828 gnd.n7105 gnd.n686 240.244
R9829 gnd.n7111 gnd.n686 240.244
R9830 gnd.n7111 gnd.n674 240.244
R9831 gnd.n7121 gnd.n674 240.244
R9832 gnd.n7121 gnd.n669 240.244
R9833 gnd.n7127 gnd.n669 240.244
R9834 gnd.n7127 gnd.n659 240.244
R9835 gnd.n7136 gnd.n659 240.244
R9836 gnd.n7136 gnd.n655 240.244
R9837 gnd.n7142 gnd.n655 240.244
R9838 gnd.n7142 gnd.n642 240.244
R9839 gnd.n7152 gnd.n642 240.244
R9840 gnd.n7152 gnd.n638 240.244
R9841 gnd.n7158 gnd.n638 240.244
R9842 gnd.n7158 gnd.n625 240.244
R9843 gnd.n7168 gnd.n625 240.244
R9844 gnd.n7168 gnd.n621 240.244
R9845 gnd.n7174 gnd.n621 240.244
R9846 gnd.n7174 gnd.n609 240.244
R9847 gnd.n7184 gnd.n609 240.244
R9848 gnd.n7184 gnd.n605 240.244
R9849 gnd.n7190 gnd.n605 240.244
R9850 gnd.n7190 gnd.n592 240.244
R9851 gnd.n7200 gnd.n592 240.244
R9852 gnd.n7200 gnd.n586 240.244
R9853 gnd.n7274 gnd.n586 240.244
R9854 gnd.n7274 gnd.n587 240.244
R9855 gnd.n587 gnd.n577 240.244
R9856 gnd.n7205 gnd.n577 240.244
R9857 gnd.n7205 gnd.n503 240.244
R9858 gnd.n1697 gnd.n1695 240.244
R9859 gnd.n1700 gnd.n1699 240.244
R9860 gnd.n1710 gnd.n1702 240.244
R9861 gnd.n1713 gnd.n1712 240.244
R9862 gnd.n1722 gnd.n1721 240.244
R9863 gnd.n1733 gnd.n1724 240.244
R9864 gnd.n1736 gnd.n1735 240.244
R9865 gnd.n1747 gnd.n1746 240.244
R9866 gnd.n5237 gnd.n2014 240.244
R9867 gnd.n5237 gnd.n2007 240.244
R9868 gnd.n5234 gnd.n2007 240.244
R9869 gnd.n5234 gnd.n1998 240.244
R9870 gnd.n5231 gnd.n1998 240.244
R9871 gnd.n5231 gnd.n1989 240.244
R9872 gnd.n5228 gnd.n1989 240.244
R9873 gnd.n5228 gnd.n1980 240.244
R9874 gnd.n2217 gnd.n1980 240.244
R9875 gnd.n2217 gnd.n1971 240.244
R9876 gnd.n2213 gnd.n1971 240.244
R9877 gnd.n2213 gnd.n1962 240.244
R9878 gnd.n1962 gnd.n1949 240.244
R9879 gnd.n5349 gnd.n1949 240.244
R9880 gnd.n5349 gnd.n1945 240.244
R9881 gnd.n5361 gnd.n1945 240.244
R9882 gnd.n5361 gnd.n1923 240.244
R9883 gnd.n5357 gnd.n1923 240.244
R9884 gnd.n5357 gnd.n1909 240.244
R9885 gnd.n5389 gnd.n1909 240.244
R9886 gnd.n5389 gnd.n1905 240.244
R9887 gnd.n5396 gnd.n1905 240.244
R9888 gnd.n5396 gnd.n1849 240.244
R9889 gnd.n5406 gnd.n1849 240.244
R9890 gnd.n5406 gnd.n1861 240.244
R9891 gnd.n1867 gnd.n1861 240.244
R9892 gnd.n5413 gnd.n1867 240.244
R9893 gnd.n5414 gnd.n5413 240.244
R9894 gnd.n5414 gnd.n1877 240.244
R9895 gnd.n1883 gnd.n1877 240.244
R9896 gnd.n5595 gnd.n1883 240.244
R9897 gnd.n5595 gnd.n1834 240.244
R9898 gnd.n5420 gnd.n1834 240.244
R9899 gnd.n5420 gnd.n1825 240.244
R9900 gnd.n5421 gnd.n1825 240.244
R9901 gnd.n5421 gnd.n1816 240.244
R9902 gnd.n5424 gnd.n1816 240.244
R9903 gnd.n5424 gnd.n1807 240.244
R9904 gnd.n5425 gnd.n1807 240.244
R9905 gnd.n5425 gnd.n1799 240.244
R9906 gnd.n5428 gnd.n1799 240.244
R9907 gnd.n5428 gnd.n1790 240.244
R9908 gnd.n5429 gnd.n1790 240.244
R9909 gnd.n5429 gnd.n1781 240.244
R9910 gnd.n5570 gnd.n1781 240.244
R9911 gnd.n5570 gnd.n1771 240.244
R9912 gnd.n1771 gnd.n1758 240.244
R9913 gnd.n5722 gnd.n1758 240.244
R9914 gnd.n5722 gnd.n1759 240.244
R9915 gnd.n1759 gnd.n1612 240.244
R9916 gnd.n5729 gnd.n1612 240.244
R9917 gnd.n5729 gnd.n1602 240.244
R9918 gnd.n5274 gnd.n5272 240.244
R9919 gnd.n5270 gnd.n2018 240.244
R9920 gnd.n5266 gnd.n5264 240.244
R9921 gnd.n5262 gnd.n2024 240.244
R9922 gnd.n5258 gnd.n5256 240.244
R9923 gnd.n5254 gnd.n2030 240.244
R9924 gnd.n5250 gnd.n5248 240.244
R9925 gnd.n5246 gnd.n2036 240.244
R9926 gnd.n5280 gnd.n2004 240.244
R9927 gnd.n5290 gnd.n2004 240.244
R9928 gnd.n5290 gnd.n2000 240.244
R9929 gnd.n5296 gnd.n2000 240.244
R9930 gnd.n5296 gnd.n1986 240.244
R9931 gnd.n5306 gnd.n1986 240.244
R9932 gnd.n5306 gnd.n1982 240.244
R9933 gnd.n5312 gnd.n1982 240.244
R9934 gnd.n5312 gnd.n1969 240.244
R9935 gnd.n5322 gnd.n1969 240.244
R9936 gnd.n5322 gnd.n1964 240.244
R9937 gnd.n5337 gnd.n1964 240.244
R9938 gnd.n5337 gnd.n1965 240.244
R9939 gnd.n1965 gnd.n1953 240.244
R9940 gnd.n5332 gnd.n1953 240.244
R9941 gnd.n5332 gnd.n1925 240.244
R9942 gnd.n5378 gnd.n1925 240.244
R9943 gnd.n5378 gnd.n1926 240.244
R9944 gnd.n5374 gnd.n1926 240.244
R9945 gnd.n5374 gnd.n1913 240.244
R9946 gnd.n1935 gnd.n1913 240.244
R9947 gnd.n1935 gnd.n1851 240.244
R9948 gnd.n5642 gnd.n1851 240.244
R9949 gnd.n5642 gnd.n1852 240.244
R9950 gnd.n5638 gnd.n1852 240.244
R9951 gnd.n5638 gnd.n1858 240.244
R9952 gnd.n5610 gnd.n1858 240.244
R9953 gnd.n5611 gnd.n5610 240.244
R9954 gnd.n5611 gnd.n1879 240.244
R9955 gnd.n5617 gnd.n1879 240.244
R9956 gnd.n5617 gnd.n1831 240.244
R9957 gnd.n5653 gnd.n1831 240.244
R9958 gnd.n5653 gnd.n1827 240.244
R9959 gnd.n5659 gnd.n1827 240.244
R9960 gnd.n5659 gnd.n1813 240.244
R9961 gnd.n5669 gnd.n1813 240.244
R9962 gnd.n5669 gnd.n1809 240.244
R9963 gnd.n5675 gnd.n1809 240.244
R9964 gnd.n5675 gnd.n1796 240.244
R9965 gnd.n5685 gnd.n1796 240.244
R9966 gnd.n5685 gnd.n1792 240.244
R9967 gnd.n5691 gnd.n1792 240.244
R9968 gnd.n5691 gnd.n1778 240.244
R9969 gnd.n5701 gnd.n1778 240.244
R9970 gnd.n5701 gnd.n1773 240.244
R9971 gnd.n5712 gnd.n1773 240.244
R9972 gnd.n5712 gnd.n1774 240.244
R9973 gnd.n1774 gnd.n1763 240.244
R9974 gnd.n1763 gnd.n1614 240.244
R9975 gnd.n5903 gnd.n1614 240.244
R9976 gnd.n5903 gnd.n1615 240.244
R9977 gnd.n1615 gnd.n1604 240.244
R9978 gnd.n3372 gnd.n2322 240.244
R9979 gnd.n3372 gnd.n2324 240.244
R9980 gnd.n3368 gnd.n2324 240.244
R9981 gnd.n3368 gnd.n2330 240.244
R9982 gnd.n3364 gnd.n2330 240.244
R9983 gnd.n3364 gnd.n2332 240.244
R9984 gnd.n3360 gnd.n2332 240.244
R9985 gnd.n3360 gnd.n2338 240.244
R9986 gnd.n3356 gnd.n2338 240.244
R9987 gnd.n3356 gnd.n2340 240.244
R9988 gnd.n3352 gnd.n2340 240.244
R9989 gnd.n3352 gnd.n2346 240.244
R9990 gnd.n3348 gnd.n2346 240.244
R9991 gnd.n3348 gnd.n2348 240.244
R9992 gnd.n3344 gnd.n2348 240.244
R9993 gnd.n3344 gnd.n2354 240.244
R9994 gnd.n3340 gnd.n2354 240.244
R9995 gnd.n3340 gnd.n2356 240.244
R9996 gnd.n3336 gnd.n2356 240.244
R9997 gnd.n3336 gnd.n2362 240.244
R9998 gnd.n3332 gnd.n2362 240.244
R9999 gnd.n3332 gnd.n2364 240.244
R10000 gnd.n3328 gnd.n2364 240.244
R10001 gnd.n3328 gnd.n2370 240.244
R10002 gnd.n3324 gnd.n2370 240.244
R10003 gnd.n3324 gnd.n2372 240.244
R10004 gnd.n3320 gnd.n2372 240.244
R10005 gnd.n3320 gnd.n2378 240.244
R10006 gnd.n3316 gnd.n2378 240.244
R10007 gnd.n3316 gnd.n2380 240.244
R10008 gnd.n3312 gnd.n2380 240.244
R10009 gnd.n3312 gnd.n2386 240.244
R10010 gnd.n3308 gnd.n2386 240.244
R10011 gnd.n3308 gnd.n2388 240.244
R10012 gnd.n3304 gnd.n2388 240.244
R10013 gnd.n3304 gnd.n2394 240.244
R10014 gnd.n3300 gnd.n2394 240.244
R10015 gnd.n3300 gnd.n2396 240.244
R10016 gnd.n3296 gnd.n2396 240.244
R10017 gnd.n3296 gnd.n2402 240.244
R10018 gnd.n3292 gnd.n2402 240.244
R10019 gnd.n3292 gnd.n2404 240.244
R10020 gnd.n3288 gnd.n2404 240.244
R10021 gnd.n3288 gnd.n2410 240.244
R10022 gnd.n3284 gnd.n2410 240.244
R10023 gnd.n3284 gnd.n2412 240.244
R10024 gnd.n3280 gnd.n2412 240.244
R10025 gnd.n3280 gnd.n2418 240.244
R10026 gnd.n3276 gnd.n2418 240.244
R10027 gnd.n3276 gnd.n2420 240.244
R10028 gnd.n3272 gnd.n2420 240.244
R10029 gnd.n3272 gnd.n2426 240.244
R10030 gnd.n3268 gnd.n2426 240.244
R10031 gnd.n3268 gnd.n2428 240.244
R10032 gnd.n3264 gnd.n2428 240.244
R10033 gnd.n3264 gnd.n2434 240.244
R10034 gnd.n3260 gnd.n2434 240.244
R10035 gnd.n3260 gnd.n2436 240.244
R10036 gnd.n3256 gnd.n2436 240.244
R10037 gnd.n3256 gnd.n2442 240.244
R10038 gnd.n3252 gnd.n2442 240.244
R10039 gnd.n3252 gnd.n2444 240.244
R10040 gnd.n3248 gnd.n2444 240.244
R10041 gnd.n3248 gnd.n2450 240.244
R10042 gnd.n3244 gnd.n2450 240.244
R10043 gnd.n3244 gnd.n2452 240.244
R10044 gnd.n3240 gnd.n2452 240.244
R10045 gnd.n3240 gnd.n2458 240.244
R10046 gnd.n3236 gnd.n2458 240.244
R10047 gnd.n3236 gnd.n2460 240.244
R10048 gnd.n3232 gnd.n2460 240.244
R10049 gnd.n3232 gnd.n2466 240.244
R10050 gnd.n3228 gnd.n2466 240.244
R10051 gnd.n3228 gnd.n2468 240.244
R10052 gnd.n3224 gnd.n2468 240.244
R10053 gnd.n3224 gnd.n2474 240.244
R10054 gnd.n3220 gnd.n2474 240.244
R10055 gnd.n3220 gnd.n2476 240.244
R10056 gnd.n3216 gnd.n2476 240.244
R10057 gnd.n3216 gnd.n2482 240.244
R10058 gnd.n3212 gnd.n2482 240.244
R10059 gnd.n3212 gnd.n2484 240.244
R10060 gnd.n3208 gnd.n2484 240.244
R10061 gnd.n3208 gnd.n2490 240.244
R10062 gnd.n3204 gnd.n2490 240.244
R10063 gnd.n3204 gnd.n2492 240.244
R10064 gnd.n3200 gnd.n2492 240.244
R10065 gnd.n3200 gnd.n2498 240.244
R10066 gnd.n3196 gnd.n2498 240.244
R10067 gnd.n3196 gnd.n2500 240.244
R10068 gnd.n3192 gnd.n2500 240.244
R10069 gnd.n3192 gnd.n2506 240.244
R10070 gnd.n3188 gnd.n2506 240.244
R10071 gnd.n3188 gnd.n2508 240.244
R10072 gnd.n3184 gnd.n2508 240.244
R10073 gnd.n3184 gnd.n2514 240.244
R10074 gnd.n3180 gnd.n2514 240.244
R10075 gnd.n3180 gnd.n2516 240.244
R10076 gnd.n3176 gnd.n2516 240.244
R10077 gnd.n3176 gnd.n2522 240.244
R10078 gnd.n3172 gnd.n2522 240.244
R10079 gnd.n3172 gnd.n2524 240.244
R10080 gnd.n3168 gnd.n2524 240.244
R10081 gnd.n3168 gnd.n2530 240.244
R10082 gnd.n3164 gnd.n2530 240.244
R10083 gnd.n3164 gnd.n2532 240.244
R10084 gnd.n3160 gnd.n2532 240.244
R10085 gnd.n3160 gnd.n2538 240.244
R10086 gnd.n3156 gnd.n2538 240.244
R10087 gnd.n3156 gnd.n2540 240.244
R10088 gnd.n3152 gnd.n2540 240.244
R10089 gnd.n3152 gnd.n2546 240.244
R10090 gnd.n3148 gnd.n2546 240.244
R10091 gnd.n3148 gnd.n2548 240.244
R10092 gnd.n3144 gnd.n2548 240.244
R10093 gnd.n3144 gnd.n2554 240.244
R10094 gnd.n3140 gnd.n2554 240.244
R10095 gnd.n3140 gnd.n2556 240.244
R10096 gnd.n3136 gnd.n2556 240.244
R10097 gnd.n3136 gnd.n2562 240.244
R10098 gnd.n3132 gnd.n2562 240.244
R10099 gnd.n3132 gnd.n2564 240.244
R10100 gnd.n3128 gnd.n2564 240.244
R10101 gnd.n3128 gnd.n2570 240.244
R10102 gnd.n3124 gnd.n2570 240.244
R10103 gnd.n3124 gnd.n2572 240.244
R10104 gnd.n3120 gnd.n2572 240.244
R10105 gnd.n3120 gnd.n2578 240.244
R10106 gnd.n3116 gnd.n2578 240.244
R10107 gnd.n3116 gnd.n2580 240.244
R10108 gnd.n3112 gnd.n2580 240.244
R10109 gnd.n3112 gnd.n2586 240.244
R10110 gnd.n3108 gnd.n2586 240.244
R10111 gnd.n3108 gnd.n2588 240.244
R10112 gnd.n3104 gnd.n2588 240.244
R10113 gnd.n3104 gnd.n2594 240.244
R10114 gnd.n3100 gnd.n2594 240.244
R10115 gnd.n3100 gnd.n2596 240.244
R10116 gnd.n3096 gnd.n2596 240.244
R10117 gnd.n3096 gnd.n2602 240.244
R10118 gnd.n3092 gnd.n2602 240.244
R10119 gnd.n3092 gnd.n2604 240.244
R10120 gnd.n3088 gnd.n2604 240.244
R10121 gnd.n3088 gnd.n2610 240.244
R10122 gnd.n3084 gnd.n2610 240.244
R10123 gnd.n3084 gnd.n2612 240.244
R10124 gnd.n3080 gnd.n2612 240.244
R10125 gnd.n3080 gnd.n2618 240.244
R10126 gnd.n3076 gnd.n2618 240.244
R10127 gnd.n3076 gnd.n2620 240.244
R10128 gnd.n3072 gnd.n2620 240.244
R10129 gnd.n3072 gnd.n2626 240.244
R10130 gnd.n3068 gnd.n2626 240.244
R10131 gnd.n3068 gnd.n2628 240.244
R10132 gnd.n3064 gnd.n2628 240.244
R10133 gnd.n3064 gnd.n2634 240.244
R10134 gnd.n3060 gnd.n2634 240.244
R10135 gnd.n3060 gnd.n2636 240.244
R10136 gnd.n3056 gnd.n2636 240.244
R10137 gnd.n3056 gnd.n2642 240.244
R10138 gnd.n3052 gnd.n2642 240.244
R10139 gnd.n3052 gnd.n2644 240.244
R10140 gnd.n3048 gnd.n2644 240.244
R10141 gnd.n3048 gnd.n2650 240.244
R10142 gnd.n3044 gnd.n2650 240.244
R10143 gnd.n3044 gnd.n2652 240.244
R10144 gnd.n3040 gnd.n2652 240.244
R10145 gnd.n3040 gnd.n2658 240.244
R10146 gnd.n3036 gnd.n2658 240.244
R10147 gnd.n3036 gnd.n2660 240.244
R10148 gnd.n3030 gnd.n2665 240.244
R10149 gnd.n3026 gnd.n2665 240.244
R10150 gnd.n3026 gnd.n2667 240.244
R10151 gnd.n3022 gnd.n2667 240.244
R10152 gnd.n3022 gnd.n2672 240.244
R10153 gnd.n3018 gnd.n2672 240.244
R10154 gnd.n3018 gnd.n2674 240.244
R10155 gnd.n3014 gnd.n2674 240.244
R10156 gnd.n3014 gnd.n2680 240.244
R10157 gnd.n3010 gnd.n2680 240.244
R10158 gnd.n3010 gnd.n2682 240.244
R10159 gnd.n3006 gnd.n2682 240.244
R10160 gnd.n3006 gnd.n2688 240.244
R10161 gnd.n3002 gnd.n2688 240.244
R10162 gnd.n3002 gnd.n2690 240.244
R10163 gnd.n2998 gnd.n2690 240.244
R10164 gnd.n2998 gnd.n2696 240.244
R10165 gnd.n2994 gnd.n2696 240.244
R10166 gnd.n2994 gnd.n2698 240.244
R10167 gnd.n2990 gnd.n2698 240.244
R10168 gnd.n2990 gnd.n2704 240.244
R10169 gnd.n2986 gnd.n2704 240.244
R10170 gnd.n2986 gnd.n2706 240.244
R10171 gnd.n2982 gnd.n2706 240.244
R10172 gnd.n2982 gnd.n2712 240.244
R10173 gnd.n2978 gnd.n2712 240.244
R10174 gnd.n2978 gnd.n2714 240.244
R10175 gnd.n2974 gnd.n2714 240.244
R10176 gnd.n2974 gnd.n2720 240.244
R10177 gnd.n2970 gnd.n2720 240.244
R10178 gnd.n2970 gnd.n2722 240.244
R10179 gnd.n2966 gnd.n2722 240.244
R10180 gnd.n2966 gnd.n2728 240.244
R10181 gnd.n2962 gnd.n2728 240.244
R10182 gnd.n2962 gnd.n2730 240.244
R10183 gnd.n2958 gnd.n2730 240.244
R10184 gnd.n2958 gnd.n2736 240.244
R10185 gnd.n2954 gnd.n2736 240.244
R10186 gnd.n2954 gnd.n2738 240.244
R10187 gnd.n2950 gnd.n2738 240.244
R10188 gnd.n2950 gnd.n2744 240.244
R10189 gnd.n2946 gnd.n2744 240.244
R10190 gnd.n2946 gnd.n2746 240.244
R10191 gnd.n2942 gnd.n2746 240.244
R10192 gnd.n2942 gnd.n2752 240.244
R10193 gnd.n2938 gnd.n2752 240.244
R10194 gnd.n2938 gnd.n2754 240.244
R10195 gnd.n2934 gnd.n2754 240.244
R10196 gnd.n2934 gnd.n2760 240.244
R10197 gnd.n2930 gnd.n2760 240.244
R10198 gnd.n2930 gnd.n2762 240.244
R10199 gnd.n2926 gnd.n2762 240.244
R10200 gnd.n2926 gnd.n2768 240.244
R10201 gnd.n2922 gnd.n2768 240.244
R10202 gnd.n2922 gnd.n2770 240.244
R10203 gnd.n2918 gnd.n2770 240.244
R10204 gnd.n2918 gnd.n2776 240.244
R10205 gnd.n2914 gnd.n2776 240.244
R10206 gnd.n2914 gnd.n2778 240.244
R10207 gnd.n2910 gnd.n2778 240.244
R10208 gnd.n2910 gnd.n2784 240.244
R10209 gnd.n2906 gnd.n2784 240.244
R10210 gnd.n2906 gnd.n2786 240.244
R10211 gnd.n2902 gnd.n2786 240.244
R10212 gnd.n2902 gnd.n2899 240.244
R10213 gnd.n2899 gnd.n2898 240.244
R10214 gnd.n5170 gnd.n5169 240.244
R10215 gnd.n5170 gnd.n2218 240.244
R10216 gnd.n5219 gnd.n2218 240.244
R10217 gnd.n5219 gnd.n2219 240.244
R10218 gnd.n5215 gnd.n2219 240.244
R10219 gnd.n5215 gnd.n5214 240.244
R10220 gnd.n5214 gnd.n5213 240.244
R10221 gnd.n5213 gnd.n5178 240.244
R10222 gnd.n5209 gnd.n5178 240.244
R10223 gnd.n5209 gnd.n5208 240.244
R10224 gnd.n5208 gnd.n5207 240.244
R10225 gnd.n5207 gnd.n5184 240.244
R10226 gnd.n5203 gnd.n5184 240.244
R10227 gnd.n5203 gnd.n5202 240.244
R10228 gnd.n5202 gnd.n5201 240.244
R10229 gnd.n5201 gnd.n5191 240.244
R10230 gnd.n5196 gnd.n5191 240.244
R10231 gnd.n5196 gnd.n5195 240.244
R10232 gnd.n5195 gnd.n1869 240.244
R10233 gnd.n5630 gnd.n1869 240.244
R10234 gnd.n5630 gnd.n1870 240.244
R10235 gnd.n5625 gnd.n1870 240.244
R10236 gnd.n5625 gnd.n1873 240.244
R10237 gnd.n5461 gnd.n1873 240.244
R10238 gnd.n5462 gnd.n5461 240.244
R10239 gnd.n5462 gnd.n5457 240.244
R10240 gnd.n5468 gnd.n5457 240.244
R10241 gnd.n5469 gnd.n5468 240.244
R10242 gnd.n5470 gnd.n5469 240.244
R10243 gnd.n5470 gnd.n5453 240.244
R10244 gnd.n5513 gnd.n5453 240.244
R10245 gnd.n5514 gnd.n5513 240.244
R10246 gnd.n5515 gnd.n5514 240.244
R10247 gnd.n5515 gnd.n5449 240.244
R10248 gnd.n5521 gnd.n5449 240.244
R10249 gnd.n5522 gnd.n5521 240.244
R10250 gnd.n5523 gnd.n5522 240.244
R10251 gnd.n5523 gnd.n5445 240.244
R10252 gnd.n5529 gnd.n5445 240.244
R10253 gnd.n5530 gnd.n5529 240.244
R10254 gnd.n5531 gnd.n5530 240.244
R10255 gnd.n5531 gnd.n5440 240.244
R10256 gnd.n5557 gnd.n5440 240.244
R10257 gnd.n5557 gnd.n5441 240.244
R10258 gnd.n5553 gnd.n5441 240.244
R10259 gnd.n5553 gnd.n5552 240.244
R10260 gnd.n5552 gnd.n5551 240.244
R10261 gnd.n5551 gnd.n5539 240.244
R10262 gnd.n5546 gnd.n5539 240.244
R10263 gnd.n5546 gnd.n1674 240.244
R10264 gnd.n5811 gnd.n1674 240.244
R10265 gnd.n5811 gnd.n1670 240.244
R10266 gnd.n5817 gnd.n1670 240.244
R10267 gnd.n5817 gnd.n1662 240.244
R10268 gnd.n5831 gnd.n1662 240.244
R10269 gnd.n5831 gnd.n1658 240.244
R10270 gnd.n5837 gnd.n1658 240.244
R10271 gnd.n5837 gnd.n1649 240.244
R10272 gnd.n5851 gnd.n1649 240.244
R10273 gnd.n5851 gnd.n1644 240.244
R10274 gnd.n5859 gnd.n1644 240.244
R10275 gnd.n5859 gnd.n1645 240.244
R10276 gnd.n1645 gnd.n1431 240.244
R10277 gnd.n6062 gnd.n1431 240.244
R10278 gnd.n6062 gnd.n1426 240.244
R10279 gnd.n6070 gnd.n1426 240.244
R10280 gnd.n6070 gnd.n1427 240.244
R10281 gnd.n1427 gnd.n1398 240.244
R10282 gnd.n6144 gnd.n1398 240.244
R10283 gnd.n6144 gnd.n1394 240.244
R10284 gnd.n6150 gnd.n1394 240.244
R10285 gnd.n6150 gnd.n1374 240.244
R10286 gnd.n6172 gnd.n1374 240.244
R10287 gnd.n6172 gnd.n1369 240.244
R10288 gnd.n6193 gnd.n1369 240.244
R10289 gnd.n6193 gnd.n1370 240.244
R10290 gnd.n6189 gnd.n1370 240.244
R10291 gnd.n6189 gnd.n6188 240.244
R10292 gnd.n6188 gnd.n6186 240.244
R10293 gnd.n6186 gnd.n6180 240.244
R10294 gnd.n6180 gnd.n1313 240.244
R10295 gnd.n6283 gnd.n1313 240.244
R10296 gnd.n6283 gnd.n1308 240.244
R10297 gnd.n6302 gnd.n1308 240.244
R10298 gnd.n6302 gnd.n1309 240.244
R10299 gnd.n6298 gnd.n1309 240.244
R10300 gnd.n6298 gnd.n6296 240.244
R10301 gnd.n6296 gnd.n6295 240.244
R10302 gnd.n6295 gnd.n1266 240.244
R10303 gnd.n6388 gnd.n1266 240.244
R10304 gnd.n6388 gnd.n1267 240.244
R10305 gnd.n6384 gnd.n1267 240.244
R10306 gnd.n6384 gnd.n1237 240.244
R10307 gnd.n6425 gnd.n1237 240.244
R10308 gnd.n6425 gnd.n1238 240.244
R10309 gnd.n6421 gnd.n1238 240.244
R10310 gnd.n6421 gnd.n1208 240.244
R10311 gnd.n6465 gnd.n1208 240.244
R10312 gnd.n6465 gnd.n1209 240.244
R10313 gnd.n6461 gnd.n1209 240.244
R10314 gnd.n6461 gnd.n1216 240.244
R10315 gnd.n1216 gnd.n1108 240.244
R10316 gnd.n6612 gnd.n1108 240.244
R10317 gnd.n6612 gnd.n1103 240.244
R10318 gnd.n6620 gnd.n1103 240.244
R10319 gnd.n6620 gnd.n1104 240.244
R10320 gnd.n1104 gnd.n1082 240.244
R10321 gnd.n6642 gnd.n1082 240.244
R10322 gnd.n6642 gnd.n1077 240.244
R10323 gnd.n6650 gnd.n1077 240.244
R10324 gnd.n6650 gnd.n1078 240.244
R10325 gnd.n1078 gnd.n1057 240.244
R10326 gnd.n6673 gnd.n1057 240.244
R10327 gnd.n6673 gnd.n1052 240.244
R10328 gnd.n6692 gnd.n1052 240.244
R10329 gnd.n6692 gnd.n1053 240.244
R10330 gnd.n6688 gnd.n1053 240.244
R10331 gnd.n6688 gnd.n6687 240.244
R10332 gnd.n6687 gnd.n6684 240.244
R10333 gnd.n6684 gnd.n972 240.244
R10334 gnd.n6714 gnd.n972 240.244
R10335 gnd.n6714 gnd.n968 240.244
R10336 gnd.n6720 gnd.n968 240.244
R10337 gnd.n6721 gnd.n6720 240.244
R10338 gnd.n6722 gnd.n6721 240.244
R10339 gnd.n6722 gnd.n964 240.244
R10340 gnd.n6728 gnd.n964 240.244
R10341 gnd.n6729 gnd.n6728 240.244
R10342 gnd.n6730 gnd.n6729 240.244
R10343 gnd.n6730 gnd.n960 240.244
R10344 gnd.n6736 gnd.n960 240.244
R10345 gnd.n6737 gnd.n6736 240.244
R10346 gnd.n6738 gnd.n6737 240.244
R10347 gnd.n6738 gnd.n956 240.244
R10348 gnd.n6744 gnd.n956 240.244
R10349 gnd.n6745 gnd.n6744 240.244
R10350 gnd.n6746 gnd.n6745 240.244
R10351 gnd.n6746 gnd.n952 240.244
R10352 gnd.n6813 gnd.n952 240.244
R10353 gnd.n6814 gnd.n6813 240.244
R10354 gnd.n6815 gnd.n6814 240.244
R10355 gnd.n6815 gnd.n948 240.244
R10356 gnd.n6821 gnd.n948 240.244
R10357 gnd.n6822 gnd.n6821 240.244
R10358 gnd.n6835 gnd.n6822 240.244
R10359 gnd.n6835 gnd.n6834 240.244
R10360 gnd.n6834 gnd.n6833 240.244
R10361 gnd.n6833 gnd.n6830 240.244
R10362 gnd.n6830 gnd.n6829 240.244
R10363 gnd.n6829 gnd.n6826 240.244
R10364 gnd.n6826 gnd.n6825 240.244
R10365 gnd.n6825 gnd.n937 240.244
R10366 gnd.n6842 gnd.n937 240.244
R10367 gnd.n6842 gnd.n938 240.244
R10368 gnd.n2807 gnd.n938 240.244
R10369 gnd.n2808 gnd.n2807 240.244
R10370 gnd.n2809 gnd.n2808 240.244
R10371 gnd.n2809 gnd.n2804 240.244
R10372 gnd.n2815 gnd.n2804 240.244
R10373 gnd.n2816 gnd.n2815 240.244
R10374 gnd.n2817 gnd.n2816 240.244
R10375 gnd.n2817 gnd.n2800 240.244
R10376 gnd.n2823 gnd.n2800 240.244
R10377 gnd.n2824 gnd.n2823 240.244
R10378 gnd.n2825 gnd.n2824 240.244
R10379 gnd.n2825 gnd.n2796 240.244
R10380 gnd.n2890 gnd.n2796 240.244
R10381 gnd.n2891 gnd.n2890 240.244
R10382 gnd.n2892 gnd.n2891 240.244
R10383 gnd.n2892 gnd.n2792 240.244
R10384 gnd.n3376 gnd.n2319 240.244
R10385 gnd.n3382 gnd.n2319 240.244
R10386 gnd.n3382 gnd.n2317 240.244
R10387 gnd.n3386 gnd.n2317 240.244
R10388 gnd.n3386 gnd.n2313 240.244
R10389 gnd.n3392 gnd.n2313 240.244
R10390 gnd.n3392 gnd.n2311 240.244
R10391 gnd.n3396 gnd.n2311 240.244
R10392 gnd.n3396 gnd.n2307 240.244
R10393 gnd.n3402 gnd.n2307 240.244
R10394 gnd.n3402 gnd.n2305 240.244
R10395 gnd.n3406 gnd.n2305 240.244
R10396 gnd.n3406 gnd.n2301 240.244
R10397 gnd.n3412 gnd.n2301 240.244
R10398 gnd.n3412 gnd.n2299 240.244
R10399 gnd.n3416 gnd.n2299 240.244
R10400 gnd.n3416 gnd.n2295 240.244
R10401 gnd.n3422 gnd.n2295 240.244
R10402 gnd.n3422 gnd.n2293 240.244
R10403 gnd.n3426 gnd.n2293 240.244
R10404 gnd.n3426 gnd.n2289 240.244
R10405 gnd.n3432 gnd.n2289 240.244
R10406 gnd.n3432 gnd.n2287 240.244
R10407 gnd.n3436 gnd.n2287 240.244
R10408 gnd.n3436 gnd.n2283 240.244
R10409 gnd.n3442 gnd.n2283 240.244
R10410 gnd.n3442 gnd.n2281 240.244
R10411 gnd.n3446 gnd.n2281 240.244
R10412 gnd.n3446 gnd.n2277 240.244
R10413 gnd.n3452 gnd.n2277 240.244
R10414 gnd.n3452 gnd.n2275 240.244
R10415 gnd.n3456 gnd.n2275 240.244
R10416 gnd.n3456 gnd.n2271 240.244
R10417 gnd.n3462 gnd.n2271 240.244
R10418 gnd.n3462 gnd.n2269 240.244
R10419 gnd.n3466 gnd.n2269 240.244
R10420 gnd.n3466 gnd.n2265 240.244
R10421 gnd.n3472 gnd.n2265 240.244
R10422 gnd.n3472 gnd.n2263 240.244
R10423 gnd.n3476 gnd.n2263 240.244
R10424 gnd.n3476 gnd.n2259 240.244
R10425 gnd.n3482 gnd.n2259 240.244
R10426 gnd.n3482 gnd.n2257 240.244
R10427 gnd.n3486 gnd.n2257 240.244
R10428 gnd.n3486 gnd.n2253 240.244
R10429 gnd.n3492 gnd.n2253 240.244
R10430 gnd.n3492 gnd.n2251 240.244
R10431 gnd.n3496 gnd.n2251 240.244
R10432 gnd.n3496 gnd.n2247 240.244
R10433 gnd.n3502 gnd.n2247 240.244
R10434 gnd.n3502 gnd.n2245 240.244
R10435 gnd.n3506 gnd.n2245 240.244
R10436 gnd.n3506 gnd.n2241 240.244
R10437 gnd.n3512 gnd.n2241 240.244
R10438 gnd.n3512 gnd.n2239 240.244
R10439 gnd.n3516 gnd.n2239 240.244
R10440 gnd.n3516 gnd.n2235 240.244
R10441 gnd.n3522 gnd.n2235 240.244
R10442 gnd.n3522 gnd.n2233 240.244
R10443 gnd.n3526 gnd.n2233 240.244
R10444 gnd.n3526 gnd.n2229 240.244
R10445 gnd.n3532 gnd.n2229 240.244
R10446 gnd.n3532 gnd.n2227 240.244
R10447 gnd.n5162 gnd.n2227 240.244
R10448 gnd.n5162 gnd.n2223 240.244
R10449 gnd.n5168 gnd.n2223 240.244
R10450 gnd.n1623 gnd.n1622 240.244
R10451 gnd.n1624 gnd.n1623 240.244
R10452 gnd.n5828 gnd.n1624 240.244
R10453 gnd.n5828 gnd.n1627 240.244
R10454 gnd.n1628 gnd.n1627 240.244
R10455 gnd.n1629 gnd.n1628 240.244
R10456 gnd.n5848 gnd.n1629 240.244
R10457 gnd.n5848 gnd.n1632 240.244
R10458 gnd.n1633 gnd.n1632 240.244
R10459 gnd.n5876 gnd.n1633 240.244
R10460 gnd.n5877 gnd.n5876 240.244
R10461 gnd.n5877 gnd.n1422 240.244
R10462 gnd.n6073 gnd.n1422 240.244
R10463 gnd.n6073 gnd.n1416 240.244
R10464 gnd.n6080 gnd.n1416 240.244
R10465 gnd.n6080 gnd.n1417 240.244
R10466 gnd.n1417 gnd.n1390 240.244
R10467 gnd.n6153 gnd.n1390 240.244
R10468 gnd.n6153 gnd.n1384 240.244
R10469 gnd.n6160 gnd.n1384 240.244
R10470 gnd.n6160 gnd.n1385 240.244
R10471 gnd.n1385 gnd.n1358 240.244
R10472 gnd.n6204 gnd.n1358 240.244
R10473 gnd.n6204 gnd.n1352 240.244
R10474 gnd.n6211 gnd.n1352 240.244
R10475 gnd.n6211 gnd.n1353 240.244
R10476 gnd.n1353 gnd.n1322 240.244
R10477 gnd.n6270 gnd.n1322 240.244
R10478 gnd.n6270 gnd.n1316 240.244
R10479 gnd.n6280 gnd.n1316 240.244
R10480 gnd.n6280 gnd.n1317 240.244
R10481 gnd.n6274 gnd.n1317 240.244
R10482 gnd.n6274 gnd.n1284 240.244
R10483 gnd.n6333 gnd.n1284 240.244
R10484 gnd.n6333 gnd.n1280 240.244
R10485 gnd.n6339 gnd.n1280 240.244
R10486 gnd.n6339 gnd.n1254 240.244
R10487 gnd.n6402 gnd.n1254 240.244
R10488 gnd.n6402 gnd.n1250 240.244
R10489 gnd.n6408 gnd.n1250 240.244
R10490 gnd.n6408 gnd.n1226 240.244
R10491 gnd.n6438 gnd.n1226 240.244
R10492 gnd.n6438 gnd.n1222 240.244
R10493 gnd.n6444 gnd.n1222 240.244
R10494 gnd.n6444 gnd.n1198 240.244
R10495 gnd.n6475 gnd.n1198 240.244
R10496 gnd.n6475 gnd.n1192 240.244
R10497 gnd.n6485 gnd.n1192 240.244
R10498 gnd.n6485 gnd.n1193 240.244
R10499 gnd.n6479 gnd.n1193 240.244
R10500 gnd.n6479 gnd.n1098 240.244
R10501 gnd.n6623 gnd.n1098 240.244
R10502 gnd.n6623 gnd.n1092 240.244
R10503 gnd.n6630 gnd.n1092 240.244
R10504 gnd.n6630 gnd.n1093 240.244
R10505 gnd.n1093 gnd.n1073 240.244
R10506 gnd.n6653 gnd.n1073 240.244
R10507 gnd.n6653 gnd.n1067 240.244
R10508 gnd.n6660 gnd.n1067 240.244
R10509 gnd.n6660 gnd.n1068 240.244
R10510 gnd.n1068 gnd.n1048 240.244
R10511 gnd.n6695 gnd.n1048 240.244
R10512 gnd.n6695 gnd.n1042 240.244
R10513 gnd.n6702 gnd.n1042 240.244
R10514 gnd.n6702 gnd.n1043 240.244
R10515 gnd.n1689 gnd.n1688 240.244
R10516 gnd.n1705 gnd.n1688 240.244
R10517 gnd.n1707 gnd.n1706 240.244
R10518 gnd.n1717 gnd.n1716 240.244
R10519 gnd.n1728 gnd.n1727 240.244
R10520 gnd.n1730 gnd.n1729 240.244
R10521 gnd.n1740 gnd.n1739 240.244
R10522 gnd.n1750 gnd.n1749 240.244
R10523 gnd.n1752 gnd.n1751 240.244
R10524 gnd.n5736 gnd.n5735 240.244
R10525 gnd.n5738 gnd.n5737 240.244
R10526 gnd.n5745 gnd.n5744 240.244
R10527 gnd.n5747 gnd.n5746 240.244
R10528 gnd.n5820 gnd.n1664 240.244
R10529 gnd.n5826 gnd.n1664 240.244
R10530 gnd.n5826 gnd.n1655 240.244
R10531 gnd.n5840 gnd.n1655 240.244
R10532 gnd.n5840 gnd.n1651 240.244
R10533 gnd.n5846 gnd.n1651 240.244
R10534 gnd.n5846 gnd.n1641 240.244
R10535 gnd.n5862 gnd.n1641 240.244
R10536 gnd.n5862 gnd.n1635 240.244
R10537 gnd.n5873 gnd.n1635 240.244
R10538 gnd.n5873 gnd.n1636 240.244
R10539 gnd.n1636 gnd.n1433 240.244
R10540 gnd.n1433 gnd.n1424 240.244
R10541 gnd.n1424 gnd.n1414 240.244
R10542 gnd.n6082 gnd.n1414 240.244
R10543 gnd.n6082 gnd.n1409 240.244
R10544 gnd.n6122 gnd.n1409 240.244
R10545 gnd.n6122 gnd.n1392 240.244
R10546 gnd.n6087 gnd.n1392 240.244
R10547 gnd.n6087 gnd.n1383 240.244
R10548 gnd.n6088 gnd.n1383 240.244
R10549 gnd.n6088 gnd.n1368 240.244
R10550 gnd.n1368 gnd.n1360 240.244
R10551 gnd.n6107 gnd.n1360 240.244
R10552 gnd.n6107 gnd.n1350 240.244
R10553 gnd.n1350 gnd.n1337 240.244
R10554 gnd.n6229 gnd.n1337 240.244
R10555 gnd.n6229 gnd.n1324 240.244
R10556 gnd.n6248 gnd.n1324 240.244
R10557 gnd.n6248 gnd.n1315 240.244
R10558 gnd.n6234 gnd.n1315 240.244
R10559 gnd.n6235 gnd.n6234 240.244
R10560 gnd.n6236 gnd.n6235 240.244
R10561 gnd.n6236 gnd.n1286 240.244
R10562 gnd.n1286 gnd.n1278 240.244
R10563 gnd.n6341 gnd.n1278 240.244
R10564 gnd.n6341 gnd.n1265 240.244
R10565 gnd.n1265 gnd.n1256 240.244
R10566 gnd.n6381 gnd.n1256 240.244
R10567 gnd.n6381 gnd.n1249 240.244
R10568 gnd.n1249 gnd.n1236 240.244
R10569 gnd.n1236 gnd.n1228 240.244
R10570 gnd.n6347 gnd.n1228 240.244
R10571 gnd.n6347 gnd.n1221 240.244
R10572 gnd.n6350 gnd.n1221 240.244
R10573 gnd.n6350 gnd.n1200 240.244
R10574 gnd.n6351 gnd.n1200 240.244
R10575 gnd.n6351 gnd.n1190 240.244
R10576 gnd.n6356 gnd.n1190 240.244
R10577 gnd.n6357 gnd.n6356 240.244
R10578 gnd.n6358 gnd.n6357 240.244
R10579 gnd.n6358 gnd.n1100 240.244
R10580 gnd.n1100 gnd.n1089 240.244
R10581 gnd.n6632 gnd.n1089 240.244
R10582 gnd.n6632 gnd.n1084 240.244
R10583 gnd.n6639 gnd.n1084 240.244
R10584 gnd.n6639 gnd.n1075 240.244
R10585 gnd.n1075 gnd.n1064 240.244
R10586 gnd.n6662 gnd.n1064 240.244
R10587 gnd.n6662 gnd.n1059 240.244
R10588 gnd.n6670 gnd.n1059 240.244
R10589 gnd.n6670 gnd.n1050 240.244
R10590 gnd.n1050 gnd.n1039 240.244
R10591 gnd.n6704 gnd.n1039 240.244
R10592 gnd.n6704 gnd.n993 240.244
R10593 gnd.n975 gnd.n796 240.244
R10594 gnd.n804 gnd.n803 240.244
R10595 gnd.n977 gnd.n811 240.244
R10596 gnd.n980 gnd.n812 240.244
R10597 gnd.n820 gnd.n819 240.244
R10598 gnd.n982 gnd.n827 240.244
R10599 gnd.n985 gnd.n828 240.244
R10600 gnd.n1009 gnd.n1008 240.244
R10601 gnd.n1004 gnd.n1003 240.244
R10602 gnd.n1024 gnd.n1023 240.244
R10603 gnd.n1000 gnd.n999 240.244
R10604 gnd.n1033 gnd.n1032 240.244
R10605 gnd.n6710 gnd.n992 240.244
R10606 gnd.n1472 gnd.n1471 240.132
R10607 gnd.n1126 gnd.n1125 240.132
R10608 gnd.n2900 gnd.n502 227.53
R10609 gnd.n3374 gnd.n3373 225.874
R10610 gnd.n3373 gnd.n2323 225.874
R10611 gnd.n3367 gnd.n2323 225.874
R10612 gnd.n3367 gnd.n3366 225.874
R10613 gnd.n3366 gnd.n3365 225.874
R10614 gnd.n3365 gnd.n2331 225.874
R10615 gnd.n3359 gnd.n2331 225.874
R10616 gnd.n3359 gnd.n3358 225.874
R10617 gnd.n3358 gnd.n3357 225.874
R10618 gnd.n3357 gnd.n2339 225.874
R10619 gnd.n3351 gnd.n2339 225.874
R10620 gnd.n3351 gnd.n3350 225.874
R10621 gnd.n3350 gnd.n3349 225.874
R10622 gnd.n3349 gnd.n2347 225.874
R10623 gnd.n3343 gnd.n2347 225.874
R10624 gnd.n3343 gnd.n3342 225.874
R10625 gnd.n3342 gnd.n3341 225.874
R10626 gnd.n3341 gnd.n2355 225.874
R10627 gnd.n3335 gnd.n2355 225.874
R10628 gnd.n3335 gnd.n3334 225.874
R10629 gnd.n3334 gnd.n3333 225.874
R10630 gnd.n3333 gnd.n2363 225.874
R10631 gnd.n3327 gnd.n2363 225.874
R10632 gnd.n3327 gnd.n3326 225.874
R10633 gnd.n3326 gnd.n3325 225.874
R10634 gnd.n3325 gnd.n2371 225.874
R10635 gnd.n3319 gnd.n2371 225.874
R10636 gnd.n3319 gnd.n3318 225.874
R10637 gnd.n3318 gnd.n3317 225.874
R10638 gnd.n3317 gnd.n2379 225.874
R10639 gnd.n3311 gnd.n2379 225.874
R10640 gnd.n3311 gnd.n3310 225.874
R10641 gnd.n3310 gnd.n3309 225.874
R10642 gnd.n3309 gnd.n2387 225.874
R10643 gnd.n3303 gnd.n2387 225.874
R10644 gnd.n3303 gnd.n3302 225.874
R10645 gnd.n3302 gnd.n3301 225.874
R10646 gnd.n3301 gnd.n2395 225.874
R10647 gnd.n3295 gnd.n2395 225.874
R10648 gnd.n3295 gnd.n3294 225.874
R10649 gnd.n3294 gnd.n3293 225.874
R10650 gnd.n3293 gnd.n2403 225.874
R10651 gnd.n3287 gnd.n2403 225.874
R10652 gnd.n3287 gnd.n3286 225.874
R10653 gnd.n3286 gnd.n3285 225.874
R10654 gnd.n3285 gnd.n2411 225.874
R10655 gnd.n3279 gnd.n2411 225.874
R10656 gnd.n3279 gnd.n3278 225.874
R10657 gnd.n3278 gnd.n3277 225.874
R10658 gnd.n3277 gnd.n2419 225.874
R10659 gnd.n3271 gnd.n2419 225.874
R10660 gnd.n3271 gnd.n3270 225.874
R10661 gnd.n3270 gnd.n3269 225.874
R10662 gnd.n3269 gnd.n2427 225.874
R10663 gnd.n3263 gnd.n2427 225.874
R10664 gnd.n3263 gnd.n3262 225.874
R10665 gnd.n3262 gnd.n3261 225.874
R10666 gnd.n3261 gnd.n2435 225.874
R10667 gnd.n3255 gnd.n2435 225.874
R10668 gnd.n3255 gnd.n3254 225.874
R10669 gnd.n3254 gnd.n3253 225.874
R10670 gnd.n3253 gnd.n2443 225.874
R10671 gnd.n3247 gnd.n2443 225.874
R10672 gnd.n3247 gnd.n3246 225.874
R10673 gnd.n3246 gnd.n3245 225.874
R10674 gnd.n3245 gnd.n2451 225.874
R10675 gnd.n3239 gnd.n2451 225.874
R10676 gnd.n3239 gnd.n3238 225.874
R10677 gnd.n3238 gnd.n3237 225.874
R10678 gnd.n3237 gnd.n2459 225.874
R10679 gnd.n3231 gnd.n2459 225.874
R10680 gnd.n3231 gnd.n3230 225.874
R10681 gnd.n3230 gnd.n3229 225.874
R10682 gnd.n3229 gnd.n2467 225.874
R10683 gnd.n3223 gnd.n2467 225.874
R10684 gnd.n3223 gnd.n3222 225.874
R10685 gnd.n3222 gnd.n3221 225.874
R10686 gnd.n3221 gnd.n2475 225.874
R10687 gnd.n3215 gnd.n2475 225.874
R10688 gnd.n3215 gnd.n3214 225.874
R10689 gnd.n3214 gnd.n3213 225.874
R10690 gnd.n3213 gnd.n2483 225.874
R10691 gnd.n3207 gnd.n2483 225.874
R10692 gnd.n3207 gnd.n3206 225.874
R10693 gnd.n3206 gnd.n3205 225.874
R10694 gnd.n3205 gnd.n2491 225.874
R10695 gnd.n3199 gnd.n2491 225.874
R10696 gnd.n3199 gnd.n3198 225.874
R10697 gnd.n3198 gnd.n3197 225.874
R10698 gnd.n3197 gnd.n2499 225.874
R10699 gnd.n3191 gnd.n2499 225.874
R10700 gnd.n3191 gnd.n3190 225.874
R10701 gnd.n3190 gnd.n3189 225.874
R10702 gnd.n3189 gnd.n2507 225.874
R10703 gnd.n3183 gnd.n2507 225.874
R10704 gnd.n3183 gnd.n3182 225.874
R10705 gnd.n3182 gnd.n3181 225.874
R10706 gnd.n3181 gnd.n2515 225.874
R10707 gnd.n3175 gnd.n2515 225.874
R10708 gnd.n3175 gnd.n3174 225.874
R10709 gnd.n3174 gnd.n3173 225.874
R10710 gnd.n3173 gnd.n2523 225.874
R10711 gnd.n3167 gnd.n2523 225.874
R10712 gnd.n3167 gnd.n3166 225.874
R10713 gnd.n3166 gnd.n3165 225.874
R10714 gnd.n3165 gnd.n2531 225.874
R10715 gnd.n3159 gnd.n2531 225.874
R10716 gnd.n3159 gnd.n3158 225.874
R10717 gnd.n3158 gnd.n3157 225.874
R10718 gnd.n3157 gnd.n2539 225.874
R10719 gnd.n3151 gnd.n2539 225.874
R10720 gnd.n3151 gnd.n3150 225.874
R10721 gnd.n3150 gnd.n3149 225.874
R10722 gnd.n3149 gnd.n2547 225.874
R10723 gnd.n3143 gnd.n2547 225.874
R10724 gnd.n3143 gnd.n3142 225.874
R10725 gnd.n3142 gnd.n3141 225.874
R10726 gnd.n3141 gnd.n2555 225.874
R10727 gnd.n3135 gnd.n2555 225.874
R10728 gnd.n3135 gnd.n3134 225.874
R10729 gnd.n3134 gnd.n3133 225.874
R10730 gnd.n3133 gnd.n2563 225.874
R10731 gnd.n3127 gnd.n2563 225.874
R10732 gnd.n3127 gnd.n3126 225.874
R10733 gnd.n3126 gnd.n3125 225.874
R10734 gnd.n3125 gnd.n2571 225.874
R10735 gnd.n3119 gnd.n2571 225.874
R10736 gnd.n3119 gnd.n3118 225.874
R10737 gnd.n3118 gnd.n3117 225.874
R10738 gnd.n3117 gnd.n2579 225.874
R10739 gnd.n3111 gnd.n2579 225.874
R10740 gnd.n3111 gnd.n3110 225.874
R10741 gnd.n3110 gnd.n3109 225.874
R10742 gnd.n3109 gnd.n2587 225.874
R10743 gnd.n3103 gnd.n2587 225.874
R10744 gnd.n3103 gnd.n3102 225.874
R10745 gnd.n3102 gnd.n3101 225.874
R10746 gnd.n3101 gnd.n2595 225.874
R10747 gnd.n3095 gnd.n2595 225.874
R10748 gnd.n3095 gnd.n3094 225.874
R10749 gnd.n3094 gnd.n3093 225.874
R10750 gnd.n3093 gnd.n2603 225.874
R10751 gnd.n3087 gnd.n2603 225.874
R10752 gnd.n3087 gnd.n3086 225.874
R10753 gnd.n3086 gnd.n3085 225.874
R10754 gnd.n3085 gnd.n2611 225.874
R10755 gnd.n3079 gnd.n2611 225.874
R10756 gnd.n3079 gnd.n3078 225.874
R10757 gnd.n3078 gnd.n3077 225.874
R10758 gnd.n3077 gnd.n2619 225.874
R10759 gnd.n3071 gnd.n2619 225.874
R10760 gnd.n3071 gnd.n3070 225.874
R10761 gnd.n3070 gnd.n3069 225.874
R10762 gnd.n3069 gnd.n2627 225.874
R10763 gnd.n3063 gnd.n2627 225.874
R10764 gnd.n3063 gnd.n3062 225.874
R10765 gnd.n3062 gnd.n3061 225.874
R10766 gnd.n3061 gnd.n2635 225.874
R10767 gnd.n3055 gnd.n2635 225.874
R10768 gnd.n3055 gnd.n3054 225.874
R10769 gnd.n3054 gnd.n3053 225.874
R10770 gnd.n3053 gnd.n2643 225.874
R10771 gnd.n3047 gnd.n2643 225.874
R10772 gnd.n3047 gnd.n3046 225.874
R10773 gnd.n3046 gnd.n3045 225.874
R10774 gnd.n3045 gnd.n2651 225.874
R10775 gnd.n3039 gnd.n2651 225.874
R10776 gnd.n3039 gnd.n3038 225.874
R10777 gnd.n3038 gnd.n3037 225.874
R10778 gnd.n3037 gnd.n2659 225.874
R10779 gnd.n5741 gnd.t206 224.174
R10780 gnd.n3971 gnd.t199 224.174
R10781 gnd.n3674 gnd.t129 224.174
R10782 gnd.n7235 gnd.t161 224.174
R10783 gnd.n6968 gnd.t137 224.174
R10784 gnd.n1743 gnd.t133 224.174
R10785 gnd.n880 gnd.t112 224.174
R10786 gnd.n900 gnd.t202 224.174
R10787 gnd.n571 gnd.t170 224.174
R10788 gnd.n535 gnd.t185 224.174
R10789 gnd.n2122 gnd.t151 224.174
R10790 gnd.n2051 gnd.t126 224.174
R10791 gnd.n5243 gnd.t154 224.174
R10792 gnd.n1594 gnd.t164 224.174
R10793 gnd.n1559 gnd.t182 224.174
R10794 gnd.n996 gnd.t212 224.174
R10795 gnd.n3029 gnd.n3028 209.825
R10796 gnd.n3028 gnd.n3027 209.825
R10797 gnd.n3027 gnd.n2666 209.825
R10798 gnd.n3021 gnd.n2666 209.825
R10799 gnd.n3021 gnd.n3020 209.825
R10800 gnd.n3020 gnd.n3019 209.825
R10801 gnd.n3019 gnd.n2673 209.825
R10802 gnd.n3013 gnd.n2673 209.825
R10803 gnd.n3013 gnd.n3012 209.825
R10804 gnd.n3012 gnd.n3011 209.825
R10805 gnd.n3011 gnd.n2681 209.825
R10806 gnd.n3005 gnd.n2681 209.825
R10807 gnd.n3005 gnd.n3004 209.825
R10808 gnd.n3004 gnd.n3003 209.825
R10809 gnd.n3003 gnd.n2689 209.825
R10810 gnd.n2997 gnd.n2689 209.825
R10811 gnd.n2997 gnd.n2996 209.825
R10812 gnd.n2996 gnd.n2995 209.825
R10813 gnd.n2995 gnd.n2697 209.825
R10814 gnd.n2989 gnd.n2697 209.825
R10815 gnd.n2989 gnd.n2988 209.825
R10816 gnd.n2988 gnd.n2987 209.825
R10817 gnd.n2987 gnd.n2705 209.825
R10818 gnd.n2981 gnd.n2705 209.825
R10819 gnd.n2981 gnd.n2980 209.825
R10820 gnd.n2980 gnd.n2979 209.825
R10821 gnd.n2979 gnd.n2713 209.825
R10822 gnd.n2973 gnd.n2713 209.825
R10823 gnd.n2973 gnd.n2972 209.825
R10824 gnd.n2972 gnd.n2971 209.825
R10825 gnd.n2971 gnd.n2721 209.825
R10826 gnd.n2965 gnd.n2721 209.825
R10827 gnd.n2965 gnd.n2964 209.825
R10828 gnd.n2964 gnd.n2963 209.825
R10829 gnd.n2963 gnd.n2729 209.825
R10830 gnd.n2957 gnd.n2729 209.825
R10831 gnd.n2957 gnd.n2956 209.825
R10832 gnd.n2956 gnd.n2955 209.825
R10833 gnd.n2955 gnd.n2737 209.825
R10834 gnd.n2949 gnd.n2737 209.825
R10835 gnd.n2949 gnd.n2948 209.825
R10836 gnd.n2948 gnd.n2947 209.825
R10837 gnd.n2947 gnd.n2745 209.825
R10838 gnd.n2941 gnd.n2745 209.825
R10839 gnd.n2941 gnd.n2940 209.825
R10840 gnd.n2940 gnd.n2939 209.825
R10841 gnd.n2939 gnd.n2753 209.825
R10842 gnd.n2933 gnd.n2753 209.825
R10843 gnd.n2933 gnd.n2932 209.825
R10844 gnd.n2932 gnd.n2931 209.825
R10845 gnd.n2931 gnd.n2761 209.825
R10846 gnd.n2925 gnd.n2761 209.825
R10847 gnd.n2925 gnd.n2924 209.825
R10848 gnd.n2924 gnd.n2923 209.825
R10849 gnd.n2923 gnd.n2769 209.825
R10850 gnd.n2917 gnd.n2769 209.825
R10851 gnd.n2917 gnd.n2916 209.825
R10852 gnd.n2916 gnd.n2915 209.825
R10853 gnd.n2915 gnd.n2777 209.825
R10854 gnd.n2909 gnd.n2777 209.825
R10855 gnd.n2909 gnd.n2908 209.825
R10856 gnd.n2908 gnd.n2907 209.825
R10857 gnd.n2907 gnd.n2785 209.825
R10858 gnd.n2901 gnd.n2785 209.825
R10859 gnd.n2901 gnd.n2900 209.825
R10860 gnd.n1490 gnd.t122 204.78
R10861 gnd.n1159 gnd.t157 204.78
R10862 gnd.n1488 gnd.t174 204.78
R10863 gnd.n1154 gnd.t188 204.78
R10864 gnd.n878 gnd.n839 199.319
R10865 gnd.n878 gnd.n840 199.319
R10866 gnd.n5927 gnd.n1561 199.319
R10867 gnd.n1566 gnd.n1561 199.319
R10868 gnd.n1473 gnd.n1470 186.49
R10869 gnd.n1127 gnd.n1124 186.49
R10870 gnd.n4293 gnd.n4292 185
R10871 gnd.n4291 gnd.n4290 185
R10872 gnd.n4270 gnd.n4269 185
R10873 gnd.n4285 gnd.n4284 185
R10874 gnd.n4283 gnd.n4282 185
R10875 gnd.n4274 gnd.n4273 185
R10876 gnd.n4277 gnd.n4276 185
R10877 gnd.n4330 gnd.n4329 185
R10878 gnd.n4328 gnd.n4327 185
R10879 gnd.n4307 gnd.n4306 185
R10880 gnd.n4322 gnd.n4321 185
R10881 gnd.n4320 gnd.n4319 185
R10882 gnd.n4311 gnd.n4310 185
R10883 gnd.n4314 gnd.n4313 185
R10884 gnd.n4154 gnd.n4153 185
R10885 gnd.n4152 gnd.n4151 185
R10886 gnd.n4131 gnd.n4130 185
R10887 gnd.n4146 gnd.n4145 185
R10888 gnd.n4144 gnd.n4143 185
R10889 gnd.n4135 gnd.n4134 185
R10890 gnd.n4138 gnd.n4137 185
R10891 gnd.n4191 gnd.n4190 185
R10892 gnd.n4189 gnd.n4188 185
R10893 gnd.n4168 gnd.n4167 185
R10894 gnd.n4183 gnd.n4182 185
R10895 gnd.n4181 gnd.n4180 185
R10896 gnd.n4172 gnd.n4171 185
R10897 gnd.n4175 gnd.n4174 185
R10898 gnd.n4223 gnd.n4222 185
R10899 gnd.n4221 gnd.n4220 185
R10900 gnd.n4200 gnd.n4199 185
R10901 gnd.n4215 gnd.n4214 185
R10902 gnd.n4213 gnd.n4212 185
R10903 gnd.n4204 gnd.n4203 185
R10904 gnd.n4207 gnd.n4206 185
R10905 gnd.n4260 gnd.n4259 185
R10906 gnd.n4258 gnd.n4257 185
R10907 gnd.n4237 gnd.n4236 185
R10908 gnd.n4252 gnd.n4251 185
R10909 gnd.n4250 gnd.n4249 185
R10910 gnd.n4241 gnd.n4240 185
R10911 gnd.n4244 gnd.n4243 185
R10912 gnd.n459 gnd.n458 185
R10913 gnd.n457 gnd.n456 185
R10914 gnd.n436 gnd.n435 185
R10915 gnd.n451 gnd.n450 185
R10916 gnd.n449 gnd.n448 185
R10917 gnd.n440 gnd.n439 185
R10918 gnd.n443 gnd.n442 185
R10919 gnd.n422 gnd.n421 185
R10920 gnd.n420 gnd.n419 185
R10921 gnd.n399 gnd.n398 185
R10922 gnd.n414 gnd.n413 185
R10923 gnd.n412 gnd.n411 185
R10924 gnd.n403 gnd.n402 185
R10925 gnd.n406 gnd.n405 185
R10926 gnd.n320 gnd.n319 185
R10927 gnd.n318 gnd.n317 185
R10928 gnd.n297 gnd.n296 185
R10929 gnd.n312 gnd.n311 185
R10930 gnd.n310 gnd.n309 185
R10931 gnd.n301 gnd.n300 185
R10932 gnd.n304 gnd.n303 185
R10933 gnd.n283 gnd.n282 185
R10934 gnd.n281 gnd.n280 185
R10935 gnd.n260 gnd.n259 185
R10936 gnd.n275 gnd.n274 185
R10937 gnd.n273 gnd.n272 185
R10938 gnd.n264 gnd.n263 185
R10939 gnd.n267 gnd.n266 185
R10940 gnd.n389 gnd.n388 185
R10941 gnd.n387 gnd.n386 185
R10942 gnd.n366 gnd.n365 185
R10943 gnd.n381 gnd.n380 185
R10944 gnd.n379 gnd.n378 185
R10945 gnd.n370 gnd.n369 185
R10946 gnd.n373 gnd.n372 185
R10947 gnd.n352 gnd.n351 185
R10948 gnd.n350 gnd.n349 185
R10949 gnd.n329 gnd.n328 185
R10950 gnd.n344 gnd.n343 185
R10951 gnd.n342 gnd.n341 185
R10952 gnd.n333 gnd.n332 185
R10953 gnd.n336 gnd.n335 185
R10954 gnd.n4996 gnd.n4995 185
R10955 gnd.n4994 gnd.n4993 185
R10956 gnd.n4973 gnd.n4972 185
R10957 gnd.n4988 gnd.n4987 185
R10958 gnd.n4986 gnd.n4985 185
R10959 gnd.n4977 gnd.n4976 185
R10960 gnd.n4980 gnd.n4979 185
R10961 gnd.n4964 gnd.n4963 185
R10962 gnd.n4962 gnd.n4961 185
R10963 gnd.n4941 gnd.n4940 185
R10964 gnd.n4956 gnd.n4955 185
R10965 gnd.n4954 gnd.n4953 185
R10966 gnd.n4945 gnd.n4944 185
R10967 gnd.n4948 gnd.n4947 185
R10968 gnd.n4932 gnd.n4931 185
R10969 gnd.n4930 gnd.n4929 185
R10970 gnd.n4909 gnd.n4908 185
R10971 gnd.n4924 gnd.n4923 185
R10972 gnd.n4922 gnd.n4921 185
R10973 gnd.n4913 gnd.n4912 185
R10974 gnd.n4916 gnd.n4915 185
R10975 gnd.n4901 gnd.n4900 185
R10976 gnd.n4899 gnd.n4898 185
R10977 gnd.n4878 gnd.n4877 185
R10978 gnd.n4893 gnd.n4892 185
R10979 gnd.n4891 gnd.n4890 185
R10980 gnd.n4882 gnd.n4881 185
R10981 gnd.n4885 gnd.n4884 185
R10982 gnd.n4869 gnd.n4868 185
R10983 gnd.n4867 gnd.n4866 185
R10984 gnd.n4846 gnd.n4845 185
R10985 gnd.n4861 gnd.n4860 185
R10986 gnd.n4859 gnd.n4858 185
R10987 gnd.n4850 gnd.n4849 185
R10988 gnd.n4853 gnd.n4852 185
R10989 gnd.n4837 gnd.n4836 185
R10990 gnd.n4835 gnd.n4834 185
R10991 gnd.n4814 gnd.n4813 185
R10992 gnd.n4829 gnd.n4828 185
R10993 gnd.n4827 gnd.n4826 185
R10994 gnd.n4818 gnd.n4817 185
R10995 gnd.n4821 gnd.n4820 185
R10996 gnd.n4805 gnd.n4804 185
R10997 gnd.n4803 gnd.n4802 185
R10998 gnd.n4782 gnd.n4781 185
R10999 gnd.n4797 gnd.n4796 185
R11000 gnd.n4795 gnd.n4794 185
R11001 gnd.n4786 gnd.n4785 185
R11002 gnd.n4789 gnd.n4788 185
R11003 gnd.n4774 gnd.n4773 185
R11004 gnd.n4772 gnd.n4771 185
R11005 gnd.n4751 gnd.n4750 185
R11006 gnd.n4766 gnd.n4765 185
R11007 gnd.n4764 gnd.n4763 185
R11008 gnd.n4755 gnd.n4754 185
R11009 gnd.n4758 gnd.n4757 185
R11010 gnd.n123 gnd.n122 185
R11011 gnd.n121 gnd.n120 185
R11012 gnd.n100 gnd.n99 185
R11013 gnd.n115 gnd.n114 185
R11014 gnd.n113 gnd.n112 185
R11015 gnd.n104 gnd.n103 185
R11016 gnd.n107 gnd.n106 185
R11017 gnd.n91 gnd.n90 185
R11018 gnd.n89 gnd.n88 185
R11019 gnd.n68 gnd.n67 185
R11020 gnd.n83 gnd.n82 185
R11021 gnd.n81 gnd.n80 185
R11022 gnd.n72 gnd.n71 185
R11023 gnd.n75 gnd.n74 185
R11024 gnd.n59 gnd.n58 185
R11025 gnd.n57 gnd.n56 185
R11026 gnd.n36 gnd.n35 185
R11027 gnd.n51 gnd.n50 185
R11028 gnd.n49 gnd.n48 185
R11029 gnd.n40 gnd.n39 185
R11030 gnd.n43 gnd.n42 185
R11031 gnd.n28 gnd.n27 185
R11032 gnd.n26 gnd.n25 185
R11033 gnd.n5 gnd.n4 185
R11034 gnd.n20 gnd.n19 185
R11035 gnd.n18 gnd.n17 185
R11036 gnd.n9 gnd.n8 185
R11037 gnd.n12 gnd.n11 185
R11038 gnd.n250 gnd.n249 185
R11039 gnd.n248 gnd.n247 185
R11040 gnd.n227 gnd.n226 185
R11041 gnd.n242 gnd.n241 185
R11042 gnd.n240 gnd.n239 185
R11043 gnd.n231 gnd.n230 185
R11044 gnd.n234 gnd.n233 185
R11045 gnd.n218 gnd.n217 185
R11046 gnd.n216 gnd.n215 185
R11047 gnd.n195 gnd.n194 185
R11048 gnd.n210 gnd.n209 185
R11049 gnd.n208 gnd.n207 185
R11050 gnd.n199 gnd.n198 185
R11051 gnd.n202 gnd.n201 185
R11052 gnd.n186 gnd.n185 185
R11053 gnd.n184 gnd.n183 185
R11054 gnd.n163 gnd.n162 185
R11055 gnd.n178 gnd.n177 185
R11056 gnd.n176 gnd.n175 185
R11057 gnd.n167 gnd.n166 185
R11058 gnd.n170 gnd.n169 185
R11059 gnd.n155 gnd.n154 185
R11060 gnd.n153 gnd.n152 185
R11061 gnd.n132 gnd.n131 185
R11062 gnd.n147 gnd.n146 185
R11063 gnd.n145 gnd.n144 185
R11064 gnd.n136 gnd.n135 185
R11065 gnd.n139 gnd.n138 185
R11066 gnd.n1491 gnd.t121 178.987
R11067 gnd.n1160 gnd.t158 178.987
R11068 gnd.n5742 gnd.t205 178.987
R11069 gnd.n1489 gnd.t173 178.987
R11070 gnd.n1155 gnd.t189 178.987
R11071 gnd.n3972 gnd.t198 178.987
R11072 gnd.n3675 gnd.t130 178.987
R11073 gnd.n7236 gnd.t162 178.987
R11074 gnd.n6969 gnd.t136 178.987
R11075 gnd.n1744 gnd.t134 178.987
R11076 gnd.n881 gnd.t111 178.987
R11077 gnd.n901 gnd.t201 178.987
R11078 gnd.n572 gnd.t171 178.987
R11079 gnd.n536 gnd.t186 178.987
R11080 gnd.n2123 gnd.t150 178.987
R11081 gnd.n2052 gnd.t125 178.987
R11082 gnd.n5244 gnd.t153 178.987
R11083 gnd.n1595 gnd.t165 178.987
R11084 gnd.n1560 gnd.t183 178.987
R11085 gnd.n997 gnd.t213 178.987
R11086 gnd.n6604 gnd.n6603 163.367
R11087 gnd.n6601 gnd.n1135 163.367
R11088 gnd.n6597 gnd.n6596 163.367
R11089 gnd.n6594 gnd.n1138 163.367
R11090 gnd.n6590 gnd.n6589 163.367
R11091 gnd.n6587 gnd.n1141 163.367
R11092 gnd.n6583 gnd.n6582 163.367
R11093 gnd.n6580 gnd.n1144 163.367
R11094 gnd.n6576 gnd.n6575 163.367
R11095 gnd.n6573 gnd.n1147 163.367
R11096 gnd.n6569 gnd.n6568 163.367
R11097 gnd.n6566 gnd.n1150 163.367
R11098 gnd.n6562 gnd.n6561 163.367
R11099 gnd.n6559 gnd.n1153 163.367
R11100 gnd.n6555 gnd.n6554 163.367
R11101 gnd.n6550 gnd.n1158 163.367
R11102 gnd.n6546 gnd.n6545 163.367
R11103 gnd.n6543 gnd.n1164 163.367
R11104 gnd.n6539 gnd.n6538 163.367
R11105 gnd.n6536 gnd.n1167 163.367
R11106 gnd.n6532 gnd.n6531 163.367
R11107 gnd.n6529 gnd.n1170 163.367
R11108 gnd.n6525 gnd.n6524 163.367
R11109 gnd.n6522 gnd.n1173 163.367
R11110 gnd.n6518 gnd.n6517 163.367
R11111 gnd.n6515 gnd.n1176 163.367
R11112 gnd.n6511 gnd.n6510 163.367
R11113 gnd.n6508 gnd.n1179 163.367
R11114 gnd.n6504 gnd.n6503 163.367
R11115 gnd.n1498 gnd.n1497 163.367
R11116 gnd.n1497 gnd.n1405 163.367
R11117 gnd.n6130 gnd.n1405 163.367
R11118 gnd.n6130 gnd.n1400 163.367
R11119 gnd.n6126 gnd.n1400 163.367
R11120 gnd.n6126 gnd.n1408 163.367
R11121 gnd.n6091 gnd.n1408 163.367
R11122 gnd.n6091 gnd.n1381 163.367
R11123 gnd.n1382 gnd.n1381 163.367
R11124 gnd.n1382 gnd.n1375 163.367
R11125 gnd.n6097 gnd.n1375 163.367
R11126 gnd.n6097 gnd.n1367 163.367
R11127 gnd.n6100 gnd.n1367 163.367
R11128 gnd.n6100 gnd.n1361 163.367
R11129 gnd.n6105 gnd.n1361 163.367
R11130 gnd.n6105 gnd.n1349 163.367
R11131 gnd.n1349 gnd.n1341 163.367
R11132 gnd.n6221 gnd.n1341 163.367
R11133 gnd.n6221 gnd.n1339 163.367
R11134 gnd.n6226 gnd.n1339 163.367
R11135 gnd.n6226 gnd.n1325 163.367
R11136 gnd.n6251 gnd.n1325 163.367
R11137 gnd.n6252 gnd.n6251 163.367
R11138 gnd.n6252 gnd.n1331 163.367
R11139 gnd.n6258 gnd.n1331 163.367
R11140 gnd.n6258 gnd.n1305 163.367
R11141 gnd.n1305 gnd.n1298 163.367
R11142 gnd.n6311 gnd.n1298 163.367
R11143 gnd.n6312 gnd.n6311 163.367
R11144 gnd.n6312 gnd.n1287 163.367
R11145 gnd.n1295 gnd.n1287 163.367
R11146 gnd.n6324 gnd.n1295 163.367
R11147 gnd.n6324 gnd.n1296 163.367
R11148 gnd.n1296 gnd.n1264 163.367
R11149 gnd.n6319 gnd.n1264 163.367
R11150 gnd.n6319 gnd.n1257 163.367
R11151 gnd.n6316 gnd.n1257 163.367
R11152 gnd.n6316 gnd.n1247 163.367
R11153 gnd.n6411 gnd.n1247 163.367
R11154 gnd.n6411 gnd.n1235 163.367
R11155 gnd.n6414 gnd.n1235 163.367
R11156 gnd.n6414 gnd.n1229 163.367
R11157 gnd.n6418 gnd.n1229 163.367
R11158 gnd.n6418 gnd.n1219 163.367
R11159 gnd.n6448 gnd.n1219 163.367
R11160 gnd.n6448 gnd.n1207 163.367
R11161 gnd.n6451 gnd.n1207 163.367
R11162 gnd.n6451 gnd.n1201 163.367
R11163 gnd.n6458 gnd.n1201 163.367
R11164 gnd.n6458 gnd.n1189 163.367
R11165 gnd.n6454 gnd.n1189 163.367
R11166 gnd.n6454 gnd.n1185 163.367
R11167 gnd.n6496 gnd.n1185 163.367
R11168 gnd.n6496 gnd.n1110 163.367
R11169 gnd.n1183 gnd.n1110 163.367
R11170 gnd.n1464 gnd.n1463 163.367
R11171 gnd.n6052 gnd.n1463 163.367
R11172 gnd.n6050 gnd.n6049 163.367
R11173 gnd.n6046 gnd.n6045 163.367
R11174 gnd.n6042 gnd.n6041 163.367
R11175 gnd.n6038 gnd.n6037 163.367
R11176 gnd.n6034 gnd.n6033 163.367
R11177 gnd.n6030 gnd.n6029 163.367
R11178 gnd.n6026 gnd.n6025 163.367
R11179 gnd.n6022 gnd.n6021 163.367
R11180 gnd.n6018 gnd.n6017 163.367
R11181 gnd.n6014 gnd.n6013 163.367
R11182 gnd.n6010 gnd.n6009 163.367
R11183 gnd.n6005 gnd.n6004 163.367
R11184 gnd.n6001 gnd.n6000 163.367
R11185 gnd.n1555 gnd.n1554 163.367
R11186 gnd.n1551 gnd.n1550 163.367
R11187 gnd.n1547 gnd.n1546 163.367
R11188 gnd.n1543 gnd.n1542 163.367
R11189 gnd.n1539 gnd.n1538 163.367
R11190 gnd.n1535 gnd.n1534 163.367
R11191 gnd.n1531 gnd.n1530 163.367
R11192 gnd.n1527 gnd.n1526 163.367
R11193 gnd.n1523 gnd.n1522 163.367
R11194 gnd.n1519 gnd.n1518 163.367
R11195 gnd.n1515 gnd.n1514 163.367
R11196 gnd.n1511 gnd.n1510 163.367
R11197 gnd.n1507 gnd.n1506 163.367
R11198 gnd.n1503 gnd.n1502 163.367
R11199 gnd.n1465 gnd.n1404 163.367
R11200 gnd.n6134 gnd.n1404 163.367
R11201 gnd.n6134 gnd.n1401 163.367
R11202 gnd.n6141 gnd.n1401 163.367
R11203 gnd.n6141 gnd.n1402 163.367
R11204 gnd.n6137 gnd.n1402 163.367
R11205 gnd.n6137 gnd.n1379 163.367
R11206 gnd.n6165 gnd.n1379 163.367
R11207 gnd.n6165 gnd.n1377 163.367
R11208 gnd.n6169 gnd.n1377 163.367
R11209 gnd.n6169 gnd.n1365 163.367
R11210 gnd.n6197 gnd.n1365 163.367
R11211 gnd.n6197 gnd.n1363 163.367
R11212 gnd.n6201 gnd.n1363 163.367
R11213 gnd.n6201 gnd.n1347 163.367
R11214 gnd.n6214 gnd.n1347 163.367
R11215 gnd.n6214 gnd.n1344 163.367
R11216 gnd.n6219 gnd.n1344 163.367
R11217 gnd.n6219 gnd.n1345 163.367
R11218 gnd.n1345 gnd.n1327 163.367
R11219 gnd.n6267 gnd.n1327 163.367
R11220 gnd.n6267 gnd.n1328 163.367
R11221 gnd.n6263 gnd.n1328 163.367
R11222 gnd.n6263 gnd.n6262 163.367
R11223 gnd.n6262 gnd.n1303 163.367
R11224 gnd.n6305 gnd.n1303 163.367
R11225 gnd.n6305 gnd.n1301 163.367
R11226 gnd.n6309 gnd.n1301 163.367
R11227 gnd.n6309 gnd.n1289 163.367
R11228 gnd.n6330 gnd.n1289 163.367
R11229 gnd.n6330 gnd.n1290 163.367
R11230 gnd.n6326 gnd.n1290 163.367
R11231 gnd.n6326 gnd.n1262 163.367
R11232 gnd.n6392 gnd.n1262 163.367
R11233 gnd.n6392 gnd.n1259 163.367
R11234 gnd.n6399 gnd.n1259 163.367
R11235 gnd.n6399 gnd.n1260 163.367
R11236 gnd.n6395 gnd.n1260 163.367
R11237 gnd.n6395 gnd.n1233 163.367
R11238 gnd.n6428 gnd.n1233 163.367
R11239 gnd.n6428 gnd.n1230 163.367
R11240 gnd.n6435 gnd.n1230 163.367
R11241 gnd.n6435 gnd.n1231 163.367
R11242 gnd.n6431 gnd.n1231 163.367
R11243 gnd.n6431 gnd.n1205 163.367
R11244 gnd.n6468 gnd.n1205 163.367
R11245 gnd.n6468 gnd.n1203 163.367
R11246 gnd.n6472 gnd.n1203 163.367
R11247 gnd.n6472 gnd.n1188 163.367
R11248 gnd.n6488 gnd.n1188 163.367
R11249 gnd.n6488 gnd.n1186 163.367
R11250 gnd.n6492 gnd.n1186 163.367
R11251 gnd.n6492 gnd.n1112 163.367
R11252 gnd.n6609 gnd.n1112 163.367
R11253 gnd.n6609 gnd.n1113 163.367
R11254 gnd.n1133 gnd.n1132 156.462
R11255 gnd.n4936 gnd.n4904 153.042
R11256 gnd.n63 gnd.n31 153.042
R11257 gnd.n5000 gnd.n4999 152.079
R11258 gnd.n4968 gnd.n4967 152.079
R11259 gnd.n4936 gnd.n4935 152.079
R11260 gnd.n127 gnd.n126 152.079
R11261 gnd.n95 gnd.n94 152.079
R11262 gnd.n63 gnd.n62 152.079
R11263 gnd.n1478 gnd.n1477 152
R11264 gnd.n1479 gnd.n1468 152
R11265 gnd.n1481 gnd.n1480 152
R11266 gnd.n1483 gnd.n1466 152
R11267 gnd.n1485 gnd.n1484 152
R11268 gnd.n1131 gnd.n1115 152
R11269 gnd.n1123 gnd.n1116 152
R11270 gnd.n1122 gnd.n1121 152
R11271 gnd.n1120 gnd.n1117 152
R11272 gnd.n1118 gnd.t207 150.546
R11273 gnd.t97 gnd.n4275 147.661
R11274 gnd.t95 gnd.n4312 147.661
R11275 gnd.t55 gnd.n4136 147.661
R11276 gnd.t76 gnd.n4173 147.661
R11277 gnd.t107 gnd.n4205 147.661
R11278 gnd.t66 gnd.n4242 147.661
R11279 gnd.t96 gnd.n441 147.661
R11280 gnd.t99 gnd.n404 147.661
R11281 gnd.t100 gnd.n302 147.661
R11282 gnd.t79 gnd.n265 147.661
R11283 gnd.t88 gnd.n371 147.661
R11284 gnd.t69 gnd.n334 147.661
R11285 gnd.t36 gnd.n4978 147.661
R11286 gnd.t34 gnd.n4946 147.661
R11287 gnd.t32 gnd.n4914 147.661
R11288 gnd.t30 gnd.n4883 147.661
R11289 gnd.t28 gnd.n4851 147.661
R11290 gnd.t40 gnd.n4819 147.661
R11291 gnd.t44 gnd.n4787 147.661
R11292 gnd.t42 gnd.n4756 147.661
R11293 gnd.t5 gnd.n105 147.661
R11294 gnd.t38 gnd.n73 147.661
R11295 gnd.t7 gnd.n41 147.661
R11296 gnd.t1 gnd.n10 147.661
R11297 gnd.t219 gnd.n232 147.661
R11298 gnd.t26 gnd.n200 147.661
R11299 gnd.t14 gnd.n168 147.661
R11300 gnd.t3 gnd.n137 147.661
R11301 gnd.n6553 gnd.n6552 143.351
R11302 gnd.n6552 gnd.n6551 143.351
R11303 gnd.n5998 gnd.n1447 143.351
R11304 gnd.n5998 gnd.n1448 143.351
R11305 gnd.n1475 gnd.t116 130.484
R11306 gnd.n1484 gnd.t178 126.766
R11307 gnd.n1482 gnd.t190 126.766
R11308 gnd.n1468 gnd.t166 126.766
R11309 gnd.n1476 gnd.t214 126.766
R11310 gnd.n1119 gnd.t138 126.766
R11311 gnd.n1121 gnd.t113 126.766
R11312 gnd.n1130 gnd.t175 126.766
R11313 gnd.n1132 gnd.t193 126.766
R11314 gnd.n6937 gnd.n877 110.912
R11315 gnd.n5999 gnd.n5997 110.912
R11316 gnd.n4292 gnd.n4291 104.615
R11317 gnd.n4291 gnd.n4269 104.615
R11318 gnd.n4284 gnd.n4269 104.615
R11319 gnd.n4284 gnd.n4283 104.615
R11320 gnd.n4283 gnd.n4273 104.615
R11321 gnd.n4276 gnd.n4273 104.615
R11322 gnd.n4329 gnd.n4328 104.615
R11323 gnd.n4328 gnd.n4306 104.615
R11324 gnd.n4321 gnd.n4306 104.615
R11325 gnd.n4321 gnd.n4320 104.615
R11326 gnd.n4320 gnd.n4310 104.615
R11327 gnd.n4313 gnd.n4310 104.615
R11328 gnd.n4153 gnd.n4152 104.615
R11329 gnd.n4152 gnd.n4130 104.615
R11330 gnd.n4145 gnd.n4130 104.615
R11331 gnd.n4145 gnd.n4144 104.615
R11332 gnd.n4144 gnd.n4134 104.615
R11333 gnd.n4137 gnd.n4134 104.615
R11334 gnd.n4190 gnd.n4189 104.615
R11335 gnd.n4189 gnd.n4167 104.615
R11336 gnd.n4182 gnd.n4167 104.615
R11337 gnd.n4182 gnd.n4181 104.615
R11338 gnd.n4181 gnd.n4171 104.615
R11339 gnd.n4174 gnd.n4171 104.615
R11340 gnd.n4222 gnd.n4221 104.615
R11341 gnd.n4221 gnd.n4199 104.615
R11342 gnd.n4214 gnd.n4199 104.615
R11343 gnd.n4214 gnd.n4213 104.615
R11344 gnd.n4213 gnd.n4203 104.615
R11345 gnd.n4206 gnd.n4203 104.615
R11346 gnd.n4259 gnd.n4258 104.615
R11347 gnd.n4258 gnd.n4236 104.615
R11348 gnd.n4251 gnd.n4236 104.615
R11349 gnd.n4251 gnd.n4250 104.615
R11350 gnd.n4250 gnd.n4240 104.615
R11351 gnd.n4243 gnd.n4240 104.615
R11352 gnd.n458 gnd.n457 104.615
R11353 gnd.n457 gnd.n435 104.615
R11354 gnd.n450 gnd.n435 104.615
R11355 gnd.n450 gnd.n449 104.615
R11356 gnd.n449 gnd.n439 104.615
R11357 gnd.n442 gnd.n439 104.615
R11358 gnd.n421 gnd.n420 104.615
R11359 gnd.n420 gnd.n398 104.615
R11360 gnd.n413 gnd.n398 104.615
R11361 gnd.n413 gnd.n412 104.615
R11362 gnd.n412 gnd.n402 104.615
R11363 gnd.n405 gnd.n402 104.615
R11364 gnd.n319 gnd.n318 104.615
R11365 gnd.n318 gnd.n296 104.615
R11366 gnd.n311 gnd.n296 104.615
R11367 gnd.n311 gnd.n310 104.615
R11368 gnd.n310 gnd.n300 104.615
R11369 gnd.n303 gnd.n300 104.615
R11370 gnd.n282 gnd.n281 104.615
R11371 gnd.n281 gnd.n259 104.615
R11372 gnd.n274 gnd.n259 104.615
R11373 gnd.n274 gnd.n273 104.615
R11374 gnd.n273 gnd.n263 104.615
R11375 gnd.n266 gnd.n263 104.615
R11376 gnd.n388 gnd.n387 104.615
R11377 gnd.n387 gnd.n365 104.615
R11378 gnd.n380 gnd.n365 104.615
R11379 gnd.n380 gnd.n379 104.615
R11380 gnd.n379 gnd.n369 104.615
R11381 gnd.n372 gnd.n369 104.615
R11382 gnd.n351 gnd.n350 104.615
R11383 gnd.n350 gnd.n328 104.615
R11384 gnd.n343 gnd.n328 104.615
R11385 gnd.n343 gnd.n342 104.615
R11386 gnd.n342 gnd.n332 104.615
R11387 gnd.n335 gnd.n332 104.615
R11388 gnd.n4995 gnd.n4994 104.615
R11389 gnd.n4994 gnd.n4972 104.615
R11390 gnd.n4987 gnd.n4972 104.615
R11391 gnd.n4987 gnd.n4986 104.615
R11392 gnd.n4986 gnd.n4976 104.615
R11393 gnd.n4979 gnd.n4976 104.615
R11394 gnd.n4963 gnd.n4962 104.615
R11395 gnd.n4962 gnd.n4940 104.615
R11396 gnd.n4955 gnd.n4940 104.615
R11397 gnd.n4955 gnd.n4954 104.615
R11398 gnd.n4954 gnd.n4944 104.615
R11399 gnd.n4947 gnd.n4944 104.615
R11400 gnd.n4931 gnd.n4930 104.615
R11401 gnd.n4930 gnd.n4908 104.615
R11402 gnd.n4923 gnd.n4908 104.615
R11403 gnd.n4923 gnd.n4922 104.615
R11404 gnd.n4922 gnd.n4912 104.615
R11405 gnd.n4915 gnd.n4912 104.615
R11406 gnd.n4900 gnd.n4899 104.615
R11407 gnd.n4899 gnd.n4877 104.615
R11408 gnd.n4892 gnd.n4877 104.615
R11409 gnd.n4892 gnd.n4891 104.615
R11410 gnd.n4891 gnd.n4881 104.615
R11411 gnd.n4884 gnd.n4881 104.615
R11412 gnd.n4868 gnd.n4867 104.615
R11413 gnd.n4867 gnd.n4845 104.615
R11414 gnd.n4860 gnd.n4845 104.615
R11415 gnd.n4860 gnd.n4859 104.615
R11416 gnd.n4859 gnd.n4849 104.615
R11417 gnd.n4852 gnd.n4849 104.615
R11418 gnd.n4836 gnd.n4835 104.615
R11419 gnd.n4835 gnd.n4813 104.615
R11420 gnd.n4828 gnd.n4813 104.615
R11421 gnd.n4828 gnd.n4827 104.615
R11422 gnd.n4827 gnd.n4817 104.615
R11423 gnd.n4820 gnd.n4817 104.615
R11424 gnd.n4804 gnd.n4803 104.615
R11425 gnd.n4803 gnd.n4781 104.615
R11426 gnd.n4796 gnd.n4781 104.615
R11427 gnd.n4796 gnd.n4795 104.615
R11428 gnd.n4795 gnd.n4785 104.615
R11429 gnd.n4788 gnd.n4785 104.615
R11430 gnd.n4773 gnd.n4772 104.615
R11431 gnd.n4772 gnd.n4750 104.615
R11432 gnd.n4765 gnd.n4750 104.615
R11433 gnd.n4765 gnd.n4764 104.615
R11434 gnd.n4764 gnd.n4754 104.615
R11435 gnd.n4757 gnd.n4754 104.615
R11436 gnd.n122 gnd.n121 104.615
R11437 gnd.n121 gnd.n99 104.615
R11438 gnd.n114 gnd.n99 104.615
R11439 gnd.n114 gnd.n113 104.615
R11440 gnd.n113 gnd.n103 104.615
R11441 gnd.n106 gnd.n103 104.615
R11442 gnd.n90 gnd.n89 104.615
R11443 gnd.n89 gnd.n67 104.615
R11444 gnd.n82 gnd.n67 104.615
R11445 gnd.n82 gnd.n81 104.615
R11446 gnd.n81 gnd.n71 104.615
R11447 gnd.n74 gnd.n71 104.615
R11448 gnd.n58 gnd.n57 104.615
R11449 gnd.n57 gnd.n35 104.615
R11450 gnd.n50 gnd.n35 104.615
R11451 gnd.n50 gnd.n49 104.615
R11452 gnd.n49 gnd.n39 104.615
R11453 gnd.n42 gnd.n39 104.615
R11454 gnd.n27 gnd.n26 104.615
R11455 gnd.n26 gnd.n4 104.615
R11456 gnd.n19 gnd.n4 104.615
R11457 gnd.n19 gnd.n18 104.615
R11458 gnd.n18 gnd.n8 104.615
R11459 gnd.n11 gnd.n8 104.615
R11460 gnd.n249 gnd.n248 104.615
R11461 gnd.n248 gnd.n226 104.615
R11462 gnd.n241 gnd.n226 104.615
R11463 gnd.n241 gnd.n240 104.615
R11464 gnd.n240 gnd.n230 104.615
R11465 gnd.n233 gnd.n230 104.615
R11466 gnd.n217 gnd.n216 104.615
R11467 gnd.n216 gnd.n194 104.615
R11468 gnd.n209 gnd.n194 104.615
R11469 gnd.n209 gnd.n208 104.615
R11470 gnd.n208 gnd.n198 104.615
R11471 gnd.n201 gnd.n198 104.615
R11472 gnd.n185 gnd.n184 104.615
R11473 gnd.n184 gnd.n162 104.615
R11474 gnd.n177 gnd.n162 104.615
R11475 gnd.n177 gnd.n176 104.615
R11476 gnd.n176 gnd.n166 104.615
R11477 gnd.n169 gnd.n166 104.615
R11478 gnd.n154 gnd.n153 104.615
R11479 gnd.n153 gnd.n131 104.615
R11480 gnd.n146 gnd.n131 104.615
R11481 gnd.n146 gnd.n145 104.615
R11482 gnd.n145 gnd.n135 104.615
R11483 gnd.n138 gnd.n135 104.615
R11484 gnd.n4396 gnd.t148 100.632
R11485 gnd.n3648 gnd.t143 100.632
R11486 gnd.n7345 gnd.n512 99.6594
R11487 gnd.n7343 gnd.n7342 99.6594
R11488 gnd.n7338 gnd.n519 99.6594
R11489 gnd.n7336 gnd.n7335 99.6594
R11490 gnd.n7331 gnd.n526 99.6594
R11491 gnd.n7329 gnd.n7328 99.6594
R11492 gnd.n7324 gnd.n533 99.6594
R11493 gnd.n7322 gnd.n7321 99.6594
R11494 gnd.n7317 gnd.n543 99.6594
R11495 gnd.n7315 gnd.n7314 99.6594
R11496 gnd.n7310 gnd.n550 99.6594
R11497 gnd.n7308 gnd.n7307 99.6594
R11498 gnd.n7303 gnd.n557 99.6594
R11499 gnd.n7301 gnd.n7300 99.6594
R11500 gnd.n7296 gnd.n564 99.6594
R11501 gnd.n7294 gnd.n7293 99.6594
R11502 gnd.n569 gnd.n568 99.6594
R11503 gnd.n6963 gnd.n785 99.6594
R11504 gnd.n6958 gnd.n834 99.6594
R11505 gnd.n6955 gnd.n835 99.6594
R11506 gnd.n6951 gnd.n836 99.6594
R11507 gnd.n6947 gnd.n837 99.6594
R11508 gnd.n6943 gnd.n838 99.6594
R11509 gnd.n6939 gnd.n839 99.6594
R11510 gnd.n6934 gnd.n841 99.6594
R11511 gnd.n6930 gnd.n842 99.6594
R11512 gnd.n6926 gnd.n843 99.6594
R11513 gnd.n6922 gnd.n844 99.6594
R11514 gnd.n6918 gnd.n845 99.6594
R11515 gnd.n6914 gnd.n846 99.6594
R11516 gnd.n6910 gnd.n847 99.6594
R11517 gnd.n6906 gnd.n848 99.6594
R11518 gnd.n899 gnd.n849 99.6594
R11519 gnd.n5950 gnd.n5949 99.6594
R11520 gnd.n5947 gnd.n5946 99.6594
R11521 gnd.n5942 gnd.n5919 99.6594
R11522 gnd.n5940 gnd.n5939 99.6594
R11523 gnd.n5935 gnd.n5926 99.6594
R11524 gnd.n5933 gnd.n5932 99.6594
R11525 gnd.n1566 gnd.n1565 99.6594
R11526 gnd.n5991 gnd.n5990 99.6594
R11527 gnd.n5988 gnd.n5987 99.6594
R11528 gnd.n5983 gnd.n1575 99.6594
R11529 gnd.n5981 gnd.n5980 99.6594
R11530 gnd.n5976 gnd.n1582 99.6594
R11531 gnd.n5974 gnd.n5973 99.6594
R11532 gnd.n5969 gnd.n1589 99.6594
R11533 gnd.n5967 gnd.n5966 99.6594
R11534 gnd.n1600 gnd.n1599 99.6594
R11535 gnd.n2086 gnd.n2011 99.6594
R11536 gnd.n2094 gnd.n2093 99.6594
R11537 gnd.n2097 gnd.n2096 99.6594
R11538 gnd.n2104 gnd.n2103 99.6594
R11539 gnd.n2107 gnd.n2106 99.6594
R11540 gnd.n2114 gnd.n2113 99.6594
R11541 gnd.n2117 gnd.n2116 99.6594
R11542 gnd.n2127 gnd.n2126 99.6594
R11543 gnd.n2130 gnd.n2129 99.6594
R11544 gnd.n2137 gnd.n2136 99.6594
R11545 gnd.n2140 gnd.n2139 99.6594
R11546 gnd.n2147 gnd.n2146 99.6594
R11547 gnd.n2150 gnd.n2149 99.6594
R11548 gnd.n2157 gnd.n2156 99.6594
R11549 gnd.n2160 gnd.n2159 99.6594
R11550 gnd.n2168 gnd.n2167 99.6594
R11551 gnd.n2171 gnd.n2170 99.6594
R11552 gnd.n5115 gnd.n5114 99.6594
R11553 gnd.n5110 gnd.n3626 99.6594
R11554 gnd.n5106 gnd.n3625 99.6594
R11555 gnd.n5102 gnd.n3624 99.6594
R11556 gnd.n5098 gnd.n3623 99.6594
R11557 gnd.n5094 gnd.n3622 99.6594
R11558 gnd.n5090 gnd.n3621 99.6594
R11559 gnd.n3646 gnd.n3620 99.6594
R11560 gnd.n4429 gnd.n4428 99.6594
R11561 gnd.n4423 gnd.n4371 99.6594
R11562 gnd.n4420 gnd.n4372 99.6594
R11563 gnd.n4416 gnd.n4373 99.6594
R11564 gnd.n4412 gnd.n4374 99.6594
R11565 gnd.n4408 gnd.n4375 99.6594
R11566 gnd.n4404 gnd.n4376 99.6594
R11567 gnd.n4400 gnd.n4377 99.6594
R11568 gnd.n5080 gnd.n3607 99.6594
R11569 gnd.n5076 gnd.n3608 99.6594
R11570 gnd.n5072 gnd.n3609 99.6594
R11571 gnd.n5068 gnd.n3610 99.6594
R11572 gnd.n5064 gnd.n3611 99.6594
R11573 gnd.n5060 gnd.n3612 99.6594
R11574 gnd.n5056 gnd.n3613 99.6594
R11575 gnd.n5052 gnd.n3614 99.6594
R11576 gnd.n5048 gnd.n3615 99.6594
R11577 gnd.n5044 gnd.n3616 99.6594
R11578 gnd.n5040 gnd.n3617 99.6594
R11579 gnd.n5036 gnd.n3618 99.6594
R11580 gnd.n5032 gnd.n3619 99.6594
R11581 gnd.n4026 gnd.n3936 99.6594
R11582 gnd.n4024 gnd.n3939 99.6594
R11583 gnd.n4020 gnd.n4019 99.6594
R11584 gnd.n4013 gnd.n3944 99.6594
R11585 gnd.n4012 gnd.n4011 99.6594
R11586 gnd.n4005 gnd.n3950 99.6594
R11587 gnd.n4004 gnd.n4003 99.6594
R11588 gnd.n3997 gnd.n3956 99.6594
R11589 gnd.n3996 gnd.n3995 99.6594
R11590 gnd.n3989 gnd.n3962 99.6594
R11591 gnd.n3988 gnd.n3987 99.6594
R11592 gnd.n3980 gnd.n3968 99.6594
R11593 gnd.n3979 gnd.n3978 99.6594
R11594 gnd.n7210 gnd.n7209 99.6594
R11595 gnd.n7215 gnd.n7214 99.6594
R11596 gnd.n7218 gnd.n7217 99.6594
R11597 gnd.n7223 gnd.n7222 99.6594
R11598 gnd.n7226 gnd.n7225 99.6594
R11599 gnd.n7231 gnd.n7230 99.6594
R11600 gnd.n7234 gnd.n7233 99.6594
R11601 gnd.n7237 gnd.n499 99.6594
R11602 gnd.n850 gnd.n790 99.6594
R11603 gnd.n852 gnd.n851 99.6594
R11604 gnd.n854 gnd.n800 99.6594
R11605 gnd.n855 gnd.n807 99.6594
R11606 gnd.n857 gnd.n856 99.6594
R11607 gnd.n859 gnd.n816 99.6594
R11608 gnd.n860 gnd.n823 99.6594
R11609 gnd.n6966 gnd.n6965 99.6594
R11610 gnd.n1699 gnd.n1698 99.6594
R11611 gnd.n1702 gnd.n1701 99.6594
R11612 gnd.n1712 gnd.n1711 99.6594
R11613 gnd.n1721 gnd.n1720 99.6594
R11614 gnd.n1724 gnd.n1723 99.6594
R11615 gnd.n1735 gnd.n1734 99.6594
R11616 gnd.n1746 gnd.n1745 99.6594
R11617 gnd.n5768 gnd.n5767 99.6594
R11618 gnd.n5273 gnd.n2015 99.6594
R11619 gnd.n5272 gnd.n5271 99.6594
R11620 gnd.n5265 gnd.n2018 99.6594
R11621 gnd.n5264 gnd.n5263 99.6594
R11622 gnd.n5257 gnd.n2024 99.6594
R11623 gnd.n5256 gnd.n5255 99.6594
R11624 gnd.n5249 gnd.n2030 99.6594
R11625 gnd.n5248 gnd.n5247 99.6594
R11626 gnd.n5274 gnd.n5273 99.6594
R11627 gnd.n5271 gnd.n5270 99.6594
R11628 gnd.n5266 gnd.n5265 99.6594
R11629 gnd.n5263 gnd.n5262 99.6594
R11630 gnd.n5258 gnd.n5257 99.6594
R11631 gnd.n5255 gnd.n5254 99.6594
R11632 gnd.n5250 gnd.n5249 99.6594
R11633 gnd.n5247 gnd.n5246 99.6594
R11634 gnd.n5767 gnd.n1747 99.6594
R11635 gnd.n1745 gnd.n1736 99.6594
R11636 gnd.n1734 gnd.n1733 99.6594
R11637 gnd.n1723 gnd.n1722 99.6594
R11638 gnd.n1720 gnd.n1713 99.6594
R11639 gnd.n1711 gnd.n1710 99.6594
R11640 gnd.n1701 gnd.n1700 99.6594
R11641 gnd.n1698 gnd.n1697 99.6594
R11642 gnd.n850 gnd.n792 99.6594
R11643 gnd.n852 gnd.n799 99.6594
R11644 gnd.n854 gnd.n853 99.6594
R11645 gnd.n855 gnd.n808 99.6594
R11646 gnd.n857 gnd.n815 99.6594
R11647 gnd.n859 gnd.n858 99.6594
R11648 gnd.n860 gnd.n824 99.6594
R11649 gnd.n6967 gnd.n6966 99.6594
R11650 gnd.n7238 gnd.n7237 99.6594
R11651 gnd.n7233 gnd.n7232 99.6594
R11652 gnd.n7230 gnd.n7229 99.6594
R11653 gnd.n7225 gnd.n7224 99.6594
R11654 gnd.n7222 gnd.n7221 99.6594
R11655 gnd.n7217 gnd.n7216 99.6594
R11656 gnd.n7214 gnd.n7213 99.6594
R11657 gnd.n7209 gnd.n7208 99.6594
R11658 gnd.n4027 gnd.n4026 99.6594
R11659 gnd.n4021 gnd.n3939 99.6594
R11660 gnd.n4019 gnd.n4018 99.6594
R11661 gnd.n4014 gnd.n4013 99.6594
R11662 gnd.n4011 gnd.n4010 99.6594
R11663 gnd.n4006 gnd.n4005 99.6594
R11664 gnd.n4003 gnd.n4002 99.6594
R11665 gnd.n3998 gnd.n3997 99.6594
R11666 gnd.n3995 gnd.n3994 99.6594
R11667 gnd.n3990 gnd.n3989 99.6594
R11668 gnd.n3987 gnd.n3986 99.6594
R11669 gnd.n3981 gnd.n3980 99.6594
R11670 gnd.n3978 gnd.n3934 99.6594
R11671 gnd.n5035 gnd.n3619 99.6594
R11672 gnd.n5039 gnd.n3618 99.6594
R11673 gnd.n5043 gnd.n3617 99.6594
R11674 gnd.n5047 gnd.n3616 99.6594
R11675 gnd.n5051 gnd.n3615 99.6594
R11676 gnd.n5055 gnd.n3614 99.6594
R11677 gnd.n5059 gnd.n3613 99.6594
R11678 gnd.n5063 gnd.n3612 99.6594
R11679 gnd.n5067 gnd.n3611 99.6594
R11680 gnd.n5071 gnd.n3610 99.6594
R11681 gnd.n5075 gnd.n3609 99.6594
R11682 gnd.n5079 gnd.n3608 99.6594
R11683 gnd.n3652 gnd.n3607 99.6594
R11684 gnd.n4429 gnd.n4379 99.6594
R11685 gnd.n4421 gnd.n4371 99.6594
R11686 gnd.n4417 gnd.n4372 99.6594
R11687 gnd.n4413 gnd.n4373 99.6594
R11688 gnd.n4409 gnd.n4374 99.6594
R11689 gnd.n4405 gnd.n4375 99.6594
R11690 gnd.n4401 gnd.n4376 99.6594
R11691 gnd.n4377 gnd.n3896 99.6594
R11692 gnd.n5089 gnd.n3620 99.6594
R11693 gnd.n5093 gnd.n3621 99.6594
R11694 gnd.n5097 gnd.n3622 99.6594
R11695 gnd.n5101 gnd.n3623 99.6594
R11696 gnd.n5105 gnd.n3624 99.6594
R11697 gnd.n5109 gnd.n3625 99.6594
R11698 gnd.n3628 gnd.n3626 99.6594
R11699 gnd.n5115 gnd.n3627 99.6594
R11700 gnd.n2087 gnd.n2086 99.6594
R11701 gnd.n2095 gnd.n2094 99.6594
R11702 gnd.n2096 gnd.n2079 99.6594
R11703 gnd.n2105 gnd.n2104 99.6594
R11704 gnd.n2106 gnd.n2075 99.6594
R11705 gnd.n2115 gnd.n2114 99.6594
R11706 gnd.n2116 gnd.n2071 99.6594
R11707 gnd.n2128 gnd.n2127 99.6594
R11708 gnd.n2129 gnd.n2067 99.6594
R11709 gnd.n2138 gnd.n2137 99.6594
R11710 gnd.n2139 gnd.n2063 99.6594
R11711 gnd.n2148 gnd.n2147 99.6594
R11712 gnd.n2149 gnd.n2059 99.6594
R11713 gnd.n2158 gnd.n2157 99.6594
R11714 gnd.n2159 gnd.n2055 99.6594
R11715 gnd.n2169 gnd.n2168 99.6594
R11716 gnd.n2172 gnd.n2171 99.6594
R11717 gnd.n1599 gnd.n1590 99.6594
R11718 gnd.n5968 gnd.n5967 99.6594
R11719 gnd.n1589 gnd.n1583 99.6594
R11720 gnd.n5975 gnd.n5974 99.6594
R11721 gnd.n1582 gnd.n1576 99.6594
R11722 gnd.n5982 gnd.n5981 99.6594
R11723 gnd.n1575 gnd.n1569 99.6594
R11724 gnd.n5989 gnd.n5988 99.6594
R11725 gnd.n5992 gnd.n5991 99.6594
R11726 gnd.n5928 gnd.n5927 99.6594
R11727 gnd.n5934 gnd.n5933 99.6594
R11728 gnd.n5926 gnd.n5920 99.6594
R11729 gnd.n5941 gnd.n5940 99.6594
R11730 gnd.n5919 gnd.n5912 99.6594
R11731 gnd.n5948 gnd.n5947 99.6594
R11732 gnd.n5951 gnd.n5950 99.6594
R11733 gnd.n6963 gnd.n6962 99.6594
R11734 gnd.n6956 gnd.n834 99.6594
R11735 gnd.n6952 gnd.n835 99.6594
R11736 gnd.n6948 gnd.n836 99.6594
R11737 gnd.n6944 gnd.n837 99.6594
R11738 gnd.n6940 gnd.n838 99.6594
R11739 gnd.n6935 gnd.n840 99.6594
R11740 gnd.n6931 gnd.n841 99.6594
R11741 gnd.n6927 gnd.n842 99.6594
R11742 gnd.n6923 gnd.n843 99.6594
R11743 gnd.n6919 gnd.n844 99.6594
R11744 gnd.n6915 gnd.n845 99.6594
R11745 gnd.n6911 gnd.n846 99.6594
R11746 gnd.n6907 gnd.n847 99.6594
R11747 gnd.n898 gnd.n848 99.6594
R11748 gnd.n6899 gnd.n849 99.6594
R11749 gnd.n568 gnd.n565 99.6594
R11750 gnd.n7295 gnd.n7294 99.6594
R11751 gnd.n564 gnd.n558 99.6594
R11752 gnd.n7302 gnd.n7301 99.6594
R11753 gnd.n557 gnd.n551 99.6594
R11754 gnd.n7309 gnd.n7308 99.6594
R11755 gnd.n550 gnd.n544 99.6594
R11756 gnd.n7316 gnd.n7315 99.6594
R11757 gnd.n543 gnd.n534 99.6594
R11758 gnd.n7323 gnd.n7322 99.6594
R11759 gnd.n533 gnd.n527 99.6594
R11760 gnd.n7330 gnd.n7329 99.6594
R11761 gnd.n526 gnd.n520 99.6594
R11762 gnd.n7337 gnd.n7336 99.6594
R11763 gnd.n519 gnd.n513 99.6594
R11764 gnd.n7344 gnd.n7343 99.6594
R11765 gnd.n512 gnd.n509 99.6594
R11766 gnd.n5808 gnd.n5807 99.6594
R11767 gnd.n1705 gnd.n1676 99.6594
R11768 gnd.n1707 gnd.n1677 99.6594
R11769 gnd.n1717 gnd.n1678 99.6594
R11770 gnd.n1728 gnd.n1679 99.6594
R11771 gnd.n1730 gnd.n1680 99.6594
R11772 gnd.n1740 gnd.n1681 99.6594
R11773 gnd.n1750 gnd.n1682 99.6594
R11774 gnd.n1752 gnd.n1683 99.6594
R11775 gnd.n5736 gnd.n1684 99.6594
R11776 gnd.n5738 gnd.n1685 99.6594
R11777 gnd.n5745 gnd.n1686 99.6594
R11778 gnd.n5747 gnd.n1687 99.6594
R11779 gnd.n5808 gnd.n1689 99.6594
R11780 gnd.n1706 gnd.n1676 99.6594
R11781 gnd.n1716 gnd.n1677 99.6594
R11782 gnd.n1727 gnd.n1678 99.6594
R11783 gnd.n1729 gnd.n1679 99.6594
R11784 gnd.n1739 gnd.n1680 99.6594
R11785 gnd.n1749 gnd.n1681 99.6594
R11786 gnd.n1751 gnd.n1682 99.6594
R11787 gnd.n5735 gnd.n1683 99.6594
R11788 gnd.n5737 gnd.n1684 99.6594
R11789 gnd.n5744 gnd.n1685 99.6594
R11790 gnd.n5746 gnd.n1686 99.6594
R11791 gnd.n1687 gnd.n1667 99.6594
R11792 gnd.n974 gnd.n796 99.6594
R11793 gnd.n976 gnd.n803 99.6594
R11794 gnd.n978 gnd.n977 99.6594
R11795 gnd.n979 gnd.n812 99.6594
R11796 gnd.n981 gnd.n819 99.6594
R11797 gnd.n983 gnd.n982 99.6594
R11798 gnd.n984 gnd.n828 99.6594
R11799 gnd.n1008 gnd.n986 99.6594
R11800 gnd.n1003 gnd.n987 99.6594
R11801 gnd.n1023 gnd.n988 99.6594
R11802 gnd.n999 gnd.n989 99.6594
R11803 gnd.n1032 gnd.n990 99.6594
R11804 gnd.n992 gnd.n991 99.6594
R11805 gnd.n1033 gnd.n991 99.6594
R11806 gnd.n1000 gnd.n990 99.6594
R11807 gnd.n1024 gnd.n989 99.6594
R11808 gnd.n1004 gnd.n988 99.6594
R11809 gnd.n1009 gnd.n987 99.6594
R11810 gnd.n986 gnd.n985 99.6594
R11811 gnd.n984 gnd.n827 99.6594
R11812 gnd.n983 gnd.n820 99.6594
R11813 gnd.n981 gnd.n980 99.6594
R11814 gnd.n979 gnd.n811 99.6594
R11815 gnd.n978 gnd.n804 99.6594
R11816 gnd.n976 gnd.n975 99.6594
R11817 gnd.n974 gnd.n795 99.6594
R11818 gnd.n1475 gnd.n1474 81.8399
R11819 gnd.n4397 gnd.t147 74.8376
R11820 gnd.n3649 gnd.t144 74.8376
R11821 gnd.n1476 gnd.n1469 72.8411
R11822 gnd.n1482 gnd.n1467 72.8411
R11823 gnd.n1130 gnd.n1129 72.8411
R11824 gnd.n6602 gnd.n6601 71.676
R11825 gnd.n6597 gnd.n1137 71.676
R11826 gnd.n6595 gnd.n6594 71.676
R11827 gnd.n6590 gnd.n1140 71.676
R11828 gnd.n6588 gnd.n6587 71.676
R11829 gnd.n6583 gnd.n1143 71.676
R11830 gnd.n6581 gnd.n6580 71.676
R11831 gnd.n6576 gnd.n1146 71.676
R11832 gnd.n6574 gnd.n6573 71.676
R11833 gnd.n6569 gnd.n1149 71.676
R11834 gnd.n6567 gnd.n6566 71.676
R11835 gnd.n6562 gnd.n1152 71.676
R11836 gnd.n6560 gnd.n6559 71.676
R11837 gnd.n6555 gnd.n1157 71.676
R11838 gnd.n6551 gnd.n6550 71.676
R11839 gnd.n6546 gnd.n1162 71.676
R11840 gnd.n6544 gnd.n6543 71.676
R11841 gnd.n6539 gnd.n1166 71.676
R11842 gnd.n6537 gnd.n6536 71.676
R11843 gnd.n6532 gnd.n1169 71.676
R11844 gnd.n6530 gnd.n6529 71.676
R11845 gnd.n6525 gnd.n1172 71.676
R11846 gnd.n6523 gnd.n6522 71.676
R11847 gnd.n6518 gnd.n1175 71.676
R11848 gnd.n6516 gnd.n6515 71.676
R11849 gnd.n6511 gnd.n1178 71.676
R11850 gnd.n6509 gnd.n6508 71.676
R11851 gnd.n6504 gnd.n1181 71.676
R11852 gnd.n6502 gnd.n6501 71.676
R11853 gnd.n6058 gnd.n6057 71.676
R11854 gnd.n6052 gnd.n1434 71.676
R11855 gnd.n6049 gnd.n1435 71.676
R11856 gnd.n6045 gnd.n1436 71.676
R11857 gnd.n6041 gnd.n1437 71.676
R11858 gnd.n6037 gnd.n1438 71.676
R11859 gnd.n6033 gnd.n1439 71.676
R11860 gnd.n6029 gnd.n1440 71.676
R11861 gnd.n6025 gnd.n1441 71.676
R11862 gnd.n6021 gnd.n1442 71.676
R11863 gnd.n6017 gnd.n1443 71.676
R11864 gnd.n6013 gnd.n1444 71.676
R11865 gnd.n6009 gnd.n1445 71.676
R11866 gnd.n6004 gnd.n1446 71.676
R11867 gnd.n6000 gnd.n1447 71.676
R11868 gnd.n1554 gnd.n1449 71.676
R11869 gnd.n1550 gnd.n1450 71.676
R11870 gnd.n1546 gnd.n1451 71.676
R11871 gnd.n1542 gnd.n1452 71.676
R11872 gnd.n1538 gnd.n1453 71.676
R11873 gnd.n1534 gnd.n1454 71.676
R11874 gnd.n1530 gnd.n1455 71.676
R11875 gnd.n1526 gnd.n1456 71.676
R11876 gnd.n1522 gnd.n1457 71.676
R11877 gnd.n1518 gnd.n1458 71.676
R11878 gnd.n1514 gnd.n1459 71.676
R11879 gnd.n1510 gnd.n1460 71.676
R11880 gnd.n1506 gnd.n1461 71.676
R11881 gnd.n1502 gnd.n1462 71.676
R11882 gnd.n6058 gnd.n1464 71.676
R11883 gnd.n6050 gnd.n1434 71.676
R11884 gnd.n6046 gnd.n1435 71.676
R11885 gnd.n6042 gnd.n1436 71.676
R11886 gnd.n6038 gnd.n1437 71.676
R11887 gnd.n6034 gnd.n1438 71.676
R11888 gnd.n6030 gnd.n1439 71.676
R11889 gnd.n6026 gnd.n1440 71.676
R11890 gnd.n6022 gnd.n1441 71.676
R11891 gnd.n6018 gnd.n1442 71.676
R11892 gnd.n6014 gnd.n1443 71.676
R11893 gnd.n6010 gnd.n1444 71.676
R11894 gnd.n6005 gnd.n1445 71.676
R11895 gnd.n6001 gnd.n1446 71.676
R11896 gnd.n1555 gnd.n1448 71.676
R11897 gnd.n1551 gnd.n1449 71.676
R11898 gnd.n1547 gnd.n1450 71.676
R11899 gnd.n1543 gnd.n1451 71.676
R11900 gnd.n1539 gnd.n1452 71.676
R11901 gnd.n1535 gnd.n1453 71.676
R11902 gnd.n1531 gnd.n1454 71.676
R11903 gnd.n1527 gnd.n1455 71.676
R11904 gnd.n1523 gnd.n1456 71.676
R11905 gnd.n1519 gnd.n1457 71.676
R11906 gnd.n1515 gnd.n1458 71.676
R11907 gnd.n1511 gnd.n1459 71.676
R11908 gnd.n1507 gnd.n1460 71.676
R11909 gnd.n1503 gnd.n1461 71.676
R11910 gnd.n1499 gnd.n1462 71.676
R11911 gnd.n6503 gnd.n6502 71.676
R11912 gnd.n1181 gnd.n1179 71.676
R11913 gnd.n6510 gnd.n6509 71.676
R11914 gnd.n1178 gnd.n1176 71.676
R11915 gnd.n6517 gnd.n6516 71.676
R11916 gnd.n1175 gnd.n1173 71.676
R11917 gnd.n6524 gnd.n6523 71.676
R11918 gnd.n1172 gnd.n1170 71.676
R11919 gnd.n6531 gnd.n6530 71.676
R11920 gnd.n1169 gnd.n1167 71.676
R11921 gnd.n6538 gnd.n6537 71.676
R11922 gnd.n1166 gnd.n1164 71.676
R11923 gnd.n6545 gnd.n6544 71.676
R11924 gnd.n1162 gnd.n1158 71.676
R11925 gnd.n6554 gnd.n6553 71.676
R11926 gnd.n1157 gnd.n1153 71.676
R11927 gnd.n6561 gnd.n6560 71.676
R11928 gnd.n1152 gnd.n1150 71.676
R11929 gnd.n6568 gnd.n6567 71.676
R11930 gnd.n1149 gnd.n1147 71.676
R11931 gnd.n6575 gnd.n6574 71.676
R11932 gnd.n1146 gnd.n1144 71.676
R11933 gnd.n6582 gnd.n6581 71.676
R11934 gnd.n1143 gnd.n1141 71.676
R11935 gnd.n6589 gnd.n6588 71.676
R11936 gnd.n1140 gnd.n1138 71.676
R11937 gnd.n6596 gnd.n6595 71.676
R11938 gnd.n1137 gnd.n1135 71.676
R11939 gnd.n6603 gnd.n6602 71.676
R11940 gnd.n4034 gnd.n3935 67.3134
R11941 gnd.n5117 gnd.n5116 59.9823
R11942 gnd.n1492 gnd.n1491 59.5399
R11943 gnd.n1161 gnd.n1160 59.5399
R11944 gnd.n6007 gnd.n1489 59.5399
R11945 gnd.n1156 gnd.n1155 59.5399
R11946 gnd.n1487 gnd.n1485 59.1804
R11947 gnd.n4298 gnd.n4297 56.1363
R11948 gnd.n4300 gnd.n4299 56.1363
R11949 gnd.n4302 gnd.n4301 56.1363
R11950 gnd.n4159 gnd.n4158 56.1363
R11951 gnd.n4161 gnd.n4160 56.1363
R11952 gnd.n4163 gnd.n4162 56.1363
R11953 gnd.n4228 gnd.n4227 56.1363
R11954 gnd.n4230 gnd.n4229 56.1363
R11955 gnd.n4232 gnd.n4231 56.1363
R11956 gnd.n431 gnd.n430 56.1363
R11957 gnd.n429 gnd.n428 56.1363
R11958 gnd.n427 gnd.n426 56.1363
R11959 gnd.n292 gnd.n291 56.1363
R11960 gnd.n290 gnd.n289 56.1363
R11961 gnd.n288 gnd.n287 56.1363
R11962 gnd.n361 gnd.n360 56.1363
R11963 gnd.n359 gnd.n358 56.1363
R11964 gnd.n357 gnd.n356 56.1363
R11965 gnd.n5281 gnd.n2012 55.3171
R11966 gnd.n7353 gnd.n502 55.3171
R11967 gnd.n1473 gnd.n1472 54.358
R11968 gnd.n1127 gnd.n1126 54.358
R11969 gnd.n1118 gnd.n1117 52.4801
R11970 gnd.n4276 gnd.t97 52.3082
R11971 gnd.n4313 gnd.t95 52.3082
R11972 gnd.n4137 gnd.t55 52.3082
R11973 gnd.n4174 gnd.t76 52.3082
R11974 gnd.n4206 gnd.t107 52.3082
R11975 gnd.n4243 gnd.t66 52.3082
R11976 gnd.n442 gnd.t96 52.3082
R11977 gnd.n405 gnd.t99 52.3082
R11978 gnd.n303 gnd.t100 52.3082
R11979 gnd.n266 gnd.t79 52.3082
R11980 gnd.n372 gnd.t88 52.3082
R11981 gnd.n335 gnd.t69 52.3082
R11982 gnd.n4979 gnd.t36 52.3082
R11983 gnd.n4947 gnd.t34 52.3082
R11984 gnd.n4915 gnd.t32 52.3082
R11985 gnd.n4884 gnd.t30 52.3082
R11986 gnd.n4852 gnd.t28 52.3082
R11987 gnd.n4820 gnd.t40 52.3082
R11988 gnd.n4788 gnd.t44 52.3082
R11989 gnd.n4757 gnd.t42 52.3082
R11990 gnd.n106 gnd.t5 52.3082
R11991 gnd.n74 gnd.t38 52.3082
R11992 gnd.n42 gnd.t7 52.3082
R11993 gnd.n11 gnd.t1 52.3082
R11994 gnd.n233 gnd.t219 52.3082
R11995 gnd.n201 gnd.t26 52.3082
R11996 gnd.n169 gnd.t14 52.3082
R11997 gnd.n138 gnd.t3 52.3082
R11998 gnd.n4809 gnd.n4777 51.4173
R11999 gnd.n190 gnd.n158 51.4173
R12000 gnd.n4873 gnd.n4872 50.455
R12001 gnd.n4841 gnd.n4840 50.455
R12002 gnd.n4809 gnd.n4808 50.455
R12003 gnd.n254 gnd.n253 50.455
R12004 gnd.n222 gnd.n221 50.455
R12005 gnd.n190 gnd.n189 50.455
R12006 gnd.n5742 gnd.n5741 45.1884
R12007 gnd.n3972 gnd.n3971 45.1884
R12008 gnd.n3675 gnd.n3674 45.1884
R12009 gnd.n7236 gnd.n7235 45.1884
R12010 gnd.n6969 gnd.n6968 45.1884
R12011 gnd.n1744 gnd.n1743 45.1884
R12012 gnd.n881 gnd.n880 45.1884
R12013 gnd.n901 gnd.n900 45.1884
R12014 gnd.n572 gnd.n571 45.1884
R12015 gnd.n536 gnd.n535 45.1884
R12016 gnd.n2123 gnd.n2122 45.1884
R12017 gnd.n2052 gnd.n2051 45.1884
R12018 gnd.n5244 gnd.n5243 45.1884
R12019 gnd.n1595 gnd.n1594 45.1884
R12020 gnd.n1560 gnd.n1559 45.1884
R12021 gnd.n997 gnd.n996 45.1884
R12022 gnd.n6606 gnd.n1133 44.3322
R12023 gnd.n1476 gnd.n1475 44.3189
R12024 gnd.n5743 gnd.n5742 42.2793
R12025 gnd.n3984 gnd.n3972 42.2793
R12026 gnd.n3676 gnd.n3675 42.2793
R12027 gnd.n4399 gnd.n4397 42.2793
R12028 gnd.n5088 gnd.n3649 42.2793
R12029 gnd.n7239 gnd.n7236 42.2793
R12030 gnd.n6970 gnd.n6969 42.2793
R12031 gnd.n5770 gnd.n1744 42.2793
R12032 gnd.n902 gnd.n901 42.2793
R12033 gnd.n7291 gnd.n572 42.2793
R12034 gnd.n537 gnd.n536 42.2793
R12035 gnd.n2124 gnd.n2123 42.2793
R12036 gnd.n2053 gnd.n2052 42.2793
R12037 gnd.n5245 gnd.n5244 42.2793
R12038 gnd.n5964 gnd.n1595 42.2793
R12039 gnd.n1030 gnd.n997 42.2793
R12040 gnd.n1474 gnd.n1473 41.6274
R12041 gnd.n1128 gnd.n1127 41.6274
R12042 gnd.n3375 gnd.n2318 41.2608
R12043 gnd.n3383 gnd.n2318 41.2608
R12044 gnd.n3384 gnd.n3383 41.2608
R12045 gnd.n3385 gnd.n3384 41.2608
R12046 gnd.n3385 gnd.n2312 41.2608
R12047 gnd.n3393 gnd.n2312 41.2608
R12048 gnd.n3394 gnd.n3393 41.2608
R12049 gnd.n3395 gnd.n3394 41.2608
R12050 gnd.n3395 gnd.n2306 41.2608
R12051 gnd.n3403 gnd.n2306 41.2608
R12052 gnd.n3404 gnd.n3403 41.2608
R12053 gnd.n3405 gnd.n3404 41.2608
R12054 gnd.n3405 gnd.n2300 41.2608
R12055 gnd.n3413 gnd.n2300 41.2608
R12056 gnd.n3414 gnd.n3413 41.2608
R12057 gnd.n3415 gnd.n3414 41.2608
R12058 gnd.n3415 gnd.n2294 41.2608
R12059 gnd.n3423 gnd.n2294 41.2608
R12060 gnd.n3424 gnd.n3423 41.2608
R12061 gnd.n3425 gnd.n3424 41.2608
R12062 gnd.n3425 gnd.n2288 41.2608
R12063 gnd.n3433 gnd.n2288 41.2608
R12064 gnd.n3434 gnd.n3433 41.2608
R12065 gnd.n3435 gnd.n3434 41.2608
R12066 gnd.n3435 gnd.n2282 41.2608
R12067 gnd.n3443 gnd.n2282 41.2608
R12068 gnd.n3444 gnd.n3443 41.2608
R12069 gnd.n3445 gnd.n3444 41.2608
R12070 gnd.n3445 gnd.n2276 41.2608
R12071 gnd.n3453 gnd.n2276 41.2608
R12072 gnd.n3454 gnd.n3453 41.2608
R12073 gnd.n3455 gnd.n3454 41.2608
R12074 gnd.n3455 gnd.n2270 41.2608
R12075 gnd.n3463 gnd.n2270 41.2608
R12076 gnd.n3464 gnd.n3463 41.2608
R12077 gnd.n3465 gnd.n3464 41.2608
R12078 gnd.n3465 gnd.n2264 41.2608
R12079 gnd.n3473 gnd.n2264 41.2608
R12080 gnd.n3474 gnd.n3473 41.2608
R12081 gnd.n3475 gnd.n3474 41.2608
R12082 gnd.n3475 gnd.n2258 41.2608
R12083 gnd.n3483 gnd.n2258 41.2608
R12084 gnd.n3484 gnd.n3483 41.2608
R12085 gnd.n3485 gnd.n3484 41.2608
R12086 gnd.n3485 gnd.n2252 41.2608
R12087 gnd.n3493 gnd.n2252 41.2608
R12088 gnd.n3494 gnd.n3493 41.2608
R12089 gnd.n3495 gnd.n3494 41.2608
R12090 gnd.n3495 gnd.n2246 41.2608
R12091 gnd.n3503 gnd.n2246 41.2608
R12092 gnd.n3504 gnd.n3503 41.2608
R12093 gnd.n3505 gnd.n3504 41.2608
R12094 gnd.n3505 gnd.n2240 41.2608
R12095 gnd.n3513 gnd.n2240 41.2608
R12096 gnd.n3514 gnd.n3513 41.2608
R12097 gnd.n3515 gnd.n3514 41.2608
R12098 gnd.n3515 gnd.n2234 41.2608
R12099 gnd.n3523 gnd.n2234 41.2608
R12100 gnd.n3524 gnd.n3523 41.2608
R12101 gnd.n3525 gnd.n3524 41.2608
R12102 gnd.n3525 gnd.n2228 41.2608
R12103 gnd.n3533 gnd.n2228 41.2608
R12104 gnd.n3534 gnd.n3533 41.2608
R12105 gnd.n5161 gnd.n3534 41.2608
R12106 gnd.n5161 gnd.n5160 41.2608
R12107 gnd.n1483 gnd.n1482 40.8975
R12108 gnd.n1131 gnd.n1130 40.8975
R12109 gnd.n4298 gnd.n4296 39.1642
R12110 gnd.n427 gnd.n425 39.1642
R12111 gnd.n4159 gnd.n4157 38.8139
R12112 gnd.n4228 gnd.n4226 38.8139
R12113 gnd.n288 gnd.n286 38.8139
R12114 gnd.n357 gnd.n355 38.8139
R12115 gnd.n4334 gnd.n4333 37.8096
R12116 gnd.n4195 gnd.n4194 37.8096
R12117 gnd.n4264 gnd.n4263 37.8096
R12118 gnd.n463 gnd.n462 37.8096
R12119 gnd.n324 gnd.n323 37.8096
R12120 gnd.n393 gnd.n392 37.8096
R12121 gnd.n6937 gnd.n881 36.9518
R12122 gnd.n5997 gnd.n1560 36.9518
R12123 gnd.n1482 gnd.n1481 35.055
R12124 gnd.n1477 gnd.n1476 35.055
R12125 gnd.n1120 gnd.n1119 35.055
R12126 gnd.n1130 gnd.n1116 35.055
R12127 gnd.n6500 gnd.n6499 33.8737
R12128 gnd.n1500 gnd.n1493 33.8737
R12129 gnd.n4034 gnd.n3930 33.3237
R12130 gnd.n4042 gnd.n3930 33.3237
R12131 gnd.n4050 gnd.n3924 33.3237
R12132 gnd.n4050 gnd.n3918 33.3237
R12133 gnd.n4058 gnd.n3918 33.3237
R12134 gnd.n4058 gnd.n3911 33.3237
R12135 gnd.n4066 gnd.n3911 33.3237
R12136 gnd.n4066 gnd.n3912 33.3237
R12137 gnd.n4440 gnd.n3897 33.3237
R12138 gnd.n5281 gnd.n2005 33.3237
R12139 gnd.n5289 gnd.n2005 33.3237
R12140 gnd.n5297 gnd.n1996 33.3237
R12141 gnd.n5305 gnd.n1987 33.3237
R12142 gnd.n5550 gnd.n1603 33.3237
R12143 gnd.n5545 gnd.n5544 33.3237
R12144 gnd.n5545 gnd.n1675 33.3237
R12145 gnd.n5810 gnd.n1668 33.3237
R12146 gnd.n6686 gnd.n973 33.3237
R12147 gnd.n6713 gnd.n6712 33.3237
R12148 gnd.n6713 gnd.n833 33.3237
R12149 gnd.n861 gnd.n786 33.3237
R12150 gnd.n7199 gnd.n596 33.3237
R12151 gnd.n7275 gnd.n585 33.3237
R12152 gnd.n7283 gnd.n500 33.3237
R12153 gnd.n7353 gnd.n500 33.3237
R12154 gnd.n5227 gnd.n1990 31.9908
R12155 gnd.n5313 gnd.n1978 31.9908
R12156 gnd.n5221 gnd.n1981 31.9908
R12157 gnd.n2212 gnd.n1972 31.9908
R12158 gnd.n5338 gnd.n1960 31.9908
R12159 gnd.n2206 gnd.n1963 31.9908
R12160 gnd.n5348 gnd.n1950 31.9908
R12161 gnd.n5362 gnd.n1944 31.9908
R12162 gnd.n5379 gnd.n1921 31.9908
R12163 gnd.n5356 gnd.n1924 31.9908
R12164 gnd.n5373 gnd.n1938 31.9908
R12165 gnd.n5388 gnd.n1910 31.9908
R12166 gnd.n1934 gnd.n1912 31.9908
R12167 gnd.n5397 gnd.n1904 31.9908
R12168 gnd.n5643 gnd.n1847 31.9908
R12169 gnd.n5637 gnd.n1859 31.9908
R12170 gnd.n5632 gnd.n1862 31.9908
R12171 gnd.n5631 gnd.n1868 31.9908
R12172 gnd.n1875 gnd.n1874 31.9908
R12173 gnd.n5618 gnd.n1878 31.9908
R12174 gnd.n5596 gnd.n1884 31.9908
R12175 gnd.n5652 gnd.n1832 31.9908
R12176 gnd.n5660 gnd.n1823 31.9908
R12177 gnd.n5484 gnd.n1826 31.9908
R12178 gnd.n5668 gnd.n1814 31.9908
R12179 gnd.n5511 gnd.n1817 31.9908
R12180 gnd.n5505 gnd.n1808 31.9908
R12181 gnd.n5684 gnd.n1797 31.9908
R12182 gnd.n5501 gnd.n1800 31.9908
R12183 gnd.n5692 gnd.n1788 31.9908
R12184 gnd.n5700 gnd.n1779 31.9908
R12185 gnd.n5569 gnd.n1782 31.9908
R12186 gnd.n5713 gnd.n1769 31.9908
R12187 gnd.n5563 gnd.n1772 31.9908
R12188 gnd.n5721 gnd.n1760 31.9908
R12189 gnd.n5559 gnd.n1762 31.9908
R12190 gnd.n5728 gnd.n1613 31.9908
R12191 gnd.n5958 gnd.n1601 31.9908
R12192 gnd.n7015 gnd.n789 31.9908
R12193 gnd.n1013 gnd.n779 31.9908
R12194 gnd.n6892 gnd.n770 31.9908
R12195 gnd.n7031 gnd.n773 31.9908
R12196 gnd.n6758 gnd.n761 31.9908
R12197 gnd.n7039 gnd.n764 31.9908
R12198 gnd.n6764 gnd.n752 31.9908
R12199 gnd.n7047 gnd.n755 31.9908
R12200 gnd.n7055 gnd.n746 31.9908
R12201 gnd.n6774 gnd.n734 31.9908
R12202 gnd.n7063 gnd.n737 31.9908
R12203 gnd.n6778 gnd.n726 31.9908
R12204 gnd.n6811 gnd.n717 31.9908
R12205 gnd.n7079 gnd.n720 31.9908
R12206 gnd.n6805 gnd.n708 31.9908
R12207 gnd.n7088 gnd.n711 31.9908
R12208 gnd.n7096 gnd.n702 31.9908
R12209 gnd.n6797 gnd.n691 31.9908
R12210 gnd.n7104 gnd.n694 31.9908
R12211 gnd.n7112 gnd.n685 31.9908
R12212 gnd.n6854 gnd.n675 31.9908
R12213 gnd.n7120 gnd.n678 31.9908
R12214 gnd.n6848 gnd.n667 31.9908
R12215 gnd.n6844 gnd.n660 31.9908
R12216 gnd.n7135 gnd.n663 31.9908
R12217 gnd.n2840 gnd.n652 31.9908
R12218 gnd.n7143 gnd.n654 31.9908
R12219 gnd.n2844 gnd.n643 31.9908
R12220 gnd.n7151 gnd.n646 31.9908
R12221 gnd.n2850 gnd.n635 31.9908
R12222 gnd.n7159 gnd.n637 31.9908
R12223 gnd.n7167 gnd.n629 31.9908
R12224 gnd.n2860 gnd.n618 31.9908
R12225 gnd.n7175 gnd.n620 31.9908
R12226 gnd.n2864 gnd.n610 31.9908
R12227 gnd.n2888 gnd.n602 31.9908
R12228 gnd.n7191 gnd.n604 31.9908
R12229 gnd.n2882 gnd.n593 31.9908
R12230 gnd.t77 gnd.n1835 31.6576
R12231 gnd.t47 gnd.n699 31.6576
R12232 gnd.n5289 gnd.t124 28.3253
R12233 gnd.n5904 gnd.t132 28.3253
R12234 gnd.n7023 gnd.t110 28.3253
R12235 gnd.n7283 gnd.t160 28.3253
R12236 gnd.n4441 gnd.n3887 25.9926
R12237 gnd.n3890 gnd.n3880 25.9926
R12238 gnd.n4471 gnd.n3873 25.9926
R12239 gnd.n4472 gnd.n3862 25.9926
R12240 gnd.n3865 gnd.n3853 25.9926
R12241 gnd.n4493 gnd.n3854 25.9926
R12242 gnd.n4514 gnd.n4513 25.9926
R12243 gnd.n3839 gnd.n3827 25.9926
R12244 gnd.n4524 gnd.n3828 25.9926
R12245 gnd.n4534 gnd.n3810 25.9926
R12246 gnd.n4545 gnd.n4544 25.9926
R12247 gnd.n4555 gnd.n3803 25.9926
R12248 gnd.n4564 gnd.n3795 25.9926
R12249 gnd.n4565 gnd.n3784 25.9926
R12250 gnd.n4576 gnd.n4575 25.9926
R12251 gnd.n4595 gnd.n3770 25.9926
R12252 gnd.n4607 gnd.n4606 25.9926
R12253 gnd.n4106 gnd.n3762 25.9926
R12254 gnd.n4617 gnd.n3752 25.9926
R12255 gnd.n4626 gnd.n3745 25.9926
R12256 gnd.n4637 gnd.n4636 25.9926
R12257 gnd.n3735 gnd.n3726 25.9926
R12258 gnd.n3717 gnd.n3710 25.9926
R12259 gnd.n4679 gnd.n4678 25.9926
R12260 gnd.n4694 gnd.n3701 25.9926
R12261 gnd.n4693 gnd.n3703 25.9926
R12262 gnd.n4669 gnd.n3537 25.9926
R12263 gnd.n5152 gnd.n3546 25.9926
R12264 gnd.n4715 gnd.n3557 25.9926
R12265 gnd.n4738 gnd.n4737 25.9926
R12266 gnd.n5138 gnd.n3568 25.9926
R12267 gnd.n4730 gnd.n3581 25.9926
R12268 gnd.n5131 gnd.n5130 25.9926
R12269 gnd.n5023 gnd.n3584 25.9926
R12270 gnd.n5016 gnd.n3604 25.9926
R12271 gnd.n1491 gnd.n1490 25.7944
R12272 gnd.n1160 gnd.n1159 25.7944
R12273 gnd.n1489 gnd.n1488 25.7944
R12274 gnd.n1155 gnd.n1154 25.7944
R12275 gnd.n4397 gnd.n4396 25.7944
R12276 gnd.n3649 gnd.n3648 25.7944
R12277 gnd.n5160 gnd.n5159 24.7567
R12278 gnd.n4462 gnd.t41 24.3265
R12279 gnd.n4452 gnd.t146 23.66
R12280 gnd.n5497 gnd.t54 22.9935
R12281 gnd.n6768 gnd.t68 22.9935
R12282 gnd.n4431 gnd.t29 22.3271
R12283 gnd.t60 gnd.n5623 22.3271
R12284 gnd.n6793 gnd.t51 22.3271
R12285 gnd.n4716 gnd.t20 21.6606
R12286 gnd.n5220 gnd.t65 21.6606
R12287 gnd.n5331 gnd.t56 21.6606
R12288 gnd.n2854 gnd.t62 21.6606
R12289 gnd.n2889 gnd.t87 21.6606
R12290 gnd.n1487 gnd.n1486 21.0737
R12291 gnd.n6607 gnd.n6606 21.0737
R12292 gnd.n4657 gnd.t221 20.9941
R12293 gnd.n1999 gnd.n1987 20.9941
R12294 gnd.t45 gnd.n1850 20.9941
R12295 gnd.n6843 gnd.t74 20.9941
R12296 gnd.n596 gnd.n583 20.9941
R12297 gnd.n5550 gnd.n1567 20.6609
R12298 gnd.n6964 gnd.n861 20.6609
R12299 gnd.t226 gnd.n3759 20.3277
R12300 gnd.n5512 gnd.t58 20.3277
R12301 gnd.n6812 gnd.t49 20.3277
R12302 gnd.n1470 gnd.t216 19.8005
R12303 gnd.n1470 gnd.t118 19.8005
R12304 gnd.n1471 gnd.t192 19.8005
R12305 gnd.n1471 gnd.t168 19.8005
R12306 gnd.n1124 gnd.t177 19.8005
R12307 gnd.n1124 gnd.t195 19.8005
R12308 gnd.n1125 gnd.t140 19.8005
R12309 gnd.n1125 gnd.t115 19.8005
R12310 gnd.t9 gnd.n3802 19.6612
R12311 gnd.n4586 gnd.t33 19.6612
R12312 gnd.n1467 gnd.n1466 19.5087
R12313 gnd.n1480 gnd.n1467 19.5087
R12314 gnd.n1478 gnd.n1469 19.5087
R12315 gnd.n1129 gnd.n1123 19.5087
R12316 gnd.n5821 gnd.n1665 19.3944
R12317 gnd.n5825 gnd.n1665 19.3944
R12318 gnd.n5825 gnd.n1654 19.3944
R12319 gnd.n5841 gnd.n1654 19.3944
R12320 gnd.n5841 gnd.n1652 19.3944
R12321 gnd.n5845 gnd.n1652 19.3944
R12322 gnd.n5845 gnd.n1640 19.3944
R12323 gnd.n5863 gnd.n1640 19.3944
R12324 gnd.n5863 gnd.n1637 19.3944
R12325 gnd.n5872 gnd.n1637 19.3944
R12326 gnd.n5872 gnd.n1638 19.3944
R12327 gnd.n5868 gnd.n1638 19.3944
R12328 gnd.n5868 gnd.n5867 19.3944
R12329 gnd.n5867 gnd.n1413 19.3944
R12330 gnd.n6083 gnd.n1413 19.3944
R12331 gnd.n6083 gnd.n1410 19.3944
R12332 gnd.n6121 gnd.n1410 19.3944
R12333 gnd.n6121 gnd.n1411 19.3944
R12334 gnd.n6117 gnd.n1411 19.3944
R12335 gnd.n6117 gnd.n6116 19.3944
R12336 gnd.n6116 gnd.n6115 19.3944
R12337 gnd.n6115 gnd.n6089 19.3944
R12338 gnd.n6111 gnd.n6089 19.3944
R12339 gnd.n6111 gnd.n6110 19.3944
R12340 gnd.n6110 gnd.n6109 19.3944
R12341 gnd.n6109 gnd.n1336 19.3944
R12342 gnd.n6230 gnd.n1336 19.3944
R12343 gnd.n6230 gnd.n1333 19.3944
R12344 gnd.n6247 gnd.n1333 19.3944
R12345 gnd.n6247 gnd.n1334 19.3944
R12346 gnd.n6243 gnd.n1334 19.3944
R12347 gnd.n6243 gnd.n6242 19.3944
R12348 gnd.n6242 gnd.n6241 19.3944
R12349 gnd.n6241 gnd.n6237 19.3944
R12350 gnd.n6237 gnd.n1277 19.3944
R12351 gnd.n6342 gnd.n1277 19.3944
R12352 gnd.n6343 gnd.n6342 19.3944
R12353 gnd.n6343 gnd.n1274 19.3944
R12354 gnd.n6380 gnd.n1274 19.3944
R12355 gnd.n6380 gnd.n1275 19.3944
R12356 gnd.n6376 gnd.n1275 19.3944
R12357 gnd.n6376 gnd.n6375 19.3944
R12358 gnd.n6375 gnd.n6374 19.3944
R12359 gnd.n6374 gnd.n6348 19.3944
R12360 gnd.n6370 gnd.n6348 19.3944
R12361 gnd.n6370 gnd.n6369 19.3944
R12362 gnd.n6369 gnd.n6368 19.3944
R12363 gnd.n6368 gnd.n6352 19.3944
R12364 gnd.n6364 gnd.n6352 19.3944
R12365 gnd.n6364 gnd.n6363 19.3944
R12366 gnd.n6363 gnd.n6362 19.3944
R12367 gnd.n6362 gnd.n6359 19.3944
R12368 gnd.n6359 gnd.n1088 19.3944
R12369 gnd.n6633 gnd.n1088 19.3944
R12370 gnd.n6633 gnd.n1085 19.3944
R12371 gnd.n6638 gnd.n1085 19.3944
R12372 gnd.n6638 gnd.n1086 19.3944
R12373 gnd.n1086 gnd.n1063 19.3944
R12374 gnd.n6663 gnd.n1063 19.3944
R12375 gnd.n6663 gnd.n1060 19.3944
R12376 gnd.n6669 gnd.n1060 19.3944
R12377 gnd.n6669 gnd.n1061 19.3944
R12378 gnd.n1061 gnd.n1038 19.3944
R12379 gnd.n6705 gnd.n1038 19.3944
R12380 gnd.n6706 gnd.n6705 19.3944
R12381 gnd.n5752 gnd.n5751 19.3944
R12382 gnd.n5751 gnd.n5750 19.3944
R12383 gnd.n5750 gnd.n5748 19.3944
R12384 gnd.n5806 gnd.n5805 19.3944
R12385 gnd.n5805 gnd.n1691 19.3944
R12386 gnd.n5798 gnd.n1691 19.3944
R12387 gnd.n5798 gnd.n5797 19.3944
R12388 gnd.n5797 gnd.n1708 19.3944
R12389 gnd.n5790 gnd.n1708 19.3944
R12390 gnd.n5790 gnd.n5789 19.3944
R12391 gnd.n5789 gnd.n1718 19.3944
R12392 gnd.n5782 gnd.n1718 19.3944
R12393 gnd.n5782 gnd.n5781 19.3944
R12394 gnd.n5781 gnd.n1731 19.3944
R12395 gnd.n5774 gnd.n1731 19.3944
R12396 gnd.n5774 gnd.n5773 19.3944
R12397 gnd.n5773 gnd.n1741 19.3944
R12398 gnd.n5764 gnd.n1741 19.3944
R12399 gnd.n5764 gnd.n5763 19.3944
R12400 gnd.n5763 gnd.n5762 19.3944
R12401 gnd.n5762 gnd.n1753 19.3944
R12402 gnd.n5758 gnd.n1753 19.3944
R12403 gnd.n5758 gnd.n5757 19.3944
R12404 gnd.n5757 gnd.n5756 19.3944
R12405 gnd.n5756 gnd.n5739 19.3944
R12406 gnd.n4029 gnd.n4028 19.3944
R12407 gnd.n4028 gnd.n3938 19.3944
R12408 gnd.n4023 gnd.n3938 19.3944
R12409 gnd.n4023 gnd.n4022 19.3944
R12410 gnd.n4022 gnd.n3943 19.3944
R12411 gnd.n4017 gnd.n3943 19.3944
R12412 gnd.n4017 gnd.n4016 19.3944
R12413 gnd.n4016 gnd.n4015 19.3944
R12414 gnd.n4015 gnd.n3949 19.3944
R12415 gnd.n4009 gnd.n3949 19.3944
R12416 gnd.n4009 gnd.n4008 19.3944
R12417 gnd.n4008 gnd.n4007 19.3944
R12418 gnd.n4007 gnd.n3955 19.3944
R12419 gnd.n4001 gnd.n3955 19.3944
R12420 gnd.n4001 gnd.n4000 19.3944
R12421 gnd.n4000 gnd.n3999 19.3944
R12422 gnd.n3999 gnd.n3961 19.3944
R12423 gnd.n3993 gnd.n3961 19.3944
R12424 gnd.n3993 gnd.n3992 19.3944
R12425 gnd.n3992 gnd.n3991 19.3944
R12426 gnd.n3991 gnd.n3967 19.3944
R12427 gnd.n3985 gnd.n3967 19.3944
R12428 gnd.n3983 gnd.n3982 19.3944
R12429 gnd.n3982 gnd.n3977 19.3944
R12430 gnd.n3977 gnd.n3975 19.3944
R12431 gnd.n5038 gnd.n5037 19.3944
R12432 gnd.n5037 gnd.n5034 19.3944
R12433 gnd.n5034 gnd.n5033 19.3944
R12434 gnd.n5083 gnd.n5082 19.3944
R12435 gnd.n5082 gnd.n5081 19.3944
R12436 gnd.n5081 gnd.n5078 19.3944
R12437 gnd.n5078 gnd.n5077 19.3944
R12438 gnd.n5077 gnd.n5074 19.3944
R12439 gnd.n5074 gnd.n5073 19.3944
R12440 gnd.n5073 gnd.n5070 19.3944
R12441 gnd.n5070 gnd.n5069 19.3944
R12442 gnd.n5069 gnd.n5066 19.3944
R12443 gnd.n5066 gnd.n5065 19.3944
R12444 gnd.n5065 gnd.n5062 19.3944
R12445 gnd.n5062 gnd.n5061 19.3944
R12446 gnd.n5061 gnd.n5058 19.3944
R12447 gnd.n5058 gnd.n5057 19.3944
R12448 gnd.n5057 gnd.n5054 19.3944
R12449 gnd.n5054 gnd.n5053 19.3944
R12450 gnd.n5053 gnd.n5050 19.3944
R12451 gnd.n5050 gnd.n5049 19.3944
R12452 gnd.n5049 gnd.n5046 19.3944
R12453 gnd.n5046 gnd.n5045 19.3944
R12454 gnd.n5045 gnd.n5042 19.3944
R12455 gnd.n5042 gnd.n5041 19.3944
R12456 gnd.n4444 gnd.n4443 19.3944
R12457 gnd.n4444 gnd.n3878 19.3944
R12458 gnd.n4464 gnd.n3878 19.3944
R12459 gnd.n4464 gnd.n3870 19.3944
R12460 gnd.n4474 gnd.n3870 19.3944
R12461 gnd.n4475 gnd.n4474 19.3944
R12462 gnd.n4475 gnd.n3851 19.3944
R12463 gnd.n4495 gnd.n3851 19.3944
R12464 gnd.n4495 gnd.n3844 19.3944
R12465 gnd.n4505 gnd.n3844 19.3944
R12466 gnd.n4506 gnd.n4505 19.3944
R12467 gnd.n4506 gnd.n3825 19.3944
R12468 gnd.n4526 gnd.n3825 19.3944
R12469 gnd.n4526 gnd.n3818 19.3944
R12470 gnd.n4536 gnd.n3818 19.3944
R12471 gnd.n4537 gnd.n4536 19.3944
R12472 gnd.n4537 gnd.n3800 19.3944
R12473 gnd.n4557 gnd.n3800 19.3944
R12474 gnd.n4557 gnd.n3792 19.3944
R12475 gnd.n4567 gnd.n3792 19.3944
R12476 gnd.n4568 gnd.n4567 19.3944
R12477 gnd.n4568 gnd.n3775 19.3944
R12478 gnd.n4588 gnd.n3775 19.3944
R12479 gnd.n4588 gnd.n3767 19.3944
R12480 gnd.n4598 gnd.n3767 19.3944
R12481 gnd.n4599 gnd.n4598 19.3944
R12482 gnd.n4599 gnd.n3750 19.3944
R12483 gnd.n4619 gnd.n3750 19.3944
R12484 gnd.n4619 gnd.n3741 19.3944
R12485 gnd.n4629 gnd.n3741 19.3944
R12486 gnd.n4630 gnd.n4629 19.3944
R12487 gnd.n4631 gnd.n4630 19.3944
R12488 gnd.n4631 gnd.n3724 19.3944
R12489 gnd.n4648 gnd.n3724 19.3944
R12490 gnd.n4651 gnd.n4648 19.3944
R12491 gnd.n4651 gnd.n4650 19.3944
R12492 gnd.n4650 gnd.n3697 19.3944
R12493 gnd.n4701 gnd.n3697 19.3944
R12494 gnd.n4701 gnd.n3694 19.3944
R12495 gnd.n4705 gnd.n3694 19.3944
R12496 gnd.n4706 gnd.n4705 19.3944
R12497 gnd.n4713 gnd.n4706 19.3944
R12498 gnd.n4713 gnd.n4712 19.3944
R12499 gnd.n4712 gnd.n3688 19.3944
R12500 gnd.n4741 gnd.n3688 19.3944
R12501 gnd.n4742 gnd.n4741 19.3944
R12502 gnd.n4742 gnd.n3686 19.3944
R12503 gnd.n5004 gnd.n3686 19.3944
R12504 gnd.n5006 gnd.n5004 19.3944
R12505 gnd.n5020 gnd.n5006 19.3944
R12506 gnd.n5020 gnd.n5019 19.3944
R12507 gnd.n5019 gnd.n5018 19.3944
R12508 gnd.n5018 gnd.n5014 19.3944
R12509 gnd.n4427 gnd.n4426 19.3944
R12510 gnd.n4426 gnd.n4425 19.3944
R12511 gnd.n4425 gnd.n4424 19.3944
R12512 gnd.n4424 gnd.n4422 19.3944
R12513 gnd.n4422 gnd.n4419 19.3944
R12514 gnd.n4419 gnd.n4418 19.3944
R12515 gnd.n4418 gnd.n4415 19.3944
R12516 gnd.n4415 gnd.n4414 19.3944
R12517 gnd.n4414 gnd.n4411 19.3944
R12518 gnd.n4411 gnd.n4410 19.3944
R12519 gnd.n4410 gnd.n4407 19.3944
R12520 gnd.n4407 gnd.n4406 19.3944
R12521 gnd.n4406 gnd.n4403 19.3944
R12522 gnd.n4403 gnd.n4402 19.3944
R12523 gnd.n4454 gnd.n3885 19.3944
R12524 gnd.n4454 gnd.n3883 19.3944
R12525 gnd.n4460 gnd.n3883 19.3944
R12526 gnd.n4460 gnd.n4459 19.3944
R12527 gnd.n4459 gnd.n3860 19.3944
R12528 gnd.n4485 gnd.n3860 19.3944
R12529 gnd.n4485 gnd.n3858 19.3944
R12530 gnd.n4491 gnd.n3858 19.3944
R12531 gnd.n4491 gnd.n4490 19.3944
R12532 gnd.n4490 gnd.n3834 19.3944
R12533 gnd.n4516 gnd.n3834 19.3944
R12534 gnd.n4516 gnd.n3832 19.3944
R12535 gnd.n4522 gnd.n3832 19.3944
R12536 gnd.n4522 gnd.n4521 19.3944
R12537 gnd.n4521 gnd.n3808 19.3944
R12538 gnd.n4547 gnd.n3808 19.3944
R12539 gnd.n4547 gnd.n3806 19.3944
R12540 gnd.n4553 gnd.n3806 19.3944
R12541 gnd.n4553 gnd.n4552 19.3944
R12542 gnd.n4552 gnd.n3782 19.3944
R12543 gnd.n4578 gnd.n3782 19.3944
R12544 gnd.n4578 gnd.n3780 19.3944
R12545 gnd.n4584 gnd.n3780 19.3944
R12546 gnd.n4584 gnd.n4583 19.3944
R12547 gnd.n4583 gnd.n3757 19.3944
R12548 gnd.n4609 gnd.n3757 19.3944
R12549 gnd.n4609 gnd.n3755 19.3944
R12550 gnd.n4615 gnd.n3755 19.3944
R12551 gnd.n4615 gnd.n4614 19.3944
R12552 gnd.n4614 gnd.n3730 19.3944
R12553 gnd.n4639 gnd.n3730 19.3944
R12554 gnd.n4639 gnd.n3728 19.3944
R12555 gnd.n4643 gnd.n3728 19.3944
R12556 gnd.n4643 gnd.n3708 19.3944
R12557 gnd.n4681 gnd.n3708 19.3944
R12558 gnd.n4681 gnd.n3706 19.3944
R12559 gnd.n4691 gnd.n3706 19.3944
R12560 gnd.n4691 gnd.n4690 19.3944
R12561 gnd.n4690 gnd.n4689 19.3944
R12562 gnd.n4689 gnd.n3551 19.3944
R12563 gnd.n5149 gnd.n3551 19.3944
R12564 gnd.n5149 gnd.n5148 19.3944
R12565 gnd.n5148 gnd.n5147 19.3944
R12566 gnd.n5147 gnd.n3555 19.3944
R12567 gnd.n3573 gnd.n3555 19.3944
R12568 gnd.n5135 gnd.n3573 19.3944
R12569 gnd.n5135 gnd.n5134 19.3944
R12570 gnd.n5134 gnd.n5133 19.3944
R12571 gnd.n5133 gnd.n3579 19.3944
R12572 gnd.n3597 gnd.n3579 19.3944
R12573 gnd.n5121 gnd.n3597 19.3944
R12574 gnd.n5121 gnd.n5120 19.3944
R12575 gnd.n5120 gnd.n5119 19.3944
R12576 gnd.n3630 gnd.n3629 19.3944
R12577 gnd.n5113 gnd.n3629 19.3944
R12578 gnd.n5113 gnd.n5112 19.3944
R12579 gnd.n5112 gnd.n5111 19.3944
R12580 gnd.n5111 gnd.n5108 19.3944
R12581 gnd.n5108 gnd.n5107 19.3944
R12582 gnd.n5107 gnd.n5104 19.3944
R12583 gnd.n5104 gnd.n5103 19.3944
R12584 gnd.n5103 gnd.n5100 19.3944
R12585 gnd.n5100 gnd.n5099 19.3944
R12586 gnd.n5099 gnd.n5096 19.3944
R12587 gnd.n5096 gnd.n5095 19.3944
R12588 gnd.n5095 gnd.n5092 19.3944
R12589 gnd.n5092 gnd.n5091 19.3944
R12590 gnd.n4036 gnd.n3932 19.3944
R12591 gnd.n4040 gnd.n3932 19.3944
R12592 gnd.n4040 gnd.n3922 19.3944
R12593 gnd.n4052 gnd.n3922 19.3944
R12594 gnd.n4052 gnd.n3920 19.3944
R12595 gnd.n4056 gnd.n3920 19.3944
R12596 gnd.n4056 gnd.n3909 19.3944
R12597 gnd.n4068 gnd.n3909 19.3944
R12598 gnd.n4068 gnd.n3907 19.3944
R12599 gnd.n4369 gnd.n3907 19.3944
R12600 gnd.n4369 gnd.n4368 19.3944
R12601 gnd.n4368 gnd.n4367 19.3944
R12602 gnd.n4367 gnd.n4366 19.3944
R12603 gnd.n4366 gnd.n4364 19.3944
R12604 gnd.n4364 gnd.n4363 19.3944
R12605 gnd.n4363 gnd.n4359 19.3944
R12606 gnd.n4359 gnd.n4358 19.3944
R12607 gnd.n4358 gnd.n4357 19.3944
R12608 gnd.n4357 gnd.n4355 19.3944
R12609 gnd.n4355 gnd.n4354 19.3944
R12610 gnd.n4354 gnd.n4351 19.3944
R12611 gnd.n4351 gnd.n4350 19.3944
R12612 gnd.n4350 gnd.n4349 19.3944
R12613 gnd.n4349 gnd.n4347 19.3944
R12614 gnd.n4347 gnd.n4346 19.3944
R12615 gnd.n4346 gnd.n4343 19.3944
R12616 gnd.n4343 gnd.n4342 19.3944
R12617 gnd.n4342 gnd.n4341 19.3944
R12618 gnd.n4341 gnd.n4339 19.3944
R12619 gnd.n4125 gnd.n4090 19.3944
R12620 gnd.n4122 gnd.n4121 19.3944
R12621 gnd.n4118 gnd.n4117 19.3944
R12622 gnd.n4113 gnd.n4112 19.3944
R12623 gnd.n4112 gnd.n4111 19.3944
R12624 gnd.n4111 gnd.n4109 19.3944
R12625 gnd.n4109 gnd.n4108 19.3944
R12626 gnd.n4108 gnd.n4104 19.3944
R12627 gnd.n4104 gnd.n4103 19.3944
R12628 gnd.n4103 gnd.n4102 19.3944
R12629 gnd.n4102 gnd.n4100 19.3944
R12630 gnd.n4100 gnd.n3715 19.3944
R12631 gnd.n4659 gnd.n3715 19.3944
R12632 gnd.n4659 gnd.n3713 19.3944
R12633 gnd.n4676 gnd.n3713 19.3944
R12634 gnd.n4676 gnd.n4675 19.3944
R12635 gnd.n4675 gnd.n4674 19.3944
R12636 gnd.n4674 gnd.n4672 19.3944
R12637 gnd.n4672 gnd.n4671 19.3944
R12638 gnd.n4671 gnd.n4668 19.3944
R12639 gnd.n4668 gnd.n3692 19.3944
R12640 gnd.n4719 gnd.n3692 19.3944
R12641 gnd.n4719 gnd.n3690 19.3944
R12642 gnd.n4735 gnd.n3690 19.3944
R12643 gnd.n4735 gnd.n4734 19.3944
R12644 gnd.n4734 gnd.n4733 19.3944
R12645 gnd.n4733 gnd.n4727 19.3944
R12646 gnd.n4727 gnd.n3684 19.3944
R12647 gnd.n5025 gnd.n3684 19.3944
R12648 gnd.n5026 gnd.n5025 19.3944
R12649 gnd.n5026 gnd.n3682 19.3944
R12650 gnd.n5030 gnd.n3682 19.3944
R12651 gnd.n4032 gnd.n3928 19.3944
R12652 gnd.n4044 gnd.n3928 19.3944
R12653 gnd.n4044 gnd.n3926 19.3944
R12654 gnd.n4048 gnd.n3926 19.3944
R12655 gnd.n4048 gnd.n3916 19.3944
R12656 gnd.n4060 gnd.n3916 19.3944
R12657 gnd.n4060 gnd.n3914 19.3944
R12658 gnd.n4064 gnd.n3914 19.3944
R12659 gnd.n4064 gnd.n3903 19.3944
R12660 gnd.n4433 gnd.n3903 19.3944
R12661 gnd.n4433 gnd.n3900 19.3944
R12662 gnd.n4438 gnd.n3900 19.3944
R12663 gnd.n4438 gnd.n3893 19.3944
R12664 gnd.n4449 gnd.n3893 19.3944
R12665 gnd.n4449 gnd.n4448 19.3944
R12666 gnd.n4448 gnd.n3876 19.3944
R12667 gnd.n4469 gnd.n3876 19.3944
R12668 gnd.n4469 gnd.n3868 19.3944
R12669 gnd.n4480 gnd.n3868 19.3944
R12670 gnd.n4480 gnd.n4479 19.3944
R12671 gnd.n4479 gnd.n3849 19.3944
R12672 gnd.n4500 gnd.n3849 19.3944
R12673 gnd.n4500 gnd.n3842 19.3944
R12674 gnd.n4511 gnd.n3842 19.3944
R12675 gnd.n4511 gnd.n4510 19.3944
R12676 gnd.n4510 gnd.n3823 19.3944
R12677 gnd.n4531 gnd.n3823 19.3944
R12678 gnd.n4531 gnd.n3816 19.3944
R12679 gnd.n4542 gnd.n3816 19.3944
R12680 gnd.n4542 gnd.n4541 19.3944
R12681 gnd.n4541 gnd.n3798 19.3944
R12682 gnd.n4562 gnd.n3798 19.3944
R12683 gnd.n4562 gnd.n3790 19.3944
R12684 gnd.n4573 gnd.n3790 19.3944
R12685 gnd.n4573 gnd.n4572 19.3944
R12686 gnd.n4572 gnd.n3773 19.3944
R12687 gnd.n4593 gnd.n3773 19.3944
R12688 gnd.n4593 gnd.n3765 19.3944
R12689 gnd.n4604 gnd.n3765 19.3944
R12690 gnd.n4604 gnd.n4603 19.3944
R12691 gnd.n4603 gnd.n3748 19.3944
R12692 gnd.n4624 gnd.n3748 19.3944
R12693 gnd.n4624 gnd.n3737 19.3944
R12694 gnd.n4634 gnd.n3737 19.3944
R12695 gnd.n4634 gnd.n3720 19.3944
R12696 gnd.n4655 gnd.n3720 19.3944
R12697 gnd.n4655 gnd.n4654 19.3944
R12698 gnd.n4654 gnd.n3699 19.3944
R12699 gnd.n4696 gnd.n3699 19.3944
R12700 gnd.n4696 gnd.n3540 19.3944
R12701 gnd.n5156 gnd.n3540 19.3944
R12702 gnd.n5156 gnd.n5155 19.3944
R12703 gnd.n5155 gnd.n5154 19.3944
R12704 gnd.n5154 gnd.n3544 19.3944
R12705 gnd.n3562 gnd.n3544 19.3944
R12706 gnd.n5142 gnd.n3562 19.3944
R12707 gnd.n5142 gnd.n5141 19.3944
R12708 gnd.n5141 gnd.n5140 19.3944
R12709 gnd.n5140 gnd.n3566 19.3944
R12710 gnd.n3587 gnd.n3566 19.3944
R12711 gnd.n5128 gnd.n3587 19.3944
R12712 gnd.n5128 gnd.n5127 19.3944
R12713 gnd.n5127 gnd.n5126 19.3944
R12714 gnd.n5126 gnd.n3591 19.3944
R12715 gnd.n5011 gnd.n3591 19.3944
R12716 gnd.n1016 gnd.n1015 19.3944
R12717 gnd.n1015 gnd.n909 19.3944
R12718 gnd.n6890 gnd.n909 19.3944
R12719 gnd.n6890 gnd.n910 19.3944
R12720 gnd.n6886 gnd.n910 19.3944
R12721 gnd.n6886 gnd.n6885 19.3944
R12722 gnd.n6885 gnd.n6884 19.3944
R12723 gnd.n6884 gnd.n915 19.3944
R12724 gnd.n6880 gnd.n915 19.3944
R12725 gnd.n6880 gnd.n6879 19.3944
R12726 gnd.n6879 gnd.n6878 19.3944
R12727 gnd.n6878 gnd.n919 19.3944
R12728 gnd.n6874 gnd.n919 19.3944
R12729 gnd.n6874 gnd.n6873 19.3944
R12730 gnd.n6873 gnd.n6872 19.3944
R12731 gnd.n6872 gnd.n923 19.3944
R12732 gnd.n6868 gnd.n923 19.3944
R12733 gnd.n6868 gnd.n6867 19.3944
R12734 gnd.n6867 gnd.n6866 19.3944
R12735 gnd.n6866 gnd.n927 19.3944
R12736 gnd.n6862 gnd.n927 19.3944
R12737 gnd.n6862 gnd.n6861 19.3944
R12738 gnd.n6861 gnd.n6860 19.3944
R12739 gnd.n6860 gnd.n6857 19.3944
R12740 gnd.n6857 gnd.n6856 19.3944
R12741 gnd.n6856 gnd.n466 19.3944
R12742 gnd.n7392 gnd.n466 19.3944
R12743 gnd.n7392 gnd.n7391 19.3944
R12744 gnd.n7391 gnd.n7390 19.3944
R12745 gnd.n7390 gnd.n471 19.3944
R12746 gnd.n7386 gnd.n471 19.3944
R12747 gnd.n7386 gnd.n7385 19.3944
R12748 gnd.n7385 gnd.n7384 19.3944
R12749 gnd.n7384 gnd.n476 19.3944
R12750 gnd.n7380 gnd.n476 19.3944
R12751 gnd.n7380 gnd.n7379 19.3944
R12752 gnd.n7379 gnd.n7378 19.3944
R12753 gnd.n7378 gnd.n481 19.3944
R12754 gnd.n7374 gnd.n481 19.3944
R12755 gnd.n7374 gnd.n7373 19.3944
R12756 gnd.n7373 gnd.n7372 19.3944
R12757 gnd.n7372 gnd.n486 19.3944
R12758 gnd.n7368 gnd.n486 19.3944
R12759 gnd.n7368 gnd.n7367 19.3944
R12760 gnd.n7367 gnd.n7366 19.3944
R12761 gnd.n7366 gnd.n491 19.3944
R12762 gnd.n7362 gnd.n491 19.3944
R12763 gnd.n7362 gnd.n7361 19.3944
R12764 gnd.n7361 gnd.n7360 19.3944
R12765 gnd.n7360 gnd.n496 19.3944
R12766 gnd.n7356 gnd.n496 19.3944
R12767 gnd.n7356 gnd.n7355 19.3944
R12768 gnd.n7264 gnd.n7263 19.3944
R12769 gnd.n7263 gnd.n7262 19.3944
R12770 gnd.n7262 gnd.n7211 19.3944
R12771 gnd.n7258 gnd.n7211 19.3944
R12772 gnd.n7258 gnd.n7257 19.3944
R12773 gnd.n7257 gnd.n7256 19.3944
R12774 gnd.n7256 gnd.n7219 19.3944
R12775 gnd.n7252 gnd.n7219 19.3944
R12776 gnd.n7252 gnd.n7251 19.3944
R12777 gnd.n7251 gnd.n7250 19.3944
R12778 gnd.n7250 gnd.n7227 19.3944
R12779 gnd.n7246 gnd.n7227 19.3944
R12780 gnd.n7246 gnd.n7245 19.3944
R12781 gnd.n7245 gnd.n7244 19.3944
R12782 gnd.n7010 gnd.n7009 19.3944
R12783 gnd.n7009 gnd.n793 19.3944
R12784 gnd.n7002 gnd.n793 19.3944
R12785 gnd.n7002 gnd.n7001 19.3944
R12786 gnd.n7001 gnd.n801 19.3944
R12787 gnd.n6994 gnd.n801 19.3944
R12788 gnd.n6994 gnd.n6993 19.3944
R12789 gnd.n6993 gnd.n809 19.3944
R12790 gnd.n6986 gnd.n809 19.3944
R12791 gnd.n6986 gnd.n6985 19.3944
R12792 gnd.n6985 gnd.n817 19.3944
R12793 gnd.n6978 gnd.n817 19.3944
R12794 gnd.n6978 gnd.n6977 19.3944
R12795 gnd.n6977 gnd.n825 19.3944
R12796 gnd.n7013 gnd.n777 19.3944
R12797 gnd.n7025 gnd.n777 19.3944
R12798 gnd.n7025 gnd.n775 19.3944
R12799 gnd.n7029 gnd.n775 19.3944
R12800 gnd.n7029 gnd.n759 19.3944
R12801 gnd.n7041 gnd.n759 19.3944
R12802 gnd.n7041 gnd.n757 19.3944
R12803 gnd.n7045 gnd.n757 19.3944
R12804 gnd.n7045 gnd.n741 19.3944
R12805 gnd.n7057 gnd.n741 19.3944
R12806 gnd.n7057 gnd.n739 19.3944
R12807 gnd.n7061 gnd.n739 19.3944
R12808 gnd.n7061 gnd.n724 19.3944
R12809 gnd.n7073 gnd.n724 19.3944
R12810 gnd.n7073 gnd.n722 19.3944
R12811 gnd.n7077 gnd.n722 19.3944
R12812 gnd.n7077 gnd.n706 19.3944
R12813 gnd.n7090 gnd.n706 19.3944
R12814 gnd.n7090 gnd.n704 19.3944
R12815 gnd.n7094 gnd.n704 19.3944
R12816 gnd.n7094 gnd.n689 19.3944
R12817 gnd.n7106 gnd.n689 19.3944
R12818 gnd.n7106 gnd.n687 19.3944
R12819 gnd.n7110 gnd.n687 19.3944
R12820 gnd.n7110 gnd.n673 19.3944
R12821 gnd.n7122 gnd.n673 19.3944
R12822 gnd.n7122 gnd.n670 19.3944
R12823 gnd.n7126 gnd.n670 19.3944
R12824 gnd.n7126 gnd.n658 19.3944
R12825 gnd.n7137 gnd.n658 19.3944
R12826 gnd.n7137 gnd.n656 19.3944
R12827 gnd.n7141 gnd.n656 19.3944
R12828 gnd.n7141 gnd.n641 19.3944
R12829 gnd.n7153 gnd.n641 19.3944
R12830 gnd.n7153 gnd.n639 19.3944
R12831 gnd.n7157 gnd.n639 19.3944
R12832 gnd.n7157 gnd.n624 19.3944
R12833 gnd.n7169 gnd.n624 19.3944
R12834 gnd.n7169 gnd.n622 19.3944
R12835 gnd.n7173 gnd.n622 19.3944
R12836 gnd.n7173 gnd.n608 19.3944
R12837 gnd.n7185 gnd.n608 19.3944
R12838 gnd.n7185 gnd.n606 19.3944
R12839 gnd.n7189 gnd.n606 19.3944
R12840 gnd.n7189 gnd.n591 19.3944
R12841 gnd.n7201 gnd.n591 19.3944
R12842 gnd.n7201 gnd.n588 19.3944
R12843 gnd.n7273 gnd.n588 19.3944
R12844 gnd.n7273 gnd.n589 19.3944
R12845 gnd.n7269 gnd.n589 19.3944
R12846 gnd.n7269 gnd.n7268 19.3944
R12847 gnd.n7268 gnd.n7267 19.3944
R12848 gnd.n1696 gnd.n1619 19.3944
R12849 gnd.n1696 gnd.n1694 19.3944
R12850 gnd.n5802 gnd.n1694 19.3944
R12851 gnd.n5802 gnd.n5801 19.3944
R12852 gnd.n5801 gnd.n1703 19.3944
R12853 gnd.n5794 gnd.n1703 19.3944
R12854 gnd.n5794 gnd.n5793 19.3944
R12855 gnd.n5793 gnd.n1714 19.3944
R12856 gnd.n5786 gnd.n1714 19.3944
R12857 gnd.n5786 gnd.n5785 19.3944
R12858 gnd.n5785 gnd.n1725 19.3944
R12859 gnd.n5778 gnd.n1725 19.3944
R12860 gnd.n5778 gnd.n5777 19.3944
R12861 gnd.n5777 gnd.n1737 19.3944
R12862 gnd.n3031 gnd.n2664 19.3944
R12863 gnd.n3025 gnd.n2664 19.3944
R12864 gnd.n3025 gnd.n3024 19.3944
R12865 gnd.n3024 gnd.n3023 19.3944
R12866 gnd.n3023 gnd.n2671 19.3944
R12867 gnd.n3017 gnd.n2671 19.3944
R12868 gnd.n3017 gnd.n3016 19.3944
R12869 gnd.n3016 gnd.n3015 19.3944
R12870 gnd.n3015 gnd.n2679 19.3944
R12871 gnd.n3009 gnd.n2679 19.3944
R12872 gnd.n3009 gnd.n3008 19.3944
R12873 gnd.n3008 gnd.n3007 19.3944
R12874 gnd.n3007 gnd.n2687 19.3944
R12875 gnd.n3001 gnd.n2687 19.3944
R12876 gnd.n3001 gnd.n3000 19.3944
R12877 gnd.n3000 gnd.n2999 19.3944
R12878 gnd.n2999 gnd.n2695 19.3944
R12879 gnd.n2993 gnd.n2695 19.3944
R12880 gnd.n2993 gnd.n2992 19.3944
R12881 gnd.n2992 gnd.n2991 19.3944
R12882 gnd.n2991 gnd.n2703 19.3944
R12883 gnd.n2985 gnd.n2703 19.3944
R12884 gnd.n2985 gnd.n2984 19.3944
R12885 gnd.n2984 gnd.n2983 19.3944
R12886 gnd.n2983 gnd.n2711 19.3944
R12887 gnd.n2977 gnd.n2711 19.3944
R12888 gnd.n2977 gnd.n2976 19.3944
R12889 gnd.n2976 gnd.n2975 19.3944
R12890 gnd.n2975 gnd.n2719 19.3944
R12891 gnd.n2969 gnd.n2719 19.3944
R12892 gnd.n2969 gnd.n2968 19.3944
R12893 gnd.n2968 gnd.n2967 19.3944
R12894 gnd.n2967 gnd.n2727 19.3944
R12895 gnd.n2961 gnd.n2727 19.3944
R12896 gnd.n2961 gnd.n2960 19.3944
R12897 gnd.n2960 gnd.n2959 19.3944
R12898 gnd.n2959 gnd.n2735 19.3944
R12899 gnd.n2953 gnd.n2735 19.3944
R12900 gnd.n2953 gnd.n2952 19.3944
R12901 gnd.n2952 gnd.n2951 19.3944
R12902 gnd.n2951 gnd.n2743 19.3944
R12903 gnd.n2945 gnd.n2743 19.3944
R12904 gnd.n2945 gnd.n2944 19.3944
R12905 gnd.n2944 gnd.n2943 19.3944
R12906 gnd.n2943 gnd.n2751 19.3944
R12907 gnd.n2937 gnd.n2751 19.3944
R12908 gnd.n2937 gnd.n2936 19.3944
R12909 gnd.n2936 gnd.n2935 19.3944
R12910 gnd.n2935 gnd.n2759 19.3944
R12911 gnd.n2929 gnd.n2759 19.3944
R12912 gnd.n2929 gnd.n2928 19.3944
R12913 gnd.n2928 gnd.n2927 19.3944
R12914 gnd.n2927 gnd.n2767 19.3944
R12915 gnd.n2921 gnd.n2767 19.3944
R12916 gnd.n2921 gnd.n2920 19.3944
R12917 gnd.n2920 gnd.n2919 19.3944
R12918 gnd.n2919 gnd.n2775 19.3944
R12919 gnd.n2913 gnd.n2775 19.3944
R12920 gnd.n2913 gnd.n2912 19.3944
R12921 gnd.n2912 gnd.n2911 19.3944
R12922 gnd.n2911 gnd.n2783 19.3944
R12923 gnd.n2905 gnd.n2783 19.3944
R12924 gnd.n2905 gnd.n2904 19.3944
R12925 gnd.n2904 gnd.n2903 19.3944
R12926 gnd.n2903 gnd.n2791 19.3944
R12927 gnd.n2897 gnd.n2791 19.3944
R12928 gnd.n3371 gnd.n2325 19.3944
R12929 gnd.n3371 gnd.n3370 19.3944
R12930 gnd.n3370 gnd.n3369 19.3944
R12931 gnd.n3369 gnd.n2329 19.3944
R12932 gnd.n3363 gnd.n2329 19.3944
R12933 gnd.n3363 gnd.n3362 19.3944
R12934 gnd.n3362 gnd.n3361 19.3944
R12935 gnd.n3361 gnd.n2337 19.3944
R12936 gnd.n3355 gnd.n2337 19.3944
R12937 gnd.n3355 gnd.n3354 19.3944
R12938 gnd.n3354 gnd.n3353 19.3944
R12939 gnd.n3353 gnd.n2345 19.3944
R12940 gnd.n3347 gnd.n2345 19.3944
R12941 gnd.n3347 gnd.n3346 19.3944
R12942 gnd.n3346 gnd.n3345 19.3944
R12943 gnd.n3345 gnd.n2353 19.3944
R12944 gnd.n3339 gnd.n2353 19.3944
R12945 gnd.n3339 gnd.n3338 19.3944
R12946 gnd.n3338 gnd.n3337 19.3944
R12947 gnd.n3337 gnd.n2361 19.3944
R12948 gnd.n3331 gnd.n2361 19.3944
R12949 gnd.n3331 gnd.n3330 19.3944
R12950 gnd.n3330 gnd.n3329 19.3944
R12951 gnd.n3329 gnd.n2369 19.3944
R12952 gnd.n3323 gnd.n2369 19.3944
R12953 gnd.n3323 gnd.n3322 19.3944
R12954 gnd.n3322 gnd.n3321 19.3944
R12955 gnd.n3321 gnd.n2377 19.3944
R12956 gnd.n3315 gnd.n2377 19.3944
R12957 gnd.n3315 gnd.n3314 19.3944
R12958 gnd.n3314 gnd.n3313 19.3944
R12959 gnd.n3313 gnd.n2385 19.3944
R12960 gnd.n3307 gnd.n2385 19.3944
R12961 gnd.n3307 gnd.n3306 19.3944
R12962 gnd.n3306 gnd.n3305 19.3944
R12963 gnd.n3305 gnd.n2393 19.3944
R12964 gnd.n3299 gnd.n2393 19.3944
R12965 gnd.n3299 gnd.n3298 19.3944
R12966 gnd.n3298 gnd.n3297 19.3944
R12967 gnd.n3297 gnd.n2401 19.3944
R12968 gnd.n3291 gnd.n2401 19.3944
R12969 gnd.n3291 gnd.n3290 19.3944
R12970 gnd.n3290 gnd.n3289 19.3944
R12971 gnd.n3289 gnd.n2409 19.3944
R12972 gnd.n3283 gnd.n2409 19.3944
R12973 gnd.n3283 gnd.n3282 19.3944
R12974 gnd.n3282 gnd.n3281 19.3944
R12975 gnd.n3281 gnd.n2417 19.3944
R12976 gnd.n3275 gnd.n2417 19.3944
R12977 gnd.n3275 gnd.n3274 19.3944
R12978 gnd.n3274 gnd.n3273 19.3944
R12979 gnd.n3273 gnd.n2425 19.3944
R12980 gnd.n3267 gnd.n2425 19.3944
R12981 gnd.n3267 gnd.n3266 19.3944
R12982 gnd.n3266 gnd.n3265 19.3944
R12983 gnd.n3265 gnd.n2433 19.3944
R12984 gnd.n3259 gnd.n2433 19.3944
R12985 gnd.n3259 gnd.n3258 19.3944
R12986 gnd.n3258 gnd.n3257 19.3944
R12987 gnd.n3257 gnd.n2441 19.3944
R12988 gnd.n3251 gnd.n2441 19.3944
R12989 gnd.n3251 gnd.n3250 19.3944
R12990 gnd.n3250 gnd.n3249 19.3944
R12991 gnd.n3249 gnd.n2449 19.3944
R12992 gnd.n3243 gnd.n2449 19.3944
R12993 gnd.n3243 gnd.n3242 19.3944
R12994 gnd.n3242 gnd.n3241 19.3944
R12995 gnd.n3241 gnd.n2457 19.3944
R12996 gnd.n3235 gnd.n2457 19.3944
R12997 gnd.n3235 gnd.n3234 19.3944
R12998 gnd.n3234 gnd.n3233 19.3944
R12999 gnd.n3233 gnd.n2465 19.3944
R13000 gnd.n3227 gnd.n2465 19.3944
R13001 gnd.n3227 gnd.n3226 19.3944
R13002 gnd.n3226 gnd.n3225 19.3944
R13003 gnd.n3225 gnd.n2473 19.3944
R13004 gnd.n3219 gnd.n2473 19.3944
R13005 gnd.n3219 gnd.n3218 19.3944
R13006 gnd.n3218 gnd.n3217 19.3944
R13007 gnd.n3217 gnd.n2481 19.3944
R13008 gnd.n3211 gnd.n2481 19.3944
R13009 gnd.n3211 gnd.n3210 19.3944
R13010 gnd.n3210 gnd.n3209 19.3944
R13011 gnd.n3209 gnd.n2489 19.3944
R13012 gnd.n3203 gnd.n2489 19.3944
R13013 gnd.n3203 gnd.n3202 19.3944
R13014 gnd.n3202 gnd.n3201 19.3944
R13015 gnd.n3201 gnd.n2497 19.3944
R13016 gnd.n3195 gnd.n2497 19.3944
R13017 gnd.n3195 gnd.n3194 19.3944
R13018 gnd.n3194 gnd.n3193 19.3944
R13019 gnd.n3193 gnd.n2505 19.3944
R13020 gnd.n3187 gnd.n2505 19.3944
R13021 gnd.n3187 gnd.n3186 19.3944
R13022 gnd.n3186 gnd.n3185 19.3944
R13023 gnd.n3185 gnd.n2513 19.3944
R13024 gnd.n3179 gnd.n2513 19.3944
R13025 gnd.n3179 gnd.n3178 19.3944
R13026 gnd.n3178 gnd.n3177 19.3944
R13027 gnd.n3177 gnd.n2521 19.3944
R13028 gnd.n3171 gnd.n2521 19.3944
R13029 gnd.n3171 gnd.n3170 19.3944
R13030 gnd.n3170 gnd.n3169 19.3944
R13031 gnd.n3169 gnd.n2529 19.3944
R13032 gnd.n3163 gnd.n2529 19.3944
R13033 gnd.n3163 gnd.n3162 19.3944
R13034 gnd.n3162 gnd.n3161 19.3944
R13035 gnd.n3161 gnd.n2537 19.3944
R13036 gnd.n3155 gnd.n2537 19.3944
R13037 gnd.n3155 gnd.n3154 19.3944
R13038 gnd.n3154 gnd.n3153 19.3944
R13039 gnd.n3153 gnd.n2545 19.3944
R13040 gnd.n3147 gnd.n2545 19.3944
R13041 gnd.n3147 gnd.n3146 19.3944
R13042 gnd.n3146 gnd.n3145 19.3944
R13043 gnd.n3145 gnd.n2553 19.3944
R13044 gnd.n3139 gnd.n2553 19.3944
R13045 gnd.n3139 gnd.n3138 19.3944
R13046 gnd.n3138 gnd.n3137 19.3944
R13047 gnd.n3137 gnd.n2561 19.3944
R13048 gnd.n3131 gnd.n2561 19.3944
R13049 gnd.n3131 gnd.n3130 19.3944
R13050 gnd.n3130 gnd.n3129 19.3944
R13051 gnd.n3129 gnd.n2569 19.3944
R13052 gnd.n3123 gnd.n2569 19.3944
R13053 gnd.n3123 gnd.n3122 19.3944
R13054 gnd.n3122 gnd.n3121 19.3944
R13055 gnd.n3121 gnd.n2577 19.3944
R13056 gnd.n3115 gnd.n2577 19.3944
R13057 gnd.n3115 gnd.n3114 19.3944
R13058 gnd.n3114 gnd.n3113 19.3944
R13059 gnd.n3113 gnd.n2585 19.3944
R13060 gnd.n3107 gnd.n2585 19.3944
R13061 gnd.n3107 gnd.n3106 19.3944
R13062 gnd.n3106 gnd.n3105 19.3944
R13063 gnd.n3105 gnd.n2593 19.3944
R13064 gnd.n3099 gnd.n2593 19.3944
R13065 gnd.n3099 gnd.n3098 19.3944
R13066 gnd.n3098 gnd.n3097 19.3944
R13067 gnd.n3097 gnd.n2601 19.3944
R13068 gnd.n3091 gnd.n2601 19.3944
R13069 gnd.n3091 gnd.n3090 19.3944
R13070 gnd.n3090 gnd.n3089 19.3944
R13071 gnd.n3089 gnd.n2609 19.3944
R13072 gnd.n3083 gnd.n2609 19.3944
R13073 gnd.n3083 gnd.n3082 19.3944
R13074 gnd.n3082 gnd.n3081 19.3944
R13075 gnd.n3081 gnd.n2617 19.3944
R13076 gnd.n3075 gnd.n2617 19.3944
R13077 gnd.n3075 gnd.n3074 19.3944
R13078 gnd.n3074 gnd.n3073 19.3944
R13079 gnd.n3073 gnd.n2625 19.3944
R13080 gnd.n3067 gnd.n2625 19.3944
R13081 gnd.n3067 gnd.n3066 19.3944
R13082 gnd.n3066 gnd.n3065 19.3944
R13083 gnd.n3065 gnd.n2633 19.3944
R13084 gnd.n3059 gnd.n2633 19.3944
R13085 gnd.n3059 gnd.n3058 19.3944
R13086 gnd.n3058 gnd.n3057 19.3944
R13087 gnd.n3057 gnd.n2641 19.3944
R13088 gnd.n3051 gnd.n2641 19.3944
R13089 gnd.n3051 gnd.n3050 19.3944
R13090 gnd.n3050 gnd.n3049 19.3944
R13091 gnd.n3049 gnd.n2649 19.3944
R13092 gnd.n3043 gnd.n2649 19.3944
R13093 gnd.n3043 gnd.n3042 19.3944
R13094 gnd.n3042 gnd.n3041 19.3944
R13095 gnd.n3041 gnd.n2657 19.3944
R13096 gnd.n3035 gnd.n2657 19.3944
R13097 gnd.n3035 gnd.n3034 19.3944
R13098 gnd.n6961 gnd.n863 19.3944
R13099 gnd.n6961 gnd.n6960 19.3944
R13100 gnd.n6960 gnd.n6959 19.3944
R13101 gnd.n6959 gnd.n6957 19.3944
R13102 gnd.n6957 gnd.n6954 19.3944
R13103 gnd.n6954 gnd.n6953 19.3944
R13104 gnd.n6953 gnd.n6950 19.3944
R13105 gnd.n6950 gnd.n6949 19.3944
R13106 gnd.n6949 gnd.n6946 19.3944
R13107 gnd.n6946 gnd.n6945 19.3944
R13108 gnd.n6945 gnd.n6942 19.3944
R13109 gnd.n6942 gnd.n6941 19.3944
R13110 gnd.n6941 gnd.n6938 19.3944
R13111 gnd.n6936 gnd.n6933 19.3944
R13112 gnd.n6933 gnd.n6932 19.3944
R13113 gnd.n6932 gnd.n6929 19.3944
R13114 gnd.n6929 gnd.n6928 19.3944
R13115 gnd.n6928 gnd.n6925 19.3944
R13116 gnd.n6925 gnd.n6924 19.3944
R13117 gnd.n6924 gnd.n6921 19.3944
R13118 gnd.n6921 gnd.n6920 19.3944
R13119 gnd.n6920 gnd.n6917 19.3944
R13120 gnd.n6917 gnd.n6916 19.3944
R13121 gnd.n6916 gnd.n6913 19.3944
R13122 gnd.n6913 gnd.n6912 19.3944
R13123 gnd.n6912 gnd.n6909 19.3944
R13124 gnd.n6909 gnd.n6908 19.3944
R13125 gnd.n6908 gnd.n6905 19.3944
R13126 gnd.n6905 gnd.n6904 19.3944
R13127 gnd.n6897 gnd.n6896 19.3944
R13128 gnd.n6896 gnd.n6895 19.3944
R13129 gnd.n6895 gnd.n6894 19.3944
R13130 gnd.n6894 gnd.n907 19.3944
R13131 gnd.n6760 gnd.n907 19.3944
R13132 gnd.n6760 gnd.n6756 19.3944
R13133 gnd.n6766 gnd.n6756 19.3944
R13134 gnd.n6767 gnd.n6766 19.3944
R13135 gnd.n6770 gnd.n6767 19.3944
R13136 gnd.n6770 gnd.n6754 19.3944
R13137 gnd.n6776 gnd.n6754 19.3944
R13138 gnd.n6777 gnd.n6776 19.3944
R13139 gnd.n6780 gnd.n6777 19.3944
R13140 gnd.n6780 gnd.n6752 19.3944
R13141 gnd.n6809 gnd.n6752 19.3944
R13142 gnd.n6809 gnd.n6808 19.3944
R13143 gnd.n6808 gnd.n6807 19.3944
R13144 gnd.n6807 gnd.n6804 19.3944
R13145 gnd.n6804 gnd.n6803 19.3944
R13146 gnd.n6803 gnd.n6800 19.3944
R13147 gnd.n6800 gnd.n6799 19.3944
R13148 gnd.n6799 gnd.n6796 19.3944
R13149 gnd.n6796 gnd.n6795 19.3944
R13150 gnd.n6795 gnd.n931 19.3944
R13151 gnd.n6852 gnd.n931 19.3944
R13152 gnd.n6852 gnd.n6851 19.3944
R13153 gnd.n6851 gnd.n6850 19.3944
R13154 gnd.n6850 gnd.n6847 19.3944
R13155 gnd.n6847 gnd.n6846 19.3944
R13156 gnd.n6846 gnd.n936 19.3944
R13157 gnd.n2842 gnd.n936 19.3944
R13158 gnd.n2843 gnd.n2842 19.3944
R13159 gnd.n2846 gnd.n2843 19.3944
R13160 gnd.n2846 gnd.n2836 19.3944
R13161 gnd.n2852 gnd.n2836 19.3944
R13162 gnd.n2853 gnd.n2852 19.3944
R13163 gnd.n2856 gnd.n2853 19.3944
R13164 gnd.n2856 gnd.n2834 19.3944
R13165 gnd.n2862 gnd.n2834 19.3944
R13166 gnd.n2863 gnd.n2862 19.3944
R13167 gnd.n2866 gnd.n2863 19.3944
R13168 gnd.n2866 gnd.n2832 19.3944
R13169 gnd.n2886 gnd.n2832 19.3944
R13170 gnd.n2886 gnd.n2885 19.3944
R13171 gnd.n2885 gnd.n2884 19.3944
R13172 gnd.n2884 gnd.n2881 19.3944
R13173 gnd.n2881 gnd.n2880 19.3944
R13174 gnd.n2880 gnd.n2878 19.3944
R13175 gnd.n2878 gnd.n2877 19.3944
R13176 gnd.n2877 gnd.n574 19.3944
R13177 gnd.n7286 gnd.n574 19.3944
R13178 gnd.n7287 gnd.n7286 19.3944
R13179 gnd.n7320 gnd.n7319 19.3944
R13180 gnd.n7319 gnd.n7318 19.3944
R13181 gnd.n7318 gnd.n542 19.3944
R13182 gnd.n7313 gnd.n542 19.3944
R13183 gnd.n7313 gnd.n7312 19.3944
R13184 gnd.n7312 gnd.n7311 19.3944
R13185 gnd.n7311 gnd.n549 19.3944
R13186 gnd.n7306 gnd.n549 19.3944
R13187 gnd.n7306 gnd.n7305 19.3944
R13188 gnd.n7305 gnd.n7304 19.3944
R13189 gnd.n7304 gnd.n556 19.3944
R13190 gnd.n7299 gnd.n556 19.3944
R13191 gnd.n7299 gnd.n7298 19.3944
R13192 gnd.n7298 gnd.n7297 19.3944
R13193 gnd.n7297 gnd.n563 19.3944
R13194 gnd.n7292 gnd.n563 19.3944
R13195 gnd.n7348 gnd.n7347 19.3944
R13196 gnd.n7347 gnd.n7346 19.3944
R13197 gnd.n7346 gnd.n511 19.3944
R13198 gnd.n7341 gnd.n511 19.3944
R13199 gnd.n7341 gnd.n7340 19.3944
R13200 gnd.n7340 gnd.n7339 19.3944
R13201 gnd.n7339 gnd.n518 19.3944
R13202 gnd.n7334 gnd.n518 19.3944
R13203 gnd.n7334 gnd.n7333 19.3944
R13204 gnd.n7333 gnd.n7332 19.3944
R13205 gnd.n7332 gnd.n525 19.3944
R13206 gnd.n7327 gnd.n525 19.3944
R13207 gnd.n7327 gnd.n7326 19.3944
R13208 gnd.n7326 gnd.n7325 19.3944
R13209 gnd.n7325 gnd.n532 19.3944
R13210 gnd.n7017 gnd.n783 19.3944
R13211 gnd.n7021 gnd.n783 19.3944
R13212 gnd.n7021 gnd.n768 19.3944
R13213 gnd.n7033 gnd.n768 19.3944
R13214 gnd.n7033 gnd.n766 19.3944
R13215 gnd.n7037 gnd.n766 19.3944
R13216 gnd.n7037 gnd.n750 19.3944
R13217 gnd.n7049 gnd.n750 19.3944
R13218 gnd.n7049 gnd.n748 19.3944
R13219 gnd.n7053 gnd.n748 19.3944
R13220 gnd.n7053 gnd.n732 19.3944
R13221 gnd.n7065 gnd.n732 19.3944
R13222 gnd.n7065 gnd.n730 19.3944
R13223 gnd.n7069 gnd.n730 19.3944
R13224 gnd.n7069 gnd.n715 19.3944
R13225 gnd.n7081 gnd.n715 19.3944
R13226 gnd.n7081 gnd.n713 19.3944
R13227 gnd.n7086 gnd.n713 19.3944
R13228 gnd.n7086 gnd.n696 19.3944
R13229 gnd.n7098 gnd.n696 19.3944
R13230 gnd.n7099 gnd.n7098 19.3944
R13231 gnd.n7102 gnd.n7101 19.3944
R13232 gnd.n7115 gnd.n7114 19.3944
R13233 gnd.n7118 gnd.n7117 19.3944
R13234 gnd.n7131 gnd.n7130 19.3944
R13235 gnd.n7133 gnd.n650 19.3944
R13236 gnd.n7145 gnd.n650 19.3944
R13237 gnd.n7145 gnd.n648 19.3944
R13238 gnd.n7149 gnd.n648 19.3944
R13239 gnd.n7149 gnd.n633 19.3944
R13240 gnd.n7161 gnd.n633 19.3944
R13241 gnd.n7161 gnd.n631 19.3944
R13242 gnd.n7165 gnd.n631 19.3944
R13243 gnd.n7165 gnd.n616 19.3944
R13244 gnd.n7177 gnd.n616 19.3944
R13245 gnd.n7177 gnd.n614 19.3944
R13246 gnd.n7181 gnd.n614 19.3944
R13247 gnd.n7181 gnd.n600 19.3944
R13248 gnd.n7193 gnd.n600 19.3944
R13249 gnd.n7193 gnd.n598 19.3944
R13250 gnd.n7197 gnd.n598 19.3944
R13251 gnd.n7197 gnd.n581 19.3944
R13252 gnd.n7277 gnd.n581 19.3944
R13253 gnd.n7277 gnd.n579 19.3944
R13254 gnd.n7281 gnd.n579 19.3944
R13255 gnd.n7281 gnd.n506 19.3944
R13256 gnd.n7351 gnd.n506 19.3944
R13257 gnd.n5171 gnd.n2222 19.3944
R13258 gnd.n5171 gnd.n2220 19.3944
R13259 gnd.n5218 gnd.n2220 19.3944
R13260 gnd.n5218 gnd.n5217 19.3944
R13261 gnd.n5217 gnd.n5216 19.3944
R13262 gnd.n5216 gnd.n5177 19.3944
R13263 gnd.n5212 gnd.n5177 19.3944
R13264 gnd.n5212 gnd.n5211 19.3944
R13265 gnd.n5211 gnd.n5210 19.3944
R13266 gnd.n5210 gnd.n5183 19.3944
R13267 gnd.n5206 gnd.n5183 19.3944
R13268 gnd.n5206 gnd.n5205 19.3944
R13269 gnd.n5205 gnd.n5204 19.3944
R13270 gnd.n5204 gnd.n5190 19.3944
R13271 gnd.n5200 gnd.n5190 19.3944
R13272 gnd.n5198 gnd.n5197 19.3944
R13273 gnd.n5194 gnd.n5193 19.3944
R13274 gnd.n5629 gnd.n5628 19.3944
R13275 gnd.n5626 gnd.n1872 19.3944
R13276 gnd.n5463 gnd.n5460 19.3944
R13277 gnd.n5463 gnd.n5458 19.3944
R13278 gnd.n5467 gnd.n5458 19.3944
R13279 gnd.n5467 gnd.n5456 19.3944
R13280 gnd.n5471 gnd.n5456 19.3944
R13281 gnd.n5471 gnd.n5454 19.3944
R13282 gnd.n5475 gnd.n5454 19.3944
R13283 gnd.n5475 gnd.n5452 19.3944
R13284 gnd.n5516 gnd.n5452 19.3944
R13285 gnd.n5516 gnd.n5450 19.3944
R13286 gnd.n5520 gnd.n5450 19.3944
R13287 gnd.n5520 gnd.n5448 19.3944
R13288 gnd.n5524 gnd.n5448 19.3944
R13289 gnd.n5524 gnd.n5446 19.3944
R13290 gnd.n5528 gnd.n5446 19.3944
R13291 gnd.n5528 gnd.n5444 19.3944
R13292 gnd.n5532 gnd.n5444 19.3944
R13293 gnd.n5532 gnd.n5442 19.3944
R13294 gnd.n5556 gnd.n5442 19.3944
R13295 gnd.n5556 gnd.n5555 19.3944
R13296 gnd.n5555 gnd.n5554 19.3944
R13297 gnd.n5554 gnd.n5538 19.3944
R13298 gnd.n5549 gnd.n5538 19.3944
R13299 gnd.n5549 gnd.n5548 19.3944
R13300 gnd.n5548 gnd.n5547 19.3944
R13301 gnd.n5547 gnd.n1673 19.3944
R13302 gnd.n5812 gnd.n1673 19.3944
R13303 gnd.n5812 gnd.n1671 19.3944
R13304 gnd.n5816 gnd.n1671 19.3944
R13305 gnd.n5816 gnd.n1661 19.3944
R13306 gnd.n5832 gnd.n1661 19.3944
R13307 gnd.n5832 gnd.n1659 19.3944
R13308 gnd.n5836 gnd.n1659 19.3944
R13309 gnd.n5836 gnd.n1648 19.3944
R13310 gnd.n5852 gnd.n1648 19.3944
R13311 gnd.n5852 gnd.n1646 19.3944
R13312 gnd.n5858 gnd.n1646 19.3944
R13313 gnd.n5858 gnd.n5857 19.3944
R13314 gnd.n5857 gnd.n1430 19.3944
R13315 gnd.n6063 gnd.n1430 19.3944
R13316 gnd.n6063 gnd.n1428 19.3944
R13317 gnd.n6069 gnd.n1428 19.3944
R13318 gnd.n6069 gnd.n6068 19.3944
R13319 gnd.n6068 gnd.n1397 19.3944
R13320 gnd.n6145 gnd.n1397 19.3944
R13321 gnd.n6145 gnd.n1395 19.3944
R13322 gnd.n6149 gnd.n1395 19.3944
R13323 gnd.n6149 gnd.n1373 19.3944
R13324 gnd.n6173 gnd.n1373 19.3944
R13325 gnd.n6173 gnd.n1371 19.3944
R13326 gnd.n6192 gnd.n1371 19.3944
R13327 gnd.n6192 gnd.n6191 19.3944
R13328 gnd.n6191 gnd.n6190 19.3944
R13329 gnd.n6190 gnd.n6179 19.3944
R13330 gnd.n6185 gnd.n6179 19.3944
R13331 gnd.n6185 gnd.n6184 19.3944
R13332 gnd.n6184 gnd.n1312 19.3944
R13333 gnd.n6284 gnd.n1312 19.3944
R13334 gnd.n6284 gnd.n1310 19.3944
R13335 gnd.n6301 gnd.n1310 19.3944
R13336 gnd.n6301 gnd.n6300 19.3944
R13337 gnd.n6300 gnd.n6299 19.3944
R13338 gnd.n6299 gnd.n6290 19.3944
R13339 gnd.n6294 gnd.n6290 19.3944
R13340 gnd.n6294 gnd.n1268 19.3944
R13341 gnd.n6387 gnd.n1268 19.3944
R13342 gnd.n6387 gnd.n6386 19.3944
R13343 gnd.n6386 gnd.n6385 19.3944
R13344 gnd.n6385 gnd.n1239 19.3944
R13345 gnd.n6424 gnd.n1239 19.3944
R13346 gnd.n6424 gnd.n6423 19.3944
R13347 gnd.n6423 gnd.n6422 19.3944
R13348 gnd.n6422 gnd.n1210 19.3944
R13349 gnd.n6464 gnd.n1210 19.3944
R13350 gnd.n6464 gnd.n6463 19.3944
R13351 gnd.n6463 gnd.n6462 19.3944
R13352 gnd.n6462 gnd.n1215 19.3944
R13353 gnd.n1215 gnd.n1107 19.3944
R13354 gnd.n6613 gnd.n1107 19.3944
R13355 gnd.n6613 gnd.n1105 19.3944
R13356 gnd.n6619 gnd.n1105 19.3944
R13357 gnd.n6619 gnd.n6618 19.3944
R13358 gnd.n6618 gnd.n1081 19.3944
R13359 gnd.n6643 gnd.n1081 19.3944
R13360 gnd.n6643 gnd.n1079 19.3944
R13361 gnd.n6649 gnd.n1079 19.3944
R13362 gnd.n6649 gnd.n6648 19.3944
R13363 gnd.n6648 gnd.n1056 19.3944
R13364 gnd.n6674 gnd.n1056 19.3944
R13365 gnd.n6674 gnd.n1054 19.3944
R13366 gnd.n6691 gnd.n1054 19.3944
R13367 gnd.n6691 gnd.n6690 19.3944
R13368 gnd.n6690 gnd.n6689 19.3944
R13369 gnd.n6689 gnd.n6680 19.3944
R13370 gnd.n6683 gnd.n6680 19.3944
R13371 gnd.n6683 gnd.n971 19.3944
R13372 gnd.n6715 gnd.n971 19.3944
R13373 gnd.n6715 gnd.n969 19.3944
R13374 gnd.n6719 gnd.n969 19.3944
R13375 gnd.n6719 gnd.n967 19.3944
R13376 gnd.n6723 gnd.n967 19.3944
R13377 gnd.n6723 gnd.n965 19.3944
R13378 gnd.n6727 gnd.n965 19.3944
R13379 gnd.n6727 gnd.n963 19.3944
R13380 gnd.n6731 gnd.n963 19.3944
R13381 gnd.n6731 gnd.n961 19.3944
R13382 gnd.n6735 gnd.n961 19.3944
R13383 gnd.n6735 gnd.n959 19.3944
R13384 gnd.n6739 gnd.n959 19.3944
R13385 gnd.n6739 gnd.n957 19.3944
R13386 gnd.n6743 gnd.n957 19.3944
R13387 gnd.n6743 gnd.n955 19.3944
R13388 gnd.n6747 gnd.n955 19.3944
R13389 gnd.n6747 gnd.n953 19.3944
R13390 gnd.n6751 gnd.n953 19.3944
R13391 gnd.n6751 gnd.n951 19.3944
R13392 gnd.n6816 gnd.n951 19.3944
R13393 gnd.n6816 gnd.n949 19.3944
R13394 gnd.n6820 gnd.n949 19.3944
R13395 gnd.n6820 gnd.n946 19.3944
R13396 gnd.n6836 gnd.n946 19.3944
R13397 gnd.n6836 gnd.n947 19.3944
R13398 gnd.n6832 gnd.n6831 19.3944
R13399 gnd.n6828 gnd.n6827 19.3944
R13400 gnd.n6824 gnd.n6823 19.3944
R13401 gnd.n6841 gnd.n6840 19.3944
R13402 gnd.n2806 gnd.n940 19.3944
R13403 gnd.n2810 gnd.n2806 19.3944
R13404 gnd.n2810 gnd.n2805 19.3944
R13405 gnd.n2814 gnd.n2805 19.3944
R13406 gnd.n2814 gnd.n2803 19.3944
R13407 gnd.n2818 gnd.n2803 19.3944
R13408 gnd.n2818 gnd.n2801 19.3944
R13409 gnd.n2822 gnd.n2801 19.3944
R13410 gnd.n2822 gnd.n2799 19.3944
R13411 gnd.n2826 gnd.n2799 19.3944
R13412 gnd.n2826 gnd.n2797 19.3944
R13413 gnd.n2831 gnd.n2797 19.3944
R13414 gnd.n2831 gnd.n2795 19.3944
R13415 gnd.n2893 gnd.n2795 19.3944
R13416 gnd.n2894 gnd.n2893 19.3944
R13417 gnd.n2088 gnd.n2085 19.3944
R13418 gnd.n2088 gnd.n2084 19.3944
R13419 gnd.n2092 gnd.n2084 19.3944
R13420 gnd.n2092 gnd.n2082 19.3944
R13421 gnd.n2098 gnd.n2082 19.3944
R13422 gnd.n2098 gnd.n2080 19.3944
R13423 gnd.n2102 gnd.n2080 19.3944
R13424 gnd.n2102 gnd.n2078 19.3944
R13425 gnd.n2108 gnd.n2078 19.3944
R13426 gnd.n2108 gnd.n2076 19.3944
R13427 gnd.n2112 gnd.n2076 19.3944
R13428 gnd.n2112 gnd.n2074 19.3944
R13429 gnd.n2118 gnd.n2074 19.3944
R13430 gnd.n2118 gnd.n2072 19.3944
R13431 gnd.n2125 gnd.n2072 19.3944
R13432 gnd.n2131 gnd.n2070 19.3944
R13433 gnd.n2131 gnd.n2068 19.3944
R13434 gnd.n2135 gnd.n2068 19.3944
R13435 gnd.n2135 gnd.n2066 19.3944
R13436 gnd.n2141 gnd.n2066 19.3944
R13437 gnd.n2141 gnd.n2064 19.3944
R13438 gnd.n2145 gnd.n2064 19.3944
R13439 gnd.n2145 gnd.n2062 19.3944
R13440 gnd.n2151 gnd.n2062 19.3944
R13441 gnd.n2151 gnd.n2060 19.3944
R13442 gnd.n2155 gnd.n2060 19.3944
R13443 gnd.n2155 gnd.n2058 19.3944
R13444 gnd.n2161 gnd.n2058 19.3944
R13445 gnd.n2161 gnd.n2056 19.3944
R13446 gnd.n2166 gnd.n2056 19.3944
R13447 gnd.n2166 gnd.n2054 19.3944
R13448 gnd.n5279 gnd.n2003 19.3944
R13449 gnd.n5291 gnd.n2003 19.3944
R13450 gnd.n5291 gnd.n2001 19.3944
R13451 gnd.n5295 gnd.n2001 19.3944
R13452 gnd.n5295 gnd.n1985 19.3944
R13453 gnd.n5307 gnd.n1985 19.3944
R13454 gnd.n5307 gnd.n1983 19.3944
R13455 gnd.n5311 gnd.n1983 19.3944
R13456 gnd.n5311 gnd.n1968 19.3944
R13457 gnd.n5323 gnd.n1968 19.3944
R13458 gnd.n5323 gnd.n1966 19.3944
R13459 gnd.n5336 gnd.n1966 19.3944
R13460 gnd.n5336 gnd.n5335 19.3944
R13461 gnd.n5335 gnd.n5334 19.3944
R13462 gnd.n5334 gnd.n5333 19.3944
R13463 gnd.n5333 gnd.n1927 19.3944
R13464 gnd.n5377 gnd.n1927 19.3944
R13465 gnd.n5377 gnd.n5376 19.3944
R13466 gnd.n5376 gnd.n5375 19.3944
R13467 gnd.n5375 gnd.n1937 19.3944
R13468 gnd.n1937 gnd.n1936 19.3944
R13469 gnd.n1936 gnd.n1853 19.3944
R13470 gnd.n5641 gnd.n1853 19.3944
R13471 gnd.n5641 gnd.n5640 19.3944
R13472 gnd.n5640 gnd.n5639 19.3944
R13473 gnd.n5639 gnd.n1857 19.3944
R13474 gnd.n5609 gnd.n1857 19.3944
R13475 gnd.n5612 gnd.n5609 19.3944
R13476 gnd.n5612 gnd.n1885 19.3944
R13477 gnd.n5616 gnd.n1885 19.3944
R13478 gnd.n5616 gnd.n1830 19.3944
R13479 gnd.n5654 gnd.n1830 19.3944
R13480 gnd.n5654 gnd.n1828 19.3944
R13481 gnd.n5658 gnd.n1828 19.3944
R13482 gnd.n5658 gnd.n1812 19.3944
R13483 gnd.n5670 gnd.n1812 19.3944
R13484 gnd.n5670 gnd.n1810 19.3944
R13485 gnd.n5674 gnd.n1810 19.3944
R13486 gnd.n5674 gnd.n1795 19.3944
R13487 gnd.n5686 gnd.n1795 19.3944
R13488 gnd.n5686 gnd.n1793 19.3944
R13489 gnd.n5690 gnd.n1793 19.3944
R13490 gnd.n5690 gnd.n1777 19.3944
R13491 gnd.n5702 gnd.n1777 19.3944
R13492 gnd.n5702 gnd.n1775 19.3944
R13493 gnd.n5711 gnd.n1775 19.3944
R13494 gnd.n5711 gnd.n5710 19.3944
R13495 gnd.n5710 gnd.n5709 19.3944
R13496 gnd.n5709 gnd.n1616 19.3944
R13497 gnd.n5902 gnd.n1616 19.3944
R13498 gnd.n5902 gnd.n5901 19.3944
R13499 gnd.n5901 gnd.n5900 19.3944
R13500 gnd.n5276 gnd.n5275 19.3944
R13501 gnd.n5275 gnd.n2017 19.3944
R13502 gnd.n5269 gnd.n2017 19.3944
R13503 gnd.n5269 gnd.n5268 19.3944
R13504 gnd.n5268 gnd.n5267 19.3944
R13505 gnd.n5267 gnd.n2023 19.3944
R13506 gnd.n5261 gnd.n2023 19.3944
R13507 gnd.n5261 gnd.n5260 19.3944
R13508 gnd.n5260 gnd.n5259 19.3944
R13509 gnd.n5259 gnd.n2029 19.3944
R13510 gnd.n5253 gnd.n2029 19.3944
R13511 gnd.n5253 gnd.n5252 19.3944
R13512 gnd.n5252 gnd.n5251 19.3944
R13513 gnd.n5251 gnd.n2035 19.3944
R13514 gnd.n5239 gnd.n5238 19.3944
R13515 gnd.n5238 gnd.n5236 19.3944
R13516 gnd.n5236 gnd.n5235 19.3944
R13517 gnd.n5235 gnd.n5233 19.3944
R13518 gnd.n5233 gnd.n5232 19.3944
R13519 gnd.n5232 gnd.n5230 19.3944
R13520 gnd.n5230 gnd.n5229 19.3944
R13521 gnd.n5229 gnd.n2046 19.3944
R13522 gnd.n2216 gnd.n2046 19.3944
R13523 gnd.n2216 gnd.n2215 19.3944
R13524 gnd.n2215 gnd.n2214 19.3944
R13525 gnd.n2214 gnd.n2198 19.3944
R13526 gnd.n2198 gnd.n1948 19.3944
R13527 gnd.n5350 gnd.n1948 19.3944
R13528 gnd.n5350 gnd.n1946 19.3944
R13529 gnd.n5360 gnd.n1946 19.3944
R13530 gnd.n5360 gnd.n5359 19.3944
R13531 gnd.n5359 gnd.n5358 19.3944
R13532 gnd.n5358 gnd.n1908 19.3944
R13533 gnd.n5390 gnd.n1908 19.3944
R13534 gnd.n5390 gnd.n1906 19.3944
R13535 gnd.n5395 gnd.n1906 19.3944
R13536 gnd.n5395 gnd.n1899 19.3944
R13537 gnd.n5407 gnd.n1899 19.3944
R13538 gnd.n5408 gnd.n5407 19.3944
R13539 gnd.n5408 gnd.n1897 19.3944
R13540 gnd.n5412 gnd.n1897 19.3944
R13541 gnd.n5415 gnd.n5412 19.3944
R13542 gnd.n5416 gnd.n5415 19.3944
R13543 gnd.n5416 gnd.n1894 19.3944
R13544 gnd.n5594 gnd.n1894 19.3944
R13545 gnd.n5594 gnd.n1895 19.3944
R13546 gnd.n5590 gnd.n1895 19.3944
R13547 gnd.n5590 gnd.n5589 19.3944
R13548 gnd.n5589 gnd.n5588 19.3944
R13549 gnd.n5588 gnd.n5422 19.3944
R13550 gnd.n5584 gnd.n5422 19.3944
R13551 gnd.n5584 gnd.n5583 19.3944
R13552 gnd.n5583 gnd.n5582 19.3944
R13553 gnd.n5582 gnd.n5426 19.3944
R13554 gnd.n5578 gnd.n5426 19.3944
R13555 gnd.n5578 gnd.n5577 19.3944
R13556 gnd.n5577 gnd.n5576 19.3944
R13557 gnd.n5576 gnd.n5430 19.3944
R13558 gnd.n5572 gnd.n5430 19.3944
R13559 gnd.n5572 gnd.n5571 19.3944
R13560 gnd.n5571 gnd.n1757 19.3944
R13561 gnd.n5723 gnd.n1757 19.3944
R13562 gnd.n5723 gnd.n1755 19.3944
R13563 gnd.n5727 gnd.n1755 19.3944
R13564 gnd.n5730 gnd.n5727 19.3944
R13565 gnd.n5731 gnd.n5730 19.3944
R13566 gnd.n2178 gnd.n2176 19.3944
R13567 gnd.n2178 gnd.n2049 19.3944
R13568 gnd.n2183 gnd.n2049 19.3944
R13569 gnd.n2184 gnd.n2183 19.3944
R13570 gnd.n2186 gnd.n2184 19.3944
R13571 gnd.n2186 gnd.n2047 19.3944
R13572 gnd.n5225 gnd.n2047 19.3944
R13573 gnd.n5225 gnd.n5224 19.3944
R13574 gnd.n5224 gnd.n5223 19.3944
R13575 gnd.n5223 gnd.n2192 19.3944
R13576 gnd.n2210 gnd.n2192 19.3944
R13577 gnd.n2210 gnd.n2209 19.3944
R13578 gnd.n2209 gnd.n2208 19.3944
R13579 gnd.n2208 gnd.n2205 19.3944
R13580 gnd.n2205 gnd.n1942 19.3944
R13581 gnd.n5364 gnd.n1942 19.3944
R13582 gnd.n5365 gnd.n5364 19.3944
R13583 gnd.n5365 gnd.n1940 19.3944
R13584 gnd.n5371 gnd.n1940 19.3944
R13585 gnd.n5371 gnd.n5370 19.3944
R13586 gnd.n5370 gnd.n1902 19.3944
R13587 gnd.n5399 gnd.n1902 19.3944
R13588 gnd.n5399 gnd.n1900 19.3944
R13589 gnd.n5403 gnd.n1900 19.3944
R13590 gnd.n5403 gnd.n1888 19.3944
R13591 gnd.n5605 gnd.n1888 19.3944
R13592 gnd.n5605 gnd.n5604 19.3944
R13593 gnd.n5604 gnd.n5601 19.3944
R13594 gnd.n5601 gnd.n5600 19.3944
R13595 gnd.n5600 gnd.n5599 19.3944
R13596 gnd.n5599 gnd.n5598 19.3944
R13597 gnd.n5598 gnd.n1893 19.3944
R13598 gnd.n5482 gnd.n1893 19.3944
R13599 gnd.n5483 gnd.n5482 19.3944
R13600 gnd.n5486 gnd.n5483 19.3944
R13601 gnd.n5486 gnd.n5476 19.3944
R13602 gnd.n5509 gnd.n5476 19.3944
R13603 gnd.n5509 gnd.n5508 19.3944
R13604 gnd.n5508 gnd.n5507 19.3944
R13605 gnd.n5507 gnd.n5504 19.3944
R13606 gnd.n5504 gnd.n5503 19.3944
R13607 gnd.n5503 gnd.n5500 19.3944
R13608 gnd.n5500 gnd.n5499 19.3944
R13609 gnd.n5499 gnd.n5432 19.3944
R13610 gnd.n5567 gnd.n5432 19.3944
R13611 gnd.n5567 gnd.n5566 19.3944
R13612 gnd.n5566 gnd.n5565 19.3944
R13613 gnd.n5565 gnd.n5562 19.3944
R13614 gnd.n5562 gnd.n5561 19.3944
R13615 gnd.n5561 gnd.n5439 19.3944
R13616 gnd.n5439 gnd.n1597 19.3944
R13617 gnd.n5960 gnd.n1597 19.3944
R13618 gnd.n5993 gnd.n1557 19.3944
R13619 gnd.n5993 gnd.n1564 19.3944
R13620 gnd.n1568 gnd.n1564 19.3944
R13621 gnd.n5986 gnd.n1568 19.3944
R13622 gnd.n5986 gnd.n5985 19.3944
R13623 gnd.n5985 gnd.n5984 19.3944
R13624 gnd.n5984 gnd.n1574 19.3944
R13625 gnd.n5979 gnd.n1574 19.3944
R13626 gnd.n5979 gnd.n5978 19.3944
R13627 gnd.n5978 gnd.n5977 19.3944
R13628 gnd.n5977 gnd.n1581 19.3944
R13629 gnd.n5972 gnd.n1581 19.3944
R13630 gnd.n5972 gnd.n5971 19.3944
R13631 gnd.n5971 gnd.n5970 19.3944
R13632 gnd.n5970 gnd.n1588 19.3944
R13633 gnd.n5965 gnd.n1588 19.3944
R13634 gnd.n5953 gnd.n5952 19.3944
R13635 gnd.n5952 gnd.n5910 19.3944
R13636 gnd.n5911 gnd.n5910 19.3944
R13637 gnd.n5945 gnd.n5911 19.3944
R13638 gnd.n5945 gnd.n5944 19.3944
R13639 gnd.n5944 gnd.n5943 19.3944
R13640 gnd.n5943 gnd.n5918 19.3944
R13641 gnd.n5938 gnd.n5918 19.3944
R13642 gnd.n5938 gnd.n5937 19.3944
R13643 gnd.n5937 gnd.n5936 19.3944
R13644 gnd.n5936 gnd.n5925 19.3944
R13645 gnd.n5931 gnd.n5925 19.3944
R13646 gnd.n5931 gnd.n1558 19.3944
R13647 gnd.n5283 gnd.n2009 19.3944
R13648 gnd.n5287 gnd.n2009 19.3944
R13649 gnd.n5287 gnd.n1994 19.3944
R13650 gnd.n5299 gnd.n1994 19.3944
R13651 gnd.n5299 gnd.n1992 19.3944
R13652 gnd.n5303 gnd.n1992 19.3944
R13653 gnd.n5303 gnd.n1976 19.3944
R13654 gnd.n5315 gnd.n1976 19.3944
R13655 gnd.n5315 gnd.n1974 19.3944
R13656 gnd.n5319 gnd.n1974 19.3944
R13657 gnd.n5319 gnd.n1958 19.3944
R13658 gnd.n5340 gnd.n1958 19.3944
R13659 gnd.n5340 gnd.n1956 19.3944
R13660 gnd.n5346 gnd.n1956 19.3944
R13661 gnd.n5346 gnd.n5345 19.3944
R13662 gnd.n5345 gnd.n1918 19.3944
R13663 gnd.n5381 gnd.n1918 19.3944
R13664 gnd.n5381 gnd.n1916 19.3944
R13665 gnd.n5385 gnd.n1916 19.3944
R13666 gnd.n5386 gnd.n5385 19.3944
R13667 gnd.n5386 gnd.n1844 19.3944
R13668 gnd.n5646 gnd.n5645 19.3944
R13669 gnd.n5635 gnd.n5634 19.3944
R13670 gnd.n1865 gnd.n1864 19.3944
R13671 gnd.n5621 gnd.n5620 19.3944
R13672 gnd.n1881 gnd.n1837 19.3944
R13673 gnd.n5650 gnd.n1837 19.3944
R13674 gnd.n5650 gnd.n1821 19.3944
R13675 gnd.n5662 gnd.n1821 19.3944
R13676 gnd.n5662 gnd.n1819 19.3944
R13677 gnd.n5666 gnd.n1819 19.3944
R13678 gnd.n5666 gnd.n1804 19.3944
R13679 gnd.n5678 gnd.n1804 19.3944
R13680 gnd.n5678 gnd.n1802 19.3944
R13681 gnd.n5682 gnd.n1802 19.3944
R13682 gnd.n5682 gnd.n1786 19.3944
R13683 gnd.n5694 gnd.n1786 19.3944
R13684 gnd.n5694 gnd.n1784 19.3944
R13685 gnd.n5698 gnd.n1784 19.3944
R13686 gnd.n5698 gnd.n1767 19.3944
R13687 gnd.n5715 gnd.n1767 19.3944
R13688 gnd.n5715 gnd.n1765 19.3944
R13689 gnd.n5719 gnd.n1765 19.3944
R13690 gnd.n5719 gnd.n1609 19.3944
R13691 gnd.n5906 gnd.n1609 19.3944
R13692 gnd.n5906 gnd.n1607 19.3944
R13693 gnd.n5956 gnd.n1607 19.3944
R13694 gnd.n3377 gnd.n2320 19.3944
R13695 gnd.n3381 gnd.n2320 19.3944
R13696 gnd.n3381 gnd.n2316 19.3944
R13697 gnd.n3387 gnd.n2316 19.3944
R13698 gnd.n3387 gnd.n2314 19.3944
R13699 gnd.n3391 gnd.n2314 19.3944
R13700 gnd.n3391 gnd.n2310 19.3944
R13701 gnd.n3397 gnd.n2310 19.3944
R13702 gnd.n3397 gnd.n2308 19.3944
R13703 gnd.n3401 gnd.n2308 19.3944
R13704 gnd.n3401 gnd.n2304 19.3944
R13705 gnd.n3407 gnd.n2304 19.3944
R13706 gnd.n3407 gnd.n2302 19.3944
R13707 gnd.n3411 gnd.n2302 19.3944
R13708 gnd.n3411 gnd.n2298 19.3944
R13709 gnd.n3417 gnd.n2298 19.3944
R13710 gnd.n3417 gnd.n2296 19.3944
R13711 gnd.n3421 gnd.n2296 19.3944
R13712 gnd.n3421 gnd.n2292 19.3944
R13713 gnd.n3427 gnd.n2292 19.3944
R13714 gnd.n3427 gnd.n2290 19.3944
R13715 gnd.n3431 gnd.n2290 19.3944
R13716 gnd.n3431 gnd.n2286 19.3944
R13717 gnd.n3437 gnd.n2286 19.3944
R13718 gnd.n3437 gnd.n2284 19.3944
R13719 gnd.n3441 gnd.n2284 19.3944
R13720 gnd.n3441 gnd.n2280 19.3944
R13721 gnd.n3447 gnd.n2280 19.3944
R13722 gnd.n3447 gnd.n2278 19.3944
R13723 gnd.n3451 gnd.n2278 19.3944
R13724 gnd.n3451 gnd.n2274 19.3944
R13725 gnd.n3457 gnd.n2274 19.3944
R13726 gnd.n3457 gnd.n2272 19.3944
R13727 gnd.n3461 gnd.n2272 19.3944
R13728 gnd.n3461 gnd.n2268 19.3944
R13729 gnd.n3467 gnd.n2268 19.3944
R13730 gnd.n3467 gnd.n2266 19.3944
R13731 gnd.n3471 gnd.n2266 19.3944
R13732 gnd.n3471 gnd.n2262 19.3944
R13733 gnd.n3477 gnd.n2262 19.3944
R13734 gnd.n3477 gnd.n2260 19.3944
R13735 gnd.n3481 gnd.n2260 19.3944
R13736 gnd.n3481 gnd.n2256 19.3944
R13737 gnd.n3487 gnd.n2256 19.3944
R13738 gnd.n3487 gnd.n2254 19.3944
R13739 gnd.n3491 gnd.n2254 19.3944
R13740 gnd.n3491 gnd.n2250 19.3944
R13741 gnd.n3497 gnd.n2250 19.3944
R13742 gnd.n3497 gnd.n2248 19.3944
R13743 gnd.n3501 gnd.n2248 19.3944
R13744 gnd.n3501 gnd.n2244 19.3944
R13745 gnd.n3507 gnd.n2244 19.3944
R13746 gnd.n3507 gnd.n2242 19.3944
R13747 gnd.n3511 gnd.n2242 19.3944
R13748 gnd.n3511 gnd.n2238 19.3944
R13749 gnd.n3517 gnd.n2238 19.3944
R13750 gnd.n3517 gnd.n2236 19.3944
R13751 gnd.n3521 gnd.n2236 19.3944
R13752 gnd.n3521 gnd.n2232 19.3944
R13753 gnd.n3527 gnd.n2232 19.3944
R13754 gnd.n3527 gnd.n2230 19.3944
R13755 gnd.n3531 gnd.n2230 19.3944
R13756 gnd.n3531 gnd.n2226 19.3944
R13757 gnd.n5163 gnd.n2226 19.3944
R13758 gnd.n5163 gnd.n2224 19.3944
R13759 gnd.n5167 gnd.n2224 19.3944
R13760 gnd.n5895 gnd.n5894 19.3944
R13761 gnd.n5894 gnd.n5893 19.3944
R13762 gnd.n5893 gnd.n1625 19.3944
R13763 gnd.n5889 gnd.n1625 19.3944
R13764 gnd.n5889 gnd.n5888 19.3944
R13765 gnd.n5888 gnd.n5887 19.3944
R13766 gnd.n5887 gnd.n1630 19.3944
R13767 gnd.n5883 gnd.n1630 19.3944
R13768 gnd.n5883 gnd.n5882 19.3944
R13769 gnd.n5882 gnd.n5881 19.3944
R13770 gnd.n5881 gnd.n5878 19.3944
R13771 gnd.n5878 gnd.n1421 19.3944
R13772 gnd.n6074 gnd.n1421 19.3944
R13773 gnd.n6074 gnd.n1418 19.3944
R13774 gnd.n6079 gnd.n1418 19.3944
R13775 gnd.n6079 gnd.n1419 19.3944
R13776 gnd.n1419 gnd.n1389 19.3944
R13777 gnd.n6154 gnd.n1389 19.3944
R13778 gnd.n6154 gnd.n1386 19.3944
R13779 gnd.n6159 gnd.n1386 19.3944
R13780 gnd.n6159 gnd.n1387 19.3944
R13781 gnd.n1387 gnd.n1357 19.3944
R13782 gnd.n6205 gnd.n1357 19.3944
R13783 gnd.n6205 gnd.n1354 19.3944
R13784 gnd.n6210 gnd.n1354 19.3944
R13785 gnd.n6210 gnd.n1355 19.3944
R13786 gnd.n1355 gnd.n1321 19.3944
R13787 gnd.n6271 gnd.n1321 19.3944
R13788 gnd.n6271 gnd.n1318 19.3944
R13789 gnd.n6279 gnd.n1318 19.3944
R13790 gnd.n6279 gnd.n1319 19.3944
R13791 gnd.n6275 gnd.n1319 19.3944
R13792 gnd.n6275 gnd.n1283 19.3944
R13793 gnd.n6334 gnd.n1283 19.3944
R13794 gnd.n6334 gnd.n1281 19.3944
R13795 gnd.n6338 gnd.n1281 19.3944
R13796 gnd.n6338 gnd.n1253 19.3944
R13797 gnd.n6403 gnd.n1253 19.3944
R13798 gnd.n6403 gnd.n1251 19.3944
R13799 gnd.n6407 gnd.n1251 19.3944
R13800 gnd.n6407 gnd.n1225 19.3944
R13801 gnd.n6439 gnd.n1225 19.3944
R13802 gnd.n6439 gnd.n1223 19.3944
R13803 gnd.n6443 gnd.n1223 19.3944
R13804 gnd.n6443 gnd.n1197 19.3944
R13805 gnd.n6476 gnd.n1197 19.3944
R13806 gnd.n6476 gnd.n1194 19.3944
R13807 gnd.n6484 gnd.n1194 19.3944
R13808 gnd.n6484 gnd.n1195 19.3944
R13809 gnd.n6480 gnd.n1195 19.3944
R13810 gnd.n6480 gnd.n1097 19.3944
R13811 gnd.n6624 gnd.n1097 19.3944
R13812 gnd.n6624 gnd.n1094 19.3944
R13813 gnd.n6629 gnd.n1094 19.3944
R13814 gnd.n6629 gnd.n1095 19.3944
R13815 gnd.n1095 gnd.n1072 19.3944
R13816 gnd.n6654 gnd.n1072 19.3944
R13817 gnd.n6654 gnd.n1069 19.3944
R13818 gnd.n6659 gnd.n1069 19.3944
R13819 gnd.n6659 gnd.n1070 19.3944
R13820 gnd.n1070 gnd.n1047 19.3944
R13821 gnd.n6696 gnd.n1047 19.3944
R13822 gnd.n6696 gnd.n1044 19.3944
R13823 gnd.n6701 gnd.n1044 19.3944
R13824 gnd.n6701 gnd.n1045 19.3944
R13825 gnd.n1034 gnd.n1031 19.3944
R13826 gnd.n1034 gnd.n994 19.3944
R13827 gnd.n6709 gnd.n994 19.3944
R13828 gnd.n7006 gnd.n7005 19.3944
R13829 gnd.n7005 gnd.n797 19.3944
R13830 gnd.n6998 gnd.n797 19.3944
R13831 gnd.n6998 gnd.n6997 19.3944
R13832 gnd.n6997 gnd.n805 19.3944
R13833 gnd.n6990 gnd.n805 19.3944
R13834 gnd.n6990 gnd.n6989 19.3944
R13835 gnd.n6989 gnd.n813 19.3944
R13836 gnd.n6982 gnd.n813 19.3944
R13837 gnd.n6982 gnd.n6981 19.3944
R13838 gnd.n6981 gnd.n821 19.3944
R13839 gnd.n6974 gnd.n821 19.3944
R13840 gnd.n6974 gnd.n6973 19.3944
R13841 gnd.n6973 gnd.n829 19.3944
R13842 gnd.n1007 gnd.n829 19.3944
R13843 gnd.n1010 gnd.n1007 19.3944
R13844 gnd.n1010 gnd.n1002 19.3944
R13845 gnd.n1021 gnd.n1002 19.3944
R13846 gnd.n1022 gnd.n1021 19.3944
R13847 gnd.n1025 gnd.n1022 19.3944
R13848 gnd.n1025 gnd.n998 19.3944
R13849 gnd.n1029 gnd.n998 19.3944
R13850 gnd.n4430 gnd.n3897 19.328
R13851 gnd.n4502 gnd.t22 18.9947
R13852 gnd.n6938 gnd.n6937 18.4247
R13853 gnd.n5997 gnd.n1558 18.4247
R13854 gnd.n4483 gnd.t10 18.3283
R13855 gnd.n7244 gnd.n7239 18.2308
R13856 gnd.n6970 gnd.n825 18.2308
R13857 gnd.n5770 gnd.n1737 18.2308
R13858 gnd.n5245 gnd.n2035 18.2308
R13859 gnd.n3830 gnd.t17 17.6618
R13860 gnd.n5810 gnd.n5809 17.3286
R13861 gnd.n6711 gnd.n973 17.3286
R13862 gnd.t197 gnd.n3924 16.9954
R13863 gnd.n3787 gnd.t225 16.9954
R13864 gnd.n5819 gnd.n1668 16.6621
R13865 gnd.n5819 gnd.n5818 16.6621
R13866 gnd.n5818 gnd.n1669 16.6621
R13867 gnd.n1669 gnd.n1663 16.6621
R13868 gnd.n5827 gnd.n1663 16.6621
R13869 gnd.n5830 gnd.n5829 16.6621
R13870 gnd.n5829 gnd.n1656 16.6621
R13871 gnd.n5839 gnd.n1656 16.6621
R13872 gnd.n5839 gnd.n5838 16.6621
R13873 gnd.n5838 gnd.n1657 16.6621
R13874 gnd.n1657 gnd.n1650 16.6621
R13875 gnd.n5847 gnd.n1650 16.6621
R13876 gnd.n5850 gnd.n5847 16.6621
R13877 gnd.n5850 gnd.n5849 16.6621
R13878 gnd.n5849 gnd.n1642 16.6621
R13879 gnd.n5861 gnd.n1642 16.6621
R13880 gnd.n5861 gnd.n5860 16.6621
R13881 gnd.n5860 gnd.n1643 16.6621
R13882 gnd.n5875 gnd.n1634 16.6621
R13883 gnd.n5875 gnd.n5874 16.6621
R13884 gnd.n5874 gnd.n1432 16.6621
R13885 gnd.n6061 gnd.n1432 16.6621
R13886 gnd.n6061 gnd.n6060 16.6621
R13887 gnd.n6072 gnd.n1423 16.6621
R13888 gnd.n6081 gnd.n1415 16.6621
R13889 gnd.n6143 gnd.n1399 16.6621
R13890 gnd.n6106 gnd.n1362 16.6621
R13891 gnd.n6106 gnd.n1348 16.6621
R13892 gnd.n6187 gnd.n1342 16.6621
R13893 gnd.n6269 gnd.n1323 16.6621
R13894 gnd.n6282 gnd.n6281 16.6621
R13895 gnd.n6303 gnd.n1307 16.6621
R13896 gnd.n6297 gnd.n1300 16.6621
R13897 gnd.n1293 gnd.n1292 16.6621
R13898 gnd.n6390 gnd.n6389 16.6621
R13899 gnd.n6383 gnd.n6382 16.6621
R13900 gnd.n6427 gnd.n1234 16.6621
R13901 gnd.n6427 gnd.n6426 16.6621
R13902 gnd.n6446 gnd.n1206 16.6621
R13903 gnd.n1217 gnd.n1202 16.6621
R13904 gnd.n6355 gnd.n6354 16.6621
R13905 gnd.n6611 gnd.n1109 16.6621
R13906 gnd.n6622 gnd.n1099 16.6621
R13907 gnd.n6622 gnd.n6621 16.6621
R13908 gnd.n1101 gnd.n1090 16.6621
R13909 gnd.n6631 gnd.n1090 16.6621
R13910 gnd.n6631 gnd.n1091 16.6621
R13911 gnd.n1091 gnd.n1083 16.6621
R13912 gnd.n6641 gnd.n1083 16.6621
R13913 gnd.n6640 gnd.n1074 16.6621
R13914 gnd.n6652 gnd.n1074 16.6621
R13915 gnd.n6652 gnd.n6651 16.6621
R13916 gnd.n6651 gnd.n1076 16.6621
R13917 gnd.n1076 gnd.n1065 16.6621
R13918 gnd.n6661 gnd.n1065 16.6621
R13919 gnd.n6661 gnd.n1066 16.6621
R13920 gnd.n1066 gnd.n1058 16.6621
R13921 gnd.n6672 gnd.n1058 16.6621
R13922 gnd.n6672 gnd.n6671 16.6621
R13923 gnd.n6671 gnd.n1049 16.6621
R13924 gnd.n6694 gnd.n1049 16.6621
R13925 gnd.n6694 gnd.n6693 16.6621
R13926 gnd.n1051 gnd.n1040 16.6621
R13927 gnd.n6703 gnd.n1040 16.6621
R13928 gnd.n6703 gnd.n1041 16.6621
R13929 gnd.n6685 gnd.n1041 16.6621
R13930 gnd.n6686 gnd.n6685 16.6621
R13931 gnd.n4042 gnd.t197 16.3289
R13932 gnd.n5124 gnd.t128 16.3289
R13933 gnd.n5015 gnd.t142 16.3289
R13934 gnd.t204 gnd.n5827 16.3289
R13935 gnd.t211 gnd.n1051 16.3289
R13936 gnd.n5809 gnd.n1675 15.9957
R13937 gnd.n1496 gnd.n1495 15.9957
R13938 gnd.n6304 gnd.n1304 15.9957
R13939 gnd.n6332 gnd.n1285 15.9957
R13940 gnd.n6486 gnd.n1191 15.9957
R13941 gnd.n6610 gnd.n1111 15.9957
R13942 gnd.n6712 gnd.n6711 15.9957
R13943 gnd.n4277 gnd.n4275 15.6674
R13944 gnd.n4314 gnd.n4312 15.6674
R13945 gnd.n4138 gnd.n4136 15.6674
R13946 gnd.n4175 gnd.n4173 15.6674
R13947 gnd.n4207 gnd.n4205 15.6674
R13948 gnd.n4244 gnd.n4242 15.6674
R13949 gnd.n443 gnd.n441 15.6674
R13950 gnd.n406 gnd.n404 15.6674
R13951 gnd.n304 gnd.n302 15.6674
R13952 gnd.n267 gnd.n265 15.6674
R13953 gnd.n373 gnd.n371 15.6674
R13954 gnd.n336 gnd.n334 15.6674
R13955 gnd.n4980 gnd.n4978 15.6674
R13956 gnd.n4948 gnd.n4946 15.6674
R13957 gnd.n4916 gnd.n4914 15.6674
R13958 gnd.n4885 gnd.n4883 15.6674
R13959 gnd.n4853 gnd.n4851 15.6674
R13960 gnd.n4821 gnd.n4819 15.6674
R13961 gnd.n4789 gnd.n4787 15.6674
R13962 gnd.n4758 gnd.n4756 15.6674
R13963 gnd.n107 gnd.n105 15.6674
R13964 gnd.n75 gnd.n73 15.6674
R13965 gnd.n43 gnd.n41 15.6674
R13966 gnd.n12 gnd.n10 15.6674
R13967 gnd.n234 gnd.n232 15.6674
R13968 gnd.n202 gnd.n200 15.6674
R13969 gnd.n170 gnd.n168 15.6674
R13970 gnd.n139 gnd.n137 15.6674
R13971 gnd.n6196 gnd.n1366 15.3292
R13972 gnd.n6220 gnd.n1343 15.3292
R13973 gnd.n1273 gnd.n1258 15.3292
R13974 gnd.n6420 gnd.n6419 15.3292
R13975 gnd.n1119 gnd.n1118 15.0827
R13976 gnd.n1474 gnd.n1469 15.0481
R13977 gnd.n1129 gnd.n1128 15.0481
R13978 gnd.n5145 gnd.t27 14.996
R13979 gnd.n5137 gnd.t11 14.996
R13980 gnd.n6060 gnd.n6059 14.996
R13981 gnd.n6072 gnd.t179 14.6627
R13982 gnd.n1393 gnd.n1380 14.6627
R13983 gnd.t31 gnd.n3836 14.3295
R13984 gnd.n4431 gnd.n4430 13.9963
R13985 gnd.n6152 gnd.t215 13.9963
R13986 gnd.n6163 gnd.n6162 13.9963
R13987 gnd.n6171 gnd.t117 13.9963
R13988 gnd.n6268 gnd.n1326 13.9963
R13989 gnd.n6391 gnd.n1263 13.9963
R13990 gnd.n6467 gnd.n6466 13.9963
R13991 gnd.n5159 gnd.n3535 13.663
R13992 gnd.n4399 gnd.n4395 13.5763
R13993 gnd.n5088 gnd.n3647 13.5763
R13994 gnd.n6904 gnd.n902 13.5763
R13995 gnd.n7292 gnd.n7291 13.5763
R13996 gnd.n2054 gnd.n2053 13.5763
R13997 gnd.n5965 gnd.n5964 13.5763
R13998 gnd.n6170 gnd.n1376 13.3298
R13999 gnd.t12 gnd.n6194 13.3298
R14000 gnd.n6228 gnd.n6227 13.3298
R14001 gnd.n6401 gnd.n1255 13.3298
R14002 gnd.t223 gnd.n1244 13.3298
R14003 gnd.n6447 gnd.n6445 13.3298
R14004 gnd.n1485 gnd.n1466 13.1884
R14005 gnd.n1480 gnd.n1479 13.1884
R14006 gnd.n1479 gnd.n1478 13.1884
R14007 gnd.n1122 gnd.n1117 13.1884
R14008 gnd.n1123 gnd.n1122 13.1884
R14009 gnd.n1481 gnd.n1468 13.146
R14010 gnd.n1477 gnd.n1468 13.146
R14011 gnd.n1121 gnd.n1120 13.146
R14012 gnd.n1121 gnd.n1116 13.146
R14013 gnd.n4278 gnd.n4274 12.8005
R14014 gnd.n4315 gnd.n4311 12.8005
R14015 gnd.n4139 gnd.n4135 12.8005
R14016 gnd.n4176 gnd.n4172 12.8005
R14017 gnd.n4208 gnd.n4204 12.8005
R14018 gnd.n4245 gnd.n4241 12.8005
R14019 gnd.n444 gnd.n440 12.8005
R14020 gnd.n407 gnd.n403 12.8005
R14021 gnd.n305 gnd.n301 12.8005
R14022 gnd.n268 gnd.n264 12.8005
R14023 gnd.n374 gnd.n370 12.8005
R14024 gnd.n337 gnd.n333 12.8005
R14025 gnd.n6056 gnd.n1487 12.8005
R14026 gnd.n6606 gnd.n6605 12.8005
R14027 gnd.n4981 gnd.n4977 12.8005
R14028 gnd.n4949 gnd.n4945 12.8005
R14029 gnd.n4917 gnd.n4913 12.8005
R14030 gnd.n4886 gnd.n4882 12.8005
R14031 gnd.n4854 gnd.n4850 12.8005
R14032 gnd.n4822 gnd.n4818 12.8005
R14033 gnd.n4790 gnd.n4786 12.8005
R14034 gnd.n4759 gnd.n4755 12.8005
R14035 gnd.n108 gnd.n104 12.8005
R14036 gnd.n76 gnd.n72 12.8005
R14037 gnd.n44 gnd.n40 12.8005
R14038 gnd.n13 gnd.n9 12.8005
R14039 gnd.n235 gnd.n231 12.8005
R14040 gnd.n203 gnd.n199 12.8005
R14041 gnd.n171 gnd.n167 12.8005
R14042 gnd.n140 gnd.n136 12.8005
R14043 gnd.n5544 gnd.n1567 12.6633
R14044 gnd.n6124 gnd.n1391 12.6633
R14045 gnd.n6261 gnd.n6260 12.6633
R14046 gnd.n1294 gnd.n1288 12.6633
R14047 gnd.t208 gnd.n6473 12.6633
R14048 gnd.n6460 gnd.n6459 12.6633
R14049 gnd.n6964 gnd.n833 12.6633
R14050 gnd.n4402 gnd.n4399 12.4126
R14051 gnd.n5091 gnd.n5088 12.4126
R14052 gnd.n6900 gnd.n902 12.4126
R14053 gnd.n7291 gnd.n570 12.4126
R14054 gnd.n2173 gnd.n2053 12.4126
R14055 gnd.n5964 gnd.n1593 12.4126
R14056 gnd.n5297 gnd.n1999 12.3301
R14057 gnd.n7275 gnd.n583 12.3301
R14058 gnd.n4282 gnd.n4281 12.0247
R14059 gnd.n4319 gnd.n4318 12.0247
R14060 gnd.n4143 gnd.n4142 12.0247
R14061 gnd.n4180 gnd.n4179 12.0247
R14062 gnd.n4212 gnd.n4211 12.0247
R14063 gnd.n4249 gnd.n4248 12.0247
R14064 gnd.n448 gnd.n447 12.0247
R14065 gnd.n411 gnd.n410 12.0247
R14066 gnd.n309 gnd.n308 12.0247
R14067 gnd.n272 gnd.n271 12.0247
R14068 gnd.n378 gnd.n377 12.0247
R14069 gnd.n341 gnd.n340 12.0247
R14070 gnd.n4985 gnd.n4984 12.0247
R14071 gnd.n4953 gnd.n4952 12.0247
R14072 gnd.n4921 gnd.n4920 12.0247
R14073 gnd.n4890 gnd.n4889 12.0247
R14074 gnd.n4858 gnd.n4857 12.0247
R14075 gnd.n4826 gnd.n4825 12.0247
R14076 gnd.n4794 gnd.n4793 12.0247
R14077 gnd.n4763 gnd.n4762 12.0247
R14078 gnd.n112 gnd.n111 12.0247
R14079 gnd.n80 gnd.n79 12.0247
R14080 gnd.n48 gnd.n47 12.0247
R14081 gnd.n17 gnd.n16 12.0247
R14082 gnd.n239 gnd.n238 12.0247
R14083 gnd.n207 gnd.n206 12.0247
R14084 gnd.n175 gnd.n174 12.0247
R14085 gnd.n144 gnd.n143 12.0247
R14086 gnd.n6203 gnd.n1359 11.9969
R14087 gnd.n6212 gnd.n1351 11.9969
R14088 gnd.n6409 gnd.n1248 11.9969
R14089 gnd.n6437 gnd.n6436 11.9969
R14090 gnd.n4503 gnd.t31 11.6636
R14091 gnd.n5676 gnd.t58 11.6636
R14092 gnd.n7071 gnd.t49 11.6636
R14093 gnd.n6133 gnd.n6132 11.3304
R14094 gnd.n6132 gnd.n6131 11.3304
R14095 gnd.n1306 gnd.n1299 11.3304
R14096 gnd.n6310 gnd.n1299 11.3304
R14097 gnd.n6495 gnd.n6494 11.3304
R14098 gnd.n4285 gnd.n4272 11.249
R14099 gnd.n4322 gnd.n4309 11.249
R14100 gnd.n4146 gnd.n4133 11.249
R14101 gnd.n4183 gnd.n4170 11.249
R14102 gnd.n4215 gnd.n4202 11.249
R14103 gnd.n4252 gnd.n4239 11.249
R14104 gnd.n451 gnd.n438 11.249
R14105 gnd.n414 gnd.n401 11.249
R14106 gnd.n312 gnd.n299 11.249
R14107 gnd.n275 gnd.n262 11.249
R14108 gnd.n381 gnd.n368 11.249
R14109 gnd.n344 gnd.n331 11.249
R14110 gnd.n4988 gnd.n4975 11.249
R14111 gnd.n4956 gnd.n4943 11.249
R14112 gnd.n4924 gnd.n4911 11.249
R14113 gnd.n4893 gnd.n4880 11.249
R14114 gnd.n4861 gnd.n4848 11.249
R14115 gnd.n4829 gnd.n4816 11.249
R14116 gnd.n4797 gnd.n4784 11.249
R14117 gnd.n4766 gnd.n4753 11.249
R14118 gnd.n115 gnd.n102 11.249
R14119 gnd.n83 gnd.n70 11.249
R14120 gnd.n51 gnd.n38 11.249
R14121 gnd.n20 gnd.n7 11.249
R14122 gnd.n242 gnd.n229 11.249
R14123 gnd.n210 gnd.n197 11.249
R14124 gnd.n178 gnd.n165 11.249
R14125 gnd.n147 gnd.n134 11.249
R14126 gnd.n3912 gnd.t29 10.9972
R14127 gnd.t27 gnd.n5144 10.9972
R14128 gnd.n4731 gnd.t11 10.9972
R14129 gnd.n5405 gnd.t45 10.9972
R14130 gnd.n1643 gnd.t0 10.9972
R14131 gnd.t218 gnd.n6640 10.9972
R14132 gnd.n7128 gnd.t74 10.9972
R14133 gnd.n6203 gnd.n6202 10.6639
R14134 gnd.n6437 gnd.n1227 10.6639
R14135 gnd.n6549 gnd.n6548 10.6151
R14136 gnd.n6548 gnd.n6547 10.6151
R14137 gnd.n6542 gnd.n1163 10.6151
R14138 gnd.n6542 gnd.n6541 10.6151
R14139 gnd.n6541 gnd.n6540 10.6151
R14140 gnd.n6540 gnd.n1165 10.6151
R14141 gnd.n6535 gnd.n1165 10.6151
R14142 gnd.n6535 gnd.n6534 10.6151
R14143 gnd.n6534 gnd.n6533 10.6151
R14144 gnd.n6533 gnd.n1168 10.6151
R14145 gnd.n6528 gnd.n1168 10.6151
R14146 gnd.n6528 gnd.n6527 10.6151
R14147 gnd.n6527 gnd.n6526 10.6151
R14148 gnd.n6526 gnd.n1171 10.6151
R14149 gnd.n6521 gnd.n1171 10.6151
R14150 gnd.n6521 gnd.n6520 10.6151
R14151 gnd.n6520 gnd.n6519 10.6151
R14152 gnd.n6519 gnd.n1174 10.6151
R14153 gnd.n6514 gnd.n1174 10.6151
R14154 gnd.n6514 gnd.n6513 10.6151
R14155 gnd.n6513 gnd.n6512 10.6151
R14156 gnd.n6512 gnd.n1177 10.6151
R14157 gnd.n6507 gnd.n1177 10.6151
R14158 gnd.n6507 gnd.n6506 10.6151
R14159 gnd.n6506 gnd.n6505 10.6151
R14160 gnd.n6505 gnd.n1180 10.6151
R14161 gnd.n6500 gnd.n1180 10.6151
R14162 gnd.n1494 gnd.n1493 10.6151
R14163 gnd.n1494 gnd.n1406 10.6151
R14164 gnd.n6129 gnd.n1406 10.6151
R14165 gnd.n6129 gnd.n6128 10.6151
R14166 gnd.n6128 gnd.n6127 10.6151
R14167 gnd.n6127 gnd.n1407 10.6151
R14168 gnd.n6092 gnd.n1407 10.6151
R14169 gnd.n6093 gnd.n6092 10.6151
R14170 gnd.n6094 gnd.n6093 10.6151
R14171 gnd.n6095 gnd.n6094 10.6151
R14172 gnd.n6098 gnd.n6095 10.6151
R14173 gnd.n6099 gnd.n6098 10.6151
R14174 gnd.n6101 gnd.n6099 10.6151
R14175 gnd.n6102 gnd.n6101 10.6151
R14176 gnd.n6104 gnd.n6102 10.6151
R14177 gnd.n6104 gnd.n6103 10.6151
R14178 gnd.n6103 gnd.n1340 10.6151
R14179 gnd.n6222 gnd.n1340 10.6151
R14180 gnd.n6223 gnd.n6222 10.6151
R14181 gnd.n6225 gnd.n6223 10.6151
R14182 gnd.n6225 gnd.n6224 10.6151
R14183 gnd.n6224 gnd.n1332 10.6151
R14184 gnd.n6253 gnd.n1332 10.6151
R14185 gnd.n6254 gnd.n6253 10.6151
R14186 gnd.n6257 gnd.n6254 10.6151
R14187 gnd.n6257 gnd.n6256 10.6151
R14188 gnd.n6256 gnd.n6255 10.6151
R14189 gnd.n6255 gnd.n1297 10.6151
R14190 gnd.n6313 gnd.n1297 10.6151
R14191 gnd.n6314 gnd.n6313 10.6151
R14192 gnd.n6315 gnd.n6314 10.6151
R14193 gnd.n6323 gnd.n6315 10.6151
R14194 gnd.n6323 gnd.n6322 10.6151
R14195 gnd.n6322 gnd.n6321 10.6151
R14196 gnd.n6321 gnd.n6320 10.6151
R14197 gnd.n6320 gnd.n6318 10.6151
R14198 gnd.n6318 gnd.n6317 10.6151
R14199 gnd.n6317 gnd.n1246 10.6151
R14200 gnd.n6412 gnd.n1246 10.6151
R14201 gnd.n6413 gnd.n6412 10.6151
R14202 gnd.n6415 gnd.n6413 10.6151
R14203 gnd.n6416 gnd.n6415 10.6151
R14204 gnd.n6417 gnd.n6416 10.6151
R14205 gnd.n6417 gnd.n1218 10.6151
R14206 gnd.n6449 gnd.n1218 10.6151
R14207 gnd.n6450 gnd.n6449 10.6151
R14208 gnd.n6452 gnd.n6450 10.6151
R14209 gnd.n6453 gnd.n6452 10.6151
R14210 gnd.n6457 gnd.n6453 10.6151
R14211 gnd.n6457 gnd.n6456 10.6151
R14212 gnd.n6456 gnd.n6455 10.6151
R14213 gnd.n6455 gnd.n1184 10.6151
R14214 gnd.n6497 gnd.n1184 10.6151
R14215 gnd.n6498 gnd.n6497 10.6151
R14216 gnd.n6499 gnd.n6498 10.6151
R14217 gnd.n1556 gnd.n1553 10.6151
R14218 gnd.n1553 gnd.n1552 10.6151
R14219 gnd.n1549 gnd.n1548 10.6151
R14220 gnd.n1548 gnd.n1545 10.6151
R14221 gnd.n1545 gnd.n1544 10.6151
R14222 gnd.n1544 gnd.n1541 10.6151
R14223 gnd.n1541 gnd.n1540 10.6151
R14224 gnd.n1540 gnd.n1537 10.6151
R14225 gnd.n1537 gnd.n1536 10.6151
R14226 gnd.n1536 gnd.n1533 10.6151
R14227 gnd.n1533 gnd.n1532 10.6151
R14228 gnd.n1532 gnd.n1529 10.6151
R14229 gnd.n1529 gnd.n1528 10.6151
R14230 gnd.n1528 gnd.n1525 10.6151
R14231 gnd.n1525 gnd.n1524 10.6151
R14232 gnd.n1524 gnd.n1521 10.6151
R14233 gnd.n1521 gnd.n1520 10.6151
R14234 gnd.n1520 gnd.n1517 10.6151
R14235 gnd.n1517 gnd.n1516 10.6151
R14236 gnd.n1516 gnd.n1513 10.6151
R14237 gnd.n1513 gnd.n1512 10.6151
R14238 gnd.n1512 gnd.n1509 10.6151
R14239 gnd.n1509 gnd.n1508 10.6151
R14240 gnd.n1508 gnd.n1505 10.6151
R14241 gnd.n1505 gnd.n1504 10.6151
R14242 gnd.n1504 gnd.n1501 10.6151
R14243 gnd.n1501 gnd.n1500 10.6151
R14244 gnd.n6056 gnd.n6055 10.6151
R14245 gnd.n6055 gnd.n6054 10.6151
R14246 gnd.n6054 gnd.n6053 10.6151
R14247 gnd.n6053 gnd.n6051 10.6151
R14248 gnd.n6051 gnd.n6048 10.6151
R14249 gnd.n6048 gnd.n6047 10.6151
R14250 gnd.n6047 gnd.n6044 10.6151
R14251 gnd.n6044 gnd.n6043 10.6151
R14252 gnd.n6043 gnd.n6040 10.6151
R14253 gnd.n6040 gnd.n6039 10.6151
R14254 gnd.n6039 gnd.n6036 10.6151
R14255 gnd.n6036 gnd.n6035 10.6151
R14256 gnd.n6035 gnd.n6032 10.6151
R14257 gnd.n6032 gnd.n6031 10.6151
R14258 gnd.n6031 gnd.n6028 10.6151
R14259 gnd.n6028 gnd.n6027 10.6151
R14260 gnd.n6027 gnd.n6024 10.6151
R14261 gnd.n6024 gnd.n6023 10.6151
R14262 gnd.n6023 gnd.n6020 10.6151
R14263 gnd.n6020 gnd.n6019 10.6151
R14264 gnd.n6019 gnd.n6016 10.6151
R14265 gnd.n6016 gnd.n6015 10.6151
R14266 gnd.n6015 gnd.n6012 10.6151
R14267 gnd.n6012 gnd.n6011 10.6151
R14268 gnd.n6011 gnd.n6008 10.6151
R14269 gnd.n6006 gnd.n6003 10.6151
R14270 gnd.n6003 gnd.n6002 10.6151
R14271 gnd.n6605 gnd.n1134 10.6151
R14272 gnd.n6600 gnd.n1134 10.6151
R14273 gnd.n6600 gnd.n6599 10.6151
R14274 gnd.n6599 gnd.n6598 10.6151
R14275 gnd.n6598 gnd.n1136 10.6151
R14276 gnd.n6593 gnd.n1136 10.6151
R14277 gnd.n6593 gnd.n6592 10.6151
R14278 gnd.n6592 gnd.n6591 10.6151
R14279 gnd.n6591 gnd.n1139 10.6151
R14280 gnd.n6586 gnd.n1139 10.6151
R14281 gnd.n6586 gnd.n6585 10.6151
R14282 gnd.n6585 gnd.n6584 10.6151
R14283 gnd.n6584 gnd.n1142 10.6151
R14284 gnd.n6579 gnd.n1142 10.6151
R14285 gnd.n6579 gnd.n6578 10.6151
R14286 gnd.n6578 gnd.n6577 10.6151
R14287 gnd.n6577 gnd.n1145 10.6151
R14288 gnd.n6572 gnd.n1145 10.6151
R14289 gnd.n6572 gnd.n6571 10.6151
R14290 gnd.n6571 gnd.n6570 10.6151
R14291 gnd.n6570 gnd.n1148 10.6151
R14292 gnd.n6565 gnd.n1148 10.6151
R14293 gnd.n6565 gnd.n6564 10.6151
R14294 gnd.n6564 gnd.n6563 10.6151
R14295 gnd.n6563 gnd.n1151 10.6151
R14296 gnd.n6558 gnd.n6557 10.6151
R14297 gnd.n6557 gnd.n6556 10.6151
R14298 gnd.n1486 gnd.n1403 10.6151
R14299 gnd.n6135 gnd.n1403 10.6151
R14300 gnd.n6136 gnd.n6135 10.6151
R14301 gnd.n6140 gnd.n6136 10.6151
R14302 gnd.n6140 gnd.n6139 10.6151
R14303 gnd.n6139 gnd.n6138 10.6151
R14304 gnd.n6138 gnd.n1378 10.6151
R14305 gnd.n6166 gnd.n1378 10.6151
R14306 gnd.n6167 gnd.n6166 10.6151
R14307 gnd.n6168 gnd.n6167 10.6151
R14308 gnd.n6168 gnd.n1364 10.6151
R14309 gnd.n6198 gnd.n1364 10.6151
R14310 gnd.n6199 gnd.n6198 10.6151
R14311 gnd.n6200 gnd.n6199 10.6151
R14312 gnd.n6200 gnd.n1346 10.6151
R14313 gnd.n6215 gnd.n1346 10.6151
R14314 gnd.n6216 gnd.n6215 10.6151
R14315 gnd.n6218 gnd.n6216 10.6151
R14316 gnd.n6218 gnd.n6217 10.6151
R14317 gnd.n6217 gnd.n1329 10.6151
R14318 gnd.n6266 gnd.n1329 10.6151
R14319 gnd.n6266 gnd.n6265 10.6151
R14320 gnd.n6265 gnd.n6264 10.6151
R14321 gnd.n6264 gnd.n1330 10.6151
R14322 gnd.n1330 gnd.n1302 10.6151
R14323 gnd.n6306 gnd.n1302 10.6151
R14324 gnd.n6307 gnd.n6306 10.6151
R14325 gnd.n6308 gnd.n6307 10.6151
R14326 gnd.n6308 gnd.n1291 10.6151
R14327 gnd.n6329 gnd.n1291 10.6151
R14328 gnd.n6329 gnd.n6328 10.6151
R14329 gnd.n6328 gnd.n6327 10.6151
R14330 gnd.n6327 gnd.n1261 10.6151
R14331 gnd.n6393 gnd.n1261 10.6151
R14332 gnd.n6394 gnd.n6393 10.6151
R14333 gnd.n6398 gnd.n6394 10.6151
R14334 gnd.n6398 gnd.n6397 10.6151
R14335 gnd.n6397 gnd.n6396 10.6151
R14336 gnd.n6396 gnd.n1232 10.6151
R14337 gnd.n6429 gnd.n1232 10.6151
R14338 gnd.n6430 gnd.n6429 10.6151
R14339 gnd.n6434 gnd.n6430 10.6151
R14340 gnd.n6434 gnd.n6433 10.6151
R14341 gnd.n6433 gnd.n6432 10.6151
R14342 gnd.n6432 gnd.n1204 10.6151
R14343 gnd.n6469 gnd.n1204 10.6151
R14344 gnd.n6470 gnd.n6469 10.6151
R14345 gnd.n6471 gnd.n6470 10.6151
R14346 gnd.n6471 gnd.n1187 10.6151
R14347 gnd.n6489 gnd.n1187 10.6151
R14348 gnd.n6490 gnd.n6489 10.6151
R14349 gnd.n6491 gnd.n6490 10.6151
R14350 gnd.n6491 gnd.n1114 10.6151
R14351 gnd.n6608 gnd.n1114 10.6151
R14352 gnd.n6608 gnd.n6607 10.6151
R14353 gnd.n4286 gnd.n4270 10.4732
R14354 gnd.n4323 gnd.n4307 10.4732
R14355 gnd.n4147 gnd.n4131 10.4732
R14356 gnd.n4184 gnd.n4168 10.4732
R14357 gnd.n4216 gnd.n4200 10.4732
R14358 gnd.n4253 gnd.n4237 10.4732
R14359 gnd.n452 gnd.n436 10.4732
R14360 gnd.n415 gnd.n399 10.4732
R14361 gnd.n313 gnd.n297 10.4732
R14362 gnd.n276 gnd.n260 10.4732
R14363 gnd.n382 gnd.n366 10.4732
R14364 gnd.n345 gnd.n329 10.4732
R14365 gnd.n4989 gnd.n4973 10.4732
R14366 gnd.n4957 gnd.n4941 10.4732
R14367 gnd.n4925 gnd.n4909 10.4732
R14368 gnd.n4894 gnd.n4878 10.4732
R14369 gnd.n4862 gnd.n4846 10.4732
R14370 gnd.n4830 gnd.n4814 10.4732
R14371 gnd.n4798 gnd.n4782 10.4732
R14372 gnd.n4767 gnd.n4751 10.4732
R14373 gnd.n116 gnd.n100 10.4732
R14374 gnd.n84 gnd.n68 10.4732
R14375 gnd.n52 gnd.n36 10.4732
R14376 gnd.n21 gnd.n5 10.4732
R14377 gnd.n243 gnd.n227 10.4732
R14378 gnd.n211 gnd.n195 10.4732
R14379 gnd.n179 gnd.n163 10.4732
R14380 gnd.n148 gnd.n132 10.4732
R14381 gnd.t222 gnd.n5158 10.3307
R14382 gnd.n5321 gnd.t65 10.3307
R14383 gnd.t56 gnd.n1952 10.3307
R14384 gnd.t62 gnd.n626 10.3307
R14385 gnd.n7183 gnd.t87 10.3307
R14386 gnd.n6071 gnd.n1425 9.99747
R14387 gnd.n6260 gnd.n6259 9.99747
R14388 gnd.n6331 gnd.n1288 9.99747
R14389 gnd.n1182 gnd.n1099 9.99747
R14390 gnd.t194 gnd.n1101 9.99747
R14391 gnd.n4290 gnd.n4289 9.69747
R14392 gnd.n4327 gnd.n4326 9.69747
R14393 gnd.n4151 gnd.n4150 9.69747
R14394 gnd.n4188 gnd.n4187 9.69747
R14395 gnd.n4220 gnd.n4219 9.69747
R14396 gnd.n4257 gnd.n4256 9.69747
R14397 gnd.n456 gnd.n455 9.69747
R14398 gnd.n419 gnd.n418 9.69747
R14399 gnd.n317 gnd.n316 9.69747
R14400 gnd.n280 gnd.n279 9.69747
R14401 gnd.n386 gnd.n385 9.69747
R14402 gnd.n349 gnd.n348 9.69747
R14403 gnd.n4993 gnd.n4992 9.69747
R14404 gnd.n4961 gnd.n4960 9.69747
R14405 gnd.n4929 gnd.n4928 9.69747
R14406 gnd.n4898 gnd.n4897 9.69747
R14407 gnd.n4866 gnd.n4865 9.69747
R14408 gnd.n4834 gnd.n4833 9.69747
R14409 gnd.n4802 gnd.n4801 9.69747
R14410 gnd.n4771 gnd.n4770 9.69747
R14411 gnd.n120 gnd.n119 9.69747
R14412 gnd.n88 gnd.n87 9.69747
R14413 gnd.n56 gnd.n55 9.69747
R14414 gnd.n25 gnd.n24 9.69747
R14415 gnd.n247 gnd.n246 9.69747
R14416 gnd.n215 gnd.n214 9.69747
R14417 gnd.n183 gnd.n182 9.69747
R14418 gnd.n152 gnd.n151 9.69747
R14419 gnd.t24 gnd.n3732 9.66424
R14420 gnd.n5022 gnd.t128 9.66424
R14421 gnd.n5123 gnd.t142 9.66424
R14422 gnd.n5624 gnd.t60 9.66424
R14423 gnd.t51 gnd.n682 9.66424
R14424 gnd.n5898 gnd.n1619 9.45599
R14425 gnd.n7011 gnd.n7010 9.45599
R14426 gnd.n4296 gnd.n4295 9.45567
R14427 gnd.n4333 gnd.n4332 9.45567
R14428 gnd.n4157 gnd.n4156 9.45567
R14429 gnd.n4194 gnd.n4193 9.45567
R14430 gnd.n4226 gnd.n4225 9.45567
R14431 gnd.n4263 gnd.n4262 9.45567
R14432 gnd.n462 gnd.n461 9.45567
R14433 gnd.n425 gnd.n424 9.45567
R14434 gnd.n323 gnd.n322 9.45567
R14435 gnd.n286 gnd.n285 9.45567
R14436 gnd.n392 gnd.n391 9.45567
R14437 gnd.n355 gnd.n354 9.45567
R14438 gnd.n4999 gnd.n4998 9.45567
R14439 gnd.n4967 gnd.n4966 9.45567
R14440 gnd.n4935 gnd.n4934 9.45567
R14441 gnd.n4904 gnd.n4903 9.45567
R14442 gnd.n4872 gnd.n4871 9.45567
R14443 gnd.n4840 gnd.n4839 9.45567
R14444 gnd.n4808 gnd.n4807 9.45567
R14445 gnd.n4777 gnd.n4776 9.45567
R14446 gnd.n126 gnd.n125 9.45567
R14447 gnd.n94 gnd.n93 9.45567
R14448 gnd.n62 gnd.n61 9.45567
R14449 gnd.n31 gnd.n30 9.45567
R14450 gnd.n253 gnd.n252 9.45567
R14451 gnd.n221 gnd.n220 9.45567
R14452 gnd.n189 gnd.n188 9.45567
R14453 gnd.n158 gnd.n157 9.45567
R14454 gnd.t39 gnd.t24 9.33101
R14455 gnd.n6096 gnd.n1376 9.33101
R14456 gnd.n6228 gnd.n1338 9.33101
R14457 gnd.n6401 gnd.n6400 9.33101
R14458 gnd.n6445 gnd.n1220 9.33101
R14459 gnd.n4295 gnd.n4294 9.3005
R14460 gnd.n4268 gnd.n4267 9.3005
R14461 gnd.n4289 gnd.n4288 9.3005
R14462 gnd.n4287 gnd.n4286 9.3005
R14463 gnd.n4272 gnd.n4271 9.3005
R14464 gnd.n4281 gnd.n4280 9.3005
R14465 gnd.n4279 gnd.n4278 9.3005
R14466 gnd.n4332 gnd.n4331 9.3005
R14467 gnd.n4305 gnd.n4304 9.3005
R14468 gnd.n4326 gnd.n4325 9.3005
R14469 gnd.n4324 gnd.n4323 9.3005
R14470 gnd.n4309 gnd.n4308 9.3005
R14471 gnd.n4318 gnd.n4317 9.3005
R14472 gnd.n4316 gnd.n4315 9.3005
R14473 gnd.n4156 gnd.n4155 9.3005
R14474 gnd.n4129 gnd.n4128 9.3005
R14475 gnd.n4150 gnd.n4149 9.3005
R14476 gnd.n4148 gnd.n4147 9.3005
R14477 gnd.n4133 gnd.n4132 9.3005
R14478 gnd.n4142 gnd.n4141 9.3005
R14479 gnd.n4140 gnd.n4139 9.3005
R14480 gnd.n4193 gnd.n4192 9.3005
R14481 gnd.n4166 gnd.n4165 9.3005
R14482 gnd.n4187 gnd.n4186 9.3005
R14483 gnd.n4185 gnd.n4184 9.3005
R14484 gnd.n4170 gnd.n4169 9.3005
R14485 gnd.n4179 gnd.n4178 9.3005
R14486 gnd.n4177 gnd.n4176 9.3005
R14487 gnd.n4225 gnd.n4224 9.3005
R14488 gnd.n4198 gnd.n4197 9.3005
R14489 gnd.n4219 gnd.n4218 9.3005
R14490 gnd.n4217 gnd.n4216 9.3005
R14491 gnd.n4202 gnd.n4201 9.3005
R14492 gnd.n4211 gnd.n4210 9.3005
R14493 gnd.n4209 gnd.n4208 9.3005
R14494 gnd.n4262 gnd.n4261 9.3005
R14495 gnd.n4235 gnd.n4234 9.3005
R14496 gnd.n4256 gnd.n4255 9.3005
R14497 gnd.n4254 gnd.n4253 9.3005
R14498 gnd.n4239 gnd.n4238 9.3005
R14499 gnd.n4248 gnd.n4247 9.3005
R14500 gnd.n4246 gnd.n4245 9.3005
R14501 gnd.n461 gnd.n460 9.3005
R14502 gnd.n434 gnd.n433 9.3005
R14503 gnd.n455 gnd.n454 9.3005
R14504 gnd.n453 gnd.n452 9.3005
R14505 gnd.n438 gnd.n437 9.3005
R14506 gnd.n447 gnd.n446 9.3005
R14507 gnd.n445 gnd.n444 9.3005
R14508 gnd.n424 gnd.n423 9.3005
R14509 gnd.n397 gnd.n396 9.3005
R14510 gnd.n418 gnd.n417 9.3005
R14511 gnd.n416 gnd.n415 9.3005
R14512 gnd.n401 gnd.n400 9.3005
R14513 gnd.n410 gnd.n409 9.3005
R14514 gnd.n408 gnd.n407 9.3005
R14515 gnd.n322 gnd.n321 9.3005
R14516 gnd.n295 gnd.n294 9.3005
R14517 gnd.n316 gnd.n315 9.3005
R14518 gnd.n314 gnd.n313 9.3005
R14519 gnd.n299 gnd.n298 9.3005
R14520 gnd.n308 gnd.n307 9.3005
R14521 gnd.n306 gnd.n305 9.3005
R14522 gnd.n285 gnd.n284 9.3005
R14523 gnd.n258 gnd.n257 9.3005
R14524 gnd.n279 gnd.n278 9.3005
R14525 gnd.n277 gnd.n276 9.3005
R14526 gnd.n262 gnd.n261 9.3005
R14527 gnd.n271 gnd.n270 9.3005
R14528 gnd.n269 gnd.n268 9.3005
R14529 gnd.n391 gnd.n390 9.3005
R14530 gnd.n364 gnd.n363 9.3005
R14531 gnd.n385 gnd.n384 9.3005
R14532 gnd.n383 gnd.n382 9.3005
R14533 gnd.n368 gnd.n367 9.3005
R14534 gnd.n377 gnd.n376 9.3005
R14535 gnd.n375 gnd.n374 9.3005
R14536 gnd.n354 gnd.n353 9.3005
R14537 gnd.n327 gnd.n326 9.3005
R14538 gnd.n348 gnd.n347 9.3005
R14539 gnd.n346 gnd.n345 9.3005
R14540 gnd.n331 gnd.n330 9.3005
R14541 gnd.n340 gnd.n339 9.3005
R14542 gnd.n338 gnd.n337 9.3005
R14543 gnd.n4998 gnd.n4997 9.3005
R14544 gnd.n4971 gnd.n4970 9.3005
R14545 gnd.n4992 gnd.n4991 9.3005
R14546 gnd.n4990 gnd.n4989 9.3005
R14547 gnd.n4975 gnd.n4974 9.3005
R14548 gnd.n4984 gnd.n4983 9.3005
R14549 gnd.n4982 gnd.n4981 9.3005
R14550 gnd.n4966 gnd.n4965 9.3005
R14551 gnd.n4939 gnd.n4938 9.3005
R14552 gnd.n4960 gnd.n4959 9.3005
R14553 gnd.n4958 gnd.n4957 9.3005
R14554 gnd.n4943 gnd.n4942 9.3005
R14555 gnd.n4952 gnd.n4951 9.3005
R14556 gnd.n4950 gnd.n4949 9.3005
R14557 gnd.n4934 gnd.n4933 9.3005
R14558 gnd.n4907 gnd.n4906 9.3005
R14559 gnd.n4928 gnd.n4927 9.3005
R14560 gnd.n4926 gnd.n4925 9.3005
R14561 gnd.n4911 gnd.n4910 9.3005
R14562 gnd.n4920 gnd.n4919 9.3005
R14563 gnd.n4918 gnd.n4917 9.3005
R14564 gnd.n4903 gnd.n4902 9.3005
R14565 gnd.n4876 gnd.n4875 9.3005
R14566 gnd.n4897 gnd.n4896 9.3005
R14567 gnd.n4895 gnd.n4894 9.3005
R14568 gnd.n4880 gnd.n4879 9.3005
R14569 gnd.n4889 gnd.n4888 9.3005
R14570 gnd.n4887 gnd.n4886 9.3005
R14571 gnd.n4871 gnd.n4870 9.3005
R14572 gnd.n4844 gnd.n4843 9.3005
R14573 gnd.n4865 gnd.n4864 9.3005
R14574 gnd.n4863 gnd.n4862 9.3005
R14575 gnd.n4848 gnd.n4847 9.3005
R14576 gnd.n4857 gnd.n4856 9.3005
R14577 gnd.n4855 gnd.n4854 9.3005
R14578 gnd.n4839 gnd.n4838 9.3005
R14579 gnd.n4812 gnd.n4811 9.3005
R14580 gnd.n4833 gnd.n4832 9.3005
R14581 gnd.n4831 gnd.n4830 9.3005
R14582 gnd.n4816 gnd.n4815 9.3005
R14583 gnd.n4825 gnd.n4824 9.3005
R14584 gnd.n4823 gnd.n4822 9.3005
R14585 gnd.n4807 gnd.n4806 9.3005
R14586 gnd.n4780 gnd.n4779 9.3005
R14587 gnd.n4801 gnd.n4800 9.3005
R14588 gnd.n4799 gnd.n4798 9.3005
R14589 gnd.n4784 gnd.n4783 9.3005
R14590 gnd.n4793 gnd.n4792 9.3005
R14591 gnd.n4791 gnd.n4790 9.3005
R14592 gnd.n4776 gnd.n4775 9.3005
R14593 gnd.n4749 gnd.n4748 9.3005
R14594 gnd.n4770 gnd.n4769 9.3005
R14595 gnd.n4768 gnd.n4767 9.3005
R14596 gnd.n4753 gnd.n4752 9.3005
R14597 gnd.n4762 gnd.n4761 9.3005
R14598 gnd.n4760 gnd.n4759 9.3005
R14599 gnd.n3632 gnd.n3629 9.3005
R14600 gnd.n5113 gnd.n3633 9.3005
R14601 gnd.n5112 gnd.n3634 9.3005
R14602 gnd.n5111 gnd.n3635 9.3005
R14603 gnd.n5108 gnd.n3636 9.3005
R14604 gnd.n5107 gnd.n3637 9.3005
R14605 gnd.n5104 gnd.n3638 9.3005
R14606 gnd.n5103 gnd.n3639 9.3005
R14607 gnd.n5100 gnd.n3640 9.3005
R14608 gnd.n5099 gnd.n3641 9.3005
R14609 gnd.n5096 gnd.n3642 9.3005
R14610 gnd.n5095 gnd.n3643 9.3005
R14611 gnd.n5092 gnd.n3644 9.3005
R14612 gnd.n5091 gnd.n3645 9.3005
R14613 gnd.n5088 gnd.n5087 9.3005
R14614 gnd.n5086 gnd.n3647 9.3005
R14615 gnd.n3631 gnd.n3630 9.3005
R14616 gnd.n4455 gnd.n4454 9.3005
R14617 gnd.n4456 gnd.n3883 9.3005
R14618 gnd.n4460 gnd.n4457 9.3005
R14619 gnd.n4459 gnd.n4458 9.3005
R14620 gnd.n3860 gnd.n3859 9.3005
R14621 gnd.n4486 gnd.n4485 9.3005
R14622 gnd.n4487 gnd.n3858 9.3005
R14623 gnd.n4491 gnd.n4488 9.3005
R14624 gnd.n4490 gnd.n4489 9.3005
R14625 gnd.n3834 gnd.n3833 9.3005
R14626 gnd.n4517 gnd.n4516 9.3005
R14627 gnd.n4518 gnd.n3832 9.3005
R14628 gnd.n4522 gnd.n4519 9.3005
R14629 gnd.n4521 gnd.n4520 9.3005
R14630 gnd.n3808 gnd.n3807 9.3005
R14631 gnd.n4548 gnd.n4547 9.3005
R14632 gnd.n4549 gnd.n3806 9.3005
R14633 gnd.n4553 gnd.n4550 9.3005
R14634 gnd.n4552 gnd.n4551 9.3005
R14635 gnd.n3782 gnd.n3781 9.3005
R14636 gnd.n4579 gnd.n4578 9.3005
R14637 gnd.n4580 gnd.n3780 9.3005
R14638 gnd.n4584 gnd.n4581 9.3005
R14639 gnd.n4583 gnd.n4582 9.3005
R14640 gnd.n3757 gnd.n3756 9.3005
R14641 gnd.n4610 gnd.n4609 9.3005
R14642 gnd.n4611 gnd.n3755 9.3005
R14643 gnd.n4615 gnd.n4612 9.3005
R14644 gnd.n4614 gnd.n4613 9.3005
R14645 gnd.n3730 gnd.n3729 9.3005
R14646 gnd.n4640 gnd.n4639 9.3005
R14647 gnd.n4641 gnd.n3728 9.3005
R14648 gnd.n4643 gnd.n4642 9.3005
R14649 gnd.n3708 gnd.n3707 9.3005
R14650 gnd.n4682 gnd.n4681 9.3005
R14651 gnd.n4683 gnd.n3706 9.3005
R14652 gnd.n4691 gnd.n4684 9.3005
R14653 gnd.n4690 gnd.n4685 9.3005
R14654 gnd.n4689 gnd.n4687 9.3005
R14655 gnd.n4686 gnd.n3551 9.3005
R14656 gnd.n5149 gnd.n3552 9.3005
R14657 gnd.n5148 gnd.n3553 9.3005
R14658 gnd.n5147 gnd.n3554 9.3005
R14659 gnd.n3574 gnd.n3555 9.3005
R14660 gnd.n3575 gnd.n3573 9.3005
R14661 gnd.n5135 gnd.n3576 9.3005
R14662 gnd.n5134 gnd.n3577 9.3005
R14663 gnd.n5133 gnd.n3578 9.3005
R14664 gnd.n3598 gnd.n3579 9.3005
R14665 gnd.n3599 gnd.n3597 9.3005
R14666 gnd.n5121 gnd.n3600 9.3005
R14667 gnd.n5120 gnd.n3601 9.3005
R14668 gnd.n5119 gnd.n3602 9.3005
R14669 gnd.n3885 gnd.n3884 9.3005
R14670 gnd.n4399 gnd.n4398 9.3005
R14671 gnd.n4402 gnd.n4394 9.3005
R14672 gnd.n4403 gnd.n4393 9.3005
R14673 gnd.n4406 gnd.n4392 9.3005
R14674 gnd.n4407 gnd.n4391 9.3005
R14675 gnd.n4410 gnd.n4390 9.3005
R14676 gnd.n4411 gnd.n4389 9.3005
R14677 gnd.n4414 gnd.n4388 9.3005
R14678 gnd.n4415 gnd.n4387 9.3005
R14679 gnd.n4418 gnd.n4386 9.3005
R14680 gnd.n4419 gnd.n4385 9.3005
R14681 gnd.n4422 gnd.n4384 9.3005
R14682 gnd.n4424 gnd.n4383 9.3005
R14683 gnd.n4425 gnd.n4382 9.3005
R14684 gnd.n4426 gnd.n4381 9.3005
R14685 gnd.n4427 gnd.n4380 9.3005
R14686 gnd.n4395 gnd.n3901 9.3005
R14687 gnd.n4445 gnd.n4444 9.3005
R14688 gnd.n4446 gnd.n3878 9.3005
R14689 gnd.n4465 gnd.n4464 9.3005
R14690 gnd.n4467 gnd.n3870 9.3005
R14691 gnd.n4474 gnd.n3871 9.3005
R14692 gnd.n4476 gnd.n4475 9.3005
R14693 gnd.n4477 gnd.n3851 9.3005
R14694 gnd.n4496 gnd.n4495 9.3005
R14695 gnd.n4498 gnd.n3844 9.3005
R14696 gnd.n4505 gnd.n3845 9.3005
R14697 gnd.n4507 gnd.n4506 9.3005
R14698 gnd.n4508 gnd.n3825 9.3005
R14699 gnd.n4527 gnd.n4526 9.3005
R14700 gnd.n4529 gnd.n3818 9.3005
R14701 gnd.n4536 gnd.n3819 9.3005
R14702 gnd.n4538 gnd.n4537 9.3005
R14703 gnd.n4539 gnd.n3800 9.3005
R14704 gnd.n4558 gnd.n4557 9.3005
R14705 gnd.n4560 gnd.n3792 9.3005
R14706 gnd.n4567 gnd.n3793 9.3005
R14707 gnd.n4569 gnd.n4568 9.3005
R14708 gnd.n4570 gnd.n3775 9.3005
R14709 gnd.n4589 gnd.n4588 9.3005
R14710 gnd.n4591 gnd.n3767 9.3005
R14711 gnd.n4598 gnd.n3768 9.3005
R14712 gnd.n4600 gnd.n4599 9.3005
R14713 gnd.n4601 gnd.n3750 9.3005
R14714 gnd.n4620 gnd.n4619 9.3005
R14715 gnd.n4622 gnd.n3741 9.3005
R14716 gnd.n4629 gnd.n3743 9.3005
R14717 gnd.n4630 gnd.n3738 9.3005
R14718 gnd.n4632 gnd.n4631 9.3005
R14719 gnd.n3739 gnd.n3724 9.3005
R14720 gnd.n4648 gnd.n3722 9.3005
R14721 gnd.n4652 gnd.n4651 9.3005
R14722 gnd.n4650 gnd.n3698 9.3005
R14723 gnd.n4698 gnd.n3697 9.3005
R14724 gnd.n4701 gnd.n4700 9.3005
R14725 gnd.n3694 gnd.n3693 9.3005
R14726 gnd.n4705 gnd.n3695 9.3005
R14727 gnd.n4707 gnd.n4706 9.3005
R14728 gnd.n4713 gnd.n4709 9.3005
R14729 gnd.n4712 gnd.n4711 9.3005
R14730 gnd.n3688 gnd.n3687 9.3005
R14731 gnd.n4741 gnd.n3689 9.3005
R14732 gnd.n4743 gnd.n4742 9.3005
R14733 gnd.n4745 gnd.n3686 9.3005
R14734 gnd.n5004 gnd.n5003 9.3005
R14735 gnd.n5006 gnd.n5005 9.3005
R14736 gnd.n5020 gnd.n5007 9.3005
R14737 gnd.n5019 gnd.n5008 9.3005
R14738 gnd.n5018 gnd.n5013 9.3005
R14739 gnd.n5014 gnd.n3650 9.3005
R14740 gnd.n4443 gnd.n3895 9.3005
R14741 gnd.n5082 gnd.n3651 9.3005
R14742 gnd.n5081 gnd.n3653 9.3005
R14743 gnd.n5078 gnd.n3654 9.3005
R14744 gnd.n5077 gnd.n3655 9.3005
R14745 gnd.n5074 gnd.n3656 9.3005
R14746 gnd.n5073 gnd.n3657 9.3005
R14747 gnd.n5070 gnd.n3658 9.3005
R14748 gnd.n5069 gnd.n3659 9.3005
R14749 gnd.n5066 gnd.n3660 9.3005
R14750 gnd.n5065 gnd.n3661 9.3005
R14751 gnd.n5062 gnd.n3662 9.3005
R14752 gnd.n5061 gnd.n3663 9.3005
R14753 gnd.n5058 gnd.n3664 9.3005
R14754 gnd.n5057 gnd.n3665 9.3005
R14755 gnd.n5054 gnd.n3666 9.3005
R14756 gnd.n5053 gnd.n3667 9.3005
R14757 gnd.n5050 gnd.n3668 9.3005
R14758 gnd.n5049 gnd.n3669 9.3005
R14759 gnd.n5046 gnd.n3670 9.3005
R14760 gnd.n5045 gnd.n3671 9.3005
R14761 gnd.n5042 gnd.n3672 9.3005
R14762 gnd.n5041 gnd.n3673 9.3005
R14763 gnd.n5038 gnd.n3677 9.3005
R14764 gnd.n5037 gnd.n3678 9.3005
R14765 gnd.n5034 gnd.n3679 9.3005
R14766 gnd.n5033 gnd.n3680 9.3005
R14767 gnd.n5084 gnd.n5083 9.3005
R14768 gnd.n4112 gnd.n4091 9.3005
R14769 gnd.n4111 gnd.n4093 9.3005
R14770 gnd.n4109 gnd.n4094 9.3005
R14771 gnd.n4108 gnd.n4095 9.3005
R14772 gnd.n4104 gnd.n4096 9.3005
R14773 gnd.n4103 gnd.n4097 9.3005
R14774 gnd.n4102 gnd.n4098 9.3005
R14775 gnd.n4100 gnd.n4099 9.3005
R14776 gnd.n3715 gnd.n3714 9.3005
R14777 gnd.n4660 gnd.n4659 9.3005
R14778 gnd.n4661 gnd.n3713 9.3005
R14779 gnd.n4676 gnd.n4662 9.3005
R14780 gnd.n4675 gnd.n4663 9.3005
R14781 gnd.n4674 gnd.n4664 9.3005
R14782 gnd.n4672 gnd.n4665 9.3005
R14783 gnd.n4671 gnd.n4666 9.3005
R14784 gnd.n4668 gnd.n4667 9.3005
R14785 gnd.n3692 gnd.n3691 9.3005
R14786 gnd.n4720 gnd.n4719 9.3005
R14787 gnd.n4721 gnd.n3690 9.3005
R14788 gnd.n4735 gnd.n4722 9.3005
R14789 gnd.n4734 gnd.n4723 9.3005
R14790 gnd.n4733 gnd.n4724 9.3005
R14791 gnd.n4727 gnd.n4726 9.3005
R14792 gnd.n4725 gnd.n3684 9.3005
R14793 gnd.n5025 gnd.n3683 9.3005
R14794 gnd.n5027 gnd.n5026 9.3005
R14795 gnd.n5028 gnd.n3682 9.3005
R14796 gnd.n5030 gnd.n5029 9.3005
R14797 gnd.n4038 gnd.n3932 9.3005
R14798 gnd.n4040 gnd.n4039 9.3005
R14799 gnd.n3922 gnd.n3921 9.3005
R14800 gnd.n4053 gnd.n4052 9.3005
R14801 gnd.n4054 gnd.n3920 9.3005
R14802 gnd.n4056 gnd.n4055 9.3005
R14803 gnd.n3909 gnd.n3908 9.3005
R14804 gnd.n4069 gnd.n4068 9.3005
R14805 gnd.n4070 gnd.n3907 9.3005
R14806 gnd.n4369 gnd.n4071 9.3005
R14807 gnd.n4368 gnd.n4072 9.3005
R14808 gnd.n4367 gnd.n4073 9.3005
R14809 gnd.n4366 gnd.n4074 9.3005
R14810 gnd.n4364 gnd.n4075 9.3005
R14811 gnd.n4363 gnd.n4076 9.3005
R14812 gnd.n4359 gnd.n4077 9.3005
R14813 gnd.n4358 gnd.n4078 9.3005
R14814 gnd.n4357 gnd.n4079 9.3005
R14815 gnd.n4355 gnd.n4080 9.3005
R14816 gnd.n4354 gnd.n4081 9.3005
R14817 gnd.n4351 gnd.n4082 9.3005
R14818 gnd.n4350 gnd.n4083 9.3005
R14819 gnd.n4349 gnd.n4084 9.3005
R14820 gnd.n4347 gnd.n4085 9.3005
R14821 gnd.n4346 gnd.n4086 9.3005
R14822 gnd.n4343 gnd.n4087 9.3005
R14823 gnd.n4342 gnd.n4088 9.3005
R14824 gnd.n4341 gnd.n4089 9.3005
R14825 gnd.n4037 gnd.n4036 9.3005
R14826 gnd.n3977 gnd.n3976 9.3005
R14827 gnd.n3982 gnd.n3974 9.3005
R14828 gnd.n3983 gnd.n3973 9.3005
R14829 gnd.n3985 gnd.n3970 9.3005
R14830 gnd.n3969 gnd.n3967 9.3005
R14831 gnd.n3991 gnd.n3966 9.3005
R14832 gnd.n3992 gnd.n3965 9.3005
R14833 gnd.n3993 gnd.n3964 9.3005
R14834 gnd.n3963 gnd.n3961 9.3005
R14835 gnd.n3999 gnd.n3960 9.3005
R14836 gnd.n4000 gnd.n3959 9.3005
R14837 gnd.n4001 gnd.n3958 9.3005
R14838 gnd.n3957 gnd.n3955 9.3005
R14839 gnd.n4007 gnd.n3954 9.3005
R14840 gnd.n4008 gnd.n3953 9.3005
R14841 gnd.n4009 gnd.n3952 9.3005
R14842 gnd.n3951 gnd.n3949 9.3005
R14843 gnd.n4015 gnd.n3948 9.3005
R14844 gnd.n4016 gnd.n3947 9.3005
R14845 gnd.n4017 gnd.n3946 9.3005
R14846 gnd.n3945 gnd.n3943 9.3005
R14847 gnd.n4022 gnd.n3942 9.3005
R14848 gnd.n4023 gnd.n3941 9.3005
R14849 gnd.n3940 gnd.n3938 9.3005
R14850 gnd.n4028 gnd.n3937 9.3005
R14851 gnd.n4030 gnd.n4029 9.3005
R14852 gnd.n3975 gnd.n3933 9.3005
R14853 gnd.n3928 gnd.n3927 9.3005
R14854 gnd.n4045 gnd.n4044 9.3005
R14855 gnd.n4046 gnd.n3926 9.3005
R14856 gnd.n4048 gnd.n4047 9.3005
R14857 gnd.n3916 gnd.n3915 9.3005
R14858 gnd.n4061 gnd.n4060 9.3005
R14859 gnd.n4062 gnd.n3914 9.3005
R14860 gnd.n4064 gnd.n4063 9.3005
R14861 gnd.n3903 gnd.n3902 9.3005
R14862 gnd.n4434 gnd.n4433 9.3005
R14863 gnd.n4436 gnd.n3900 9.3005
R14864 gnd.n4438 gnd.n4437 9.3005
R14865 gnd.n3894 gnd.n3893 9.3005
R14866 gnd.n4449 gnd.n4447 9.3005
R14867 gnd.n4448 gnd.n3877 9.3005
R14868 gnd.n4466 gnd.n3876 9.3005
R14869 gnd.n4469 gnd.n4468 9.3005
R14870 gnd.n3869 gnd.n3868 9.3005
R14871 gnd.n4480 gnd.n4478 9.3005
R14872 gnd.n4479 gnd.n3850 9.3005
R14873 gnd.n4497 gnd.n3849 9.3005
R14874 gnd.n4500 gnd.n4499 9.3005
R14875 gnd.n3843 gnd.n3842 9.3005
R14876 gnd.n4511 gnd.n4509 9.3005
R14877 gnd.n4510 gnd.n3824 9.3005
R14878 gnd.n4528 gnd.n3823 9.3005
R14879 gnd.n4531 gnd.n4530 9.3005
R14880 gnd.n3817 gnd.n3816 9.3005
R14881 gnd.n4542 gnd.n4540 9.3005
R14882 gnd.n4541 gnd.n3799 9.3005
R14883 gnd.n4559 gnd.n3798 9.3005
R14884 gnd.n4562 gnd.n4561 9.3005
R14885 gnd.n3791 gnd.n3790 9.3005
R14886 gnd.n4573 gnd.n4571 9.3005
R14887 gnd.n4572 gnd.n3774 9.3005
R14888 gnd.n4590 gnd.n3773 9.3005
R14889 gnd.n4593 gnd.n4592 9.3005
R14890 gnd.n3766 gnd.n3765 9.3005
R14891 gnd.n4604 gnd.n4602 9.3005
R14892 gnd.n4603 gnd.n3749 9.3005
R14893 gnd.n4621 gnd.n3748 9.3005
R14894 gnd.n4624 gnd.n4623 9.3005
R14895 gnd.n3742 gnd.n3737 9.3005
R14896 gnd.n4634 gnd.n4633 9.3005
R14897 gnd.n3740 gnd.n3720 9.3005
R14898 gnd.n4655 gnd.n3721 9.3005
R14899 gnd.n4654 gnd.n4653 9.3005
R14900 gnd.n3723 gnd.n3699 9.3005
R14901 gnd.n4697 gnd.n4696 9.3005
R14902 gnd.n4699 gnd.n3540 9.3005
R14903 gnd.n5156 gnd.n3541 9.3005
R14904 gnd.n5155 gnd.n3542 9.3005
R14905 gnd.n5154 gnd.n3543 9.3005
R14906 gnd.n4708 gnd.n3544 9.3005
R14907 gnd.n4710 gnd.n3562 9.3005
R14908 gnd.n5142 gnd.n3563 9.3005
R14909 gnd.n5141 gnd.n3564 9.3005
R14910 gnd.n5140 gnd.n3565 9.3005
R14911 gnd.n4744 gnd.n3566 9.3005
R14912 gnd.n4746 gnd.n3587 9.3005
R14913 gnd.n5128 gnd.n3588 9.3005
R14914 gnd.n5127 gnd.n3589 9.3005
R14915 gnd.n5126 gnd.n3590 9.3005
R14916 gnd.n5009 gnd.n3591 9.3005
R14917 gnd.n5012 gnd.n5011 9.3005
R14918 gnd.n4032 gnd.n4031 9.3005
R14919 gnd.n2325 gnd.n2321 9.3005
R14920 gnd.n3371 gnd.n2326 9.3005
R14921 gnd.n3370 gnd.n2327 9.3005
R14922 gnd.n3369 gnd.n2328 9.3005
R14923 gnd.n2333 gnd.n2329 9.3005
R14924 gnd.n3363 gnd.n2334 9.3005
R14925 gnd.n3362 gnd.n2335 9.3005
R14926 gnd.n3361 gnd.n2336 9.3005
R14927 gnd.n2341 gnd.n2337 9.3005
R14928 gnd.n3355 gnd.n2342 9.3005
R14929 gnd.n3354 gnd.n2343 9.3005
R14930 gnd.n3353 gnd.n2344 9.3005
R14931 gnd.n2349 gnd.n2345 9.3005
R14932 gnd.n3347 gnd.n2350 9.3005
R14933 gnd.n3346 gnd.n2351 9.3005
R14934 gnd.n3345 gnd.n2352 9.3005
R14935 gnd.n2357 gnd.n2353 9.3005
R14936 gnd.n3339 gnd.n2358 9.3005
R14937 gnd.n3338 gnd.n2359 9.3005
R14938 gnd.n3337 gnd.n2360 9.3005
R14939 gnd.n2365 gnd.n2361 9.3005
R14940 gnd.n3331 gnd.n2366 9.3005
R14941 gnd.n3330 gnd.n2367 9.3005
R14942 gnd.n3329 gnd.n2368 9.3005
R14943 gnd.n2373 gnd.n2369 9.3005
R14944 gnd.n3323 gnd.n2374 9.3005
R14945 gnd.n3322 gnd.n2375 9.3005
R14946 gnd.n3321 gnd.n2376 9.3005
R14947 gnd.n2381 gnd.n2377 9.3005
R14948 gnd.n3315 gnd.n2382 9.3005
R14949 gnd.n3314 gnd.n2383 9.3005
R14950 gnd.n3313 gnd.n2384 9.3005
R14951 gnd.n2389 gnd.n2385 9.3005
R14952 gnd.n3307 gnd.n2390 9.3005
R14953 gnd.n3306 gnd.n2391 9.3005
R14954 gnd.n3305 gnd.n2392 9.3005
R14955 gnd.n2397 gnd.n2393 9.3005
R14956 gnd.n3299 gnd.n2398 9.3005
R14957 gnd.n3298 gnd.n2399 9.3005
R14958 gnd.n3297 gnd.n2400 9.3005
R14959 gnd.n2405 gnd.n2401 9.3005
R14960 gnd.n3291 gnd.n2406 9.3005
R14961 gnd.n3290 gnd.n2407 9.3005
R14962 gnd.n3289 gnd.n2408 9.3005
R14963 gnd.n2413 gnd.n2409 9.3005
R14964 gnd.n3283 gnd.n2414 9.3005
R14965 gnd.n3282 gnd.n2415 9.3005
R14966 gnd.n3281 gnd.n2416 9.3005
R14967 gnd.n2421 gnd.n2417 9.3005
R14968 gnd.n3275 gnd.n2422 9.3005
R14969 gnd.n3274 gnd.n2423 9.3005
R14970 gnd.n3273 gnd.n2424 9.3005
R14971 gnd.n2429 gnd.n2425 9.3005
R14972 gnd.n3267 gnd.n2430 9.3005
R14973 gnd.n3266 gnd.n2431 9.3005
R14974 gnd.n3265 gnd.n2432 9.3005
R14975 gnd.n2437 gnd.n2433 9.3005
R14976 gnd.n3259 gnd.n2438 9.3005
R14977 gnd.n3258 gnd.n2439 9.3005
R14978 gnd.n3257 gnd.n2440 9.3005
R14979 gnd.n2445 gnd.n2441 9.3005
R14980 gnd.n3251 gnd.n2446 9.3005
R14981 gnd.n3250 gnd.n2447 9.3005
R14982 gnd.n3249 gnd.n2448 9.3005
R14983 gnd.n2453 gnd.n2449 9.3005
R14984 gnd.n3243 gnd.n2454 9.3005
R14985 gnd.n3242 gnd.n2455 9.3005
R14986 gnd.n3241 gnd.n2456 9.3005
R14987 gnd.n2461 gnd.n2457 9.3005
R14988 gnd.n3235 gnd.n2462 9.3005
R14989 gnd.n3234 gnd.n2463 9.3005
R14990 gnd.n3233 gnd.n2464 9.3005
R14991 gnd.n2469 gnd.n2465 9.3005
R14992 gnd.n3227 gnd.n2470 9.3005
R14993 gnd.n3226 gnd.n2471 9.3005
R14994 gnd.n3225 gnd.n2472 9.3005
R14995 gnd.n2477 gnd.n2473 9.3005
R14996 gnd.n3219 gnd.n2478 9.3005
R14997 gnd.n3218 gnd.n2479 9.3005
R14998 gnd.n3217 gnd.n2480 9.3005
R14999 gnd.n2485 gnd.n2481 9.3005
R15000 gnd.n3211 gnd.n2486 9.3005
R15001 gnd.n3210 gnd.n2487 9.3005
R15002 gnd.n3209 gnd.n2488 9.3005
R15003 gnd.n2493 gnd.n2489 9.3005
R15004 gnd.n3203 gnd.n2494 9.3005
R15005 gnd.n3202 gnd.n2495 9.3005
R15006 gnd.n3201 gnd.n2496 9.3005
R15007 gnd.n2501 gnd.n2497 9.3005
R15008 gnd.n3195 gnd.n2502 9.3005
R15009 gnd.n3194 gnd.n2503 9.3005
R15010 gnd.n3193 gnd.n2504 9.3005
R15011 gnd.n2509 gnd.n2505 9.3005
R15012 gnd.n3187 gnd.n2510 9.3005
R15013 gnd.n3186 gnd.n2511 9.3005
R15014 gnd.n3185 gnd.n2512 9.3005
R15015 gnd.n2517 gnd.n2513 9.3005
R15016 gnd.n3179 gnd.n2518 9.3005
R15017 gnd.n3178 gnd.n2519 9.3005
R15018 gnd.n3177 gnd.n2520 9.3005
R15019 gnd.n2525 gnd.n2521 9.3005
R15020 gnd.n3171 gnd.n2526 9.3005
R15021 gnd.n3170 gnd.n2527 9.3005
R15022 gnd.n3169 gnd.n2528 9.3005
R15023 gnd.n2533 gnd.n2529 9.3005
R15024 gnd.n3163 gnd.n2534 9.3005
R15025 gnd.n3162 gnd.n2535 9.3005
R15026 gnd.n3161 gnd.n2536 9.3005
R15027 gnd.n2541 gnd.n2537 9.3005
R15028 gnd.n3155 gnd.n2542 9.3005
R15029 gnd.n3154 gnd.n2543 9.3005
R15030 gnd.n3153 gnd.n2544 9.3005
R15031 gnd.n2549 gnd.n2545 9.3005
R15032 gnd.n3147 gnd.n2550 9.3005
R15033 gnd.n3146 gnd.n2551 9.3005
R15034 gnd.n3145 gnd.n2552 9.3005
R15035 gnd.n2557 gnd.n2553 9.3005
R15036 gnd.n3139 gnd.n2558 9.3005
R15037 gnd.n3138 gnd.n2559 9.3005
R15038 gnd.n3137 gnd.n2560 9.3005
R15039 gnd.n2565 gnd.n2561 9.3005
R15040 gnd.n3131 gnd.n2566 9.3005
R15041 gnd.n3130 gnd.n2567 9.3005
R15042 gnd.n3129 gnd.n2568 9.3005
R15043 gnd.n2573 gnd.n2569 9.3005
R15044 gnd.n3123 gnd.n2574 9.3005
R15045 gnd.n3122 gnd.n2575 9.3005
R15046 gnd.n3121 gnd.n2576 9.3005
R15047 gnd.n2581 gnd.n2577 9.3005
R15048 gnd.n3115 gnd.n2582 9.3005
R15049 gnd.n3114 gnd.n2583 9.3005
R15050 gnd.n3113 gnd.n2584 9.3005
R15051 gnd.n2589 gnd.n2585 9.3005
R15052 gnd.n3107 gnd.n2590 9.3005
R15053 gnd.n3106 gnd.n2591 9.3005
R15054 gnd.n3105 gnd.n2592 9.3005
R15055 gnd.n2597 gnd.n2593 9.3005
R15056 gnd.n3099 gnd.n2598 9.3005
R15057 gnd.n3098 gnd.n2599 9.3005
R15058 gnd.n3097 gnd.n2600 9.3005
R15059 gnd.n2605 gnd.n2601 9.3005
R15060 gnd.n3091 gnd.n2606 9.3005
R15061 gnd.n3090 gnd.n2607 9.3005
R15062 gnd.n3089 gnd.n2608 9.3005
R15063 gnd.n2613 gnd.n2609 9.3005
R15064 gnd.n3083 gnd.n2614 9.3005
R15065 gnd.n3082 gnd.n2615 9.3005
R15066 gnd.n3081 gnd.n2616 9.3005
R15067 gnd.n2621 gnd.n2617 9.3005
R15068 gnd.n3075 gnd.n2622 9.3005
R15069 gnd.n3074 gnd.n2623 9.3005
R15070 gnd.n3073 gnd.n2624 9.3005
R15071 gnd.n2629 gnd.n2625 9.3005
R15072 gnd.n3067 gnd.n2630 9.3005
R15073 gnd.n3066 gnd.n2631 9.3005
R15074 gnd.n3065 gnd.n2632 9.3005
R15075 gnd.n2637 gnd.n2633 9.3005
R15076 gnd.n3059 gnd.n2638 9.3005
R15077 gnd.n3058 gnd.n2639 9.3005
R15078 gnd.n3057 gnd.n2640 9.3005
R15079 gnd.n2645 gnd.n2641 9.3005
R15080 gnd.n3051 gnd.n2646 9.3005
R15081 gnd.n3050 gnd.n2647 9.3005
R15082 gnd.n3049 gnd.n2648 9.3005
R15083 gnd.n2653 gnd.n2649 9.3005
R15084 gnd.n3043 gnd.n2654 9.3005
R15085 gnd.n3042 gnd.n2655 9.3005
R15086 gnd.n3041 gnd.n2656 9.3005
R15087 gnd.n2661 gnd.n2657 9.3005
R15088 gnd.n3035 gnd.n2662 9.3005
R15089 gnd.n3034 gnd.n3033 9.3005
R15090 gnd.n2664 gnd.n2663 9.3005
R15091 gnd.n3025 gnd.n2668 9.3005
R15092 gnd.n3024 gnd.n2669 9.3005
R15093 gnd.n3023 gnd.n2670 9.3005
R15094 gnd.n2675 gnd.n2671 9.3005
R15095 gnd.n3017 gnd.n2676 9.3005
R15096 gnd.n3016 gnd.n2677 9.3005
R15097 gnd.n3015 gnd.n2678 9.3005
R15098 gnd.n2683 gnd.n2679 9.3005
R15099 gnd.n3009 gnd.n2684 9.3005
R15100 gnd.n3008 gnd.n2685 9.3005
R15101 gnd.n3007 gnd.n2686 9.3005
R15102 gnd.n2691 gnd.n2687 9.3005
R15103 gnd.n3001 gnd.n2692 9.3005
R15104 gnd.n3000 gnd.n2693 9.3005
R15105 gnd.n2999 gnd.n2694 9.3005
R15106 gnd.n2699 gnd.n2695 9.3005
R15107 gnd.n2993 gnd.n2700 9.3005
R15108 gnd.n2992 gnd.n2701 9.3005
R15109 gnd.n2991 gnd.n2702 9.3005
R15110 gnd.n2707 gnd.n2703 9.3005
R15111 gnd.n2985 gnd.n2708 9.3005
R15112 gnd.n2984 gnd.n2709 9.3005
R15113 gnd.n2983 gnd.n2710 9.3005
R15114 gnd.n2715 gnd.n2711 9.3005
R15115 gnd.n2977 gnd.n2716 9.3005
R15116 gnd.n2976 gnd.n2717 9.3005
R15117 gnd.n2975 gnd.n2718 9.3005
R15118 gnd.n2723 gnd.n2719 9.3005
R15119 gnd.n2969 gnd.n2724 9.3005
R15120 gnd.n2968 gnd.n2725 9.3005
R15121 gnd.n2967 gnd.n2726 9.3005
R15122 gnd.n2731 gnd.n2727 9.3005
R15123 gnd.n2961 gnd.n2732 9.3005
R15124 gnd.n2960 gnd.n2733 9.3005
R15125 gnd.n2959 gnd.n2734 9.3005
R15126 gnd.n2739 gnd.n2735 9.3005
R15127 gnd.n2953 gnd.n2740 9.3005
R15128 gnd.n2952 gnd.n2741 9.3005
R15129 gnd.n2951 gnd.n2742 9.3005
R15130 gnd.n2747 gnd.n2743 9.3005
R15131 gnd.n2945 gnd.n2748 9.3005
R15132 gnd.n2944 gnd.n2749 9.3005
R15133 gnd.n2943 gnd.n2750 9.3005
R15134 gnd.n2755 gnd.n2751 9.3005
R15135 gnd.n2937 gnd.n2756 9.3005
R15136 gnd.n2936 gnd.n2757 9.3005
R15137 gnd.n2935 gnd.n2758 9.3005
R15138 gnd.n2763 gnd.n2759 9.3005
R15139 gnd.n2929 gnd.n2764 9.3005
R15140 gnd.n2928 gnd.n2765 9.3005
R15141 gnd.n2927 gnd.n2766 9.3005
R15142 gnd.n2771 gnd.n2767 9.3005
R15143 gnd.n2921 gnd.n2772 9.3005
R15144 gnd.n2920 gnd.n2773 9.3005
R15145 gnd.n2919 gnd.n2774 9.3005
R15146 gnd.n2779 gnd.n2775 9.3005
R15147 gnd.n2913 gnd.n2780 9.3005
R15148 gnd.n2912 gnd.n2781 9.3005
R15149 gnd.n2911 gnd.n2782 9.3005
R15150 gnd.n2787 gnd.n2783 9.3005
R15151 gnd.n2905 gnd.n2788 9.3005
R15152 gnd.n2904 gnd.n2789 9.3005
R15153 gnd.n2903 gnd.n2790 9.3005
R15154 gnd.n2793 gnd.n2791 9.3005
R15155 gnd.n2897 gnd.n2896 9.3005
R15156 gnd.n3032 gnd.n3031 9.3005
R15157 gnd.n7347 gnd.n508 9.3005
R15158 gnd.n7346 gnd.n510 9.3005
R15159 gnd.n514 gnd.n511 9.3005
R15160 gnd.n7341 gnd.n515 9.3005
R15161 gnd.n7340 gnd.n516 9.3005
R15162 gnd.n7339 gnd.n517 9.3005
R15163 gnd.n521 gnd.n518 9.3005
R15164 gnd.n7334 gnd.n522 9.3005
R15165 gnd.n7333 gnd.n523 9.3005
R15166 gnd.n7332 gnd.n524 9.3005
R15167 gnd.n528 gnd.n525 9.3005
R15168 gnd.n7327 gnd.n529 9.3005
R15169 gnd.n7326 gnd.n530 9.3005
R15170 gnd.n7325 gnd.n531 9.3005
R15171 gnd.n538 gnd.n532 9.3005
R15172 gnd.n7320 gnd.n539 9.3005
R15173 gnd.n7319 gnd.n540 9.3005
R15174 gnd.n7318 gnd.n541 9.3005
R15175 gnd.n545 gnd.n542 9.3005
R15176 gnd.n7313 gnd.n546 9.3005
R15177 gnd.n7312 gnd.n547 9.3005
R15178 gnd.n7311 gnd.n548 9.3005
R15179 gnd.n552 gnd.n549 9.3005
R15180 gnd.n7306 gnd.n553 9.3005
R15181 gnd.n7305 gnd.n554 9.3005
R15182 gnd.n7304 gnd.n555 9.3005
R15183 gnd.n559 gnd.n556 9.3005
R15184 gnd.n7299 gnd.n560 9.3005
R15185 gnd.n7298 gnd.n561 9.3005
R15186 gnd.n7297 gnd.n562 9.3005
R15187 gnd.n566 gnd.n563 9.3005
R15188 gnd.n7292 gnd.n567 9.3005
R15189 gnd.n7291 gnd.n7290 9.3005
R15190 gnd.n7289 gnd.n570 9.3005
R15191 gnd.n7349 gnd.n7348 9.3005
R15192 gnd.n6896 gnd.n903 9.3005
R15193 gnd.n6895 gnd.n905 9.3005
R15194 gnd.n6894 gnd.n906 9.3005
R15195 gnd.n6757 gnd.n907 9.3005
R15196 gnd.n6761 gnd.n6760 9.3005
R15197 gnd.n6762 gnd.n6756 9.3005
R15198 gnd.n6766 gnd.n6763 9.3005
R15199 gnd.n6767 gnd.n6755 9.3005
R15200 gnd.n6771 gnd.n6770 9.3005
R15201 gnd.n6772 gnd.n6754 9.3005
R15202 gnd.n6776 gnd.n6773 9.3005
R15203 gnd.n6777 gnd.n6753 9.3005
R15204 gnd.n6781 gnd.n6780 9.3005
R15205 gnd.n6782 gnd.n6752 9.3005
R15206 gnd.n6809 gnd.n6783 9.3005
R15207 gnd.n6808 gnd.n6784 9.3005
R15208 gnd.n6807 gnd.n6785 9.3005
R15209 gnd.n6804 gnd.n6786 9.3005
R15210 gnd.n6803 gnd.n6787 9.3005
R15211 gnd.n6800 gnd.n6788 9.3005
R15212 gnd.n6799 gnd.n6789 9.3005
R15213 gnd.n6796 gnd.n6790 9.3005
R15214 gnd.n6795 gnd.n6792 9.3005
R15215 gnd.n6791 gnd.n931 9.3005
R15216 gnd.n6852 gnd.n932 9.3005
R15217 gnd.n6851 gnd.n671 9.3005
R15218 gnd.n6850 gnd.n933 9.3005
R15219 gnd.n6847 gnd.n934 9.3005
R15220 gnd.n6846 gnd.n935 9.3005
R15221 gnd.n2838 gnd.n936 9.3005
R15222 gnd.n2842 gnd.n2839 9.3005
R15223 gnd.n2843 gnd.n2837 9.3005
R15224 gnd.n2847 gnd.n2846 9.3005
R15225 gnd.n2848 gnd.n2836 9.3005
R15226 gnd.n2852 gnd.n2849 9.3005
R15227 gnd.n2853 gnd.n2835 9.3005
R15228 gnd.n2857 gnd.n2856 9.3005
R15229 gnd.n2858 gnd.n2834 9.3005
R15230 gnd.n2862 gnd.n2859 9.3005
R15231 gnd.n2863 gnd.n2833 9.3005
R15232 gnd.n2867 gnd.n2866 9.3005
R15233 gnd.n2868 gnd.n2832 9.3005
R15234 gnd.n2886 gnd.n2869 9.3005
R15235 gnd.n2885 gnd.n2870 9.3005
R15236 gnd.n2884 gnd.n2871 9.3005
R15237 gnd.n2881 gnd.n2872 9.3005
R15238 gnd.n2880 gnd.n2873 9.3005
R15239 gnd.n2878 gnd.n2874 9.3005
R15240 gnd.n2877 gnd.n2876 9.3005
R15241 gnd.n2875 gnd.n574 9.3005
R15242 gnd.n7286 gnd.n573 9.3005
R15243 gnd.n7288 gnd.n7287 9.3005
R15244 gnd.n6898 gnd.n6897 9.3005
R15245 gnd.n6904 gnd.n6903 9.3005
R15246 gnd.n6905 gnd.n897 9.3005
R15247 gnd.n6908 gnd.n896 9.3005
R15248 gnd.n6909 gnd.n895 9.3005
R15249 gnd.n6912 gnd.n894 9.3005
R15250 gnd.n6913 gnd.n893 9.3005
R15251 gnd.n6916 gnd.n892 9.3005
R15252 gnd.n6917 gnd.n891 9.3005
R15253 gnd.n6920 gnd.n890 9.3005
R15254 gnd.n6921 gnd.n889 9.3005
R15255 gnd.n6924 gnd.n888 9.3005
R15256 gnd.n6925 gnd.n887 9.3005
R15257 gnd.n6928 gnd.n886 9.3005
R15258 gnd.n6929 gnd.n885 9.3005
R15259 gnd.n6932 gnd.n884 9.3005
R15260 gnd.n6933 gnd.n883 9.3005
R15261 gnd.n6936 gnd.n882 9.3005
R15262 gnd.n6938 gnd.n876 9.3005
R15263 gnd.n6941 gnd.n875 9.3005
R15264 gnd.n6942 gnd.n874 9.3005
R15265 gnd.n6945 gnd.n873 9.3005
R15266 gnd.n6946 gnd.n872 9.3005
R15267 gnd.n6949 gnd.n871 9.3005
R15268 gnd.n6950 gnd.n870 9.3005
R15269 gnd.n6953 gnd.n869 9.3005
R15270 gnd.n6954 gnd.n868 9.3005
R15271 gnd.n6957 gnd.n867 9.3005
R15272 gnd.n6959 gnd.n866 9.3005
R15273 gnd.n6960 gnd.n865 9.3005
R15274 gnd.n6961 gnd.n864 9.3005
R15275 gnd.n863 gnd.n784 9.3005
R15276 gnd.n6902 gnd.n902 9.3005
R15277 gnd.n6901 gnd.n6900 9.3005
R15278 gnd.n7019 gnd.n783 9.3005
R15279 gnd.n7021 gnd.n7020 9.3005
R15280 gnd.n768 gnd.n767 9.3005
R15281 gnd.n7034 gnd.n7033 9.3005
R15282 gnd.n7035 gnd.n766 9.3005
R15283 gnd.n7037 gnd.n7036 9.3005
R15284 gnd.n750 gnd.n749 9.3005
R15285 gnd.n7050 gnd.n7049 9.3005
R15286 gnd.n7051 gnd.n748 9.3005
R15287 gnd.n7053 gnd.n7052 9.3005
R15288 gnd.n732 gnd.n731 9.3005
R15289 gnd.n7066 gnd.n7065 9.3005
R15290 gnd.n7067 gnd.n730 9.3005
R15291 gnd.n7069 gnd.n7068 9.3005
R15292 gnd.n715 gnd.n714 9.3005
R15293 gnd.n7082 gnd.n7081 9.3005
R15294 gnd.n7083 gnd.n713 9.3005
R15295 gnd.n7086 gnd.n7085 9.3005
R15296 gnd.n7084 gnd.n696 9.3005
R15297 gnd.n7098 gnd.n697 9.3005
R15298 gnd.n7146 gnd.n7145 9.3005
R15299 gnd.n7147 gnd.n648 9.3005
R15300 gnd.n7149 gnd.n7148 9.3005
R15301 gnd.n633 gnd.n632 9.3005
R15302 gnd.n7162 gnd.n7161 9.3005
R15303 gnd.n7163 gnd.n631 9.3005
R15304 gnd.n7165 gnd.n7164 9.3005
R15305 gnd.n616 gnd.n615 9.3005
R15306 gnd.n7178 gnd.n7177 9.3005
R15307 gnd.n7179 gnd.n614 9.3005
R15308 gnd.n7181 gnd.n7180 9.3005
R15309 gnd.n600 gnd.n599 9.3005
R15310 gnd.n7194 gnd.n7193 9.3005
R15311 gnd.n7195 gnd.n598 9.3005
R15312 gnd.n7197 gnd.n7196 9.3005
R15313 gnd.n581 gnd.n580 9.3005
R15314 gnd.n7278 gnd.n7277 9.3005
R15315 gnd.n7279 gnd.n579 9.3005
R15316 gnd.n7281 gnd.n7280 9.3005
R15317 gnd.n507 gnd.n506 9.3005
R15318 gnd.n7351 gnd.n7350 9.3005
R15319 gnd.n7018 gnd.n7017 9.3005
R15320 gnd.n650 gnd.n649 9.3005
R15321 gnd.n5464 gnd.n5463 9.3005
R15322 gnd.n5465 gnd.n5458 9.3005
R15323 gnd.n5467 gnd.n5466 9.3005
R15324 gnd.n5456 gnd.n5455 9.3005
R15325 gnd.n5472 gnd.n5471 9.3005
R15326 gnd.n5473 gnd.n5454 9.3005
R15327 gnd.n5475 gnd.n5474 9.3005
R15328 gnd.n5452 gnd.n5451 9.3005
R15329 gnd.n5517 gnd.n5516 9.3005
R15330 gnd.n5518 gnd.n5450 9.3005
R15331 gnd.n5520 gnd.n5519 9.3005
R15332 gnd.n5448 gnd.n5447 9.3005
R15333 gnd.n5525 gnd.n5524 9.3005
R15334 gnd.n5526 gnd.n5446 9.3005
R15335 gnd.n5528 gnd.n5527 9.3005
R15336 gnd.n5444 gnd.n5443 9.3005
R15337 gnd.n5533 gnd.n5532 9.3005
R15338 gnd.n5534 gnd.n5442 9.3005
R15339 gnd.n5556 gnd.n5535 9.3005
R15340 gnd.n5555 gnd.n5536 9.3005
R15341 gnd.n5554 gnd.n5537 9.3005
R15342 gnd.n5540 gnd.n5538 9.3005
R15343 gnd.n5549 gnd.n5541 9.3005
R15344 gnd.n5548 gnd.n5542 9.3005
R15345 gnd.n5547 gnd.n5543 9.3005
R15346 gnd.n1673 gnd.n1672 9.3005
R15347 gnd.n5813 gnd.n5812 9.3005
R15348 gnd.n5814 gnd.n1671 9.3005
R15349 gnd.n5816 gnd.n5815 9.3005
R15350 gnd.n1661 gnd.n1660 9.3005
R15351 gnd.n5833 gnd.n5832 9.3005
R15352 gnd.n5834 gnd.n1659 9.3005
R15353 gnd.n5836 gnd.n5835 9.3005
R15354 gnd.n1648 gnd.n1647 9.3005
R15355 gnd.n5853 gnd.n5852 9.3005
R15356 gnd.n5854 gnd.n1646 9.3005
R15357 gnd.n5858 gnd.n5855 9.3005
R15358 gnd.n5857 gnd.n5856 9.3005
R15359 gnd.n1430 gnd.n1429 9.3005
R15360 gnd.n6064 gnd.n6063 9.3005
R15361 gnd.n6065 gnd.n1428 9.3005
R15362 gnd.n6069 gnd.n6066 9.3005
R15363 gnd.n6068 gnd.n6067 9.3005
R15364 gnd.n1397 gnd.n1396 9.3005
R15365 gnd.n6146 gnd.n6145 9.3005
R15366 gnd.n6147 gnd.n1395 9.3005
R15367 gnd.n6149 gnd.n6148 9.3005
R15368 gnd.n1373 gnd.n1372 9.3005
R15369 gnd.n6174 gnd.n6173 9.3005
R15370 gnd.n6175 gnd.n1371 9.3005
R15371 gnd.n6192 gnd.n6176 9.3005
R15372 gnd.n6191 gnd.n6177 9.3005
R15373 gnd.n6190 gnd.n6178 9.3005
R15374 gnd.n6181 gnd.n6179 9.3005
R15375 gnd.n6185 gnd.n6182 9.3005
R15376 gnd.n6184 gnd.n6183 9.3005
R15377 gnd.n1312 gnd.n1311 9.3005
R15378 gnd.n6285 gnd.n6284 9.3005
R15379 gnd.n6286 gnd.n1310 9.3005
R15380 gnd.n6301 gnd.n6287 9.3005
R15381 gnd.n6300 gnd.n6288 9.3005
R15382 gnd.n6299 gnd.n6289 9.3005
R15383 gnd.n6291 gnd.n6290 9.3005
R15384 gnd.n6294 gnd.n6293 9.3005
R15385 gnd.n6292 gnd.n1268 9.3005
R15386 gnd.n6387 gnd.n1269 9.3005
R15387 gnd.n6386 gnd.n1270 9.3005
R15388 gnd.n6385 gnd.n1272 9.3005
R15389 gnd.n1271 gnd.n1239 9.3005
R15390 gnd.n6424 gnd.n1240 9.3005
R15391 gnd.n6423 gnd.n1241 9.3005
R15392 gnd.n6422 gnd.n1243 9.3005
R15393 gnd.n1242 gnd.n1210 9.3005
R15394 gnd.n6464 gnd.n1211 9.3005
R15395 gnd.n6463 gnd.n1212 9.3005
R15396 gnd.n6462 gnd.n1213 9.3005
R15397 gnd.n1215 gnd.n1214 9.3005
R15398 gnd.n1107 gnd.n1106 9.3005
R15399 gnd.n6614 gnd.n6613 9.3005
R15400 gnd.n6615 gnd.n1105 9.3005
R15401 gnd.n6619 gnd.n6616 9.3005
R15402 gnd.n6618 gnd.n6617 9.3005
R15403 gnd.n1081 gnd.n1080 9.3005
R15404 gnd.n6644 gnd.n6643 9.3005
R15405 gnd.n6645 gnd.n1079 9.3005
R15406 gnd.n6649 gnd.n6646 9.3005
R15407 gnd.n6648 gnd.n6647 9.3005
R15408 gnd.n1056 gnd.n1055 9.3005
R15409 gnd.n6675 gnd.n6674 9.3005
R15410 gnd.n6676 gnd.n1054 9.3005
R15411 gnd.n6691 gnd.n6677 9.3005
R15412 gnd.n6690 gnd.n6678 9.3005
R15413 gnd.n6689 gnd.n6679 9.3005
R15414 gnd.n6681 gnd.n6680 9.3005
R15415 gnd.n6683 gnd.n6682 9.3005
R15416 gnd.n971 gnd.n970 9.3005
R15417 gnd.n6716 gnd.n6715 9.3005
R15418 gnd.n6717 gnd.n969 9.3005
R15419 gnd.n6719 gnd.n6718 9.3005
R15420 gnd.n967 gnd.n966 9.3005
R15421 gnd.n6724 gnd.n6723 9.3005
R15422 gnd.n6725 gnd.n965 9.3005
R15423 gnd.n6727 gnd.n6726 9.3005
R15424 gnd.n963 gnd.n962 9.3005
R15425 gnd.n6732 gnd.n6731 9.3005
R15426 gnd.n6733 gnd.n961 9.3005
R15427 gnd.n6735 gnd.n6734 9.3005
R15428 gnd.n959 gnd.n958 9.3005
R15429 gnd.n6740 gnd.n6739 9.3005
R15430 gnd.n6741 gnd.n957 9.3005
R15431 gnd.n6743 gnd.n6742 9.3005
R15432 gnd.n955 gnd.n954 9.3005
R15433 gnd.n6748 gnd.n6747 9.3005
R15434 gnd.n6749 gnd.n953 9.3005
R15435 gnd.n6751 gnd.n6750 9.3005
R15436 gnd.n951 gnd.n950 9.3005
R15437 gnd.n6817 gnd.n6816 9.3005
R15438 gnd.n6818 gnd.n949 9.3005
R15439 gnd.n6820 gnd.n6819 9.3005
R15440 gnd.n946 gnd.n945 9.3005
R15441 gnd.n6837 gnd.n6836 9.3005
R15442 gnd.n2806 gnd.n941 9.3005
R15443 gnd.n2811 gnd.n2810 9.3005
R15444 gnd.n2812 gnd.n2805 9.3005
R15445 gnd.n2814 gnd.n2813 9.3005
R15446 gnd.n2803 gnd.n2802 9.3005
R15447 gnd.n2819 gnd.n2818 9.3005
R15448 gnd.n2820 gnd.n2801 9.3005
R15449 gnd.n2822 gnd.n2821 9.3005
R15450 gnd.n2799 gnd.n2798 9.3005
R15451 gnd.n2827 gnd.n2826 9.3005
R15452 gnd.n2828 gnd.n2797 9.3005
R15453 gnd.n2831 gnd.n2830 9.3005
R15454 gnd.n2829 gnd.n2795 9.3005
R15455 gnd.n2893 gnd.n2794 9.3005
R15456 gnd.n2895 gnd.n2894 9.3005
R15457 gnd.n5410 gnd.n1897 9.3005
R15458 gnd.n5238 gnd.n2039 9.3005
R15459 gnd.n5236 gnd.n2040 9.3005
R15460 gnd.n5235 gnd.n2041 9.3005
R15461 gnd.n5233 gnd.n2042 9.3005
R15462 gnd.n5232 gnd.n2043 9.3005
R15463 gnd.n5230 gnd.n2044 9.3005
R15464 gnd.n5229 gnd.n2045 9.3005
R15465 gnd.n2193 gnd.n2046 9.3005
R15466 gnd.n2216 gnd.n2194 9.3005
R15467 gnd.n2215 gnd.n2195 9.3005
R15468 gnd.n2214 gnd.n2196 9.3005
R15469 gnd.n2198 gnd.n2197 9.3005
R15470 gnd.n1948 gnd.n1947 9.3005
R15471 gnd.n5351 gnd.n5350 9.3005
R15472 gnd.n5352 gnd.n1946 9.3005
R15473 gnd.n5360 gnd.n5353 9.3005
R15474 gnd.n5359 gnd.n5354 9.3005
R15475 gnd.n5358 gnd.n5355 9.3005
R15476 gnd.n1908 gnd.n1907 9.3005
R15477 gnd.n5391 gnd.n5390 9.3005
R15478 gnd.n5392 gnd.n1906 9.3005
R15479 gnd.n5395 gnd.n5394 9.3005
R15480 gnd.n5393 gnd.n1899 9.3005
R15481 gnd.n5407 gnd.n1898 9.3005
R15482 gnd.n5409 gnd.n5408 9.3005
R15483 gnd.n5240 gnd.n5239 9.3005
R15484 gnd.n2038 gnd.n2035 9.3005
R15485 gnd.n5251 gnd.n2034 9.3005
R15486 gnd.n5252 gnd.n2033 9.3005
R15487 gnd.n5253 gnd.n2032 9.3005
R15488 gnd.n2031 gnd.n2029 9.3005
R15489 gnd.n5259 gnd.n2028 9.3005
R15490 gnd.n5260 gnd.n2027 9.3005
R15491 gnd.n5261 gnd.n2026 9.3005
R15492 gnd.n2025 gnd.n2023 9.3005
R15493 gnd.n5267 gnd.n2022 9.3005
R15494 gnd.n5268 gnd.n2021 9.3005
R15495 gnd.n5269 gnd.n2020 9.3005
R15496 gnd.n2019 gnd.n2017 9.3005
R15497 gnd.n5275 gnd.n2016 9.3005
R15498 gnd.n5277 gnd.n5276 9.3005
R15499 gnd.n5245 gnd.n5242 9.3005
R15500 gnd.n5241 gnd.n2037 9.3005
R15501 gnd.n2003 gnd.n2002 9.3005
R15502 gnd.n5292 gnd.n5291 9.3005
R15503 gnd.n5293 gnd.n2001 9.3005
R15504 gnd.n5295 gnd.n5294 9.3005
R15505 gnd.n1985 gnd.n1984 9.3005
R15506 gnd.n5308 gnd.n5307 9.3005
R15507 gnd.n5309 gnd.n1983 9.3005
R15508 gnd.n5311 gnd.n5310 9.3005
R15509 gnd.n1968 gnd.n1967 9.3005
R15510 gnd.n5324 gnd.n5323 9.3005
R15511 gnd.n5325 gnd.n1966 9.3005
R15512 gnd.n5336 gnd.n5326 9.3005
R15513 gnd.n5335 gnd.n5327 9.3005
R15514 gnd.n5334 gnd.n5328 9.3005
R15515 gnd.n5333 gnd.n5330 9.3005
R15516 gnd.n5329 gnd.n1927 9.3005
R15517 gnd.n5377 gnd.n1928 9.3005
R15518 gnd.n5376 gnd.n1929 9.3005
R15519 gnd.n5375 gnd.n1930 9.3005
R15520 gnd.n1937 gnd.n1931 9.3005
R15521 gnd.n1936 gnd.n1933 9.3005
R15522 gnd.n1932 gnd.n1853 9.3005
R15523 gnd.n5641 gnd.n1854 9.3005
R15524 gnd.n5640 gnd.n1855 9.3005
R15525 gnd.n5639 gnd.n1856 9.3005
R15526 gnd.n5607 gnd.n1857 9.3005
R15527 gnd.n5609 gnd.n5608 9.3005
R15528 gnd.n5613 gnd.n5612 9.3005
R15529 gnd.n5614 gnd.n1885 9.3005
R15530 gnd.n5616 gnd.n5615 9.3005
R15531 gnd.n1830 gnd.n1829 9.3005
R15532 gnd.n5655 gnd.n5654 9.3005
R15533 gnd.n5656 gnd.n1828 9.3005
R15534 gnd.n5658 gnd.n5657 9.3005
R15535 gnd.n1812 gnd.n1811 9.3005
R15536 gnd.n5671 gnd.n5670 9.3005
R15537 gnd.n5672 gnd.n1810 9.3005
R15538 gnd.n5674 gnd.n5673 9.3005
R15539 gnd.n1795 gnd.n1794 9.3005
R15540 gnd.n5687 gnd.n5686 9.3005
R15541 gnd.n5688 gnd.n1793 9.3005
R15542 gnd.n5690 gnd.n5689 9.3005
R15543 gnd.n1777 gnd.n1776 9.3005
R15544 gnd.n5703 gnd.n5702 9.3005
R15545 gnd.n5704 gnd.n1775 9.3005
R15546 gnd.n5711 gnd.n5705 9.3005
R15547 gnd.n5710 gnd.n5706 9.3005
R15548 gnd.n5709 gnd.n5708 9.3005
R15549 gnd.n5707 gnd.n1616 9.3005
R15550 gnd.n5902 gnd.n1617 9.3005
R15551 gnd.n5901 gnd.n1618 9.3005
R15552 gnd.n5900 gnd.n5899 9.3005
R15553 gnd.n5279 gnd.n5278 9.3005
R15554 gnd.n1562 gnd.n1558 9.3005
R15555 gnd.n5931 gnd.n5930 9.3005
R15556 gnd.n5929 gnd.n5925 9.3005
R15557 gnd.n5936 gnd.n5924 9.3005
R15558 gnd.n5937 gnd.n5923 9.3005
R15559 gnd.n5938 gnd.n5922 9.3005
R15560 gnd.n5921 gnd.n5918 9.3005
R15561 gnd.n5943 gnd.n5917 9.3005
R15562 gnd.n5944 gnd.n5916 9.3005
R15563 gnd.n5945 gnd.n5915 9.3005
R15564 gnd.n5914 gnd.n5911 9.3005
R15565 gnd.n5913 gnd.n5910 9.3005
R15566 gnd.n5952 gnd.n5909 9.3005
R15567 gnd.n5954 gnd.n5953 9.3005
R15568 gnd.n5994 gnd.n5993 9.3005
R15569 gnd.n1564 gnd.n1563 9.3005
R15570 gnd.n1570 gnd.n1568 9.3005
R15571 gnd.n5986 gnd.n1571 9.3005
R15572 gnd.n5985 gnd.n1572 9.3005
R15573 gnd.n5984 gnd.n1573 9.3005
R15574 gnd.n1577 gnd.n1574 9.3005
R15575 gnd.n5979 gnd.n1578 9.3005
R15576 gnd.n5978 gnd.n1579 9.3005
R15577 gnd.n5977 gnd.n1580 9.3005
R15578 gnd.n1584 gnd.n1581 9.3005
R15579 gnd.n5972 gnd.n1585 9.3005
R15580 gnd.n5971 gnd.n1586 9.3005
R15581 gnd.n5970 gnd.n1587 9.3005
R15582 gnd.n1591 gnd.n1588 9.3005
R15583 gnd.n5965 gnd.n1592 9.3005
R15584 gnd.n5964 gnd.n5963 9.3005
R15585 gnd.n5962 gnd.n1593 9.3005
R15586 gnd.n5995 gnd.n1557 9.3005
R15587 gnd.n2179 gnd.n2178 9.3005
R15588 gnd.n2180 gnd.n2049 9.3005
R15589 gnd.n2183 gnd.n2181 9.3005
R15590 gnd.n2184 gnd.n2048 9.3005
R15591 gnd.n2187 gnd.n2186 9.3005
R15592 gnd.n2188 gnd.n2047 9.3005
R15593 gnd.n5225 gnd.n2189 9.3005
R15594 gnd.n5224 gnd.n2190 9.3005
R15595 gnd.n5223 gnd.n2191 9.3005
R15596 gnd.n2199 gnd.n2192 9.3005
R15597 gnd.n2210 gnd.n2200 9.3005
R15598 gnd.n2209 gnd.n2201 9.3005
R15599 gnd.n2208 gnd.n2202 9.3005
R15600 gnd.n2205 gnd.n2204 9.3005
R15601 gnd.n2203 gnd.n1942 9.3005
R15602 gnd.n5364 gnd.n1941 9.3005
R15603 gnd.n5366 gnd.n5365 9.3005
R15604 gnd.n5367 gnd.n1940 9.3005
R15605 gnd.n5371 gnd.n5368 9.3005
R15606 gnd.n5370 gnd.n5369 9.3005
R15607 gnd.n1902 gnd.n1901 9.3005
R15608 gnd.n5400 gnd.n5399 9.3005
R15609 gnd.n5401 gnd.n1900 9.3005
R15610 gnd.n5403 gnd.n5402 9.3005
R15611 gnd.n1888 gnd.n1886 9.3005
R15612 gnd.n5606 gnd.n5605 9.3005
R15613 gnd.n5604 gnd.n1887 9.3005
R15614 gnd.n5601 gnd.n1889 9.3005
R15615 gnd.n5600 gnd.n1890 9.3005
R15616 gnd.n5599 gnd.n1891 9.3005
R15617 gnd.n5598 gnd.n1892 9.3005
R15618 gnd.n5478 gnd.n1893 9.3005
R15619 gnd.n5482 gnd.n5479 9.3005
R15620 gnd.n5483 gnd.n5477 9.3005
R15621 gnd.n5487 gnd.n5486 9.3005
R15622 gnd.n5488 gnd.n5476 9.3005
R15623 gnd.n5509 gnd.n5489 9.3005
R15624 gnd.n5508 gnd.n5490 9.3005
R15625 gnd.n5507 gnd.n5491 9.3005
R15626 gnd.n5504 gnd.n5492 9.3005
R15627 gnd.n5503 gnd.n5493 9.3005
R15628 gnd.n5500 gnd.n5494 9.3005
R15629 gnd.n5499 gnd.n5496 9.3005
R15630 gnd.n5495 gnd.n5432 9.3005
R15631 gnd.n5567 gnd.n5433 9.3005
R15632 gnd.n5566 gnd.n5434 9.3005
R15633 gnd.n5565 gnd.n5435 9.3005
R15634 gnd.n5562 gnd.n5436 9.3005
R15635 gnd.n5561 gnd.n5437 9.3005
R15636 gnd.n5439 gnd.n5438 9.3005
R15637 gnd.n1597 gnd.n1596 9.3005
R15638 gnd.n5961 gnd.n5960 9.3005
R15639 gnd.n2176 gnd.n2175 9.3005
R15640 gnd.n2164 gnd.n2054 9.3005
R15641 gnd.n2166 gnd.n2165 9.3005
R15642 gnd.n2163 gnd.n2056 9.3005
R15643 gnd.n2162 gnd.n2161 9.3005
R15644 gnd.n2058 gnd.n2057 9.3005
R15645 gnd.n2155 gnd.n2154 9.3005
R15646 gnd.n2153 gnd.n2060 9.3005
R15647 gnd.n2152 gnd.n2151 9.3005
R15648 gnd.n2062 gnd.n2061 9.3005
R15649 gnd.n2145 gnd.n2144 9.3005
R15650 gnd.n2143 gnd.n2064 9.3005
R15651 gnd.n2142 gnd.n2141 9.3005
R15652 gnd.n2066 gnd.n2065 9.3005
R15653 gnd.n2135 gnd.n2134 9.3005
R15654 gnd.n2133 gnd.n2068 9.3005
R15655 gnd.n2132 gnd.n2131 9.3005
R15656 gnd.n2070 gnd.n2069 9.3005
R15657 gnd.n2125 gnd.n2121 9.3005
R15658 gnd.n2120 gnd.n2072 9.3005
R15659 gnd.n2119 gnd.n2118 9.3005
R15660 gnd.n2074 gnd.n2073 9.3005
R15661 gnd.n2112 gnd.n2111 9.3005
R15662 gnd.n2110 gnd.n2076 9.3005
R15663 gnd.n2109 gnd.n2108 9.3005
R15664 gnd.n2078 gnd.n2077 9.3005
R15665 gnd.n2102 gnd.n2101 9.3005
R15666 gnd.n2100 gnd.n2080 9.3005
R15667 gnd.n2099 gnd.n2098 9.3005
R15668 gnd.n2082 gnd.n2081 9.3005
R15669 gnd.n2092 gnd.n2091 9.3005
R15670 gnd.n2090 gnd.n2084 9.3005
R15671 gnd.n2089 gnd.n2088 9.3005
R15672 gnd.n2085 gnd.n2010 9.3005
R15673 gnd.n2053 gnd.n2050 9.3005
R15674 gnd.n2174 gnd.n2173 9.3005
R15675 gnd.n5285 gnd.n2009 9.3005
R15676 gnd.n5287 gnd.n5286 9.3005
R15677 gnd.n1994 gnd.n1993 9.3005
R15678 gnd.n5300 gnd.n5299 9.3005
R15679 gnd.n5301 gnd.n1992 9.3005
R15680 gnd.n5303 gnd.n5302 9.3005
R15681 gnd.n1976 gnd.n1975 9.3005
R15682 gnd.n5316 gnd.n5315 9.3005
R15683 gnd.n5317 gnd.n1974 9.3005
R15684 gnd.n5319 gnd.n5318 9.3005
R15685 gnd.n1958 gnd.n1957 9.3005
R15686 gnd.n5341 gnd.n5340 9.3005
R15687 gnd.n5342 gnd.n1956 9.3005
R15688 gnd.n5346 gnd.n5343 9.3005
R15689 gnd.n5345 gnd.n5344 9.3005
R15690 gnd.n1918 gnd.n1917 9.3005
R15691 gnd.n5382 gnd.n5381 9.3005
R15692 gnd.n5383 gnd.n1916 9.3005
R15693 gnd.n5385 gnd.n5384 9.3005
R15694 gnd.n5386 gnd.n1838 9.3005
R15695 gnd.n5650 gnd.n5649 9.3005
R15696 gnd.n1821 gnd.n1820 9.3005
R15697 gnd.n5663 gnd.n5662 9.3005
R15698 gnd.n5664 gnd.n1819 9.3005
R15699 gnd.n5666 gnd.n5665 9.3005
R15700 gnd.n1804 gnd.n1803 9.3005
R15701 gnd.n5679 gnd.n5678 9.3005
R15702 gnd.n5680 gnd.n1802 9.3005
R15703 gnd.n5682 gnd.n5681 9.3005
R15704 gnd.n1786 gnd.n1785 9.3005
R15705 gnd.n5695 gnd.n5694 9.3005
R15706 gnd.n5696 gnd.n1784 9.3005
R15707 gnd.n5698 gnd.n5697 9.3005
R15708 gnd.n1767 gnd.n1766 9.3005
R15709 gnd.n5716 gnd.n5715 9.3005
R15710 gnd.n5717 gnd.n1765 9.3005
R15711 gnd.n5719 gnd.n5718 9.3005
R15712 gnd.n1609 gnd.n1608 9.3005
R15713 gnd.n5907 gnd.n5906 9.3005
R15714 gnd.n5908 gnd.n1607 9.3005
R15715 gnd.n5956 gnd.n5955 9.3005
R15716 gnd.n5284 gnd.n5283 9.3005
R15717 gnd.n5648 gnd.n1837 9.3005
R15718 gnd.n5172 gnd.n5171 9.3005
R15719 gnd.n5173 gnd.n2220 9.3005
R15720 gnd.n5218 gnd.n5174 9.3005
R15721 gnd.n5217 gnd.n5175 9.3005
R15722 gnd.n5216 gnd.n5176 9.3005
R15723 gnd.n5179 gnd.n5177 9.3005
R15724 gnd.n5212 gnd.n5180 9.3005
R15725 gnd.n5211 gnd.n5181 9.3005
R15726 gnd.n5210 gnd.n5182 9.3005
R15727 gnd.n5185 gnd.n5183 9.3005
R15728 gnd.n5206 gnd.n5186 9.3005
R15729 gnd.n5205 gnd.n5187 9.3005
R15730 gnd.n5204 gnd.n5188 9.3005
R15731 gnd.n5190 gnd.n5189 9.3005
R15732 gnd.n2222 gnd.n2221 9.3005
R15733 gnd.n5165 gnd.n2224 9.3005
R15734 gnd.n5164 gnd.n5163 9.3005
R15735 gnd.n2226 gnd.n2225 9.3005
R15736 gnd.n3531 gnd.n3530 9.3005
R15737 gnd.n3529 gnd.n2230 9.3005
R15738 gnd.n3528 gnd.n3527 9.3005
R15739 gnd.n2232 gnd.n2231 9.3005
R15740 gnd.n3521 gnd.n3520 9.3005
R15741 gnd.n3519 gnd.n2236 9.3005
R15742 gnd.n3518 gnd.n3517 9.3005
R15743 gnd.n2238 gnd.n2237 9.3005
R15744 gnd.n3511 gnd.n3510 9.3005
R15745 gnd.n3509 gnd.n2242 9.3005
R15746 gnd.n3508 gnd.n3507 9.3005
R15747 gnd.n2244 gnd.n2243 9.3005
R15748 gnd.n3501 gnd.n3500 9.3005
R15749 gnd.n3499 gnd.n2248 9.3005
R15750 gnd.n3498 gnd.n3497 9.3005
R15751 gnd.n2250 gnd.n2249 9.3005
R15752 gnd.n3491 gnd.n3490 9.3005
R15753 gnd.n3489 gnd.n2254 9.3005
R15754 gnd.n3488 gnd.n3487 9.3005
R15755 gnd.n2256 gnd.n2255 9.3005
R15756 gnd.n3481 gnd.n3480 9.3005
R15757 gnd.n3479 gnd.n2260 9.3005
R15758 gnd.n3478 gnd.n3477 9.3005
R15759 gnd.n2262 gnd.n2261 9.3005
R15760 gnd.n3471 gnd.n3470 9.3005
R15761 gnd.n3469 gnd.n2266 9.3005
R15762 gnd.n3468 gnd.n3467 9.3005
R15763 gnd.n2268 gnd.n2267 9.3005
R15764 gnd.n3461 gnd.n3460 9.3005
R15765 gnd.n3459 gnd.n2272 9.3005
R15766 gnd.n3458 gnd.n3457 9.3005
R15767 gnd.n2274 gnd.n2273 9.3005
R15768 gnd.n3451 gnd.n3450 9.3005
R15769 gnd.n3449 gnd.n2278 9.3005
R15770 gnd.n3448 gnd.n3447 9.3005
R15771 gnd.n2280 gnd.n2279 9.3005
R15772 gnd.n3441 gnd.n3440 9.3005
R15773 gnd.n3439 gnd.n2284 9.3005
R15774 gnd.n3438 gnd.n3437 9.3005
R15775 gnd.n2286 gnd.n2285 9.3005
R15776 gnd.n3431 gnd.n3430 9.3005
R15777 gnd.n3429 gnd.n2290 9.3005
R15778 gnd.n3428 gnd.n3427 9.3005
R15779 gnd.n2292 gnd.n2291 9.3005
R15780 gnd.n3421 gnd.n3420 9.3005
R15781 gnd.n3419 gnd.n2296 9.3005
R15782 gnd.n3418 gnd.n3417 9.3005
R15783 gnd.n2298 gnd.n2297 9.3005
R15784 gnd.n3411 gnd.n3410 9.3005
R15785 gnd.n3409 gnd.n2302 9.3005
R15786 gnd.n3408 gnd.n3407 9.3005
R15787 gnd.n2304 gnd.n2303 9.3005
R15788 gnd.n3401 gnd.n3400 9.3005
R15789 gnd.n3399 gnd.n2308 9.3005
R15790 gnd.n3398 gnd.n3397 9.3005
R15791 gnd.n2310 gnd.n2309 9.3005
R15792 gnd.n3391 gnd.n3390 9.3005
R15793 gnd.n3389 gnd.n2314 9.3005
R15794 gnd.n3388 gnd.n3387 9.3005
R15795 gnd.n2316 gnd.n2315 9.3005
R15796 gnd.n3381 gnd.n3380 9.3005
R15797 gnd.n3379 gnd.n2320 9.3005
R15798 gnd.n3378 gnd.n3377 9.3005
R15799 gnd.n5167 gnd.n5166 9.3005
R15800 gnd.n7005 gnd.n7004 9.3005
R15801 gnd.n798 gnd.n797 9.3005
R15802 gnd.n6999 gnd.n6998 9.3005
R15803 gnd.n6997 gnd.n6996 9.3005
R15804 gnd.n806 gnd.n805 9.3005
R15805 gnd.n6991 gnd.n6990 9.3005
R15806 gnd.n6989 gnd.n6988 9.3005
R15807 gnd.n814 gnd.n813 9.3005
R15808 gnd.n6983 gnd.n6982 9.3005
R15809 gnd.n6981 gnd.n6980 9.3005
R15810 gnd.n822 gnd.n821 9.3005
R15811 gnd.n6975 gnd.n6974 9.3005
R15812 gnd.n6973 gnd.n6972 9.3005
R15813 gnd.n830 gnd.n829 9.3005
R15814 gnd.n1007 gnd.n1006 9.3005
R15815 gnd.n1011 gnd.n1010 9.3005
R15816 gnd.n7007 gnd.n7006 9.3005
R15817 gnd.n826 gnd.n825 9.3005
R15818 gnd.n6977 gnd.n6976 9.3005
R15819 gnd.n6979 gnd.n6978 9.3005
R15820 gnd.n818 gnd.n817 9.3005
R15821 gnd.n6985 gnd.n6984 9.3005
R15822 gnd.n6987 gnd.n6986 9.3005
R15823 gnd.n810 gnd.n809 9.3005
R15824 gnd.n6993 gnd.n6992 9.3005
R15825 gnd.n6995 gnd.n6994 9.3005
R15826 gnd.n802 gnd.n801 9.3005
R15827 gnd.n7001 gnd.n7000 9.3005
R15828 gnd.n7003 gnd.n7002 9.3005
R15829 gnd.n794 gnd.n793 9.3005
R15830 gnd.n7009 gnd.n7008 9.3005
R15831 gnd.n6971 gnd.n6970 9.3005
R15832 gnd.n1005 gnd.n831 9.3005
R15833 gnd.n1019 gnd.n1002 9.3005
R15834 gnd.n1021 gnd.n1020 9.3005
R15835 gnd.n1022 gnd.n1001 9.3005
R15836 gnd.n1026 gnd.n1025 9.3005
R15837 gnd.n1027 gnd.n998 9.3005
R15838 gnd.n1029 gnd.n1028 9.3005
R15839 gnd.n1031 gnd.n995 9.3005
R15840 gnd.n1035 gnd.n1034 9.3005
R15841 gnd.n1036 gnd.n994 9.3005
R15842 gnd.n6709 gnd.n6708 9.3005
R15843 gnd.n5823 gnd.n1665 9.3005
R15844 gnd.n5825 gnd.n5824 9.3005
R15845 gnd.n1654 gnd.n1653 9.3005
R15846 gnd.n5842 gnd.n5841 9.3005
R15847 gnd.n5843 gnd.n1652 9.3005
R15848 gnd.n5845 gnd.n5844 9.3005
R15849 gnd.n1640 gnd.n1639 9.3005
R15850 gnd.n5864 gnd.n5863 9.3005
R15851 gnd.n5865 gnd.n1637 9.3005
R15852 gnd.n5872 gnd.n5871 9.3005
R15853 gnd.n5870 gnd.n1638 9.3005
R15854 gnd.n5869 gnd.n5868 9.3005
R15855 gnd.n5867 gnd.n5866 9.3005
R15856 gnd.n1413 gnd.n1412 9.3005
R15857 gnd.n6084 gnd.n6083 9.3005
R15858 gnd.n6085 gnd.n1410 9.3005
R15859 gnd.n6121 gnd.n6120 9.3005
R15860 gnd.n6119 gnd.n1411 9.3005
R15861 gnd.n6118 gnd.n6117 9.3005
R15862 gnd.n6116 gnd.n6086 9.3005
R15863 gnd.n6115 gnd.n6114 9.3005
R15864 gnd.n6113 gnd.n6089 9.3005
R15865 gnd.n6112 gnd.n6111 9.3005
R15866 gnd.n6110 gnd.n6090 9.3005
R15867 gnd.n6109 gnd.n6108 9.3005
R15868 gnd.n1336 gnd.n1335 9.3005
R15869 gnd.n6231 gnd.n6230 9.3005
R15870 gnd.n6232 gnd.n1333 9.3005
R15871 gnd.n6247 gnd.n6246 9.3005
R15872 gnd.n6245 gnd.n1334 9.3005
R15873 gnd.n6244 gnd.n6243 9.3005
R15874 gnd.n6242 gnd.n6233 9.3005
R15875 gnd.n6241 gnd.n6240 9.3005
R15876 gnd.n6239 gnd.n6237 9.3005
R15877 gnd.n6238 gnd.n1277 9.3005
R15878 gnd.n6342 gnd.n1276 9.3005
R15879 gnd.n6344 gnd.n6343 9.3005
R15880 gnd.n6345 gnd.n1274 9.3005
R15881 gnd.n6380 gnd.n6379 9.3005
R15882 gnd.n6378 gnd.n1275 9.3005
R15883 gnd.n6377 gnd.n6376 9.3005
R15884 gnd.n6375 gnd.n6346 9.3005
R15885 gnd.n6374 gnd.n6373 9.3005
R15886 gnd.n6372 gnd.n6348 9.3005
R15887 gnd.n6371 gnd.n6370 9.3005
R15888 gnd.n6369 gnd.n6349 9.3005
R15889 gnd.n6368 gnd.n6367 9.3005
R15890 gnd.n6366 gnd.n6352 9.3005
R15891 gnd.n6365 gnd.n6364 9.3005
R15892 gnd.n6363 gnd.n6353 9.3005
R15893 gnd.n6362 gnd.n6361 9.3005
R15894 gnd.n6360 gnd.n6359 9.3005
R15895 gnd.n1088 gnd.n1087 9.3005
R15896 gnd.n6634 gnd.n6633 9.3005
R15897 gnd.n6635 gnd.n1085 9.3005
R15898 gnd.n6638 gnd.n6637 9.3005
R15899 gnd.n6636 gnd.n1086 9.3005
R15900 gnd.n1063 gnd.n1062 9.3005
R15901 gnd.n6664 gnd.n6663 9.3005
R15902 gnd.n6665 gnd.n1060 9.3005
R15903 gnd.n6669 gnd.n6668 9.3005
R15904 gnd.n6667 gnd.n1061 9.3005
R15905 gnd.n6666 gnd.n1038 9.3005
R15906 gnd.n6705 gnd.n1037 9.3005
R15907 gnd.n6707 gnd.n6706 9.3005
R15908 gnd.n5822 gnd.n5821 9.3005
R15909 gnd.n5750 gnd.n5749 9.3005
R15910 gnd.n5751 gnd.n5740 9.3005
R15911 gnd.n5753 gnd.n5752 9.3005
R15912 gnd.n5754 gnd.n5739 9.3005
R15913 gnd.n5756 gnd.n5755 9.3005
R15914 gnd.n5757 gnd.n5734 9.3005
R15915 gnd.n5759 gnd.n5758 9.3005
R15916 gnd.n5760 gnd.n1753 9.3005
R15917 gnd.n5762 gnd.n5761 9.3005
R15918 gnd.n5748 gnd.n1666 9.3005
R15919 gnd.n5412 gnd.n5411 9.3005
R15920 gnd.n5415 gnd.n1896 9.3005
R15921 gnd.n5417 gnd.n5416 9.3005
R15922 gnd.n5418 gnd.n1894 9.3005
R15923 gnd.n5594 gnd.n5593 9.3005
R15924 gnd.n5592 gnd.n1895 9.3005
R15925 gnd.n5591 gnd.n5590 9.3005
R15926 gnd.n5589 gnd.n5419 9.3005
R15927 gnd.n5588 gnd.n5587 9.3005
R15928 gnd.n5586 gnd.n5422 9.3005
R15929 gnd.n5585 gnd.n5584 9.3005
R15930 gnd.n5583 gnd.n5423 9.3005
R15931 gnd.n5582 gnd.n5581 9.3005
R15932 gnd.n5580 gnd.n5426 9.3005
R15933 gnd.n5579 gnd.n5578 9.3005
R15934 gnd.n5577 gnd.n5427 9.3005
R15935 gnd.n5576 gnd.n5575 9.3005
R15936 gnd.n5574 gnd.n5430 9.3005
R15937 gnd.n5573 gnd.n5572 9.3005
R15938 gnd.n5571 gnd.n5431 9.3005
R15939 gnd.n1757 gnd.n1756 9.3005
R15940 gnd.n5724 gnd.n5723 9.3005
R15941 gnd.n5725 gnd.n1755 9.3005
R15942 gnd.n5727 gnd.n5726 9.3005
R15943 gnd.n5730 gnd.n1754 9.3005
R15944 gnd.n5732 gnd.n5731 9.3005
R15945 gnd.n5763 gnd.n1748 9.3005
R15946 gnd.n5765 gnd.n5764 9.3005
R15947 gnd.n1742 gnd.n1741 9.3005
R15948 gnd.n5773 gnd.n5772 9.3005
R15949 gnd.n5775 gnd.n5774 9.3005
R15950 gnd.n1732 gnd.n1731 9.3005
R15951 gnd.n5781 gnd.n5780 9.3005
R15952 gnd.n5783 gnd.n5782 9.3005
R15953 gnd.n1719 gnd.n1718 9.3005
R15954 gnd.n5789 gnd.n5788 9.3005
R15955 gnd.n5791 gnd.n5790 9.3005
R15956 gnd.n1709 gnd.n1708 9.3005
R15957 gnd.n5797 gnd.n5796 9.3005
R15958 gnd.n5799 gnd.n5798 9.3005
R15959 gnd.n1693 gnd.n1691 9.3005
R15960 gnd.n5805 gnd.n5804 9.3005
R15961 gnd.n5806 gnd.n1690 9.3005
R15962 gnd.n1696 gnd.n1620 9.3005
R15963 gnd.n1694 gnd.n1692 9.3005
R15964 gnd.n5803 gnd.n5802 9.3005
R15965 gnd.n5801 gnd.n5800 9.3005
R15966 gnd.n1704 gnd.n1703 9.3005
R15967 gnd.n5795 gnd.n5794 9.3005
R15968 gnd.n5793 gnd.n5792 9.3005
R15969 gnd.n1715 gnd.n1714 9.3005
R15970 gnd.n5787 gnd.n5786 9.3005
R15971 gnd.n5785 gnd.n5784 9.3005
R15972 gnd.n1726 gnd.n1725 9.3005
R15973 gnd.n5779 gnd.n5778 9.3005
R15974 gnd.n5777 gnd.n5776 9.3005
R15975 gnd.n1738 gnd.n1737 9.3005
R15976 gnd.n5771 gnd.n5770 9.3005
R15977 gnd.n5769 gnd.n5766 9.3005
R15978 gnd.n5894 gnd.n1621 9.3005
R15979 gnd.n5893 gnd.n5892 9.3005
R15980 gnd.n5891 gnd.n1625 9.3005
R15981 gnd.n5890 gnd.n5889 9.3005
R15982 gnd.n5888 gnd.n1626 9.3005
R15983 gnd.n5887 gnd.n5886 9.3005
R15984 gnd.n5885 gnd.n1630 9.3005
R15985 gnd.n5884 gnd.n5883 9.3005
R15986 gnd.n5882 gnd.n1631 9.3005
R15987 gnd.n5881 gnd.n5880 9.3005
R15988 gnd.n5879 gnd.n5878 9.3005
R15989 gnd.n1421 gnd.n1420 9.3005
R15990 gnd.n6075 gnd.n6074 9.3005
R15991 gnd.n6076 gnd.n1418 9.3005
R15992 gnd.n6079 gnd.n6078 9.3005
R15993 gnd.n6077 gnd.n1419 9.3005
R15994 gnd.n1389 gnd.n1388 9.3005
R15995 gnd.n6155 gnd.n6154 9.3005
R15996 gnd.n6156 gnd.n1386 9.3005
R15997 gnd.n6159 gnd.n6158 9.3005
R15998 gnd.n6157 gnd.n1387 9.3005
R15999 gnd.n1357 gnd.n1356 9.3005
R16000 gnd.n6206 gnd.n6205 9.3005
R16001 gnd.n6207 gnd.n1354 9.3005
R16002 gnd.n6210 gnd.n6209 9.3005
R16003 gnd.n6208 gnd.n1355 9.3005
R16004 gnd.n1321 gnd.n1320 9.3005
R16005 gnd.n6272 gnd.n6271 9.3005
R16006 gnd.n6273 gnd.n1318 9.3005
R16007 gnd.n6279 gnd.n6278 9.3005
R16008 gnd.n6277 gnd.n1319 9.3005
R16009 gnd.n6276 gnd.n6275 9.3005
R16010 gnd.n1283 gnd.n1282 9.3005
R16011 gnd.n6335 gnd.n6334 9.3005
R16012 gnd.n6336 gnd.n1281 9.3005
R16013 gnd.n6338 gnd.n6337 9.3005
R16014 gnd.n1253 gnd.n1252 9.3005
R16015 gnd.n6404 gnd.n6403 9.3005
R16016 gnd.n6405 gnd.n1251 9.3005
R16017 gnd.n6407 gnd.n6406 9.3005
R16018 gnd.n1225 gnd.n1224 9.3005
R16019 gnd.n6440 gnd.n6439 9.3005
R16020 gnd.n6441 gnd.n1223 9.3005
R16021 gnd.n6443 gnd.n6442 9.3005
R16022 gnd.n1197 gnd.n1196 9.3005
R16023 gnd.n6477 gnd.n6476 9.3005
R16024 gnd.n6478 gnd.n1194 9.3005
R16025 gnd.n6484 gnd.n6483 9.3005
R16026 gnd.n6482 gnd.n1195 9.3005
R16027 gnd.n6481 gnd.n6480 9.3005
R16028 gnd.n1097 gnd.n1096 9.3005
R16029 gnd.n6625 gnd.n6624 9.3005
R16030 gnd.n6626 gnd.n1094 9.3005
R16031 gnd.n6629 gnd.n6628 9.3005
R16032 gnd.n6627 gnd.n1095 9.3005
R16033 gnd.n1072 gnd.n1071 9.3005
R16034 gnd.n6655 gnd.n6654 9.3005
R16035 gnd.n6656 gnd.n1069 9.3005
R16036 gnd.n6659 gnd.n6658 9.3005
R16037 gnd.n6657 gnd.n1070 9.3005
R16038 gnd.n1047 gnd.n1046 9.3005
R16039 gnd.n6697 gnd.n6696 9.3005
R16040 gnd.n6698 gnd.n1044 9.3005
R16041 gnd.n6701 gnd.n6700 9.3005
R16042 gnd.n6699 gnd.n1045 9.3005
R16043 gnd.n5896 gnd.n5895 9.3005
R16044 gnd.n777 gnd.n776 9.3005
R16045 gnd.n7026 gnd.n7025 9.3005
R16046 gnd.n7027 gnd.n775 9.3005
R16047 gnd.n7029 gnd.n7028 9.3005
R16048 gnd.n759 gnd.n758 9.3005
R16049 gnd.n7042 gnd.n7041 9.3005
R16050 gnd.n7043 gnd.n757 9.3005
R16051 gnd.n7045 gnd.n7044 9.3005
R16052 gnd.n741 gnd.n740 9.3005
R16053 gnd.n7058 gnd.n7057 9.3005
R16054 gnd.n7059 gnd.n739 9.3005
R16055 gnd.n7061 gnd.n7060 9.3005
R16056 gnd.n724 gnd.n723 9.3005
R16057 gnd.n7074 gnd.n7073 9.3005
R16058 gnd.n7075 gnd.n722 9.3005
R16059 gnd.n7077 gnd.n7076 9.3005
R16060 gnd.n706 gnd.n705 9.3005
R16061 gnd.n7091 gnd.n7090 9.3005
R16062 gnd.n7092 gnd.n704 9.3005
R16063 gnd.n7094 gnd.n7093 9.3005
R16064 gnd.n689 gnd.n688 9.3005
R16065 gnd.n7107 gnd.n7106 9.3005
R16066 gnd.n7108 gnd.n687 9.3005
R16067 gnd.n7110 gnd.n7109 9.3005
R16068 gnd.n673 gnd.n672 9.3005
R16069 gnd.n7123 gnd.n7122 9.3005
R16070 gnd.n7124 gnd.n670 9.3005
R16071 gnd.n7126 gnd.n7125 9.3005
R16072 gnd.n658 gnd.n657 9.3005
R16073 gnd.n7138 gnd.n7137 9.3005
R16074 gnd.n7139 gnd.n656 9.3005
R16075 gnd.n7141 gnd.n7140 9.3005
R16076 gnd.n641 gnd.n640 9.3005
R16077 gnd.n7154 gnd.n7153 9.3005
R16078 gnd.n7155 gnd.n639 9.3005
R16079 gnd.n7157 gnd.n7156 9.3005
R16080 gnd.n624 gnd.n623 9.3005
R16081 gnd.n7170 gnd.n7169 9.3005
R16082 gnd.n7171 gnd.n622 9.3005
R16083 gnd.n7173 gnd.n7172 9.3005
R16084 gnd.n608 gnd.n607 9.3005
R16085 gnd.n7186 gnd.n7185 9.3005
R16086 gnd.n7187 gnd.n606 9.3005
R16087 gnd.n7189 gnd.n7188 9.3005
R16088 gnd.n591 gnd.n590 9.3005
R16089 gnd.n7202 gnd.n7201 9.3005
R16090 gnd.n7203 gnd.n588 9.3005
R16091 gnd.n7273 gnd.n7272 9.3005
R16092 gnd.n7271 gnd.n589 9.3005
R16093 gnd.n7270 gnd.n7269 9.3005
R16094 gnd.n7268 gnd.n7204 9.3005
R16095 gnd.n7267 gnd.n7266 9.3005
R16096 gnd.n7013 gnd.n7012 9.3005
R16097 gnd.n7263 gnd.n7206 9.3005
R16098 gnd.n7262 gnd.n7261 9.3005
R16099 gnd.n7260 gnd.n7211 9.3005
R16100 gnd.n7259 gnd.n7258 9.3005
R16101 gnd.n7257 gnd.n7212 9.3005
R16102 gnd.n7256 gnd.n7255 9.3005
R16103 gnd.n7254 gnd.n7219 9.3005
R16104 gnd.n7253 gnd.n7252 9.3005
R16105 gnd.n7251 gnd.n7220 9.3005
R16106 gnd.n7250 gnd.n7249 9.3005
R16107 gnd.n7248 gnd.n7227 9.3005
R16108 gnd.n7247 gnd.n7246 9.3005
R16109 gnd.n7245 gnd.n7228 9.3005
R16110 gnd.n7244 gnd.n7243 9.3005
R16111 gnd.n7242 gnd.n7239 9.3005
R16112 gnd.n7241 gnd.n7240 9.3005
R16113 gnd.n7265 gnd.n7264 9.3005
R16114 gnd.n1015 gnd.n1012 9.3005
R16115 gnd.n911 gnd.n909 9.3005
R16116 gnd.n6890 gnd.n6889 9.3005
R16117 gnd.n6888 gnd.n910 9.3005
R16118 gnd.n6887 gnd.n6886 9.3005
R16119 gnd.n6885 gnd.n912 9.3005
R16120 gnd.n6884 gnd.n6883 9.3005
R16121 gnd.n6882 gnd.n915 9.3005
R16122 gnd.n6881 gnd.n6880 9.3005
R16123 gnd.n6879 gnd.n916 9.3005
R16124 gnd.n6878 gnd.n6877 9.3005
R16125 gnd.n6876 gnd.n919 9.3005
R16126 gnd.n6875 gnd.n6874 9.3005
R16127 gnd.n6873 gnd.n920 9.3005
R16128 gnd.n6872 gnd.n6871 9.3005
R16129 gnd.n6870 gnd.n923 9.3005
R16130 gnd.n6869 gnd.n6868 9.3005
R16131 gnd.n6867 gnd.n924 9.3005
R16132 gnd.n6866 gnd.n6865 9.3005
R16133 gnd.n6864 gnd.n927 9.3005
R16134 gnd.n6863 gnd.n6862 9.3005
R16135 gnd.n6861 gnd.n928 9.3005
R16136 gnd.n6860 gnd.n6859 9.3005
R16137 gnd.n6858 gnd.n6857 9.3005
R16138 gnd.n6856 gnd.n465 9.3005
R16139 gnd.n7394 gnd.n466 9.3005
R16140 gnd.n7393 gnd.n7392 9.3005
R16141 gnd.n7391 gnd.n467 9.3005
R16142 gnd.n7390 gnd.n7389 9.3005
R16143 gnd.n7388 gnd.n471 9.3005
R16144 gnd.n7387 gnd.n7386 9.3005
R16145 gnd.n7385 gnd.n472 9.3005
R16146 gnd.n7384 gnd.n7383 9.3005
R16147 gnd.n7382 gnd.n476 9.3005
R16148 gnd.n7381 gnd.n7380 9.3005
R16149 gnd.n7379 gnd.n477 9.3005
R16150 gnd.n7378 gnd.n7377 9.3005
R16151 gnd.n7376 gnd.n481 9.3005
R16152 gnd.n7375 gnd.n7374 9.3005
R16153 gnd.n7373 gnd.n482 9.3005
R16154 gnd.n7372 gnd.n7371 9.3005
R16155 gnd.n7370 gnd.n486 9.3005
R16156 gnd.n7369 gnd.n7368 9.3005
R16157 gnd.n7367 gnd.n487 9.3005
R16158 gnd.n7366 gnd.n7365 9.3005
R16159 gnd.n7364 gnd.n491 9.3005
R16160 gnd.n7363 gnd.n7362 9.3005
R16161 gnd.n7361 gnd.n492 9.3005
R16162 gnd.n7360 gnd.n7359 9.3005
R16163 gnd.n7358 gnd.n496 9.3005
R16164 gnd.n7357 gnd.n7356 9.3005
R16165 gnd.n7355 gnd.n497 9.3005
R16166 gnd.n1017 gnd.n1016 9.3005
R16167 gnd.n125 gnd.n124 9.3005
R16168 gnd.n98 gnd.n97 9.3005
R16169 gnd.n119 gnd.n118 9.3005
R16170 gnd.n117 gnd.n116 9.3005
R16171 gnd.n102 gnd.n101 9.3005
R16172 gnd.n111 gnd.n110 9.3005
R16173 gnd.n109 gnd.n108 9.3005
R16174 gnd.n93 gnd.n92 9.3005
R16175 gnd.n66 gnd.n65 9.3005
R16176 gnd.n87 gnd.n86 9.3005
R16177 gnd.n85 gnd.n84 9.3005
R16178 gnd.n70 gnd.n69 9.3005
R16179 gnd.n79 gnd.n78 9.3005
R16180 gnd.n77 gnd.n76 9.3005
R16181 gnd.n61 gnd.n60 9.3005
R16182 gnd.n34 gnd.n33 9.3005
R16183 gnd.n55 gnd.n54 9.3005
R16184 gnd.n53 gnd.n52 9.3005
R16185 gnd.n38 gnd.n37 9.3005
R16186 gnd.n47 gnd.n46 9.3005
R16187 gnd.n45 gnd.n44 9.3005
R16188 gnd.n30 gnd.n29 9.3005
R16189 gnd.n3 gnd.n2 9.3005
R16190 gnd.n24 gnd.n23 9.3005
R16191 gnd.n22 gnd.n21 9.3005
R16192 gnd.n7 gnd.n6 9.3005
R16193 gnd.n16 gnd.n15 9.3005
R16194 gnd.n14 gnd.n13 9.3005
R16195 gnd.n252 gnd.n251 9.3005
R16196 gnd.n225 gnd.n224 9.3005
R16197 gnd.n246 gnd.n245 9.3005
R16198 gnd.n244 gnd.n243 9.3005
R16199 gnd.n229 gnd.n228 9.3005
R16200 gnd.n238 gnd.n237 9.3005
R16201 gnd.n236 gnd.n235 9.3005
R16202 gnd.n220 gnd.n219 9.3005
R16203 gnd.n193 gnd.n192 9.3005
R16204 gnd.n214 gnd.n213 9.3005
R16205 gnd.n212 gnd.n211 9.3005
R16206 gnd.n197 gnd.n196 9.3005
R16207 gnd.n206 gnd.n205 9.3005
R16208 gnd.n204 gnd.n203 9.3005
R16209 gnd.n188 gnd.n187 9.3005
R16210 gnd.n161 gnd.n160 9.3005
R16211 gnd.n182 gnd.n181 9.3005
R16212 gnd.n180 gnd.n179 9.3005
R16213 gnd.n165 gnd.n164 9.3005
R16214 gnd.n174 gnd.n173 9.3005
R16215 gnd.n172 gnd.n171 9.3005
R16216 gnd.n157 gnd.n156 9.3005
R16217 gnd.n130 gnd.n129 9.3005
R16218 gnd.n151 gnd.n150 9.3005
R16219 gnd.n149 gnd.n148 9.3005
R16220 gnd.n134 gnd.n133 9.3005
R16221 gnd.n143 gnd.n142 9.3005
R16222 gnd.n141 gnd.n140 9.3005
R16223 gnd.n7395 gnd.n464 9.29925
R16224 gnd.n4336 gnd.n4335 9.0033
R16225 gnd.t225 gnd.n3777 8.99777
R16226 gnd.t54 gnd.n1791 8.99777
R16227 gnd.t68 gnd.n743 8.99777
R16228 gnd.n4293 gnd.n4268 8.92171
R16229 gnd.n4330 gnd.n4305 8.92171
R16230 gnd.n4154 gnd.n4129 8.92171
R16231 gnd.n4191 gnd.n4166 8.92171
R16232 gnd.n4223 gnd.n4198 8.92171
R16233 gnd.n4260 gnd.n4235 8.92171
R16234 gnd.n459 gnd.n434 8.92171
R16235 gnd.n422 gnd.n397 8.92171
R16236 gnd.n320 gnd.n295 8.92171
R16237 gnd.n283 gnd.n258 8.92171
R16238 gnd.n389 gnd.n364 8.92171
R16239 gnd.n352 gnd.n327 8.92171
R16240 gnd.n4996 gnd.n4971 8.92171
R16241 gnd.n4964 gnd.n4939 8.92171
R16242 gnd.n4932 gnd.n4907 8.92171
R16243 gnd.n4901 gnd.n4876 8.92171
R16244 gnd.n4869 gnd.n4844 8.92171
R16245 gnd.n4837 gnd.n4812 8.92171
R16246 gnd.n4805 gnd.n4780 8.92171
R16247 gnd.n4774 gnd.n4749 8.92171
R16248 gnd.n123 gnd.n98 8.92171
R16249 gnd.n91 gnd.n66 8.92171
R16250 gnd.n59 gnd.n34 8.92171
R16251 gnd.n28 gnd.n3 8.92171
R16252 gnd.n250 gnd.n225 8.92171
R16253 gnd.n218 gnd.n193 8.92171
R16254 gnd.n186 gnd.n161 8.92171
R16255 gnd.n155 gnd.n130 8.92171
R16256 gnd.n1133 gnd.n1115 8.72777
R16257 gnd.n6164 gnd.n6163 8.66454
R16258 gnd.n6250 gnd.n1326 8.66454
R16259 gnd.n1279 gnd.n1263 8.66454
R16260 gnd.n6466 gnd.n1199 8.66454
R16261 gnd.n5410 gnd.n0 8.41206
R16262 gnd.n7395 gnd.n7394 8.41206
R16263 gnd.n4533 gnd.t17 8.33131
R16264 gnd.t13 gnd.n1314 8.33131
R16265 gnd.n6325 gnd.t37 8.33131
R16266 gnd.n4294 gnd.n4266 8.14595
R16267 gnd.n4331 gnd.n4303 8.14595
R16268 gnd.n4155 gnd.n4127 8.14595
R16269 gnd.n4192 gnd.n4164 8.14595
R16270 gnd.n4224 gnd.n4196 8.14595
R16271 gnd.n4261 gnd.n4233 8.14595
R16272 gnd.n460 gnd.n432 8.14595
R16273 gnd.n423 gnd.n395 8.14595
R16274 gnd.n321 gnd.n293 8.14595
R16275 gnd.n284 gnd.n256 8.14595
R16276 gnd.n390 gnd.n362 8.14595
R16277 gnd.n353 gnd.n325 8.14595
R16278 gnd.n4997 gnd.n4969 8.14595
R16279 gnd.n4965 gnd.n4937 8.14595
R16280 gnd.n4933 gnd.n4905 8.14595
R16281 gnd.n4902 gnd.n4874 8.14595
R16282 gnd.n4870 gnd.n4842 8.14595
R16283 gnd.n4838 gnd.n4810 8.14595
R16284 gnd.n4806 gnd.n4778 8.14595
R16285 gnd.n4775 gnd.n4747 8.14595
R16286 gnd.n124 gnd.n96 8.14595
R16287 gnd.n92 gnd.n64 8.14595
R16288 gnd.n60 gnd.n32 8.14595
R16289 gnd.n29 gnd.n1 8.14595
R16290 gnd.n251 gnd.n223 8.14595
R16291 gnd.n219 gnd.n191 8.14595
R16292 gnd.n187 gnd.n159 8.14595
R16293 gnd.n156 gnd.n128 8.14595
R16294 gnd.n4265 gnd.n4195 8.05588
R16295 gnd.n394 gnd.n324 8.05588
R16296 gnd.n6142 gnd.t167 7.99808
R16297 gnd.n6123 gnd.t167 7.99808
R16298 gnd.t120 gnd.n6124 7.99808
R16299 gnd.n6164 gnd.n1380 7.99808
R16300 gnd.t8 gnd.n6212 7.99808
R16301 gnd.n6250 gnd.n6249 7.99808
R16302 gnd.n6340 gnd.n1279 7.99808
R16303 gnd.t21 gnd.n6409 7.99808
R16304 gnd.n6474 gnd.n1199 7.99808
R16305 gnd.n5002 gnd.n5001 7.97301
R16306 gnd.n7240 gnd.n7239 7.75808
R16307 gnd.n6970 gnd.n831 7.75808
R16308 gnd.n5770 gnd.n5769 7.75808
R16309 gnd.n5245 gnd.n2037 7.75808
R16310 gnd.t10 gnd.n4482 7.66484
R16311 gnd.n4441 gnd.n4440 7.33161
R16312 gnd.n4452 gnd.n3887 7.33161
R16313 gnd.n4451 gnd.n3890 7.33161
R16314 gnd.n4462 gnd.n3880 7.33161
R16315 gnd.n4360 gnd.n3873 7.33161
R16316 gnd.n4472 gnd.n4471 7.33161
R16317 gnd.n4483 gnd.n3862 7.33161
R16318 gnd.n4482 gnd.n3865 7.33161
R16319 gnd.n4493 gnd.n3853 7.33161
R16320 gnd.n3856 gnd.n3854 7.33161
R16321 gnd.n4503 gnd.n4502 7.33161
R16322 gnd.n4514 gnd.n3836 7.33161
R16323 gnd.n4524 gnd.n3827 7.33161
R16324 gnd.n3830 gnd.n3828 7.33161
R16325 gnd.n4534 gnd.n4533 7.33161
R16326 gnd.n4545 gnd.n3810 7.33161
R16327 gnd.n4555 gnd.n3802 7.33161
R16328 gnd.n3803 gnd.n3795 7.33161
R16329 gnd.n4576 gnd.n3784 7.33161
R16330 gnd.n4575 gnd.n3787 7.33161
R16331 gnd.n4586 gnd.n3777 7.33161
R16332 gnd.n4114 gnd.n3770 7.33161
R16333 gnd.n4596 gnd.n4595 7.33161
R16334 gnd.n4607 gnd.n3759 7.33161
R16335 gnd.n4606 gnd.n3762 7.33161
R16336 gnd.n3752 gnd.n3745 7.33161
R16337 gnd.n4627 gnd.n4626 7.33161
R16338 gnd.n4637 gnd.n3732 7.33161
R16339 gnd.n4636 gnd.n3735 7.33161
R16340 gnd.n4645 gnd.n3726 7.33161
R16341 gnd.n4657 gnd.n3717 7.33161
R16342 gnd.n4679 gnd.n3710 7.33161
R16343 gnd.n3703 gnd.n3535 7.33161
R16344 gnd.n5158 gnd.n3537 7.33161
R16345 gnd.n4669 gnd.n3546 7.33161
R16346 gnd.n5152 gnd.n5151 7.33161
R16347 gnd.n4716 gnd.n4715 7.33161
R16348 gnd.n5145 gnd.n3557 7.33161
R16349 gnd.n4737 gnd.n3568 7.33161
R16350 gnd.n5138 gnd.n5137 7.33161
R16351 gnd.n4731 gnd.n4730 7.33161
R16352 gnd.n5131 gnd.n3581 7.33161
R16353 gnd.n5130 gnd.n3584 7.33161
R16354 gnd.n5023 gnd.n5022 7.33161
R16355 gnd.n5124 gnd.n5123 7.33161
R16356 gnd.n5016 gnd.n5015 7.33161
R16357 gnd.n5117 gnd.n3604 7.33161
R16358 gnd.n6096 gnd.n1366 7.33161
R16359 gnd.n1343 gnd.n1338 7.33161
R16360 gnd.n6400 gnd.n1258 7.33161
R16361 gnd.n6420 gnd.n1220 7.33161
R16362 gnd.n6460 gnd.t139 7.33161
R16363 gnd.t114 gnd.n6493 7.33161
R16364 gnd.n1484 gnd.n1483 7.30353
R16365 gnd.n1132 gnd.n1131 7.30353
R16366 gnd.n3856 gnd.t22 6.99838
R16367 gnd.n4627 gnd.t39 6.99838
R16368 gnd.n4738 gnd.t227 6.99838
R16369 gnd.n1495 gnd.n1425 6.66515
R16370 gnd.n6125 gnd.n6123 6.66515
R16371 gnd.n6259 gnd.n1304 6.66515
R16372 gnd.n6332 gnd.n6331 6.66515
R16373 gnd.n6487 gnd.n6486 6.66515
R16374 gnd.n6547 gnd.n1161 6.5566
R16375 gnd.n1552 gnd.n1492 6.5566
R16376 gnd.n6007 gnd.n6006 6.5566
R16377 gnd.n6558 gnd.n1156 6.5566
R16378 gnd.n4544 gnd.t43 6.33191
R16379 gnd.n3813 gnd.t9 6.33191
R16380 gnd.n4114 gnd.t33 6.33191
R16381 gnd.t16 gnd.n3701 6.33191
R16382 gnd.n6249 gnd.t13 6.33191
R16383 gnd.n6340 gnd.t37 6.33191
R16384 gnd.n7320 gnd.n537 6.20656
R16385 gnd.n2124 gnd.n2070 6.20656
R16386 gnd.n6202 gnd.n1362 5.99868
R16387 gnd.n6213 gnd.n1348 5.99868
R16388 gnd.n6410 gnd.n1234 5.99868
R16389 gnd.n6426 gnd.n1227 5.99868
R16390 gnd.n4296 gnd.n4266 5.81868
R16391 gnd.n4333 gnd.n4303 5.81868
R16392 gnd.n4157 gnd.n4127 5.81868
R16393 gnd.n4194 gnd.n4164 5.81868
R16394 gnd.n4226 gnd.n4196 5.81868
R16395 gnd.n4263 gnd.n4233 5.81868
R16396 gnd.n462 gnd.n432 5.81868
R16397 gnd.n425 gnd.n395 5.81868
R16398 gnd.n323 gnd.n293 5.81868
R16399 gnd.n286 gnd.n256 5.81868
R16400 gnd.n392 gnd.n362 5.81868
R16401 gnd.n355 gnd.n325 5.81868
R16402 gnd.n4999 gnd.n4969 5.81868
R16403 gnd.n4967 gnd.n4937 5.81868
R16404 gnd.n4935 gnd.n4905 5.81868
R16405 gnd.n4904 gnd.n4874 5.81868
R16406 gnd.n4872 gnd.n4842 5.81868
R16407 gnd.n4840 gnd.n4810 5.81868
R16408 gnd.n4808 gnd.n4778 5.81868
R16409 gnd.n4777 gnd.n4747 5.81868
R16410 gnd.n126 gnd.n96 5.81868
R16411 gnd.n94 gnd.n64 5.81868
R16412 gnd.n62 gnd.n32 5.81868
R16413 gnd.n31 gnd.n1 5.81868
R16414 gnd.n253 gnd.n223 5.81868
R16415 gnd.n221 gnd.n191 5.81868
R16416 gnd.n189 gnd.n159 5.81868
R16417 gnd.n158 gnd.n128 5.81868
R16418 gnd.n4596 gnd.t226 5.66545
R16419 gnd.n4617 gnd.t23 5.66545
R16420 gnd.t35 gnd.n4693 5.66545
R16421 gnd.t0 gnd.n1634 5.66545
R16422 gnd.n6641 gnd.t218 5.66545
R16423 gnd.n6549 gnd.n877 5.62001
R16424 gnd.n5999 gnd.n1556 5.62001
R16425 gnd.n6002 gnd.n5999 5.62001
R16426 gnd.n6556 gnd.n877 5.62001
R16427 gnd.n5752 gnd.n5743 5.4308
R16428 gnd.n3984 gnd.n3983 5.4308
R16429 gnd.n5038 gnd.n3676 5.4308
R16430 gnd.n1031 gnd.n1030 5.4308
R16431 gnd.n1307 gnd.n1306 5.33222
R16432 gnd.n6310 gnd.n1300 5.33222
R16433 gnd.n6495 gnd.n1109 5.33222
R16434 gnd.n1182 gnd.t176 5.33222
R16435 gnd.n4294 gnd.n4293 5.04292
R16436 gnd.n4331 gnd.n4330 5.04292
R16437 gnd.n4155 gnd.n4154 5.04292
R16438 gnd.n4192 gnd.n4191 5.04292
R16439 gnd.n4224 gnd.n4223 5.04292
R16440 gnd.n4261 gnd.n4260 5.04292
R16441 gnd.n460 gnd.n459 5.04292
R16442 gnd.n423 gnd.n422 5.04292
R16443 gnd.n321 gnd.n320 5.04292
R16444 gnd.n284 gnd.n283 5.04292
R16445 gnd.n390 gnd.n389 5.04292
R16446 gnd.n353 gnd.n352 5.04292
R16447 gnd.n4997 gnd.n4996 5.04292
R16448 gnd.n4965 gnd.n4964 5.04292
R16449 gnd.n4933 gnd.n4932 5.04292
R16450 gnd.n4902 gnd.n4901 5.04292
R16451 gnd.n4870 gnd.n4869 5.04292
R16452 gnd.n4838 gnd.n4837 5.04292
R16453 gnd.n4806 gnd.n4805 5.04292
R16454 gnd.n4775 gnd.n4774 5.04292
R16455 gnd.n124 gnd.n123 5.04292
R16456 gnd.n92 gnd.n91 5.04292
R16457 gnd.n60 gnd.n59 5.04292
R16458 gnd.n29 gnd.n28 5.04292
R16459 gnd.n251 gnd.n250 5.04292
R16460 gnd.n219 gnd.n218 5.04292
R16461 gnd.n187 gnd.n186 5.04292
R16462 gnd.n156 gnd.n155 5.04292
R16463 gnd.n4565 gnd.t19 4.99899
R16464 gnd.n4645 gnd.t221 4.99899
R16465 gnd.t124 gnd.n1996 4.99899
R16466 gnd.n1102 gnd.t194 4.99899
R16467 gnd.n585 gnd.t160 4.99899
R16468 gnd.n4335 gnd.n4334 4.82753
R16469 gnd.n464 gnd.n463 4.82753
R16470 gnd.n4339 gnd.n4338 4.74817
R16471 gnd.n4126 gnd.n4122 4.74817
R16472 gnd.n4119 gnd.n4118 4.74817
R16473 gnd.n4113 gnd.n4092 4.74817
R16474 gnd.n4338 gnd.n4090 4.74817
R16475 gnd.n4126 gnd.n4125 4.74817
R16476 gnd.n4121 gnd.n4119 4.74817
R16477 gnd.n4117 gnd.n4092 4.74817
R16478 gnd.n7102 gnd.n7100 4.74817
R16479 gnd.n7114 gnd.n680 4.74817
R16480 gnd.n7118 gnd.n7116 4.74817
R16481 gnd.n7130 gnd.n665 4.74817
R16482 gnd.n7133 gnd.n7132 4.74817
R16483 gnd.n7100 gnd.n7099 4.74817
R16484 gnd.n7101 gnd.n680 4.74817
R16485 gnd.n7116 gnd.n7115 4.74817
R16486 gnd.n7117 gnd.n665 4.74817
R16487 gnd.n7132 gnd.n7131 4.74817
R16488 gnd.n5200 gnd.n5199 4.74817
R16489 gnd.n5194 gnd.n5192 4.74817
R16490 gnd.n5629 gnd.n1871 4.74817
R16491 gnd.n5627 gnd.n5626 4.74817
R16492 gnd.n5460 gnd.n5459 4.74817
R16493 gnd.n6832 gnd.n944 4.74817
R16494 gnd.n6828 gnd.n943 4.74817
R16495 gnd.n6824 gnd.n942 4.74817
R16496 gnd.n6841 gnd.n939 4.74817
R16497 gnd.n6839 gnd.n940 4.74817
R16498 gnd.n947 gnd.n944 4.74817
R16499 gnd.n6831 gnd.n943 4.74817
R16500 gnd.n6827 gnd.n942 4.74817
R16501 gnd.n6823 gnd.n939 4.74817
R16502 gnd.n6840 gnd.n6839 4.74817
R16503 gnd.n5647 gnd.n5646 4.74817
R16504 gnd.n5634 gnd.n1843 4.74817
R16505 gnd.n1865 gnd.n1842 4.74817
R16506 gnd.n5620 gnd.n1841 4.74817
R16507 gnd.n1881 gnd.n1840 4.74817
R16508 gnd.n5647 gnd.n1844 4.74817
R16509 gnd.n5645 gnd.n1843 4.74817
R16510 gnd.n5635 gnd.n1842 4.74817
R16511 gnd.n1864 gnd.n1841 4.74817
R16512 gnd.n5621 gnd.n1840 4.74817
R16513 gnd.n5199 gnd.n5198 4.74817
R16514 gnd.n5197 gnd.n5192 4.74817
R16515 gnd.n5193 gnd.n1871 4.74817
R16516 gnd.n5628 gnd.n5627 4.74817
R16517 gnd.n5459 gnd.n1872 4.74817
R16518 gnd.n4265 gnd.n4264 4.7074
R16519 gnd.n394 gnd.n393 4.7074
R16520 gnd.n6187 gnd.n1351 4.66575
R16521 gnd.n6383 gnd.n1248 4.66575
R16522 gnd.n6937 gnd.n879 4.6132
R16523 gnd.n5997 gnd.n5996 4.6132
R16524 gnd.n1128 gnd.n1115 4.46111
R16525 gnd.n4279 gnd.n4275 4.38594
R16526 gnd.n4316 gnd.n4312 4.38594
R16527 gnd.n4140 gnd.n4136 4.38594
R16528 gnd.n4177 gnd.n4173 4.38594
R16529 gnd.n4209 gnd.n4205 4.38594
R16530 gnd.n4246 gnd.n4242 4.38594
R16531 gnd.n445 gnd.n441 4.38594
R16532 gnd.n408 gnd.n404 4.38594
R16533 gnd.n306 gnd.n302 4.38594
R16534 gnd.n269 gnd.n265 4.38594
R16535 gnd.n375 gnd.n371 4.38594
R16536 gnd.n338 gnd.n334 4.38594
R16537 gnd.n4982 gnd.n4978 4.38594
R16538 gnd.n4950 gnd.n4946 4.38594
R16539 gnd.n4918 gnd.n4914 4.38594
R16540 gnd.n4887 gnd.n4883 4.38594
R16541 gnd.n4855 gnd.n4851 4.38594
R16542 gnd.n4823 gnd.n4819 4.38594
R16543 gnd.n4791 gnd.n4787 4.38594
R16544 gnd.n4760 gnd.n4756 4.38594
R16545 gnd.n109 gnd.n105 4.38594
R16546 gnd.n77 gnd.n73 4.38594
R16547 gnd.n45 gnd.n41 4.38594
R16548 gnd.n14 gnd.n10 4.38594
R16549 gnd.n236 gnd.n232 4.38594
R16550 gnd.n204 gnd.n200 4.38594
R16551 gnd.n172 gnd.n168 4.38594
R16552 gnd.n141 gnd.n137 4.38594
R16553 gnd.t220 gnd.n3839 4.33252
R16554 gnd.n5151 gnd.t20 4.33252
R16555 gnd.n4335 gnd.n4265 4.2808
R16556 gnd.n464 gnd.n394 4.2808
R16557 gnd.n4290 gnd.n4268 4.26717
R16558 gnd.n4327 gnd.n4305 4.26717
R16559 gnd.n4151 gnd.n4129 4.26717
R16560 gnd.n4188 gnd.n4166 4.26717
R16561 gnd.n4220 gnd.n4198 4.26717
R16562 gnd.n4257 gnd.n4235 4.26717
R16563 gnd.n456 gnd.n434 4.26717
R16564 gnd.n419 gnd.n397 4.26717
R16565 gnd.n317 gnd.n295 4.26717
R16566 gnd.n280 gnd.n258 4.26717
R16567 gnd.n386 gnd.n364 4.26717
R16568 gnd.n349 gnd.n327 4.26717
R16569 gnd.n4993 gnd.n4971 4.26717
R16570 gnd.n4961 gnd.n4939 4.26717
R16571 gnd.n4929 gnd.n4907 4.26717
R16572 gnd.n4898 gnd.n4876 4.26717
R16573 gnd.n4866 gnd.n4844 4.26717
R16574 gnd.n4834 gnd.n4812 4.26717
R16575 gnd.n4802 gnd.n4780 4.26717
R16576 gnd.n4771 gnd.n4749 4.26717
R16577 gnd.n120 gnd.n98 4.26717
R16578 gnd.n88 gnd.n66 4.26717
R16579 gnd.n56 gnd.n34 4.26717
R16580 gnd.n25 gnd.n3 4.26717
R16581 gnd.n247 gnd.n225 4.26717
R16582 gnd.n215 gnd.n193 4.26717
R16583 gnd.n183 gnd.n161 4.26717
R16584 gnd.n152 gnd.n130 4.26717
R16585 gnd.n255 gnd.n127 4.14478
R16586 gnd.n5001 gnd.n5000 4.08274
R16587 gnd.n1163 gnd.n1161 4.05904
R16588 gnd.n1549 gnd.n1492 4.05904
R16589 gnd.n6008 gnd.n6007 4.05904
R16590 gnd.n1156 gnd.n1151 4.05904
R16591 gnd.n6152 gnd.n1391 3.99929
R16592 gnd.n6459 gnd.n1217 3.99929
R16593 gnd.n6494 gnd.t114 3.99929
R16594 gnd.n5001 gnd.n4873 3.70378
R16595 gnd.n5558 gnd.t132 3.66606
R16596 gnd.n6131 gnd.t2 3.66606
R16597 gnd.n6493 gnd.t4 3.66606
R16598 gnd.n908 gnd.t110 3.66606
R16599 gnd.n255 gnd.n254 3.60163
R16600 gnd.n4337 gnd.n4336 3.58001
R16601 gnd.n4289 gnd.n4270 3.49141
R16602 gnd.n4326 gnd.n4307 3.49141
R16603 gnd.n4150 gnd.n4131 3.49141
R16604 gnd.n4187 gnd.n4168 3.49141
R16605 gnd.n4219 gnd.n4200 3.49141
R16606 gnd.n4256 gnd.n4237 3.49141
R16607 gnd.n455 gnd.n436 3.49141
R16608 gnd.n418 gnd.n399 3.49141
R16609 gnd.n316 gnd.n297 3.49141
R16610 gnd.n279 gnd.n260 3.49141
R16611 gnd.n385 gnd.n366 3.49141
R16612 gnd.n348 gnd.n329 3.49141
R16613 gnd.n4992 gnd.n4973 3.49141
R16614 gnd.n4960 gnd.n4941 3.49141
R16615 gnd.n4928 gnd.n4909 3.49141
R16616 gnd.n4897 gnd.n4878 3.49141
R16617 gnd.n4865 gnd.n4846 3.49141
R16618 gnd.n4833 gnd.n4814 3.49141
R16619 gnd.n4801 gnd.n4782 3.49141
R16620 gnd.n4770 gnd.n4751 3.49141
R16621 gnd.n119 gnd.n100 3.49141
R16622 gnd.n87 gnd.n68 3.49141
R16623 gnd.n55 gnd.n36 3.49141
R16624 gnd.n24 gnd.n5 3.49141
R16625 gnd.n246 gnd.n227 3.49141
R16626 gnd.n214 gnd.n195 3.49141
R16627 gnd.n182 gnd.n163 3.49141
R16628 gnd.n151 gnd.n132 3.49141
R16629 gnd.n6081 gnd.t191 3.33282
R16630 gnd.n6171 gnd.n6170 3.33282
R16631 gnd.n6195 gnd.t12 3.33282
R16632 gnd.n1245 gnd.t223 3.33282
R16633 gnd.n6447 gnd.n6446 3.33282
R16634 gnd.n4297 gnd.t93 3.3005
R16635 gnd.n4297 gnd.t64 3.3005
R16636 gnd.n4299 gnd.t46 3.3005
R16637 gnd.n4299 gnd.t90 3.3005
R16638 gnd.n4301 gnd.t67 3.3005
R16639 gnd.n4301 gnd.t86 3.3005
R16640 gnd.n4158 gnd.t84 3.3005
R16641 gnd.n4158 gnd.t70 3.3005
R16642 gnd.n4160 gnd.t104 3.3005
R16643 gnd.n4160 gnd.t71 3.3005
R16644 gnd.n4162 gnd.t57 3.3005
R16645 gnd.n4162 gnd.t101 3.3005
R16646 gnd.n4227 gnd.t78 3.3005
R16647 gnd.n4227 gnd.t59 3.3005
R16648 gnd.n4229 gnd.t92 3.3005
R16649 gnd.n4229 gnd.t61 3.3005
R16650 gnd.n4231 gnd.t108 3.3005
R16651 gnd.n4231 gnd.t89 3.3005
R16652 gnd.n430 gnd.t80 3.3005
R16653 gnd.n430 gnd.t63 3.3005
R16654 gnd.n428 gnd.t83 3.3005
R16655 gnd.n428 gnd.t106 3.3005
R16656 gnd.n426 gnd.t53 3.3005
R16657 gnd.n426 gnd.t94 3.3005
R16658 gnd.n291 gnd.t81 3.3005
R16659 gnd.n291 gnd.t102 3.3005
R16660 gnd.n289 gnd.t52 3.3005
R16661 gnd.n289 gnd.t82 3.3005
R16662 gnd.n287 gnd.t50 3.3005
R16663 gnd.n287 gnd.t48 3.3005
R16664 gnd.n360 gnd.t73 3.3005
R16665 gnd.n360 gnd.t91 3.3005
R16666 gnd.n358 gnd.t105 3.3005
R16667 gnd.n358 gnd.t75 3.3005
R16668 gnd.n356 gnd.t103 3.3005
R16669 gnd.n356 gnd.t98 3.3005
R16670 gnd.n4513 gnd.t220 2.99959
R16671 gnd.n4286 gnd.n4285 2.71565
R16672 gnd.n4323 gnd.n4322 2.71565
R16673 gnd.n4147 gnd.n4146 2.71565
R16674 gnd.n4184 gnd.n4183 2.71565
R16675 gnd.n4216 gnd.n4215 2.71565
R16676 gnd.n4253 gnd.n4252 2.71565
R16677 gnd.n452 gnd.n451 2.71565
R16678 gnd.n415 gnd.n414 2.71565
R16679 gnd.n313 gnd.n312 2.71565
R16680 gnd.n276 gnd.n275 2.71565
R16681 gnd.n382 gnd.n381 2.71565
R16682 gnd.n345 gnd.n344 2.71565
R16683 gnd.n4989 gnd.n4988 2.71565
R16684 gnd.n4957 gnd.n4956 2.71565
R16685 gnd.n4925 gnd.n4924 2.71565
R16686 gnd.n4894 gnd.n4893 2.71565
R16687 gnd.n4862 gnd.n4861 2.71565
R16688 gnd.n4830 gnd.n4829 2.71565
R16689 gnd.n4798 gnd.n4797 2.71565
R16690 gnd.n4767 gnd.n4766 2.71565
R16691 gnd.n116 gnd.n115 2.71565
R16692 gnd.n84 gnd.n83 2.71565
R16693 gnd.n52 gnd.n51 2.71565
R16694 gnd.n21 gnd.n20 2.71565
R16695 gnd.n243 gnd.n242 2.71565
R16696 gnd.n211 gnd.n210 2.71565
R16697 gnd.n179 gnd.n178 2.71565
R16698 gnd.n148 gnd.n147 2.71565
R16699 gnd.t215 gnd.n6151 2.66636
R16700 gnd.n6162 gnd.n6161 2.66636
R16701 gnd.n6161 gnd.t117 2.66636
R16702 gnd.n6213 gnd.t8 2.66636
R16703 gnd.t18 gnd.n1323 2.66636
R16704 gnd.n6269 gnd.n6268 2.66636
R16705 gnd.n6281 gnd.t217 2.66636
R16706 gnd.t224 gnd.n1293 2.66636
R16707 gnd.n6391 gnd.n6390 2.66636
R16708 gnd.n6389 gnd.t15 2.66636
R16709 gnd.n6410 gnd.t21 2.66636
R16710 gnd.n6467 gnd.n1206 2.66636
R16711 gnd.t146 gnd.n4451 2.33313
R16712 gnd.t19 gnd.n4564 2.33313
R16713 gnd.n6194 gnd.t6 2.33313
R16714 gnd.t6 gnd.n1359 2.33313
R16715 gnd.n6436 gnd.t25 2.33313
R16716 gnd.n1244 gnd.t25 2.33313
R16717 gnd.n4338 gnd.n4337 2.27742
R16718 gnd.n4337 gnd.n4126 2.27742
R16719 gnd.n4337 gnd.n4119 2.27742
R16720 gnd.n4337 gnd.n4092 2.27742
R16721 gnd.n7100 gnd.n649 2.27742
R16722 gnd.n680 gnd.n649 2.27742
R16723 gnd.n7116 gnd.n649 2.27742
R16724 gnd.n665 gnd.n649 2.27742
R16725 gnd.n7132 gnd.n649 2.27742
R16726 gnd.n6838 gnd.n944 2.27742
R16727 gnd.n6838 gnd.n943 2.27742
R16728 gnd.n6838 gnd.n942 2.27742
R16729 gnd.n6838 gnd.n939 2.27742
R16730 gnd.n6839 gnd.n6838 2.27742
R16731 gnd.n5648 gnd.n5647 2.27742
R16732 gnd.n5648 gnd.n1843 2.27742
R16733 gnd.n5648 gnd.n1842 2.27742
R16734 gnd.n5648 gnd.n1841 2.27742
R16735 gnd.n5648 gnd.n1840 2.27742
R16736 gnd.n5199 gnd.n1839 2.27742
R16737 gnd.n5192 gnd.n1839 2.27742
R16738 gnd.n1871 gnd.n1839 2.27742
R16739 gnd.n5627 gnd.n1839 2.27742
R16740 gnd.n5459 gnd.n1839 2.27742
R16741 gnd.n5159 gnd.t222 1.99989
R16742 gnd.t179 gnd.n6071 1.99989
R16743 gnd.n6133 gnd.t191 1.99989
R16744 gnd.n6125 gnd.t120 1.99989
R16745 gnd.n6151 gnd.n1393 1.99989
R16746 gnd.n6282 gnd.n1314 1.99989
R16747 gnd.n6325 gnd.n1292 1.99989
R16748 gnd.n6474 gnd.t208 1.99989
R16749 gnd.n6473 gnd.n1202 1.99989
R16750 gnd.n6487 gnd.t156 1.99989
R16751 gnd.n4282 gnd.n4272 1.93989
R16752 gnd.n4319 gnd.n4309 1.93989
R16753 gnd.n4143 gnd.n4133 1.93989
R16754 gnd.n4180 gnd.n4170 1.93989
R16755 gnd.n4212 gnd.n4202 1.93989
R16756 gnd.n4249 gnd.n4239 1.93989
R16757 gnd.n448 gnd.n438 1.93989
R16758 gnd.n411 gnd.n401 1.93989
R16759 gnd.n309 gnd.n299 1.93989
R16760 gnd.n272 gnd.n262 1.93989
R16761 gnd.n378 gnd.n368 1.93989
R16762 gnd.n341 gnd.n331 1.93989
R16763 gnd.n4985 gnd.n4975 1.93989
R16764 gnd.n4953 gnd.n4943 1.93989
R16765 gnd.n4921 gnd.n4911 1.93989
R16766 gnd.n4890 gnd.n4880 1.93989
R16767 gnd.n4858 gnd.n4848 1.93989
R16768 gnd.n4826 gnd.n4816 1.93989
R16769 gnd.n4794 gnd.n4784 1.93989
R16770 gnd.n4763 gnd.n4753 1.93989
R16771 gnd.n112 gnd.n102 1.93989
R16772 gnd.n80 gnd.n70 1.93989
R16773 gnd.n48 gnd.n38 1.93989
R16774 gnd.n17 gnd.n7 1.93989
R16775 gnd.n239 gnd.n229 1.93989
R16776 gnd.n207 gnd.n197 1.93989
R16777 gnd.n175 gnd.n165 1.93989
R16778 gnd.n144 gnd.n134 1.93989
R16779 gnd.n4360 gnd.t41 1.66666
R16780 gnd.n4106 gnd.t23 1.66666
R16781 gnd.n4694 gnd.t35 1.66666
R16782 gnd.n6059 gnd.n1423 1.66666
R16783 gnd.t2 gnd.n1399 1.66666
R16784 gnd.n6355 gnd.t4 1.66666
R16785 gnd.n6621 gnd.n1102 1.66666
R16786 gnd.n4302 gnd.n4300 1.35515
R16787 gnd.n431 gnd.n429 1.35515
R16788 gnd.n4334 gnd.n4302 1.35515
R16789 gnd.n4300 gnd.n4298 1.35515
R16790 gnd.n429 gnd.n427 1.35515
R16791 gnd.n463 gnd.n431 1.35515
R16792 gnd.n5305 gnd.n1990 1.33343
R16793 gnd.n5227 gnd.n1978 1.33343
R16794 gnd.n5313 gnd.n1981 1.33343
R16795 gnd.n5221 gnd.n5220 1.33343
R16796 gnd.n5321 gnd.n1972 1.33343
R16797 gnd.n2212 gnd.n1960 1.33343
R16798 gnd.n5338 gnd.n1963 1.33343
R16799 gnd.n2206 gnd.n1950 1.33343
R16800 gnd.n5348 gnd.n1952 1.33343
R16801 gnd.n5331 gnd.n1944 1.33343
R16802 gnd.n5362 gnd.n1921 1.33343
R16803 gnd.n5379 gnd.n1924 1.33343
R16804 gnd.n5356 gnd.n1938 1.33343
R16805 gnd.n5388 gnd.n1912 1.33343
R16806 gnd.n1934 gnd.n1904 1.33343
R16807 gnd.n5397 gnd.n1847 1.33343
R16808 gnd.n5643 gnd.n1850 1.33343
R16809 gnd.n5405 gnd.n1859 1.33343
R16810 gnd.n5637 gnd.n1862 1.33343
R16811 gnd.n5632 gnd.n5631 1.33343
R16812 gnd.n1874 gnd.n1868 1.33343
R16813 gnd.n5624 gnd.n1875 1.33343
R16814 gnd.n5623 gnd.n1878 1.33343
R16815 gnd.n5618 gnd.n1884 1.33343
R16816 gnd.n5596 gnd.n1832 1.33343
R16817 gnd.n5652 gnd.n1835 1.33343
R16818 gnd.n5480 gnd.n1823 1.33343
R16819 gnd.n5660 gnd.n1826 1.33343
R16820 gnd.n5484 gnd.n1814 1.33343
R16821 gnd.n5668 gnd.n1817 1.33343
R16822 gnd.n5512 gnd.n5511 1.33343
R16823 gnd.n5676 gnd.n1808 1.33343
R16824 gnd.n5505 gnd.n1797 1.33343
R16825 gnd.n5684 gnd.n1800 1.33343
R16826 gnd.n5501 gnd.n1788 1.33343
R16827 gnd.n5692 gnd.n1791 1.33343
R16828 gnd.n5497 gnd.n1779 1.33343
R16829 gnd.n5700 gnd.n1782 1.33343
R16830 gnd.n5569 gnd.n1769 1.33343
R16831 gnd.n5713 gnd.n1772 1.33343
R16832 gnd.n5563 gnd.n1760 1.33343
R16833 gnd.n5721 gnd.n1762 1.33343
R16834 gnd.n5559 gnd.n5558 1.33343
R16835 gnd.n5904 gnd.n1613 1.33343
R16836 gnd.n5728 gnd.n1601 1.33343
R16837 gnd.n5958 gnd.n1603 1.33343
R16838 gnd.n6196 gnd.n6195 1.33343
R16839 gnd.n6220 gnd.n1342 1.33343
R16840 gnd.n6261 gnd.t217 1.33343
R16841 gnd.n1294 gnd.t224 1.33343
R16842 gnd.n6382 gnd.n1273 1.33343
R16843 gnd.n6419 gnd.n1245 1.33343
R16844 gnd.t176 gnd.n1111 1.33343
R16845 gnd.n7015 gnd.n786 1.33343
R16846 gnd.n1013 gnd.n789 1.33343
R16847 gnd.n7023 gnd.n779 1.33343
R16848 gnd.n6892 gnd.n908 1.33343
R16849 gnd.n7031 gnd.n770 1.33343
R16850 gnd.n6758 gnd.n773 1.33343
R16851 gnd.n7039 gnd.n761 1.33343
R16852 gnd.n6764 gnd.n764 1.33343
R16853 gnd.n7047 gnd.n752 1.33343
R16854 gnd.n6768 gnd.n755 1.33343
R16855 gnd.n7055 gnd.n743 1.33343
R16856 gnd.n6774 gnd.n746 1.33343
R16857 gnd.n7063 gnd.n734 1.33343
R16858 gnd.n6778 gnd.n737 1.33343
R16859 gnd.n7071 gnd.n726 1.33343
R16860 gnd.n6812 gnd.n6811 1.33343
R16861 gnd.n7079 gnd.n717 1.33343
R16862 gnd.n6805 gnd.n720 1.33343
R16863 gnd.n7088 gnd.n708 1.33343
R16864 gnd.n6801 gnd.n711 1.33343
R16865 gnd.n7096 gnd.n699 1.33343
R16866 gnd.n6797 gnd.n702 1.33343
R16867 gnd.n7104 gnd.n691 1.33343
R16868 gnd.n6793 gnd.n694 1.33343
R16869 gnd.n7112 gnd.n682 1.33343
R16870 gnd.n6854 gnd.n685 1.33343
R16871 gnd.n7120 gnd.n675 1.33343
R16872 gnd.n6848 gnd.n678 1.33343
R16873 gnd.n7128 gnd.n667 1.33343
R16874 gnd.n6844 gnd.n6843 1.33343
R16875 gnd.n7135 gnd.n660 1.33343
R16876 gnd.n2840 gnd.n663 1.33343
R16877 gnd.n7143 gnd.n652 1.33343
R16878 gnd.n7151 gnd.n643 1.33343
R16879 gnd.n2850 gnd.n646 1.33343
R16880 gnd.n7159 gnd.n635 1.33343
R16881 gnd.n2854 gnd.n637 1.33343
R16882 gnd.n7167 gnd.n626 1.33343
R16883 gnd.n2860 gnd.n629 1.33343
R16884 gnd.n7175 gnd.n618 1.33343
R16885 gnd.n2864 gnd.n620 1.33343
R16886 gnd.n7183 gnd.n610 1.33343
R16887 gnd.n2889 gnd.n2888 1.33343
R16888 gnd.n7191 gnd.n602 1.33343
R16889 gnd.n2882 gnd.n604 1.33343
R16890 gnd.n7199 gnd.n593 1.33343
R16891 gnd.n4281 gnd.n4274 1.16414
R16892 gnd.n4318 gnd.n4311 1.16414
R16893 gnd.n4142 gnd.n4135 1.16414
R16894 gnd.n4179 gnd.n4172 1.16414
R16895 gnd.n4211 gnd.n4204 1.16414
R16896 gnd.n4248 gnd.n4241 1.16414
R16897 gnd.n447 gnd.n440 1.16414
R16898 gnd.n410 gnd.n403 1.16414
R16899 gnd.n308 gnd.n301 1.16414
R16900 gnd.n271 gnd.n264 1.16414
R16901 gnd.n377 gnd.n370 1.16414
R16902 gnd.n340 gnd.n333 1.16414
R16903 gnd.n5743 gnd.n5739 1.16414
R16904 gnd.n3985 gnd.n3984 1.16414
R16905 gnd.n5041 gnd.n3676 1.16414
R16906 gnd.n4984 gnd.n4977 1.16414
R16907 gnd.n4952 gnd.n4945 1.16414
R16908 gnd.n4920 gnd.n4913 1.16414
R16909 gnd.n4889 gnd.n4882 1.16414
R16910 gnd.n4857 gnd.n4850 1.16414
R16911 gnd.n4825 gnd.n4818 1.16414
R16912 gnd.n4793 gnd.n4786 1.16414
R16913 gnd.n4762 gnd.n4755 1.16414
R16914 gnd.n1030 gnd.n1029 1.16414
R16915 gnd.n111 gnd.n104 1.16414
R16916 gnd.n79 gnd.n72 1.16414
R16917 gnd.n47 gnd.n40 1.16414
R16918 gnd.n16 gnd.n9 1.16414
R16919 gnd.n238 gnd.n231 1.16414
R16920 gnd.n206 gnd.n199 1.16414
R16921 gnd.n174 gnd.n167 1.16414
R16922 gnd.n143 gnd.n136 1.16414
R16923 gnd.n4195 gnd.n4163 1.00481
R16924 gnd.n4163 gnd.n4161 1.00481
R16925 gnd.n4161 gnd.n4159 1.00481
R16926 gnd.n4264 gnd.n4232 1.00481
R16927 gnd.n4232 gnd.n4230 1.00481
R16928 gnd.n4230 gnd.n4228 1.00481
R16929 gnd.n290 gnd.n288 1.00481
R16930 gnd.n292 gnd.n290 1.00481
R16931 gnd.n324 gnd.n292 1.00481
R16932 gnd.n359 gnd.n357 1.00481
R16933 gnd.n361 gnd.n359 1.00481
R16934 gnd.n393 gnd.n361 1.00481
R16935 gnd.t43 gnd.n3813 1.0002
R16936 gnd.n4678 gnd.t16 1.0002
R16937 gnd.t85 gnd.n1910 1.0002
R16938 gnd.t72 gnd.n654 1.0002
R16939 gnd.n6937 gnd.n6936 0.970197
R16940 gnd.n5997 gnd.n1557 0.970197
R16941 gnd.n4968 gnd.n4936 0.962709
R16942 gnd.n5000 gnd.n4968 0.962709
R16943 gnd.n4841 gnd.n4809 0.962709
R16944 gnd.n4873 gnd.n4841 0.962709
R16945 gnd.n95 gnd.n63 0.962709
R16946 gnd.n127 gnd.n95 0.962709
R16947 gnd.n222 gnd.n190 0.962709
R16948 gnd.n254 gnd.n222 0.962709
R16949 gnd.n1496 gnd.n1415 0.666965
R16950 gnd.n6143 gnd.n6142 0.666965
R16951 gnd.n6227 gnd.t18 0.666965
R16952 gnd.n6304 gnd.n6303 0.666965
R16953 gnd.n6297 gnd.n1285 0.666965
R16954 gnd.t15 gnd.n1255 0.666965
R16955 gnd.t139 gnd.t156 0.666965
R16956 gnd.n6354 gnd.n1191 0.666965
R16957 gnd.n6611 gnd.n6610 0.666965
R16958 gnd.n7396 gnd.n7395 0.57484
R16959 gnd.n6838 gnd.n649 0.549125
R16960 gnd.n5648 gnd.n1839 0.549125
R16961 gnd.n5897 gnd.n5896 0.526415
R16962 gnd.n6699 gnd.n791 0.526415
R16963 gnd gnd.n0 0.52173
R16964 gnd.n5029 gnd.n3680 0.486781
R16965 gnd.n4037 gnd.n3933 0.48678
R16966 gnd.n6708 gnd.n6707 0.48678
R16967 gnd.n5822 gnd.n1666 0.48678
R16968 gnd.n5241 gnd.n5240 0.483732
R16969 gnd.n5278 gnd.n5277 0.483732
R16970 gnd.n7266 gnd.n7265 0.483732
R16971 gnd.n7241 gnd.n497 0.483732
R16972 gnd.n3631 gnd.n3602 0.480683
R16973 gnd.n4380 gnd.n3884 0.480683
R16974 gnd.n7350 gnd.n7349 0.471537
R16975 gnd.n7289 gnd.n7288 0.471537
R16976 gnd.n6901 gnd.n6898 0.471537
R16977 gnd.n7018 gnd.n784 0.471537
R16978 gnd.n5955 gnd.n5954 0.471537
R16979 gnd.n5962 gnd.n5961 0.471537
R16980 gnd.n2175 gnd.n2174 0.471537
R16981 gnd.n5284 gnd.n2010 0.471537
R16982 gnd.n3378 gnd.n2321 0.438
R16983 gnd.n3033 gnd.n3032 0.438
R16984 gnd.n2896 gnd.n2895 0.438
R16985 gnd.n5166 gnd.n2221 0.438
R16986 gnd.n4278 gnd.n4277 0.388379
R16987 gnd.n4315 gnd.n4314 0.388379
R16988 gnd.n4139 gnd.n4138 0.388379
R16989 gnd.n4176 gnd.n4175 0.388379
R16990 gnd.n4208 gnd.n4207 0.388379
R16991 gnd.n4245 gnd.n4244 0.388379
R16992 gnd.n444 gnd.n443 0.388379
R16993 gnd.n407 gnd.n406 0.388379
R16994 gnd.n305 gnd.n304 0.388379
R16995 gnd.n268 gnd.n267 0.388379
R16996 gnd.n374 gnd.n373 0.388379
R16997 gnd.n337 gnd.n336 0.388379
R16998 gnd.n4981 gnd.n4980 0.388379
R16999 gnd.n4949 gnd.n4948 0.388379
R17000 gnd.n4917 gnd.n4916 0.388379
R17001 gnd.n4886 gnd.n4885 0.388379
R17002 gnd.n4854 gnd.n4853 0.388379
R17003 gnd.n4822 gnd.n4821 0.388379
R17004 gnd.n4790 gnd.n4789 0.388379
R17005 gnd.n4759 gnd.n4758 0.388379
R17006 gnd.n537 gnd.n532 0.388379
R17007 gnd.n2125 gnd.n2124 0.388379
R17008 gnd.n108 gnd.n107 0.388379
R17009 gnd.n76 gnd.n75 0.388379
R17010 gnd.n44 gnd.n43 0.388379
R17011 gnd.n13 gnd.n12 0.388379
R17012 gnd.n235 gnd.n234 0.388379
R17013 gnd.n203 gnd.n202 0.388379
R17014 gnd.n171 gnd.n170 0.388379
R17015 gnd.n140 gnd.n139 0.388379
R17016 gnd.n5899 gnd.n5898 0.383651
R17017 gnd.n7012 gnd.n7011 0.383651
R17018 gnd.n7396 gnd.n255 0.341877
R17019 gnd.n5144 gnd.t227 0.333732
R17020 gnd.n5373 gnd.t85 0.333732
R17021 gnd.n5480 gnd.t77 0.333732
R17022 gnd.n5830 gnd.t204 0.333732
R17023 gnd.n6693 gnd.t211 0.333732
R17024 gnd.n6801 gnd.t47 0.333732
R17025 gnd.n2844 gnd.t72 0.333732
R17026 gnd.n4031 gnd.n4030 0.311721
R17027 gnd.n5086 gnd.n5085 0.268793
R17028 gnd.n5733 gnd.n5732 0.253549
R17029 gnd.n1018 gnd.n1017 0.253549
R17030 gnd.n5085 gnd.n5084 0.241354
R17031 gnd.n879 gnd.n876 0.229039
R17032 gnd.n882 gnd.n879 0.229039
R17033 gnd.n5996 gnd.n1562 0.229039
R17034 gnd.n5996 gnd.n5995 0.229039
R17035 gnd gnd.n7396 0.213018
R17036 gnd.n4435 gnd.n3901 0.206293
R17037 gnd.n4295 gnd.n4267 0.155672
R17038 gnd.n4288 gnd.n4267 0.155672
R17039 gnd.n4288 gnd.n4287 0.155672
R17040 gnd.n4287 gnd.n4271 0.155672
R17041 gnd.n4280 gnd.n4271 0.155672
R17042 gnd.n4280 gnd.n4279 0.155672
R17043 gnd.n4332 gnd.n4304 0.155672
R17044 gnd.n4325 gnd.n4304 0.155672
R17045 gnd.n4325 gnd.n4324 0.155672
R17046 gnd.n4324 gnd.n4308 0.155672
R17047 gnd.n4317 gnd.n4308 0.155672
R17048 gnd.n4317 gnd.n4316 0.155672
R17049 gnd.n4156 gnd.n4128 0.155672
R17050 gnd.n4149 gnd.n4128 0.155672
R17051 gnd.n4149 gnd.n4148 0.155672
R17052 gnd.n4148 gnd.n4132 0.155672
R17053 gnd.n4141 gnd.n4132 0.155672
R17054 gnd.n4141 gnd.n4140 0.155672
R17055 gnd.n4193 gnd.n4165 0.155672
R17056 gnd.n4186 gnd.n4165 0.155672
R17057 gnd.n4186 gnd.n4185 0.155672
R17058 gnd.n4185 gnd.n4169 0.155672
R17059 gnd.n4178 gnd.n4169 0.155672
R17060 gnd.n4178 gnd.n4177 0.155672
R17061 gnd.n4225 gnd.n4197 0.155672
R17062 gnd.n4218 gnd.n4197 0.155672
R17063 gnd.n4218 gnd.n4217 0.155672
R17064 gnd.n4217 gnd.n4201 0.155672
R17065 gnd.n4210 gnd.n4201 0.155672
R17066 gnd.n4210 gnd.n4209 0.155672
R17067 gnd.n4262 gnd.n4234 0.155672
R17068 gnd.n4255 gnd.n4234 0.155672
R17069 gnd.n4255 gnd.n4254 0.155672
R17070 gnd.n4254 gnd.n4238 0.155672
R17071 gnd.n4247 gnd.n4238 0.155672
R17072 gnd.n4247 gnd.n4246 0.155672
R17073 gnd.n461 gnd.n433 0.155672
R17074 gnd.n454 gnd.n433 0.155672
R17075 gnd.n454 gnd.n453 0.155672
R17076 gnd.n453 gnd.n437 0.155672
R17077 gnd.n446 gnd.n437 0.155672
R17078 gnd.n446 gnd.n445 0.155672
R17079 gnd.n424 gnd.n396 0.155672
R17080 gnd.n417 gnd.n396 0.155672
R17081 gnd.n417 gnd.n416 0.155672
R17082 gnd.n416 gnd.n400 0.155672
R17083 gnd.n409 gnd.n400 0.155672
R17084 gnd.n409 gnd.n408 0.155672
R17085 gnd.n322 gnd.n294 0.155672
R17086 gnd.n315 gnd.n294 0.155672
R17087 gnd.n315 gnd.n314 0.155672
R17088 gnd.n314 gnd.n298 0.155672
R17089 gnd.n307 gnd.n298 0.155672
R17090 gnd.n307 gnd.n306 0.155672
R17091 gnd.n285 gnd.n257 0.155672
R17092 gnd.n278 gnd.n257 0.155672
R17093 gnd.n278 gnd.n277 0.155672
R17094 gnd.n277 gnd.n261 0.155672
R17095 gnd.n270 gnd.n261 0.155672
R17096 gnd.n270 gnd.n269 0.155672
R17097 gnd.n391 gnd.n363 0.155672
R17098 gnd.n384 gnd.n363 0.155672
R17099 gnd.n384 gnd.n383 0.155672
R17100 gnd.n383 gnd.n367 0.155672
R17101 gnd.n376 gnd.n367 0.155672
R17102 gnd.n376 gnd.n375 0.155672
R17103 gnd.n354 gnd.n326 0.155672
R17104 gnd.n347 gnd.n326 0.155672
R17105 gnd.n347 gnd.n346 0.155672
R17106 gnd.n346 gnd.n330 0.155672
R17107 gnd.n339 gnd.n330 0.155672
R17108 gnd.n339 gnd.n338 0.155672
R17109 gnd.n4998 gnd.n4970 0.155672
R17110 gnd.n4991 gnd.n4970 0.155672
R17111 gnd.n4991 gnd.n4990 0.155672
R17112 gnd.n4990 gnd.n4974 0.155672
R17113 gnd.n4983 gnd.n4974 0.155672
R17114 gnd.n4983 gnd.n4982 0.155672
R17115 gnd.n4966 gnd.n4938 0.155672
R17116 gnd.n4959 gnd.n4938 0.155672
R17117 gnd.n4959 gnd.n4958 0.155672
R17118 gnd.n4958 gnd.n4942 0.155672
R17119 gnd.n4951 gnd.n4942 0.155672
R17120 gnd.n4951 gnd.n4950 0.155672
R17121 gnd.n4934 gnd.n4906 0.155672
R17122 gnd.n4927 gnd.n4906 0.155672
R17123 gnd.n4927 gnd.n4926 0.155672
R17124 gnd.n4926 gnd.n4910 0.155672
R17125 gnd.n4919 gnd.n4910 0.155672
R17126 gnd.n4919 gnd.n4918 0.155672
R17127 gnd.n4903 gnd.n4875 0.155672
R17128 gnd.n4896 gnd.n4875 0.155672
R17129 gnd.n4896 gnd.n4895 0.155672
R17130 gnd.n4895 gnd.n4879 0.155672
R17131 gnd.n4888 gnd.n4879 0.155672
R17132 gnd.n4888 gnd.n4887 0.155672
R17133 gnd.n4871 gnd.n4843 0.155672
R17134 gnd.n4864 gnd.n4843 0.155672
R17135 gnd.n4864 gnd.n4863 0.155672
R17136 gnd.n4863 gnd.n4847 0.155672
R17137 gnd.n4856 gnd.n4847 0.155672
R17138 gnd.n4856 gnd.n4855 0.155672
R17139 gnd.n4839 gnd.n4811 0.155672
R17140 gnd.n4832 gnd.n4811 0.155672
R17141 gnd.n4832 gnd.n4831 0.155672
R17142 gnd.n4831 gnd.n4815 0.155672
R17143 gnd.n4824 gnd.n4815 0.155672
R17144 gnd.n4824 gnd.n4823 0.155672
R17145 gnd.n4807 gnd.n4779 0.155672
R17146 gnd.n4800 gnd.n4779 0.155672
R17147 gnd.n4800 gnd.n4799 0.155672
R17148 gnd.n4799 gnd.n4783 0.155672
R17149 gnd.n4792 gnd.n4783 0.155672
R17150 gnd.n4792 gnd.n4791 0.155672
R17151 gnd.n4776 gnd.n4748 0.155672
R17152 gnd.n4769 gnd.n4748 0.155672
R17153 gnd.n4769 gnd.n4768 0.155672
R17154 gnd.n4768 gnd.n4752 0.155672
R17155 gnd.n4761 gnd.n4752 0.155672
R17156 gnd.n4761 gnd.n4760 0.155672
R17157 gnd.n125 gnd.n97 0.155672
R17158 gnd.n118 gnd.n97 0.155672
R17159 gnd.n118 gnd.n117 0.155672
R17160 gnd.n117 gnd.n101 0.155672
R17161 gnd.n110 gnd.n101 0.155672
R17162 gnd.n110 gnd.n109 0.155672
R17163 gnd.n93 gnd.n65 0.155672
R17164 gnd.n86 gnd.n65 0.155672
R17165 gnd.n86 gnd.n85 0.155672
R17166 gnd.n85 gnd.n69 0.155672
R17167 gnd.n78 gnd.n69 0.155672
R17168 gnd.n78 gnd.n77 0.155672
R17169 gnd.n61 gnd.n33 0.155672
R17170 gnd.n54 gnd.n33 0.155672
R17171 gnd.n54 gnd.n53 0.155672
R17172 gnd.n53 gnd.n37 0.155672
R17173 gnd.n46 gnd.n37 0.155672
R17174 gnd.n46 gnd.n45 0.155672
R17175 gnd.n30 gnd.n2 0.155672
R17176 gnd.n23 gnd.n2 0.155672
R17177 gnd.n23 gnd.n22 0.155672
R17178 gnd.n22 gnd.n6 0.155672
R17179 gnd.n15 gnd.n6 0.155672
R17180 gnd.n15 gnd.n14 0.155672
R17181 gnd.n252 gnd.n224 0.155672
R17182 gnd.n245 gnd.n224 0.155672
R17183 gnd.n245 gnd.n244 0.155672
R17184 gnd.n244 gnd.n228 0.155672
R17185 gnd.n237 gnd.n228 0.155672
R17186 gnd.n237 gnd.n236 0.155672
R17187 gnd.n220 gnd.n192 0.155672
R17188 gnd.n213 gnd.n192 0.155672
R17189 gnd.n213 gnd.n212 0.155672
R17190 gnd.n212 gnd.n196 0.155672
R17191 gnd.n205 gnd.n196 0.155672
R17192 gnd.n205 gnd.n204 0.155672
R17193 gnd.n188 gnd.n160 0.155672
R17194 gnd.n181 gnd.n160 0.155672
R17195 gnd.n181 gnd.n180 0.155672
R17196 gnd.n180 gnd.n164 0.155672
R17197 gnd.n173 gnd.n164 0.155672
R17198 gnd.n173 gnd.n172 0.155672
R17199 gnd.n157 gnd.n129 0.155672
R17200 gnd.n150 gnd.n129 0.155672
R17201 gnd.n150 gnd.n149 0.155672
R17202 gnd.n149 gnd.n133 0.155672
R17203 gnd.n142 gnd.n133 0.155672
R17204 gnd.n142 gnd.n141 0.155672
R17205 gnd.n3632 gnd.n3631 0.152939
R17206 gnd.n3633 gnd.n3632 0.152939
R17207 gnd.n3634 gnd.n3633 0.152939
R17208 gnd.n3635 gnd.n3634 0.152939
R17209 gnd.n3636 gnd.n3635 0.152939
R17210 gnd.n3637 gnd.n3636 0.152939
R17211 gnd.n3638 gnd.n3637 0.152939
R17212 gnd.n3639 gnd.n3638 0.152939
R17213 gnd.n3640 gnd.n3639 0.152939
R17214 gnd.n3641 gnd.n3640 0.152939
R17215 gnd.n3642 gnd.n3641 0.152939
R17216 gnd.n3643 gnd.n3642 0.152939
R17217 gnd.n3644 gnd.n3643 0.152939
R17218 gnd.n3645 gnd.n3644 0.152939
R17219 gnd.n5087 gnd.n3645 0.152939
R17220 gnd.n5087 gnd.n5086 0.152939
R17221 gnd.n4455 gnd.n3884 0.152939
R17222 gnd.n4456 gnd.n4455 0.152939
R17223 gnd.n4457 gnd.n4456 0.152939
R17224 gnd.n4458 gnd.n4457 0.152939
R17225 gnd.n4458 gnd.n3859 0.152939
R17226 gnd.n4486 gnd.n3859 0.152939
R17227 gnd.n4487 gnd.n4486 0.152939
R17228 gnd.n4488 gnd.n4487 0.152939
R17229 gnd.n4489 gnd.n4488 0.152939
R17230 gnd.n4489 gnd.n3833 0.152939
R17231 gnd.n4517 gnd.n3833 0.152939
R17232 gnd.n4518 gnd.n4517 0.152939
R17233 gnd.n4519 gnd.n4518 0.152939
R17234 gnd.n4520 gnd.n4519 0.152939
R17235 gnd.n4520 gnd.n3807 0.152939
R17236 gnd.n4548 gnd.n3807 0.152939
R17237 gnd.n4549 gnd.n4548 0.152939
R17238 gnd.n4550 gnd.n4549 0.152939
R17239 gnd.n4551 gnd.n4550 0.152939
R17240 gnd.n4551 gnd.n3781 0.152939
R17241 gnd.n4579 gnd.n3781 0.152939
R17242 gnd.n4580 gnd.n4579 0.152939
R17243 gnd.n4581 gnd.n4580 0.152939
R17244 gnd.n4582 gnd.n4581 0.152939
R17245 gnd.n4582 gnd.n3756 0.152939
R17246 gnd.n4610 gnd.n3756 0.152939
R17247 gnd.n4611 gnd.n4610 0.152939
R17248 gnd.n4612 gnd.n4611 0.152939
R17249 gnd.n4613 gnd.n4612 0.152939
R17250 gnd.n4613 gnd.n3729 0.152939
R17251 gnd.n4640 gnd.n3729 0.152939
R17252 gnd.n4641 gnd.n4640 0.152939
R17253 gnd.n4642 gnd.n4641 0.152939
R17254 gnd.n4642 gnd.n3707 0.152939
R17255 gnd.n4682 gnd.n3707 0.152939
R17256 gnd.n4683 gnd.n4682 0.152939
R17257 gnd.n4684 gnd.n4683 0.152939
R17258 gnd.n4685 gnd.n4684 0.152939
R17259 gnd.n4687 gnd.n4685 0.152939
R17260 gnd.n4687 gnd.n4686 0.152939
R17261 gnd.n4686 gnd.n3552 0.152939
R17262 gnd.n3553 gnd.n3552 0.152939
R17263 gnd.n3554 gnd.n3553 0.152939
R17264 gnd.n3574 gnd.n3554 0.152939
R17265 gnd.n3575 gnd.n3574 0.152939
R17266 gnd.n3576 gnd.n3575 0.152939
R17267 gnd.n3577 gnd.n3576 0.152939
R17268 gnd.n3578 gnd.n3577 0.152939
R17269 gnd.n3598 gnd.n3578 0.152939
R17270 gnd.n3599 gnd.n3598 0.152939
R17271 gnd.n3600 gnd.n3599 0.152939
R17272 gnd.n3601 gnd.n3600 0.152939
R17273 gnd.n3602 gnd.n3601 0.152939
R17274 gnd.n4381 gnd.n4380 0.152939
R17275 gnd.n4382 gnd.n4381 0.152939
R17276 gnd.n4383 gnd.n4382 0.152939
R17277 gnd.n4384 gnd.n4383 0.152939
R17278 gnd.n4385 gnd.n4384 0.152939
R17279 gnd.n4386 gnd.n4385 0.152939
R17280 gnd.n4387 gnd.n4386 0.152939
R17281 gnd.n4388 gnd.n4387 0.152939
R17282 gnd.n4389 gnd.n4388 0.152939
R17283 gnd.n4390 gnd.n4389 0.152939
R17284 gnd.n4391 gnd.n4390 0.152939
R17285 gnd.n4392 gnd.n4391 0.152939
R17286 gnd.n4393 gnd.n4392 0.152939
R17287 gnd.n4394 gnd.n4393 0.152939
R17288 gnd.n4398 gnd.n4394 0.152939
R17289 gnd.n4398 gnd.n3901 0.152939
R17290 gnd.n5084 gnd.n3651 0.152939
R17291 gnd.n3653 gnd.n3651 0.152939
R17292 gnd.n3654 gnd.n3653 0.152939
R17293 gnd.n3655 gnd.n3654 0.152939
R17294 gnd.n3656 gnd.n3655 0.152939
R17295 gnd.n3657 gnd.n3656 0.152939
R17296 gnd.n3658 gnd.n3657 0.152939
R17297 gnd.n3659 gnd.n3658 0.152939
R17298 gnd.n3660 gnd.n3659 0.152939
R17299 gnd.n3661 gnd.n3660 0.152939
R17300 gnd.n3662 gnd.n3661 0.152939
R17301 gnd.n3663 gnd.n3662 0.152939
R17302 gnd.n3664 gnd.n3663 0.152939
R17303 gnd.n3665 gnd.n3664 0.152939
R17304 gnd.n3666 gnd.n3665 0.152939
R17305 gnd.n3667 gnd.n3666 0.152939
R17306 gnd.n3668 gnd.n3667 0.152939
R17307 gnd.n3669 gnd.n3668 0.152939
R17308 gnd.n3670 gnd.n3669 0.152939
R17309 gnd.n3671 gnd.n3670 0.152939
R17310 gnd.n3672 gnd.n3671 0.152939
R17311 gnd.n3673 gnd.n3672 0.152939
R17312 gnd.n3677 gnd.n3673 0.152939
R17313 gnd.n3678 gnd.n3677 0.152939
R17314 gnd.n3679 gnd.n3678 0.152939
R17315 gnd.n3680 gnd.n3679 0.152939
R17316 gnd.n4093 gnd.n4091 0.152939
R17317 gnd.n4094 gnd.n4093 0.152939
R17318 gnd.n4095 gnd.n4094 0.152939
R17319 gnd.n4096 gnd.n4095 0.152939
R17320 gnd.n4097 gnd.n4096 0.152939
R17321 gnd.n4098 gnd.n4097 0.152939
R17322 gnd.n4099 gnd.n4098 0.152939
R17323 gnd.n4099 gnd.n3714 0.152939
R17324 gnd.n4660 gnd.n3714 0.152939
R17325 gnd.n4661 gnd.n4660 0.152939
R17326 gnd.n4662 gnd.n4661 0.152939
R17327 gnd.n4663 gnd.n4662 0.152939
R17328 gnd.n4664 gnd.n4663 0.152939
R17329 gnd.n4665 gnd.n4664 0.152939
R17330 gnd.n4666 gnd.n4665 0.152939
R17331 gnd.n4667 gnd.n4666 0.152939
R17332 gnd.n4667 gnd.n3691 0.152939
R17333 gnd.n4720 gnd.n3691 0.152939
R17334 gnd.n4721 gnd.n4720 0.152939
R17335 gnd.n4722 gnd.n4721 0.152939
R17336 gnd.n4723 gnd.n4722 0.152939
R17337 gnd.n4724 gnd.n4723 0.152939
R17338 gnd.n4726 gnd.n4724 0.152939
R17339 gnd.n4726 gnd.n4725 0.152939
R17340 gnd.n4725 gnd.n3683 0.152939
R17341 gnd.n5027 gnd.n3683 0.152939
R17342 gnd.n5028 gnd.n5027 0.152939
R17343 gnd.n5029 gnd.n5028 0.152939
R17344 gnd.n4038 gnd.n4037 0.152939
R17345 gnd.n4039 gnd.n4038 0.152939
R17346 gnd.n4039 gnd.n3921 0.152939
R17347 gnd.n4053 gnd.n3921 0.152939
R17348 gnd.n4054 gnd.n4053 0.152939
R17349 gnd.n4055 gnd.n4054 0.152939
R17350 gnd.n4055 gnd.n3908 0.152939
R17351 gnd.n4069 gnd.n3908 0.152939
R17352 gnd.n4070 gnd.n4069 0.152939
R17353 gnd.n4071 gnd.n4070 0.152939
R17354 gnd.n4072 gnd.n4071 0.152939
R17355 gnd.n4073 gnd.n4072 0.152939
R17356 gnd.n4074 gnd.n4073 0.152939
R17357 gnd.n4075 gnd.n4074 0.152939
R17358 gnd.n4076 gnd.n4075 0.152939
R17359 gnd.n4077 gnd.n4076 0.152939
R17360 gnd.n4078 gnd.n4077 0.152939
R17361 gnd.n4079 gnd.n4078 0.152939
R17362 gnd.n4080 gnd.n4079 0.152939
R17363 gnd.n4081 gnd.n4080 0.152939
R17364 gnd.n4082 gnd.n4081 0.152939
R17365 gnd.n4083 gnd.n4082 0.152939
R17366 gnd.n4084 gnd.n4083 0.152939
R17367 gnd.n4085 gnd.n4084 0.152939
R17368 gnd.n4086 gnd.n4085 0.152939
R17369 gnd.n4087 gnd.n4086 0.152939
R17370 gnd.n4088 gnd.n4087 0.152939
R17371 gnd.n4089 gnd.n4088 0.152939
R17372 gnd.n4030 gnd.n3937 0.152939
R17373 gnd.n3940 gnd.n3937 0.152939
R17374 gnd.n3941 gnd.n3940 0.152939
R17375 gnd.n3942 gnd.n3941 0.152939
R17376 gnd.n3945 gnd.n3942 0.152939
R17377 gnd.n3946 gnd.n3945 0.152939
R17378 gnd.n3947 gnd.n3946 0.152939
R17379 gnd.n3948 gnd.n3947 0.152939
R17380 gnd.n3951 gnd.n3948 0.152939
R17381 gnd.n3952 gnd.n3951 0.152939
R17382 gnd.n3953 gnd.n3952 0.152939
R17383 gnd.n3954 gnd.n3953 0.152939
R17384 gnd.n3957 gnd.n3954 0.152939
R17385 gnd.n3958 gnd.n3957 0.152939
R17386 gnd.n3959 gnd.n3958 0.152939
R17387 gnd.n3960 gnd.n3959 0.152939
R17388 gnd.n3963 gnd.n3960 0.152939
R17389 gnd.n3964 gnd.n3963 0.152939
R17390 gnd.n3965 gnd.n3964 0.152939
R17391 gnd.n3966 gnd.n3965 0.152939
R17392 gnd.n3969 gnd.n3966 0.152939
R17393 gnd.n3970 gnd.n3969 0.152939
R17394 gnd.n3973 gnd.n3970 0.152939
R17395 gnd.n3974 gnd.n3973 0.152939
R17396 gnd.n3976 gnd.n3974 0.152939
R17397 gnd.n3976 gnd.n3933 0.152939
R17398 gnd.n2326 gnd.n2321 0.152939
R17399 gnd.n2327 gnd.n2326 0.152939
R17400 gnd.n2328 gnd.n2327 0.152939
R17401 gnd.n2333 gnd.n2328 0.152939
R17402 gnd.n2334 gnd.n2333 0.152939
R17403 gnd.n2335 gnd.n2334 0.152939
R17404 gnd.n2336 gnd.n2335 0.152939
R17405 gnd.n2341 gnd.n2336 0.152939
R17406 gnd.n2342 gnd.n2341 0.152939
R17407 gnd.n2343 gnd.n2342 0.152939
R17408 gnd.n2344 gnd.n2343 0.152939
R17409 gnd.n2349 gnd.n2344 0.152939
R17410 gnd.n2350 gnd.n2349 0.152939
R17411 gnd.n2351 gnd.n2350 0.152939
R17412 gnd.n2352 gnd.n2351 0.152939
R17413 gnd.n2357 gnd.n2352 0.152939
R17414 gnd.n2358 gnd.n2357 0.152939
R17415 gnd.n2359 gnd.n2358 0.152939
R17416 gnd.n2360 gnd.n2359 0.152939
R17417 gnd.n2365 gnd.n2360 0.152939
R17418 gnd.n2366 gnd.n2365 0.152939
R17419 gnd.n2367 gnd.n2366 0.152939
R17420 gnd.n2368 gnd.n2367 0.152939
R17421 gnd.n2373 gnd.n2368 0.152939
R17422 gnd.n2374 gnd.n2373 0.152939
R17423 gnd.n2375 gnd.n2374 0.152939
R17424 gnd.n2376 gnd.n2375 0.152939
R17425 gnd.n2381 gnd.n2376 0.152939
R17426 gnd.n2382 gnd.n2381 0.152939
R17427 gnd.n2383 gnd.n2382 0.152939
R17428 gnd.n2384 gnd.n2383 0.152939
R17429 gnd.n2389 gnd.n2384 0.152939
R17430 gnd.n2390 gnd.n2389 0.152939
R17431 gnd.n2391 gnd.n2390 0.152939
R17432 gnd.n2392 gnd.n2391 0.152939
R17433 gnd.n2397 gnd.n2392 0.152939
R17434 gnd.n2398 gnd.n2397 0.152939
R17435 gnd.n2399 gnd.n2398 0.152939
R17436 gnd.n2400 gnd.n2399 0.152939
R17437 gnd.n2405 gnd.n2400 0.152939
R17438 gnd.n2406 gnd.n2405 0.152939
R17439 gnd.n2407 gnd.n2406 0.152939
R17440 gnd.n2408 gnd.n2407 0.152939
R17441 gnd.n2413 gnd.n2408 0.152939
R17442 gnd.n2414 gnd.n2413 0.152939
R17443 gnd.n2415 gnd.n2414 0.152939
R17444 gnd.n2416 gnd.n2415 0.152939
R17445 gnd.n2421 gnd.n2416 0.152939
R17446 gnd.n2422 gnd.n2421 0.152939
R17447 gnd.n2423 gnd.n2422 0.152939
R17448 gnd.n2424 gnd.n2423 0.152939
R17449 gnd.n2429 gnd.n2424 0.152939
R17450 gnd.n2430 gnd.n2429 0.152939
R17451 gnd.n2431 gnd.n2430 0.152939
R17452 gnd.n2432 gnd.n2431 0.152939
R17453 gnd.n2437 gnd.n2432 0.152939
R17454 gnd.n2438 gnd.n2437 0.152939
R17455 gnd.n2439 gnd.n2438 0.152939
R17456 gnd.n2440 gnd.n2439 0.152939
R17457 gnd.n2445 gnd.n2440 0.152939
R17458 gnd.n2446 gnd.n2445 0.152939
R17459 gnd.n2447 gnd.n2446 0.152939
R17460 gnd.n2448 gnd.n2447 0.152939
R17461 gnd.n2453 gnd.n2448 0.152939
R17462 gnd.n2454 gnd.n2453 0.152939
R17463 gnd.n2455 gnd.n2454 0.152939
R17464 gnd.n2456 gnd.n2455 0.152939
R17465 gnd.n2461 gnd.n2456 0.152939
R17466 gnd.n2462 gnd.n2461 0.152939
R17467 gnd.n2463 gnd.n2462 0.152939
R17468 gnd.n2464 gnd.n2463 0.152939
R17469 gnd.n2469 gnd.n2464 0.152939
R17470 gnd.n2470 gnd.n2469 0.152939
R17471 gnd.n2471 gnd.n2470 0.152939
R17472 gnd.n2472 gnd.n2471 0.152939
R17473 gnd.n2477 gnd.n2472 0.152939
R17474 gnd.n2478 gnd.n2477 0.152939
R17475 gnd.n2479 gnd.n2478 0.152939
R17476 gnd.n2480 gnd.n2479 0.152939
R17477 gnd.n2485 gnd.n2480 0.152939
R17478 gnd.n2486 gnd.n2485 0.152939
R17479 gnd.n2487 gnd.n2486 0.152939
R17480 gnd.n2488 gnd.n2487 0.152939
R17481 gnd.n2493 gnd.n2488 0.152939
R17482 gnd.n2494 gnd.n2493 0.152939
R17483 gnd.n2495 gnd.n2494 0.152939
R17484 gnd.n2496 gnd.n2495 0.152939
R17485 gnd.n2501 gnd.n2496 0.152939
R17486 gnd.n2502 gnd.n2501 0.152939
R17487 gnd.n2503 gnd.n2502 0.152939
R17488 gnd.n2504 gnd.n2503 0.152939
R17489 gnd.n2509 gnd.n2504 0.152939
R17490 gnd.n2510 gnd.n2509 0.152939
R17491 gnd.n2511 gnd.n2510 0.152939
R17492 gnd.n2512 gnd.n2511 0.152939
R17493 gnd.n2517 gnd.n2512 0.152939
R17494 gnd.n2518 gnd.n2517 0.152939
R17495 gnd.n2519 gnd.n2518 0.152939
R17496 gnd.n2520 gnd.n2519 0.152939
R17497 gnd.n2525 gnd.n2520 0.152939
R17498 gnd.n2526 gnd.n2525 0.152939
R17499 gnd.n2527 gnd.n2526 0.152939
R17500 gnd.n2528 gnd.n2527 0.152939
R17501 gnd.n2533 gnd.n2528 0.152939
R17502 gnd.n2534 gnd.n2533 0.152939
R17503 gnd.n2535 gnd.n2534 0.152939
R17504 gnd.n2536 gnd.n2535 0.152939
R17505 gnd.n2541 gnd.n2536 0.152939
R17506 gnd.n2542 gnd.n2541 0.152939
R17507 gnd.n2543 gnd.n2542 0.152939
R17508 gnd.n2544 gnd.n2543 0.152939
R17509 gnd.n2549 gnd.n2544 0.152939
R17510 gnd.n2550 gnd.n2549 0.152939
R17511 gnd.n2551 gnd.n2550 0.152939
R17512 gnd.n2552 gnd.n2551 0.152939
R17513 gnd.n2557 gnd.n2552 0.152939
R17514 gnd.n2558 gnd.n2557 0.152939
R17515 gnd.n2559 gnd.n2558 0.152939
R17516 gnd.n2560 gnd.n2559 0.152939
R17517 gnd.n2565 gnd.n2560 0.152939
R17518 gnd.n2566 gnd.n2565 0.152939
R17519 gnd.n2567 gnd.n2566 0.152939
R17520 gnd.n2568 gnd.n2567 0.152939
R17521 gnd.n2573 gnd.n2568 0.152939
R17522 gnd.n2574 gnd.n2573 0.152939
R17523 gnd.n2575 gnd.n2574 0.152939
R17524 gnd.n2576 gnd.n2575 0.152939
R17525 gnd.n2581 gnd.n2576 0.152939
R17526 gnd.n2582 gnd.n2581 0.152939
R17527 gnd.n2583 gnd.n2582 0.152939
R17528 gnd.n2584 gnd.n2583 0.152939
R17529 gnd.n2589 gnd.n2584 0.152939
R17530 gnd.n2590 gnd.n2589 0.152939
R17531 gnd.n2591 gnd.n2590 0.152939
R17532 gnd.n2592 gnd.n2591 0.152939
R17533 gnd.n2597 gnd.n2592 0.152939
R17534 gnd.n2598 gnd.n2597 0.152939
R17535 gnd.n2599 gnd.n2598 0.152939
R17536 gnd.n2600 gnd.n2599 0.152939
R17537 gnd.n2605 gnd.n2600 0.152939
R17538 gnd.n2606 gnd.n2605 0.152939
R17539 gnd.n2607 gnd.n2606 0.152939
R17540 gnd.n2608 gnd.n2607 0.152939
R17541 gnd.n2613 gnd.n2608 0.152939
R17542 gnd.n2614 gnd.n2613 0.152939
R17543 gnd.n2615 gnd.n2614 0.152939
R17544 gnd.n2616 gnd.n2615 0.152939
R17545 gnd.n2621 gnd.n2616 0.152939
R17546 gnd.n2622 gnd.n2621 0.152939
R17547 gnd.n2623 gnd.n2622 0.152939
R17548 gnd.n2624 gnd.n2623 0.152939
R17549 gnd.n2629 gnd.n2624 0.152939
R17550 gnd.n2630 gnd.n2629 0.152939
R17551 gnd.n2631 gnd.n2630 0.152939
R17552 gnd.n2632 gnd.n2631 0.152939
R17553 gnd.n2637 gnd.n2632 0.152939
R17554 gnd.n2638 gnd.n2637 0.152939
R17555 gnd.n2639 gnd.n2638 0.152939
R17556 gnd.n2640 gnd.n2639 0.152939
R17557 gnd.n2645 gnd.n2640 0.152939
R17558 gnd.n2646 gnd.n2645 0.152939
R17559 gnd.n2647 gnd.n2646 0.152939
R17560 gnd.n2648 gnd.n2647 0.152939
R17561 gnd.n2653 gnd.n2648 0.152939
R17562 gnd.n2654 gnd.n2653 0.152939
R17563 gnd.n2655 gnd.n2654 0.152939
R17564 gnd.n2656 gnd.n2655 0.152939
R17565 gnd.n2661 gnd.n2656 0.152939
R17566 gnd.n2662 gnd.n2661 0.152939
R17567 gnd.n3033 gnd.n2662 0.152939
R17568 gnd.n3032 gnd.n2663 0.152939
R17569 gnd.n2668 gnd.n2663 0.152939
R17570 gnd.n2669 gnd.n2668 0.152939
R17571 gnd.n2670 gnd.n2669 0.152939
R17572 gnd.n2675 gnd.n2670 0.152939
R17573 gnd.n2676 gnd.n2675 0.152939
R17574 gnd.n2677 gnd.n2676 0.152939
R17575 gnd.n2678 gnd.n2677 0.152939
R17576 gnd.n2683 gnd.n2678 0.152939
R17577 gnd.n2684 gnd.n2683 0.152939
R17578 gnd.n2685 gnd.n2684 0.152939
R17579 gnd.n2686 gnd.n2685 0.152939
R17580 gnd.n2691 gnd.n2686 0.152939
R17581 gnd.n2692 gnd.n2691 0.152939
R17582 gnd.n2693 gnd.n2692 0.152939
R17583 gnd.n2694 gnd.n2693 0.152939
R17584 gnd.n2699 gnd.n2694 0.152939
R17585 gnd.n2700 gnd.n2699 0.152939
R17586 gnd.n2701 gnd.n2700 0.152939
R17587 gnd.n2702 gnd.n2701 0.152939
R17588 gnd.n2707 gnd.n2702 0.152939
R17589 gnd.n2708 gnd.n2707 0.152939
R17590 gnd.n2709 gnd.n2708 0.152939
R17591 gnd.n2710 gnd.n2709 0.152939
R17592 gnd.n2715 gnd.n2710 0.152939
R17593 gnd.n2716 gnd.n2715 0.152939
R17594 gnd.n2717 gnd.n2716 0.152939
R17595 gnd.n2718 gnd.n2717 0.152939
R17596 gnd.n2723 gnd.n2718 0.152939
R17597 gnd.n2724 gnd.n2723 0.152939
R17598 gnd.n2725 gnd.n2724 0.152939
R17599 gnd.n2726 gnd.n2725 0.152939
R17600 gnd.n2731 gnd.n2726 0.152939
R17601 gnd.n2732 gnd.n2731 0.152939
R17602 gnd.n2733 gnd.n2732 0.152939
R17603 gnd.n2734 gnd.n2733 0.152939
R17604 gnd.n2739 gnd.n2734 0.152939
R17605 gnd.n2740 gnd.n2739 0.152939
R17606 gnd.n2741 gnd.n2740 0.152939
R17607 gnd.n2742 gnd.n2741 0.152939
R17608 gnd.n2747 gnd.n2742 0.152939
R17609 gnd.n2748 gnd.n2747 0.152939
R17610 gnd.n2749 gnd.n2748 0.152939
R17611 gnd.n2750 gnd.n2749 0.152939
R17612 gnd.n2755 gnd.n2750 0.152939
R17613 gnd.n2756 gnd.n2755 0.152939
R17614 gnd.n2757 gnd.n2756 0.152939
R17615 gnd.n2758 gnd.n2757 0.152939
R17616 gnd.n2763 gnd.n2758 0.152939
R17617 gnd.n2764 gnd.n2763 0.152939
R17618 gnd.n2765 gnd.n2764 0.152939
R17619 gnd.n2766 gnd.n2765 0.152939
R17620 gnd.n2771 gnd.n2766 0.152939
R17621 gnd.n2772 gnd.n2771 0.152939
R17622 gnd.n2773 gnd.n2772 0.152939
R17623 gnd.n2774 gnd.n2773 0.152939
R17624 gnd.n2779 gnd.n2774 0.152939
R17625 gnd.n2780 gnd.n2779 0.152939
R17626 gnd.n2781 gnd.n2780 0.152939
R17627 gnd.n2782 gnd.n2781 0.152939
R17628 gnd.n2787 gnd.n2782 0.152939
R17629 gnd.n2788 gnd.n2787 0.152939
R17630 gnd.n2789 gnd.n2788 0.152939
R17631 gnd.n2790 gnd.n2789 0.152939
R17632 gnd.n2793 gnd.n2790 0.152939
R17633 gnd.n2896 gnd.n2793 0.152939
R17634 gnd.n2811 gnd.n941 0.152939
R17635 gnd.n2812 gnd.n2811 0.152939
R17636 gnd.n2813 gnd.n2812 0.152939
R17637 gnd.n2813 gnd.n2802 0.152939
R17638 gnd.n2819 gnd.n2802 0.152939
R17639 gnd.n2820 gnd.n2819 0.152939
R17640 gnd.n2821 gnd.n2820 0.152939
R17641 gnd.n2821 gnd.n2798 0.152939
R17642 gnd.n2827 gnd.n2798 0.152939
R17643 gnd.n2828 gnd.n2827 0.152939
R17644 gnd.n2830 gnd.n2828 0.152939
R17645 gnd.n2830 gnd.n2829 0.152939
R17646 gnd.n2829 gnd.n2794 0.152939
R17647 gnd.n2895 gnd.n2794 0.152939
R17648 gnd.n7146 gnd.n649 0.152939
R17649 gnd.n7147 gnd.n7146 0.152939
R17650 gnd.n7148 gnd.n7147 0.152939
R17651 gnd.n7148 gnd.n632 0.152939
R17652 gnd.n7162 gnd.n632 0.152939
R17653 gnd.n7163 gnd.n7162 0.152939
R17654 gnd.n7164 gnd.n7163 0.152939
R17655 gnd.n7164 gnd.n615 0.152939
R17656 gnd.n7178 gnd.n615 0.152939
R17657 gnd.n7179 gnd.n7178 0.152939
R17658 gnd.n7180 gnd.n7179 0.152939
R17659 gnd.n7180 gnd.n599 0.152939
R17660 gnd.n7194 gnd.n599 0.152939
R17661 gnd.n7195 gnd.n7194 0.152939
R17662 gnd.n7196 gnd.n7195 0.152939
R17663 gnd.n7196 gnd.n580 0.152939
R17664 gnd.n7278 gnd.n580 0.152939
R17665 gnd.n7279 gnd.n7278 0.152939
R17666 gnd.n7280 gnd.n7279 0.152939
R17667 gnd.n7280 gnd.n507 0.152939
R17668 gnd.n7350 gnd.n507 0.152939
R17669 gnd.n7349 gnd.n508 0.152939
R17670 gnd.n510 gnd.n508 0.152939
R17671 gnd.n514 gnd.n510 0.152939
R17672 gnd.n515 gnd.n514 0.152939
R17673 gnd.n516 gnd.n515 0.152939
R17674 gnd.n517 gnd.n516 0.152939
R17675 gnd.n521 gnd.n517 0.152939
R17676 gnd.n522 gnd.n521 0.152939
R17677 gnd.n523 gnd.n522 0.152939
R17678 gnd.n524 gnd.n523 0.152939
R17679 gnd.n528 gnd.n524 0.152939
R17680 gnd.n529 gnd.n528 0.152939
R17681 gnd.n530 gnd.n529 0.152939
R17682 gnd.n531 gnd.n530 0.152939
R17683 gnd.n538 gnd.n531 0.152939
R17684 gnd.n539 gnd.n538 0.152939
R17685 gnd.n540 gnd.n539 0.152939
R17686 gnd.n541 gnd.n540 0.152939
R17687 gnd.n545 gnd.n541 0.152939
R17688 gnd.n546 gnd.n545 0.152939
R17689 gnd.n547 gnd.n546 0.152939
R17690 gnd.n548 gnd.n547 0.152939
R17691 gnd.n552 gnd.n548 0.152939
R17692 gnd.n553 gnd.n552 0.152939
R17693 gnd.n554 gnd.n553 0.152939
R17694 gnd.n555 gnd.n554 0.152939
R17695 gnd.n559 gnd.n555 0.152939
R17696 gnd.n560 gnd.n559 0.152939
R17697 gnd.n561 gnd.n560 0.152939
R17698 gnd.n562 gnd.n561 0.152939
R17699 gnd.n566 gnd.n562 0.152939
R17700 gnd.n567 gnd.n566 0.152939
R17701 gnd.n7290 gnd.n567 0.152939
R17702 gnd.n7290 gnd.n7289 0.152939
R17703 gnd.n6898 gnd.n903 0.152939
R17704 gnd.n905 gnd.n903 0.152939
R17705 gnd.n906 gnd.n905 0.152939
R17706 gnd.n6757 gnd.n906 0.152939
R17707 gnd.n6761 gnd.n6757 0.152939
R17708 gnd.n6762 gnd.n6761 0.152939
R17709 gnd.n6763 gnd.n6762 0.152939
R17710 gnd.n6763 gnd.n6755 0.152939
R17711 gnd.n6771 gnd.n6755 0.152939
R17712 gnd.n6772 gnd.n6771 0.152939
R17713 gnd.n6773 gnd.n6772 0.152939
R17714 gnd.n6773 gnd.n6753 0.152939
R17715 gnd.n6781 gnd.n6753 0.152939
R17716 gnd.n6782 gnd.n6781 0.152939
R17717 gnd.n6783 gnd.n6782 0.152939
R17718 gnd.n6784 gnd.n6783 0.152939
R17719 gnd.n6785 gnd.n6784 0.152939
R17720 gnd.n6786 gnd.n6785 0.152939
R17721 gnd.n6787 gnd.n6786 0.152939
R17722 gnd.n6788 gnd.n6787 0.152939
R17723 gnd.n6789 gnd.n6788 0.152939
R17724 gnd.n6790 gnd.n6789 0.152939
R17725 gnd.n6792 gnd.n6790 0.152939
R17726 gnd.n6792 gnd.n6791 0.152939
R17727 gnd.n6791 gnd.n932 0.152939
R17728 gnd.n932 gnd.n671 0.152939
R17729 gnd.n933 gnd.n671 0.152939
R17730 gnd.n934 gnd.n933 0.152939
R17731 gnd.n935 gnd.n934 0.152939
R17732 gnd.n2838 gnd.n935 0.152939
R17733 gnd.n2839 gnd.n2838 0.152939
R17734 gnd.n2839 gnd.n2837 0.152939
R17735 gnd.n2847 gnd.n2837 0.152939
R17736 gnd.n2848 gnd.n2847 0.152939
R17737 gnd.n2849 gnd.n2848 0.152939
R17738 gnd.n2849 gnd.n2835 0.152939
R17739 gnd.n2857 gnd.n2835 0.152939
R17740 gnd.n2858 gnd.n2857 0.152939
R17741 gnd.n2859 gnd.n2858 0.152939
R17742 gnd.n2859 gnd.n2833 0.152939
R17743 gnd.n2867 gnd.n2833 0.152939
R17744 gnd.n2868 gnd.n2867 0.152939
R17745 gnd.n2869 gnd.n2868 0.152939
R17746 gnd.n2870 gnd.n2869 0.152939
R17747 gnd.n2871 gnd.n2870 0.152939
R17748 gnd.n2872 gnd.n2871 0.152939
R17749 gnd.n2873 gnd.n2872 0.152939
R17750 gnd.n2874 gnd.n2873 0.152939
R17751 gnd.n2876 gnd.n2874 0.152939
R17752 gnd.n2876 gnd.n2875 0.152939
R17753 gnd.n2875 gnd.n573 0.152939
R17754 gnd.n7288 gnd.n573 0.152939
R17755 gnd.n864 gnd.n784 0.152939
R17756 gnd.n865 gnd.n864 0.152939
R17757 gnd.n866 gnd.n865 0.152939
R17758 gnd.n867 gnd.n866 0.152939
R17759 gnd.n868 gnd.n867 0.152939
R17760 gnd.n869 gnd.n868 0.152939
R17761 gnd.n870 gnd.n869 0.152939
R17762 gnd.n871 gnd.n870 0.152939
R17763 gnd.n872 gnd.n871 0.152939
R17764 gnd.n873 gnd.n872 0.152939
R17765 gnd.n874 gnd.n873 0.152939
R17766 gnd.n875 gnd.n874 0.152939
R17767 gnd.n876 gnd.n875 0.152939
R17768 gnd.n883 gnd.n882 0.152939
R17769 gnd.n884 gnd.n883 0.152939
R17770 gnd.n885 gnd.n884 0.152939
R17771 gnd.n886 gnd.n885 0.152939
R17772 gnd.n887 gnd.n886 0.152939
R17773 gnd.n888 gnd.n887 0.152939
R17774 gnd.n889 gnd.n888 0.152939
R17775 gnd.n890 gnd.n889 0.152939
R17776 gnd.n891 gnd.n890 0.152939
R17777 gnd.n892 gnd.n891 0.152939
R17778 gnd.n893 gnd.n892 0.152939
R17779 gnd.n894 gnd.n893 0.152939
R17780 gnd.n895 gnd.n894 0.152939
R17781 gnd.n896 gnd.n895 0.152939
R17782 gnd.n897 gnd.n896 0.152939
R17783 gnd.n6903 gnd.n897 0.152939
R17784 gnd.n6903 gnd.n6902 0.152939
R17785 gnd.n6902 gnd.n6901 0.152939
R17786 gnd.n7019 gnd.n7018 0.152939
R17787 gnd.n7020 gnd.n7019 0.152939
R17788 gnd.n7020 gnd.n767 0.152939
R17789 gnd.n7034 gnd.n767 0.152939
R17790 gnd.n7035 gnd.n7034 0.152939
R17791 gnd.n7036 gnd.n7035 0.152939
R17792 gnd.n7036 gnd.n749 0.152939
R17793 gnd.n7050 gnd.n749 0.152939
R17794 gnd.n7051 gnd.n7050 0.152939
R17795 gnd.n7052 gnd.n7051 0.152939
R17796 gnd.n7052 gnd.n731 0.152939
R17797 gnd.n7066 gnd.n731 0.152939
R17798 gnd.n7067 gnd.n7066 0.152939
R17799 gnd.n7068 gnd.n7067 0.152939
R17800 gnd.n7068 gnd.n714 0.152939
R17801 gnd.n7082 gnd.n714 0.152939
R17802 gnd.n7083 gnd.n7082 0.152939
R17803 gnd.n7085 gnd.n7083 0.152939
R17804 gnd.n7085 gnd.n7084 0.152939
R17805 gnd.n7084 gnd.n697 0.152939
R17806 gnd.n697 gnd.n649 0.152939
R17807 gnd.n5465 gnd.n5464 0.152939
R17808 gnd.n5466 gnd.n5465 0.152939
R17809 gnd.n5466 gnd.n5455 0.152939
R17810 gnd.n5472 gnd.n5455 0.152939
R17811 gnd.n5473 gnd.n5472 0.152939
R17812 gnd.n5474 gnd.n5473 0.152939
R17813 gnd.n5474 gnd.n5451 0.152939
R17814 gnd.n5517 gnd.n5451 0.152939
R17815 gnd.n5518 gnd.n5517 0.152939
R17816 gnd.n5519 gnd.n5518 0.152939
R17817 gnd.n5519 gnd.n5447 0.152939
R17818 gnd.n5525 gnd.n5447 0.152939
R17819 gnd.n5526 gnd.n5525 0.152939
R17820 gnd.n5527 gnd.n5526 0.152939
R17821 gnd.n5527 gnd.n5443 0.152939
R17822 gnd.n5533 gnd.n5443 0.152939
R17823 gnd.n5534 gnd.n5533 0.152939
R17824 gnd.n5535 gnd.n5534 0.152939
R17825 gnd.n5536 gnd.n5535 0.152939
R17826 gnd.n5537 gnd.n5536 0.152939
R17827 gnd.n5540 gnd.n5537 0.152939
R17828 gnd.n5541 gnd.n5540 0.152939
R17829 gnd.n5542 gnd.n5541 0.152939
R17830 gnd.n5543 gnd.n5542 0.152939
R17831 gnd.n5543 gnd.n1672 0.152939
R17832 gnd.n5813 gnd.n1672 0.152939
R17833 gnd.n5814 gnd.n5813 0.152939
R17834 gnd.n5815 gnd.n5814 0.152939
R17835 gnd.n5815 gnd.n1660 0.152939
R17836 gnd.n5833 gnd.n1660 0.152939
R17837 gnd.n5834 gnd.n5833 0.152939
R17838 gnd.n5835 gnd.n5834 0.152939
R17839 gnd.n5835 gnd.n1647 0.152939
R17840 gnd.n5853 gnd.n1647 0.152939
R17841 gnd.n5854 gnd.n5853 0.152939
R17842 gnd.n5855 gnd.n5854 0.152939
R17843 gnd.n5856 gnd.n5855 0.152939
R17844 gnd.n5856 gnd.n1429 0.152939
R17845 gnd.n6064 gnd.n1429 0.152939
R17846 gnd.n6065 gnd.n6064 0.152939
R17847 gnd.n6066 gnd.n6065 0.152939
R17848 gnd.n6067 gnd.n6066 0.152939
R17849 gnd.n6067 gnd.n1396 0.152939
R17850 gnd.n6146 gnd.n1396 0.152939
R17851 gnd.n6147 gnd.n6146 0.152939
R17852 gnd.n6148 gnd.n6147 0.152939
R17853 gnd.n6148 gnd.n1372 0.152939
R17854 gnd.n6174 gnd.n1372 0.152939
R17855 gnd.n6175 gnd.n6174 0.152939
R17856 gnd.n6176 gnd.n6175 0.152939
R17857 gnd.n6177 gnd.n6176 0.152939
R17858 gnd.n6178 gnd.n6177 0.152939
R17859 gnd.n6181 gnd.n6178 0.152939
R17860 gnd.n6182 gnd.n6181 0.152939
R17861 gnd.n6183 gnd.n6182 0.152939
R17862 gnd.n6183 gnd.n1311 0.152939
R17863 gnd.n6285 gnd.n1311 0.152939
R17864 gnd.n6286 gnd.n6285 0.152939
R17865 gnd.n6287 gnd.n6286 0.152939
R17866 gnd.n6288 gnd.n6287 0.152939
R17867 gnd.n6289 gnd.n6288 0.152939
R17868 gnd.n6291 gnd.n6289 0.152939
R17869 gnd.n6293 gnd.n6291 0.152939
R17870 gnd.n6293 gnd.n6292 0.152939
R17871 gnd.n6292 gnd.n1269 0.152939
R17872 gnd.n1270 gnd.n1269 0.152939
R17873 gnd.n1272 gnd.n1270 0.152939
R17874 gnd.n1272 gnd.n1271 0.152939
R17875 gnd.n1271 gnd.n1240 0.152939
R17876 gnd.n1241 gnd.n1240 0.152939
R17877 gnd.n1243 gnd.n1241 0.152939
R17878 gnd.n1243 gnd.n1242 0.152939
R17879 gnd.n1242 gnd.n1211 0.152939
R17880 gnd.n1212 gnd.n1211 0.152939
R17881 gnd.n1213 gnd.n1212 0.152939
R17882 gnd.n1214 gnd.n1213 0.152939
R17883 gnd.n1214 gnd.n1106 0.152939
R17884 gnd.n6614 gnd.n1106 0.152939
R17885 gnd.n6615 gnd.n6614 0.152939
R17886 gnd.n6616 gnd.n6615 0.152939
R17887 gnd.n6617 gnd.n6616 0.152939
R17888 gnd.n6617 gnd.n1080 0.152939
R17889 gnd.n6644 gnd.n1080 0.152939
R17890 gnd.n6645 gnd.n6644 0.152939
R17891 gnd.n6646 gnd.n6645 0.152939
R17892 gnd.n6647 gnd.n6646 0.152939
R17893 gnd.n6647 gnd.n1055 0.152939
R17894 gnd.n6675 gnd.n1055 0.152939
R17895 gnd.n6676 gnd.n6675 0.152939
R17896 gnd.n6677 gnd.n6676 0.152939
R17897 gnd.n6678 gnd.n6677 0.152939
R17898 gnd.n6679 gnd.n6678 0.152939
R17899 gnd.n6681 gnd.n6679 0.152939
R17900 gnd.n6682 gnd.n6681 0.152939
R17901 gnd.n6682 gnd.n970 0.152939
R17902 gnd.n6716 gnd.n970 0.152939
R17903 gnd.n6717 gnd.n6716 0.152939
R17904 gnd.n6718 gnd.n6717 0.152939
R17905 gnd.n6718 gnd.n966 0.152939
R17906 gnd.n6724 gnd.n966 0.152939
R17907 gnd.n6725 gnd.n6724 0.152939
R17908 gnd.n6726 gnd.n6725 0.152939
R17909 gnd.n6726 gnd.n962 0.152939
R17910 gnd.n6732 gnd.n962 0.152939
R17911 gnd.n6733 gnd.n6732 0.152939
R17912 gnd.n6734 gnd.n6733 0.152939
R17913 gnd.n6734 gnd.n958 0.152939
R17914 gnd.n6740 gnd.n958 0.152939
R17915 gnd.n6741 gnd.n6740 0.152939
R17916 gnd.n6742 gnd.n6741 0.152939
R17917 gnd.n6742 gnd.n954 0.152939
R17918 gnd.n6748 gnd.n954 0.152939
R17919 gnd.n6749 gnd.n6748 0.152939
R17920 gnd.n6750 gnd.n6749 0.152939
R17921 gnd.n6750 gnd.n950 0.152939
R17922 gnd.n6817 gnd.n950 0.152939
R17923 gnd.n6818 gnd.n6817 0.152939
R17924 gnd.n6819 gnd.n6818 0.152939
R17925 gnd.n6819 gnd.n945 0.152939
R17926 gnd.n6837 gnd.n945 0.152939
R17927 gnd.n5240 gnd.n2039 0.152939
R17928 gnd.n2040 gnd.n2039 0.152939
R17929 gnd.n2041 gnd.n2040 0.152939
R17930 gnd.n2042 gnd.n2041 0.152939
R17931 gnd.n2043 gnd.n2042 0.152939
R17932 gnd.n2044 gnd.n2043 0.152939
R17933 gnd.n2045 gnd.n2044 0.152939
R17934 gnd.n2193 gnd.n2045 0.152939
R17935 gnd.n2194 gnd.n2193 0.152939
R17936 gnd.n2195 gnd.n2194 0.152939
R17937 gnd.n2196 gnd.n2195 0.152939
R17938 gnd.n2197 gnd.n2196 0.152939
R17939 gnd.n2197 gnd.n1947 0.152939
R17940 gnd.n5351 gnd.n1947 0.152939
R17941 gnd.n5352 gnd.n5351 0.152939
R17942 gnd.n5353 gnd.n5352 0.152939
R17943 gnd.n5354 gnd.n5353 0.152939
R17944 gnd.n5355 gnd.n5354 0.152939
R17945 gnd.n5355 gnd.n1907 0.152939
R17946 gnd.n5391 gnd.n1907 0.152939
R17947 gnd.n5392 gnd.n5391 0.152939
R17948 gnd.n5394 gnd.n5392 0.152939
R17949 gnd.n5394 gnd.n5393 0.152939
R17950 gnd.n5393 gnd.n1898 0.152939
R17951 gnd.n5409 gnd.n1898 0.152939
R17952 gnd.n5277 gnd.n2016 0.152939
R17953 gnd.n2019 gnd.n2016 0.152939
R17954 gnd.n2020 gnd.n2019 0.152939
R17955 gnd.n2021 gnd.n2020 0.152939
R17956 gnd.n2022 gnd.n2021 0.152939
R17957 gnd.n2025 gnd.n2022 0.152939
R17958 gnd.n2026 gnd.n2025 0.152939
R17959 gnd.n2027 gnd.n2026 0.152939
R17960 gnd.n2028 gnd.n2027 0.152939
R17961 gnd.n2031 gnd.n2028 0.152939
R17962 gnd.n2032 gnd.n2031 0.152939
R17963 gnd.n2033 gnd.n2032 0.152939
R17964 gnd.n2034 gnd.n2033 0.152939
R17965 gnd.n2038 gnd.n2034 0.152939
R17966 gnd.n5242 gnd.n2038 0.152939
R17967 gnd.n5242 gnd.n5241 0.152939
R17968 gnd.n5278 gnd.n2002 0.152939
R17969 gnd.n5292 gnd.n2002 0.152939
R17970 gnd.n5293 gnd.n5292 0.152939
R17971 gnd.n5294 gnd.n5293 0.152939
R17972 gnd.n5294 gnd.n1984 0.152939
R17973 gnd.n5308 gnd.n1984 0.152939
R17974 gnd.n5309 gnd.n5308 0.152939
R17975 gnd.n5310 gnd.n5309 0.152939
R17976 gnd.n5310 gnd.n1967 0.152939
R17977 gnd.n5324 gnd.n1967 0.152939
R17978 gnd.n5325 gnd.n5324 0.152939
R17979 gnd.n5326 gnd.n5325 0.152939
R17980 gnd.n5327 gnd.n5326 0.152939
R17981 gnd.n5328 gnd.n5327 0.152939
R17982 gnd.n5330 gnd.n5328 0.152939
R17983 gnd.n5330 gnd.n5329 0.152939
R17984 gnd.n5329 gnd.n1928 0.152939
R17985 gnd.n1929 gnd.n1928 0.152939
R17986 gnd.n1930 gnd.n1929 0.152939
R17987 gnd.n1931 gnd.n1930 0.152939
R17988 gnd.n1933 gnd.n1931 0.152939
R17989 gnd.n1933 gnd.n1932 0.152939
R17990 gnd.n1932 gnd.n1854 0.152939
R17991 gnd.n1855 gnd.n1854 0.152939
R17992 gnd.n1856 gnd.n1855 0.152939
R17993 gnd.n5607 gnd.n1856 0.152939
R17994 gnd.n5608 gnd.n5607 0.152939
R17995 gnd.n5613 gnd.n5608 0.152939
R17996 gnd.n5614 gnd.n5613 0.152939
R17997 gnd.n5615 gnd.n5614 0.152939
R17998 gnd.n5615 gnd.n1829 0.152939
R17999 gnd.n5655 gnd.n1829 0.152939
R18000 gnd.n5656 gnd.n5655 0.152939
R18001 gnd.n5657 gnd.n5656 0.152939
R18002 gnd.n5657 gnd.n1811 0.152939
R18003 gnd.n5671 gnd.n1811 0.152939
R18004 gnd.n5672 gnd.n5671 0.152939
R18005 gnd.n5673 gnd.n5672 0.152939
R18006 gnd.n5673 gnd.n1794 0.152939
R18007 gnd.n5687 gnd.n1794 0.152939
R18008 gnd.n5688 gnd.n5687 0.152939
R18009 gnd.n5689 gnd.n5688 0.152939
R18010 gnd.n5689 gnd.n1776 0.152939
R18011 gnd.n5703 gnd.n1776 0.152939
R18012 gnd.n5704 gnd.n5703 0.152939
R18013 gnd.n5705 gnd.n5704 0.152939
R18014 gnd.n5706 gnd.n5705 0.152939
R18015 gnd.n5708 gnd.n5706 0.152939
R18016 gnd.n5708 gnd.n5707 0.152939
R18017 gnd.n5707 gnd.n1617 0.152939
R18018 gnd.n1618 gnd.n1617 0.152939
R18019 gnd.n5899 gnd.n1618 0.152939
R18020 gnd.n5649 gnd.n5648 0.152939
R18021 gnd.n5649 gnd.n1820 0.152939
R18022 gnd.n5663 gnd.n1820 0.152939
R18023 gnd.n5664 gnd.n5663 0.152939
R18024 gnd.n5665 gnd.n5664 0.152939
R18025 gnd.n5665 gnd.n1803 0.152939
R18026 gnd.n5679 gnd.n1803 0.152939
R18027 gnd.n5680 gnd.n5679 0.152939
R18028 gnd.n5681 gnd.n5680 0.152939
R18029 gnd.n5681 gnd.n1785 0.152939
R18030 gnd.n5695 gnd.n1785 0.152939
R18031 gnd.n5696 gnd.n5695 0.152939
R18032 gnd.n5697 gnd.n5696 0.152939
R18033 gnd.n5697 gnd.n1766 0.152939
R18034 gnd.n5716 gnd.n1766 0.152939
R18035 gnd.n5717 gnd.n5716 0.152939
R18036 gnd.n5718 gnd.n5717 0.152939
R18037 gnd.n5718 gnd.n1608 0.152939
R18038 gnd.n5907 gnd.n1608 0.152939
R18039 gnd.n5908 gnd.n5907 0.152939
R18040 gnd.n5955 gnd.n5908 0.152939
R18041 gnd.n5954 gnd.n5909 0.152939
R18042 gnd.n5913 gnd.n5909 0.152939
R18043 gnd.n5914 gnd.n5913 0.152939
R18044 gnd.n5915 gnd.n5914 0.152939
R18045 gnd.n5916 gnd.n5915 0.152939
R18046 gnd.n5917 gnd.n5916 0.152939
R18047 gnd.n5921 gnd.n5917 0.152939
R18048 gnd.n5922 gnd.n5921 0.152939
R18049 gnd.n5923 gnd.n5922 0.152939
R18050 gnd.n5924 gnd.n5923 0.152939
R18051 gnd.n5929 gnd.n5924 0.152939
R18052 gnd.n5930 gnd.n5929 0.152939
R18053 gnd.n5930 gnd.n1562 0.152939
R18054 gnd.n5995 gnd.n5994 0.152939
R18055 gnd.n5994 gnd.n1563 0.152939
R18056 gnd.n1570 gnd.n1563 0.152939
R18057 gnd.n1571 gnd.n1570 0.152939
R18058 gnd.n1572 gnd.n1571 0.152939
R18059 gnd.n1573 gnd.n1572 0.152939
R18060 gnd.n1577 gnd.n1573 0.152939
R18061 gnd.n1578 gnd.n1577 0.152939
R18062 gnd.n1579 gnd.n1578 0.152939
R18063 gnd.n1580 gnd.n1579 0.152939
R18064 gnd.n1584 gnd.n1580 0.152939
R18065 gnd.n1585 gnd.n1584 0.152939
R18066 gnd.n1586 gnd.n1585 0.152939
R18067 gnd.n1587 gnd.n1586 0.152939
R18068 gnd.n1591 gnd.n1587 0.152939
R18069 gnd.n1592 gnd.n1591 0.152939
R18070 gnd.n5963 gnd.n1592 0.152939
R18071 gnd.n5963 gnd.n5962 0.152939
R18072 gnd.n2179 gnd.n2175 0.152939
R18073 gnd.n2180 gnd.n2179 0.152939
R18074 gnd.n2181 gnd.n2180 0.152939
R18075 gnd.n2181 gnd.n2048 0.152939
R18076 gnd.n2187 gnd.n2048 0.152939
R18077 gnd.n2188 gnd.n2187 0.152939
R18078 gnd.n2189 gnd.n2188 0.152939
R18079 gnd.n2190 gnd.n2189 0.152939
R18080 gnd.n2191 gnd.n2190 0.152939
R18081 gnd.n2199 gnd.n2191 0.152939
R18082 gnd.n2200 gnd.n2199 0.152939
R18083 gnd.n2201 gnd.n2200 0.152939
R18084 gnd.n2202 gnd.n2201 0.152939
R18085 gnd.n2204 gnd.n2202 0.152939
R18086 gnd.n2204 gnd.n2203 0.152939
R18087 gnd.n2203 gnd.n1941 0.152939
R18088 gnd.n5366 gnd.n1941 0.152939
R18089 gnd.n5367 gnd.n5366 0.152939
R18090 gnd.n5368 gnd.n5367 0.152939
R18091 gnd.n5369 gnd.n5368 0.152939
R18092 gnd.n5369 gnd.n1901 0.152939
R18093 gnd.n5400 gnd.n1901 0.152939
R18094 gnd.n5401 gnd.n5400 0.152939
R18095 gnd.n5402 gnd.n5401 0.152939
R18096 gnd.n5402 gnd.n1886 0.152939
R18097 gnd.n5606 gnd.n1886 0.152939
R18098 gnd.n5606 gnd.n1887 0.152939
R18099 gnd.n1889 gnd.n1887 0.152939
R18100 gnd.n1890 gnd.n1889 0.152939
R18101 gnd.n1891 gnd.n1890 0.152939
R18102 gnd.n1892 gnd.n1891 0.152939
R18103 gnd.n5478 gnd.n1892 0.152939
R18104 gnd.n5479 gnd.n5478 0.152939
R18105 gnd.n5479 gnd.n5477 0.152939
R18106 gnd.n5487 gnd.n5477 0.152939
R18107 gnd.n5488 gnd.n5487 0.152939
R18108 gnd.n5489 gnd.n5488 0.152939
R18109 gnd.n5490 gnd.n5489 0.152939
R18110 gnd.n5491 gnd.n5490 0.152939
R18111 gnd.n5492 gnd.n5491 0.152939
R18112 gnd.n5493 gnd.n5492 0.152939
R18113 gnd.n5494 gnd.n5493 0.152939
R18114 gnd.n5496 gnd.n5494 0.152939
R18115 gnd.n5496 gnd.n5495 0.152939
R18116 gnd.n5495 gnd.n5433 0.152939
R18117 gnd.n5434 gnd.n5433 0.152939
R18118 gnd.n5435 gnd.n5434 0.152939
R18119 gnd.n5436 gnd.n5435 0.152939
R18120 gnd.n5437 gnd.n5436 0.152939
R18121 gnd.n5438 gnd.n5437 0.152939
R18122 gnd.n5438 gnd.n1596 0.152939
R18123 gnd.n5961 gnd.n1596 0.152939
R18124 gnd.n2089 gnd.n2010 0.152939
R18125 gnd.n2090 gnd.n2089 0.152939
R18126 gnd.n2091 gnd.n2090 0.152939
R18127 gnd.n2091 gnd.n2081 0.152939
R18128 gnd.n2099 gnd.n2081 0.152939
R18129 gnd.n2100 gnd.n2099 0.152939
R18130 gnd.n2101 gnd.n2100 0.152939
R18131 gnd.n2101 gnd.n2077 0.152939
R18132 gnd.n2109 gnd.n2077 0.152939
R18133 gnd.n2110 gnd.n2109 0.152939
R18134 gnd.n2111 gnd.n2110 0.152939
R18135 gnd.n2111 gnd.n2073 0.152939
R18136 gnd.n2119 gnd.n2073 0.152939
R18137 gnd.n2120 gnd.n2119 0.152939
R18138 gnd.n2121 gnd.n2120 0.152939
R18139 gnd.n2121 gnd.n2069 0.152939
R18140 gnd.n2132 gnd.n2069 0.152939
R18141 gnd.n2133 gnd.n2132 0.152939
R18142 gnd.n2134 gnd.n2133 0.152939
R18143 gnd.n2134 gnd.n2065 0.152939
R18144 gnd.n2142 gnd.n2065 0.152939
R18145 gnd.n2143 gnd.n2142 0.152939
R18146 gnd.n2144 gnd.n2143 0.152939
R18147 gnd.n2144 gnd.n2061 0.152939
R18148 gnd.n2152 gnd.n2061 0.152939
R18149 gnd.n2153 gnd.n2152 0.152939
R18150 gnd.n2154 gnd.n2153 0.152939
R18151 gnd.n2154 gnd.n2057 0.152939
R18152 gnd.n2162 gnd.n2057 0.152939
R18153 gnd.n2163 gnd.n2162 0.152939
R18154 gnd.n2165 gnd.n2163 0.152939
R18155 gnd.n2165 gnd.n2164 0.152939
R18156 gnd.n2164 gnd.n2050 0.152939
R18157 gnd.n2174 gnd.n2050 0.152939
R18158 gnd.n5285 gnd.n5284 0.152939
R18159 gnd.n5286 gnd.n5285 0.152939
R18160 gnd.n5286 gnd.n1993 0.152939
R18161 gnd.n5300 gnd.n1993 0.152939
R18162 gnd.n5301 gnd.n5300 0.152939
R18163 gnd.n5302 gnd.n5301 0.152939
R18164 gnd.n5302 gnd.n1975 0.152939
R18165 gnd.n5316 gnd.n1975 0.152939
R18166 gnd.n5317 gnd.n5316 0.152939
R18167 gnd.n5318 gnd.n5317 0.152939
R18168 gnd.n5318 gnd.n1957 0.152939
R18169 gnd.n5341 gnd.n1957 0.152939
R18170 gnd.n5342 gnd.n5341 0.152939
R18171 gnd.n5343 gnd.n5342 0.152939
R18172 gnd.n5344 gnd.n5343 0.152939
R18173 gnd.n5344 gnd.n1917 0.152939
R18174 gnd.n5382 gnd.n1917 0.152939
R18175 gnd.n5383 gnd.n5382 0.152939
R18176 gnd.n5384 gnd.n5383 0.152939
R18177 gnd.n5384 gnd.n1838 0.152939
R18178 gnd.n5648 gnd.n1838 0.152939
R18179 gnd.n5172 gnd.n2221 0.152939
R18180 gnd.n5173 gnd.n5172 0.152939
R18181 gnd.n5174 gnd.n5173 0.152939
R18182 gnd.n5175 gnd.n5174 0.152939
R18183 gnd.n5176 gnd.n5175 0.152939
R18184 gnd.n5179 gnd.n5176 0.152939
R18185 gnd.n5180 gnd.n5179 0.152939
R18186 gnd.n5181 gnd.n5180 0.152939
R18187 gnd.n5182 gnd.n5181 0.152939
R18188 gnd.n5185 gnd.n5182 0.152939
R18189 gnd.n5186 gnd.n5185 0.152939
R18190 gnd.n5187 gnd.n5186 0.152939
R18191 gnd.n5188 gnd.n5187 0.152939
R18192 gnd.n5189 gnd.n5188 0.152939
R18193 gnd.n3379 gnd.n3378 0.152939
R18194 gnd.n3380 gnd.n3379 0.152939
R18195 gnd.n3380 gnd.n2315 0.152939
R18196 gnd.n3388 gnd.n2315 0.152939
R18197 gnd.n3389 gnd.n3388 0.152939
R18198 gnd.n3390 gnd.n3389 0.152939
R18199 gnd.n3390 gnd.n2309 0.152939
R18200 gnd.n3398 gnd.n2309 0.152939
R18201 gnd.n3399 gnd.n3398 0.152939
R18202 gnd.n3400 gnd.n3399 0.152939
R18203 gnd.n3400 gnd.n2303 0.152939
R18204 gnd.n3408 gnd.n2303 0.152939
R18205 gnd.n3409 gnd.n3408 0.152939
R18206 gnd.n3410 gnd.n3409 0.152939
R18207 gnd.n3410 gnd.n2297 0.152939
R18208 gnd.n3418 gnd.n2297 0.152939
R18209 gnd.n3419 gnd.n3418 0.152939
R18210 gnd.n3420 gnd.n3419 0.152939
R18211 gnd.n3420 gnd.n2291 0.152939
R18212 gnd.n3428 gnd.n2291 0.152939
R18213 gnd.n3429 gnd.n3428 0.152939
R18214 gnd.n3430 gnd.n3429 0.152939
R18215 gnd.n3430 gnd.n2285 0.152939
R18216 gnd.n3438 gnd.n2285 0.152939
R18217 gnd.n3439 gnd.n3438 0.152939
R18218 gnd.n3440 gnd.n3439 0.152939
R18219 gnd.n3440 gnd.n2279 0.152939
R18220 gnd.n3448 gnd.n2279 0.152939
R18221 gnd.n3449 gnd.n3448 0.152939
R18222 gnd.n3450 gnd.n3449 0.152939
R18223 gnd.n3450 gnd.n2273 0.152939
R18224 gnd.n3458 gnd.n2273 0.152939
R18225 gnd.n3459 gnd.n3458 0.152939
R18226 gnd.n3460 gnd.n3459 0.152939
R18227 gnd.n3460 gnd.n2267 0.152939
R18228 gnd.n3468 gnd.n2267 0.152939
R18229 gnd.n3469 gnd.n3468 0.152939
R18230 gnd.n3470 gnd.n3469 0.152939
R18231 gnd.n3470 gnd.n2261 0.152939
R18232 gnd.n3478 gnd.n2261 0.152939
R18233 gnd.n3479 gnd.n3478 0.152939
R18234 gnd.n3480 gnd.n3479 0.152939
R18235 gnd.n3480 gnd.n2255 0.152939
R18236 gnd.n3488 gnd.n2255 0.152939
R18237 gnd.n3489 gnd.n3488 0.152939
R18238 gnd.n3490 gnd.n3489 0.152939
R18239 gnd.n3490 gnd.n2249 0.152939
R18240 gnd.n3498 gnd.n2249 0.152939
R18241 gnd.n3499 gnd.n3498 0.152939
R18242 gnd.n3500 gnd.n3499 0.152939
R18243 gnd.n3500 gnd.n2243 0.152939
R18244 gnd.n3508 gnd.n2243 0.152939
R18245 gnd.n3509 gnd.n3508 0.152939
R18246 gnd.n3510 gnd.n3509 0.152939
R18247 gnd.n3510 gnd.n2237 0.152939
R18248 gnd.n3518 gnd.n2237 0.152939
R18249 gnd.n3519 gnd.n3518 0.152939
R18250 gnd.n3520 gnd.n3519 0.152939
R18251 gnd.n3520 gnd.n2231 0.152939
R18252 gnd.n3528 gnd.n2231 0.152939
R18253 gnd.n3529 gnd.n3528 0.152939
R18254 gnd.n3530 gnd.n3529 0.152939
R18255 gnd.n3530 gnd.n2225 0.152939
R18256 gnd.n5164 gnd.n2225 0.152939
R18257 gnd.n5165 gnd.n5164 0.152939
R18258 gnd.n5166 gnd.n5165 0.152939
R18259 gnd.n1020 gnd.n1019 0.152939
R18260 gnd.n1020 gnd.n1001 0.152939
R18261 gnd.n1026 gnd.n1001 0.152939
R18262 gnd.n1027 gnd.n1026 0.152939
R18263 gnd.n1028 gnd.n1027 0.152939
R18264 gnd.n1028 gnd.n995 0.152939
R18265 gnd.n1035 gnd.n995 0.152939
R18266 gnd.n1036 gnd.n1035 0.152939
R18267 gnd.n6708 gnd.n1036 0.152939
R18268 gnd.n5823 gnd.n5822 0.152939
R18269 gnd.n5824 gnd.n5823 0.152939
R18270 gnd.n5824 gnd.n1653 0.152939
R18271 gnd.n5842 gnd.n1653 0.152939
R18272 gnd.n5843 gnd.n5842 0.152939
R18273 gnd.n5844 gnd.n5843 0.152939
R18274 gnd.n5844 gnd.n1639 0.152939
R18275 gnd.n5864 gnd.n1639 0.152939
R18276 gnd.n5865 gnd.n5864 0.152939
R18277 gnd.n5871 gnd.n5865 0.152939
R18278 gnd.n5871 gnd.n5870 0.152939
R18279 gnd.n5870 gnd.n5869 0.152939
R18280 gnd.n5869 gnd.n5866 0.152939
R18281 gnd.n5866 gnd.n1412 0.152939
R18282 gnd.n6084 gnd.n1412 0.152939
R18283 gnd.n6085 gnd.n6084 0.152939
R18284 gnd.n6120 gnd.n6085 0.152939
R18285 gnd.n6120 gnd.n6119 0.152939
R18286 gnd.n6119 gnd.n6118 0.152939
R18287 gnd.n6118 gnd.n6086 0.152939
R18288 gnd.n6114 gnd.n6086 0.152939
R18289 gnd.n6114 gnd.n6113 0.152939
R18290 gnd.n6113 gnd.n6112 0.152939
R18291 gnd.n6112 gnd.n6090 0.152939
R18292 gnd.n6108 gnd.n6090 0.152939
R18293 gnd.n6108 gnd.n1335 0.152939
R18294 gnd.n6231 gnd.n1335 0.152939
R18295 gnd.n6232 gnd.n6231 0.152939
R18296 gnd.n6246 gnd.n6232 0.152939
R18297 gnd.n6246 gnd.n6245 0.152939
R18298 gnd.n6245 gnd.n6244 0.152939
R18299 gnd.n6244 gnd.n6233 0.152939
R18300 gnd.n6240 gnd.n6233 0.152939
R18301 gnd.n6240 gnd.n6239 0.152939
R18302 gnd.n6239 gnd.n6238 0.152939
R18303 gnd.n6238 gnd.n1276 0.152939
R18304 gnd.n6344 gnd.n1276 0.152939
R18305 gnd.n6345 gnd.n6344 0.152939
R18306 gnd.n6379 gnd.n6345 0.152939
R18307 gnd.n6379 gnd.n6378 0.152939
R18308 gnd.n6378 gnd.n6377 0.152939
R18309 gnd.n6377 gnd.n6346 0.152939
R18310 gnd.n6373 gnd.n6346 0.152939
R18311 gnd.n6373 gnd.n6372 0.152939
R18312 gnd.n6372 gnd.n6371 0.152939
R18313 gnd.n6371 gnd.n6349 0.152939
R18314 gnd.n6367 gnd.n6349 0.152939
R18315 gnd.n6367 gnd.n6366 0.152939
R18316 gnd.n6366 gnd.n6365 0.152939
R18317 gnd.n6365 gnd.n6353 0.152939
R18318 gnd.n6361 gnd.n6353 0.152939
R18319 gnd.n6361 gnd.n6360 0.152939
R18320 gnd.n6360 gnd.n1087 0.152939
R18321 gnd.n6634 gnd.n1087 0.152939
R18322 gnd.n6635 gnd.n6634 0.152939
R18323 gnd.n6637 gnd.n6635 0.152939
R18324 gnd.n6637 gnd.n6636 0.152939
R18325 gnd.n6636 gnd.n1062 0.152939
R18326 gnd.n6664 gnd.n1062 0.152939
R18327 gnd.n6665 gnd.n6664 0.152939
R18328 gnd.n6668 gnd.n6665 0.152939
R18329 gnd.n6668 gnd.n6667 0.152939
R18330 gnd.n6667 gnd.n6666 0.152939
R18331 gnd.n6666 gnd.n1037 0.152939
R18332 gnd.n6707 gnd.n1037 0.152939
R18333 gnd.n5761 gnd.n5760 0.152939
R18334 gnd.n5760 gnd.n5759 0.152939
R18335 gnd.n5759 gnd.n5734 0.152939
R18336 gnd.n5755 gnd.n5734 0.152939
R18337 gnd.n5755 gnd.n5754 0.152939
R18338 gnd.n5754 gnd.n5753 0.152939
R18339 gnd.n5753 gnd.n5740 0.152939
R18340 gnd.n5749 gnd.n5740 0.152939
R18341 gnd.n5749 gnd.n1666 0.152939
R18342 gnd.n5411 gnd.n1896 0.152939
R18343 gnd.n5417 gnd.n1896 0.152939
R18344 gnd.n5418 gnd.n5417 0.152939
R18345 gnd.n5593 gnd.n5418 0.152939
R18346 gnd.n5593 gnd.n5592 0.152939
R18347 gnd.n5592 gnd.n5591 0.152939
R18348 gnd.n5591 gnd.n5419 0.152939
R18349 gnd.n5587 gnd.n5419 0.152939
R18350 gnd.n5587 gnd.n5586 0.152939
R18351 gnd.n5586 gnd.n5585 0.152939
R18352 gnd.n5585 gnd.n5423 0.152939
R18353 gnd.n5581 gnd.n5423 0.152939
R18354 gnd.n5581 gnd.n5580 0.152939
R18355 gnd.n5580 gnd.n5579 0.152939
R18356 gnd.n5579 gnd.n5427 0.152939
R18357 gnd.n5575 gnd.n5427 0.152939
R18358 gnd.n5575 gnd.n5574 0.152939
R18359 gnd.n5574 gnd.n5573 0.152939
R18360 gnd.n5573 gnd.n5431 0.152939
R18361 gnd.n5431 gnd.n1756 0.152939
R18362 gnd.n5724 gnd.n1756 0.152939
R18363 gnd.n5725 gnd.n5724 0.152939
R18364 gnd.n5726 gnd.n5725 0.152939
R18365 gnd.n5726 gnd.n1754 0.152939
R18366 gnd.n5732 gnd.n1754 0.152939
R18367 gnd.n5896 gnd.n1621 0.152939
R18368 gnd.n5892 gnd.n1621 0.152939
R18369 gnd.n5892 gnd.n5891 0.152939
R18370 gnd.n5891 gnd.n5890 0.152939
R18371 gnd.n5890 gnd.n1626 0.152939
R18372 gnd.n5886 gnd.n1626 0.152939
R18373 gnd.n5886 gnd.n5885 0.152939
R18374 gnd.n5885 gnd.n5884 0.152939
R18375 gnd.n5884 gnd.n1631 0.152939
R18376 gnd.n5880 gnd.n1631 0.152939
R18377 gnd.n5880 gnd.n5879 0.152939
R18378 gnd.n5879 gnd.n1420 0.152939
R18379 gnd.n6075 gnd.n1420 0.152939
R18380 gnd.n6076 gnd.n6075 0.152939
R18381 gnd.n6078 gnd.n6076 0.152939
R18382 gnd.n6078 gnd.n6077 0.152939
R18383 gnd.n6077 gnd.n1388 0.152939
R18384 gnd.n6155 gnd.n1388 0.152939
R18385 gnd.n6156 gnd.n6155 0.152939
R18386 gnd.n6158 gnd.n6156 0.152939
R18387 gnd.n6158 gnd.n6157 0.152939
R18388 gnd.n6157 gnd.n1356 0.152939
R18389 gnd.n6206 gnd.n1356 0.152939
R18390 gnd.n6207 gnd.n6206 0.152939
R18391 gnd.n6209 gnd.n6207 0.152939
R18392 gnd.n6209 gnd.n6208 0.152939
R18393 gnd.n6208 gnd.n1320 0.152939
R18394 gnd.n6272 gnd.n1320 0.152939
R18395 gnd.n6273 gnd.n6272 0.152939
R18396 gnd.n6278 gnd.n6273 0.152939
R18397 gnd.n6278 gnd.n6277 0.152939
R18398 gnd.n6277 gnd.n6276 0.152939
R18399 gnd.n6276 gnd.n1282 0.152939
R18400 gnd.n6335 gnd.n1282 0.152939
R18401 gnd.n6336 gnd.n6335 0.152939
R18402 gnd.n6337 gnd.n6336 0.152939
R18403 gnd.n6337 gnd.n1252 0.152939
R18404 gnd.n6404 gnd.n1252 0.152939
R18405 gnd.n6405 gnd.n6404 0.152939
R18406 gnd.n6406 gnd.n6405 0.152939
R18407 gnd.n6406 gnd.n1224 0.152939
R18408 gnd.n6440 gnd.n1224 0.152939
R18409 gnd.n6441 gnd.n6440 0.152939
R18410 gnd.n6442 gnd.n6441 0.152939
R18411 gnd.n6442 gnd.n1196 0.152939
R18412 gnd.n6477 gnd.n1196 0.152939
R18413 gnd.n6478 gnd.n6477 0.152939
R18414 gnd.n6483 gnd.n6478 0.152939
R18415 gnd.n6483 gnd.n6482 0.152939
R18416 gnd.n6482 gnd.n6481 0.152939
R18417 gnd.n6481 gnd.n1096 0.152939
R18418 gnd.n6625 gnd.n1096 0.152939
R18419 gnd.n6626 gnd.n6625 0.152939
R18420 gnd.n6628 gnd.n6626 0.152939
R18421 gnd.n6628 gnd.n6627 0.152939
R18422 gnd.n6627 gnd.n1071 0.152939
R18423 gnd.n6655 gnd.n1071 0.152939
R18424 gnd.n6656 gnd.n6655 0.152939
R18425 gnd.n6658 gnd.n6656 0.152939
R18426 gnd.n6658 gnd.n6657 0.152939
R18427 gnd.n6657 gnd.n1046 0.152939
R18428 gnd.n6697 gnd.n1046 0.152939
R18429 gnd.n6698 gnd.n6697 0.152939
R18430 gnd.n6700 gnd.n6698 0.152939
R18431 gnd.n6700 gnd.n6699 0.152939
R18432 gnd.n7012 gnd.n776 0.152939
R18433 gnd.n7026 gnd.n776 0.152939
R18434 gnd.n7027 gnd.n7026 0.152939
R18435 gnd.n7028 gnd.n7027 0.152939
R18436 gnd.n7028 gnd.n758 0.152939
R18437 gnd.n7042 gnd.n758 0.152939
R18438 gnd.n7043 gnd.n7042 0.152939
R18439 gnd.n7044 gnd.n7043 0.152939
R18440 gnd.n7044 gnd.n740 0.152939
R18441 gnd.n7058 gnd.n740 0.152939
R18442 gnd.n7059 gnd.n7058 0.152939
R18443 gnd.n7060 gnd.n7059 0.152939
R18444 gnd.n7060 gnd.n723 0.152939
R18445 gnd.n7074 gnd.n723 0.152939
R18446 gnd.n7075 gnd.n7074 0.152939
R18447 gnd.n7076 gnd.n7075 0.152939
R18448 gnd.n7076 gnd.n705 0.152939
R18449 gnd.n7091 gnd.n705 0.152939
R18450 gnd.n7092 gnd.n7091 0.152939
R18451 gnd.n7093 gnd.n7092 0.152939
R18452 gnd.n7093 gnd.n688 0.152939
R18453 gnd.n7107 gnd.n688 0.152939
R18454 gnd.n7108 gnd.n7107 0.152939
R18455 gnd.n7109 gnd.n7108 0.152939
R18456 gnd.n7109 gnd.n672 0.152939
R18457 gnd.n7123 gnd.n672 0.152939
R18458 gnd.n7124 gnd.n7123 0.152939
R18459 gnd.n7125 gnd.n7124 0.152939
R18460 gnd.n7125 gnd.n657 0.152939
R18461 gnd.n7138 gnd.n657 0.152939
R18462 gnd.n7139 gnd.n7138 0.152939
R18463 gnd.n7140 gnd.n7139 0.152939
R18464 gnd.n7140 gnd.n640 0.152939
R18465 gnd.n7154 gnd.n640 0.152939
R18466 gnd.n7155 gnd.n7154 0.152939
R18467 gnd.n7156 gnd.n7155 0.152939
R18468 gnd.n7156 gnd.n623 0.152939
R18469 gnd.n7170 gnd.n623 0.152939
R18470 gnd.n7171 gnd.n7170 0.152939
R18471 gnd.n7172 gnd.n7171 0.152939
R18472 gnd.n7172 gnd.n607 0.152939
R18473 gnd.n7186 gnd.n607 0.152939
R18474 gnd.n7187 gnd.n7186 0.152939
R18475 gnd.n7188 gnd.n7187 0.152939
R18476 gnd.n7188 gnd.n590 0.152939
R18477 gnd.n7202 gnd.n590 0.152939
R18478 gnd.n7203 gnd.n7202 0.152939
R18479 gnd.n7272 gnd.n7203 0.152939
R18480 gnd.n7272 gnd.n7271 0.152939
R18481 gnd.n7271 gnd.n7270 0.152939
R18482 gnd.n7270 gnd.n7204 0.152939
R18483 gnd.n7266 gnd.n7204 0.152939
R18484 gnd.n7265 gnd.n7206 0.152939
R18485 gnd.n7261 gnd.n7206 0.152939
R18486 gnd.n7261 gnd.n7260 0.152939
R18487 gnd.n7260 gnd.n7259 0.152939
R18488 gnd.n7259 gnd.n7212 0.152939
R18489 gnd.n7255 gnd.n7212 0.152939
R18490 gnd.n7255 gnd.n7254 0.152939
R18491 gnd.n7254 gnd.n7253 0.152939
R18492 gnd.n7253 gnd.n7220 0.152939
R18493 gnd.n7249 gnd.n7220 0.152939
R18494 gnd.n7249 gnd.n7248 0.152939
R18495 gnd.n7248 gnd.n7247 0.152939
R18496 gnd.n7247 gnd.n7228 0.152939
R18497 gnd.n7243 gnd.n7228 0.152939
R18498 gnd.n7243 gnd.n7242 0.152939
R18499 gnd.n7242 gnd.n7241 0.152939
R18500 gnd.n1017 gnd.n1012 0.152939
R18501 gnd.n1012 gnd.n911 0.152939
R18502 gnd.n6889 gnd.n911 0.152939
R18503 gnd.n6889 gnd.n6888 0.152939
R18504 gnd.n6888 gnd.n6887 0.152939
R18505 gnd.n6887 gnd.n912 0.152939
R18506 gnd.n6883 gnd.n912 0.152939
R18507 gnd.n6883 gnd.n6882 0.152939
R18508 gnd.n6882 gnd.n6881 0.152939
R18509 gnd.n6881 gnd.n916 0.152939
R18510 gnd.n6877 gnd.n916 0.152939
R18511 gnd.n6877 gnd.n6876 0.152939
R18512 gnd.n6876 gnd.n6875 0.152939
R18513 gnd.n6875 gnd.n920 0.152939
R18514 gnd.n6871 gnd.n920 0.152939
R18515 gnd.n6871 gnd.n6870 0.152939
R18516 gnd.n6870 gnd.n6869 0.152939
R18517 gnd.n6869 gnd.n924 0.152939
R18518 gnd.n6865 gnd.n924 0.152939
R18519 gnd.n6865 gnd.n6864 0.152939
R18520 gnd.n6864 gnd.n6863 0.152939
R18521 gnd.n6863 gnd.n928 0.152939
R18522 gnd.n6859 gnd.n928 0.152939
R18523 gnd.n6859 gnd.n6858 0.152939
R18524 gnd.n6858 gnd.n465 0.152939
R18525 gnd.n7394 gnd.n465 0.152939
R18526 gnd.n7394 gnd.n7393 0.152939
R18527 gnd.n7393 gnd.n467 0.152939
R18528 gnd.n7389 gnd.n467 0.152939
R18529 gnd.n7389 gnd.n7388 0.152939
R18530 gnd.n7388 gnd.n7387 0.152939
R18531 gnd.n7387 gnd.n472 0.152939
R18532 gnd.n7383 gnd.n472 0.152939
R18533 gnd.n7383 gnd.n7382 0.152939
R18534 gnd.n7382 gnd.n7381 0.152939
R18535 gnd.n7381 gnd.n477 0.152939
R18536 gnd.n7377 gnd.n477 0.152939
R18537 gnd.n7377 gnd.n7376 0.152939
R18538 gnd.n7376 gnd.n7375 0.152939
R18539 gnd.n7375 gnd.n482 0.152939
R18540 gnd.n7371 gnd.n482 0.152939
R18541 gnd.n7371 gnd.n7370 0.152939
R18542 gnd.n7370 gnd.n7369 0.152939
R18543 gnd.n7369 gnd.n487 0.152939
R18544 gnd.n7365 gnd.n487 0.152939
R18545 gnd.n7365 gnd.n7364 0.152939
R18546 gnd.n7364 gnd.n7363 0.152939
R18547 gnd.n7363 gnd.n492 0.152939
R18548 gnd.n7359 gnd.n492 0.152939
R18549 gnd.n7359 gnd.n7358 0.152939
R18550 gnd.n7358 gnd.n7357 0.152939
R18551 gnd.n7357 gnd.n497 0.152939
R18552 gnd.n4336 gnd.n0 0.148472
R18553 gnd.n6838 gnd.n941 0.146841
R18554 gnd.n5189 gnd.n1839 0.146841
R18555 gnd.n5410 gnd.n5409 0.145814
R18556 gnd.n5411 gnd.n5410 0.145814
R18557 gnd.n1019 gnd.n1018 0.145317
R18558 gnd.n5761 gnd.n5733 0.145317
R18559 gnd.n4337 gnd.n4091 0.0767195
R18560 gnd.n4337 gnd.n4089 0.0767195
R18561 gnd.n5898 gnd.n5897 0.063
R18562 gnd.n7011 gnd.n791 0.063
R18563 gnd.n5085 gnd.n3650 0.0477147
R18564 gnd.n4031 gnd.n3927 0.0442063
R18565 gnd.n4045 gnd.n3927 0.0442063
R18566 gnd.n4046 gnd.n4045 0.0442063
R18567 gnd.n4047 gnd.n4046 0.0442063
R18568 gnd.n4047 gnd.n3915 0.0442063
R18569 gnd.n4061 gnd.n3915 0.0442063
R18570 gnd.n4062 gnd.n4061 0.0442063
R18571 gnd.n4063 gnd.n4062 0.0442063
R18572 gnd.n4063 gnd.n3902 0.0442063
R18573 gnd.n4434 gnd.n3902 0.0442063
R18574 gnd.n4437 gnd.n4436 0.0344674
R18575 gnd.n1011 gnd.n1006 0.0344674
R18576 gnd.n5765 gnd.n1748 0.0344674
R18577 gnd.n3895 gnd.n3894 0.0269946
R18578 gnd.n4447 gnd.n4445 0.0269946
R18579 gnd.n4446 gnd.n3877 0.0269946
R18580 gnd.n4466 gnd.n4465 0.0269946
R18581 gnd.n4468 gnd.n4467 0.0269946
R18582 gnd.n3871 gnd.n3869 0.0269946
R18583 gnd.n4478 gnd.n4476 0.0269946
R18584 gnd.n4477 gnd.n3850 0.0269946
R18585 gnd.n4497 gnd.n4496 0.0269946
R18586 gnd.n4499 gnd.n4498 0.0269946
R18587 gnd.n3845 gnd.n3843 0.0269946
R18588 gnd.n4509 gnd.n4507 0.0269946
R18589 gnd.n4508 gnd.n3824 0.0269946
R18590 gnd.n4528 gnd.n4527 0.0269946
R18591 gnd.n4530 gnd.n4529 0.0269946
R18592 gnd.n3819 gnd.n3817 0.0269946
R18593 gnd.n4540 gnd.n4538 0.0269946
R18594 gnd.n4539 gnd.n3799 0.0269946
R18595 gnd.n4559 gnd.n4558 0.0269946
R18596 gnd.n4561 gnd.n4560 0.0269946
R18597 gnd.n3793 gnd.n3791 0.0269946
R18598 gnd.n4571 gnd.n4569 0.0269946
R18599 gnd.n4570 gnd.n3774 0.0269946
R18600 gnd.n4590 gnd.n4589 0.0269946
R18601 gnd.n4592 gnd.n4591 0.0269946
R18602 gnd.n3768 gnd.n3766 0.0269946
R18603 gnd.n4602 gnd.n4600 0.0269946
R18604 gnd.n4601 gnd.n3749 0.0269946
R18605 gnd.n4621 gnd.n4620 0.0269946
R18606 gnd.n4623 gnd.n4622 0.0269946
R18607 gnd.n3743 gnd.n3742 0.0269946
R18608 gnd.n4633 gnd.n3738 0.0269946
R18609 gnd.n4632 gnd.n3740 0.0269946
R18610 gnd.n3739 gnd.n3721 0.0269946
R18611 gnd.n4653 gnd.n3722 0.0269946
R18612 gnd.n4652 gnd.n3723 0.0269946
R18613 gnd.n4697 gnd.n3698 0.0269946
R18614 gnd.n4699 gnd.n4698 0.0269946
R18615 gnd.n4700 gnd.n3541 0.0269946
R18616 gnd.n3693 gnd.n3542 0.0269946
R18617 gnd.n3695 gnd.n3543 0.0269946
R18618 gnd.n4708 gnd.n4707 0.0269946
R18619 gnd.n4710 gnd.n4709 0.0269946
R18620 gnd.n4711 gnd.n3563 0.0269946
R18621 gnd.n3687 gnd.n3564 0.0269946
R18622 gnd.n3689 gnd.n3565 0.0269946
R18623 gnd.n4744 gnd.n4743 0.0269946
R18624 gnd.n4746 gnd.n4745 0.0269946
R18625 gnd.n5005 gnd.n3589 0.0269946
R18626 gnd.n5007 gnd.n3590 0.0269946
R18627 gnd.n5009 gnd.n5008 0.0269946
R18628 gnd.n5013 gnd.n5012 0.0269946
R18629 gnd.n7008 gnd.n791 0.0246168
R18630 gnd.n5897 gnd.n1620 0.0246168
R18631 gnd.n4436 gnd.n4435 0.0202011
R18632 gnd.n7007 gnd.n794 0.0188424
R18633 gnd.n7004 gnd.n7003 0.0188424
R18634 gnd.n7000 gnd.n798 0.0188424
R18635 gnd.n6999 gnd.n802 0.0188424
R18636 gnd.n6996 gnd.n6995 0.0188424
R18637 gnd.n6992 gnd.n806 0.0188424
R18638 gnd.n6991 gnd.n810 0.0188424
R18639 gnd.n6988 gnd.n6987 0.0188424
R18640 gnd.n6984 gnd.n814 0.0188424
R18641 gnd.n6983 gnd.n818 0.0188424
R18642 gnd.n6980 gnd.n6979 0.0188424
R18643 gnd.n6976 gnd.n822 0.0188424
R18644 gnd.n6975 gnd.n826 0.0188424
R18645 gnd.n6972 gnd.n6971 0.0188424
R18646 gnd.n1005 gnd.n830 0.0188424
R18647 gnd.n1692 gnd.n1690 0.0188424
R18648 gnd.n5804 gnd.n5803 0.0188424
R18649 gnd.n5800 gnd.n1693 0.0188424
R18650 gnd.n5799 gnd.n1704 0.0188424
R18651 gnd.n5796 gnd.n5795 0.0188424
R18652 gnd.n5792 gnd.n1709 0.0188424
R18653 gnd.n5791 gnd.n1715 0.0188424
R18654 gnd.n5788 gnd.n5787 0.0188424
R18655 gnd.n5784 gnd.n1719 0.0188424
R18656 gnd.n5783 gnd.n1726 0.0188424
R18657 gnd.n5780 gnd.n5779 0.0188424
R18658 gnd.n5776 gnd.n1732 0.0188424
R18659 gnd.n5775 gnd.n1738 0.0188424
R18660 gnd.n5772 gnd.n5771 0.0188424
R18661 gnd.n5766 gnd.n1742 0.0188424
R18662 gnd.n7008 gnd.n7007 0.016125
R18663 gnd.n7004 gnd.n794 0.016125
R18664 gnd.n7003 gnd.n798 0.016125
R18665 gnd.n7000 gnd.n6999 0.016125
R18666 gnd.n6996 gnd.n802 0.016125
R18667 gnd.n6995 gnd.n806 0.016125
R18668 gnd.n6992 gnd.n6991 0.016125
R18669 gnd.n6988 gnd.n810 0.016125
R18670 gnd.n6987 gnd.n814 0.016125
R18671 gnd.n6984 gnd.n6983 0.016125
R18672 gnd.n6980 gnd.n818 0.016125
R18673 gnd.n6979 gnd.n822 0.016125
R18674 gnd.n6976 gnd.n6975 0.016125
R18675 gnd.n6972 gnd.n826 0.016125
R18676 gnd.n6971 gnd.n830 0.016125
R18677 gnd.n1006 gnd.n1005 0.016125
R18678 gnd.n1690 gnd.n1620 0.016125
R18679 gnd.n5804 gnd.n1692 0.016125
R18680 gnd.n5803 gnd.n1693 0.016125
R18681 gnd.n5800 gnd.n5799 0.016125
R18682 gnd.n5796 gnd.n1704 0.016125
R18683 gnd.n5795 gnd.n1709 0.016125
R18684 gnd.n5792 gnd.n5791 0.016125
R18685 gnd.n5788 gnd.n1715 0.016125
R18686 gnd.n5787 gnd.n1719 0.016125
R18687 gnd.n5784 gnd.n5783 0.016125
R18688 gnd.n5780 gnd.n1726 0.016125
R18689 gnd.n5779 gnd.n1732 0.016125
R18690 gnd.n5776 gnd.n5775 0.016125
R18691 gnd.n5772 gnd.n1738 0.016125
R18692 gnd.n5771 gnd.n1742 0.016125
R18693 gnd.n5766 gnd.n5765 0.016125
R18694 gnd.n4435 gnd.n4434 0.0148637
R18695 gnd.n5003 gnd.n5002 0.0144266
R18696 gnd.n5002 gnd.n3588 0.0130679
R18697 gnd.n4437 gnd.n3895 0.00797283
R18698 gnd.n4445 gnd.n3894 0.00797283
R18699 gnd.n4447 gnd.n4446 0.00797283
R18700 gnd.n4465 gnd.n3877 0.00797283
R18701 gnd.n4467 gnd.n4466 0.00797283
R18702 gnd.n4468 gnd.n3871 0.00797283
R18703 gnd.n4476 gnd.n3869 0.00797283
R18704 gnd.n4478 gnd.n4477 0.00797283
R18705 gnd.n4496 gnd.n3850 0.00797283
R18706 gnd.n4498 gnd.n4497 0.00797283
R18707 gnd.n4499 gnd.n3845 0.00797283
R18708 gnd.n4507 gnd.n3843 0.00797283
R18709 gnd.n4509 gnd.n4508 0.00797283
R18710 gnd.n4527 gnd.n3824 0.00797283
R18711 gnd.n4529 gnd.n4528 0.00797283
R18712 gnd.n4530 gnd.n3819 0.00797283
R18713 gnd.n4538 gnd.n3817 0.00797283
R18714 gnd.n4540 gnd.n4539 0.00797283
R18715 gnd.n4558 gnd.n3799 0.00797283
R18716 gnd.n4560 gnd.n4559 0.00797283
R18717 gnd.n4561 gnd.n3793 0.00797283
R18718 gnd.n4569 gnd.n3791 0.00797283
R18719 gnd.n4571 gnd.n4570 0.00797283
R18720 gnd.n4589 gnd.n3774 0.00797283
R18721 gnd.n4591 gnd.n4590 0.00797283
R18722 gnd.n4592 gnd.n3768 0.00797283
R18723 gnd.n4600 gnd.n3766 0.00797283
R18724 gnd.n4602 gnd.n4601 0.00797283
R18725 gnd.n4620 gnd.n3749 0.00797283
R18726 gnd.n4622 gnd.n4621 0.00797283
R18727 gnd.n4623 gnd.n3743 0.00797283
R18728 gnd.n3742 gnd.n3738 0.00797283
R18729 gnd.n4633 gnd.n4632 0.00797283
R18730 gnd.n3740 gnd.n3739 0.00797283
R18731 gnd.n3722 gnd.n3721 0.00797283
R18732 gnd.n4653 gnd.n4652 0.00797283
R18733 gnd.n3723 gnd.n3698 0.00797283
R18734 gnd.n4698 gnd.n4697 0.00797283
R18735 gnd.n4700 gnd.n4699 0.00797283
R18736 gnd.n3693 gnd.n3541 0.00797283
R18737 gnd.n3695 gnd.n3542 0.00797283
R18738 gnd.n4707 gnd.n3543 0.00797283
R18739 gnd.n4709 gnd.n4708 0.00797283
R18740 gnd.n4711 gnd.n4710 0.00797283
R18741 gnd.n3687 gnd.n3563 0.00797283
R18742 gnd.n3689 gnd.n3564 0.00797283
R18743 gnd.n4743 gnd.n3565 0.00797283
R18744 gnd.n4745 gnd.n4744 0.00797283
R18745 gnd.n5003 gnd.n4746 0.00797283
R18746 gnd.n5005 gnd.n3588 0.00797283
R18747 gnd.n5007 gnd.n3589 0.00797283
R18748 gnd.n5008 gnd.n3590 0.00797283
R18749 gnd.n5013 gnd.n5009 0.00797283
R18750 gnd.n5012 gnd.n3650 0.00797283
R18751 gnd.n5464 gnd.n1839 0.00659756
R18752 gnd.n6838 gnd.n6837 0.00659756
R18753 gnd.n7123 gnd.n671 0.0051789
R18754 gnd.n5607 gnd.n5606 0.0051789
R18755 gnd.n1018 gnd.n1011 0.00219837
R18756 gnd.n5733 gnd.n1748 0.00219837
R18757 CSoutput.n19 CSoutput.t94 184.661
R18758 CSoutput.n78 CSoutput.n77 165.8
R18759 CSoutput.n76 CSoutput.n0 165.8
R18760 CSoutput.n75 CSoutput.n74 165.8
R18761 CSoutput.n73 CSoutput.n72 165.8
R18762 CSoutput.n71 CSoutput.n2 165.8
R18763 CSoutput.n69 CSoutput.n68 165.8
R18764 CSoutput.n67 CSoutput.n3 165.8
R18765 CSoutput.n66 CSoutput.n65 165.8
R18766 CSoutput.n63 CSoutput.n4 165.8
R18767 CSoutput.n61 CSoutput.n60 165.8
R18768 CSoutput.n59 CSoutput.n5 165.8
R18769 CSoutput.n58 CSoutput.n57 165.8
R18770 CSoutput.n55 CSoutput.n6 165.8
R18771 CSoutput.n54 CSoutput.n53 165.8
R18772 CSoutput.n52 CSoutput.n51 165.8
R18773 CSoutput.n50 CSoutput.n8 165.8
R18774 CSoutput.n48 CSoutput.n47 165.8
R18775 CSoutput.n46 CSoutput.n9 165.8
R18776 CSoutput.n45 CSoutput.n44 165.8
R18777 CSoutput.n42 CSoutput.n10 165.8
R18778 CSoutput.n41 CSoutput.n40 165.8
R18779 CSoutput.n39 CSoutput.n38 165.8
R18780 CSoutput.n37 CSoutput.n12 165.8
R18781 CSoutput.n35 CSoutput.n34 165.8
R18782 CSoutput.n33 CSoutput.n13 165.8
R18783 CSoutput.n32 CSoutput.n31 165.8
R18784 CSoutput.n29 CSoutput.n14 165.8
R18785 CSoutput.n28 CSoutput.n27 165.8
R18786 CSoutput.n26 CSoutput.n25 165.8
R18787 CSoutput.n24 CSoutput.n16 165.8
R18788 CSoutput.n22 CSoutput.n21 165.8
R18789 CSoutput.n20 CSoutput.n17 165.8
R18790 CSoutput.n77 CSoutput.t95 162.194
R18791 CSoutput.n18 CSoutput.t111 120.501
R18792 CSoutput.n23 CSoutput.t105 120.501
R18793 CSoutput.n15 CSoutput.t101 120.501
R18794 CSoutput.n30 CSoutput.t96 120.501
R18795 CSoutput.n36 CSoutput.t108 120.501
R18796 CSoutput.n11 CSoutput.t102 120.501
R18797 CSoutput.n43 CSoutput.t103 120.501
R18798 CSoutput.n49 CSoutput.t112 120.501
R18799 CSoutput.n7 CSoutput.t113 120.501
R18800 CSoutput.n56 CSoutput.t107 120.501
R18801 CSoutput.n62 CSoutput.t100 120.501
R18802 CSoutput.n64 CSoutput.t92 120.501
R18803 CSoutput.n70 CSoutput.t110 120.501
R18804 CSoutput.n1 CSoutput.t104 120.501
R18805 CSoutput.n280 CSoutput.n278 102.66
R18806 CSoutput.n270 CSoutput.n268 102.66
R18807 CSoutput.n261 CSoutput.n259 102.66
R18808 CSoutput.n100 CSoutput.n98 102.66
R18809 CSoutput.n90 CSoutput.n88 102.66
R18810 CSoutput.n81 CSoutput.n79 102.66
R18811 CSoutput.n284 CSoutput.n283 102.088
R18812 CSoutput.n282 CSoutput.n281 102.088
R18813 CSoutput.n280 CSoutput.n279 102.088
R18814 CSoutput.n276 CSoutput.n275 102.088
R18815 CSoutput.n274 CSoutput.n273 102.088
R18816 CSoutput.n272 CSoutput.n271 102.088
R18817 CSoutput.n270 CSoutput.n269 102.088
R18818 CSoutput.n267 CSoutput.n266 102.088
R18819 CSoutput.n265 CSoutput.n264 102.088
R18820 CSoutput.n263 CSoutput.n262 102.088
R18821 CSoutput.n261 CSoutput.n260 102.088
R18822 CSoutput.n100 CSoutput.n99 102.088
R18823 CSoutput.n102 CSoutput.n101 102.088
R18824 CSoutput.n104 CSoutput.n103 102.088
R18825 CSoutput.n106 CSoutput.n105 102.088
R18826 CSoutput.n90 CSoutput.n89 102.088
R18827 CSoutput.n92 CSoutput.n91 102.088
R18828 CSoutput.n94 CSoutput.n93 102.088
R18829 CSoutput.n96 CSoutput.n95 102.088
R18830 CSoutput.n81 CSoutput.n80 102.088
R18831 CSoutput.n83 CSoutput.n82 102.088
R18832 CSoutput.n85 CSoutput.n84 102.088
R18833 CSoutput.n87 CSoutput.n86 102.088
R18834 CSoutput.n286 CSoutput.n285 102.088
R18835 CSoutput.n298 CSoutput.n296 85.0679
R18836 CSoutput.n291 CSoutput.n289 85.0679
R18837 CSoutput.n314 CSoutput.n312 85.0679
R18838 CSoutput.n307 CSoutput.n305 85.0679
R18839 CSoutput.n302 CSoutput.n301 84.0635
R18840 CSoutput.n300 CSoutput.n299 84.0635
R18841 CSoutput.n298 CSoutput.n297 84.0635
R18842 CSoutput.n295 CSoutput.n294 84.0635
R18843 CSoutput.n293 CSoutput.n292 84.0635
R18844 CSoutput.n291 CSoutput.n290 84.0635
R18845 CSoutput.n314 CSoutput.n313 84.0635
R18846 CSoutput.n316 CSoutput.n315 84.0635
R18847 CSoutput.n318 CSoutput.n317 84.0635
R18848 CSoutput.n307 CSoutput.n306 84.0635
R18849 CSoutput.n309 CSoutput.n308 84.0635
R18850 CSoutput.n311 CSoutput.n310 84.0635
R18851 CSoutput.n25 CSoutput.n24 48.1486
R18852 CSoutput.n69 CSoutput.n3 48.1486
R18853 CSoutput.n38 CSoutput.n37 48.1486
R18854 CSoutput.n42 CSoutput.n41 48.1486
R18855 CSoutput.n51 CSoutput.n50 48.1486
R18856 CSoutput.n55 CSoutput.n54 48.1486
R18857 CSoutput.n22 CSoutput.n17 46.462
R18858 CSoutput.n72 CSoutput.n71 46.462
R18859 CSoutput.n20 CSoutput.n19 44.9055
R18860 CSoutput.n29 CSoutput.n28 43.7635
R18861 CSoutput.n65 CSoutput.n63 43.7635
R18862 CSoutput.n35 CSoutput.n13 41.7396
R18863 CSoutput.n57 CSoutput.n5 41.7396
R18864 CSoutput.n44 CSoutput.n9 37.0171
R18865 CSoutput.n48 CSoutput.n9 37.0171
R18866 CSoutput.n76 CSoutput.n75 34.9932
R18867 CSoutput.n31 CSoutput.n13 32.2947
R18868 CSoutput.n61 CSoutput.n5 32.2947
R18869 CSoutput.n30 CSoutput.n29 29.6014
R18870 CSoutput.n63 CSoutput.n62 29.6014
R18871 CSoutput.n19 CSoutput.n18 28.4085
R18872 CSoutput.n18 CSoutput.n17 25.1176
R18873 CSoutput.n72 CSoutput.n1 25.1176
R18874 CSoutput.n43 CSoutput.n42 22.0922
R18875 CSoutput.n50 CSoutput.n49 22.0922
R18876 CSoutput.n77 CSoutput.n76 21.8586
R18877 CSoutput.n37 CSoutput.n36 18.9681
R18878 CSoutput.n56 CSoutput.n55 18.9681
R18879 CSoutput.n25 CSoutput.n15 17.6292
R18880 CSoutput.n64 CSoutput.n3 17.6292
R18881 CSoutput.n24 CSoutput.n23 15.844
R18882 CSoutput.n70 CSoutput.n69 15.844
R18883 CSoutput.n38 CSoutput.n11 14.5051
R18884 CSoutput.n54 CSoutput.n7 14.5051
R18885 CSoutput.n321 CSoutput.n78 11.6139
R18886 CSoutput.n41 CSoutput.n11 11.3811
R18887 CSoutput.n51 CSoutput.n7 11.3811
R18888 CSoutput.n23 CSoutput.n22 10.0422
R18889 CSoutput.n71 CSoutput.n70 10.0422
R18890 CSoutput.n277 CSoutput.n267 8.98182
R18891 CSoutput.n97 CSoutput.n87 8.98182
R18892 CSoutput.n303 CSoutput.n295 8.81666
R18893 CSoutput.n319 CSoutput.n311 8.81666
R18894 CSoutput.n304 CSoutput.n288 8.44388
R18895 CSoutput.n28 CSoutput.n15 8.25698
R18896 CSoutput.n65 CSoutput.n64 8.25698
R18897 CSoutput.n304 CSoutput.n303 7.89345
R18898 CSoutput.n320 CSoutput.n319 7.89345
R18899 CSoutput.n36 CSoutput.n35 6.91809
R18900 CSoutput.n57 CSoutput.n56 6.91809
R18901 CSoutput.n288 CSoutput.n287 5.99005
R18902 CSoutput.n108 CSoutput.n107 5.99005
R18903 CSoutput.n303 CSoutput.n302 5.46817
R18904 CSoutput.n319 CSoutput.n318 5.46817
R18905 CSoutput.n287 CSoutput.n286 5.25266
R18906 CSoutput.n277 CSoutput.n276 5.25266
R18907 CSoutput.n107 CSoutput.n106 5.25266
R18908 CSoutput.n97 CSoutput.n96 5.25266
R18909 CSoutput.n321 CSoutput.n108 4.82011
R18910 CSoutput.n285 CSoutput.t9 4.64407
R18911 CSoutput.n285 CSoutput.t22 4.64407
R18912 CSoutput.n283 CSoutput.t6 4.64407
R18913 CSoutput.n283 CSoutput.t38 4.64407
R18914 CSoutput.n281 CSoutput.t28 4.64407
R18915 CSoutput.n281 CSoutput.t0 4.64407
R18916 CSoutput.n279 CSoutput.t31 4.64407
R18917 CSoutput.n279 CSoutput.t72 4.64407
R18918 CSoutput.n278 CSoutput.t10 4.64407
R18919 CSoutput.n278 CSoutput.t2 4.64407
R18920 CSoutput.n275 CSoutput.t89 4.64407
R18921 CSoutput.n275 CSoutput.t78 4.64407
R18922 CSoutput.n273 CSoutput.t5 4.64407
R18923 CSoutput.n273 CSoutput.t3 4.64407
R18924 CSoutput.n271 CSoutput.t79 4.64407
R18925 CSoutput.n271 CSoutput.t87 4.64407
R18926 CSoutput.n269 CSoutput.t8 4.64407
R18927 CSoutput.n269 CSoutput.t83 4.64407
R18928 CSoutput.n268 CSoutput.t33 4.64407
R18929 CSoutput.n268 CSoutput.t25 4.64407
R18930 CSoutput.n266 CSoutput.t88 4.64407
R18931 CSoutput.n266 CSoutput.t35 4.64407
R18932 CSoutput.n264 CSoutput.t26 4.64407
R18933 CSoutput.n264 CSoutput.t1 4.64407
R18934 CSoutput.n262 CSoutput.t32 4.64407
R18935 CSoutput.n262 CSoutput.t23 4.64407
R18936 CSoutput.n260 CSoutput.t90 4.64407
R18937 CSoutput.n260 CSoutput.t36 4.64407
R18938 CSoutput.n259 CSoutput.t84 4.64407
R18939 CSoutput.n259 CSoutput.t30 4.64407
R18940 CSoutput.n98 CSoutput.t85 4.64407
R18941 CSoutput.n98 CSoutput.t34 4.64407
R18942 CSoutput.n99 CSoutput.t76 4.64407
R18943 CSoutput.n99 CSoutput.t74 4.64407
R18944 CSoutput.n101 CSoutput.t11 4.64407
R18945 CSoutput.n101 CSoutput.t24 4.64407
R18946 CSoutput.n103 CSoutput.t18 4.64407
R18947 CSoutput.n103 CSoutput.t77 4.64407
R18948 CSoutput.n105 CSoutput.t4 4.64407
R18949 CSoutput.n105 CSoutput.t86 4.64407
R18950 CSoutput.n88 CSoutput.t15 4.64407
R18951 CSoutput.n88 CSoutput.t82 4.64407
R18952 CSoutput.n89 CSoutput.t21 4.64407
R18953 CSoutput.n89 CSoutput.t73 4.64407
R18954 CSoutput.n91 CSoutput.t37 4.64407
R18955 CSoutput.n91 CSoutput.t17 4.64407
R18956 CSoutput.n93 CSoutput.t91 4.64407
R18957 CSoutput.n93 CSoutput.t14 4.64407
R18958 CSoutput.n95 CSoutput.t27 4.64407
R18959 CSoutput.n95 CSoutput.t75 4.64407
R18960 CSoutput.n79 CSoutput.t80 4.64407
R18961 CSoutput.n79 CSoutput.t16 4.64407
R18962 CSoutput.n80 CSoutput.t39 4.64407
R18963 CSoutput.n80 CSoutput.t12 4.64407
R18964 CSoutput.n82 CSoutput.t7 4.64407
R18965 CSoutput.n82 CSoutput.t29 4.64407
R18966 CSoutput.n84 CSoutput.t19 4.64407
R18967 CSoutput.n84 CSoutput.t20 4.64407
R18968 CSoutput.n86 CSoutput.t13 4.64407
R18969 CSoutput.n86 CSoutput.t81 4.64407
R18970 CSoutput.n199 CSoutput.n152 4.5005
R18971 CSoutput.n168 CSoutput.n152 4.5005
R18972 CSoutput.n163 CSoutput.n147 4.5005
R18973 CSoutput.n163 CSoutput.n149 4.5005
R18974 CSoutput.n163 CSoutput.n146 4.5005
R18975 CSoutput.n163 CSoutput.n150 4.5005
R18976 CSoutput.n163 CSoutput.n145 4.5005
R18977 CSoutput.n163 CSoutput.t109 4.5005
R18978 CSoutput.n163 CSoutput.n144 4.5005
R18979 CSoutput.n163 CSoutput.n151 4.5005
R18980 CSoutput.n163 CSoutput.n152 4.5005
R18981 CSoutput.n161 CSoutput.n147 4.5005
R18982 CSoutput.n161 CSoutput.n149 4.5005
R18983 CSoutput.n161 CSoutput.n146 4.5005
R18984 CSoutput.n161 CSoutput.n150 4.5005
R18985 CSoutput.n161 CSoutput.n145 4.5005
R18986 CSoutput.n161 CSoutput.t109 4.5005
R18987 CSoutput.n161 CSoutput.n144 4.5005
R18988 CSoutput.n161 CSoutput.n151 4.5005
R18989 CSoutput.n161 CSoutput.n152 4.5005
R18990 CSoutput.n160 CSoutput.n147 4.5005
R18991 CSoutput.n160 CSoutput.n149 4.5005
R18992 CSoutput.n160 CSoutput.n146 4.5005
R18993 CSoutput.n160 CSoutput.n150 4.5005
R18994 CSoutput.n160 CSoutput.n145 4.5005
R18995 CSoutput.n160 CSoutput.t109 4.5005
R18996 CSoutput.n160 CSoutput.n144 4.5005
R18997 CSoutput.n160 CSoutput.n151 4.5005
R18998 CSoutput.n160 CSoutput.n152 4.5005
R18999 CSoutput.n245 CSoutput.n147 4.5005
R19000 CSoutput.n245 CSoutput.n149 4.5005
R19001 CSoutput.n245 CSoutput.n146 4.5005
R19002 CSoutput.n245 CSoutput.n150 4.5005
R19003 CSoutput.n245 CSoutput.n145 4.5005
R19004 CSoutput.n245 CSoutput.t109 4.5005
R19005 CSoutput.n245 CSoutput.n144 4.5005
R19006 CSoutput.n245 CSoutput.n151 4.5005
R19007 CSoutput.n245 CSoutput.n152 4.5005
R19008 CSoutput.n243 CSoutput.n147 4.5005
R19009 CSoutput.n243 CSoutput.n149 4.5005
R19010 CSoutput.n243 CSoutput.n146 4.5005
R19011 CSoutput.n243 CSoutput.n150 4.5005
R19012 CSoutput.n243 CSoutput.n145 4.5005
R19013 CSoutput.n243 CSoutput.t109 4.5005
R19014 CSoutput.n243 CSoutput.n144 4.5005
R19015 CSoutput.n243 CSoutput.n151 4.5005
R19016 CSoutput.n241 CSoutput.n147 4.5005
R19017 CSoutput.n241 CSoutput.n149 4.5005
R19018 CSoutput.n241 CSoutput.n146 4.5005
R19019 CSoutput.n241 CSoutput.n150 4.5005
R19020 CSoutput.n241 CSoutput.n145 4.5005
R19021 CSoutput.n241 CSoutput.t109 4.5005
R19022 CSoutput.n241 CSoutput.n144 4.5005
R19023 CSoutput.n241 CSoutput.n151 4.5005
R19024 CSoutput.n171 CSoutput.n147 4.5005
R19025 CSoutput.n171 CSoutput.n149 4.5005
R19026 CSoutput.n171 CSoutput.n146 4.5005
R19027 CSoutput.n171 CSoutput.n150 4.5005
R19028 CSoutput.n171 CSoutput.n145 4.5005
R19029 CSoutput.n171 CSoutput.t109 4.5005
R19030 CSoutput.n171 CSoutput.n144 4.5005
R19031 CSoutput.n171 CSoutput.n151 4.5005
R19032 CSoutput.n171 CSoutput.n152 4.5005
R19033 CSoutput.n170 CSoutput.n147 4.5005
R19034 CSoutput.n170 CSoutput.n149 4.5005
R19035 CSoutput.n170 CSoutput.n146 4.5005
R19036 CSoutput.n170 CSoutput.n150 4.5005
R19037 CSoutput.n170 CSoutput.n145 4.5005
R19038 CSoutput.n170 CSoutput.t109 4.5005
R19039 CSoutput.n170 CSoutput.n144 4.5005
R19040 CSoutput.n170 CSoutput.n151 4.5005
R19041 CSoutput.n170 CSoutput.n152 4.5005
R19042 CSoutput.n174 CSoutput.n147 4.5005
R19043 CSoutput.n174 CSoutput.n149 4.5005
R19044 CSoutput.n174 CSoutput.n146 4.5005
R19045 CSoutput.n174 CSoutput.n150 4.5005
R19046 CSoutput.n174 CSoutput.n145 4.5005
R19047 CSoutput.n174 CSoutput.t109 4.5005
R19048 CSoutput.n174 CSoutput.n144 4.5005
R19049 CSoutput.n174 CSoutput.n151 4.5005
R19050 CSoutput.n174 CSoutput.n152 4.5005
R19051 CSoutput.n173 CSoutput.n147 4.5005
R19052 CSoutput.n173 CSoutput.n149 4.5005
R19053 CSoutput.n173 CSoutput.n146 4.5005
R19054 CSoutput.n173 CSoutput.n150 4.5005
R19055 CSoutput.n173 CSoutput.n145 4.5005
R19056 CSoutput.n173 CSoutput.t109 4.5005
R19057 CSoutput.n173 CSoutput.n144 4.5005
R19058 CSoutput.n173 CSoutput.n151 4.5005
R19059 CSoutput.n173 CSoutput.n152 4.5005
R19060 CSoutput.n156 CSoutput.n147 4.5005
R19061 CSoutput.n156 CSoutput.n149 4.5005
R19062 CSoutput.n156 CSoutput.n146 4.5005
R19063 CSoutput.n156 CSoutput.n150 4.5005
R19064 CSoutput.n156 CSoutput.n145 4.5005
R19065 CSoutput.n156 CSoutput.t109 4.5005
R19066 CSoutput.n156 CSoutput.n144 4.5005
R19067 CSoutput.n156 CSoutput.n151 4.5005
R19068 CSoutput.n156 CSoutput.n152 4.5005
R19069 CSoutput.n248 CSoutput.n147 4.5005
R19070 CSoutput.n248 CSoutput.n149 4.5005
R19071 CSoutput.n248 CSoutput.n146 4.5005
R19072 CSoutput.n248 CSoutput.n150 4.5005
R19073 CSoutput.n248 CSoutput.n145 4.5005
R19074 CSoutput.n248 CSoutput.t109 4.5005
R19075 CSoutput.n248 CSoutput.n144 4.5005
R19076 CSoutput.n248 CSoutput.n151 4.5005
R19077 CSoutput.n248 CSoutput.n152 4.5005
R19078 CSoutput.n235 CSoutput.n206 4.5005
R19079 CSoutput.n235 CSoutput.n212 4.5005
R19080 CSoutput.n193 CSoutput.n182 4.5005
R19081 CSoutput.n193 CSoutput.n184 4.5005
R19082 CSoutput.n193 CSoutput.n181 4.5005
R19083 CSoutput.n193 CSoutput.n185 4.5005
R19084 CSoutput.n193 CSoutput.n180 4.5005
R19085 CSoutput.n193 CSoutput.t99 4.5005
R19086 CSoutput.n193 CSoutput.n179 4.5005
R19087 CSoutput.n193 CSoutput.n186 4.5005
R19088 CSoutput.n235 CSoutput.n193 4.5005
R19089 CSoutput.n214 CSoutput.n182 4.5005
R19090 CSoutput.n214 CSoutput.n184 4.5005
R19091 CSoutput.n214 CSoutput.n181 4.5005
R19092 CSoutput.n214 CSoutput.n185 4.5005
R19093 CSoutput.n214 CSoutput.n180 4.5005
R19094 CSoutput.n214 CSoutput.t99 4.5005
R19095 CSoutput.n214 CSoutput.n179 4.5005
R19096 CSoutput.n214 CSoutput.n186 4.5005
R19097 CSoutput.n235 CSoutput.n214 4.5005
R19098 CSoutput.n192 CSoutput.n182 4.5005
R19099 CSoutput.n192 CSoutput.n184 4.5005
R19100 CSoutput.n192 CSoutput.n181 4.5005
R19101 CSoutput.n192 CSoutput.n185 4.5005
R19102 CSoutput.n192 CSoutput.n180 4.5005
R19103 CSoutput.n192 CSoutput.t99 4.5005
R19104 CSoutput.n192 CSoutput.n179 4.5005
R19105 CSoutput.n192 CSoutput.n186 4.5005
R19106 CSoutput.n235 CSoutput.n192 4.5005
R19107 CSoutput.n216 CSoutput.n182 4.5005
R19108 CSoutput.n216 CSoutput.n184 4.5005
R19109 CSoutput.n216 CSoutput.n181 4.5005
R19110 CSoutput.n216 CSoutput.n185 4.5005
R19111 CSoutput.n216 CSoutput.n180 4.5005
R19112 CSoutput.n216 CSoutput.t99 4.5005
R19113 CSoutput.n216 CSoutput.n179 4.5005
R19114 CSoutput.n216 CSoutput.n186 4.5005
R19115 CSoutput.n235 CSoutput.n216 4.5005
R19116 CSoutput.n182 CSoutput.n177 4.5005
R19117 CSoutput.n184 CSoutput.n177 4.5005
R19118 CSoutput.n181 CSoutput.n177 4.5005
R19119 CSoutput.n185 CSoutput.n177 4.5005
R19120 CSoutput.n180 CSoutput.n177 4.5005
R19121 CSoutput.t99 CSoutput.n177 4.5005
R19122 CSoutput.n179 CSoutput.n177 4.5005
R19123 CSoutput.n186 CSoutput.n177 4.5005
R19124 CSoutput.n238 CSoutput.n182 4.5005
R19125 CSoutput.n238 CSoutput.n184 4.5005
R19126 CSoutput.n238 CSoutput.n181 4.5005
R19127 CSoutput.n238 CSoutput.n185 4.5005
R19128 CSoutput.n238 CSoutput.n180 4.5005
R19129 CSoutput.n238 CSoutput.t99 4.5005
R19130 CSoutput.n238 CSoutput.n179 4.5005
R19131 CSoutput.n238 CSoutput.n186 4.5005
R19132 CSoutput.n236 CSoutput.n182 4.5005
R19133 CSoutput.n236 CSoutput.n184 4.5005
R19134 CSoutput.n236 CSoutput.n181 4.5005
R19135 CSoutput.n236 CSoutput.n185 4.5005
R19136 CSoutput.n236 CSoutput.n180 4.5005
R19137 CSoutput.n236 CSoutput.t99 4.5005
R19138 CSoutput.n236 CSoutput.n179 4.5005
R19139 CSoutput.n236 CSoutput.n186 4.5005
R19140 CSoutput.n236 CSoutput.n235 4.5005
R19141 CSoutput.n218 CSoutput.n182 4.5005
R19142 CSoutput.n218 CSoutput.n184 4.5005
R19143 CSoutput.n218 CSoutput.n181 4.5005
R19144 CSoutput.n218 CSoutput.n185 4.5005
R19145 CSoutput.n218 CSoutput.n180 4.5005
R19146 CSoutput.n218 CSoutput.t99 4.5005
R19147 CSoutput.n218 CSoutput.n179 4.5005
R19148 CSoutput.n218 CSoutput.n186 4.5005
R19149 CSoutput.n235 CSoutput.n218 4.5005
R19150 CSoutput.n190 CSoutput.n182 4.5005
R19151 CSoutput.n190 CSoutput.n184 4.5005
R19152 CSoutput.n190 CSoutput.n181 4.5005
R19153 CSoutput.n190 CSoutput.n185 4.5005
R19154 CSoutput.n190 CSoutput.n180 4.5005
R19155 CSoutput.n190 CSoutput.t99 4.5005
R19156 CSoutput.n190 CSoutput.n179 4.5005
R19157 CSoutput.n190 CSoutput.n186 4.5005
R19158 CSoutput.n235 CSoutput.n190 4.5005
R19159 CSoutput.n220 CSoutput.n182 4.5005
R19160 CSoutput.n220 CSoutput.n184 4.5005
R19161 CSoutput.n220 CSoutput.n181 4.5005
R19162 CSoutput.n220 CSoutput.n185 4.5005
R19163 CSoutput.n220 CSoutput.n180 4.5005
R19164 CSoutput.n220 CSoutput.t99 4.5005
R19165 CSoutput.n220 CSoutput.n179 4.5005
R19166 CSoutput.n220 CSoutput.n186 4.5005
R19167 CSoutput.n235 CSoutput.n220 4.5005
R19168 CSoutput.n189 CSoutput.n182 4.5005
R19169 CSoutput.n189 CSoutput.n184 4.5005
R19170 CSoutput.n189 CSoutput.n181 4.5005
R19171 CSoutput.n189 CSoutput.n185 4.5005
R19172 CSoutput.n189 CSoutput.n180 4.5005
R19173 CSoutput.n189 CSoutput.t99 4.5005
R19174 CSoutput.n189 CSoutput.n179 4.5005
R19175 CSoutput.n189 CSoutput.n186 4.5005
R19176 CSoutput.n235 CSoutput.n189 4.5005
R19177 CSoutput.n234 CSoutput.n182 4.5005
R19178 CSoutput.n234 CSoutput.n184 4.5005
R19179 CSoutput.n234 CSoutput.n181 4.5005
R19180 CSoutput.n234 CSoutput.n185 4.5005
R19181 CSoutput.n234 CSoutput.n180 4.5005
R19182 CSoutput.n234 CSoutput.t99 4.5005
R19183 CSoutput.n234 CSoutput.n179 4.5005
R19184 CSoutput.n234 CSoutput.n186 4.5005
R19185 CSoutput.n235 CSoutput.n234 4.5005
R19186 CSoutput.n233 CSoutput.n118 4.5005
R19187 CSoutput.n134 CSoutput.n118 4.5005
R19188 CSoutput.n129 CSoutput.n113 4.5005
R19189 CSoutput.n129 CSoutput.n115 4.5005
R19190 CSoutput.n129 CSoutput.n112 4.5005
R19191 CSoutput.n129 CSoutput.n116 4.5005
R19192 CSoutput.n129 CSoutput.n111 4.5005
R19193 CSoutput.n129 CSoutput.t106 4.5005
R19194 CSoutput.n129 CSoutput.n110 4.5005
R19195 CSoutput.n129 CSoutput.n117 4.5005
R19196 CSoutput.n129 CSoutput.n118 4.5005
R19197 CSoutput.n127 CSoutput.n113 4.5005
R19198 CSoutput.n127 CSoutput.n115 4.5005
R19199 CSoutput.n127 CSoutput.n112 4.5005
R19200 CSoutput.n127 CSoutput.n116 4.5005
R19201 CSoutput.n127 CSoutput.n111 4.5005
R19202 CSoutput.n127 CSoutput.t106 4.5005
R19203 CSoutput.n127 CSoutput.n110 4.5005
R19204 CSoutput.n127 CSoutput.n117 4.5005
R19205 CSoutput.n127 CSoutput.n118 4.5005
R19206 CSoutput.n126 CSoutput.n113 4.5005
R19207 CSoutput.n126 CSoutput.n115 4.5005
R19208 CSoutput.n126 CSoutput.n112 4.5005
R19209 CSoutput.n126 CSoutput.n116 4.5005
R19210 CSoutput.n126 CSoutput.n111 4.5005
R19211 CSoutput.n126 CSoutput.t106 4.5005
R19212 CSoutput.n126 CSoutput.n110 4.5005
R19213 CSoutput.n126 CSoutput.n117 4.5005
R19214 CSoutput.n126 CSoutput.n118 4.5005
R19215 CSoutput.n255 CSoutput.n113 4.5005
R19216 CSoutput.n255 CSoutput.n115 4.5005
R19217 CSoutput.n255 CSoutput.n112 4.5005
R19218 CSoutput.n255 CSoutput.n116 4.5005
R19219 CSoutput.n255 CSoutput.n111 4.5005
R19220 CSoutput.n255 CSoutput.t106 4.5005
R19221 CSoutput.n255 CSoutput.n110 4.5005
R19222 CSoutput.n255 CSoutput.n117 4.5005
R19223 CSoutput.n255 CSoutput.n118 4.5005
R19224 CSoutput.n253 CSoutput.n113 4.5005
R19225 CSoutput.n253 CSoutput.n115 4.5005
R19226 CSoutput.n253 CSoutput.n112 4.5005
R19227 CSoutput.n253 CSoutput.n116 4.5005
R19228 CSoutput.n253 CSoutput.n111 4.5005
R19229 CSoutput.n253 CSoutput.t106 4.5005
R19230 CSoutput.n253 CSoutput.n110 4.5005
R19231 CSoutput.n253 CSoutput.n117 4.5005
R19232 CSoutput.n251 CSoutput.n113 4.5005
R19233 CSoutput.n251 CSoutput.n115 4.5005
R19234 CSoutput.n251 CSoutput.n112 4.5005
R19235 CSoutput.n251 CSoutput.n116 4.5005
R19236 CSoutput.n251 CSoutput.n111 4.5005
R19237 CSoutput.n251 CSoutput.t106 4.5005
R19238 CSoutput.n251 CSoutput.n110 4.5005
R19239 CSoutput.n251 CSoutput.n117 4.5005
R19240 CSoutput.n137 CSoutput.n113 4.5005
R19241 CSoutput.n137 CSoutput.n115 4.5005
R19242 CSoutput.n137 CSoutput.n112 4.5005
R19243 CSoutput.n137 CSoutput.n116 4.5005
R19244 CSoutput.n137 CSoutput.n111 4.5005
R19245 CSoutput.n137 CSoutput.t106 4.5005
R19246 CSoutput.n137 CSoutput.n110 4.5005
R19247 CSoutput.n137 CSoutput.n117 4.5005
R19248 CSoutput.n137 CSoutput.n118 4.5005
R19249 CSoutput.n136 CSoutput.n113 4.5005
R19250 CSoutput.n136 CSoutput.n115 4.5005
R19251 CSoutput.n136 CSoutput.n112 4.5005
R19252 CSoutput.n136 CSoutput.n116 4.5005
R19253 CSoutput.n136 CSoutput.n111 4.5005
R19254 CSoutput.n136 CSoutput.t106 4.5005
R19255 CSoutput.n136 CSoutput.n110 4.5005
R19256 CSoutput.n136 CSoutput.n117 4.5005
R19257 CSoutput.n136 CSoutput.n118 4.5005
R19258 CSoutput.n140 CSoutput.n113 4.5005
R19259 CSoutput.n140 CSoutput.n115 4.5005
R19260 CSoutput.n140 CSoutput.n112 4.5005
R19261 CSoutput.n140 CSoutput.n116 4.5005
R19262 CSoutput.n140 CSoutput.n111 4.5005
R19263 CSoutput.n140 CSoutput.t106 4.5005
R19264 CSoutput.n140 CSoutput.n110 4.5005
R19265 CSoutput.n140 CSoutput.n117 4.5005
R19266 CSoutput.n140 CSoutput.n118 4.5005
R19267 CSoutput.n139 CSoutput.n113 4.5005
R19268 CSoutput.n139 CSoutput.n115 4.5005
R19269 CSoutput.n139 CSoutput.n112 4.5005
R19270 CSoutput.n139 CSoutput.n116 4.5005
R19271 CSoutput.n139 CSoutput.n111 4.5005
R19272 CSoutput.n139 CSoutput.t106 4.5005
R19273 CSoutput.n139 CSoutput.n110 4.5005
R19274 CSoutput.n139 CSoutput.n117 4.5005
R19275 CSoutput.n139 CSoutput.n118 4.5005
R19276 CSoutput.n122 CSoutput.n113 4.5005
R19277 CSoutput.n122 CSoutput.n115 4.5005
R19278 CSoutput.n122 CSoutput.n112 4.5005
R19279 CSoutput.n122 CSoutput.n116 4.5005
R19280 CSoutput.n122 CSoutput.n111 4.5005
R19281 CSoutput.n122 CSoutput.t106 4.5005
R19282 CSoutput.n122 CSoutput.n110 4.5005
R19283 CSoutput.n122 CSoutput.n117 4.5005
R19284 CSoutput.n122 CSoutput.n118 4.5005
R19285 CSoutput.n258 CSoutput.n113 4.5005
R19286 CSoutput.n258 CSoutput.n115 4.5005
R19287 CSoutput.n258 CSoutput.n112 4.5005
R19288 CSoutput.n258 CSoutput.n116 4.5005
R19289 CSoutput.n258 CSoutput.n111 4.5005
R19290 CSoutput.n258 CSoutput.t106 4.5005
R19291 CSoutput.n258 CSoutput.n110 4.5005
R19292 CSoutput.n258 CSoutput.n117 4.5005
R19293 CSoutput.n258 CSoutput.n118 4.5005
R19294 CSoutput.n44 CSoutput.n43 3.79402
R19295 CSoutput.n49 CSoutput.n48 3.79402
R19296 CSoutput.n287 CSoutput.n277 3.72967
R19297 CSoutput.n107 CSoutput.n97 3.72967
R19298 CSoutput.n321 CSoutput.n320 3.60477
R19299 CSoutput.n301 CSoutput.t66 3.3005
R19300 CSoutput.n301 CSoutput.t64 3.3005
R19301 CSoutput.n299 CSoutput.t57 3.3005
R19302 CSoutput.n299 CSoutput.t56 3.3005
R19303 CSoutput.n297 CSoutput.t40 3.3005
R19304 CSoutput.n297 CSoutput.t42 3.3005
R19305 CSoutput.n296 CSoutput.t55 3.3005
R19306 CSoutput.n296 CSoutput.t41 3.3005
R19307 CSoutput.n294 CSoutput.t61 3.3005
R19308 CSoutput.n294 CSoutput.t59 3.3005
R19309 CSoutput.n292 CSoutput.t52 3.3005
R19310 CSoutput.n292 CSoutput.t51 3.3005
R19311 CSoutput.n290 CSoutput.t63 3.3005
R19312 CSoutput.n290 CSoutput.t68 3.3005
R19313 CSoutput.n289 CSoutput.t48 3.3005
R19314 CSoutput.n289 CSoutput.t67 3.3005
R19315 CSoutput.n312 CSoutput.t49 3.3005
R19316 CSoutput.n312 CSoutput.t43 3.3005
R19317 CSoutput.n313 CSoutput.t50 3.3005
R19318 CSoutput.n313 CSoutput.t58 3.3005
R19319 CSoutput.n315 CSoutput.t65 3.3005
R19320 CSoutput.n315 CSoutput.t69 3.3005
R19321 CSoutput.n317 CSoutput.t53 3.3005
R19322 CSoutput.n317 CSoutput.t44 3.3005
R19323 CSoutput.n305 CSoutput.t45 3.3005
R19324 CSoutput.n305 CSoutput.t70 3.3005
R19325 CSoutput.n306 CSoutput.t46 3.3005
R19326 CSoutput.n306 CSoutput.t54 3.3005
R19327 CSoutput.n308 CSoutput.t60 3.3005
R19328 CSoutput.n308 CSoutput.t62 3.3005
R19329 CSoutput.n310 CSoutput.t47 3.3005
R19330 CSoutput.n310 CSoutput.t71 3.3005
R19331 CSoutput.n320 CSoutput.n304 2.72117
R19332 CSoutput.n288 CSoutput.n108 2.58832
R19333 CSoutput.n75 CSoutput.n1 2.45513
R19334 CSoutput.n199 CSoutput.n197 2.251
R19335 CSoutput.n199 CSoutput.n196 2.251
R19336 CSoutput.n199 CSoutput.n195 2.251
R19337 CSoutput.n199 CSoutput.n194 2.251
R19338 CSoutput.n168 CSoutput.n167 2.251
R19339 CSoutput.n168 CSoutput.n166 2.251
R19340 CSoutput.n168 CSoutput.n165 2.251
R19341 CSoutput.n168 CSoutput.n164 2.251
R19342 CSoutput.n241 CSoutput.n240 2.251
R19343 CSoutput.n206 CSoutput.n204 2.251
R19344 CSoutput.n206 CSoutput.n203 2.251
R19345 CSoutput.n206 CSoutput.n202 2.251
R19346 CSoutput.n224 CSoutput.n206 2.251
R19347 CSoutput.n212 CSoutput.n211 2.251
R19348 CSoutput.n212 CSoutput.n210 2.251
R19349 CSoutput.n212 CSoutput.n209 2.251
R19350 CSoutput.n212 CSoutput.n208 2.251
R19351 CSoutput.n238 CSoutput.n178 2.251
R19352 CSoutput.n233 CSoutput.n231 2.251
R19353 CSoutput.n233 CSoutput.n230 2.251
R19354 CSoutput.n233 CSoutput.n229 2.251
R19355 CSoutput.n233 CSoutput.n228 2.251
R19356 CSoutput.n134 CSoutput.n133 2.251
R19357 CSoutput.n134 CSoutput.n132 2.251
R19358 CSoutput.n134 CSoutput.n131 2.251
R19359 CSoutput.n134 CSoutput.n130 2.251
R19360 CSoutput.n251 CSoutput.n250 2.251
R19361 CSoutput.n168 CSoutput.n148 2.2505
R19362 CSoutput.n163 CSoutput.n148 2.2505
R19363 CSoutput.n161 CSoutput.n148 2.2505
R19364 CSoutput.n160 CSoutput.n148 2.2505
R19365 CSoutput.n245 CSoutput.n148 2.2505
R19366 CSoutput.n243 CSoutput.n148 2.2505
R19367 CSoutput.n241 CSoutput.n148 2.2505
R19368 CSoutput.n171 CSoutput.n148 2.2505
R19369 CSoutput.n170 CSoutput.n148 2.2505
R19370 CSoutput.n174 CSoutput.n148 2.2505
R19371 CSoutput.n173 CSoutput.n148 2.2505
R19372 CSoutput.n156 CSoutput.n148 2.2505
R19373 CSoutput.n248 CSoutput.n148 2.2505
R19374 CSoutput.n248 CSoutput.n247 2.2505
R19375 CSoutput.n212 CSoutput.n183 2.2505
R19376 CSoutput.n193 CSoutput.n183 2.2505
R19377 CSoutput.n214 CSoutput.n183 2.2505
R19378 CSoutput.n192 CSoutput.n183 2.2505
R19379 CSoutput.n216 CSoutput.n183 2.2505
R19380 CSoutput.n183 CSoutput.n177 2.2505
R19381 CSoutput.n238 CSoutput.n183 2.2505
R19382 CSoutput.n236 CSoutput.n183 2.2505
R19383 CSoutput.n218 CSoutput.n183 2.2505
R19384 CSoutput.n190 CSoutput.n183 2.2505
R19385 CSoutput.n220 CSoutput.n183 2.2505
R19386 CSoutput.n189 CSoutput.n183 2.2505
R19387 CSoutput.n234 CSoutput.n183 2.2505
R19388 CSoutput.n234 CSoutput.n187 2.2505
R19389 CSoutput.n134 CSoutput.n114 2.2505
R19390 CSoutput.n129 CSoutput.n114 2.2505
R19391 CSoutput.n127 CSoutput.n114 2.2505
R19392 CSoutput.n126 CSoutput.n114 2.2505
R19393 CSoutput.n255 CSoutput.n114 2.2505
R19394 CSoutput.n253 CSoutput.n114 2.2505
R19395 CSoutput.n251 CSoutput.n114 2.2505
R19396 CSoutput.n137 CSoutput.n114 2.2505
R19397 CSoutput.n136 CSoutput.n114 2.2505
R19398 CSoutput.n140 CSoutput.n114 2.2505
R19399 CSoutput.n139 CSoutput.n114 2.2505
R19400 CSoutput.n122 CSoutput.n114 2.2505
R19401 CSoutput.n258 CSoutput.n114 2.2505
R19402 CSoutput.n258 CSoutput.n257 2.2505
R19403 CSoutput.n176 CSoutput.n169 2.25024
R19404 CSoutput.n176 CSoutput.n162 2.25024
R19405 CSoutput.n244 CSoutput.n176 2.25024
R19406 CSoutput.n176 CSoutput.n172 2.25024
R19407 CSoutput.n176 CSoutput.n175 2.25024
R19408 CSoutput.n176 CSoutput.n143 2.25024
R19409 CSoutput.n226 CSoutput.n223 2.25024
R19410 CSoutput.n226 CSoutput.n222 2.25024
R19411 CSoutput.n226 CSoutput.n221 2.25024
R19412 CSoutput.n226 CSoutput.n188 2.25024
R19413 CSoutput.n226 CSoutput.n225 2.25024
R19414 CSoutput.n227 CSoutput.n226 2.25024
R19415 CSoutput.n142 CSoutput.n135 2.25024
R19416 CSoutput.n142 CSoutput.n128 2.25024
R19417 CSoutput.n254 CSoutput.n142 2.25024
R19418 CSoutput.n142 CSoutput.n138 2.25024
R19419 CSoutput.n142 CSoutput.n141 2.25024
R19420 CSoutput.n142 CSoutput.n109 2.25024
R19421 CSoutput.n243 CSoutput.n153 1.50111
R19422 CSoutput.n191 CSoutput.n177 1.50111
R19423 CSoutput.n253 CSoutput.n119 1.50111
R19424 CSoutput.n199 CSoutput.n198 1.501
R19425 CSoutput.n206 CSoutput.n205 1.501
R19426 CSoutput.n233 CSoutput.n232 1.501
R19427 CSoutput.n247 CSoutput.n158 1.12536
R19428 CSoutput.n247 CSoutput.n159 1.12536
R19429 CSoutput.n247 CSoutput.n246 1.12536
R19430 CSoutput.n207 CSoutput.n187 1.12536
R19431 CSoutput.n213 CSoutput.n187 1.12536
R19432 CSoutput.n215 CSoutput.n187 1.12536
R19433 CSoutput.n257 CSoutput.n124 1.12536
R19434 CSoutput.n257 CSoutput.n125 1.12536
R19435 CSoutput.n257 CSoutput.n256 1.12536
R19436 CSoutput.n247 CSoutput.n154 1.12536
R19437 CSoutput.n247 CSoutput.n155 1.12536
R19438 CSoutput.n247 CSoutput.n157 1.12536
R19439 CSoutput.n237 CSoutput.n187 1.12536
R19440 CSoutput.n217 CSoutput.n187 1.12536
R19441 CSoutput.n219 CSoutput.n187 1.12536
R19442 CSoutput.n257 CSoutput.n120 1.12536
R19443 CSoutput.n257 CSoutput.n121 1.12536
R19444 CSoutput.n257 CSoutput.n123 1.12536
R19445 CSoutput.n300 CSoutput.n298 1.00481
R19446 CSoutput.n302 CSoutput.n300 1.00481
R19447 CSoutput.n293 CSoutput.n291 1.00481
R19448 CSoutput.n295 CSoutput.n293 1.00481
R19449 CSoutput.n318 CSoutput.n316 1.00481
R19450 CSoutput.n316 CSoutput.n314 1.00481
R19451 CSoutput.n311 CSoutput.n309 1.00481
R19452 CSoutput.n309 CSoutput.n307 1.00481
R19453 CSoutput.n31 CSoutput.n30 0.669944
R19454 CSoutput.n62 CSoutput.n61 0.669944
R19455 CSoutput.n282 CSoutput.n280 0.573776
R19456 CSoutput.n284 CSoutput.n282 0.573776
R19457 CSoutput.n286 CSoutput.n284 0.573776
R19458 CSoutput.n272 CSoutput.n270 0.573776
R19459 CSoutput.n274 CSoutput.n272 0.573776
R19460 CSoutput.n276 CSoutput.n274 0.573776
R19461 CSoutput.n263 CSoutput.n261 0.573776
R19462 CSoutput.n265 CSoutput.n263 0.573776
R19463 CSoutput.n267 CSoutput.n265 0.573776
R19464 CSoutput.n106 CSoutput.n104 0.573776
R19465 CSoutput.n104 CSoutput.n102 0.573776
R19466 CSoutput.n102 CSoutput.n100 0.573776
R19467 CSoutput.n96 CSoutput.n94 0.573776
R19468 CSoutput.n94 CSoutput.n92 0.573776
R19469 CSoutput.n92 CSoutput.n90 0.573776
R19470 CSoutput.n87 CSoutput.n85 0.573776
R19471 CSoutput.n85 CSoutput.n83 0.573776
R19472 CSoutput.n83 CSoutput.n81 0.573776
R19473 CSoutput.n321 CSoutput.n258 0.534733
R19474 CSoutput.n21 CSoutput.n20 0.169105
R19475 CSoutput.n21 CSoutput.n16 0.169105
R19476 CSoutput.n26 CSoutput.n16 0.169105
R19477 CSoutput.n27 CSoutput.n26 0.169105
R19478 CSoutput.n27 CSoutput.n14 0.169105
R19479 CSoutput.n32 CSoutput.n14 0.169105
R19480 CSoutput.n33 CSoutput.n32 0.169105
R19481 CSoutput.n34 CSoutput.n33 0.169105
R19482 CSoutput.n34 CSoutput.n12 0.169105
R19483 CSoutput.n39 CSoutput.n12 0.169105
R19484 CSoutput.n40 CSoutput.n39 0.169105
R19485 CSoutput.n40 CSoutput.n10 0.169105
R19486 CSoutput.n45 CSoutput.n10 0.169105
R19487 CSoutput.n46 CSoutput.n45 0.169105
R19488 CSoutput.n47 CSoutput.n46 0.169105
R19489 CSoutput.n47 CSoutput.n8 0.169105
R19490 CSoutput.n52 CSoutput.n8 0.169105
R19491 CSoutput.n53 CSoutput.n52 0.169105
R19492 CSoutput.n53 CSoutput.n6 0.169105
R19493 CSoutput.n58 CSoutput.n6 0.169105
R19494 CSoutput.n59 CSoutput.n58 0.169105
R19495 CSoutput.n60 CSoutput.n59 0.169105
R19496 CSoutput.n60 CSoutput.n4 0.169105
R19497 CSoutput.n66 CSoutput.n4 0.169105
R19498 CSoutput.n67 CSoutput.n66 0.169105
R19499 CSoutput.n68 CSoutput.n67 0.169105
R19500 CSoutput.n68 CSoutput.n2 0.169105
R19501 CSoutput.n73 CSoutput.n2 0.169105
R19502 CSoutput.n74 CSoutput.n73 0.169105
R19503 CSoutput.n74 CSoutput.n0 0.169105
R19504 CSoutput.n78 CSoutput.n0 0.169105
R19505 CSoutput.n201 CSoutput.n200 0.0910737
R19506 CSoutput.n252 CSoutput.n249 0.0723685
R19507 CSoutput.n206 CSoutput.n201 0.0522944
R19508 CSoutput.n249 CSoutput.n248 0.0499135
R19509 CSoutput.n200 CSoutput.n199 0.0499135
R19510 CSoutput.n234 CSoutput.n233 0.0464294
R19511 CSoutput.n242 CSoutput.n239 0.0391444
R19512 CSoutput.n201 CSoutput.t93 0.023435
R19513 CSoutput.n249 CSoutput.t97 0.02262
R19514 CSoutput.n200 CSoutput.t98 0.02262
R19515 CSoutput CSoutput.n321 0.0052
R19516 CSoutput.n171 CSoutput.n154 0.00365111
R19517 CSoutput.n174 CSoutput.n155 0.00365111
R19518 CSoutput.n157 CSoutput.n156 0.00365111
R19519 CSoutput.n199 CSoutput.n158 0.00365111
R19520 CSoutput.n163 CSoutput.n159 0.00365111
R19521 CSoutput.n246 CSoutput.n160 0.00365111
R19522 CSoutput.n237 CSoutput.n236 0.00365111
R19523 CSoutput.n217 CSoutput.n190 0.00365111
R19524 CSoutput.n219 CSoutput.n189 0.00365111
R19525 CSoutput.n207 CSoutput.n206 0.00365111
R19526 CSoutput.n213 CSoutput.n193 0.00365111
R19527 CSoutput.n215 CSoutput.n192 0.00365111
R19528 CSoutput.n137 CSoutput.n120 0.00365111
R19529 CSoutput.n140 CSoutput.n121 0.00365111
R19530 CSoutput.n123 CSoutput.n122 0.00365111
R19531 CSoutput.n233 CSoutput.n124 0.00365111
R19532 CSoutput.n129 CSoutput.n125 0.00365111
R19533 CSoutput.n256 CSoutput.n126 0.00365111
R19534 CSoutput.n168 CSoutput.n158 0.00340054
R19535 CSoutput.n161 CSoutput.n159 0.00340054
R19536 CSoutput.n246 CSoutput.n245 0.00340054
R19537 CSoutput.n241 CSoutput.n154 0.00340054
R19538 CSoutput.n170 CSoutput.n155 0.00340054
R19539 CSoutput.n173 CSoutput.n157 0.00340054
R19540 CSoutput.n212 CSoutput.n207 0.00340054
R19541 CSoutput.n214 CSoutput.n213 0.00340054
R19542 CSoutput.n216 CSoutput.n215 0.00340054
R19543 CSoutput.n238 CSoutput.n237 0.00340054
R19544 CSoutput.n218 CSoutput.n217 0.00340054
R19545 CSoutput.n220 CSoutput.n219 0.00340054
R19546 CSoutput.n134 CSoutput.n124 0.00340054
R19547 CSoutput.n127 CSoutput.n125 0.00340054
R19548 CSoutput.n256 CSoutput.n255 0.00340054
R19549 CSoutput.n251 CSoutput.n120 0.00340054
R19550 CSoutput.n136 CSoutput.n121 0.00340054
R19551 CSoutput.n139 CSoutput.n123 0.00340054
R19552 CSoutput.n169 CSoutput.n163 0.00252698
R19553 CSoutput.n162 CSoutput.n160 0.00252698
R19554 CSoutput.n244 CSoutput.n243 0.00252698
R19555 CSoutput.n172 CSoutput.n170 0.00252698
R19556 CSoutput.n175 CSoutput.n173 0.00252698
R19557 CSoutput.n248 CSoutput.n143 0.00252698
R19558 CSoutput.n169 CSoutput.n168 0.00252698
R19559 CSoutput.n162 CSoutput.n161 0.00252698
R19560 CSoutput.n245 CSoutput.n244 0.00252698
R19561 CSoutput.n172 CSoutput.n171 0.00252698
R19562 CSoutput.n175 CSoutput.n174 0.00252698
R19563 CSoutput.n156 CSoutput.n143 0.00252698
R19564 CSoutput.n223 CSoutput.n193 0.00252698
R19565 CSoutput.n222 CSoutput.n192 0.00252698
R19566 CSoutput.n221 CSoutput.n177 0.00252698
R19567 CSoutput.n218 CSoutput.n188 0.00252698
R19568 CSoutput.n225 CSoutput.n220 0.00252698
R19569 CSoutput.n234 CSoutput.n227 0.00252698
R19570 CSoutput.n223 CSoutput.n212 0.00252698
R19571 CSoutput.n222 CSoutput.n214 0.00252698
R19572 CSoutput.n221 CSoutput.n216 0.00252698
R19573 CSoutput.n236 CSoutput.n188 0.00252698
R19574 CSoutput.n225 CSoutput.n190 0.00252698
R19575 CSoutput.n227 CSoutput.n189 0.00252698
R19576 CSoutput.n135 CSoutput.n129 0.00252698
R19577 CSoutput.n128 CSoutput.n126 0.00252698
R19578 CSoutput.n254 CSoutput.n253 0.00252698
R19579 CSoutput.n138 CSoutput.n136 0.00252698
R19580 CSoutput.n141 CSoutput.n139 0.00252698
R19581 CSoutput.n258 CSoutput.n109 0.00252698
R19582 CSoutput.n135 CSoutput.n134 0.00252698
R19583 CSoutput.n128 CSoutput.n127 0.00252698
R19584 CSoutput.n255 CSoutput.n254 0.00252698
R19585 CSoutput.n138 CSoutput.n137 0.00252698
R19586 CSoutput.n141 CSoutput.n140 0.00252698
R19587 CSoutput.n122 CSoutput.n109 0.00252698
R19588 CSoutput.n243 CSoutput.n242 0.0020275
R19589 CSoutput.n242 CSoutput.n241 0.0020275
R19590 CSoutput.n239 CSoutput.n177 0.0020275
R19591 CSoutput.n239 CSoutput.n238 0.0020275
R19592 CSoutput.n253 CSoutput.n252 0.0020275
R19593 CSoutput.n252 CSoutput.n251 0.0020275
R19594 CSoutput.n153 CSoutput.n152 0.00166668
R19595 CSoutput.n235 CSoutput.n191 0.00166668
R19596 CSoutput.n119 CSoutput.n118 0.00166668
R19597 CSoutput.n257 CSoutput.n119 0.00133328
R19598 CSoutput.n191 CSoutput.n187 0.00133328
R19599 CSoutput.n247 CSoutput.n153 0.00133328
R19600 CSoutput.n250 CSoutput.n142 0.001
R19601 CSoutput.n228 CSoutput.n142 0.001
R19602 CSoutput.n130 CSoutput.n110 0.001
R19603 CSoutput.n229 CSoutput.n110 0.001
R19604 CSoutput.n131 CSoutput.n111 0.001
R19605 CSoutput.n230 CSoutput.n111 0.001
R19606 CSoutput.n132 CSoutput.n112 0.001
R19607 CSoutput.n231 CSoutput.n112 0.001
R19608 CSoutput.n133 CSoutput.n113 0.001
R19609 CSoutput.n232 CSoutput.n113 0.001
R19610 CSoutput.n226 CSoutput.n178 0.001
R19611 CSoutput.n226 CSoutput.n224 0.001
R19612 CSoutput.n208 CSoutput.n179 0.001
R19613 CSoutput.n202 CSoutput.n179 0.001
R19614 CSoutput.n209 CSoutput.n180 0.001
R19615 CSoutput.n203 CSoutput.n180 0.001
R19616 CSoutput.n210 CSoutput.n181 0.001
R19617 CSoutput.n204 CSoutput.n181 0.001
R19618 CSoutput.n211 CSoutput.n182 0.001
R19619 CSoutput.n205 CSoutput.n182 0.001
R19620 CSoutput.n240 CSoutput.n176 0.001
R19621 CSoutput.n194 CSoutput.n176 0.001
R19622 CSoutput.n164 CSoutput.n144 0.001
R19623 CSoutput.n195 CSoutput.n144 0.001
R19624 CSoutput.n165 CSoutput.n145 0.001
R19625 CSoutput.n196 CSoutput.n145 0.001
R19626 CSoutput.n166 CSoutput.n146 0.001
R19627 CSoutput.n197 CSoutput.n146 0.001
R19628 CSoutput.n167 CSoutput.n147 0.001
R19629 CSoutput.n198 CSoutput.n147 0.001
R19630 CSoutput.n198 CSoutput.n148 0.001
R19631 CSoutput.n197 CSoutput.n149 0.001
R19632 CSoutput.n196 CSoutput.n150 0.001
R19633 CSoutput.n195 CSoutput.t109 0.001
R19634 CSoutput.n194 CSoutput.n151 0.001
R19635 CSoutput.n167 CSoutput.n149 0.001
R19636 CSoutput.n166 CSoutput.n150 0.001
R19637 CSoutput.n165 CSoutput.t109 0.001
R19638 CSoutput.n164 CSoutput.n151 0.001
R19639 CSoutput.n240 CSoutput.n152 0.001
R19640 CSoutput.n205 CSoutput.n183 0.001
R19641 CSoutput.n204 CSoutput.n184 0.001
R19642 CSoutput.n203 CSoutput.n185 0.001
R19643 CSoutput.n202 CSoutput.t99 0.001
R19644 CSoutput.n224 CSoutput.n186 0.001
R19645 CSoutput.n211 CSoutput.n184 0.001
R19646 CSoutput.n210 CSoutput.n185 0.001
R19647 CSoutput.n209 CSoutput.t99 0.001
R19648 CSoutput.n208 CSoutput.n186 0.001
R19649 CSoutput.n235 CSoutput.n178 0.001
R19650 CSoutput.n232 CSoutput.n114 0.001
R19651 CSoutput.n231 CSoutput.n115 0.001
R19652 CSoutput.n230 CSoutput.n116 0.001
R19653 CSoutput.n229 CSoutput.t106 0.001
R19654 CSoutput.n228 CSoutput.n117 0.001
R19655 CSoutput.n133 CSoutput.n115 0.001
R19656 CSoutput.n132 CSoutput.n116 0.001
R19657 CSoutput.n131 CSoutput.t106 0.001
R19658 CSoutput.n130 CSoutput.n117 0.001
R19659 CSoutput.n250 CSoutput.n118 0.001
R19660 a_n7677_7899.n153 a_n7677_7899.t76 223.136
R19661 a_n7677_7899.n164 a_n7677_7899.t48 223.136
R19662 a_n7677_7899.n176 a_n7677_7899.t21 223.136
R19663 a_n7677_7899.n108 a_n7677_7899.t58 223.136
R19664 a_n7677_7899.n122 a_n7677_7899.t31 223.136
R19665 a_n7677_7899.n137 a_n7677_7899.t39 223.136
R19666 a_n7677_7899.n11 a_n7677_7899.t40 223.097
R19667 a_n7677_7899.n10 a_n7677_7899.t65 223.097
R19668 a_n7677_7899.n9 a_n7677_7899.t74 223.097
R19669 a_n7677_7899.n117 a_n7677_7899.t20 207.983
R19670 a_n7677_7899.n131 a_n7677_7899.t50 207.983
R19671 a_n7677_7899.n146 a_n7677_7899.t32 207.983
R19672 a_n7677_7899.n159 a_n7677_7899.t36 168.701
R19673 a_n7677_7899.n158 a_n7677_7899.t69 168.701
R19674 a_n7677_7899.n149 a_n7677_7899.t24 168.701
R19675 a_n7677_7899.n155 a_n7677_7899.t78 168.701
R19676 a_n7677_7899.n154 a_n7677_7899.t56 168.701
R19677 a_n7677_7899.n150 a_n7677_7899.t34 168.701
R19678 a_n7677_7899.n151 a_n7677_7899.t62 168.701
R19679 a_n7677_7899.n152 a_n7677_7899.t43 168.701
R19680 a_n7677_7899.n170 a_n7677_7899.t61 168.701
R19681 a_n7677_7899.n169 a_n7677_7899.t42 168.701
R19682 a_n7677_7899.n160 a_n7677_7899.t51 168.701
R19683 a_n7677_7899.n166 a_n7677_7899.t49 168.701
R19684 a_n7677_7899.n165 a_n7677_7899.t29 168.701
R19685 a_n7677_7899.n161 a_n7677_7899.t59 168.701
R19686 a_n7677_7899.n162 a_n7677_7899.t37 168.701
R19687 a_n7677_7899.n163 a_n7677_7899.t71 168.701
R19688 a_n7677_7899.n182 a_n7677_7899.t68 168.701
R19689 a_n7677_7899.n181 a_n7677_7899.t22 168.701
R19690 a_n7677_7899.n172 a_n7677_7899.t66 168.701
R19691 a_n7677_7899.n180 a_n7677_7899.t64 168.701
R19692 a_n7677_7899.n179 a_n7677_7899.t77 168.701
R19693 a_n7677_7899.n173 a_n7677_7899.t30 168.701
R19694 a_n7677_7899.n174 a_n7677_7899.t57 168.701
R19695 a_n7677_7899.n175 a_n7677_7899.t70 168.701
R19696 a_n7677_7899.n107 a_n7677_7899.t28 168.701
R19697 a_n7677_7899.n106 a_n7677_7899.t52 168.701
R19698 a_n7677_7899.n105 a_n7677_7899.t73 168.701
R19699 a_n7677_7899.n111 a_n7677_7899.t41 168.701
R19700 a_n7677_7899.n112 a_n7677_7899.t60 168.701
R19701 a_n7677_7899.n23 a_n7677_7899.t72 168.701
R19702 a_n7677_7899.n114 a_n7677_7899.t54 168.701
R19703 a_n7677_7899.n115 a_n7677_7899.t75 168.701
R19704 a_n7677_7899.n121 a_n7677_7899.t55 168.701
R19705 a_n7677_7899.n120 a_n7677_7899.t23 168.701
R19706 a_n7677_7899.n119 a_n7677_7899.t46 168.701
R19707 a_n7677_7899.n125 a_n7677_7899.t67 168.701
R19708 a_n7677_7899.n126 a_n7677_7899.t33 168.701
R19709 a_n7677_7899.n25 a_n7677_7899.t45 168.701
R19710 a_n7677_7899.n128 a_n7677_7899.t25 168.701
R19711 a_n7677_7899.n129 a_n7677_7899.t47 168.701
R19712 a_n7677_7899.n136 a_n7677_7899.t27 168.701
R19713 a_n7677_7899.n135 a_n7677_7899.t53 168.701
R19714 a_n7677_7899.n134 a_n7677_7899.t44 168.701
R19715 a_n7677_7899.n140 a_n7677_7899.t35 168.701
R19716 a_n7677_7899.n141 a_n7677_7899.t79 168.701
R19717 a_n7677_7899.n27 a_n7677_7899.t63 168.701
R19718 a_n7677_7899.n143 a_n7677_7899.t38 168.701
R19719 a_n7677_7899.n144 a_n7677_7899.t26 168.701
R19720 a_n7677_7899.n19 a_n7677_7899.n0 39.6376
R19721 a_n7677_7899.n5 a_n7677_7899.n0 39.7274
R19722 a_n7677_7899.n29 a_n7677_7899.n0 68.6201
R19723 a_n7677_7899.n20 a_n7677_7899.n0 39.6373
R19724 a_n7677_7899.n156 a_n7677_7899.n0 161.3
R19725 a_n7677_7899.n1 a_n7677_7899.n157 161.3
R19726 a_n7677_7899.n21 a_n7677_7899.n1 39.7274
R19727 a_n7677_7899.n22 a_n7677_7899.n1 39.6376
R19728 a_n7677_7899.n15 a_n7677_7899.n2 39.6376
R19729 a_n7677_7899.n6 a_n7677_7899.n2 39.7274
R19730 a_n7677_7899.n30 a_n7677_7899.n2 68.6201
R19731 a_n7677_7899.n16 a_n7677_7899.n2 39.6373
R19732 a_n7677_7899.n167 a_n7677_7899.n2 161.3
R19733 a_n7677_7899.n3 a_n7677_7899.n168 161.3
R19734 a_n7677_7899.n17 a_n7677_7899.n3 39.7274
R19735 a_n7677_7899.n18 a_n7677_7899.n3 39.6376
R19736 a_n7677_7899.n35 a_n7677_7899.n33 71.8318
R19737 a_n7677_7899.n34 a_n7677_7899.n177 161.3
R19738 a_n7677_7899.n178 a_n7677_7899.n34 161.3
R19739 a_n7677_7899.n32 a_n7677_7899.n7 74.8341
R19740 a_n7677_7899.n31 a_n7677_7899.n4 68.6201
R19741 a_n7677_7899.n12 a_n7677_7899.n4 39.6373
R19742 a_n7677_7899.n4 a_n7677_7899.n8 68.6201
R19743 a_n7677_7899.n13 a_n7677_7899.n4 39.7274
R19744 a_n7677_7899.n14 a_n7677_7899.n4 39.6376
R19745 a_n7677_7899.n116 a_n7677_7899.n53 161.3
R19746 a_n7677_7899.n50 a_n7677_7899.n53 161.3
R19747 a_n7677_7899.n52 a_n7677_7899.n51 71.4497
R19748 a_n7677_7899.n49 a_n7677_7899.n48 68.7078
R19749 a_n7677_7899.n24 a_n7677_7899.n23 11.426
R19750 a_n7677_7899.n47 a_n7677_7899.n24 74.9385
R19751 a_n7677_7899.n113 a_n7677_7899.n46 161.3
R19752 a_n7677_7899.n43 a_n7677_7899.n46 161.3
R19753 a_n7677_7899.n45 a_n7677_7899.n44 71.6402
R19754 a_n7677_7899.n42 a_n7677_7899.n41 68.6201
R19755 a_n7677_7899.n38 a_n7677_7899.n40 74.8341
R19756 a_n7677_7899.n110 a_n7677_7899.n39 161.3
R19757 a_n7677_7899.n39 a_n7677_7899.n109 161.3
R19758 a_n7677_7899.n37 a_n7677_7899.n36 71.8318
R19759 a_n7677_7899.n130 a_n7677_7899.n71 161.3
R19760 a_n7677_7899.n68 a_n7677_7899.n71 161.3
R19761 a_n7677_7899.n70 a_n7677_7899.n69 71.4497
R19762 a_n7677_7899.n67 a_n7677_7899.n66 68.7078
R19763 a_n7677_7899.n26 a_n7677_7899.n25 11.426
R19764 a_n7677_7899.n65 a_n7677_7899.n26 74.9385
R19765 a_n7677_7899.n127 a_n7677_7899.n64 161.3
R19766 a_n7677_7899.n61 a_n7677_7899.n64 161.3
R19767 a_n7677_7899.n63 a_n7677_7899.n62 71.6402
R19768 a_n7677_7899.n60 a_n7677_7899.n59 68.6201
R19769 a_n7677_7899.n56 a_n7677_7899.n58 74.8341
R19770 a_n7677_7899.n124 a_n7677_7899.n57 161.3
R19771 a_n7677_7899.n57 a_n7677_7899.n123 161.3
R19772 a_n7677_7899.n55 a_n7677_7899.n54 71.8318
R19773 a_n7677_7899.n145 a_n7677_7899.n89 161.3
R19774 a_n7677_7899.n86 a_n7677_7899.n89 161.3
R19775 a_n7677_7899.n88 a_n7677_7899.n87 71.4497
R19776 a_n7677_7899.n85 a_n7677_7899.n84 68.7078
R19777 a_n7677_7899.n28 a_n7677_7899.n27 11.426
R19778 a_n7677_7899.n83 a_n7677_7899.n28 74.9385
R19779 a_n7677_7899.n142 a_n7677_7899.n82 161.3
R19780 a_n7677_7899.n79 a_n7677_7899.n82 161.3
R19781 a_n7677_7899.n81 a_n7677_7899.n80 71.6402
R19782 a_n7677_7899.n78 a_n7677_7899.n77 68.6201
R19783 a_n7677_7899.n74 a_n7677_7899.n76 74.8341
R19784 a_n7677_7899.n139 a_n7677_7899.n75 161.3
R19785 a_n7677_7899.n75 a_n7677_7899.n138 161.3
R19786 a_n7677_7899.n73 a_n7677_7899.n72 71.8318
R19787 a_n7677_7899.n92 a_n7677_7899.n90 109.74
R19788 a_n7677_7899.n95 a_n7677_7899.n93 109.74
R19789 a_n7677_7899.n92 a_n7677_7899.n91 109.166
R19790 a_n7677_7899.n95 a_n7677_7899.n94 109.166
R19791 a_n7677_7899.n97 a_n7677_7899.n96 109.166
R19792 a_n7677_7899.n188 a_n7677_7899.n187 109.166
R19793 a_n7677_7899.n104 a_n7677_7899.n98 84.3502
R19794 a_n7677_7899.n101 a_n7677_7899.n100 84.35
R19795 a_n7677_7899.n101 a_n7677_7899.n99 84.35
R19796 a_n7677_7899.n103 a_n7677_7899.n102 84.0635
R19797 a_n7677_7899.n1 a_n7677_7899.n11 43.6696
R19798 a_n7677_7899.n3 a_n7677_7899.n10 43.6696
R19799 a_n7677_7899.n4 a_n7677_7899.n9 43.6696
R19800 a_n7677_7899.n118 a_n7677_7899.n117 80.6037
R19801 a_n7677_7899.n132 a_n7677_7899.n131 80.6037
R19802 a_n7677_7899.n147 a_n7677_7899.n146 80.6037
R19803 a_n7677_7899.n157 a_n7677_7899.n156 56.5617
R19804 a_n7677_7899.n29 a_n7677_7899.n150 48.4088
R19805 a_n7677_7899.n168 a_n7677_7899.n167 56.5617
R19806 a_n7677_7899.n30 a_n7677_7899.n161 48.4088
R19807 a_n7677_7899.n31 a_n7677_7899.n173 48.4088
R19808 a_n7677_7899.n111 a_n7677_7899.n42 40.5394
R19809 a_n7677_7899.n24 a_n7677_7899.n113 67.9872
R19810 a_n7677_7899.n125 a_n7677_7899.n60 40.5394
R19811 a_n7677_7899.n26 a_n7677_7899.n127 67.9872
R19812 a_n7677_7899.n140 a_n7677_7899.n78 40.5394
R19813 a_n7677_7899.n28 a_n7677_7899.n142 67.9872
R19814 a_n7677_7899.n158 a_n7677_7899.n21 51.9316
R19815 a_n7677_7899.n169 a_n7677_7899.n17 51.9316
R19816 a_n7677_7899.n181 a_n7677_7899.n13 51.9316
R19817 a_n7677_7899.n40 a_n7677_7899.n110 67.7116
R19818 a_n7677_7899.n114 a_n7677_7899.n49 39.872
R19819 a_n7677_7899.n58 a_n7677_7899.n124 67.7116
R19820 a_n7677_7899.n128 a_n7677_7899.n67 39.872
R19821 a_n7677_7899.n76 a_n7677_7899.n139 67.7116
R19822 a_n7677_7899.n143 a_n7677_7899.n85 39.872
R19823 a_n7677_7899.n117 a_n7677_7899.n116 55.824
R19824 a_n7677_7899.n131 a_n7677_7899.n130 55.824
R19825 a_n7677_7899.n146 a_n7677_7899.n145 55.824
R19826 a_n7677_7899.n153 a_n7677_7899.n152 47.1841
R19827 a_n7677_7899.n164 a_n7677_7899.n163 47.1841
R19828 a_n7677_7899.n176 a_n7677_7899.n175 47.1841
R19829 a_n7677_7899.n108 a_n7677_7899.n107 47.1841
R19830 a_n7677_7899.n122 a_n7677_7899.n121 47.1841
R19831 a_n7677_7899.n137 a_n7677_7899.n136 47.1841
R19832 a_n7677_7899.n36 a_n7677_7899.n108 43.9713
R19833 a_n7677_7899.n54 a_n7677_7899.n122 43.9713
R19834 a_n7677_7899.n72 a_n7677_7899.n137 43.9713
R19835 a_n7677_7899.n0 a_n7677_7899.n153 43.9713
R19836 a_n7677_7899.n2 a_n7677_7899.n164 43.9713
R19837 a_n7677_7899.n33 a_n7677_7899.n176 43.9713
R19838 a_n7677_7899.n158 a_n7677_7899.n22 41.2665
R19839 a_n7677_7899.n169 a_n7677_7899.n18 41.2665
R19840 a_n7677_7899.n181 a_n7677_7899.n14 41.2665
R19841 a_n7677_7899.n177 a_n7677_7899.n35 59.1846
R19842 a_n7677_7899.n109 a_n7677_7899.n37 59.1846
R19843 a_n7677_7899.n51 a_n7677_7899.n50 58.0115
R19844 a_n7677_7899.n123 a_n7677_7899.n55 59.1846
R19845 a_n7677_7899.n69 a_n7677_7899.n68 58.0115
R19846 a_n7677_7899.n138 a_n7677_7899.n73 59.1846
R19847 a_n7677_7899.n87 a_n7677_7899.n86 58.0115
R19848 a_n7677_7899.n154 a_n7677_7899.n20 40.5378
R19849 a_n7677_7899.n165 a_n7677_7899.n16 40.5378
R19850 a_n7677_7899.n179 a_n7677_7899.n12 40.5378
R19851 a_n7677_7899.n44 a_n7677_7899.n43 58.5991
R19852 a_n7677_7899.n62 a_n7677_7899.n61 58.5991
R19853 a_n7677_7899.n80 a_n7677_7899.n79 58.5991
R19854 a_n7677_7899.n19 a_n7677_7899.n152 39.8067
R19855 a_n7677_7899.n15 a_n7677_7899.n163 39.8067
R19856 a_n7677_7899.n35 a_n7677_7899.n175 25.2628
R19857 a_n7677_7899.n103 a_n7677_7899.n101 30.5791
R19858 a_n7677_7899.n186 a_n7677_7899.n97 27.4144
R19859 a_n7677_7899.n5 a_n7677_7899.n151 51.931
R19860 a_n7677_7899.n6 a_n7677_7899.n162 51.931
R19861 a_n7677_7899.n32 a_n7677_7899.n178 67.7116
R19862 a_n7677_7899.n105 a_n7677_7899.n40 11.8807
R19863 a_n7677_7899.n49 a_n7677_7899.n23 48.9635
R19864 a_n7677_7899.n119 a_n7677_7899.n58 11.8807
R19865 a_n7677_7899.n67 a_n7677_7899.n25 48.9635
R19866 a_n7677_7899.n134 a_n7677_7899.n76 11.8807
R19867 a_n7677_7899.n85 a_n7677_7899.n27 48.9635
R19868 a_n7677_7899.n157 a_n7677_7899.n149 24.3464
R19869 a_n7677_7899.n168 a_n7677_7899.n160 24.3464
R19870 a_n7677_7899.n8 a_n7677_7899.n172 48.4088
R19871 a_n7677_7899.n42 a_n7677_7899.n105 48.4088
R19872 a_n7677_7899.n60 a_n7677_7899.n119 48.4088
R19873 a_n7677_7899.n78 a_n7677_7899.n134 48.4088
R19874 a_n7677_7899.n187 a_n7677_7899.n186 17.7829
R19875 a_n7677_7899.n11 a_n7677_7899.n159 47.213
R19876 a_n7677_7899.n10 a_n7677_7899.n170 47.213
R19877 a_n7677_7899.n9 a_n7677_7899.n182 47.213
R19878 a_n7677_7899.n116 a_n7677_7899.n115 16.9689
R19879 a_n7677_7899.n130 a_n7677_7899.n129 16.9689
R19880 a_n7677_7899.n145 a_n7677_7899.n144 16.9689
R19881 a_n7677_7899.n156 a_n7677_7899.n155 16.477
R19882 a_n7677_7899.n154 a_n7677_7899.n29 40.5394
R19883 a_n7677_7899.n167 a_n7677_7899.n166 16.477
R19884 a_n7677_7899.n165 a_n7677_7899.n30 40.5394
R19885 a_n7677_7899.n8 a_n7677_7899.n180 40.5394
R19886 a_n7677_7899.n179 a_n7677_7899.n31 40.5394
R19887 a_n7677_7899.n113 a_n7677_7899.n112 16.477
R19888 a_n7677_7899.n127 a_n7677_7899.n126 16.477
R19889 a_n7677_7899.n142 a_n7677_7899.n141 16.477
R19890 a_n7677_7899.n178 a_n7677_7899.n174 15.9852
R19891 a_n7677_7899.n110 a_n7677_7899.n106 15.9852
R19892 a_n7677_7899.n124 a_n7677_7899.n120 15.9852
R19893 a_n7677_7899.n139 a_n7677_7899.n135 15.9852
R19894 a_n7677_7899.n185 a_n7677_7899.n104 12.3349
R19895 a_n7677_7899.n186 a_n7677_7899.n185 11.4887
R19896 a_n7677_7899.n171 a_n7677_7899.n1 8.79829
R19897 a_n7677_7899.n133 a_n7677_7899.n118 8.79829
R19898 a_n7677_7899.n19 a_n7677_7899.n151 41.266
R19899 a_n7677_7899.n15 a_n7677_7899.n162 41.266
R19900 a_n7677_7899.n177 a_n7677_7899.n174 8.60764
R19901 a_n7677_7899.n109 a_n7677_7899.n106 8.60764
R19902 a_n7677_7899.n51 a_n7677_7899.n114 27.0108
R19903 a_n7677_7899.n123 a_n7677_7899.n120 8.60764
R19904 a_n7677_7899.n69 a_n7677_7899.n128 27.0108
R19905 a_n7677_7899.n138 a_n7677_7899.n135 8.60764
R19906 a_n7677_7899.n87 a_n7677_7899.n143 27.0108
R19907 a_n7677_7899.n155 a_n7677_7899.n20 40.5373
R19908 a_n7677_7899.n166 a_n7677_7899.n16 40.5373
R19909 a_n7677_7899.n180 a_n7677_7899.n12 40.5373
R19910 a_n7677_7899.n44 a_n7677_7899.n111 26.1378
R19911 a_n7677_7899.n112 a_n7677_7899.n43 8.11581
R19912 a_n7677_7899.n62 a_n7677_7899.n125 26.1378
R19913 a_n7677_7899.n126 a_n7677_7899.n61 8.11581
R19914 a_n7677_7899.n80 a_n7677_7899.n140 26.1378
R19915 a_n7677_7899.n141 a_n7677_7899.n79 8.11581
R19916 a_n7677_7899.n159 a_n7677_7899.n22 39.8062
R19917 a_n7677_7899.n170 a_n7677_7899.n18 39.8062
R19918 a_n7677_7899.n182 a_n7677_7899.n14 39.8062
R19919 a_n7677_7899.n37 a_n7677_7899.n107 25.2628
R19920 a_n7677_7899.n115 a_n7677_7899.n50 7.62397
R19921 a_n7677_7899.n55 a_n7677_7899.n121 25.2628
R19922 a_n7677_7899.n129 a_n7677_7899.n68 7.62397
R19923 a_n7677_7899.n73 a_n7677_7899.n136 25.2628
R19924 a_n7677_7899.n144 a_n7677_7899.n86 7.62397
R19925 a_n7677_7899.n184 a_n7677_7899.n148 5.76529
R19926 a_n7677_7899.n184 a_n7677_7899.n183 5.56444
R19927 a_n7677_7899.n91 a_n7677_7899.t4 5.418
R19928 a_n7677_7899.n91 a_n7677_7899.t19 5.418
R19929 a_n7677_7899.n90 a_n7677_7899.t5 5.418
R19930 a_n7677_7899.n90 a_n7677_7899.t13 5.418
R19931 a_n7677_7899.n93 a_n7677_7899.t9 5.418
R19932 a_n7677_7899.n93 a_n7677_7899.t10 5.418
R19933 a_n7677_7899.n94 a_n7677_7899.t12 5.418
R19934 a_n7677_7899.n94 a_n7677_7899.t6 5.418
R19935 a_n7677_7899.n96 a_n7677_7899.t11 5.418
R19936 a_n7677_7899.n96 a_n7677_7899.t8 5.418
R19937 a_n7677_7899.n188 a_n7677_7899.t7 5.418
R19938 a_n7677_7899.t0 a_n7677_7899.n188 5.418
R19939 a_n7677_7899.n171 a_n7677_7899.n3 5.06913
R19940 a_n7677_7899.n183 a_n7677_7899.n4 5.06913
R19941 a_n7677_7899.n133 a_n7677_7899.n132 5.06913
R19942 a_n7677_7899.n148 a_n7677_7899.n147 5.06913
R19943 a_n7677_7899.n183 a_n7677_7899.n171 3.72967
R19944 a_n7677_7899.n148 a_n7677_7899.n133 3.72967
R19945 a_n7677_7899.n185 a_n7677_7899.n184 3.4105
R19946 a_n7677_7899.n102 a_n7677_7899.t17 3.3005
R19947 a_n7677_7899.n102 a_n7677_7899.t16 3.3005
R19948 a_n7677_7899.n98 a_n7677_7899.t18 3.3005
R19949 a_n7677_7899.n98 a_n7677_7899.t15 3.3005
R19950 a_n7677_7899.n100 a_n7677_7899.t3 3.3005
R19951 a_n7677_7899.n100 a_n7677_7899.t14 3.3005
R19952 a_n7677_7899.n99 a_n7677_7899.t2 3.3005
R19953 a_n7677_7899.n99 a_n7677_7899.t1 3.3005
R19954 a_n7677_7899.n97 a_n7677_7899.n95 0.573776
R19955 a_n7677_7899.n187 a_n7677_7899.n92 0.573776
R19956 a_n7677_7899.n75 a_n7677_7899.n72 0.568682
R19957 a_n7677_7899.n57 a_n7677_7899.n54 0.568682
R19958 a_n7677_7899.n39 a_n7677_7899.n36 0.568682
R19959 a_n7677_7899.n89 a_n7677_7899.n88 0.379288
R19960 a_n7677_7899.n88 a_n7677_7899.n84 0.379288
R19961 a_n7677_7899.n84 a_n7677_7899.n83 0.379288
R19962 a_n7677_7899.n83 a_n7677_7899.n82 0.379288
R19963 a_n7677_7899.n82 a_n7677_7899.n81 0.379288
R19964 a_n7677_7899.n81 a_n7677_7899.n77 0.379288
R19965 a_n7677_7899.n77 a_n7677_7899.n74 0.379288
R19966 a_n7677_7899.n75 a_n7677_7899.n74 0.379288
R19967 a_n7677_7899.n71 a_n7677_7899.n70 0.379288
R19968 a_n7677_7899.n70 a_n7677_7899.n66 0.379288
R19969 a_n7677_7899.n66 a_n7677_7899.n65 0.379288
R19970 a_n7677_7899.n65 a_n7677_7899.n64 0.379288
R19971 a_n7677_7899.n64 a_n7677_7899.n63 0.379288
R19972 a_n7677_7899.n63 a_n7677_7899.n59 0.379288
R19973 a_n7677_7899.n59 a_n7677_7899.n56 0.379288
R19974 a_n7677_7899.n57 a_n7677_7899.n56 0.379288
R19975 a_n7677_7899.n53 a_n7677_7899.n52 0.379288
R19976 a_n7677_7899.n52 a_n7677_7899.n48 0.379288
R19977 a_n7677_7899.n48 a_n7677_7899.n47 0.379288
R19978 a_n7677_7899.n47 a_n7677_7899.n46 0.379288
R19979 a_n7677_7899.n46 a_n7677_7899.n45 0.379288
R19980 a_n7677_7899.n45 a_n7677_7899.n41 0.379288
R19981 a_n7677_7899.n41 a_n7677_7899.n38 0.379288
R19982 a_n7677_7899.n39 a_n7677_7899.n38 0.379288
R19983 a_n7677_7899.n34 a_n7677_7899.n33 0.379288
R19984 a_n7677_7899.n34 a_n7677_7899.n7 0.379288
R19985 a_n7677_7899.n104 a_n7677_7899.n103 0.287138
R19986 a_n7677_7899.n118 a_n7677_7899.n53 0.285035
R19987 a_n7677_7899.n132 a_n7677_7899.n71 0.285035
R19988 a_n7677_7899.n147 a_n7677_7899.n89 0.285035
R19989 a_n7677_7899.n149 a_n7677_7899.n21 28.5572
R19990 a_n7677_7899.n5 a_n7677_7899.n150 28.5577
R19991 a_n7677_7899.n160 a_n7677_7899.n17 28.5572
R19992 a_n7677_7899.n6 a_n7677_7899.n161 28.5577
R19993 a_n7677_7899.n172 a_n7677_7899.n13 28.5572
R19994 a_n7677_7899.n32 a_n7677_7899.n173 11.8807
R19995 a_n7677_7899.n3 a_n7677_7899.n2 3.88352
R19996 a_n7677_7899.n1 a_n7677_7899.n0 3.88352
R19997 a_n7677_7899.n4 a_n7677_7899.n7 3.12594
R19998 plus.n28 plus.t0 243.97
R19999 plus.n28 plus.n27 223.454
R20000 plus.n30 plus.n29 223.454
R20001 plus.n15 plus.t7 199.144
R20002 plus.n2 plus.t5 199.144
R20003 plus.n24 plus.t10 183.883
R20004 plus.n11 plus.t9 183.883
R20005 plus.n23 plus.n13 161.3
R20006 plus.n21 plus.n20 161.3
R20007 plus.n19 plus.n14 161.3
R20008 plus.n18 plus.n17 161.3
R20009 plus.n5 plus.n4 161.3
R20010 plus.n6 plus.n1 161.3
R20011 plus.n8 plus.n7 161.3
R20012 plus.n10 plus.n0 161.3
R20013 plus.n16 plus.t6 144.601
R20014 plus.n22 plus.t11 144.601
R20015 plus.n9 plus.t8 144.601
R20016 plus.n3 plus.t12 144.601
R20017 plus.n25 plus.n24 80.6037
R20018 plus.n12 plus.n11 80.6037
R20019 plus.n24 plus.n23 56.3158
R20020 plus.n11 plus.n10 56.3158
R20021 plus.n16 plus.n15 46.9082
R20022 plus.n3 plus.n2 46.9082
R20023 plus.n18 plus.n15 43.8991
R20024 plus.n5 plus.n2 43.8991
R20025 plus.n17 plus.n14 40.577
R20026 plus.n21 plus.n14 40.577
R20027 plus.n8 plus.n1 40.577
R20028 plus.n4 plus.n1 40.577
R20029 plus.n26 plus.n25 27.893
R20030 plus.n27 plus.t1 19.8005
R20031 plus.n27 plus.t4 19.8005
R20032 plus.n29 plus.t2 19.8005
R20033 plus.n29 plus.t3 19.8005
R20034 plus.n23 plus.n22 16.477
R20035 plus.n10 plus.n9 16.477
R20036 plus plus.n31 13.8471
R20037 plus.n26 plus.n12 11.6998
R20038 plus.n17 plus.n16 8.11581
R20039 plus.n22 plus.n21 8.11581
R20040 plus.n9 plus.n8 8.11581
R20041 plus.n4 plus.n3 8.11581
R20042 plus.n31 plus.n30 5.40567
R20043 plus.n31 plus.n26 1.188
R20044 plus.n30 plus.n28 0.716017
R20045 plus.n25 plus.n13 0.285035
R20046 plus.n12 plus.n0 0.285035
R20047 plus.n19 plus.n18 0.189894
R20048 plus.n20 plus.n19 0.189894
R20049 plus.n20 plus.n13 0.189894
R20050 plus.n7 plus.n0 0.189894
R20051 plus.n7 plus.n6 0.189894
R20052 plus.n6 plus.n5 0.189894
R20053 a_n1455_n3628.n308 a_n1455_n3628.n288 289.615
R20054 a_n1455_n3628.n335 a_n1455_n3628.n315 289.615
R20055 a_n1455_n3628.n177 a_n1455_n3628.n157 289.615
R20056 a_n1455_n3628.n281 a_n1455_n3628.n261 289.615
R20057 a_n1455_n3628.n255 a_n1455_n3628.n235 289.615
R20058 a_n1455_n3628.n229 a_n1455_n3628.n209 289.615
R20059 a_n1455_n3628.n203 a_n1455_n3628.n183 289.615
R20060 a_n1455_n3628.n69 a_n1455_n3628.n49 289.615
R20061 a_n1455_n3628.n97 a_n1455_n3628.n77 289.615
R20062 a_n1455_n3628.n123 a_n1455_n3628.n103 289.615
R20063 a_n1455_n3628.n151 a_n1455_n3628.n131 289.615
R20064 a_n1455_n3628.n344 a_n1455_n3628.n46 289.615
R20065 a_n1455_n3628.n208 a_n1455_n3628.n207 196.838
R20066 a_n1455_n3628.n286 a_n1455_n3628.n285 196.298
R20067 a_n1455_n3628.n260 a_n1455_n3628.n259 196.298
R20068 a_n1455_n3628.n234 a_n1455_n3628.n233 196.298
R20069 a_n1455_n3628.n297 a_n1455_n3628.n296 185
R20070 a_n1455_n3628.n294 a_n1455_n3628.n293 185
R20071 a_n1455_n3628.n301 a_n1455_n3628.n300 185
R20072 a_n1455_n3628.n303 a_n1455_n3628.n302 185
R20073 a_n1455_n3628.n291 a_n1455_n3628.n290 185
R20074 a_n1455_n3628.n307 a_n1455_n3628.n306 185
R20075 a_n1455_n3628.n309 a_n1455_n3628.n308 185
R20076 a_n1455_n3628.n324 a_n1455_n3628.n323 185
R20077 a_n1455_n3628.n321 a_n1455_n3628.n320 185
R20078 a_n1455_n3628.n328 a_n1455_n3628.n327 185
R20079 a_n1455_n3628.n330 a_n1455_n3628.n329 185
R20080 a_n1455_n3628.n318 a_n1455_n3628.n317 185
R20081 a_n1455_n3628.n334 a_n1455_n3628.n333 185
R20082 a_n1455_n3628.n336 a_n1455_n3628.n335 185
R20083 a_n1455_n3628.n166 a_n1455_n3628.n165 185
R20084 a_n1455_n3628.n163 a_n1455_n3628.n162 185
R20085 a_n1455_n3628.n170 a_n1455_n3628.n169 185
R20086 a_n1455_n3628.n172 a_n1455_n3628.n171 185
R20087 a_n1455_n3628.n160 a_n1455_n3628.n159 185
R20088 a_n1455_n3628.n176 a_n1455_n3628.n175 185
R20089 a_n1455_n3628.n178 a_n1455_n3628.n177 185
R20090 a_n1455_n3628.n282 a_n1455_n3628.n281 185
R20091 a_n1455_n3628.n280 a_n1455_n3628.n279 185
R20092 a_n1455_n3628.n264 a_n1455_n3628.n263 185
R20093 a_n1455_n3628.n276 a_n1455_n3628.n275 185
R20094 a_n1455_n3628.n274 a_n1455_n3628.n273 185
R20095 a_n1455_n3628.n267 a_n1455_n3628.n266 185
R20096 a_n1455_n3628.n270 a_n1455_n3628.n269 185
R20097 a_n1455_n3628.n256 a_n1455_n3628.n255 185
R20098 a_n1455_n3628.n254 a_n1455_n3628.n253 185
R20099 a_n1455_n3628.n238 a_n1455_n3628.n237 185
R20100 a_n1455_n3628.n250 a_n1455_n3628.n249 185
R20101 a_n1455_n3628.n248 a_n1455_n3628.n247 185
R20102 a_n1455_n3628.n241 a_n1455_n3628.n240 185
R20103 a_n1455_n3628.n244 a_n1455_n3628.n243 185
R20104 a_n1455_n3628.n230 a_n1455_n3628.n229 185
R20105 a_n1455_n3628.n228 a_n1455_n3628.n227 185
R20106 a_n1455_n3628.n212 a_n1455_n3628.n211 185
R20107 a_n1455_n3628.n224 a_n1455_n3628.n223 185
R20108 a_n1455_n3628.n222 a_n1455_n3628.n221 185
R20109 a_n1455_n3628.n215 a_n1455_n3628.n214 185
R20110 a_n1455_n3628.n218 a_n1455_n3628.n217 185
R20111 a_n1455_n3628.n204 a_n1455_n3628.n203 185
R20112 a_n1455_n3628.n202 a_n1455_n3628.n201 185
R20113 a_n1455_n3628.n186 a_n1455_n3628.n185 185
R20114 a_n1455_n3628.n198 a_n1455_n3628.n197 185
R20115 a_n1455_n3628.n196 a_n1455_n3628.n195 185
R20116 a_n1455_n3628.n189 a_n1455_n3628.n188 185
R20117 a_n1455_n3628.n192 a_n1455_n3628.n191 185
R20118 a_n1455_n3628.n70 a_n1455_n3628.n69 185
R20119 a_n1455_n3628.n68 a_n1455_n3628.n67 185
R20120 a_n1455_n3628.n52 a_n1455_n3628.n51 185
R20121 a_n1455_n3628.n64 a_n1455_n3628.n63 185
R20122 a_n1455_n3628.n62 a_n1455_n3628.n61 185
R20123 a_n1455_n3628.n55 a_n1455_n3628.n54 185
R20124 a_n1455_n3628.n58 a_n1455_n3628.n57 185
R20125 a_n1455_n3628.n98 a_n1455_n3628.n97 185
R20126 a_n1455_n3628.n96 a_n1455_n3628.n95 185
R20127 a_n1455_n3628.n80 a_n1455_n3628.n79 185
R20128 a_n1455_n3628.n92 a_n1455_n3628.n91 185
R20129 a_n1455_n3628.n90 a_n1455_n3628.n89 185
R20130 a_n1455_n3628.n83 a_n1455_n3628.n82 185
R20131 a_n1455_n3628.n86 a_n1455_n3628.n85 185
R20132 a_n1455_n3628.n124 a_n1455_n3628.n123 185
R20133 a_n1455_n3628.n122 a_n1455_n3628.n121 185
R20134 a_n1455_n3628.n106 a_n1455_n3628.n105 185
R20135 a_n1455_n3628.n118 a_n1455_n3628.n117 185
R20136 a_n1455_n3628.n116 a_n1455_n3628.n115 185
R20137 a_n1455_n3628.n109 a_n1455_n3628.n108 185
R20138 a_n1455_n3628.n112 a_n1455_n3628.n111 185
R20139 a_n1455_n3628.n152 a_n1455_n3628.n151 185
R20140 a_n1455_n3628.n150 a_n1455_n3628.n149 185
R20141 a_n1455_n3628.n134 a_n1455_n3628.n133 185
R20142 a_n1455_n3628.n146 a_n1455_n3628.n145 185
R20143 a_n1455_n3628.n144 a_n1455_n3628.n143 185
R20144 a_n1455_n3628.n137 a_n1455_n3628.n136 185
R20145 a_n1455_n3628.n140 a_n1455_n3628.n139 185
R20146 a_n1455_n3628.n357 a_n1455_n3628.n356 185
R20147 a_n1455_n3628.n41 a_n1455_n3628.n40 185
R20148 a_n1455_n3628.n352 a_n1455_n3628.n351 185
R20149 a_n1455_n3628.n350 a_n1455_n3628.n349 185
R20150 a_n1455_n3628.n44 a_n1455_n3628.n43 185
R20151 a_n1455_n3628.n346 a_n1455_n3628.n345 185
R20152 a_n1455_n3628.n344 a_n1455_n3628.n343 185
R20153 a_n1455_n3628.t19 a_n1455_n3628.n295 147.661
R20154 a_n1455_n3628.t18 a_n1455_n3628.n322 147.661
R20155 a_n1455_n3628.t9 a_n1455_n3628.n164 147.661
R20156 a_n1455_n3628.t1 a_n1455_n3628.n268 147.661
R20157 a_n1455_n3628.t14 a_n1455_n3628.n242 147.661
R20158 a_n1455_n3628.t2 a_n1455_n3628.n216 147.661
R20159 a_n1455_n3628.t0 a_n1455_n3628.n190 147.661
R20160 a_n1455_n3628.t8 a_n1455_n3628.n56 147.661
R20161 a_n1455_n3628.t11 a_n1455_n3628.n84 147.661
R20162 a_n1455_n3628.t15 a_n1455_n3628.n110 147.661
R20163 a_n1455_n3628.t16 a_n1455_n3628.n138 147.661
R20164 a_n1455_n3628.t13 a_n1455_n3628.n39 147.661
R20165 a_n1455_n3628.n296 a_n1455_n3628.n293 104.615
R20166 a_n1455_n3628.n301 a_n1455_n3628.n293 104.615
R20167 a_n1455_n3628.n302 a_n1455_n3628.n301 104.615
R20168 a_n1455_n3628.n302 a_n1455_n3628.n290 104.615
R20169 a_n1455_n3628.n307 a_n1455_n3628.n290 104.615
R20170 a_n1455_n3628.n308 a_n1455_n3628.n307 104.615
R20171 a_n1455_n3628.n323 a_n1455_n3628.n320 104.615
R20172 a_n1455_n3628.n328 a_n1455_n3628.n320 104.615
R20173 a_n1455_n3628.n329 a_n1455_n3628.n328 104.615
R20174 a_n1455_n3628.n329 a_n1455_n3628.n317 104.615
R20175 a_n1455_n3628.n334 a_n1455_n3628.n317 104.615
R20176 a_n1455_n3628.n335 a_n1455_n3628.n334 104.615
R20177 a_n1455_n3628.n165 a_n1455_n3628.n162 104.615
R20178 a_n1455_n3628.n170 a_n1455_n3628.n162 104.615
R20179 a_n1455_n3628.n171 a_n1455_n3628.n170 104.615
R20180 a_n1455_n3628.n171 a_n1455_n3628.n159 104.615
R20181 a_n1455_n3628.n176 a_n1455_n3628.n159 104.615
R20182 a_n1455_n3628.n177 a_n1455_n3628.n176 104.615
R20183 a_n1455_n3628.n281 a_n1455_n3628.n280 104.615
R20184 a_n1455_n3628.n280 a_n1455_n3628.n263 104.615
R20185 a_n1455_n3628.n275 a_n1455_n3628.n263 104.615
R20186 a_n1455_n3628.n275 a_n1455_n3628.n274 104.615
R20187 a_n1455_n3628.n274 a_n1455_n3628.n266 104.615
R20188 a_n1455_n3628.n269 a_n1455_n3628.n266 104.615
R20189 a_n1455_n3628.n255 a_n1455_n3628.n254 104.615
R20190 a_n1455_n3628.n254 a_n1455_n3628.n237 104.615
R20191 a_n1455_n3628.n249 a_n1455_n3628.n237 104.615
R20192 a_n1455_n3628.n249 a_n1455_n3628.n248 104.615
R20193 a_n1455_n3628.n248 a_n1455_n3628.n240 104.615
R20194 a_n1455_n3628.n243 a_n1455_n3628.n240 104.615
R20195 a_n1455_n3628.n229 a_n1455_n3628.n228 104.615
R20196 a_n1455_n3628.n228 a_n1455_n3628.n211 104.615
R20197 a_n1455_n3628.n223 a_n1455_n3628.n211 104.615
R20198 a_n1455_n3628.n223 a_n1455_n3628.n222 104.615
R20199 a_n1455_n3628.n222 a_n1455_n3628.n214 104.615
R20200 a_n1455_n3628.n217 a_n1455_n3628.n214 104.615
R20201 a_n1455_n3628.n203 a_n1455_n3628.n202 104.615
R20202 a_n1455_n3628.n202 a_n1455_n3628.n185 104.615
R20203 a_n1455_n3628.n197 a_n1455_n3628.n185 104.615
R20204 a_n1455_n3628.n197 a_n1455_n3628.n196 104.615
R20205 a_n1455_n3628.n196 a_n1455_n3628.n188 104.615
R20206 a_n1455_n3628.n191 a_n1455_n3628.n188 104.615
R20207 a_n1455_n3628.n69 a_n1455_n3628.n68 104.615
R20208 a_n1455_n3628.n68 a_n1455_n3628.n51 104.615
R20209 a_n1455_n3628.n63 a_n1455_n3628.n51 104.615
R20210 a_n1455_n3628.n63 a_n1455_n3628.n62 104.615
R20211 a_n1455_n3628.n62 a_n1455_n3628.n54 104.615
R20212 a_n1455_n3628.n57 a_n1455_n3628.n54 104.615
R20213 a_n1455_n3628.n97 a_n1455_n3628.n96 104.615
R20214 a_n1455_n3628.n96 a_n1455_n3628.n79 104.615
R20215 a_n1455_n3628.n91 a_n1455_n3628.n79 104.615
R20216 a_n1455_n3628.n91 a_n1455_n3628.n90 104.615
R20217 a_n1455_n3628.n90 a_n1455_n3628.n82 104.615
R20218 a_n1455_n3628.n85 a_n1455_n3628.n82 104.615
R20219 a_n1455_n3628.n123 a_n1455_n3628.n122 104.615
R20220 a_n1455_n3628.n122 a_n1455_n3628.n105 104.615
R20221 a_n1455_n3628.n117 a_n1455_n3628.n105 104.615
R20222 a_n1455_n3628.n117 a_n1455_n3628.n116 104.615
R20223 a_n1455_n3628.n116 a_n1455_n3628.n108 104.615
R20224 a_n1455_n3628.n111 a_n1455_n3628.n108 104.615
R20225 a_n1455_n3628.n151 a_n1455_n3628.n150 104.615
R20226 a_n1455_n3628.n150 a_n1455_n3628.n133 104.615
R20227 a_n1455_n3628.n145 a_n1455_n3628.n133 104.615
R20228 a_n1455_n3628.n145 a_n1455_n3628.n144 104.615
R20229 a_n1455_n3628.n144 a_n1455_n3628.n136 104.615
R20230 a_n1455_n3628.n139 a_n1455_n3628.n136 104.615
R20231 a_n1455_n3628.n357 a_n1455_n3628.n40 104.615
R20232 a_n1455_n3628.n351 a_n1455_n3628.n40 104.615
R20233 a_n1455_n3628.n351 a_n1455_n3628.n350 104.615
R20234 a_n1455_n3628.n350 a_n1455_n3628.n43 104.615
R20235 a_n1455_n3628.n345 a_n1455_n3628.n43 104.615
R20236 a_n1455_n3628.n345 a_n1455_n3628.n344 104.615
R20237 a_n1455_n3628.n76 a_n1455_n3628.n75 56.1363
R20238 a_n1455_n3628.n130 a_n1455_n3628.n129 56.1363
R20239 a_n1455_n3628.n314 a_n1455_n3628.n313 56.1361
R20240 a_n1455_n3628.n48 a_n1455_n3628.n47 56.1361
R20241 a_n1455_n3628.n296 a_n1455_n3628.t19 52.3082
R20242 a_n1455_n3628.n323 a_n1455_n3628.t18 52.3082
R20243 a_n1455_n3628.n165 a_n1455_n3628.t9 52.3082
R20244 a_n1455_n3628.n269 a_n1455_n3628.t1 52.3082
R20245 a_n1455_n3628.n243 a_n1455_n3628.t14 52.3082
R20246 a_n1455_n3628.n217 a_n1455_n3628.t2 52.3082
R20247 a_n1455_n3628.n191 a_n1455_n3628.t0 52.3082
R20248 a_n1455_n3628.n57 a_n1455_n3628.t8 52.3082
R20249 a_n1455_n3628.n85 a_n1455_n3628.t11 52.3082
R20250 a_n1455_n3628.n111 a_n1455_n3628.t15 52.3082
R20251 a_n1455_n3628.n139 a_n1455_n3628.t16 52.3082
R20252 a_n1455_n3628.t13 a_n1455_n3628.n357 52.3082
R20253 a_n1455_n3628.n312 a_n1455_n3628.n311 37.8096
R20254 a_n1455_n3628.n339 a_n1455_n3628.n338 37.8096
R20255 a_n1455_n3628.n181 a_n1455_n3628.n180 37.8096
R20256 a_n1455_n3628.n74 a_n1455_n3628.n73 37.8096
R20257 a_n1455_n3628.n102 a_n1455_n3628.n101 37.8096
R20258 a_n1455_n3628.n128 a_n1455_n3628.n127 37.8096
R20259 a_n1455_n3628.n156 a_n1455_n3628.n155 37.8096
R20260 a_n1455_n3628.n341 a_n1455_n3628.n340 37.8096
R20261 a_n1455_n3628.n297 a_n1455_n3628.n295 15.6674
R20262 a_n1455_n3628.n324 a_n1455_n3628.n322 15.6674
R20263 a_n1455_n3628.n166 a_n1455_n3628.n164 15.6674
R20264 a_n1455_n3628.n270 a_n1455_n3628.n268 15.6674
R20265 a_n1455_n3628.n244 a_n1455_n3628.n242 15.6674
R20266 a_n1455_n3628.n218 a_n1455_n3628.n216 15.6674
R20267 a_n1455_n3628.n192 a_n1455_n3628.n190 15.6674
R20268 a_n1455_n3628.n58 a_n1455_n3628.n56 15.6674
R20269 a_n1455_n3628.n86 a_n1455_n3628.n84 15.6674
R20270 a_n1455_n3628.n112 a_n1455_n3628.n110 15.6674
R20271 a_n1455_n3628.n140 a_n1455_n3628.n138 15.6674
R20272 a_n1455_n3628.n356 a_n1455_n3628.n39 15.6674
R20273 a_n1455_n3628.n298 a_n1455_n3628.n294 12.8005
R20274 a_n1455_n3628.n325 a_n1455_n3628.n321 12.8005
R20275 a_n1455_n3628.n167 a_n1455_n3628.n163 12.8005
R20276 a_n1455_n3628.n271 a_n1455_n3628.n267 12.8005
R20277 a_n1455_n3628.n245 a_n1455_n3628.n241 12.8005
R20278 a_n1455_n3628.n219 a_n1455_n3628.n215 12.8005
R20279 a_n1455_n3628.n193 a_n1455_n3628.n189 12.8005
R20280 a_n1455_n3628.n59 a_n1455_n3628.n55 12.8005
R20281 a_n1455_n3628.n87 a_n1455_n3628.n83 12.8005
R20282 a_n1455_n3628.n113 a_n1455_n3628.n109 12.8005
R20283 a_n1455_n3628.n141 a_n1455_n3628.n137 12.8005
R20284 a_n1455_n3628.n355 a_n1455_n3628.n41 12.8005
R20285 a_n1455_n3628.n300 a_n1455_n3628.n299 12.0247
R20286 a_n1455_n3628.n327 a_n1455_n3628.n326 12.0247
R20287 a_n1455_n3628.n169 a_n1455_n3628.n168 12.0247
R20288 a_n1455_n3628.n273 a_n1455_n3628.n272 12.0247
R20289 a_n1455_n3628.n247 a_n1455_n3628.n246 12.0247
R20290 a_n1455_n3628.n221 a_n1455_n3628.n220 12.0247
R20291 a_n1455_n3628.n195 a_n1455_n3628.n194 12.0247
R20292 a_n1455_n3628.n61 a_n1455_n3628.n60 12.0247
R20293 a_n1455_n3628.n89 a_n1455_n3628.n88 12.0247
R20294 a_n1455_n3628.n115 a_n1455_n3628.n114 12.0247
R20295 a_n1455_n3628.n143 a_n1455_n3628.n142 12.0247
R20296 a_n1455_n3628.n353 a_n1455_n3628.n352 12.0247
R20297 a_n1455_n3628.n182 a_n1455_n3628.n156 11.5057
R20298 a_n1455_n3628.n287 a_n1455_n3628.n74 11.5057
R20299 a_n1455_n3628.n303 a_n1455_n3628.n292 11.249
R20300 a_n1455_n3628.n330 a_n1455_n3628.n319 11.249
R20301 a_n1455_n3628.n172 a_n1455_n3628.n161 11.249
R20302 a_n1455_n3628.n276 a_n1455_n3628.n265 11.249
R20303 a_n1455_n3628.n250 a_n1455_n3628.n239 11.249
R20304 a_n1455_n3628.n224 a_n1455_n3628.n213 11.249
R20305 a_n1455_n3628.n198 a_n1455_n3628.n187 11.249
R20306 a_n1455_n3628.n64 a_n1455_n3628.n53 11.249
R20307 a_n1455_n3628.n92 a_n1455_n3628.n81 11.249
R20308 a_n1455_n3628.n118 a_n1455_n3628.n107 11.249
R20309 a_n1455_n3628.n146 a_n1455_n3628.n135 11.249
R20310 a_n1455_n3628.n349 a_n1455_n3628.n42 11.249
R20311 a_n1455_n3628.n304 a_n1455_n3628.n291 10.4732
R20312 a_n1455_n3628.n331 a_n1455_n3628.n318 10.4732
R20313 a_n1455_n3628.n173 a_n1455_n3628.n160 10.4732
R20314 a_n1455_n3628.n277 a_n1455_n3628.n264 10.4732
R20315 a_n1455_n3628.n251 a_n1455_n3628.n238 10.4732
R20316 a_n1455_n3628.n225 a_n1455_n3628.n212 10.4732
R20317 a_n1455_n3628.n199 a_n1455_n3628.n186 10.4732
R20318 a_n1455_n3628.n65 a_n1455_n3628.n52 10.4732
R20319 a_n1455_n3628.n93 a_n1455_n3628.n80 10.4732
R20320 a_n1455_n3628.n119 a_n1455_n3628.n106 10.4732
R20321 a_n1455_n3628.n147 a_n1455_n3628.n134 10.4732
R20322 a_n1455_n3628.n348 a_n1455_n3628.n44 10.4732
R20323 a_n1455_n3628.n306 a_n1455_n3628.n305 9.69747
R20324 a_n1455_n3628.n333 a_n1455_n3628.n332 9.69747
R20325 a_n1455_n3628.n175 a_n1455_n3628.n174 9.69747
R20326 a_n1455_n3628.n279 a_n1455_n3628.n278 9.69747
R20327 a_n1455_n3628.n253 a_n1455_n3628.n252 9.69747
R20328 a_n1455_n3628.n227 a_n1455_n3628.n226 9.69747
R20329 a_n1455_n3628.n201 a_n1455_n3628.n200 9.69747
R20330 a_n1455_n3628.n67 a_n1455_n3628.n66 9.69747
R20331 a_n1455_n3628.n95 a_n1455_n3628.n94 9.69747
R20332 a_n1455_n3628.n121 a_n1455_n3628.n120 9.69747
R20333 a_n1455_n3628.n149 a_n1455_n3628.n148 9.69747
R20334 a_n1455_n3628.n347 a_n1455_n3628.n346 9.69747
R20335 a_n1455_n3628.n1 a_n1455_n3628.n341 9.45567
R20336 a_n1455_n3628.n311 a_n1455_n3628.n5 9.45567
R20337 a_n1455_n3628.n338 a_n1455_n3628.n9 9.45567
R20338 a_n1455_n3628.n180 a_n1455_n3628.n13 9.45567
R20339 a_n1455_n3628.n285 a_n1455_n3628.n284 9.45567
R20340 a_n1455_n3628.n259 a_n1455_n3628.n258 9.45567
R20341 a_n1455_n3628.n233 a_n1455_n3628.n232 9.45567
R20342 a_n1455_n3628.n207 a_n1455_n3628.n206 9.45567
R20343 a_n1455_n3628.n73 a_n1455_n3628.n72 9.45567
R20344 a_n1455_n3628.n101 a_n1455_n3628.n100 9.45567
R20345 a_n1455_n3628.n127 a_n1455_n3628.n126 9.45567
R20346 a_n1455_n3628.n155 a_n1455_n3628.n154 9.45567
R20347 a_n1455_n3628.n5 a_n1455_n3628.n310 9.3005
R20348 a_n1455_n3628.n289 a_n1455_n3628.n5 9.3005
R20349 a_n1455_n3628.n305 a_n1455_n3628.n6 9.3005
R20350 a_n1455_n3628.n6 a_n1455_n3628.n304 9.3005
R20351 a_n1455_n3628.n292 a_n1455_n3628.n4 9.3005
R20352 a_n1455_n3628.n299 a_n1455_n3628.n4 9.3005
R20353 a_n1455_n3628.n3 a_n1455_n3628.n298 9.3005
R20354 a_n1455_n3628.n9 a_n1455_n3628.n337 9.3005
R20355 a_n1455_n3628.n316 a_n1455_n3628.n9 9.3005
R20356 a_n1455_n3628.n332 a_n1455_n3628.n10 9.3005
R20357 a_n1455_n3628.n10 a_n1455_n3628.n331 9.3005
R20358 a_n1455_n3628.n319 a_n1455_n3628.n8 9.3005
R20359 a_n1455_n3628.n326 a_n1455_n3628.n8 9.3005
R20360 a_n1455_n3628.n7 a_n1455_n3628.n325 9.3005
R20361 a_n1455_n3628.n13 a_n1455_n3628.n179 9.3005
R20362 a_n1455_n3628.n158 a_n1455_n3628.n13 9.3005
R20363 a_n1455_n3628.n174 a_n1455_n3628.n14 9.3005
R20364 a_n1455_n3628.n14 a_n1455_n3628.n173 9.3005
R20365 a_n1455_n3628.n161 a_n1455_n3628.n12 9.3005
R20366 a_n1455_n3628.n168 a_n1455_n3628.n12 9.3005
R20367 a_n1455_n3628.n11 a_n1455_n3628.n167 9.3005
R20368 a_n1455_n3628.n284 a_n1455_n3628.n283 9.3005
R20369 a_n1455_n3628.n262 a_n1455_n3628.n16 9.3005
R20370 a_n1455_n3628.n278 a_n1455_n3628.n16 9.3005
R20371 a_n1455_n3628.n15 a_n1455_n3628.n277 9.3005
R20372 a_n1455_n3628.n265 a_n1455_n3628.n15 9.3005
R20373 a_n1455_n3628.n272 a_n1455_n3628.n17 9.3005
R20374 a_n1455_n3628.n17 a_n1455_n3628.n271 9.3005
R20375 a_n1455_n3628.n258 a_n1455_n3628.n257 9.3005
R20376 a_n1455_n3628.n236 a_n1455_n3628.n19 9.3005
R20377 a_n1455_n3628.n252 a_n1455_n3628.n19 9.3005
R20378 a_n1455_n3628.n18 a_n1455_n3628.n251 9.3005
R20379 a_n1455_n3628.n239 a_n1455_n3628.n18 9.3005
R20380 a_n1455_n3628.n246 a_n1455_n3628.n20 9.3005
R20381 a_n1455_n3628.n20 a_n1455_n3628.n245 9.3005
R20382 a_n1455_n3628.n232 a_n1455_n3628.n231 9.3005
R20383 a_n1455_n3628.n210 a_n1455_n3628.n22 9.3005
R20384 a_n1455_n3628.n226 a_n1455_n3628.n22 9.3005
R20385 a_n1455_n3628.n21 a_n1455_n3628.n225 9.3005
R20386 a_n1455_n3628.n213 a_n1455_n3628.n21 9.3005
R20387 a_n1455_n3628.n220 a_n1455_n3628.n23 9.3005
R20388 a_n1455_n3628.n23 a_n1455_n3628.n219 9.3005
R20389 a_n1455_n3628.n206 a_n1455_n3628.n205 9.3005
R20390 a_n1455_n3628.n184 a_n1455_n3628.n25 9.3005
R20391 a_n1455_n3628.n200 a_n1455_n3628.n25 9.3005
R20392 a_n1455_n3628.n24 a_n1455_n3628.n199 9.3005
R20393 a_n1455_n3628.n187 a_n1455_n3628.n24 9.3005
R20394 a_n1455_n3628.n194 a_n1455_n3628.n26 9.3005
R20395 a_n1455_n3628.n26 a_n1455_n3628.n193 9.3005
R20396 a_n1455_n3628.n72 a_n1455_n3628.n71 9.3005
R20397 a_n1455_n3628.n50 a_n1455_n3628.n28 9.3005
R20398 a_n1455_n3628.n66 a_n1455_n3628.n28 9.3005
R20399 a_n1455_n3628.n27 a_n1455_n3628.n65 9.3005
R20400 a_n1455_n3628.n53 a_n1455_n3628.n27 9.3005
R20401 a_n1455_n3628.n60 a_n1455_n3628.n29 9.3005
R20402 a_n1455_n3628.n29 a_n1455_n3628.n59 9.3005
R20403 a_n1455_n3628.n100 a_n1455_n3628.n99 9.3005
R20404 a_n1455_n3628.n78 a_n1455_n3628.n31 9.3005
R20405 a_n1455_n3628.n94 a_n1455_n3628.n31 9.3005
R20406 a_n1455_n3628.n30 a_n1455_n3628.n93 9.3005
R20407 a_n1455_n3628.n81 a_n1455_n3628.n30 9.3005
R20408 a_n1455_n3628.n88 a_n1455_n3628.n32 9.3005
R20409 a_n1455_n3628.n32 a_n1455_n3628.n87 9.3005
R20410 a_n1455_n3628.n126 a_n1455_n3628.n125 9.3005
R20411 a_n1455_n3628.n104 a_n1455_n3628.n34 9.3005
R20412 a_n1455_n3628.n120 a_n1455_n3628.n34 9.3005
R20413 a_n1455_n3628.n33 a_n1455_n3628.n119 9.3005
R20414 a_n1455_n3628.n107 a_n1455_n3628.n33 9.3005
R20415 a_n1455_n3628.n114 a_n1455_n3628.n35 9.3005
R20416 a_n1455_n3628.n35 a_n1455_n3628.n113 9.3005
R20417 a_n1455_n3628.n154 a_n1455_n3628.n153 9.3005
R20418 a_n1455_n3628.n132 a_n1455_n3628.n37 9.3005
R20419 a_n1455_n3628.n148 a_n1455_n3628.n37 9.3005
R20420 a_n1455_n3628.n36 a_n1455_n3628.n147 9.3005
R20421 a_n1455_n3628.n135 a_n1455_n3628.n36 9.3005
R20422 a_n1455_n3628.n142 a_n1455_n3628.n38 9.3005
R20423 a_n1455_n3628.n38 a_n1455_n3628.n141 9.3005
R20424 a_n1455_n3628.n342 a_n1455_n3628.n1 9.3005
R20425 a_n1455_n3628.n45 a_n1455_n3628.n1 9.3005
R20426 a_n1455_n3628.n2 a_n1455_n3628.n347 9.3005
R20427 a_n1455_n3628.n348 a_n1455_n3628.n2 9.3005
R20428 a_n1455_n3628.n42 a_n1455_n3628.n0 9.3005
R20429 a_n1455_n3628.n0 a_n1455_n3628.n353 9.3005
R20430 a_n1455_n3628.n355 a_n1455_n3628.n354 9.3005
R20431 a_n1455_n3628.n309 a_n1455_n3628.n289 8.92171
R20432 a_n1455_n3628.n336 a_n1455_n3628.n316 8.92171
R20433 a_n1455_n3628.n178 a_n1455_n3628.n158 8.92171
R20434 a_n1455_n3628.n282 a_n1455_n3628.n262 8.92171
R20435 a_n1455_n3628.n256 a_n1455_n3628.n236 8.92171
R20436 a_n1455_n3628.n230 a_n1455_n3628.n210 8.92171
R20437 a_n1455_n3628.n204 a_n1455_n3628.n184 8.92171
R20438 a_n1455_n3628.n70 a_n1455_n3628.n50 8.92171
R20439 a_n1455_n3628.n98 a_n1455_n3628.n78 8.92171
R20440 a_n1455_n3628.n124 a_n1455_n3628.n104 8.92171
R20441 a_n1455_n3628.n152 a_n1455_n3628.n132 8.92171
R20442 a_n1455_n3628.n343 a_n1455_n3628.n45 8.92171
R20443 a_n1455_n3628.n310 a_n1455_n3628.n288 8.14595
R20444 a_n1455_n3628.n337 a_n1455_n3628.n315 8.14595
R20445 a_n1455_n3628.n179 a_n1455_n3628.n157 8.14595
R20446 a_n1455_n3628.n283 a_n1455_n3628.n261 8.14595
R20447 a_n1455_n3628.n257 a_n1455_n3628.n235 8.14595
R20448 a_n1455_n3628.n231 a_n1455_n3628.n209 8.14595
R20449 a_n1455_n3628.n205 a_n1455_n3628.n183 8.14595
R20450 a_n1455_n3628.n71 a_n1455_n3628.n49 8.14595
R20451 a_n1455_n3628.n99 a_n1455_n3628.n77 8.14595
R20452 a_n1455_n3628.n125 a_n1455_n3628.n103 8.14595
R20453 a_n1455_n3628.n153 a_n1455_n3628.n131 8.14595
R20454 a_n1455_n3628.n342 a_n1455_n3628.n46 8.14595
R20455 a_n1455_n3628.n311 a_n1455_n3628.n288 5.81868
R20456 a_n1455_n3628.n338 a_n1455_n3628.n315 5.81868
R20457 a_n1455_n3628.n180 a_n1455_n3628.n157 5.81868
R20458 a_n1455_n3628.n285 a_n1455_n3628.n261 5.81868
R20459 a_n1455_n3628.n259 a_n1455_n3628.n235 5.81868
R20460 a_n1455_n3628.n233 a_n1455_n3628.n209 5.81868
R20461 a_n1455_n3628.n207 a_n1455_n3628.n183 5.81868
R20462 a_n1455_n3628.n73 a_n1455_n3628.n49 5.81868
R20463 a_n1455_n3628.n101 a_n1455_n3628.n77 5.81868
R20464 a_n1455_n3628.n127 a_n1455_n3628.n103 5.81868
R20465 a_n1455_n3628.n155 a_n1455_n3628.n131 5.81868
R20466 a_n1455_n3628.n341 a_n1455_n3628.n46 5.81868
R20467 a_n1455_n3628.n182 a_n1455_n3628.n181 5.18369
R20468 a_n1455_n3628.n312 a_n1455_n3628.n287 5.18369
R20469 a_n1455_n3628.n310 a_n1455_n3628.n309 5.04292
R20470 a_n1455_n3628.n337 a_n1455_n3628.n336 5.04292
R20471 a_n1455_n3628.n179 a_n1455_n3628.n178 5.04292
R20472 a_n1455_n3628.n283 a_n1455_n3628.n282 5.04292
R20473 a_n1455_n3628.n257 a_n1455_n3628.n256 5.04292
R20474 a_n1455_n3628.n231 a_n1455_n3628.n230 5.04292
R20475 a_n1455_n3628.n205 a_n1455_n3628.n204 5.04292
R20476 a_n1455_n3628.n71 a_n1455_n3628.n70 5.04292
R20477 a_n1455_n3628.n99 a_n1455_n3628.n98 5.04292
R20478 a_n1455_n3628.n125 a_n1455_n3628.n124 5.04292
R20479 a_n1455_n3628.n153 a_n1455_n3628.n152 5.04292
R20480 a_n1455_n3628.n343 a_n1455_n3628.n342 5.04292
R20481 a_n1455_n3628.n354 a_n1455_n3628.n39 4.38594
R20482 a_n1455_n3628.n3 a_n1455_n3628.n295 4.38594
R20483 a_n1455_n3628.n7 a_n1455_n3628.n322 4.38594
R20484 a_n1455_n3628.n11 a_n1455_n3628.n164 4.38594
R20485 a_n1455_n3628.n17 a_n1455_n3628.n268 4.38594
R20486 a_n1455_n3628.n20 a_n1455_n3628.n242 4.38594
R20487 a_n1455_n3628.n23 a_n1455_n3628.n216 4.38594
R20488 a_n1455_n3628.n26 a_n1455_n3628.n190 4.38594
R20489 a_n1455_n3628.n29 a_n1455_n3628.n56 4.38594
R20490 a_n1455_n3628.n32 a_n1455_n3628.n84 4.38594
R20491 a_n1455_n3628.n35 a_n1455_n3628.n110 4.38594
R20492 a_n1455_n3628.n38 a_n1455_n3628.n138 4.38594
R20493 a_n1455_n3628.n306 a_n1455_n3628.n289 4.26717
R20494 a_n1455_n3628.n333 a_n1455_n3628.n316 4.26717
R20495 a_n1455_n3628.n175 a_n1455_n3628.n158 4.26717
R20496 a_n1455_n3628.n279 a_n1455_n3628.n262 4.26717
R20497 a_n1455_n3628.n253 a_n1455_n3628.n236 4.26717
R20498 a_n1455_n3628.n227 a_n1455_n3628.n210 4.26717
R20499 a_n1455_n3628.n201 a_n1455_n3628.n184 4.26717
R20500 a_n1455_n3628.n67 a_n1455_n3628.n50 4.26717
R20501 a_n1455_n3628.n95 a_n1455_n3628.n78 4.26717
R20502 a_n1455_n3628.n121 a_n1455_n3628.n104 4.26717
R20503 a_n1455_n3628.n149 a_n1455_n3628.n132 4.26717
R20504 a_n1455_n3628.n346 a_n1455_n3628.n45 4.26717
R20505 a_n1455_n3628.n305 a_n1455_n3628.n291 3.49141
R20506 a_n1455_n3628.n332 a_n1455_n3628.n318 3.49141
R20507 a_n1455_n3628.n174 a_n1455_n3628.n160 3.49141
R20508 a_n1455_n3628.n278 a_n1455_n3628.n264 3.49141
R20509 a_n1455_n3628.n252 a_n1455_n3628.n238 3.49141
R20510 a_n1455_n3628.n226 a_n1455_n3628.n212 3.49141
R20511 a_n1455_n3628.n200 a_n1455_n3628.n186 3.49141
R20512 a_n1455_n3628.n66 a_n1455_n3628.n52 3.49141
R20513 a_n1455_n3628.n94 a_n1455_n3628.n80 3.49141
R20514 a_n1455_n3628.n120 a_n1455_n3628.n106 3.49141
R20515 a_n1455_n3628.n148 a_n1455_n3628.n134 3.49141
R20516 a_n1455_n3628.n347 a_n1455_n3628.n44 3.49141
R20517 a_n1455_n3628.n313 a_n1455_n3628.t3 3.3005
R20518 a_n1455_n3628.n313 a_n1455_n3628.t5 3.3005
R20519 a_n1455_n3628.n47 a_n1455_n3628.t10 3.3005
R20520 a_n1455_n3628.n47 a_n1455_n3628.t6 3.3005
R20521 a_n1455_n3628.n75 a_n1455_n3628.t12 3.3005
R20522 a_n1455_n3628.n75 a_n1455_n3628.t7 3.3005
R20523 a_n1455_n3628.n129 a_n1455_n3628.t17 3.3005
R20524 a_n1455_n3628.n129 a_n1455_n3628.t4 3.3005
R20525 a_n1455_n3628.n304 a_n1455_n3628.n303 2.71565
R20526 a_n1455_n3628.n331 a_n1455_n3628.n330 2.71565
R20527 a_n1455_n3628.n173 a_n1455_n3628.n172 2.71565
R20528 a_n1455_n3628.n277 a_n1455_n3628.n276 2.71565
R20529 a_n1455_n3628.n251 a_n1455_n3628.n250 2.71565
R20530 a_n1455_n3628.n225 a_n1455_n3628.n224 2.71565
R20531 a_n1455_n3628.n199 a_n1455_n3628.n198 2.71565
R20532 a_n1455_n3628.n65 a_n1455_n3628.n64 2.71565
R20533 a_n1455_n3628.n93 a_n1455_n3628.n92 2.71565
R20534 a_n1455_n3628.n119 a_n1455_n3628.n118 2.71565
R20535 a_n1455_n3628.n147 a_n1455_n3628.n146 2.71565
R20536 a_n1455_n3628.n349 a_n1455_n3628.n348 2.71565
R20537 a_n1455_n3628.n287 a_n1455_n3628.n286 2.23674
R20538 a_n1455_n3628.n208 a_n1455_n3628.n182 1.95694
R20539 a_n1455_n3628.n300 a_n1455_n3628.n292 1.93989
R20540 a_n1455_n3628.n327 a_n1455_n3628.n319 1.93989
R20541 a_n1455_n3628.n169 a_n1455_n3628.n161 1.93989
R20542 a_n1455_n3628.n273 a_n1455_n3628.n265 1.93989
R20543 a_n1455_n3628.n247 a_n1455_n3628.n239 1.93989
R20544 a_n1455_n3628.n221 a_n1455_n3628.n213 1.93989
R20545 a_n1455_n3628.n195 a_n1455_n3628.n187 1.93989
R20546 a_n1455_n3628.n61 a_n1455_n3628.n53 1.93989
R20547 a_n1455_n3628.n89 a_n1455_n3628.n81 1.93989
R20548 a_n1455_n3628.n115 a_n1455_n3628.n107 1.93989
R20549 a_n1455_n3628.n143 a_n1455_n3628.n135 1.93989
R20550 a_n1455_n3628.n352 a_n1455_n3628.n42 1.93989
R20551 a_n1455_n3628.n299 a_n1455_n3628.n294 1.16414
R20552 a_n1455_n3628.n326 a_n1455_n3628.n321 1.16414
R20553 a_n1455_n3628.n168 a_n1455_n3628.n163 1.16414
R20554 a_n1455_n3628.n272 a_n1455_n3628.n267 1.16414
R20555 a_n1455_n3628.n246 a_n1455_n3628.n241 1.16414
R20556 a_n1455_n3628.n220 a_n1455_n3628.n215 1.16414
R20557 a_n1455_n3628.n194 a_n1455_n3628.n189 1.16414
R20558 a_n1455_n3628.n60 a_n1455_n3628.n55 1.16414
R20559 a_n1455_n3628.n88 a_n1455_n3628.n83 1.16414
R20560 a_n1455_n3628.n114 a_n1455_n3628.n109 1.16414
R20561 a_n1455_n3628.n142 a_n1455_n3628.n137 1.16414
R20562 a_n1455_n3628.n353 a_n1455_n3628.n41 1.16414
R20563 a_n1455_n3628.n260 a_n1455_n3628.n234 0.962709
R20564 a_n1455_n3628.n286 a_n1455_n3628.n260 0.962709
R20565 a_n1455_n3628.n156 a_n1455_n3628.n130 0.573776
R20566 a_n1455_n3628.n130 a_n1455_n3628.n128 0.573776
R20567 a_n1455_n3628.n102 a_n1455_n3628.n76 0.573776
R20568 a_n1455_n3628.n76 a_n1455_n3628.n74 0.573776
R20569 a_n1455_n3628.n181 a_n1455_n3628.n48 0.573776
R20570 a_n1455_n3628.n340 a_n1455_n3628.n48 0.573776
R20571 a_n1455_n3628.n339 a_n1455_n3628.n314 0.573776
R20572 a_n1455_n3628.n314 a_n1455_n3628.n312 0.573776
R20573 a_n1455_n3628.n234 a_n1455_n3628.n208 0.422738
R20574 a_n1455_n3628.n298 a_n1455_n3628.n297 0.388379
R20575 a_n1455_n3628.n325 a_n1455_n3628.n324 0.388379
R20576 a_n1455_n3628.n167 a_n1455_n3628.n166 0.388379
R20577 a_n1455_n3628.n271 a_n1455_n3628.n270 0.388379
R20578 a_n1455_n3628.n245 a_n1455_n3628.n244 0.388379
R20579 a_n1455_n3628.n219 a_n1455_n3628.n218 0.388379
R20580 a_n1455_n3628.n193 a_n1455_n3628.n192 0.388379
R20581 a_n1455_n3628.n59 a_n1455_n3628.n58 0.388379
R20582 a_n1455_n3628.n87 a_n1455_n3628.n86 0.388379
R20583 a_n1455_n3628.n113 a_n1455_n3628.n112 0.388379
R20584 a_n1455_n3628.n141 a_n1455_n3628.n140 0.388379
R20585 a_n1455_n3628.n356 a_n1455_n3628.n355 0.388379
R20586 a_n1455_n3628.n38 a_n1455_n3628.n36 0.310845
R20587 a_n1455_n3628.n37 a_n1455_n3628.n36 0.310845
R20588 a_n1455_n3628.n154 a_n1455_n3628.n37 0.310845
R20589 a_n1455_n3628.n35 a_n1455_n3628.n33 0.310845
R20590 a_n1455_n3628.n34 a_n1455_n3628.n33 0.310845
R20591 a_n1455_n3628.n126 a_n1455_n3628.n34 0.310845
R20592 a_n1455_n3628.n32 a_n1455_n3628.n30 0.310845
R20593 a_n1455_n3628.n31 a_n1455_n3628.n30 0.310845
R20594 a_n1455_n3628.n100 a_n1455_n3628.n31 0.310845
R20595 a_n1455_n3628.n29 a_n1455_n3628.n27 0.310845
R20596 a_n1455_n3628.n28 a_n1455_n3628.n27 0.310845
R20597 a_n1455_n3628.n72 a_n1455_n3628.n28 0.310845
R20598 a_n1455_n3628.n26 a_n1455_n3628.n24 0.310845
R20599 a_n1455_n3628.n25 a_n1455_n3628.n24 0.310845
R20600 a_n1455_n3628.n206 a_n1455_n3628.n25 0.310845
R20601 a_n1455_n3628.n23 a_n1455_n3628.n21 0.310845
R20602 a_n1455_n3628.n22 a_n1455_n3628.n21 0.310845
R20603 a_n1455_n3628.n232 a_n1455_n3628.n22 0.310845
R20604 a_n1455_n3628.n20 a_n1455_n3628.n18 0.310845
R20605 a_n1455_n3628.n19 a_n1455_n3628.n18 0.310845
R20606 a_n1455_n3628.n258 a_n1455_n3628.n19 0.310845
R20607 a_n1455_n3628.n17 a_n1455_n3628.n15 0.310845
R20608 a_n1455_n3628.n16 a_n1455_n3628.n15 0.310845
R20609 a_n1455_n3628.n284 a_n1455_n3628.n16 0.310845
R20610 a_n1455_n3628.n14 a_n1455_n3628.n13 0.310845
R20611 a_n1455_n3628.n14 a_n1455_n3628.n12 0.310845
R20612 a_n1455_n3628.n12 a_n1455_n3628.n11 0.310845
R20613 a_n1455_n3628.n10 a_n1455_n3628.n9 0.310845
R20614 a_n1455_n3628.n10 a_n1455_n3628.n8 0.310845
R20615 a_n1455_n3628.n8 a_n1455_n3628.n7 0.310845
R20616 a_n1455_n3628.n6 a_n1455_n3628.n5 0.310845
R20617 a_n1455_n3628.n6 a_n1455_n3628.n4 0.310845
R20618 a_n1455_n3628.n4 a_n1455_n3628.n3 0.310845
R20619 a_n1455_n3628.n2 a_n1455_n3628.n1 0.310845
R20620 a_n1455_n3628.n2 a_n1455_n3628.n0 0.310845
R20621 a_n1455_n3628.n354 a_n1455_n3628.n0 0.310845
R20622 a_n1455_n3628.n128 a_n1455_n3628.n102 0.235414
R20623 a_n1455_n3628.n340 a_n1455_n3628.n339 0.235414
R20624 a_n2686_12378.n115 a_n2686_12378.n95 756.745
R20625 a_n2686_12378.n86 a_n2686_12378.n66 756.745
R20626 a_n2686_12378.n163 a_n2686_12378.n143 756.745
R20627 a_n2686_12378.n192 a_n2686_12378.n172 756.745
R20628 a_n2686_12378.n116 a_n2686_12378.n115 585
R20629 a_n2686_12378.n114 a_n2686_12378.n113 585
R20630 a_n2686_12378.n98 a_n2686_12378.n97 585
R20631 a_n2686_12378.n110 a_n2686_12378.n109 585
R20632 a_n2686_12378.n108 a_n2686_12378.n107 585
R20633 a_n2686_12378.n101 a_n2686_12378.n100 585
R20634 a_n2686_12378.n104 a_n2686_12378.n103 585
R20635 a_n2686_12378.n87 a_n2686_12378.n86 585
R20636 a_n2686_12378.n85 a_n2686_12378.n84 585
R20637 a_n2686_12378.n69 a_n2686_12378.n68 585
R20638 a_n2686_12378.n81 a_n2686_12378.n80 585
R20639 a_n2686_12378.n79 a_n2686_12378.n78 585
R20640 a_n2686_12378.n72 a_n2686_12378.n71 585
R20641 a_n2686_12378.n75 a_n2686_12378.n74 585
R20642 a_n2686_12378.n164 a_n2686_12378.n163 585
R20643 a_n2686_12378.n162 a_n2686_12378.n161 585
R20644 a_n2686_12378.n146 a_n2686_12378.n145 585
R20645 a_n2686_12378.n158 a_n2686_12378.n157 585
R20646 a_n2686_12378.n156 a_n2686_12378.n155 585
R20647 a_n2686_12378.n149 a_n2686_12378.n148 585
R20648 a_n2686_12378.n152 a_n2686_12378.n151 585
R20649 a_n2686_12378.n193 a_n2686_12378.n192 585
R20650 a_n2686_12378.n191 a_n2686_12378.n190 585
R20651 a_n2686_12378.n175 a_n2686_12378.n174 585
R20652 a_n2686_12378.n187 a_n2686_12378.n186 585
R20653 a_n2686_12378.n185 a_n2686_12378.n184 585
R20654 a_n2686_12378.n178 a_n2686_12378.n177 585
R20655 a_n2686_12378.n181 a_n2686_12378.n180 585
R20656 a_n2686_12378.t6 a_n2686_12378.n102 327.601
R20657 a_n2686_12378.t16 a_n2686_12378.n73 327.601
R20658 a_n2686_12378.t4 a_n2686_12378.n150 327.601
R20659 a_n2686_12378.t20 a_n2686_12378.n179 327.601
R20660 a_n2686_12378.n141 a_n2686_12378.t19 183.883
R20661 a_n2686_12378.n133 a_n2686_12378.t3 183.883
R20662 a_n2686_12378.n225 a_n2686_12378.t56 183.883
R20663 a_n2686_12378.n230 a_n2686_12378.t47 183.883
R20664 a_n2686_12378.n217 a_n2686_12378.t48 183.883
R20665 a_n2686_12378.n222 a_n2686_12378.t39 183.883
R20666 a_n2686_12378.n209 a_n2686_12378.t33 183.883
R20667 a_n2686_12378.n214 a_n2686_12378.t43 183.883
R20668 a_n2686_12378.n201 a_n2686_12378.t36 183.883
R20669 a_n2686_12378.n206 a_n2686_12378.t45 183.883
R20670 a_n2686_12378.n10 a_n2686_12378.t15 206.089
R20671 a_n2686_12378.n8 a_n2686_12378.t52 206.089
R20672 a_n2686_12378.n12 a_n2686_12378.t40 206.089
R20673 a_n2686_12378.n115 a_n2686_12378.n114 171.744
R20674 a_n2686_12378.n114 a_n2686_12378.n97 171.744
R20675 a_n2686_12378.n109 a_n2686_12378.n97 171.744
R20676 a_n2686_12378.n109 a_n2686_12378.n108 171.744
R20677 a_n2686_12378.n108 a_n2686_12378.n100 171.744
R20678 a_n2686_12378.n103 a_n2686_12378.n100 171.744
R20679 a_n2686_12378.n86 a_n2686_12378.n85 171.744
R20680 a_n2686_12378.n85 a_n2686_12378.n68 171.744
R20681 a_n2686_12378.n80 a_n2686_12378.n68 171.744
R20682 a_n2686_12378.n80 a_n2686_12378.n79 171.744
R20683 a_n2686_12378.n79 a_n2686_12378.n71 171.744
R20684 a_n2686_12378.n74 a_n2686_12378.n71 171.744
R20685 a_n2686_12378.n163 a_n2686_12378.n162 171.744
R20686 a_n2686_12378.n162 a_n2686_12378.n145 171.744
R20687 a_n2686_12378.n157 a_n2686_12378.n145 171.744
R20688 a_n2686_12378.n157 a_n2686_12378.n156 171.744
R20689 a_n2686_12378.n156 a_n2686_12378.n148 171.744
R20690 a_n2686_12378.n151 a_n2686_12378.n148 171.744
R20691 a_n2686_12378.n192 a_n2686_12378.n191 171.744
R20692 a_n2686_12378.n191 a_n2686_12378.n174 171.744
R20693 a_n2686_12378.n186 a_n2686_12378.n174 171.744
R20694 a_n2686_12378.n186 a_n2686_12378.n185 171.744
R20695 a_n2686_12378.n185 a_n2686_12378.n177 171.744
R20696 a_n2686_12378.n180 a_n2686_12378.n177 171.744
R20697 a_n2686_12378.n17 a_n2686_12378.n5 68.6201
R20698 a_n2686_12378.n5 a_n2686_12378.n16 71.6402
R20699 a_n2686_12378.n129 a_n2686_12378.n7 161.3
R20700 a_n2686_12378.n7 a_n2686_12378.n15 68.6201
R20701 a_n2686_12378.n19 a_n2686_12378.n3 68.6201
R20702 a_n2686_12378.n3 a_n2686_12378.n18 71.6402
R20703 a_n2686_12378.n126 a_n2686_12378.n9 161.3
R20704 a_n2686_12378.n9 a_n2686_12378.n14 68.6201
R20705 a_n2686_12378.n21 a_n2686_12378.n0 68.6201
R20706 a_n2686_12378.n0 a_n2686_12378.n20 71.6402
R20707 a_n2686_12378.n234 a_n2686_12378.n11 161.3
R20708 a_n2686_12378.n11 a_n2686_12378.n13 68.6201
R20709 a_n2686_12378.n205 a_n2686_12378.n26 161.3
R20710 a_n2686_12378.n22 a_n2686_12378.n26 161.3
R20711 a_n2686_12378.n25 a_n2686_12378.n23 71.6402
R20712 a_n2686_12378.n202 a_n2686_12378.n24 161.3
R20713 a_n2686_12378.n213 a_n2686_12378.n31 161.3
R20714 a_n2686_12378.n27 a_n2686_12378.n31 161.3
R20715 a_n2686_12378.n30 a_n2686_12378.n28 71.6402
R20716 a_n2686_12378.n210 a_n2686_12378.n29 161.3
R20717 a_n2686_12378.n221 a_n2686_12378.n36 161.3
R20718 a_n2686_12378.n32 a_n2686_12378.n36 161.3
R20719 a_n2686_12378.n35 a_n2686_12378.n33 71.6402
R20720 a_n2686_12378.n218 a_n2686_12378.n34 161.3
R20721 a_n2686_12378.n229 a_n2686_12378.n41 161.3
R20722 a_n2686_12378.n37 a_n2686_12378.n41 161.3
R20723 a_n2686_12378.n40 a_n2686_12378.n38 71.6402
R20724 a_n2686_12378.n226 a_n2686_12378.n39 161.3
R20725 a_n2686_12378.n51 a_n2686_12378.n48 74.8341
R20726 a_n2686_12378.n49 a_n2686_12378.n46 68.6201
R20727 a_n2686_12378.n45 a_n2686_12378.n47 71.6402
R20728 a_n2686_12378.n135 a_n2686_12378.n42 161.3
R20729 a_n2686_12378.n137 a_n2686_12378.n42 161.3
R20730 a_n2686_12378.n44 a_n2686_12378.n138 161.3
R20731 a_n2686_12378.n139 a_n2686_12378.n44 161.3
R20732 a_n2686_12378.n140 a_n2686_12378.n43 161.3
R20733 a_n2686_12378.n131 a_n2686_12378.t13 144.601
R20734 a_n2686_12378.n136 a_n2686_12378.t23 144.601
R20735 a_n2686_12378.n134 a_n2686_12378.t25 144.601
R20736 a_n2686_12378.n132 a_n2686_12378.t11 144.601
R20737 a_n2686_12378.n227 a_n2686_12378.t42 144.601
R20738 a_n2686_12378.n228 a_n2686_12378.t59 144.601
R20739 a_n2686_12378.n219 a_n2686_12378.t58 144.601
R20740 a_n2686_12378.n220 a_n2686_12378.t55 144.601
R20741 a_n2686_12378.n211 a_n2686_12378.t50 144.601
R20742 a_n2686_12378.n212 a_n2686_12378.t54 144.601
R20743 a_n2686_12378.n203 a_n2686_12378.t53 144.601
R20744 a_n2686_12378.n204 a_n2686_12378.t34 144.601
R20745 a_n2686_12378.n123 a_n2686_12378.t7 144.601
R20746 a_n2686_12378.n127 a_n2686_12378.t9 144.601
R20747 a_n2686_12378.n125 a_n2686_12378.t21 144.601
R20748 a_n2686_12378.n124 a_n2686_12378.t17 144.601
R20749 a_n2686_12378.n121 a_n2686_12378.t57 144.601
R20750 a_n2686_12378.n130 a_n2686_12378.t35 144.601
R20751 a_n2686_12378.n128 a_n2686_12378.t51 144.601
R20752 a_n2686_12378.n122 a_n2686_12378.t32 144.601
R20753 a_n2686_12378.n64 a_n2686_12378.t49 144.601
R20754 a_n2686_12378.n235 a_n2686_12378.t46 144.601
R20755 a_n2686_12378.n233 a_n2686_12378.t37 144.601
R20756 a_n2686_12378.n65 a_n2686_12378.t44 144.601
R20757 a_n2686_12378.n103 a_n2686_12378.t6 85.8723
R20758 a_n2686_12378.n74 a_n2686_12378.t16 85.8723
R20759 a_n2686_12378.n151 a_n2686_12378.t4 85.8723
R20760 a_n2686_12378.n180 a_n2686_12378.t20 85.8723
R20761 a_n2686_12378.n243 a_n2686_12378.n242 84.3504
R20762 a_n2686_12378.n238 a_n2686_12378.n237 84.3502
R20763 a_n2686_12378.n242 a_n2686_12378.n241 84.35
R20764 a_n2686_12378.n240 a_n2686_12378.n239 84.0635
R20765 a_n2686_12378.n94 a_n2686_12378.n93 81.2397
R20766 a_n2686_12378.n92 a_n2686_12378.n91 81.2397
R20767 a_n2686_12378.n169 a_n2686_12378.n168 81.2397
R20768 a_n2686_12378.n171 a_n2686_12378.n170 81.2397
R20769 a_n2686_12378.n6 a_n2686_12378.n5 28.1161
R20770 a_n2686_12378.n7 a_n2686_12378.n8 28.1161
R20771 a_n2686_12378.n4 a_n2686_12378.n3 28.1161
R20772 a_n2686_12378.n9 a_n2686_12378.n10 28.1161
R20773 a_n2686_12378.n1 a_n2686_12378.n0 28.1161
R20774 a_n2686_12378.n11 a_n2686_12378.n12 28.1161
R20775 a_n2686_12378.n207 a_n2686_12378.n206 80.6037
R20776 a_n2686_12378.n201 a_n2686_12378.n200 80.6037
R20777 a_n2686_12378.n215 a_n2686_12378.n214 80.6037
R20778 a_n2686_12378.n209 a_n2686_12378.n208 80.6037
R20779 a_n2686_12378.n223 a_n2686_12378.n222 80.6037
R20780 a_n2686_12378.n217 a_n2686_12378.n216 80.6037
R20781 a_n2686_12378.n231 a_n2686_12378.n230 80.6037
R20782 a_n2686_12378.n225 a_n2686_12378.n224 80.6037
R20783 a_n2686_12378.n133 a_n2686_12378.n50 80.6037
R20784 a_n2686_12378.n142 a_n2686_12378.n141 80.6037
R20785 a_n2686_12378.n138 a_n2686_12378.n137 56.5617
R20786 a_n2686_12378.n49 a_n2686_12378.n132 48.4088
R20787 a_n2686_12378.n19 a_n2686_12378.n124 48.4088
R20788 a_n2686_12378.n17 a_n2686_12378.n122 48.4088
R20789 a_n2686_12378.n21 a_n2686_12378.n65 48.4088
R20790 a_n2686_12378.n226 a_n2686_12378.n225 56.3158
R20791 a_n2686_12378.n230 a_n2686_12378.n229 56.3158
R20792 a_n2686_12378.n218 a_n2686_12378.n217 56.3158
R20793 a_n2686_12378.n222 a_n2686_12378.n221 56.3158
R20794 a_n2686_12378.n210 a_n2686_12378.n209 56.3158
R20795 a_n2686_12378.n214 a_n2686_12378.n213 56.3158
R20796 a_n2686_12378.n202 a_n2686_12378.n201 56.3158
R20797 a_n2686_12378.n206 a_n2686_12378.n205 56.3158
R20798 a_n2686_12378.n141 a_n2686_12378.n140 47.4702
R20799 a_n2686_12378.n135 a_n2686_12378.n47 58.5991
R20800 a_n2686_12378.n134 a_n2686_12378.n47 26.1378
R20801 a_n2686_12378.n38 a_n2686_12378.n37 58.5991
R20802 a_n2686_12378.n33 a_n2686_12378.n32 58.5991
R20803 a_n2686_12378.n28 a_n2686_12378.n27 58.5991
R20804 a_n2686_12378.n23 a_n2686_12378.n22 58.5991
R20805 a_n2686_12378.n126 a_n2686_12378.n18 58.5991
R20806 a_n2686_12378.n125 a_n2686_12378.n18 26.1378
R20807 a_n2686_12378.n129 a_n2686_12378.n16 58.5991
R20808 a_n2686_12378.n128 a_n2686_12378.n16 26.1378
R20809 a_n2686_12378.n234 a_n2686_12378.n20 58.5991
R20810 a_n2686_12378.n233 a_n2686_12378.n20 26.1378
R20811 a_n2686_12378.n92 a_n2686_12378.n90 38.3829
R20812 a_n2686_12378.n169 a_n2686_12378.n167 38.3829
R20813 a_n2686_12378.n120 a_n2686_12378.n119 37.8096
R20814 a_n2686_12378.n197 a_n2686_12378.n196 37.8096
R20815 a_n2686_12378.n242 a_n2686_12378.n240 29.8404
R20816 a_n2686_12378.n140 a_n2686_12378.n139 25.0767
R20817 a_n2686_12378.n51 a_n2686_12378.n133 59.1045
R20818 a_n2686_12378.n10 a_n2686_12378.n123 32.4972
R20819 a_n2686_12378.n4 a_n2686_12378.t5 206.089
R20820 a_n2686_12378.n8 a_n2686_12378.n121 32.4972
R20821 a_n2686_12378.n6 a_n2686_12378.t38 206.089
R20822 a_n2686_12378.n12 a_n2686_12378.n64 32.4972
R20823 a_n2686_12378.n1 a_n2686_12378.t41 206.089
R20824 a_n2686_12378.n138 a_n2686_12378.n131 24.3464
R20825 a_n2686_12378.n14 a_n2686_12378.n123 48.4088
R20826 a_n2686_12378.n15 a_n2686_12378.n121 48.4088
R20827 a_n2686_12378.n13 a_n2686_12378.n64 48.4088
R20828 a_n2686_12378.n238 a_n2686_12378.n236 23.892
R20829 a_n2686_12378.n137 a_n2686_12378.n136 16.477
R20830 a_n2686_12378.n134 a_n2686_12378.n49 40.5394
R20831 a_n2686_12378.n227 a_n2686_12378.n226 16.477
R20832 a_n2686_12378.n229 a_n2686_12378.n228 16.477
R20833 a_n2686_12378.n219 a_n2686_12378.n218 16.477
R20834 a_n2686_12378.n221 a_n2686_12378.n220 16.477
R20835 a_n2686_12378.n211 a_n2686_12378.n210 16.477
R20836 a_n2686_12378.n213 a_n2686_12378.n212 16.477
R20837 a_n2686_12378.n203 a_n2686_12378.n202 16.477
R20838 a_n2686_12378.n205 a_n2686_12378.n204 16.477
R20839 a_n2686_12378.n14 a_n2686_12378.n127 40.5394
R20840 a_n2686_12378.n125 a_n2686_12378.n19 40.5394
R20841 a_n2686_12378.n15 a_n2686_12378.n130 40.5394
R20842 a_n2686_12378.n128 a_n2686_12378.n17 40.5394
R20843 a_n2686_12378.n13 a_n2686_12378.n235 40.5394
R20844 a_n2686_12378.n233 a_n2686_12378.n21 40.5394
R20845 a_n2686_12378.n104 a_n2686_12378.n102 16.3865
R20846 a_n2686_12378.n75 a_n2686_12378.n73 16.3865
R20847 a_n2686_12378.n152 a_n2686_12378.n150 16.3865
R20848 a_n2686_12378.n181 a_n2686_12378.n179 16.3865
R20849 a_n2686_12378.n105 a_n2686_12378.n101 12.8005
R20850 a_n2686_12378.n76 a_n2686_12378.n72 12.8005
R20851 a_n2686_12378.n153 a_n2686_12378.n149 12.8005
R20852 a_n2686_12378.n182 a_n2686_12378.n178 12.8005
R20853 a_n2686_12378.n107 a_n2686_12378.n106 12.0247
R20854 a_n2686_12378.n78 a_n2686_12378.n77 12.0247
R20855 a_n2686_12378.n155 a_n2686_12378.n154 12.0247
R20856 a_n2686_12378.n184 a_n2686_12378.n183 12.0247
R20857 a_n2686_12378.n110 a_n2686_12378.n99 11.249
R20858 a_n2686_12378.n81 a_n2686_12378.n70 11.249
R20859 a_n2686_12378.n158 a_n2686_12378.n147 11.249
R20860 a_n2686_12378.n187 a_n2686_12378.n176 11.249
R20861 a_n2686_12378.n199 a_n2686_12378.n7 10.8153
R20862 a_n2686_12378.n0 a_n2686_12378.n232 10.6108
R20863 a_n2686_12378.n111 a_n2686_12378.n98 10.4732
R20864 a_n2686_12378.n82 a_n2686_12378.n69 10.4732
R20865 a_n2686_12378.n159 a_n2686_12378.n146 10.4732
R20866 a_n2686_12378.n188 a_n2686_12378.n175 10.4732
R20867 a_n2686_12378.n113 a_n2686_12378.n112 9.69747
R20868 a_n2686_12378.n84 a_n2686_12378.n83 9.69747
R20869 a_n2686_12378.n161 a_n2686_12378.n160 9.69747
R20870 a_n2686_12378.n190 a_n2686_12378.n189 9.69747
R20871 a_n2686_12378.n119 a_n2686_12378.n118 9.45567
R20872 a_n2686_12378.n90 a_n2686_12378.n89 9.45567
R20873 a_n2686_12378.n167 a_n2686_12378.n166 9.45567
R20874 a_n2686_12378.n196 a_n2686_12378.n195 9.45567
R20875 a_n2686_12378.n198 a_n2686_12378.n142 9.30587
R20876 a_n2686_12378.n118 a_n2686_12378.n117 9.3005
R20877 a_n2686_12378.n96 a_n2686_12378.n53 9.3005
R20878 a_n2686_12378.n112 a_n2686_12378.n53 9.3005
R20879 a_n2686_12378.n52 a_n2686_12378.n111 9.3005
R20880 a_n2686_12378.n99 a_n2686_12378.n52 9.3005
R20881 a_n2686_12378.n106 a_n2686_12378.n54 9.3005
R20882 a_n2686_12378.n54 a_n2686_12378.n105 9.3005
R20883 a_n2686_12378.n89 a_n2686_12378.n88 9.3005
R20884 a_n2686_12378.n67 a_n2686_12378.n56 9.3005
R20885 a_n2686_12378.n83 a_n2686_12378.n56 9.3005
R20886 a_n2686_12378.n55 a_n2686_12378.n82 9.3005
R20887 a_n2686_12378.n70 a_n2686_12378.n55 9.3005
R20888 a_n2686_12378.n77 a_n2686_12378.n57 9.3005
R20889 a_n2686_12378.n57 a_n2686_12378.n76 9.3005
R20890 a_n2686_12378.n166 a_n2686_12378.n165 9.3005
R20891 a_n2686_12378.n144 a_n2686_12378.n59 9.3005
R20892 a_n2686_12378.n160 a_n2686_12378.n59 9.3005
R20893 a_n2686_12378.n58 a_n2686_12378.n159 9.3005
R20894 a_n2686_12378.n147 a_n2686_12378.n58 9.3005
R20895 a_n2686_12378.n154 a_n2686_12378.n60 9.3005
R20896 a_n2686_12378.n60 a_n2686_12378.n153 9.3005
R20897 a_n2686_12378.n195 a_n2686_12378.n194 9.3005
R20898 a_n2686_12378.n173 a_n2686_12378.n62 9.3005
R20899 a_n2686_12378.n189 a_n2686_12378.n62 9.3005
R20900 a_n2686_12378.n61 a_n2686_12378.n188 9.3005
R20901 a_n2686_12378.n176 a_n2686_12378.n61 9.3005
R20902 a_n2686_12378.n183 a_n2686_12378.n63 9.3005
R20903 a_n2686_12378.n63 a_n2686_12378.n182 9.3005
R20904 a_n2686_12378.n116 a_n2686_12378.n96 8.92171
R20905 a_n2686_12378.n87 a_n2686_12378.n67 8.92171
R20906 a_n2686_12378.n164 a_n2686_12378.n144 8.92171
R20907 a_n2686_12378.n193 a_n2686_12378.n173 8.92171
R20908 a_n2686_12378.n2 a_n2686_12378.n120 8.2571
R20909 a_n2686_12378.n117 a_n2686_12378.n95 8.14595
R20910 a_n2686_12378.n88 a_n2686_12378.n66 8.14595
R20911 a_n2686_12378.n165 a_n2686_12378.n143 8.14595
R20912 a_n2686_12378.n194 a_n2686_12378.n172 8.14595
R20913 a_n2686_12378.n136 a_n2686_12378.n135 8.11581
R20914 a_n2686_12378.n38 a_n2686_12378.n227 26.1378
R20915 a_n2686_12378.n228 a_n2686_12378.n37 8.11581
R20916 a_n2686_12378.n33 a_n2686_12378.n219 26.1378
R20917 a_n2686_12378.n220 a_n2686_12378.n32 8.11581
R20918 a_n2686_12378.n28 a_n2686_12378.n211 26.1378
R20919 a_n2686_12378.n212 a_n2686_12378.n27 8.11581
R20920 a_n2686_12378.n23 a_n2686_12378.n203 26.1378
R20921 a_n2686_12378.n204 a_n2686_12378.n22 8.11581
R20922 a_n2686_12378.n127 a_n2686_12378.n126 8.11581
R20923 a_n2686_12378.n130 a_n2686_12378.n129 8.11581
R20924 a_n2686_12378.n235 a_n2686_12378.n234 8.11581
R20925 a_n2686_12378.n232 a_n2686_12378.n231 7.00284
R20926 a_n2686_12378.n200 a_n2686_12378.n199 7.00284
R20927 a_n2686_12378.n3 a_n2686_12378.n2 6.60701
R20928 a_n2686_12378.n119 a_n2686_12378.n95 5.81868
R20929 a_n2686_12378.n90 a_n2686_12378.n66 5.81868
R20930 a_n2686_12378.n167 a_n2686_12378.n143 5.81868
R20931 a_n2686_12378.n196 a_n2686_12378.n172 5.81868
R20932 a_n2686_12378.n198 a_n2686_12378.n197 5.55007
R20933 a_n2686_12378.n93 a_n2686_12378.t22 5.418
R20934 a_n2686_12378.n93 a_n2686_12378.t18 5.418
R20935 a_n2686_12378.n91 a_n2686_12378.t8 5.418
R20936 a_n2686_12378.n91 a_n2686_12378.t10 5.418
R20937 a_n2686_12378.n168 a_n2686_12378.t26 5.418
R20938 a_n2686_12378.n168 a_n2686_12378.t12 5.418
R20939 a_n2686_12378.n170 a_n2686_12378.t14 5.418
R20940 a_n2686_12378.n170 a_n2686_12378.t24 5.418
R20941 a_n2686_12378.n117 a_n2686_12378.n116 5.04292
R20942 a_n2686_12378.n88 a_n2686_12378.n87 5.04292
R20943 a_n2686_12378.n165 a_n2686_12378.n164 5.04292
R20944 a_n2686_12378.n194 a_n2686_12378.n193 5.04292
R20945 a_n2686_12378.n5 a_n2686_12378.n9 4.52033
R20946 a_n2686_12378.n113 a_n2686_12378.n96 4.26717
R20947 a_n2686_12378.n84 a_n2686_12378.n67 4.26717
R20948 a_n2686_12378.n161 a_n2686_12378.n144 4.26717
R20949 a_n2686_12378.n190 a_n2686_12378.n173 4.26717
R20950 a_n2686_12378.n232 a_n2686_12378.n2 4.20883
R20951 a_n2686_12378.n54 a_n2686_12378.n102 3.71286
R20952 a_n2686_12378.n57 a_n2686_12378.n73 3.71286
R20953 a_n2686_12378.n60 a_n2686_12378.n150 3.71286
R20954 a_n2686_12378.n63 a_n2686_12378.n179 3.71286
R20955 a_n2686_12378.n112 a_n2686_12378.n98 3.49141
R20956 a_n2686_12378.n83 a_n2686_12378.n69 3.49141
R20957 a_n2686_12378.n160 a_n2686_12378.n146 3.49141
R20958 a_n2686_12378.n189 a_n2686_12378.n175 3.49141
R20959 a_n2686_12378.n236 a_n2686_12378.n11 3.45549
R20960 a_n2686_12378.n241 a_n2686_12378.t2 3.3005
R20961 a_n2686_12378.n241 a_n2686_12378.t31 3.3005
R20962 a_n2686_12378.n237 a_n2686_12378.t1 3.3005
R20963 a_n2686_12378.n237 a_n2686_12378.t27 3.3005
R20964 a_n2686_12378.n239 a_n2686_12378.t28 3.3005
R20965 a_n2686_12378.n239 a_n2686_12378.t29 3.3005
R20966 a_n2686_12378.n243 a_n2686_12378.t30 3.3005
R20967 a_n2686_12378.t0 a_n2686_12378.n243 3.3005
R20968 a_n2686_12378.n111 a_n2686_12378.n110 2.71565
R20969 a_n2686_12378.n82 a_n2686_12378.n81 2.71565
R20970 a_n2686_12378.n159 a_n2686_12378.n158 2.71565
R20971 a_n2686_12378.n188 a_n2686_12378.n187 2.71565
R20972 a_n2686_12378.n107 a_n2686_12378.n99 1.93989
R20973 a_n2686_12378.n78 a_n2686_12378.n70 1.93989
R20974 a_n2686_12378.n155 a_n2686_12378.n147 1.93989
R20975 a_n2686_12378.n184 a_n2686_12378.n176 1.93989
R20976 a_n2686_12378.n216 a_n2686_12378.n215 1.42563
R20977 a_n2686_12378.n199 a_n2686_12378.n198 1.30542
R20978 a_n2686_12378.n106 a_n2686_12378.n101 1.16414
R20979 a_n2686_12378.n77 a_n2686_12378.n72 1.16414
R20980 a_n2686_12378.n154 a_n2686_12378.n149 1.16414
R20981 a_n2686_12378.n183 a_n2686_12378.n178 1.16414
R20982 a_n2686_12378.n236 a_n2686_12378.n50 1.02746
R20983 a_n2686_12378.n208 a_n2686_12378.n207 0.96351
R20984 a_n2686_12378.n224 a_n2686_12378.n223 0.96351
R20985 a_n2686_12378.n94 a_n2686_12378.n92 0.573776
R20986 a_n2686_12378.n120 a_n2686_12378.n94 0.573776
R20987 a_n2686_12378.n197 a_n2686_12378.n171 0.573776
R20988 a_n2686_12378.n171 a_n2686_12378.n169 0.573776
R20989 a_n2686_12378.n105 a_n2686_12378.n104 0.388379
R20990 a_n2686_12378.n76 a_n2686_12378.n75 0.388379
R20991 a_n2686_12378.n153 a_n2686_12378.n152 0.388379
R20992 a_n2686_12378.n182 a_n2686_12378.n181 0.388379
R20993 a_n2686_12378.n46 a_n2686_12378.n48 0.379288
R20994 a_n2686_12378.n63 a_n2686_12378.n61 0.310845
R20995 a_n2686_12378.n62 a_n2686_12378.n61 0.310845
R20996 a_n2686_12378.n195 a_n2686_12378.n62 0.310845
R20997 a_n2686_12378.n60 a_n2686_12378.n58 0.310845
R20998 a_n2686_12378.n59 a_n2686_12378.n58 0.310845
R20999 a_n2686_12378.n166 a_n2686_12378.n59 0.310845
R21000 a_n2686_12378.n57 a_n2686_12378.n55 0.310845
R21001 a_n2686_12378.n56 a_n2686_12378.n55 0.310845
R21002 a_n2686_12378.n89 a_n2686_12378.n56 0.310845
R21003 a_n2686_12378.n54 a_n2686_12378.n52 0.310845
R21004 a_n2686_12378.n53 a_n2686_12378.n52 0.310845
R21005 a_n2686_12378.n118 a_n2686_12378.n53 0.310845
R21006 a_n2686_12378.n240 a_n2686_12378.n238 0.287138
R21007 a_n2686_12378.n200 a_n2686_12378.n24 0.285035
R21008 a_n2686_12378.n207 a_n2686_12378.n26 0.285035
R21009 a_n2686_12378.n208 a_n2686_12378.n29 0.285035
R21010 a_n2686_12378.n215 a_n2686_12378.n31 0.285035
R21011 a_n2686_12378.n216 a_n2686_12378.n34 0.285035
R21012 a_n2686_12378.n223 a_n2686_12378.n36 0.285035
R21013 a_n2686_12378.n224 a_n2686_12378.n39 0.285035
R21014 a_n2686_12378.n231 a_n2686_12378.n41 0.285035
R21015 a_n2686_12378.n142 a_n2686_12378.n43 0.285035
R21016 a_n2686_12378.n48 a_n2686_12378.n50 0.285035
R21017 a_n2686_12378.n139 a_n2686_12378.n131 0.246418
R21018 a_n2686_12378.n51 a_n2686_12378.n132 11.8807
R21019 a_n2686_12378.n45 a_n2686_12378.n46 0.379288
R21020 a_n2686_12378.n42 a_n2686_12378.n45 0.379288
R21021 a_n2686_12378.n44 a_n2686_12378.n42 0.379288
R21022 a_n2686_12378.n44 a_n2686_12378.n43 0.379288
R21023 a_n2686_12378.n41 a_n2686_12378.n40 0.379288
R21024 a_n2686_12378.n40 a_n2686_12378.n39 0.379288
R21025 a_n2686_12378.n36 a_n2686_12378.n35 0.379288
R21026 a_n2686_12378.n35 a_n2686_12378.n34 0.379288
R21027 a_n2686_12378.n31 a_n2686_12378.n30 0.379288
R21028 a_n2686_12378.n30 a_n2686_12378.n29 0.379288
R21029 a_n2686_12378.n26 a_n2686_12378.n25 0.379288
R21030 a_n2686_12378.n25 a_n2686_12378.n24 0.379288
R21031 a_n2686_12378.n4 a_n2686_12378.n124 32.4972
R21032 a_n2686_12378.n6 a_n2686_12378.n122 32.4972
R21033 a_n2686_12378.n1 a_n2686_12378.n65 32.4972
R21034 a_n2686_12378.n7 a_n2686_12378.n5 2.46351
R21035 a_n2686_12378.n9 a_n2686_12378.n3 2.46351
R21036 a_n2686_12378.n11 a_n2686_12378.n0 2.46351
R21037 a_n2511_10156.n133 a_n2511_10156.n107 756.745
R21038 a_n2511_10156.n99 a_n2511_10156.n73 756.745
R21039 a_n2511_10156.n67 a_n2511_10156.n41 756.745
R21040 a_n2511_10156.n34 a_n2511_10156.n8 756.745
R21041 a_n2511_10156.n134 a_n2511_10156.n133 585
R21042 a_n2511_10156.n132 a_n2511_10156.n131 585
R21043 a_n2511_10156.n111 a_n2511_10156.n110 585
R21044 a_n2511_10156.n126 a_n2511_10156.n125 585
R21045 a_n2511_10156.n124 a_n2511_10156.n123 585
R21046 a_n2511_10156.n115 a_n2511_10156.n114 585
R21047 a_n2511_10156.n118 a_n2511_10156.n117 585
R21048 a_n2511_10156.n100 a_n2511_10156.n99 585
R21049 a_n2511_10156.n98 a_n2511_10156.n97 585
R21050 a_n2511_10156.n77 a_n2511_10156.n76 585
R21051 a_n2511_10156.n92 a_n2511_10156.n91 585
R21052 a_n2511_10156.n90 a_n2511_10156.n89 585
R21053 a_n2511_10156.n81 a_n2511_10156.n80 585
R21054 a_n2511_10156.n84 a_n2511_10156.n83 585
R21055 a_n2511_10156.n68 a_n2511_10156.n67 585
R21056 a_n2511_10156.n66 a_n2511_10156.n65 585
R21057 a_n2511_10156.n45 a_n2511_10156.n44 585
R21058 a_n2511_10156.n60 a_n2511_10156.n59 585
R21059 a_n2511_10156.n58 a_n2511_10156.n57 585
R21060 a_n2511_10156.n49 a_n2511_10156.n48 585
R21061 a_n2511_10156.n52 a_n2511_10156.n51 585
R21062 a_n2511_10156.n35 a_n2511_10156.n34 585
R21063 a_n2511_10156.n33 a_n2511_10156.n32 585
R21064 a_n2511_10156.n12 a_n2511_10156.n11 585
R21065 a_n2511_10156.n27 a_n2511_10156.n26 585
R21066 a_n2511_10156.n25 a_n2511_10156.n24 585
R21067 a_n2511_10156.n16 a_n2511_10156.n15 585
R21068 a_n2511_10156.n19 a_n2511_10156.n18 585
R21069 a_n2511_10156.t5 a_n2511_10156.n116 327.601
R21070 a_n2511_10156.t2 a_n2511_10156.n82 327.601
R21071 a_n2511_10156.t7 a_n2511_10156.n50 327.601
R21072 a_n2511_10156.t4 a_n2511_10156.n17 327.601
R21073 a_n2511_10156.n133 a_n2511_10156.n132 171.744
R21074 a_n2511_10156.n132 a_n2511_10156.n110 171.744
R21075 a_n2511_10156.n125 a_n2511_10156.n110 171.744
R21076 a_n2511_10156.n125 a_n2511_10156.n124 171.744
R21077 a_n2511_10156.n124 a_n2511_10156.n114 171.744
R21078 a_n2511_10156.n117 a_n2511_10156.n114 171.744
R21079 a_n2511_10156.n99 a_n2511_10156.n98 171.744
R21080 a_n2511_10156.n98 a_n2511_10156.n76 171.744
R21081 a_n2511_10156.n91 a_n2511_10156.n76 171.744
R21082 a_n2511_10156.n91 a_n2511_10156.n90 171.744
R21083 a_n2511_10156.n90 a_n2511_10156.n80 171.744
R21084 a_n2511_10156.n83 a_n2511_10156.n80 171.744
R21085 a_n2511_10156.n67 a_n2511_10156.n66 171.744
R21086 a_n2511_10156.n66 a_n2511_10156.n44 171.744
R21087 a_n2511_10156.n59 a_n2511_10156.n44 171.744
R21088 a_n2511_10156.n59 a_n2511_10156.n58 171.744
R21089 a_n2511_10156.n58 a_n2511_10156.n48 171.744
R21090 a_n2511_10156.n51 a_n2511_10156.n48 171.744
R21091 a_n2511_10156.n34 a_n2511_10156.n33 171.744
R21092 a_n2511_10156.n33 a_n2511_10156.n11 171.744
R21093 a_n2511_10156.n26 a_n2511_10156.n11 171.744
R21094 a_n2511_10156.n26 a_n2511_10156.n25 171.744
R21095 a_n2511_10156.n25 a_n2511_10156.n15 171.744
R21096 a_n2511_10156.n18 a_n2511_10156.n15 171.744
R21097 a_n2511_10156.n2 a_n2511_10156.n0 109.74
R21098 a_n2511_10156.n5 a_n2511_10156.n3 109.401
R21099 a_n2511_10156.n2 a_n2511_10156.n1 109.166
R21100 a_n2511_10156.n7 a_n2511_10156.n6 109.166
R21101 a_n2511_10156.n5 a_n2511_10156.n4 109.166
R21102 a_n2511_10156.n141 a_n2511_10156.n140 109.166
R21103 a_n2511_10156.n117 a_n2511_10156.t5 85.8723
R21104 a_n2511_10156.n83 a_n2511_10156.t2 85.8723
R21105 a_n2511_10156.n51 a_n2511_10156.t7 85.8723
R21106 a_n2511_10156.n18 a_n2511_10156.t4 85.8723
R21107 a_n2511_10156.n106 a_n2511_10156.n105 81.2397
R21108 a_n2511_10156.n40 a_n2511_10156.n39 81.2397
R21109 a_n2511_10156.n40 a_n2511_10156.n38 38.3829
R21110 a_n2511_10156.n138 a_n2511_10156.n137 37.8096
R21111 a_n2511_10156.n104 a_n2511_10156.n103 37.8096
R21112 a_n2511_10156.n72 a_n2511_10156.n71 37.8096
R21113 a_n2511_10156.n118 a_n2511_10156.n116 16.3865
R21114 a_n2511_10156.n84 a_n2511_10156.n82 16.3865
R21115 a_n2511_10156.n52 a_n2511_10156.n50 16.3865
R21116 a_n2511_10156.n19 a_n2511_10156.n17 16.3865
R21117 a_n2511_10156.n139 a_n2511_10156.n7 13.2313
R21118 a_n2511_10156.n119 a_n2511_10156.n115 12.8005
R21119 a_n2511_10156.n85 a_n2511_10156.n81 12.8005
R21120 a_n2511_10156.n53 a_n2511_10156.n49 12.8005
R21121 a_n2511_10156.n20 a_n2511_10156.n16 12.8005
R21122 a_n2511_10156.n123 a_n2511_10156.n122 12.0247
R21123 a_n2511_10156.n89 a_n2511_10156.n88 12.0247
R21124 a_n2511_10156.n57 a_n2511_10156.n56 12.0247
R21125 a_n2511_10156.n24 a_n2511_10156.n23 12.0247
R21126 a_n2511_10156.n126 a_n2511_10156.n113 11.249
R21127 a_n2511_10156.n92 a_n2511_10156.n79 11.249
R21128 a_n2511_10156.n60 a_n2511_10156.n47 11.249
R21129 a_n2511_10156.n27 a_n2511_10156.n14 11.249
R21130 a_n2511_10156.n127 a_n2511_10156.n111 10.4732
R21131 a_n2511_10156.n93 a_n2511_10156.n77 10.4732
R21132 a_n2511_10156.n61 a_n2511_10156.n45 10.4732
R21133 a_n2511_10156.n28 a_n2511_10156.n12 10.4732
R21134 a_n2511_10156.n140 a_n2511_10156.n139 10.4398
R21135 a_n2511_10156.n131 a_n2511_10156.n130 9.69747
R21136 a_n2511_10156.n97 a_n2511_10156.n96 9.69747
R21137 a_n2511_10156.n65 a_n2511_10156.n64 9.69747
R21138 a_n2511_10156.n32 a_n2511_10156.n31 9.69747
R21139 a_n2511_10156.n137 a_n2511_10156.n136 9.45567
R21140 a_n2511_10156.n103 a_n2511_10156.n102 9.45567
R21141 a_n2511_10156.n71 a_n2511_10156.n70 9.45567
R21142 a_n2511_10156.n38 a_n2511_10156.n37 9.45567
R21143 a_n2511_10156.n136 a_n2511_10156.n135 9.3005
R21144 a_n2511_10156.n109 a_n2511_10156.n108 9.3005
R21145 a_n2511_10156.n130 a_n2511_10156.n129 9.3005
R21146 a_n2511_10156.n128 a_n2511_10156.n127 9.3005
R21147 a_n2511_10156.n113 a_n2511_10156.n112 9.3005
R21148 a_n2511_10156.n122 a_n2511_10156.n121 9.3005
R21149 a_n2511_10156.n120 a_n2511_10156.n119 9.3005
R21150 a_n2511_10156.n102 a_n2511_10156.n101 9.3005
R21151 a_n2511_10156.n75 a_n2511_10156.n74 9.3005
R21152 a_n2511_10156.n96 a_n2511_10156.n95 9.3005
R21153 a_n2511_10156.n94 a_n2511_10156.n93 9.3005
R21154 a_n2511_10156.n79 a_n2511_10156.n78 9.3005
R21155 a_n2511_10156.n88 a_n2511_10156.n87 9.3005
R21156 a_n2511_10156.n86 a_n2511_10156.n85 9.3005
R21157 a_n2511_10156.n70 a_n2511_10156.n69 9.3005
R21158 a_n2511_10156.n43 a_n2511_10156.n42 9.3005
R21159 a_n2511_10156.n64 a_n2511_10156.n63 9.3005
R21160 a_n2511_10156.n62 a_n2511_10156.n61 9.3005
R21161 a_n2511_10156.n47 a_n2511_10156.n46 9.3005
R21162 a_n2511_10156.n56 a_n2511_10156.n55 9.3005
R21163 a_n2511_10156.n54 a_n2511_10156.n53 9.3005
R21164 a_n2511_10156.n37 a_n2511_10156.n36 9.3005
R21165 a_n2511_10156.n10 a_n2511_10156.n9 9.3005
R21166 a_n2511_10156.n31 a_n2511_10156.n30 9.3005
R21167 a_n2511_10156.n29 a_n2511_10156.n28 9.3005
R21168 a_n2511_10156.n14 a_n2511_10156.n13 9.3005
R21169 a_n2511_10156.n23 a_n2511_10156.n22 9.3005
R21170 a_n2511_10156.n21 a_n2511_10156.n20 9.3005
R21171 a_n2511_10156.n134 a_n2511_10156.n109 8.92171
R21172 a_n2511_10156.n100 a_n2511_10156.n75 8.92171
R21173 a_n2511_10156.n68 a_n2511_10156.n43 8.92171
R21174 a_n2511_10156.n35 a_n2511_10156.n10 8.92171
R21175 a_n2511_10156.n135 a_n2511_10156.n107 8.14595
R21176 a_n2511_10156.n101 a_n2511_10156.n73 8.14595
R21177 a_n2511_10156.n69 a_n2511_10156.n41 8.14595
R21178 a_n2511_10156.n36 a_n2511_10156.n8 8.14595
R21179 a_n2511_10156.n139 a_n2511_10156.n138 5.91753
R21180 a_n2511_10156.n137 a_n2511_10156.n107 5.81868
R21181 a_n2511_10156.n103 a_n2511_10156.n73 5.81868
R21182 a_n2511_10156.n71 a_n2511_10156.n41 5.81868
R21183 a_n2511_10156.n38 a_n2511_10156.n8 5.81868
R21184 a_n2511_10156.n1 a_n2511_10156.t16 5.418
R21185 a_n2511_10156.n1 a_n2511_10156.t14 5.418
R21186 a_n2511_10156.n0 a_n2511_10156.t12 5.418
R21187 a_n2511_10156.n0 a_n2511_10156.t15 5.418
R21188 a_n2511_10156.n105 a_n2511_10156.t6 5.418
R21189 a_n2511_10156.n105 a_n2511_10156.t0 5.418
R21190 a_n2511_10156.n39 a_n2511_10156.t1 5.418
R21191 a_n2511_10156.n39 a_n2511_10156.t3 5.418
R21192 a_n2511_10156.n6 a_n2511_10156.t9 5.418
R21193 a_n2511_10156.n6 a_n2511_10156.t13 5.418
R21194 a_n2511_10156.n4 a_n2511_10156.t17 5.418
R21195 a_n2511_10156.n4 a_n2511_10156.t19 5.418
R21196 a_n2511_10156.n3 a_n2511_10156.t11 5.418
R21197 a_n2511_10156.n3 a_n2511_10156.t10 5.418
R21198 a_n2511_10156.t18 a_n2511_10156.n141 5.418
R21199 a_n2511_10156.n141 a_n2511_10156.t8 5.418
R21200 a_n2511_10156.n135 a_n2511_10156.n134 5.04292
R21201 a_n2511_10156.n101 a_n2511_10156.n100 5.04292
R21202 a_n2511_10156.n69 a_n2511_10156.n68 5.04292
R21203 a_n2511_10156.n36 a_n2511_10156.n35 5.04292
R21204 a_n2511_10156.n131 a_n2511_10156.n109 4.26717
R21205 a_n2511_10156.n97 a_n2511_10156.n75 4.26717
R21206 a_n2511_10156.n65 a_n2511_10156.n43 4.26717
R21207 a_n2511_10156.n32 a_n2511_10156.n10 4.26717
R21208 a_n2511_10156.n120 a_n2511_10156.n116 3.71286
R21209 a_n2511_10156.n86 a_n2511_10156.n82 3.71286
R21210 a_n2511_10156.n54 a_n2511_10156.n50 3.71286
R21211 a_n2511_10156.n21 a_n2511_10156.n17 3.71286
R21212 a_n2511_10156.n130 a_n2511_10156.n111 3.49141
R21213 a_n2511_10156.n96 a_n2511_10156.n77 3.49141
R21214 a_n2511_10156.n64 a_n2511_10156.n45 3.49141
R21215 a_n2511_10156.n31 a_n2511_10156.n12 3.49141
R21216 a_n2511_10156.n127 a_n2511_10156.n126 2.71565
R21217 a_n2511_10156.n93 a_n2511_10156.n92 2.71565
R21218 a_n2511_10156.n61 a_n2511_10156.n60 2.71565
R21219 a_n2511_10156.n28 a_n2511_10156.n27 2.71565
R21220 a_n2511_10156.n123 a_n2511_10156.n113 1.93989
R21221 a_n2511_10156.n89 a_n2511_10156.n79 1.93989
R21222 a_n2511_10156.n57 a_n2511_10156.n47 1.93989
R21223 a_n2511_10156.n24 a_n2511_10156.n14 1.93989
R21224 a_n2511_10156.n122 a_n2511_10156.n115 1.16414
R21225 a_n2511_10156.n88 a_n2511_10156.n81 1.16414
R21226 a_n2511_10156.n56 a_n2511_10156.n49 1.16414
R21227 a_n2511_10156.n23 a_n2511_10156.n16 1.16414
R21228 a_n2511_10156.n72 a_n2511_10156.n40 0.573776
R21229 a_n2511_10156.n106 a_n2511_10156.n104 0.573776
R21230 a_n2511_10156.n138 a_n2511_10156.n106 0.573776
R21231 a_n2511_10156.n140 a_n2511_10156.n2 0.573776
R21232 a_n2511_10156.n119 a_n2511_10156.n118 0.388379
R21233 a_n2511_10156.n85 a_n2511_10156.n84 0.388379
R21234 a_n2511_10156.n53 a_n2511_10156.n52 0.388379
R21235 a_n2511_10156.n20 a_n2511_10156.n19 0.388379
R21236 a_n2511_10156.n7 a_n2511_10156.n5 0.234655
R21237 a_n2511_10156.n136 a_n2511_10156.n108 0.155672
R21238 a_n2511_10156.n129 a_n2511_10156.n108 0.155672
R21239 a_n2511_10156.n129 a_n2511_10156.n128 0.155672
R21240 a_n2511_10156.n128 a_n2511_10156.n112 0.155672
R21241 a_n2511_10156.n121 a_n2511_10156.n112 0.155672
R21242 a_n2511_10156.n121 a_n2511_10156.n120 0.155672
R21243 a_n2511_10156.n102 a_n2511_10156.n74 0.155672
R21244 a_n2511_10156.n95 a_n2511_10156.n74 0.155672
R21245 a_n2511_10156.n95 a_n2511_10156.n94 0.155672
R21246 a_n2511_10156.n94 a_n2511_10156.n78 0.155672
R21247 a_n2511_10156.n87 a_n2511_10156.n78 0.155672
R21248 a_n2511_10156.n87 a_n2511_10156.n86 0.155672
R21249 a_n2511_10156.n70 a_n2511_10156.n42 0.155672
R21250 a_n2511_10156.n63 a_n2511_10156.n42 0.155672
R21251 a_n2511_10156.n63 a_n2511_10156.n62 0.155672
R21252 a_n2511_10156.n62 a_n2511_10156.n46 0.155672
R21253 a_n2511_10156.n55 a_n2511_10156.n46 0.155672
R21254 a_n2511_10156.n55 a_n2511_10156.n54 0.155672
R21255 a_n2511_10156.n37 a_n2511_10156.n9 0.155672
R21256 a_n2511_10156.n30 a_n2511_10156.n9 0.155672
R21257 a_n2511_10156.n30 a_n2511_10156.n29 0.155672
R21258 a_n2511_10156.n29 a_n2511_10156.n13 0.155672
R21259 a_n2511_10156.n22 a_n2511_10156.n13 0.155672
R21260 a_n2511_10156.n22 a_n2511_10156.n21 0.155672
R21261 a_n2511_10156.n104 a_n2511_10156.n72 0.155672
R21262 a_n2686_8022.n260 a_n2686_8022.n234 756.745
R21263 a_n2686_8022.n226 a_n2686_8022.n200 756.745
R21264 a_n2686_8022.n93 a_n2686_8022.n67 756.745
R21265 a_n2686_8022.n126 a_n2686_8022.n100 756.745
R21266 a_n2686_8022.n158 a_n2686_8022.n132 756.745
R21267 a_n2686_8022.n192 a_n2686_8022.n166 756.745
R21268 a_n2686_8022.n26 a_n2686_8022.n0 756.745
R21269 a_n2686_8022.n61 a_n2686_8022.n35 756.745
R21270 a_n2686_8022.n261 a_n2686_8022.n260 585
R21271 a_n2686_8022.n259 a_n2686_8022.n258 585
R21272 a_n2686_8022.n238 a_n2686_8022.n237 585
R21273 a_n2686_8022.n253 a_n2686_8022.n252 585
R21274 a_n2686_8022.n251 a_n2686_8022.n250 585
R21275 a_n2686_8022.n242 a_n2686_8022.n241 585
R21276 a_n2686_8022.n245 a_n2686_8022.n244 585
R21277 a_n2686_8022.n227 a_n2686_8022.n226 585
R21278 a_n2686_8022.n225 a_n2686_8022.n224 585
R21279 a_n2686_8022.n204 a_n2686_8022.n203 585
R21280 a_n2686_8022.n219 a_n2686_8022.n218 585
R21281 a_n2686_8022.n217 a_n2686_8022.n216 585
R21282 a_n2686_8022.n208 a_n2686_8022.n207 585
R21283 a_n2686_8022.n211 a_n2686_8022.n210 585
R21284 a_n2686_8022.n94 a_n2686_8022.n93 585
R21285 a_n2686_8022.n92 a_n2686_8022.n91 585
R21286 a_n2686_8022.n71 a_n2686_8022.n70 585
R21287 a_n2686_8022.n86 a_n2686_8022.n85 585
R21288 a_n2686_8022.n84 a_n2686_8022.n83 585
R21289 a_n2686_8022.n75 a_n2686_8022.n74 585
R21290 a_n2686_8022.n78 a_n2686_8022.n77 585
R21291 a_n2686_8022.n127 a_n2686_8022.n126 585
R21292 a_n2686_8022.n125 a_n2686_8022.n124 585
R21293 a_n2686_8022.n104 a_n2686_8022.n103 585
R21294 a_n2686_8022.n119 a_n2686_8022.n118 585
R21295 a_n2686_8022.n117 a_n2686_8022.n116 585
R21296 a_n2686_8022.n108 a_n2686_8022.n107 585
R21297 a_n2686_8022.n111 a_n2686_8022.n110 585
R21298 a_n2686_8022.n159 a_n2686_8022.n158 585
R21299 a_n2686_8022.n157 a_n2686_8022.n156 585
R21300 a_n2686_8022.n136 a_n2686_8022.n135 585
R21301 a_n2686_8022.n151 a_n2686_8022.n150 585
R21302 a_n2686_8022.n149 a_n2686_8022.n148 585
R21303 a_n2686_8022.n140 a_n2686_8022.n139 585
R21304 a_n2686_8022.n143 a_n2686_8022.n142 585
R21305 a_n2686_8022.n193 a_n2686_8022.n192 585
R21306 a_n2686_8022.n191 a_n2686_8022.n190 585
R21307 a_n2686_8022.n170 a_n2686_8022.n169 585
R21308 a_n2686_8022.n185 a_n2686_8022.n184 585
R21309 a_n2686_8022.n183 a_n2686_8022.n182 585
R21310 a_n2686_8022.n174 a_n2686_8022.n173 585
R21311 a_n2686_8022.n177 a_n2686_8022.n176 585
R21312 a_n2686_8022.n27 a_n2686_8022.n26 585
R21313 a_n2686_8022.n25 a_n2686_8022.n24 585
R21314 a_n2686_8022.n4 a_n2686_8022.n3 585
R21315 a_n2686_8022.n19 a_n2686_8022.n18 585
R21316 a_n2686_8022.n17 a_n2686_8022.n16 585
R21317 a_n2686_8022.n8 a_n2686_8022.n7 585
R21318 a_n2686_8022.n11 a_n2686_8022.n10 585
R21319 a_n2686_8022.n62 a_n2686_8022.n61 585
R21320 a_n2686_8022.n60 a_n2686_8022.n59 585
R21321 a_n2686_8022.n39 a_n2686_8022.n38 585
R21322 a_n2686_8022.n54 a_n2686_8022.n53 585
R21323 a_n2686_8022.n52 a_n2686_8022.n51 585
R21324 a_n2686_8022.n43 a_n2686_8022.n42 585
R21325 a_n2686_8022.n46 a_n2686_8022.n45 585
R21326 a_n2686_8022.t9 a_n2686_8022.n243 327.601
R21327 a_n2686_8022.t2 a_n2686_8022.n209 327.601
R21328 a_n2686_8022.t17 a_n2686_8022.n76 327.601
R21329 a_n2686_8022.t20 a_n2686_8022.n109 327.601
R21330 a_n2686_8022.t16 a_n2686_8022.n141 327.601
R21331 a_n2686_8022.t18 a_n2686_8022.n175 327.601
R21332 a_n2686_8022.t7 a_n2686_8022.n9 327.601
R21333 a_n2686_8022.t8 a_n2686_8022.n44 327.601
R21334 a_n2686_8022.n260 a_n2686_8022.n259 171.744
R21335 a_n2686_8022.n259 a_n2686_8022.n237 171.744
R21336 a_n2686_8022.n252 a_n2686_8022.n237 171.744
R21337 a_n2686_8022.n252 a_n2686_8022.n251 171.744
R21338 a_n2686_8022.n251 a_n2686_8022.n241 171.744
R21339 a_n2686_8022.n244 a_n2686_8022.n241 171.744
R21340 a_n2686_8022.n226 a_n2686_8022.n225 171.744
R21341 a_n2686_8022.n225 a_n2686_8022.n203 171.744
R21342 a_n2686_8022.n218 a_n2686_8022.n203 171.744
R21343 a_n2686_8022.n218 a_n2686_8022.n217 171.744
R21344 a_n2686_8022.n217 a_n2686_8022.n207 171.744
R21345 a_n2686_8022.n210 a_n2686_8022.n207 171.744
R21346 a_n2686_8022.n93 a_n2686_8022.n92 171.744
R21347 a_n2686_8022.n92 a_n2686_8022.n70 171.744
R21348 a_n2686_8022.n85 a_n2686_8022.n70 171.744
R21349 a_n2686_8022.n85 a_n2686_8022.n84 171.744
R21350 a_n2686_8022.n84 a_n2686_8022.n74 171.744
R21351 a_n2686_8022.n77 a_n2686_8022.n74 171.744
R21352 a_n2686_8022.n126 a_n2686_8022.n125 171.744
R21353 a_n2686_8022.n125 a_n2686_8022.n103 171.744
R21354 a_n2686_8022.n118 a_n2686_8022.n103 171.744
R21355 a_n2686_8022.n118 a_n2686_8022.n117 171.744
R21356 a_n2686_8022.n117 a_n2686_8022.n107 171.744
R21357 a_n2686_8022.n110 a_n2686_8022.n107 171.744
R21358 a_n2686_8022.n158 a_n2686_8022.n157 171.744
R21359 a_n2686_8022.n157 a_n2686_8022.n135 171.744
R21360 a_n2686_8022.n150 a_n2686_8022.n135 171.744
R21361 a_n2686_8022.n150 a_n2686_8022.n149 171.744
R21362 a_n2686_8022.n149 a_n2686_8022.n139 171.744
R21363 a_n2686_8022.n142 a_n2686_8022.n139 171.744
R21364 a_n2686_8022.n192 a_n2686_8022.n191 171.744
R21365 a_n2686_8022.n191 a_n2686_8022.n169 171.744
R21366 a_n2686_8022.n184 a_n2686_8022.n169 171.744
R21367 a_n2686_8022.n184 a_n2686_8022.n183 171.744
R21368 a_n2686_8022.n183 a_n2686_8022.n173 171.744
R21369 a_n2686_8022.n176 a_n2686_8022.n173 171.744
R21370 a_n2686_8022.n26 a_n2686_8022.n25 171.744
R21371 a_n2686_8022.n25 a_n2686_8022.n3 171.744
R21372 a_n2686_8022.n18 a_n2686_8022.n3 171.744
R21373 a_n2686_8022.n18 a_n2686_8022.n17 171.744
R21374 a_n2686_8022.n17 a_n2686_8022.n7 171.744
R21375 a_n2686_8022.n10 a_n2686_8022.n7 171.744
R21376 a_n2686_8022.n61 a_n2686_8022.n60 171.744
R21377 a_n2686_8022.n60 a_n2686_8022.n38 171.744
R21378 a_n2686_8022.n53 a_n2686_8022.n38 171.744
R21379 a_n2686_8022.n53 a_n2686_8022.n52 171.744
R21380 a_n2686_8022.n52 a_n2686_8022.n42 171.744
R21381 a_n2686_8022.n45 a_n2686_8022.n42 171.744
R21382 a_n2686_8022.n244 a_n2686_8022.t9 85.8723
R21383 a_n2686_8022.n210 a_n2686_8022.t2 85.8723
R21384 a_n2686_8022.n77 a_n2686_8022.t17 85.8723
R21385 a_n2686_8022.n110 a_n2686_8022.t20 85.8723
R21386 a_n2686_8022.n142 a_n2686_8022.t16 85.8723
R21387 a_n2686_8022.n176 a_n2686_8022.t18 85.8723
R21388 a_n2686_8022.n10 a_n2686_8022.t7 85.8723
R21389 a_n2686_8022.n45 a_n2686_8022.t8 85.8723
R21390 a_n2686_8022.n233 a_n2686_8022.n232 81.2397
R21391 a_n2686_8022.n99 a_n2686_8022.n98 81.2397
R21392 a_n2686_8022.n165 a_n2686_8022.n164 81.2397
R21393 a_n2686_8022.n32 a_n2686_8022.n31 81.2397
R21394 a_n2686_8022.n34 a_n2686_8022.n33 81.2397
R21395 a_n2686_8022.n266 a_n2686_8022.n265 81.2397
R21396 a_n2686_8022.n265 a_n2686_8022.n264 38.3829
R21397 a_n2686_8022.n99 a_n2686_8022.n97 38.3829
R21398 a_n2686_8022.n32 a_n2686_8022.n30 38.3829
R21399 a_n2686_8022.n231 a_n2686_8022.n230 37.8096
R21400 a_n2686_8022.n131 a_n2686_8022.n130 37.8096
R21401 a_n2686_8022.n163 a_n2686_8022.n162 37.8096
R21402 a_n2686_8022.n197 a_n2686_8022.n196 37.8096
R21403 a_n2686_8022.n66 a_n2686_8022.n65 37.8096
R21404 a_n2686_8022.n198 a_n2686_8022.n66 22.3736
R21405 a_n2686_8022.n245 a_n2686_8022.n243 16.3865
R21406 a_n2686_8022.n211 a_n2686_8022.n209 16.3865
R21407 a_n2686_8022.n78 a_n2686_8022.n76 16.3865
R21408 a_n2686_8022.n111 a_n2686_8022.n109 16.3865
R21409 a_n2686_8022.n143 a_n2686_8022.n141 16.3865
R21410 a_n2686_8022.n177 a_n2686_8022.n175 16.3865
R21411 a_n2686_8022.n11 a_n2686_8022.n9 16.3865
R21412 a_n2686_8022.n46 a_n2686_8022.n44 16.3865
R21413 a_n2686_8022.n246 a_n2686_8022.n242 12.8005
R21414 a_n2686_8022.n212 a_n2686_8022.n208 12.8005
R21415 a_n2686_8022.n79 a_n2686_8022.n75 12.8005
R21416 a_n2686_8022.n112 a_n2686_8022.n108 12.8005
R21417 a_n2686_8022.n144 a_n2686_8022.n140 12.8005
R21418 a_n2686_8022.n178 a_n2686_8022.n174 12.8005
R21419 a_n2686_8022.n12 a_n2686_8022.n8 12.8005
R21420 a_n2686_8022.n47 a_n2686_8022.n43 12.8005
R21421 a_n2686_8022.n250 a_n2686_8022.n249 12.0247
R21422 a_n2686_8022.n216 a_n2686_8022.n215 12.0247
R21423 a_n2686_8022.n83 a_n2686_8022.n82 12.0247
R21424 a_n2686_8022.n116 a_n2686_8022.n115 12.0247
R21425 a_n2686_8022.n148 a_n2686_8022.n147 12.0247
R21426 a_n2686_8022.n182 a_n2686_8022.n181 12.0247
R21427 a_n2686_8022.n16 a_n2686_8022.n15 12.0247
R21428 a_n2686_8022.n51 a_n2686_8022.n50 12.0247
R21429 a_n2686_8022.n253 a_n2686_8022.n240 11.249
R21430 a_n2686_8022.n219 a_n2686_8022.n206 11.249
R21431 a_n2686_8022.n86 a_n2686_8022.n73 11.249
R21432 a_n2686_8022.n119 a_n2686_8022.n106 11.249
R21433 a_n2686_8022.n151 a_n2686_8022.n138 11.249
R21434 a_n2686_8022.n185 a_n2686_8022.n172 11.249
R21435 a_n2686_8022.n19 a_n2686_8022.n6 11.249
R21436 a_n2686_8022.n54 a_n2686_8022.n41 11.249
R21437 a_n2686_8022.n254 a_n2686_8022.n238 10.4732
R21438 a_n2686_8022.n220 a_n2686_8022.n204 10.4732
R21439 a_n2686_8022.n87 a_n2686_8022.n71 10.4732
R21440 a_n2686_8022.n120 a_n2686_8022.n104 10.4732
R21441 a_n2686_8022.n152 a_n2686_8022.n136 10.4732
R21442 a_n2686_8022.n186 a_n2686_8022.n170 10.4732
R21443 a_n2686_8022.n20 a_n2686_8022.n4 10.4732
R21444 a_n2686_8022.n55 a_n2686_8022.n39 10.4732
R21445 a_n2686_8022.n258 a_n2686_8022.n257 9.69747
R21446 a_n2686_8022.n224 a_n2686_8022.n223 9.69747
R21447 a_n2686_8022.n91 a_n2686_8022.n90 9.69747
R21448 a_n2686_8022.n124 a_n2686_8022.n123 9.69747
R21449 a_n2686_8022.n156 a_n2686_8022.n155 9.69747
R21450 a_n2686_8022.n190 a_n2686_8022.n189 9.69747
R21451 a_n2686_8022.n24 a_n2686_8022.n23 9.69747
R21452 a_n2686_8022.n59 a_n2686_8022.n58 9.69747
R21453 a_n2686_8022.n264 a_n2686_8022.n263 9.45567
R21454 a_n2686_8022.n230 a_n2686_8022.n229 9.45567
R21455 a_n2686_8022.n97 a_n2686_8022.n96 9.45567
R21456 a_n2686_8022.n130 a_n2686_8022.n129 9.45567
R21457 a_n2686_8022.n162 a_n2686_8022.n161 9.45567
R21458 a_n2686_8022.n196 a_n2686_8022.n195 9.45567
R21459 a_n2686_8022.n30 a_n2686_8022.n29 9.45567
R21460 a_n2686_8022.n65 a_n2686_8022.n64 9.45567
R21461 a_n2686_8022.n263 a_n2686_8022.n262 9.3005
R21462 a_n2686_8022.n236 a_n2686_8022.n235 9.3005
R21463 a_n2686_8022.n257 a_n2686_8022.n256 9.3005
R21464 a_n2686_8022.n255 a_n2686_8022.n254 9.3005
R21465 a_n2686_8022.n240 a_n2686_8022.n239 9.3005
R21466 a_n2686_8022.n249 a_n2686_8022.n248 9.3005
R21467 a_n2686_8022.n247 a_n2686_8022.n246 9.3005
R21468 a_n2686_8022.n229 a_n2686_8022.n228 9.3005
R21469 a_n2686_8022.n202 a_n2686_8022.n201 9.3005
R21470 a_n2686_8022.n223 a_n2686_8022.n222 9.3005
R21471 a_n2686_8022.n221 a_n2686_8022.n220 9.3005
R21472 a_n2686_8022.n206 a_n2686_8022.n205 9.3005
R21473 a_n2686_8022.n215 a_n2686_8022.n214 9.3005
R21474 a_n2686_8022.n213 a_n2686_8022.n212 9.3005
R21475 a_n2686_8022.n96 a_n2686_8022.n95 9.3005
R21476 a_n2686_8022.n69 a_n2686_8022.n68 9.3005
R21477 a_n2686_8022.n90 a_n2686_8022.n89 9.3005
R21478 a_n2686_8022.n88 a_n2686_8022.n87 9.3005
R21479 a_n2686_8022.n73 a_n2686_8022.n72 9.3005
R21480 a_n2686_8022.n82 a_n2686_8022.n81 9.3005
R21481 a_n2686_8022.n80 a_n2686_8022.n79 9.3005
R21482 a_n2686_8022.n129 a_n2686_8022.n128 9.3005
R21483 a_n2686_8022.n102 a_n2686_8022.n101 9.3005
R21484 a_n2686_8022.n123 a_n2686_8022.n122 9.3005
R21485 a_n2686_8022.n121 a_n2686_8022.n120 9.3005
R21486 a_n2686_8022.n106 a_n2686_8022.n105 9.3005
R21487 a_n2686_8022.n115 a_n2686_8022.n114 9.3005
R21488 a_n2686_8022.n113 a_n2686_8022.n112 9.3005
R21489 a_n2686_8022.n161 a_n2686_8022.n160 9.3005
R21490 a_n2686_8022.n134 a_n2686_8022.n133 9.3005
R21491 a_n2686_8022.n155 a_n2686_8022.n154 9.3005
R21492 a_n2686_8022.n153 a_n2686_8022.n152 9.3005
R21493 a_n2686_8022.n138 a_n2686_8022.n137 9.3005
R21494 a_n2686_8022.n147 a_n2686_8022.n146 9.3005
R21495 a_n2686_8022.n145 a_n2686_8022.n144 9.3005
R21496 a_n2686_8022.n195 a_n2686_8022.n194 9.3005
R21497 a_n2686_8022.n168 a_n2686_8022.n167 9.3005
R21498 a_n2686_8022.n189 a_n2686_8022.n188 9.3005
R21499 a_n2686_8022.n187 a_n2686_8022.n186 9.3005
R21500 a_n2686_8022.n172 a_n2686_8022.n171 9.3005
R21501 a_n2686_8022.n181 a_n2686_8022.n180 9.3005
R21502 a_n2686_8022.n179 a_n2686_8022.n178 9.3005
R21503 a_n2686_8022.n29 a_n2686_8022.n28 9.3005
R21504 a_n2686_8022.n2 a_n2686_8022.n1 9.3005
R21505 a_n2686_8022.n23 a_n2686_8022.n22 9.3005
R21506 a_n2686_8022.n21 a_n2686_8022.n20 9.3005
R21507 a_n2686_8022.n6 a_n2686_8022.n5 9.3005
R21508 a_n2686_8022.n15 a_n2686_8022.n14 9.3005
R21509 a_n2686_8022.n13 a_n2686_8022.n12 9.3005
R21510 a_n2686_8022.n64 a_n2686_8022.n63 9.3005
R21511 a_n2686_8022.n37 a_n2686_8022.n36 9.3005
R21512 a_n2686_8022.n58 a_n2686_8022.n57 9.3005
R21513 a_n2686_8022.n56 a_n2686_8022.n55 9.3005
R21514 a_n2686_8022.n41 a_n2686_8022.n40 9.3005
R21515 a_n2686_8022.n50 a_n2686_8022.n49 9.3005
R21516 a_n2686_8022.n48 a_n2686_8022.n47 9.3005
R21517 a_n2686_8022.n261 a_n2686_8022.n236 8.92171
R21518 a_n2686_8022.n227 a_n2686_8022.n202 8.92171
R21519 a_n2686_8022.n94 a_n2686_8022.n69 8.92171
R21520 a_n2686_8022.n127 a_n2686_8022.n102 8.92171
R21521 a_n2686_8022.n159 a_n2686_8022.n134 8.92171
R21522 a_n2686_8022.n193 a_n2686_8022.n168 8.92171
R21523 a_n2686_8022.n27 a_n2686_8022.n2 8.92171
R21524 a_n2686_8022.n62 a_n2686_8022.n37 8.92171
R21525 a_n2686_8022.n199 a_n2686_8022.t0 8.43517
R21526 a_n2686_8022.n262 a_n2686_8022.n234 8.14595
R21527 a_n2686_8022.n228 a_n2686_8022.n200 8.14595
R21528 a_n2686_8022.n95 a_n2686_8022.n67 8.14595
R21529 a_n2686_8022.n128 a_n2686_8022.n100 8.14595
R21530 a_n2686_8022.n160 a_n2686_8022.n132 8.14595
R21531 a_n2686_8022.n194 a_n2686_8022.n166 8.14595
R21532 a_n2686_8022.n28 a_n2686_8022.n0 8.14595
R21533 a_n2686_8022.n63 a_n2686_8022.n35 8.14595
R21534 a_n2686_8022.n198 a_n2686_8022.n197 5.91753
R21535 a_n2686_8022.n264 a_n2686_8022.n234 5.81868
R21536 a_n2686_8022.n230 a_n2686_8022.n200 5.81868
R21537 a_n2686_8022.n97 a_n2686_8022.n67 5.81868
R21538 a_n2686_8022.n130 a_n2686_8022.n100 5.81868
R21539 a_n2686_8022.n162 a_n2686_8022.n132 5.81868
R21540 a_n2686_8022.n196 a_n2686_8022.n166 5.81868
R21541 a_n2686_8022.n30 a_n2686_8022.n0 5.81868
R21542 a_n2686_8022.n65 a_n2686_8022.n35 5.81868
R21543 a_n2686_8022.n231 a_n2686_8022.n199 5.72895
R21544 a_n2686_8022.n232 a_n2686_8022.t1 5.418
R21545 a_n2686_8022.n232 a_n2686_8022.t11 5.418
R21546 a_n2686_8022.n98 a_n2686_8022.t15 5.418
R21547 a_n2686_8022.n98 a_n2686_8022.t13 5.418
R21548 a_n2686_8022.n164 a_n2686_8022.t14 5.418
R21549 a_n2686_8022.n164 a_n2686_8022.t19 5.418
R21550 a_n2686_8022.n31 a_n2686_8022.t10 5.418
R21551 a_n2686_8022.n31 a_n2686_8022.t6 5.418
R21552 a_n2686_8022.n33 a_n2686_8022.t4 5.418
R21553 a_n2686_8022.n33 a_n2686_8022.t5 5.418
R21554 a_n2686_8022.n266 a_n2686_8022.t3 5.418
R21555 a_n2686_8022.t12 a_n2686_8022.n266 5.418
R21556 a_n2686_8022.n262 a_n2686_8022.n261 5.04292
R21557 a_n2686_8022.n228 a_n2686_8022.n227 5.04292
R21558 a_n2686_8022.n95 a_n2686_8022.n94 5.04292
R21559 a_n2686_8022.n128 a_n2686_8022.n127 5.04292
R21560 a_n2686_8022.n160 a_n2686_8022.n159 5.04292
R21561 a_n2686_8022.n194 a_n2686_8022.n193 5.04292
R21562 a_n2686_8022.n28 a_n2686_8022.n27 5.04292
R21563 a_n2686_8022.n63 a_n2686_8022.n62 5.04292
R21564 a_n2686_8022.n258 a_n2686_8022.n236 4.26717
R21565 a_n2686_8022.n224 a_n2686_8022.n202 4.26717
R21566 a_n2686_8022.n91 a_n2686_8022.n69 4.26717
R21567 a_n2686_8022.n124 a_n2686_8022.n102 4.26717
R21568 a_n2686_8022.n156 a_n2686_8022.n134 4.26717
R21569 a_n2686_8022.n190 a_n2686_8022.n168 4.26717
R21570 a_n2686_8022.n24 a_n2686_8022.n2 4.26717
R21571 a_n2686_8022.n59 a_n2686_8022.n37 4.26717
R21572 a_n2686_8022.n199 a_n2686_8022.n198 4.20883
R21573 a_n2686_8022.n247 a_n2686_8022.n243 3.71286
R21574 a_n2686_8022.n213 a_n2686_8022.n209 3.71286
R21575 a_n2686_8022.n80 a_n2686_8022.n76 3.71286
R21576 a_n2686_8022.n113 a_n2686_8022.n109 3.71286
R21577 a_n2686_8022.n145 a_n2686_8022.n141 3.71286
R21578 a_n2686_8022.n179 a_n2686_8022.n175 3.71286
R21579 a_n2686_8022.n13 a_n2686_8022.n9 3.71286
R21580 a_n2686_8022.n48 a_n2686_8022.n44 3.71286
R21581 a_n2686_8022.n257 a_n2686_8022.n238 3.49141
R21582 a_n2686_8022.n223 a_n2686_8022.n204 3.49141
R21583 a_n2686_8022.n90 a_n2686_8022.n71 3.49141
R21584 a_n2686_8022.n123 a_n2686_8022.n104 3.49141
R21585 a_n2686_8022.n155 a_n2686_8022.n136 3.49141
R21586 a_n2686_8022.n189 a_n2686_8022.n170 3.49141
R21587 a_n2686_8022.n23 a_n2686_8022.n4 3.49141
R21588 a_n2686_8022.n58 a_n2686_8022.n39 3.49141
R21589 a_n2686_8022.n254 a_n2686_8022.n253 2.71565
R21590 a_n2686_8022.n220 a_n2686_8022.n219 2.71565
R21591 a_n2686_8022.n87 a_n2686_8022.n86 2.71565
R21592 a_n2686_8022.n120 a_n2686_8022.n119 2.71565
R21593 a_n2686_8022.n152 a_n2686_8022.n151 2.71565
R21594 a_n2686_8022.n186 a_n2686_8022.n185 2.71565
R21595 a_n2686_8022.n20 a_n2686_8022.n19 2.71565
R21596 a_n2686_8022.n55 a_n2686_8022.n54 2.71565
R21597 a_n2686_8022.n250 a_n2686_8022.n240 1.93989
R21598 a_n2686_8022.n216 a_n2686_8022.n206 1.93989
R21599 a_n2686_8022.n83 a_n2686_8022.n73 1.93989
R21600 a_n2686_8022.n116 a_n2686_8022.n106 1.93989
R21601 a_n2686_8022.n148 a_n2686_8022.n138 1.93989
R21602 a_n2686_8022.n182 a_n2686_8022.n172 1.93989
R21603 a_n2686_8022.n16 a_n2686_8022.n6 1.93989
R21604 a_n2686_8022.n51 a_n2686_8022.n41 1.93989
R21605 a_n2686_8022.n249 a_n2686_8022.n242 1.16414
R21606 a_n2686_8022.n215 a_n2686_8022.n208 1.16414
R21607 a_n2686_8022.n82 a_n2686_8022.n75 1.16414
R21608 a_n2686_8022.n115 a_n2686_8022.n108 1.16414
R21609 a_n2686_8022.n147 a_n2686_8022.n140 1.16414
R21610 a_n2686_8022.n181 a_n2686_8022.n174 1.16414
R21611 a_n2686_8022.n15 a_n2686_8022.n8 1.16414
R21612 a_n2686_8022.n50 a_n2686_8022.n43 1.16414
R21613 a_n2686_8022.n197 a_n2686_8022.n165 0.573776
R21614 a_n2686_8022.n165 a_n2686_8022.n163 0.573776
R21615 a_n2686_8022.n131 a_n2686_8022.n99 0.573776
R21616 a_n2686_8022.n66 a_n2686_8022.n34 0.573776
R21617 a_n2686_8022.n34 a_n2686_8022.n32 0.573776
R21618 a_n2686_8022.n233 a_n2686_8022.n231 0.573776
R21619 a_n2686_8022.n265 a_n2686_8022.n233 0.573776
R21620 a_n2686_8022.n246 a_n2686_8022.n245 0.388379
R21621 a_n2686_8022.n212 a_n2686_8022.n211 0.388379
R21622 a_n2686_8022.n79 a_n2686_8022.n78 0.388379
R21623 a_n2686_8022.n112 a_n2686_8022.n111 0.388379
R21624 a_n2686_8022.n144 a_n2686_8022.n143 0.388379
R21625 a_n2686_8022.n178 a_n2686_8022.n177 0.388379
R21626 a_n2686_8022.n12 a_n2686_8022.n11 0.388379
R21627 a_n2686_8022.n47 a_n2686_8022.n46 0.388379
R21628 a_n2686_8022.n263 a_n2686_8022.n235 0.155672
R21629 a_n2686_8022.n256 a_n2686_8022.n235 0.155672
R21630 a_n2686_8022.n256 a_n2686_8022.n255 0.155672
R21631 a_n2686_8022.n255 a_n2686_8022.n239 0.155672
R21632 a_n2686_8022.n248 a_n2686_8022.n239 0.155672
R21633 a_n2686_8022.n248 a_n2686_8022.n247 0.155672
R21634 a_n2686_8022.n229 a_n2686_8022.n201 0.155672
R21635 a_n2686_8022.n222 a_n2686_8022.n201 0.155672
R21636 a_n2686_8022.n222 a_n2686_8022.n221 0.155672
R21637 a_n2686_8022.n221 a_n2686_8022.n205 0.155672
R21638 a_n2686_8022.n214 a_n2686_8022.n205 0.155672
R21639 a_n2686_8022.n214 a_n2686_8022.n213 0.155672
R21640 a_n2686_8022.n96 a_n2686_8022.n68 0.155672
R21641 a_n2686_8022.n89 a_n2686_8022.n68 0.155672
R21642 a_n2686_8022.n89 a_n2686_8022.n88 0.155672
R21643 a_n2686_8022.n88 a_n2686_8022.n72 0.155672
R21644 a_n2686_8022.n81 a_n2686_8022.n72 0.155672
R21645 a_n2686_8022.n81 a_n2686_8022.n80 0.155672
R21646 a_n2686_8022.n129 a_n2686_8022.n101 0.155672
R21647 a_n2686_8022.n122 a_n2686_8022.n101 0.155672
R21648 a_n2686_8022.n122 a_n2686_8022.n121 0.155672
R21649 a_n2686_8022.n121 a_n2686_8022.n105 0.155672
R21650 a_n2686_8022.n114 a_n2686_8022.n105 0.155672
R21651 a_n2686_8022.n114 a_n2686_8022.n113 0.155672
R21652 a_n2686_8022.n161 a_n2686_8022.n133 0.155672
R21653 a_n2686_8022.n154 a_n2686_8022.n133 0.155672
R21654 a_n2686_8022.n154 a_n2686_8022.n153 0.155672
R21655 a_n2686_8022.n153 a_n2686_8022.n137 0.155672
R21656 a_n2686_8022.n146 a_n2686_8022.n137 0.155672
R21657 a_n2686_8022.n146 a_n2686_8022.n145 0.155672
R21658 a_n2686_8022.n195 a_n2686_8022.n167 0.155672
R21659 a_n2686_8022.n188 a_n2686_8022.n167 0.155672
R21660 a_n2686_8022.n188 a_n2686_8022.n187 0.155672
R21661 a_n2686_8022.n187 a_n2686_8022.n171 0.155672
R21662 a_n2686_8022.n180 a_n2686_8022.n171 0.155672
R21663 a_n2686_8022.n180 a_n2686_8022.n179 0.155672
R21664 a_n2686_8022.n163 a_n2686_8022.n131 0.155672
R21665 a_n2686_8022.n29 a_n2686_8022.n1 0.155672
R21666 a_n2686_8022.n22 a_n2686_8022.n1 0.155672
R21667 a_n2686_8022.n22 a_n2686_8022.n21 0.155672
R21668 a_n2686_8022.n21 a_n2686_8022.n5 0.155672
R21669 a_n2686_8022.n14 a_n2686_8022.n5 0.155672
R21670 a_n2686_8022.n14 a_n2686_8022.n13 0.155672
R21671 a_n2686_8022.n64 a_n2686_8022.n36 0.155672
R21672 a_n2686_8022.n57 a_n2686_8022.n36 0.155672
R21673 a_n2686_8022.n57 a_n2686_8022.n56 0.155672
R21674 a_n2686_8022.n56 a_n2686_8022.n40 0.155672
R21675 a_n2686_8022.n49 a_n2686_8022.n40 0.155672
R21676 a_n2686_8022.n49 a_n2686_8022.n48 0.155672
R21677 output.n41 output.n15 289.615
R21678 output.n72 output.n46 289.615
R21679 output.n104 output.n78 289.615
R21680 output.n136 output.n110 289.615
R21681 output.n77 output.n45 197.26
R21682 output.n77 output.n76 196.298
R21683 output.n109 output.n108 196.298
R21684 output.n141 output.n140 196.298
R21685 output.n42 output.n41 185
R21686 output.n40 output.n39 185
R21687 output.n19 output.n18 185
R21688 output.n34 output.n33 185
R21689 output.n32 output.n31 185
R21690 output.n23 output.n22 185
R21691 output.n26 output.n25 185
R21692 output.n73 output.n72 185
R21693 output.n71 output.n70 185
R21694 output.n50 output.n49 185
R21695 output.n65 output.n64 185
R21696 output.n63 output.n62 185
R21697 output.n54 output.n53 185
R21698 output.n57 output.n56 185
R21699 output.n105 output.n104 185
R21700 output.n103 output.n102 185
R21701 output.n82 output.n81 185
R21702 output.n97 output.n96 185
R21703 output.n95 output.n94 185
R21704 output.n86 output.n85 185
R21705 output.n89 output.n88 185
R21706 output.n137 output.n136 185
R21707 output.n135 output.n134 185
R21708 output.n114 output.n113 185
R21709 output.n129 output.n128 185
R21710 output.n127 output.n126 185
R21711 output.n118 output.n117 185
R21712 output.n121 output.n120 185
R21713 output.t19 output.n24 147.661
R21714 output.t18 output.n55 147.661
R21715 output.t17 output.n87 147.661
R21716 output.t16 output.n119 147.661
R21717 output.n41 output.n40 104.615
R21718 output.n40 output.n18 104.615
R21719 output.n33 output.n18 104.615
R21720 output.n33 output.n32 104.615
R21721 output.n32 output.n22 104.615
R21722 output.n25 output.n22 104.615
R21723 output.n72 output.n71 104.615
R21724 output.n71 output.n49 104.615
R21725 output.n64 output.n49 104.615
R21726 output.n64 output.n63 104.615
R21727 output.n63 output.n53 104.615
R21728 output.n56 output.n53 104.615
R21729 output.n104 output.n103 104.615
R21730 output.n103 output.n81 104.615
R21731 output.n96 output.n81 104.615
R21732 output.n96 output.n95 104.615
R21733 output.n95 output.n85 104.615
R21734 output.n88 output.n85 104.615
R21735 output.n136 output.n135 104.615
R21736 output.n135 output.n113 104.615
R21737 output.n128 output.n113 104.615
R21738 output.n128 output.n127 104.615
R21739 output.n127 output.n117 104.615
R21740 output.n120 output.n117 104.615
R21741 output.n1 output.t13 77.056
R21742 output.n14 output.t14 76.6694
R21743 output.n1 output.n0 72.7095
R21744 output.n3 output.n2 72.7095
R21745 output.n5 output.n4 72.7095
R21746 output.n7 output.n6 72.7095
R21747 output.n9 output.n8 72.7095
R21748 output.n11 output.n10 72.7095
R21749 output.n13 output.n12 72.7095
R21750 output.n25 output.t19 52.3082
R21751 output.n56 output.t18 52.3082
R21752 output.n88 output.t17 52.3082
R21753 output.n120 output.t16 52.3082
R21754 output.n26 output.n24 15.6674
R21755 output.n57 output.n55 15.6674
R21756 output.n89 output.n87 15.6674
R21757 output.n121 output.n119 15.6674
R21758 output.n27 output.n23 12.8005
R21759 output.n58 output.n54 12.8005
R21760 output.n90 output.n86 12.8005
R21761 output.n122 output.n118 12.8005
R21762 output.n31 output.n30 12.0247
R21763 output.n62 output.n61 12.0247
R21764 output.n94 output.n93 12.0247
R21765 output.n126 output.n125 12.0247
R21766 output.n34 output.n21 11.249
R21767 output.n65 output.n52 11.249
R21768 output.n97 output.n84 11.249
R21769 output.n129 output.n116 11.249
R21770 output.n35 output.n19 10.4732
R21771 output.n66 output.n50 10.4732
R21772 output.n98 output.n82 10.4732
R21773 output.n130 output.n114 10.4732
R21774 output.n39 output.n38 9.69747
R21775 output.n70 output.n69 9.69747
R21776 output.n102 output.n101 9.69747
R21777 output.n134 output.n133 9.69747
R21778 output.n45 output.n44 9.45567
R21779 output.n76 output.n75 9.45567
R21780 output.n108 output.n107 9.45567
R21781 output.n140 output.n139 9.45567
R21782 output.n44 output.n43 9.3005
R21783 output.n17 output.n16 9.3005
R21784 output.n38 output.n37 9.3005
R21785 output.n36 output.n35 9.3005
R21786 output.n21 output.n20 9.3005
R21787 output.n30 output.n29 9.3005
R21788 output.n28 output.n27 9.3005
R21789 output.n75 output.n74 9.3005
R21790 output.n48 output.n47 9.3005
R21791 output.n69 output.n68 9.3005
R21792 output.n67 output.n66 9.3005
R21793 output.n52 output.n51 9.3005
R21794 output.n61 output.n60 9.3005
R21795 output.n59 output.n58 9.3005
R21796 output.n107 output.n106 9.3005
R21797 output.n80 output.n79 9.3005
R21798 output.n101 output.n100 9.3005
R21799 output.n99 output.n98 9.3005
R21800 output.n84 output.n83 9.3005
R21801 output.n93 output.n92 9.3005
R21802 output.n91 output.n90 9.3005
R21803 output.n139 output.n138 9.3005
R21804 output.n112 output.n111 9.3005
R21805 output.n133 output.n132 9.3005
R21806 output.n131 output.n130 9.3005
R21807 output.n116 output.n115 9.3005
R21808 output.n125 output.n124 9.3005
R21809 output.n123 output.n122 9.3005
R21810 output.n42 output.n17 8.92171
R21811 output.n73 output.n48 8.92171
R21812 output.n105 output.n80 8.92171
R21813 output.n137 output.n112 8.92171
R21814 output output.n141 8.15037
R21815 output.n43 output.n15 8.14595
R21816 output.n74 output.n46 8.14595
R21817 output.n106 output.n78 8.14595
R21818 output.n138 output.n110 8.14595
R21819 output.n45 output.n15 5.81868
R21820 output.n76 output.n46 5.81868
R21821 output.n108 output.n78 5.81868
R21822 output.n140 output.n110 5.81868
R21823 output.n43 output.n42 5.04292
R21824 output.n74 output.n73 5.04292
R21825 output.n106 output.n105 5.04292
R21826 output.n138 output.n137 5.04292
R21827 output.n28 output.n24 4.38594
R21828 output.n59 output.n55 4.38594
R21829 output.n91 output.n87 4.38594
R21830 output.n123 output.n119 4.38594
R21831 output.n39 output.n17 4.26717
R21832 output.n70 output.n48 4.26717
R21833 output.n102 output.n80 4.26717
R21834 output.n134 output.n112 4.26717
R21835 output.n0 output.t3 3.9605
R21836 output.n0 output.t7 3.9605
R21837 output.n2 output.t11 3.9605
R21838 output.n2 output.t15 3.9605
R21839 output.n4 output.t0 3.9605
R21840 output.n4 output.t5 3.9605
R21841 output.n6 output.t8 3.9605
R21842 output.n6 output.t1 3.9605
R21843 output.n8 output.t4 3.9605
R21844 output.n8 output.t9 3.9605
R21845 output.n10 output.t10 3.9605
R21846 output.n10 output.t12 3.9605
R21847 output.n12 output.t2 3.9605
R21848 output.n12 output.t6 3.9605
R21849 output.n38 output.n19 3.49141
R21850 output.n69 output.n50 3.49141
R21851 output.n101 output.n82 3.49141
R21852 output.n133 output.n114 3.49141
R21853 output.n35 output.n34 2.71565
R21854 output.n66 output.n65 2.71565
R21855 output.n98 output.n97 2.71565
R21856 output.n130 output.n129 2.71565
R21857 output.n31 output.n21 1.93989
R21858 output.n62 output.n52 1.93989
R21859 output.n94 output.n84 1.93989
R21860 output.n126 output.n116 1.93989
R21861 output.n30 output.n23 1.16414
R21862 output.n61 output.n54 1.16414
R21863 output.n93 output.n86 1.16414
R21864 output.n125 output.n118 1.16414
R21865 output.n141 output.n109 0.962709
R21866 output.n109 output.n77 0.962709
R21867 output.n27 output.n26 0.388379
R21868 output.n58 output.n57 0.388379
R21869 output.n90 output.n89 0.388379
R21870 output.n122 output.n121 0.388379
R21871 output.n14 output.n13 0.387128
R21872 output.n13 output.n11 0.387128
R21873 output.n11 output.n9 0.387128
R21874 output.n9 output.n7 0.387128
R21875 output.n7 output.n5 0.387128
R21876 output.n5 output.n3 0.387128
R21877 output.n3 output.n1 0.387128
R21878 output.n44 output.n16 0.155672
R21879 output.n37 output.n16 0.155672
R21880 output.n37 output.n36 0.155672
R21881 output.n36 output.n20 0.155672
R21882 output.n29 output.n20 0.155672
R21883 output.n29 output.n28 0.155672
R21884 output.n75 output.n47 0.155672
R21885 output.n68 output.n47 0.155672
R21886 output.n68 output.n67 0.155672
R21887 output.n67 output.n51 0.155672
R21888 output.n60 output.n51 0.155672
R21889 output.n60 output.n59 0.155672
R21890 output.n107 output.n79 0.155672
R21891 output.n100 output.n79 0.155672
R21892 output.n100 output.n99 0.155672
R21893 output.n99 output.n83 0.155672
R21894 output.n92 output.n83 0.155672
R21895 output.n92 output.n91 0.155672
R21896 output.n139 output.n111 0.155672
R21897 output.n132 output.n111 0.155672
R21898 output.n132 output.n131 0.155672
R21899 output.n131 output.n115 0.155672
R21900 output.n124 output.n115 0.155672
R21901 output.n124 output.n123 0.155672
R21902 output output.n14 0.126227
R21903 minus.n30 minus.t3 243.255
R21904 minus.n29 minus.n27 224.169
R21905 minus.n29 minus.n28 223.454
R21906 minus.n15 minus.t9 199.144
R21907 minus.n2 minus.t11 199.144
R21908 minus.n24 minus.t7 183.883
R21909 minus.n11 minus.t5 183.883
R21910 minus.n18 minus.n17 161.3
R21911 minus.n19 minus.n14 161.3
R21912 minus.n21 minus.n20 161.3
R21913 minus.n23 minus.n13 161.3
R21914 minus.n10 minus.n0 161.3
R21915 minus.n8 minus.n7 161.3
R21916 minus.n6 minus.n1 161.3
R21917 minus.n5 minus.n4 161.3
R21918 minus.n22 minus.t12 144.601
R21919 minus.n16 minus.t8 144.601
R21920 minus.n3 minus.t10 144.601
R21921 minus.n9 minus.t6 144.601
R21922 minus.n25 minus.n24 80.6037
R21923 minus.n12 minus.n11 80.6037
R21924 minus.n24 minus.n23 56.3158
R21925 minus.n11 minus.n10 56.3158
R21926 minus.n16 minus.n15 46.9082
R21927 minus.n3 minus.n2 46.9082
R21928 minus.n5 minus.n2 43.8991
R21929 minus.n18 minus.n15 43.8991
R21930 minus.n21 minus.n14 40.577
R21931 minus.n17 minus.n14 40.577
R21932 minus.n4 minus.n1 40.577
R21933 minus.n8 minus.n1 40.577
R21934 minus.n26 minus.n25 28.1089
R21935 minus.n28 minus.t0 19.8005
R21936 minus.n28 minus.t2 19.8005
R21937 minus.n27 minus.t4 19.8005
R21938 minus.n27 minus.t1 19.8005
R21939 minus.n23 minus.n22 16.477
R21940 minus.n10 minus.n9 16.477
R21941 minus.n26 minus.n12 11.9157
R21942 minus minus.n31 11.5274
R21943 minus.n22 minus.n21 8.11581
R21944 minus.n17 minus.n16 8.11581
R21945 minus.n4 minus.n3 8.11581
R21946 minus.n9 minus.n8 8.11581
R21947 minus.n31 minus.n30 4.80222
R21948 minus.n31 minus.n26 0.972091
R21949 minus.n30 minus.n29 0.716017
R21950 minus.n25 minus.n13 0.285035
R21951 minus.n12 minus.n0 0.285035
R21952 minus.n20 minus.n13 0.189894
R21953 minus.n20 minus.n19 0.189894
R21954 minus.n19 minus.n18 0.189894
R21955 minus.n6 minus.n5 0.189894
R21956 minus.n7 minus.n6 0.189894
R21957 minus.n7 minus.n0 0.189894
R21958 diffpairibias.n27 diffpairibias.n1 289.615
R21959 diffpairibias.n58 diffpairibias.n32 289.615
R21960 diffpairibias.n90 diffpairibias.n64 289.615
R21961 diffpairibias.n122 diffpairibias.n96 289.615
R21962 diffpairibias.n28 diffpairibias.n27 185
R21963 diffpairibias.n26 diffpairibias.n25 185
R21964 diffpairibias.n5 diffpairibias.n4 185
R21965 diffpairibias.n20 diffpairibias.n19 185
R21966 diffpairibias.n18 diffpairibias.n17 185
R21967 diffpairibias.n9 diffpairibias.n8 185
R21968 diffpairibias.n12 diffpairibias.n11 185
R21969 diffpairibias.n59 diffpairibias.n58 185
R21970 diffpairibias.n57 diffpairibias.n56 185
R21971 diffpairibias.n36 diffpairibias.n35 185
R21972 diffpairibias.n51 diffpairibias.n50 185
R21973 diffpairibias.n49 diffpairibias.n48 185
R21974 diffpairibias.n40 diffpairibias.n39 185
R21975 diffpairibias.n43 diffpairibias.n42 185
R21976 diffpairibias.n91 diffpairibias.n90 185
R21977 diffpairibias.n89 diffpairibias.n88 185
R21978 diffpairibias.n68 diffpairibias.n67 185
R21979 diffpairibias.n83 diffpairibias.n82 185
R21980 diffpairibias.n81 diffpairibias.n80 185
R21981 diffpairibias.n72 diffpairibias.n71 185
R21982 diffpairibias.n75 diffpairibias.n74 185
R21983 diffpairibias.n123 diffpairibias.n122 185
R21984 diffpairibias.n121 diffpairibias.n120 185
R21985 diffpairibias.n100 diffpairibias.n99 185
R21986 diffpairibias.n115 diffpairibias.n114 185
R21987 diffpairibias.n113 diffpairibias.n112 185
R21988 diffpairibias.n104 diffpairibias.n103 185
R21989 diffpairibias.n107 diffpairibias.n106 185
R21990 diffpairibias.n0 diffpairibias.t9 178.945
R21991 diffpairibias.n133 diffpairibias.t10 177.018
R21992 diffpairibias.n132 diffpairibias.t11 177.018
R21993 diffpairibias.n0 diffpairibias.t8 177.018
R21994 diffpairibias.t1 diffpairibias.n10 147.661
R21995 diffpairibias.t3 diffpairibias.n41 147.661
R21996 diffpairibias.t5 diffpairibias.n73 147.661
R21997 diffpairibias.t7 diffpairibias.n105 147.661
R21998 diffpairibias.n128 diffpairibias.t0 132.363
R21999 diffpairibias.n128 diffpairibias.t2 130.436
R22000 diffpairibias.n129 diffpairibias.t4 130.436
R22001 diffpairibias.n130 diffpairibias.t6 130.436
R22002 diffpairibias.n27 diffpairibias.n26 104.615
R22003 diffpairibias.n26 diffpairibias.n4 104.615
R22004 diffpairibias.n19 diffpairibias.n4 104.615
R22005 diffpairibias.n19 diffpairibias.n18 104.615
R22006 diffpairibias.n18 diffpairibias.n8 104.615
R22007 diffpairibias.n11 diffpairibias.n8 104.615
R22008 diffpairibias.n58 diffpairibias.n57 104.615
R22009 diffpairibias.n57 diffpairibias.n35 104.615
R22010 diffpairibias.n50 diffpairibias.n35 104.615
R22011 diffpairibias.n50 diffpairibias.n49 104.615
R22012 diffpairibias.n49 diffpairibias.n39 104.615
R22013 diffpairibias.n42 diffpairibias.n39 104.615
R22014 diffpairibias.n90 diffpairibias.n89 104.615
R22015 diffpairibias.n89 diffpairibias.n67 104.615
R22016 diffpairibias.n82 diffpairibias.n67 104.615
R22017 diffpairibias.n82 diffpairibias.n81 104.615
R22018 diffpairibias.n81 diffpairibias.n71 104.615
R22019 diffpairibias.n74 diffpairibias.n71 104.615
R22020 diffpairibias.n122 diffpairibias.n121 104.615
R22021 diffpairibias.n121 diffpairibias.n99 104.615
R22022 diffpairibias.n114 diffpairibias.n99 104.615
R22023 diffpairibias.n114 diffpairibias.n113 104.615
R22024 diffpairibias.n113 diffpairibias.n103 104.615
R22025 diffpairibias.n106 diffpairibias.n103 104.615
R22026 diffpairibias.n63 diffpairibias.n31 95.6354
R22027 diffpairibias.n63 diffpairibias.n62 94.6732
R22028 diffpairibias.n95 diffpairibias.n94 94.6732
R22029 diffpairibias.n127 diffpairibias.n126 94.6732
R22030 diffpairibias.n11 diffpairibias.t1 52.3082
R22031 diffpairibias.n42 diffpairibias.t3 52.3082
R22032 diffpairibias.n74 diffpairibias.t5 52.3082
R22033 diffpairibias.n106 diffpairibias.t7 52.3082
R22034 diffpairibias.n12 diffpairibias.n10 15.6674
R22035 diffpairibias.n43 diffpairibias.n41 15.6674
R22036 diffpairibias.n75 diffpairibias.n73 15.6674
R22037 diffpairibias.n107 diffpairibias.n105 15.6674
R22038 diffpairibias.n13 diffpairibias.n9 12.8005
R22039 diffpairibias.n44 diffpairibias.n40 12.8005
R22040 diffpairibias.n76 diffpairibias.n72 12.8005
R22041 diffpairibias.n108 diffpairibias.n104 12.8005
R22042 diffpairibias.n17 diffpairibias.n16 12.0247
R22043 diffpairibias.n48 diffpairibias.n47 12.0247
R22044 diffpairibias.n80 diffpairibias.n79 12.0247
R22045 diffpairibias.n112 diffpairibias.n111 12.0247
R22046 diffpairibias.n20 diffpairibias.n7 11.249
R22047 diffpairibias.n51 diffpairibias.n38 11.249
R22048 diffpairibias.n83 diffpairibias.n70 11.249
R22049 diffpairibias.n115 diffpairibias.n102 11.249
R22050 diffpairibias.n21 diffpairibias.n5 10.4732
R22051 diffpairibias.n52 diffpairibias.n36 10.4732
R22052 diffpairibias.n84 diffpairibias.n68 10.4732
R22053 diffpairibias.n116 diffpairibias.n100 10.4732
R22054 diffpairibias.n25 diffpairibias.n24 9.69747
R22055 diffpairibias.n56 diffpairibias.n55 9.69747
R22056 diffpairibias.n88 diffpairibias.n87 9.69747
R22057 diffpairibias.n120 diffpairibias.n119 9.69747
R22058 diffpairibias.n31 diffpairibias.n30 9.45567
R22059 diffpairibias.n62 diffpairibias.n61 9.45567
R22060 diffpairibias.n94 diffpairibias.n93 9.45567
R22061 diffpairibias.n126 diffpairibias.n125 9.45567
R22062 diffpairibias.n30 diffpairibias.n29 9.3005
R22063 diffpairibias.n3 diffpairibias.n2 9.3005
R22064 diffpairibias.n24 diffpairibias.n23 9.3005
R22065 diffpairibias.n22 diffpairibias.n21 9.3005
R22066 diffpairibias.n7 diffpairibias.n6 9.3005
R22067 diffpairibias.n16 diffpairibias.n15 9.3005
R22068 diffpairibias.n14 diffpairibias.n13 9.3005
R22069 diffpairibias.n61 diffpairibias.n60 9.3005
R22070 diffpairibias.n34 diffpairibias.n33 9.3005
R22071 diffpairibias.n55 diffpairibias.n54 9.3005
R22072 diffpairibias.n53 diffpairibias.n52 9.3005
R22073 diffpairibias.n38 diffpairibias.n37 9.3005
R22074 diffpairibias.n47 diffpairibias.n46 9.3005
R22075 diffpairibias.n45 diffpairibias.n44 9.3005
R22076 diffpairibias.n93 diffpairibias.n92 9.3005
R22077 diffpairibias.n66 diffpairibias.n65 9.3005
R22078 diffpairibias.n87 diffpairibias.n86 9.3005
R22079 diffpairibias.n85 diffpairibias.n84 9.3005
R22080 diffpairibias.n70 diffpairibias.n69 9.3005
R22081 diffpairibias.n79 diffpairibias.n78 9.3005
R22082 diffpairibias.n77 diffpairibias.n76 9.3005
R22083 diffpairibias.n125 diffpairibias.n124 9.3005
R22084 diffpairibias.n98 diffpairibias.n97 9.3005
R22085 diffpairibias.n119 diffpairibias.n118 9.3005
R22086 diffpairibias.n117 diffpairibias.n116 9.3005
R22087 diffpairibias.n102 diffpairibias.n101 9.3005
R22088 diffpairibias.n111 diffpairibias.n110 9.3005
R22089 diffpairibias.n109 diffpairibias.n108 9.3005
R22090 diffpairibias.n28 diffpairibias.n3 8.92171
R22091 diffpairibias.n59 diffpairibias.n34 8.92171
R22092 diffpairibias.n91 diffpairibias.n66 8.92171
R22093 diffpairibias.n123 diffpairibias.n98 8.92171
R22094 diffpairibias.n29 diffpairibias.n1 8.14595
R22095 diffpairibias.n60 diffpairibias.n32 8.14595
R22096 diffpairibias.n92 diffpairibias.n64 8.14595
R22097 diffpairibias.n124 diffpairibias.n96 8.14595
R22098 diffpairibias.n31 diffpairibias.n1 5.81868
R22099 diffpairibias.n62 diffpairibias.n32 5.81868
R22100 diffpairibias.n94 diffpairibias.n64 5.81868
R22101 diffpairibias.n126 diffpairibias.n96 5.81868
R22102 diffpairibias.n131 diffpairibias.n130 5.20947
R22103 diffpairibias.n29 diffpairibias.n28 5.04292
R22104 diffpairibias.n60 diffpairibias.n59 5.04292
R22105 diffpairibias.n92 diffpairibias.n91 5.04292
R22106 diffpairibias.n124 diffpairibias.n123 5.04292
R22107 diffpairibias.n131 diffpairibias.n127 4.42209
R22108 diffpairibias.n14 diffpairibias.n10 4.38594
R22109 diffpairibias.n45 diffpairibias.n41 4.38594
R22110 diffpairibias.n77 diffpairibias.n73 4.38594
R22111 diffpairibias.n109 diffpairibias.n105 4.38594
R22112 diffpairibias.n132 diffpairibias.n131 4.28454
R22113 diffpairibias.n25 diffpairibias.n3 4.26717
R22114 diffpairibias.n56 diffpairibias.n34 4.26717
R22115 diffpairibias.n88 diffpairibias.n66 4.26717
R22116 diffpairibias.n120 diffpairibias.n98 4.26717
R22117 diffpairibias.n24 diffpairibias.n5 3.49141
R22118 diffpairibias.n55 diffpairibias.n36 3.49141
R22119 diffpairibias.n87 diffpairibias.n68 3.49141
R22120 diffpairibias.n119 diffpairibias.n100 3.49141
R22121 diffpairibias.n21 diffpairibias.n20 2.71565
R22122 diffpairibias.n52 diffpairibias.n51 2.71565
R22123 diffpairibias.n84 diffpairibias.n83 2.71565
R22124 diffpairibias.n116 diffpairibias.n115 2.71565
R22125 diffpairibias.n17 diffpairibias.n7 1.93989
R22126 diffpairibias.n48 diffpairibias.n38 1.93989
R22127 diffpairibias.n80 diffpairibias.n70 1.93989
R22128 diffpairibias.n112 diffpairibias.n102 1.93989
R22129 diffpairibias.n130 diffpairibias.n129 1.9266
R22130 diffpairibias.n129 diffpairibias.n128 1.9266
R22131 diffpairibias.n133 diffpairibias.n132 1.92658
R22132 diffpairibias.n134 diffpairibias.n133 1.29913
R22133 diffpairibias.n16 diffpairibias.n9 1.16414
R22134 diffpairibias.n47 diffpairibias.n40 1.16414
R22135 diffpairibias.n79 diffpairibias.n72 1.16414
R22136 diffpairibias.n111 diffpairibias.n104 1.16414
R22137 diffpairibias.n127 diffpairibias.n95 0.962709
R22138 diffpairibias.n95 diffpairibias.n63 0.962709
R22139 diffpairibias diffpairibias.n134 0.684875
R22140 diffpairibias.n13 diffpairibias.n12 0.388379
R22141 diffpairibias.n44 diffpairibias.n43 0.388379
R22142 diffpairibias.n76 diffpairibias.n75 0.388379
R22143 diffpairibias.n108 diffpairibias.n107 0.388379
R22144 diffpairibias.n134 diffpairibias.n0 0.337251
R22145 diffpairibias.n30 diffpairibias.n2 0.155672
R22146 diffpairibias.n23 diffpairibias.n2 0.155672
R22147 diffpairibias.n23 diffpairibias.n22 0.155672
R22148 diffpairibias.n22 diffpairibias.n6 0.155672
R22149 diffpairibias.n15 diffpairibias.n6 0.155672
R22150 diffpairibias.n15 diffpairibias.n14 0.155672
R22151 diffpairibias.n61 diffpairibias.n33 0.155672
R22152 diffpairibias.n54 diffpairibias.n33 0.155672
R22153 diffpairibias.n54 diffpairibias.n53 0.155672
R22154 diffpairibias.n53 diffpairibias.n37 0.155672
R22155 diffpairibias.n46 diffpairibias.n37 0.155672
R22156 diffpairibias.n46 diffpairibias.n45 0.155672
R22157 diffpairibias.n93 diffpairibias.n65 0.155672
R22158 diffpairibias.n86 diffpairibias.n65 0.155672
R22159 diffpairibias.n86 diffpairibias.n85 0.155672
R22160 diffpairibias.n85 diffpairibias.n69 0.155672
R22161 diffpairibias.n78 diffpairibias.n69 0.155672
R22162 diffpairibias.n78 diffpairibias.n77 0.155672
R22163 diffpairibias.n125 diffpairibias.n97 0.155672
R22164 diffpairibias.n118 diffpairibias.n97 0.155672
R22165 diffpairibias.n118 diffpairibias.n117 0.155672
R22166 diffpairibias.n117 diffpairibias.n101 0.155672
R22167 diffpairibias.n110 diffpairibias.n101 0.155672
R22168 diffpairibias.n110 diffpairibias.n109 0.155672
R22169 outputibias.n27 outputibias.n1 289.615
R22170 outputibias.n58 outputibias.n32 289.615
R22171 outputibias.n90 outputibias.n64 289.615
R22172 outputibias.n122 outputibias.n96 289.615
R22173 outputibias.n28 outputibias.n27 185
R22174 outputibias.n26 outputibias.n25 185
R22175 outputibias.n5 outputibias.n4 185
R22176 outputibias.n20 outputibias.n19 185
R22177 outputibias.n18 outputibias.n17 185
R22178 outputibias.n9 outputibias.n8 185
R22179 outputibias.n12 outputibias.n11 185
R22180 outputibias.n59 outputibias.n58 185
R22181 outputibias.n57 outputibias.n56 185
R22182 outputibias.n36 outputibias.n35 185
R22183 outputibias.n51 outputibias.n50 185
R22184 outputibias.n49 outputibias.n48 185
R22185 outputibias.n40 outputibias.n39 185
R22186 outputibias.n43 outputibias.n42 185
R22187 outputibias.n91 outputibias.n90 185
R22188 outputibias.n89 outputibias.n88 185
R22189 outputibias.n68 outputibias.n67 185
R22190 outputibias.n83 outputibias.n82 185
R22191 outputibias.n81 outputibias.n80 185
R22192 outputibias.n72 outputibias.n71 185
R22193 outputibias.n75 outputibias.n74 185
R22194 outputibias.n123 outputibias.n122 185
R22195 outputibias.n121 outputibias.n120 185
R22196 outputibias.n100 outputibias.n99 185
R22197 outputibias.n115 outputibias.n114 185
R22198 outputibias.n113 outputibias.n112 185
R22199 outputibias.n104 outputibias.n103 185
R22200 outputibias.n107 outputibias.n106 185
R22201 outputibias.n0 outputibias.t8 178.945
R22202 outputibias.n133 outputibias.t10 177.018
R22203 outputibias.n132 outputibias.t11 177.018
R22204 outputibias.n0 outputibias.t9 177.018
R22205 outputibias.t7 outputibias.n10 147.661
R22206 outputibias.t5 outputibias.n41 147.661
R22207 outputibias.t1 outputibias.n73 147.661
R22208 outputibias.t3 outputibias.n105 147.661
R22209 outputibias.n128 outputibias.t6 132.363
R22210 outputibias.n128 outputibias.t4 130.436
R22211 outputibias.n129 outputibias.t0 130.436
R22212 outputibias.n130 outputibias.t2 130.436
R22213 outputibias.n27 outputibias.n26 104.615
R22214 outputibias.n26 outputibias.n4 104.615
R22215 outputibias.n19 outputibias.n4 104.615
R22216 outputibias.n19 outputibias.n18 104.615
R22217 outputibias.n18 outputibias.n8 104.615
R22218 outputibias.n11 outputibias.n8 104.615
R22219 outputibias.n58 outputibias.n57 104.615
R22220 outputibias.n57 outputibias.n35 104.615
R22221 outputibias.n50 outputibias.n35 104.615
R22222 outputibias.n50 outputibias.n49 104.615
R22223 outputibias.n49 outputibias.n39 104.615
R22224 outputibias.n42 outputibias.n39 104.615
R22225 outputibias.n90 outputibias.n89 104.615
R22226 outputibias.n89 outputibias.n67 104.615
R22227 outputibias.n82 outputibias.n67 104.615
R22228 outputibias.n82 outputibias.n81 104.615
R22229 outputibias.n81 outputibias.n71 104.615
R22230 outputibias.n74 outputibias.n71 104.615
R22231 outputibias.n122 outputibias.n121 104.615
R22232 outputibias.n121 outputibias.n99 104.615
R22233 outputibias.n114 outputibias.n99 104.615
R22234 outputibias.n114 outputibias.n113 104.615
R22235 outputibias.n113 outputibias.n103 104.615
R22236 outputibias.n106 outputibias.n103 104.615
R22237 outputibias.n63 outputibias.n31 95.6354
R22238 outputibias.n63 outputibias.n62 94.6732
R22239 outputibias.n95 outputibias.n94 94.6732
R22240 outputibias.n127 outputibias.n126 94.6732
R22241 outputibias.n11 outputibias.t7 52.3082
R22242 outputibias.n42 outputibias.t5 52.3082
R22243 outputibias.n74 outputibias.t1 52.3082
R22244 outputibias.n106 outputibias.t3 52.3082
R22245 outputibias.n12 outputibias.n10 15.6674
R22246 outputibias.n43 outputibias.n41 15.6674
R22247 outputibias.n75 outputibias.n73 15.6674
R22248 outputibias.n107 outputibias.n105 15.6674
R22249 outputibias.n13 outputibias.n9 12.8005
R22250 outputibias.n44 outputibias.n40 12.8005
R22251 outputibias.n76 outputibias.n72 12.8005
R22252 outputibias.n108 outputibias.n104 12.8005
R22253 outputibias.n17 outputibias.n16 12.0247
R22254 outputibias.n48 outputibias.n47 12.0247
R22255 outputibias.n80 outputibias.n79 12.0247
R22256 outputibias.n112 outputibias.n111 12.0247
R22257 outputibias.n20 outputibias.n7 11.249
R22258 outputibias.n51 outputibias.n38 11.249
R22259 outputibias.n83 outputibias.n70 11.249
R22260 outputibias.n115 outputibias.n102 11.249
R22261 outputibias.n21 outputibias.n5 10.4732
R22262 outputibias.n52 outputibias.n36 10.4732
R22263 outputibias.n84 outputibias.n68 10.4732
R22264 outputibias.n116 outputibias.n100 10.4732
R22265 outputibias.n25 outputibias.n24 9.69747
R22266 outputibias.n56 outputibias.n55 9.69747
R22267 outputibias.n88 outputibias.n87 9.69747
R22268 outputibias.n120 outputibias.n119 9.69747
R22269 outputibias.n31 outputibias.n30 9.45567
R22270 outputibias.n62 outputibias.n61 9.45567
R22271 outputibias.n94 outputibias.n93 9.45567
R22272 outputibias.n126 outputibias.n125 9.45567
R22273 outputibias.n30 outputibias.n29 9.3005
R22274 outputibias.n3 outputibias.n2 9.3005
R22275 outputibias.n24 outputibias.n23 9.3005
R22276 outputibias.n22 outputibias.n21 9.3005
R22277 outputibias.n7 outputibias.n6 9.3005
R22278 outputibias.n16 outputibias.n15 9.3005
R22279 outputibias.n14 outputibias.n13 9.3005
R22280 outputibias.n61 outputibias.n60 9.3005
R22281 outputibias.n34 outputibias.n33 9.3005
R22282 outputibias.n55 outputibias.n54 9.3005
R22283 outputibias.n53 outputibias.n52 9.3005
R22284 outputibias.n38 outputibias.n37 9.3005
R22285 outputibias.n47 outputibias.n46 9.3005
R22286 outputibias.n45 outputibias.n44 9.3005
R22287 outputibias.n93 outputibias.n92 9.3005
R22288 outputibias.n66 outputibias.n65 9.3005
R22289 outputibias.n87 outputibias.n86 9.3005
R22290 outputibias.n85 outputibias.n84 9.3005
R22291 outputibias.n70 outputibias.n69 9.3005
R22292 outputibias.n79 outputibias.n78 9.3005
R22293 outputibias.n77 outputibias.n76 9.3005
R22294 outputibias.n125 outputibias.n124 9.3005
R22295 outputibias.n98 outputibias.n97 9.3005
R22296 outputibias.n119 outputibias.n118 9.3005
R22297 outputibias.n117 outputibias.n116 9.3005
R22298 outputibias.n102 outputibias.n101 9.3005
R22299 outputibias.n111 outputibias.n110 9.3005
R22300 outputibias.n109 outputibias.n108 9.3005
R22301 outputibias.n28 outputibias.n3 8.92171
R22302 outputibias.n59 outputibias.n34 8.92171
R22303 outputibias.n91 outputibias.n66 8.92171
R22304 outputibias.n123 outputibias.n98 8.92171
R22305 outputibias.n29 outputibias.n1 8.14595
R22306 outputibias.n60 outputibias.n32 8.14595
R22307 outputibias.n92 outputibias.n64 8.14595
R22308 outputibias.n124 outputibias.n96 8.14595
R22309 outputibias.n31 outputibias.n1 5.81868
R22310 outputibias.n62 outputibias.n32 5.81868
R22311 outputibias.n94 outputibias.n64 5.81868
R22312 outputibias.n126 outputibias.n96 5.81868
R22313 outputibias.n131 outputibias.n130 5.20947
R22314 outputibias.n29 outputibias.n28 5.04292
R22315 outputibias.n60 outputibias.n59 5.04292
R22316 outputibias.n92 outputibias.n91 5.04292
R22317 outputibias.n124 outputibias.n123 5.04292
R22318 outputibias.n131 outputibias.n127 4.42209
R22319 outputibias.n14 outputibias.n10 4.38594
R22320 outputibias.n45 outputibias.n41 4.38594
R22321 outputibias.n77 outputibias.n73 4.38594
R22322 outputibias.n109 outputibias.n105 4.38594
R22323 outputibias.n132 outputibias.n131 4.28454
R22324 outputibias.n25 outputibias.n3 4.26717
R22325 outputibias.n56 outputibias.n34 4.26717
R22326 outputibias.n88 outputibias.n66 4.26717
R22327 outputibias.n120 outputibias.n98 4.26717
R22328 outputibias.n24 outputibias.n5 3.49141
R22329 outputibias.n55 outputibias.n36 3.49141
R22330 outputibias.n87 outputibias.n68 3.49141
R22331 outputibias.n119 outputibias.n100 3.49141
R22332 outputibias.n21 outputibias.n20 2.71565
R22333 outputibias.n52 outputibias.n51 2.71565
R22334 outputibias.n84 outputibias.n83 2.71565
R22335 outputibias.n116 outputibias.n115 2.71565
R22336 outputibias.n17 outputibias.n7 1.93989
R22337 outputibias.n48 outputibias.n38 1.93989
R22338 outputibias.n80 outputibias.n70 1.93989
R22339 outputibias.n112 outputibias.n102 1.93989
R22340 outputibias.n130 outputibias.n129 1.9266
R22341 outputibias.n129 outputibias.n128 1.9266
R22342 outputibias.n133 outputibias.n132 1.92658
R22343 outputibias.n134 outputibias.n133 1.29913
R22344 outputibias.n16 outputibias.n9 1.16414
R22345 outputibias.n47 outputibias.n40 1.16414
R22346 outputibias.n79 outputibias.n72 1.16414
R22347 outputibias.n111 outputibias.n104 1.16414
R22348 outputibias.n127 outputibias.n95 0.962709
R22349 outputibias.n95 outputibias.n63 0.962709
R22350 outputibias.n13 outputibias.n12 0.388379
R22351 outputibias.n44 outputibias.n43 0.388379
R22352 outputibias.n76 outputibias.n75 0.388379
R22353 outputibias.n108 outputibias.n107 0.388379
R22354 outputibias.n134 outputibias.n0 0.337251
R22355 outputibias outputibias.n134 0.302375
R22356 outputibias.n30 outputibias.n2 0.155672
R22357 outputibias.n23 outputibias.n2 0.155672
R22358 outputibias.n23 outputibias.n22 0.155672
R22359 outputibias.n22 outputibias.n6 0.155672
R22360 outputibias.n15 outputibias.n6 0.155672
R22361 outputibias.n15 outputibias.n14 0.155672
R22362 outputibias.n61 outputibias.n33 0.155672
R22363 outputibias.n54 outputibias.n33 0.155672
R22364 outputibias.n54 outputibias.n53 0.155672
R22365 outputibias.n53 outputibias.n37 0.155672
R22366 outputibias.n46 outputibias.n37 0.155672
R22367 outputibias.n46 outputibias.n45 0.155672
R22368 outputibias.n93 outputibias.n65 0.155672
R22369 outputibias.n86 outputibias.n65 0.155672
R22370 outputibias.n86 outputibias.n85 0.155672
R22371 outputibias.n85 outputibias.n69 0.155672
R22372 outputibias.n78 outputibias.n69 0.155672
R22373 outputibias.n78 outputibias.n77 0.155672
R22374 outputibias.n125 outputibias.n97 0.155672
R22375 outputibias.n118 outputibias.n97 0.155672
R22376 outputibias.n118 outputibias.n117 0.155672
R22377 outputibias.n117 outputibias.n101 0.155672
R22378 outputibias.n110 outputibias.n101 0.155672
R22379 outputibias.n110 outputibias.n109 0.155672
C0 CSoutput output 6.13571f
C1 CSoutput outputibias 0.032386f
C2 vdd CSoutput 61.8363f
C3 commonsourceibias output 0.006808f
C4 minus diffpairibias 2.16e-19
C5 CSoutput minus 2.74686f
C6 vdd plus 0.073825f
C7 plus diffpairibias 2.16e-19
C8 commonsourceibias outputibias 0.003832f
C9 CSoutput plus 0.804612f
C10 vdd commonsourceibias 0.004218f
C11 commonsourceibias diffpairibias 0.008433f
C12 CSoutput commonsourceibias 23.9697f
C13 minus plus 7.84338f
C14 minus commonsourceibias 0.306594f
C15 plus commonsourceibias 0.266289f
C16 output outputibias 2.34152f
C17 vdd output 7.23429f
C18 diffpairibias gnd 32.797302f
C19 outputibias gnd 32.467567f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.111895p
C22 plus gnd 25.75477f
C23 minus gnd 22.45568f
C24 CSoutput gnd 73.111244f
C25 vdd gnd 0.352424p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t5 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t3 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t2 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t4 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t10 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t8 gnd 0.108432f
C174 diffpairibias.t9 gnd 0.109185f
C175 diffpairibias.n0 gnd 0.122922f
C176 diffpairibias.n1 gnd 0.001296f
C177 diffpairibias.n2 gnd 9.22e-19
C178 diffpairibias.n3 gnd 4.95e-19
C179 diffpairibias.n4 gnd 0.001171f
C180 diffpairibias.n5 gnd 5.25e-19
C181 diffpairibias.n6 gnd 9.22e-19
C182 diffpairibias.n7 gnd 4.95e-19
C183 diffpairibias.n8 gnd 0.001171f
C184 diffpairibias.n9 gnd 5.25e-19
C185 diffpairibias.n10 gnd 0.003945f
C186 diffpairibias.t1 gnd 0.001909f
C187 diffpairibias.n11 gnd 8.78e-19
C188 diffpairibias.n12 gnd 6.92e-19
C189 diffpairibias.n13 gnd 4.95e-19
C190 diffpairibias.n14 gnd 0.021937f
C191 diffpairibias.n15 gnd 9.22e-19
C192 diffpairibias.n16 gnd 4.95e-19
C193 diffpairibias.n17 gnd 5.25e-19
C194 diffpairibias.n18 gnd 0.001171f
C195 diffpairibias.n19 gnd 0.001171f
C196 diffpairibias.n20 gnd 5.25e-19
C197 diffpairibias.n21 gnd 4.95e-19
C198 diffpairibias.n22 gnd 9.22e-19
C199 diffpairibias.n23 gnd 9.22e-19
C200 diffpairibias.n24 gnd 4.95e-19
C201 diffpairibias.n25 gnd 5.25e-19
C202 diffpairibias.n26 gnd 0.001171f
C203 diffpairibias.n27 gnd 0.002535f
C204 diffpairibias.n28 gnd 5.25e-19
C205 diffpairibias.n29 gnd 4.95e-19
C206 diffpairibias.n30 gnd 0.002131f
C207 diffpairibias.n31 gnd 0.005461f
C208 diffpairibias.n32 gnd 0.001296f
C209 diffpairibias.n33 gnd 9.22e-19
C210 diffpairibias.n34 gnd 4.95e-19
C211 diffpairibias.n35 gnd 0.001171f
C212 diffpairibias.n36 gnd 5.25e-19
C213 diffpairibias.n37 gnd 9.22e-19
C214 diffpairibias.n38 gnd 4.95e-19
C215 diffpairibias.n39 gnd 0.001171f
C216 diffpairibias.n40 gnd 5.25e-19
C217 diffpairibias.n41 gnd 0.003945f
C218 diffpairibias.t3 gnd 0.001909f
C219 diffpairibias.n42 gnd 8.78e-19
C220 diffpairibias.n43 gnd 6.92e-19
C221 diffpairibias.n44 gnd 4.95e-19
C222 diffpairibias.n45 gnd 0.021937f
C223 diffpairibias.n46 gnd 9.22e-19
C224 diffpairibias.n47 gnd 4.95e-19
C225 diffpairibias.n48 gnd 5.25e-19
C226 diffpairibias.n49 gnd 0.001171f
C227 diffpairibias.n50 gnd 0.001171f
C228 diffpairibias.n51 gnd 5.25e-19
C229 diffpairibias.n52 gnd 4.95e-19
C230 diffpairibias.n53 gnd 9.22e-19
C231 diffpairibias.n54 gnd 9.22e-19
C232 diffpairibias.n55 gnd 4.95e-19
C233 diffpairibias.n56 gnd 5.25e-19
C234 diffpairibias.n57 gnd 0.001171f
C235 diffpairibias.n58 gnd 0.002535f
C236 diffpairibias.n59 gnd 5.25e-19
C237 diffpairibias.n60 gnd 4.95e-19
C238 diffpairibias.n61 gnd 0.002131f
C239 diffpairibias.n62 gnd 0.00491f
C240 diffpairibias.n63 gnd 0.11516f
C241 diffpairibias.n64 gnd 0.001296f
C242 diffpairibias.n65 gnd 9.22e-19
C243 diffpairibias.n66 gnd 4.95e-19
C244 diffpairibias.n67 gnd 0.001171f
C245 diffpairibias.n68 gnd 5.25e-19
C246 diffpairibias.n69 gnd 9.22e-19
C247 diffpairibias.n70 gnd 4.95e-19
C248 diffpairibias.n71 gnd 0.001171f
C249 diffpairibias.n72 gnd 5.25e-19
C250 diffpairibias.n73 gnd 0.003945f
C251 diffpairibias.t5 gnd 0.001909f
C252 diffpairibias.n74 gnd 8.78e-19
C253 diffpairibias.n75 gnd 6.92e-19
C254 diffpairibias.n76 gnd 4.95e-19
C255 diffpairibias.n77 gnd 0.021937f
C256 diffpairibias.n78 gnd 9.22e-19
C257 diffpairibias.n79 gnd 4.95e-19
C258 diffpairibias.n80 gnd 5.25e-19
C259 diffpairibias.n81 gnd 0.001171f
C260 diffpairibias.n82 gnd 0.001171f
C261 diffpairibias.n83 gnd 5.25e-19
C262 diffpairibias.n84 gnd 4.95e-19
C263 diffpairibias.n85 gnd 9.22e-19
C264 diffpairibias.n86 gnd 9.22e-19
C265 diffpairibias.n87 gnd 4.95e-19
C266 diffpairibias.n88 gnd 5.25e-19
C267 diffpairibias.n89 gnd 0.001171f
C268 diffpairibias.n90 gnd 0.002535f
C269 diffpairibias.n91 gnd 5.25e-19
C270 diffpairibias.n92 gnd 4.95e-19
C271 diffpairibias.n93 gnd 0.002131f
C272 diffpairibias.n94 gnd 0.00491f
C273 diffpairibias.n95 gnd 0.06095f
C274 diffpairibias.n96 gnd 0.001296f
C275 diffpairibias.n97 gnd 9.22e-19
C276 diffpairibias.n98 gnd 4.95e-19
C277 diffpairibias.n99 gnd 0.001171f
C278 diffpairibias.n100 gnd 5.25e-19
C279 diffpairibias.n101 gnd 9.22e-19
C280 diffpairibias.n102 gnd 4.95e-19
C281 diffpairibias.n103 gnd 0.001171f
C282 diffpairibias.n104 gnd 5.25e-19
C283 diffpairibias.n105 gnd 0.003945f
C284 diffpairibias.t7 gnd 0.001909f
C285 diffpairibias.n106 gnd 8.78e-19
C286 diffpairibias.n107 gnd 6.92e-19
C287 diffpairibias.n108 gnd 4.95e-19
C288 diffpairibias.n109 gnd 0.021937f
C289 diffpairibias.n110 gnd 9.22e-19
C290 diffpairibias.n111 gnd 4.95e-19
C291 diffpairibias.n112 gnd 5.25e-19
C292 diffpairibias.n113 gnd 0.001171f
C293 diffpairibias.n114 gnd 0.001171f
C294 diffpairibias.n115 gnd 5.25e-19
C295 diffpairibias.n116 gnd 4.95e-19
C296 diffpairibias.n117 gnd 9.22e-19
C297 diffpairibias.n118 gnd 9.22e-19
C298 diffpairibias.n119 gnd 4.95e-19
C299 diffpairibias.n120 gnd 5.25e-19
C300 diffpairibias.n121 gnd 0.001171f
C301 diffpairibias.n122 gnd 0.002535f
C302 diffpairibias.n123 gnd 5.25e-19
C303 diffpairibias.n124 gnd 4.95e-19
C304 diffpairibias.n125 gnd 0.002131f
C305 diffpairibias.n126 gnd 0.00491f
C306 diffpairibias.n127 gnd 0.08013f
C307 diffpairibias.t6 gnd 0.102337f
C308 diffpairibias.t4 gnd 0.102337f
C309 diffpairibias.t2 gnd 0.102337f
C310 diffpairibias.t0 gnd 0.103205f
C311 diffpairibias.n128 gnd 0.127236f
C312 diffpairibias.n129 gnd 0.068439f
C313 diffpairibias.n130 gnd 0.07541f
C314 diffpairibias.n131 gnd 0.155794f
C315 diffpairibias.t11 gnd 0.108432f
C316 diffpairibias.n132 gnd 0.063754f
C317 diffpairibias.t10 gnd 0.108432f
C318 diffpairibias.n133 gnd 0.061519f
C319 diffpairibias.n134 gnd 0.040079f
C320 minus.n0 gnd 0.037196f
C321 minus.t6 gnd 0.442682f
C322 minus.n1 gnd 0.022514f
C323 minus.t11 gnd 0.502376f
C324 minus.n2 gnd 0.221655f
C325 minus.t10 gnd 0.442682f
C326 minus.n3 gnd 0.206565f
C327 minus.n4 gnd 0.038013f
C328 minus.n5 gnd 0.119334f
C329 minus.n6 gnd 0.027876f
C330 minus.n7 gnd 0.027876f
C331 minus.n8 gnd 0.038013f
C332 minus.n9 gnd 0.18176f
C333 minus.n10 gnd 0.038235f
C334 minus.t5 gnd 0.485128f
C335 minus.n11 gnd 0.224883f
C336 minus.n12 gnd 0.333286f
C337 minus.n13 gnd 0.037196f
C338 minus.t7 gnd 0.485128f
C339 minus.t12 gnd 0.442682f
C340 minus.n14 gnd 0.022514f
C341 minus.t9 gnd 0.502376f
C342 minus.n15 gnd 0.221655f
C343 minus.t8 gnd 0.442682f
C344 minus.n16 gnd 0.206565f
C345 minus.n17 gnd 0.038013f
C346 minus.n18 gnd 0.119335f
C347 minus.n19 gnd 0.027876f
C348 minus.n20 gnd 0.027876f
C349 minus.n21 gnd 0.038013f
C350 minus.n22 gnd 0.18176f
C351 minus.n23 gnd 0.038235f
C352 minus.n24 gnd 0.224883f
C353 minus.n25 gnd 0.737722f
C354 minus.n26 gnd 1.10137f
C355 minus.t4 gnd 0.008593f
C356 minus.t1 gnd 0.008593f
C357 minus.n27 gnd 0.028257f
C358 minus.t0 gnd 0.008593f
C359 minus.t2 gnd 0.008593f
C360 minus.n28 gnd 0.027869f
C361 minus.n29 gnd 0.237852f
C362 minus.t3 gnd 0.047829f
C363 minus.n30 gnd 0.129794f
C364 minus.n31 gnd 1.74358f
C365 output.t13 gnd 0.464308f
C366 output.t3 gnd 0.044422f
C367 output.t7 gnd 0.044422f
C368 output.n0 gnd 0.364624f
C369 output.n1 gnd 0.614102f
C370 output.t11 gnd 0.044422f
C371 output.t15 gnd 0.044422f
C372 output.n2 gnd 0.364624f
C373 output.n3 gnd 0.350265f
C374 output.t0 gnd 0.044422f
C375 output.t5 gnd 0.044422f
C376 output.n4 gnd 0.364624f
C377 output.n5 gnd 0.350265f
C378 output.t8 gnd 0.044422f
C379 output.t1 gnd 0.044422f
C380 output.n6 gnd 0.364624f
C381 output.n7 gnd 0.350265f
C382 output.t4 gnd 0.044422f
C383 output.t9 gnd 0.044422f
C384 output.n8 gnd 0.364624f
C385 output.n9 gnd 0.350265f
C386 output.t10 gnd 0.044422f
C387 output.t12 gnd 0.044422f
C388 output.n10 gnd 0.364624f
C389 output.n11 gnd 0.350265f
C390 output.t2 gnd 0.044422f
C391 output.t6 gnd 0.044422f
C392 output.n12 gnd 0.364624f
C393 output.n13 gnd 0.350265f
C394 output.t14 gnd 0.462979f
C395 output.n14 gnd 0.28994f
C396 output.n15 gnd 0.015803f
C397 output.n16 gnd 0.011243f
C398 output.n17 gnd 0.006041f
C399 output.n18 gnd 0.01428f
C400 output.n19 gnd 0.006397f
C401 output.n20 gnd 0.011243f
C402 output.n21 gnd 0.006041f
C403 output.n22 gnd 0.01428f
C404 output.n23 gnd 0.006397f
C405 output.n24 gnd 0.048111f
C406 output.t19 gnd 0.023274f
C407 output.n25 gnd 0.01071f
C408 output.n26 gnd 0.008435f
C409 output.n27 gnd 0.006041f
C410 output.n28 gnd 0.267512f
C411 output.n29 gnd 0.011243f
C412 output.n30 gnd 0.006041f
C413 output.n31 gnd 0.006397f
C414 output.n32 gnd 0.01428f
C415 output.n33 gnd 0.01428f
C416 output.n34 gnd 0.006397f
C417 output.n35 gnd 0.006041f
C418 output.n36 gnd 0.011243f
C419 output.n37 gnd 0.011243f
C420 output.n38 gnd 0.006041f
C421 output.n39 gnd 0.006397f
C422 output.n40 gnd 0.01428f
C423 output.n41 gnd 0.030913f
C424 output.n42 gnd 0.006397f
C425 output.n43 gnd 0.006041f
C426 output.n44 gnd 0.025987f
C427 output.n45 gnd 0.097665f
C428 output.n46 gnd 0.015803f
C429 output.n47 gnd 0.011243f
C430 output.n48 gnd 0.006041f
C431 output.n49 gnd 0.01428f
C432 output.n50 gnd 0.006397f
C433 output.n51 gnd 0.011243f
C434 output.n52 gnd 0.006041f
C435 output.n53 gnd 0.01428f
C436 output.n54 gnd 0.006397f
C437 output.n55 gnd 0.048111f
C438 output.t18 gnd 0.023274f
C439 output.n56 gnd 0.01071f
C440 output.n57 gnd 0.008435f
C441 output.n58 gnd 0.006041f
C442 output.n59 gnd 0.267512f
C443 output.n60 gnd 0.011243f
C444 output.n61 gnd 0.006041f
C445 output.n62 gnd 0.006397f
C446 output.n63 gnd 0.01428f
C447 output.n64 gnd 0.01428f
C448 output.n65 gnd 0.006397f
C449 output.n66 gnd 0.006041f
C450 output.n67 gnd 0.011243f
C451 output.n68 gnd 0.011243f
C452 output.n69 gnd 0.006041f
C453 output.n70 gnd 0.006397f
C454 output.n71 gnd 0.01428f
C455 output.n72 gnd 0.030913f
C456 output.n73 gnd 0.006397f
C457 output.n74 gnd 0.006041f
C458 output.n75 gnd 0.025987f
C459 output.n76 gnd 0.09306f
C460 output.n77 gnd 1.65264f
C461 output.n78 gnd 0.015803f
C462 output.n79 gnd 0.011243f
C463 output.n80 gnd 0.006041f
C464 output.n81 gnd 0.01428f
C465 output.n82 gnd 0.006397f
C466 output.n83 gnd 0.011243f
C467 output.n84 gnd 0.006041f
C468 output.n85 gnd 0.01428f
C469 output.n86 gnd 0.006397f
C470 output.n87 gnd 0.048111f
C471 output.t17 gnd 0.023274f
C472 output.n88 gnd 0.01071f
C473 output.n89 gnd 0.008435f
C474 output.n90 gnd 0.006041f
C475 output.n91 gnd 0.267512f
C476 output.n92 gnd 0.011243f
C477 output.n93 gnd 0.006041f
C478 output.n94 gnd 0.006397f
C479 output.n95 gnd 0.01428f
C480 output.n96 gnd 0.01428f
C481 output.n97 gnd 0.006397f
C482 output.n98 gnd 0.006041f
C483 output.n99 gnd 0.011243f
C484 output.n100 gnd 0.011243f
C485 output.n101 gnd 0.006041f
C486 output.n102 gnd 0.006397f
C487 output.n103 gnd 0.01428f
C488 output.n104 gnd 0.030913f
C489 output.n105 gnd 0.006397f
C490 output.n106 gnd 0.006041f
C491 output.n107 gnd 0.025987f
C492 output.n108 gnd 0.09306f
C493 output.n109 gnd 0.713089f
C494 output.n110 gnd 0.015803f
C495 output.n111 gnd 0.011243f
C496 output.n112 gnd 0.006041f
C497 output.n113 gnd 0.01428f
C498 output.n114 gnd 0.006397f
C499 output.n115 gnd 0.011243f
C500 output.n116 gnd 0.006041f
C501 output.n117 gnd 0.01428f
C502 output.n118 gnd 0.006397f
C503 output.n119 gnd 0.048111f
C504 output.t16 gnd 0.023274f
C505 output.n120 gnd 0.01071f
C506 output.n121 gnd 0.008435f
C507 output.n122 gnd 0.006041f
C508 output.n123 gnd 0.267512f
C509 output.n124 gnd 0.011243f
C510 output.n125 gnd 0.006041f
C511 output.n126 gnd 0.006397f
C512 output.n127 gnd 0.01428f
C513 output.n128 gnd 0.01428f
C514 output.n129 gnd 0.006397f
C515 output.n130 gnd 0.006041f
C516 output.n131 gnd 0.011243f
C517 output.n132 gnd 0.011243f
C518 output.n133 gnd 0.006041f
C519 output.n134 gnd 0.006397f
C520 output.n135 gnd 0.01428f
C521 output.n136 gnd 0.030913f
C522 output.n137 gnd 0.006397f
C523 output.n138 gnd 0.006041f
C524 output.n139 gnd 0.025987f
C525 output.n140 gnd 0.09306f
C526 output.n141 gnd 1.67353f
C527 a_n2686_8022.t0 gnd 0.120343p
C528 a_n2686_8022.t3 gnd 0.060238f
C529 a_n2686_8022.n0 gnd 0.013907f
C530 a_n2686_8022.n1 gnd 0.012705f
C531 a_n2686_8022.n2 gnd 0.006827f
C532 a_n2686_8022.n3 gnd 0.016136f
C533 a_n2686_8022.n4 gnd 0.007229f
C534 a_n2686_8022.n5 gnd 0.012705f
C535 a_n2686_8022.n6 gnd 0.006827f
C536 a_n2686_8022.n7 gnd 0.016136f
C537 a_n2686_8022.n8 gnd 0.007229f
C538 a_n2686_8022.n9 gnd 0.056174f
C539 a_n2686_8022.t7 gnd 0.034625f
C540 a_n2686_8022.n10 gnd 0.012102f
C541 a_n2686_8022.n11 gnd 0.01026f
C542 a_n2686_8022.n12 gnd 0.006827f
C543 a_n2686_8022.n13 gnd 0.291437f
C544 a_n2686_8022.n14 gnd 0.012705f
C545 a_n2686_8022.n15 gnd 0.006827f
C546 a_n2686_8022.n16 gnd 0.007229f
C547 a_n2686_8022.n17 gnd 0.016136f
C548 a_n2686_8022.n18 gnd 0.016136f
C549 a_n2686_8022.n19 gnd 0.007229f
C550 a_n2686_8022.n20 gnd 0.006827f
C551 a_n2686_8022.n21 gnd 0.012705f
C552 a_n2686_8022.n22 gnd 0.012705f
C553 a_n2686_8022.n23 gnd 0.006827f
C554 a_n2686_8022.n24 gnd 0.007229f
C555 a_n2686_8022.n25 gnd 0.016136f
C556 a_n2686_8022.n26 gnd 0.038884f
C557 a_n2686_8022.n27 gnd 0.007229f
C558 a_n2686_8022.n28 gnd 0.006827f
C559 a_n2686_8022.n29 gnd 0.029366f
C560 a_n2686_8022.n30 gnd 0.024277f
C561 a_n2686_8022.t10 gnd 0.060238f
C562 a_n2686_8022.t6 gnd 0.060238f
C563 a_n2686_8022.n31 gnd 0.370839f
C564 a_n2686_8022.n32 gnd 0.527012f
C565 a_n2686_8022.t4 gnd 0.060238f
C566 a_n2686_8022.t5 gnd 0.060238f
C567 a_n2686_8022.n33 gnd 0.370839f
C568 a_n2686_8022.n34 gnd 0.410962f
C569 a_n2686_8022.n35 gnd 0.013907f
C570 a_n2686_8022.n36 gnd 0.012705f
C571 a_n2686_8022.n37 gnd 0.006827f
C572 a_n2686_8022.n38 gnd 0.016136f
C573 a_n2686_8022.n39 gnd 0.007229f
C574 a_n2686_8022.n40 gnd 0.012705f
C575 a_n2686_8022.n41 gnd 0.006827f
C576 a_n2686_8022.n42 gnd 0.016136f
C577 a_n2686_8022.n43 gnd 0.007229f
C578 a_n2686_8022.n44 gnd 0.056174f
C579 a_n2686_8022.t8 gnd 0.034625f
C580 a_n2686_8022.n45 gnd 0.012102f
C581 a_n2686_8022.n46 gnd 0.01026f
C582 a_n2686_8022.n47 gnd 0.006827f
C583 a_n2686_8022.n48 gnd 0.291437f
C584 a_n2686_8022.n49 gnd 0.012705f
C585 a_n2686_8022.n50 gnd 0.006827f
C586 a_n2686_8022.n51 gnd 0.007229f
C587 a_n2686_8022.n52 gnd 0.016136f
C588 a_n2686_8022.n53 gnd 0.016136f
C589 a_n2686_8022.n54 gnd 0.007229f
C590 a_n2686_8022.n55 gnd 0.006827f
C591 a_n2686_8022.n56 gnd 0.012705f
C592 a_n2686_8022.n57 gnd 0.012705f
C593 a_n2686_8022.n58 gnd 0.006827f
C594 a_n2686_8022.n59 gnd 0.007229f
C595 a_n2686_8022.n60 gnd 0.016136f
C596 a_n2686_8022.n61 gnd 0.038884f
C597 a_n2686_8022.n62 gnd 0.007229f
C598 a_n2686_8022.n63 gnd 0.006827f
C599 a_n2686_8022.n64 gnd 0.029366f
C600 a_n2686_8022.n65 gnd 0.022518f
C601 a_n2686_8022.n66 gnd 1.17289f
C602 a_n2686_8022.n67 gnd 0.013907f
C603 a_n2686_8022.n68 gnd 0.012705f
C604 a_n2686_8022.n69 gnd 0.006827f
C605 a_n2686_8022.n70 gnd 0.016136f
C606 a_n2686_8022.n71 gnd 0.007229f
C607 a_n2686_8022.n72 gnd 0.012705f
C608 a_n2686_8022.n73 gnd 0.006827f
C609 a_n2686_8022.n74 gnd 0.016136f
C610 a_n2686_8022.n75 gnd 0.007229f
C611 a_n2686_8022.n76 gnd 0.056174f
C612 a_n2686_8022.t17 gnd 0.034625f
C613 a_n2686_8022.n77 gnd 0.012102f
C614 a_n2686_8022.n78 gnd 0.01026f
C615 a_n2686_8022.n79 gnd 0.006827f
C616 a_n2686_8022.n80 gnd 0.291437f
C617 a_n2686_8022.n81 gnd 0.012705f
C618 a_n2686_8022.n82 gnd 0.006827f
C619 a_n2686_8022.n83 gnd 0.007229f
C620 a_n2686_8022.n84 gnd 0.016136f
C621 a_n2686_8022.n85 gnd 0.016136f
C622 a_n2686_8022.n86 gnd 0.007229f
C623 a_n2686_8022.n87 gnd 0.006827f
C624 a_n2686_8022.n88 gnd 0.012705f
C625 a_n2686_8022.n89 gnd 0.012705f
C626 a_n2686_8022.n90 gnd 0.006827f
C627 a_n2686_8022.n91 gnd 0.007229f
C628 a_n2686_8022.n92 gnd 0.016136f
C629 a_n2686_8022.n93 gnd 0.038884f
C630 a_n2686_8022.n94 gnd 0.007229f
C631 a_n2686_8022.n95 gnd 0.006827f
C632 a_n2686_8022.n96 gnd 0.029366f
C633 a_n2686_8022.n97 gnd 0.024277f
C634 a_n2686_8022.t15 gnd 0.060238f
C635 a_n2686_8022.t13 gnd 0.060238f
C636 a_n2686_8022.n98 gnd 0.370839f
C637 a_n2686_8022.n99 gnd 0.527012f
C638 a_n2686_8022.n100 gnd 0.013907f
C639 a_n2686_8022.n101 gnd 0.012705f
C640 a_n2686_8022.n102 gnd 0.006827f
C641 a_n2686_8022.n103 gnd 0.016136f
C642 a_n2686_8022.n104 gnd 0.007229f
C643 a_n2686_8022.n105 gnd 0.012705f
C644 a_n2686_8022.n106 gnd 0.006827f
C645 a_n2686_8022.n107 gnd 0.016136f
C646 a_n2686_8022.n108 gnd 0.007229f
C647 a_n2686_8022.n109 gnd 0.056174f
C648 a_n2686_8022.t20 gnd 0.034625f
C649 a_n2686_8022.n110 gnd 0.012102f
C650 a_n2686_8022.n111 gnd 0.01026f
C651 a_n2686_8022.n112 gnd 0.006827f
C652 a_n2686_8022.n113 gnd 0.291437f
C653 a_n2686_8022.n114 gnd 0.012705f
C654 a_n2686_8022.n115 gnd 0.006827f
C655 a_n2686_8022.n116 gnd 0.007229f
C656 a_n2686_8022.n117 gnd 0.016136f
C657 a_n2686_8022.n118 gnd 0.016136f
C658 a_n2686_8022.n119 gnd 0.007229f
C659 a_n2686_8022.n120 gnd 0.006827f
C660 a_n2686_8022.n121 gnd 0.012705f
C661 a_n2686_8022.n122 gnd 0.012705f
C662 a_n2686_8022.n123 gnd 0.006827f
C663 a_n2686_8022.n124 gnd 0.007229f
C664 a_n2686_8022.n125 gnd 0.016136f
C665 a_n2686_8022.n126 gnd 0.038884f
C666 a_n2686_8022.n127 gnd 0.007229f
C667 a_n2686_8022.n128 gnd 0.006827f
C668 a_n2686_8022.n129 gnd 0.029366f
C669 a_n2686_8022.n130 gnd 0.022518f
C670 a_n2686_8022.n131 gnd 0.132985f
C671 a_n2686_8022.n132 gnd 0.013907f
C672 a_n2686_8022.n133 gnd 0.012705f
C673 a_n2686_8022.n134 gnd 0.006827f
C674 a_n2686_8022.n135 gnd 0.016136f
C675 a_n2686_8022.n136 gnd 0.007229f
C676 a_n2686_8022.n137 gnd 0.012705f
C677 a_n2686_8022.n138 gnd 0.006827f
C678 a_n2686_8022.n139 gnd 0.016136f
C679 a_n2686_8022.n140 gnd 0.007229f
C680 a_n2686_8022.n141 gnd 0.056174f
C681 a_n2686_8022.t16 gnd 0.034625f
C682 a_n2686_8022.n142 gnd 0.012102f
C683 a_n2686_8022.n143 gnd 0.01026f
C684 a_n2686_8022.n144 gnd 0.006827f
C685 a_n2686_8022.n145 gnd 0.291437f
C686 a_n2686_8022.n146 gnd 0.012705f
C687 a_n2686_8022.n147 gnd 0.006827f
C688 a_n2686_8022.n148 gnd 0.007229f
C689 a_n2686_8022.n149 gnd 0.016136f
C690 a_n2686_8022.n150 gnd 0.016136f
C691 a_n2686_8022.n151 gnd 0.007229f
C692 a_n2686_8022.n152 gnd 0.006827f
C693 a_n2686_8022.n153 gnd 0.012705f
C694 a_n2686_8022.n154 gnd 0.012705f
C695 a_n2686_8022.n155 gnd 0.006827f
C696 a_n2686_8022.n156 gnd 0.007229f
C697 a_n2686_8022.n157 gnd 0.016136f
C698 a_n2686_8022.n158 gnd 0.038884f
C699 a_n2686_8022.n159 gnd 0.007229f
C700 a_n2686_8022.n160 gnd 0.006827f
C701 a_n2686_8022.n161 gnd 0.029366f
C702 a_n2686_8022.n162 gnd 0.022518f
C703 a_n2686_8022.n163 gnd 0.132985f
C704 a_n2686_8022.t14 gnd 0.060238f
C705 a_n2686_8022.t19 gnd 0.060238f
C706 a_n2686_8022.n164 gnd 0.370839f
C707 a_n2686_8022.n165 gnd 0.410962f
C708 a_n2686_8022.n166 gnd 0.013907f
C709 a_n2686_8022.n167 gnd 0.012705f
C710 a_n2686_8022.n168 gnd 0.006827f
C711 a_n2686_8022.n169 gnd 0.016136f
C712 a_n2686_8022.n170 gnd 0.007229f
C713 a_n2686_8022.n171 gnd 0.012705f
C714 a_n2686_8022.n172 gnd 0.006827f
C715 a_n2686_8022.n173 gnd 0.016136f
C716 a_n2686_8022.n174 gnd 0.007229f
C717 a_n2686_8022.n175 gnd 0.056174f
C718 a_n2686_8022.t18 gnd 0.034625f
C719 a_n2686_8022.n176 gnd 0.012102f
C720 a_n2686_8022.n177 gnd 0.01026f
C721 a_n2686_8022.n178 gnd 0.006827f
C722 a_n2686_8022.n179 gnd 0.291437f
C723 a_n2686_8022.n180 gnd 0.012705f
C724 a_n2686_8022.n181 gnd 0.006827f
C725 a_n2686_8022.n182 gnd 0.007229f
C726 a_n2686_8022.n183 gnd 0.016136f
C727 a_n2686_8022.n184 gnd 0.016136f
C728 a_n2686_8022.n185 gnd 0.007229f
C729 a_n2686_8022.n186 gnd 0.006827f
C730 a_n2686_8022.n187 gnd 0.012705f
C731 a_n2686_8022.n188 gnd 0.012705f
C732 a_n2686_8022.n189 gnd 0.006827f
C733 a_n2686_8022.n190 gnd 0.007229f
C734 a_n2686_8022.n191 gnd 0.016136f
C735 a_n2686_8022.n192 gnd 0.038884f
C736 a_n2686_8022.n193 gnd 0.007229f
C737 a_n2686_8022.n194 gnd 0.006827f
C738 a_n2686_8022.n195 gnd 0.029366f
C739 a_n2686_8022.n196 gnd 0.022518f
C740 a_n2686_8022.n197 gnd 0.527622f
C741 a_n2686_8022.n198 gnd 1.52338f
C742 a_n2686_8022.n199 gnd 1.76384f
C743 a_n2686_8022.n200 gnd 0.013907f
C744 a_n2686_8022.n201 gnd 0.012705f
C745 a_n2686_8022.n202 gnd 0.006827f
C746 a_n2686_8022.n203 gnd 0.016136f
C747 a_n2686_8022.n204 gnd 0.007229f
C748 a_n2686_8022.n205 gnd 0.012705f
C749 a_n2686_8022.n206 gnd 0.006827f
C750 a_n2686_8022.n207 gnd 0.016136f
C751 a_n2686_8022.n208 gnd 0.007229f
C752 a_n2686_8022.n209 gnd 0.056174f
C753 a_n2686_8022.t2 gnd 0.034625f
C754 a_n2686_8022.n210 gnd 0.012102f
C755 a_n2686_8022.n211 gnd 0.01026f
C756 a_n2686_8022.n212 gnd 0.006827f
C757 a_n2686_8022.n213 gnd 0.291437f
C758 a_n2686_8022.n214 gnd 0.012705f
C759 a_n2686_8022.n215 gnd 0.006827f
C760 a_n2686_8022.n216 gnd 0.007229f
C761 a_n2686_8022.n217 gnd 0.016136f
C762 a_n2686_8022.n218 gnd 0.016136f
C763 a_n2686_8022.n219 gnd 0.007229f
C764 a_n2686_8022.n220 gnd 0.006827f
C765 a_n2686_8022.n221 gnd 0.012705f
C766 a_n2686_8022.n222 gnd 0.012705f
C767 a_n2686_8022.n223 gnd 0.006827f
C768 a_n2686_8022.n224 gnd 0.007229f
C769 a_n2686_8022.n225 gnd 0.016136f
C770 a_n2686_8022.n226 gnd 0.038884f
C771 a_n2686_8022.n227 gnd 0.007229f
C772 a_n2686_8022.n228 gnd 0.006827f
C773 a_n2686_8022.n229 gnd 0.029366f
C774 a_n2686_8022.n230 gnd 0.022518f
C775 a_n2686_8022.n231 gnd 0.478674f
C776 a_n2686_8022.t1 gnd 0.060238f
C777 a_n2686_8022.t11 gnd 0.060238f
C778 a_n2686_8022.n232 gnd 0.370839f
C779 a_n2686_8022.n233 gnd 0.410962f
C780 a_n2686_8022.n234 gnd 0.013907f
C781 a_n2686_8022.n235 gnd 0.012705f
C782 a_n2686_8022.n236 gnd 0.006827f
C783 a_n2686_8022.n237 gnd 0.016136f
C784 a_n2686_8022.n238 gnd 0.007229f
C785 a_n2686_8022.n239 gnd 0.012705f
C786 a_n2686_8022.n240 gnd 0.006827f
C787 a_n2686_8022.n241 gnd 0.016136f
C788 a_n2686_8022.n242 gnd 0.007229f
C789 a_n2686_8022.n243 gnd 0.056174f
C790 a_n2686_8022.t9 gnd 0.034625f
C791 a_n2686_8022.n244 gnd 0.012102f
C792 a_n2686_8022.n245 gnd 0.01026f
C793 a_n2686_8022.n246 gnd 0.006827f
C794 a_n2686_8022.n247 gnd 0.291437f
C795 a_n2686_8022.n248 gnd 0.012705f
C796 a_n2686_8022.n249 gnd 0.006827f
C797 a_n2686_8022.n250 gnd 0.007229f
C798 a_n2686_8022.n251 gnd 0.016136f
C799 a_n2686_8022.n252 gnd 0.016136f
C800 a_n2686_8022.n253 gnd 0.007229f
C801 a_n2686_8022.n254 gnd 0.006827f
C802 a_n2686_8022.n255 gnd 0.012705f
C803 a_n2686_8022.n256 gnd 0.012705f
C804 a_n2686_8022.n257 gnd 0.006827f
C805 a_n2686_8022.n258 gnd 0.007229f
C806 a_n2686_8022.n259 gnd 0.016136f
C807 a_n2686_8022.n260 gnd 0.038884f
C808 a_n2686_8022.n261 gnd 0.007229f
C809 a_n2686_8022.n262 gnd 0.006827f
C810 a_n2686_8022.n263 gnd 0.029366f
C811 a_n2686_8022.n264 gnd 0.024277f
C812 a_n2686_8022.n265 gnd 0.527012f
C813 a_n2686_8022.n266 gnd 0.370839f
C814 a_n2686_8022.t12 gnd 0.060238f
C815 a_n2511_10156.t8 gnd 0.115035f
C816 a_n2511_10156.t12 gnd 0.115035f
C817 a_n2511_10156.t15 gnd 0.115035f
C818 a_n2511_10156.n0 gnd 0.831205f
C819 a_n2511_10156.t16 gnd 0.115035f
C820 a_n2511_10156.t14 gnd 0.115035f
C821 a_n2511_10156.n1 gnd 0.827337f
C822 a_n2511_10156.n2 gnd 1.45743f
C823 a_n2511_10156.t11 gnd 0.115035f
C824 a_n2511_10156.t10 gnd 0.115035f
C825 a_n2511_10156.n3 gnd 0.830094f
C826 a_n2511_10156.t17 gnd 0.115035f
C827 a_n2511_10156.t19 gnd 0.115035f
C828 a_n2511_10156.n4 gnd 0.827337f
C829 a_n2511_10156.n5 gnd 2.52538f
C830 a_n2511_10156.t9 gnd 0.115035f
C831 a_n2511_10156.t13 gnd 0.115035f
C832 a_n2511_10156.n6 gnd 0.827337f
C833 a_n2511_10156.n7 gnd 3.96056f
C834 a_n2511_10156.n8 gnd 0.026557f
C835 a_n2511_10156.n9 gnd 0.024262f
C836 a_n2511_10156.n10 gnd 0.013037f
C837 a_n2511_10156.n11 gnd 0.030816f
C838 a_n2511_10156.n12 gnd 0.013804f
C839 a_n2511_10156.n13 gnd 0.024262f
C840 a_n2511_10156.n14 gnd 0.013037f
C841 a_n2511_10156.n15 gnd 0.030816f
C842 a_n2511_10156.n16 gnd 0.013804f
C843 a_n2511_10156.n17 gnd 0.107274f
C844 a_n2511_10156.t4 gnd 0.066122f
C845 a_n2511_10156.n18 gnd 0.023112f
C846 a_n2511_10156.n19 gnd 0.019593f
C847 a_n2511_10156.n20 gnd 0.013037f
C848 a_n2511_10156.n21 gnd 0.556554f
C849 a_n2511_10156.n22 gnd 0.024262f
C850 a_n2511_10156.n23 gnd 0.013037f
C851 a_n2511_10156.n24 gnd 0.013804f
C852 a_n2511_10156.n25 gnd 0.030816f
C853 a_n2511_10156.n26 gnd 0.030816f
C854 a_n2511_10156.n27 gnd 0.013804f
C855 a_n2511_10156.n28 gnd 0.013037f
C856 a_n2511_10156.n29 gnd 0.024262f
C857 a_n2511_10156.n30 gnd 0.024262f
C858 a_n2511_10156.n31 gnd 0.013037f
C859 a_n2511_10156.n32 gnd 0.013804f
C860 a_n2511_10156.n33 gnd 0.030816f
C861 a_n2511_10156.n34 gnd 0.074256f
C862 a_n2511_10156.n35 gnd 0.013804f
C863 a_n2511_10156.n36 gnd 0.013037f
C864 a_n2511_10156.n37 gnd 0.056081f
C865 a_n2511_10156.n38 gnd 0.046363f
C866 a_n2511_10156.t1 gnd 0.115035f
C867 a_n2511_10156.t3 gnd 0.115035f
C868 a_n2511_10156.n39 gnd 0.708188f
C869 a_n2511_10156.n40 gnd 1.00643f
C870 a_n2511_10156.n41 gnd 0.026557f
C871 a_n2511_10156.n42 gnd 0.024262f
C872 a_n2511_10156.n43 gnd 0.013037f
C873 a_n2511_10156.n44 gnd 0.030816f
C874 a_n2511_10156.n45 gnd 0.013804f
C875 a_n2511_10156.n46 gnd 0.024262f
C876 a_n2511_10156.n47 gnd 0.013037f
C877 a_n2511_10156.n48 gnd 0.030816f
C878 a_n2511_10156.n49 gnd 0.013804f
C879 a_n2511_10156.n50 gnd 0.107274f
C880 a_n2511_10156.t7 gnd 0.066122f
C881 a_n2511_10156.n51 gnd 0.023112f
C882 a_n2511_10156.n52 gnd 0.019593f
C883 a_n2511_10156.n53 gnd 0.013037f
C884 a_n2511_10156.n54 gnd 0.556554f
C885 a_n2511_10156.n55 gnd 0.024262f
C886 a_n2511_10156.n56 gnd 0.013037f
C887 a_n2511_10156.n57 gnd 0.013804f
C888 a_n2511_10156.n58 gnd 0.030816f
C889 a_n2511_10156.n59 gnd 0.030816f
C890 a_n2511_10156.n60 gnd 0.013804f
C891 a_n2511_10156.n61 gnd 0.013037f
C892 a_n2511_10156.n62 gnd 0.024262f
C893 a_n2511_10156.n63 gnd 0.024262f
C894 a_n2511_10156.n64 gnd 0.013037f
C895 a_n2511_10156.n65 gnd 0.013804f
C896 a_n2511_10156.n66 gnd 0.030816f
C897 a_n2511_10156.n67 gnd 0.074256f
C898 a_n2511_10156.n68 gnd 0.013804f
C899 a_n2511_10156.n69 gnd 0.013037f
C900 a_n2511_10156.n70 gnd 0.056081f
C901 a_n2511_10156.n71 gnd 0.043002f
C902 a_n2511_10156.n72 gnd 0.25396f
C903 a_n2511_10156.n73 gnd 0.026557f
C904 a_n2511_10156.n74 gnd 0.024262f
C905 a_n2511_10156.n75 gnd 0.013037f
C906 a_n2511_10156.n76 gnd 0.030816f
C907 a_n2511_10156.n77 gnd 0.013804f
C908 a_n2511_10156.n78 gnd 0.024262f
C909 a_n2511_10156.n79 gnd 0.013037f
C910 a_n2511_10156.n80 gnd 0.030816f
C911 a_n2511_10156.n81 gnd 0.013804f
C912 a_n2511_10156.n82 gnd 0.107274f
C913 a_n2511_10156.t2 gnd 0.066122f
C914 a_n2511_10156.n83 gnd 0.023112f
C915 a_n2511_10156.n84 gnd 0.019593f
C916 a_n2511_10156.n85 gnd 0.013037f
C917 a_n2511_10156.n86 gnd 0.556554f
C918 a_n2511_10156.n87 gnd 0.024262f
C919 a_n2511_10156.n88 gnd 0.013037f
C920 a_n2511_10156.n89 gnd 0.013804f
C921 a_n2511_10156.n90 gnd 0.030816f
C922 a_n2511_10156.n91 gnd 0.030816f
C923 a_n2511_10156.n92 gnd 0.013804f
C924 a_n2511_10156.n93 gnd 0.013037f
C925 a_n2511_10156.n94 gnd 0.024262f
C926 a_n2511_10156.n95 gnd 0.024262f
C927 a_n2511_10156.n96 gnd 0.013037f
C928 a_n2511_10156.n97 gnd 0.013804f
C929 a_n2511_10156.n98 gnd 0.030816f
C930 a_n2511_10156.n99 gnd 0.074256f
C931 a_n2511_10156.n100 gnd 0.013804f
C932 a_n2511_10156.n101 gnd 0.013037f
C933 a_n2511_10156.n102 gnd 0.056081f
C934 a_n2511_10156.n103 gnd 0.043002f
C935 a_n2511_10156.n104 gnd 0.25396f
C936 a_n2511_10156.t6 gnd 0.115035f
C937 a_n2511_10156.t0 gnd 0.115035f
C938 a_n2511_10156.n105 gnd 0.708188f
C939 a_n2511_10156.n106 gnd 0.78481f
C940 a_n2511_10156.n107 gnd 0.026557f
C941 a_n2511_10156.n108 gnd 0.024262f
C942 a_n2511_10156.n109 gnd 0.013037f
C943 a_n2511_10156.n110 gnd 0.030816f
C944 a_n2511_10156.n111 gnd 0.013804f
C945 a_n2511_10156.n112 gnd 0.024262f
C946 a_n2511_10156.n113 gnd 0.013037f
C947 a_n2511_10156.n114 gnd 0.030816f
C948 a_n2511_10156.n115 gnd 0.013804f
C949 a_n2511_10156.n116 gnd 0.107274f
C950 a_n2511_10156.t5 gnd 0.066122f
C951 a_n2511_10156.n117 gnd 0.023112f
C952 a_n2511_10156.n118 gnd 0.019593f
C953 a_n2511_10156.n119 gnd 0.013037f
C954 a_n2511_10156.n120 gnd 0.556554f
C955 a_n2511_10156.n121 gnd 0.024262f
C956 a_n2511_10156.n122 gnd 0.013037f
C957 a_n2511_10156.n123 gnd 0.013804f
C958 a_n2511_10156.n124 gnd 0.030816f
C959 a_n2511_10156.n125 gnd 0.030816f
C960 a_n2511_10156.n126 gnd 0.013804f
C961 a_n2511_10156.n127 gnd 0.013037f
C962 a_n2511_10156.n128 gnd 0.024262f
C963 a_n2511_10156.n129 gnd 0.024262f
C964 a_n2511_10156.n130 gnd 0.013037f
C965 a_n2511_10156.n131 gnd 0.013804f
C966 a_n2511_10156.n132 gnd 0.030816f
C967 a_n2511_10156.n133 gnd 0.074256f
C968 a_n2511_10156.n134 gnd 0.013804f
C969 a_n2511_10156.n135 gnd 0.013037f
C970 a_n2511_10156.n136 gnd 0.056081f
C971 a_n2511_10156.n137 gnd 0.043002f
C972 a_n2511_10156.n138 gnd 1.00759f
C973 a_n2511_10156.n139 gnd 2.19047f
C974 a_n2511_10156.n140 gnd 1.64036f
C975 a_n2511_10156.n141 gnd 0.827337f
C976 a_n2511_10156.t18 gnd 0.115035f
C977 a_n2686_12378.n0 gnd 0.76127f
C978 a_n2686_12378.n1 gnd 0.353754f
C979 a_n2686_12378.n2 gnd 0.758272f
C980 a_n2686_12378.n3 gnd 0.622246f
C981 a_n2686_12378.n4 gnd 0.353754f
C982 a_n2686_12378.n5 gnd 0.680802f
C983 a_n2686_12378.n6 gnd 0.353754f
C984 a_n2686_12378.n7 gnd 0.725401f
C985 a_n2686_12378.n8 gnd 0.353754f
C986 a_n2686_12378.n9 gnd 0.634611f
C987 a_n2686_12378.n10 gnd 0.353754f
C988 a_n2686_12378.n11 gnd 0.553928f
C989 a_n2686_12378.n12 gnd 0.353754f
C990 a_n2686_12378.n13 gnd 0.054189f
C991 a_n2686_12378.n14 gnd 0.054189f
C992 a_n2686_12378.n15 gnd 0.054189f
C993 a_n2686_12378.n16 gnd 0.04539f
C994 a_n2686_12378.n17 gnd 0.054189f
C995 a_n2686_12378.n18 gnd 0.04539f
C996 a_n2686_12378.n19 gnd 0.054189f
C997 a_n2686_12378.n20 gnd 0.04539f
C998 a_n2686_12378.n21 gnd 0.054189f
C999 a_n2686_12378.n22 gnd 0.074463f
C1000 a_n2686_12378.n23 gnd 0.04539f
C1001 a_n2686_12378.n24 gnd 0.061636f
C1002 a_n2686_12378.n25 gnd 0.092382f
C1003 a_n2686_12378.n26 gnd 0.107827f
C1004 a_n2686_12378.n27 gnd 0.074463f
C1005 a_n2686_12378.n28 gnd 0.04539f
C1006 a_n2686_12378.n29 gnd 0.061636f
C1007 a_n2686_12378.n30 gnd 0.092382f
C1008 a_n2686_12378.n31 gnd 0.107827f
C1009 a_n2686_12378.n32 gnd 0.074463f
C1010 a_n2686_12378.n33 gnd 0.04539f
C1011 a_n2686_12378.n34 gnd 0.061636f
C1012 a_n2686_12378.n35 gnd 0.092382f
C1013 a_n2686_12378.n36 gnd 0.107827f
C1014 a_n2686_12378.n37 gnd 0.074463f
C1015 a_n2686_12378.n38 gnd 0.04539f
C1016 a_n2686_12378.n39 gnd 0.061636f
C1017 a_n2686_12378.n40 gnd 0.092382f
C1018 a_n2686_12378.n41 gnd 0.107827f
C1019 a_n2686_12378.n42 gnd 0.092382f
C1020 a_n2686_12378.n43 gnd 0.061636f
C1021 a_n2686_12378.n44 gnd 0.092382f
C1022 a_n2686_12378.n45 gnd 0.092382f
C1023 a_n2686_12378.n46 gnd 0.092382f
C1024 a_n2686_12378.n47 gnd 0.04539f
C1025 a_n2686_12378.n48 gnd 0.107827f
C1026 a_n2686_12378.n49 gnd 0.054189f
C1027 a_n2686_12378.n50 gnd 0.123504f
C1028 a_n2686_12378.n51 gnd 0.042097f
C1029 a_n2686_12378.n52 gnd 0.036039f
C1030 a_n2686_12378.n53 gnd 0.036039f
C1031 a_n2686_12378.n54 gnd 0.431369f
C1032 a_n2686_12378.n55 gnd 0.036039f
C1033 a_n2686_12378.n56 gnd 0.036039f
C1034 a_n2686_12378.n57 gnd 0.431369f
C1035 a_n2686_12378.n58 gnd 0.036039f
C1036 a_n2686_12378.n59 gnd 0.036039f
C1037 a_n2686_12378.n60 gnd 0.431369f
C1038 a_n2686_12378.n61 gnd 0.036039f
C1039 a_n2686_12378.n62 gnd 0.036039f
C1040 a_n2686_12378.n63 gnd 0.431369f
C1041 a_n2686_12378.t30 gnd 0.085436f
C1042 a_n2686_12378.t40 gnd 0.84474f
C1043 a_n2686_12378.t49 gnd 0.733544f
C1044 a_n2686_12378.n64 gnd 0.399646f
C1045 a_n2686_12378.t46 gnd 0.733544f
C1046 a_n2686_12378.t37 gnd 0.733544f
C1047 a_n2686_12378.t44 gnd 0.733544f
C1048 a_n2686_12378.n65 gnd 0.399646f
C1049 a_n2686_12378.t41 gnd 0.84474f
C1050 a_n2686_12378.n66 gnd 0.019724f
C1051 a_n2686_12378.n67 gnd 0.009683f
C1052 a_n2686_12378.n68 gnd 0.022887f
C1053 a_n2686_12378.n69 gnd 0.010252f
C1054 a_n2686_12378.n70 gnd 0.009683f
C1055 a_n2686_12378.n71 gnd 0.022887f
C1056 a_n2686_12378.n72 gnd 0.010252f
C1057 a_n2686_12378.n73 gnd 0.079672f
C1058 a_n2686_12378.t16 gnd 0.049109f
C1059 a_n2686_12378.n74 gnd 0.017165f
C1060 a_n2686_12378.n75 gnd 0.014552f
C1061 a_n2686_12378.n76 gnd 0.009683f
C1062 a_n2686_12378.n77 gnd 0.009683f
C1063 a_n2686_12378.n78 gnd 0.010252f
C1064 a_n2686_12378.n79 gnd 0.022887f
C1065 a_n2686_12378.n80 gnd 0.022887f
C1066 a_n2686_12378.n81 gnd 0.010252f
C1067 a_n2686_12378.n82 gnd 0.009683f
C1068 a_n2686_12378.n83 gnd 0.009683f
C1069 a_n2686_12378.n84 gnd 0.010252f
C1070 a_n2686_12378.n85 gnd 0.022887f
C1071 a_n2686_12378.n86 gnd 0.055149f
C1072 a_n2686_12378.n87 gnd 0.010252f
C1073 a_n2686_12378.n88 gnd 0.009683f
C1074 a_n2686_12378.n89 gnd 0.041651f
C1075 a_n2686_12378.n90 gnd 0.034433f
C1076 a_n2686_12378.t8 gnd 0.085436f
C1077 a_n2686_12378.t10 gnd 0.085436f
C1078 a_n2686_12378.n91 gnd 0.525968f
C1079 a_n2686_12378.n92 gnd 0.747471f
C1080 a_n2686_12378.t22 gnd 0.085436f
C1081 a_n2686_12378.t18 gnd 0.085436f
C1082 a_n2686_12378.n93 gnd 0.525968f
C1083 a_n2686_12378.n94 gnd 0.582875f
C1084 a_n2686_12378.n95 gnd 0.019724f
C1085 a_n2686_12378.n96 gnd 0.009683f
C1086 a_n2686_12378.n97 gnd 0.022887f
C1087 a_n2686_12378.n98 gnd 0.010252f
C1088 a_n2686_12378.n99 gnd 0.009683f
C1089 a_n2686_12378.n100 gnd 0.022887f
C1090 a_n2686_12378.n101 gnd 0.010252f
C1091 a_n2686_12378.n102 gnd 0.079672f
C1092 a_n2686_12378.t6 gnd 0.049109f
C1093 a_n2686_12378.n103 gnd 0.017165f
C1094 a_n2686_12378.n104 gnd 0.014552f
C1095 a_n2686_12378.n105 gnd 0.009683f
C1096 a_n2686_12378.n106 gnd 0.009683f
C1097 a_n2686_12378.n107 gnd 0.010252f
C1098 a_n2686_12378.n108 gnd 0.022887f
C1099 a_n2686_12378.n109 gnd 0.022887f
C1100 a_n2686_12378.n110 gnd 0.010252f
C1101 a_n2686_12378.n111 gnd 0.009683f
C1102 a_n2686_12378.n112 gnd 0.009683f
C1103 a_n2686_12378.n113 gnd 0.010252f
C1104 a_n2686_12378.n114 gnd 0.022887f
C1105 a_n2686_12378.n115 gnd 0.055149f
C1106 a_n2686_12378.n116 gnd 0.010252f
C1107 a_n2686_12378.n117 gnd 0.009683f
C1108 a_n2686_12378.n118 gnd 0.041651f
C1109 a_n2686_12378.n119 gnd 0.031937f
C1110 a_n2686_12378.n120 gnd 0.69539f
C1111 a_n2686_12378.t59 gnd 0.733544f
C1112 a_n2686_12378.t42 gnd 0.733544f
C1113 a_n2686_12378.t56 gnd 0.803878f
C1114 a_n2686_12378.t55 gnd 0.733544f
C1115 a_n2686_12378.t58 gnd 0.733544f
C1116 a_n2686_12378.t48 gnd 0.803878f
C1117 a_n2686_12378.t54 gnd 0.733544f
C1118 a_n2686_12378.t50 gnd 0.733544f
C1119 a_n2686_12378.t33 gnd 0.803878f
C1120 a_n2686_12378.t34 gnd 0.733544f
C1121 a_n2686_12378.t53 gnd 0.733544f
C1122 a_n2686_12378.t36 gnd 0.803878f
C1123 a_n2686_12378.t52 gnd 0.84474f
C1124 a_n2686_12378.t57 gnd 0.733544f
C1125 a_n2686_12378.n121 gnd 0.399646f
C1126 a_n2686_12378.t35 gnd 0.733544f
C1127 a_n2686_12378.t51 gnd 0.733544f
C1128 a_n2686_12378.t32 gnd 0.733544f
C1129 a_n2686_12378.n122 gnd 0.399646f
C1130 a_n2686_12378.t38 gnd 0.84474f
C1131 a_n2686_12378.t15 gnd 0.84474f
C1132 a_n2686_12378.t7 gnd 0.733544f
C1133 a_n2686_12378.n123 gnd 0.399646f
C1134 a_n2686_12378.t9 gnd 0.733544f
C1135 a_n2686_12378.t21 gnd 0.733544f
C1136 a_n2686_12378.t17 gnd 0.733544f
C1137 a_n2686_12378.n124 gnd 0.399646f
C1138 a_n2686_12378.t5 gnd 0.84474f
C1139 a_n2686_12378.n125 gnd 0.382257f
C1140 a_n2686_12378.n126 gnd 0.074463f
C1141 a_n2686_12378.n127 gnd 0.338826f
C1142 a_n2686_12378.n128 gnd 0.382257f
C1143 a_n2686_12378.n129 gnd 0.074463f
C1144 a_n2686_12378.n130 gnd 0.338826f
C1145 a_n2686_12378.t19 gnd 0.803878f
C1146 a_n2686_12378.t13 gnd 0.733544f
C1147 a_n2686_12378.n131 gnd 0.301185f
C1148 a_n2686_12378.t23 gnd 0.733544f
C1149 a_n2686_12378.t25 gnd 0.733544f
C1150 a_n2686_12378.t11 gnd 0.733544f
C1151 a_n2686_12378.n132 gnd 0.37294f
C1152 a_n2686_12378.t3 gnd 0.803878f
C1153 a_n2686_12378.n133 gnd 0.379225f
C1154 a_n2686_12378.n134 gnd 0.382257f
C1155 a_n2686_12378.n135 gnd 0.074463f
C1156 a_n2686_12378.n136 gnd 0.301185f
C1157 a_n2686_12378.n137 gnd 0.063415f
C1158 a_n2686_12378.n138 gnd 0.056499f
C1159 a_n2686_12378.n139 gnd 0.044594f
C1160 a_n2686_12378.n140 gnd 0.051265f
C1161 a_n2686_12378.n141 gnd 0.369134f
C1162 a_n2686_12378.n142 gnd 0.408054f
C1163 a_n2686_12378.n143 gnd 0.019724f
C1164 a_n2686_12378.n144 gnd 0.009683f
C1165 a_n2686_12378.n145 gnd 0.022887f
C1166 a_n2686_12378.n146 gnd 0.010252f
C1167 a_n2686_12378.n147 gnd 0.009683f
C1168 a_n2686_12378.n148 gnd 0.022887f
C1169 a_n2686_12378.n149 gnd 0.010252f
C1170 a_n2686_12378.n150 gnd 0.079672f
C1171 a_n2686_12378.t4 gnd 0.049109f
C1172 a_n2686_12378.n151 gnd 0.017165f
C1173 a_n2686_12378.n152 gnd 0.014552f
C1174 a_n2686_12378.n153 gnd 0.009683f
C1175 a_n2686_12378.n154 gnd 0.009683f
C1176 a_n2686_12378.n155 gnd 0.010252f
C1177 a_n2686_12378.n156 gnd 0.022887f
C1178 a_n2686_12378.n157 gnd 0.022887f
C1179 a_n2686_12378.n158 gnd 0.010252f
C1180 a_n2686_12378.n159 gnd 0.009683f
C1181 a_n2686_12378.n160 gnd 0.009683f
C1182 a_n2686_12378.n161 gnd 0.010252f
C1183 a_n2686_12378.n162 gnd 0.022887f
C1184 a_n2686_12378.n163 gnd 0.055149f
C1185 a_n2686_12378.n164 gnd 0.010252f
C1186 a_n2686_12378.n165 gnd 0.009683f
C1187 a_n2686_12378.n166 gnd 0.041651f
C1188 a_n2686_12378.n167 gnd 0.034433f
C1189 a_n2686_12378.t26 gnd 0.085436f
C1190 a_n2686_12378.t12 gnd 0.085436f
C1191 a_n2686_12378.n168 gnd 0.525968f
C1192 a_n2686_12378.n169 gnd 0.747471f
C1193 a_n2686_12378.t14 gnd 0.085436f
C1194 a_n2686_12378.t24 gnd 0.085436f
C1195 a_n2686_12378.n170 gnd 0.525968f
C1196 a_n2686_12378.n171 gnd 0.582875f
C1197 a_n2686_12378.n172 gnd 0.019724f
C1198 a_n2686_12378.n173 gnd 0.009683f
C1199 a_n2686_12378.n174 gnd 0.022887f
C1200 a_n2686_12378.n175 gnd 0.010252f
C1201 a_n2686_12378.n176 gnd 0.009683f
C1202 a_n2686_12378.n177 gnd 0.022887f
C1203 a_n2686_12378.n178 gnd 0.010252f
C1204 a_n2686_12378.n179 gnd 0.079672f
C1205 a_n2686_12378.t20 gnd 0.049109f
C1206 a_n2686_12378.n180 gnd 0.017165f
C1207 a_n2686_12378.n181 gnd 0.014552f
C1208 a_n2686_12378.n182 gnd 0.009683f
C1209 a_n2686_12378.n183 gnd 0.009683f
C1210 a_n2686_12378.n184 gnd 0.010252f
C1211 a_n2686_12378.n185 gnd 0.022887f
C1212 a_n2686_12378.n186 gnd 0.022887f
C1213 a_n2686_12378.n187 gnd 0.010252f
C1214 a_n2686_12378.n188 gnd 0.009683f
C1215 a_n2686_12378.n189 gnd 0.009683f
C1216 a_n2686_12378.n190 gnd 0.010252f
C1217 a_n2686_12378.n191 gnd 0.022887f
C1218 a_n2686_12378.n192 gnd 0.055149f
C1219 a_n2686_12378.n193 gnd 0.010252f
C1220 a_n2686_12378.n194 gnd 0.009683f
C1221 a_n2686_12378.n195 gnd 0.041651f
C1222 a_n2686_12378.n196 gnd 0.031937f
C1223 a_n2686_12378.n197 gnd 0.606936f
C1224 a_n2686_12378.n198 gnd 0.542054f
C1225 a_n2686_12378.n199 gnd 0.724548f
C1226 a_n2686_12378.n200 gnd 0.371593f
C1227 a_n2686_12378.n201 gnd 0.372641f
C1228 a_n2686_12378.n202 gnd 0.063358f
C1229 a_n2686_12378.n203 gnd 0.344616f
C1230 a_n2686_12378.n204 gnd 0.301185f
C1231 a_n2686_12378.n205 gnd 0.063358f
C1232 a_n2686_12378.t45 gnd 0.803878f
C1233 a_n2686_12378.n206 gnd 0.372641f
C1234 a_n2686_12378.n207 gnd 0.120794f
C1235 a_n2686_12378.n208 gnd 0.120794f
C1236 a_n2686_12378.n209 gnd 0.372641f
C1237 a_n2686_12378.n210 gnd 0.063358f
C1238 a_n2686_12378.n211 gnd 0.344616f
C1239 a_n2686_12378.n212 gnd 0.301185f
C1240 a_n2686_12378.n213 gnd 0.063358f
C1241 a_n2686_12378.t43 gnd 0.803878f
C1242 a_n2686_12378.n214 gnd 0.372641f
C1243 a_n2686_12378.n215 gnd 0.155538f
C1244 a_n2686_12378.n216 gnd 0.155538f
C1245 a_n2686_12378.n217 gnd 0.372641f
C1246 a_n2686_12378.n218 gnd 0.063358f
C1247 a_n2686_12378.n219 gnd 0.344616f
C1248 a_n2686_12378.n220 gnd 0.301185f
C1249 a_n2686_12378.n221 gnd 0.063358f
C1250 a_n2686_12378.t39 gnd 0.803878f
C1251 a_n2686_12378.n222 gnd 0.372641f
C1252 a_n2686_12378.n223 gnd 0.120794f
C1253 a_n2686_12378.n224 gnd 0.120794f
C1254 a_n2686_12378.n225 gnd 0.372641f
C1255 a_n2686_12378.n226 gnd 0.063358f
C1256 a_n2686_12378.n227 gnd 0.344616f
C1257 a_n2686_12378.n228 gnd 0.301185f
C1258 a_n2686_12378.n229 gnd 0.063358f
C1259 a_n2686_12378.t47 gnd 0.803878f
C1260 a_n2686_12378.n230 gnd 0.372641f
C1261 a_n2686_12378.n231 gnd 0.371593f
C1262 a_n2686_12378.n232 gnd 0.922404f
C1263 a_n2686_12378.n233 gnd 0.382257f
C1264 a_n2686_12378.n234 gnd 0.074463f
C1265 a_n2686_12378.n235 gnd 0.338826f
C1266 a_n2686_12378.n236 gnd 2.62959f
C1267 a_n2686_12378.t1 gnd 0.085436f
C1268 a_n2686_12378.t27 gnd 0.085436f
C1269 a_n2686_12378.n237 gnd 0.747348f
C1270 a_n2686_12378.n238 gnd 2.77836f
C1271 a_n2686_12378.t28 gnd 0.085436f
C1272 a_n2686_12378.t29 gnd 0.085436f
C1273 a_n2686_12378.n239 gnd 0.746153f
C1274 a_n2686_12378.n240 gnd 2.02743f
C1275 a_n2686_12378.t2 gnd 0.085436f
C1276 a_n2686_12378.t31 gnd 0.085436f
C1277 a_n2686_12378.n241 gnd 0.747345f
C1278 a_n2686_12378.n242 gnd 2.16299f
C1279 a_n2686_12378.n243 gnd 0.747345f
C1280 a_n2686_12378.t0 gnd 0.085436f
C1281 a_n1455_n3628.n0 gnd 0.029433f
C1282 a_n1455_n3628.n1 gnd 0.048734f
C1283 a_n1455_n3628.n2 gnd 0.029433f
C1284 a_n1455_n3628.n3 gnd 0.350169f
C1285 a_n1455_n3628.n4 gnd 0.029433f
C1286 a_n1455_n3628.n5 gnd 0.048734f
C1287 a_n1455_n3628.n6 gnd 0.029433f
C1288 a_n1455_n3628.n7 gnd 0.350169f
C1289 a_n1455_n3628.n8 gnd 0.029433f
C1290 a_n1455_n3628.n9 gnd 0.048734f
C1291 a_n1455_n3628.n10 gnd 0.029433f
C1292 a_n1455_n3628.n11 gnd 0.350169f
C1293 a_n1455_n3628.n12 gnd 0.029433f
C1294 a_n1455_n3628.n13 gnd 0.048734f
C1295 a_n1455_n3628.n14 gnd 0.029433f
C1296 a_n1455_n3628.n15 gnd 0.029433f
C1297 a_n1455_n3628.n16 gnd 0.029433f
C1298 a_n1455_n3628.n17 gnd 0.364885f
C1299 a_n1455_n3628.n18 gnd 0.029433f
C1300 a_n1455_n3628.n19 gnd 0.029433f
C1301 a_n1455_n3628.n20 gnd 0.364885f
C1302 a_n1455_n3628.n21 gnd 0.029433f
C1303 a_n1455_n3628.n22 gnd 0.029433f
C1304 a_n1455_n3628.n23 gnd 0.364885f
C1305 a_n1455_n3628.n24 gnd 0.029433f
C1306 a_n1455_n3628.n25 gnd 0.029433f
C1307 a_n1455_n3628.n26 gnd 0.364885f
C1308 a_n1455_n3628.n27 gnd 0.029433f
C1309 a_n1455_n3628.n28 gnd 0.029433f
C1310 a_n1455_n3628.n29 gnd 0.364885f
C1311 a_n1455_n3628.n30 gnd 0.029433f
C1312 a_n1455_n3628.n31 gnd 0.029433f
C1313 a_n1455_n3628.n32 gnd 0.364885f
C1314 a_n1455_n3628.n33 gnd 0.029433f
C1315 a_n1455_n3628.n34 gnd 0.029433f
C1316 a_n1455_n3628.n35 gnd 0.364885f
C1317 a_n1455_n3628.n36 gnd 0.029433f
C1318 a_n1455_n3628.n37 gnd 0.029433f
C1319 a_n1455_n3628.n38 gnd 0.364885f
C1320 a_n1455_n3628.n39 gnd 0.062977f
C1321 a_n1455_n3628.n40 gnd 0.018692f
C1322 a_n1455_n3628.n41 gnd 0.008373f
C1323 a_n1455_n3628.n42 gnd 0.007908f
C1324 a_n1455_n3628.n43 gnd 0.018692f
C1325 a_n1455_n3628.n44 gnd 0.008373f
C1326 a_n1455_n3628.n45 gnd 0.007908f
C1327 a_n1455_n3628.n46 gnd 0.020686f
C1328 a_n1455_n3628.t10 gnd 0.069777f
C1329 a_n1455_n3628.t6 gnd 0.069777f
C1330 a_n1455_n3628.n47 gnd 0.558309f
C1331 a_n1455_n3628.n48 gnd 0.347302f
C1332 a_n1455_n3628.n49 gnd 0.020686f
C1333 a_n1455_n3628.n50 gnd 0.007908f
C1334 a_n1455_n3628.n51 gnd 0.018692f
C1335 a_n1455_n3628.n52 gnd 0.008373f
C1336 a_n1455_n3628.n53 gnd 0.007908f
C1337 a_n1455_n3628.n54 gnd 0.018692f
C1338 a_n1455_n3628.n55 gnd 0.008373f
C1339 a_n1455_n3628.n56 gnd 0.062977f
C1340 a_n1455_n3628.t8 gnd 0.030465f
C1341 a_n1455_n3628.n57 gnd 0.014019f
C1342 a_n1455_n3628.n58 gnd 0.011041f
C1343 a_n1455_n3628.n59 gnd 0.007908f
C1344 a_n1455_n3628.n60 gnd 0.007908f
C1345 a_n1455_n3628.n61 gnd 0.008373f
C1346 a_n1455_n3628.n62 gnd 0.018692f
C1347 a_n1455_n3628.n63 gnd 0.018692f
C1348 a_n1455_n3628.n64 gnd 0.008373f
C1349 a_n1455_n3628.n65 gnd 0.007908f
C1350 a_n1455_n3628.n66 gnd 0.007908f
C1351 a_n1455_n3628.n67 gnd 0.008373f
C1352 a_n1455_n3628.n68 gnd 0.018692f
C1353 a_n1455_n3628.n69 gnd 0.040465f
C1354 a_n1455_n3628.n70 gnd 0.008373f
C1355 a_n1455_n3628.n71 gnd 0.007908f
C1356 a_n1455_n3628.n72 gnd 0.034017f
C1357 a_n1455_n3628.n73 gnd 0.026084f
C1358 a_n1455_n3628.n74 gnd 0.610154f
C1359 a_n1455_n3628.t12 gnd 0.069777f
C1360 a_n1455_n3628.t7 gnd 0.069777f
C1361 a_n1455_n3628.n75 gnd 0.558312f
C1362 a_n1455_n3628.n76 gnd 0.347298f
C1363 a_n1455_n3628.n77 gnd 0.020686f
C1364 a_n1455_n3628.n78 gnd 0.007908f
C1365 a_n1455_n3628.n79 gnd 0.018692f
C1366 a_n1455_n3628.n80 gnd 0.008373f
C1367 a_n1455_n3628.n81 gnd 0.007908f
C1368 a_n1455_n3628.n82 gnd 0.018692f
C1369 a_n1455_n3628.n83 gnd 0.008373f
C1370 a_n1455_n3628.n84 gnd 0.062977f
C1371 a_n1455_n3628.t11 gnd 0.030465f
C1372 a_n1455_n3628.n85 gnd 0.014019f
C1373 a_n1455_n3628.n86 gnd 0.011041f
C1374 a_n1455_n3628.n87 gnd 0.007908f
C1375 a_n1455_n3628.n88 gnd 0.007908f
C1376 a_n1455_n3628.n89 gnd 0.008373f
C1377 a_n1455_n3628.n90 gnd 0.018692f
C1378 a_n1455_n3628.n91 gnd 0.018692f
C1379 a_n1455_n3628.n92 gnd 0.008373f
C1380 a_n1455_n3628.n93 gnd 0.007908f
C1381 a_n1455_n3628.n94 gnd 0.007908f
C1382 a_n1455_n3628.n95 gnd 0.008373f
C1383 a_n1455_n3628.n96 gnd 0.018692f
C1384 a_n1455_n3628.n97 gnd 0.040465f
C1385 a_n1455_n3628.n98 gnd 0.008373f
C1386 a_n1455_n3628.n99 gnd 0.007908f
C1387 a_n1455_n3628.n100 gnd 0.034017f
C1388 a_n1455_n3628.n101 gnd 0.026084f
C1389 a_n1455_n3628.n102 gnd 0.16917f
C1390 a_n1455_n3628.n103 gnd 0.020686f
C1391 a_n1455_n3628.n104 gnd 0.007908f
C1392 a_n1455_n3628.n105 gnd 0.018692f
C1393 a_n1455_n3628.n106 gnd 0.008373f
C1394 a_n1455_n3628.n107 gnd 0.007908f
C1395 a_n1455_n3628.n108 gnd 0.018692f
C1396 a_n1455_n3628.n109 gnd 0.008373f
C1397 a_n1455_n3628.n110 gnd 0.062977f
C1398 a_n1455_n3628.t15 gnd 0.030465f
C1399 a_n1455_n3628.n111 gnd 0.014019f
C1400 a_n1455_n3628.n112 gnd 0.011041f
C1401 a_n1455_n3628.n113 gnd 0.007908f
C1402 a_n1455_n3628.n114 gnd 0.007908f
C1403 a_n1455_n3628.n115 gnd 0.008373f
C1404 a_n1455_n3628.n116 gnd 0.018692f
C1405 a_n1455_n3628.n117 gnd 0.018692f
C1406 a_n1455_n3628.n118 gnd 0.008373f
C1407 a_n1455_n3628.n119 gnd 0.007908f
C1408 a_n1455_n3628.n120 gnd 0.007908f
C1409 a_n1455_n3628.n121 gnd 0.008373f
C1410 a_n1455_n3628.n122 gnd 0.018692f
C1411 a_n1455_n3628.n123 gnd 0.040465f
C1412 a_n1455_n3628.n124 gnd 0.008373f
C1413 a_n1455_n3628.n125 gnd 0.007908f
C1414 a_n1455_n3628.n126 gnd 0.034017f
C1415 a_n1455_n3628.n127 gnd 0.026084f
C1416 a_n1455_n3628.n128 gnd 0.16917f
C1417 a_n1455_n3628.t17 gnd 0.069777f
C1418 a_n1455_n3628.t4 gnd 0.069777f
C1419 a_n1455_n3628.n129 gnd 0.558312f
C1420 a_n1455_n3628.n130 gnd 0.347298f
C1421 a_n1455_n3628.n131 gnd 0.020686f
C1422 a_n1455_n3628.n132 gnd 0.007908f
C1423 a_n1455_n3628.n133 gnd 0.018692f
C1424 a_n1455_n3628.n134 gnd 0.008373f
C1425 a_n1455_n3628.n135 gnd 0.007908f
C1426 a_n1455_n3628.n136 gnd 0.018692f
C1427 a_n1455_n3628.n137 gnd 0.008373f
C1428 a_n1455_n3628.n138 gnd 0.062977f
C1429 a_n1455_n3628.t16 gnd 0.030465f
C1430 a_n1455_n3628.n139 gnd 0.014019f
C1431 a_n1455_n3628.n140 gnd 0.011041f
C1432 a_n1455_n3628.n141 gnd 0.007908f
C1433 a_n1455_n3628.n142 gnd 0.007908f
C1434 a_n1455_n3628.n143 gnd 0.008373f
C1435 a_n1455_n3628.n144 gnd 0.018692f
C1436 a_n1455_n3628.n145 gnd 0.018692f
C1437 a_n1455_n3628.n146 gnd 0.008373f
C1438 a_n1455_n3628.n147 gnd 0.007908f
C1439 a_n1455_n3628.n148 gnd 0.007908f
C1440 a_n1455_n3628.n149 gnd 0.008373f
C1441 a_n1455_n3628.n150 gnd 0.018692f
C1442 a_n1455_n3628.n151 gnd 0.040465f
C1443 a_n1455_n3628.n152 gnd 0.008373f
C1444 a_n1455_n3628.n153 gnd 0.007908f
C1445 a_n1455_n3628.n154 gnd 0.034017f
C1446 a_n1455_n3628.n155 gnd 0.026084f
C1447 a_n1455_n3628.n156 gnd 0.610154f
C1448 a_n1455_n3628.n157 gnd 0.020686f
C1449 a_n1455_n3628.n158 gnd 0.007908f
C1450 a_n1455_n3628.n159 gnd 0.018692f
C1451 a_n1455_n3628.n160 gnd 0.008373f
C1452 a_n1455_n3628.n161 gnd 0.007908f
C1453 a_n1455_n3628.n162 gnd 0.018692f
C1454 a_n1455_n3628.n163 gnd 0.008373f
C1455 a_n1455_n3628.n164 gnd 0.062977f
C1456 a_n1455_n3628.t9 gnd 0.030465f
C1457 a_n1455_n3628.n165 gnd 0.014019f
C1458 a_n1455_n3628.n166 gnd 0.011041f
C1459 a_n1455_n3628.n167 gnd 0.007908f
C1460 a_n1455_n3628.n168 gnd 0.007908f
C1461 a_n1455_n3628.n169 gnd 0.008373f
C1462 a_n1455_n3628.n170 gnd 0.018692f
C1463 a_n1455_n3628.n171 gnd 0.018692f
C1464 a_n1455_n3628.n172 gnd 0.008373f
C1465 a_n1455_n3628.n173 gnd 0.007908f
C1466 a_n1455_n3628.n174 gnd 0.007908f
C1467 a_n1455_n3628.n175 gnd 0.008373f
C1468 a_n1455_n3628.n176 gnd 0.018692f
C1469 a_n1455_n3628.n177 gnd 0.040465f
C1470 a_n1455_n3628.n178 gnd 0.008373f
C1471 a_n1455_n3628.n179 gnd 0.007908f
C1472 a_n1455_n3628.n180 gnd 0.026084f
C1473 a_n1455_n3628.n181 gnd 0.381969f
C1474 a_n1455_n3628.n182 gnd 0.714807f
C1475 a_n1455_n3628.n183 gnd 0.020686f
C1476 a_n1455_n3628.n184 gnd 0.007908f
C1477 a_n1455_n3628.n185 gnd 0.018692f
C1478 a_n1455_n3628.n186 gnd 0.008373f
C1479 a_n1455_n3628.n187 gnd 0.007908f
C1480 a_n1455_n3628.n188 gnd 0.018692f
C1481 a_n1455_n3628.n189 gnd 0.008373f
C1482 a_n1455_n3628.n190 gnd 0.062977f
C1483 a_n1455_n3628.t0 gnd 0.030465f
C1484 a_n1455_n3628.n191 gnd 0.014019f
C1485 a_n1455_n3628.n192 gnd 0.011041f
C1486 a_n1455_n3628.n193 gnd 0.007908f
C1487 a_n1455_n3628.n194 gnd 0.007908f
C1488 a_n1455_n3628.n195 gnd 0.008373f
C1489 a_n1455_n3628.n196 gnd 0.018692f
C1490 a_n1455_n3628.n197 gnd 0.018692f
C1491 a_n1455_n3628.n198 gnd 0.008373f
C1492 a_n1455_n3628.n199 gnd 0.007908f
C1493 a_n1455_n3628.n200 gnd 0.007908f
C1494 a_n1455_n3628.n201 gnd 0.008373f
C1495 a_n1455_n3628.n202 gnd 0.018692f
C1496 a_n1455_n3628.n203 gnd 0.040465f
C1497 a_n1455_n3628.n204 gnd 0.008373f
C1498 a_n1455_n3628.n205 gnd 0.007908f
C1499 a_n1455_n3628.n206 gnd 0.034017f
C1500 a_n1455_n3628.n207 gnd 0.122845f
C1501 a_n1455_n3628.n208 gnd 0.89644f
C1502 a_n1455_n3628.n209 gnd 0.020686f
C1503 a_n1455_n3628.n210 gnd 0.007908f
C1504 a_n1455_n3628.n211 gnd 0.018692f
C1505 a_n1455_n3628.n212 gnd 0.008373f
C1506 a_n1455_n3628.n213 gnd 0.007908f
C1507 a_n1455_n3628.n214 gnd 0.018692f
C1508 a_n1455_n3628.n215 gnd 0.008373f
C1509 a_n1455_n3628.n216 gnd 0.062977f
C1510 a_n1455_n3628.t2 gnd 0.030465f
C1511 a_n1455_n3628.n217 gnd 0.014019f
C1512 a_n1455_n3628.n218 gnd 0.011041f
C1513 a_n1455_n3628.n219 gnd 0.007908f
C1514 a_n1455_n3628.n220 gnd 0.007908f
C1515 a_n1455_n3628.n221 gnd 0.008373f
C1516 a_n1455_n3628.n222 gnd 0.018692f
C1517 a_n1455_n3628.n223 gnd 0.018692f
C1518 a_n1455_n3628.n224 gnd 0.008373f
C1519 a_n1455_n3628.n225 gnd 0.007908f
C1520 a_n1455_n3628.n226 gnd 0.007908f
C1521 a_n1455_n3628.n227 gnd 0.008373f
C1522 a_n1455_n3628.n228 gnd 0.018692f
C1523 a_n1455_n3628.n229 gnd 0.040465f
C1524 a_n1455_n3628.n230 gnd 0.008373f
C1525 a_n1455_n3628.n231 gnd 0.007908f
C1526 a_n1455_n3628.n232 gnd 0.034017f
C1527 a_n1455_n3628.n233 gnd 0.121814f
C1528 a_n1455_n3628.n234 gnd 0.708238f
C1529 a_n1455_n3628.n235 gnd 0.020686f
C1530 a_n1455_n3628.n236 gnd 0.007908f
C1531 a_n1455_n3628.n237 gnd 0.018692f
C1532 a_n1455_n3628.n238 gnd 0.008373f
C1533 a_n1455_n3628.n239 gnd 0.007908f
C1534 a_n1455_n3628.n240 gnd 0.018692f
C1535 a_n1455_n3628.n241 gnd 0.008373f
C1536 a_n1455_n3628.n242 gnd 0.062977f
C1537 a_n1455_n3628.t14 gnd 0.030465f
C1538 a_n1455_n3628.n243 gnd 0.014019f
C1539 a_n1455_n3628.n244 gnd 0.011041f
C1540 a_n1455_n3628.n245 gnd 0.007908f
C1541 a_n1455_n3628.n246 gnd 0.007908f
C1542 a_n1455_n3628.n247 gnd 0.008373f
C1543 a_n1455_n3628.n248 gnd 0.018692f
C1544 a_n1455_n3628.n249 gnd 0.018692f
C1545 a_n1455_n3628.n250 gnd 0.008373f
C1546 a_n1455_n3628.n251 gnd 0.007908f
C1547 a_n1455_n3628.n252 gnd 0.007908f
C1548 a_n1455_n3628.n253 gnd 0.008373f
C1549 a_n1455_n3628.n254 gnd 0.018692f
C1550 a_n1455_n3628.n255 gnd 0.040465f
C1551 a_n1455_n3628.n256 gnd 0.008373f
C1552 a_n1455_n3628.n257 gnd 0.007908f
C1553 a_n1455_n3628.n258 gnd 0.034017f
C1554 a_n1455_n3628.n259 gnd 0.121814f
C1555 a_n1455_n3628.n260 gnd 0.933421f
C1556 a_n1455_n3628.n261 gnd 0.020686f
C1557 a_n1455_n3628.n262 gnd 0.007908f
C1558 a_n1455_n3628.n263 gnd 0.018692f
C1559 a_n1455_n3628.n264 gnd 0.008373f
C1560 a_n1455_n3628.n265 gnd 0.007908f
C1561 a_n1455_n3628.n266 gnd 0.018692f
C1562 a_n1455_n3628.n267 gnd 0.008373f
C1563 a_n1455_n3628.n268 gnd 0.062977f
C1564 a_n1455_n3628.t1 gnd 0.030465f
C1565 a_n1455_n3628.n269 gnd 0.014019f
C1566 a_n1455_n3628.n270 gnd 0.011041f
C1567 a_n1455_n3628.n271 gnd 0.007908f
C1568 a_n1455_n3628.n272 gnd 0.007908f
C1569 a_n1455_n3628.n273 gnd 0.008373f
C1570 a_n1455_n3628.n274 gnd 0.018692f
C1571 a_n1455_n3628.n275 gnd 0.018692f
C1572 a_n1455_n3628.n276 gnd 0.008373f
C1573 a_n1455_n3628.n277 gnd 0.007908f
C1574 a_n1455_n3628.n278 gnd 0.007908f
C1575 a_n1455_n3628.n279 gnd 0.008373f
C1576 a_n1455_n3628.n280 gnd 0.018692f
C1577 a_n1455_n3628.n281 gnd 0.040465f
C1578 a_n1455_n3628.n282 gnd 0.008373f
C1579 a_n1455_n3628.n283 gnd 0.007908f
C1580 a_n1455_n3628.n284 gnd 0.034017f
C1581 a_n1455_n3628.n285 gnd 0.121814f
C1582 a_n1455_n3628.n286 gnd 1.26754f
C1583 a_n1455_n3628.n287 gnd 0.80329f
C1584 a_n1455_n3628.n288 gnd 0.020686f
C1585 a_n1455_n3628.n289 gnd 0.007908f
C1586 a_n1455_n3628.n290 gnd 0.018692f
C1587 a_n1455_n3628.n291 gnd 0.008373f
C1588 a_n1455_n3628.n292 gnd 0.007908f
C1589 a_n1455_n3628.n293 gnd 0.018692f
C1590 a_n1455_n3628.n294 gnd 0.008373f
C1591 a_n1455_n3628.n295 gnd 0.062977f
C1592 a_n1455_n3628.t19 gnd 0.030465f
C1593 a_n1455_n3628.n296 gnd 0.014019f
C1594 a_n1455_n3628.n297 gnd 0.011041f
C1595 a_n1455_n3628.n298 gnd 0.007908f
C1596 a_n1455_n3628.n299 gnd 0.007908f
C1597 a_n1455_n3628.n300 gnd 0.008373f
C1598 a_n1455_n3628.n301 gnd 0.018692f
C1599 a_n1455_n3628.n302 gnd 0.018692f
C1600 a_n1455_n3628.n303 gnd 0.008373f
C1601 a_n1455_n3628.n304 gnd 0.007908f
C1602 a_n1455_n3628.n305 gnd 0.007908f
C1603 a_n1455_n3628.n306 gnd 0.008373f
C1604 a_n1455_n3628.n307 gnd 0.018692f
C1605 a_n1455_n3628.n308 gnd 0.040465f
C1606 a_n1455_n3628.n309 gnd 0.008373f
C1607 a_n1455_n3628.n310 gnd 0.007908f
C1608 a_n1455_n3628.n311 gnd 0.026084f
C1609 a_n1455_n3628.n312 gnd 0.381969f
C1610 a_n1455_n3628.t3 gnd 0.069777f
C1611 a_n1455_n3628.t5 gnd 0.069777f
C1612 a_n1455_n3628.n313 gnd 0.558309f
C1613 a_n1455_n3628.n314 gnd 0.347302f
C1614 a_n1455_n3628.n315 gnd 0.020686f
C1615 a_n1455_n3628.n316 gnd 0.007908f
C1616 a_n1455_n3628.n317 gnd 0.018692f
C1617 a_n1455_n3628.n318 gnd 0.008373f
C1618 a_n1455_n3628.n319 gnd 0.007908f
C1619 a_n1455_n3628.n320 gnd 0.018692f
C1620 a_n1455_n3628.n321 gnd 0.008373f
C1621 a_n1455_n3628.n322 gnd 0.062977f
C1622 a_n1455_n3628.t18 gnd 0.030465f
C1623 a_n1455_n3628.n323 gnd 0.014019f
C1624 a_n1455_n3628.n324 gnd 0.011041f
C1625 a_n1455_n3628.n325 gnd 0.007908f
C1626 a_n1455_n3628.n326 gnd 0.007908f
C1627 a_n1455_n3628.n327 gnd 0.008373f
C1628 a_n1455_n3628.n328 gnd 0.018692f
C1629 a_n1455_n3628.n329 gnd 0.018692f
C1630 a_n1455_n3628.n330 gnd 0.008373f
C1631 a_n1455_n3628.n331 gnd 0.007908f
C1632 a_n1455_n3628.n332 gnd 0.007908f
C1633 a_n1455_n3628.n333 gnd 0.008373f
C1634 a_n1455_n3628.n334 gnd 0.018692f
C1635 a_n1455_n3628.n335 gnd 0.040465f
C1636 a_n1455_n3628.n336 gnd 0.008373f
C1637 a_n1455_n3628.n337 gnd 0.007908f
C1638 a_n1455_n3628.n338 gnd 0.026084f
C1639 a_n1455_n3628.n339 gnd 0.16917f
C1640 a_n1455_n3628.n340 gnd 0.16917f
C1641 a_n1455_n3628.n341 gnd 0.026084f
C1642 a_n1455_n3628.n342 gnd 0.007908f
C1643 a_n1455_n3628.n343 gnd 0.008373f
C1644 a_n1455_n3628.n344 gnd 0.040465f
C1645 a_n1455_n3628.n345 gnd 0.018692f
C1646 a_n1455_n3628.n346 gnd 0.008373f
C1647 a_n1455_n3628.n347 gnd 0.007908f
C1648 a_n1455_n3628.n348 gnd 0.007908f
C1649 a_n1455_n3628.n349 gnd 0.008373f
C1650 a_n1455_n3628.n350 gnd 0.018692f
C1651 a_n1455_n3628.n351 gnd 0.018692f
C1652 a_n1455_n3628.n352 gnd 0.008373f
C1653 a_n1455_n3628.n353 gnd 0.007908f
C1654 a_n1455_n3628.n354 gnd 0.350169f
C1655 a_n1455_n3628.n355 gnd 0.007908f
C1656 a_n1455_n3628.n356 gnd 0.011041f
C1657 a_n1455_n3628.n357 gnd 0.014019f
C1658 a_n1455_n3628.t13 gnd 0.030465f
C1659 plus.n0 gnd 0.02619f
C1660 plus.t9 gnd 0.34158f
C1661 plus.t8 gnd 0.311694f
C1662 plus.n1 gnd 0.015852f
C1663 plus.t5 gnd 0.353724f
C1664 plus.n2 gnd 0.156068f
C1665 plus.t12 gnd 0.311694f
C1666 plus.n3 gnd 0.145443f
C1667 plus.n4 gnd 0.026765f
C1668 plus.n5 gnd 0.084024f
C1669 plus.n6 gnd 0.019627f
C1670 plus.n7 gnd 0.019627f
C1671 plus.n8 gnd 0.026765f
C1672 plus.n9 gnd 0.127978f
C1673 plus.n10 gnd 0.026922f
C1674 plus.n11 gnd 0.158341f
C1675 plus.n12 gnd 0.229753f
C1676 plus.n13 gnd 0.02619f
C1677 plus.t11 gnd 0.311694f
C1678 plus.n14 gnd 0.015852f
C1679 plus.t7 gnd 0.353724f
C1680 plus.n15 gnd 0.156068f
C1681 plus.t6 gnd 0.311694f
C1682 plus.n16 gnd 0.145443f
C1683 plus.n17 gnd 0.026765f
C1684 plus.n18 gnd 0.084024f
C1685 plus.n19 gnd 0.019627f
C1686 plus.n20 gnd 0.019627f
C1687 plus.n21 gnd 0.026765f
C1688 plus.n22 gnd 0.127978f
C1689 plus.n23 gnd 0.026922f
C1690 plus.t10 gnd 0.34158f
C1691 plus.n24 gnd 0.158341f
C1692 plus.n25 gnd 0.511565f
C1693 plus.n26 gnd 0.767569f
C1694 plus.t0 gnd 0.033882f
C1695 plus.t1 gnd 0.006051f
C1696 plus.t4 gnd 0.006051f
C1697 plus.n27 gnd 0.019623f
C1698 plus.n28 gnd 0.152334f
C1699 plus.t2 gnd 0.006051f
C1700 plus.t3 gnd 0.006051f
C1701 plus.n29 gnd 0.019623f
C1702 plus.n30 gnd 0.114345f
C1703 plus.n31 gnd 1.87645f
C1704 a_n7677_7899.n0 gnd 0.657706f
C1705 a_n7677_7899.n1 gnd 0.615244f
C1706 a_n7677_7899.n2 gnd 0.657706f
C1707 a_n7677_7899.n3 gnd 0.49764f
C1708 a_n7677_7899.n4 gnd 0.756092f
C1709 a_n7677_7899.n5 gnd 0.039021f
C1710 a_n7677_7899.n6 gnd 0.039021f
C1711 a_n7677_7899.n7 gnd 0.08615f
C1712 a_n7677_7899.n8 gnd 0.050534f
C1713 a_n7677_7899.n9 gnd 0.382272f
C1714 a_n7677_7899.n10 gnd 0.382272f
C1715 a_n7677_7899.n11 gnd 0.382272f
C1716 a_n7677_7899.n12 gnd 0.041194f
C1717 a_n7677_7899.n13 gnd 0.03902f
C1718 a_n7677_7899.n14 gnd 0.041186f
C1719 a_n7677_7899.n15 gnd 0.041186f
C1720 a_n7677_7899.n16 gnd 0.041194f
C1721 a_n7677_7899.n17 gnd 0.03902f
C1722 a_n7677_7899.n18 gnd 0.041186f
C1723 a_n7677_7899.n19 gnd 0.041186f
C1724 a_n7677_7899.n20 gnd 0.041194f
C1725 a_n7677_7899.n21 gnd 0.03902f
C1726 a_n7677_7899.n22 gnd 0.041186f
C1727 a_n7677_7899.n23 gnd 0.387695f
C1728 a_n7677_7899.n24 gnd 0.043833f
C1729 a_n7677_7899.n25 gnd 0.387695f
C1730 a_n7677_7899.n26 gnd 0.043833f
C1731 a_n7677_7899.n27 gnd 0.387695f
C1732 a_n7677_7899.n28 gnd 0.043833f
C1733 a_n7677_7899.n29 gnd 0.050534f
C1734 a_n7677_7899.n30 gnd 0.050534f
C1735 a_n7677_7899.n31 gnd 0.050534f
C1736 a_n7677_7899.n32 gnd 0.043305f
C1737 a_n7677_7899.n33 gnd 0.226953f
C1738 a_n7677_7899.n34 gnd 0.08615f
C1739 a_n7677_7899.n35 gnd 0.042069f
C1740 a_n7677_7899.n36 gnd 0.226953f
C1741 a_n7677_7899.n37 gnd 0.042069f
C1742 a_n7677_7899.n38 gnd 0.08615f
C1743 a_n7677_7899.n39 gnd 0.08615f
C1744 a_n7677_7899.n40 gnd 0.043305f
C1745 a_n7677_7899.n41 gnd 0.08615f
C1746 a_n7677_7899.n42 gnd 0.050534f
C1747 a_n7677_7899.n43 gnd 0.06944f
C1748 a_n7677_7899.n44 gnd 0.042329f
C1749 a_n7677_7899.n45 gnd 0.08615f
C1750 a_n7677_7899.n46 gnd 0.08615f
C1751 a_n7677_7899.n47 gnd 0.08615f
C1752 a_n7677_7899.n48 gnd 0.08615f
C1753 a_n7677_7899.n49 gnd 0.050075f
C1754 a_n7677_7899.n50 gnd 0.069405f
C1755 a_n7677_7899.n51 gnd 0.042616f
C1756 a_n7677_7899.n52 gnd 0.08615f
C1757 a_n7677_7899.n53 gnd 0.100554f
C1758 a_n7677_7899.n54 gnd 0.226953f
C1759 a_n7677_7899.n55 gnd 0.042069f
C1760 a_n7677_7899.n56 gnd 0.08615f
C1761 a_n7677_7899.n57 gnd 0.08615f
C1762 a_n7677_7899.n58 gnd 0.043305f
C1763 a_n7677_7899.n59 gnd 0.08615f
C1764 a_n7677_7899.n60 gnd 0.050534f
C1765 a_n7677_7899.n61 gnd 0.06944f
C1766 a_n7677_7899.n62 gnd 0.042329f
C1767 a_n7677_7899.n63 gnd 0.08615f
C1768 a_n7677_7899.n64 gnd 0.08615f
C1769 a_n7677_7899.n65 gnd 0.08615f
C1770 a_n7677_7899.n66 gnd 0.08615f
C1771 a_n7677_7899.n67 gnd 0.050075f
C1772 a_n7677_7899.n68 gnd 0.069405f
C1773 a_n7677_7899.n69 gnd 0.042616f
C1774 a_n7677_7899.n70 gnd 0.08615f
C1775 a_n7677_7899.n71 gnd 0.100554f
C1776 a_n7677_7899.n72 gnd 0.226953f
C1777 a_n7677_7899.n73 gnd 0.042069f
C1778 a_n7677_7899.n74 gnd 0.08615f
C1779 a_n7677_7899.n75 gnd 0.08615f
C1780 a_n7677_7899.n76 gnd 0.043305f
C1781 a_n7677_7899.n77 gnd 0.08615f
C1782 a_n7677_7899.n78 gnd 0.050534f
C1783 a_n7677_7899.n79 gnd 0.06944f
C1784 a_n7677_7899.n80 gnd 0.042329f
C1785 a_n7677_7899.n81 gnd 0.08615f
C1786 a_n7677_7899.n82 gnd 0.08615f
C1787 a_n7677_7899.n83 gnd 0.08615f
C1788 a_n7677_7899.n84 gnd 0.08615f
C1789 a_n7677_7899.n85 gnd 0.050075f
C1790 a_n7677_7899.n86 gnd 0.069405f
C1791 a_n7677_7899.n87 gnd 0.042616f
C1792 a_n7677_7899.n88 gnd 0.08615f
C1793 a_n7677_7899.n89 gnd 0.100554f
C1794 a_n7677_7899.t7 gnd 0.079673f
C1795 a_n7677_7899.t5 gnd 0.079673f
C1796 a_n7677_7899.t13 gnd 0.079673f
C1797 a_n7677_7899.n90 gnd 0.57569f
C1798 a_n7677_7899.t4 gnd 0.079673f
C1799 a_n7677_7899.t19 gnd 0.079673f
C1800 a_n7677_7899.n91 gnd 0.573011f
C1801 a_n7677_7899.n92 gnd 1.00941f
C1802 a_n7677_7899.t9 gnd 0.079673f
C1803 a_n7677_7899.t10 gnd 0.079673f
C1804 a_n7677_7899.n93 gnd 0.575688f
C1805 a_n7677_7899.t12 gnd 0.079673f
C1806 a_n7677_7899.t6 gnd 0.079673f
C1807 a_n7677_7899.n94 gnd 0.573011f
C1808 a_n7677_7899.n95 gnd 1.00942f
C1809 a_n7677_7899.t11 gnd 0.079673f
C1810 a_n7677_7899.t8 gnd 0.079673f
C1811 a_n7677_7899.n96 gnd 0.573011f
C1812 a_n7677_7899.n97 gnd 2.26042f
C1813 a_n7677_7899.t18 gnd 0.079673f
C1814 a_n7677_7899.t15 gnd 0.079673f
C1815 a_n7677_7899.n98 gnd 0.696936f
C1816 a_n7677_7899.t2 gnd 0.079673f
C1817 a_n7677_7899.t1 gnd 0.079673f
C1818 a_n7677_7899.n99 gnd 0.696933f
C1819 a_n7677_7899.t3 gnd 0.079673f
C1820 a_n7677_7899.t14 gnd 0.079673f
C1821 a_n7677_7899.n100 gnd 0.696933f
C1822 a_n7677_7899.n101 gnd 2.06f
C1823 a_n7677_7899.t17 gnd 0.079673f
C1824 a_n7677_7899.t16 gnd 0.079673f
C1825 a_n7677_7899.n102 gnd 0.695821f
C1826 a_n7677_7899.n103 gnd 1.93461f
C1827 a_n7677_7899.n104 gnd 0.745095f
C1828 a_n7677_7899.t75 gnd 0.80478f
C1829 a_n7677_7899.t54 gnd 0.80478f
C1830 a_n7677_7899.t60 gnd 0.80478f
C1831 a_n7677_7899.t41 gnd 0.80478f
C1832 a_n7677_7899.t73 gnd 0.80478f
C1833 a_n7677_7899.n105 gnd 0.388022f
C1834 a_n7677_7899.t52 gnd 0.80478f
C1835 a_n7677_7899.n106 gnd 0.321107f
C1836 a_n7677_7899.t28 gnd 0.80478f
C1837 a_n7677_7899.n107 gnd 0.399354f
C1838 a_n7677_7899.t58 gnd 0.896702f
C1839 a_n7677_7899.n108 gnd 0.383108f
C1840 a_n7677_7899.n109 gnd 0.069459f
C1841 a_n7677_7899.n110 gnd 0.068241f
C1842 a_n7677_7899.n111 gnd 0.396711f
C1843 a_n7677_7899.n112 gnd 0.321107f
C1844 a_n7677_7899.n113 gnd 0.067992f
C1845 a_n7677_7899.t72 gnd 0.80478f
C1846 a_n7677_7899.n114 gnd 0.396964f
C1847 a_n7677_7899.n115 gnd 0.321107f
C1848 a_n7677_7899.n116 gnd 0.058567f
C1849 a_n7677_7899.t20 gnd 0.87037f
C1850 a_n7677_7899.n117 gnd 0.387472f
C1851 a_n7677_7899.n118 gnd 0.256239f
C1852 a_n7677_7899.t47 gnd 0.80478f
C1853 a_n7677_7899.t25 gnd 0.80478f
C1854 a_n7677_7899.t33 gnd 0.80478f
C1855 a_n7677_7899.t67 gnd 0.80478f
C1856 a_n7677_7899.t46 gnd 0.80478f
C1857 a_n7677_7899.n119 gnd 0.388022f
C1858 a_n7677_7899.t23 gnd 0.80478f
C1859 a_n7677_7899.n120 gnd 0.321107f
C1860 a_n7677_7899.t55 gnd 0.80478f
C1861 a_n7677_7899.n121 gnd 0.399354f
C1862 a_n7677_7899.t31 gnd 0.896702f
C1863 a_n7677_7899.n122 gnd 0.383108f
C1864 a_n7677_7899.n123 gnd 0.069459f
C1865 a_n7677_7899.n124 gnd 0.068241f
C1866 a_n7677_7899.n125 gnd 0.396711f
C1867 a_n7677_7899.n126 gnd 0.321107f
C1868 a_n7677_7899.n127 gnd 0.067992f
C1869 a_n7677_7899.t45 gnd 0.80478f
C1870 a_n7677_7899.n128 gnd 0.396964f
C1871 a_n7677_7899.n129 gnd 0.321107f
C1872 a_n7677_7899.n130 gnd 0.058567f
C1873 a_n7677_7899.t50 gnd 0.87037f
C1874 a_n7677_7899.n131 gnd 0.387472f
C1875 a_n7677_7899.n132 gnd 0.138635f
C1876 a_n7677_7899.n133 gnd 0.689992f
C1877 a_n7677_7899.t26 gnd 0.80478f
C1878 a_n7677_7899.t38 gnd 0.80478f
C1879 a_n7677_7899.t79 gnd 0.80478f
C1880 a_n7677_7899.t35 gnd 0.80478f
C1881 a_n7677_7899.t44 gnd 0.80478f
C1882 a_n7677_7899.n134 gnd 0.388022f
C1883 a_n7677_7899.t53 gnd 0.80478f
C1884 a_n7677_7899.n135 gnd 0.321107f
C1885 a_n7677_7899.t27 gnd 0.80478f
C1886 a_n7677_7899.n136 gnd 0.399354f
C1887 a_n7677_7899.t39 gnd 0.896702f
C1888 a_n7677_7899.n137 gnd 0.383108f
C1889 a_n7677_7899.n138 gnd 0.069459f
C1890 a_n7677_7899.n139 gnd 0.068241f
C1891 a_n7677_7899.n140 gnd 0.396711f
C1892 a_n7677_7899.n141 gnd 0.321107f
C1893 a_n7677_7899.n142 gnd 0.067992f
C1894 a_n7677_7899.t63 gnd 0.80478f
C1895 a_n7677_7899.n143 gnd 0.396964f
C1896 a_n7677_7899.n144 gnd 0.321107f
C1897 a_n7677_7899.n145 gnd 0.058567f
C1898 a_n7677_7899.t32 gnd 0.87037f
C1899 a_n7677_7899.n146 gnd 0.387472f
C1900 a_n7677_7899.n147 gnd 0.138635f
C1901 a_n7677_7899.n148 gnd 1.22705f
C1902 a_n7677_7899.t40 gnd 0.896619f
C1903 a_n7677_7899.t36 gnd 0.80478f
C1904 a_n7677_7899.t69 gnd 0.80478f
C1905 a_n7677_7899.t24 gnd 0.80478f
C1906 a_n7677_7899.n149 gnd 0.387122f
C1907 a_n7677_7899.t78 gnd 0.80478f
C1908 a_n7677_7899.t56 gnd 0.80478f
C1909 a_n7677_7899.t34 gnd 0.80478f
C1910 a_n7677_7899.n150 gnd 0.413311f
C1911 a_n7677_7899.t62 gnd 0.80478f
C1912 a_n7677_7899.n151 gnd 0.423315f
C1913 a_n7677_7899.t43 gnd 0.80478f
C1914 a_n7677_7899.n152 gnd 0.414725f
C1915 a_n7677_7899.t76 gnd 0.896702f
C1916 a_n7677_7899.n153 gnd 0.383107f
C1917 a_n7677_7899.n154 gnd 0.411747f
C1918 a_n7677_7899.n155 gnd 0.376646f
C1919 a_n7677_7899.n156 gnd 0.059137f
C1920 a_n7677_7899.n157 gnd 0.052688f
C1921 a_n7677_7899.n158 gnd 0.423315f
C1922 a_n7677_7899.n159 gnd 0.414738f
C1923 a_n7677_7899.t65 gnd 0.896619f
C1924 a_n7677_7899.t61 gnd 0.80478f
C1925 a_n7677_7899.t42 gnd 0.80478f
C1926 a_n7677_7899.t51 gnd 0.80478f
C1927 a_n7677_7899.n160 gnd 0.387122f
C1928 a_n7677_7899.t49 gnd 0.80478f
C1929 a_n7677_7899.t29 gnd 0.80478f
C1930 a_n7677_7899.t59 gnd 0.80478f
C1931 a_n7677_7899.n161 gnd 0.413311f
C1932 a_n7677_7899.t37 gnd 0.80478f
C1933 a_n7677_7899.n162 gnd 0.423315f
C1934 a_n7677_7899.t71 gnd 0.80478f
C1935 a_n7677_7899.n163 gnd 0.414725f
C1936 a_n7677_7899.t48 gnd 0.896702f
C1937 a_n7677_7899.n164 gnd 0.383107f
C1938 a_n7677_7899.n165 gnd 0.411747f
C1939 a_n7677_7899.n166 gnd 0.376646f
C1940 a_n7677_7899.n167 gnd 0.059137f
C1941 a_n7677_7899.n168 gnd 0.052688f
C1942 a_n7677_7899.n169 gnd 0.423315f
C1943 a_n7677_7899.n170 gnd 0.414738f
C1944 a_n7677_7899.n171 gnd 0.689992f
C1945 a_n7677_7899.t74 gnd 0.896619f
C1946 a_n7677_7899.t68 gnd 0.80478f
C1947 a_n7677_7899.t22 gnd 0.80478f
C1948 a_n7677_7899.t66 gnd 0.80478f
C1949 a_n7677_7899.n172 gnd 0.413312f
C1950 a_n7677_7899.t64 gnd 0.80478f
C1951 a_n7677_7899.t77 gnd 0.80478f
C1952 a_n7677_7899.t30 gnd 0.80478f
C1953 a_n7677_7899.n173 gnd 0.388022f
C1954 a_n7677_7899.t57 gnd 0.80478f
C1955 a_n7677_7899.n174 gnd 0.321107f
C1956 a_n7677_7899.t70 gnd 0.80478f
C1957 a_n7677_7899.n175 gnd 0.399354f
C1958 a_n7677_7899.t21 gnd 0.896702f
C1959 a_n7677_7899.n176 gnd 0.383107f
C1960 a_n7677_7899.n177 gnd 0.069459f
C1961 a_n7677_7899.n178 gnd 0.068241f
C1962 a_n7677_7899.n179 gnd 0.411747f
C1963 a_n7677_7899.n180 gnd 0.411747f
C1964 a_n7677_7899.n181 gnd 0.423315f
C1965 a_n7677_7899.n182 gnd 0.414738f
C1966 a_n7677_7899.n183 gnd 1.02545f
C1967 a_n7677_7899.n184 gnd 11.371099f
C1968 a_n7677_7899.n185 gnd 3.62931f
C1969 a_n7677_7899.n186 gnd 4.84333f
C1970 a_n7677_7899.n187 gnd 1.55922f
C1971 a_n7677_7899.n188 gnd 0.573011f
C1972 a_n7677_7899.t0 gnd 0.079673f
C1973 CSoutput.n0 gnd 0.037226f
C1974 CSoutput.t104 gnd 0.246243f
C1975 CSoutput.n1 gnd 0.111191f
C1976 CSoutput.n2 gnd 0.037226f
C1977 CSoutput.t110 gnd 0.246243f
C1978 CSoutput.n3 gnd 0.029505f
C1979 CSoutput.n4 gnd 0.037226f
C1980 CSoutput.t100 gnd 0.246243f
C1981 CSoutput.n5 gnd 0.025442f
C1982 CSoutput.n6 gnd 0.037226f
C1983 CSoutput.t107 gnd 0.246243f
C1984 CSoutput.t113 gnd 0.246243f
C1985 CSoutput.n7 gnd 0.109979f
C1986 CSoutput.n8 gnd 0.037226f
C1987 CSoutput.t112 gnd 0.246243f
C1988 CSoutput.n9 gnd 0.024258f
C1989 CSoutput.n10 gnd 0.037226f
C1990 CSoutput.t103 gnd 0.246243f
C1991 CSoutput.t102 gnd 0.246243f
C1992 CSoutput.n11 gnd 0.109979f
C1993 CSoutput.n12 gnd 0.037226f
C1994 CSoutput.t108 gnd 0.246243f
C1995 CSoutput.n13 gnd 0.025442f
C1996 CSoutput.n14 gnd 0.037226f
C1997 CSoutput.t96 gnd 0.246243f
C1998 CSoutput.t101 gnd 0.246243f
C1999 CSoutput.n15 gnd 0.109979f
C2000 CSoutput.n16 gnd 0.037226f
C2001 CSoutput.t105 gnd 0.246243f
C2002 CSoutput.n17 gnd 0.027174f
C2003 CSoutput.t94 gnd 0.294267f
C2004 CSoutput.t111 gnd 0.246243f
C2005 CSoutput.n18 gnd 0.140401f
C2006 CSoutput.n19 gnd 0.136237f
C2007 CSoutput.n20 gnd 0.158052f
C2008 CSoutput.n21 gnd 0.037226f
C2009 CSoutput.n22 gnd 0.031069f
C2010 CSoutput.n23 gnd 0.109979f
C2011 CSoutput.n24 gnd 0.02995f
C2012 CSoutput.n25 gnd 0.029505f
C2013 CSoutput.n26 gnd 0.037226f
C2014 CSoutput.n27 gnd 0.037226f
C2015 CSoutput.n28 gnd 0.030831f
C2016 CSoutput.n29 gnd 0.026176f
C2017 CSoutput.n30 gnd 0.112428f
C2018 CSoutput.n31 gnd 0.026536f
C2019 CSoutput.n32 gnd 0.037226f
C2020 CSoutput.n33 gnd 0.037226f
C2021 CSoutput.n34 gnd 0.037226f
C2022 CSoutput.n35 gnd 0.030502f
C2023 CSoutput.n36 gnd 0.109979f
C2024 CSoutput.n37 gnd 0.029171f
C2025 CSoutput.n38 gnd 0.030284f
C2026 CSoutput.n39 gnd 0.037226f
C2027 CSoutput.n40 gnd 0.037226f
C2028 CSoutput.n41 gnd 0.031063f
C2029 CSoutput.n42 gnd 0.028392f
C2030 CSoutput.n43 gnd 0.109979f
C2031 CSoutput.n44 gnd 0.029112f
C2032 CSoutput.n45 gnd 0.037226f
C2033 CSoutput.n46 gnd 0.037226f
C2034 CSoutput.n47 gnd 0.037226f
C2035 CSoutput.n48 gnd 0.029112f
C2036 CSoutput.n49 gnd 0.109979f
C2037 CSoutput.n50 gnd 0.028392f
C2038 CSoutput.n51 gnd 0.031063f
C2039 CSoutput.n52 gnd 0.037226f
C2040 CSoutput.n53 gnd 0.037226f
C2041 CSoutput.n54 gnd 0.030284f
C2042 CSoutput.n55 gnd 0.029171f
C2043 CSoutput.n56 gnd 0.109979f
C2044 CSoutput.n57 gnd 0.030502f
C2045 CSoutput.n58 gnd 0.037226f
C2046 CSoutput.n59 gnd 0.037226f
C2047 CSoutput.n60 gnd 0.037226f
C2048 CSoutput.n61 gnd 0.026536f
C2049 CSoutput.n62 gnd 0.112428f
C2050 CSoutput.n63 gnd 0.026176f
C2051 CSoutput.t92 gnd 0.246243f
C2052 CSoutput.n64 gnd 0.109979f
C2053 CSoutput.n65 gnd 0.030831f
C2054 CSoutput.n66 gnd 0.037226f
C2055 CSoutput.n67 gnd 0.037226f
C2056 CSoutput.n68 gnd 0.037226f
C2057 CSoutput.n69 gnd 0.02995f
C2058 CSoutput.n70 gnd 0.109979f
C2059 CSoutput.n71 gnd 0.031069f
C2060 CSoutput.n72 gnd 0.027174f
C2061 CSoutput.n73 gnd 0.037226f
C2062 CSoutput.n74 gnd 0.037226f
C2063 CSoutput.n75 gnd 0.028181f
C2064 CSoutput.n76 gnd 0.016737f
C2065 CSoutput.t95 gnd 0.276672f
C2066 CSoutput.n77 gnd 0.137439f
C2067 CSoutput.n78 gnd 0.588091f
C2068 CSoutput.t80 gnd 0.04063f
C2069 CSoutput.t16 gnd 0.04063f
C2070 CSoutput.n79 gnd 0.303036f
C2071 CSoutput.t39 gnd 0.04063f
C2072 CSoutput.t12 gnd 0.04063f
C2073 CSoutput.n80 gnd 0.301763f
C2074 CSoutput.n81 gnd 0.448989f
C2075 CSoutput.t7 gnd 0.04063f
C2076 CSoutput.t29 gnd 0.04063f
C2077 CSoutput.n82 gnd 0.301763f
C2078 CSoutput.n83 gnd 0.222173f
C2079 CSoutput.t19 gnd 0.04063f
C2080 CSoutput.t20 gnd 0.04063f
C2081 CSoutput.n84 gnd 0.301763f
C2082 CSoutput.n85 gnd 0.222173f
C2083 CSoutput.t13 gnd 0.04063f
C2084 CSoutput.t81 gnd 0.04063f
C2085 CSoutput.n86 gnd 0.301763f
C2086 CSoutput.n87 gnd 0.361433f
C2087 CSoutput.t15 gnd 0.04063f
C2088 CSoutput.t82 gnd 0.04063f
C2089 CSoutput.n88 gnd 0.303036f
C2090 CSoutput.t21 gnd 0.04063f
C2091 CSoutput.t73 gnd 0.04063f
C2092 CSoutput.n89 gnd 0.301763f
C2093 CSoutput.n90 gnd 0.448989f
C2094 CSoutput.t37 gnd 0.04063f
C2095 CSoutput.t17 gnd 0.04063f
C2096 CSoutput.n91 gnd 0.301763f
C2097 CSoutput.n92 gnd 0.222173f
C2098 CSoutput.t91 gnd 0.04063f
C2099 CSoutput.t14 gnd 0.04063f
C2100 CSoutput.n93 gnd 0.301763f
C2101 CSoutput.n94 gnd 0.222173f
C2102 CSoutput.t27 gnd 0.04063f
C2103 CSoutput.t75 gnd 0.04063f
C2104 CSoutput.n95 gnd 0.301763f
C2105 CSoutput.n96 gnd 0.307633f
C2106 CSoutput.n97 gnd 0.315799f
C2107 CSoutput.t85 gnd 0.04063f
C2108 CSoutput.t34 gnd 0.04063f
C2109 CSoutput.n98 gnd 0.303036f
C2110 CSoutput.t76 gnd 0.04063f
C2111 CSoutput.t74 gnd 0.04063f
C2112 CSoutput.n99 gnd 0.301763f
C2113 CSoutput.n100 gnd 0.448989f
C2114 CSoutput.t11 gnd 0.04063f
C2115 CSoutput.t24 gnd 0.04063f
C2116 CSoutput.n101 gnd 0.301763f
C2117 CSoutput.n102 gnd 0.222173f
C2118 CSoutput.t18 gnd 0.04063f
C2119 CSoutput.t77 gnd 0.04063f
C2120 CSoutput.n103 gnd 0.301763f
C2121 CSoutput.n104 gnd 0.222173f
C2122 CSoutput.t4 gnd 0.04063f
C2123 CSoutput.t86 gnd 0.04063f
C2124 CSoutput.n105 gnd 0.301763f
C2125 CSoutput.n106 gnd 0.307633f
C2126 CSoutput.n107 gnd 0.338139f
C2127 CSoutput.n108 gnd 6.21298f
C2128 CSoutput.n110 gnd 0.658525f
C2129 CSoutput.n111 gnd 0.493894f
C2130 CSoutput.n112 gnd 0.658525f
C2131 CSoutput.n113 gnd 0.658525f
C2132 CSoutput.n114 gnd 1.77295f
C2133 CSoutput.n115 gnd 0.658525f
C2134 CSoutput.n116 gnd 0.658525f
C2135 CSoutput.t106 gnd 0.823156f
C2136 CSoutput.n117 gnd 0.658525f
C2137 CSoutput.n118 gnd 0.658525f
C2138 CSoutput.n122 gnd 0.658525f
C2139 CSoutput.n126 gnd 0.658525f
C2140 CSoutput.n127 gnd 0.658525f
C2141 CSoutput.n129 gnd 0.658525f
C2142 CSoutput.n134 gnd 0.658525f
C2143 CSoutput.n136 gnd 0.658525f
C2144 CSoutput.n137 gnd 0.658525f
C2145 CSoutput.n139 gnd 0.658525f
C2146 CSoutput.n140 gnd 0.658525f
C2147 CSoutput.n142 gnd 0.658525f
C2148 CSoutput.t97 gnd 11.003901f
C2149 CSoutput.n144 gnd 0.658525f
C2150 CSoutput.n145 gnd 0.493894f
C2151 CSoutput.n146 gnd 0.658525f
C2152 CSoutput.n147 gnd 0.658525f
C2153 CSoutput.n148 gnd 1.77295f
C2154 CSoutput.n149 gnd 0.658525f
C2155 CSoutput.n150 gnd 0.658525f
C2156 CSoutput.t109 gnd 0.823156f
C2157 CSoutput.n151 gnd 0.658525f
C2158 CSoutput.n152 gnd 0.658525f
C2159 CSoutput.n156 gnd 0.658525f
C2160 CSoutput.n160 gnd 0.658525f
C2161 CSoutput.n161 gnd 0.658525f
C2162 CSoutput.n163 gnd 0.658525f
C2163 CSoutput.n168 gnd 0.658525f
C2164 CSoutput.n170 gnd 0.658525f
C2165 CSoutput.n171 gnd 0.658525f
C2166 CSoutput.n173 gnd 0.658525f
C2167 CSoutput.n174 gnd 0.658525f
C2168 CSoutput.n176 gnd 0.658525f
C2169 CSoutput.n177 gnd 0.493894f
C2170 CSoutput.n179 gnd 0.658525f
C2171 CSoutput.n180 gnd 0.493894f
C2172 CSoutput.n181 gnd 0.658525f
C2173 CSoutput.n182 gnd 0.658525f
C2174 CSoutput.n183 gnd 1.77295f
C2175 CSoutput.n184 gnd 0.658525f
C2176 CSoutput.n185 gnd 0.658525f
C2177 CSoutput.t99 gnd 0.823156f
C2178 CSoutput.n186 gnd 0.658525f
C2179 CSoutput.n187 gnd 1.77295f
C2180 CSoutput.n189 gnd 0.658525f
C2181 CSoutput.n190 gnd 0.658525f
C2182 CSoutput.n192 gnd 0.658525f
C2183 CSoutput.n193 gnd 0.658525f
C2184 CSoutput.t93 gnd 10.8246f
C2185 CSoutput.t98 gnd 11.003901f
C2186 CSoutput.n199 gnd 2.06589f
C2187 CSoutput.n200 gnd 8.41568f
C2188 CSoutput.n201 gnd 8.76783f
C2189 CSoutput.n206 gnd 2.23792f
C2190 CSoutput.n212 gnd 0.658525f
C2191 CSoutput.n214 gnd 0.658525f
C2192 CSoutput.n216 gnd 0.658525f
C2193 CSoutput.n218 gnd 0.658525f
C2194 CSoutput.n220 gnd 0.658525f
C2195 CSoutput.n226 gnd 0.658525f
C2196 CSoutput.n233 gnd 1.20814f
C2197 CSoutput.n234 gnd 1.20814f
C2198 CSoutput.n235 gnd 0.658525f
C2199 CSoutput.n236 gnd 0.658525f
C2200 CSoutput.n238 gnd 0.493894f
C2201 CSoutput.n239 gnd 0.422976f
C2202 CSoutput.n241 gnd 0.493894f
C2203 CSoutput.n242 gnd 0.422976f
C2204 CSoutput.n243 gnd 0.493894f
C2205 CSoutput.n245 gnd 0.658525f
C2206 CSoutput.n247 gnd 1.77295f
C2207 CSoutput.n248 gnd 2.06589f
C2208 CSoutput.n249 gnd 7.74026f
C2209 CSoutput.n251 gnd 0.493894f
C2210 CSoutput.n252 gnd 1.27082f
C2211 CSoutput.n253 gnd 0.493894f
C2212 CSoutput.n255 gnd 0.658525f
C2213 CSoutput.n257 gnd 1.77295f
C2214 CSoutput.n258 gnd 3.86436f
C2215 CSoutput.t84 gnd 0.04063f
C2216 CSoutput.t30 gnd 0.04063f
C2217 CSoutput.n259 gnd 0.303036f
C2218 CSoutput.t90 gnd 0.04063f
C2219 CSoutput.t36 gnd 0.04063f
C2220 CSoutput.n260 gnd 0.301763f
C2221 CSoutput.n261 gnd 0.448989f
C2222 CSoutput.t32 gnd 0.04063f
C2223 CSoutput.t23 gnd 0.04063f
C2224 CSoutput.n262 gnd 0.301763f
C2225 CSoutput.n263 gnd 0.222173f
C2226 CSoutput.t26 gnd 0.04063f
C2227 CSoutput.t1 gnd 0.04063f
C2228 CSoutput.n264 gnd 0.301763f
C2229 CSoutput.n265 gnd 0.222173f
C2230 CSoutput.t88 gnd 0.04063f
C2231 CSoutput.t35 gnd 0.04063f
C2232 CSoutput.n266 gnd 0.301763f
C2233 CSoutput.n267 gnd 0.361433f
C2234 CSoutput.t33 gnd 0.04063f
C2235 CSoutput.t25 gnd 0.04063f
C2236 CSoutput.n268 gnd 0.303036f
C2237 CSoutput.t8 gnd 0.04063f
C2238 CSoutput.t83 gnd 0.04063f
C2239 CSoutput.n269 gnd 0.301763f
C2240 CSoutput.n270 gnd 0.448989f
C2241 CSoutput.t79 gnd 0.04063f
C2242 CSoutput.t87 gnd 0.04063f
C2243 CSoutput.n271 gnd 0.301763f
C2244 CSoutput.n272 gnd 0.222173f
C2245 CSoutput.t5 gnd 0.04063f
C2246 CSoutput.t3 gnd 0.04063f
C2247 CSoutput.n273 gnd 0.301763f
C2248 CSoutput.n274 gnd 0.222173f
C2249 CSoutput.t89 gnd 0.04063f
C2250 CSoutput.t78 gnd 0.04063f
C2251 CSoutput.n275 gnd 0.301763f
C2252 CSoutput.n276 gnd 0.307633f
C2253 CSoutput.n277 gnd 0.315799f
C2254 CSoutput.t10 gnd 0.04063f
C2255 CSoutput.t2 gnd 0.04063f
C2256 CSoutput.n278 gnd 0.303036f
C2257 CSoutput.t31 gnd 0.04063f
C2258 CSoutput.t72 gnd 0.04063f
C2259 CSoutput.n279 gnd 0.301763f
C2260 CSoutput.n280 gnd 0.448989f
C2261 CSoutput.t28 gnd 0.04063f
C2262 CSoutput.t0 gnd 0.04063f
C2263 CSoutput.n281 gnd 0.301763f
C2264 CSoutput.n282 gnd 0.222173f
C2265 CSoutput.t6 gnd 0.04063f
C2266 CSoutput.t38 gnd 0.04063f
C2267 CSoutput.n283 gnd 0.301763f
C2268 CSoutput.n284 gnd 0.222173f
C2269 CSoutput.t9 gnd 0.04063f
C2270 CSoutput.t22 gnd 0.04063f
C2271 CSoutput.n285 gnd 0.301762f
C2272 CSoutput.n286 gnd 0.307634f
C2273 CSoutput.n287 gnd 0.338139f
C2274 CSoutput.n288 gnd 8.902969f
C2275 CSoutput.t48 gnd 0.034826f
C2276 CSoutput.t67 gnd 0.034826f
C2277 CSoutput.n289 gnd 0.307125f
C2278 CSoutput.t63 gnd 0.034826f
C2279 CSoutput.t68 gnd 0.034826f
C2280 CSoutput.n290 gnd 0.304149f
C2281 CSoutput.n291 gnd 0.495279f
C2282 CSoutput.t52 gnd 0.034826f
C2283 CSoutput.t51 gnd 0.034826f
C2284 CSoutput.n292 gnd 0.304149f
C2285 CSoutput.n293 gnd 0.246169f
C2286 CSoutput.t61 gnd 0.034826f
C2287 CSoutput.t59 gnd 0.034826f
C2288 CSoutput.n294 gnd 0.304149f
C2289 CSoutput.n295 gnd 0.372497f
C2290 CSoutput.t55 gnd 0.034826f
C2291 CSoutput.t41 gnd 0.034826f
C2292 CSoutput.n296 gnd 0.307125f
C2293 CSoutput.t40 gnd 0.034826f
C2294 CSoutput.t42 gnd 0.034826f
C2295 CSoutput.n297 gnd 0.304149f
C2296 CSoutput.n298 gnd 0.495279f
C2297 CSoutput.t57 gnd 0.034826f
C2298 CSoutput.t56 gnd 0.034826f
C2299 CSoutput.n299 gnd 0.304149f
C2300 CSoutput.n300 gnd 0.246169f
C2301 CSoutput.t66 gnd 0.034826f
C2302 CSoutput.t64 gnd 0.034826f
C2303 CSoutput.n301 gnd 0.304149f
C2304 CSoutput.n302 gnd 0.325318f
C2305 CSoutput.n303 gnd 0.461201f
C2306 CSoutput.n304 gnd 9.03697f
C2307 CSoutput.t45 gnd 0.034826f
C2308 CSoutput.t70 gnd 0.034826f
C2309 CSoutput.n305 gnd 0.307125f
C2310 CSoutput.t46 gnd 0.034826f
C2311 CSoutput.t54 gnd 0.034826f
C2312 CSoutput.n306 gnd 0.304149f
C2313 CSoutput.n307 gnd 0.495279f
C2314 CSoutput.t60 gnd 0.034826f
C2315 CSoutput.t62 gnd 0.034826f
C2316 CSoutput.n308 gnd 0.304149f
C2317 CSoutput.n309 gnd 0.246169f
C2318 CSoutput.t47 gnd 0.034826f
C2319 CSoutput.t71 gnd 0.034826f
C2320 CSoutput.n310 gnd 0.304149f
C2321 CSoutput.n311 gnd 0.372497f
C2322 CSoutput.t49 gnd 0.034826f
C2323 CSoutput.t43 gnd 0.034826f
C2324 CSoutput.n312 gnd 0.307125f
C2325 CSoutput.t50 gnd 0.034826f
C2326 CSoutput.t58 gnd 0.034826f
C2327 CSoutput.n313 gnd 0.304149f
C2328 CSoutput.n314 gnd 0.495279f
C2329 CSoutput.t65 gnd 0.034826f
C2330 CSoutput.t69 gnd 0.034826f
C2331 CSoutput.n315 gnd 0.304149f
C2332 CSoutput.n316 gnd 0.246169f
C2333 CSoutput.t53 gnd 0.034826f
C2334 CSoutput.t44 gnd 0.034826f
C2335 CSoutput.n317 gnd 0.304149f
C2336 CSoutput.n318 gnd 0.325318f
C2337 CSoutput.n319 gnd 0.461201f
C2338 CSoutput.n320 gnd 5.45873f
C2339 CSoutput.n321 gnd 10.9191f
C2340 commonsourceibias.n0 gnd 0.00802f
C2341 commonsourceibias.t55 gnd 0.193208f
C2342 commonsourceibias.n1 gnd 0.008674f
C2343 commonsourceibias.n2 gnd 0.006083f
C2344 commonsourceibias.t36 gnd 0.193208f
C2345 commonsourceibias.n3 gnd 0.005572f
C2346 commonsourceibias.n4 gnd 0.006083f
C2347 commonsourceibias.t40 gnd 0.193208f
C2348 commonsourceibias.n5 gnd 0.011335f
C2349 commonsourceibias.n6 gnd 0.006083f
C2350 commonsourceibias.t35 gnd 0.193208f
C2351 commonsourceibias.n7 gnd 0.07376f
C2352 commonsourceibias.n8 gnd 0.005314f
C2353 commonsourceibias.n9 gnd 0.010334f
C2354 commonsourceibias.n10 gnd 0.00802f
C2355 commonsourceibias.t30 gnd 0.193208f
C2356 commonsourceibias.n11 gnd 0.008674f
C2357 commonsourceibias.n12 gnd 0.006083f
C2358 commonsourceibias.t16 gnd 0.193208f
C2359 commonsourceibias.n13 gnd 0.005572f
C2360 commonsourceibias.n14 gnd 0.006083f
C2361 commonsourceibias.t22 gnd 0.193208f
C2362 commonsourceibias.n15 gnd 0.011335f
C2363 commonsourceibias.n16 gnd 0.006083f
C2364 commonsourceibias.t18 gnd 0.193208f
C2365 commonsourceibias.n17 gnd 0.07376f
C2366 commonsourceibias.n18 gnd 0.006083f
C2367 commonsourceibias.n19 gnd 0.010334f
C2368 commonsourceibias.n20 gnd 0.006083f
C2369 commonsourceibias.t4 gnd 0.193208f
C2370 commonsourceibias.n21 gnd 0.07376f
C2371 commonsourceibias.n22 gnd 0.011335f
C2372 commonsourceibias.n23 gnd 0.006083f
C2373 commonsourceibias.t10 gnd 0.193208f
C2374 commonsourceibias.n24 gnd 0.005572f
C2375 commonsourceibias.n25 gnd 0.045538f
C2376 commonsourceibias.t12 gnd 0.193208f
C2377 commonsourceibias.t26 gnd 0.223789f
C2378 commonsourceibias.n26 gnd 0.088589f
C2379 commonsourceibias.n27 gnd 0.086415f
C2380 commonsourceibias.n28 gnd 0.006547f
C2381 commonsourceibias.n29 gnd 0.01217f
C2382 commonsourceibias.n30 gnd 0.006083f
C2383 commonsourceibias.n31 gnd 0.006083f
C2384 commonsourceibias.n32 gnd 0.006083f
C2385 commonsourceibias.n33 gnd 0.011225f
C2386 commonsourceibias.n34 gnd 0.008552f
C2387 commonsourceibias.n35 gnd 0.07376f
C2388 commonsourceibias.n36 gnd 0.00844f
C2389 commonsourceibias.n37 gnd 0.006083f
C2390 commonsourceibias.n38 gnd 0.006083f
C2391 commonsourceibias.n39 gnd 0.006083f
C2392 commonsourceibias.n40 gnd 0.005428f
C2393 commonsourceibias.n41 gnd 0.012203f
C2394 commonsourceibias.n42 gnd 0.006658f
C2395 commonsourceibias.n43 gnd 0.006083f
C2396 commonsourceibias.n44 gnd 0.006083f
C2397 commonsourceibias.n45 gnd 0.006083f
C2398 commonsourceibias.n46 gnd 0.008843f
C2399 commonsourceibias.n47 gnd 0.008843f
C2400 commonsourceibias.n48 gnd 0.010334f
C2401 commonsourceibias.n49 gnd 0.006083f
C2402 commonsourceibias.n50 gnd 0.006083f
C2403 commonsourceibias.n51 gnd 0.006658f
C2404 commonsourceibias.n52 gnd 0.012203f
C2405 commonsourceibias.n53 gnd 0.005428f
C2406 commonsourceibias.n54 gnd 0.006083f
C2407 commonsourceibias.n55 gnd 0.006083f
C2408 commonsourceibias.n56 gnd 0.006083f
C2409 commonsourceibias.n57 gnd 0.00844f
C2410 commonsourceibias.n58 gnd 0.07376f
C2411 commonsourceibias.n59 gnd 0.008552f
C2412 commonsourceibias.n60 gnd 0.011225f
C2413 commonsourceibias.n61 gnd 0.006083f
C2414 commonsourceibias.n62 gnd 0.006083f
C2415 commonsourceibias.n63 gnd 0.006083f
C2416 commonsourceibias.n64 gnd 0.01217f
C2417 commonsourceibias.n65 gnd 0.006547f
C2418 commonsourceibias.n66 gnd 0.07376f
C2419 commonsourceibias.n67 gnd 0.010445f
C2420 commonsourceibias.n68 gnd 0.006083f
C2421 commonsourceibias.n69 gnd 0.006083f
C2422 commonsourceibias.n70 gnd 0.006083f
C2423 commonsourceibias.n71 gnd 0.009011f
C2424 commonsourceibias.n72 gnd 0.010223f
C2425 commonsourceibias.n73 gnd 0.09231f
C2426 commonsourceibias.n74 gnd 0.061098f
C2427 commonsourceibias.t31 gnd 0.011251f
C2428 commonsourceibias.t17 gnd 0.011251f
C2429 commonsourceibias.n75 gnd 0.098265f
C2430 commonsourceibias.n76 gnd 0.121797f
C2431 commonsourceibias.t23 gnd 0.011251f
C2432 commonsourceibias.t19 gnd 0.011251f
C2433 commonsourceibias.n77 gnd 0.098265f
C2434 commonsourceibias.n78 gnd 0.064174f
C2435 commonsourceibias.t13 gnd 0.011251f
C2436 commonsourceibias.t27 gnd 0.011251f
C2437 commonsourceibias.n79 gnd 0.099226f
C2438 commonsourceibias.t5 gnd 0.011251f
C2439 commonsourceibias.t11 gnd 0.011251f
C2440 commonsourceibias.n80 gnd 0.098265f
C2441 commonsourceibias.n81 gnd 0.144656f
C2442 commonsourceibias.n82 gnd 0.067084f
C2443 commonsourceibias.n83 gnd 0.03937f
C2444 commonsourceibias.n84 gnd 0.006083f
C2445 commonsourceibias.t51 gnd 0.193208f
C2446 commonsourceibias.n85 gnd 0.07376f
C2447 commonsourceibias.n86 gnd 0.011335f
C2448 commonsourceibias.n87 gnd 0.006083f
C2449 commonsourceibias.t52 gnd 0.193208f
C2450 commonsourceibias.n88 gnd 0.005572f
C2451 commonsourceibias.n89 gnd 0.045538f
C2452 commonsourceibias.t42 gnd 0.193208f
C2453 commonsourceibias.t44 gnd 0.223789f
C2454 commonsourceibias.n90 gnd 0.088589f
C2455 commonsourceibias.n91 gnd 0.086415f
C2456 commonsourceibias.n92 gnd 0.006547f
C2457 commonsourceibias.n93 gnd 0.01217f
C2458 commonsourceibias.n94 gnd 0.006083f
C2459 commonsourceibias.n95 gnd 0.006083f
C2460 commonsourceibias.n96 gnd 0.006083f
C2461 commonsourceibias.n97 gnd 0.011225f
C2462 commonsourceibias.n98 gnd 0.008552f
C2463 commonsourceibias.n99 gnd 0.07376f
C2464 commonsourceibias.n100 gnd 0.00844f
C2465 commonsourceibias.n101 gnd 0.006083f
C2466 commonsourceibias.n102 gnd 0.006083f
C2467 commonsourceibias.n103 gnd 0.006083f
C2468 commonsourceibias.n104 gnd 0.005428f
C2469 commonsourceibias.n105 gnd 0.012203f
C2470 commonsourceibias.n106 gnd 0.006658f
C2471 commonsourceibias.n107 gnd 0.006083f
C2472 commonsourceibias.n108 gnd 0.006083f
C2473 commonsourceibias.n109 gnd 0.005314f
C2474 commonsourceibias.n110 gnd 0.008843f
C2475 commonsourceibias.n111 gnd 0.008843f
C2476 commonsourceibias.n112 gnd 0.010334f
C2477 commonsourceibias.n113 gnd 0.006083f
C2478 commonsourceibias.n114 gnd 0.006083f
C2479 commonsourceibias.n115 gnd 0.006658f
C2480 commonsourceibias.n116 gnd 0.012203f
C2481 commonsourceibias.n117 gnd 0.005428f
C2482 commonsourceibias.n118 gnd 0.006083f
C2483 commonsourceibias.n119 gnd 0.006083f
C2484 commonsourceibias.n120 gnd 0.006083f
C2485 commonsourceibias.n121 gnd 0.00844f
C2486 commonsourceibias.n122 gnd 0.07376f
C2487 commonsourceibias.n123 gnd 0.008552f
C2488 commonsourceibias.n124 gnd 0.011225f
C2489 commonsourceibias.n125 gnd 0.006083f
C2490 commonsourceibias.n126 gnd 0.006083f
C2491 commonsourceibias.n127 gnd 0.006083f
C2492 commonsourceibias.n128 gnd 0.01217f
C2493 commonsourceibias.n129 gnd 0.006547f
C2494 commonsourceibias.n130 gnd 0.07376f
C2495 commonsourceibias.n131 gnd 0.010445f
C2496 commonsourceibias.n132 gnd 0.006083f
C2497 commonsourceibias.n133 gnd 0.006083f
C2498 commonsourceibias.n134 gnd 0.006083f
C2499 commonsourceibias.n135 gnd 0.009011f
C2500 commonsourceibias.n136 gnd 0.010223f
C2501 commonsourceibias.n137 gnd 0.09231f
C2502 commonsourceibias.n138 gnd 0.036167f
C2503 commonsourceibias.n139 gnd 0.00802f
C2504 commonsourceibias.t48 gnd 0.193208f
C2505 commonsourceibias.n140 gnd 0.008674f
C2506 commonsourceibias.n141 gnd 0.006083f
C2507 commonsourceibias.t62 gnd 0.193208f
C2508 commonsourceibias.n142 gnd 0.005572f
C2509 commonsourceibias.n143 gnd 0.006083f
C2510 commonsourceibias.t63 gnd 0.193208f
C2511 commonsourceibias.n144 gnd 0.011335f
C2512 commonsourceibias.n145 gnd 0.006083f
C2513 commonsourceibias.t61 gnd 0.193208f
C2514 commonsourceibias.n146 gnd 0.07376f
C2515 commonsourceibias.n147 gnd 0.006083f
C2516 commonsourceibias.n148 gnd 0.010334f
C2517 commonsourceibias.n149 gnd 0.006083f
C2518 commonsourceibias.t46 gnd 0.193208f
C2519 commonsourceibias.n150 gnd 0.07376f
C2520 commonsourceibias.n151 gnd 0.011335f
C2521 commonsourceibias.n152 gnd 0.006083f
C2522 commonsourceibias.t47 gnd 0.193208f
C2523 commonsourceibias.n153 gnd 0.005572f
C2524 commonsourceibias.n154 gnd 0.045538f
C2525 commonsourceibias.t37 gnd 0.193208f
C2526 commonsourceibias.t39 gnd 0.223789f
C2527 commonsourceibias.n155 gnd 0.088589f
C2528 commonsourceibias.n156 gnd 0.086415f
C2529 commonsourceibias.n157 gnd 0.006547f
C2530 commonsourceibias.n158 gnd 0.01217f
C2531 commonsourceibias.n159 gnd 0.006083f
C2532 commonsourceibias.n160 gnd 0.006083f
C2533 commonsourceibias.n161 gnd 0.006083f
C2534 commonsourceibias.n162 gnd 0.011225f
C2535 commonsourceibias.n163 gnd 0.008552f
C2536 commonsourceibias.n164 gnd 0.07376f
C2537 commonsourceibias.n165 gnd 0.00844f
C2538 commonsourceibias.n166 gnd 0.006083f
C2539 commonsourceibias.n167 gnd 0.006083f
C2540 commonsourceibias.n168 gnd 0.006083f
C2541 commonsourceibias.n169 gnd 0.005428f
C2542 commonsourceibias.n170 gnd 0.012203f
C2543 commonsourceibias.n171 gnd 0.006658f
C2544 commonsourceibias.n172 gnd 0.006083f
C2545 commonsourceibias.n173 gnd 0.006083f
C2546 commonsourceibias.n174 gnd 0.006083f
C2547 commonsourceibias.n175 gnd 0.008843f
C2548 commonsourceibias.n176 gnd 0.008843f
C2549 commonsourceibias.n177 gnd 0.010334f
C2550 commonsourceibias.n178 gnd 0.006083f
C2551 commonsourceibias.n179 gnd 0.006083f
C2552 commonsourceibias.n180 gnd 0.006658f
C2553 commonsourceibias.n181 gnd 0.012203f
C2554 commonsourceibias.n182 gnd 0.005428f
C2555 commonsourceibias.n183 gnd 0.006083f
C2556 commonsourceibias.n184 gnd 0.006083f
C2557 commonsourceibias.n185 gnd 0.006083f
C2558 commonsourceibias.n186 gnd 0.00844f
C2559 commonsourceibias.n187 gnd 0.07376f
C2560 commonsourceibias.n188 gnd 0.008552f
C2561 commonsourceibias.n189 gnd 0.011225f
C2562 commonsourceibias.n190 gnd 0.006083f
C2563 commonsourceibias.n191 gnd 0.006083f
C2564 commonsourceibias.n192 gnd 0.006083f
C2565 commonsourceibias.n193 gnd 0.01217f
C2566 commonsourceibias.n194 gnd 0.006547f
C2567 commonsourceibias.n195 gnd 0.07376f
C2568 commonsourceibias.n196 gnd 0.010445f
C2569 commonsourceibias.n197 gnd 0.006083f
C2570 commonsourceibias.n198 gnd 0.006083f
C2571 commonsourceibias.n199 gnd 0.006083f
C2572 commonsourceibias.n200 gnd 0.009011f
C2573 commonsourceibias.n201 gnd 0.010223f
C2574 commonsourceibias.n202 gnd 0.09231f
C2575 commonsourceibias.n203 gnd 0.022047f
C2576 commonsourceibias.n204 gnd 0.272706f
C2577 commonsourceibias.n205 gnd 0.00802f
C2578 commonsourceibias.t33 gnd 0.193208f
C2579 commonsourceibias.n206 gnd 0.008674f
C2580 commonsourceibias.n207 gnd 0.006083f
C2581 commonsourceibias.t58 gnd 0.193208f
C2582 commonsourceibias.n208 gnd 0.005572f
C2583 commonsourceibias.n209 gnd 0.006083f
C2584 commonsourceibias.t49 gnd 0.193208f
C2585 commonsourceibias.n210 gnd 0.011335f
C2586 commonsourceibias.n211 gnd 0.006083f
C2587 commonsourceibias.t57 gnd 0.193208f
C2588 commonsourceibias.n212 gnd 0.07376f
C2589 commonsourceibias.n213 gnd 0.005314f
C2590 commonsourceibias.n214 gnd 0.010334f
C2591 commonsourceibias.n215 gnd 0.006083f
C2592 commonsourceibias.n216 gnd 0.011335f
C2593 commonsourceibias.n217 gnd 0.006083f
C2594 commonsourceibias.t43 gnd 0.193208f
C2595 commonsourceibias.n218 gnd 0.005572f
C2596 commonsourceibias.n219 gnd 0.045538f
C2597 commonsourceibias.t32 gnd 0.193208f
C2598 commonsourceibias.t56 gnd 0.223789f
C2599 commonsourceibias.n220 gnd 0.088589f
C2600 commonsourceibias.n221 gnd 0.086415f
C2601 commonsourceibias.n222 gnd 0.006547f
C2602 commonsourceibias.n223 gnd 0.01217f
C2603 commonsourceibias.n224 gnd 0.006083f
C2604 commonsourceibias.n225 gnd 0.006083f
C2605 commonsourceibias.n226 gnd 0.006083f
C2606 commonsourceibias.n227 gnd 0.011225f
C2607 commonsourceibias.n228 gnd 0.008552f
C2608 commonsourceibias.n229 gnd 0.07376f
C2609 commonsourceibias.n230 gnd 0.00844f
C2610 commonsourceibias.n231 gnd 0.006083f
C2611 commonsourceibias.n232 gnd 0.006083f
C2612 commonsourceibias.n233 gnd 0.006083f
C2613 commonsourceibias.n234 gnd 0.005428f
C2614 commonsourceibias.n235 gnd 0.012203f
C2615 commonsourceibias.t41 gnd 0.193208f
C2616 commonsourceibias.n236 gnd 0.07376f
C2617 commonsourceibias.n237 gnd 0.006658f
C2618 commonsourceibias.n238 gnd 0.006083f
C2619 commonsourceibias.n239 gnd 0.006083f
C2620 commonsourceibias.t25 gnd 0.011251f
C2621 commonsourceibias.t7 gnd 0.011251f
C2622 commonsourceibias.n240 gnd 0.099226f
C2623 commonsourceibias.t21 gnd 0.011251f
C2624 commonsourceibias.t9 gnd 0.011251f
C2625 commonsourceibias.n241 gnd 0.098265f
C2626 commonsourceibias.n242 gnd 0.144656f
C2627 commonsourceibias.n243 gnd 0.00802f
C2628 commonsourceibias.t28 gnd 0.193208f
C2629 commonsourceibias.n244 gnd 0.008674f
C2630 commonsourceibias.n245 gnd 0.006083f
C2631 commonsourceibias.t14 gnd 0.193208f
C2632 commonsourceibias.n246 gnd 0.005572f
C2633 commonsourceibias.n247 gnd 0.006083f
C2634 commonsourceibias.t2 gnd 0.193208f
C2635 commonsourceibias.n248 gnd 0.011335f
C2636 commonsourceibias.n249 gnd 0.006083f
C2637 commonsourceibias.t0 gnd 0.193208f
C2638 commonsourceibias.n250 gnd 0.07376f
C2639 commonsourceibias.n251 gnd 0.006083f
C2640 commonsourceibias.n252 gnd 0.010334f
C2641 commonsourceibias.n253 gnd 0.006083f
C2642 commonsourceibias.n254 gnd 0.011335f
C2643 commonsourceibias.n255 gnd 0.006083f
C2644 commonsourceibias.t20 gnd 0.193208f
C2645 commonsourceibias.n256 gnd 0.005572f
C2646 commonsourceibias.n257 gnd 0.045538f
C2647 commonsourceibias.t6 gnd 0.193208f
C2648 commonsourceibias.t24 gnd 0.223789f
C2649 commonsourceibias.n258 gnd 0.088589f
C2650 commonsourceibias.n259 gnd 0.086415f
C2651 commonsourceibias.n260 gnd 0.006547f
C2652 commonsourceibias.n261 gnd 0.01217f
C2653 commonsourceibias.n262 gnd 0.006083f
C2654 commonsourceibias.n263 gnd 0.006083f
C2655 commonsourceibias.n264 gnd 0.006083f
C2656 commonsourceibias.n265 gnd 0.011225f
C2657 commonsourceibias.n266 gnd 0.008552f
C2658 commonsourceibias.n267 gnd 0.07376f
C2659 commonsourceibias.n268 gnd 0.00844f
C2660 commonsourceibias.n269 gnd 0.006083f
C2661 commonsourceibias.n270 gnd 0.006083f
C2662 commonsourceibias.n271 gnd 0.006083f
C2663 commonsourceibias.n272 gnd 0.005428f
C2664 commonsourceibias.n273 gnd 0.012203f
C2665 commonsourceibias.t8 gnd 0.193208f
C2666 commonsourceibias.n274 gnd 0.07376f
C2667 commonsourceibias.n275 gnd 0.006658f
C2668 commonsourceibias.n276 gnd 0.006083f
C2669 commonsourceibias.n277 gnd 0.006083f
C2670 commonsourceibias.n278 gnd 0.006083f
C2671 commonsourceibias.n279 gnd 0.008843f
C2672 commonsourceibias.n280 gnd 0.008843f
C2673 commonsourceibias.n281 gnd 0.010334f
C2674 commonsourceibias.n282 gnd 0.006083f
C2675 commonsourceibias.n283 gnd 0.006083f
C2676 commonsourceibias.n284 gnd 0.006658f
C2677 commonsourceibias.n285 gnd 0.012203f
C2678 commonsourceibias.n286 gnd 0.005428f
C2679 commonsourceibias.n287 gnd 0.006083f
C2680 commonsourceibias.n288 gnd 0.006083f
C2681 commonsourceibias.n289 gnd 0.006083f
C2682 commonsourceibias.n290 gnd 0.00844f
C2683 commonsourceibias.n291 gnd 0.07376f
C2684 commonsourceibias.n292 gnd 0.008552f
C2685 commonsourceibias.n293 gnd 0.011225f
C2686 commonsourceibias.n294 gnd 0.006083f
C2687 commonsourceibias.n295 gnd 0.006083f
C2688 commonsourceibias.n296 gnd 0.006083f
C2689 commonsourceibias.n297 gnd 0.01217f
C2690 commonsourceibias.n298 gnd 0.006547f
C2691 commonsourceibias.n299 gnd 0.07376f
C2692 commonsourceibias.n300 gnd 0.010445f
C2693 commonsourceibias.n301 gnd 0.006083f
C2694 commonsourceibias.n302 gnd 0.006083f
C2695 commonsourceibias.n303 gnd 0.006083f
C2696 commonsourceibias.n304 gnd 0.009011f
C2697 commonsourceibias.n305 gnd 0.010223f
C2698 commonsourceibias.n306 gnd 0.09231f
C2699 commonsourceibias.n307 gnd 0.061098f
C2700 commonsourceibias.t15 gnd 0.011251f
C2701 commonsourceibias.t29 gnd 0.011251f
C2702 commonsourceibias.n308 gnd 0.098265f
C2703 commonsourceibias.n309 gnd 0.121797f
C2704 commonsourceibias.t1 gnd 0.011251f
C2705 commonsourceibias.t3 gnd 0.011251f
C2706 commonsourceibias.n310 gnd 0.098265f
C2707 commonsourceibias.n311 gnd 0.064174f
C2708 commonsourceibias.n312 gnd 0.067084f
C2709 commonsourceibias.n313 gnd 0.03937f
C2710 commonsourceibias.n314 gnd 0.005314f
C2711 commonsourceibias.n315 gnd 0.008843f
C2712 commonsourceibias.n316 gnd 0.008843f
C2713 commonsourceibias.n317 gnd 0.010334f
C2714 commonsourceibias.n318 gnd 0.006083f
C2715 commonsourceibias.n319 gnd 0.006083f
C2716 commonsourceibias.n320 gnd 0.006658f
C2717 commonsourceibias.n321 gnd 0.012203f
C2718 commonsourceibias.n322 gnd 0.005428f
C2719 commonsourceibias.n323 gnd 0.006083f
C2720 commonsourceibias.n324 gnd 0.006083f
C2721 commonsourceibias.n325 gnd 0.006083f
C2722 commonsourceibias.n326 gnd 0.00844f
C2723 commonsourceibias.n327 gnd 0.07376f
C2724 commonsourceibias.n328 gnd 0.008552f
C2725 commonsourceibias.n329 gnd 0.011225f
C2726 commonsourceibias.n330 gnd 0.006083f
C2727 commonsourceibias.n331 gnd 0.006083f
C2728 commonsourceibias.n332 gnd 0.006083f
C2729 commonsourceibias.n333 gnd 0.01217f
C2730 commonsourceibias.n334 gnd 0.006547f
C2731 commonsourceibias.n335 gnd 0.07376f
C2732 commonsourceibias.n336 gnd 0.010445f
C2733 commonsourceibias.n337 gnd 0.006083f
C2734 commonsourceibias.n338 gnd 0.006083f
C2735 commonsourceibias.n339 gnd 0.006083f
C2736 commonsourceibias.n340 gnd 0.009011f
C2737 commonsourceibias.n341 gnd 0.010223f
C2738 commonsourceibias.n342 gnd 0.09231f
C2739 commonsourceibias.n343 gnd 0.036167f
C2740 commonsourceibias.n344 gnd 0.00802f
C2741 commonsourceibias.t60 gnd 0.193208f
C2742 commonsourceibias.n345 gnd 0.008674f
C2743 commonsourceibias.n346 gnd 0.006083f
C2744 commonsourceibias.t54 gnd 0.193208f
C2745 commonsourceibias.n347 gnd 0.005572f
C2746 commonsourceibias.n348 gnd 0.006083f
C2747 commonsourceibias.t45 gnd 0.193208f
C2748 commonsourceibias.n349 gnd 0.011335f
C2749 commonsourceibias.n350 gnd 0.006083f
C2750 commonsourceibias.t53 gnd 0.193208f
C2751 commonsourceibias.n351 gnd 0.07376f
C2752 commonsourceibias.n352 gnd 0.006083f
C2753 commonsourceibias.n353 gnd 0.010334f
C2754 commonsourceibias.n354 gnd 0.006083f
C2755 commonsourceibias.n355 gnd 0.011335f
C2756 commonsourceibias.n356 gnd 0.006083f
C2757 commonsourceibias.t38 gnd 0.193208f
C2758 commonsourceibias.n357 gnd 0.005572f
C2759 commonsourceibias.n358 gnd 0.045538f
C2760 commonsourceibias.t59 gnd 0.193208f
C2761 commonsourceibias.t50 gnd 0.223789f
C2762 commonsourceibias.n359 gnd 0.088589f
C2763 commonsourceibias.n360 gnd 0.086415f
C2764 commonsourceibias.n361 gnd 0.006547f
C2765 commonsourceibias.n362 gnd 0.01217f
C2766 commonsourceibias.n363 gnd 0.006083f
C2767 commonsourceibias.n364 gnd 0.006083f
C2768 commonsourceibias.n365 gnd 0.006083f
C2769 commonsourceibias.n366 gnd 0.011225f
C2770 commonsourceibias.n367 gnd 0.008552f
C2771 commonsourceibias.n368 gnd 0.07376f
C2772 commonsourceibias.n369 gnd 0.00844f
C2773 commonsourceibias.n370 gnd 0.006083f
C2774 commonsourceibias.n371 gnd 0.006083f
C2775 commonsourceibias.n372 gnd 0.006083f
C2776 commonsourceibias.n373 gnd 0.005428f
C2777 commonsourceibias.n374 gnd 0.012203f
C2778 commonsourceibias.t34 gnd 0.193208f
C2779 commonsourceibias.n375 gnd 0.07376f
C2780 commonsourceibias.n376 gnd 0.006658f
C2781 commonsourceibias.n377 gnd 0.006083f
C2782 commonsourceibias.n378 gnd 0.006083f
C2783 commonsourceibias.n379 gnd 0.006083f
C2784 commonsourceibias.n380 gnd 0.008843f
C2785 commonsourceibias.n381 gnd 0.008843f
C2786 commonsourceibias.n382 gnd 0.010334f
C2787 commonsourceibias.n383 gnd 0.006083f
C2788 commonsourceibias.n384 gnd 0.006083f
C2789 commonsourceibias.n385 gnd 0.006658f
C2790 commonsourceibias.n386 gnd 0.012203f
C2791 commonsourceibias.n387 gnd 0.005428f
C2792 commonsourceibias.n388 gnd 0.006083f
C2793 commonsourceibias.n389 gnd 0.006083f
C2794 commonsourceibias.n390 gnd 0.006083f
C2795 commonsourceibias.n391 gnd 0.00844f
C2796 commonsourceibias.n392 gnd 0.07376f
C2797 commonsourceibias.n393 gnd 0.008552f
C2798 commonsourceibias.n394 gnd 0.011225f
C2799 commonsourceibias.n395 gnd 0.006083f
C2800 commonsourceibias.n396 gnd 0.006083f
C2801 commonsourceibias.n397 gnd 0.006083f
C2802 commonsourceibias.n398 gnd 0.01217f
C2803 commonsourceibias.n399 gnd 0.006547f
C2804 commonsourceibias.n400 gnd 0.07376f
C2805 commonsourceibias.n401 gnd 0.010445f
C2806 commonsourceibias.n402 gnd 0.006083f
C2807 commonsourceibias.n403 gnd 0.006083f
C2808 commonsourceibias.n404 gnd 0.006083f
C2809 commonsourceibias.n405 gnd 0.009011f
C2810 commonsourceibias.n406 gnd 0.010223f
C2811 commonsourceibias.n407 gnd 0.09231f
C2812 commonsourceibias.n408 gnd 0.022047f
C2813 commonsourceibias.n409 gnd 0.159609f
C2814 commonsourceibias.n410 gnd 3.00565f
C2815 vdd.t136 gnd 0.022905f
C2816 vdd.t195 gnd 0.022905f
C2817 vdd.n0 gnd 0.165504f
C2818 vdd.t143 gnd 0.022905f
C2819 vdd.t202 gnd 0.022905f
C2820 vdd.n1 gnd 0.164733f
C2821 vdd.n2 gnd 0.299855f
C2822 vdd.t139 gnd 0.022905f
C2823 vdd.t123 gnd 0.022905f
C2824 vdd.n3 gnd 0.164733f
C2825 vdd.n4 gnd 0.153198f
C2826 vdd.t182 gnd 0.022905f
C2827 vdd.t166 gnd 0.022905f
C2828 vdd.n5 gnd 0.164733f
C2829 vdd.n6 gnd 0.138705f
C2830 vdd.t141 gnd 0.022905f
C2831 vdd.t125 gnd 0.022905f
C2832 vdd.n7 gnd 0.165504f
C2833 vdd.t180 gnd 0.022905f
C2834 vdd.t178 gnd 0.022905f
C2835 vdd.n8 gnd 0.164733f
C2836 vdd.n9 gnd 0.299855f
C2837 vdd.t2 gnd 0.022905f
C2838 vdd.t146 gnd 0.022905f
C2839 vdd.n10 gnd 0.164733f
C2840 vdd.n11 gnd 0.153198f
C2841 vdd.t175 gnd 0.022905f
C2842 vdd.t215 gnd 0.022905f
C2843 vdd.n12 gnd 0.164733f
C2844 vdd.n13 gnd 0.138705f
C2845 vdd.n14 gnd 0.091946f
C2846 vdd.t209 gnd 0.019088f
C2847 vdd.t13 gnd 0.019088f
C2848 vdd.n15 gnd 0.175693f
C2849 vdd.t198 gnd 0.019088f
C2850 vdd.t109 gnd 0.019088f
C2851 vdd.n16 gnd 0.175179f
C2852 vdd.n17 gnd 0.304865f
C2853 vdd.t197 gnd 0.019088f
C2854 vdd.t106 gnd 0.019088f
C2855 vdd.n18 gnd 0.175179f
C2856 vdd.n19 gnd 0.126127f
C2857 vdd.t12 gnd 0.019088f
C2858 vdd.t126 gnd 0.019088f
C2859 vdd.n20 gnd 0.175693f
C2860 vdd.t196 gnd 0.019088f
C2861 vdd.t107 gnd 0.019088f
C2862 vdd.n21 gnd 0.175179f
C2863 vdd.n22 gnd 0.304865f
C2864 vdd.t8 gnd 0.019088f
C2865 vdd.t108 gnd 0.019088f
C2866 vdd.n23 gnd 0.175179f
C2867 vdd.n24 gnd 0.126127f
C2868 vdd.t207 gnd 0.019088f
C2869 vdd.t208 gnd 0.019088f
C2870 vdd.n25 gnd 0.175179f
C2871 vdd.t127 gnd 0.019088f
C2872 vdd.t128 gnd 0.019088f
C2873 vdd.n26 gnd 0.175179f
C2874 vdd.n27 gnd 18.204899f
C2875 vdd.n28 gnd 6.93796f
C2876 vdd.t203 gnd 0.232594f
C2877 vdd.t159 gnd 0.026723f
C2878 vdd.t212 gnd 0.026723f
C2879 vdd.n29 gnd 0.171507f
C2880 vdd.n30 gnd 0.304174f
C2881 vdd.t168 gnd 0.026723f
C2882 vdd.t161 gnd 0.026723f
C2883 vdd.n31 gnd 0.171507f
C2884 vdd.n32 gnd 0.162092f
C2885 vdd.t149 gnd 0.026723f
C2886 vdd.t152 gnd 0.026723f
C2887 vdd.n33 gnd 0.171507f
C2888 vdd.n34 gnd 0.162092f
C2889 vdd.t7 gnd 0.026723f
C2890 vdd.t210 gnd 0.026723f
C2891 vdd.n35 gnd 0.171507f
C2892 vdd.n36 gnd 0.162092f
C2893 vdd.t164 gnd 0.23156f
C2894 vdd.n37 gnd 0.204642f
C2895 vdd.t162 gnd 0.232594f
C2896 vdd.t151 gnd 0.026723f
C2897 vdd.t24 gnd 0.026723f
C2898 vdd.n38 gnd 0.171507f
C2899 vdd.n39 gnd 0.304174f
C2900 vdd.t200 gnd 0.026723f
C2901 vdd.t191 gnd 0.026723f
C2902 vdd.n40 gnd 0.171507f
C2903 vdd.n41 gnd 0.162092f
C2904 vdd.t206 gnd 0.026723f
C2905 vdd.t17 gnd 0.026723f
C2906 vdd.n42 gnd 0.171507f
C2907 vdd.n43 gnd 0.162092f
C2908 vdd.t11 gnd 0.026723f
C2909 vdd.t211 gnd 0.026723f
C2910 vdd.n44 gnd 0.171507f
C2911 vdd.n45 gnd 0.162092f
C2912 vdd.t190 gnd 0.23156f
C2913 vdd.n46 gnd 0.169939f
C2914 vdd.n47 gnd 0.194956f
C2915 vdd.t104 gnd 0.232594f
C2916 vdd.t10 gnd 0.026723f
C2917 vdd.t160 gnd 0.026723f
C2918 vdd.n48 gnd 0.171507f
C2919 vdd.n49 gnd 0.304174f
C2920 vdd.t183 gnd 0.026723f
C2921 vdd.t157 gnd 0.026723f
C2922 vdd.n50 gnd 0.171507f
C2923 vdd.n51 gnd 0.162092f
C2924 vdd.t5 gnd 0.026723f
C2925 vdd.t18 gnd 0.026723f
C2926 vdd.n52 gnd 0.171507f
C2927 vdd.n53 gnd 0.162092f
C2928 vdd.t170 gnd 0.026723f
C2929 vdd.t26 gnd 0.026723f
C2930 vdd.n54 gnd 0.171507f
C2931 vdd.n55 gnd 0.162092f
C2932 vdd.t148 gnd 0.23156f
C2933 vdd.n56 gnd 0.169939f
C2934 vdd.n57 gnd 0.213388f
C2935 vdd.n58 gnd 0.007291f
C2936 vdd.n59 gnd 0.009486f
C2937 vdd.n60 gnd 0.007635f
C2938 vdd.n61 gnd 0.007635f
C2939 vdd.n62 gnd 0.009486f
C2940 vdd.n63 gnd 0.009486f
C2941 vdd.n64 gnd 0.696487f
C2942 vdd.n65 gnd 0.009486f
C2943 vdd.n66 gnd 0.009486f
C2944 vdd.n67 gnd 0.009486f
C2945 vdd.n68 gnd 0.567085f
C2946 vdd.n69 gnd 0.009486f
C2947 vdd.n70 gnd 0.009486f
C2948 vdd.n71 gnd 0.009486f
C2949 vdd.n72 gnd 0.009486f
C2950 vdd.n73 gnd 0.007635f
C2951 vdd.n74 gnd 0.009486f
C2952 vdd.t16 gnd 0.380594f
C2953 vdd.n75 gnd 0.009486f
C2954 vdd.n76 gnd 0.009486f
C2955 vdd.n77 gnd 0.009486f
C2956 vdd.t6 gnd 0.380594f
C2957 vdd.n78 gnd 0.009486f
C2958 vdd.n79 gnd 0.009486f
C2959 vdd.n80 gnd 0.009486f
C2960 vdd.n81 gnd 0.009486f
C2961 vdd.n82 gnd 0.009486f
C2962 vdd.n83 gnd 0.007635f
C2963 vdd.n84 gnd 0.009486f
C2964 vdd.n85 gnd 0.704099f
C2965 vdd.n86 gnd 0.009486f
C2966 vdd.n87 gnd 0.009486f
C2967 vdd.n88 gnd 0.009486f
C2968 vdd.n89 gnd 0.559473f
C2969 vdd.n90 gnd 0.009486f
C2970 vdd.n91 gnd 0.009486f
C2971 vdd.n92 gnd 0.009486f
C2972 vdd.n93 gnd 0.009486f
C2973 vdd.n94 gnd 0.009486f
C2974 vdd.n95 gnd 0.007635f
C2975 vdd.n96 gnd 0.009486f
C2976 vdd.t147 gnd 0.380594f
C2977 vdd.n97 gnd 0.009486f
C2978 vdd.n98 gnd 0.009486f
C2979 vdd.n99 gnd 0.009486f
C2980 vdd.n100 gnd 0.761188f
C2981 vdd.n101 gnd 0.009486f
C2982 vdd.n102 gnd 0.009486f
C2983 vdd.n103 gnd 0.009486f
C2984 vdd.n104 gnd 0.009486f
C2985 vdd.n105 gnd 0.009486f
C2986 vdd.n106 gnd 0.007635f
C2987 vdd.n107 gnd 0.009486f
C2988 vdd.n108 gnd 0.009486f
C2989 vdd.n109 gnd 0.009486f
C2990 vdd.n110 gnd 0.021312f
C2991 vdd.n111 gnd 1.65558f
C2992 vdd.n112 gnd 0.021375f
C2993 vdd.n113 gnd 0.009486f
C2994 vdd.n114 gnd 0.009486f
C2995 vdd.n116 gnd 0.009486f
C2996 vdd.n117 gnd 0.009486f
C2997 vdd.n118 gnd 0.007635f
C2998 vdd.n119 gnd 0.007635f
C2999 vdd.n120 gnd 0.009486f
C3000 vdd.n121 gnd 0.009486f
C3001 vdd.n122 gnd 0.009486f
C3002 vdd.n123 gnd 0.009486f
C3003 vdd.n124 gnd 0.009486f
C3004 vdd.n125 gnd 0.009486f
C3005 vdd.n126 gnd 0.007635f
C3006 vdd.n128 gnd 0.009486f
C3007 vdd.n129 gnd 0.009486f
C3008 vdd.n130 gnd 0.009486f
C3009 vdd.n131 gnd 0.009486f
C3010 vdd.n132 gnd 0.009486f
C3011 vdd.n133 gnd 0.007635f
C3012 vdd.n135 gnd 0.009486f
C3013 vdd.n136 gnd 0.009486f
C3014 vdd.n137 gnd 0.009486f
C3015 vdd.n138 gnd 0.009486f
C3016 vdd.n139 gnd 0.009486f
C3017 vdd.n140 gnd 0.006375f
C3018 vdd.n142 gnd 0.009486f
C3019 vdd.n143 gnd 0.006375f
C3020 vdd.t73 gnd 0.194308f
C3021 vdd.t72 gnd 0.203627f
C3022 vdd.t71 gnd 0.283884f
C3023 vdd.n144 gnd 0.096222f
C3024 vdd.n145 gnd 0.055169f
C3025 vdd.n146 gnd 0.009486f
C3026 vdd.n147 gnd 0.009486f
C3027 vdd.n148 gnd 0.007635f
C3028 vdd.n150 gnd 0.009486f
C3029 vdd.n151 gnd 0.009486f
C3030 vdd.n152 gnd 0.009486f
C3031 vdd.n153 gnd 0.009486f
C3032 vdd.n154 gnd 0.007635f
C3033 vdd.n156 gnd 0.009486f
C3034 vdd.n157 gnd 0.009486f
C3035 vdd.n158 gnd 0.009486f
C3036 vdd.n159 gnd 0.009486f
C3037 vdd.n160 gnd 0.009486f
C3038 vdd.n161 gnd 0.007635f
C3039 vdd.n163 gnd 0.009486f
C3040 vdd.n164 gnd 0.009486f
C3041 vdd.n165 gnd 0.009486f
C3042 vdd.n166 gnd 0.009486f
C3043 vdd.n167 gnd 0.009486f
C3044 vdd.n168 gnd 0.007635f
C3045 vdd.n170 gnd 0.009486f
C3046 vdd.n171 gnd 0.009486f
C3047 vdd.n172 gnd 0.009486f
C3048 vdd.n173 gnd 0.009486f
C3049 vdd.n174 gnd 0.009486f
C3050 vdd.n175 gnd 0.005192f
C3051 vdd.n177 gnd 0.009486f
C3052 vdd.n178 gnd 0.007559f
C3053 vdd.t41 gnd 0.194308f
C3054 vdd.t40 gnd 0.203627f
C3055 vdd.t39 gnd 0.283884f
C3056 vdd.n179 gnd 0.096222f
C3057 vdd.n180 gnd 0.055169f
C3058 vdd.n181 gnd 0.009486f
C3059 vdd.n182 gnd 0.009486f
C3060 vdd.n183 gnd 0.007635f
C3061 vdd.n185 gnd 0.009486f
C3062 vdd.n186 gnd 0.009486f
C3063 vdd.n187 gnd 0.009486f
C3064 vdd.n188 gnd 0.009486f
C3065 vdd.n189 gnd 0.007635f
C3066 vdd.n191 gnd 0.009486f
C3067 vdd.n192 gnd 0.009486f
C3068 vdd.n193 gnd 0.009486f
C3069 vdd.n194 gnd 0.009486f
C3070 vdd.n195 gnd 0.009486f
C3071 vdd.n196 gnd 0.007635f
C3072 vdd.n198 gnd 0.009486f
C3073 vdd.n199 gnd 0.009486f
C3074 vdd.n200 gnd 0.009486f
C3075 vdd.n201 gnd 0.009486f
C3076 vdd.n202 gnd 0.009486f
C3077 vdd.n203 gnd 0.007635f
C3078 vdd.n205 gnd 0.009486f
C3079 vdd.n206 gnd 0.009486f
C3080 vdd.n207 gnd 0.009486f
C3081 vdd.n208 gnd 0.009486f
C3082 vdd.n209 gnd 0.009486f
C3083 vdd.n210 gnd 0.004008f
C3084 vdd.t30 gnd 0.194308f
C3085 vdd.t29 gnd 0.203627f
C3086 vdd.t27 gnd 0.283884f
C3087 vdd.n212 gnd 0.096222f
C3088 vdd.n213 gnd 0.055169f
C3089 vdd.n214 gnd 0.011796f
C3090 vdd.n215 gnd 0.009486f
C3091 vdd.n216 gnd 0.009486f
C3092 vdd.n217 gnd 0.009486f
C3093 vdd.n218 gnd 0.007635f
C3094 vdd.n219 gnd 0.009486f
C3095 vdd.n220 gnd 0.009486f
C3096 vdd.n221 gnd 0.007635f
C3097 vdd.n222 gnd 0.009486f
C3098 vdd.n223 gnd 0.009486f
C3099 vdd.n224 gnd 0.007635f
C3100 vdd.n225 gnd 0.009486f
C3101 vdd.n226 gnd 0.009486f
C3102 vdd.n227 gnd 0.007635f
C3103 vdd.n228 gnd 0.009486f
C3104 vdd.n229 gnd 0.007635f
C3105 vdd.n230 gnd 0.009486f
C3106 vdd.n231 gnd 0.007635f
C3107 vdd.n232 gnd 0.009486f
C3108 vdd.n233 gnd 0.009486f
C3109 vdd.n234 gnd 0.761188f
C3110 vdd.t156 gnd 0.380594f
C3111 vdd.n235 gnd 0.009486f
C3112 vdd.n236 gnd 0.007635f
C3113 vdd.n237 gnd 0.009486f
C3114 vdd.n238 gnd 0.007635f
C3115 vdd.n239 gnd 0.009486f
C3116 vdd.t167 gnd 0.380594f
C3117 vdd.n240 gnd 0.009486f
C3118 vdd.n241 gnd 0.007635f
C3119 vdd.n242 gnd 0.009486f
C3120 vdd.n243 gnd 0.007635f
C3121 vdd.n244 gnd 0.009486f
C3122 vdd.n245 gnd 0.437683f
C3123 vdd.n246 gnd 0.574697f
C3124 vdd.n247 gnd 0.009486f
C3125 vdd.n248 gnd 0.007635f
C3126 vdd.n249 gnd 0.009486f
C3127 vdd.n250 gnd 0.007635f
C3128 vdd.n251 gnd 0.009486f
C3129 vdd.n252 gnd 0.688875f
C3130 vdd.n253 gnd 0.009486f
C3131 vdd.n254 gnd 0.007635f
C3132 vdd.n255 gnd 0.009486f
C3133 vdd.n256 gnd 0.007635f
C3134 vdd.n257 gnd 0.009486f
C3135 vdd.n258 gnd 0.761188f
C3136 vdd.t9 gnd 0.380594f
C3137 vdd.n259 gnd 0.009486f
C3138 vdd.n260 gnd 0.007635f
C3139 vdd.n261 gnd 0.009486f
C3140 vdd.n262 gnd 0.007635f
C3141 vdd.n263 gnd 0.009486f
C3142 vdd.t103 gnd 0.380594f
C3143 vdd.n264 gnd 0.009486f
C3144 vdd.n265 gnd 0.007635f
C3145 vdd.n266 gnd 0.009486f
C3146 vdd.n267 gnd 0.007635f
C3147 vdd.n268 gnd 0.009486f
C3148 vdd.n269 gnd 0.761188f
C3149 vdd.n270 gnd 0.582309f
C3150 vdd.n271 gnd 0.009486f
C3151 vdd.n272 gnd 0.007635f
C3152 vdd.n273 gnd 0.009486f
C3153 vdd.n274 gnd 0.007635f
C3154 vdd.n275 gnd 0.009486f
C3155 vdd.n276 gnd 0.498578f
C3156 vdd.n277 gnd 0.009486f
C3157 vdd.n278 gnd 0.007635f
C3158 vdd.n279 gnd 0.021312f
C3159 vdd.n280 gnd 0.006337f
C3160 vdd.n281 gnd 0.021312f
C3161 vdd.n282 gnd 0.978126f
C3162 vdd.t36 gnd 0.380594f
C3163 vdd.n283 gnd 0.021312f
C3164 vdd.n284 gnd 0.006337f
C3165 vdd.n285 gnd 0.009486f
C3166 vdd.n286 gnd 0.007635f
C3167 vdd.n287 gnd 0.009486f
C3168 vdd.n288 gnd 4.45295f
C3169 vdd.n316 gnd 0.021375f
C3170 vdd.n317 gnd 0.009486f
C3171 vdd.n318 gnd 0.009486f
C3172 vdd.n319 gnd 0.009486f
C3173 vdd.n320 gnd 0.008158f
C3174 vdd.n321 gnd 0.007635f
C3175 vdd.n322 gnd 0.006071f
C3176 vdd.n323 gnd 0.008999f
C3177 vdd.n324 gnd 0.009486f
C3178 vdd.n325 gnd 0.009486f
C3179 vdd.n326 gnd 0.007635f
C3180 vdd.n327 gnd 0.009486f
C3181 vdd.n328 gnd 0.009486f
C3182 vdd.n329 gnd 0.009486f
C3183 vdd.n330 gnd 0.009486f
C3184 vdd.n331 gnd 0.009486f
C3185 vdd.n332 gnd 0.009486f
C3186 vdd.n333 gnd 0.009486f
C3187 vdd.n334 gnd 0.009486f
C3188 vdd.n335 gnd 0.006375f
C3189 vdd.n336 gnd 0.009486f
C3190 vdd.n337 gnd 0.009486f
C3191 vdd.n338 gnd 0.009486f
C3192 vdd.n339 gnd 0.009486f
C3193 vdd.n340 gnd 0.009486f
C3194 vdd.n341 gnd 0.009486f
C3195 vdd.n342 gnd 0.009486f
C3196 vdd.n343 gnd 0.009486f
C3197 vdd.n344 gnd 0.009486f
C3198 vdd.n345 gnd 0.009486f
C3199 vdd.n346 gnd 0.009486f
C3200 vdd.n347 gnd 0.009486f
C3201 vdd.n348 gnd 0.009486f
C3202 vdd.n349 gnd 0.009486f
C3203 vdd.n350 gnd 0.009486f
C3204 vdd.n351 gnd 0.009486f
C3205 vdd.n352 gnd 0.009486f
C3206 vdd.n353 gnd 0.007559f
C3207 vdd.t82 gnd 0.194308f
C3208 vdd.t83 gnd 0.203627f
C3209 vdd.t81 gnd 0.283884f
C3210 vdd.n354 gnd 0.096222f
C3211 vdd.n355 gnd 0.055169f
C3212 vdd.n356 gnd 0.009486f
C3213 vdd.n357 gnd 0.009486f
C3214 vdd.n358 gnd 0.009486f
C3215 vdd.n359 gnd 0.009486f
C3216 vdd.n360 gnd 0.009486f
C3217 vdd.n361 gnd 0.009486f
C3218 vdd.n362 gnd 0.009486f
C3219 vdd.n363 gnd 0.009486f
C3220 vdd.n364 gnd 0.006071f
C3221 vdd.n365 gnd 0.007635f
C3222 vdd.n366 gnd 0.008158f
C3223 vdd.n367 gnd 0.004838f
C3224 vdd.n368 gnd 0.00645f
C3225 vdd.n370 gnd 0.00645f
C3226 vdd.n371 gnd 0.00645f
C3227 vdd.n373 gnd 0.00645f
C3228 vdd.n374 gnd 0.00498f
C3229 vdd.n376 gnd 0.00645f
C3230 vdd.t63 gnd 0.082471f
C3231 vdd.t62 gnd 0.093776f
C3232 vdd.t60 gnd 0.246066f
C3233 vdd.n377 gnd 0.164301f
C3234 vdd.n378 gnd 0.132315f
C3235 vdd.n379 gnd 0.009219f
C3236 vdd.n380 gnd 0.015119f
C3237 vdd.n382 gnd 0.00645f
C3238 vdd.n383 gnd 0.517608f
C3239 vdd.n384 gnd 0.014326f
C3240 vdd.n385 gnd 0.014326f
C3241 vdd.n386 gnd 0.00645f
C3242 vdd.n387 gnd 0.015081f
C3243 vdd.n388 gnd 0.00645f
C3244 vdd.n389 gnd 0.00645f
C3245 vdd.n391 gnd 0.00645f
C3246 vdd.n392 gnd 0.00645f
C3247 vdd.n394 gnd 0.00645f
C3248 vdd.n395 gnd 0.00645f
C3249 vdd.n397 gnd 0.00645f
C3250 vdd.n398 gnd 0.00645f
C3251 vdd.n400 gnd 0.00645f
C3252 vdd.n401 gnd 0.00645f
C3253 vdd.n403 gnd 0.00645f
C3254 vdd.t96 gnd 0.082471f
C3255 vdd.t95 gnd 0.093776f
C3256 vdd.t94 gnd 0.246066f
C3257 vdd.n404 gnd 0.164301f
C3258 vdd.n405 gnd 0.132315f
C3259 vdd.n406 gnd 0.00645f
C3260 vdd.n408 gnd 0.00645f
C3261 vdd.n409 gnd 0.00645f
C3262 vdd.n410 gnd 0.285445f
C3263 vdd.n411 gnd 0.00645f
C3264 vdd.n412 gnd 0.00645f
C3265 vdd.n413 gnd 0.00645f
C3266 vdd.n414 gnd 0.00645f
C3267 vdd.n415 gnd 0.00645f
C3268 vdd.n416 gnd 0.433877f
C3269 vdd.n417 gnd 0.00645f
C3270 vdd.n418 gnd 0.00645f
C3271 vdd.t61 gnd 0.258804f
C3272 vdd.n419 gnd 0.00645f
C3273 vdd.n420 gnd 0.00645f
C3274 vdd.t76 gnd 0.093776f
C3275 vdd.t74 gnd 0.246066f
C3276 vdd.t77 gnd 0.093776f
C3277 vdd.n421 gnd 0.297299f
C3278 vdd.n422 gnd 0.00645f
C3279 vdd.n423 gnd 0.00645f
C3280 vdd.n424 gnd 0.517608f
C3281 vdd.n425 gnd 0.00645f
C3282 vdd.n426 gnd 0.00645f
C3283 vdd.t75 gnd 0.258804f
C3284 vdd.n427 gnd 0.00645f
C3285 vdd.n428 gnd 0.00645f
C3286 vdd.n429 gnd 0.00645f
C3287 vdd.n430 gnd 0.517608f
C3288 vdd.n431 gnd 0.00645f
C3289 vdd.n432 gnd 0.00645f
C3290 vdd.n433 gnd 0.00645f
C3291 vdd.n434 gnd 0.00645f
C3292 vdd.n435 gnd 0.00645f
C3293 vdd.t0 gnd 0.258804f
C3294 vdd.n436 gnd 0.00645f
C3295 vdd.n437 gnd 0.00645f
C3296 vdd.n438 gnd 0.00645f
C3297 vdd.n439 gnd 0.00645f
C3298 vdd.n440 gnd 0.00645f
C3299 vdd.t124 gnd 0.258804f
C3300 vdd.n441 gnd 0.00645f
C3301 vdd.n442 gnd 0.00645f
C3302 vdd.n443 gnd 0.460519f
C3303 vdd.n444 gnd 0.00645f
C3304 vdd.n445 gnd 0.00645f
C3305 vdd.n446 gnd 0.00645f
C3306 vdd.t155 gnd 0.258804f
C3307 vdd.n447 gnd 0.00645f
C3308 vdd.n448 gnd 0.00645f
C3309 vdd.n449 gnd 0.312087f
C3310 vdd.n450 gnd 0.00645f
C3311 vdd.n451 gnd 0.00645f
C3312 vdd.n452 gnd 0.00645f
C3313 vdd.t140 gnd 0.258804f
C3314 vdd.n453 gnd 0.00645f
C3315 vdd.n454 gnd 0.00645f
C3316 vdd.n455 gnd 0.483354f
C3317 vdd.n456 gnd 0.00645f
C3318 vdd.n457 gnd 0.00645f
C3319 vdd.n458 gnd 0.00645f
C3320 vdd.t21 gnd 0.258804f
C3321 vdd.n459 gnd 0.00645f
C3322 vdd.n460 gnd 0.00645f
C3323 vdd.n461 gnd 0.334923f
C3324 vdd.n462 gnd 0.00645f
C3325 vdd.n463 gnd 0.00645f
C3326 vdd.n464 gnd 0.00645f
C3327 vdd.t177 gnd 0.258804f
C3328 vdd.n465 gnd 0.00645f
C3329 vdd.n466 gnd 0.00645f
C3330 vdd.n467 gnd 0.50619f
C3331 vdd.n468 gnd 0.00645f
C3332 vdd.n469 gnd 0.00645f
C3333 vdd.n470 gnd 0.00645f
C3334 vdd.n471 gnd 0.517608f
C3335 vdd.n472 gnd 0.00645f
C3336 vdd.n473 gnd 0.00645f
C3337 vdd.t137 gnd 0.258804f
C3338 vdd.n474 gnd 0.00645f
C3339 vdd.n475 gnd 0.00645f
C3340 vdd.n476 gnd 0.00645f
C3341 vdd.t179 gnd 0.258804f
C3342 vdd.n477 gnd 0.00645f
C3343 vdd.n478 gnd 0.00645f
C3344 vdd.n479 gnd 0.00645f
C3345 vdd.n480 gnd 0.00645f
C3346 vdd.n481 gnd 0.00645f
C3347 vdd.n482 gnd 0.517608f
C3348 vdd.n483 gnd 0.00645f
C3349 vdd.n484 gnd 0.00645f
C3350 vdd.t176 gnd 0.258804f
C3351 vdd.n485 gnd 0.00645f
C3352 vdd.n486 gnd 0.00645f
C3353 vdd.n487 gnd 0.00645f
C3354 vdd.n488 gnd 0.460519f
C3355 vdd.n489 gnd 0.00645f
C3356 vdd.n490 gnd 0.00645f
C3357 vdd.n491 gnd 0.00645f
C3358 vdd.n492 gnd 0.00645f
C3359 vdd.n493 gnd 0.00645f
C3360 vdd.t145 gnd 0.258804f
C3361 vdd.n494 gnd 0.00645f
C3362 vdd.n495 gnd 0.00645f
C3363 vdd.t113 gnd 0.258804f
C3364 vdd.n496 gnd 0.00645f
C3365 vdd.n497 gnd 0.00645f
C3366 vdd.n498 gnd 0.00645f
C3367 vdd.n499 gnd 0.517608f
C3368 vdd.n500 gnd 0.00645f
C3369 vdd.n501 gnd 0.00645f
C3370 vdd.n502 gnd 0.372982f
C3371 vdd.n503 gnd 0.00645f
C3372 vdd.n504 gnd 0.00645f
C3373 vdd.n505 gnd 0.00645f
C3374 vdd.t1 gnd 0.258804f
C3375 vdd.n506 gnd 0.00645f
C3376 vdd.n507 gnd 0.00645f
C3377 vdd.n508 gnd 0.00645f
C3378 vdd.n509 gnd 0.00645f
C3379 vdd.n510 gnd 0.00645f
C3380 vdd.t47 gnd 0.258804f
C3381 vdd.n511 gnd 0.00645f
C3382 vdd.n512 gnd 0.00645f
C3383 vdd.n513 gnd 0.395818f
C3384 vdd.n514 gnd 0.00645f
C3385 vdd.n515 gnd 0.00645f
C3386 vdd.n516 gnd 0.00645f
C3387 vdd.t214 gnd 0.258804f
C3388 vdd.n517 gnd 0.00645f
C3389 vdd.n518 gnd 0.00645f
C3390 vdd.n519 gnd 0.285445f
C3391 vdd.n520 gnd 0.00645f
C3392 vdd.n521 gnd 0.015081f
C3393 vdd.n522 gnd 0.015081f
C3394 vdd.n523 gnd 0.715516f
C3395 vdd.n549 gnd 0.015081f
C3396 vdd.n550 gnd 0.014326f
C3397 vdd.n551 gnd 0.00645f
C3398 vdd.n552 gnd 0.014326f
C3399 vdd.t80 gnd 0.082471f
C3400 vdd.t79 gnd 0.093776f
C3401 vdd.t78 gnd 0.246066f
C3402 vdd.n553 gnd 0.164301f
C3403 vdd.n554 gnd 0.132315f
C3404 vdd.n555 gnd 0.009219f
C3405 vdd.n556 gnd 0.00645f
C3406 vdd.n557 gnd 0.00645f
C3407 vdd.t181 gnd 0.258804f
C3408 vdd.n558 gnd 0.00645f
C3409 vdd.n559 gnd 0.00645f
C3410 vdd.n560 gnd 0.00645f
C3411 vdd.n561 gnd 0.014326f
C3412 vdd.n562 gnd 0.00645f
C3413 vdd.t56 gnd 0.082471f
C3414 vdd.t55 gnd 0.093776f
C3415 vdd.t53 gnd 0.246066f
C3416 vdd.n563 gnd 0.164301f
C3417 vdd.n564 gnd 0.132315f
C3418 vdd.n565 gnd 0.00645f
C3419 vdd.n566 gnd 0.00645f
C3420 vdd.n567 gnd 0.285445f
C3421 vdd.n568 gnd 0.00645f
C3422 vdd.n569 gnd 0.00645f
C3423 vdd.n570 gnd 0.00645f
C3424 vdd.n571 gnd 0.395818f
C3425 vdd.n572 gnd 0.00645f
C3426 vdd.n573 gnd 0.00645f
C3427 vdd.t54 gnd 0.258804f
C3428 vdd.n574 gnd 0.00645f
C3429 vdd.n575 gnd 0.00645f
C3430 vdd.n576 gnd 0.00645f
C3431 vdd.n577 gnd 0.00645f
C3432 vdd.n578 gnd 0.517608f
C3433 vdd.n579 gnd 0.00645f
C3434 vdd.n580 gnd 0.00645f
C3435 vdd.t122 gnd 0.258804f
C3436 vdd.n581 gnd 0.00645f
C3437 vdd.n582 gnd 0.00645f
C3438 vdd.n583 gnd 0.00645f
C3439 vdd.n584 gnd 0.372982f
C3440 vdd.n585 gnd 0.00645f
C3441 vdd.n586 gnd 0.00645f
C3442 vdd.n587 gnd 0.00645f
C3443 vdd.n588 gnd 0.00645f
C3444 vdd.n589 gnd 0.00645f
C3445 vdd.t173 gnd 0.258804f
C3446 vdd.n590 gnd 0.00645f
C3447 vdd.n591 gnd 0.00645f
C3448 vdd.t138 gnd 0.258804f
C3449 vdd.n592 gnd 0.00645f
C3450 vdd.n593 gnd 0.00645f
C3451 vdd.n594 gnd 0.00645f
C3452 vdd.n595 gnd 0.517608f
C3453 vdd.n596 gnd 0.00645f
C3454 vdd.n597 gnd 0.00645f
C3455 vdd.n598 gnd 0.460519f
C3456 vdd.n599 gnd 0.00645f
C3457 vdd.n600 gnd 0.00645f
C3458 vdd.n601 gnd 0.00645f
C3459 vdd.t22 gnd 0.258804f
C3460 vdd.n602 gnd 0.00645f
C3461 vdd.n603 gnd 0.00645f
C3462 vdd.n604 gnd 0.00645f
C3463 vdd.n605 gnd 0.00645f
C3464 vdd.n606 gnd 0.00645f
C3465 vdd.n607 gnd 0.517608f
C3466 vdd.n608 gnd 0.00645f
C3467 vdd.n609 gnd 0.00645f
C3468 vdd.t201 gnd 0.258804f
C3469 vdd.n610 gnd 0.00645f
C3470 vdd.n611 gnd 0.00645f
C3471 vdd.n612 gnd 0.00645f
C3472 vdd.t144 gnd 0.258804f
C3473 vdd.n613 gnd 0.00645f
C3474 vdd.n614 gnd 0.00645f
C3475 vdd.n615 gnd 0.00645f
C3476 vdd.n616 gnd 0.00645f
C3477 vdd.n617 gnd 0.00645f
C3478 vdd.n618 gnd 0.50619f
C3479 vdd.n619 gnd 0.00645f
C3480 vdd.n620 gnd 0.00645f
C3481 vdd.t142 gnd 0.258804f
C3482 vdd.n621 gnd 0.00645f
C3483 vdd.n622 gnd 0.00645f
C3484 vdd.n623 gnd 0.00645f
C3485 vdd.n624 gnd 0.334923f
C3486 vdd.n625 gnd 0.00645f
C3487 vdd.n626 gnd 0.00645f
C3488 vdd.t172 gnd 0.258804f
C3489 vdd.n627 gnd 0.00645f
C3490 vdd.n628 gnd 0.00645f
C3491 vdd.n629 gnd 0.00645f
C3492 vdd.n630 gnd 0.483354f
C3493 vdd.n631 gnd 0.00645f
C3494 vdd.n632 gnd 0.00645f
C3495 vdd.t194 gnd 0.258804f
C3496 vdd.n633 gnd 0.00645f
C3497 vdd.n634 gnd 0.00645f
C3498 vdd.n635 gnd 0.00645f
C3499 vdd.n636 gnd 0.312087f
C3500 vdd.n637 gnd 0.00645f
C3501 vdd.n638 gnd 0.00645f
C3502 vdd.t154 gnd 0.258804f
C3503 vdd.n639 gnd 0.00645f
C3504 vdd.n640 gnd 0.00645f
C3505 vdd.n641 gnd 0.00645f
C3506 vdd.n642 gnd 0.460519f
C3507 vdd.n643 gnd 0.00645f
C3508 vdd.n644 gnd 0.00645f
C3509 vdd.t135 gnd 0.258804f
C3510 vdd.n645 gnd 0.00645f
C3511 vdd.n646 gnd 0.00645f
C3512 vdd.n647 gnd 0.00645f
C3513 vdd.n648 gnd 0.517608f
C3514 vdd.n649 gnd 0.00645f
C3515 vdd.n650 gnd 0.00645f
C3516 vdd.t3 gnd 0.258804f
C3517 vdd.n651 gnd 0.00645f
C3518 vdd.n652 gnd 0.00645f
C3519 vdd.n653 gnd 0.00645f
C3520 vdd.n654 gnd 0.517608f
C3521 vdd.n655 gnd 0.00645f
C3522 vdd.n656 gnd 0.00645f
C3523 vdd.n657 gnd 0.00645f
C3524 vdd.n658 gnd 0.00645f
C3525 vdd.n659 gnd 0.00645f
C3526 vdd.t91 gnd 0.258804f
C3527 vdd.n660 gnd 0.00645f
C3528 vdd.n661 gnd 0.00645f
C3529 vdd.n662 gnd 0.00645f
C3530 vdd.t92 gnd 0.093776f
C3531 vdd.t90 gnd 0.246066f
C3532 vdd.t93 gnd 0.093776f
C3533 vdd.n663 gnd 0.297299f
C3534 vdd.n664 gnd 0.00645f
C3535 vdd.n665 gnd 0.00645f
C3536 vdd.t32 gnd 0.258804f
C3537 vdd.n666 gnd 0.00645f
C3538 vdd.n667 gnd 0.00645f
C3539 vdd.n668 gnd 0.433877f
C3540 vdd.n669 gnd 0.00645f
C3541 vdd.n670 gnd 0.00645f
C3542 vdd.n671 gnd 0.00645f
C3543 vdd.n672 gnd 0.517608f
C3544 vdd.n673 gnd 0.00645f
C3545 vdd.n674 gnd 0.00645f
C3546 vdd.n675 gnd 0.285445f
C3547 vdd.n676 gnd 0.00645f
C3548 vdd.n677 gnd 0.015081f
C3549 vdd.n678 gnd 0.015081f
C3550 vdd.n679 gnd 4.45295f
C3551 vdd.n680 gnd 0.014326f
C3552 vdd.n681 gnd 0.014326f
C3553 vdd.n682 gnd 0.015081f
C3554 vdd.n683 gnd 0.00645f
C3555 vdd.n685 gnd 0.00645f
C3556 vdd.n686 gnd 0.00645f
C3557 vdd.n687 gnd 0.00645f
C3558 vdd.n688 gnd 0.00645f
C3559 vdd.n689 gnd 0.012762f
C3560 vdd.n691 gnd 0.00645f
C3561 vdd.n692 gnd 0.00645f
C3562 vdd.n693 gnd 0.00645f
C3563 vdd.n694 gnd 0.00645f
C3564 vdd.t33 gnd 0.082471f
C3565 vdd.t34 gnd 0.093776f
C3566 vdd.t31 gnd 0.246066f
C3567 vdd.n695 gnd 0.164301f
C3568 vdd.n696 gnd 0.132315f
C3569 vdd.n697 gnd 0.009219f
C3570 vdd.n699 gnd 0.00645f
C3571 vdd.n700 gnd 0.00645f
C3572 vdd.n701 gnd 0.00645f
C3573 vdd.t65 gnd 0.082471f
C3574 vdd.t66 gnd 0.093776f
C3575 vdd.t64 gnd 0.246066f
C3576 vdd.n702 gnd 0.164301f
C3577 vdd.n703 gnd 0.132315f
C3578 vdd.n704 gnd 0.00645f
C3579 vdd.n705 gnd 0.00645f
C3580 vdd.n706 gnd 0.00645f
C3581 vdd.n707 gnd 0.00645f
C3582 vdd.n708 gnd 0.006071f
C3583 vdd.n711 gnd 0.009486f
C3584 vdd.n712 gnd 0.007635f
C3585 vdd.n713 gnd 0.009486f
C3586 vdd.n714 gnd 0.009486f
C3587 vdd.n715 gnd 0.009486f
C3588 vdd.n716 gnd 0.004008f
C3589 vdd.n717 gnd 0.021312f
C3590 vdd.t89 gnd 0.194308f
C3591 vdd.t88 gnd 0.203627f
C3592 vdd.t87 gnd 0.283884f
C3593 vdd.n718 gnd 0.096222f
C3594 vdd.n719 gnd 0.055169f
C3595 vdd.n720 gnd 0.011796f
C3596 vdd.n721 gnd 0.009486f
C3597 vdd.n723 gnd 0.009486f
C3598 vdd.n724 gnd 0.006337f
C3599 vdd.n725 gnd 0.643204f
C3600 vdd.n727 gnd 4.59377f
C3601 vdd.n728 gnd 0.009486f
C3602 vdd.n729 gnd 0.021375f
C3603 vdd.n730 gnd 0.007635f
C3604 vdd.n731 gnd 0.009486f
C3605 vdd.n732 gnd 0.007635f
C3606 vdd.n733 gnd 0.009486f
C3607 vdd.n734 gnd 0.761188f
C3608 vdd.n735 gnd 0.009486f
C3609 vdd.n736 gnd 0.007635f
C3610 vdd.n737 gnd 0.007635f
C3611 vdd.n738 gnd 0.009486f
C3612 vdd.n739 gnd 0.007635f
C3613 vdd.n740 gnd 0.009486f
C3614 vdd.n741 gnd 0.761188f
C3615 vdd.n742 gnd 0.009486f
C3616 vdd.n743 gnd 0.007635f
C3617 vdd.n744 gnd 0.009486f
C3618 vdd.n745 gnd 0.007635f
C3619 vdd.n746 gnd 0.009486f
C3620 vdd.t118 gnd 0.380594f
C3621 vdd.n747 gnd 0.009486f
C3622 vdd.n748 gnd 0.007635f
C3623 vdd.n749 gnd 0.009486f
C3624 vdd.n750 gnd 0.007635f
C3625 vdd.n751 gnd 0.009486f
C3626 vdd.n752 gnd 0.452907f
C3627 vdd.n753 gnd 0.559473f
C3628 vdd.n754 gnd 0.009486f
C3629 vdd.n755 gnd 0.007635f
C3630 vdd.n756 gnd 0.009486f
C3631 vdd.n757 gnd 0.007635f
C3632 vdd.n758 gnd 0.009486f
C3633 vdd.n759 gnd 0.704099f
C3634 vdd.n760 gnd 0.009486f
C3635 vdd.n761 gnd 0.007635f
C3636 vdd.n762 gnd 0.009486f
C3637 vdd.n763 gnd 0.007635f
C3638 vdd.n764 gnd 0.009486f
C3639 vdd.n765 gnd 0.761188f
C3640 vdd.t110 gnd 0.380594f
C3641 vdd.n766 gnd 0.009486f
C3642 vdd.n767 gnd 0.007635f
C3643 vdd.n768 gnd 0.009486f
C3644 vdd.n769 gnd 0.007635f
C3645 vdd.n770 gnd 0.009486f
C3646 vdd.t133 gnd 0.380594f
C3647 vdd.n771 gnd 0.009486f
C3648 vdd.n772 gnd 0.007635f
C3649 vdd.n773 gnd 0.009486f
C3650 vdd.n774 gnd 0.007635f
C3651 vdd.n775 gnd 0.009486f
C3652 vdd.n776 gnd 0.445295f
C3653 vdd.n777 gnd 0.567085f
C3654 vdd.n778 gnd 0.009486f
C3655 vdd.n779 gnd 0.007635f
C3656 vdd.t119 gnd 0.232594f
C3657 vdd.t111 gnd 0.026723f
C3658 vdd.t192 gnd 0.026723f
C3659 vdd.n780 gnd 0.171507f
C3660 vdd.n781 gnd 0.304174f
C3661 vdd.t158 gnd 0.026723f
C3662 vdd.t171 gnd 0.026723f
C3663 vdd.n782 gnd 0.171507f
C3664 vdd.n783 gnd 0.162092f
C3665 vdd.t132 gnd 0.026723f
C3666 vdd.t20 gnd 0.026723f
C3667 vdd.n784 gnd 0.171507f
C3668 vdd.n785 gnd 0.162092f
C3669 vdd.t193 gnd 0.026723f
C3670 vdd.t131 gnd 0.026723f
C3671 vdd.n786 gnd 0.171507f
C3672 vdd.n787 gnd 0.162092f
C3673 vdd.t112 gnd 0.23156f
C3674 vdd.n788 gnd 0.204642f
C3675 vdd.t199 gnd 0.232594f
C3676 vdd.t184 gnd 0.026723f
C3677 vdd.t117 gnd 0.026723f
C3678 vdd.n789 gnd 0.171507f
C3679 vdd.n790 gnd 0.304174f
C3680 vdd.t121 gnd 0.026723f
C3681 vdd.t134 gnd 0.026723f
C3682 vdd.n791 gnd 0.171507f
C3683 vdd.n792 gnd 0.162092f
C3684 vdd.t115 gnd 0.026723f
C3685 vdd.t169 gnd 0.026723f
C3686 vdd.n793 gnd 0.171507f
C3687 vdd.n794 gnd 0.162092f
C3688 vdd.t187 gnd 0.026723f
C3689 vdd.t213 gnd 0.026723f
C3690 vdd.n795 gnd 0.171507f
C3691 vdd.n796 gnd 0.162092f
C3692 vdd.t153 gnd 0.23156f
C3693 vdd.n797 gnd 0.169939f
C3694 vdd.n798 gnd 0.194956f
C3695 vdd.t163 gnd 0.232594f
C3696 vdd.t185 gnd 0.026723f
C3697 vdd.t204 gnd 0.026723f
C3698 vdd.n799 gnd 0.171507f
C3699 vdd.n800 gnd 0.304174f
C3700 vdd.t150 gnd 0.026723f
C3701 vdd.t188 gnd 0.026723f
C3702 vdd.n801 gnd 0.171507f
C3703 vdd.n802 gnd 0.162092f
C3704 vdd.t189 gnd 0.026723f
C3705 vdd.t105 gnd 0.026723f
C3706 vdd.n803 gnd 0.171507f
C3707 vdd.n804 gnd 0.162092f
C3708 vdd.t205 gnd 0.026723f
C3709 vdd.t130 gnd 0.026723f
C3710 vdd.n805 gnd 0.171507f
C3711 vdd.n806 gnd 0.162092f
C3712 vdd.t15 gnd 0.23156f
C3713 vdd.n807 gnd 0.169939f
C3714 vdd.n808 gnd 0.213388f
C3715 vdd.n809 gnd 1.97048f
C3716 vdd.n810 gnd 0.2589f
C3717 vdd.n811 gnd 0.007635f
C3718 vdd.n812 gnd 0.009486f
C3719 vdd.n813 gnd 0.696487f
C3720 vdd.n814 gnd 0.009486f
C3721 vdd.n815 gnd 0.007635f
C3722 vdd.n816 gnd 0.009486f
C3723 vdd.n817 gnd 0.007635f
C3724 vdd.n818 gnd 0.009486f
C3725 vdd.n819 gnd 0.761188f
C3726 vdd.t19 gnd 0.380594f
C3727 vdd.n820 gnd 0.009486f
C3728 vdd.n821 gnd 0.007635f
C3729 vdd.n822 gnd 0.009486f
C3730 vdd.n823 gnd 0.007635f
C3731 vdd.n824 gnd 0.009486f
C3732 vdd.t114 gnd 0.380594f
C3733 vdd.n825 gnd 0.009486f
C3734 vdd.n826 gnd 0.007635f
C3735 vdd.n827 gnd 0.009486f
C3736 vdd.n828 gnd 0.007635f
C3737 vdd.n829 gnd 0.009486f
C3738 vdd.n830 gnd 0.437683f
C3739 vdd.n831 gnd 0.574697f
C3740 vdd.n832 gnd 0.009486f
C3741 vdd.n833 gnd 0.007635f
C3742 vdd.n834 gnd 0.009486f
C3743 vdd.n835 gnd 0.007635f
C3744 vdd.n836 gnd 0.009486f
C3745 vdd.n837 gnd 0.688875f
C3746 vdd.n838 gnd 0.009486f
C3747 vdd.n839 gnd 0.007635f
C3748 vdd.n840 gnd 0.009486f
C3749 vdd.n841 gnd 0.007635f
C3750 vdd.n842 gnd 0.009486f
C3751 vdd.n843 gnd 0.761188f
C3752 vdd.t186 gnd 0.380594f
C3753 vdd.n844 gnd 0.009486f
C3754 vdd.n845 gnd 0.007635f
C3755 vdd.n846 gnd 0.009486f
C3756 vdd.n847 gnd 0.007635f
C3757 vdd.n848 gnd 0.009486f
C3758 vdd.t14 gnd 0.380594f
C3759 vdd.n849 gnd 0.009486f
C3760 vdd.n850 gnd 0.007635f
C3761 vdd.n851 gnd 0.009486f
C3762 vdd.n852 gnd 0.007635f
C3763 vdd.n853 gnd 0.009486f
C3764 vdd.n854 gnd 0.761188f
C3765 vdd.n855 gnd 0.582309f
C3766 vdd.n856 gnd 0.009486f
C3767 vdd.n857 gnd 0.007635f
C3768 vdd.n858 gnd 0.009486f
C3769 vdd.n859 gnd 0.007635f
C3770 vdd.n860 gnd 0.009486f
C3771 vdd.n861 gnd 0.498578f
C3772 vdd.n862 gnd 0.009486f
C3773 vdd.n863 gnd 0.007635f
C3774 vdd.n864 gnd 0.021312f
C3775 vdd.n865 gnd 0.006337f
C3776 vdd.n866 gnd 0.021312f
C3777 vdd.n867 gnd 0.978126f
C3778 vdd.t43 gnd 0.380594f
C3779 vdd.n868 gnd 0.021312f
C3780 vdd.n869 gnd 0.006337f
C3781 vdd.n870 gnd 0.009486f
C3782 vdd.n871 gnd 0.007635f
C3783 vdd.n872 gnd 0.009486f
C3784 vdd.n900 gnd 0.021375f
C3785 vdd.n901 gnd 0.009486f
C3786 vdd.n902 gnd 0.007635f
C3787 vdd.n903 gnd 0.009486f
C3788 vdd.n904 gnd 0.009486f
C3789 vdd.n905 gnd 0.009486f
C3790 vdd.n906 gnd 0.009486f
C3791 vdd.n907 gnd 0.009486f
C3792 vdd.n908 gnd 0.007635f
C3793 vdd.n909 gnd 0.009486f
C3794 vdd.n910 gnd 0.009486f
C3795 vdd.n911 gnd 0.009486f
C3796 vdd.n912 gnd 0.009486f
C3797 vdd.n913 gnd 0.009486f
C3798 vdd.n914 gnd 0.007635f
C3799 vdd.n915 gnd 0.009486f
C3800 vdd.n916 gnd 0.009486f
C3801 vdd.n917 gnd 0.009486f
C3802 vdd.n918 gnd 0.009486f
C3803 vdd.n919 gnd 0.009486f
C3804 vdd.n920 gnd 0.007635f
C3805 vdd.n921 gnd 0.009486f
C3806 vdd.n922 gnd 0.009486f
C3807 vdd.n923 gnd 0.009486f
C3808 vdd.n924 gnd 0.009486f
C3809 vdd.n925 gnd 0.007635f
C3810 vdd.n926 gnd 0.009486f
C3811 vdd.n927 gnd 0.009486f
C3812 vdd.n928 gnd 0.009486f
C3813 vdd.n929 gnd 0.009486f
C3814 vdd.n930 gnd 0.009486f
C3815 vdd.n931 gnd 0.007635f
C3816 vdd.n932 gnd 0.009486f
C3817 vdd.n933 gnd 0.009486f
C3818 vdd.n934 gnd 0.009486f
C3819 vdd.n935 gnd 0.009486f
C3820 vdd.n936 gnd 0.009486f
C3821 vdd.n937 gnd 0.007635f
C3822 vdd.n938 gnd 0.009486f
C3823 vdd.n939 gnd 0.009486f
C3824 vdd.n940 gnd 0.009486f
C3825 vdd.n941 gnd 0.009486f
C3826 vdd.n942 gnd 0.009486f
C3827 vdd.n943 gnd 0.007635f
C3828 vdd.n944 gnd 0.009486f
C3829 vdd.n945 gnd 0.009486f
C3830 vdd.n946 gnd 0.009486f
C3831 vdd.n947 gnd 0.009486f
C3832 vdd.n948 gnd 0.009486f
C3833 vdd.n949 gnd 0.007635f
C3834 vdd.n950 gnd 0.009486f
C3835 vdd.n951 gnd 0.009486f
C3836 vdd.n952 gnd 0.009486f
C3837 vdd.n953 gnd 0.009486f
C3838 vdd.n954 gnd 0.007635f
C3839 vdd.n955 gnd 0.009486f
C3840 vdd.n956 gnd 0.009486f
C3841 vdd.n957 gnd 0.009486f
C3842 vdd.n958 gnd 0.009486f
C3843 vdd.n959 gnd 0.009486f
C3844 vdd.n960 gnd 0.007635f
C3845 vdd.n961 gnd 0.009486f
C3846 vdd.n962 gnd 0.009486f
C3847 vdd.n963 gnd 0.009486f
C3848 vdd.n964 gnd 0.009486f
C3849 vdd.n965 gnd 0.009486f
C3850 vdd.n966 gnd 0.007635f
C3851 vdd.n967 gnd 0.009486f
C3852 vdd.n968 gnd 0.009486f
C3853 vdd.n969 gnd 0.009486f
C3854 vdd.n970 gnd 0.009486f
C3855 vdd.n971 gnd 0.009486f
C3856 vdd.n972 gnd 0.007635f
C3857 vdd.n973 gnd 0.009486f
C3858 vdd.n974 gnd 0.009486f
C3859 vdd.n975 gnd 0.009486f
C3860 vdd.n976 gnd 0.009486f
C3861 vdd.n977 gnd 0.009486f
C3862 vdd.n978 gnd 0.007635f
C3863 vdd.n979 gnd 0.021375f
C3864 vdd.n980 gnd 0.009486f
C3865 vdd.n981 gnd 0.003627f
C3866 vdd.t44 gnd 0.194308f
C3867 vdd.t45 gnd 0.203627f
C3868 vdd.t42 gnd 0.283884f
C3869 vdd.n982 gnd 0.096222f
C3870 vdd.n983 gnd 0.055169f
C3871 vdd.n984 gnd 0.011796f
C3872 vdd.n985 gnd 0.004008f
C3873 vdd.n986 gnd 0.009486f
C3874 vdd.n987 gnd 0.009486f
C3875 vdd.n988 gnd 0.009486f
C3876 vdd.n989 gnd 0.007635f
C3877 vdd.n990 gnd 0.007635f
C3878 vdd.n991 gnd 0.007635f
C3879 vdd.n992 gnd 0.009486f
C3880 vdd.n993 gnd 0.009486f
C3881 vdd.n994 gnd 0.009486f
C3882 vdd.n995 gnd 0.007635f
C3883 vdd.n996 gnd 0.007635f
C3884 vdd.n997 gnd 0.007635f
C3885 vdd.n998 gnd 0.009486f
C3886 vdd.n999 gnd 0.009486f
C3887 vdd.n1000 gnd 0.009486f
C3888 vdd.n1001 gnd 0.007635f
C3889 vdd.n1002 gnd 0.007635f
C3890 vdd.n1003 gnd 0.007635f
C3891 vdd.n1004 gnd 0.009486f
C3892 vdd.n1005 gnd 0.009486f
C3893 vdd.n1006 gnd 0.009486f
C3894 vdd.n1007 gnd 0.007635f
C3895 vdd.n1008 gnd 0.007635f
C3896 vdd.n1009 gnd 0.007635f
C3897 vdd.n1010 gnd 0.009486f
C3898 vdd.n1011 gnd 0.009486f
C3899 vdd.n1012 gnd 0.009486f
C3900 vdd.n1013 gnd 0.007559f
C3901 vdd.n1014 gnd 0.009486f
C3902 vdd.t58 gnd 0.194308f
C3903 vdd.t59 gnd 0.203627f
C3904 vdd.t57 gnd 0.283884f
C3905 vdd.n1015 gnd 0.096222f
C3906 vdd.n1016 gnd 0.055169f
C3907 vdd.n1017 gnd 0.015614f
C3908 vdd.n1018 gnd 0.005192f
C3909 vdd.n1019 gnd 0.009486f
C3910 vdd.n1020 gnd 0.009486f
C3911 vdd.n1021 gnd 0.009486f
C3912 vdd.n1022 gnd 0.007635f
C3913 vdd.n1023 gnd 0.007635f
C3914 vdd.n1024 gnd 0.007635f
C3915 vdd.n1025 gnd 0.009486f
C3916 vdd.n1026 gnd 0.009486f
C3917 vdd.n1027 gnd 0.009486f
C3918 vdd.n1028 gnd 0.007635f
C3919 vdd.n1029 gnd 0.007635f
C3920 vdd.n1030 gnd 0.007635f
C3921 vdd.n1031 gnd 0.009486f
C3922 vdd.n1032 gnd 0.009486f
C3923 vdd.n1033 gnd 0.009486f
C3924 vdd.n1034 gnd 0.007635f
C3925 vdd.n1035 gnd 0.007635f
C3926 vdd.n1036 gnd 0.007635f
C3927 vdd.n1037 gnd 0.009486f
C3928 vdd.n1038 gnd 0.009486f
C3929 vdd.n1039 gnd 0.009486f
C3930 vdd.n1040 gnd 0.007635f
C3931 vdd.n1041 gnd 0.007635f
C3932 vdd.n1042 gnd 0.007635f
C3933 vdd.n1043 gnd 0.009486f
C3934 vdd.n1044 gnd 0.009486f
C3935 vdd.n1045 gnd 0.009486f
C3936 vdd.n1046 gnd 0.006375f
C3937 vdd.n1047 gnd 0.009486f
C3938 vdd.t85 gnd 0.194308f
C3939 vdd.t86 gnd 0.203627f
C3940 vdd.t84 gnd 0.283884f
C3941 vdd.n1048 gnd 0.096222f
C3942 vdd.n1049 gnd 0.055169f
C3943 vdd.n1050 gnd 0.015614f
C3944 vdd.n1051 gnd 0.006375f
C3945 vdd.n1052 gnd 0.009486f
C3946 vdd.n1053 gnd 0.009486f
C3947 vdd.n1054 gnd 0.009486f
C3948 vdd.n1055 gnd 0.007635f
C3949 vdd.n1056 gnd 0.007635f
C3950 vdd.n1057 gnd 0.007635f
C3951 vdd.n1058 gnd 0.009486f
C3952 vdd.n1059 gnd 0.009486f
C3953 vdd.n1060 gnd 0.009486f
C3954 vdd.n1061 gnd 0.007635f
C3955 vdd.n1062 gnd 0.007635f
C3956 vdd.n1063 gnd 0.007635f
C3957 vdd.n1064 gnd 0.009486f
C3958 vdd.n1065 gnd 0.009486f
C3959 vdd.n1066 gnd 0.009486f
C3960 vdd.n1067 gnd 0.007635f
C3961 vdd.n1068 gnd 0.007635f
C3962 vdd.n1069 gnd 0.007635f
C3963 vdd.n1070 gnd 0.009486f
C3964 vdd.n1071 gnd 0.009486f
C3965 vdd.n1072 gnd 0.009486f
C3966 vdd.n1073 gnd 0.007635f
C3967 vdd.n1074 gnd 0.009486f
C3968 vdd.n1075 gnd 1.65558f
C3969 vdd.n1077 gnd 0.021375f
C3970 vdd.n1078 gnd 0.006337f
C3971 vdd.n1079 gnd 0.021375f
C3972 vdd.n1080 gnd 0.021312f
C3973 vdd.n1081 gnd 0.009486f
C3974 vdd.n1082 gnd 0.007635f
C3975 vdd.n1083 gnd 0.009486f
C3976 vdd.n1084 gnd 0.643204f
C3977 vdd.n1085 gnd 0.009486f
C3978 vdd.n1086 gnd 0.007635f
C3979 vdd.n1087 gnd 0.009486f
C3980 vdd.n1088 gnd 0.009486f
C3981 vdd.n1089 gnd 0.009486f
C3982 vdd.n1090 gnd 0.007635f
C3983 vdd.n1091 gnd 0.009486f
C3984 vdd.n1092 gnd 0.761188f
C3985 vdd.n1093 gnd 0.009486f
C3986 vdd.n1094 gnd 0.007635f
C3987 vdd.n1095 gnd 0.009486f
C3988 vdd.n1096 gnd 0.009486f
C3989 vdd.n1097 gnd 0.009486f
C3990 vdd.n1098 gnd 0.007635f
C3991 vdd.n1099 gnd 0.009486f
C3992 vdd.n1100 gnd 0.761188f
C3993 vdd.n1101 gnd 0.009486f
C3994 vdd.n1102 gnd 0.007635f
C3995 vdd.n1103 gnd 0.009486f
C3996 vdd.n1104 gnd 0.009486f
C3997 vdd.n1105 gnd 0.009486f
C3998 vdd.n1106 gnd 0.007635f
C3999 vdd.n1107 gnd 0.009486f
C4000 vdd.n1108 gnd 0.559473f
C4001 vdd.n1109 gnd 0.009486f
C4002 vdd.n1110 gnd 0.007635f
C4003 vdd.n1111 gnd 0.009486f
C4004 vdd.n1112 gnd 0.009486f
C4005 vdd.n1113 gnd 0.009486f
C4006 vdd.n1114 gnd 0.007635f
C4007 vdd.n1115 gnd 0.009486f
C4008 vdd.n1116 gnd 0.452907f
C4009 vdd.n1117 gnd 0.009486f
C4010 vdd.n1118 gnd 0.007635f
C4011 vdd.n1119 gnd 0.009486f
C4012 vdd.n1120 gnd 0.009486f
C4013 vdd.n1121 gnd 0.009486f
C4014 vdd.n1122 gnd 0.007635f
C4015 vdd.n1123 gnd 0.009486f
C4016 vdd.t129 gnd 0.380594f
C4017 vdd.n1124 gnd 0.704099f
C4018 vdd.n1125 gnd 0.009486f
C4019 vdd.n1126 gnd 0.007635f
C4020 vdd.n1127 gnd 0.009486f
C4021 vdd.n1128 gnd 0.009486f
C4022 vdd.n1129 gnd 0.009486f
C4023 vdd.n1130 gnd 0.007635f
C4024 vdd.n1131 gnd 0.009486f
C4025 vdd.n1132 gnd 0.761188f
C4026 vdd.n1133 gnd 0.009486f
C4027 vdd.n1134 gnd 0.007635f
C4028 vdd.n1135 gnd 0.009486f
C4029 vdd.n1136 gnd 0.009486f
C4030 vdd.n1137 gnd 0.009486f
C4031 vdd.n1138 gnd 0.007635f
C4032 vdd.n1139 gnd 0.009486f
C4033 vdd.n1140 gnd 0.567085f
C4034 vdd.n1141 gnd 0.009486f
C4035 vdd.n1142 gnd 0.007635f
C4036 vdd.n1143 gnd 0.009486f
C4037 vdd.n1144 gnd 0.009486f
C4038 vdd.n1145 gnd 0.007291f
C4039 vdd.n1146 gnd 0.009486f
C4040 vdd.n1147 gnd 0.007635f
C4041 vdd.n1148 gnd 0.009486f
C4042 vdd.n1149 gnd 0.445295f
C4043 vdd.n1150 gnd 0.009486f
C4044 vdd.n1151 gnd 0.007635f
C4045 vdd.n1152 gnd 0.009486f
C4046 vdd.n1153 gnd 0.009486f
C4047 vdd.n1154 gnd 0.009486f
C4048 vdd.n1155 gnd 0.007635f
C4049 vdd.n1156 gnd 0.009486f
C4050 vdd.t120 gnd 0.380594f
C4051 vdd.n1157 gnd 0.696487f
C4052 vdd.n1158 gnd 0.009486f
C4053 vdd.n1159 gnd 0.007635f
C4054 vdd.n1160 gnd 0.007291f
C4055 vdd.n1161 gnd 0.009486f
C4056 vdd.n1162 gnd 0.009486f
C4057 vdd.n1163 gnd 0.007635f
C4058 vdd.n1164 gnd 0.009486f
C4059 vdd.n1165 gnd 0.761188f
C4060 vdd.n1166 gnd 0.009486f
C4061 vdd.n1167 gnd 0.007635f
C4062 vdd.n1168 gnd 0.009486f
C4063 vdd.n1169 gnd 0.009486f
C4064 vdd.n1170 gnd 0.009486f
C4065 vdd.n1171 gnd 0.007635f
C4066 vdd.n1172 gnd 0.009486f
C4067 vdd.n1173 gnd 0.574697f
C4068 vdd.n1174 gnd 0.009486f
C4069 vdd.n1175 gnd 0.007635f
C4070 vdd.n1176 gnd 0.009486f
C4071 vdd.n1177 gnd 0.009486f
C4072 vdd.n1178 gnd 0.009486f
C4073 vdd.n1179 gnd 0.007635f
C4074 vdd.n1180 gnd 0.009486f
C4075 vdd.n1181 gnd 0.437683f
C4076 vdd.n1182 gnd 0.009486f
C4077 vdd.n1183 gnd 0.007635f
C4078 vdd.n1184 gnd 0.009486f
C4079 vdd.n1185 gnd 0.009486f
C4080 vdd.n1186 gnd 0.009486f
C4081 vdd.n1187 gnd 0.007635f
C4082 vdd.n1188 gnd 0.009486f
C4083 vdd.t116 gnd 0.380594f
C4084 vdd.n1189 gnd 0.688875f
C4085 vdd.n1190 gnd 0.009486f
C4086 vdd.n1191 gnd 0.007635f
C4087 vdd.n1192 gnd 0.009486f
C4088 vdd.n1193 gnd 0.009486f
C4089 vdd.n1194 gnd 0.009486f
C4090 vdd.n1195 gnd 0.007635f
C4091 vdd.n1196 gnd 0.009486f
C4092 vdd.n1197 gnd 0.761188f
C4093 vdd.n1198 gnd 0.009486f
C4094 vdd.n1199 gnd 0.007635f
C4095 vdd.n1200 gnd 0.009486f
C4096 vdd.n1201 gnd 0.009486f
C4097 vdd.n1202 gnd 0.009486f
C4098 vdd.n1203 gnd 0.007635f
C4099 vdd.n1204 gnd 0.009486f
C4100 vdd.n1205 gnd 0.582309f
C4101 vdd.n1206 gnd 0.009486f
C4102 vdd.n1207 gnd 0.007635f
C4103 vdd.n1208 gnd 0.009486f
C4104 vdd.n1209 gnd 0.009486f
C4105 vdd.n1210 gnd 0.009486f
C4106 vdd.n1211 gnd 0.007635f
C4107 vdd.n1212 gnd 0.009486f
C4108 vdd.n1213 gnd 0.761188f
C4109 vdd.n1214 gnd 0.009486f
C4110 vdd.n1215 gnd 0.007635f
C4111 vdd.n1216 gnd 0.009486f
C4112 vdd.n1217 gnd 0.009486f
C4113 vdd.n1218 gnd 0.009486f
C4114 vdd.n1219 gnd 0.009486f
C4115 vdd.n1220 gnd 0.007635f
C4116 vdd.n1221 gnd 0.009486f
C4117 vdd.t68 gnd 0.380594f
C4118 vdd.n1222 gnd 0.498578f
C4119 vdd.n1223 gnd 0.009486f
C4120 vdd.n1224 gnd 0.007635f
C4121 vdd.n1225 gnd 0.009486f
C4122 vdd.n1226 gnd 0.009486f
C4123 vdd.n1227 gnd 0.009486f
C4124 vdd.n1228 gnd 0.007635f
C4125 vdd.n1230 gnd 0.009486f
C4126 vdd.n1231 gnd 0.009486f
C4127 vdd.n1232 gnd 0.009486f
C4128 vdd.n1233 gnd 0.008158f
C4129 vdd.n1235 gnd 0.009486f
C4130 vdd.n1236 gnd 0.007635f
C4131 vdd.n1237 gnd 0.006071f
C4132 vdd.n1238 gnd 0.007635f
C4133 vdd.n1239 gnd 0.009486f
C4134 vdd.n1241 gnd 0.009486f
C4135 vdd.n1242 gnd 0.009486f
C4136 vdd.n1243 gnd 0.009486f
C4137 vdd.n1244 gnd 0.007635f
C4138 vdd.n1246 gnd 0.009486f
C4139 vdd.n1247 gnd 0.009486f
C4140 vdd.n1248 gnd 0.009486f
C4141 vdd.n1249 gnd 0.009486f
C4142 vdd.n1250 gnd 0.009486f
C4143 vdd.n1251 gnd 0.006375f
C4144 vdd.n1253 gnd 0.009486f
C4145 vdd.n1254 gnd 0.006375f
C4146 vdd.t70 gnd 0.194308f
C4147 vdd.t69 gnd 0.203627f
C4148 vdd.t67 gnd 0.283884f
C4149 vdd.n1255 gnd 0.096222f
C4150 vdd.n1256 gnd 0.055169f
C4151 vdd.n1257 gnd 0.009486f
C4152 vdd.n1258 gnd 0.009486f
C4153 vdd.n1259 gnd 0.007635f
C4154 vdd.n1261 gnd 0.009486f
C4155 vdd.n1262 gnd 0.009486f
C4156 vdd.n1263 gnd 0.009486f
C4157 vdd.n1264 gnd 0.009486f
C4158 vdd.n1265 gnd 0.007635f
C4159 vdd.n1267 gnd 0.009486f
C4160 vdd.n1268 gnd 0.009486f
C4161 vdd.n1269 gnd 0.009486f
C4162 vdd.n1270 gnd 0.009486f
C4163 vdd.n1271 gnd 0.009486f
C4164 vdd.n1272 gnd 0.007635f
C4165 vdd.n1274 gnd 0.009486f
C4166 vdd.n1275 gnd 0.009486f
C4167 vdd.n1276 gnd 0.009486f
C4168 vdd.n1277 gnd 0.009486f
C4169 vdd.n1278 gnd 0.009486f
C4170 vdd.n1279 gnd 0.007635f
C4171 vdd.n1281 gnd 0.009486f
C4172 vdd.n1282 gnd 0.009486f
C4173 vdd.n1283 gnd 0.009486f
C4174 vdd.n1284 gnd 0.009486f
C4175 vdd.n1285 gnd 0.009486f
C4176 vdd.n1286 gnd 0.005192f
C4177 vdd.n1288 gnd 0.009486f
C4178 vdd.n1289 gnd 0.007559f
C4179 vdd.t99 gnd 0.194308f
C4180 vdd.t98 gnd 0.203627f
C4181 vdd.t97 gnd 0.283884f
C4182 vdd.n1290 gnd 0.096222f
C4183 vdd.n1291 gnd 0.055169f
C4184 vdd.n1292 gnd 0.009486f
C4185 vdd.n1293 gnd 0.009486f
C4186 vdd.n1294 gnd 0.007635f
C4187 vdd.n1296 gnd 0.009486f
C4188 vdd.n1297 gnd 0.009486f
C4189 vdd.n1298 gnd 0.009486f
C4190 vdd.n1299 gnd 0.009486f
C4191 vdd.n1300 gnd 0.007635f
C4192 vdd.n1302 gnd 0.009486f
C4193 vdd.n1303 gnd 0.009486f
C4194 vdd.n1304 gnd 0.009486f
C4195 vdd.n1305 gnd 0.009486f
C4196 vdd.n1306 gnd 0.009486f
C4197 vdd.n1307 gnd 0.007635f
C4198 vdd.n1309 gnd 0.007635f
C4199 vdd.n1311 gnd 0.009486f
C4200 vdd.n1312 gnd 0.007635f
C4201 vdd.n1313 gnd 0.009486f
C4202 vdd.n1315 gnd 0.009486f
C4203 vdd.n1316 gnd 0.007635f
C4204 vdd.n1317 gnd 0.009486f
C4205 vdd.n1319 gnd 0.009486f
C4206 vdd.n1320 gnd 0.009486f
C4207 vdd.n1321 gnd 0.007635f
C4208 vdd.n1322 gnd 0.007635f
C4209 vdd.n1323 gnd 0.007635f
C4210 vdd.n1324 gnd 0.009486f
C4211 vdd.n1326 gnd 0.009486f
C4212 vdd.n1327 gnd 0.009486f
C4213 vdd.n1328 gnd 0.007635f
C4214 vdd.n1329 gnd 0.007635f
C4215 vdd.n1330 gnd 0.007635f
C4216 vdd.n1331 gnd 0.009486f
C4217 vdd.n1333 gnd 0.009486f
C4218 vdd.n1334 gnd 0.009486f
C4219 vdd.n1335 gnd 0.007635f
C4220 vdd.n1336 gnd 0.009486f
C4221 vdd.n1337 gnd 0.009486f
C4222 vdd.n1338 gnd 0.009486f
C4223 vdd.n1339 gnd 0.015614f
C4224 vdd.n1340 gnd 0.009486f
C4225 vdd.n1342 gnd 0.009486f
C4226 vdd.n1343 gnd 0.009486f
C4227 vdd.n1344 gnd 0.007635f
C4228 vdd.n1345 gnd 0.007635f
C4229 vdd.n1346 gnd 0.007635f
C4230 vdd.n1347 gnd 0.009486f
C4231 vdd.n1349 gnd 0.009486f
C4232 vdd.n1350 gnd 0.009486f
C4233 vdd.n1351 gnd 0.007635f
C4234 vdd.n1352 gnd 0.007635f
C4235 vdd.n1353 gnd 0.007635f
C4236 vdd.n1354 gnd 0.009486f
C4237 vdd.n1356 gnd 0.009486f
C4238 vdd.n1357 gnd 0.009486f
C4239 vdd.n1358 gnd 0.007635f
C4240 vdd.n1359 gnd 0.007635f
C4241 vdd.n1360 gnd 0.007635f
C4242 vdd.n1361 gnd 0.009486f
C4243 vdd.n1363 gnd 0.009486f
C4244 vdd.n1364 gnd 0.009486f
C4245 vdd.n1365 gnd 0.007635f
C4246 vdd.n1366 gnd 0.007635f
C4247 vdd.n1367 gnd 0.007635f
C4248 vdd.n1368 gnd 0.009486f
C4249 vdd.n1370 gnd 0.009486f
C4250 vdd.n1371 gnd 0.009486f
C4251 vdd.n1372 gnd 0.007635f
C4252 vdd.n1373 gnd 0.009486f
C4253 vdd.n1374 gnd 0.009486f
C4254 vdd.n1375 gnd 0.009486f
C4255 vdd.n1376 gnd 0.015614f
C4256 vdd.n1377 gnd 0.009486f
C4257 vdd.n1379 gnd 0.009486f
C4258 vdd.n1380 gnd 0.009486f
C4259 vdd.n1381 gnd 0.007635f
C4260 vdd.n1382 gnd 0.007635f
C4261 vdd.n1383 gnd 0.007635f
C4262 vdd.n1384 gnd 0.009486f
C4263 vdd.n1386 gnd 0.009486f
C4264 vdd.n1387 gnd 0.009486f
C4265 vdd.n1388 gnd 0.007635f
C4266 vdd.n1389 gnd 0.007635f
C4267 vdd.n1390 gnd 0.007635f
C4268 vdd.n1391 gnd 0.009486f
C4269 vdd.n1393 gnd 0.009486f
C4270 vdd.n1394 gnd 0.009486f
C4271 vdd.n1395 gnd 0.007635f
C4272 vdd.n1397 gnd 0.48107f
C4273 vdd.n1399 gnd 0.007635f
C4274 vdd.n1400 gnd 0.007635f
C4275 vdd.n1401 gnd 0.007635f
C4276 vdd.n1402 gnd 0.009486f
C4277 vdd.n1404 gnd 0.009486f
C4278 vdd.n1405 gnd 0.009486f
C4279 vdd.n1406 gnd 0.007635f
C4280 vdd.n1407 gnd 0.006337f
C4281 vdd.n1408 gnd 0.021375f
C4282 vdd.n1409 gnd 0.021312f
C4283 vdd.n1410 gnd 0.006337f
C4284 vdd.n1411 gnd 0.021312f
C4285 vdd.n1412 gnd 0.978126f
C4286 vdd.n1413 gnd 0.021312f
C4287 vdd.n1414 gnd 0.021375f
C4288 vdd.n1415 gnd 0.003627f
C4289 vdd.n1416 gnd 0.021375f
C4290 vdd.n1417 gnd 0.009486f
C4291 vdd.n1418 gnd 0.009486f
C4292 vdd.n1419 gnd 0.007635f
C4293 vdd.n1420 gnd 0.007635f
C4294 vdd.n1421 gnd 0.007635f
C4295 vdd.n1422 gnd 0.008158f
C4296 vdd.n1423 gnd 0.48107f
C4297 vdd.n1424 gnd 0.012762f
C4298 vdd.n1425 gnd 0.004838f
C4299 vdd.n1426 gnd 0.00645f
C4300 vdd.n1427 gnd 0.00645f
C4301 vdd.n1428 gnd 0.00645f
C4302 vdd.n1429 gnd 0.00645f
C4303 vdd.n1430 gnd 0.00645f
C4304 vdd.n1432 gnd 0.00645f
C4305 vdd.n1433 gnd 0.00645f
C4306 vdd.n1434 gnd 0.00645f
C4307 vdd.n1435 gnd 0.00645f
C4308 vdd.n1436 gnd 0.00645f
C4309 vdd.n1438 gnd 0.00645f
C4310 vdd.n1440 gnd 0.00645f
C4311 vdd.n1441 gnd 0.00645f
C4312 vdd.n1442 gnd 0.00645f
C4313 vdd.n1443 gnd 0.00645f
C4314 vdd.n1444 gnd 0.00645f
C4315 vdd.n1446 gnd 0.00645f
C4316 vdd.n1448 gnd 0.00645f
C4317 vdd.n1449 gnd 0.00645f
C4318 vdd.n1450 gnd 0.00645f
C4319 vdd.n1451 gnd 0.00645f
C4320 vdd.n1452 gnd 0.00645f
C4321 vdd.n1454 gnd 0.00645f
C4322 vdd.n1456 gnd 0.00645f
C4323 vdd.n1457 gnd 0.004838f
C4324 vdd.n1458 gnd 0.00645f
C4325 vdd.n1459 gnd 0.00645f
C4326 vdd.n1460 gnd 0.00645f
C4327 vdd.n1462 gnd 0.00645f
C4328 vdd.n1464 gnd 0.00645f
C4329 vdd.n1465 gnd 0.00645f
C4330 vdd.n1466 gnd 0.00645f
C4331 vdd.n1467 gnd 0.00645f
C4332 vdd.n1468 gnd 0.00645f
C4333 vdd.n1470 gnd 0.00645f
C4334 vdd.n1472 gnd 0.00645f
C4335 vdd.n1473 gnd 0.00645f
C4336 vdd.n1474 gnd 0.00498f
C4337 vdd.n1475 gnd 0.009219f
C4338 vdd.n1476 gnd 0.004696f
C4339 vdd.n1477 gnd 0.00645f
C4340 vdd.n1479 gnd 0.00645f
C4341 vdd.n1480 gnd 0.015081f
C4342 vdd.n1481 gnd 0.015081f
C4343 vdd.n1482 gnd 0.014326f
C4344 vdd.n1483 gnd 0.00645f
C4345 vdd.n1484 gnd 0.00645f
C4346 vdd.n1485 gnd 0.00645f
C4347 vdd.n1486 gnd 0.00645f
C4348 vdd.n1487 gnd 0.00645f
C4349 vdd.n1488 gnd 0.00645f
C4350 vdd.n1489 gnd 0.00645f
C4351 vdd.n1490 gnd 0.00645f
C4352 vdd.n1491 gnd 0.00645f
C4353 vdd.n1492 gnd 0.00645f
C4354 vdd.n1493 gnd 0.00645f
C4355 vdd.n1494 gnd 0.00645f
C4356 vdd.n1495 gnd 0.00645f
C4357 vdd.n1496 gnd 0.00645f
C4358 vdd.n1497 gnd 0.00645f
C4359 vdd.n1498 gnd 0.00645f
C4360 vdd.n1499 gnd 0.00645f
C4361 vdd.n1500 gnd 0.00645f
C4362 vdd.n1501 gnd 0.00645f
C4363 vdd.n1502 gnd 0.00645f
C4364 vdd.n1503 gnd 0.00645f
C4365 vdd.n1504 gnd 0.00645f
C4366 vdd.n1505 gnd 0.00645f
C4367 vdd.n1506 gnd 0.00645f
C4368 vdd.n1507 gnd 0.00645f
C4369 vdd.n1508 gnd 0.00645f
C4370 vdd.n1509 gnd 0.00645f
C4371 vdd.n1510 gnd 0.00645f
C4372 vdd.n1511 gnd 0.00645f
C4373 vdd.n1512 gnd 0.00645f
C4374 vdd.n1513 gnd 0.00645f
C4375 vdd.n1514 gnd 0.00645f
C4376 vdd.n1515 gnd 0.00645f
C4377 vdd.n1516 gnd 0.00645f
C4378 vdd.n1517 gnd 0.00645f
C4379 vdd.n1518 gnd 0.00645f
C4380 vdd.n1519 gnd 0.00645f
C4381 vdd.n1520 gnd 0.00645f
C4382 vdd.n1521 gnd 0.00645f
C4383 vdd.n1522 gnd 0.00645f
C4384 vdd.n1523 gnd 0.00645f
C4385 vdd.n1524 gnd 0.00645f
C4386 vdd.n1525 gnd 0.00645f
C4387 vdd.n1526 gnd 0.00645f
C4388 vdd.n1527 gnd 0.00645f
C4389 vdd.n1528 gnd 0.00645f
C4390 vdd.n1529 gnd 0.00645f
C4391 vdd.n1530 gnd 0.00645f
C4392 vdd.n1531 gnd 0.00645f
C4393 vdd.n1532 gnd 0.00645f
C4394 vdd.n1533 gnd 0.00645f
C4395 vdd.n1534 gnd 0.00645f
C4396 vdd.n1535 gnd 0.00645f
C4397 vdd.n1536 gnd 0.00645f
C4398 vdd.n1537 gnd 0.00645f
C4399 vdd.n1538 gnd 0.00645f
C4400 vdd.n1539 gnd 0.00645f
C4401 vdd.n1540 gnd 0.00645f
C4402 vdd.n1541 gnd 0.00645f
C4403 vdd.n1542 gnd 0.00645f
C4404 vdd.n1543 gnd 0.00645f
C4405 vdd.n1544 gnd 0.00645f
C4406 vdd.n1545 gnd 0.00645f
C4407 vdd.n1546 gnd 0.00645f
C4408 vdd.n1547 gnd 0.00645f
C4409 vdd.n1548 gnd 0.00645f
C4410 vdd.n1549 gnd 0.00645f
C4411 vdd.n1550 gnd 0.00645f
C4412 vdd.n1551 gnd 0.00645f
C4413 vdd.n1552 gnd 0.00645f
C4414 vdd.n1553 gnd 0.34634f
C4415 vdd.n1554 gnd 0.00645f
C4416 vdd.n1555 gnd 0.00645f
C4417 vdd.n1556 gnd 0.00645f
C4418 vdd.n1557 gnd 0.00645f
C4419 vdd.n1558 gnd 0.00645f
C4420 vdd.n1559 gnd 0.00645f
C4421 vdd.n1560 gnd 0.00645f
C4422 vdd.n1561 gnd 0.00645f
C4423 vdd.n1562 gnd 0.34634f
C4424 vdd.n1563 gnd 0.00645f
C4425 vdd.n1564 gnd 0.00645f
C4426 vdd.n1565 gnd 0.00645f
C4427 vdd.n1566 gnd 0.00645f
C4428 vdd.n1567 gnd 0.00645f
C4429 vdd.n1568 gnd 0.00645f
C4430 vdd.n1569 gnd 0.00645f
C4431 vdd.n1570 gnd 0.00645f
C4432 vdd.n1571 gnd 0.00645f
C4433 vdd.n1572 gnd 0.00645f
C4434 vdd.n1573 gnd 0.00645f
C4435 vdd.n1574 gnd 0.00645f
C4436 vdd.n1575 gnd 0.00645f
C4437 vdd.n1576 gnd 0.00645f
C4438 vdd.n1577 gnd 0.00645f
C4439 vdd.n1578 gnd 0.00645f
C4440 vdd.n1579 gnd 0.00645f
C4441 vdd.n1580 gnd 0.00645f
C4442 vdd.n1581 gnd 0.00645f
C4443 vdd.n1582 gnd 0.00645f
C4444 vdd.n1583 gnd 0.00645f
C4445 vdd.n1584 gnd 0.00645f
C4446 vdd.n1585 gnd 0.00645f
C4447 vdd.n1586 gnd 0.00645f
C4448 vdd.n1587 gnd 0.00645f
C4449 vdd.n1588 gnd 0.00645f
C4450 vdd.n1589 gnd 0.00645f
C4451 vdd.n1590 gnd 0.00645f
C4452 vdd.n1591 gnd 0.00645f
C4453 vdd.n1592 gnd 0.00645f
C4454 vdd.n1593 gnd 0.00645f
C4455 vdd.n1594 gnd 0.00645f
C4456 vdd.n1595 gnd 0.014326f
C4457 vdd.n1596 gnd 0.015081f
C4458 vdd.n1597 gnd 0.015081f
C4459 vdd.n1598 gnd 0.00645f
C4460 vdd.n1599 gnd 0.00645f
C4461 vdd.n1600 gnd 0.004696f
C4462 vdd.n1601 gnd 0.00645f
C4463 vdd.n1603 gnd 0.00645f
C4464 vdd.n1604 gnd 0.00498f
C4465 vdd.n1605 gnd 0.00645f
C4466 vdd.n1606 gnd 0.00645f
C4467 vdd.n1607 gnd 0.00645f
C4468 vdd.n1609 gnd 0.00645f
C4469 vdd.n1611 gnd 0.00645f
C4470 vdd.n1612 gnd 0.00645f
C4471 vdd.n1613 gnd 0.00645f
C4472 vdd.n1614 gnd 0.00645f
C4473 vdd.n1615 gnd 0.00645f
C4474 vdd.n1617 gnd 0.00645f
C4475 vdd.n1618 gnd 0.00645f
C4476 vdd.n1619 gnd 0.00645f
C4477 vdd.n1620 gnd 0.004838f
C4478 vdd.n1621 gnd 0.00645f
C4479 vdd.n1623 gnd 0.00645f
C4480 vdd.n1624 gnd 0.004838f
C4481 vdd.n1625 gnd 0.00645f
C4482 vdd.n1626 gnd 0.00645f
C4483 vdd.n1627 gnd 0.00645f
C4484 vdd.n1629 gnd 0.00645f
C4485 vdd.n1631 gnd 0.00645f
C4486 vdd.n1632 gnd 0.00645f
C4487 vdd.n1633 gnd 0.00645f
C4488 vdd.n1634 gnd 0.00645f
C4489 vdd.n1635 gnd 0.00645f
C4490 vdd.n1637 gnd 0.00645f
C4491 vdd.n1638 gnd 0.00645f
C4492 vdd.n1639 gnd 0.00645f
C4493 vdd.n1640 gnd 0.00645f
C4494 vdd.n1641 gnd 0.00645f
C4495 vdd.n1642 gnd 0.00645f
C4496 vdd.n1644 gnd 0.00645f
C4497 vdd.n1645 gnd 0.00645f
C4498 vdd.n1646 gnd 0.015081f
C4499 vdd.n1647 gnd 0.014326f
C4500 vdd.n1648 gnd 0.014326f
C4501 vdd.n1649 gnd 0.715516f
C4502 vdd.n1650 gnd 0.014326f
C4503 vdd.n1651 gnd 0.014326f
C4504 vdd.n1652 gnd 0.00645f
C4505 vdd.n1653 gnd 0.00645f
C4506 vdd.n1654 gnd 0.00645f
C4507 vdd.n1655 gnd 0.517608f
C4508 vdd.n1656 gnd 0.00645f
C4509 vdd.n1657 gnd 0.00645f
C4510 vdd.n1658 gnd 0.00645f
C4511 vdd.n1659 gnd 0.00645f
C4512 vdd.n1660 gnd 0.00645f
C4513 vdd.n1661 gnd 0.490966f
C4514 vdd.n1662 gnd 0.00645f
C4515 vdd.n1663 gnd 0.00645f
C4516 vdd.n1664 gnd 0.005407f
C4517 vdd.n1665 gnd 0.018686f
C4518 vdd.n1666 gnd 0.004269f
C4519 vdd.n1667 gnd 0.00645f
C4520 vdd.n1668 gnd 0.342534f
C4521 vdd.n1669 gnd 0.00645f
C4522 vdd.n1670 gnd 0.00645f
C4523 vdd.n1671 gnd 0.00645f
C4524 vdd.n1672 gnd 0.00645f
C4525 vdd.n1673 gnd 0.00645f
C4526 vdd.n1674 gnd 0.517608f
C4527 vdd.n1675 gnd 0.00645f
C4528 vdd.n1676 gnd 0.00645f
C4529 vdd.n1677 gnd 0.00645f
C4530 vdd.n1678 gnd 0.00645f
C4531 vdd.n1679 gnd 0.00645f
C4532 vdd.n1680 gnd 0.315893f
C4533 vdd.n1681 gnd 0.00645f
C4534 vdd.n1682 gnd 0.00645f
C4535 vdd.n1683 gnd 0.00645f
C4536 vdd.n1684 gnd 0.00645f
C4537 vdd.n1685 gnd 0.00645f
C4538 vdd.n1686 gnd 0.464324f
C4539 vdd.n1687 gnd 0.00645f
C4540 vdd.n1688 gnd 0.00645f
C4541 vdd.n1689 gnd 0.00645f
C4542 vdd.n1690 gnd 0.00645f
C4543 vdd.n1691 gnd 0.00645f
C4544 vdd.n1692 gnd 0.293057f
C4545 vdd.n1693 gnd 0.00645f
C4546 vdd.n1694 gnd 0.00645f
C4547 vdd.n1695 gnd 0.00645f
C4548 vdd.n1696 gnd 0.00645f
C4549 vdd.n1697 gnd 0.00645f
C4550 vdd.n1698 gnd 0.441489f
C4551 vdd.n1699 gnd 0.00645f
C4552 vdd.n1700 gnd 0.00645f
C4553 vdd.n1701 gnd 0.00645f
C4554 vdd.n1702 gnd 0.00645f
C4555 vdd.n1703 gnd 0.00645f
C4556 vdd.n1704 gnd 0.270222f
C4557 vdd.n1705 gnd 0.00645f
C4558 vdd.n1706 gnd 0.00645f
C4559 vdd.n1707 gnd 0.00645f
C4560 vdd.n1708 gnd 0.00645f
C4561 vdd.n1709 gnd 0.00645f
C4562 vdd.n1710 gnd 0.418653f
C4563 vdd.n1711 gnd 0.00645f
C4564 vdd.n1712 gnd 0.00645f
C4565 vdd.n1713 gnd 0.00645f
C4566 vdd.n1714 gnd 0.00645f
C4567 vdd.n1715 gnd 0.00645f
C4568 vdd.n1716 gnd 0.270222f
C4569 vdd.n1717 gnd 0.00645f
C4570 vdd.n1718 gnd 0.00645f
C4571 vdd.n1719 gnd 0.00645f
C4572 vdd.n1720 gnd 0.00645f
C4573 vdd.n1721 gnd 0.00645f
C4574 vdd.n1722 gnd 0.395818f
C4575 vdd.n1723 gnd 0.00645f
C4576 vdd.n1724 gnd 0.00645f
C4577 vdd.n1725 gnd 0.00645f
C4578 vdd.n1726 gnd 0.00645f
C4579 vdd.n1727 gnd 0.00645f
C4580 vdd.n1728 gnd 0.293057f
C4581 vdd.n1729 gnd 0.00645f
C4582 vdd.n1730 gnd 0.00645f
C4583 vdd.n1731 gnd 0.00645f
C4584 vdd.n1732 gnd 0.00645f
C4585 vdd.n1733 gnd 0.00645f
C4586 vdd.n1734 gnd 0.517608f
C4587 vdd.n1735 gnd 0.00645f
C4588 vdd.n1736 gnd 0.00645f
C4589 vdd.n1737 gnd 0.00645f
C4590 vdd.n1738 gnd 0.00645f
C4591 vdd.n1739 gnd 0.00645f
C4592 vdd.n1740 gnd 0.201715f
C4593 vdd.n1741 gnd 0.00645f
C4594 vdd.n1742 gnd 0.00645f
C4595 vdd.n1743 gnd 0.00645f
C4596 vdd.n1744 gnd 0.00645f
C4597 vdd.n1745 gnd 0.00645f
C4598 vdd.n1746 gnd 0.517608f
C4599 vdd.n1747 gnd 0.00645f
C4600 vdd.n1748 gnd 0.00645f
C4601 vdd.n1749 gnd 0.00645f
C4602 vdd.n1750 gnd 0.00645f
C4603 vdd.n1751 gnd 0.00645f
C4604 vdd.n1752 gnd 0.380594f
C4605 vdd.n1753 gnd 0.00645f
C4606 vdd.n1754 gnd 0.00645f
C4607 vdd.n1755 gnd 0.00645f
C4608 vdd.n1756 gnd 0.00645f
C4609 vdd.n1757 gnd 0.00645f
C4610 vdd.n1758 gnd 0.00645f
C4611 vdd.n1759 gnd 0.490966f
C4612 vdd.n1760 gnd 0.00645f
C4613 vdd.n1761 gnd 0.00645f
C4614 vdd.n1762 gnd 0.00645f
C4615 vdd.n1763 gnd 0.00645f
C4616 vdd.n1764 gnd 0.00645f
C4617 vdd.n1765 gnd 0.00645f
C4618 vdd.n1766 gnd 0.357758f
C4619 vdd.n1767 gnd 0.00645f
C4620 vdd.n1768 gnd 0.00645f
C4621 vdd.n1769 gnd 0.00645f
C4622 vdd.n1770 gnd 0.015119f
C4623 vdd.n1771 gnd 0.014326f
C4624 vdd.n1772 gnd 0.015081f
C4625 vdd.n1773 gnd 0.014287f
C4626 vdd.n1774 gnd 0.00645f
C4627 vdd.n1775 gnd 0.00645f
C4628 vdd.n1776 gnd 0.00645f
C4629 vdd.n1777 gnd 0.004696f
C4630 vdd.n1778 gnd 0.009219f
C4631 vdd.n1779 gnd 0.00498f
C4632 vdd.n1780 gnd 0.00645f
C4633 vdd.n1781 gnd 0.00645f
C4634 vdd.n1782 gnd 0.00645f
C4635 vdd.n1783 gnd 0.00645f
C4636 vdd.n1784 gnd 0.00645f
C4637 vdd.n1785 gnd 0.00645f
C4638 vdd.n1786 gnd 0.00645f
C4639 vdd.n1787 gnd 0.00645f
C4640 vdd.n1788 gnd 0.00645f
C4641 vdd.n1789 gnd 0.00645f
C4642 vdd.n1790 gnd 0.00645f
C4643 vdd.n1791 gnd 0.00645f
C4644 vdd.n1792 gnd 0.00645f
C4645 vdd.n1793 gnd 0.00645f
C4646 vdd.n1794 gnd 0.00645f
C4647 vdd.n1795 gnd 0.00645f
C4648 vdd.n1796 gnd 0.00645f
C4649 vdd.n1797 gnd 0.00645f
C4650 vdd.n1798 gnd 0.00645f
C4651 vdd.n1799 gnd 0.00645f
C4652 vdd.n1800 gnd 0.00645f
C4653 vdd.n1801 gnd 0.00645f
C4654 vdd.n1802 gnd 0.00645f
C4655 vdd.n1803 gnd 0.00645f
C4656 vdd.n1804 gnd 0.00645f
C4657 vdd.n1805 gnd 0.00645f
C4658 vdd.n1806 gnd 0.00645f
C4659 vdd.n1807 gnd 0.00645f
C4660 vdd.n1808 gnd 0.00645f
C4661 vdd.n1809 gnd 0.00645f
C4662 vdd.n1810 gnd 0.00645f
C4663 vdd.n1811 gnd 0.00645f
C4664 vdd.n1812 gnd 0.00645f
C4665 vdd.n1813 gnd 0.00645f
C4666 vdd.n1814 gnd 0.00645f
C4667 vdd.n1815 gnd 0.00645f
C4668 vdd.n1816 gnd 0.00645f
C4669 vdd.n1817 gnd 0.00645f
C4670 vdd.n1818 gnd 0.00645f
C4671 vdd.n1819 gnd 0.00645f
C4672 vdd.n1820 gnd 0.00645f
C4673 vdd.n1821 gnd 0.00645f
C4674 vdd.n1822 gnd 0.00645f
C4675 vdd.n1823 gnd 0.015081f
C4676 vdd.n1824 gnd 0.015081f
C4677 vdd.n1825 gnd 0.014326f
C4678 vdd.n1826 gnd 0.00645f
C4679 vdd.n1827 gnd 0.00645f
C4680 vdd.n1828 gnd 0.418653f
C4681 vdd.n1829 gnd 0.00645f
C4682 vdd.n1830 gnd 0.014326f
C4683 vdd.n1831 gnd 0.015119f
C4684 vdd.n1832 gnd 0.014287f
C4685 vdd.n1833 gnd 0.00645f
C4686 vdd.n1834 gnd 0.00645f
C4687 vdd.n1835 gnd 0.004696f
C4688 vdd.n1836 gnd 0.00645f
C4689 vdd.n1837 gnd 0.00645f
C4690 vdd.n1838 gnd 0.00498f
C4691 vdd.n1839 gnd 0.00645f
C4692 vdd.n1840 gnd 0.00645f
C4693 vdd.n1841 gnd 0.00645f
C4694 vdd.n1842 gnd 0.00645f
C4695 vdd.n1843 gnd 0.00645f
C4696 vdd.n1844 gnd 0.00645f
C4697 vdd.n1845 gnd 0.00645f
C4698 vdd.n1846 gnd 0.00645f
C4699 vdd.n1847 gnd 0.00645f
C4700 vdd.n1848 gnd 0.00645f
C4701 vdd.n1849 gnd 0.00645f
C4702 vdd.n1850 gnd 0.00645f
C4703 vdd.n1851 gnd 0.00645f
C4704 vdd.n1852 gnd 0.00645f
C4705 vdd.n1853 gnd 0.00645f
C4706 vdd.n1854 gnd 0.00645f
C4707 vdd.n1855 gnd 0.00645f
C4708 vdd.n1856 gnd 0.00645f
C4709 vdd.n1857 gnd 0.00645f
C4710 vdd.n1858 gnd 0.00645f
C4711 vdd.n1859 gnd 0.00645f
C4712 vdd.n1860 gnd 0.00645f
C4713 vdd.n1861 gnd 0.00645f
C4714 vdd.n1862 gnd 0.00645f
C4715 vdd.n1863 gnd 0.00645f
C4716 vdd.n1864 gnd 0.00645f
C4717 vdd.n1865 gnd 0.00645f
C4718 vdd.n1866 gnd 0.00645f
C4719 vdd.n1867 gnd 0.00645f
C4720 vdd.n1868 gnd 0.00645f
C4721 vdd.n1869 gnd 0.00645f
C4722 vdd.n1870 gnd 0.00645f
C4723 vdd.n1871 gnd 0.00645f
C4724 vdd.n1872 gnd 0.00645f
C4725 vdd.n1873 gnd 0.00645f
C4726 vdd.n1874 gnd 0.00645f
C4727 vdd.n1875 gnd 0.00645f
C4728 vdd.n1876 gnd 0.00645f
C4729 vdd.n1877 gnd 0.00645f
C4730 vdd.n1878 gnd 0.00645f
C4731 vdd.n1879 gnd 0.00645f
C4732 vdd.n1880 gnd 0.015081f
C4733 vdd.n1881 gnd 0.015081f
C4734 vdd.n1882 gnd 0.593726f
C4735 vdd.t165 gnd 2.6261f
C4736 vdd.t174 gnd 2.6261f
C4737 vdd.n1883 gnd 0.593726f
C4738 vdd.n1884 gnd 0.014326f
C4739 vdd.n1885 gnd 0.014326f
C4740 vdd.n1886 gnd 0.418653f
C4741 vdd.n1887 gnd 0.015081f
C4742 vdd.n1888 gnd 0.00645f
C4743 vdd.n1889 gnd 0.00645f
C4744 vdd.n1890 gnd 0.00645f
C4745 vdd.n1891 gnd 0.00645f
C4746 vdd.n1892 gnd 0.00645f
C4747 vdd.n1893 gnd 0.00645f
C4748 vdd.n1894 gnd 0.00645f
C4749 vdd.n1895 gnd 0.00645f
C4750 vdd.n1896 gnd 0.00645f
C4751 vdd.n1897 gnd 0.00645f
C4752 vdd.n1898 gnd 0.00498f
C4753 vdd.n1899 gnd 0.00645f
C4754 vdd.t101 gnd 0.082471f
C4755 vdd.t102 gnd 0.093776f
C4756 vdd.t100 gnd 0.246066f
C4757 vdd.n1900 gnd 0.164301f
C4758 vdd.n1901 gnd 0.132315f
C4759 vdd.n1902 gnd 0.009219f
C4760 vdd.n1903 gnd 0.00645f
C4761 vdd.n1904 gnd 0.00645f
C4762 vdd.n1905 gnd 0.00645f
C4763 vdd.t48 gnd 0.082471f
C4764 vdd.t49 gnd 0.093776f
C4765 vdd.t46 gnd 0.246066f
C4766 vdd.n1906 gnd 0.164301f
C4767 vdd.n1907 gnd 0.132315f
C4768 vdd.n1908 gnd 0.00645f
C4769 vdd.n1909 gnd 0.00645f
C4770 vdd.n1910 gnd 0.00645f
C4771 vdd.n1911 gnd 0.00645f
C4772 vdd.n1912 gnd 0.00645f
C4773 vdd.n1913 gnd 0.00645f
C4774 vdd.n1914 gnd 0.00645f
C4775 vdd.n1915 gnd 0.00645f
C4776 vdd.n1916 gnd 0.00645f
C4777 vdd.n1917 gnd 0.00645f
C4778 vdd.n1919 gnd 0.00645f
C4779 vdd.n1920 gnd 0.00645f
C4780 vdd.n1921 gnd 0.00645f
C4781 vdd.n1922 gnd 0.00645f
C4782 vdd.n1923 gnd 0.00645f
C4783 vdd.n1925 gnd 0.00645f
C4784 vdd.n1927 gnd 0.00645f
C4785 vdd.n1928 gnd 0.00645f
C4786 vdd.n1929 gnd 0.00645f
C4787 vdd.n1930 gnd 0.00645f
C4788 vdd.n1931 gnd 0.00645f
C4789 vdd.n1933 gnd 0.00645f
C4790 vdd.n1935 gnd 0.00645f
C4791 vdd.n1936 gnd 0.00645f
C4792 vdd.n1937 gnd 0.00645f
C4793 vdd.n1938 gnd 0.00645f
C4794 vdd.n1939 gnd 0.00645f
C4795 vdd.n1941 gnd 0.00645f
C4796 vdd.n1943 gnd 0.00645f
C4797 vdd.n1944 gnd 0.00645f
C4798 vdd.n1945 gnd 0.00645f
C4799 vdd.n1946 gnd 0.00645f
C4800 vdd.n1947 gnd 0.00645f
C4801 vdd.n1949 gnd 0.00645f
C4802 vdd.n1951 gnd 0.00645f
C4803 vdd.n1952 gnd 0.00645f
C4804 vdd.n1953 gnd 0.00645f
C4805 vdd.n1954 gnd 0.00645f
C4806 vdd.n1955 gnd 0.00645f
C4807 vdd.n1957 gnd 0.00645f
C4808 vdd.n1959 gnd 0.00645f
C4809 vdd.n1960 gnd 0.00645f
C4810 vdd.n1961 gnd 0.00498f
C4811 vdd.n1962 gnd 0.009219f
C4812 vdd.n1963 gnd 0.004696f
C4813 vdd.n1964 gnd 0.00645f
C4814 vdd.n1966 gnd 0.00645f
C4815 vdd.n1967 gnd 0.015081f
C4816 vdd.n1968 gnd 0.015081f
C4817 vdd.n1969 gnd 0.014326f
C4818 vdd.n1970 gnd 0.00645f
C4819 vdd.n1971 gnd 0.00645f
C4820 vdd.n1972 gnd 0.00645f
C4821 vdd.n1973 gnd 0.00645f
C4822 vdd.n1974 gnd 0.00645f
C4823 vdd.n1975 gnd 0.00645f
C4824 vdd.n1976 gnd 0.00645f
C4825 vdd.n1977 gnd 0.00645f
C4826 vdd.n1978 gnd 0.00645f
C4827 vdd.n1979 gnd 0.00645f
C4828 vdd.n1980 gnd 0.00645f
C4829 vdd.n1981 gnd 0.00645f
C4830 vdd.n1982 gnd 0.00645f
C4831 vdd.n1983 gnd 0.00645f
C4832 vdd.n1984 gnd 0.00645f
C4833 vdd.n1985 gnd 0.00645f
C4834 vdd.n1986 gnd 0.00645f
C4835 vdd.n1987 gnd 0.00645f
C4836 vdd.n1988 gnd 0.00645f
C4837 vdd.n1989 gnd 0.00645f
C4838 vdd.n1990 gnd 0.00645f
C4839 vdd.n1991 gnd 0.00645f
C4840 vdd.n1992 gnd 0.00645f
C4841 vdd.n1993 gnd 0.00645f
C4842 vdd.n1994 gnd 0.00645f
C4843 vdd.n1995 gnd 0.00645f
C4844 vdd.n1996 gnd 0.00645f
C4845 vdd.n1997 gnd 0.00645f
C4846 vdd.n1998 gnd 0.00645f
C4847 vdd.n1999 gnd 0.00645f
C4848 vdd.n2000 gnd 0.00645f
C4849 vdd.n2001 gnd 0.00645f
C4850 vdd.n2002 gnd 0.00645f
C4851 vdd.n2003 gnd 0.00645f
C4852 vdd.n2004 gnd 0.00645f
C4853 vdd.n2005 gnd 0.00645f
C4854 vdd.n2006 gnd 0.00645f
C4855 vdd.n2007 gnd 0.00645f
C4856 vdd.n2008 gnd 0.00645f
C4857 vdd.n2009 gnd 0.00645f
C4858 vdd.n2010 gnd 0.00645f
C4859 vdd.n2011 gnd 0.00645f
C4860 vdd.n2012 gnd 0.00645f
C4861 vdd.n2013 gnd 0.00645f
C4862 vdd.n2014 gnd 0.00645f
C4863 vdd.n2015 gnd 0.00645f
C4864 vdd.n2016 gnd 0.00645f
C4865 vdd.n2017 gnd 0.00645f
C4866 vdd.n2018 gnd 0.00645f
C4867 vdd.n2019 gnd 0.00645f
C4868 vdd.n2020 gnd 0.00645f
C4869 vdd.n2021 gnd 0.00645f
C4870 vdd.n2022 gnd 0.00645f
C4871 vdd.n2023 gnd 0.00645f
C4872 vdd.n2024 gnd 0.00645f
C4873 vdd.n2025 gnd 0.00645f
C4874 vdd.n2026 gnd 0.00645f
C4875 vdd.n2027 gnd 0.00645f
C4876 vdd.n2028 gnd 0.00645f
C4877 vdd.n2029 gnd 0.00645f
C4878 vdd.n2030 gnd 0.00645f
C4879 vdd.n2031 gnd 0.00645f
C4880 vdd.n2032 gnd 0.00645f
C4881 vdd.n2033 gnd 0.00645f
C4882 vdd.n2034 gnd 0.00645f
C4883 vdd.n2035 gnd 0.00645f
C4884 vdd.n2036 gnd 0.00645f
C4885 vdd.n2037 gnd 0.00645f
C4886 vdd.n2038 gnd 0.00645f
C4887 vdd.n2039 gnd 0.00645f
C4888 vdd.n2040 gnd 0.00645f
C4889 vdd.n2041 gnd 0.00645f
C4890 vdd.n2042 gnd 0.00645f
C4891 vdd.n2043 gnd 0.00645f
C4892 vdd.n2044 gnd 0.00645f
C4893 vdd.n2045 gnd 0.00645f
C4894 vdd.n2046 gnd 0.00645f
C4895 vdd.n2047 gnd 0.00645f
C4896 vdd.n2048 gnd 0.00645f
C4897 vdd.n2049 gnd 0.00645f
C4898 vdd.n2050 gnd 0.00645f
C4899 vdd.n2051 gnd 0.34634f
C4900 vdd.n2052 gnd 0.00645f
C4901 vdd.n2053 gnd 0.00645f
C4902 vdd.n2054 gnd 0.00645f
C4903 vdd.n2055 gnd 0.00645f
C4904 vdd.n2056 gnd 0.00645f
C4905 vdd.n2057 gnd 0.00645f
C4906 vdd.n2058 gnd 0.00645f
C4907 vdd.n2059 gnd 0.00645f
C4908 vdd.n2060 gnd 0.34634f
C4909 vdd.n2061 gnd 0.00645f
C4910 vdd.n2062 gnd 0.00645f
C4911 vdd.n2063 gnd 0.00645f
C4912 vdd.n2064 gnd 0.00645f
C4913 vdd.n2065 gnd 0.00645f
C4914 vdd.n2066 gnd 0.00645f
C4915 vdd.n2067 gnd 0.00645f
C4916 vdd.n2068 gnd 0.00645f
C4917 vdd.n2069 gnd 0.00645f
C4918 vdd.n2070 gnd 0.00645f
C4919 vdd.n2071 gnd 0.00645f
C4920 vdd.n2072 gnd 0.00645f
C4921 vdd.n2073 gnd 0.00645f
C4922 vdd.n2074 gnd 0.00645f
C4923 vdd.n2075 gnd 0.00645f
C4924 vdd.n2076 gnd 0.00645f
C4925 vdd.n2077 gnd 0.00645f
C4926 vdd.n2078 gnd 0.00645f
C4927 vdd.n2079 gnd 0.00645f
C4928 vdd.n2080 gnd 0.00645f
C4929 vdd.n2081 gnd 0.00645f
C4930 vdd.n2082 gnd 0.00645f
C4931 vdd.n2083 gnd 0.00645f
C4932 vdd.n2084 gnd 0.014326f
C4933 vdd.n2086 gnd 0.015081f
C4934 vdd.n2087 gnd 0.015081f
C4935 vdd.n2088 gnd 0.00645f
C4936 vdd.n2089 gnd 0.004696f
C4937 vdd.n2090 gnd 0.00645f
C4938 vdd.n2092 gnd 0.00645f
C4939 vdd.n2094 gnd 0.00645f
C4940 vdd.n2095 gnd 0.00645f
C4941 vdd.n2096 gnd 0.00645f
C4942 vdd.n2097 gnd 0.00645f
C4943 vdd.n2098 gnd 0.00645f
C4944 vdd.n2100 gnd 0.00645f
C4945 vdd.n2102 gnd 0.00645f
C4946 vdd.n2103 gnd 0.00645f
C4947 vdd.n2104 gnd 0.00645f
C4948 vdd.n2105 gnd 0.00645f
C4949 vdd.n2106 gnd 0.00645f
C4950 vdd.n2108 gnd 0.00645f
C4951 vdd.n2110 gnd 0.00645f
C4952 vdd.n2111 gnd 0.00645f
C4953 vdd.n2112 gnd 0.00645f
C4954 vdd.n2113 gnd 0.00645f
C4955 vdd.n2114 gnd 0.00645f
C4956 vdd.n2116 gnd 0.00645f
C4957 vdd.n2118 gnd 0.00645f
C4958 vdd.n2119 gnd 0.00645f
C4959 vdd.n2120 gnd 0.00645f
C4960 vdd.n2121 gnd 0.00645f
C4961 vdd.n2122 gnd 0.00645f
C4962 vdd.n2124 gnd 0.00645f
C4963 vdd.n2126 gnd 0.00645f
C4964 vdd.n2127 gnd 0.00645f
C4965 vdd.n2128 gnd 0.00645f
C4966 vdd.n2129 gnd 0.00645f
C4967 vdd.n2130 gnd 0.00645f
C4968 vdd.n2132 gnd 0.00645f
C4969 vdd.n2134 gnd 0.00645f
C4970 vdd.n2135 gnd 0.00645f
C4971 vdd.n2136 gnd 0.015081f
C4972 vdd.n2137 gnd 0.014326f
C4973 vdd.n2138 gnd 0.014326f
C4974 vdd.n2139 gnd 0.715516f
C4975 vdd.n2140 gnd 0.014326f
C4976 vdd.n2141 gnd 0.014326f
C4977 vdd.n2142 gnd 0.00645f
C4978 vdd.n2143 gnd 0.00645f
C4979 vdd.n2144 gnd 0.00645f
C4980 vdd.n2145 gnd 0.357758f
C4981 vdd.n2146 gnd 0.00645f
C4982 vdd.n2147 gnd 0.00645f
C4983 vdd.n2148 gnd 0.00645f
C4984 vdd.n2149 gnd 0.00645f
C4985 vdd.n2150 gnd 0.00645f
C4986 vdd.n2151 gnd 0.490966f
C4987 vdd.n2152 gnd 0.00645f
C4988 vdd.n2153 gnd 0.00645f
C4989 vdd.n2154 gnd 0.00645f
C4990 vdd.n2155 gnd 0.00645f
C4991 vdd.n2156 gnd 0.00645f
C4992 vdd.n2157 gnd 0.380594f
C4993 vdd.n2158 gnd 0.00645f
C4994 vdd.n2159 gnd 0.00645f
C4995 vdd.n2160 gnd 0.00645f
C4996 vdd.n2161 gnd 0.00645f
C4997 vdd.n2162 gnd 0.00645f
C4998 vdd.n2163 gnd 0.517608f
C4999 vdd.n2164 gnd 0.00645f
C5000 vdd.n2165 gnd 0.00645f
C5001 vdd.n2166 gnd 0.00645f
C5002 vdd.n2167 gnd 0.00645f
C5003 vdd.n2168 gnd 0.00645f
C5004 vdd.n2169 gnd 0.201715f
C5005 vdd.n2170 gnd 0.00645f
C5006 vdd.n2171 gnd 0.00645f
C5007 vdd.n2172 gnd 0.00645f
C5008 vdd.n2173 gnd 0.00645f
C5009 vdd.n2174 gnd 0.00645f
C5010 vdd.n2175 gnd 0.517608f
C5011 vdd.n2176 gnd 0.00645f
C5012 vdd.n2177 gnd 0.00645f
C5013 vdd.n2178 gnd 0.00645f
C5014 vdd.n2179 gnd 0.00645f
C5015 vdd.n2180 gnd 0.00645f
C5016 vdd.n2181 gnd 0.293057f
C5017 vdd.n2182 gnd 0.00645f
C5018 vdd.n2183 gnd 0.00645f
C5019 vdd.n2184 gnd 0.00645f
C5020 vdd.n2185 gnd 0.00645f
C5021 vdd.n2186 gnd 0.00645f
C5022 vdd.n2187 gnd 0.395818f
C5023 vdd.n2188 gnd 0.00645f
C5024 vdd.n2189 gnd 0.00645f
C5025 vdd.n2190 gnd 0.00645f
C5026 vdd.n2191 gnd 0.00645f
C5027 vdd.n2192 gnd 0.00645f
C5028 vdd.n2193 gnd 0.270222f
C5029 vdd.n2194 gnd 0.00645f
C5030 vdd.n2195 gnd 0.00645f
C5031 vdd.n2196 gnd 0.00645f
C5032 vdd.n2197 gnd 0.00645f
C5033 vdd.n2198 gnd 0.00645f
C5034 vdd.n2199 gnd 0.418653f
C5035 vdd.n2200 gnd 0.00645f
C5036 vdd.n2201 gnd 0.00645f
C5037 vdd.n2202 gnd 0.00645f
C5038 vdd.n2203 gnd 0.00645f
C5039 vdd.n2204 gnd 0.00645f
C5040 vdd.n2205 gnd 0.270222f
C5041 vdd.n2206 gnd 0.00645f
C5042 vdd.n2207 gnd 0.00645f
C5043 vdd.n2208 gnd 0.00645f
C5044 vdd.n2209 gnd 0.00645f
C5045 vdd.n2210 gnd 0.00645f
C5046 vdd.n2211 gnd 0.441489f
C5047 vdd.n2212 gnd 0.00645f
C5048 vdd.n2213 gnd 0.00645f
C5049 vdd.n2214 gnd 0.00645f
C5050 vdd.n2215 gnd 0.00645f
C5051 vdd.n2216 gnd 0.00645f
C5052 vdd.n2217 gnd 0.293057f
C5053 vdd.n2218 gnd 0.00645f
C5054 vdd.n2219 gnd 0.00645f
C5055 vdd.n2220 gnd 0.00645f
C5056 vdd.n2221 gnd 0.00645f
C5057 vdd.n2222 gnd 0.00645f
C5058 vdd.n2223 gnd 0.464324f
C5059 vdd.n2224 gnd 0.00645f
C5060 vdd.n2225 gnd 0.00645f
C5061 vdd.n2226 gnd 0.00645f
C5062 vdd.n2227 gnd 0.00645f
C5063 vdd.n2228 gnd 0.00645f
C5064 vdd.n2229 gnd 0.315893f
C5065 vdd.n2230 gnd 0.00645f
C5066 vdd.n2231 gnd 0.00645f
C5067 vdd.n2232 gnd 0.00645f
C5068 vdd.n2233 gnd 0.00645f
C5069 vdd.n2234 gnd 0.00645f
C5070 vdd.n2235 gnd 0.517608f
C5071 vdd.n2236 gnd 0.00645f
C5072 vdd.n2237 gnd 0.00645f
C5073 vdd.n2238 gnd 0.00645f
C5074 vdd.n2239 gnd 0.00645f
C5075 vdd.n2240 gnd 0.00645f
C5076 vdd.n2241 gnd 0.342534f
C5077 vdd.n2242 gnd 0.00645f
C5078 vdd.n2243 gnd 0.004269f
C5079 vdd.n2244 gnd 0.018686f
C5080 vdd.n2245 gnd 0.005407f
C5081 vdd.n2246 gnd 0.00645f
C5082 vdd.n2247 gnd 0.00645f
C5083 vdd.n2248 gnd 0.00645f
C5084 vdd.n2249 gnd 0.00645f
C5085 vdd.n2251 gnd 0.00645f
C5086 vdd.n2252 gnd 0.00645f
C5087 vdd.n2254 gnd 0.00645f
C5088 vdd.n2255 gnd 0.00645f
C5089 vdd.n2256 gnd 0.00645f
C5090 vdd.n2258 gnd 0.00645f
C5091 vdd.n2259 gnd 0.00645f
C5092 vdd.n2260 gnd 0.00645f
C5093 vdd.n2261 gnd 0.00645f
C5094 vdd.n2262 gnd 0.00645f
C5095 vdd.n2263 gnd 0.00645f
C5096 vdd.n2265 gnd 0.00645f
C5097 vdd.n2266 gnd 0.00645f
C5098 vdd.n2267 gnd 0.00645f
C5099 vdd.n2268 gnd 0.00645f
C5100 vdd.n2269 gnd 0.00645f
C5101 vdd.n2270 gnd 0.00645f
C5102 vdd.n2272 gnd 0.00645f
C5103 vdd.n2273 gnd 0.00645f
C5104 vdd.n2275 gnd 0.015081f
C5105 vdd.n2276 gnd 0.015081f
C5106 vdd.n2277 gnd 0.014326f
C5107 vdd.n2278 gnd 0.00645f
C5108 vdd.n2279 gnd 0.00645f
C5109 vdd.n2280 gnd 0.00645f
C5110 vdd.n2281 gnd 0.00645f
C5111 vdd.n2282 gnd 0.00645f
C5112 vdd.n2283 gnd 0.00645f
C5113 vdd.n2284 gnd 0.490966f
C5114 vdd.n2285 gnd 0.00645f
C5115 vdd.n2286 gnd 0.00645f
C5116 vdd.n2287 gnd 0.00645f
C5117 vdd.n2288 gnd 0.00645f
C5118 vdd.n2289 gnd 0.00645f
C5119 vdd.n2290 gnd 0.517608f
C5120 vdd.n2291 gnd 0.00645f
C5121 vdd.n2292 gnd 0.00645f
C5122 vdd.n2293 gnd 0.00645f
C5123 vdd.n2294 gnd 0.015119f
C5124 vdd.n2295 gnd 0.014287f
C5125 vdd.n2296 gnd 0.015081f
C5126 vdd.n2298 gnd 0.00645f
C5127 vdd.n2299 gnd 0.00645f
C5128 vdd.n2300 gnd 0.004696f
C5129 vdd.n2301 gnd 0.009219f
C5130 vdd.n2302 gnd 0.00498f
C5131 vdd.n2303 gnd 0.00645f
C5132 vdd.n2304 gnd 0.00645f
C5133 vdd.n2306 gnd 0.00645f
C5134 vdd.n2307 gnd 0.00645f
C5135 vdd.n2308 gnd 0.00645f
C5136 vdd.n2309 gnd 0.00645f
C5137 vdd.n2310 gnd 0.00645f
C5138 vdd.n2311 gnd 0.00645f
C5139 vdd.n2313 gnd 0.00645f
C5140 vdd.n2314 gnd 0.00645f
C5141 vdd.n2315 gnd 0.00645f
C5142 vdd.n2316 gnd 0.00645f
C5143 vdd.n2317 gnd 0.004838f
C5144 vdd.n2318 gnd 0.00645f
C5145 vdd.n2320 gnd 0.00645f
C5146 vdd.n2321 gnd 0.004838f
C5147 vdd.n2322 gnd 0.00645f
C5148 vdd.n2323 gnd 0.00645f
C5149 vdd.n2325 gnd 0.00645f
C5150 vdd.n2326 gnd 0.00645f
C5151 vdd.n2327 gnd 0.00645f
C5152 vdd.n2328 gnd 0.00645f
C5153 vdd.n2329 gnd 0.00645f
C5154 vdd.n2330 gnd 0.00645f
C5155 vdd.n2332 gnd 0.00645f
C5156 vdd.n2333 gnd 0.00645f
C5157 vdd.n2334 gnd 0.00645f
C5158 vdd.n2335 gnd 0.00645f
C5159 vdd.n2336 gnd 0.00645f
C5160 vdd.n2337 gnd 0.00645f
C5161 vdd.n2339 gnd 0.00645f
C5162 vdd.n2340 gnd 0.00645f
C5163 vdd.n2341 gnd 0.00645f
C5164 vdd.n2342 gnd 0.015081f
C5165 vdd.n2343 gnd 0.014326f
C5166 vdd.n2344 gnd 0.014326f
C5167 vdd.n2345 gnd 0.715516f
C5168 vdd.n2346 gnd 0.014326f
C5169 vdd.n2347 gnd 0.015081f
C5170 vdd.n2348 gnd 0.014287f
C5171 vdd.n2349 gnd 0.00645f
C5172 vdd.n2350 gnd 0.004696f
C5173 vdd.n2351 gnd 0.00645f
C5174 vdd.n2353 gnd 0.00645f
C5175 vdd.n2354 gnd 0.00645f
C5176 vdd.n2355 gnd 0.00645f
C5177 vdd.n2356 gnd 0.00645f
C5178 vdd.n2357 gnd 0.00645f
C5179 vdd.n2358 gnd 0.00645f
C5180 vdd.n2360 gnd 0.00645f
C5181 vdd.n2361 gnd 0.00645f
C5182 vdd.n2362 gnd 0.00645f
C5183 vdd.n2363 gnd 0.00645f
C5184 vdd.n2364 gnd 0.00645f
C5185 vdd.n2365 gnd 0.00645f
C5186 vdd.n2367 gnd 0.00645f
C5187 vdd.n2368 gnd 0.00645f
C5188 vdd.n2369 gnd 0.004838f
C5189 vdd.n2370 gnd 0.008999f
C5190 vdd.n2371 gnd 0.009486f
C5191 vdd.n2372 gnd 0.009486f
C5192 vdd.n2373 gnd 0.007635f
C5193 vdd.n2374 gnd 0.009486f
C5194 vdd.n2375 gnd 0.009486f
C5195 vdd.n2376 gnd 0.009486f
C5196 vdd.n2377 gnd 0.009486f
C5197 vdd.n2378 gnd 0.021375f
C5198 vdd.n2379 gnd 0.003627f
C5199 vdd.t37 gnd 0.194308f
C5200 vdd.t38 gnd 0.203627f
C5201 vdd.t35 gnd 0.283884f
C5202 vdd.n2380 gnd 0.096222f
C5203 vdd.n2381 gnd 0.055169f
C5204 vdd.n2382 gnd 0.011796f
C5205 vdd.n2383 gnd 0.009486f
C5206 vdd.n2384 gnd 0.004008f
C5207 vdd.n2385 gnd 0.007635f
C5208 vdd.n2386 gnd 0.009486f
C5209 vdd.n2387 gnd 0.009486f
C5210 vdd.n2388 gnd 0.007635f
C5211 vdd.n2389 gnd 0.009486f
C5212 vdd.n2390 gnd 0.007635f
C5213 vdd.n2391 gnd 0.007635f
C5214 vdd.n2393 gnd 0.484834f
C5215 vdd.n2395 gnd 0.007635f
C5216 vdd.n2396 gnd 0.009486f
C5217 vdd.n2397 gnd 0.009486f
C5218 vdd.n2398 gnd 0.007635f
C5219 vdd.n2399 gnd 0.007635f
C5220 vdd.n2400 gnd 0.009486f
C5221 vdd.n2401 gnd 0.009486f
C5222 vdd.n2402 gnd 0.007635f
C5223 vdd.n2403 gnd 0.007635f
C5224 vdd.n2404 gnd 0.009486f
C5225 vdd.n2405 gnd 0.009486f
C5226 vdd.n2406 gnd 0.007635f
C5227 vdd.n2407 gnd 0.007635f
C5228 vdd.n2408 gnd 0.009486f
C5229 vdd.n2409 gnd 0.009486f
C5230 vdd.n2410 gnd 0.007635f
C5231 vdd.n2411 gnd 0.007635f
C5232 vdd.n2412 gnd 0.009486f
C5233 vdd.n2413 gnd 0.009486f
C5234 vdd.n2414 gnd 0.007635f
C5235 vdd.n2415 gnd 0.009486f
C5236 vdd.n2416 gnd 0.009486f
C5237 vdd.n2417 gnd 0.007635f
C5238 vdd.n2418 gnd 0.009486f
C5239 vdd.n2419 gnd 0.009486f
C5240 vdd.n2420 gnd 0.009486f
C5241 vdd.n2421 gnd 0.015614f
C5242 vdd.n2422 gnd 0.009486f
C5243 vdd.n2423 gnd 0.009486f
C5244 vdd.n2424 gnd 0.005192f
C5245 vdd.n2425 gnd 0.007635f
C5246 vdd.n2426 gnd 0.009486f
C5247 vdd.n2427 gnd 0.009486f
C5248 vdd.n2428 gnd 0.007635f
C5249 vdd.n2429 gnd 0.007635f
C5250 vdd.n2430 gnd 0.009486f
C5251 vdd.n2431 gnd 0.009486f
C5252 vdd.n2432 gnd 0.007635f
C5253 vdd.n2433 gnd 0.007635f
C5254 vdd.n2434 gnd 0.009486f
C5255 vdd.n2435 gnd 0.009486f
C5256 vdd.n2436 gnd 0.007635f
C5257 vdd.n2437 gnd 0.007635f
C5258 vdd.n2438 gnd 0.009486f
C5259 vdd.n2439 gnd 0.009486f
C5260 vdd.n2440 gnd 0.007635f
C5261 vdd.n2441 gnd 0.007635f
C5262 vdd.n2442 gnd 0.009486f
C5263 vdd.n2443 gnd 0.009486f
C5264 vdd.n2444 gnd 0.007635f
C5265 vdd.n2445 gnd 0.007635f
C5266 vdd.n2446 gnd 0.009486f
C5267 vdd.n2447 gnd 0.009486f
C5268 vdd.n2448 gnd 0.007635f
C5269 vdd.n2449 gnd 0.007635f
C5270 vdd.n2450 gnd 0.009486f
C5271 vdd.n2451 gnd 0.009486f
C5272 vdd.n2452 gnd 0.007635f
C5273 vdd.n2453 gnd 0.007635f
C5274 vdd.n2454 gnd 0.009486f
C5275 vdd.n2455 gnd 0.009486f
C5276 vdd.n2456 gnd 0.007635f
C5277 vdd.n2457 gnd 0.009486f
C5278 vdd.n2458 gnd 0.009486f
C5279 vdd.n2459 gnd 0.007635f
C5280 vdd.n2460 gnd 0.009486f
C5281 vdd.n2461 gnd 0.009486f
C5282 vdd.n2462 gnd 0.009486f
C5283 vdd.t51 gnd 0.194308f
C5284 vdd.t52 gnd 0.203627f
C5285 vdd.t50 gnd 0.283884f
C5286 vdd.n2463 gnd 0.096222f
C5287 vdd.n2464 gnd 0.055169f
C5288 vdd.n2465 gnd 0.015614f
C5289 vdd.n2466 gnd 0.009486f
C5290 vdd.n2467 gnd 0.009486f
C5291 vdd.n2468 gnd 0.006375f
C5292 vdd.n2469 gnd 0.007635f
C5293 vdd.n2470 gnd 0.009486f
C5294 vdd.n2471 gnd 0.009486f
C5295 vdd.n2472 gnd 0.007635f
C5296 vdd.n2473 gnd 0.007635f
C5297 vdd.n2474 gnd 0.009486f
C5298 vdd.n2475 gnd 0.009486f
C5299 vdd.n2476 gnd 0.007635f
C5300 vdd.n2477 gnd 0.007635f
C5301 vdd.n2478 gnd 0.009486f
C5302 vdd.n2479 gnd 0.009486f
C5303 vdd.n2480 gnd 0.007635f
C5304 vdd.n2481 gnd 0.009486f
C5305 vdd.n2482 gnd 0.007635f
C5306 vdd.n2483 gnd 0.007635f
C5307 vdd.n2485 gnd 0.484834f
C5308 vdd.n2487 gnd 0.007635f
C5309 vdd.n2488 gnd 0.009486f
C5310 vdd.n2489 gnd 0.009486f
C5311 vdd.n2490 gnd 0.007635f
C5312 vdd.n2491 gnd 0.007635f
C5313 vdd.n2492 gnd 0.007635f
C5314 vdd.n2493 gnd 0.009486f
C5315 vdd.n2494 gnd 4.59377f
C5316 vdd.n2496 gnd 0.021375f
C5317 vdd.n2497 gnd 0.006337f
C5318 vdd.n2498 gnd 0.021375f
C5319 vdd.n2499 gnd 0.021312f
C5320 vdd.n2500 gnd 0.009486f
C5321 vdd.n2501 gnd 0.007635f
C5322 vdd.n2502 gnd 0.009486f
C5323 vdd.n2503 gnd 0.643204f
C5324 vdd.n2504 gnd 0.009486f
C5325 vdd.n2505 gnd 0.007635f
C5326 vdd.n2506 gnd 0.009486f
C5327 vdd.n2507 gnd 0.009486f
C5328 vdd.n2508 gnd 0.009486f
C5329 vdd.n2509 gnd 0.007635f
C5330 vdd.n2510 gnd 0.009486f
C5331 vdd.n2511 gnd 0.761188f
C5332 vdd.n2512 gnd 0.009486f
C5333 vdd.n2513 gnd 0.007635f
C5334 vdd.n2514 gnd 0.009486f
C5335 vdd.n2515 gnd 0.009486f
C5336 vdd.n2516 gnd 0.009486f
C5337 vdd.n2517 gnd 0.007635f
C5338 vdd.n2518 gnd 0.009486f
C5339 vdd.n2519 gnd 0.761188f
C5340 vdd.n2520 gnd 0.009486f
C5341 vdd.n2521 gnd 0.007635f
C5342 vdd.n2522 gnd 0.009486f
C5343 vdd.n2523 gnd 0.009486f
C5344 vdd.n2524 gnd 0.009486f
C5345 vdd.n2525 gnd 0.007635f
C5346 vdd.n2526 gnd 0.009486f
C5347 vdd.n2527 gnd 0.559473f
C5348 vdd.n2528 gnd 0.009486f
C5349 vdd.n2529 gnd 0.007635f
C5350 vdd.n2530 gnd 0.009486f
C5351 vdd.n2531 gnd 0.009486f
C5352 vdd.n2532 gnd 0.009486f
C5353 vdd.n2533 gnd 0.007635f
C5354 vdd.n2534 gnd 0.009486f
C5355 vdd.n2535 gnd 0.452907f
C5356 vdd.n2536 gnd 0.009486f
C5357 vdd.n2537 gnd 0.007635f
C5358 vdd.n2538 gnd 0.009486f
C5359 vdd.n2539 gnd 0.009486f
C5360 vdd.n2540 gnd 0.009486f
C5361 vdd.n2541 gnd 0.007635f
C5362 vdd.n2542 gnd 0.009486f
C5363 vdd.t23 gnd 0.380594f
C5364 vdd.n2543 gnd 0.704099f
C5365 vdd.n2544 gnd 0.009486f
C5366 vdd.n2545 gnd 0.007635f
C5367 vdd.n2546 gnd 0.009486f
C5368 vdd.n2547 gnd 0.009486f
C5369 vdd.n2548 gnd 0.009486f
C5370 vdd.n2549 gnd 0.007635f
C5371 vdd.n2550 gnd 0.009486f
C5372 vdd.n2551 gnd 0.761188f
C5373 vdd.n2552 gnd 0.009486f
C5374 vdd.n2553 gnd 0.007635f
C5375 vdd.n2554 gnd 0.009486f
C5376 vdd.n2555 gnd 0.009486f
C5377 vdd.n2556 gnd 0.009486f
C5378 vdd.n2557 gnd 0.007635f
C5379 vdd.n2558 gnd 0.009486f
C5380 vdd.n2559 gnd 0.567085f
C5381 vdd.n2560 gnd 0.009486f
C5382 vdd.n2561 gnd 0.007635f
C5383 vdd.n2562 gnd 0.009486f
C5384 vdd.n2563 gnd 0.009486f
C5385 vdd.n2564 gnd 0.009486f
C5386 vdd.n2565 gnd 0.007635f
C5387 vdd.n2566 gnd 0.009486f
C5388 vdd.n2567 gnd 0.445295f
C5389 vdd.n2568 gnd 0.009486f
C5390 vdd.n2569 gnd 0.007635f
C5391 vdd.n2570 gnd 0.009486f
C5392 vdd.n2571 gnd 0.009486f
C5393 vdd.n2572 gnd 0.009486f
C5394 vdd.n2573 gnd 0.007635f
C5395 vdd.n2574 gnd 0.007635f
C5396 vdd.n2575 gnd 0.007635f
C5397 vdd.n2576 gnd 0.009486f
C5398 vdd.n2577 gnd 0.009486f
C5399 vdd.n2578 gnd 0.009486f
C5400 vdd.n2579 gnd 0.007635f
C5401 vdd.n2580 gnd 0.007635f
C5402 vdd.n2581 gnd 0.007635f
C5403 vdd.n2582 gnd 0.009486f
C5404 vdd.n2583 gnd 0.009486f
C5405 vdd.n2584 gnd 0.009486f
C5406 vdd.n2585 gnd 0.007635f
C5407 vdd.n2586 gnd 0.007635f
C5408 vdd.n2587 gnd 0.007635f
C5409 vdd.n2588 gnd 0.009486f
C5410 vdd.n2589 gnd 0.009486f
C5411 vdd.n2590 gnd 0.009486f
C5412 vdd.n2591 gnd 0.007635f
C5413 vdd.n2592 gnd 0.007635f
C5414 vdd.n2593 gnd 0.007635f
C5415 vdd.n2594 gnd 0.009486f
C5416 vdd.n2595 gnd 0.009486f
C5417 vdd.n2596 gnd 0.009486f
C5418 vdd.n2597 gnd 0.007635f
C5419 vdd.n2598 gnd 0.007635f
C5420 vdd.n2599 gnd 0.006337f
C5421 vdd.n2600 gnd 0.021312f
C5422 vdd.n2601 gnd 0.021375f
C5423 vdd.n2602 gnd 0.003627f
C5424 vdd.n2603 gnd 0.021375f
C5425 vdd.n2605 gnd 0.009486f
C5426 vdd.n2606 gnd 0.009486f
C5427 vdd.n2607 gnd 0.007635f
C5428 vdd.n2608 gnd 0.007635f
C5429 vdd.n2609 gnd 0.007635f
C5430 vdd.n2610 gnd 0.009486f
C5431 vdd.n2612 gnd 0.009486f
C5432 vdd.n2613 gnd 0.009486f
C5433 vdd.n2614 gnd 0.007635f
C5434 vdd.n2615 gnd 0.007635f
C5435 vdd.n2616 gnd 0.007635f
C5436 vdd.n2617 gnd 0.009486f
C5437 vdd.n2619 gnd 0.009486f
C5438 vdd.n2620 gnd 0.009486f
C5439 vdd.n2621 gnd 0.007635f
C5440 vdd.n2622 gnd 0.007635f
C5441 vdd.n2623 gnd 0.007635f
C5442 vdd.n2624 gnd 0.009486f
C5443 vdd.n2626 gnd 0.009486f
C5444 vdd.n2627 gnd 0.009486f
C5445 vdd.n2628 gnd 0.007635f
C5446 vdd.n2629 gnd 0.007635f
C5447 vdd.n2630 gnd 0.007635f
C5448 vdd.n2631 gnd 0.009486f
C5449 vdd.n2633 gnd 0.009486f
C5450 vdd.n2634 gnd 0.009486f
C5451 vdd.n2635 gnd 0.007635f
C5452 vdd.n2636 gnd 0.009486f
C5453 vdd.n2637 gnd 0.009486f
C5454 vdd.n2638 gnd 0.009486f
C5455 vdd.n2639 gnd 0.015614f
C5456 vdd.n2640 gnd 0.009486f
C5457 vdd.n2642 gnd 0.009486f
C5458 vdd.n2643 gnd 0.009486f
C5459 vdd.n2644 gnd 0.007635f
C5460 vdd.n2645 gnd 0.007635f
C5461 vdd.n2646 gnd 0.007635f
C5462 vdd.n2647 gnd 0.009486f
C5463 vdd.n2649 gnd 0.009486f
C5464 vdd.n2650 gnd 0.009486f
C5465 vdd.n2651 gnd 0.007635f
C5466 vdd.n2652 gnd 0.007635f
C5467 vdd.n2653 gnd 0.007635f
C5468 vdd.n2654 gnd 0.009486f
C5469 vdd.n2656 gnd 0.009486f
C5470 vdd.n2657 gnd 0.009486f
C5471 vdd.n2658 gnd 0.007635f
C5472 vdd.n2659 gnd 0.007635f
C5473 vdd.n2660 gnd 0.007635f
C5474 vdd.n2661 gnd 0.009486f
C5475 vdd.n2663 gnd 0.009486f
C5476 vdd.n2664 gnd 0.009486f
C5477 vdd.n2665 gnd 0.007635f
C5478 vdd.n2666 gnd 0.007635f
C5479 vdd.n2667 gnd 0.007635f
C5480 vdd.n2668 gnd 0.009486f
C5481 vdd.n2670 gnd 0.009486f
C5482 vdd.n2671 gnd 0.009486f
C5483 vdd.n2672 gnd 0.007635f
C5484 vdd.n2673 gnd 0.009486f
C5485 vdd.n2674 gnd 0.009486f
C5486 vdd.n2675 gnd 0.009486f
C5487 vdd.n2676 gnd 0.015614f
C5488 vdd.n2677 gnd 0.009486f
C5489 vdd.n2679 gnd 0.009486f
C5490 vdd.n2680 gnd 0.009486f
C5491 vdd.n2681 gnd 0.007635f
C5492 vdd.n2682 gnd 0.007635f
C5493 vdd.n2683 gnd 0.007635f
C5494 vdd.n2684 gnd 0.009486f
C5495 vdd.n2686 gnd 0.009486f
C5496 vdd.n2687 gnd 0.009486f
C5497 vdd.n2688 gnd 0.007635f
C5498 vdd.n2689 gnd 0.007635f
C5499 vdd.n2690 gnd 0.007635f
C5500 vdd.n2691 gnd 0.009486f
C5501 vdd.n2693 gnd 0.009486f
C5502 vdd.n2694 gnd 0.009486f
C5503 vdd.n2695 gnd 0.007635f
C5504 vdd.n2696 gnd 0.007635f
C5505 vdd.n2697 gnd 0.007635f
C5506 vdd.n2698 gnd 0.009486f
C5507 vdd.n2700 gnd 0.009486f
C5508 vdd.n2701 gnd 0.009486f
C5509 vdd.n2703 gnd 0.009486f
C5510 vdd.n2704 gnd 0.007635f
C5511 vdd.n2705 gnd 0.007635f
C5512 vdd.n2706 gnd 0.006337f
C5513 vdd.n2707 gnd 0.021375f
C5514 vdd.n2708 gnd 0.021312f
C5515 vdd.n2709 gnd 0.006337f
C5516 vdd.n2710 gnd 0.021312f
C5517 vdd.n2711 gnd 0.978126f
C5518 vdd.n2712 gnd 0.643204f
C5519 vdd.t28 gnd 0.380594f
C5520 vdd.n2713 gnd 0.498578f
C5521 vdd.n2714 gnd 0.009486f
C5522 vdd.n2715 gnd 0.007635f
C5523 vdd.n2716 gnd 0.007635f
C5524 vdd.n2717 gnd 0.007635f
C5525 vdd.n2718 gnd 0.009486f
C5526 vdd.n2719 gnd 0.761188f
C5527 vdd.n2720 gnd 0.761188f
C5528 vdd.n2721 gnd 0.582309f
C5529 vdd.n2722 gnd 0.009486f
C5530 vdd.n2723 gnd 0.007635f
C5531 vdd.n2724 gnd 0.007635f
C5532 vdd.n2725 gnd 0.007635f
C5533 vdd.n2726 gnd 0.009486f
C5534 vdd.n2727 gnd 0.761188f
C5535 vdd.n2728 gnd 0.452907f
C5536 vdd.t25 gnd 0.380594f
C5537 vdd.n2729 gnd 0.688875f
C5538 vdd.n2730 gnd 0.009486f
C5539 vdd.n2731 gnd 0.007635f
C5540 vdd.n2732 gnd 0.007635f
C5541 vdd.n2733 gnd 0.007635f
C5542 vdd.n2734 gnd 0.009486f
C5543 vdd.n2735 gnd 0.437683f
C5544 vdd.n2736 gnd 0.761188f
C5545 vdd.n2737 gnd 0.574697f
C5546 vdd.n2738 gnd 0.009486f
C5547 vdd.n2739 gnd 0.007635f
C5548 vdd.n2740 gnd 0.007635f
C5549 vdd.n2741 gnd 0.007635f
C5550 vdd.n2742 gnd 0.009486f
C5551 vdd.n2743 gnd 0.761188f
C5552 vdd.n2744 gnd 0.445295f
C5553 vdd.t4 gnd 0.380594f
C5554 vdd.n2745 gnd 0.696487f
C5555 vdd.n2746 gnd 0.009486f
C5556 vdd.n2747 gnd 0.007635f
C5557 vdd.n2748 gnd 0.007291f
C5558 vdd.n2749 gnd 0.2589f
C5559 vdd.n2750 gnd 1.95992f
.ends

