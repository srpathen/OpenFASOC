* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 vdd.t183 a_n5644_8799.t36 CSoutput.t91 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 a_n1986_8322.t11 a_n2848_n452.t48 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n1808_13878.t19 a_n2848_n452.t30 a_n2848_n452.t31 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X3 a_n5644_8799.t19 plus.t5 a_n3827_n3924.t23 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X4 gnd.t196 gnd.t193 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X5 outputibias.t7 outputibias.t6 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X6 a_n3827_n3924.t22 plus.t6 a_n5644_8799.t6 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X7 gnd.t192 gnd.t190 gnd.t191 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 gnd.t17 commonsourceibias.t80 CSoutput.t5 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 a_n3827_n3924.t27 diffpairibias.t20 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 commonsourceibias.t79 commonsourceibias.t78 gnd.t303 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X11 a_n2848_n452.t33 a_n2848_n452.t32 a_n1808_13878.t18 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 a_n1808_13878.t17 a_n2848_n452.t28 a_n2848_n452.t29 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 vdd.t107 vdd.t105 vdd.t106 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X14 a_n1808_13878.t7 a_n2848_n452.t49 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 gnd.t189 gnd.t187 gnd.t188 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X16 commonsourceibias.t77 commonsourceibias.t76 gnd.t333 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t68 a_n5644_8799.t37 vdd.t182 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 CSoutput.t6 commonsourceibias.t81 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t186 gnd.t184 gnd.t185 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X20 vdd.t104 vdd.t102 vdd.t103 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X21 gnd.t183 gnd.t181 gnd.t182 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X22 gnd.t225 commonsourceibias.t74 commonsourceibias.t75 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t57 commonsourceibias.t82 gnd.t301 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 a_n1986_8322.t23 a_n2848_n452.t50 a_n5644_8799.t22 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 a_n2848_n452.t5 minus.t5 a_n3827_n3924.t34 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 a_n5644_8799.t5 plus.t7 a_n3827_n3924.t21 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 commonsourceibias.t73 commonsourceibias.t72 gnd.t294 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 plus.t0 gnd.t178 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 CSoutput.t58 commonsourceibias.t83 gnd.t302 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n2848_n452.t4 minus.t6 a_n3827_n3924.t33 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 output.t19 CSoutput.t128 vdd.t16 gnd.t279 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X32 commonsourceibias.t71 commonsourceibias.t70 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 CSoutput.t67 a_n5644_8799.t38 vdd.t181 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 vdd.t180 a_n5644_8799.t39 CSoutput.t66 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n3827_n3924.t20 plus.t8 a_n5644_8799.t14 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X36 a_n5644_8799.t23 a_n2848_n452.t51 a_n1986_8322.t22 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X37 CSoutput.t65 a_n5644_8799.t40 vdd.t179 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X38 vdd.t178 a_n5644_8799.t41 CSoutput.t64 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 a_n3827_n3924.t32 minus.t7 a_n2848_n452.t3 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X40 CSoutput.t10 commonsourceibias.t84 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n3827_n3924.t54 diffpairibias.t21 gnd.t346 gnd.t345 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 gnd.t177 gnd.t175 gnd.t176 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X43 gnd.t357 commonsourceibias.t68 commonsourceibias.t69 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 gnd.t38 commonsourceibias.t85 CSoutput.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 CSoutput.t86 a_n5644_8799.t42 vdd.t177 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 vdd.t101 vdd.t99 vdd.t100 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X47 gnd.t7 commonsourceibias.t86 CSoutput.t1 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 commonsourceibias.t67 commonsourceibias.t66 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 gnd.t9 commonsourceibias.t87 CSoutput.t2 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 vdd.t15 CSoutput.t129 output.t18 gnd.t278 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X51 gnd.t331 commonsourceibias.t88 CSoutput.t62 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 gnd.t174 gnd.t172 gnd.t173 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X53 a_n3827_n3924.t19 plus.t9 a_n5644_8799.t13 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X54 gnd.t11 commonsourceibias.t64 commonsourceibias.t65 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 a_n1808_13878.t16 a_n2848_n452.t42 a_n2848_n452.t43 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X56 vdd.t176 a_n5644_8799.t43 CSoutput.t85 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 a_n3827_n3924.t18 plus.t10 a_n5644_8799.t26 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X58 a_n3827_n3924.t31 minus.t8 a_n2848_n452.t2 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X59 commonsourceibias.t63 commonsourceibias.t62 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 diffpairibias.t19 diffpairibias.t18 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 a_n2848_n452.t35 a_n2848_n452.t34 a_n1808_13878.t15 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X62 CSoutput.t84 a_n5644_8799.t44 vdd.t175 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 output.t17 CSoutput.t130 vdd.t10 gnd.t277 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X64 vdd.t98 vdd.t96 vdd.t97 vdd.t65 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X65 commonsourceibias.t61 commonsourceibias.t60 gnd.t344 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 gnd.t326 commonsourceibias.t58 commonsourceibias.t59 gnd.t292 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 diffpairibias.t17 diffpairibias.t16 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X68 gnd.t171 gnd.t168 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X69 vdd.t95 vdd.t93 vdd.t94 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X70 CSoutput.t63 commonsourceibias.t89 gnd.t332 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 vdd.t174 a_n5644_8799.t45 CSoutput.t83 vdd.t173 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 CSoutput.t42 commonsourceibias.t90 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 vdd.t172 a_n5644_8799.t46 CSoutput.t96 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t95 a_n5644_8799.t47 vdd.t171 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X75 a_n3827_n3924.t30 minus.t9 a_n2848_n452.t1 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X76 gnd.t304 commonsourceibias.t56 commonsourceibias.t57 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 CSoutput.t43 commonsourceibias.t91 gnd.t257 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 a_n3827_n3924.t17 plus.t11 a_n5644_8799.t16 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X79 CSoutput.t124 commonsourceibias.t92 gnd.t355 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t170 a_n5644_8799.t48 CSoutput.t94 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t125 commonsourceibias.t93 gnd.t356 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 a_n5644_8799.t21 plus.t12 a_n3827_n3924.t16 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X83 vdd.t18 CSoutput.t131 output.t16 gnd.t276 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X84 output.t15 CSoutput.t132 vdd.t12 gnd.t275 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X85 CSoutput.t93 a_n5644_8799.t49 vdd.t169 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 CSoutput.t92 a_n5644_8799.t50 vdd.t168 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 CSoutput.t8 commonsourceibias.t94 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 a_n3827_n3924.t24 diffpairibias.t22 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X89 CSoutput.t77 a_n5644_8799.t51 vdd.t167 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n3827_n3924.t15 plus.t13 a_n5644_8799.t29 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X91 vdd.t166 a_n5644_8799.t52 CSoutput.t76 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 gnd.t197 commonsourceibias.t54 commonsourceibias.t55 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t327 commonsourceibias.t52 commonsourceibias.t53 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 gnd.t305 commonsourceibias.t50 commonsourceibias.t51 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 a_n2848_n452.t27 a_n2848_n452.t26 a_n1808_13878.t14 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X96 output.t3 outputibias.t8 gnd.t352 gnd.t351 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X97 a_n2848_n452.t39 a_n2848_n452.t38 a_n1808_13878.t13 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t165 a_n5644_8799.t53 CSoutput.t75 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n5644_8799.t30 a_n2848_n452.t52 a_n1986_8322.t21 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 CSoutput.t133 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X101 vdd.t164 a_n5644_8799.t54 CSoutput.t74 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n2848_n452.t6 minus.t10 a_n3827_n3924.t35 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X103 gnd.t167 gnd.t164 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X104 diffpairibias.t15 diffpairibias.t14 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X105 output.t2 outputibias.t9 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X106 gnd.t31 commonsourceibias.t95 CSoutput.t9 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 gnd.t291 commonsourceibias.t96 CSoutput.t51 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t293 commonsourceibias.t97 CSoutput.t52 gnd.t292 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t222 commonsourceibias.t98 CSoutput.t26 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t92 vdd.t90 vdd.t91 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X111 gnd.t223 commonsourceibias.t99 CSoutput.t27 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 vdd.t163 a_n5644_8799.t55 CSoutput.t73 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 vdd.t89 vdd.t87 vdd.t88 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t252 commonsourceibias.t100 CSoutput.t40 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X115 gnd.t163 gnd.t161 gnd.t162 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X116 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 vdd.t13 CSoutput.t134 output.t14 gnd.t274 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X118 a_n3827_n3924.t26 diffpairibias.t23 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X119 vdd.t82 vdd.t79 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 gnd.t160 gnd.t158 minus.t4 gnd.t159 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X121 CSoutput.t41 commonsourceibias.t101 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X122 gnd.t157 gnd.t155 gnd.t156 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X123 gnd.t198 commonsourceibias.t48 commonsourceibias.t49 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t185 a_n2848_n452.t53 a_n1986_8322.t10 vdd.t184 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 vdd.t78 vdd.t76 vdd.t77 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 CSoutput.t99 a_n5644_8799.t56 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 a_n1986_8322.t9 a_n2848_n452.t54 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 gnd.t299 commonsourceibias.t102 CSoutput.t55 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 vdd.t160 a_n5644_8799.t57 CSoutput.t98 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 vdd.t117 a_n2848_n452.t55 a_n1808_13878.t6 vdd.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X131 gnd.t154 gnd.t152 plus.t3 gnd.t153 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X132 gnd.t328 commonsourceibias.t46 commonsourceibias.t47 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 a_n2848_n452.t12 minus.t11 a_n3827_n3924.t41 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X134 a_n5644_8799.t1 plus.t14 a_n3827_n3924.t14 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X135 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 a_n5644_8799.t0 plus.t15 a_n3827_n3924.t13 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 a_n2848_n452.t15 minus.t12 a_n3827_n3924.t44 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X138 CSoutput.t135 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X139 diffpairibias.t13 diffpairibias.t12 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X140 CSoutput.t56 commonsourceibias.t103 gnd.t300 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t71 vdd.t68 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 vdd.t158 a_n5644_8799.t58 CSoutput.t97 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X143 CSoutput.t53 commonsourceibias.t104 gnd.t297 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 commonsourceibias.t45 commonsourceibias.t44 gnd.t199 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 CSoutput.t54 commonsourceibias.t105 gnd.t298 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 a_n5644_8799.t31 a_n2848_n452.t56 a_n1986_8322.t20 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 a_n1986_8322.t8 a_n2848_n452.t57 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X148 vdd.t67 vdd.t64 vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X149 CSoutput.t38 commonsourceibias.t106 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 gnd.t251 commonsourceibias.t107 CSoutput.t39 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X151 a_n2848_n452.t45 a_n2848_n452.t44 a_n1808_13878.t12 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 CSoutput.t36 commonsourceibias.t108 gnd.t246 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n3827_n3924.t40 minus.t13 a_n2848_n452.t11 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X154 a_n5644_8799.t27 a_n2848_n452.t58 a_n1986_8322.t19 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 gnd.t247 commonsourceibias.t109 CSoutput.t37 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 gnd.t78 commonsourceibias.t42 commonsourceibias.t43 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 a_n1808_13878.t11 a_n2848_n452.t46 a_n2848_n452.t47 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 gnd.t244 commonsourceibias.t110 CSoutput.t34 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n3827_n3924.t12 plus.t16 a_n5644_8799.t4 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X160 a_n2848_n452.t10 minus.t14 a_n3827_n3924.t39 gnd.t64 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 commonsourceibias.t41 commonsourceibias.t40 gnd.t308 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 gnd.t208 commonsourceibias.t38 commonsourceibias.t39 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 vdd.t113 a_n2848_n452.t59 a_n1986_8322.t7 vdd.t112 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X164 gnd.t258 commonsourceibias.t36 commonsourceibias.t37 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 vdd.t63 vdd.t61 vdd.t62 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X166 a_n3827_n3924.t25 diffpairibias.t24 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X167 commonsourceibias.t35 commonsourceibias.t34 gnd.t209 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 CSoutput.t90 a_n5644_8799.t59 vdd.t156 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 a_n5644_8799.t2 plus.t17 a_n3827_n3924.t11 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X170 gnd.t245 commonsourceibias.t111 CSoutput.t35 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n3827_n3924.t46 diffpairibias.t25 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X172 vdd.t155 a_n5644_8799.t60 CSoutput.t89 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X173 gnd.t242 commonsourceibias.t112 CSoutput.t32 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 gnd.t243 commonsourceibias.t113 CSoutput.t33 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t342 commonsourceibias.t114 CSoutput.t120 gnd.t292 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 gnd.t343 commonsourceibias.t115 CSoutput.t121 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X177 a_n5644_8799.t17 plus.t18 a_n3827_n3924.t10 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X178 vdd.t154 a_n5644_8799.t61 CSoutput.t88 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 CSoutput.t118 commonsourceibias.t116 gnd.t340 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 vdd.t4 CSoutput.t136 output.t13 gnd.t273 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X181 CSoutput.t137 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X182 commonsourceibias.t33 commonsourceibias.t32 gnd.t259 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 minus.t3 gnd.t149 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X184 gnd.t341 commonsourceibias.t117 CSoutput.t119 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 CSoutput.t116 commonsourceibias.t118 gnd.t338 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X186 CSoutput.t138 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X187 CSoutput.t117 commonsourceibias.t119 gnd.t339 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 diffpairibias.t11 diffpairibias.t10 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 gnd.t148 gnd.t146 gnd.t147 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X190 gnd.t334 commonsourceibias.t120 CSoutput.t112 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n2848_n452.t9 minus.t15 a_n3827_n3924.t38 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 output.t1 outputibias.t10 gnd.t330 gnd.t329 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X193 a_n3827_n3924.t9 plus.t19 a_n5644_8799.t11 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X194 gnd.t309 commonsourceibias.t30 commonsourceibias.t31 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X195 gnd.t310 commonsourceibias.t28 commonsourceibias.t29 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t87 a_n5644_8799.t62 vdd.t153 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t115 commonsourceibias.t121 gnd.t337 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 commonsourceibias.t27 commonsourceibias.t26 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 vdd.t60 vdd.t58 vdd.t59 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 a_n1808_13878.t5 a_n2848_n452.t60 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 vdd.t189 a_n2848_n452.t61 a_n1808_13878.t4 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 diffpairibias.t9 diffpairibias.t8 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X204 a_n3827_n3924.t37 minus.t16 a_n2848_n452.t8 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X205 CSoutput.t114 commonsourceibias.t122 gnd.t336 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X206 gnd.t79 commonsourceibias.t24 commonsourceibias.t25 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias.t7 diffpairibias.t6 gnd.t348 gnd.t347 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 CSoutput.t102 a_n5644_8799.t63 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd.t286 commonsourceibias.t123 CSoutput.t46 gnd.t250 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X210 vdd.t150 a_n5644_8799.t64 CSoutput.t101 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput.t113 commonsourceibias.t124 gnd.t335 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 a_n3827_n3924.t36 minus.t17 a_n2848_n452.t7 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 a_n3827_n3924.t8 plus.t20 a_n5644_8799.t25 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X214 CSoutput.t21 commonsourceibias.t125 gnd.t84 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n1986_8322.t18 a_n2848_n452.t62 a_n5644_8799.t28 vdd.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 gnd.t76 commonsourceibias.t126 CSoutput.t17 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 a_n3827_n3924.t45 minus.t18 a_n2848_n452.t16 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X218 gnd.t145 gnd.t142 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X219 vdd.t149 a_n5644_8799.t65 CSoutput.t100 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 CSoutput.t82 a_n5644_8799.t66 vdd.t147 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 CSoutput.t20 commonsourceibias.t127 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 gnd.t74 commonsourceibias.t128 CSoutput.t16 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 vdd.t5 CSoutput.t139 output.t12 gnd.t272 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X224 gnd.t141 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X225 vdd.t146 a_n5644_8799.t67 CSoutput.t81 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 vdd.t119 a_n2848_n452.t63 a_n1986_8322.t6 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X227 CSoutput.t19 commonsourceibias.t129 gnd.t81 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 commonsourceibias.t23 commonsourceibias.t22 gnd.t311 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 gnd.t137 gnd.t134 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X230 a_n1808_13878.t3 a_n2848_n452.t64 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X231 gnd.t133 gnd.t131 gnd.t132 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X232 minus.t2 gnd.t128 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X233 a_n3827_n3924.t28 diffpairibias.t26 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 CSoutput.t80 a_n5644_8799.t68 vdd.t145 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 a_n5644_8799.t24 plus.t21 a_n3827_n3924.t7 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X236 a_n2848_n452.t19 minus.t19 a_n3827_n3924.t49 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X237 gnd.t72 commonsourceibias.t130 CSoutput.t15 gnd.t71 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 CSoutput.t79 a_n5644_8799.t69 vdd.t144 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X239 a_n3827_n3924.t48 minus.t20 a_n2848_n452.t18 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X240 vdd.t53 vdd.t51 vdd.t52 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X241 CSoutput.t47 commonsourceibias.t131 gnd.t287 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 gnd.t288 commonsourceibias.t132 CSoutput.t48 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 a_n1986_8322.t17 a_n2848_n452.t65 a_n5644_8799.t32 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X244 vdd.t195 a_n2848_n452.t66 a_n1986_8322.t5 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 vdd.t143 a_n5644_8799.t70 CSoutput.t78 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 CSoutput.t71 a_n5644_8799.t71 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 a_n3827_n3924.t47 minus.t21 a_n2848_n452.t17 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X248 CSoutput.t44 commonsourceibias.t133 gnd.t284 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 gnd.t325 commonsourceibias.t134 CSoutput.t61 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 a_n3827_n3924.t53 minus.t22 a_n2848_n452.t23 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X251 gnd.t324 commonsourceibias.t135 CSoutput.t60 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 CSoutput.t59 commonsourceibias.t136 gnd.t323 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 diffpairibias.t5 diffpairibias.t4 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X254 vdd.t50 vdd.t47 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X255 gnd.t354 commonsourceibias.t137 CSoutput.t123 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X256 output.t11 CSoutput.t140 vdd.t3 gnd.t271 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X257 commonsourceibias.t21 commonsourceibias.t20 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 vdd.t46 vdd.t43 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X259 CSoutput.t127 commonsourceibias.t138 gnd.t363 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 gnd.t260 commonsourceibias.t18 commonsourceibias.t19 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 a_n1808_13878.t10 a_n2848_n452.t24 a_n2848_n452.t25 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X262 CSoutput.t50 commonsourceibias.t139 gnd.t290 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 a_n3827_n3924.t57 diffpairibias.t27 gnd.t361 gnd.t360 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X264 a_n1986_8322.t16 a_n2848_n452.t67 a_n5644_8799.t33 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X265 CSoutput.t141 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X266 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X267 a_n3827_n3924.t29 minus.t23 a_n2848_n452.t0 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X268 CSoutput.t45 commonsourceibias.t140 gnd.t285 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X269 output.t0 outputibias.t11 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X270 gnd.t312 commonsourceibias.t16 commonsourceibias.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 CSoutput.t70 a_n5644_8799.t72 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X272 a_n1986_8322.t4 a_n2848_n452.t68 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X273 gnd.t241 commonsourceibias.t141 CSoutput.t31 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 CSoutput.t14 commonsourceibias.t142 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd.t123 gnd.t121 plus.t4 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X276 gnd.t120 gnd.t117 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X277 output.t10 CSoutput.t142 vdd.t14 gnd.t270 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X278 CSoutput.t30 commonsourceibias.t143 gnd.t240 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 vdd.t199 a_n2848_n452.t69 a_n1808_13878.t2 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X280 CSoutput.t25 commonsourceibias.t144 gnd.t206 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 commonsourceibias.t15 commonsourceibias.t14 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 commonsourceibias.t13 commonsourceibias.t12 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X283 CSoutput.t4 commonsourceibias.t145 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 gnd.t68 commonsourceibias.t146 CSoutput.t13 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 gnd.t215 commonsourceibias.t10 commonsourceibias.t11 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 vdd.t42 vdd.t39 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X287 vdd.t9 CSoutput.t143 output.t9 gnd.t269 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X288 output.t8 CSoutput.t144 vdd.t8 gnd.t268 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X289 a_n1986_8322.t15 a_n2848_n452.t70 a_n5644_8799.t34 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X290 gnd.t116 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X291 a_n3827_n3924.t6 plus.t22 a_n5644_8799.t3 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X292 vdd.t38 vdd.t36 vdd.t37 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X293 a_n5644_8799.t35 a_n2848_n452.t71 a_n1986_8322.t14 vdd.t110 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X294 a_n1808_13878.t1 a_n2848_n452.t72 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X295 vdd.t138 a_n5644_8799.t73 CSoutput.t69 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t105 a_n5644_8799.t74 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 gnd.t112 gnd.t110 minus.t1 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X298 a_n2848_n452.t14 minus.t24 a_n3827_n3924.t43 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X299 a_n5644_8799.t15 plus.t23 a_n3827_n3924.t5 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X300 commonsourceibias.t9 commonsourceibias.t8 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 a_n2848_n452.t13 minus.t25 a_n3827_n3924.t42 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X302 gnd.t263 commonsourceibias.t6 commonsourceibias.t7 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 CSoutput.t24 commonsourceibias.t147 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 commonsourceibias.t5 commonsourceibias.t4 gnd.t313 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 gnd.t27 commonsourceibias.t148 CSoutput.t7 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 CSoutput.t145 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X307 gnd.t80 commonsourceibias.t149 CSoutput.t18 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 CSoutput.t104 a_n5644_8799.t75 vdd.t134 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 a_n1808_13878.t9 a_n2848_n452.t36 a_n2848_n452.t37 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 a_n3827_n3924.t50 minus.t26 a_n2848_n452.t20 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X311 a_n3827_n3924.t55 diffpairibias.t28 gnd.t350 gnd.t349 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X312 gnd.t66 commonsourceibias.t150 CSoutput.t12 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X314 output.t7 CSoutput.t146 vdd.t7 gnd.t267 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 gnd.t13 commonsourceibias.t151 CSoutput.t3 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 a_n5644_8799.t7 plus.t24 a_n3827_n3924.t4 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X317 CSoutput.t103 a_n5644_8799.t76 vdd.t133 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t22 commonsourceibias.t152 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 CSoutput.t0 commonsourceibias.t153 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 commonsourceibias.t3 commonsourceibias.t2 gnd.t314 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 gnd.t105 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X322 vdd.t132 a_n5644_8799.t77 CSoutput.t108 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 output.t6 CSoutput.t147 vdd.t6 gnd.t266 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X324 outputibias.t5 outputibias.t4 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X325 diffpairibias.t3 diffpairibias.t2 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X326 a_n5644_8799.t12 a_n2848_n452.t73 a_n1986_8322.t13 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X327 a_n2848_n452.t41 a_n2848_n452.t40 a_n1808_13878.t8 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X328 gnd.t101 gnd.t99 plus.t2 gnd.t100 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X329 a_n2848_n452.t22 minus.t27 a_n3827_n3924.t52 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X330 vdd.t131 a_n5644_8799.t78 CSoutput.t107 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 outputibias.t3 outputibias.t2 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X332 vdd.t35 vdd.t32 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X333 diffpairibias.t1 diffpairibias.t0 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X334 gnd.t353 commonsourceibias.t154 CSoutput.t122 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 outputibias.t1 outputibias.t0 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X336 CSoutput.t126 commonsourceibias.t155 gnd.t362 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 plus.t1 gnd.t96 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X338 CSoutput.t49 commonsourceibias.t156 gnd.t289 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 gnd.t95 gnd.t93 minus.t0 gnd.t94 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X340 gnd.t92 gnd.t89 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X341 a_n5644_8799.t9 plus.t25 a_n3827_n3924.t3 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X342 gnd.t239 commonsourceibias.t157 CSoutput.t29 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 vdd.t17 CSoutput.t148 output.t5 gnd.t265 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X344 vdd.t20 a_n2848_n452.t74 a_n1808_13878.t0 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X345 CSoutput.t106 a_n5644_8799.t79 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 a_n5644_8799.t20 plus.t26 a_n3827_n3924.t2 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X347 a_n2848_n452.t21 minus.t28 a_n3827_n3924.t51 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X348 gnd.t238 commonsourceibias.t158 CSoutput.t28 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 CSoutput.t111 a_n5644_8799.t80 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 gnd.t203 commonsourceibias.t159 CSoutput.t23 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 vdd.t11 CSoutput.t149 output.t4 gnd.t264 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X352 vdd.t125 a_n5644_8799.t81 CSoutput.t110 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 a_n1986_8322.t12 a_n2848_n452.t75 a_n5644_8799.t10 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X354 a_n3827_n3924.t1 plus.t27 a_n5644_8799.t8 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X355 commonsourceibias.t1 commonsourceibias.t0 gnd.t218 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 vdd.t123 a_n5644_8799.t82 CSoutput.t109 vdd.t122 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X357 CSoutput.t72 a_n5644_8799.t83 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X358 a_n3827_n3924.t0 plus.t28 a_n5644_8799.t18 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X359 a_n3827_n3924.t56 diffpairibias.t29 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 a_n5644_8799.n99 a_n5644_8799.t69 485.149
R1 a_n5644_8799.n106 a_n5644_8799.t72 485.149
R2 a_n5644_8799.n114 a_n5644_8799.t38 485.149
R3 a_n5644_8799.n75 a_n5644_8799.t53 485.149
R4 a_n5644_8799.n82 a_n5644_8799.t58 485.149
R5 a_n5644_8799.n90 a_n5644_8799.t39 485.149
R6 a_n5644_8799.n24 a_n5644_8799.t60 485.135
R7 a_n5644_8799.n103 a_n5644_8799.t59 464.166
R8 a_n5644_8799.n97 a_n5644_8799.t46 464.166
R9 a_n5644_8799.n102 a_n5644_8799.t76 464.166
R10 a_n5644_8799.n101 a_n5644_8799.t61 464.166
R11 a_n5644_8799.n98 a_n5644_8799.t51 464.166
R12 a_n5644_8799.n100 a_n5644_8799.t78 464.166
R13 a_n5644_8799.n29 a_n5644_8799.t64 485.135
R14 a_n5644_8799.n110 a_n5644_8799.t63 464.166
R15 a_n5644_8799.n104 a_n5644_8799.t55 464.166
R16 a_n5644_8799.n109 a_n5644_8799.t80 464.166
R17 a_n5644_8799.n108 a_n5644_8799.t67 464.166
R18 a_n5644_8799.n105 a_n5644_8799.t56 464.166
R19 a_n5644_8799.n107 a_n5644_8799.t36 464.166
R20 a_n5644_8799.n34 a_n5644_8799.t82 485.135
R21 a_n5644_8799.n118 a_n5644_8799.t44 464.166
R22 a_n5644_8799.n112 a_n5644_8799.t65 464.166
R23 a_n5644_8799.n117 a_n5644_8799.t37 464.166
R24 a_n5644_8799.n116 a_n5644_8799.t73 464.166
R25 a_n5644_8799.n113 a_n5644_8799.t50 464.166
R26 a_n5644_8799.n115 a_n5644_8799.t70 464.166
R27 a_n5644_8799.n76 a_n5644_8799.t62 464.166
R28 a_n5644_8799.n77 a_n5644_8799.t77 464.166
R29 a_n5644_8799.n78 a_n5644_8799.t42 464.166
R30 a_n5644_8799.n79 a_n5644_8799.t52 464.166
R31 a_n5644_8799.n74 a_n5644_8799.t75 464.166
R32 a_n5644_8799.n80 a_n5644_8799.t41 464.166
R33 a_n5644_8799.n83 a_n5644_8799.t68 464.166
R34 a_n5644_8799.n84 a_n5644_8799.t81 464.166
R35 a_n5644_8799.n85 a_n5644_8799.t49 464.166
R36 a_n5644_8799.n86 a_n5644_8799.t57 464.166
R37 a_n5644_8799.n81 a_n5644_8799.t79 464.166
R38 a_n5644_8799.n87 a_n5644_8799.t45 464.166
R39 a_n5644_8799.n91 a_n5644_8799.t71 464.166
R40 a_n5644_8799.n92 a_n5644_8799.t48 464.166
R41 a_n5644_8799.n93 a_n5644_8799.t74 464.166
R42 a_n5644_8799.n94 a_n5644_8799.t54 464.166
R43 a_n5644_8799.n89 a_n5644_8799.t66 464.166
R44 a_n5644_8799.n95 a_n5644_8799.t43 464.166
R45 a_n5644_8799.n16 a_n5644_8799.n28 72.3034
R46 a_n5644_8799.n28 a_n5644_8799.n98 16.6962
R47 a_n5644_8799.n27 a_n5644_8799.n16 77.6622
R48 a_n5644_8799.n101 a_n5644_8799.n27 5.97853
R49 a_n5644_8799.n26 a_n5644_8799.n15 77.6622
R50 a_n5644_8799.n15 a_n5644_8799.n25 72.3034
R51 a_n5644_8799.n103 a_n5644_8799.n24 20.9683
R52 a_n5644_8799.n17 a_n5644_8799.n24 70.1674
R53 a_n5644_8799.n13 a_n5644_8799.n33 72.3034
R54 a_n5644_8799.n33 a_n5644_8799.n105 16.6962
R55 a_n5644_8799.n32 a_n5644_8799.n13 77.6622
R56 a_n5644_8799.n108 a_n5644_8799.n32 5.97853
R57 a_n5644_8799.n31 a_n5644_8799.n12 77.6622
R58 a_n5644_8799.n12 a_n5644_8799.n30 72.3034
R59 a_n5644_8799.n110 a_n5644_8799.n29 20.9683
R60 a_n5644_8799.n14 a_n5644_8799.n29 70.1674
R61 a_n5644_8799.n10 a_n5644_8799.n38 72.3034
R62 a_n5644_8799.n38 a_n5644_8799.n113 16.6962
R63 a_n5644_8799.n37 a_n5644_8799.n10 77.6622
R64 a_n5644_8799.n116 a_n5644_8799.n37 5.97853
R65 a_n5644_8799.n36 a_n5644_8799.n9 77.6622
R66 a_n5644_8799.n9 a_n5644_8799.n35 72.3034
R67 a_n5644_8799.n118 a_n5644_8799.n34 20.9683
R68 a_n5644_8799.n11 a_n5644_8799.n34 70.1674
R69 a_n5644_8799.n7 a_n5644_8799.n43 70.1674
R70 a_n5644_8799.n80 a_n5644_8799.n43 20.9683
R71 a_n5644_8799.n42 a_n5644_8799.n7 72.3034
R72 a_n5644_8799.n42 a_n5644_8799.n74 16.6962
R73 a_n5644_8799.n6 a_n5644_8799.n41 77.6622
R74 a_n5644_8799.n79 a_n5644_8799.n41 5.97853
R75 a_n5644_8799.n40 a_n5644_8799.n6 77.6622
R76 a_n5644_8799.n39 a_n5644_8799.n77 16.6962
R77 a_n5644_8799.n39 a_n5644_8799.n8 72.3034
R78 a_n5644_8799.n4 a_n5644_8799.n48 70.1674
R79 a_n5644_8799.n87 a_n5644_8799.n48 20.9683
R80 a_n5644_8799.n47 a_n5644_8799.n4 72.3034
R81 a_n5644_8799.n47 a_n5644_8799.n81 16.6962
R82 a_n5644_8799.n3 a_n5644_8799.n46 77.6622
R83 a_n5644_8799.n86 a_n5644_8799.n46 5.97853
R84 a_n5644_8799.n45 a_n5644_8799.n3 77.6622
R85 a_n5644_8799.n44 a_n5644_8799.n84 16.6962
R86 a_n5644_8799.n44 a_n5644_8799.n5 72.3034
R87 a_n5644_8799.n1 a_n5644_8799.n53 70.1674
R88 a_n5644_8799.n95 a_n5644_8799.n53 20.9683
R89 a_n5644_8799.n52 a_n5644_8799.n1 72.3034
R90 a_n5644_8799.n52 a_n5644_8799.n89 16.6962
R91 a_n5644_8799.n0 a_n5644_8799.n51 77.6622
R92 a_n5644_8799.n94 a_n5644_8799.n51 5.97853
R93 a_n5644_8799.n50 a_n5644_8799.n0 77.6622
R94 a_n5644_8799.n49 a_n5644_8799.n92 16.6962
R95 a_n5644_8799.n49 a_n5644_8799.n2 72.3034
R96 a_n5644_8799.n125 a_n5644_8799.n19 98.9632
R97 a_n5644_8799.n18 a_n5644_8799.n54 98.9631
R98 a_n5644_8799.n19 a_n5644_8799.n123 98.6055
R99 a_n5644_8799.n19 a_n5644_8799.n124 98.6055
R100 a_n5644_8799.n18 a_n5644_8799.n55 98.6055
R101 a_n5644_8799.n18 a_n5644_8799.n56 98.6055
R102 a_n5644_8799.n59 a_n5644_8799.n57 81.4626
R103 a_n5644_8799.n67 a_n5644_8799.n65 81.4626
R104 a_n5644_8799.n63 a_n5644_8799.n61 81.4626
R105 a_n5644_8799.n70 a_n5644_8799.n69 80.9324
R106 a_n5644_8799.n72 a_n5644_8799.n71 80.9324
R107 a_n5644_8799.n23 a_n5644_8799.n73 80.9324
R108 a_n5644_8799.n22 a_n5644_8799.n60 80.9324
R109 a_n5644_8799.n59 a_n5644_8799.n58 80.9324
R110 a_n5644_8799.n67 a_n5644_8799.n66 80.9324
R111 a_n5644_8799.n21 a_n5644_8799.n68 80.9324
R112 a_n5644_8799.n20 a_n5644_8799.n64 80.9324
R113 a_n5644_8799.n63 a_n5644_8799.n62 80.9324
R114 a_n5644_8799.n16 a_n5644_8799.n99 70.4033
R115 a_n5644_8799.n13 a_n5644_8799.n106 70.4033
R116 a_n5644_8799.n10 a_n5644_8799.n114 70.4033
R117 a_n5644_8799.n75 a_n5644_8799.n8 70.4033
R118 a_n5644_8799.n82 a_n5644_8799.n5 70.4033
R119 a_n5644_8799.n90 a_n5644_8799.n2 70.4033
R120 a_n5644_8799.n102 a_n5644_8799.n101 48.2005
R121 a_n5644_8799.n109 a_n5644_8799.n108 48.2005
R122 a_n5644_8799.n117 a_n5644_8799.n116 48.2005
R123 a_n5644_8799.n79 a_n5644_8799.n78 48.2005
R124 a_n5644_8799.t40 a_n5644_8799.n43 485.135
R125 a_n5644_8799.n86 a_n5644_8799.n85 48.2005
R126 a_n5644_8799.t47 a_n5644_8799.n48 485.135
R127 a_n5644_8799.n94 a_n5644_8799.n93 48.2005
R128 a_n5644_8799.t83 a_n5644_8799.n53 485.135
R129 a_n5644_8799.n25 a_n5644_8799.n97 16.6962
R130 a_n5644_8799.n100 a_n5644_8799.n28 27.6507
R131 a_n5644_8799.n30 a_n5644_8799.n104 16.6962
R132 a_n5644_8799.n107 a_n5644_8799.n33 27.6507
R133 a_n5644_8799.n35 a_n5644_8799.n112 16.6962
R134 a_n5644_8799.n115 a_n5644_8799.n38 27.6507
R135 a_n5644_8799.n80 a_n5644_8799.n42 27.6507
R136 a_n5644_8799.n87 a_n5644_8799.n47 27.6507
R137 a_n5644_8799.n95 a_n5644_8799.n52 27.6507
R138 a_n5644_8799.n26 a_n5644_8799.n97 41.7634
R139 a_n5644_8799.n31 a_n5644_8799.n104 41.7634
R140 a_n5644_8799.n36 a_n5644_8799.n112 41.7634
R141 a_n5644_8799.n77 a_n5644_8799.n40 41.7634
R142 a_n5644_8799.n84 a_n5644_8799.n45 41.7634
R143 a_n5644_8799.n92 a_n5644_8799.n50 41.7634
R144 a_n5644_8799.n70 a_n5644_8799.n21 34.3237
R145 a_n5644_8799.n100 a_n5644_8799.n99 20.9576
R146 a_n5644_8799.n107 a_n5644_8799.n106 20.9576
R147 a_n5644_8799.n115 a_n5644_8799.n114 20.9576
R148 a_n5644_8799.n76 a_n5644_8799.n75 20.9576
R149 a_n5644_8799.n83 a_n5644_8799.n82 20.9576
R150 a_n5644_8799.n91 a_n5644_8799.n90 20.9576
R151 a_n5644_8799.n26 a_n5644_8799.n102 5.97853
R152 a_n5644_8799.n27 a_n5644_8799.n98 41.7634
R153 a_n5644_8799.n31 a_n5644_8799.n109 5.97853
R154 a_n5644_8799.n32 a_n5644_8799.n105 41.7634
R155 a_n5644_8799.n36 a_n5644_8799.n117 5.97853
R156 a_n5644_8799.n37 a_n5644_8799.n113 41.7634
R157 a_n5644_8799.n78 a_n5644_8799.n40 5.97853
R158 a_n5644_8799.n74 a_n5644_8799.n41 41.7634
R159 a_n5644_8799.n85 a_n5644_8799.n45 5.97853
R160 a_n5644_8799.n81 a_n5644_8799.n46 41.7634
R161 a_n5644_8799.n93 a_n5644_8799.n50 5.97853
R162 a_n5644_8799.n89 a_n5644_8799.n51 41.7634
R163 a_n5644_8799.n122 a_n5644_8799.n18 31.5519
R164 a_n5644_8799.n121 a_n5644_8799.n23 12.3339
R165 a_n5644_8799.n122 a_n5644_8799.n121 11.4887
R166 a_n5644_8799.n103 a_n5644_8799.n25 27.6507
R167 a_n5644_8799.n110 a_n5644_8799.n30 27.6507
R168 a_n5644_8799.n118 a_n5644_8799.n35 27.6507
R169 a_n5644_8799.n39 a_n5644_8799.n76 27.6507
R170 a_n5644_8799.n44 a_n5644_8799.n83 27.6507
R171 a_n5644_8799.n49 a_n5644_8799.n91 27.6507
R172 a_n5644_8799.n19 a_n5644_8799.n122 17.6132
R173 a_n5644_8799.n111 a_n5644_8799.n17 9.05164
R174 a_n5644_8799.n88 a_n5644_8799.n7 9.05164
R175 a_n5644_8799.n120 a_n5644_8799.n96 6.93972
R176 a_n5644_8799.n120 a_n5644_8799.n119 6.44309
R177 a_n5644_8799.n111 a_n5644_8799.n14 4.94368
R178 a_n5644_8799.n119 a_n5644_8799.n11 4.94368
R179 a_n5644_8799.n88 a_n5644_8799.n4 4.94368
R180 a_n5644_8799.n96 a_n5644_8799.n1 4.94368
R181 a_n5644_8799.n119 a_n5644_8799.n111 4.10845
R182 a_n5644_8799.n96 a_n5644_8799.n88 4.10845
R183 a_n5644_8799.n123 a_n5644_8799.t33 3.61217
R184 a_n5644_8799.n123 a_n5644_8799.t12 3.61217
R185 a_n5644_8799.n124 a_n5644_8799.t28 3.61217
R186 a_n5644_8799.n124 a_n5644_8799.t30 3.61217
R187 a_n5644_8799.n54 a_n5644_8799.t32 3.61217
R188 a_n5644_8799.n54 a_n5644_8799.t23 3.61217
R189 a_n5644_8799.n55 a_n5644_8799.t22 3.61217
R190 a_n5644_8799.n55 a_n5644_8799.t31 3.61217
R191 a_n5644_8799.n56 a_n5644_8799.t34 3.61217
R192 a_n5644_8799.n56 a_n5644_8799.t35 3.61217
R193 a_n5644_8799.t10 a_n5644_8799.n125 3.61217
R194 a_n5644_8799.n125 a_n5644_8799.t27 3.61217
R195 a_n5644_8799.n121 a_n5644_8799.n120 3.4105
R196 a_n5644_8799.n69 a_n5644_8799.t18 2.82907
R197 a_n5644_8799.n69 a_n5644_8799.t7 2.82907
R198 a_n5644_8799.n71 a_n5644_8799.t26 2.82907
R199 a_n5644_8799.n71 a_n5644_8799.t20 2.82907
R200 a_n5644_8799.n73 a_n5644_8799.t29 2.82907
R201 a_n5644_8799.n73 a_n5644_8799.t0 2.82907
R202 a_n5644_8799.n60 a_n5644_8799.t4 2.82907
R203 a_n5644_8799.n60 a_n5644_8799.t2 2.82907
R204 a_n5644_8799.n58 a_n5644_8799.t3 2.82907
R205 a_n5644_8799.n58 a_n5644_8799.t24 2.82907
R206 a_n5644_8799.n57 a_n5644_8799.t16 2.82907
R207 a_n5644_8799.n57 a_n5644_8799.t19 2.82907
R208 a_n5644_8799.n65 a_n5644_8799.t13 2.82907
R209 a_n5644_8799.n65 a_n5644_8799.t1 2.82907
R210 a_n5644_8799.n66 a_n5644_8799.t8 2.82907
R211 a_n5644_8799.n66 a_n5644_8799.t9 2.82907
R212 a_n5644_8799.n68 a_n5644_8799.t11 2.82907
R213 a_n5644_8799.n68 a_n5644_8799.t17 2.82907
R214 a_n5644_8799.n64 a_n5644_8799.t14 2.82907
R215 a_n5644_8799.n64 a_n5644_8799.t5 2.82907
R216 a_n5644_8799.n62 a_n5644_8799.t6 2.82907
R217 a_n5644_8799.n62 a_n5644_8799.t21 2.82907
R218 a_n5644_8799.n61 a_n5644_8799.t25 2.82907
R219 a_n5644_8799.n61 a_n5644_8799.t15 2.82907
R220 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R221 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R222 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R223 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R224 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R225 a_n5644_8799.n1 a_n5644_8799.n0 1.13686
R226 a_n5644_8799.n0 a_n5644_8799.n2 0.568682
R227 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R228 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R229 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R230 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R231 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R232 a_n5644_8799.n20 a_n5644_8799.n63 0.530672
R233 a_n5644_8799.n21 a_n5644_8799.n67 0.530672
R234 a_n5644_8799.n22 a_n5644_8799.n59 0.530672
R235 a_n5644_8799.n23 a_n5644_8799.n72 0.530672
R236 a_n5644_8799.n72 a_n5644_8799.n70 0.530672
R237 a_n5644_8799.n23 a_n5644_8799.n22 0.530672
R238 a_n5644_8799.n21 a_n5644_8799.n20 0.530672
R239 CSoutput.n19 CSoutput.t130 184.661
R240 CSoutput.n78 CSoutput.n77 165.8
R241 CSoutput.n76 CSoutput.n0 165.8
R242 CSoutput.n75 CSoutput.n74 165.8
R243 CSoutput.n73 CSoutput.n72 165.8
R244 CSoutput.n71 CSoutput.n2 165.8
R245 CSoutput.n69 CSoutput.n68 165.8
R246 CSoutput.n67 CSoutput.n3 165.8
R247 CSoutput.n66 CSoutput.n65 165.8
R248 CSoutput.n63 CSoutput.n4 165.8
R249 CSoutput.n61 CSoutput.n60 165.8
R250 CSoutput.n59 CSoutput.n5 165.8
R251 CSoutput.n58 CSoutput.n57 165.8
R252 CSoutput.n55 CSoutput.n6 165.8
R253 CSoutput.n54 CSoutput.n53 165.8
R254 CSoutput.n52 CSoutput.n51 165.8
R255 CSoutput.n50 CSoutput.n8 165.8
R256 CSoutput.n48 CSoutput.n47 165.8
R257 CSoutput.n46 CSoutput.n9 165.8
R258 CSoutput.n45 CSoutput.n44 165.8
R259 CSoutput.n42 CSoutput.n10 165.8
R260 CSoutput.n41 CSoutput.n40 165.8
R261 CSoutput.n39 CSoutput.n38 165.8
R262 CSoutput.n37 CSoutput.n12 165.8
R263 CSoutput.n35 CSoutput.n34 165.8
R264 CSoutput.n33 CSoutput.n13 165.8
R265 CSoutput.n32 CSoutput.n31 165.8
R266 CSoutput.n29 CSoutput.n14 165.8
R267 CSoutput.n28 CSoutput.n27 165.8
R268 CSoutput.n26 CSoutput.n25 165.8
R269 CSoutput.n24 CSoutput.n16 165.8
R270 CSoutput.n22 CSoutput.n21 165.8
R271 CSoutput.n20 CSoutput.n17 165.8
R272 CSoutput.n77 CSoutput.t131 162.194
R273 CSoutput.n18 CSoutput.t149 120.501
R274 CSoutput.n23 CSoutput.t144 120.501
R275 CSoutput.n15 CSoutput.t139 120.501
R276 CSoutput.n30 CSoutput.t128 120.501
R277 CSoutput.n36 CSoutput.t129 120.501
R278 CSoutput.n11 CSoutput.t140 120.501
R279 CSoutput.n43 CSoutput.t136 120.501
R280 CSoutput.n49 CSoutput.t132 120.501
R281 CSoutput.n7 CSoutput.t143 120.501
R282 CSoutput.n56 CSoutput.t146 120.501
R283 CSoutput.n62 CSoutput.t134 120.501
R284 CSoutput.n64 CSoutput.t147 120.501
R285 CSoutput.n70 CSoutput.t148 120.501
R286 CSoutput.n1 CSoutput.t142 120.501
R287 CSoutput.n270 CSoutput.n268 103.469
R288 CSoutput.n262 CSoutput.n260 103.469
R289 CSoutput.n255 CSoutput.n253 103.469
R290 CSoutput.n96 CSoutput.n94 103.469
R291 CSoutput.n88 CSoutput.n86 103.469
R292 CSoutput.n81 CSoutput.n79 103.469
R293 CSoutput.n272 CSoutput.n271 103.111
R294 CSoutput.n270 CSoutput.n269 103.111
R295 CSoutput.n266 CSoutput.n265 103.111
R296 CSoutput.n264 CSoutput.n263 103.111
R297 CSoutput.n262 CSoutput.n261 103.111
R298 CSoutput.n259 CSoutput.n258 103.111
R299 CSoutput.n257 CSoutput.n256 103.111
R300 CSoutput.n255 CSoutput.n254 103.111
R301 CSoutput.n96 CSoutput.n95 103.111
R302 CSoutput.n98 CSoutput.n97 103.111
R303 CSoutput.n100 CSoutput.n99 103.111
R304 CSoutput.n88 CSoutput.n87 103.111
R305 CSoutput.n90 CSoutput.n89 103.111
R306 CSoutput.n92 CSoutput.n91 103.111
R307 CSoutput.n81 CSoutput.n80 103.111
R308 CSoutput.n83 CSoutput.n82 103.111
R309 CSoutput.n85 CSoutput.n84 103.111
R310 CSoutput.n274 CSoutput.n273 103.111
R311 CSoutput.n298 CSoutput.n296 81.5057
R312 CSoutput.n279 CSoutput.n277 81.5057
R313 CSoutput.n338 CSoutput.n336 81.5057
R314 CSoutput.n319 CSoutput.n317 81.5057
R315 CSoutput.n314 CSoutput.n313 80.9324
R316 CSoutput.n312 CSoutput.n311 80.9324
R317 CSoutput.n310 CSoutput.n309 80.9324
R318 CSoutput.n308 CSoutput.n307 80.9324
R319 CSoutput.n306 CSoutput.n305 80.9324
R320 CSoutput.n304 CSoutput.n303 80.9324
R321 CSoutput.n302 CSoutput.n301 80.9324
R322 CSoutput.n300 CSoutput.n299 80.9324
R323 CSoutput.n298 CSoutput.n297 80.9324
R324 CSoutput.n295 CSoutput.n294 80.9324
R325 CSoutput.n293 CSoutput.n292 80.9324
R326 CSoutput.n291 CSoutput.n290 80.9324
R327 CSoutput.n289 CSoutput.n288 80.9324
R328 CSoutput.n287 CSoutput.n286 80.9324
R329 CSoutput.n285 CSoutput.n284 80.9324
R330 CSoutput.n283 CSoutput.n282 80.9324
R331 CSoutput.n281 CSoutput.n280 80.9324
R332 CSoutput.n279 CSoutput.n278 80.9324
R333 CSoutput.n338 CSoutput.n337 80.9324
R334 CSoutput.n340 CSoutput.n339 80.9324
R335 CSoutput.n342 CSoutput.n341 80.9324
R336 CSoutput.n344 CSoutput.n343 80.9324
R337 CSoutput.n346 CSoutput.n345 80.9324
R338 CSoutput.n348 CSoutput.n347 80.9324
R339 CSoutput.n350 CSoutput.n349 80.9324
R340 CSoutput.n352 CSoutput.n351 80.9324
R341 CSoutput.n354 CSoutput.n353 80.9324
R342 CSoutput.n319 CSoutput.n318 80.9324
R343 CSoutput.n321 CSoutput.n320 80.9324
R344 CSoutput.n323 CSoutput.n322 80.9324
R345 CSoutput.n325 CSoutput.n324 80.9324
R346 CSoutput.n327 CSoutput.n326 80.9324
R347 CSoutput.n329 CSoutput.n328 80.9324
R348 CSoutput.n331 CSoutput.n330 80.9324
R349 CSoutput.n333 CSoutput.n332 80.9324
R350 CSoutput.n335 CSoutput.n334 80.9324
R351 CSoutput.n25 CSoutput.n24 48.1486
R352 CSoutput.n69 CSoutput.n3 48.1486
R353 CSoutput.n38 CSoutput.n37 48.1486
R354 CSoutput.n42 CSoutput.n41 48.1486
R355 CSoutput.n51 CSoutput.n50 48.1486
R356 CSoutput.n55 CSoutput.n54 48.1486
R357 CSoutput.n22 CSoutput.n17 46.462
R358 CSoutput.n72 CSoutput.n71 46.462
R359 CSoutput.n20 CSoutput.n19 44.9055
R360 CSoutput.n29 CSoutput.n28 43.7635
R361 CSoutput.n65 CSoutput.n63 43.7635
R362 CSoutput.n35 CSoutput.n13 41.7396
R363 CSoutput.n57 CSoutput.n5 41.7396
R364 CSoutput.n44 CSoutput.n9 37.0171
R365 CSoutput.n48 CSoutput.n9 37.0171
R366 CSoutput.n76 CSoutput.n75 34.9932
R367 CSoutput.n31 CSoutput.n13 32.2947
R368 CSoutput.n61 CSoutput.n5 32.2947
R369 CSoutput.n30 CSoutput.n29 29.6014
R370 CSoutput.n63 CSoutput.n62 29.6014
R371 CSoutput.n19 CSoutput.n18 28.4085
R372 CSoutput.n18 CSoutput.n17 25.1176
R373 CSoutput.n72 CSoutput.n1 25.1176
R374 CSoutput.n43 CSoutput.n42 22.0922
R375 CSoutput.n50 CSoutput.n49 22.0922
R376 CSoutput.n77 CSoutput.n76 21.8586
R377 CSoutput.n37 CSoutput.n36 18.9681
R378 CSoutput.n56 CSoutput.n55 18.9681
R379 CSoutput.n25 CSoutput.n15 17.6292
R380 CSoutput.n64 CSoutput.n3 17.6292
R381 CSoutput.n24 CSoutput.n23 15.844
R382 CSoutput.n70 CSoutput.n69 15.844
R383 CSoutput.n38 CSoutput.n11 14.5051
R384 CSoutput.n54 CSoutput.n7 14.5051
R385 CSoutput.n357 CSoutput.n78 11.6139
R386 CSoutput.n41 CSoutput.n11 11.3811
R387 CSoutput.n51 CSoutput.n7 11.3811
R388 CSoutput.n23 CSoutput.n22 10.0422
R389 CSoutput.n71 CSoutput.n70 10.0422
R390 CSoutput.n316 CSoutput.n276 9.40675
R391 CSoutput.n267 CSoutput.n259 9.25285
R392 CSoutput.n93 CSoutput.n85 9.25285
R393 CSoutput.n315 CSoutput.n295 8.97993
R394 CSoutput.n355 CSoutput.n335 8.97993
R395 CSoutput.n28 CSoutput.n15 8.25698
R396 CSoutput.n65 CSoutput.n64 8.25698
R397 CSoutput.n316 CSoutput.n315 7.89345
R398 CSoutput.n356 CSoutput.n355 7.89345
R399 CSoutput.n276 CSoutput.n275 7.12641
R400 CSoutput.n102 CSoutput.n101 7.12641
R401 CSoutput.n36 CSoutput.n35 6.91809
R402 CSoutput.n57 CSoutput.n56 6.91809
R403 CSoutput.n357 CSoutput.n102 5.81432
R404 CSoutput.n315 CSoutput.n314 5.25266
R405 CSoutput.n355 CSoutput.n354 5.25266
R406 CSoutput.n275 CSoutput.n274 5.1449
R407 CSoutput.n267 CSoutput.n266 5.1449
R408 CSoutput.n101 CSoutput.n100 5.1449
R409 CSoutput.n93 CSoutput.n92 5.1449
R410 CSoutput.n193 CSoutput.n146 4.5005
R411 CSoutput.n162 CSoutput.n146 4.5005
R412 CSoutput.n157 CSoutput.n141 4.5005
R413 CSoutput.n157 CSoutput.n143 4.5005
R414 CSoutput.n157 CSoutput.n140 4.5005
R415 CSoutput.n157 CSoutput.n144 4.5005
R416 CSoutput.n157 CSoutput.n139 4.5005
R417 CSoutput.n157 CSoutput.t135 4.5005
R418 CSoutput.n157 CSoutput.n138 4.5005
R419 CSoutput.n157 CSoutput.n145 4.5005
R420 CSoutput.n157 CSoutput.n146 4.5005
R421 CSoutput.n155 CSoutput.n141 4.5005
R422 CSoutput.n155 CSoutput.n143 4.5005
R423 CSoutput.n155 CSoutput.n140 4.5005
R424 CSoutput.n155 CSoutput.n144 4.5005
R425 CSoutput.n155 CSoutput.n139 4.5005
R426 CSoutput.n155 CSoutput.t135 4.5005
R427 CSoutput.n155 CSoutput.n138 4.5005
R428 CSoutput.n155 CSoutput.n145 4.5005
R429 CSoutput.n155 CSoutput.n146 4.5005
R430 CSoutput.n154 CSoutput.n141 4.5005
R431 CSoutput.n154 CSoutput.n143 4.5005
R432 CSoutput.n154 CSoutput.n140 4.5005
R433 CSoutput.n154 CSoutput.n144 4.5005
R434 CSoutput.n154 CSoutput.n139 4.5005
R435 CSoutput.n154 CSoutput.t135 4.5005
R436 CSoutput.n154 CSoutput.n138 4.5005
R437 CSoutput.n154 CSoutput.n145 4.5005
R438 CSoutput.n154 CSoutput.n146 4.5005
R439 CSoutput.n239 CSoutput.n141 4.5005
R440 CSoutput.n239 CSoutput.n143 4.5005
R441 CSoutput.n239 CSoutput.n140 4.5005
R442 CSoutput.n239 CSoutput.n144 4.5005
R443 CSoutput.n239 CSoutput.n139 4.5005
R444 CSoutput.n239 CSoutput.t135 4.5005
R445 CSoutput.n239 CSoutput.n138 4.5005
R446 CSoutput.n239 CSoutput.n145 4.5005
R447 CSoutput.n239 CSoutput.n146 4.5005
R448 CSoutput.n237 CSoutput.n141 4.5005
R449 CSoutput.n237 CSoutput.n143 4.5005
R450 CSoutput.n237 CSoutput.n140 4.5005
R451 CSoutput.n237 CSoutput.n144 4.5005
R452 CSoutput.n237 CSoutput.n139 4.5005
R453 CSoutput.n237 CSoutput.t135 4.5005
R454 CSoutput.n237 CSoutput.n138 4.5005
R455 CSoutput.n237 CSoutput.n145 4.5005
R456 CSoutput.n235 CSoutput.n141 4.5005
R457 CSoutput.n235 CSoutput.n143 4.5005
R458 CSoutput.n235 CSoutput.n140 4.5005
R459 CSoutput.n235 CSoutput.n144 4.5005
R460 CSoutput.n235 CSoutput.n139 4.5005
R461 CSoutput.n235 CSoutput.t135 4.5005
R462 CSoutput.n235 CSoutput.n138 4.5005
R463 CSoutput.n235 CSoutput.n145 4.5005
R464 CSoutput.n165 CSoutput.n141 4.5005
R465 CSoutput.n165 CSoutput.n143 4.5005
R466 CSoutput.n165 CSoutput.n140 4.5005
R467 CSoutput.n165 CSoutput.n144 4.5005
R468 CSoutput.n165 CSoutput.n139 4.5005
R469 CSoutput.n165 CSoutput.t135 4.5005
R470 CSoutput.n165 CSoutput.n138 4.5005
R471 CSoutput.n165 CSoutput.n145 4.5005
R472 CSoutput.n165 CSoutput.n146 4.5005
R473 CSoutput.n164 CSoutput.n141 4.5005
R474 CSoutput.n164 CSoutput.n143 4.5005
R475 CSoutput.n164 CSoutput.n140 4.5005
R476 CSoutput.n164 CSoutput.n144 4.5005
R477 CSoutput.n164 CSoutput.n139 4.5005
R478 CSoutput.n164 CSoutput.t135 4.5005
R479 CSoutput.n164 CSoutput.n138 4.5005
R480 CSoutput.n164 CSoutput.n145 4.5005
R481 CSoutput.n164 CSoutput.n146 4.5005
R482 CSoutput.n168 CSoutput.n141 4.5005
R483 CSoutput.n168 CSoutput.n143 4.5005
R484 CSoutput.n168 CSoutput.n140 4.5005
R485 CSoutput.n168 CSoutput.n144 4.5005
R486 CSoutput.n168 CSoutput.n139 4.5005
R487 CSoutput.n168 CSoutput.t135 4.5005
R488 CSoutput.n168 CSoutput.n138 4.5005
R489 CSoutput.n168 CSoutput.n145 4.5005
R490 CSoutput.n168 CSoutput.n146 4.5005
R491 CSoutput.n167 CSoutput.n141 4.5005
R492 CSoutput.n167 CSoutput.n143 4.5005
R493 CSoutput.n167 CSoutput.n140 4.5005
R494 CSoutput.n167 CSoutput.n144 4.5005
R495 CSoutput.n167 CSoutput.n139 4.5005
R496 CSoutput.n167 CSoutput.t135 4.5005
R497 CSoutput.n167 CSoutput.n138 4.5005
R498 CSoutput.n167 CSoutput.n145 4.5005
R499 CSoutput.n167 CSoutput.n146 4.5005
R500 CSoutput.n150 CSoutput.n141 4.5005
R501 CSoutput.n150 CSoutput.n143 4.5005
R502 CSoutput.n150 CSoutput.n140 4.5005
R503 CSoutput.n150 CSoutput.n144 4.5005
R504 CSoutput.n150 CSoutput.n139 4.5005
R505 CSoutput.n150 CSoutput.t135 4.5005
R506 CSoutput.n150 CSoutput.n138 4.5005
R507 CSoutput.n150 CSoutput.n145 4.5005
R508 CSoutput.n150 CSoutput.n146 4.5005
R509 CSoutput.n242 CSoutput.n141 4.5005
R510 CSoutput.n242 CSoutput.n143 4.5005
R511 CSoutput.n242 CSoutput.n140 4.5005
R512 CSoutput.n242 CSoutput.n144 4.5005
R513 CSoutput.n242 CSoutput.n139 4.5005
R514 CSoutput.n242 CSoutput.t135 4.5005
R515 CSoutput.n242 CSoutput.n138 4.5005
R516 CSoutput.n242 CSoutput.n145 4.5005
R517 CSoutput.n242 CSoutput.n146 4.5005
R518 CSoutput.n229 CSoutput.n200 4.5005
R519 CSoutput.n229 CSoutput.n206 4.5005
R520 CSoutput.n187 CSoutput.n176 4.5005
R521 CSoutput.n187 CSoutput.n178 4.5005
R522 CSoutput.n187 CSoutput.n175 4.5005
R523 CSoutput.n187 CSoutput.n179 4.5005
R524 CSoutput.n187 CSoutput.n174 4.5005
R525 CSoutput.n187 CSoutput.t137 4.5005
R526 CSoutput.n187 CSoutput.n173 4.5005
R527 CSoutput.n187 CSoutput.n180 4.5005
R528 CSoutput.n229 CSoutput.n187 4.5005
R529 CSoutput.n208 CSoutput.n176 4.5005
R530 CSoutput.n208 CSoutput.n178 4.5005
R531 CSoutput.n208 CSoutput.n175 4.5005
R532 CSoutput.n208 CSoutput.n179 4.5005
R533 CSoutput.n208 CSoutput.n174 4.5005
R534 CSoutput.n208 CSoutput.t137 4.5005
R535 CSoutput.n208 CSoutput.n173 4.5005
R536 CSoutput.n208 CSoutput.n180 4.5005
R537 CSoutput.n229 CSoutput.n208 4.5005
R538 CSoutput.n186 CSoutput.n176 4.5005
R539 CSoutput.n186 CSoutput.n178 4.5005
R540 CSoutput.n186 CSoutput.n175 4.5005
R541 CSoutput.n186 CSoutput.n179 4.5005
R542 CSoutput.n186 CSoutput.n174 4.5005
R543 CSoutput.n186 CSoutput.t137 4.5005
R544 CSoutput.n186 CSoutput.n173 4.5005
R545 CSoutput.n186 CSoutput.n180 4.5005
R546 CSoutput.n229 CSoutput.n186 4.5005
R547 CSoutput.n210 CSoutput.n176 4.5005
R548 CSoutput.n210 CSoutput.n178 4.5005
R549 CSoutput.n210 CSoutput.n175 4.5005
R550 CSoutput.n210 CSoutput.n179 4.5005
R551 CSoutput.n210 CSoutput.n174 4.5005
R552 CSoutput.n210 CSoutput.t137 4.5005
R553 CSoutput.n210 CSoutput.n173 4.5005
R554 CSoutput.n210 CSoutput.n180 4.5005
R555 CSoutput.n229 CSoutput.n210 4.5005
R556 CSoutput.n176 CSoutput.n171 4.5005
R557 CSoutput.n178 CSoutput.n171 4.5005
R558 CSoutput.n175 CSoutput.n171 4.5005
R559 CSoutput.n179 CSoutput.n171 4.5005
R560 CSoutput.n174 CSoutput.n171 4.5005
R561 CSoutput.t137 CSoutput.n171 4.5005
R562 CSoutput.n173 CSoutput.n171 4.5005
R563 CSoutput.n180 CSoutput.n171 4.5005
R564 CSoutput.n232 CSoutput.n176 4.5005
R565 CSoutput.n232 CSoutput.n178 4.5005
R566 CSoutput.n232 CSoutput.n175 4.5005
R567 CSoutput.n232 CSoutput.n179 4.5005
R568 CSoutput.n232 CSoutput.n174 4.5005
R569 CSoutput.n232 CSoutput.t137 4.5005
R570 CSoutput.n232 CSoutput.n173 4.5005
R571 CSoutput.n232 CSoutput.n180 4.5005
R572 CSoutput.n230 CSoutput.n176 4.5005
R573 CSoutput.n230 CSoutput.n178 4.5005
R574 CSoutput.n230 CSoutput.n175 4.5005
R575 CSoutput.n230 CSoutput.n179 4.5005
R576 CSoutput.n230 CSoutput.n174 4.5005
R577 CSoutput.n230 CSoutput.t137 4.5005
R578 CSoutput.n230 CSoutput.n173 4.5005
R579 CSoutput.n230 CSoutput.n180 4.5005
R580 CSoutput.n230 CSoutput.n229 4.5005
R581 CSoutput.n212 CSoutput.n176 4.5005
R582 CSoutput.n212 CSoutput.n178 4.5005
R583 CSoutput.n212 CSoutput.n175 4.5005
R584 CSoutput.n212 CSoutput.n179 4.5005
R585 CSoutput.n212 CSoutput.n174 4.5005
R586 CSoutput.n212 CSoutput.t137 4.5005
R587 CSoutput.n212 CSoutput.n173 4.5005
R588 CSoutput.n212 CSoutput.n180 4.5005
R589 CSoutput.n229 CSoutput.n212 4.5005
R590 CSoutput.n184 CSoutput.n176 4.5005
R591 CSoutput.n184 CSoutput.n178 4.5005
R592 CSoutput.n184 CSoutput.n175 4.5005
R593 CSoutput.n184 CSoutput.n179 4.5005
R594 CSoutput.n184 CSoutput.n174 4.5005
R595 CSoutput.n184 CSoutput.t137 4.5005
R596 CSoutput.n184 CSoutput.n173 4.5005
R597 CSoutput.n184 CSoutput.n180 4.5005
R598 CSoutput.n229 CSoutput.n184 4.5005
R599 CSoutput.n214 CSoutput.n176 4.5005
R600 CSoutput.n214 CSoutput.n178 4.5005
R601 CSoutput.n214 CSoutput.n175 4.5005
R602 CSoutput.n214 CSoutput.n179 4.5005
R603 CSoutput.n214 CSoutput.n174 4.5005
R604 CSoutput.n214 CSoutput.t137 4.5005
R605 CSoutput.n214 CSoutput.n173 4.5005
R606 CSoutput.n214 CSoutput.n180 4.5005
R607 CSoutput.n229 CSoutput.n214 4.5005
R608 CSoutput.n183 CSoutput.n176 4.5005
R609 CSoutput.n183 CSoutput.n178 4.5005
R610 CSoutput.n183 CSoutput.n175 4.5005
R611 CSoutput.n183 CSoutput.n179 4.5005
R612 CSoutput.n183 CSoutput.n174 4.5005
R613 CSoutput.n183 CSoutput.t137 4.5005
R614 CSoutput.n183 CSoutput.n173 4.5005
R615 CSoutput.n183 CSoutput.n180 4.5005
R616 CSoutput.n229 CSoutput.n183 4.5005
R617 CSoutput.n228 CSoutput.n176 4.5005
R618 CSoutput.n228 CSoutput.n178 4.5005
R619 CSoutput.n228 CSoutput.n175 4.5005
R620 CSoutput.n228 CSoutput.n179 4.5005
R621 CSoutput.n228 CSoutput.n174 4.5005
R622 CSoutput.n228 CSoutput.t137 4.5005
R623 CSoutput.n228 CSoutput.n173 4.5005
R624 CSoutput.n228 CSoutput.n180 4.5005
R625 CSoutput.n229 CSoutput.n228 4.5005
R626 CSoutput.n227 CSoutput.n112 4.5005
R627 CSoutput.n128 CSoutput.n112 4.5005
R628 CSoutput.n123 CSoutput.n107 4.5005
R629 CSoutput.n123 CSoutput.n109 4.5005
R630 CSoutput.n123 CSoutput.n106 4.5005
R631 CSoutput.n123 CSoutput.n110 4.5005
R632 CSoutput.n123 CSoutput.n105 4.5005
R633 CSoutput.n123 CSoutput.t138 4.5005
R634 CSoutput.n123 CSoutput.n104 4.5005
R635 CSoutput.n123 CSoutput.n111 4.5005
R636 CSoutput.n123 CSoutput.n112 4.5005
R637 CSoutput.n121 CSoutput.n107 4.5005
R638 CSoutput.n121 CSoutput.n109 4.5005
R639 CSoutput.n121 CSoutput.n106 4.5005
R640 CSoutput.n121 CSoutput.n110 4.5005
R641 CSoutput.n121 CSoutput.n105 4.5005
R642 CSoutput.n121 CSoutput.t138 4.5005
R643 CSoutput.n121 CSoutput.n104 4.5005
R644 CSoutput.n121 CSoutput.n111 4.5005
R645 CSoutput.n121 CSoutput.n112 4.5005
R646 CSoutput.n120 CSoutput.n107 4.5005
R647 CSoutput.n120 CSoutput.n109 4.5005
R648 CSoutput.n120 CSoutput.n106 4.5005
R649 CSoutput.n120 CSoutput.n110 4.5005
R650 CSoutput.n120 CSoutput.n105 4.5005
R651 CSoutput.n120 CSoutput.t138 4.5005
R652 CSoutput.n120 CSoutput.n104 4.5005
R653 CSoutput.n120 CSoutput.n111 4.5005
R654 CSoutput.n120 CSoutput.n112 4.5005
R655 CSoutput.n249 CSoutput.n107 4.5005
R656 CSoutput.n249 CSoutput.n109 4.5005
R657 CSoutput.n249 CSoutput.n106 4.5005
R658 CSoutput.n249 CSoutput.n110 4.5005
R659 CSoutput.n249 CSoutput.n105 4.5005
R660 CSoutput.n249 CSoutput.t138 4.5005
R661 CSoutput.n249 CSoutput.n104 4.5005
R662 CSoutput.n249 CSoutput.n111 4.5005
R663 CSoutput.n249 CSoutput.n112 4.5005
R664 CSoutput.n247 CSoutput.n107 4.5005
R665 CSoutput.n247 CSoutput.n109 4.5005
R666 CSoutput.n247 CSoutput.n106 4.5005
R667 CSoutput.n247 CSoutput.n110 4.5005
R668 CSoutput.n247 CSoutput.n105 4.5005
R669 CSoutput.n247 CSoutput.t138 4.5005
R670 CSoutput.n247 CSoutput.n104 4.5005
R671 CSoutput.n247 CSoutput.n111 4.5005
R672 CSoutput.n245 CSoutput.n107 4.5005
R673 CSoutput.n245 CSoutput.n109 4.5005
R674 CSoutput.n245 CSoutput.n106 4.5005
R675 CSoutput.n245 CSoutput.n110 4.5005
R676 CSoutput.n245 CSoutput.n105 4.5005
R677 CSoutput.n245 CSoutput.t138 4.5005
R678 CSoutput.n245 CSoutput.n104 4.5005
R679 CSoutput.n245 CSoutput.n111 4.5005
R680 CSoutput.n131 CSoutput.n107 4.5005
R681 CSoutput.n131 CSoutput.n109 4.5005
R682 CSoutput.n131 CSoutput.n106 4.5005
R683 CSoutput.n131 CSoutput.n110 4.5005
R684 CSoutput.n131 CSoutput.n105 4.5005
R685 CSoutput.n131 CSoutput.t138 4.5005
R686 CSoutput.n131 CSoutput.n104 4.5005
R687 CSoutput.n131 CSoutput.n111 4.5005
R688 CSoutput.n131 CSoutput.n112 4.5005
R689 CSoutput.n130 CSoutput.n107 4.5005
R690 CSoutput.n130 CSoutput.n109 4.5005
R691 CSoutput.n130 CSoutput.n106 4.5005
R692 CSoutput.n130 CSoutput.n110 4.5005
R693 CSoutput.n130 CSoutput.n105 4.5005
R694 CSoutput.n130 CSoutput.t138 4.5005
R695 CSoutput.n130 CSoutput.n104 4.5005
R696 CSoutput.n130 CSoutput.n111 4.5005
R697 CSoutput.n130 CSoutput.n112 4.5005
R698 CSoutput.n134 CSoutput.n107 4.5005
R699 CSoutput.n134 CSoutput.n109 4.5005
R700 CSoutput.n134 CSoutput.n106 4.5005
R701 CSoutput.n134 CSoutput.n110 4.5005
R702 CSoutput.n134 CSoutput.n105 4.5005
R703 CSoutput.n134 CSoutput.t138 4.5005
R704 CSoutput.n134 CSoutput.n104 4.5005
R705 CSoutput.n134 CSoutput.n111 4.5005
R706 CSoutput.n134 CSoutput.n112 4.5005
R707 CSoutput.n133 CSoutput.n107 4.5005
R708 CSoutput.n133 CSoutput.n109 4.5005
R709 CSoutput.n133 CSoutput.n106 4.5005
R710 CSoutput.n133 CSoutput.n110 4.5005
R711 CSoutput.n133 CSoutput.n105 4.5005
R712 CSoutput.n133 CSoutput.t138 4.5005
R713 CSoutput.n133 CSoutput.n104 4.5005
R714 CSoutput.n133 CSoutput.n111 4.5005
R715 CSoutput.n133 CSoutput.n112 4.5005
R716 CSoutput.n116 CSoutput.n107 4.5005
R717 CSoutput.n116 CSoutput.n109 4.5005
R718 CSoutput.n116 CSoutput.n106 4.5005
R719 CSoutput.n116 CSoutput.n110 4.5005
R720 CSoutput.n116 CSoutput.n105 4.5005
R721 CSoutput.n116 CSoutput.t138 4.5005
R722 CSoutput.n116 CSoutput.n104 4.5005
R723 CSoutput.n116 CSoutput.n111 4.5005
R724 CSoutput.n116 CSoutput.n112 4.5005
R725 CSoutput.n252 CSoutput.n107 4.5005
R726 CSoutput.n252 CSoutput.n109 4.5005
R727 CSoutput.n252 CSoutput.n106 4.5005
R728 CSoutput.n252 CSoutput.n110 4.5005
R729 CSoutput.n252 CSoutput.n105 4.5005
R730 CSoutput.n252 CSoutput.t138 4.5005
R731 CSoutput.n252 CSoutput.n104 4.5005
R732 CSoutput.n252 CSoutput.n111 4.5005
R733 CSoutput.n252 CSoutput.n112 4.5005
R734 CSoutput.n275 CSoutput.n267 4.10845
R735 CSoutput.n101 CSoutput.n93 4.10845
R736 CSoutput.n273 CSoutput.t107 4.06363
R737 CSoutput.n273 CSoutput.t79 4.06363
R738 CSoutput.n271 CSoutput.t88 4.06363
R739 CSoutput.n271 CSoutput.t77 4.06363
R740 CSoutput.n269 CSoutput.t96 4.06363
R741 CSoutput.n269 CSoutput.t103 4.06363
R742 CSoutput.n268 CSoutput.t89 4.06363
R743 CSoutput.n268 CSoutput.t90 4.06363
R744 CSoutput.n265 CSoutput.t91 4.06363
R745 CSoutput.n265 CSoutput.t70 4.06363
R746 CSoutput.n263 CSoutput.t81 4.06363
R747 CSoutput.n263 CSoutput.t99 4.06363
R748 CSoutput.n261 CSoutput.t73 4.06363
R749 CSoutput.n261 CSoutput.t111 4.06363
R750 CSoutput.n260 CSoutput.t101 4.06363
R751 CSoutput.n260 CSoutput.t102 4.06363
R752 CSoutput.n258 CSoutput.t78 4.06363
R753 CSoutput.n258 CSoutput.t67 4.06363
R754 CSoutput.n256 CSoutput.t69 4.06363
R755 CSoutput.n256 CSoutput.t92 4.06363
R756 CSoutput.n254 CSoutput.t100 4.06363
R757 CSoutput.n254 CSoutput.t68 4.06363
R758 CSoutput.n253 CSoutput.t109 4.06363
R759 CSoutput.n253 CSoutput.t84 4.06363
R760 CSoutput.n94 CSoutput.t64 4.06363
R761 CSoutput.n94 CSoutput.t65 4.06363
R762 CSoutput.n95 CSoutput.t76 4.06363
R763 CSoutput.n95 CSoutput.t104 4.06363
R764 CSoutput.n97 CSoutput.t108 4.06363
R765 CSoutput.n97 CSoutput.t86 4.06363
R766 CSoutput.n99 CSoutput.t75 4.06363
R767 CSoutput.n99 CSoutput.t87 4.06363
R768 CSoutput.n86 CSoutput.t83 4.06363
R769 CSoutput.n86 CSoutput.t95 4.06363
R770 CSoutput.n87 CSoutput.t98 4.06363
R771 CSoutput.n87 CSoutput.t106 4.06363
R772 CSoutput.n89 CSoutput.t110 4.06363
R773 CSoutput.n89 CSoutput.t93 4.06363
R774 CSoutput.n91 CSoutput.t97 4.06363
R775 CSoutput.n91 CSoutput.t80 4.06363
R776 CSoutput.n79 CSoutput.t85 4.06363
R777 CSoutput.n79 CSoutput.t72 4.06363
R778 CSoutput.n80 CSoutput.t74 4.06363
R779 CSoutput.n80 CSoutput.t82 4.06363
R780 CSoutput.n82 CSoutput.t94 4.06363
R781 CSoutput.n82 CSoutput.t105 4.06363
R782 CSoutput.n84 CSoutput.t66 4.06363
R783 CSoutput.n84 CSoutput.t71 4.06363
R784 CSoutput.n44 CSoutput.n43 3.79402
R785 CSoutput.n49 CSoutput.n48 3.79402
R786 CSoutput.n356 CSoutput.n316 3.71319
R787 CSoutput.n357 CSoutput.n356 3.57343
R788 CSoutput.n313 CSoutput.t2 2.82907
R789 CSoutput.n313 CSoutput.t41 2.82907
R790 CSoutput.n311 CSoutput.t34 2.82907
R791 CSoutput.n311 CSoutput.t19 2.82907
R792 CSoutput.n309 CSoutput.t9 2.82907
R793 CSoutput.n309 CSoutput.t125 2.82907
R794 CSoutput.n307 CSoutput.t55 2.82907
R795 CSoutput.n307 CSoutput.t115 2.82907
R796 CSoutput.n305 CSoutput.t23 2.82907
R797 CSoutput.n305 CSoutput.t36 2.82907
R798 CSoutput.n303 CSoutput.t119 2.82907
R799 CSoutput.n303 CSoutput.t127 2.82907
R800 CSoutput.n301 CSoutput.t1 2.82907
R801 CSoutput.n301 CSoutput.t58 2.82907
R802 CSoutput.n299 CSoutput.t37 2.82907
R803 CSoutput.n299 CSoutput.t20 2.82907
R804 CSoutput.n297 CSoutput.t123 2.82907
R805 CSoutput.n297 CSoutput.t43 2.82907
R806 CSoutput.n296 CSoutput.t40 2.82907
R807 CSoutput.n296 CSoutput.t117 2.82907
R808 CSoutput.n294 CSoutput.t27 2.82907
R809 CSoutput.n294 CSoutput.t116 2.82907
R810 CSoutput.n292 CSoutput.t16 2.82907
R811 CSoutput.n292 CSoutput.t4 2.82907
R812 CSoutput.n290 CSoutput.t32 2.82907
R813 CSoutput.n290 CSoutput.t38 2.82907
R814 CSoutput.n288 CSoutput.t112 2.82907
R815 CSoutput.n288 CSoutput.t50 2.82907
R816 CSoutput.n286 CSoutput.t62 2.82907
R817 CSoutput.n286 CSoutput.t113 2.82907
R818 CSoutput.n284 CSoutput.t61 2.82907
R819 CSoutput.n284 CSoutput.t22 2.82907
R820 CSoutput.n282 CSoutput.t51 2.82907
R821 CSoutput.n282 CSoutput.t8 2.82907
R822 CSoutput.n280 CSoutput.t17 2.82907
R823 CSoutput.n280 CSoutput.t25 2.82907
R824 CSoutput.n278 CSoutput.t3 2.82907
R825 CSoutput.n278 CSoutput.t53 2.82907
R826 CSoutput.n277 CSoutput.t121 2.82907
R827 CSoutput.n277 CSoutput.t59 2.82907
R828 CSoutput.n336 CSoutput.t31 2.82907
R829 CSoutput.n336 CSoutput.t114 2.82907
R830 CSoutput.n337 CSoutput.t35 2.82907
R831 CSoutput.n337 CSoutput.t49 2.82907
R832 CSoutput.n339 CSoutput.t18 2.82907
R833 CSoutput.n339 CSoutput.t47 2.82907
R834 CSoutput.n341 CSoutput.t52 2.82907
R835 CSoutput.n341 CSoutput.t6 2.82907
R836 CSoutput.n343 CSoutput.t29 2.82907
R837 CSoutput.n343 CSoutput.t14 2.82907
R838 CSoutput.n345 CSoutput.t48 2.82907
R839 CSoutput.n345 CSoutput.t0 2.82907
R840 CSoutput.n347 CSoutput.t13 2.82907
R841 CSoutput.n347 CSoutput.t21 2.82907
R842 CSoutput.n349 CSoutput.t26 2.82907
R843 CSoutput.n349 CSoutput.t124 2.82907
R844 CSoutput.n351 CSoutput.t60 2.82907
R845 CSoutput.n351 CSoutput.t118 2.82907
R846 CSoutput.n353 CSoutput.t39 2.82907
R847 CSoutput.n353 CSoutput.t42 2.82907
R848 CSoutput.n317 CSoutput.t122 2.82907
R849 CSoutput.n317 CSoutput.t45 2.82907
R850 CSoutput.n318 CSoutput.t15 2.82907
R851 CSoutput.n318 CSoutput.t10 2.82907
R852 CSoutput.n320 CSoutput.t5 2.82907
R853 CSoutput.n320 CSoutput.t24 2.82907
R854 CSoutput.n322 CSoutput.t120 2.82907
R855 CSoutput.n322 CSoutput.t63 2.82907
R856 CSoutput.n324 CSoutput.t11 2.82907
R857 CSoutput.n324 CSoutput.t126 2.82907
R858 CSoutput.n326 CSoutput.t7 2.82907
R859 CSoutput.n326 CSoutput.t57 2.82907
R860 CSoutput.n328 CSoutput.t28 2.82907
R861 CSoutput.n328 CSoutput.t30 2.82907
R862 CSoutput.n330 CSoutput.t33 2.82907
R863 CSoutput.n330 CSoutput.t54 2.82907
R864 CSoutput.n332 CSoutput.t12 2.82907
R865 CSoutput.n332 CSoutput.t44 2.82907
R866 CSoutput.n334 CSoutput.t46 2.82907
R867 CSoutput.n334 CSoutput.t56 2.82907
R868 CSoutput.n75 CSoutput.n1 2.45513
R869 CSoutput.n193 CSoutput.n191 2.251
R870 CSoutput.n193 CSoutput.n190 2.251
R871 CSoutput.n193 CSoutput.n189 2.251
R872 CSoutput.n193 CSoutput.n188 2.251
R873 CSoutput.n162 CSoutput.n161 2.251
R874 CSoutput.n162 CSoutput.n160 2.251
R875 CSoutput.n162 CSoutput.n159 2.251
R876 CSoutput.n162 CSoutput.n158 2.251
R877 CSoutput.n235 CSoutput.n234 2.251
R878 CSoutput.n200 CSoutput.n198 2.251
R879 CSoutput.n200 CSoutput.n197 2.251
R880 CSoutput.n200 CSoutput.n196 2.251
R881 CSoutput.n218 CSoutput.n200 2.251
R882 CSoutput.n206 CSoutput.n205 2.251
R883 CSoutput.n206 CSoutput.n204 2.251
R884 CSoutput.n206 CSoutput.n203 2.251
R885 CSoutput.n206 CSoutput.n202 2.251
R886 CSoutput.n232 CSoutput.n172 2.251
R887 CSoutput.n227 CSoutput.n225 2.251
R888 CSoutput.n227 CSoutput.n224 2.251
R889 CSoutput.n227 CSoutput.n223 2.251
R890 CSoutput.n227 CSoutput.n222 2.251
R891 CSoutput.n128 CSoutput.n127 2.251
R892 CSoutput.n128 CSoutput.n126 2.251
R893 CSoutput.n128 CSoutput.n125 2.251
R894 CSoutput.n128 CSoutput.n124 2.251
R895 CSoutput.n245 CSoutput.n244 2.251
R896 CSoutput.n162 CSoutput.n142 2.2505
R897 CSoutput.n157 CSoutput.n142 2.2505
R898 CSoutput.n155 CSoutput.n142 2.2505
R899 CSoutput.n154 CSoutput.n142 2.2505
R900 CSoutput.n239 CSoutput.n142 2.2505
R901 CSoutput.n237 CSoutput.n142 2.2505
R902 CSoutput.n235 CSoutput.n142 2.2505
R903 CSoutput.n165 CSoutput.n142 2.2505
R904 CSoutput.n164 CSoutput.n142 2.2505
R905 CSoutput.n168 CSoutput.n142 2.2505
R906 CSoutput.n167 CSoutput.n142 2.2505
R907 CSoutput.n150 CSoutput.n142 2.2505
R908 CSoutput.n242 CSoutput.n142 2.2505
R909 CSoutput.n242 CSoutput.n241 2.2505
R910 CSoutput.n206 CSoutput.n177 2.2505
R911 CSoutput.n187 CSoutput.n177 2.2505
R912 CSoutput.n208 CSoutput.n177 2.2505
R913 CSoutput.n186 CSoutput.n177 2.2505
R914 CSoutput.n210 CSoutput.n177 2.2505
R915 CSoutput.n177 CSoutput.n171 2.2505
R916 CSoutput.n232 CSoutput.n177 2.2505
R917 CSoutput.n230 CSoutput.n177 2.2505
R918 CSoutput.n212 CSoutput.n177 2.2505
R919 CSoutput.n184 CSoutput.n177 2.2505
R920 CSoutput.n214 CSoutput.n177 2.2505
R921 CSoutput.n183 CSoutput.n177 2.2505
R922 CSoutput.n228 CSoutput.n177 2.2505
R923 CSoutput.n228 CSoutput.n181 2.2505
R924 CSoutput.n128 CSoutput.n108 2.2505
R925 CSoutput.n123 CSoutput.n108 2.2505
R926 CSoutput.n121 CSoutput.n108 2.2505
R927 CSoutput.n120 CSoutput.n108 2.2505
R928 CSoutput.n249 CSoutput.n108 2.2505
R929 CSoutput.n247 CSoutput.n108 2.2505
R930 CSoutput.n245 CSoutput.n108 2.2505
R931 CSoutput.n131 CSoutput.n108 2.2505
R932 CSoutput.n130 CSoutput.n108 2.2505
R933 CSoutput.n134 CSoutput.n108 2.2505
R934 CSoutput.n133 CSoutput.n108 2.2505
R935 CSoutput.n116 CSoutput.n108 2.2505
R936 CSoutput.n252 CSoutput.n108 2.2505
R937 CSoutput.n252 CSoutput.n251 2.2505
R938 CSoutput.n170 CSoutput.n163 2.25024
R939 CSoutput.n170 CSoutput.n156 2.25024
R940 CSoutput.n238 CSoutput.n170 2.25024
R941 CSoutput.n170 CSoutput.n166 2.25024
R942 CSoutput.n170 CSoutput.n169 2.25024
R943 CSoutput.n170 CSoutput.n137 2.25024
R944 CSoutput.n220 CSoutput.n217 2.25024
R945 CSoutput.n220 CSoutput.n216 2.25024
R946 CSoutput.n220 CSoutput.n215 2.25024
R947 CSoutput.n220 CSoutput.n182 2.25024
R948 CSoutput.n220 CSoutput.n219 2.25024
R949 CSoutput.n221 CSoutput.n220 2.25024
R950 CSoutput.n136 CSoutput.n129 2.25024
R951 CSoutput.n136 CSoutput.n122 2.25024
R952 CSoutput.n248 CSoutput.n136 2.25024
R953 CSoutput.n136 CSoutput.n132 2.25024
R954 CSoutput.n136 CSoutput.n135 2.25024
R955 CSoutput.n136 CSoutput.n103 2.25024
R956 CSoutput.n276 CSoutput.n102 1.95131
R957 CSoutput.n237 CSoutput.n147 1.50111
R958 CSoutput.n185 CSoutput.n171 1.50111
R959 CSoutput.n247 CSoutput.n113 1.50111
R960 CSoutput.n193 CSoutput.n192 1.501
R961 CSoutput.n200 CSoutput.n199 1.501
R962 CSoutput.n227 CSoutput.n226 1.501
R963 CSoutput.n241 CSoutput.n152 1.12536
R964 CSoutput.n241 CSoutput.n153 1.12536
R965 CSoutput.n241 CSoutput.n240 1.12536
R966 CSoutput.n201 CSoutput.n181 1.12536
R967 CSoutput.n207 CSoutput.n181 1.12536
R968 CSoutput.n209 CSoutput.n181 1.12536
R969 CSoutput.n251 CSoutput.n118 1.12536
R970 CSoutput.n251 CSoutput.n119 1.12536
R971 CSoutput.n251 CSoutput.n250 1.12536
R972 CSoutput.n241 CSoutput.n148 1.12536
R973 CSoutput.n241 CSoutput.n149 1.12536
R974 CSoutput.n241 CSoutput.n151 1.12536
R975 CSoutput.n231 CSoutput.n181 1.12536
R976 CSoutput.n211 CSoutput.n181 1.12536
R977 CSoutput.n213 CSoutput.n181 1.12536
R978 CSoutput.n251 CSoutput.n114 1.12536
R979 CSoutput.n251 CSoutput.n115 1.12536
R980 CSoutput.n251 CSoutput.n117 1.12536
R981 CSoutput.n31 CSoutput.n30 0.669944
R982 CSoutput.n62 CSoutput.n61 0.669944
R983 CSoutput.n300 CSoutput.n298 0.573776
R984 CSoutput.n302 CSoutput.n300 0.573776
R985 CSoutput.n304 CSoutput.n302 0.573776
R986 CSoutput.n306 CSoutput.n304 0.573776
R987 CSoutput.n308 CSoutput.n306 0.573776
R988 CSoutput.n310 CSoutput.n308 0.573776
R989 CSoutput.n312 CSoutput.n310 0.573776
R990 CSoutput.n314 CSoutput.n312 0.573776
R991 CSoutput.n281 CSoutput.n279 0.573776
R992 CSoutput.n283 CSoutput.n281 0.573776
R993 CSoutput.n285 CSoutput.n283 0.573776
R994 CSoutput.n287 CSoutput.n285 0.573776
R995 CSoutput.n289 CSoutput.n287 0.573776
R996 CSoutput.n291 CSoutput.n289 0.573776
R997 CSoutput.n293 CSoutput.n291 0.573776
R998 CSoutput.n295 CSoutput.n293 0.573776
R999 CSoutput.n354 CSoutput.n352 0.573776
R1000 CSoutput.n352 CSoutput.n350 0.573776
R1001 CSoutput.n350 CSoutput.n348 0.573776
R1002 CSoutput.n348 CSoutput.n346 0.573776
R1003 CSoutput.n346 CSoutput.n344 0.573776
R1004 CSoutput.n344 CSoutput.n342 0.573776
R1005 CSoutput.n342 CSoutput.n340 0.573776
R1006 CSoutput.n340 CSoutput.n338 0.573776
R1007 CSoutput.n335 CSoutput.n333 0.573776
R1008 CSoutput.n333 CSoutput.n331 0.573776
R1009 CSoutput.n331 CSoutput.n329 0.573776
R1010 CSoutput.n329 CSoutput.n327 0.573776
R1011 CSoutput.n327 CSoutput.n325 0.573776
R1012 CSoutput.n325 CSoutput.n323 0.573776
R1013 CSoutput.n323 CSoutput.n321 0.573776
R1014 CSoutput.n321 CSoutput.n319 0.573776
R1015 CSoutput.n357 CSoutput.n252 0.53442
R1016 CSoutput.n272 CSoutput.n270 0.358259
R1017 CSoutput.n274 CSoutput.n272 0.358259
R1018 CSoutput.n264 CSoutput.n262 0.358259
R1019 CSoutput.n266 CSoutput.n264 0.358259
R1020 CSoutput.n257 CSoutput.n255 0.358259
R1021 CSoutput.n259 CSoutput.n257 0.358259
R1022 CSoutput.n100 CSoutput.n98 0.358259
R1023 CSoutput.n98 CSoutput.n96 0.358259
R1024 CSoutput.n92 CSoutput.n90 0.358259
R1025 CSoutput.n90 CSoutput.n88 0.358259
R1026 CSoutput.n85 CSoutput.n83 0.358259
R1027 CSoutput.n83 CSoutput.n81 0.358259
R1028 CSoutput.n21 CSoutput.n20 0.169105
R1029 CSoutput.n21 CSoutput.n16 0.169105
R1030 CSoutput.n26 CSoutput.n16 0.169105
R1031 CSoutput.n27 CSoutput.n26 0.169105
R1032 CSoutput.n27 CSoutput.n14 0.169105
R1033 CSoutput.n32 CSoutput.n14 0.169105
R1034 CSoutput.n33 CSoutput.n32 0.169105
R1035 CSoutput.n34 CSoutput.n33 0.169105
R1036 CSoutput.n34 CSoutput.n12 0.169105
R1037 CSoutput.n39 CSoutput.n12 0.169105
R1038 CSoutput.n40 CSoutput.n39 0.169105
R1039 CSoutput.n40 CSoutput.n10 0.169105
R1040 CSoutput.n45 CSoutput.n10 0.169105
R1041 CSoutput.n46 CSoutput.n45 0.169105
R1042 CSoutput.n47 CSoutput.n46 0.169105
R1043 CSoutput.n47 CSoutput.n8 0.169105
R1044 CSoutput.n52 CSoutput.n8 0.169105
R1045 CSoutput.n53 CSoutput.n52 0.169105
R1046 CSoutput.n53 CSoutput.n6 0.169105
R1047 CSoutput.n58 CSoutput.n6 0.169105
R1048 CSoutput.n59 CSoutput.n58 0.169105
R1049 CSoutput.n60 CSoutput.n59 0.169105
R1050 CSoutput.n60 CSoutput.n4 0.169105
R1051 CSoutput.n66 CSoutput.n4 0.169105
R1052 CSoutput.n67 CSoutput.n66 0.169105
R1053 CSoutput.n68 CSoutput.n67 0.169105
R1054 CSoutput.n68 CSoutput.n2 0.169105
R1055 CSoutput.n73 CSoutput.n2 0.169105
R1056 CSoutput.n74 CSoutput.n73 0.169105
R1057 CSoutput.n74 CSoutput.n0 0.169105
R1058 CSoutput.n78 CSoutput.n0 0.169105
R1059 CSoutput.n195 CSoutput.n194 0.0910737
R1060 CSoutput.n246 CSoutput.n243 0.0723685
R1061 CSoutput.n200 CSoutput.n195 0.0522944
R1062 CSoutput.n243 CSoutput.n242 0.0499135
R1063 CSoutput.n194 CSoutput.n193 0.0499135
R1064 CSoutput.n228 CSoutput.n227 0.0464294
R1065 CSoutput.n236 CSoutput.n233 0.0391444
R1066 CSoutput.n195 CSoutput.t145 0.023435
R1067 CSoutput.n243 CSoutput.t133 0.02262
R1068 CSoutput.n194 CSoutput.t141 0.02262
R1069 CSoutput CSoutput.n357 0.0052
R1070 CSoutput.n165 CSoutput.n148 0.00365111
R1071 CSoutput.n168 CSoutput.n149 0.00365111
R1072 CSoutput.n151 CSoutput.n150 0.00365111
R1073 CSoutput.n193 CSoutput.n152 0.00365111
R1074 CSoutput.n157 CSoutput.n153 0.00365111
R1075 CSoutput.n240 CSoutput.n154 0.00365111
R1076 CSoutput.n231 CSoutput.n230 0.00365111
R1077 CSoutput.n211 CSoutput.n184 0.00365111
R1078 CSoutput.n213 CSoutput.n183 0.00365111
R1079 CSoutput.n201 CSoutput.n200 0.00365111
R1080 CSoutput.n207 CSoutput.n187 0.00365111
R1081 CSoutput.n209 CSoutput.n186 0.00365111
R1082 CSoutput.n131 CSoutput.n114 0.00365111
R1083 CSoutput.n134 CSoutput.n115 0.00365111
R1084 CSoutput.n117 CSoutput.n116 0.00365111
R1085 CSoutput.n227 CSoutput.n118 0.00365111
R1086 CSoutput.n123 CSoutput.n119 0.00365111
R1087 CSoutput.n250 CSoutput.n120 0.00365111
R1088 CSoutput.n162 CSoutput.n152 0.00340054
R1089 CSoutput.n155 CSoutput.n153 0.00340054
R1090 CSoutput.n240 CSoutput.n239 0.00340054
R1091 CSoutput.n235 CSoutput.n148 0.00340054
R1092 CSoutput.n164 CSoutput.n149 0.00340054
R1093 CSoutput.n167 CSoutput.n151 0.00340054
R1094 CSoutput.n206 CSoutput.n201 0.00340054
R1095 CSoutput.n208 CSoutput.n207 0.00340054
R1096 CSoutput.n210 CSoutput.n209 0.00340054
R1097 CSoutput.n232 CSoutput.n231 0.00340054
R1098 CSoutput.n212 CSoutput.n211 0.00340054
R1099 CSoutput.n214 CSoutput.n213 0.00340054
R1100 CSoutput.n128 CSoutput.n118 0.00340054
R1101 CSoutput.n121 CSoutput.n119 0.00340054
R1102 CSoutput.n250 CSoutput.n249 0.00340054
R1103 CSoutput.n245 CSoutput.n114 0.00340054
R1104 CSoutput.n130 CSoutput.n115 0.00340054
R1105 CSoutput.n133 CSoutput.n117 0.00340054
R1106 CSoutput.n163 CSoutput.n157 0.00252698
R1107 CSoutput.n156 CSoutput.n154 0.00252698
R1108 CSoutput.n238 CSoutput.n237 0.00252698
R1109 CSoutput.n166 CSoutput.n164 0.00252698
R1110 CSoutput.n169 CSoutput.n167 0.00252698
R1111 CSoutput.n242 CSoutput.n137 0.00252698
R1112 CSoutput.n163 CSoutput.n162 0.00252698
R1113 CSoutput.n156 CSoutput.n155 0.00252698
R1114 CSoutput.n239 CSoutput.n238 0.00252698
R1115 CSoutput.n166 CSoutput.n165 0.00252698
R1116 CSoutput.n169 CSoutput.n168 0.00252698
R1117 CSoutput.n150 CSoutput.n137 0.00252698
R1118 CSoutput.n217 CSoutput.n187 0.00252698
R1119 CSoutput.n216 CSoutput.n186 0.00252698
R1120 CSoutput.n215 CSoutput.n171 0.00252698
R1121 CSoutput.n212 CSoutput.n182 0.00252698
R1122 CSoutput.n219 CSoutput.n214 0.00252698
R1123 CSoutput.n228 CSoutput.n221 0.00252698
R1124 CSoutput.n217 CSoutput.n206 0.00252698
R1125 CSoutput.n216 CSoutput.n208 0.00252698
R1126 CSoutput.n215 CSoutput.n210 0.00252698
R1127 CSoutput.n230 CSoutput.n182 0.00252698
R1128 CSoutput.n219 CSoutput.n184 0.00252698
R1129 CSoutput.n221 CSoutput.n183 0.00252698
R1130 CSoutput.n129 CSoutput.n123 0.00252698
R1131 CSoutput.n122 CSoutput.n120 0.00252698
R1132 CSoutput.n248 CSoutput.n247 0.00252698
R1133 CSoutput.n132 CSoutput.n130 0.00252698
R1134 CSoutput.n135 CSoutput.n133 0.00252698
R1135 CSoutput.n252 CSoutput.n103 0.00252698
R1136 CSoutput.n129 CSoutput.n128 0.00252698
R1137 CSoutput.n122 CSoutput.n121 0.00252698
R1138 CSoutput.n249 CSoutput.n248 0.00252698
R1139 CSoutput.n132 CSoutput.n131 0.00252698
R1140 CSoutput.n135 CSoutput.n134 0.00252698
R1141 CSoutput.n116 CSoutput.n103 0.00252698
R1142 CSoutput.n237 CSoutput.n236 0.0020275
R1143 CSoutput.n236 CSoutput.n235 0.0020275
R1144 CSoutput.n233 CSoutput.n171 0.0020275
R1145 CSoutput.n233 CSoutput.n232 0.0020275
R1146 CSoutput.n247 CSoutput.n246 0.0020275
R1147 CSoutput.n246 CSoutput.n245 0.0020275
R1148 CSoutput.n147 CSoutput.n146 0.00166668
R1149 CSoutput.n229 CSoutput.n185 0.00166668
R1150 CSoutput.n113 CSoutput.n112 0.00166668
R1151 CSoutput.n251 CSoutput.n113 0.00133328
R1152 CSoutput.n185 CSoutput.n181 0.00133328
R1153 CSoutput.n241 CSoutput.n147 0.00133328
R1154 CSoutput.n244 CSoutput.n136 0.001
R1155 CSoutput.n222 CSoutput.n136 0.001
R1156 CSoutput.n124 CSoutput.n104 0.001
R1157 CSoutput.n223 CSoutput.n104 0.001
R1158 CSoutput.n125 CSoutput.n105 0.001
R1159 CSoutput.n224 CSoutput.n105 0.001
R1160 CSoutput.n126 CSoutput.n106 0.001
R1161 CSoutput.n225 CSoutput.n106 0.001
R1162 CSoutput.n127 CSoutput.n107 0.001
R1163 CSoutput.n226 CSoutput.n107 0.001
R1164 CSoutput.n220 CSoutput.n172 0.001
R1165 CSoutput.n220 CSoutput.n218 0.001
R1166 CSoutput.n202 CSoutput.n173 0.001
R1167 CSoutput.n196 CSoutput.n173 0.001
R1168 CSoutput.n203 CSoutput.n174 0.001
R1169 CSoutput.n197 CSoutput.n174 0.001
R1170 CSoutput.n204 CSoutput.n175 0.001
R1171 CSoutput.n198 CSoutput.n175 0.001
R1172 CSoutput.n205 CSoutput.n176 0.001
R1173 CSoutput.n199 CSoutput.n176 0.001
R1174 CSoutput.n234 CSoutput.n170 0.001
R1175 CSoutput.n188 CSoutput.n170 0.001
R1176 CSoutput.n158 CSoutput.n138 0.001
R1177 CSoutput.n189 CSoutput.n138 0.001
R1178 CSoutput.n159 CSoutput.n139 0.001
R1179 CSoutput.n190 CSoutput.n139 0.001
R1180 CSoutput.n160 CSoutput.n140 0.001
R1181 CSoutput.n191 CSoutput.n140 0.001
R1182 CSoutput.n161 CSoutput.n141 0.001
R1183 CSoutput.n192 CSoutput.n141 0.001
R1184 CSoutput.n192 CSoutput.n142 0.001
R1185 CSoutput.n191 CSoutput.n143 0.001
R1186 CSoutput.n190 CSoutput.n144 0.001
R1187 CSoutput.n189 CSoutput.t135 0.001
R1188 CSoutput.n188 CSoutput.n145 0.001
R1189 CSoutput.n161 CSoutput.n143 0.001
R1190 CSoutput.n160 CSoutput.n144 0.001
R1191 CSoutput.n159 CSoutput.t135 0.001
R1192 CSoutput.n158 CSoutput.n145 0.001
R1193 CSoutput.n234 CSoutput.n146 0.001
R1194 CSoutput.n199 CSoutput.n177 0.001
R1195 CSoutput.n198 CSoutput.n178 0.001
R1196 CSoutput.n197 CSoutput.n179 0.001
R1197 CSoutput.n196 CSoutput.t137 0.001
R1198 CSoutput.n218 CSoutput.n180 0.001
R1199 CSoutput.n205 CSoutput.n178 0.001
R1200 CSoutput.n204 CSoutput.n179 0.001
R1201 CSoutput.n203 CSoutput.t137 0.001
R1202 CSoutput.n202 CSoutput.n180 0.001
R1203 CSoutput.n229 CSoutput.n172 0.001
R1204 CSoutput.n226 CSoutput.n108 0.001
R1205 CSoutput.n225 CSoutput.n109 0.001
R1206 CSoutput.n224 CSoutput.n110 0.001
R1207 CSoutput.n223 CSoutput.t138 0.001
R1208 CSoutput.n222 CSoutput.n111 0.001
R1209 CSoutput.n127 CSoutput.n109 0.001
R1210 CSoutput.n126 CSoutput.n110 0.001
R1211 CSoutput.n125 CSoutput.t138 0.001
R1212 CSoutput.n124 CSoutput.n111 0.001
R1213 CSoutput.n244 CSoutput.n112 0.001
R1214 vdd.n291 vdd.n255 756.745
R1215 vdd.n244 vdd.n208 756.745
R1216 vdd.n201 vdd.n165 756.745
R1217 vdd.n154 vdd.n118 756.745
R1218 vdd.n112 vdd.n76 756.745
R1219 vdd.n65 vdd.n29 756.745
R1220 vdd.n1106 vdd.n1070 756.745
R1221 vdd.n1153 vdd.n1117 756.745
R1222 vdd.n1016 vdd.n980 756.745
R1223 vdd.n1063 vdd.n1027 756.745
R1224 vdd.n927 vdd.n891 756.745
R1225 vdd.n974 vdd.n938 756.745
R1226 vdd.n1791 vdd.t79 640.208
R1227 vdd.n755 vdd.t64 640.208
R1228 vdd.n1765 vdd.t105 640.208
R1229 vdd.n747 vdd.t96 640.208
R1230 vdd.n2536 vdd.t47 640.208
R1231 vdd.n2256 vdd.t87 640.208
R1232 vdd.n622 vdd.t68 640.208
R1233 vdd.n2253 vdd.t72 640.208
R1234 vdd.n589 vdd.t76 640.208
R1235 vdd.n817 vdd.t83 640.208
R1236 vdd.n1320 vdd.t43 592.009
R1237 vdd.n1358 vdd.t90 592.009
R1238 vdd.n1254 vdd.t93 592.009
R1239 vdd.n1947 vdd.t39 592.009
R1240 vdd.n1584 vdd.t51 592.009
R1241 vdd.n1544 vdd.t58 592.009
R1242 vdd.n2908 vdd.t102 592.009
R1243 vdd.n405 vdd.t54 592.009
R1244 vdd.n365 vdd.t61 592.009
R1245 vdd.n557 vdd.t32 592.009
R1246 vdd.n2804 vdd.t36 592.009
R1247 vdd.n2711 vdd.t99 592.009
R1248 vdd.n292 vdd.n291 585
R1249 vdd.n290 vdd.n257 585
R1250 vdd.n289 vdd.n288 585
R1251 vdd.n260 vdd.n258 585
R1252 vdd.n283 vdd.n282 585
R1253 vdd.n281 vdd.n280 585
R1254 vdd.n264 vdd.n263 585
R1255 vdd.n275 vdd.n274 585
R1256 vdd.n273 vdd.n272 585
R1257 vdd.n268 vdd.n267 585
R1258 vdd.n245 vdd.n244 585
R1259 vdd.n243 vdd.n210 585
R1260 vdd.n242 vdd.n241 585
R1261 vdd.n213 vdd.n211 585
R1262 vdd.n236 vdd.n235 585
R1263 vdd.n234 vdd.n233 585
R1264 vdd.n217 vdd.n216 585
R1265 vdd.n228 vdd.n227 585
R1266 vdd.n226 vdd.n225 585
R1267 vdd.n221 vdd.n220 585
R1268 vdd.n202 vdd.n201 585
R1269 vdd.n200 vdd.n167 585
R1270 vdd.n199 vdd.n198 585
R1271 vdd.n170 vdd.n168 585
R1272 vdd.n193 vdd.n192 585
R1273 vdd.n191 vdd.n190 585
R1274 vdd.n174 vdd.n173 585
R1275 vdd.n185 vdd.n184 585
R1276 vdd.n183 vdd.n182 585
R1277 vdd.n178 vdd.n177 585
R1278 vdd.n155 vdd.n154 585
R1279 vdd.n153 vdd.n120 585
R1280 vdd.n152 vdd.n151 585
R1281 vdd.n123 vdd.n121 585
R1282 vdd.n146 vdd.n145 585
R1283 vdd.n144 vdd.n143 585
R1284 vdd.n127 vdd.n126 585
R1285 vdd.n138 vdd.n137 585
R1286 vdd.n136 vdd.n135 585
R1287 vdd.n131 vdd.n130 585
R1288 vdd.n113 vdd.n112 585
R1289 vdd.n111 vdd.n78 585
R1290 vdd.n110 vdd.n109 585
R1291 vdd.n81 vdd.n79 585
R1292 vdd.n104 vdd.n103 585
R1293 vdd.n102 vdd.n101 585
R1294 vdd.n85 vdd.n84 585
R1295 vdd.n96 vdd.n95 585
R1296 vdd.n94 vdd.n93 585
R1297 vdd.n89 vdd.n88 585
R1298 vdd.n66 vdd.n65 585
R1299 vdd.n64 vdd.n31 585
R1300 vdd.n63 vdd.n62 585
R1301 vdd.n34 vdd.n32 585
R1302 vdd.n57 vdd.n56 585
R1303 vdd.n55 vdd.n54 585
R1304 vdd.n38 vdd.n37 585
R1305 vdd.n49 vdd.n48 585
R1306 vdd.n47 vdd.n46 585
R1307 vdd.n42 vdd.n41 585
R1308 vdd.n1107 vdd.n1106 585
R1309 vdd.n1105 vdd.n1072 585
R1310 vdd.n1104 vdd.n1103 585
R1311 vdd.n1075 vdd.n1073 585
R1312 vdd.n1098 vdd.n1097 585
R1313 vdd.n1096 vdd.n1095 585
R1314 vdd.n1079 vdd.n1078 585
R1315 vdd.n1090 vdd.n1089 585
R1316 vdd.n1088 vdd.n1087 585
R1317 vdd.n1083 vdd.n1082 585
R1318 vdd.n1154 vdd.n1153 585
R1319 vdd.n1152 vdd.n1119 585
R1320 vdd.n1151 vdd.n1150 585
R1321 vdd.n1122 vdd.n1120 585
R1322 vdd.n1145 vdd.n1144 585
R1323 vdd.n1143 vdd.n1142 585
R1324 vdd.n1126 vdd.n1125 585
R1325 vdd.n1137 vdd.n1136 585
R1326 vdd.n1135 vdd.n1134 585
R1327 vdd.n1130 vdd.n1129 585
R1328 vdd.n1017 vdd.n1016 585
R1329 vdd.n1015 vdd.n982 585
R1330 vdd.n1014 vdd.n1013 585
R1331 vdd.n985 vdd.n983 585
R1332 vdd.n1008 vdd.n1007 585
R1333 vdd.n1006 vdd.n1005 585
R1334 vdd.n989 vdd.n988 585
R1335 vdd.n1000 vdd.n999 585
R1336 vdd.n998 vdd.n997 585
R1337 vdd.n993 vdd.n992 585
R1338 vdd.n1064 vdd.n1063 585
R1339 vdd.n1062 vdd.n1029 585
R1340 vdd.n1061 vdd.n1060 585
R1341 vdd.n1032 vdd.n1030 585
R1342 vdd.n1055 vdd.n1054 585
R1343 vdd.n1053 vdd.n1052 585
R1344 vdd.n1036 vdd.n1035 585
R1345 vdd.n1047 vdd.n1046 585
R1346 vdd.n1045 vdd.n1044 585
R1347 vdd.n1040 vdd.n1039 585
R1348 vdd.n928 vdd.n927 585
R1349 vdd.n926 vdd.n893 585
R1350 vdd.n925 vdd.n924 585
R1351 vdd.n896 vdd.n894 585
R1352 vdd.n919 vdd.n918 585
R1353 vdd.n917 vdd.n916 585
R1354 vdd.n900 vdd.n899 585
R1355 vdd.n911 vdd.n910 585
R1356 vdd.n909 vdd.n908 585
R1357 vdd.n904 vdd.n903 585
R1358 vdd.n975 vdd.n974 585
R1359 vdd.n973 vdd.n940 585
R1360 vdd.n972 vdd.n971 585
R1361 vdd.n943 vdd.n941 585
R1362 vdd.n966 vdd.n965 585
R1363 vdd.n964 vdd.n963 585
R1364 vdd.n947 vdd.n946 585
R1365 vdd.n958 vdd.n957 585
R1366 vdd.n956 vdd.n955 585
R1367 vdd.n951 vdd.n950 585
R1368 vdd.n3024 vdd.n330 515.122
R1369 vdd.n2906 vdd.n328 515.122
R1370 vdd.n515 vdd.n478 515.122
R1371 vdd.n2842 vdd.n479 515.122
R1372 vdd.n1942 vdd.n865 515.122
R1373 vdd.n1945 vdd.n1944 515.122
R1374 vdd.n1227 vdd.n1191 515.122
R1375 vdd.n1423 vdd.n1192 515.122
R1376 vdd.n269 vdd.t144 329.043
R1377 vdd.n222 vdd.t155 329.043
R1378 vdd.n179 vdd.t140 329.043
R1379 vdd.n132 vdd.t150 329.043
R1380 vdd.n90 vdd.t181 329.043
R1381 vdd.n43 vdd.t123 329.043
R1382 vdd.n1084 vdd.t179 329.043
R1383 vdd.n1131 vdd.t165 329.043
R1384 vdd.n994 vdd.t171 329.043
R1385 vdd.n1041 vdd.t158 329.043
R1386 vdd.n905 vdd.t121 329.043
R1387 vdd.n952 vdd.t180 329.043
R1388 vdd.n1320 vdd.t46 319.788
R1389 vdd.n1358 vdd.t92 319.788
R1390 vdd.n1254 vdd.t95 319.788
R1391 vdd.n1947 vdd.t41 319.788
R1392 vdd.n1584 vdd.t52 319.788
R1393 vdd.n1544 vdd.t59 319.788
R1394 vdd.n2908 vdd.t103 319.788
R1395 vdd.n405 vdd.t56 319.788
R1396 vdd.n365 vdd.t62 319.788
R1397 vdd.n557 vdd.t35 319.788
R1398 vdd.n2804 vdd.t38 319.788
R1399 vdd.n2711 vdd.t101 319.788
R1400 vdd.n1321 vdd.t45 303.69
R1401 vdd.n1359 vdd.t91 303.69
R1402 vdd.n1255 vdd.t94 303.69
R1403 vdd.n1948 vdd.t42 303.69
R1404 vdd.n1585 vdd.t53 303.69
R1405 vdd.n1545 vdd.t60 303.69
R1406 vdd.n2909 vdd.t104 303.69
R1407 vdd.n406 vdd.t57 303.69
R1408 vdd.n366 vdd.t63 303.69
R1409 vdd.n558 vdd.t34 303.69
R1410 vdd.n2805 vdd.t37 303.69
R1411 vdd.n2712 vdd.t100 303.69
R1412 vdd.n2479 vdd.n703 297.074
R1413 vdd.n2672 vdd.n599 297.074
R1414 vdd.n2609 vdd.n596 297.074
R1415 vdd.n2402 vdd.n704 297.074
R1416 vdd.n2217 vdd.n744 297.074
R1417 vdd.n2148 vdd.n2147 297.074
R1418 vdd.n1894 vdd.n840 297.074
R1419 vdd.n1990 vdd.n838 297.074
R1420 vdd.n2588 vdd.n597 297.074
R1421 vdd.n2675 vdd.n2674 297.074
R1422 vdd.n2251 vdd.n705 297.074
R1423 vdd.n2477 vdd.n706 297.074
R1424 vdd.n2145 vdd.n753 297.074
R1425 vdd.n751 vdd.n726 297.074
R1426 vdd.n1831 vdd.n841 297.074
R1427 vdd.n1988 vdd.n842 297.074
R1428 vdd.n2590 vdd.n597 185
R1429 vdd.n2673 vdd.n597 185
R1430 vdd.n2592 vdd.n2591 185
R1431 vdd.n2591 vdd.n595 185
R1432 vdd.n2593 vdd.n629 185
R1433 vdd.n2603 vdd.n629 185
R1434 vdd.n2594 vdd.n638 185
R1435 vdd.n638 vdd.n636 185
R1436 vdd.n2596 vdd.n2595 185
R1437 vdd.n2597 vdd.n2596 185
R1438 vdd.n2549 vdd.n637 185
R1439 vdd.n637 vdd.n633 185
R1440 vdd.n2548 vdd.n2547 185
R1441 vdd.n2547 vdd.n2546 185
R1442 vdd.n640 vdd.n639 185
R1443 vdd.n641 vdd.n640 185
R1444 vdd.n2539 vdd.n2538 185
R1445 vdd.n2540 vdd.n2539 185
R1446 vdd.n2535 vdd.n650 185
R1447 vdd.n650 vdd.n647 185
R1448 vdd.n2534 vdd.n2533 185
R1449 vdd.n2533 vdd.n2532 185
R1450 vdd.n652 vdd.n651 185
R1451 vdd.n660 vdd.n652 185
R1452 vdd.n2525 vdd.n2524 185
R1453 vdd.n2526 vdd.n2525 185
R1454 vdd.n2523 vdd.n661 185
R1455 vdd.n2374 vdd.n661 185
R1456 vdd.n2522 vdd.n2521 185
R1457 vdd.n2521 vdd.n2520 185
R1458 vdd.n663 vdd.n662 185
R1459 vdd.n664 vdd.n663 185
R1460 vdd.n2513 vdd.n2512 185
R1461 vdd.n2514 vdd.n2513 185
R1462 vdd.n2511 vdd.n673 185
R1463 vdd.n673 vdd.n670 185
R1464 vdd.n2510 vdd.n2509 185
R1465 vdd.n2509 vdd.n2508 185
R1466 vdd.n675 vdd.n674 185
R1467 vdd.n683 vdd.n675 185
R1468 vdd.n2501 vdd.n2500 185
R1469 vdd.n2502 vdd.n2501 185
R1470 vdd.n2499 vdd.n684 185
R1471 vdd.n690 vdd.n684 185
R1472 vdd.n2498 vdd.n2497 185
R1473 vdd.n2497 vdd.n2496 185
R1474 vdd.n686 vdd.n685 185
R1475 vdd.n687 vdd.n686 185
R1476 vdd.n2489 vdd.n2488 185
R1477 vdd.n2490 vdd.n2489 185
R1478 vdd.n2487 vdd.n696 185
R1479 vdd.n2395 vdd.n696 185
R1480 vdd.n2486 vdd.n2485 185
R1481 vdd.n2485 vdd.n2484 185
R1482 vdd.n698 vdd.n697 185
R1483 vdd.t186 vdd.n698 185
R1484 vdd.n2477 vdd.n2476 185
R1485 vdd.n2478 vdd.n2477 185
R1486 vdd.n2475 vdd.n706 185
R1487 vdd.n2474 vdd.n2473 185
R1488 vdd.n708 vdd.n707 185
R1489 vdd.n2260 vdd.n2259 185
R1490 vdd.n2262 vdd.n2261 185
R1491 vdd.n2264 vdd.n2263 185
R1492 vdd.n2266 vdd.n2265 185
R1493 vdd.n2268 vdd.n2267 185
R1494 vdd.n2270 vdd.n2269 185
R1495 vdd.n2272 vdd.n2271 185
R1496 vdd.n2274 vdd.n2273 185
R1497 vdd.n2276 vdd.n2275 185
R1498 vdd.n2278 vdd.n2277 185
R1499 vdd.n2280 vdd.n2279 185
R1500 vdd.n2282 vdd.n2281 185
R1501 vdd.n2284 vdd.n2283 185
R1502 vdd.n2286 vdd.n2285 185
R1503 vdd.n2288 vdd.n2287 185
R1504 vdd.n2290 vdd.n2289 185
R1505 vdd.n2292 vdd.n2291 185
R1506 vdd.n2294 vdd.n2293 185
R1507 vdd.n2296 vdd.n2295 185
R1508 vdd.n2298 vdd.n2297 185
R1509 vdd.n2300 vdd.n2299 185
R1510 vdd.n2302 vdd.n2301 185
R1511 vdd.n2304 vdd.n2303 185
R1512 vdd.n2306 vdd.n2305 185
R1513 vdd.n2308 vdd.n2307 185
R1514 vdd.n2310 vdd.n2309 185
R1515 vdd.n2312 vdd.n2311 185
R1516 vdd.n2314 vdd.n2313 185
R1517 vdd.n2316 vdd.n2315 185
R1518 vdd.n2318 vdd.n2317 185
R1519 vdd.n2320 vdd.n2319 185
R1520 vdd.n2321 vdd.n2251 185
R1521 vdd.n2471 vdd.n2251 185
R1522 vdd.n2676 vdd.n2675 185
R1523 vdd.n2677 vdd.n588 185
R1524 vdd.n2679 vdd.n2678 185
R1525 vdd.n2681 vdd.n586 185
R1526 vdd.n2683 vdd.n2682 185
R1527 vdd.n2684 vdd.n585 185
R1528 vdd.n2686 vdd.n2685 185
R1529 vdd.n2688 vdd.n583 185
R1530 vdd.n2690 vdd.n2689 185
R1531 vdd.n2691 vdd.n582 185
R1532 vdd.n2693 vdd.n2692 185
R1533 vdd.n2695 vdd.n580 185
R1534 vdd.n2697 vdd.n2696 185
R1535 vdd.n2698 vdd.n579 185
R1536 vdd.n2700 vdd.n2699 185
R1537 vdd.n2702 vdd.n578 185
R1538 vdd.n2703 vdd.n576 185
R1539 vdd.n2706 vdd.n2705 185
R1540 vdd.n577 vdd.n575 185
R1541 vdd.n2562 vdd.n2561 185
R1542 vdd.n2564 vdd.n2563 185
R1543 vdd.n2566 vdd.n2558 185
R1544 vdd.n2568 vdd.n2567 185
R1545 vdd.n2569 vdd.n2557 185
R1546 vdd.n2571 vdd.n2570 185
R1547 vdd.n2573 vdd.n2555 185
R1548 vdd.n2575 vdd.n2574 185
R1549 vdd.n2576 vdd.n2554 185
R1550 vdd.n2578 vdd.n2577 185
R1551 vdd.n2580 vdd.n2552 185
R1552 vdd.n2582 vdd.n2581 185
R1553 vdd.n2583 vdd.n2551 185
R1554 vdd.n2585 vdd.n2584 185
R1555 vdd.n2587 vdd.n2550 185
R1556 vdd.n2589 vdd.n2588 185
R1557 vdd.n2588 vdd.n484 185
R1558 vdd.n2674 vdd.n592 185
R1559 vdd.n2674 vdd.n2673 185
R1560 vdd.n2326 vdd.n594 185
R1561 vdd.n595 vdd.n594 185
R1562 vdd.n2327 vdd.n628 185
R1563 vdd.n2603 vdd.n628 185
R1564 vdd.n2329 vdd.n2328 185
R1565 vdd.n2328 vdd.n636 185
R1566 vdd.n2330 vdd.n635 185
R1567 vdd.n2597 vdd.n635 185
R1568 vdd.n2332 vdd.n2331 185
R1569 vdd.n2331 vdd.n633 185
R1570 vdd.n2333 vdd.n643 185
R1571 vdd.n2546 vdd.n643 185
R1572 vdd.n2335 vdd.n2334 185
R1573 vdd.n2334 vdd.n641 185
R1574 vdd.n2336 vdd.n649 185
R1575 vdd.n2540 vdd.n649 185
R1576 vdd.n2338 vdd.n2337 185
R1577 vdd.n2337 vdd.n647 185
R1578 vdd.n2339 vdd.n654 185
R1579 vdd.n2532 vdd.n654 185
R1580 vdd.n2341 vdd.n2340 185
R1581 vdd.n2340 vdd.n660 185
R1582 vdd.n2342 vdd.n659 185
R1583 vdd.n2526 vdd.n659 185
R1584 vdd.n2376 vdd.n2375 185
R1585 vdd.n2375 vdd.n2374 185
R1586 vdd.n2377 vdd.n666 185
R1587 vdd.n2520 vdd.n666 185
R1588 vdd.n2379 vdd.n2378 185
R1589 vdd.n2378 vdd.n664 185
R1590 vdd.n2380 vdd.n672 185
R1591 vdd.n2514 vdd.n672 185
R1592 vdd.n2382 vdd.n2381 185
R1593 vdd.n2381 vdd.n670 185
R1594 vdd.n2383 vdd.n677 185
R1595 vdd.n2508 vdd.n677 185
R1596 vdd.n2385 vdd.n2384 185
R1597 vdd.n2384 vdd.n683 185
R1598 vdd.n2386 vdd.n682 185
R1599 vdd.n2502 vdd.n682 185
R1600 vdd.n2388 vdd.n2387 185
R1601 vdd.n2387 vdd.n690 185
R1602 vdd.n2389 vdd.n689 185
R1603 vdd.n2496 vdd.n689 185
R1604 vdd.n2391 vdd.n2390 185
R1605 vdd.n2390 vdd.n687 185
R1606 vdd.n2392 vdd.n695 185
R1607 vdd.n2490 vdd.n695 185
R1608 vdd.n2394 vdd.n2393 185
R1609 vdd.n2395 vdd.n2394 185
R1610 vdd.n2325 vdd.n700 185
R1611 vdd.n2484 vdd.n700 185
R1612 vdd.n2324 vdd.n2323 185
R1613 vdd.n2323 vdd.t186 185
R1614 vdd.n2322 vdd.n705 185
R1615 vdd.n2478 vdd.n705 185
R1616 vdd.n1942 vdd.n1941 185
R1617 vdd.n1943 vdd.n1942 185
R1618 vdd.n866 vdd.n864 185
R1619 vdd.n1508 vdd.n864 185
R1620 vdd.n1511 vdd.n1510 185
R1621 vdd.n1510 vdd.n1509 185
R1622 vdd.n869 vdd.n868 185
R1623 vdd.n870 vdd.n869 185
R1624 vdd.n1497 vdd.n1496 185
R1625 vdd.n1498 vdd.n1497 185
R1626 vdd.n878 vdd.n877 185
R1627 vdd.n1489 vdd.n877 185
R1628 vdd.n1492 vdd.n1491 185
R1629 vdd.n1491 vdd.n1490 185
R1630 vdd.n881 vdd.n880 185
R1631 vdd.n888 vdd.n881 185
R1632 vdd.n1480 vdd.n1479 185
R1633 vdd.n1481 vdd.n1480 185
R1634 vdd.n890 vdd.n889 185
R1635 vdd.n889 vdd.n887 185
R1636 vdd.n1475 vdd.n1474 185
R1637 vdd.n1474 vdd.n1473 185
R1638 vdd.n1163 vdd.n1162 185
R1639 vdd.n1164 vdd.n1163 185
R1640 vdd.n1464 vdd.n1463 185
R1641 vdd.n1465 vdd.n1464 185
R1642 vdd.n1171 vdd.n1170 185
R1643 vdd.n1455 vdd.n1170 185
R1644 vdd.n1458 vdd.n1457 185
R1645 vdd.n1457 vdd.n1456 185
R1646 vdd.n1174 vdd.n1173 185
R1647 vdd.n1180 vdd.n1174 185
R1648 vdd.n1446 vdd.n1445 185
R1649 vdd.n1447 vdd.n1446 185
R1650 vdd.n1182 vdd.n1181 185
R1651 vdd.n1438 vdd.n1181 185
R1652 vdd.n1441 vdd.n1440 185
R1653 vdd.n1440 vdd.n1439 185
R1654 vdd.n1185 vdd.n1184 185
R1655 vdd.n1186 vdd.n1185 185
R1656 vdd.n1429 vdd.n1428 185
R1657 vdd.n1430 vdd.n1429 185
R1658 vdd.n1193 vdd.n1192 185
R1659 vdd.n1228 vdd.n1192 185
R1660 vdd.n1424 vdd.n1423 185
R1661 vdd.n1196 vdd.n1195 185
R1662 vdd.n1420 vdd.n1419 185
R1663 vdd.n1421 vdd.n1420 185
R1664 vdd.n1230 vdd.n1229 185
R1665 vdd.n1415 vdd.n1232 185
R1666 vdd.n1414 vdd.n1233 185
R1667 vdd.n1413 vdd.n1234 185
R1668 vdd.n1236 vdd.n1235 185
R1669 vdd.n1409 vdd.n1238 185
R1670 vdd.n1408 vdd.n1239 185
R1671 vdd.n1407 vdd.n1240 185
R1672 vdd.n1242 vdd.n1241 185
R1673 vdd.n1403 vdd.n1244 185
R1674 vdd.n1402 vdd.n1245 185
R1675 vdd.n1401 vdd.n1246 185
R1676 vdd.n1248 vdd.n1247 185
R1677 vdd.n1397 vdd.n1250 185
R1678 vdd.n1396 vdd.n1251 185
R1679 vdd.n1395 vdd.n1252 185
R1680 vdd.n1256 vdd.n1253 185
R1681 vdd.n1391 vdd.n1258 185
R1682 vdd.n1390 vdd.n1259 185
R1683 vdd.n1389 vdd.n1260 185
R1684 vdd.n1262 vdd.n1261 185
R1685 vdd.n1385 vdd.n1264 185
R1686 vdd.n1384 vdd.n1265 185
R1687 vdd.n1383 vdd.n1266 185
R1688 vdd.n1268 vdd.n1267 185
R1689 vdd.n1379 vdd.n1270 185
R1690 vdd.n1378 vdd.n1271 185
R1691 vdd.n1377 vdd.n1272 185
R1692 vdd.n1274 vdd.n1273 185
R1693 vdd.n1373 vdd.n1276 185
R1694 vdd.n1372 vdd.n1277 185
R1695 vdd.n1371 vdd.n1278 185
R1696 vdd.n1280 vdd.n1279 185
R1697 vdd.n1367 vdd.n1282 185
R1698 vdd.n1366 vdd.n1283 185
R1699 vdd.n1365 vdd.n1284 185
R1700 vdd.n1286 vdd.n1285 185
R1701 vdd.n1361 vdd.n1288 185
R1702 vdd.n1360 vdd.n1357 185
R1703 vdd.n1356 vdd.n1289 185
R1704 vdd.n1291 vdd.n1290 185
R1705 vdd.n1352 vdd.n1293 185
R1706 vdd.n1351 vdd.n1294 185
R1707 vdd.n1350 vdd.n1295 185
R1708 vdd.n1297 vdd.n1296 185
R1709 vdd.n1346 vdd.n1299 185
R1710 vdd.n1345 vdd.n1300 185
R1711 vdd.n1344 vdd.n1301 185
R1712 vdd.n1303 vdd.n1302 185
R1713 vdd.n1340 vdd.n1305 185
R1714 vdd.n1339 vdd.n1306 185
R1715 vdd.n1338 vdd.n1307 185
R1716 vdd.n1309 vdd.n1308 185
R1717 vdd.n1334 vdd.n1311 185
R1718 vdd.n1333 vdd.n1312 185
R1719 vdd.n1332 vdd.n1313 185
R1720 vdd.n1315 vdd.n1314 185
R1721 vdd.n1328 vdd.n1317 185
R1722 vdd.n1327 vdd.n1318 185
R1723 vdd.n1326 vdd.n1319 185
R1724 vdd.n1323 vdd.n1227 185
R1725 vdd.n1421 vdd.n1227 185
R1726 vdd.n1946 vdd.n1945 185
R1727 vdd.n1950 vdd.n859 185
R1728 vdd.n1613 vdd.n858 185
R1729 vdd.n1616 vdd.n1615 185
R1730 vdd.n1618 vdd.n1617 185
R1731 vdd.n1621 vdd.n1620 185
R1732 vdd.n1623 vdd.n1622 185
R1733 vdd.n1625 vdd.n1611 185
R1734 vdd.n1627 vdd.n1626 185
R1735 vdd.n1628 vdd.n1605 185
R1736 vdd.n1630 vdd.n1629 185
R1737 vdd.n1632 vdd.n1603 185
R1738 vdd.n1634 vdd.n1633 185
R1739 vdd.n1635 vdd.n1598 185
R1740 vdd.n1637 vdd.n1636 185
R1741 vdd.n1639 vdd.n1596 185
R1742 vdd.n1641 vdd.n1640 185
R1743 vdd.n1642 vdd.n1592 185
R1744 vdd.n1644 vdd.n1643 185
R1745 vdd.n1646 vdd.n1589 185
R1746 vdd.n1648 vdd.n1647 185
R1747 vdd.n1590 vdd.n1583 185
R1748 vdd.n1652 vdd.n1587 185
R1749 vdd.n1653 vdd.n1579 185
R1750 vdd.n1655 vdd.n1654 185
R1751 vdd.n1657 vdd.n1577 185
R1752 vdd.n1659 vdd.n1658 185
R1753 vdd.n1660 vdd.n1572 185
R1754 vdd.n1662 vdd.n1661 185
R1755 vdd.n1664 vdd.n1570 185
R1756 vdd.n1666 vdd.n1665 185
R1757 vdd.n1667 vdd.n1565 185
R1758 vdd.n1669 vdd.n1668 185
R1759 vdd.n1671 vdd.n1563 185
R1760 vdd.n1673 vdd.n1672 185
R1761 vdd.n1674 vdd.n1558 185
R1762 vdd.n1676 vdd.n1675 185
R1763 vdd.n1678 vdd.n1556 185
R1764 vdd.n1680 vdd.n1679 185
R1765 vdd.n1681 vdd.n1552 185
R1766 vdd.n1683 vdd.n1682 185
R1767 vdd.n1685 vdd.n1549 185
R1768 vdd.n1687 vdd.n1686 185
R1769 vdd.n1550 vdd.n1543 185
R1770 vdd.n1691 vdd.n1547 185
R1771 vdd.n1692 vdd.n1539 185
R1772 vdd.n1694 vdd.n1693 185
R1773 vdd.n1696 vdd.n1537 185
R1774 vdd.n1698 vdd.n1697 185
R1775 vdd.n1699 vdd.n1532 185
R1776 vdd.n1701 vdd.n1700 185
R1777 vdd.n1703 vdd.n1530 185
R1778 vdd.n1705 vdd.n1704 185
R1779 vdd.n1706 vdd.n1525 185
R1780 vdd.n1708 vdd.n1707 185
R1781 vdd.n1710 vdd.n1524 185
R1782 vdd.n1711 vdd.n1521 185
R1783 vdd.n1714 vdd.n1713 185
R1784 vdd.n1523 vdd.n1519 185
R1785 vdd.n1931 vdd.n1517 185
R1786 vdd.n1933 vdd.n1932 185
R1787 vdd.n1935 vdd.n1515 185
R1788 vdd.n1937 vdd.n1936 185
R1789 vdd.n1938 vdd.n865 185
R1790 vdd.n1944 vdd.n862 185
R1791 vdd.n1944 vdd.n1943 185
R1792 vdd.n873 vdd.n861 185
R1793 vdd.n1508 vdd.n861 185
R1794 vdd.n1507 vdd.n1506 185
R1795 vdd.n1509 vdd.n1507 185
R1796 vdd.n872 vdd.n871 185
R1797 vdd.n871 vdd.n870 185
R1798 vdd.n1500 vdd.n1499 185
R1799 vdd.n1499 vdd.n1498 185
R1800 vdd.n876 vdd.n875 185
R1801 vdd.n1489 vdd.n876 185
R1802 vdd.n1488 vdd.n1487 185
R1803 vdd.n1490 vdd.n1488 185
R1804 vdd.n883 vdd.n882 185
R1805 vdd.n888 vdd.n882 185
R1806 vdd.n1483 vdd.n1482 185
R1807 vdd.n1482 vdd.n1481 185
R1808 vdd.n886 vdd.n885 185
R1809 vdd.n887 vdd.n886 185
R1810 vdd.n1472 vdd.n1471 185
R1811 vdd.n1473 vdd.n1472 185
R1812 vdd.n1166 vdd.n1165 185
R1813 vdd.n1165 vdd.n1164 185
R1814 vdd.n1467 vdd.n1466 185
R1815 vdd.n1466 vdd.n1465 185
R1816 vdd.n1169 vdd.n1168 185
R1817 vdd.n1455 vdd.n1169 185
R1818 vdd.n1454 vdd.n1453 185
R1819 vdd.n1456 vdd.n1454 185
R1820 vdd.n1176 vdd.n1175 185
R1821 vdd.n1180 vdd.n1175 185
R1822 vdd.n1449 vdd.n1448 185
R1823 vdd.n1448 vdd.n1447 185
R1824 vdd.n1179 vdd.n1178 185
R1825 vdd.n1438 vdd.n1179 185
R1826 vdd.n1437 vdd.n1436 185
R1827 vdd.n1439 vdd.n1437 185
R1828 vdd.n1188 vdd.n1187 185
R1829 vdd.n1187 vdd.n1186 185
R1830 vdd.n1432 vdd.n1431 185
R1831 vdd.n1431 vdd.n1430 185
R1832 vdd.n1191 vdd.n1190 185
R1833 vdd.n1228 vdd.n1191 185
R1834 vdd.n746 vdd.n744 185
R1835 vdd.n2146 vdd.n744 185
R1836 vdd.n2068 vdd.n763 185
R1837 vdd.n763 vdd.t184 185
R1838 vdd.n2070 vdd.n2069 185
R1839 vdd.n2071 vdd.n2070 185
R1840 vdd.n2067 vdd.n762 185
R1841 vdd.n1770 vdd.n762 185
R1842 vdd.n2066 vdd.n2065 185
R1843 vdd.n2065 vdd.n2064 185
R1844 vdd.n765 vdd.n764 185
R1845 vdd.n766 vdd.n765 185
R1846 vdd.n2055 vdd.n2054 185
R1847 vdd.n2056 vdd.n2055 185
R1848 vdd.n2053 vdd.n776 185
R1849 vdd.n776 vdd.n773 185
R1850 vdd.n2052 vdd.n2051 185
R1851 vdd.n2051 vdd.n2050 185
R1852 vdd.n778 vdd.n777 185
R1853 vdd.n779 vdd.n778 185
R1854 vdd.n2043 vdd.n2042 185
R1855 vdd.n2044 vdd.n2043 185
R1856 vdd.n2041 vdd.n787 185
R1857 vdd.n792 vdd.n787 185
R1858 vdd.n2040 vdd.n2039 185
R1859 vdd.n2039 vdd.n2038 185
R1860 vdd.n789 vdd.n788 185
R1861 vdd.n798 vdd.n789 185
R1862 vdd.n2031 vdd.n2030 185
R1863 vdd.n2032 vdd.n2031 185
R1864 vdd.n2029 vdd.n799 185
R1865 vdd.n1871 vdd.n799 185
R1866 vdd.n2028 vdd.n2027 185
R1867 vdd.n2027 vdd.n2026 185
R1868 vdd.n801 vdd.n800 185
R1869 vdd.n802 vdd.n801 185
R1870 vdd.n2019 vdd.n2018 185
R1871 vdd.n2020 vdd.n2019 185
R1872 vdd.n2017 vdd.n811 185
R1873 vdd.n811 vdd.n808 185
R1874 vdd.n2016 vdd.n2015 185
R1875 vdd.n2015 vdd.n2014 185
R1876 vdd.n813 vdd.n812 185
R1877 vdd.n823 vdd.n813 185
R1878 vdd.n2006 vdd.n2005 185
R1879 vdd.n2007 vdd.n2006 185
R1880 vdd.n2004 vdd.n824 185
R1881 vdd.n824 vdd.n820 185
R1882 vdd.n2003 vdd.n2002 185
R1883 vdd.n2002 vdd.n2001 185
R1884 vdd.n826 vdd.n825 185
R1885 vdd.n827 vdd.n826 185
R1886 vdd.n1994 vdd.n1993 185
R1887 vdd.n1995 vdd.n1994 185
R1888 vdd.n1992 vdd.n836 185
R1889 vdd.n836 vdd.n833 185
R1890 vdd.n1991 vdd.n1990 185
R1891 vdd.n1990 vdd.n1989 185
R1892 vdd.n838 vdd.n837 185
R1893 vdd.n1726 vdd.n1725 185
R1894 vdd.n1727 vdd.n1723 185
R1895 vdd.n1723 vdd.n839 185
R1896 vdd.n1729 vdd.n1728 185
R1897 vdd.n1731 vdd.n1722 185
R1898 vdd.n1734 vdd.n1733 185
R1899 vdd.n1735 vdd.n1721 185
R1900 vdd.n1737 vdd.n1736 185
R1901 vdd.n1739 vdd.n1720 185
R1902 vdd.n1742 vdd.n1741 185
R1903 vdd.n1743 vdd.n1719 185
R1904 vdd.n1745 vdd.n1744 185
R1905 vdd.n1747 vdd.n1718 185
R1906 vdd.n1750 vdd.n1749 185
R1907 vdd.n1751 vdd.n1717 185
R1908 vdd.n1753 vdd.n1752 185
R1909 vdd.n1755 vdd.n1716 185
R1910 vdd.n1928 vdd.n1756 185
R1911 vdd.n1927 vdd.n1926 185
R1912 vdd.n1924 vdd.n1757 185
R1913 vdd.n1922 vdd.n1921 185
R1914 vdd.n1920 vdd.n1758 185
R1915 vdd.n1919 vdd.n1918 185
R1916 vdd.n1916 vdd.n1759 185
R1917 vdd.n1914 vdd.n1913 185
R1918 vdd.n1912 vdd.n1760 185
R1919 vdd.n1911 vdd.n1910 185
R1920 vdd.n1908 vdd.n1761 185
R1921 vdd.n1906 vdd.n1905 185
R1922 vdd.n1904 vdd.n1762 185
R1923 vdd.n1903 vdd.n1902 185
R1924 vdd.n1900 vdd.n1763 185
R1925 vdd.n1898 vdd.n1897 185
R1926 vdd.n1896 vdd.n1764 185
R1927 vdd.n1895 vdd.n1894 185
R1928 vdd.n2149 vdd.n2148 185
R1929 vdd.n2151 vdd.n2150 185
R1930 vdd.n2153 vdd.n2152 185
R1931 vdd.n2156 vdd.n2155 185
R1932 vdd.n2158 vdd.n2157 185
R1933 vdd.n2160 vdd.n2159 185
R1934 vdd.n2162 vdd.n2161 185
R1935 vdd.n2164 vdd.n2163 185
R1936 vdd.n2166 vdd.n2165 185
R1937 vdd.n2168 vdd.n2167 185
R1938 vdd.n2170 vdd.n2169 185
R1939 vdd.n2172 vdd.n2171 185
R1940 vdd.n2174 vdd.n2173 185
R1941 vdd.n2176 vdd.n2175 185
R1942 vdd.n2178 vdd.n2177 185
R1943 vdd.n2180 vdd.n2179 185
R1944 vdd.n2182 vdd.n2181 185
R1945 vdd.n2184 vdd.n2183 185
R1946 vdd.n2186 vdd.n2185 185
R1947 vdd.n2188 vdd.n2187 185
R1948 vdd.n2190 vdd.n2189 185
R1949 vdd.n2192 vdd.n2191 185
R1950 vdd.n2194 vdd.n2193 185
R1951 vdd.n2196 vdd.n2195 185
R1952 vdd.n2198 vdd.n2197 185
R1953 vdd.n2200 vdd.n2199 185
R1954 vdd.n2202 vdd.n2201 185
R1955 vdd.n2204 vdd.n2203 185
R1956 vdd.n2206 vdd.n2205 185
R1957 vdd.n2208 vdd.n2207 185
R1958 vdd.n2210 vdd.n2209 185
R1959 vdd.n2212 vdd.n2211 185
R1960 vdd.n2214 vdd.n2213 185
R1961 vdd.n2215 vdd.n745 185
R1962 vdd.n2217 vdd.n2216 185
R1963 vdd.n2218 vdd.n2217 185
R1964 vdd.n2147 vdd.n749 185
R1965 vdd.n2147 vdd.n2146 185
R1966 vdd.n1768 vdd.n750 185
R1967 vdd.t184 vdd.n750 185
R1968 vdd.n1769 vdd.n760 185
R1969 vdd.n2071 vdd.n760 185
R1970 vdd.n1772 vdd.n1771 185
R1971 vdd.n1771 vdd.n1770 185
R1972 vdd.n1773 vdd.n767 185
R1973 vdd.n2064 vdd.n767 185
R1974 vdd.n1775 vdd.n1774 185
R1975 vdd.n1774 vdd.n766 185
R1976 vdd.n1776 vdd.n774 185
R1977 vdd.n2056 vdd.n774 185
R1978 vdd.n1778 vdd.n1777 185
R1979 vdd.n1777 vdd.n773 185
R1980 vdd.n1779 vdd.n780 185
R1981 vdd.n2050 vdd.n780 185
R1982 vdd.n1781 vdd.n1780 185
R1983 vdd.n1780 vdd.n779 185
R1984 vdd.n1782 vdd.n785 185
R1985 vdd.n2044 vdd.n785 185
R1986 vdd.n1784 vdd.n1783 185
R1987 vdd.n1783 vdd.n792 185
R1988 vdd.n1785 vdd.n790 185
R1989 vdd.n2038 vdd.n790 185
R1990 vdd.n1787 vdd.n1786 185
R1991 vdd.n1786 vdd.n798 185
R1992 vdd.n1788 vdd.n796 185
R1993 vdd.n2032 vdd.n796 185
R1994 vdd.n1873 vdd.n1872 185
R1995 vdd.n1872 vdd.n1871 185
R1996 vdd.n1874 vdd.n803 185
R1997 vdd.n2026 vdd.n803 185
R1998 vdd.n1876 vdd.n1875 185
R1999 vdd.n1875 vdd.n802 185
R2000 vdd.n1877 vdd.n809 185
R2001 vdd.n2020 vdd.n809 185
R2002 vdd.n1879 vdd.n1878 185
R2003 vdd.n1878 vdd.n808 185
R2004 vdd.n1880 vdd.n814 185
R2005 vdd.n2014 vdd.n814 185
R2006 vdd.n1882 vdd.n1881 185
R2007 vdd.n1881 vdd.n823 185
R2008 vdd.n1883 vdd.n821 185
R2009 vdd.n2007 vdd.n821 185
R2010 vdd.n1885 vdd.n1884 185
R2011 vdd.n1884 vdd.n820 185
R2012 vdd.n1886 vdd.n828 185
R2013 vdd.n2001 vdd.n828 185
R2014 vdd.n1888 vdd.n1887 185
R2015 vdd.n1887 vdd.n827 185
R2016 vdd.n1889 vdd.n834 185
R2017 vdd.n1995 vdd.n834 185
R2018 vdd.n1891 vdd.n1890 185
R2019 vdd.n1890 vdd.n833 185
R2020 vdd.n1892 vdd.n840 185
R2021 vdd.n1989 vdd.n840 185
R2022 vdd.n3024 vdd.n3023 185
R2023 vdd.n3025 vdd.n3024 185
R2024 vdd.n325 vdd.n324 185
R2025 vdd.n3026 vdd.n325 185
R2026 vdd.n3029 vdd.n3028 185
R2027 vdd.n3028 vdd.n3027 185
R2028 vdd.n3030 vdd.n319 185
R2029 vdd.n319 vdd.n318 185
R2030 vdd.n3032 vdd.n3031 185
R2031 vdd.n3033 vdd.n3032 185
R2032 vdd.n314 vdd.n313 185
R2033 vdd.n3034 vdd.n314 185
R2034 vdd.n3037 vdd.n3036 185
R2035 vdd.n3036 vdd.n3035 185
R2036 vdd.n3038 vdd.n309 185
R2037 vdd.n309 vdd.n308 185
R2038 vdd.n3040 vdd.n3039 185
R2039 vdd.n3041 vdd.n3040 185
R2040 vdd.n303 vdd.n301 185
R2041 vdd.n3042 vdd.n303 185
R2042 vdd.n3045 vdd.n3044 185
R2043 vdd.n3044 vdd.n3043 185
R2044 vdd.n302 vdd.n300 185
R2045 vdd.n304 vdd.n302 185
R2046 vdd.n2881 vdd.n2880 185
R2047 vdd.n2882 vdd.n2881 185
R2048 vdd.n458 vdd.n457 185
R2049 vdd.n457 vdd.n456 185
R2050 vdd.n2876 vdd.n2875 185
R2051 vdd.n2875 vdd.n2874 185
R2052 vdd.n461 vdd.n460 185
R2053 vdd.n467 vdd.n461 185
R2054 vdd.n2865 vdd.n2864 185
R2055 vdd.n2866 vdd.n2865 185
R2056 vdd.n469 vdd.n468 185
R2057 vdd.n2857 vdd.n468 185
R2058 vdd.n2860 vdd.n2859 185
R2059 vdd.n2859 vdd.n2858 185
R2060 vdd.n472 vdd.n471 185
R2061 vdd.n473 vdd.n472 185
R2062 vdd.n2848 vdd.n2847 185
R2063 vdd.n2849 vdd.n2848 185
R2064 vdd.n480 vdd.n479 185
R2065 vdd.n516 vdd.n479 185
R2066 vdd.n2843 vdd.n2842 185
R2067 vdd.n483 vdd.n482 185
R2068 vdd.n2839 vdd.n2838 185
R2069 vdd.n2840 vdd.n2839 185
R2070 vdd.n518 vdd.n517 185
R2071 vdd.n522 vdd.n521 185
R2072 vdd.n2834 vdd.n523 185
R2073 vdd.n2833 vdd.n2832 185
R2074 vdd.n2831 vdd.n2830 185
R2075 vdd.n2829 vdd.n2828 185
R2076 vdd.n2827 vdd.n2826 185
R2077 vdd.n2825 vdd.n2824 185
R2078 vdd.n2823 vdd.n2822 185
R2079 vdd.n2821 vdd.n2820 185
R2080 vdd.n2819 vdd.n2818 185
R2081 vdd.n2817 vdd.n2816 185
R2082 vdd.n2815 vdd.n2814 185
R2083 vdd.n2813 vdd.n2812 185
R2084 vdd.n2811 vdd.n2810 185
R2085 vdd.n2809 vdd.n2808 185
R2086 vdd.n2807 vdd.n2806 185
R2087 vdd.n2798 vdd.n536 185
R2088 vdd.n2800 vdd.n2799 185
R2089 vdd.n2797 vdd.n2796 185
R2090 vdd.n2795 vdd.n2794 185
R2091 vdd.n2793 vdd.n2792 185
R2092 vdd.n2791 vdd.n2790 185
R2093 vdd.n2789 vdd.n2788 185
R2094 vdd.n2787 vdd.n2786 185
R2095 vdd.n2785 vdd.n2784 185
R2096 vdd.n2783 vdd.n2782 185
R2097 vdd.n2781 vdd.n2780 185
R2098 vdd.n2779 vdd.n2778 185
R2099 vdd.n2777 vdd.n2776 185
R2100 vdd.n2775 vdd.n2774 185
R2101 vdd.n2773 vdd.n2772 185
R2102 vdd.n2771 vdd.n2770 185
R2103 vdd.n2769 vdd.n2768 185
R2104 vdd.n2767 vdd.n2766 185
R2105 vdd.n2765 vdd.n2764 185
R2106 vdd.n2763 vdd.n2762 185
R2107 vdd.n2761 vdd.n2760 185
R2108 vdd.n2759 vdd.n2758 185
R2109 vdd.n2752 vdd.n556 185
R2110 vdd.n2754 vdd.n2753 185
R2111 vdd.n2751 vdd.n2750 185
R2112 vdd.n2749 vdd.n2748 185
R2113 vdd.n2747 vdd.n2746 185
R2114 vdd.n2745 vdd.n2744 185
R2115 vdd.n2743 vdd.n2742 185
R2116 vdd.n2741 vdd.n2740 185
R2117 vdd.n2739 vdd.n2738 185
R2118 vdd.n2737 vdd.n2736 185
R2119 vdd.n2735 vdd.n2734 185
R2120 vdd.n2733 vdd.n2732 185
R2121 vdd.n2731 vdd.n2730 185
R2122 vdd.n2729 vdd.n2728 185
R2123 vdd.n2727 vdd.n2726 185
R2124 vdd.n2725 vdd.n2724 185
R2125 vdd.n2723 vdd.n2722 185
R2126 vdd.n2721 vdd.n2720 185
R2127 vdd.n2719 vdd.n2718 185
R2128 vdd.n2717 vdd.n2716 185
R2129 vdd.n2715 vdd.n2714 185
R2130 vdd.n2710 vdd.n515 185
R2131 vdd.n2840 vdd.n515 185
R2132 vdd.n2907 vdd.n2906 185
R2133 vdd.n2911 vdd.n440 185
R2134 vdd.n2913 vdd.n2912 185
R2135 vdd.n2915 vdd.n438 185
R2136 vdd.n2917 vdd.n2916 185
R2137 vdd.n2918 vdd.n433 185
R2138 vdd.n2920 vdd.n2919 185
R2139 vdd.n2922 vdd.n431 185
R2140 vdd.n2924 vdd.n2923 185
R2141 vdd.n2925 vdd.n426 185
R2142 vdd.n2927 vdd.n2926 185
R2143 vdd.n2929 vdd.n424 185
R2144 vdd.n2931 vdd.n2930 185
R2145 vdd.n2932 vdd.n419 185
R2146 vdd.n2934 vdd.n2933 185
R2147 vdd.n2936 vdd.n417 185
R2148 vdd.n2938 vdd.n2937 185
R2149 vdd.n2939 vdd.n413 185
R2150 vdd.n2941 vdd.n2940 185
R2151 vdd.n2943 vdd.n410 185
R2152 vdd.n2945 vdd.n2944 185
R2153 vdd.n411 vdd.n404 185
R2154 vdd.n2949 vdd.n408 185
R2155 vdd.n2950 vdd.n400 185
R2156 vdd.n2952 vdd.n2951 185
R2157 vdd.n2954 vdd.n398 185
R2158 vdd.n2956 vdd.n2955 185
R2159 vdd.n2957 vdd.n393 185
R2160 vdd.n2959 vdd.n2958 185
R2161 vdd.n2961 vdd.n391 185
R2162 vdd.n2963 vdd.n2962 185
R2163 vdd.n2964 vdd.n386 185
R2164 vdd.n2966 vdd.n2965 185
R2165 vdd.n2968 vdd.n384 185
R2166 vdd.n2970 vdd.n2969 185
R2167 vdd.n2971 vdd.n379 185
R2168 vdd.n2973 vdd.n2972 185
R2169 vdd.n2975 vdd.n377 185
R2170 vdd.n2977 vdd.n2976 185
R2171 vdd.n2978 vdd.n373 185
R2172 vdd.n2980 vdd.n2979 185
R2173 vdd.n2982 vdd.n370 185
R2174 vdd.n2984 vdd.n2983 185
R2175 vdd.n371 vdd.n364 185
R2176 vdd.n2988 vdd.n368 185
R2177 vdd.n2989 vdd.n360 185
R2178 vdd.n2991 vdd.n2990 185
R2179 vdd.n2993 vdd.n358 185
R2180 vdd.n2995 vdd.n2994 185
R2181 vdd.n2996 vdd.n353 185
R2182 vdd.n2998 vdd.n2997 185
R2183 vdd.n3000 vdd.n351 185
R2184 vdd.n3002 vdd.n3001 185
R2185 vdd.n3003 vdd.n346 185
R2186 vdd.n3005 vdd.n3004 185
R2187 vdd.n3007 vdd.n344 185
R2188 vdd.n3009 vdd.n3008 185
R2189 vdd.n3010 vdd.n338 185
R2190 vdd.n3012 vdd.n3011 185
R2191 vdd.n3014 vdd.n337 185
R2192 vdd.n3015 vdd.n336 185
R2193 vdd.n3018 vdd.n3017 185
R2194 vdd.n3019 vdd.n334 185
R2195 vdd.n3020 vdd.n330 185
R2196 vdd.n2902 vdd.n328 185
R2197 vdd.n3025 vdd.n328 185
R2198 vdd.n2901 vdd.n327 185
R2199 vdd.n3026 vdd.n327 185
R2200 vdd.n2900 vdd.n326 185
R2201 vdd.n3027 vdd.n326 185
R2202 vdd.n446 vdd.n445 185
R2203 vdd.n445 vdd.n318 185
R2204 vdd.n2896 vdd.n317 185
R2205 vdd.n3033 vdd.n317 185
R2206 vdd.n2895 vdd.n316 185
R2207 vdd.n3034 vdd.n316 185
R2208 vdd.n2894 vdd.n315 185
R2209 vdd.n3035 vdd.n315 185
R2210 vdd.n449 vdd.n448 185
R2211 vdd.n448 vdd.n308 185
R2212 vdd.n2890 vdd.n307 185
R2213 vdd.n3041 vdd.n307 185
R2214 vdd.n2889 vdd.n306 185
R2215 vdd.n3042 vdd.n306 185
R2216 vdd.n2888 vdd.n305 185
R2217 vdd.n3043 vdd.n305 185
R2218 vdd.n455 vdd.n451 185
R2219 vdd.n455 vdd.n304 185
R2220 vdd.n2884 vdd.n2883 185
R2221 vdd.n2883 vdd.n2882 185
R2222 vdd.n454 vdd.n453 185
R2223 vdd.n456 vdd.n454 185
R2224 vdd.n2873 vdd.n2872 185
R2225 vdd.n2874 vdd.n2873 185
R2226 vdd.n463 vdd.n462 185
R2227 vdd.n467 vdd.n462 185
R2228 vdd.n2868 vdd.n2867 185
R2229 vdd.n2867 vdd.n2866 185
R2230 vdd.n466 vdd.n465 185
R2231 vdd.n2857 vdd.n466 185
R2232 vdd.n2856 vdd.n2855 185
R2233 vdd.n2858 vdd.n2856 185
R2234 vdd.n475 vdd.n474 185
R2235 vdd.n474 vdd.n473 185
R2236 vdd.n2851 vdd.n2850 185
R2237 vdd.n2850 vdd.n2849 185
R2238 vdd.n478 vdd.n477 185
R2239 vdd.n516 vdd.n478 185
R2240 vdd.n703 vdd.n702 185
R2241 vdd.n2469 vdd.n2468 185
R2242 vdd.n2467 vdd.n2252 185
R2243 vdd.n2471 vdd.n2252 185
R2244 vdd.n2466 vdd.n2465 185
R2245 vdd.n2464 vdd.n2463 185
R2246 vdd.n2462 vdd.n2461 185
R2247 vdd.n2460 vdd.n2459 185
R2248 vdd.n2458 vdd.n2457 185
R2249 vdd.n2456 vdd.n2455 185
R2250 vdd.n2454 vdd.n2453 185
R2251 vdd.n2452 vdd.n2451 185
R2252 vdd.n2450 vdd.n2449 185
R2253 vdd.n2448 vdd.n2447 185
R2254 vdd.n2446 vdd.n2445 185
R2255 vdd.n2444 vdd.n2443 185
R2256 vdd.n2442 vdd.n2441 185
R2257 vdd.n2440 vdd.n2439 185
R2258 vdd.n2438 vdd.n2437 185
R2259 vdd.n2436 vdd.n2435 185
R2260 vdd.n2434 vdd.n2433 185
R2261 vdd.n2432 vdd.n2431 185
R2262 vdd.n2430 vdd.n2429 185
R2263 vdd.n2428 vdd.n2427 185
R2264 vdd.n2426 vdd.n2425 185
R2265 vdd.n2424 vdd.n2423 185
R2266 vdd.n2422 vdd.n2421 185
R2267 vdd.n2420 vdd.n2419 185
R2268 vdd.n2418 vdd.n2417 185
R2269 vdd.n2416 vdd.n2415 185
R2270 vdd.n2414 vdd.n2413 185
R2271 vdd.n2412 vdd.n2411 185
R2272 vdd.n2410 vdd.n2409 185
R2273 vdd.n2407 vdd.n2406 185
R2274 vdd.n2405 vdd.n2404 185
R2275 vdd.n2403 vdd.n2402 185
R2276 vdd.n2609 vdd.n2608 185
R2277 vdd.n2611 vdd.n624 185
R2278 vdd.n2613 vdd.n2612 185
R2279 vdd.n2615 vdd.n621 185
R2280 vdd.n2617 vdd.n2616 185
R2281 vdd.n2619 vdd.n619 185
R2282 vdd.n2621 vdd.n2620 185
R2283 vdd.n2622 vdd.n618 185
R2284 vdd.n2624 vdd.n2623 185
R2285 vdd.n2626 vdd.n616 185
R2286 vdd.n2628 vdd.n2627 185
R2287 vdd.n2629 vdd.n615 185
R2288 vdd.n2631 vdd.n2630 185
R2289 vdd.n2633 vdd.n613 185
R2290 vdd.n2635 vdd.n2634 185
R2291 vdd.n2636 vdd.n612 185
R2292 vdd.n2638 vdd.n2637 185
R2293 vdd.n2640 vdd.n520 185
R2294 vdd.n2642 vdd.n2641 185
R2295 vdd.n2644 vdd.n610 185
R2296 vdd.n2646 vdd.n2645 185
R2297 vdd.n2647 vdd.n609 185
R2298 vdd.n2649 vdd.n2648 185
R2299 vdd.n2651 vdd.n607 185
R2300 vdd.n2653 vdd.n2652 185
R2301 vdd.n2654 vdd.n606 185
R2302 vdd.n2656 vdd.n2655 185
R2303 vdd.n2658 vdd.n604 185
R2304 vdd.n2660 vdd.n2659 185
R2305 vdd.n2661 vdd.n603 185
R2306 vdd.n2663 vdd.n2662 185
R2307 vdd.n2665 vdd.n602 185
R2308 vdd.n2666 vdd.n601 185
R2309 vdd.n2669 vdd.n2668 185
R2310 vdd.n2670 vdd.n599 185
R2311 vdd.n599 vdd.n484 185
R2312 vdd.n2607 vdd.n596 185
R2313 vdd.n2673 vdd.n596 185
R2314 vdd.n2606 vdd.n2605 185
R2315 vdd.n2605 vdd.n595 185
R2316 vdd.n2604 vdd.n626 185
R2317 vdd.n2604 vdd.n2603 185
R2318 vdd.n2358 vdd.n627 185
R2319 vdd.n636 vdd.n627 185
R2320 vdd.n2359 vdd.n634 185
R2321 vdd.n2597 vdd.n634 185
R2322 vdd.n2361 vdd.n2360 185
R2323 vdd.n2360 vdd.n633 185
R2324 vdd.n2362 vdd.n642 185
R2325 vdd.n2546 vdd.n642 185
R2326 vdd.n2364 vdd.n2363 185
R2327 vdd.n2363 vdd.n641 185
R2328 vdd.n2365 vdd.n648 185
R2329 vdd.n2540 vdd.n648 185
R2330 vdd.n2367 vdd.n2366 185
R2331 vdd.n2366 vdd.n647 185
R2332 vdd.n2368 vdd.n653 185
R2333 vdd.n2532 vdd.n653 185
R2334 vdd.n2370 vdd.n2369 185
R2335 vdd.n2369 vdd.n660 185
R2336 vdd.n2371 vdd.n658 185
R2337 vdd.n2526 vdd.n658 185
R2338 vdd.n2373 vdd.n2372 185
R2339 vdd.n2374 vdd.n2373 185
R2340 vdd.n2357 vdd.n665 185
R2341 vdd.n2520 vdd.n665 185
R2342 vdd.n2356 vdd.n2355 185
R2343 vdd.n2355 vdd.n664 185
R2344 vdd.n2354 vdd.n671 185
R2345 vdd.n2514 vdd.n671 185
R2346 vdd.n2353 vdd.n2352 185
R2347 vdd.n2352 vdd.n670 185
R2348 vdd.n2351 vdd.n676 185
R2349 vdd.n2508 vdd.n676 185
R2350 vdd.n2350 vdd.n2349 185
R2351 vdd.n2349 vdd.n683 185
R2352 vdd.n2348 vdd.n681 185
R2353 vdd.n2502 vdd.n681 185
R2354 vdd.n2347 vdd.n2346 185
R2355 vdd.n2346 vdd.n690 185
R2356 vdd.n2345 vdd.n688 185
R2357 vdd.n2496 vdd.n688 185
R2358 vdd.n2344 vdd.n2343 185
R2359 vdd.n2343 vdd.n687 185
R2360 vdd.n2255 vdd.n694 185
R2361 vdd.n2490 vdd.n694 185
R2362 vdd.n2397 vdd.n2396 185
R2363 vdd.n2396 vdd.n2395 185
R2364 vdd.n2398 vdd.n699 185
R2365 vdd.n2484 vdd.n699 185
R2366 vdd.n2400 vdd.n2399 185
R2367 vdd.n2399 vdd.t186 185
R2368 vdd.n2401 vdd.n704 185
R2369 vdd.n2478 vdd.n704 185
R2370 vdd.n2480 vdd.n2479 185
R2371 vdd.n2479 vdd.n2478 185
R2372 vdd.n2481 vdd.n701 185
R2373 vdd.n701 vdd.t186 185
R2374 vdd.n2483 vdd.n2482 185
R2375 vdd.n2484 vdd.n2483 185
R2376 vdd.n693 vdd.n692 185
R2377 vdd.n2395 vdd.n693 185
R2378 vdd.n2492 vdd.n2491 185
R2379 vdd.n2491 vdd.n2490 185
R2380 vdd.n2493 vdd.n691 185
R2381 vdd.n691 vdd.n687 185
R2382 vdd.n2495 vdd.n2494 185
R2383 vdd.n2496 vdd.n2495 185
R2384 vdd.n680 vdd.n679 185
R2385 vdd.n690 vdd.n680 185
R2386 vdd.n2504 vdd.n2503 185
R2387 vdd.n2503 vdd.n2502 185
R2388 vdd.n2505 vdd.n678 185
R2389 vdd.n683 vdd.n678 185
R2390 vdd.n2507 vdd.n2506 185
R2391 vdd.n2508 vdd.n2507 185
R2392 vdd.n669 vdd.n668 185
R2393 vdd.n670 vdd.n669 185
R2394 vdd.n2516 vdd.n2515 185
R2395 vdd.n2515 vdd.n2514 185
R2396 vdd.n2517 vdd.n667 185
R2397 vdd.n667 vdd.n664 185
R2398 vdd.n2519 vdd.n2518 185
R2399 vdd.n2520 vdd.n2519 185
R2400 vdd.n657 vdd.n656 185
R2401 vdd.n2374 vdd.n657 185
R2402 vdd.n2528 vdd.n2527 185
R2403 vdd.n2527 vdd.n2526 185
R2404 vdd.n2529 vdd.n655 185
R2405 vdd.n660 vdd.n655 185
R2406 vdd.n2531 vdd.n2530 185
R2407 vdd.n2532 vdd.n2531 185
R2408 vdd.n646 vdd.n645 185
R2409 vdd.n647 vdd.n646 185
R2410 vdd.n2542 vdd.n2541 185
R2411 vdd.n2541 vdd.n2540 185
R2412 vdd.n2543 vdd.n644 185
R2413 vdd.n644 vdd.n641 185
R2414 vdd.n2545 vdd.n2544 185
R2415 vdd.n2546 vdd.n2545 185
R2416 vdd.n632 vdd.n631 185
R2417 vdd.n633 vdd.n632 185
R2418 vdd.n2599 vdd.n2598 185
R2419 vdd.n2598 vdd.n2597 185
R2420 vdd.n2600 vdd.n630 185
R2421 vdd.n636 vdd.n630 185
R2422 vdd.n2602 vdd.n2601 185
R2423 vdd.n2603 vdd.n2602 185
R2424 vdd.n600 vdd.n598 185
R2425 vdd.n598 vdd.n595 185
R2426 vdd.n2672 vdd.n2671 185
R2427 vdd.n2673 vdd.n2672 185
R2428 vdd.n2145 vdd.n2144 185
R2429 vdd.n2146 vdd.n2145 185
R2430 vdd.n754 vdd.n752 185
R2431 vdd.n752 vdd.t184 185
R2432 vdd.n2060 vdd.n761 185
R2433 vdd.n2071 vdd.n761 185
R2434 vdd.n2061 vdd.n770 185
R2435 vdd.n1770 vdd.n770 185
R2436 vdd.n2063 vdd.n2062 185
R2437 vdd.n2064 vdd.n2063 185
R2438 vdd.n2059 vdd.n769 185
R2439 vdd.n769 vdd.n766 185
R2440 vdd.n2058 vdd.n2057 185
R2441 vdd.n2057 vdd.n2056 185
R2442 vdd.n772 vdd.n771 185
R2443 vdd.n773 vdd.n772 185
R2444 vdd.n2049 vdd.n2048 185
R2445 vdd.n2050 vdd.n2049 185
R2446 vdd.n2047 vdd.n782 185
R2447 vdd.n782 vdd.n779 185
R2448 vdd.n2046 vdd.n2045 185
R2449 vdd.n2045 vdd.n2044 185
R2450 vdd.n784 vdd.n783 185
R2451 vdd.n792 vdd.n784 185
R2452 vdd.n2037 vdd.n2036 185
R2453 vdd.n2038 vdd.n2037 185
R2454 vdd.n2035 vdd.n793 185
R2455 vdd.n798 vdd.n793 185
R2456 vdd.n2034 vdd.n2033 185
R2457 vdd.n2033 vdd.n2032 185
R2458 vdd.n795 vdd.n794 185
R2459 vdd.n1871 vdd.n795 185
R2460 vdd.n2025 vdd.n2024 185
R2461 vdd.n2026 vdd.n2025 185
R2462 vdd.n2023 vdd.n805 185
R2463 vdd.n805 vdd.n802 185
R2464 vdd.n2022 vdd.n2021 185
R2465 vdd.n2021 vdd.n2020 185
R2466 vdd.n807 vdd.n806 185
R2467 vdd.n808 vdd.n807 185
R2468 vdd.n2013 vdd.n2012 185
R2469 vdd.n2014 vdd.n2013 185
R2470 vdd.n2010 vdd.n816 185
R2471 vdd.n823 vdd.n816 185
R2472 vdd.n2009 vdd.n2008 185
R2473 vdd.n2008 vdd.n2007 185
R2474 vdd.n819 vdd.n818 185
R2475 vdd.n820 vdd.n819 185
R2476 vdd.n2000 vdd.n1999 185
R2477 vdd.n2001 vdd.n2000 185
R2478 vdd.n1998 vdd.n830 185
R2479 vdd.n830 vdd.n827 185
R2480 vdd.n1997 vdd.n1996 185
R2481 vdd.n1996 vdd.n1995 185
R2482 vdd.n832 vdd.n831 185
R2483 vdd.n833 vdd.n832 185
R2484 vdd.n1988 vdd.n1987 185
R2485 vdd.n1989 vdd.n1988 185
R2486 vdd.n2076 vdd.n726 185
R2487 vdd.n2218 vdd.n726 185
R2488 vdd.n2078 vdd.n2077 185
R2489 vdd.n2080 vdd.n2079 185
R2490 vdd.n2082 vdd.n2081 185
R2491 vdd.n2084 vdd.n2083 185
R2492 vdd.n2086 vdd.n2085 185
R2493 vdd.n2088 vdd.n2087 185
R2494 vdd.n2090 vdd.n2089 185
R2495 vdd.n2092 vdd.n2091 185
R2496 vdd.n2094 vdd.n2093 185
R2497 vdd.n2096 vdd.n2095 185
R2498 vdd.n2098 vdd.n2097 185
R2499 vdd.n2100 vdd.n2099 185
R2500 vdd.n2102 vdd.n2101 185
R2501 vdd.n2104 vdd.n2103 185
R2502 vdd.n2106 vdd.n2105 185
R2503 vdd.n2108 vdd.n2107 185
R2504 vdd.n2110 vdd.n2109 185
R2505 vdd.n2112 vdd.n2111 185
R2506 vdd.n2114 vdd.n2113 185
R2507 vdd.n2116 vdd.n2115 185
R2508 vdd.n2118 vdd.n2117 185
R2509 vdd.n2120 vdd.n2119 185
R2510 vdd.n2122 vdd.n2121 185
R2511 vdd.n2124 vdd.n2123 185
R2512 vdd.n2126 vdd.n2125 185
R2513 vdd.n2128 vdd.n2127 185
R2514 vdd.n2130 vdd.n2129 185
R2515 vdd.n2132 vdd.n2131 185
R2516 vdd.n2134 vdd.n2133 185
R2517 vdd.n2136 vdd.n2135 185
R2518 vdd.n2138 vdd.n2137 185
R2519 vdd.n2140 vdd.n2139 185
R2520 vdd.n2142 vdd.n2141 185
R2521 vdd.n2143 vdd.n753 185
R2522 vdd.n2075 vdd.n751 185
R2523 vdd.n2146 vdd.n751 185
R2524 vdd.n2074 vdd.n2073 185
R2525 vdd.n2073 vdd.t184 185
R2526 vdd.n2072 vdd.n758 185
R2527 vdd.n2072 vdd.n2071 185
R2528 vdd.n1852 vdd.n759 185
R2529 vdd.n1770 vdd.n759 185
R2530 vdd.n1853 vdd.n768 185
R2531 vdd.n2064 vdd.n768 185
R2532 vdd.n1855 vdd.n1854 185
R2533 vdd.n1854 vdd.n766 185
R2534 vdd.n1856 vdd.n775 185
R2535 vdd.n2056 vdd.n775 185
R2536 vdd.n1858 vdd.n1857 185
R2537 vdd.n1857 vdd.n773 185
R2538 vdd.n1859 vdd.n781 185
R2539 vdd.n2050 vdd.n781 185
R2540 vdd.n1861 vdd.n1860 185
R2541 vdd.n1860 vdd.n779 185
R2542 vdd.n1862 vdd.n786 185
R2543 vdd.n2044 vdd.n786 185
R2544 vdd.n1864 vdd.n1863 185
R2545 vdd.n1863 vdd.n792 185
R2546 vdd.n1865 vdd.n791 185
R2547 vdd.n2038 vdd.n791 185
R2548 vdd.n1867 vdd.n1866 185
R2549 vdd.n1866 vdd.n798 185
R2550 vdd.n1868 vdd.n797 185
R2551 vdd.n2032 vdd.n797 185
R2552 vdd.n1870 vdd.n1869 185
R2553 vdd.n1871 vdd.n1870 185
R2554 vdd.n1851 vdd.n804 185
R2555 vdd.n2026 vdd.n804 185
R2556 vdd.n1850 vdd.n1849 185
R2557 vdd.n1849 vdd.n802 185
R2558 vdd.n1848 vdd.n810 185
R2559 vdd.n2020 vdd.n810 185
R2560 vdd.n1847 vdd.n1846 185
R2561 vdd.n1846 vdd.n808 185
R2562 vdd.n1845 vdd.n815 185
R2563 vdd.n2014 vdd.n815 185
R2564 vdd.n1844 vdd.n1843 185
R2565 vdd.n1843 vdd.n823 185
R2566 vdd.n1842 vdd.n822 185
R2567 vdd.n2007 vdd.n822 185
R2568 vdd.n1841 vdd.n1840 185
R2569 vdd.n1840 vdd.n820 185
R2570 vdd.n1839 vdd.n829 185
R2571 vdd.n2001 vdd.n829 185
R2572 vdd.n1838 vdd.n1837 185
R2573 vdd.n1837 vdd.n827 185
R2574 vdd.n1836 vdd.n835 185
R2575 vdd.n1995 vdd.n835 185
R2576 vdd.n1835 vdd.n1834 185
R2577 vdd.n1834 vdd.n833 185
R2578 vdd.n1833 vdd.n841 185
R2579 vdd.n1989 vdd.n841 185
R2580 vdd.n1986 vdd.n842 185
R2581 vdd.n1985 vdd.n1984 185
R2582 vdd.n1982 vdd.n843 185
R2583 vdd.n1980 vdd.n1979 185
R2584 vdd.n1978 vdd.n844 185
R2585 vdd.n1977 vdd.n1976 185
R2586 vdd.n1974 vdd.n845 185
R2587 vdd.n1972 vdd.n1971 185
R2588 vdd.n1970 vdd.n846 185
R2589 vdd.n1969 vdd.n1968 185
R2590 vdd.n1966 vdd.n847 185
R2591 vdd.n1964 vdd.n1963 185
R2592 vdd.n1962 vdd.n848 185
R2593 vdd.n1961 vdd.n1960 185
R2594 vdd.n1958 vdd.n849 185
R2595 vdd.n1956 vdd.n1955 185
R2596 vdd.n1954 vdd.n850 185
R2597 vdd.n1953 vdd.n852 185
R2598 vdd.n1798 vdd.n853 185
R2599 vdd.n1801 vdd.n1800 185
R2600 vdd.n1803 vdd.n1802 185
R2601 vdd.n1805 vdd.n1797 185
R2602 vdd.n1808 vdd.n1807 185
R2603 vdd.n1809 vdd.n1796 185
R2604 vdd.n1811 vdd.n1810 185
R2605 vdd.n1813 vdd.n1795 185
R2606 vdd.n1816 vdd.n1815 185
R2607 vdd.n1817 vdd.n1794 185
R2608 vdd.n1819 vdd.n1818 185
R2609 vdd.n1821 vdd.n1793 185
R2610 vdd.n1824 vdd.n1823 185
R2611 vdd.n1825 vdd.n1790 185
R2612 vdd.n1828 vdd.n1827 185
R2613 vdd.n1830 vdd.n1789 185
R2614 vdd.n1832 vdd.n1831 185
R2615 vdd.n1831 vdd.n839 185
R2616 vdd.n291 vdd.n290 171.744
R2617 vdd.n290 vdd.n289 171.744
R2618 vdd.n289 vdd.n258 171.744
R2619 vdd.n282 vdd.n258 171.744
R2620 vdd.n282 vdd.n281 171.744
R2621 vdd.n281 vdd.n263 171.744
R2622 vdd.n274 vdd.n263 171.744
R2623 vdd.n274 vdd.n273 171.744
R2624 vdd.n273 vdd.n267 171.744
R2625 vdd.n244 vdd.n243 171.744
R2626 vdd.n243 vdd.n242 171.744
R2627 vdd.n242 vdd.n211 171.744
R2628 vdd.n235 vdd.n211 171.744
R2629 vdd.n235 vdd.n234 171.744
R2630 vdd.n234 vdd.n216 171.744
R2631 vdd.n227 vdd.n216 171.744
R2632 vdd.n227 vdd.n226 171.744
R2633 vdd.n226 vdd.n220 171.744
R2634 vdd.n201 vdd.n200 171.744
R2635 vdd.n200 vdd.n199 171.744
R2636 vdd.n199 vdd.n168 171.744
R2637 vdd.n192 vdd.n168 171.744
R2638 vdd.n192 vdd.n191 171.744
R2639 vdd.n191 vdd.n173 171.744
R2640 vdd.n184 vdd.n173 171.744
R2641 vdd.n184 vdd.n183 171.744
R2642 vdd.n183 vdd.n177 171.744
R2643 vdd.n154 vdd.n153 171.744
R2644 vdd.n153 vdd.n152 171.744
R2645 vdd.n152 vdd.n121 171.744
R2646 vdd.n145 vdd.n121 171.744
R2647 vdd.n145 vdd.n144 171.744
R2648 vdd.n144 vdd.n126 171.744
R2649 vdd.n137 vdd.n126 171.744
R2650 vdd.n137 vdd.n136 171.744
R2651 vdd.n136 vdd.n130 171.744
R2652 vdd.n112 vdd.n111 171.744
R2653 vdd.n111 vdd.n110 171.744
R2654 vdd.n110 vdd.n79 171.744
R2655 vdd.n103 vdd.n79 171.744
R2656 vdd.n103 vdd.n102 171.744
R2657 vdd.n102 vdd.n84 171.744
R2658 vdd.n95 vdd.n84 171.744
R2659 vdd.n95 vdd.n94 171.744
R2660 vdd.n94 vdd.n88 171.744
R2661 vdd.n65 vdd.n64 171.744
R2662 vdd.n64 vdd.n63 171.744
R2663 vdd.n63 vdd.n32 171.744
R2664 vdd.n56 vdd.n32 171.744
R2665 vdd.n56 vdd.n55 171.744
R2666 vdd.n55 vdd.n37 171.744
R2667 vdd.n48 vdd.n37 171.744
R2668 vdd.n48 vdd.n47 171.744
R2669 vdd.n47 vdd.n41 171.744
R2670 vdd.n1106 vdd.n1105 171.744
R2671 vdd.n1105 vdd.n1104 171.744
R2672 vdd.n1104 vdd.n1073 171.744
R2673 vdd.n1097 vdd.n1073 171.744
R2674 vdd.n1097 vdd.n1096 171.744
R2675 vdd.n1096 vdd.n1078 171.744
R2676 vdd.n1089 vdd.n1078 171.744
R2677 vdd.n1089 vdd.n1088 171.744
R2678 vdd.n1088 vdd.n1082 171.744
R2679 vdd.n1153 vdd.n1152 171.744
R2680 vdd.n1152 vdd.n1151 171.744
R2681 vdd.n1151 vdd.n1120 171.744
R2682 vdd.n1144 vdd.n1120 171.744
R2683 vdd.n1144 vdd.n1143 171.744
R2684 vdd.n1143 vdd.n1125 171.744
R2685 vdd.n1136 vdd.n1125 171.744
R2686 vdd.n1136 vdd.n1135 171.744
R2687 vdd.n1135 vdd.n1129 171.744
R2688 vdd.n1016 vdd.n1015 171.744
R2689 vdd.n1015 vdd.n1014 171.744
R2690 vdd.n1014 vdd.n983 171.744
R2691 vdd.n1007 vdd.n983 171.744
R2692 vdd.n1007 vdd.n1006 171.744
R2693 vdd.n1006 vdd.n988 171.744
R2694 vdd.n999 vdd.n988 171.744
R2695 vdd.n999 vdd.n998 171.744
R2696 vdd.n998 vdd.n992 171.744
R2697 vdd.n1063 vdd.n1062 171.744
R2698 vdd.n1062 vdd.n1061 171.744
R2699 vdd.n1061 vdd.n1030 171.744
R2700 vdd.n1054 vdd.n1030 171.744
R2701 vdd.n1054 vdd.n1053 171.744
R2702 vdd.n1053 vdd.n1035 171.744
R2703 vdd.n1046 vdd.n1035 171.744
R2704 vdd.n1046 vdd.n1045 171.744
R2705 vdd.n1045 vdd.n1039 171.744
R2706 vdd.n927 vdd.n926 171.744
R2707 vdd.n926 vdd.n925 171.744
R2708 vdd.n925 vdd.n894 171.744
R2709 vdd.n918 vdd.n894 171.744
R2710 vdd.n918 vdd.n917 171.744
R2711 vdd.n917 vdd.n899 171.744
R2712 vdd.n910 vdd.n899 171.744
R2713 vdd.n910 vdd.n909 171.744
R2714 vdd.n909 vdd.n903 171.744
R2715 vdd.n974 vdd.n973 171.744
R2716 vdd.n973 vdd.n972 171.744
R2717 vdd.n972 vdd.n941 171.744
R2718 vdd.n965 vdd.n941 171.744
R2719 vdd.n965 vdd.n964 171.744
R2720 vdd.n964 vdd.n946 171.744
R2721 vdd.n957 vdd.n946 171.744
R2722 vdd.n957 vdd.n956 171.744
R2723 vdd.n956 vdd.n950 171.744
R2724 vdd.n3017 vdd.n334 146.341
R2725 vdd.n3015 vdd.n3014 146.341
R2726 vdd.n3012 vdd.n338 146.341
R2727 vdd.n3008 vdd.n3007 146.341
R2728 vdd.n3005 vdd.n346 146.341
R2729 vdd.n3001 vdd.n3000 146.341
R2730 vdd.n2998 vdd.n353 146.341
R2731 vdd.n2994 vdd.n2993 146.341
R2732 vdd.n2991 vdd.n360 146.341
R2733 vdd.n371 vdd.n368 146.341
R2734 vdd.n2983 vdd.n2982 146.341
R2735 vdd.n2980 vdd.n373 146.341
R2736 vdd.n2976 vdd.n2975 146.341
R2737 vdd.n2973 vdd.n379 146.341
R2738 vdd.n2969 vdd.n2968 146.341
R2739 vdd.n2966 vdd.n386 146.341
R2740 vdd.n2962 vdd.n2961 146.341
R2741 vdd.n2959 vdd.n393 146.341
R2742 vdd.n2955 vdd.n2954 146.341
R2743 vdd.n2952 vdd.n400 146.341
R2744 vdd.n411 vdd.n408 146.341
R2745 vdd.n2944 vdd.n2943 146.341
R2746 vdd.n2941 vdd.n413 146.341
R2747 vdd.n2937 vdd.n2936 146.341
R2748 vdd.n2934 vdd.n419 146.341
R2749 vdd.n2930 vdd.n2929 146.341
R2750 vdd.n2927 vdd.n426 146.341
R2751 vdd.n2923 vdd.n2922 146.341
R2752 vdd.n2920 vdd.n433 146.341
R2753 vdd.n2916 vdd.n2915 146.341
R2754 vdd.n2913 vdd.n440 146.341
R2755 vdd.n2850 vdd.n478 146.341
R2756 vdd.n2850 vdd.n474 146.341
R2757 vdd.n2856 vdd.n474 146.341
R2758 vdd.n2856 vdd.n466 146.341
R2759 vdd.n2867 vdd.n466 146.341
R2760 vdd.n2867 vdd.n462 146.341
R2761 vdd.n2873 vdd.n462 146.341
R2762 vdd.n2873 vdd.n454 146.341
R2763 vdd.n2883 vdd.n454 146.341
R2764 vdd.n2883 vdd.n455 146.341
R2765 vdd.n455 vdd.n305 146.341
R2766 vdd.n306 vdd.n305 146.341
R2767 vdd.n307 vdd.n306 146.341
R2768 vdd.n448 vdd.n307 146.341
R2769 vdd.n448 vdd.n315 146.341
R2770 vdd.n316 vdd.n315 146.341
R2771 vdd.n317 vdd.n316 146.341
R2772 vdd.n445 vdd.n317 146.341
R2773 vdd.n445 vdd.n326 146.341
R2774 vdd.n327 vdd.n326 146.341
R2775 vdd.n328 vdd.n327 146.341
R2776 vdd.n2839 vdd.n483 146.341
R2777 vdd.n2839 vdd.n517 146.341
R2778 vdd.n523 vdd.n522 146.341
R2779 vdd.n2832 vdd.n2831 146.341
R2780 vdd.n2828 vdd.n2827 146.341
R2781 vdd.n2824 vdd.n2823 146.341
R2782 vdd.n2820 vdd.n2819 146.341
R2783 vdd.n2816 vdd.n2815 146.341
R2784 vdd.n2812 vdd.n2811 146.341
R2785 vdd.n2808 vdd.n2807 146.341
R2786 vdd.n2799 vdd.n2798 146.341
R2787 vdd.n2796 vdd.n2795 146.341
R2788 vdd.n2792 vdd.n2791 146.341
R2789 vdd.n2788 vdd.n2787 146.341
R2790 vdd.n2784 vdd.n2783 146.341
R2791 vdd.n2780 vdd.n2779 146.341
R2792 vdd.n2776 vdd.n2775 146.341
R2793 vdd.n2772 vdd.n2771 146.341
R2794 vdd.n2768 vdd.n2767 146.341
R2795 vdd.n2764 vdd.n2763 146.341
R2796 vdd.n2760 vdd.n2759 146.341
R2797 vdd.n2753 vdd.n2752 146.341
R2798 vdd.n2750 vdd.n2749 146.341
R2799 vdd.n2746 vdd.n2745 146.341
R2800 vdd.n2742 vdd.n2741 146.341
R2801 vdd.n2738 vdd.n2737 146.341
R2802 vdd.n2734 vdd.n2733 146.341
R2803 vdd.n2730 vdd.n2729 146.341
R2804 vdd.n2726 vdd.n2725 146.341
R2805 vdd.n2722 vdd.n2721 146.341
R2806 vdd.n2718 vdd.n2717 146.341
R2807 vdd.n2714 vdd.n515 146.341
R2808 vdd.n2848 vdd.n479 146.341
R2809 vdd.n2848 vdd.n472 146.341
R2810 vdd.n2859 vdd.n472 146.341
R2811 vdd.n2859 vdd.n468 146.341
R2812 vdd.n2865 vdd.n468 146.341
R2813 vdd.n2865 vdd.n461 146.341
R2814 vdd.n2875 vdd.n461 146.341
R2815 vdd.n2875 vdd.n457 146.341
R2816 vdd.n2881 vdd.n457 146.341
R2817 vdd.n2881 vdd.n302 146.341
R2818 vdd.n3044 vdd.n302 146.341
R2819 vdd.n3044 vdd.n303 146.341
R2820 vdd.n3040 vdd.n303 146.341
R2821 vdd.n3040 vdd.n309 146.341
R2822 vdd.n3036 vdd.n309 146.341
R2823 vdd.n3036 vdd.n314 146.341
R2824 vdd.n3032 vdd.n314 146.341
R2825 vdd.n3032 vdd.n319 146.341
R2826 vdd.n3028 vdd.n319 146.341
R2827 vdd.n3028 vdd.n325 146.341
R2828 vdd.n3024 vdd.n325 146.341
R2829 vdd.n1936 vdd.n1935 146.341
R2830 vdd.n1933 vdd.n1517 146.341
R2831 vdd.n1713 vdd.n1523 146.341
R2832 vdd.n1711 vdd.n1710 146.341
R2833 vdd.n1708 vdd.n1525 146.341
R2834 vdd.n1704 vdd.n1703 146.341
R2835 vdd.n1701 vdd.n1532 146.341
R2836 vdd.n1697 vdd.n1696 146.341
R2837 vdd.n1694 vdd.n1539 146.341
R2838 vdd.n1550 vdd.n1547 146.341
R2839 vdd.n1686 vdd.n1685 146.341
R2840 vdd.n1683 vdd.n1552 146.341
R2841 vdd.n1679 vdd.n1678 146.341
R2842 vdd.n1676 vdd.n1558 146.341
R2843 vdd.n1672 vdd.n1671 146.341
R2844 vdd.n1669 vdd.n1565 146.341
R2845 vdd.n1665 vdd.n1664 146.341
R2846 vdd.n1662 vdd.n1572 146.341
R2847 vdd.n1658 vdd.n1657 146.341
R2848 vdd.n1655 vdd.n1579 146.341
R2849 vdd.n1590 vdd.n1587 146.341
R2850 vdd.n1647 vdd.n1646 146.341
R2851 vdd.n1644 vdd.n1592 146.341
R2852 vdd.n1640 vdd.n1639 146.341
R2853 vdd.n1637 vdd.n1598 146.341
R2854 vdd.n1633 vdd.n1632 146.341
R2855 vdd.n1630 vdd.n1605 146.341
R2856 vdd.n1626 vdd.n1625 146.341
R2857 vdd.n1623 vdd.n1620 146.341
R2858 vdd.n1618 vdd.n1615 146.341
R2859 vdd.n1613 vdd.n859 146.341
R2860 vdd.n1431 vdd.n1191 146.341
R2861 vdd.n1431 vdd.n1187 146.341
R2862 vdd.n1437 vdd.n1187 146.341
R2863 vdd.n1437 vdd.n1179 146.341
R2864 vdd.n1448 vdd.n1179 146.341
R2865 vdd.n1448 vdd.n1175 146.341
R2866 vdd.n1454 vdd.n1175 146.341
R2867 vdd.n1454 vdd.n1169 146.341
R2868 vdd.n1466 vdd.n1169 146.341
R2869 vdd.n1466 vdd.n1165 146.341
R2870 vdd.n1472 vdd.n1165 146.341
R2871 vdd.n1472 vdd.n886 146.341
R2872 vdd.n1482 vdd.n886 146.341
R2873 vdd.n1482 vdd.n882 146.341
R2874 vdd.n1488 vdd.n882 146.341
R2875 vdd.n1488 vdd.n876 146.341
R2876 vdd.n1499 vdd.n876 146.341
R2877 vdd.n1499 vdd.n871 146.341
R2878 vdd.n1507 vdd.n871 146.341
R2879 vdd.n1507 vdd.n861 146.341
R2880 vdd.n1944 vdd.n861 146.341
R2881 vdd.n1420 vdd.n1196 146.341
R2882 vdd.n1420 vdd.n1229 146.341
R2883 vdd.n1233 vdd.n1232 146.341
R2884 vdd.n1235 vdd.n1234 146.341
R2885 vdd.n1239 vdd.n1238 146.341
R2886 vdd.n1241 vdd.n1240 146.341
R2887 vdd.n1245 vdd.n1244 146.341
R2888 vdd.n1247 vdd.n1246 146.341
R2889 vdd.n1251 vdd.n1250 146.341
R2890 vdd.n1253 vdd.n1252 146.341
R2891 vdd.n1259 vdd.n1258 146.341
R2892 vdd.n1261 vdd.n1260 146.341
R2893 vdd.n1265 vdd.n1264 146.341
R2894 vdd.n1267 vdd.n1266 146.341
R2895 vdd.n1271 vdd.n1270 146.341
R2896 vdd.n1273 vdd.n1272 146.341
R2897 vdd.n1277 vdd.n1276 146.341
R2898 vdd.n1279 vdd.n1278 146.341
R2899 vdd.n1283 vdd.n1282 146.341
R2900 vdd.n1285 vdd.n1284 146.341
R2901 vdd.n1357 vdd.n1288 146.341
R2902 vdd.n1290 vdd.n1289 146.341
R2903 vdd.n1294 vdd.n1293 146.341
R2904 vdd.n1296 vdd.n1295 146.341
R2905 vdd.n1300 vdd.n1299 146.341
R2906 vdd.n1302 vdd.n1301 146.341
R2907 vdd.n1306 vdd.n1305 146.341
R2908 vdd.n1308 vdd.n1307 146.341
R2909 vdd.n1312 vdd.n1311 146.341
R2910 vdd.n1314 vdd.n1313 146.341
R2911 vdd.n1318 vdd.n1317 146.341
R2912 vdd.n1319 vdd.n1227 146.341
R2913 vdd.n1429 vdd.n1192 146.341
R2914 vdd.n1429 vdd.n1185 146.341
R2915 vdd.n1440 vdd.n1185 146.341
R2916 vdd.n1440 vdd.n1181 146.341
R2917 vdd.n1446 vdd.n1181 146.341
R2918 vdd.n1446 vdd.n1174 146.341
R2919 vdd.n1457 vdd.n1174 146.341
R2920 vdd.n1457 vdd.n1170 146.341
R2921 vdd.n1464 vdd.n1170 146.341
R2922 vdd.n1464 vdd.n1163 146.341
R2923 vdd.n1474 vdd.n1163 146.341
R2924 vdd.n1474 vdd.n889 146.341
R2925 vdd.n1480 vdd.n889 146.341
R2926 vdd.n1480 vdd.n881 146.341
R2927 vdd.n1491 vdd.n881 146.341
R2928 vdd.n1491 vdd.n877 146.341
R2929 vdd.n1497 vdd.n877 146.341
R2930 vdd.n1497 vdd.n869 146.341
R2931 vdd.n1510 vdd.n869 146.341
R2932 vdd.n1510 vdd.n864 146.341
R2933 vdd.n1942 vdd.n864 146.341
R2934 vdd.n863 vdd.n839 141.707
R2935 vdd.n2840 vdd.n484 141.707
R2936 vdd.n1791 vdd.t82 127.284
R2937 vdd.n755 vdd.t66 127.284
R2938 vdd.n1765 vdd.t107 127.284
R2939 vdd.n747 vdd.t97 127.284
R2940 vdd.n2536 vdd.t49 127.284
R2941 vdd.n2536 vdd.t50 127.284
R2942 vdd.n2256 vdd.t89 127.284
R2943 vdd.n622 vdd.t70 127.284
R2944 vdd.n2253 vdd.t75 127.284
R2945 vdd.n589 vdd.t77 127.284
R2946 vdd.n817 vdd.t85 127.284
R2947 vdd.n817 vdd.t86 127.284
R2948 vdd.n22 vdd.n20 117.314
R2949 vdd.n17 vdd.n15 117.314
R2950 vdd.n27 vdd.n26 116.927
R2951 vdd.n24 vdd.n23 116.927
R2952 vdd.n22 vdd.n21 116.927
R2953 vdd.n17 vdd.n16 116.927
R2954 vdd.n19 vdd.n18 116.927
R2955 vdd.n27 vdd.n25 116.927
R2956 vdd.n1792 vdd.t81 111.188
R2957 vdd.n756 vdd.t67 111.188
R2958 vdd.n1766 vdd.t106 111.188
R2959 vdd.n748 vdd.t98 111.188
R2960 vdd.n2257 vdd.t88 111.188
R2961 vdd.n623 vdd.t71 111.188
R2962 vdd.n2254 vdd.t74 111.188
R2963 vdd.n590 vdd.t78 111.188
R2964 vdd.n2479 vdd.n701 99.5127
R2965 vdd.n2483 vdd.n701 99.5127
R2966 vdd.n2483 vdd.n693 99.5127
R2967 vdd.n2491 vdd.n693 99.5127
R2968 vdd.n2491 vdd.n691 99.5127
R2969 vdd.n2495 vdd.n691 99.5127
R2970 vdd.n2495 vdd.n680 99.5127
R2971 vdd.n2503 vdd.n680 99.5127
R2972 vdd.n2503 vdd.n678 99.5127
R2973 vdd.n2507 vdd.n678 99.5127
R2974 vdd.n2507 vdd.n669 99.5127
R2975 vdd.n2515 vdd.n669 99.5127
R2976 vdd.n2515 vdd.n667 99.5127
R2977 vdd.n2519 vdd.n667 99.5127
R2978 vdd.n2519 vdd.n657 99.5127
R2979 vdd.n2527 vdd.n657 99.5127
R2980 vdd.n2527 vdd.n655 99.5127
R2981 vdd.n2531 vdd.n655 99.5127
R2982 vdd.n2531 vdd.n646 99.5127
R2983 vdd.n2541 vdd.n646 99.5127
R2984 vdd.n2541 vdd.n644 99.5127
R2985 vdd.n2545 vdd.n644 99.5127
R2986 vdd.n2545 vdd.n632 99.5127
R2987 vdd.n2598 vdd.n632 99.5127
R2988 vdd.n2598 vdd.n630 99.5127
R2989 vdd.n2602 vdd.n630 99.5127
R2990 vdd.n2602 vdd.n598 99.5127
R2991 vdd.n2672 vdd.n598 99.5127
R2992 vdd.n2668 vdd.n599 99.5127
R2993 vdd.n2666 vdd.n2665 99.5127
R2994 vdd.n2663 vdd.n603 99.5127
R2995 vdd.n2659 vdd.n2658 99.5127
R2996 vdd.n2656 vdd.n606 99.5127
R2997 vdd.n2652 vdd.n2651 99.5127
R2998 vdd.n2649 vdd.n609 99.5127
R2999 vdd.n2645 vdd.n2644 99.5127
R3000 vdd.n2642 vdd.n2640 99.5127
R3001 vdd.n2638 vdd.n612 99.5127
R3002 vdd.n2634 vdd.n2633 99.5127
R3003 vdd.n2631 vdd.n615 99.5127
R3004 vdd.n2627 vdd.n2626 99.5127
R3005 vdd.n2624 vdd.n618 99.5127
R3006 vdd.n2620 vdd.n2619 99.5127
R3007 vdd.n2617 vdd.n621 99.5127
R3008 vdd.n2612 vdd.n2611 99.5127
R3009 vdd.n2399 vdd.n704 99.5127
R3010 vdd.n2399 vdd.n699 99.5127
R3011 vdd.n2396 vdd.n699 99.5127
R3012 vdd.n2396 vdd.n694 99.5127
R3013 vdd.n2343 vdd.n694 99.5127
R3014 vdd.n2343 vdd.n688 99.5127
R3015 vdd.n2346 vdd.n688 99.5127
R3016 vdd.n2346 vdd.n681 99.5127
R3017 vdd.n2349 vdd.n681 99.5127
R3018 vdd.n2349 vdd.n676 99.5127
R3019 vdd.n2352 vdd.n676 99.5127
R3020 vdd.n2352 vdd.n671 99.5127
R3021 vdd.n2355 vdd.n671 99.5127
R3022 vdd.n2355 vdd.n665 99.5127
R3023 vdd.n2373 vdd.n665 99.5127
R3024 vdd.n2373 vdd.n658 99.5127
R3025 vdd.n2369 vdd.n658 99.5127
R3026 vdd.n2369 vdd.n653 99.5127
R3027 vdd.n2366 vdd.n653 99.5127
R3028 vdd.n2366 vdd.n648 99.5127
R3029 vdd.n2363 vdd.n648 99.5127
R3030 vdd.n2363 vdd.n642 99.5127
R3031 vdd.n2360 vdd.n642 99.5127
R3032 vdd.n2360 vdd.n634 99.5127
R3033 vdd.n634 vdd.n627 99.5127
R3034 vdd.n2604 vdd.n627 99.5127
R3035 vdd.n2605 vdd.n2604 99.5127
R3036 vdd.n2605 vdd.n596 99.5127
R3037 vdd.n2469 vdd.n2252 99.5127
R3038 vdd.n2465 vdd.n2252 99.5127
R3039 vdd.n2463 vdd.n2462 99.5127
R3040 vdd.n2459 vdd.n2458 99.5127
R3041 vdd.n2455 vdd.n2454 99.5127
R3042 vdd.n2451 vdd.n2450 99.5127
R3043 vdd.n2447 vdd.n2446 99.5127
R3044 vdd.n2443 vdd.n2442 99.5127
R3045 vdd.n2439 vdd.n2438 99.5127
R3046 vdd.n2435 vdd.n2434 99.5127
R3047 vdd.n2431 vdd.n2430 99.5127
R3048 vdd.n2427 vdd.n2426 99.5127
R3049 vdd.n2423 vdd.n2422 99.5127
R3050 vdd.n2419 vdd.n2418 99.5127
R3051 vdd.n2415 vdd.n2414 99.5127
R3052 vdd.n2411 vdd.n2410 99.5127
R3053 vdd.n2406 vdd.n2405 99.5127
R3054 vdd.n2217 vdd.n745 99.5127
R3055 vdd.n2213 vdd.n2212 99.5127
R3056 vdd.n2209 vdd.n2208 99.5127
R3057 vdd.n2205 vdd.n2204 99.5127
R3058 vdd.n2201 vdd.n2200 99.5127
R3059 vdd.n2197 vdd.n2196 99.5127
R3060 vdd.n2193 vdd.n2192 99.5127
R3061 vdd.n2189 vdd.n2188 99.5127
R3062 vdd.n2185 vdd.n2184 99.5127
R3063 vdd.n2181 vdd.n2180 99.5127
R3064 vdd.n2177 vdd.n2176 99.5127
R3065 vdd.n2173 vdd.n2172 99.5127
R3066 vdd.n2169 vdd.n2168 99.5127
R3067 vdd.n2165 vdd.n2164 99.5127
R3068 vdd.n2161 vdd.n2160 99.5127
R3069 vdd.n2157 vdd.n2156 99.5127
R3070 vdd.n2152 vdd.n2151 99.5127
R3071 vdd.n1890 vdd.n840 99.5127
R3072 vdd.n1890 vdd.n834 99.5127
R3073 vdd.n1887 vdd.n834 99.5127
R3074 vdd.n1887 vdd.n828 99.5127
R3075 vdd.n1884 vdd.n828 99.5127
R3076 vdd.n1884 vdd.n821 99.5127
R3077 vdd.n1881 vdd.n821 99.5127
R3078 vdd.n1881 vdd.n814 99.5127
R3079 vdd.n1878 vdd.n814 99.5127
R3080 vdd.n1878 vdd.n809 99.5127
R3081 vdd.n1875 vdd.n809 99.5127
R3082 vdd.n1875 vdd.n803 99.5127
R3083 vdd.n1872 vdd.n803 99.5127
R3084 vdd.n1872 vdd.n796 99.5127
R3085 vdd.n1786 vdd.n796 99.5127
R3086 vdd.n1786 vdd.n790 99.5127
R3087 vdd.n1783 vdd.n790 99.5127
R3088 vdd.n1783 vdd.n785 99.5127
R3089 vdd.n1780 vdd.n785 99.5127
R3090 vdd.n1780 vdd.n780 99.5127
R3091 vdd.n1777 vdd.n780 99.5127
R3092 vdd.n1777 vdd.n774 99.5127
R3093 vdd.n1774 vdd.n774 99.5127
R3094 vdd.n1774 vdd.n767 99.5127
R3095 vdd.n1771 vdd.n767 99.5127
R3096 vdd.n1771 vdd.n760 99.5127
R3097 vdd.n760 vdd.n750 99.5127
R3098 vdd.n2147 vdd.n750 99.5127
R3099 vdd.n1725 vdd.n1723 99.5127
R3100 vdd.n1729 vdd.n1723 99.5127
R3101 vdd.n1733 vdd.n1731 99.5127
R3102 vdd.n1737 vdd.n1721 99.5127
R3103 vdd.n1741 vdd.n1739 99.5127
R3104 vdd.n1745 vdd.n1719 99.5127
R3105 vdd.n1749 vdd.n1747 99.5127
R3106 vdd.n1753 vdd.n1717 99.5127
R3107 vdd.n1756 vdd.n1755 99.5127
R3108 vdd.n1926 vdd.n1924 99.5127
R3109 vdd.n1922 vdd.n1758 99.5127
R3110 vdd.n1918 vdd.n1916 99.5127
R3111 vdd.n1914 vdd.n1760 99.5127
R3112 vdd.n1910 vdd.n1908 99.5127
R3113 vdd.n1906 vdd.n1762 99.5127
R3114 vdd.n1902 vdd.n1900 99.5127
R3115 vdd.n1898 vdd.n1764 99.5127
R3116 vdd.n1990 vdd.n836 99.5127
R3117 vdd.n1994 vdd.n836 99.5127
R3118 vdd.n1994 vdd.n826 99.5127
R3119 vdd.n2002 vdd.n826 99.5127
R3120 vdd.n2002 vdd.n824 99.5127
R3121 vdd.n2006 vdd.n824 99.5127
R3122 vdd.n2006 vdd.n813 99.5127
R3123 vdd.n2015 vdd.n813 99.5127
R3124 vdd.n2015 vdd.n811 99.5127
R3125 vdd.n2019 vdd.n811 99.5127
R3126 vdd.n2019 vdd.n801 99.5127
R3127 vdd.n2027 vdd.n801 99.5127
R3128 vdd.n2027 vdd.n799 99.5127
R3129 vdd.n2031 vdd.n799 99.5127
R3130 vdd.n2031 vdd.n789 99.5127
R3131 vdd.n2039 vdd.n789 99.5127
R3132 vdd.n2039 vdd.n787 99.5127
R3133 vdd.n2043 vdd.n787 99.5127
R3134 vdd.n2043 vdd.n778 99.5127
R3135 vdd.n2051 vdd.n778 99.5127
R3136 vdd.n2051 vdd.n776 99.5127
R3137 vdd.n2055 vdd.n776 99.5127
R3138 vdd.n2055 vdd.n765 99.5127
R3139 vdd.n2065 vdd.n765 99.5127
R3140 vdd.n2065 vdd.n762 99.5127
R3141 vdd.n2070 vdd.n762 99.5127
R3142 vdd.n2070 vdd.n763 99.5127
R3143 vdd.n763 vdd.n744 99.5127
R3144 vdd.n2588 vdd.n2587 99.5127
R3145 vdd.n2585 vdd.n2551 99.5127
R3146 vdd.n2581 vdd.n2580 99.5127
R3147 vdd.n2578 vdd.n2554 99.5127
R3148 vdd.n2574 vdd.n2573 99.5127
R3149 vdd.n2571 vdd.n2557 99.5127
R3150 vdd.n2567 vdd.n2566 99.5127
R3151 vdd.n2564 vdd.n2561 99.5127
R3152 vdd.n2705 vdd.n577 99.5127
R3153 vdd.n2703 vdd.n2702 99.5127
R3154 vdd.n2700 vdd.n579 99.5127
R3155 vdd.n2696 vdd.n2695 99.5127
R3156 vdd.n2693 vdd.n582 99.5127
R3157 vdd.n2689 vdd.n2688 99.5127
R3158 vdd.n2686 vdd.n585 99.5127
R3159 vdd.n2682 vdd.n2681 99.5127
R3160 vdd.n2679 vdd.n588 99.5127
R3161 vdd.n2323 vdd.n705 99.5127
R3162 vdd.n2323 vdd.n700 99.5127
R3163 vdd.n2394 vdd.n700 99.5127
R3164 vdd.n2394 vdd.n695 99.5127
R3165 vdd.n2390 vdd.n695 99.5127
R3166 vdd.n2390 vdd.n689 99.5127
R3167 vdd.n2387 vdd.n689 99.5127
R3168 vdd.n2387 vdd.n682 99.5127
R3169 vdd.n2384 vdd.n682 99.5127
R3170 vdd.n2384 vdd.n677 99.5127
R3171 vdd.n2381 vdd.n677 99.5127
R3172 vdd.n2381 vdd.n672 99.5127
R3173 vdd.n2378 vdd.n672 99.5127
R3174 vdd.n2378 vdd.n666 99.5127
R3175 vdd.n2375 vdd.n666 99.5127
R3176 vdd.n2375 vdd.n659 99.5127
R3177 vdd.n2340 vdd.n659 99.5127
R3178 vdd.n2340 vdd.n654 99.5127
R3179 vdd.n2337 vdd.n654 99.5127
R3180 vdd.n2337 vdd.n649 99.5127
R3181 vdd.n2334 vdd.n649 99.5127
R3182 vdd.n2334 vdd.n643 99.5127
R3183 vdd.n2331 vdd.n643 99.5127
R3184 vdd.n2331 vdd.n635 99.5127
R3185 vdd.n2328 vdd.n635 99.5127
R3186 vdd.n2328 vdd.n628 99.5127
R3187 vdd.n628 vdd.n594 99.5127
R3188 vdd.n2674 vdd.n594 99.5127
R3189 vdd.n2473 vdd.n708 99.5127
R3190 vdd.n2261 vdd.n2260 99.5127
R3191 vdd.n2265 vdd.n2264 99.5127
R3192 vdd.n2269 vdd.n2268 99.5127
R3193 vdd.n2273 vdd.n2272 99.5127
R3194 vdd.n2277 vdd.n2276 99.5127
R3195 vdd.n2281 vdd.n2280 99.5127
R3196 vdd.n2285 vdd.n2284 99.5127
R3197 vdd.n2289 vdd.n2288 99.5127
R3198 vdd.n2293 vdd.n2292 99.5127
R3199 vdd.n2297 vdd.n2296 99.5127
R3200 vdd.n2301 vdd.n2300 99.5127
R3201 vdd.n2305 vdd.n2304 99.5127
R3202 vdd.n2309 vdd.n2308 99.5127
R3203 vdd.n2313 vdd.n2312 99.5127
R3204 vdd.n2317 vdd.n2316 99.5127
R3205 vdd.n2319 vdd.n2251 99.5127
R3206 vdd.n2477 vdd.n698 99.5127
R3207 vdd.n2485 vdd.n698 99.5127
R3208 vdd.n2485 vdd.n696 99.5127
R3209 vdd.n2489 vdd.n696 99.5127
R3210 vdd.n2489 vdd.n686 99.5127
R3211 vdd.n2497 vdd.n686 99.5127
R3212 vdd.n2497 vdd.n684 99.5127
R3213 vdd.n2501 vdd.n684 99.5127
R3214 vdd.n2501 vdd.n675 99.5127
R3215 vdd.n2509 vdd.n675 99.5127
R3216 vdd.n2509 vdd.n673 99.5127
R3217 vdd.n2513 vdd.n673 99.5127
R3218 vdd.n2513 vdd.n663 99.5127
R3219 vdd.n2521 vdd.n663 99.5127
R3220 vdd.n2521 vdd.n661 99.5127
R3221 vdd.n2525 vdd.n661 99.5127
R3222 vdd.n2525 vdd.n652 99.5127
R3223 vdd.n2533 vdd.n652 99.5127
R3224 vdd.n2533 vdd.n650 99.5127
R3225 vdd.n2539 vdd.n650 99.5127
R3226 vdd.n2539 vdd.n640 99.5127
R3227 vdd.n2547 vdd.n640 99.5127
R3228 vdd.n2547 vdd.n637 99.5127
R3229 vdd.n2596 vdd.n637 99.5127
R3230 vdd.n2596 vdd.n638 99.5127
R3231 vdd.n638 vdd.n629 99.5127
R3232 vdd.n2591 vdd.n629 99.5127
R3233 vdd.n2591 vdd.n597 99.5127
R3234 vdd.n2141 vdd.n2140 99.5127
R3235 vdd.n2137 vdd.n2136 99.5127
R3236 vdd.n2133 vdd.n2132 99.5127
R3237 vdd.n2129 vdd.n2128 99.5127
R3238 vdd.n2125 vdd.n2124 99.5127
R3239 vdd.n2121 vdd.n2120 99.5127
R3240 vdd.n2117 vdd.n2116 99.5127
R3241 vdd.n2113 vdd.n2112 99.5127
R3242 vdd.n2109 vdd.n2108 99.5127
R3243 vdd.n2105 vdd.n2104 99.5127
R3244 vdd.n2101 vdd.n2100 99.5127
R3245 vdd.n2097 vdd.n2096 99.5127
R3246 vdd.n2093 vdd.n2092 99.5127
R3247 vdd.n2089 vdd.n2088 99.5127
R3248 vdd.n2085 vdd.n2084 99.5127
R3249 vdd.n2081 vdd.n2080 99.5127
R3250 vdd.n2077 vdd.n726 99.5127
R3251 vdd.n1834 vdd.n841 99.5127
R3252 vdd.n1834 vdd.n835 99.5127
R3253 vdd.n1837 vdd.n835 99.5127
R3254 vdd.n1837 vdd.n829 99.5127
R3255 vdd.n1840 vdd.n829 99.5127
R3256 vdd.n1840 vdd.n822 99.5127
R3257 vdd.n1843 vdd.n822 99.5127
R3258 vdd.n1843 vdd.n815 99.5127
R3259 vdd.n1846 vdd.n815 99.5127
R3260 vdd.n1846 vdd.n810 99.5127
R3261 vdd.n1849 vdd.n810 99.5127
R3262 vdd.n1849 vdd.n804 99.5127
R3263 vdd.n1870 vdd.n804 99.5127
R3264 vdd.n1870 vdd.n797 99.5127
R3265 vdd.n1866 vdd.n797 99.5127
R3266 vdd.n1866 vdd.n791 99.5127
R3267 vdd.n1863 vdd.n791 99.5127
R3268 vdd.n1863 vdd.n786 99.5127
R3269 vdd.n1860 vdd.n786 99.5127
R3270 vdd.n1860 vdd.n781 99.5127
R3271 vdd.n1857 vdd.n781 99.5127
R3272 vdd.n1857 vdd.n775 99.5127
R3273 vdd.n1854 vdd.n775 99.5127
R3274 vdd.n1854 vdd.n768 99.5127
R3275 vdd.n768 vdd.n759 99.5127
R3276 vdd.n2072 vdd.n759 99.5127
R3277 vdd.n2073 vdd.n2072 99.5127
R3278 vdd.n2073 vdd.n751 99.5127
R3279 vdd.n1984 vdd.n1982 99.5127
R3280 vdd.n1980 vdd.n844 99.5127
R3281 vdd.n1976 vdd.n1974 99.5127
R3282 vdd.n1972 vdd.n846 99.5127
R3283 vdd.n1968 vdd.n1966 99.5127
R3284 vdd.n1964 vdd.n848 99.5127
R3285 vdd.n1960 vdd.n1958 99.5127
R3286 vdd.n1956 vdd.n850 99.5127
R3287 vdd.n1798 vdd.n852 99.5127
R3288 vdd.n1803 vdd.n1800 99.5127
R3289 vdd.n1807 vdd.n1805 99.5127
R3290 vdd.n1811 vdd.n1796 99.5127
R3291 vdd.n1815 vdd.n1813 99.5127
R3292 vdd.n1819 vdd.n1794 99.5127
R3293 vdd.n1823 vdd.n1821 99.5127
R3294 vdd.n1828 vdd.n1790 99.5127
R3295 vdd.n1831 vdd.n1830 99.5127
R3296 vdd.n1988 vdd.n832 99.5127
R3297 vdd.n1996 vdd.n832 99.5127
R3298 vdd.n1996 vdd.n830 99.5127
R3299 vdd.n2000 vdd.n830 99.5127
R3300 vdd.n2000 vdd.n819 99.5127
R3301 vdd.n2008 vdd.n819 99.5127
R3302 vdd.n2008 vdd.n816 99.5127
R3303 vdd.n2013 vdd.n816 99.5127
R3304 vdd.n2013 vdd.n807 99.5127
R3305 vdd.n2021 vdd.n807 99.5127
R3306 vdd.n2021 vdd.n805 99.5127
R3307 vdd.n2025 vdd.n805 99.5127
R3308 vdd.n2025 vdd.n795 99.5127
R3309 vdd.n2033 vdd.n795 99.5127
R3310 vdd.n2033 vdd.n793 99.5127
R3311 vdd.n2037 vdd.n793 99.5127
R3312 vdd.n2037 vdd.n784 99.5127
R3313 vdd.n2045 vdd.n784 99.5127
R3314 vdd.n2045 vdd.n782 99.5127
R3315 vdd.n2049 vdd.n782 99.5127
R3316 vdd.n2049 vdd.n772 99.5127
R3317 vdd.n2057 vdd.n772 99.5127
R3318 vdd.n2057 vdd.n769 99.5127
R3319 vdd.n2063 vdd.n769 99.5127
R3320 vdd.n2063 vdd.n770 99.5127
R3321 vdd.n770 vdd.n761 99.5127
R3322 vdd.n761 vdd.n752 99.5127
R3323 vdd.n2145 vdd.n752 99.5127
R3324 vdd.n9 vdd.n7 98.9633
R3325 vdd.n2 vdd.n0 98.9633
R3326 vdd.n9 vdd.n8 98.6055
R3327 vdd.n11 vdd.n10 98.6055
R3328 vdd.n13 vdd.n12 98.6055
R3329 vdd.n6 vdd.n5 98.6055
R3330 vdd.n4 vdd.n3 98.6055
R3331 vdd.n2 vdd.n1 98.6055
R3332 vdd.t144 vdd.n267 85.8723
R3333 vdd.t155 vdd.n220 85.8723
R3334 vdd.t140 vdd.n177 85.8723
R3335 vdd.t150 vdd.n130 85.8723
R3336 vdd.t181 vdd.n88 85.8723
R3337 vdd.t123 vdd.n41 85.8723
R3338 vdd.t179 vdd.n1082 85.8723
R3339 vdd.t165 vdd.n1129 85.8723
R3340 vdd.t171 vdd.n992 85.8723
R3341 vdd.t158 vdd.n1039 85.8723
R3342 vdd.t121 vdd.n903 85.8723
R3343 vdd.t180 vdd.n950 85.8723
R3344 vdd.n2537 vdd.n2536 78.546
R3345 vdd.n2011 vdd.n817 78.546
R3346 vdd.n254 vdd.n253 75.1835
R3347 vdd.n252 vdd.n251 75.1835
R3348 vdd.n250 vdd.n249 75.1835
R3349 vdd.n164 vdd.n163 75.1835
R3350 vdd.n162 vdd.n161 75.1835
R3351 vdd.n160 vdd.n159 75.1835
R3352 vdd.n75 vdd.n74 75.1835
R3353 vdd.n73 vdd.n72 75.1835
R3354 vdd.n71 vdd.n70 75.1835
R3355 vdd.n1112 vdd.n1111 75.1835
R3356 vdd.n1114 vdd.n1113 75.1835
R3357 vdd.n1116 vdd.n1115 75.1835
R3358 vdd.n1022 vdd.n1021 75.1835
R3359 vdd.n1024 vdd.n1023 75.1835
R3360 vdd.n1026 vdd.n1025 75.1835
R3361 vdd.n933 vdd.n932 75.1835
R3362 vdd.n935 vdd.n934 75.1835
R3363 vdd.n937 vdd.n936 75.1835
R3364 vdd.n2472 vdd.n2471 72.8958
R3365 vdd.n2471 vdd.n2235 72.8958
R3366 vdd.n2471 vdd.n2236 72.8958
R3367 vdd.n2471 vdd.n2237 72.8958
R3368 vdd.n2471 vdd.n2238 72.8958
R3369 vdd.n2471 vdd.n2239 72.8958
R3370 vdd.n2471 vdd.n2240 72.8958
R3371 vdd.n2471 vdd.n2241 72.8958
R3372 vdd.n2471 vdd.n2242 72.8958
R3373 vdd.n2471 vdd.n2243 72.8958
R3374 vdd.n2471 vdd.n2244 72.8958
R3375 vdd.n2471 vdd.n2245 72.8958
R3376 vdd.n2471 vdd.n2246 72.8958
R3377 vdd.n2471 vdd.n2247 72.8958
R3378 vdd.n2471 vdd.n2248 72.8958
R3379 vdd.n2471 vdd.n2249 72.8958
R3380 vdd.n2471 vdd.n2250 72.8958
R3381 vdd.n593 vdd.n484 72.8958
R3382 vdd.n2680 vdd.n484 72.8958
R3383 vdd.n587 vdd.n484 72.8958
R3384 vdd.n2687 vdd.n484 72.8958
R3385 vdd.n584 vdd.n484 72.8958
R3386 vdd.n2694 vdd.n484 72.8958
R3387 vdd.n581 vdd.n484 72.8958
R3388 vdd.n2701 vdd.n484 72.8958
R3389 vdd.n2704 vdd.n484 72.8958
R3390 vdd.n2560 vdd.n484 72.8958
R3391 vdd.n2565 vdd.n484 72.8958
R3392 vdd.n2559 vdd.n484 72.8958
R3393 vdd.n2572 vdd.n484 72.8958
R3394 vdd.n2556 vdd.n484 72.8958
R3395 vdd.n2579 vdd.n484 72.8958
R3396 vdd.n2553 vdd.n484 72.8958
R3397 vdd.n2586 vdd.n484 72.8958
R3398 vdd.n1724 vdd.n839 72.8958
R3399 vdd.n1730 vdd.n839 72.8958
R3400 vdd.n1732 vdd.n839 72.8958
R3401 vdd.n1738 vdd.n839 72.8958
R3402 vdd.n1740 vdd.n839 72.8958
R3403 vdd.n1746 vdd.n839 72.8958
R3404 vdd.n1748 vdd.n839 72.8958
R3405 vdd.n1754 vdd.n839 72.8958
R3406 vdd.n1925 vdd.n839 72.8958
R3407 vdd.n1923 vdd.n839 72.8958
R3408 vdd.n1917 vdd.n839 72.8958
R3409 vdd.n1915 vdd.n839 72.8958
R3410 vdd.n1909 vdd.n839 72.8958
R3411 vdd.n1907 vdd.n839 72.8958
R3412 vdd.n1901 vdd.n839 72.8958
R3413 vdd.n1899 vdd.n839 72.8958
R3414 vdd.n1893 vdd.n839 72.8958
R3415 vdd.n2218 vdd.n727 72.8958
R3416 vdd.n2218 vdd.n728 72.8958
R3417 vdd.n2218 vdd.n729 72.8958
R3418 vdd.n2218 vdd.n730 72.8958
R3419 vdd.n2218 vdd.n731 72.8958
R3420 vdd.n2218 vdd.n732 72.8958
R3421 vdd.n2218 vdd.n733 72.8958
R3422 vdd.n2218 vdd.n734 72.8958
R3423 vdd.n2218 vdd.n735 72.8958
R3424 vdd.n2218 vdd.n736 72.8958
R3425 vdd.n2218 vdd.n737 72.8958
R3426 vdd.n2218 vdd.n738 72.8958
R3427 vdd.n2218 vdd.n739 72.8958
R3428 vdd.n2218 vdd.n740 72.8958
R3429 vdd.n2218 vdd.n741 72.8958
R3430 vdd.n2218 vdd.n742 72.8958
R3431 vdd.n2218 vdd.n743 72.8958
R3432 vdd.n2471 vdd.n2470 72.8958
R3433 vdd.n2471 vdd.n2219 72.8958
R3434 vdd.n2471 vdd.n2220 72.8958
R3435 vdd.n2471 vdd.n2221 72.8958
R3436 vdd.n2471 vdd.n2222 72.8958
R3437 vdd.n2471 vdd.n2223 72.8958
R3438 vdd.n2471 vdd.n2224 72.8958
R3439 vdd.n2471 vdd.n2225 72.8958
R3440 vdd.n2471 vdd.n2226 72.8958
R3441 vdd.n2471 vdd.n2227 72.8958
R3442 vdd.n2471 vdd.n2228 72.8958
R3443 vdd.n2471 vdd.n2229 72.8958
R3444 vdd.n2471 vdd.n2230 72.8958
R3445 vdd.n2471 vdd.n2231 72.8958
R3446 vdd.n2471 vdd.n2232 72.8958
R3447 vdd.n2471 vdd.n2233 72.8958
R3448 vdd.n2471 vdd.n2234 72.8958
R3449 vdd.n2610 vdd.n484 72.8958
R3450 vdd.n625 vdd.n484 72.8958
R3451 vdd.n2618 vdd.n484 72.8958
R3452 vdd.n620 vdd.n484 72.8958
R3453 vdd.n2625 vdd.n484 72.8958
R3454 vdd.n617 vdd.n484 72.8958
R3455 vdd.n2632 vdd.n484 72.8958
R3456 vdd.n614 vdd.n484 72.8958
R3457 vdd.n2639 vdd.n484 72.8958
R3458 vdd.n2643 vdd.n484 72.8958
R3459 vdd.n611 vdd.n484 72.8958
R3460 vdd.n2650 vdd.n484 72.8958
R3461 vdd.n608 vdd.n484 72.8958
R3462 vdd.n2657 vdd.n484 72.8958
R3463 vdd.n605 vdd.n484 72.8958
R3464 vdd.n2664 vdd.n484 72.8958
R3465 vdd.n2667 vdd.n484 72.8958
R3466 vdd.n2218 vdd.n725 72.8958
R3467 vdd.n2218 vdd.n724 72.8958
R3468 vdd.n2218 vdd.n723 72.8958
R3469 vdd.n2218 vdd.n722 72.8958
R3470 vdd.n2218 vdd.n721 72.8958
R3471 vdd.n2218 vdd.n720 72.8958
R3472 vdd.n2218 vdd.n719 72.8958
R3473 vdd.n2218 vdd.n718 72.8958
R3474 vdd.n2218 vdd.n717 72.8958
R3475 vdd.n2218 vdd.n716 72.8958
R3476 vdd.n2218 vdd.n715 72.8958
R3477 vdd.n2218 vdd.n714 72.8958
R3478 vdd.n2218 vdd.n713 72.8958
R3479 vdd.n2218 vdd.n712 72.8958
R3480 vdd.n2218 vdd.n711 72.8958
R3481 vdd.n2218 vdd.n710 72.8958
R3482 vdd.n2218 vdd.n709 72.8958
R3483 vdd.n1983 vdd.n839 72.8958
R3484 vdd.n1981 vdd.n839 72.8958
R3485 vdd.n1975 vdd.n839 72.8958
R3486 vdd.n1973 vdd.n839 72.8958
R3487 vdd.n1967 vdd.n839 72.8958
R3488 vdd.n1965 vdd.n839 72.8958
R3489 vdd.n1959 vdd.n839 72.8958
R3490 vdd.n1957 vdd.n839 72.8958
R3491 vdd.n851 vdd.n839 72.8958
R3492 vdd.n1799 vdd.n839 72.8958
R3493 vdd.n1804 vdd.n839 72.8958
R3494 vdd.n1806 vdd.n839 72.8958
R3495 vdd.n1812 vdd.n839 72.8958
R3496 vdd.n1814 vdd.n839 72.8958
R3497 vdd.n1820 vdd.n839 72.8958
R3498 vdd.n1822 vdd.n839 72.8958
R3499 vdd.n1829 vdd.n839 72.8958
R3500 vdd.n1422 vdd.n1421 66.2847
R3501 vdd.n1421 vdd.n1197 66.2847
R3502 vdd.n1421 vdd.n1198 66.2847
R3503 vdd.n1421 vdd.n1199 66.2847
R3504 vdd.n1421 vdd.n1200 66.2847
R3505 vdd.n1421 vdd.n1201 66.2847
R3506 vdd.n1421 vdd.n1202 66.2847
R3507 vdd.n1421 vdd.n1203 66.2847
R3508 vdd.n1421 vdd.n1204 66.2847
R3509 vdd.n1421 vdd.n1205 66.2847
R3510 vdd.n1421 vdd.n1206 66.2847
R3511 vdd.n1421 vdd.n1207 66.2847
R3512 vdd.n1421 vdd.n1208 66.2847
R3513 vdd.n1421 vdd.n1209 66.2847
R3514 vdd.n1421 vdd.n1210 66.2847
R3515 vdd.n1421 vdd.n1211 66.2847
R3516 vdd.n1421 vdd.n1212 66.2847
R3517 vdd.n1421 vdd.n1213 66.2847
R3518 vdd.n1421 vdd.n1214 66.2847
R3519 vdd.n1421 vdd.n1215 66.2847
R3520 vdd.n1421 vdd.n1216 66.2847
R3521 vdd.n1421 vdd.n1217 66.2847
R3522 vdd.n1421 vdd.n1218 66.2847
R3523 vdd.n1421 vdd.n1219 66.2847
R3524 vdd.n1421 vdd.n1220 66.2847
R3525 vdd.n1421 vdd.n1221 66.2847
R3526 vdd.n1421 vdd.n1222 66.2847
R3527 vdd.n1421 vdd.n1223 66.2847
R3528 vdd.n1421 vdd.n1224 66.2847
R3529 vdd.n1421 vdd.n1225 66.2847
R3530 vdd.n1421 vdd.n1226 66.2847
R3531 vdd.n863 vdd.n860 66.2847
R3532 vdd.n1614 vdd.n863 66.2847
R3533 vdd.n1619 vdd.n863 66.2847
R3534 vdd.n1624 vdd.n863 66.2847
R3535 vdd.n1612 vdd.n863 66.2847
R3536 vdd.n1631 vdd.n863 66.2847
R3537 vdd.n1604 vdd.n863 66.2847
R3538 vdd.n1638 vdd.n863 66.2847
R3539 vdd.n1597 vdd.n863 66.2847
R3540 vdd.n1645 vdd.n863 66.2847
R3541 vdd.n1591 vdd.n863 66.2847
R3542 vdd.n1586 vdd.n863 66.2847
R3543 vdd.n1656 vdd.n863 66.2847
R3544 vdd.n1578 vdd.n863 66.2847
R3545 vdd.n1663 vdd.n863 66.2847
R3546 vdd.n1571 vdd.n863 66.2847
R3547 vdd.n1670 vdd.n863 66.2847
R3548 vdd.n1564 vdd.n863 66.2847
R3549 vdd.n1677 vdd.n863 66.2847
R3550 vdd.n1557 vdd.n863 66.2847
R3551 vdd.n1684 vdd.n863 66.2847
R3552 vdd.n1551 vdd.n863 66.2847
R3553 vdd.n1546 vdd.n863 66.2847
R3554 vdd.n1695 vdd.n863 66.2847
R3555 vdd.n1538 vdd.n863 66.2847
R3556 vdd.n1702 vdd.n863 66.2847
R3557 vdd.n1531 vdd.n863 66.2847
R3558 vdd.n1709 vdd.n863 66.2847
R3559 vdd.n1712 vdd.n863 66.2847
R3560 vdd.n1522 vdd.n863 66.2847
R3561 vdd.n1934 vdd.n863 66.2847
R3562 vdd.n1516 vdd.n863 66.2847
R3563 vdd.n2841 vdd.n2840 66.2847
R3564 vdd.n2840 vdd.n485 66.2847
R3565 vdd.n2840 vdd.n486 66.2847
R3566 vdd.n2840 vdd.n487 66.2847
R3567 vdd.n2840 vdd.n488 66.2847
R3568 vdd.n2840 vdd.n489 66.2847
R3569 vdd.n2840 vdd.n490 66.2847
R3570 vdd.n2840 vdd.n491 66.2847
R3571 vdd.n2840 vdd.n492 66.2847
R3572 vdd.n2840 vdd.n493 66.2847
R3573 vdd.n2840 vdd.n494 66.2847
R3574 vdd.n2840 vdd.n495 66.2847
R3575 vdd.n2840 vdd.n496 66.2847
R3576 vdd.n2840 vdd.n497 66.2847
R3577 vdd.n2840 vdd.n498 66.2847
R3578 vdd.n2840 vdd.n499 66.2847
R3579 vdd.n2840 vdd.n500 66.2847
R3580 vdd.n2840 vdd.n501 66.2847
R3581 vdd.n2840 vdd.n502 66.2847
R3582 vdd.n2840 vdd.n503 66.2847
R3583 vdd.n2840 vdd.n504 66.2847
R3584 vdd.n2840 vdd.n505 66.2847
R3585 vdd.n2840 vdd.n506 66.2847
R3586 vdd.n2840 vdd.n507 66.2847
R3587 vdd.n2840 vdd.n508 66.2847
R3588 vdd.n2840 vdd.n509 66.2847
R3589 vdd.n2840 vdd.n510 66.2847
R3590 vdd.n2840 vdd.n511 66.2847
R3591 vdd.n2840 vdd.n512 66.2847
R3592 vdd.n2840 vdd.n513 66.2847
R3593 vdd.n2840 vdd.n514 66.2847
R3594 vdd.n2905 vdd.n329 66.2847
R3595 vdd.n2914 vdd.n329 66.2847
R3596 vdd.n439 vdd.n329 66.2847
R3597 vdd.n2921 vdd.n329 66.2847
R3598 vdd.n432 vdd.n329 66.2847
R3599 vdd.n2928 vdd.n329 66.2847
R3600 vdd.n425 vdd.n329 66.2847
R3601 vdd.n2935 vdd.n329 66.2847
R3602 vdd.n418 vdd.n329 66.2847
R3603 vdd.n2942 vdd.n329 66.2847
R3604 vdd.n412 vdd.n329 66.2847
R3605 vdd.n407 vdd.n329 66.2847
R3606 vdd.n2953 vdd.n329 66.2847
R3607 vdd.n399 vdd.n329 66.2847
R3608 vdd.n2960 vdd.n329 66.2847
R3609 vdd.n392 vdd.n329 66.2847
R3610 vdd.n2967 vdd.n329 66.2847
R3611 vdd.n385 vdd.n329 66.2847
R3612 vdd.n2974 vdd.n329 66.2847
R3613 vdd.n378 vdd.n329 66.2847
R3614 vdd.n2981 vdd.n329 66.2847
R3615 vdd.n372 vdd.n329 66.2847
R3616 vdd.n367 vdd.n329 66.2847
R3617 vdd.n2992 vdd.n329 66.2847
R3618 vdd.n359 vdd.n329 66.2847
R3619 vdd.n2999 vdd.n329 66.2847
R3620 vdd.n352 vdd.n329 66.2847
R3621 vdd.n3006 vdd.n329 66.2847
R3622 vdd.n345 vdd.n329 66.2847
R3623 vdd.n3013 vdd.n329 66.2847
R3624 vdd.n3016 vdd.n329 66.2847
R3625 vdd.n333 vdd.n329 66.2847
R3626 vdd.n334 vdd.n333 52.4337
R3627 vdd.n3016 vdd.n3015 52.4337
R3628 vdd.n3013 vdd.n3012 52.4337
R3629 vdd.n3008 vdd.n345 52.4337
R3630 vdd.n3006 vdd.n3005 52.4337
R3631 vdd.n3001 vdd.n352 52.4337
R3632 vdd.n2999 vdd.n2998 52.4337
R3633 vdd.n2994 vdd.n359 52.4337
R3634 vdd.n2992 vdd.n2991 52.4337
R3635 vdd.n368 vdd.n367 52.4337
R3636 vdd.n2983 vdd.n372 52.4337
R3637 vdd.n2981 vdd.n2980 52.4337
R3638 vdd.n2976 vdd.n378 52.4337
R3639 vdd.n2974 vdd.n2973 52.4337
R3640 vdd.n2969 vdd.n385 52.4337
R3641 vdd.n2967 vdd.n2966 52.4337
R3642 vdd.n2962 vdd.n392 52.4337
R3643 vdd.n2960 vdd.n2959 52.4337
R3644 vdd.n2955 vdd.n399 52.4337
R3645 vdd.n2953 vdd.n2952 52.4337
R3646 vdd.n408 vdd.n407 52.4337
R3647 vdd.n2944 vdd.n412 52.4337
R3648 vdd.n2942 vdd.n2941 52.4337
R3649 vdd.n2937 vdd.n418 52.4337
R3650 vdd.n2935 vdd.n2934 52.4337
R3651 vdd.n2930 vdd.n425 52.4337
R3652 vdd.n2928 vdd.n2927 52.4337
R3653 vdd.n2923 vdd.n432 52.4337
R3654 vdd.n2921 vdd.n2920 52.4337
R3655 vdd.n2916 vdd.n439 52.4337
R3656 vdd.n2914 vdd.n2913 52.4337
R3657 vdd.n2906 vdd.n2905 52.4337
R3658 vdd.n2842 vdd.n2841 52.4337
R3659 vdd.n517 vdd.n485 52.4337
R3660 vdd.n523 vdd.n486 52.4337
R3661 vdd.n2831 vdd.n487 52.4337
R3662 vdd.n2827 vdd.n488 52.4337
R3663 vdd.n2823 vdd.n489 52.4337
R3664 vdd.n2819 vdd.n490 52.4337
R3665 vdd.n2815 vdd.n491 52.4337
R3666 vdd.n2811 vdd.n492 52.4337
R3667 vdd.n2807 vdd.n493 52.4337
R3668 vdd.n2799 vdd.n494 52.4337
R3669 vdd.n2795 vdd.n495 52.4337
R3670 vdd.n2791 vdd.n496 52.4337
R3671 vdd.n2787 vdd.n497 52.4337
R3672 vdd.n2783 vdd.n498 52.4337
R3673 vdd.n2779 vdd.n499 52.4337
R3674 vdd.n2775 vdd.n500 52.4337
R3675 vdd.n2771 vdd.n501 52.4337
R3676 vdd.n2767 vdd.n502 52.4337
R3677 vdd.n2763 vdd.n503 52.4337
R3678 vdd.n2759 vdd.n504 52.4337
R3679 vdd.n2753 vdd.n505 52.4337
R3680 vdd.n2749 vdd.n506 52.4337
R3681 vdd.n2745 vdd.n507 52.4337
R3682 vdd.n2741 vdd.n508 52.4337
R3683 vdd.n2737 vdd.n509 52.4337
R3684 vdd.n2733 vdd.n510 52.4337
R3685 vdd.n2729 vdd.n511 52.4337
R3686 vdd.n2725 vdd.n512 52.4337
R3687 vdd.n2721 vdd.n513 52.4337
R3688 vdd.n2717 vdd.n514 52.4337
R3689 vdd.n1936 vdd.n1516 52.4337
R3690 vdd.n1934 vdd.n1933 52.4337
R3691 vdd.n1523 vdd.n1522 52.4337
R3692 vdd.n1712 vdd.n1711 52.4337
R3693 vdd.n1709 vdd.n1708 52.4337
R3694 vdd.n1704 vdd.n1531 52.4337
R3695 vdd.n1702 vdd.n1701 52.4337
R3696 vdd.n1697 vdd.n1538 52.4337
R3697 vdd.n1695 vdd.n1694 52.4337
R3698 vdd.n1547 vdd.n1546 52.4337
R3699 vdd.n1686 vdd.n1551 52.4337
R3700 vdd.n1684 vdd.n1683 52.4337
R3701 vdd.n1679 vdd.n1557 52.4337
R3702 vdd.n1677 vdd.n1676 52.4337
R3703 vdd.n1672 vdd.n1564 52.4337
R3704 vdd.n1670 vdd.n1669 52.4337
R3705 vdd.n1665 vdd.n1571 52.4337
R3706 vdd.n1663 vdd.n1662 52.4337
R3707 vdd.n1658 vdd.n1578 52.4337
R3708 vdd.n1656 vdd.n1655 52.4337
R3709 vdd.n1587 vdd.n1586 52.4337
R3710 vdd.n1647 vdd.n1591 52.4337
R3711 vdd.n1645 vdd.n1644 52.4337
R3712 vdd.n1640 vdd.n1597 52.4337
R3713 vdd.n1638 vdd.n1637 52.4337
R3714 vdd.n1633 vdd.n1604 52.4337
R3715 vdd.n1631 vdd.n1630 52.4337
R3716 vdd.n1626 vdd.n1612 52.4337
R3717 vdd.n1624 vdd.n1623 52.4337
R3718 vdd.n1619 vdd.n1618 52.4337
R3719 vdd.n1614 vdd.n1613 52.4337
R3720 vdd.n1945 vdd.n860 52.4337
R3721 vdd.n1423 vdd.n1422 52.4337
R3722 vdd.n1229 vdd.n1197 52.4337
R3723 vdd.n1233 vdd.n1198 52.4337
R3724 vdd.n1235 vdd.n1199 52.4337
R3725 vdd.n1239 vdd.n1200 52.4337
R3726 vdd.n1241 vdd.n1201 52.4337
R3727 vdd.n1245 vdd.n1202 52.4337
R3728 vdd.n1247 vdd.n1203 52.4337
R3729 vdd.n1251 vdd.n1204 52.4337
R3730 vdd.n1253 vdd.n1205 52.4337
R3731 vdd.n1259 vdd.n1206 52.4337
R3732 vdd.n1261 vdd.n1207 52.4337
R3733 vdd.n1265 vdd.n1208 52.4337
R3734 vdd.n1267 vdd.n1209 52.4337
R3735 vdd.n1271 vdd.n1210 52.4337
R3736 vdd.n1273 vdd.n1211 52.4337
R3737 vdd.n1277 vdd.n1212 52.4337
R3738 vdd.n1279 vdd.n1213 52.4337
R3739 vdd.n1283 vdd.n1214 52.4337
R3740 vdd.n1285 vdd.n1215 52.4337
R3741 vdd.n1357 vdd.n1216 52.4337
R3742 vdd.n1290 vdd.n1217 52.4337
R3743 vdd.n1294 vdd.n1218 52.4337
R3744 vdd.n1296 vdd.n1219 52.4337
R3745 vdd.n1300 vdd.n1220 52.4337
R3746 vdd.n1302 vdd.n1221 52.4337
R3747 vdd.n1306 vdd.n1222 52.4337
R3748 vdd.n1308 vdd.n1223 52.4337
R3749 vdd.n1312 vdd.n1224 52.4337
R3750 vdd.n1314 vdd.n1225 52.4337
R3751 vdd.n1318 vdd.n1226 52.4337
R3752 vdd.n1422 vdd.n1196 52.4337
R3753 vdd.n1232 vdd.n1197 52.4337
R3754 vdd.n1234 vdd.n1198 52.4337
R3755 vdd.n1238 vdd.n1199 52.4337
R3756 vdd.n1240 vdd.n1200 52.4337
R3757 vdd.n1244 vdd.n1201 52.4337
R3758 vdd.n1246 vdd.n1202 52.4337
R3759 vdd.n1250 vdd.n1203 52.4337
R3760 vdd.n1252 vdd.n1204 52.4337
R3761 vdd.n1258 vdd.n1205 52.4337
R3762 vdd.n1260 vdd.n1206 52.4337
R3763 vdd.n1264 vdd.n1207 52.4337
R3764 vdd.n1266 vdd.n1208 52.4337
R3765 vdd.n1270 vdd.n1209 52.4337
R3766 vdd.n1272 vdd.n1210 52.4337
R3767 vdd.n1276 vdd.n1211 52.4337
R3768 vdd.n1278 vdd.n1212 52.4337
R3769 vdd.n1282 vdd.n1213 52.4337
R3770 vdd.n1284 vdd.n1214 52.4337
R3771 vdd.n1288 vdd.n1215 52.4337
R3772 vdd.n1289 vdd.n1216 52.4337
R3773 vdd.n1293 vdd.n1217 52.4337
R3774 vdd.n1295 vdd.n1218 52.4337
R3775 vdd.n1299 vdd.n1219 52.4337
R3776 vdd.n1301 vdd.n1220 52.4337
R3777 vdd.n1305 vdd.n1221 52.4337
R3778 vdd.n1307 vdd.n1222 52.4337
R3779 vdd.n1311 vdd.n1223 52.4337
R3780 vdd.n1313 vdd.n1224 52.4337
R3781 vdd.n1317 vdd.n1225 52.4337
R3782 vdd.n1319 vdd.n1226 52.4337
R3783 vdd.n860 vdd.n859 52.4337
R3784 vdd.n1615 vdd.n1614 52.4337
R3785 vdd.n1620 vdd.n1619 52.4337
R3786 vdd.n1625 vdd.n1624 52.4337
R3787 vdd.n1612 vdd.n1605 52.4337
R3788 vdd.n1632 vdd.n1631 52.4337
R3789 vdd.n1604 vdd.n1598 52.4337
R3790 vdd.n1639 vdd.n1638 52.4337
R3791 vdd.n1597 vdd.n1592 52.4337
R3792 vdd.n1646 vdd.n1645 52.4337
R3793 vdd.n1591 vdd.n1590 52.4337
R3794 vdd.n1586 vdd.n1579 52.4337
R3795 vdd.n1657 vdd.n1656 52.4337
R3796 vdd.n1578 vdd.n1572 52.4337
R3797 vdd.n1664 vdd.n1663 52.4337
R3798 vdd.n1571 vdd.n1565 52.4337
R3799 vdd.n1671 vdd.n1670 52.4337
R3800 vdd.n1564 vdd.n1558 52.4337
R3801 vdd.n1678 vdd.n1677 52.4337
R3802 vdd.n1557 vdd.n1552 52.4337
R3803 vdd.n1685 vdd.n1684 52.4337
R3804 vdd.n1551 vdd.n1550 52.4337
R3805 vdd.n1546 vdd.n1539 52.4337
R3806 vdd.n1696 vdd.n1695 52.4337
R3807 vdd.n1538 vdd.n1532 52.4337
R3808 vdd.n1703 vdd.n1702 52.4337
R3809 vdd.n1531 vdd.n1525 52.4337
R3810 vdd.n1710 vdd.n1709 52.4337
R3811 vdd.n1713 vdd.n1712 52.4337
R3812 vdd.n1522 vdd.n1517 52.4337
R3813 vdd.n1935 vdd.n1934 52.4337
R3814 vdd.n1516 vdd.n865 52.4337
R3815 vdd.n2841 vdd.n483 52.4337
R3816 vdd.n522 vdd.n485 52.4337
R3817 vdd.n2832 vdd.n486 52.4337
R3818 vdd.n2828 vdd.n487 52.4337
R3819 vdd.n2824 vdd.n488 52.4337
R3820 vdd.n2820 vdd.n489 52.4337
R3821 vdd.n2816 vdd.n490 52.4337
R3822 vdd.n2812 vdd.n491 52.4337
R3823 vdd.n2808 vdd.n492 52.4337
R3824 vdd.n2798 vdd.n493 52.4337
R3825 vdd.n2796 vdd.n494 52.4337
R3826 vdd.n2792 vdd.n495 52.4337
R3827 vdd.n2788 vdd.n496 52.4337
R3828 vdd.n2784 vdd.n497 52.4337
R3829 vdd.n2780 vdd.n498 52.4337
R3830 vdd.n2776 vdd.n499 52.4337
R3831 vdd.n2772 vdd.n500 52.4337
R3832 vdd.n2768 vdd.n501 52.4337
R3833 vdd.n2764 vdd.n502 52.4337
R3834 vdd.n2760 vdd.n503 52.4337
R3835 vdd.n2752 vdd.n504 52.4337
R3836 vdd.n2750 vdd.n505 52.4337
R3837 vdd.n2746 vdd.n506 52.4337
R3838 vdd.n2742 vdd.n507 52.4337
R3839 vdd.n2738 vdd.n508 52.4337
R3840 vdd.n2734 vdd.n509 52.4337
R3841 vdd.n2730 vdd.n510 52.4337
R3842 vdd.n2726 vdd.n511 52.4337
R3843 vdd.n2722 vdd.n512 52.4337
R3844 vdd.n2718 vdd.n513 52.4337
R3845 vdd.n2714 vdd.n514 52.4337
R3846 vdd.n2905 vdd.n440 52.4337
R3847 vdd.n2915 vdd.n2914 52.4337
R3848 vdd.n439 vdd.n433 52.4337
R3849 vdd.n2922 vdd.n2921 52.4337
R3850 vdd.n432 vdd.n426 52.4337
R3851 vdd.n2929 vdd.n2928 52.4337
R3852 vdd.n425 vdd.n419 52.4337
R3853 vdd.n2936 vdd.n2935 52.4337
R3854 vdd.n418 vdd.n413 52.4337
R3855 vdd.n2943 vdd.n2942 52.4337
R3856 vdd.n412 vdd.n411 52.4337
R3857 vdd.n407 vdd.n400 52.4337
R3858 vdd.n2954 vdd.n2953 52.4337
R3859 vdd.n399 vdd.n393 52.4337
R3860 vdd.n2961 vdd.n2960 52.4337
R3861 vdd.n392 vdd.n386 52.4337
R3862 vdd.n2968 vdd.n2967 52.4337
R3863 vdd.n385 vdd.n379 52.4337
R3864 vdd.n2975 vdd.n2974 52.4337
R3865 vdd.n378 vdd.n373 52.4337
R3866 vdd.n2982 vdd.n2981 52.4337
R3867 vdd.n372 vdd.n371 52.4337
R3868 vdd.n367 vdd.n360 52.4337
R3869 vdd.n2993 vdd.n2992 52.4337
R3870 vdd.n359 vdd.n353 52.4337
R3871 vdd.n3000 vdd.n2999 52.4337
R3872 vdd.n352 vdd.n346 52.4337
R3873 vdd.n3007 vdd.n3006 52.4337
R3874 vdd.n345 vdd.n338 52.4337
R3875 vdd.n3014 vdd.n3013 52.4337
R3876 vdd.n3017 vdd.n3016 52.4337
R3877 vdd.n333 vdd.n330 52.4337
R3878 vdd.t22 vdd.t118 51.4683
R3879 vdd.n250 vdd.n248 42.0461
R3880 vdd.n160 vdd.n158 42.0461
R3881 vdd.n71 vdd.n69 42.0461
R3882 vdd.n1112 vdd.n1110 42.0461
R3883 vdd.n1022 vdd.n1020 42.0461
R3884 vdd.n933 vdd.n931 42.0461
R3885 vdd.n296 vdd.n295 41.6884
R3886 vdd.n206 vdd.n205 41.6884
R3887 vdd.n117 vdd.n116 41.6884
R3888 vdd.n1158 vdd.n1157 41.6884
R3889 vdd.n1068 vdd.n1067 41.6884
R3890 vdd.n979 vdd.n978 41.6884
R3891 vdd.n1322 vdd.n1321 41.1157
R3892 vdd.n1360 vdd.n1359 41.1157
R3893 vdd.n1256 vdd.n1255 41.1157
R3894 vdd.n2910 vdd.n2909 41.1157
R3895 vdd.n2949 vdd.n406 41.1157
R3896 vdd.n2988 vdd.n366 41.1157
R3897 vdd.n2667 vdd.n2666 39.2114
R3898 vdd.n2664 vdd.n2663 39.2114
R3899 vdd.n2659 vdd.n605 39.2114
R3900 vdd.n2657 vdd.n2656 39.2114
R3901 vdd.n2652 vdd.n608 39.2114
R3902 vdd.n2650 vdd.n2649 39.2114
R3903 vdd.n2645 vdd.n611 39.2114
R3904 vdd.n2643 vdd.n2642 39.2114
R3905 vdd.n2639 vdd.n2638 39.2114
R3906 vdd.n2634 vdd.n614 39.2114
R3907 vdd.n2632 vdd.n2631 39.2114
R3908 vdd.n2627 vdd.n617 39.2114
R3909 vdd.n2625 vdd.n2624 39.2114
R3910 vdd.n2620 vdd.n620 39.2114
R3911 vdd.n2618 vdd.n2617 39.2114
R3912 vdd.n2612 vdd.n625 39.2114
R3913 vdd.n2610 vdd.n2609 39.2114
R3914 vdd.n2470 vdd.n703 39.2114
R3915 vdd.n2465 vdd.n2219 39.2114
R3916 vdd.n2462 vdd.n2220 39.2114
R3917 vdd.n2458 vdd.n2221 39.2114
R3918 vdd.n2454 vdd.n2222 39.2114
R3919 vdd.n2450 vdd.n2223 39.2114
R3920 vdd.n2446 vdd.n2224 39.2114
R3921 vdd.n2442 vdd.n2225 39.2114
R3922 vdd.n2438 vdd.n2226 39.2114
R3923 vdd.n2434 vdd.n2227 39.2114
R3924 vdd.n2430 vdd.n2228 39.2114
R3925 vdd.n2426 vdd.n2229 39.2114
R3926 vdd.n2422 vdd.n2230 39.2114
R3927 vdd.n2418 vdd.n2231 39.2114
R3928 vdd.n2414 vdd.n2232 39.2114
R3929 vdd.n2410 vdd.n2233 39.2114
R3930 vdd.n2405 vdd.n2234 39.2114
R3931 vdd.n2213 vdd.n743 39.2114
R3932 vdd.n2209 vdd.n742 39.2114
R3933 vdd.n2205 vdd.n741 39.2114
R3934 vdd.n2201 vdd.n740 39.2114
R3935 vdd.n2197 vdd.n739 39.2114
R3936 vdd.n2193 vdd.n738 39.2114
R3937 vdd.n2189 vdd.n737 39.2114
R3938 vdd.n2185 vdd.n736 39.2114
R3939 vdd.n2181 vdd.n735 39.2114
R3940 vdd.n2177 vdd.n734 39.2114
R3941 vdd.n2173 vdd.n733 39.2114
R3942 vdd.n2169 vdd.n732 39.2114
R3943 vdd.n2165 vdd.n731 39.2114
R3944 vdd.n2161 vdd.n730 39.2114
R3945 vdd.n2157 vdd.n729 39.2114
R3946 vdd.n2152 vdd.n728 39.2114
R3947 vdd.n2148 vdd.n727 39.2114
R3948 vdd.n1724 vdd.n838 39.2114
R3949 vdd.n1730 vdd.n1729 39.2114
R3950 vdd.n1733 vdd.n1732 39.2114
R3951 vdd.n1738 vdd.n1737 39.2114
R3952 vdd.n1741 vdd.n1740 39.2114
R3953 vdd.n1746 vdd.n1745 39.2114
R3954 vdd.n1749 vdd.n1748 39.2114
R3955 vdd.n1754 vdd.n1753 39.2114
R3956 vdd.n1925 vdd.n1756 39.2114
R3957 vdd.n1924 vdd.n1923 39.2114
R3958 vdd.n1917 vdd.n1758 39.2114
R3959 vdd.n1916 vdd.n1915 39.2114
R3960 vdd.n1909 vdd.n1760 39.2114
R3961 vdd.n1908 vdd.n1907 39.2114
R3962 vdd.n1901 vdd.n1762 39.2114
R3963 vdd.n1900 vdd.n1899 39.2114
R3964 vdd.n1893 vdd.n1764 39.2114
R3965 vdd.n2586 vdd.n2585 39.2114
R3966 vdd.n2581 vdd.n2553 39.2114
R3967 vdd.n2579 vdd.n2578 39.2114
R3968 vdd.n2574 vdd.n2556 39.2114
R3969 vdd.n2572 vdd.n2571 39.2114
R3970 vdd.n2567 vdd.n2559 39.2114
R3971 vdd.n2565 vdd.n2564 39.2114
R3972 vdd.n2560 vdd.n577 39.2114
R3973 vdd.n2704 vdd.n2703 39.2114
R3974 vdd.n2701 vdd.n2700 39.2114
R3975 vdd.n2696 vdd.n581 39.2114
R3976 vdd.n2694 vdd.n2693 39.2114
R3977 vdd.n2689 vdd.n584 39.2114
R3978 vdd.n2687 vdd.n2686 39.2114
R3979 vdd.n2682 vdd.n587 39.2114
R3980 vdd.n2680 vdd.n2679 39.2114
R3981 vdd.n2675 vdd.n593 39.2114
R3982 vdd.n2472 vdd.n706 39.2114
R3983 vdd.n2235 vdd.n708 39.2114
R3984 vdd.n2261 vdd.n2236 39.2114
R3985 vdd.n2265 vdd.n2237 39.2114
R3986 vdd.n2269 vdd.n2238 39.2114
R3987 vdd.n2273 vdd.n2239 39.2114
R3988 vdd.n2277 vdd.n2240 39.2114
R3989 vdd.n2281 vdd.n2241 39.2114
R3990 vdd.n2285 vdd.n2242 39.2114
R3991 vdd.n2289 vdd.n2243 39.2114
R3992 vdd.n2293 vdd.n2244 39.2114
R3993 vdd.n2297 vdd.n2245 39.2114
R3994 vdd.n2301 vdd.n2246 39.2114
R3995 vdd.n2305 vdd.n2247 39.2114
R3996 vdd.n2309 vdd.n2248 39.2114
R3997 vdd.n2313 vdd.n2249 39.2114
R3998 vdd.n2317 vdd.n2250 39.2114
R3999 vdd.n2473 vdd.n2472 39.2114
R4000 vdd.n2260 vdd.n2235 39.2114
R4001 vdd.n2264 vdd.n2236 39.2114
R4002 vdd.n2268 vdd.n2237 39.2114
R4003 vdd.n2272 vdd.n2238 39.2114
R4004 vdd.n2276 vdd.n2239 39.2114
R4005 vdd.n2280 vdd.n2240 39.2114
R4006 vdd.n2284 vdd.n2241 39.2114
R4007 vdd.n2288 vdd.n2242 39.2114
R4008 vdd.n2292 vdd.n2243 39.2114
R4009 vdd.n2296 vdd.n2244 39.2114
R4010 vdd.n2300 vdd.n2245 39.2114
R4011 vdd.n2304 vdd.n2246 39.2114
R4012 vdd.n2308 vdd.n2247 39.2114
R4013 vdd.n2312 vdd.n2248 39.2114
R4014 vdd.n2316 vdd.n2249 39.2114
R4015 vdd.n2319 vdd.n2250 39.2114
R4016 vdd.n593 vdd.n588 39.2114
R4017 vdd.n2681 vdd.n2680 39.2114
R4018 vdd.n587 vdd.n585 39.2114
R4019 vdd.n2688 vdd.n2687 39.2114
R4020 vdd.n584 vdd.n582 39.2114
R4021 vdd.n2695 vdd.n2694 39.2114
R4022 vdd.n581 vdd.n579 39.2114
R4023 vdd.n2702 vdd.n2701 39.2114
R4024 vdd.n2705 vdd.n2704 39.2114
R4025 vdd.n2561 vdd.n2560 39.2114
R4026 vdd.n2566 vdd.n2565 39.2114
R4027 vdd.n2559 vdd.n2557 39.2114
R4028 vdd.n2573 vdd.n2572 39.2114
R4029 vdd.n2556 vdd.n2554 39.2114
R4030 vdd.n2580 vdd.n2579 39.2114
R4031 vdd.n2553 vdd.n2551 39.2114
R4032 vdd.n2587 vdd.n2586 39.2114
R4033 vdd.n1725 vdd.n1724 39.2114
R4034 vdd.n1731 vdd.n1730 39.2114
R4035 vdd.n1732 vdd.n1721 39.2114
R4036 vdd.n1739 vdd.n1738 39.2114
R4037 vdd.n1740 vdd.n1719 39.2114
R4038 vdd.n1747 vdd.n1746 39.2114
R4039 vdd.n1748 vdd.n1717 39.2114
R4040 vdd.n1755 vdd.n1754 39.2114
R4041 vdd.n1926 vdd.n1925 39.2114
R4042 vdd.n1923 vdd.n1922 39.2114
R4043 vdd.n1918 vdd.n1917 39.2114
R4044 vdd.n1915 vdd.n1914 39.2114
R4045 vdd.n1910 vdd.n1909 39.2114
R4046 vdd.n1907 vdd.n1906 39.2114
R4047 vdd.n1902 vdd.n1901 39.2114
R4048 vdd.n1899 vdd.n1898 39.2114
R4049 vdd.n1894 vdd.n1893 39.2114
R4050 vdd.n2151 vdd.n727 39.2114
R4051 vdd.n2156 vdd.n728 39.2114
R4052 vdd.n2160 vdd.n729 39.2114
R4053 vdd.n2164 vdd.n730 39.2114
R4054 vdd.n2168 vdd.n731 39.2114
R4055 vdd.n2172 vdd.n732 39.2114
R4056 vdd.n2176 vdd.n733 39.2114
R4057 vdd.n2180 vdd.n734 39.2114
R4058 vdd.n2184 vdd.n735 39.2114
R4059 vdd.n2188 vdd.n736 39.2114
R4060 vdd.n2192 vdd.n737 39.2114
R4061 vdd.n2196 vdd.n738 39.2114
R4062 vdd.n2200 vdd.n739 39.2114
R4063 vdd.n2204 vdd.n740 39.2114
R4064 vdd.n2208 vdd.n741 39.2114
R4065 vdd.n2212 vdd.n742 39.2114
R4066 vdd.n745 vdd.n743 39.2114
R4067 vdd.n2470 vdd.n2469 39.2114
R4068 vdd.n2463 vdd.n2219 39.2114
R4069 vdd.n2459 vdd.n2220 39.2114
R4070 vdd.n2455 vdd.n2221 39.2114
R4071 vdd.n2451 vdd.n2222 39.2114
R4072 vdd.n2447 vdd.n2223 39.2114
R4073 vdd.n2443 vdd.n2224 39.2114
R4074 vdd.n2439 vdd.n2225 39.2114
R4075 vdd.n2435 vdd.n2226 39.2114
R4076 vdd.n2431 vdd.n2227 39.2114
R4077 vdd.n2427 vdd.n2228 39.2114
R4078 vdd.n2423 vdd.n2229 39.2114
R4079 vdd.n2419 vdd.n2230 39.2114
R4080 vdd.n2415 vdd.n2231 39.2114
R4081 vdd.n2411 vdd.n2232 39.2114
R4082 vdd.n2406 vdd.n2233 39.2114
R4083 vdd.n2402 vdd.n2234 39.2114
R4084 vdd.n2611 vdd.n2610 39.2114
R4085 vdd.n625 vdd.n621 39.2114
R4086 vdd.n2619 vdd.n2618 39.2114
R4087 vdd.n620 vdd.n618 39.2114
R4088 vdd.n2626 vdd.n2625 39.2114
R4089 vdd.n617 vdd.n615 39.2114
R4090 vdd.n2633 vdd.n2632 39.2114
R4091 vdd.n614 vdd.n612 39.2114
R4092 vdd.n2640 vdd.n2639 39.2114
R4093 vdd.n2644 vdd.n2643 39.2114
R4094 vdd.n611 vdd.n609 39.2114
R4095 vdd.n2651 vdd.n2650 39.2114
R4096 vdd.n608 vdd.n606 39.2114
R4097 vdd.n2658 vdd.n2657 39.2114
R4098 vdd.n605 vdd.n603 39.2114
R4099 vdd.n2665 vdd.n2664 39.2114
R4100 vdd.n2668 vdd.n2667 39.2114
R4101 vdd.n753 vdd.n709 39.2114
R4102 vdd.n2140 vdd.n710 39.2114
R4103 vdd.n2136 vdd.n711 39.2114
R4104 vdd.n2132 vdd.n712 39.2114
R4105 vdd.n2128 vdd.n713 39.2114
R4106 vdd.n2124 vdd.n714 39.2114
R4107 vdd.n2120 vdd.n715 39.2114
R4108 vdd.n2116 vdd.n716 39.2114
R4109 vdd.n2112 vdd.n717 39.2114
R4110 vdd.n2108 vdd.n718 39.2114
R4111 vdd.n2104 vdd.n719 39.2114
R4112 vdd.n2100 vdd.n720 39.2114
R4113 vdd.n2096 vdd.n721 39.2114
R4114 vdd.n2092 vdd.n722 39.2114
R4115 vdd.n2088 vdd.n723 39.2114
R4116 vdd.n2084 vdd.n724 39.2114
R4117 vdd.n2080 vdd.n725 39.2114
R4118 vdd.n1983 vdd.n842 39.2114
R4119 vdd.n1982 vdd.n1981 39.2114
R4120 vdd.n1975 vdd.n844 39.2114
R4121 vdd.n1974 vdd.n1973 39.2114
R4122 vdd.n1967 vdd.n846 39.2114
R4123 vdd.n1966 vdd.n1965 39.2114
R4124 vdd.n1959 vdd.n848 39.2114
R4125 vdd.n1958 vdd.n1957 39.2114
R4126 vdd.n851 vdd.n850 39.2114
R4127 vdd.n1799 vdd.n1798 39.2114
R4128 vdd.n1804 vdd.n1803 39.2114
R4129 vdd.n1807 vdd.n1806 39.2114
R4130 vdd.n1812 vdd.n1811 39.2114
R4131 vdd.n1815 vdd.n1814 39.2114
R4132 vdd.n1820 vdd.n1819 39.2114
R4133 vdd.n1823 vdd.n1822 39.2114
R4134 vdd.n1829 vdd.n1828 39.2114
R4135 vdd.n2077 vdd.n725 39.2114
R4136 vdd.n2081 vdd.n724 39.2114
R4137 vdd.n2085 vdd.n723 39.2114
R4138 vdd.n2089 vdd.n722 39.2114
R4139 vdd.n2093 vdd.n721 39.2114
R4140 vdd.n2097 vdd.n720 39.2114
R4141 vdd.n2101 vdd.n719 39.2114
R4142 vdd.n2105 vdd.n718 39.2114
R4143 vdd.n2109 vdd.n717 39.2114
R4144 vdd.n2113 vdd.n716 39.2114
R4145 vdd.n2117 vdd.n715 39.2114
R4146 vdd.n2121 vdd.n714 39.2114
R4147 vdd.n2125 vdd.n713 39.2114
R4148 vdd.n2129 vdd.n712 39.2114
R4149 vdd.n2133 vdd.n711 39.2114
R4150 vdd.n2137 vdd.n710 39.2114
R4151 vdd.n2141 vdd.n709 39.2114
R4152 vdd.n1984 vdd.n1983 39.2114
R4153 vdd.n1981 vdd.n1980 39.2114
R4154 vdd.n1976 vdd.n1975 39.2114
R4155 vdd.n1973 vdd.n1972 39.2114
R4156 vdd.n1968 vdd.n1967 39.2114
R4157 vdd.n1965 vdd.n1964 39.2114
R4158 vdd.n1960 vdd.n1959 39.2114
R4159 vdd.n1957 vdd.n1956 39.2114
R4160 vdd.n852 vdd.n851 39.2114
R4161 vdd.n1800 vdd.n1799 39.2114
R4162 vdd.n1805 vdd.n1804 39.2114
R4163 vdd.n1806 vdd.n1796 39.2114
R4164 vdd.n1813 vdd.n1812 39.2114
R4165 vdd.n1814 vdd.n1794 39.2114
R4166 vdd.n1821 vdd.n1820 39.2114
R4167 vdd.n1822 vdd.n1790 39.2114
R4168 vdd.n1830 vdd.n1829 39.2114
R4169 vdd.n1949 vdd.n1948 37.2369
R4170 vdd.n1652 vdd.n1585 37.2369
R4171 vdd.n1691 vdd.n1545 37.2369
R4172 vdd.n2758 vdd.n558 37.2369
R4173 vdd.n2806 vdd.n2805 37.2369
R4174 vdd.n2713 vdd.n2712 37.2369
R4175 vdd.n1991 vdd.n837 31.6883
R4176 vdd.n2216 vdd.n746 31.6883
R4177 vdd.n2149 vdd.n749 31.6883
R4178 vdd.n1895 vdd.n1892 31.6883
R4179 vdd.n2403 vdd.n2401 31.6883
R4180 vdd.n2608 vdd.n2607 31.6883
R4181 vdd.n2480 vdd.n702 31.6883
R4182 vdd.n2671 vdd.n2670 31.6883
R4183 vdd.n2590 vdd.n2589 31.6883
R4184 vdd.n2676 vdd.n592 31.6883
R4185 vdd.n2322 vdd.n2321 31.6883
R4186 vdd.n2476 vdd.n2475 31.6883
R4187 vdd.n1987 vdd.n1986 31.6883
R4188 vdd.n2144 vdd.n2143 31.6883
R4189 vdd.n2076 vdd.n2075 31.6883
R4190 vdd.n1833 vdd.n1832 31.6883
R4191 vdd.n1826 vdd.n1792 30.449
R4192 vdd.n757 vdd.n756 30.449
R4193 vdd.n1767 vdd.n1766 30.449
R4194 vdd.n2154 vdd.n748 30.449
R4195 vdd.n2258 vdd.n2257 30.449
R4196 vdd.n2614 vdd.n623 30.449
R4197 vdd.n2408 vdd.n2254 30.449
R4198 vdd.n591 vdd.n590 30.449
R4199 vdd.n1421 vdd.n1228 22.6735
R4200 vdd.n1943 vdd.n863 22.6735
R4201 vdd.n2840 vdd.n516 22.6735
R4202 vdd.n3025 vdd.n329 22.6735
R4203 vdd.n1432 vdd.n1190 19.3944
R4204 vdd.n1432 vdd.n1188 19.3944
R4205 vdd.n1436 vdd.n1188 19.3944
R4206 vdd.n1436 vdd.n1178 19.3944
R4207 vdd.n1449 vdd.n1178 19.3944
R4208 vdd.n1449 vdd.n1176 19.3944
R4209 vdd.n1453 vdd.n1176 19.3944
R4210 vdd.n1453 vdd.n1168 19.3944
R4211 vdd.n1467 vdd.n1168 19.3944
R4212 vdd.n1467 vdd.n1166 19.3944
R4213 vdd.n1471 vdd.n1166 19.3944
R4214 vdd.n1471 vdd.n885 19.3944
R4215 vdd.n1483 vdd.n885 19.3944
R4216 vdd.n1483 vdd.n883 19.3944
R4217 vdd.n1487 vdd.n883 19.3944
R4218 vdd.n1487 vdd.n875 19.3944
R4219 vdd.n1500 vdd.n875 19.3944
R4220 vdd.n1500 vdd.n872 19.3944
R4221 vdd.n1506 vdd.n872 19.3944
R4222 vdd.n1506 vdd.n873 19.3944
R4223 vdd.n873 vdd.n862 19.3944
R4224 vdd.n1356 vdd.n1291 19.3944
R4225 vdd.n1352 vdd.n1291 19.3944
R4226 vdd.n1352 vdd.n1351 19.3944
R4227 vdd.n1351 vdd.n1350 19.3944
R4228 vdd.n1350 vdd.n1297 19.3944
R4229 vdd.n1346 vdd.n1297 19.3944
R4230 vdd.n1346 vdd.n1345 19.3944
R4231 vdd.n1345 vdd.n1344 19.3944
R4232 vdd.n1344 vdd.n1303 19.3944
R4233 vdd.n1340 vdd.n1303 19.3944
R4234 vdd.n1340 vdd.n1339 19.3944
R4235 vdd.n1339 vdd.n1338 19.3944
R4236 vdd.n1338 vdd.n1309 19.3944
R4237 vdd.n1334 vdd.n1309 19.3944
R4238 vdd.n1334 vdd.n1333 19.3944
R4239 vdd.n1333 vdd.n1332 19.3944
R4240 vdd.n1332 vdd.n1315 19.3944
R4241 vdd.n1328 vdd.n1315 19.3944
R4242 vdd.n1328 vdd.n1327 19.3944
R4243 vdd.n1327 vdd.n1326 19.3944
R4244 vdd.n1391 vdd.n1390 19.3944
R4245 vdd.n1390 vdd.n1389 19.3944
R4246 vdd.n1389 vdd.n1262 19.3944
R4247 vdd.n1385 vdd.n1262 19.3944
R4248 vdd.n1385 vdd.n1384 19.3944
R4249 vdd.n1384 vdd.n1383 19.3944
R4250 vdd.n1383 vdd.n1268 19.3944
R4251 vdd.n1379 vdd.n1268 19.3944
R4252 vdd.n1379 vdd.n1378 19.3944
R4253 vdd.n1378 vdd.n1377 19.3944
R4254 vdd.n1377 vdd.n1274 19.3944
R4255 vdd.n1373 vdd.n1274 19.3944
R4256 vdd.n1373 vdd.n1372 19.3944
R4257 vdd.n1372 vdd.n1371 19.3944
R4258 vdd.n1371 vdd.n1280 19.3944
R4259 vdd.n1367 vdd.n1280 19.3944
R4260 vdd.n1367 vdd.n1366 19.3944
R4261 vdd.n1366 vdd.n1365 19.3944
R4262 vdd.n1365 vdd.n1286 19.3944
R4263 vdd.n1361 vdd.n1286 19.3944
R4264 vdd.n1424 vdd.n1195 19.3944
R4265 vdd.n1419 vdd.n1195 19.3944
R4266 vdd.n1419 vdd.n1230 19.3944
R4267 vdd.n1415 vdd.n1230 19.3944
R4268 vdd.n1415 vdd.n1414 19.3944
R4269 vdd.n1414 vdd.n1413 19.3944
R4270 vdd.n1413 vdd.n1236 19.3944
R4271 vdd.n1409 vdd.n1236 19.3944
R4272 vdd.n1409 vdd.n1408 19.3944
R4273 vdd.n1408 vdd.n1407 19.3944
R4274 vdd.n1407 vdd.n1242 19.3944
R4275 vdd.n1403 vdd.n1242 19.3944
R4276 vdd.n1403 vdd.n1402 19.3944
R4277 vdd.n1402 vdd.n1401 19.3944
R4278 vdd.n1401 vdd.n1248 19.3944
R4279 vdd.n1397 vdd.n1248 19.3944
R4280 vdd.n1397 vdd.n1396 19.3944
R4281 vdd.n1396 vdd.n1395 19.3944
R4282 vdd.n1648 vdd.n1583 19.3944
R4283 vdd.n1648 vdd.n1589 19.3944
R4284 vdd.n1643 vdd.n1589 19.3944
R4285 vdd.n1643 vdd.n1642 19.3944
R4286 vdd.n1642 vdd.n1641 19.3944
R4287 vdd.n1641 vdd.n1596 19.3944
R4288 vdd.n1636 vdd.n1596 19.3944
R4289 vdd.n1636 vdd.n1635 19.3944
R4290 vdd.n1635 vdd.n1634 19.3944
R4291 vdd.n1634 vdd.n1603 19.3944
R4292 vdd.n1629 vdd.n1603 19.3944
R4293 vdd.n1629 vdd.n1628 19.3944
R4294 vdd.n1628 vdd.n1627 19.3944
R4295 vdd.n1627 vdd.n1611 19.3944
R4296 vdd.n1622 vdd.n1611 19.3944
R4297 vdd.n1622 vdd.n1621 19.3944
R4298 vdd.n1617 vdd.n1616 19.3944
R4299 vdd.n1950 vdd.n858 19.3944
R4300 vdd.n1687 vdd.n1543 19.3944
R4301 vdd.n1687 vdd.n1549 19.3944
R4302 vdd.n1682 vdd.n1549 19.3944
R4303 vdd.n1682 vdd.n1681 19.3944
R4304 vdd.n1681 vdd.n1680 19.3944
R4305 vdd.n1680 vdd.n1556 19.3944
R4306 vdd.n1675 vdd.n1556 19.3944
R4307 vdd.n1675 vdd.n1674 19.3944
R4308 vdd.n1674 vdd.n1673 19.3944
R4309 vdd.n1673 vdd.n1563 19.3944
R4310 vdd.n1668 vdd.n1563 19.3944
R4311 vdd.n1668 vdd.n1667 19.3944
R4312 vdd.n1667 vdd.n1666 19.3944
R4313 vdd.n1666 vdd.n1570 19.3944
R4314 vdd.n1661 vdd.n1570 19.3944
R4315 vdd.n1661 vdd.n1660 19.3944
R4316 vdd.n1660 vdd.n1659 19.3944
R4317 vdd.n1659 vdd.n1577 19.3944
R4318 vdd.n1654 vdd.n1577 19.3944
R4319 vdd.n1654 vdd.n1653 19.3944
R4320 vdd.n1938 vdd.n1937 19.3944
R4321 vdd.n1937 vdd.n1515 19.3944
R4322 vdd.n1932 vdd.n1931 19.3944
R4323 vdd.n1714 vdd.n1519 19.3944
R4324 vdd.n1714 vdd.n1521 19.3944
R4325 vdd.n1524 vdd.n1521 19.3944
R4326 vdd.n1707 vdd.n1524 19.3944
R4327 vdd.n1707 vdd.n1706 19.3944
R4328 vdd.n1706 vdd.n1705 19.3944
R4329 vdd.n1705 vdd.n1530 19.3944
R4330 vdd.n1700 vdd.n1530 19.3944
R4331 vdd.n1700 vdd.n1699 19.3944
R4332 vdd.n1699 vdd.n1698 19.3944
R4333 vdd.n1698 vdd.n1537 19.3944
R4334 vdd.n1693 vdd.n1537 19.3944
R4335 vdd.n1693 vdd.n1692 19.3944
R4336 vdd.n1428 vdd.n1193 19.3944
R4337 vdd.n1428 vdd.n1184 19.3944
R4338 vdd.n1441 vdd.n1184 19.3944
R4339 vdd.n1441 vdd.n1182 19.3944
R4340 vdd.n1445 vdd.n1182 19.3944
R4341 vdd.n1445 vdd.n1173 19.3944
R4342 vdd.n1458 vdd.n1173 19.3944
R4343 vdd.n1458 vdd.n1171 19.3944
R4344 vdd.n1463 vdd.n1171 19.3944
R4345 vdd.n1463 vdd.n1162 19.3944
R4346 vdd.n1475 vdd.n1162 19.3944
R4347 vdd.n1475 vdd.n890 19.3944
R4348 vdd.n1479 vdd.n890 19.3944
R4349 vdd.n1479 vdd.n880 19.3944
R4350 vdd.n1492 vdd.n880 19.3944
R4351 vdd.n1492 vdd.n878 19.3944
R4352 vdd.n1496 vdd.n878 19.3944
R4353 vdd.n1496 vdd.n868 19.3944
R4354 vdd.n1511 vdd.n868 19.3944
R4355 vdd.n1511 vdd.n866 19.3944
R4356 vdd.n1941 vdd.n866 19.3944
R4357 vdd.n2851 vdd.n477 19.3944
R4358 vdd.n2851 vdd.n475 19.3944
R4359 vdd.n2855 vdd.n475 19.3944
R4360 vdd.n2855 vdd.n465 19.3944
R4361 vdd.n2868 vdd.n465 19.3944
R4362 vdd.n2868 vdd.n463 19.3944
R4363 vdd.n2872 vdd.n463 19.3944
R4364 vdd.n2872 vdd.n453 19.3944
R4365 vdd.n2884 vdd.n453 19.3944
R4366 vdd.n2884 vdd.n451 19.3944
R4367 vdd.n2888 vdd.n451 19.3944
R4368 vdd.n2889 vdd.n2888 19.3944
R4369 vdd.n2890 vdd.n2889 19.3944
R4370 vdd.n2890 vdd.n449 19.3944
R4371 vdd.n2894 vdd.n449 19.3944
R4372 vdd.n2895 vdd.n2894 19.3944
R4373 vdd.n2896 vdd.n2895 19.3944
R4374 vdd.n2896 vdd.n446 19.3944
R4375 vdd.n2900 vdd.n446 19.3944
R4376 vdd.n2901 vdd.n2900 19.3944
R4377 vdd.n2902 vdd.n2901 19.3944
R4378 vdd.n2945 vdd.n404 19.3944
R4379 vdd.n2945 vdd.n410 19.3944
R4380 vdd.n2940 vdd.n410 19.3944
R4381 vdd.n2940 vdd.n2939 19.3944
R4382 vdd.n2939 vdd.n2938 19.3944
R4383 vdd.n2938 vdd.n417 19.3944
R4384 vdd.n2933 vdd.n417 19.3944
R4385 vdd.n2933 vdd.n2932 19.3944
R4386 vdd.n2932 vdd.n2931 19.3944
R4387 vdd.n2931 vdd.n424 19.3944
R4388 vdd.n2926 vdd.n424 19.3944
R4389 vdd.n2926 vdd.n2925 19.3944
R4390 vdd.n2925 vdd.n2924 19.3944
R4391 vdd.n2924 vdd.n431 19.3944
R4392 vdd.n2919 vdd.n431 19.3944
R4393 vdd.n2919 vdd.n2918 19.3944
R4394 vdd.n2918 vdd.n2917 19.3944
R4395 vdd.n2917 vdd.n438 19.3944
R4396 vdd.n2912 vdd.n438 19.3944
R4397 vdd.n2912 vdd.n2911 19.3944
R4398 vdd.n2984 vdd.n364 19.3944
R4399 vdd.n2984 vdd.n370 19.3944
R4400 vdd.n2979 vdd.n370 19.3944
R4401 vdd.n2979 vdd.n2978 19.3944
R4402 vdd.n2978 vdd.n2977 19.3944
R4403 vdd.n2977 vdd.n377 19.3944
R4404 vdd.n2972 vdd.n377 19.3944
R4405 vdd.n2972 vdd.n2971 19.3944
R4406 vdd.n2971 vdd.n2970 19.3944
R4407 vdd.n2970 vdd.n384 19.3944
R4408 vdd.n2965 vdd.n384 19.3944
R4409 vdd.n2965 vdd.n2964 19.3944
R4410 vdd.n2964 vdd.n2963 19.3944
R4411 vdd.n2963 vdd.n391 19.3944
R4412 vdd.n2958 vdd.n391 19.3944
R4413 vdd.n2958 vdd.n2957 19.3944
R4414 vdd.n2957 vdd.n2956 19.3944
R4415 vdd.n2956 vdd.n398 19.3944
R4416 vdd.n2951 vdd.n398 19.3944
R4417 vdd.n2951 vdd.n2950 19.3944
R4418 vdd.n3020 vdd.n3019 19.3944
R4419 vdd.n3019 vdd.n3018 19.3944
R4420 vdd.n3018 vdd.n336 19.3944
R4421 vdd.n337 vdd.n336 19.3944
R4422 vdd.n3011 vdd.n337 19.3944
R4423 vdd.n3011 vdd.n3010 19.3944
R4424 vdd.n3010 vdd.n3009 19.3944
R4425 vdd.n3009 vdd.n344 19.3944
R4426 vdd.n3004 vdd.n344 19.3944
R4427 vdd.n3004 vdd.n3003 19.3944
R4428 vdd.n3003 vdd.n3002 19.3944
R4429 vdd.n3002 vdd.n351 19.3944
R4430 vdd.n2997 vdd.n351 19.3944
R4431 vdd.n2997 vdd.n2996 19.3944
R4432 vdd.n2996 vdd.n2995 19.3944
R4433 vdd.n2995 vdd.n358 19.3944
R4434 vdd.n2990 vdd.n358 19.3944
R4435 vdd.n2990 vdd.n2989 19.3944
R4436 vdd.n2847 vdd.n480 19.3944
R4437 vdd.n2847 vdd.n471 19.3944
R4438 vdd.n2860 vdd.n471 19.3944
R4439 vdd.n2860 vdd.n469 19.3944
R4440 vdd.n2864 vdd.n469 19.3944
R4441 vdd.n2864 vdd.n460 19.3944
R4442 vdd.n2876 vdd.n460 19.3944
R4443 vdd.n2876 vdd.n458 19.3944
R4444 vdd.n2880 vdd.n458 19.3944
R4445 vdd.n2880 vdd.n300 19.3944
R4446 vdd.n3045 vdd.n300 19.3944
R4447 vdd.n3045 vdd.n301 19.3944
R4448 vdd.n3039 vdd.n301 19.3944
R4449 vdd.n3039 vdd.n3038 19.3944
R4450 vdd.n3038 vdd.n3037 19.3944
R4451 vdd.n3037 vdd.n313 19.3944
R4452 vdd.n3031 vdd.n313 19.3944
R4453 vdd.n3031 vdd.n3030 19.3944
R4454 vdd.n3030 vdd.n3029 19.3944
R4455 vdd.n3029 vdd.n324 19.3944
R4456 vdd.n3023 vdd.n324 19.3944
R4457 vdd.n2800 vdd.n536 19.3944
R4458 vdd.n2800 vdd.n2797 19.3944
R4459 vdd.n2797 vdd.n2794 19.3944
R4460 vdd.n2794 vdd.n2793 19.3944
R4461 vdd.n2793 vdd.n2790 19.3944
R4462 vdd.n2790 vdd.n2789 19.3944
R4463 vdd.n2789 vdd.n2786 19.3944
R4464 vdd.n2786 vdd.n2785 19.3944
R4465 vdd.n2785 vdd.n2782 19.3944
R4466 vdd.n2782 vdd.n2781 19.3944
R4467 vdd.n2781 vdd.n2778 19.3944
R4468 vdd.n2778 vdd.n2777 19.3944
R4469 vdd.n2777 vdd.n2774 19.3944
R4470 vdd.n2774 vdd.n2773 19.3944
R4471 vdd.n2773 vdd.n2770 19.3944
R4472 vdd.n2770 vdd.n2769 19.3944
R4473 vdd.n2769 vdd.n2766 19.3944
R4474 vdd.n2766 vdd.n2765 19.3944
R4475 vdd.n2765 vdd.n2762 19.3944
R4476 vdd.n2762 vdd.n2761 19.3944
R4477 vdd.n2843 vdd.n482 19.3944
R4478 vdd.n2838 vdd.n482 19.3944
R4479 vdd.n521 vdd.n518 19.3944
R4480 vdd.n2834 vdd.n2833 19.3944
R4481 vdd.n2833 vdd.n2830 19.3944
R4482 vdd.n2830 vdd.n2829 19.3944
R4483 vdd.n2829 vdd.n2826 19.3944
R4484 vdd.n2826 vdd.n2825 19.3944
R4485 vdd.n2825 vdd.n2822 19.3944
R4486 vdd.n2822 vdd.n2821 19.3944
R4487 vdd.n2821 vdd.n2818 19.3944
R4488 vdd.n2818 vdd.n2817 19.3944
R4489 vdd.n2817 vdd.n2814 19.3944
R4490 vdd.n2814 vdd.n2813 19.3944
R4491 vdd.n2813 vdd.n2810 19.3944
R4492 vdd.n2810 vdd.n2809 19.3944
R4493 vdd.n2754 vdd.n556 19.3944
R4494 vdd.n2754 vdd.n2751 19.3944
R4495 vdd.n2751 vdd.n2748 19.3944
R4496 vdd.n2748 vdd.n2747 19.3944
R4497 vdd.n2747 vdd.n2744 19.3944
R4498 vdd.n2744 vdd.n2743 19.3944
R4499 vdd.n2743 vdd.n2740 19.3944
R4500 vdd.n2740 vdd.n2739 19.3944
R4501 vdd.n2739 vdd.n2736 19.3944
R4502 vdd.n2736 vdd.n2735 19.3944
R4503 vdd.n2735 vdd.n2732 19.3944
R4504 vdd.n2732 vdd.n2731 19.3944
R4505 vdd.n2731 vdd.n2728 19.3944
R4506 vdd.n2728 vdd.n2727 19.3944
R4507 vdd.n2727 vdd.n2724 19.3944
R4508 vdd.n2724 vdd.n2723 19.3944
R4509 vdd.n2720 vdd.n2719 19.3944
R4510 vdd.n2716 vdd.n2715 19.3944
R4511 vdd.n1360 vdd.n1356 19.0066
R4512 vdd.n1652 vdd.n1583 19.0066
R4513 vdd.n2949 vdd.n404 19.0066
R4514 vdd.n2758 vdd.n556 19.0066
R4515 vdd.n1792 vdd.n1791 16.0975
R4516 vdd.n756 vdd.n755 16.0975
R4517 vdd.n1321 vdd.n1320 16.0975
R4518 vdd.n1359 vdd.n1358 16.0975
R4519 vdd.n1255 vdd.n1254 16.0975
R4520 vdd.n1948 vdd.n1947 16.0975
R4521 vdd.n1585 vdd.n1584 16.0975
R4522 vdd.n1545 vdd.n1544 16.0975
R4523 vdd.n1766 vdd.n1765 16.0975
R4524 vdd.n748 vdd.n747 16.0975
R4525 vdd.n2257 vdd.n2256 16.0975
R4526 vdd.n2909 vdd.n2908 16.0975
R4527 vdd.n406 vdd.n405 16.0975
R4528 vdd.n366 vdd.n365 16.0975
R4529 vdd.n558 vdd.n557 16.0975
R4530 vdd.n2805 vdd.n2804 16.0975
R4531 vdd.n623 vdd.n622 16.0975
R4532 vdd.n2254 vdd.n2253 16.0975
R4533 vdd.n2712 vdd.n2711 16.0975
R4534 vdd.n590 vdd.n589 16.0975
R4535 vdd.t118 vdd.n2218 15.4182
R4536 vdd.n2471 vdd.t22 15.4182
R4537 vdd.n28 vdd.n27 15.0023
R4538 vdd.n1989 vdd.n839 14.5112
R4539 vdd.n2673 vdd.n484 14.5112
R4540 vdd.n292 vdd.n257 13.1884
R4541 vdd.n245 vdd.n210 13.1884
R4542 vdd.n202 vdd.n167 13.1884
R4543 vdd.n155 vdd.n120 13.1884
R4544 vdd.n113 vdd.n78 13.1884
R4545 vdd.n66 vdd.n31 13.1884
R4546 vdd.n1107 vdd.n1072 13.1884
R4547 vdd.n1154 vdd.n1119 13.1884
R4548 vdd.n1017 vdd.n982 13.1884
R4549 vdd.n1064 vdd.n1029 13.1884
R4550 vdd.n928 vdd.n893 13.1884
R4551 vdd.n975 vdd.n940 13.1884
R4552 vdd.n1391 vdd.n1256 12.9944
R4553 vdd.n1395 vdd.n1256 12.9944
R4554 vdd.n1691 vdd.n1543 12.9944
R4555 vdd.n1692 vdd.n1691 12.9944
R4556 vdd.n2988 vdd.n364 12.9944
R4557 vdd.n2989 vdd.n2988 12.9944
R4558 vdd.n2806 vdd.n536 12.9944
R4559 vdd.n2809 vdd.n2806 12.9944
R4560 vdd.n293 vdd.n255 12.8005
R4561 vdd.n288 vdd.n259 12.8005
R4562 vdd.n246 vdd.n208 12.8005
R4563 vdd.n241 vdd.n212 12.8005
R4564 vdd.n203 vdd.n165 12.8005
R4565 vdd.n198 vdd.n169 12.8005
R4566 vdd.n156 vdd.n118 12.8005
R4567 vdd.n151 vdd.n122 12.8005
R4568 vdd.n114 vdd.n76 12.8005
R4569 vdd.n109 vdd.n80 12.8005
R4570 vdd.n67 vdd.n29 12.8005
R4571 vdd.n62 vdd.n33 12.8005
R4572 vdd.n1108 vdd.n1070 12.8005
R4573 vdd.n1103 vdd.n1074 12.8005
R4574 vdd.n1155 vdd.n1117 12.8005
R4575 vdd.n1150 vdd.n1121 12.8005
R4576 vdd.n1018 vdd.n980 12.8005
R4577 vdd.n1013 vdd.n984 12.8005
R4578 vdd.n1065 vdd.n1027 12.8005
R4579 vdd.n1060 vdd.n1031 12.8005
R4580 vdd.n929 vdd.n891 12.8005
R4581 vdd.n924 vdd.n895 12.8005
R4582 vdd.n976 vdd.n938 12.8005
R4583 vdd.n971 vdd.n942 12.8005
R4584 vdd.n287 vdd.n260 12.0247
R4585 vdd.n240 vdd.n213 12.0247
R4586 vdd.n197 vdd.n170 12.0247
R4587 vdd.n150 vdd.n123 12.0247
R4588 vdd.n108 vdd.n81 12.0247
R4589 vdd.n61 vdd.n34 12.0247
R4590 vdd.n1102 vdd.n1075 12.0247
R4591 vdd.n1149 vdd.n1122 12.0247
R4592 vdd.n1012 vdd.n985 12.0247
R4593 vdd.n1059 vdd.n1032 12.0247
R4594 vdd.n923 vdd.n896 12.0247
R4595 vdd.n970 vdd.n943 12.0247
R4596 vdd.n1430 vdd.n1186 11.337
R4597 vdd.n1439 vdd.n1186 11.337
R4598 vdd.n1439 vdd.n1438 11.337
R4599 vdd.n1447 vdd.n1180 11.337
R4600 vdd.n1456 vdd.n1455 11.337
R4601 vdd.n1473 vdd.n1164 11.337
R4602 vdd.n1481 vdd.n887 11.337
R4603 vdd.n1490 vdd.n1489 11.337
R4604 vdd.n1498 vdd.n870 11.337
R4605 vdd.n1509 vdd.n870 11.337
R4606 vdd.n1509 vdd.n1508 11.337
R4607 vdd.n2849 vdd.n473 11.337
R4608 vdd.n2858 vdd.n473 11.337
R4609 vdd.n2858 vdd.n2857 11.337
R4610 vdd.n2866 vdd.n467 11.337
R4611 vdd.n2882 vdd.n456 11.337
R4612 vdd.n3043 vdd.n304 11.337
R4613 vdd.n3041 vdd.n308 11.337
R4614 vdd.n3035 vdd.n3034 11.337
R4615 vdd.n3033 vdd.n318 11.337
R4616 vdd.n3027 vdd.n318 11.337
R4617 vdd.n3027 vdd.n3026 11.337
R4618 vdd.n284 vdd.n283 11.249
R4619 vdd.n237 vdd.n236 11.249
R4620 vdd.n194 vdd.n193 11.249
R4621 vdd.n147 vdd.n146 11.249
R4622 vdd.n105 vdd.n104 11.249
R4623 vdd.n58 vdd.n57 11.249
R4624 vdd.n1099 vdd.n1098 11.249
R4625 vdd.n1146 vdd.n1145 11.249
R4626 vdd.n1009 vdd.n1008 11.249
R4627 vdd.n1056 vdd.n1055 11.249
R4628 vdd.n920 vdd.n919 11.249
R4629 vdd.n967 vdd.n966 11.249
R4630 vdd.n2146 vdd.t114 11.1103
R4631 vdd.n2478 vdd.t188 11.1103
R4632 vdd.n1228 vdd.t44 10.7702
R4633 vdd.t55 vdd.n3025 10.7702
R4634 vdd.n269 vdd.n268 10.7238
R4635 vdd.n222 vdd.n221 10.7238
R4636 vdd.n179 vdd.n178 10.7238
R4637 vdd.n132 vdd.n131 10.7238
R4638 vdd.n90 vdd.n89 10.7238
R4639 vdd.n43 vdd.n42 10.7238
R4640 vdd.n1084 vdd.n1083 10.7238
R4641 vdd.n1131 vdd.n1130 10.7238
R4642 vdd.n994 vdd.n993 10.7238
R4643 vdd.n1041 vdd.n1040 10.7238
R4644 vdd.n905 vdd.n904 10.7238
R4645 vdd.n952 vdd.n951 10.7238
R4646 vdd.n1992 vdd.n1991 10.6151
R4647 vdd.n1993 vdd.n1992 10.6151
R4648 vdd.n1993 vdd.n825 10.6151
R4649 vdd.n2003 vdd.n825 10.6151
R4650 vdd.n2004 vdd.n2003 10.6151
R4651 vdd.n2005 vdd.n2004 10.6151
R4652 vdd.n2005 vdd.n812 10.6151
R4653 vdd.n2016 vdd.n812 10.6151
R4654 vdd.n2017 vdd.n2016 10.6151
R4655 vdd.n2018 vdd.n2017 10.6151
R4656 vdd.n2018 vdd.n800 10.6151
R4657 vdd.n2028 vdd.n800 10.6151
R4658 vdd.n2029 vdd.n2028 10.6151
R4659 vdd.n2030 vdd.n2029 10.6151
R4660 vdd.n2030 vdd.n788 10.6151
R4661 vdd.n2040 vdd.n788 10.6151
R4662 vdd.n2041 vdd.n2040 10.6151
R4663 vdd.n2042 vdd.n2041 10.6151
R4664 vdd.n2042 vdd.n777 10.6151
R4665 vdd.n2052 vdd.n777 10.6151
R4666 vdd.n2053 vdd.n2052 10.6151
R4667 vdd.n2054 vdd.n2053 10.6151
R4668 vdd.n2054 vdd.n764 10.6151
R4669 vdd.n2066 vdd.n764 10.6151
R4670 vdd.n2067 vdd.n2066 10.6151
R4671 vdd.n2069 vdd.n2067 10.6151
R4672 vdd.n2069 vdd.n2068 10.6151
R4673 vdd.n2068 vdd.n746 10.6151
R4674 vdd.n2216 vdd.n2215 10.6151
R4675 vdd.n2215 vdd.n2214 10.6151
R4676 vdd.n2214 vdd.n2211 10.6151
R4677 vdd.n2211 vdd.n2210 10.6151
R4678 vdd.n2210 vdd.n2207 10.6151
R4679 vdd.n2207 vdd.n2206 10.6151
R4680 vdd.n2206 vdd.n2203 10.6151
R4681 vdd.n2203 vdd.n2202 10.6151
R4682 vdd.n2202 vdd.n2199 10.6151
R4683 vdd.n2199 vdd.n2198 10.6151
R4684 vdd.n2198 vdd.n2195 10.6151
R4685 vdd.n2195 vdd.n2194 10.6151
R4686 vdd.n2194 vdd.n2191 10.6151
R4687 vdd.n2191 vdd.n2190 10.6151
R4688 vdd.n2190 vdd.n2187 10.6151
R4689 vdd.n2187 vdd.n2186 10.6151
R4690 vdd.n2186 vdd.n2183 10.6151
R4691 vdd.n2183 vdd.n2182 10.6151
R4692 vdd.n2182 vdd.n2179 10.6151
R4693 vdd.n2179 vdd.n2178 10.6151
R4694 vdd.n2178 vdd.n2175 10.6151
R4695 vdd.n2175 vdd.n2174 10.6151
R4696 vdd.n2174 vdd.n2171 10.6151
R4697 vdd.n2171 vdd.n2170 10.6151
R4698 vdd.n2170 vdd.n2167 10.6151
R4699 vdd.n2167 vdd.n2166 10.6151
R4700 vdd.n2166 vdd.n2163 10.6151
R4701 vdd.n2163 vdd.n2162 10.6151
R4702 vdd.n2162 vdd.n2159 10.6151
R4703 vdd.n2159 vdd.n2158 10.6151
R4704 vdd.n2158 vdd.n2155 10.6151
R4705 vdd.n2153 vdd.n2150 10.6151
R4706 vdd.n2150 vdd.n2149 10.6151
R4707 vdd.n1892 vdd.n1891 10.6151
R4708 vdd.n1891 vdd.n1889 10.6151
R4709 vdd.n1889 vdd.n1888 10.6151
R4710 vdd.n1888 vdd.n1886 10.6151
R4711 vdd.n1886 vdd.n1885 10.6151
R4712 vdd.n1885 vdd.n1883 10.6151
R4713 vdd.n1883 vdd.n1882 10.6151
R4714 vdd.n1882 vdd.n1880 10.6151
R4715 vdd.n1880 vdd.n1879 10.6151
R4716 vdd.n1879 vdd.n1877 10.6151
R4717 vdd.n1877 vdd.n1876 10.6151
R4718 vdd.n1876 vdd.n1874 10.6151
R4719 vdd.n1874 vdd.n1873 10.6151
R4720 vdd.n1873 vdd.n1788 10.6151
R4721 vdd.n1788 vdd.n1787 10.6151
R4722 vdd.n1787 vdd.n1785 10.6151
R4723 vdd.n1785 vdd.n1784 10.6151
R4724 vdd.n1784 vdd.n1782 10.6151
R4725 vdd.n1782 vdd.n1781 10.6151
R4726 vdd.n1781 vdd.n1779 10.6151
R4727 vdd.n1779 vdd.n1778 10.6151
R4728 vdd.n1778 vdd.n1776 10.6151
R4729 vdd.n1776 vdd.n1775 10.6151
R4730 vdd.n1775 vdd.n1773 10.6151
R4731 vdd.n1773 vdd.n1772 10.6151
R4732 vdd.n1772 vdd.n1769 10.6151
R4733 vdd.n1769 vdd.n1768 10.6151
R4734 vdd.n1768 vdd.n749 10.6151
R4735 vdd.n1726 vdd.n837 10.6151
R4736 vdd.n1727 vdd.n1726 10.6151
R4737 vdd.n1728 vdd.n1727 10.6151
R4738 vdd.n1728 vdd.n1722 10.6151
R4739 vdd.n1734 vdd.n1722 10.6151
R4740 vdd.n1735 vdd.n1734 10.6151
R4741 vdd.n1736 vdd.n1735 10.6151
R4742 vdd.n1736 vdd.n1720 10.6151
R4743 vdd.n1742 vdd.n1720 10.6151
R4744 vdd.n1743 vdd.n1742 10.6151
R4745 vdd.n1744 vdd.n1743 10.6151
R4746 vdd.n1744 vdd.n1718 10.6151
R4747 vdd.n1750 vdd.n1718 10.6151
R4748 vdd.n1751 vdd.n1750 10.6151
R4749 vdd.n1752 vdd.n1751 10.6151
R4750 vdd.n1752 vdd.n1716 10.6151
R4751 vdd.n1928 vdd.n1716 10.6151
R4752 vdd.n1928 vdd.n1927 10.6151
R4753 vdd.n1927 vdd.n1757 10.6151
R4754 vdd.n1921 vdd.n1757 10.6151
R4755 vdd.n1921 vdd.n1920 10.6151
R4756 vdd.n1920 vdd.n1919 10.6151
R4757 vdd.n1919 vdd.n1759 10.6151
R4758 vdd.n1913 vdd.n1759 10.6151
R4759 vdd.n1913 vdd.n1912 10.6151
R4760 vdd.n1912 vdd.n1911 10.6151
R4761 vdd.n1911 vdd.n1761 10.6151
R4762 vdd.n1905 vdd.n1761 10.6151
R4763 vdd.n1905 vdd.n1904 10.6151
R4764 vdd.n1904 vdd.n1903 10.6151
R4765 vdd.n1903 vdd.n1763 10.6151
R4766 vdd.n1897 vdd.n1896 10.6151
R4767 vdd.n1896 vdd.n1895 10.6151
R4768 vdd.n2401 vdd.n2400 10.6151
R4769 vdd.n2400 vdd.n2398 10.6151
R4770 vdd.n2398 vdd.n2397 10.6151
R4771 vdd.n2397 vdd.n2255 10.6151
R4772 vdd.n2344 vdd.n2255 10.6151
R4773 vdd.n2345 vdd.n2344 10.6151
R4774 vdd.n2347 vdd.n2345 10.6151
R4775 vdd.n2348 vdd.n2347 10.6151
R4776 vdd.n2350 vdd.n2348 10.6151
R4777 vdd.n2351 vdd.n2350 10.6151
R4778 vdd.n2353 vdd.n2351 10.6151
R4779 vdd.n2354 vdd.n2353 10.6151
R4780 vdd.n2356 vdd.n2354 10.6151
R4781 vdd.n2357 vdd.n2356 10.6151
R4782 vdd.n2372 vdd.n2357 10.6151
R4783 vdd.n2372 vdd.n2371 10.6151
R4784 vdd.n2371 vdd.n2370 10.6151
R4785 vdd.n2370 vdd.n2368 10.6151
R4786 vdd.n2368 vdd.n2367 10.6151
R4787 vdd.n2367 vdd.n2365 10.6151
R4788 vdd.n2365 vdd.n2364 10.6151
R4789 vdd.n2364 vdd.n2362 10.6151
R4790 vdd.n2362 vdd.n2361 10.6151
R4791 vdd.n2361 vdd.n2359 10.6151
R4792 vdd.n2359 vdd.n2358 10.6151
R4793 vdd.n2358 vdd.n626 10.6151
R4794 vdd.n2606 vdd.n626 10.6151
R4795 vdd.n2607 vdd.n2606 10.6151
R4796 vdd.n2468 vdd.n702 10.6151
R4797 vdd.n2468 vdd.n2467 10.6151
R4798 vdd.n2467 vdd.n2466 10.6151
R4799 vdd.n2466 vdd.n2464 10.6151
R4800 vdd.n2464 vdd.n2461 10.6151
R4801 vdd.n2461 vdd.n2460 10.6151
R4802 vdd.n2460 vdd.n2457 10.6151
R4803 vdd.n2457 vdd.n2456 10.6151
R4804 vdd.n2456 vdd.n2453 10.6151
R4805 vdd.n2453 vdd.n2452 10.6151
R4806 vdd.n2452 vdd.n2449 10.6151
R4807 vdd.n2449 vdd.n2448 10.6151
R4808 vdd.n2448 vdd.n2445 10.6151
R4809 vdd.n2445 vdd.n2444 10.6151
R4810 vdd.n2444 vdd.n2441 10.6151
R4811 vdd.n2441 vdd.n2440 10.6151
R4812 vdd.n2440 vdd.n2437 10.6151
R4813 vdd.n2437 vdd.n2436 10.6151
R4814 vdd.n2436 vdd.n2433 10.6151
R4815 vdd.n2433 vdd.n2432 10.6151
R4816 vdd.n2432 vdd.n2429 10.6151
R4817 vdd.n2429 vdd.n2428 10.6151
R4818 vdd.n2428 vdd.n2425 10.6151
R4819 vdd.n2425 vdd.n2424 10.6151
R4820 vdd.n2424 vdd.n2421 10.6151
R4821 vdd.n2421 vdd.n2420 10.6151
R4822 vdd.n2420 vdd.n2417 10.6151
R4823 vdd.n2417 vdd.n2416 10.6151
R4824 vdd.n2416 vdd.n2413 10.6151
R4825 vdd.n2413 vdd.n2412 10.6151
R4826 vdd.n2412 vdd.n2409 10.6151
R4827 vdd.n2407 vdd.n2404 10.6151
R4828 vdd.n2404 vdd.n2403 10.6151
R4829 vdd.n2481 vdd.n2480 10.6151
R4830 vdd.n2482 vdd.n2481 10.6151
R4831 vdd.n2482 vdd.n692 10.6151
R4832 vdd.n2492 vdd.n692 10.6151
R4833 vdd.n2493 vdd.n2492 10.6151
R4834 vdd.n2494 vdd.n2493 10.6151
R4835 vdd.n2494 vdd.n679 10.6151
R4836 vdd.n2504 vdd.n679 10.6151
R4837 vdd.n2505 vdd.n2504 10.6151
R4838 vdd.n2506 vdd.n2505 10.6151
R4839 vdd.n2506 vdd.n668 10.6151
R4840 vdd.n2516 vdd.n668 10.6151
R4841 vdd.n2517 vdd.n2516 10.6151
R4842 vdd.n2518 vdd.n2517 10.6151
R4843 vdd.n2518 vdd.n656 10.6151
R4844 vdd.n2528 vdd.n656 10.6151
R4845 vdd.n2529 vdd.n2528 10.6151
R4846 vdd.n2530 vdd.n2529 10.6151
R4847 vdd.n2530 vdd.n645 10.6151
R4848 vdd.n2542 vdd.n645 10.6151
R4849 vdd.n2543 vdd.n2542 10.6151
R4850 vdd.n2544 vdd.n2543 10.6151
R4851 vdd.n2544 vdd.n631 10.6151
R4852 vdd.n2599 vdd.n631 10.6151
R4853 vdd.n2600 vdd.n2599 10.6151
R4854 vdd.n2601 vdd.n2600 10.6151
R4855 vdd.n2601 vdd.n600 10.6151
R4856 vdd.n2671 vdd.n600 10.6151
R4857 vdd.n2670 vdd.n2669 10.6151
R4858 vdd.n2669 vdd.n601 10.6151
R4859 vdd.n602 vdd.n601 10.6151
R4860 vdd.n2662 vdd.n602 10.6151
R4861 vdd.n2662 vdd.n2661 10.6151
R4862 vdd.n2661 vdd.n2660 10.6151
R4863 vdd.n2660 vdd.n604 10.6151
R4864 vdd.n2655 vdd.n604 10.6151
R4865 vdd.n2655 vdd.n2654 10.6151
R4866 vdd.n2654 vdd.n2653 10.6151
R4867 vdd.n2653 vdd.n607 10.6151
R4868 vdd.n2648 vdd.n607 10.6151
R4869 vdd.n2648 vdd.n2647 10.6151
R4870 vdd.n2647 vdd.n2646 10.6151
R4871 vdd.n2646 vdd.n610 10.6151
R4872 vdd.n2641 vdd.n610 10.6151
R4873 vdd.n2641 vdd.n520 10.6151
R4874 vdd.n2637 vdd.n520 10.6151
R4875 vdd.n2637 vdd.n2636 10.6151
R4876 vdd.n2636 vdd.n2635 10.6151
R4877 vdd.n2635 vdd.n613 10.6151
R4878 vdd.n2630 vdd.n613 10.6151
R4879 vdd.n2630 vdd.n2629 10.6151
R4880 vdd.n2629 vdd.n2628 10.6151
R4881 vdd.n2628 vdd.n616 10.6151
R4882 vdd.n2623 vdd.n616 10.6151
R4883 vdd.n2623 vdd.n2622 10.6151
R4884 vdd.n2622 vdd.n2621 10.6151
R4885 vdd.n2621 vdd.n619 10.6151
R4886 vdd.n2616 vdd.n619 10.6151
R4887 vdd.n2616 vdd.n2615 10.6151
R4888 vdd.n2613 vdd.n624 10.6151
R4889 vdd.n2608 vdd.n624 10.6151
R4890 vdd.n2589 vdd.n2550 10.6151
R4891 vdd.n2584 vdd.n2550 10.6151
R4892 vdd.n2584 vdd.n2583 10.6151
R4893 vdd.n2583 vdd.n2582 10.6151
R4894 vdd.n2582 vdd.n2552 10.6151
R4895 vdd.n2577 vdd.n2552 10.6151
R4896 vdd.n2577 vdd.n2576 10.6151
R4897 vdd.n2576 vdd.n2575 10.6151
R4898 vdd.n2575 vdd.n2555 10.6151
R4899 vdd.n2570 vdd.n2555 10.6151
R4900 vdd.n2570 vdd.n2569 10.6151
R4901 vdd.n2569 vdd.n2568 10.6151
R4902 vdd.n2568 vdd.n2558 10.6151
R4903 vdd.n2563 vdd.n2558 10.6151
R4904 vdd.n2563 vdd.n2562 10.6151
R4905 vdd.n2562 vdd.n575 10.6151
R4906 vdd.n2706 vdd.n575 10.6151
R4907 vdd.n2706 vdd.n576 10.6151
R4908 vdd.n578 vdd.n576 10.6151
R4909 vdd.n2699 vdd.n578 10.6151
R4910 vdd.n2699 vdd.n2698 10.6151
R4911 vdd.n2698 vdd.n2697 10.6151
R4912 vdd.n2697 vdd.n580 10.6151
R4913 vdd.n2692 vdd.n580 10.6151
R4914 vdd.n2692 vdd.n2691 10.6151
R4915 vdd.n2691 vdd.n2690 10.6151
R4916 vdd.n2690 vdd.n583 10.6151
R4917 vdd.n2685 vdd.n583 10.6151
R4918 vdd.n2685 vdd.n2684 10.6151
R4919 vdd.n2684 vdd.n2683 10.6151
R4920 vdd.n2683 vdd.n586 10.6151
R4921 vdd.n2678 vdd.n2677 10.6151
R4922 vdd.n2677 vdd.n2676 10.6151
R4923 vdd.n2324 vdd.n2322 10.6151
R4924 vdd.n2325 vdd.n2324 10.6151
R4925 vdd.n2393 vdd.n2325 10.6151
R4926 vdd.n2393 vdd.n2392 10.6151
R4927 vdd.n2392 vdd.n2391 10.6151
R4928 vdd.n2391 vdd.n2389 10.6151
R4929 vdd.n2389 vdd.n2388 10.6151
R4930 vdd.n2388 vdd.n2386 10.6151
R4931 vdd.n2386 vdd.n2385 10.6151
R4932 vdd.n2385 vdd.n2383 10.6151
R4933 vdd.n2383 vdd.n2382 10.6151
R4934 vdd.n2382 vdd.n2380 10.6151
R4935 vdd.n2380 vdd.n2379 10.6151
R4936 vdd.n2379 vdd.n2377 10.6151
R4937 vdd.n2377 vdd.n2376 10.6151
R4938 vdd.n2376 vdd.n2342 10.6151
R4939 vdd.n2342 vdd.n2341 10.6151
R4940 vdd.n2341 vdd.n2339 10.6151
R4941 vdd.n2339 vdd.n2338 10.6151
R4942 vdd.n2338 vdd.n2336 10.6151
R4943 vdd.n2336 vdd.n2335 10.6151
R4944 vdd.n2335 vdd.n2333 10.6151
R4945 vdd.n2333 vdd.n2332 10.6151
R4946 vdd.n2332 vdd.n2330 10.6151
R4947 vdd.n2330 vdd.n2329 10.6151
R4948 vdd.n2329 vdd.n2327 10.6151
R4949 vdd.n2327 vdd.n2326 10.6151
R4950 vdd.n2326 vdd.n592 10.6151
R4951 vdd.n2475 vdd.n2474 10.6151
R4952 vdd.n2474 vdd.n707 10.6151
R4953 vdd.n2259 vdd.n707 10.6151
R4954 vdd.n2262 vdd.n2259 10.6151
R4955 vdd.n2263 vdd.n2262 10.6151
R4956 vdd.n2266 vdd.n2263 10.6151
R4957 vdd.n2267 vdd.n2266 10.6151
R4958 vdd.n2270 vdd.n2267 10.6151
R4959 vdd.n2271 vdd.n2270 10.6151
R4960 vdd.n2274 vdd.n2271 10.6151
R4961 vdd.n2275 vdd.n2274 10.6151
R4962 vdd.n2278 vdd.n2275 10.6151
R4963 vdd.n2279 vdd.n2278 10.6151
R4964 vdd.n2282 vdd.n2279 10.6151
R4965 vdd.n2283 vdd.n2282 10.6151
R4966 vdd.n2286 vdd.n2283 10.6151
R4967 vdd.n2287 vdd.n2286 10.6151
R4968 vdd.n2290 vdd.n2287 10.6151
R4969 vdd.n2291 vdd.n2290 10.6151
R4970 vdd.n2294 vdd.n2291 10.6151
R4971 vdd.n2295 vdd.n2294 10.6151
R4972 vdd.n2298 vdd.n2295 10.6151
R4973 vdd.n2299 vdd.n2298 10.6151
R4974 vdd.n2302 vdd.n2299 10.6151
R4975 vdd.n2303 vdd.n2302 10.6151
R4976 vdd.n2306 vdd.n2303 10.6151
R4977 vdd.n2307 vdd.n2306 10.6151
R4978 vdd.n2310 vdd.n2307 10.6151
R4979 vdd.n2311 vdd.n2310 10.6151
R4980 vdd.n2314 vdd.n2311 10.6151
R4981 vdd.n2315 vdd.n2314 10.6151
R4982 vdd.n2320 vdd.n2318 10.6151
R4983 vdd.n2321 vdd.n2320 10.6151
R4984 vdd.n2476 vdd.n697 10.6151
R4985 vdd.n2486 vdd.n697 10.6151
R4986 vdd.n2487 vdd.n2486 10.6151
R4987 vdd.n2488 vdd.n2487 10.6151
R4988 vdd.n2488 vdd.n685 10.6151
R4989 vdd.n2498 vdd.n685 10.6151
R4990 vdd.n2499 vdd.n2498 10.6151
R4991 vdd.n2500 vdd.n2499 10.6151
R4992 vdd.n2500 vdd.n674 10.6151
R4993 vdd.n2510 vdd.n674 10.6151
R4994 vdd.n2511 vdd.n2510 10.6151
R4995 vdd.n2512 vdd.n2511 10.6151
R4996 vdd.n2512 vdd.n662 10.6151
R4997 vdd.n2522 vdd.n662 10.6151
R4998 vdd.n2523 vdd.n2522 10.6151
R4999 vdd.n2524 vdd.n2523 10.6151
R5000 vdd.n2524 vdd.n651 10.6151
R5001 vdd.n2534 vdd.n651 10.6151
R5002 vdd.n2535 vdd.n2534 10.6151
R5003 vdd.n2538 vdd.n2535 10.6151
R5004 vdd.n2548 vdd.n639 10.6151
R5005 vdd.n2549 vdd.n2548 10.6151
R5006 vdd.n2595 vdd.n2549 10.6151
R5007 vdd.n2595 vdd.n2594 10.6151
R5008 vdd.n2594 vdd.n2593 10.6151
R5009 vdd.n2593 vdd.n2592 10.6151
R5010 vdd.n2592 vdd.n2590 10.6151
R5011 vdd.n1987 vdd.n831 10.6151
R5012 vdd.n1997 vdd.n831 10.6151
R5013 vdd.n1998 vdd.n1997 10.6151
R5014 vdd.n1999 vdd.n1998 10.6151
R5015 vdd.n1999 vdd.n818 10.6151
R5016 vdd.n2009 vdd.n818 10.6151
R5017 vdd.n2010 vdd.n2009 10.6151
R5018 vdd.n2012 vdd.n806 10.6151
R5019 vdd.n2022 vdd.n806 10.6151
R5020 vdd.n2023 vdd.n2022 10.6151
R5021 vdd.n2024 vdd.n2023 10.6151
R5022 vdd.n2024 vdd.n794 10.6151
R5023 vdd.n2034 vdd.n794 10.6151
R5024 vdd.n2035 vdd.n2034 10.6151
R5025 vdd.n2036 vdd.n2035 10.6151
R5026 vdd.n2036 vdd.n783 10.6151
R5027 vdd.n2046 vdd.n783 10.6151
R5028 vdd.n2047 vdd.n2046 10.6151
R5029 vdd.n2048 vdd.n2047 10.6151
R5030 vdd.n2048 vdd.n771 10.6151
R5031 vdd.n2058 vdd.n771 10.6151
R5032 vdd.n2059 vdd.n2058 10.6151
R5033 vdd.n2062 vdd.n2059 10.6151
R5034 vdd.n2062 vdd.n2061 10.6151
R5035 vdd.n2061 vdd.n2060 10.6151
R5036 vdd.n2060 vdd.n754 10.6151
R5037 vdd.n2144 vdd.n754 10.6151
R5038 vdd.n2143 vdd.n2142 10.6151
R5039 vdd.n2142 vdd.n2139 10.6151
R5040 vdd.n2139 vdd.n2138 10.6151
R5041 vdd.n2138 vdd.n2135 10.6151
R5042 vdd.n2135 vdd.n2134 10.6151
R5043 vdd.n2134 vdd.n2131 10.6151
R5044 vdd.n2131 vdd.n2130 10.6151
R5045 vdd.n2130 vdd.n2127 10.6151
R5046 vdd.n2127 vdd.n2126 10.6151
R5047 vdd.n2126 vdd.n2123 10.6151
R5048 vdd.n2123 vdd.n2122 10.6151
R5049 vdd.n2122 vdd.n2119 10.6151
R5050 vdd.n2119 vdd.n2118 10.6151
R5051 vdd.n2118 vdd.n2115 10.6151
R5052 vdd.n2115 vdd.n2114 10.6151
R5053 vdd.n2114 vdd.n2111 10.6151
R5054 vdd.n2111 vdd.n2110 10.6151
R5055 vdd.n2110 vdd.n2107 10.6151
R5056 vdd.n2107 vdd.n2106 10.6151
R5057 vdd.n2106 vdd.n2103 10.6151
R5058 vdd.n2103 vdd.n2102 10.6151
R5059 vdd.n2102 vdd.n2099 10.6151
R5060 vdd.n2099 vdd.n2098 10.6151
R5061 vdd.n2098 vdd.n2095 10.6151
R5062 vdd.n2095 vdd.n2094 10.6151
R5063 vdd.n2094 vdd.n2091 10.6151
R5064 vdd.n2091 vdd.n2090 10.6151
R5065 vdd.n2090 vdd.n2087 10.6151
R5066 vdd.n2087 vdd.n2086 10.6151
R5067 vdd.n2086 vdd.n2083 10.6151
R5068 vdd.n2083 vdd.n2082 10.6151
R5069 vdd.n2079 vdd.n2078 10.6151
R5070 vdd.n2078 vdd.n2076 10.6151
R5071 vdd.n1835 vdd.n1833 10.6151
R5072 vdd.n1836 vdd.n1835 10.6151
R5073 vdd.n1838 vdd.n1836 10.6151
R5074 vdd.n1839 vdd.n1838 10.6151
R5075 vdd.n1841 vdd.n1839 10.6151
R5076 vdd.n1842 vdd.n1841 10.6151
R5077 vdd.n1844 vdd.n1842 10.6151
R5078 vdd.n1845 vdd.n1844 10.6151
R5079 vdd.n1847 vdd.n1845 10.6151
R5080 vdd.n1848 vdd.n1847 10.6151
R5081 vdd.n1850 vdd.n1848 10.6151
R5082 vdd.n1851 vdd.n1850 10.6151
R5083 vdd.n1869 vdd.n1851 10.6151
R5084 vdd.n1869 vdd.n1868 10.6151
R5085 vdd.n1868 vdd.n1867 10.6151
R5086 vdd.n1867 vdd.n1865 10.6151
R5087 vdd.n1865 vdd.n1864 10.6151
R5088 vdd.n1864 vdd.n1862 10.6151
R5089 vdd.n1862 vdd.n1861 10.6151
R5090 vdd.n1861 vdd.n1859 10.6151
R5091 vdd.n1859 vdd.n1858 10.6151
R5092 vdd.n1858 vdd.n1856 10.6151
R5093 vdd.n1856 vdd.n1855 10.6151
R5094 vdd.n1855 vdd.n1853 10.6151
R5095 vdd.n1853 vdd.n1852 10.6151
R5096 vdd.n1852 vdd.n758 10.6151
R5097 vdd.n2074 vdd.n758 10.6151
R5098 vdd.n2075 vdd.n2074 10.6151
R5099 vdd.n1986 vdd.n1985 10.6151
R5100 vdd.n1985 vdd.n843 10.6151
R5101 vdd.n1979 vdd.n843 10.6151
R5102 vdd.n1979 vdd.n1978 10.6151
R5103 vdd.n1978 vdd.n1977 10.6151
R5104 vdd.n1977 vdd.n845 10.6151
R5105 vdd.n1971 vdd.n845 10.6151
R5106 vdd.n1971 vdd.n1970 10.6151
R5107 vdd.n1970 vdd.n1969 10.6151
R5108 vdd.n1969 vdd.n847 10.6151
R5109 vdd.n1963 vdd.n847 10.6151
R5110 vdd.n1963 vdd.n1962 10.6151
R5111 vdd.n1962 vdd.n1961 10.6151
R5112 vdd.n1961 vdd.n849 10.6151
R5113 vdd.n1955 vdd.n849 10.6151
R5114 vdd.n1955 vdd.n1954 10.6151
R5115 vdd.n1954 vdd.n1953 10.6151
R5116 vdd.n1953 vdd.n853 10.6151
R5117 vdd.n1801 vdd.n853 10.6151
R5118 vdd.n1802 vdd.n1801 10.6151
R5119 vdd.n1802 vdd.n1797 10.6151
R5120 vdd.n1808 vdd.n1797 10.6151
R5121 vdd.n1809 vdd.n1808 10.6151
R5122 vdd.n1810 vdd.n1809 10.6151
R5123 vdd.n1810 vdd.n1795 10.6151
R5124 vdd.n1816 vdd.n1795 10.6151
R5125 vdd.n1817 vdd.n1816 10.6151
R5126 vdd.n1818 vdd.n1817 10.6151
R5127 vdd.n1818 vdd.n1793 10.6151
R5128 vdd.n1824 vdd.n1793 10.6151
R5129 vdd.n1825 vdd.n1824 10.6151
R5130 vdd.n1827 vdd.n1789 10.6151
R5131 vdd.n1832 vdd.n1789 10.6151
R5132 vdd.n280 vdd.n262 10.4732
R5133 vdd.n233 vdd.n215 10.4732
R5134 vdd.n190 vdd.n172 10.4732
R5135 vdd.n143 vdd.n125 10.4732
R5136 vdd.n101 vdd.n83 10.4732
R5137 vdd.n54 vdd.n36 10.4732
R5138 vdd.n1095 vdd.n1077 10.4732
R5139 vdd.n1142 vdd.n1124 10.4732
R5140 vdd.n1005 vdd.n987 10.4732
R5141 vdd.n1052 vdd.n1034 10.4732
R5142 vdd.n916 vdd.n898 10.4732
R5143 vdd.n963 vdd.n945 10.4732
R5144 vdd.t128 vdd.n888 10.3167
R5145 vdd.n2874 vdd.t148 10.3167
R5146 vdd.n1465 vdd.t124 10.09
R5147 vdd.n3042 vdd.t161 10.09
R5148 vdd.n279 vdd.n264 9.69747
R5149 vdd.n232 vdd.n217 9.69747
R5150 vdd.n189 vdd.n174 9.69747
R5151 vdd.n142 vdd.n127 9.69747
R5152 vdd.n100 vdd.n85 9.69747
R5153 vdd.n53 vdd.n38 9.69747
R5154 vdd.n1094 vdd.n1079 9.69747
R5155 vdd.n1141 vdd.n1126 9.69747
R5156 vdd.n1004 vdd.n989 9.69747
R5157 vdd.n1051 vdd.n1036 9.69747
R5158 vdd.n915 vdd.n900 9.69747
R5159 vdd.n962 vdd.n947 9.69747
R5160 vdd.n1929 vdd.n1928 9.67831
R5161 vdd.n2836 vdd.n520 9.67831
R5162 vdd.n2707 vdd.n2706 9.67831
R5163 vdd.n1953 vdd.n1952 9.67831
R5164 vdd.n295 vdd.n294 9.45567
R5165 vdd.n248 vdd.n247 9.45567
R5166 vdd.n205 vdd.n204 9.45567
R5167 vdd.n158 vdd.n157 9.45567
R5168 vdd.n116 vdd.n115 9.45567
R5169 vdd.n69 vdd.n68 9.45567
R5170 vdd.n1110 vdd.n1109 9.45567
R5171 vdd.n1157 vdd.n1156 9.45567
R5172 vdd.n1020 vdd.n1019 9.45567
R5173 vdd.n1067 vdd.n1066 9.45567
R5174 vdd.n931 vdd.n930 9.45567
R5175 vdd.n978 vdd.n977 9.45567
R5176 vdd.n1689 vdd.n1543 9.3005
R5177 vdd.n1688 vdd.n1687 9.3005
R5178 vdd.n1549 vdd.n1548 9.3005
R5179 vdd.n1682 vdd.n1553 9.3005
R5180 vdd.n1681 vdd.n1554 9.3005
R5181 vdd.n1680 vdd.n1555 9.3005
R5182 vdd.n1559 vdd.n1556 9.3005
R5183 vdd.n1675 vdd.n1560 9.3005
R5184 vdd.n1674 vdd.n1561 9.3005
R5185 vdd.n1673 vdd.n1562 9.3005
R5186 vdd.n1566 vdd.n1563 9.3005
R5187 vdd.n1668 vdd.n1567 9.3005
R5188 vdd.n1667 vdd.n1568 9.3005
R5189 vdd.n1666 vdd.n1569 9.3005
R5190 vdd.n1573 vdd.n1570 9.3005
R5191 vdd.n1661 vdd.n1574 9.3005
R5192 vdd.n1660 vdd.n1575 9.3005
R5193 vdd.n1659 vdd.n1576 9.3005
R5194 vdd.n1580 vdd.n1577 9.3005
R5195 vdd.n1654 vdd.n1581 9.3005
R5196 vdd.n1653 vdd.n1582 9.3005
R5197 vdd.n1652 vdd.n1651 9.3005
R5198 vdd.n1650 vdd.n1583 9.3005
R5199 vdd.n1649 vdd.n1648 9.3005
R5200 vdd.n1589 vdd.n1588 9.3005
R5201 vdd.n1643 vdd.n1593 9.3005
R5202 vdd.n1642 vdd.n1594 9.3005
R5203 vdd.n1641 vdd.n1595 9.3005
R5204 vdd.n1599 vdd.n1596 9.3005
R5205 vdd.n1636 vdd.n1600 9.3005
R5206 vdd.n1635 vdd.n1601 9.3005
R5207 vdd.n1634 vdd.n1602 9.3005
R5208 vdd.n1606 vdd.n1603 9.3005
R5209 vdd.n1629 vdd.n1607 9.3005
R5210 vdd.n1628 vdd.n1608 9.3005
R5211 vdd.n1627 vdd.n1609 9.3005
R5212 vdd.n1611 vdd.n1610 9.3005
R5213 vdd.n1622 vdd.n854 9.3005
R5214 vdd.n1691 vdd.n1690 9.3005
R5215 vdd.n1715 vdd.n1714 9.3005
R5216 vdd.n1521 vdd.n1520 9.3005
R5217 vdd.n1526 vdd.n1524 9.3005
R5218 vdd.n1707 vdd.n1527 9.3005
R5219 vdd.n1706 vdd.n1528 9.3005
R5220 vdd.n1705 vdd.n1529 9.3005
R5221 vdd.n1533 vdd.n1530 9.3005
R5222 vdd.n1700 vdd.n1534 9.3005
R5223 vdd.n1699 vdd.n1535 9.3005
R5224 vdd.n1698 vdd.n1536 9.3005
R5225 vdd.n1540 vdd.n1537 9.3005
R5226 vdd.n1693 vdd.n1541 9.3005
R5227 vdd.n1692 vdd.n1542 9.3005
R5228 vdd.n1937 vdd.n1514 9.3005
R5229 vdd.n1939 vdd.n1938 9.3005
R5230 vdd.n1476 vdd.n1475 9.3005
R5231 vdd.n1477 vdd.n890 9.3005
R5232 vdd.n1479 vdd.n1478 9.3005
R5233 vdd.n880 vdd.n879 9.3005
R5234 vdd.n1493 vdd.n1492 9.3005
R5235 vdd.n1494 vdd.n878 9.3005
R5236 vdd.n1496 vdd.n1495 9.3005
R5237 vdd.n868 vdd.n867 9.3005
R5238 vdd.n1512 vdd.n1511 9.3005
R5239 vdd.n1513 vdd.n866 9.3005
R5240 vdd.n1941 vdd.n1940 9.3005
R5241 vdd.n271 vdd.n270 9.3005
R5242 vdd.n266 vdd.n265 9.3005
R5243 vdd.n277 vdd.n276 9.3005
R5244 vdd.n279 vdd.n278 9.3005
R5245 vdd.n262 vdd.n261 9.3005
R5246 vdd.n285 vdd.n284 9.3005
R5247 vdd.n287 vdd.n286 9.3005
R5248 vdd.n259 vdd.n256 9.3005
R5249 vdd.n294 vdd.n293 9.3005
R5250 vdd.n224 vdd.n223 9.3005
R5251 vdd.n219 vdd.n218 9.3005
R5252 vdd.n230 vdd.n229 9.3005
R5253 vdd.n232 vdd.n231 9.3005
R5254 vdd.n215 vdd.n214 9.3005
R5255 vdd.n238 vdd.n237 9.3005
R5256 vdd.n240 vdd.n239 9.3005
R5257 vdd.n212 vdd.n209 9.3005
R5258 vdd.n247 vdd.n246 9.3005
R5259 vdd.n181 vdd.n180 9.3005
R5260 vdd.n176 vdd.n175 9.3005
R5261 vdd.n187 vdd.n186 9.3005
R5262 vdd.n189 vdd.n188 9.3005
R5263 vdd.n172 vdd.n171 9.3005
R5264 vdd.n195 vdd.n194 9.3005
R5265 vdd.n197 vdd.n196 9.3005
R5266 vdd.n169 vdd.n166 9.3005
R5267 vdd.n204 vdd.n203 9.3005
R5268 vdd.n134 vdd.n133 9.3005
R5269 vdd.n129 vdd.n128 9.3005
R5270 vdd.n140 vdd.n139 9.3005
R5271 vdd.n142 vdd.n141 9.3005
R5272 vdd.n125 vdd.n124 9.3005
R5273 vdd.n148 vdd.n147 9.3005
R5274 vdd.n150 vdd.n149 9.3005
R5275 vdd.n122 vdd.n119 9.3005
R5276 vdd.n157 vdd.n156 9.3005
R5277 vdd.n92 vdd.n91 9.3005
R5278 vdd.n87 vdd.n86 9.3005
R5279 vdd.n98 vdd.n97 9.3005
R5280 vdd.n100 vdd.n99 9.3005
R5281 vdd.n83 vdd.n82 9.3005
R5282 vdd.n106 vdd.n105 9.3005
R5283 vdd.n108 vdd.n107 9.3005
R5284 vdd.n80 vdd.n77 9.3005
R5285 vdd.n115 vdd.n114 9.3005
R5286 vdd.n45 vdd.n44 9.3005
R5287 vdd.n40 vdd.n39 9.3005
R5288 vdd.n51 vdd.n50 9.3005
R5289 vdd.n53 vdd.n52 9.3005
R5290 vdd.n36 vdd.n35 9.3005
R5291 vdd.n59 vdd.n58 9.3005
R5292 vdd.n61 vdd.n60 9.3005
R5293 vdd.n33 vdd.n30 9.3005
R5294 vdd.n68 vdd.n67 9.3005
R5295 vdd.n2758 vdd.n2757 9.3005
R5296 vdd.n2761 vdd.n555 9.3005
R5297 vdd.n2762 vdd.n554 9.3005
R5298 vdd.n2765 vdd.n553 9.3005
R5299 vdd.n2766 vdd.n552 9.3005
R5300 vdd.n2769 vdd.n551 9.3005
R5301 vdd.n2770 vdd.n550 9.3005
R5302 vdd.n2773 vdd.n549 9.3005
R5303 vdd.n2774 vdd.n548 9.3005
R5304 vdd.n2777 vdd.n547 9.3005
R5305 vdd.n2778 vdd.n546 9.3005
R5306 vdd.n2781 vdd.n545 9.3005
R5307 vdd.n2782 vdd.n544 9.3005
R5308 vdd.n2785 vdd.n543 9.3005
R5309 vdd.n2786 vdd.n542 9.3005
R5310 vdd.n2789 vdd.n541 9.3005
R5311 vdd.n2790 vdd.n540 9.3005
R5312 vdd.n2793 vdd.n539 9.3005
R5313 vdd.n2794 vdd.n538 9.3005
R5314 vdd.n2797 vdd.n537 9.3005
R5315 vdd.n2801 vdd.n2800 9.3005
R5316 vdd.n2802 vdd.n536 9.3005
R5317 vdd.n2806 vdd.n2803 9.3005
R5318 vdd.n2809 vdd.n535 9.3005
R5319 vdd.n2810 vdd.n534 9.3005
R5320 vdd.n2813 vdd.n533 9.3005
R5321 vdd.n2814 vdd.n532 9.3005
R5322 vdd.n2817 vdd.n531 9.3005
R5323 vdd.n2818 vdd.n530 9.3005
R5324 vdd.n2821 vdd.n529 9.3005
R5325 vdd.n2822 vdd.n528 9.3005
R5326 vdd.n2825 vdd.n527 9.3005
R5327 vdd.n2826 vdd.n526 9.3005
R5328 vdd.n2829 vdd.n525 9.3005
R5329 vdd.n2830 vdd.n524 9.3005
R5330 vdd.n2833 vdd.n519 9.3005
R5331 vdd.n482 vdd.n481 9.3005
R5332 vdd.n2844 vdd.n2843 9.3005
R5333 vdd.n2847 vdd.n2846 9.3005
R5334 vdd.n471 vdd.n470 9.3005
R5335 vdd.n2861 vdd.n2860 9.3005
R5336 vdd.n2862 vdd.n469 9.3005
R5337 vdd.n2864 vdd.n2863 9.3005
R5338 vdd.n460 vdd.n459 9.3005
R5339 vdd.n2877 vdd.n2876 9.3005
R5340 vdd.n2878 vdd.n458 9.3005
R5341 vdd.n2880 vdd.n2879 9.3005
R5342 vdd.n300 vdd.n298 9.3005
R5343 vdd.n2845 vdd.n480 9.3005
R5344 vdd.n3046 vdd.n3045 9.3005
R5345 vdd.n301 vdd.n299 9.3005
R5346 vdd.n3039 vdd.n310 9.3005
R5347 vdd.n3038 vdd.n311 9.3005
R5348 vdd.n3037 vdd.n312 9.3005
R5349 vdd.n320 vdd.n313 9.3005
R5350 vdd.n3031 vdd.n321 9.3005
R5351 vdd.n3030 vdd.n322 9.3005
R5352 vdd.n3029 vdd.n323 9.3005
R5353 vdd.n331 vdd.n324 9.3005
R5354 vdd.n3023 vdd.n3022 9.3005
R5355 vdd.n3019 vdd.n332 9.3005
R5356 vdd.n3018 vdd.n335 9.3005
R5357 vdd.n339 vdd.n336 9.3005
R5358 vdd.n340 vdd.n337 9.3005
R5359 vdd.n3011 vdd.n341 9.3005
R5360 vdd.n3010 vdd.n342 9.3005
R5361 vdd.n3009 vdd.n343 9.3005
R5362 vdd.n347 vdd.n344 9.3005
R5363 vdd.n3004 vdd.n348 9.3005
R5364 vdd.n3003 vdd.n349 9.3005
R5365 vdd.n3002 vdd.n350 9.3005
R5366 vdd.n354 vdd.n351 9.3005
R5367 vdd.n2997 vdd.n355 9.3005
R5368 vdd.n2996 vdd.n356 9.3005
R5369 vdd.n2995 vdd.n357 9.3005
R5370 vdd.n361 vdd.n358 9.3005
R5371 vdd.n2990 vdd.n362 9.3005
R5372 vdd.n2989 vdd.n363 9.3005
R5373 vdd.n2988 vdd.n2987 9.3005
R5374 vdd.n2986 vdd.n364 9.3005
R5375 vdd.n2985 vdd.n2984 9.3005
R5376 vdd.n370 vdd.n369 9.3005
R5377 vdd.n2979 vdd.n374 9.3005
R5378 vdd.n2978 vdd.n375 9.3005
R5379 vdd.n2977 vdd.n376 9.3005
R5380 vdd.n380 vdd.n377 9.3005
R5381 vdd.n2972 vdd.n381 9.3005
R5382 vdd.n2971 vdd.n382 9.3005
R5383 vdd.n2970 vdd.n383 9.3005
R5384 vdd.n387 vdd.n384 9.3005
R5385 vdd.n2965 vdd.n388 9.3005
R5386 vdd.n2964 vdd.n389 9.3005
R5387 vdd.n2963 vdd.n390 9.3005
R5388 vdd.n394 vdd.n391 9.3005
R5389 vdd.n2958 vdd.n395 9.3005
R5390 vdd.n2957 vdd.n396 9.3005
R5391 vdd.n2956 vdd.n397 9.3005
R5392 vdd.n401 vdd.n398 9.3005
R5393 vdd.n2951 vdd.n402 9.3005
R5394 vdd.n2950 vdd.n403 9.3005
R5395 vdd.n2949 vdd.n2948 9.3005
R5396 vdd.n2947 vdd.n404 9.3005
R5397 vdd.n2946 vdd.n2945 9.3005
R5398 vdd.n410 vdd.n409 9.3005
R5399 vdd.n2940 vdd.n414 9.3005
R5400 vdd.n2939 vdd.n415 9.3005
R5401 vdd.n2938 vdd.n416 9.3005
R5402 vdd.n420 vdd.n417 9.3005
R5403 vdd.n2933 vdd.n421 9.3005
R5404 vdd.n2932 vdd.n422 9.3005
R5405 vdd.n2931 vdd.n423 9.3005
R5406 vdd.n427 vdd.n424 9.3005
R5407 vdd.n2926 vdd.n428 9.3005
R5408 vdd.n2925 vdd.n429 9.3005
R5409 vdd.n2924 vdd.n430 9.3005
R5410 vdd.n434 vdd.n431 9.3005
R5411 vdd.n2919 vdd.n435 9.3005
R5412 vdd.n2918 vdd.n436 9.3005
R5413 vdd.n2917 vdd.n437 9.3005
R5414 vdd.n441 vdd.n438 9.3005
R5415 vdd.n2912 vdd.n442 9.3005
R5416 vdd.n2911 vdd.n443 9.3005
R5417 vdd.n2907 vdd.n2904 9.3005
R5418 vdd.n3021 vdd.n3020 9.3005
R5419 vdd.n2852 vdd.n2851 9.3005
R5420 vdd.n2853 vdd.n475 9.3005
R5421 vdd.n2855 vdd.n2854 9.3005
R5422 vdd.n465 vdd.n464 9.3005
R5423 vdd.n2869 vdd.n2868 9.3005
R5424 vdd.n2870 vdd.n463 9.3005
R5425 vdd.n2872 vdd.n2871 9.3005
R5426 vdd.n453 vdd.n452 9.3005
R5427 vdd.n2885 vdd.n2884 9.3005
R5428 vdd.n2886 vdd.n451 9.3005
R5429 vdd.n2888 vdd.n2887 9.3005
R5430 vdd.n2889 vdd.n450 9.3005
R5431 vdd.n2891 vdd.n2890 9.3005
R5432 vdd.n2892 vdd.n449 9.3005
R5433 vdd.n2894 vdd.n2893 9.3005
R5434 vdd.n2895 vdd.n447 9.3005
R5435 vdd.n2897 vdd.n2896 9.3005
R5436 vdd.n2898 vdd.n446 9.3005
R5437 vdd.n2900 vdd.n2899 9.3005
R5438 vdd.n2901 vdd.n444 9.3005
R5439 vdd.n2903 vdd.n2902 9.3005
R5440 vdd.n477 vdd.n476 9.3005
R5441 vdd.n2710 vdd.n2709 9.3005
R5442 vdd.n2715 vdd.n2708 9.3005
R5443 vdd.n2724 vdd.n572 9.3005
R5444 vdd.n2727 vdd.n571 9.3005
R5445 vdd.n2728 vdd.n570 9.3005
R5446 vdd.n2731 vdd.n569 9.3005
R5447 vdd.n2732 vdd.n568 9.3005
R5448 vdd.n2735 vdd.n567 9.3005
R5449 vdd.n2736 vdd.n566 9.3005
R5450 vdd.n2739 vdd.n565 9.3005
R5451 vdd.n2740 vdd.n564 9.3005
R5452 vdd.n2743 vdd.n563 9.3005
R5453 vdd.n2744 vdd.n562 9.3005
R5454 vdd.n2747 vdd.n561 9.3005
R5455 vdd.n2748 vdd.n560 9.3005
R5456 vdd.n2751 vdd.n559 9.3005
R5457 vdd.n2755 vdd.n2754 9.3005
R5458 vdd.n2756 vdd.n556 9.3005
R5459 vdd.n1951 vdd.n1950 9.3005
R5460 vdd.n1946 vdd.n857 9.3005
R5461 vdd.n1433 vdd.n1432 9.3005
R5462 vdd.n1434 vdd.n1188 9.3005
R5463 vdd.n1436 vdd.n1435 9.3005
R5464 vdd.n1178 vdd.n1177 9.3005
R5465 vdd.n1450 vdd.n1449 9.3005
R5466 vdd.n1451 vdd.n1176 9.3005
R5467 vdd.n1453 vdd.n1452 9.3005
R5468 vdd.n1168 vdd.n1167 9.3005
R5469 vdd.n1468 vdd.n1467 9.3005
R5470 vdd.n1469 vdd.n1166 9.3005
R5471 vdd.n1471 vdd.n1470 9.3005
R5472 vdd.n885 vdd.n884 9.3005
R5473 vdd.n1484 vdd.n1483 9.3005
R5474 vdd.n1485 vdd.n883 9.3005
R5475 vdd.n1487 vdd.n1486 9.3005
R5476 vdd.n875 vdd.n874 9.3005
R5477 vdd.n1501 vdd.n1500 9.3005
R5478 vdd.n1502 vdd.n872 9.3005
R5479 vdd.n1506 vdd.n1505 9.3005
R5480 vdd.n1504 vdd.n873 9.3005
R5481 vdd.n1503 vdd.n862 9.3005
R5482 vdd.n1190 vdd.n1189 9.3005
R5483 vdd.n1326 vdd.n1325 9.3005
R5484 vdd.n1327 vdd.n1316 9.3005
R5485 vdd.n1329 vdd.n1328 9.3005
R5486 vdd.n1330 vdd.n1315 9.3005
R5487 vdd.n1332 vdd.n1331 9.3005
R5488 vdd.n1333 vdd.n1310 9.3005
R5489 vdd.n1335 vdd.n1334 9.3005
R5490 vdd.n1336 vdd.n1309 9.3005
R5491 vdd.n1338 vdd.n1337 9.3005
R5492 vdd.n1339 vdd.n1304 9.3005
R5493 vdd.n1341 vdd.n1340 9.3005
R5494 vdd.n1342 vdd.n1303 9.3005
R5495 vdd.n1344 vdd.n1343 9.3005
R5496 vdd.n1345 vdd.n1298 9.3005
R5497 vdd.n1347 vdd.n1346 9.3005
R5498 vdd.n1348 vdd.n1297 9.3005
R5499 vdd.n1350 vdd.n1349 9.3005
R5500 vdd.n1351 vdd.n1292 9.3005
R5501 vdd.n1353 vdd.n1352 9.3005
R5502 vdd.n1354 vdd.n1291 9.3005
R5503 vdd.n1356 vdd.n1355 9.3005
R5504 vdd.n1360 vdd.n1287 9.3005
R5505 vdd.n1362 vdd.n1361 9.3005
R5506 vdd.n1363 vdd.n1286 9.3005
R5507 vdd.n1365 vdd.n1364 9.3005
R5508 vdd.n1366 vdd.n1281 9.3005
R5509 vdd.n1368 vdd.n1367 9.3005
R5510 vdd.n1369 vdd.n1280 9.3005
R5511 vdd.n1371 vdd.n1370 9.3005
R5512 vdd.n1372 vdd.n1275 9.3005
R5513 vdd.n1374 vdd.n1373 9.3005
R5514 vdd.n1375 vdd.n1274 9.3005
R5515 vdd.n1377 vdd.n1376 9.3005
R5516 vdd.n1378 vdd.n1269 9.3005
R5517 vdd.n1380 vdd.n1379 9.3005
R5518 vdd.n1381 vdd.n1268 9.3005
R5519 vdd.n1383 vdd.n1382 9.3005
R5520 vdd.n1384 vdd.n1263 9.3005
R5521 vdd.n1386 vdd.n1385 9.3005
R5522 vdd.n1387 vdd.n1262 9.3005
R5523 vdd.n1389 vdd.n1388 9.3005
R5524 vdd.n1390 vdd.n1257 9.3005
R5525 vdd.n1392 vdd.n1391 9.3005
R5526 vdd.n1393 vdd.n1256 9.3005
R5527 vdd.n1395 vdd.n1394 9.3005
R5528 vdd.n1396 vdd.n1249 9.3005
R5529 vdd.n1398 vdd.n1397 9.3005
R5530 vdd.n1399 vdd.n1248 9.3005
R5531 vdd.n1401 vdd.n1400 9.3005
R5532 vdd.n1402 vdd.n1243 9.3005
R5533 vdd.n1404 vdd.n1403 9.3005
R5534 vdd.n1405 vdd.n1242 9.3005
R5535 vdd.n1407 vdd.n1406 9.3005
R5536 vdd.n1408 vdd.n1237 9.3005
R5537 vdd.n1410 vdd.n1409 9.3005
R5538 vdd.n1411 vdd.n1236 9.3005
R5539 vdd.n1413 vdd.n1412 9.3005
R5540 vdd.n1414 vdd.n1231 9.3005
R5541 vdd.n1416 vdd.n1415 9.3005
R5542 vdd.n1417 vdd.n1230 9.3005
R5543 vdd.n1419 vdd.n1418 9.3005
R5544 vdd.n1195 vdd.n1194 9.3005
R5545 vdd.n1425 vdd.n1424 9.3005
R5546 vdd.n1324 vdd.n1323 9.3005
R5547 vdd.n1428 vdd.n1427 9.3005
R5548 vdd.n1184 vdd.n1183 9.3005
R5549 vdd.n1442 vdd.n1441 9.3005
R5550 vdd.n1443 vdd.n1182 9.3005
R5551 vdd.n1445 vdd.n1444 9.3005
R5552 vdd.n1173 vdd.n1172 9.3005
R5553 vdd.n1459 vdd.n1458 9.3005
R5554 vdd.n1460 vdd.n1171 9.3005
R5555 vdd.n1463 vdd.n1462 9.3005
R5556 vdd.n1461 vdd.n1162 9.3005
R5557 vdd.n1426 vdd.n1193 9.3005
R5558 vdd.n1086 vdd.n1085 9.3005
R5559 vdd.n1081 vdd.n1080 9.3005
R5560 vdd.n1092 vdd.n1091 9.3005
R5561 vdd.n1094 vdd.n1093 9.3005
R5562 vdd.n1077 vdd.n1076 9.3005
R5563 vdd.n1100 vdd.n1099 9.3005
R5564 vdd.n1102 vdd.n1101 9.3005
R5565 vdd.n1074 vdd.n1071 9.3005
R5566 vdd.n1109 vdd.n1108 9.3005
R5567 vdd.n1133 vdd.n1132 9.3005
R5568 vdd.n1128 vdd.n1127 9.3005
R5569 vdd.n1139 vdd.n1138 9.3005
R5570 vdd.n1141 vdd.n1140 9.3005
R5571 vdd.n1124 vdd.n1123 9.3005
R5572 vdd.n1147 vdd.n1146 9.3005
R5573 vdd.n1149 vdd.n1148 9.3005
R5574 vdd.n1121 vdd.n1118 9.3005
R5575 vdd.n1156 vdd.n1155 9.3005
R5576 vdd.n996 vdd.n995 9.3005
R5577 vdd.n991 vdd.n990 9.3005
R5578 vdd.n1002 vdd.n1001 9.3005
R5579 vdd.n1004 vdd.n1003 9.3005
R5580 vdd.n987 vdd.n986 9.3005
R5581 vdd.n1010 vdd.n1009 9.3005
R5582 vdd.n1012 vdd.n1011 9.3005
R5583 vdd.n984 vdd.n981 9.3005
R5584 vdd.n1019 vdd.n1018 9.3005
R5585 vdd.n1043 vdd.n1042 9.3005
R5586 vdd.n1038 vdd.n1037 9.3005
R5587 vdd.n1049 vdd.n1048 9.3005
R5588 vdd.n1051 vdd.n1050 9.3005
R5589 vdd.n1034 vdd.n1033 9.3005
R5590 vdd.n1057 vdd.n1056 9.3005
R5591 vdd.n1059 vdd.n1058 9.3005
R5592 vdd.n1031 vdd.n1028 9.3005
R5593 vdd.n1066 vdd.n1065 9.3005
R5594 vdd.n907 vdd.n906 9.3005
R5595 vdd.n902 vdd.n901 9.3005
R5596 vdd.n913 vdd.n912 9.3005
R5597 vdd.n915 vdd.n914 9.3005
R5598 vdd.n898 vdd.n897 9.3005
R5599 vdd.n921 vdd.n920 9.3005
R5600 vdd.n923 vdd.n922 9.3005
R5601 vdd.n895 vdd.n892 9.3005
R5602 vdd.n930 vdd.n929 9.3005
R5603 vdd.n954 vdd.n953 9.3005
R5604 vdd.n949 vdd.n948 9.3005
R5605 vdd.n960 vdd.n959 9.3005
R5606 vdd.n962 vdd.n961 9.3005
R5607 vdd.n945 vdd.n944 9.3005
R5608 vdd.n968 vdd.n967 9.3005
R5609 vdd.n970 vdd.n969 9.3005
R5610 vdd.n942 vdd.n939 9.3005
R5611 vdd.n977 vdd.n976 9.3005
R5612 vdd.n1438 vdd.t157 8.95635
R5613 vdd.t139 vdd.n3033 8.95635
R5614 vdd.n276 vdd.n275 8.92171
R5615 vdd.n229 vdd.n228 8.92171
R5616 vdd.n186 vdd.n185 8.92171
R5617 vdd.n139 vdd.n138 8.92171
R5618 vdd.n97 vdd.n96 8.92171
R5619 vdd.n50 vdd.n49 8.92171
R5620 vdd.n1091 vdd.n1090 8.92171
R5621 vdd.n1138 vdd.n1137 8.92171
R5622 vdd.n1001 vdd.n1000 8.92171
R5623 vdd.n1048 vdd.n1047 8.92171
R5624 vdd.n912 vdd.n911 8.92171
R5625 vdd.n959 vdd.n958 8.92171
R5626 vdd.n207 vdd.n117 8.81535
R5627 vdd.n1069 vdd.n979 8.81535
R5628 vdd.n1465 vdd.t135 8.72962
R5629 vdd.t137 vdd.n3042 8.72962
R5630 vdd.n888 vdd.t173 8.50289
R5631 vdd.n1943 vdd.t40 8.50289
R5632 vdd.n516 vdd.t33 8.50289
R5633 vdd.n2874 vdd.t151 8.50289
R5634 vdd.n28 vdd.n14 8.42249
R5635 vdd.n3048 vdd.n3047 8.16225
R5636 vdd.n1161 vdd.n1160 8.16225
R5637 vdd.n272 vdd.n266 8.14595
R5638 vdd.n225 vdd.n219 8.14595
R5639 vdd.n182 vdd.n176 8.14595
R5640 vdd.n135 vdd.n129 8.14595
R5641 vdd.n93 vdd.n87 8.14595
R5642 vdd.n46 vdd.n40 8.14595
R5643 vdd.n1087 vdd.n1081 8.14595
R5644 vdd.n1134 vdd.n1128 8.14595
R5645 vdd.n997 vdd.n991 8.14595
R5646 vdd.n1044 vdd.n1038 8.14595
R5647 vdd.n908 vdd.n902 8.14595
R5648 vdd.n955 vdd.n949 8.14595
R5649 vdd.n2537 vdd.n639 8.11757
R5650 vdd.n2011 vdd.n2010 8.11757
R5651 vdd.n1989 vdd.n833 7.70933
R5652 vdd.n1995 vdd.n833 7.70933
R5653 vdd.n2001 vdd.n827 7.70933
R5654 vdd.n2001 vdd.n820 7.70933
R5655 vdd.n2007 vdd.n820 7.70933
R5656 vdd.n2007 vdd.n823 7.70933
R5657 vdd.n2014 vdd.n808 7.70933
R5658 vdd.n2020 vdd.n808 7.70933
R5659 vdd.n2026 vdd.n802 7.70933
R5660 vdd.n2032 vdd.n798 7.70933
R5661 vdd.n2038 vdd.n792 7.70933
R5662 vdd.n2050 vdd.n779 7.70933
R5663 vdd.n2056 vdd.n773 7.70933
R5664 vdd.n2056 vdd.n766 7.70933
R5665 vdd.n2064 vdd.n766 7.70933
R5666 vdd.n2071 vdd.t184 7.70933
R5667 vdd.n2146 vdd.t184 7.70933
R5668 vdd.n2478 vdd.t186 7.70933
R5669 vdd.n2484 vdd.t186 7.70933
R5670 vdd.n2490 vdd.n687 7.70933
R5671 vdd.n2496 vdd.n687 7.70933
R5672 vdd.n2496 vdd.n690 7.70933
R5673 vdd.n2502 vdd.n683 7.70933
R5674 vdd.n2514 vdd.n670 7.70933
R5675 vdd.n2520 vdd.n664 7.70933
R5676 vdd.n2526 vdd.n660 7.70933
R5677 vdd.n2532 vdd.n647 7.70933
R5678 vdd.n2540 vdd.n647 7.70933
R5679 vdd.n2546 vdd.n641 7.70933
R5680 vdd.n2546 vdd.n633 7.70933
R5681 vdd.n2597 vdd.n633 7.70933
R5682 vdd.n2597 vdd.n636 7.70933
R5683 vdd.n2603 vdd.n595 7.70933
R5684 vdd.n2673 vdd.n595 7.70933
R5685 vdd.n271 vdd.n268 7.3702
R5686 vdd.n224 vdd.n221 7.3702
R5687 vdd.n181 vdd.n178 7.3702
R5688 vdd.n134 vdd.n131 7.3702
R5689 vdd.n92 vdd.n89 7.3702
R5690 vdd.n45 vdd.n42 7.3702
R5691 vdd.n1086 vdd.n1083 7.3702
R5692 vdd.n1133 vdd.n1130 7.3702
R5693 vdd.n996 vdd.n993 7.3702
R5694 vdd.n1043 vdd.n1040 7.3702
R5695 vdd.n907 vdd.n904 7.3702
R5696 vdd.n954 vdd.n951 7.3702
R5697 vdd.n1361 vdd.n1360 6.98232
R5698 vdd.n1653 vdd.n1652 6.98232
R5699 vdd.n2950 vdd.n2949 6.98232
R5700 vdd.n2761 vdd.n2758 6.98232
R5701 vdd.n1498 vdd.t120 6.68904
R5702 vdd.n2857 vdd.t122 6.68904
R5703 vdd.t159 vdd.n887 6.46231
R5704 vdd.n2882 vdd.t126 6.46231
R5705 vdd.n1456 vdd.t141 6.23558
R5706 vdd.t130 vdd.n308 6.23558
R5707 vdd.n3048 vdd.n297 6.22547
R5708 vdd.n1160 vdd.n1159 6.22547
R5709 vdd.n2026 vdd.t0 6.00885
R5710 vdd.n2526 vdd.t26 6.00885
R5711 vdd.n823 vdd.t84 5.89549
R5712 vdd.t48 vdd.n641 5.89549
R5713 vdd.n272 vdd.n271 5.81868
R5714 vdd.n225 vdd.n224 5.81868
R5715 vdd.n182 vdd.n181 5.81868
R5716 vdd.n135 vdd.n134 5.81868
R5717 vdd.n93 vdd.n92 5.81868
R5718 vdd.n46 vdd.n45 5.81868
R5719 vdd.n1087 vdd.n1086 5.81868
R5720 vdd.n1134 vdd.n1133 5.81868
R5721 vdd.n997 vdd.n996 5.81868
R5722 vdd.n1044 vdd.n1043 5.81868
R5723 vdd.n908 vdd.n907 5.81868
R5724 vdd.n955 vdd.n954 5.81868
R5725 vdd.t80 vdd.n827 5.78212
R5726 vdd.n1770 vdd.t65 5.78212
R5727 vdd.n2395 vdd.t73 5.78212
R5728 vdd.n636 vdd.t69 5.78212
R5729 vdd.n2154 vdd.n2153 5.77611
R5730 vdd.n1897 vdd.n1767 5.77611
R5731 vdd.n2408 vdd.n2407 5.77611
R5732 vdd.n2614 vdd.n2613 5.77611
R5733 vdd.n2678 vdd.n591 5.77611
R5734 vdd.n2318 vdd.n2258 5.77611
R5735 vdd.n2079 vdd.n757 5.77611
R5736 vdd.n1827 vdd.n1826 5.77611
R5737 vdd.n1323 vdd.n1322 5.62474
R5738 vdd.n1949 vdd.n1946 5.62474
R5739 vdd.n2910 vdd.n2907 5.62474
R5740 vdd.n2713 vdd.n2710 5.62474
R5741 vdd.t27 vdd.n779 5.44203
R5742 vdd.n683 vdd.t116 5.44203
R5743 vdd.n1180 vdd.t141 5.10193
R5744 vdd.t110 vdd.n802 5.10193
R5745 vdd.n792 vdd.t25 5.10193
R5746 vdd.t1 vdd.n670 5.10193
R5747 vdd.n660 vdd.t2 5.10193
R5748 vdd.n3035 vdd.t130 5.10193
R5749 vdd.n275 vdd.n266 5.04292
R5750 vdd.n228 vdd.n219 5.04292
R5751 vdd.n185 vdd.n176 5.04292
R5752 vdd.n138 vdd.n129 5.04292
R5753 vdd.n96 vdd.n87 5.04292
R5754 vdd.n49 vdd.n40 5.04292
R5755 vdd.n1090 vdd.n1081 5.04292
R5756 vdd.n1137 vdd.n1128 5.04292
R5757 vdd.n1000 vdd.n991 5.04292
R5758 vdd.n1047 vdd.n1038 5.04292
R5759 vdd.n911 vdd.n902 5.04292
R5760 vdd.n958 vdd.n949 5.04292
R5761 vdd.n1473 vdd.t159 4.8752
R5762 vdd.t31 vdd.t194 4.8752
R5763 vdd.t111 vdd.t112 4.8752
R5764 vdd.t192 vdd.t21 4.8752
R5765 vdd.t29 vdd.t108 4.8752
R5766 vdd.t126 vdd.n304 4.8752
R5767 vdd.n2155 vdd.n2154 4.83952
R5768 vdd.n1767 vdd.n1763 4.83952
R5769 vdd.n2409 vdd.n2408 4.83952
R5770 vdd.n2615 vdd.n2614 4.83952
R5771 vdd.n591 vdd.n586 4.83952
R5772 vdd.n2315 vdd.n2258 4.83952
R5773 vdd.n2082 vdd.n757 4.83952
R5774 vdd.n1826 vdd.n1825 4.83952
R5775 vdd.n1621 vdd.n855 4.74817
R5776 vdd.n1616 vdd.n856 4.74817
R5777 vdd.n1518 vdd.n1515 4.74817
R5778 vdd.n1930 vdd.n1519 4.74817
R5779 vdd.n1932 vdd.n1518 4.74817
R5780 vdd.n1931 vdd.n1930 4.74817
R5781 vdd.n2838 vdd.n2837 4.74817
R5782 vdd.n2835 vdd.n2834 4.74817
R5783 vdd.n2835 vdd.n521 4.74817
R5784 vdd.n2837 vdd.n518 4.74817
R5785 vdd.n2720 vdd.n573 4.74817
R5786 vdd.n2716 vdd.n574 4.74817
R5787 vdd.n2719 vdd.n574 4.74817
R5788 vdd.n2723 vdd.n573 4.74817
R5789 vdd.n1617 vdd.n855 4.74817
R5790 vdd.n858 vdd.n856 4.74817
R5791 vdd.n297 vdd.n296 4.7074
R5792 vdd.n207 vdd.n206 4.7074
R5793 vdd.n1159 vdd.n1158 4.7074
R5794 vdd.n1069 vdd.n1068 4.7074
R5795 vdd.n1489 vdd.t120 4.64847
R5796 vdd.n2866 vdd.t122 4.64847
R5797 vdd.n2032 vdd.t190 4.53511
R5798 vdd.n2520 vdd.t198 4.53511
R5799 vdd.n2064 vdd.t196 4.30838
R5800 vdd.n2490 vdd.t19 4.30838
R5801 vdd.n276 vdd.n264 4.26717
R5802 vdd.n229 vdd.n217 4.26717
R5803 vdd.n186 vdd.n174 4.26717
R5804 vdd.n139 vdd.n127 4.26717
R5805 vdd.n97 vdd.n85 4.26717
R5806 vdd.n50 vdd.n38 4.26717
R5807 vdd.n1091 vdd.n1079 4.26717
R5808 vdd.n1138 vdd.n1126 4.26717
R5809 vdd.n1001 vdd.n989 4.26717
R5810 vdd.n1048 vdd.n1036 4.26717
R5811 vdd.n912 vdd.n900 4.26717
R5812 vdd.n959 vdd.n947 4.26717
R5813 vdd.n297 vdd.n207 4.10845
R5814 vdd.n1159 vdd.n1069 4.10845
R5815 vdd.n253 vdd.t167 4.06363
R5816 vdd.n253 vdd.t131 4.06363
R5817 vdd.n251 vdd.t133 4.06363
R5818 vdd.n251 vdd.t154 4.06363
R5819 vdd.n249 vdd.t156 4.06363
R5820 vdd.n249 vdd.t172 4.06363
R5821 vdd.n163 vdd.t162 4.06363
R5822 vdd.n163 vdd.t183 4.06363
R5823 vdd.n161 vdd.t127 4.06363
R5824 vdd.n161 vdd.t146 4.06363
R5825 vdd.n159 vdd.t152 4.06363
R5826 vdd.n159 vdd.t163 4.06363
R5827 vdd.n74 vdd.t168 4.06363
R5828 vdd.n74 vdd.t143 4.06363
R5829 vdd.n72 vdd.t182 4.06363
R5830 vdd.n72 vdd.t138 4.06363
R5831 vdd.n70 vdd.t175 4.06363
R5832 vdd.n70 vdd.t149 4.06363
R5833 vdd.n1111 vdd.t134 4.06363
R5834 vdd.n1111 vdd.t178 4.06363
R5835 vdd.n1113 vdd.t177 4.06363
R5836 vdd.n1113 vdd.t166 4.06363
R5837 vdd.n1115 vdd.t153 4.06363
R5838 vdd.n1115 vdd.t132 4.06363
R5839 vdd.n1021 vdd.t129 4.06363
R5840 vdd.n1021 vdd.t174 4.06363
R5841 vdd.n1023 vdd.t169 4.06363
R5842 vdd.n1023 vdd.t160 4.06363
R5843 vdd.n1025 vdd.t145 4.06363
R5844 vdd.n1025 vdd.t125 4.06363
R5845 vdd.n932 vdd.t147 4.06363
R5846 vdd.n932 vdd.t176 4.06363
R5847 vdd.n934 vdd.t136 4.06363
R5848 vdd.n934 vdd.t164 4.06363
R5849 vdd.n936 vdd.t142 4.06363
R5850 vdd.n936 vdd.t170 4.06363
R5851 vdd.n26 vdd.t12 3.9605
R5852 vdd.n26 vdd.t9 3.9605
R5853 vdd.n23 vdd.t16 3.9605
R5854 vdd.n23 vdd.t15 3.9605
R5855 vdd.n21 vdd.t8 3.9605
R5856 vdd.n21 vdd.t5 3.9605
R5857 vdd.n20 vdd.t10 3.9605
R5858 vdd.n20 vdd.t11 3.9605
R5859 vdd.n15 vdd.t14 3.9605
R5860 vdd.n15 vdd.t18 3.9605
R5861 vdd.n16 vdd.t6 3.9605
R5862 vdd.n16 vdd.t17 3.9605
R5863 vdd.n18 vdd.t7 3.9605
R5864 vdd.n18 vdd.t13 3.9605
R5865 vdd.n25 vdd.t3 3.9605
R5866 vdd.n25 vdd.t4 3.9605
R5867 vdd.n7 vdd.t30 3.61217
R5868 vdd.n7 vdd.t199 3.61217
R5869 vdd.n8 vdd.t193 3.61217
R5870 vdd.n8 vdd.t117 3.61217
R5871 vdd.n10 vdd.t187 3.61217
R5872 vdd.n10 vdd.t20 3.61217
R5873 vdd.n12 vdd.t23 3.61217
R5874 vdd.n12 vdd.t189 3.61217
R5875 vdd.n5 vdd.t115 3.61217
R5876 vdd.n5 vdd.t119 3.61217
R5877 vdd.n3 vdd.t197 3.61217
R5878 vdd.n3 vdd.t185 3.61217
R5879 vdd.n1 vdd.t28 3.61217
R5880 vdd.n1 vdd.t113 3.61217
R5881 vdd.n0 vdd.t191 3.61217
R5882 vdd.n0 vdd.t195 3.61217
R5883 vdd.n280 vdd.n279 3.49141
R5884 vdd.n233 vdd.n232 3.49141
R5885 vdd.n190 vdd.n189 3.49141
R5886 vdd.n143 vdd.n142 3.49141
R5887 vdd.n101 vdd.n100 3.49141
R5888 vdd.n54 vdd.n53 3.49141
R5889 vdd.n1095 vdd.n1094 3.49141
R5890 vdd.n1142 vdd.n1141 3.49141
R5891 vdd.n1005 vdd.n1004 3.49141
R5892 vdd.n1052 vdd.n1051 3.49141
R5893 vdd.n916 vdd.n915 3.49141
R5894 vdd.n963 vdd.n962 3.49141
R5895 vdd.n1770 vdd.t196 3.40145
R5896 vdd.n2218 vdd.t114 3.40145
R5897 vdd.n2471 vdd.t188 3.40145
R5898 vdd.n2395 vdd.t19 3.40145
R5899 vdd.n1871 vdd.t190 3.17472
R5900 vdd.n2374 vdd.t198 3.17472
R5901 vdd.n1490 vdd.t173 2.83463
R5902 vdd.n1508 vdd.t40 2.83463
R5903 vdd.n2849 vdd.t33 2.83463
R5904 vdd.n467 vdd.t151 2.83463
R5905 vdd.n283 vdd.n262 2.71565
R5906 vdd.n236 vdd.n215 2.71565
R5907 vdd.n193 vdd.n172 2.71565
R5908 vdd.n146 vdd.n125 2.71565
R5909 vdd.n104 vdd.n83 2.71565
R5910 vdd.n57 vdd.n36 2.71565
R5911 vdd.n1098 vdd.n1077 2.71565
R5912 vdd.n1145 vdd.n1124 2.71565
R5913 vdd.n1008 vdd.n987 2.71565
R5914 vdd.n1055 vdd.n1034 2.71565
R5915 vdd.n919 vdd.n898 2.71565
R5916 vdd.n966 vdd.n945 2.71565
R5917 vdd.t135 vdd.n1164 2.6079
R5918 vdd.n2020 vdd.t110 2.6079
R5919 vdd.n2044 vdd.t25 2.6079
R5920 vdd.n2508 vdd.t1 2.6079
R5921 vdd.n2532 vdd.t2 2.6079
R5922 vdd.n3043 vdd.t137 2.6079
R5923 vdd.n2538 vdd.n2537 2.49806
R5924 vdd.n2012 vdd.n2011 2.49806
R5925 vdd.n270 vdd.n269 2.4129
R5926 vdd.n223 vdd.n222 2.4129
R5927 vdd.n180 vdd.n179 2.4129
R5928 vdd.n133 vdd.n132 2.4129
R5929 vdd.n91 vdd.n90 2.4129
R5930 vdd.n44 vdd.n43 2.4129
R5931 vdd.n1085 vdd.n1084 2.4129
R5932 vdd.n1132 vdd.n1131 2.4129
R5933 vdd.n995 vdd.n994 2.4129
R5934 vdd.n1042 vdd.n1041 2.4129
R5935 vdd.n906 vdd.n905 2.4129
R5936 vdd.n953 vdd.n952 2.4129
R5937 vdd.n1447 vdd.t157 2.38117
R5938 vdd.n3034 vdd.t139 2.38117
R5939 vdd.n1929 vdd.n1518 2.27742
R5940 vdd.n1930 vdd.n1929 2.27742
R5941 vdd.n2836 vdd.n2835 2.27742
R5942 vdd.n2837 vdd.n2836 2.27742
R5943 vdd.n2707 vdd.n574 2.27742
R5944 vdd.n2707 vdd.n573 2.27742
R5945 vdd.n1952 vdd.n855 2.27742
R5946 vdd.n1952 vdd.n856 2.27742
R5947 vdd.n2044 vdd.t27 2.2678
R5948 vdd.n2508 vdd.t116 2.2678
R5949 vdd.t112 vdd.n773 2.04107
R5950 vdd.n690 vdd.t192 2.04107
R5951 vdd.n284 vdd.n260 1.93989
R5952 vdd.n237 vdd.n213 1.93989
R5953 vdd.n194 vdd.n170 1.93989
R5954 vdd.n147 vdd.n123 1.93989
R5955 vdd.n105 vdd.n81 1.93989
R5956 vdd.n58 vdd.n34 1.93989
R5957 vdd.n1099 vdd.n1075 1.93989
R5958 vdd.n1146 vdd.n1122 1.93989
R5959 vdd.n1009 vdd.n985 1.93989
R5960 vdd.n1056 vdd.n1032 1.93989
R5961 vdd.n920 vdd.n896 1.93989
R5962 vdd.n967 vdd.n943 1.93989
R5963 vdd.n1995 vdd.t80 1.92771
R5964 vdd.n2071 vdd.t65 1.92771
R5965 vdd.n2484 vdd.t73 1.92771
R5966 vdd.n2603 vdd.t69 1.92771
R5967 vdd.n1871 vdd.t0 1.70098
R5968 vdd.n798 vdd.t31 1.70098
R5969 vdd.t108 vdd.n664 1.70098
R5970 vdd.n2374 vdd.t26 1.70098
R5971 vdd.n1455 vdd.t124 1.24752
R5972 vdd.t161 vdd.n3041 1.24752
R5973 vdd.n295 vdd.n255 1.16414
R5974 vdd.n288 vdd.n287 1.16414
R5975 vdd.n248 vdd.n208 1.16414
R5976 vdd.n241 vdd.n240 1.16414
R5977 vdd.n205 vdd.n165 1.16414
R5978 vdd.n198 vdd.n197 1.16414
R5979 vdd.n158 vdd.n118 1.16414
R5980 vdd.n151 vdd.n150 1.16414
R5981 vdd.n116 vdd.n76 1.16414
R5982 vdd.n109 vdd.n108 1.16414
R5983 vdd.n69 vdd.n29 1.16414
R5984 vdd.n62 vdd.n61 1.16414
R5985 vdd.n1110 vdd.n1070 1.16414
R5986 vdd.n1103 vdd.n1102 1.16414
R5987 vdd.n1157 vdd.n1117 1.16414
R5988 vdd.n1150 vdd.n1149 1.16414
R5989 vdd.n1020 vdd.n980 1.16414
R5990 vdd.n1013 vdd.n1012 1.16414
R5991 vdd.n1067 vdd.n1027 1.16414
R5992 vdd.n1060 vdd.n1059 1.16414
R5993 vdd.n931 vdd.n891 1.16414
R5994 vdd.n924 vdd.n923 1.16414
R5995 vdd.n978 vdd.n938 1.16414
R5996 vdd.n971 vdd.n970 1.16414
R5997 vdd.n2038 vdd.t194 1.13415
R5998 vdd.n2514 vdd.t29 1.13415
R5999 vdd.n1481 vdd.t128 1.02079
R6000 vdd.t84 vdd.t109 1.02079
R6001 vdd.t24 vdd.t48 1.02079
R6002 vdd.t148 vdd.n456 1.02079
R6003 vdd.n1326 vdd.n1322 0.970197
R6004 vdd.n1950 vdd.n1949 0.970197
R6005 vdd.n2911 vdd.n2910 0.970197
R6006 vdd.n2715 vdd.n2713 0.970197
R6007 vdd.n2014 vdd.t109 0.794056
R6008 vdd.n2050 vdd.t111 0.794056
R6009 vdd.n2502 vdd.t21 0.794056
R6010 vdd.n2540 vdd.t24 0.794056
R6011 vdd.n1160 vdd.n28 0.74827
R6012 vdd vdd.n3048 0.740437
R6013 vdd.n1430 vdd.t44 0.567326
R6014 vdd.n3026 vdd.t55 0.567326
R6015 vdd.n1940 vdd.n1939 0.537085
R6016 vdd.n2845 vdd.n2844 0.537085
R6017 vdd.n3022 vdd.n3021 0.537085
R6018 vdd.n2904 vdd.n2903 0.537085
R6019 vdd.n2709 vdd.n476 0.537085
R6020 vdd.n1503 vdd.n857 0.537085
R6021 vdd.n1324 vdd.n1189 0.537085
R6022 vdd.n1426 vdd.n1425 0.537085
R6023 vdd.n4 vdd.n2 0.459552
R6024 vdd.n11 vdd.n9 0.459552
R6025 vdd.n293 vdd.n292 0.388379
R6026 vdd.n259 vdd.n257 0.388379
R6027 vdd.n246 vdd.n245 0.388379
R6028 vdd.n212 vdd.n210 0.388379
R6029 vdd.n203 vdd.n202 0.388379
R6030 vdd.n169 vdd.n167 0.388379
R6031 vdd.n156 vdd.n155 0.388379
R6032 vdd.n122 vdd.n120 0.388379
R6033 vdd.n114 vdd.n113 0.388379
R6034 vdd.n80 vdd.n78 0.388379
R6035 vdd.n67 vdd.n66 0.388379
R6036 vdd.n33 vdd.n31 0.388379
R6037 vdd.n1108 vdd.n1107 0.388379
R6038 vdd.n1074 vdd.n1072 0.388379
R6039 vdd.n1155 vdd.n1154 0.388379
R6040 vdd.n1121 vdd.n1119 0.388379
R6041 vdd.n1018 vdd.n1017 0.388379
R6042 vdd.n984 vdd.n982 0.388379
R6043 vdd.n1065 vdd.n1064 0.388379
R6044 vdd.n1031 vdd.n1029 0.388379
R6045 vdd.n929 vdd.n928 0.388379
R6046 vdd.n895 vdd.n893 0.388379
R6047 vdd.n976 vdd.n975 0.388379
R6048 vdd.n942 vdd.n940 0.388379
R6049 vdd.n19 vdd.n17 0.387128
R6050 vdd.n24 vdd.n22 0.387128
R6051 vdd.n6 vdd.n4 0.358259
R6052 vdd.n13 vdd.n11 0.358259
R6053 vdd.n252 vdd.n250 0.358259
R6054 vdd.n254 vdd.n252 0.358259
R6055 vdd.n296 vdd.n254 0.358259
R6056 vdd.n162 vdd.n160 0.358259
R6057 vdd.n164 vdd.n162 0.358259
R6058 vdd.n206 vdd.n164 0.358259
R6059 vdd.n73 vdd.n71 0.358259
R6060 vdd.n75 vdd.n73 0.358259
R6061 vdd.n117 vdd.n75 0.358259
R6062 vdd.n1158 vdd.n1116 0.358259
R6063 vdd.n1116 vdd.n1114 0.358259
R6064 vdd.n1114 vdd.n1112 0.358259
R6065 vdd.n1068 vdd.n1026 0.358259
R6066 vdd.n1026 vdd.n1024 0.358259
R6067 vdd.n1024 vdd.n1022 0.358259
R6068 vdd.n979 vdd.n937 0.358259
R6069 vdd.n937 vdd.n935 0.358259
R6070 vdd.n935 vdd.n933 0.358259
R6071 vdd.n14 vdd.n6 0.334552
R6072 vdd.n14 vdd.n13 0.334552
R6073 vdd.n27 vdd.n19 0.21707
R6074 vdd.n27 vdd.n24 0.21707
R6075 vdd.n294 vdd.n256 0.155672
R6076 vdd.n286 vdd.n256 0.155672
R6077 vdd.n286 vdd.n285 0.155672
R6078 vdd.n285 vdd.n261 0.155672
R6079 vdd.n278 vdd.n261 0.155672
R6080 vdd.n278 vdd.n277 0.155672
R6081 vdd.n277 vdd.n265 0.155672
R6082 vdd.n270 vdd.n265 0.155672
R6083 vdd.n247 vdd.n209 0.155672
R6084 vdd.n239 vdd.n209 0.155672
R6085 vdd.n239 vdd.n238 0.155672
R6086 vdd.n238 vdd.n214 0.155672
R6087 vdd.n231 vdd.n214 0.155672
R6088 vdd.n231 vdd.n230 0.155672
R6089 vdd.n230 vdd.n218 0.155672
R6090 vdd.n223 vdd.n218 0.155672
R6091 vdd.n204 vdd.n166 0.155672
R6092 vdd.n196 vdd.n166 0.155672
R6093 vdd.n196 vdd.n195 0.155672
R6094 vdd.n195 vdd.n171 0.155672
R6095 vdd.n188 vdd.n171 0.155672
R6096 vdd.n188 vdd.n187 0.155672
R6097 vdd.n187 vdd.n175 0.155672
R6098 vdd.n180 vdd.n175 0.155672
R6099 vdd.n157 vdd.n119 0.155672
R6100 vdd.n149 vdd.n119 0.155672
R6101 vdd.n149 vdd.n148 0.155672
R6102 vdd.n148 vdd.n124 0.155672
R6103 vdd.n141 vdd.n124 0.155672
R6104 vdd.n141 vdd.n140 0.155672
R6105 vdd.n140 vdd.n128 0.155672
R6106 vdd.n133 vdd.n128 0.155672
R6107 vdd.n115 vdd.n77 0.155672
R6108 vdd.n107 vdd.n77 0.155672
R6109 vdd.n107 vdd.n106 0.155672
R6110 vdd.n106 vdd.n82 0.155672
R6111 vdd.n99 vdd.n82 0.155672
R6112 vdd.n99 vdd.n98 0.155672
R6113 vdd.n98 vdd.n86 0.155672
R6114 vdd.n91 vdd.n86 0.155672
R6115 vdd.n68 vdd.n30 0.155672
R6116 vdd.n60 vdd.n30 0.155672
R6117 vdd.n60 vdd.n59 0.155672
R6118 vdd.n59 vdd.n35 0.155672
R6119 vdd.n52 vdd.n35 0.155672
R6120 vdd.n52 vdd.n51 0.155672
R6121 vdd.n51 vdd.n39 0.155672
R6122 vdd.n44 vdd.n39 0.155672
R6123 vdd.n1109 vdd.n1071 0.155672
R6124 vdd.n1101 vdd.n1071 0.155672
R6125 vdd.n1101 vdd.n1100 0.155672
R6126 vdd.n1100 vdd.n1076 0.155672
R6127 vdd.n1093 vdd.n1076 0.155672
R6128 vdd.n1093 vdd.n1092 0.155672
R6129 vdd.n1092 vdd.n1080 0.155672
R6130 vdd.n1085 vdd.n1080 0.155672
R6131 vdd.n1156 vdd.n1118 0.155672
R6132 vdd.n1148 vdd.n1118 0.155672
R6133 vdd.n1148 vdd.n1147 0.155672
R6134 vdd.n1147 vdd.n1123 0.155672
R6135 vdd.n1140 vdd.n1123 0.155672
R6136 vdd.n1140 vdd.n1139 0.155672
R6137 vdd.n1139 vdd.n1127 0.155672
R6138 vdd.n1132 vdd.n1127 0.155672
R6139 vdd.n1019 vdd.n981 0.155672
R6140 vdd.n1011 vdd.n981 0.155672
R6141 vdd.n1011 vdd.n1010 0.155672
R6142 vdd.n1010 vdd.n986 0.155672
R6143 vdd.n1003 vdd.n986 0.155672
R6144 vdd.n1003 vdd.n1002 0.155672
R6145 vdd.n1002 vdd.n990 0.155672
R6146 vdd.n995 vdd.n990 0.155672
R6147 vdd.n1066 vdd.n1028 0.155672
R6148 vdd.n1058 vdd.n1028 0.155672
R6149 vdd.n1058 vdd.n1057 0.155672
R6150 vdd.n1057 vdd.n1033 0.155672
R6151 vdd.n1050 vdd.n1033 0.155672
R6152 vdd.n1050 vdd.n1049 0.155672
R6153 vdd.n1049 vdd.n1037 0.155672
R6154 vdd.n1042 vdd.n1037 0.155672
R6155 vdd.n930 vdd.n892 0.155672
R6156 vdd.n922 vdd.n892 0.155672
R6157 vdd.n922 vdd.n921 0.155672
R6158 vdd.n921 vdd.n897 0.155672
R6159 vdd.n914 vdd.n897 0.155672
R6160 vdd.n914 vdd.n913 0.155672
R6161 vdd.n913 vdd.n901 0.155672
R6162 vdd.n906 vdd.n901 0.155672
R6163 vdd.n977 vdd.n939 0.155672
R6164 vdd.n969 vdd.n939 0.155672
R6165 vdd.n969 vdd.n968 0.155672
R6166 vdd.n968 vdd.n944 0.155672
R6167 vdd.n961 vdd.n944 0.155672
R6168 vdd.n961 vdd.n960 0.155672
R6169 vdd.n960 vdd.n948 0.155672
R6170 vdd.n953 vdd.n948 0.155672
R6171 vdd.n1715 vdd.n1520 0.152939
R6172 vdd.n1526 vdd.n1520 0.152939
R6173 vdd.n1527 vdd.n1526 0.152939
R6174 vdd.n1528 vdd.n1527 0.152939
R6175 vdd.n1529 vdd.n1528 0.152939
R6176 vdd.n1533 vdd.n1529 0.152939
R6177 vdd.n1534 vdd.n1533 0.152939
R6178 vdd.n1535 vdd.n1534 0.152939
R6179 vdd.n1536 vdd.n1535 0.152939
R6180 vdd.n1540 vdd.n1536 0.152939
R6181 vdd.n1541 vdd.n1540 0.152939
R6182 vdd.n1542 vdd.n1541 0.152939
R6183 vdd.n1690 vdd.n1542 0.152939
R6184 vdd.n1690 vdd.n1689 0.152939
R6185 vdd.n1689 vdd.n1688 0.152939
R6186 vdd.n1688 vdd.n1548 0.152939
R6187 vdd.n1553 vdd.n1548 0.152939
R6188 vdd.n1554 vdd.n1553 0.152939
R6189 vdd.n1555 vdd.n1554 0.152939
R6190 vdd.n1559 vdd.n1555 0.152939
R6191 vdd.n1560 vdd.n1559 0.152939
R6192 vdd.n1561 vdd.n1560 0.152939
R6193 vdd.n1562 vdd.n1561 0.152939
R6194 vdd.n1566 vdd.n1562 0.152939
R6195 vdd.n1567 vdd.n1566 0.152939
R6196 vdd.n1568 vdd.n1567 0.152939
R6197 vdd.n1569 vdd.n1568 0.152939
R6198 vdd.n1573 vdd.n1569 0.152939
R6199 vdd.n1574 vdd.n1573 0.152939
R6200 vdd.n1575 vdd.n1574 0.152939
R6201 vdd.n1576 vdd.n1575 0.152939
R6202 vdd.n1580 vdd.n1576 0.152939
R6203 vdd.n1581 vdd.n1580 0.152939
R6204 vdd.n1582 vdd.n1581 0.152939
R6205 vdd.n1651 vdd.n1582 0.152939
R6206 vdd.n1651 vdd.n1650 0.152939
R6207 vdd.n1650 vdd.n1649 0.152939
R6208 vdd.n1649 vdd.n1588 0.152939
R6209 vdd.n1593 vdd.n1588 0.152939
R6210 vdd.n1594 vdd.n1593 0.152939
R6211 vdd.n1595 vdd.n1594 0.152939
R6212 vdd.n1599 vdd.n1595 0.152939
R6213 vdd.n1600 vdd.n1599 0.152939
R6214 vdd.n1601 vdd.n1600 0.152939
R6215 vdd.n1602 vdd.n1601 0.152939
R6216 vdd.n1606 vdd.n1602 0.152939
R6217 vdd.n1607 vdd.n1606 0.152939
R6218 vdd.n1608 vdd.n1607 0.152939
R6219 vdd.n1609 vdd.n1608 0.152939
R6220 vdd.n1610 vdd.n1609 0.152939
R6221 vdd.n1610 vdd.n854 0.152939
R6222 vdd.n1939 vdd.n1514 0.152939
R6223 vdd.n1477 vdd.n1476 0.152939
R6224 vdd.n1478 vdd.n1477 0.152939
R6225 vdd.n1478 vdd.n879 0.152939
R6226 vdd.n1493 vdd.n879 0.152939
R6227 vdd.n1494 vdd.n1493 0.152939
R6228 vdd.n1495 vdd.n1494 0.152939
R6229 vdd.n1495 vdd.n867 0.152939
R6230 vdd.n1512 vdd.n867 0.152939
R6231 vdd.n1513 vdd.n1512 0.152939
R6232 vdd.n1940 vdd.n1513 0.152939
R6233 vdd.n524 vdd.n519 0.152939
R6234 vdd.n525 vdd.n524 0.152939
R6235 vdd.n526 vdd.n525 0.152939
R6236 vdd.n527 vdd.n526 0.152939
R6237 vdd.n528 vdd.n527 0.152939
R6238 vdd.n529 vdd.n528 0.152939
R6239 vdd.n530 vdd.n529 0.152939
R6240 vdd.n531 vdd.n530 0.152939
R6241 vdd.n532 vdd.n531 0.152939
R6242 vdd.n533 vdd.n532 0.152939
R6243 vdd.n534 vdd.n533 0.152939
R6244 vdd.n535 vdd.n534 0.152939
R6245 vdd.n2803 vdd.n535 0.152939
R6246 vdd.n2803 vdd.n2802 0.152939
R6247 vdd.n2802 vdd.n2801 0.152939
R6248 vdd.n2801 vdd.n537 0.152939
R6249 vdd.n538 vdd.n537 0.152939
R6250 vdd.n539 vdd.n538 0.152939
R6251 vdd.n540 vdd.n539 0.152939
R6252 vdd.n541 vdd.n540 0.152939
R6253 vdd.n542 vdd.n541 0.152939
R6254 vdd.n543 vdd.n542 0.152939
R6255 vdd.n544 vdd.n543 0.152939
R6256 vdd.n545 vdd.n544 0.152939
R6257 vdd.n546 vdd.n545 0.152939
R6258 vdd.n547 vdd.n546 0.152939
R6259 vdd.n548 vdd.n547 0.152939
R6260 vdd.n549 vdd.n548 0.152939
R6261 vdd.n550 vdd.n549 0.152939
R6262 vdd.n551 vdd.n550 0.152939
R6263 vdd.n552 vdd.n551 0.152939
R6264 vdd.n553 vdd.n552 0.152939
R6265 vdd.n554 vdd.n553 0.152939
R6266 vdd.n555 vdd.n554 0.152939
R6267 vdd.n2757 vdd.n555 0.152939
R6268 vdd.n2757 vdd.n2756 0.152939
R6269 vdd.n2756 vdd.n2755 0.152939
R6270 vdd.n2755 vdd.n559 0.152939
R6271 vdd.n560 vdd.n559 0.152939
R6272 vdd.n561 vdd.n560 0.152939
R6273 vdd.n562 vdd.n561 0.152939
R6274 vdd.n563 vdd.n562 0.152939
R6275 vdd.n564 vdd.n563 0.152939
R6276 vdd.n565 vdd.n564 0.152939
R6277 vdd.n566 vdd.n565 0.152939
R6278 vdd.n567 vdd.n566 0.152939
R6279 vdd.n568 vdd.n567 0.152939
R6280 vdd.n569 vdd.n568 0.152939
R6281 vdd.n570 vdd.n569 0.152939
R6282 vdd.n571 vdd.n570 0.152939
R6283 vdd.n572 vdd.n571 0.152939
R6284 vdd.n2844 vdd.n481 0.152939
R6285 vdd.n2846 vdd.n2845 0.152939
R6286 vdd.n2846 vdd.n470 0.152939
R6287 vdd.n2861 vdd.n470 0.152939
R6288 vdd.n2862 vdd.n2861 0.152939
R6289 vdd.n2863 vdd.n2862 0.152939
R6290 vdd.n2863 vdd.n459 0.152939
R6291 vdd.n2877 vdd.n459 0.152939
R6292 vdd.n2878 vdd.n2877 0.152939
R6293 vdd.n2879 vdd.n2878 0.152939
R6294 vdd.n2879 vdd.n298 0.152939
R6295 vdd.n3046 vdd.n299 0.152939
R6296 vdd.n310 vdd.n299 0.152939
R6297 vdd.n311 vdd.n310 0.152939
R6298 vdd.n312 vdd.n311 0.152939
R6299 vdd.n320 vdd.n312 0.152939
R6300 vdd.n321 vdd.n320 0.152939
R6301 vdd.n322 vdd.n321 0.152939
R6302 vdd.n323 vdd.n322 0.152939
R6303 vdd.n331 vdd.n323 0.152939
R6304 vdd.n3022 vdd.n331 0.152939
R6305 vdd.n3021 vdd.n332 0.152939
R6306 vdd.n335 vdd.n332 0.152939
R6307 vdd.n339 vdd.n335 0.152939
R6308 vdd.n340 vdd.n339 0.152939
R6309 vdd.n341 vdd.n340 0.152939
R6310 vdd.n342 vdd.n341 0.152939
R6311 vdd.n343 vdd.n342 0.152939
R6312 vdd.n347 vdd.n343 0.152939
R6313 vdd.n348 vdd.n347 0.152939
R6314 vdd.n349 vdd.n348 0.152939
R6315 vdd.n350 vdd.n349 0.152939
R6316 vdd.n354 vdd.n350 0.152939
R6317 vdd.n355 vdd.n354 0.152939
R6318 vdd.n356 vdd.n355 0.152939
R6319 vdd.n357 vdd.n356 0.152939
R6320 vdd.n361 vdd.n357 0.152939
R6321 vdd.n362 vdd.n361 0.152939
R6322 vdd.n363 vdd.n362 0.152939
R6323 vdd.n2987 vdd.n363 0.152939
R6324 vdd.n2987 vdd.n2986 0.152939
R6325 vdd.n2986 vdd.n2985 0.152939
R6326 vdd.n2985 vdd.n369 0.152939
R6327 vdd.n374 vdd.n369 0.152939
R6328 vdd.n375 vdd.n374 0.152939
R6329 vdd.n376 vdd.n375 0.152939
R6330 vdd.n380 vdd.n376 0.152939
R6331 vdd.n381 vdd.n380 0.152939
R6332 vdd.n382 vdd.n381 0.152939
R6333 vdd.n383 vdd.n382 0.152939
R6334 vdd.n387 vdd.n383 0.152939
R6335 vdd.n388 vdd.n387 0.152939
R6336 vdd.n389 vdd.n388 0.152939
R6337 vdd.n390 vdd.n389 0.152939
R6338 vdd.n394 vdd.n390 0.152939
R6339 vdd.n395 vdd.n394 0.152939
R6340 vdd.n396 vdd.n395 0.152939
R6341 vdd.n397 vdd.n396 0.152939
R6342 vdd.n401 vdd.n397 0.152939
R6343 vdd.n402 vdd.n401 0.152939
R6344 vdd.n403 vdd.n402 0.152939
R6345 vdd.n2948 vdd.n403 0.152939
R6346 vdd.n2948 vdd.n2947 0.152939
R6347 vdd.n2947 vdd.n2946 0.152939
R6348 vdd.n2946 vdd.n409 0.152939
R6349 vdd.n414 vdd.n409 0.152939
R6350 vdd.n415 vdd.n414 0.152939
R6351 vdd.n416 vdd.n415 0.152939
R6352 vdd.n420 vdd.n416 0.152939
R6353 vdd.n421 vdd.n420 0.152939
R6354 vdd.n422 vdd.n421 0.152939
R6355 vdd.n423 vdd.n422 0.152939
R6356 vdd.n427 vdd.n423 0.152939
R6357 vdd.n428 vdd.n427 0.152939
R6358 vdd.n429 vdd.n428 0.152939
R6359 vdd.n430 vdd.n429 0.152939
R6360 vdd.n434 vdd.n430 0.152939
R6361 vdd.n435 vdd.n434 0.152939
R6362 vdd.n436 vdd.n435 0.152939
R6363 vdd.n437 vdd.n436 0.152939
R6364 vdd.n441 vdd.n437 0.152939
R6365 vdd.n442 vdd.n441 0.152939
R6366 vdd.n443 vdd.n442 0.152939
R6367 vdd.n2904 vdd.n443 0.152939
R6368 vdd.n2852 vdd.n476 0.152939
R6369 vdd.n2853 vdd.n2852 0.152939
R6370 vdd.n2854 vdd.n2853 0.152939
R6371 vdd.n2854 vdd.n464 0.152939
R6372 vdd.n2869 vdd.n464 0.152939
R6373 vdd.n2870 vdd.n2869 0.152939
R6374 vdd.n2871 vdd.n2870 0.152939
R6375 vdd.n2871 vdd.n452 0.152939
R6376 vdd.n2885 vdd.n452 0.152939
R6377 vdd.n2886 vdd.n2885 0.152939
R6378 vdd.n2887 vdd.n2886 0.152939
R6379 vdd.n2887 vdd.n450 0.152939
R6380 vdd.n2891 vdd.n450 0.152939
R6381 vdd.n2892 vdd.n2891 0.152939
R6382 vdd.n2893 vdd.n2892 0.152939
R6383 vdd.n2893 vdd.n447 0.152939
R6384 vdd.n2897 vdd.n447 0.152939
R6385 vdd.n2898 vdd.n2897 0.152939
R6386 vdd.n2899 vdd.n2898 0.152939
R6387 vdd.n2899 vdd.n444 0.152939
R6388 vdd.n2903 vdd.n444 0.152939
R6389 vdd.n2709 vdd.n2708 0.152939
R6390 vdd.n1951 vdd.n857 0.152939
R6391 vdd.n1433 vdd.n1189 0.152939
R6392 vdd.n1434 vdd.n1433 0.152939
R6393 vdd.n1435 vdd.n1434 0.152939
R6394 vdd.n1435 vdd.n1177 0.152939
R6395 vdd.n1450 vdd.n1177 0.152939
R6396 vdd.n1451 vdd.n1450 0.152939
R6397 vdd.n1452 vdd.n1451 0.152939
R6398 vdd.n1452 vdd.n1167 0.152939
R6399 vdd.n1468 vdd.n1167 0.152939
R6400 vdd.n1469 vdd.n1468 0.152939
R6401 vdd.n1470 vdd.n1469 0.152939
R6402 vdd.n1470 vdd.n884 0.152939
R6403 vdd.n1484 vdd.n884 0.152939
R6404 vdd.n1485 vdd.n1484 0.152939
R6405 vdd.n1486 vdd.n1485 0.152939
R6406 vdd.n1486 vdd.n874 0.152939
R6407 vdd.n1501 vdd.n874 0.152939
R6408 vdd.n1502 vdd.n1501 0.152939
R6409 vdd.n1505 vdd.n1502 0.152939
R6410 vdd.n1505 vdd.n1504 0.152939
R6411 vdd.n1504 vdd.n1503 0.152939
R6412 vdd.n1425 vdd.n1194 0.152939
R6413 vdd.n1418 vdd.n1194 0.152939
R6414 vdd.n1418 vdd.n1417 0.152939
R6415 vdd.n1417 vdd.n1416 0.152939
R6416 vdd.n1416 vdd.n1231 0.152939
R6417 vdd.n1412 vdd.n1231 0.152939
R6418 vdd.n1412 vdd.n1411 0.152939
R6419 vdd.n1411 vdd.n1410 0.152939
R6420 vdd.n1410 vdd.n1237 0.152939
R6421 vdd.n1406 vdd.n1237 0.152939
R6422 vdd.n1406 vdd.n1405 0.152939
R6423 vdd.n1405 vdd.n1404 0.152939
R6424 vdd.n1404 vdd.n1243 0.152939
R6425 vdd.n1400 vdd.n1243 0.152939
R6426 vdd.n1400 vdd.n1399 0.152939
R6427 vdd.n1399 vdd.n1398 0.152939
R6428 vdd.n1398 vdd.n1249 0.152939
R6429 vdd.n1394 vdd.n1249 0.152939
R6430 vdd.n1394 vdd.n1393 0.152939
R6431 vdd.n1393 vdd.n1392 0.152939
R6432 vdd.n1392 vdd.n1257 0.152939
R6433 vdd.n1388 vdd.n1257 0.152939
R6434 vdd.n1388 vdd.n1387 0.152939
R6435 vdd.n1387 vdd.n1386 0.152939
R6436 vdd.n1386 vdd.n1263 0.152939
R6437 vdd.n1382 vdd.n1263 0.152939
R6438 vdd.n1382 vdd.n1381 0.152939
R6439 vdd.n1381 vdd.n1380 0.152939
R6440 vdd.n1380 vdd.n1269 0.152939
R6441 vdd.n1376 vdd.n1269 0.152939
R6442 vdd.n1376 vdd.n1375 0.152939
R6443 vdd.n1375 vdd.n1374 0.152939
R6444 vdd.n1374 vdd.n1275 0.152939
R6445 vdd.n1370 vdd.n1275 0.152939
R6446 vdd.n1370 vdd.n1369 0.152939
R6447 vdd.n1369 vdd.n1368 0.152939
R6448 vdd.n1368 vdd.n1281 0.152939
R6449 vdd.n1364 vdd.n1281 0.152939
R6450 vdd.n1364 vdd.n1363 0.152939
R6451 vdd.n1363 vdd.n1362 0.152939
R6452 vdd.n1362 vdd.n1287 0.152939
R6453 vdd.n1355 vdd.n1287 0.152939
R6454 vdd.n1355 vdd.n1354 0.152939
R6455 vdd.n1354 vdd.n1353 0.152939
R6456 vdd.n1353 vdd.n1292 0.152939
R6457 vdd.n1349 vdd.n1292 0.152939
R6458 vdd.n1349 vdd.n1348 0.152939
R6459 vdd.n1348 vdd.n1347 0.152939
R6460 vdd.n1347 vdd.n1298 0.152939
R6461 vdd.n1343 vdd.n1298 0.152939
R6462 vdd.n1343 vdd.n1342 0.152939
R6463 vdd.n1342 vdd.n1341 0.152939
R6464 vdd.n1341 vdd.n1304 0.152939
R6465 vdd.n1337 vdd.n1304 0.152939
R6466 vdd.n1337 vdd.n1336 0.152939
R6467 vdd.n1336 vdd.n1335 0.152939
R6468 vdd.n1335 vdd.n1310 0.152939
R6469 vdd.n1331 vdd.n1310 0.152939
R6470 vdd.n1331 vdd.n1330 0.152939
R6471 vdd.n1330 vdd.n1329 0.152939
R6472 vdd.n1329 vdd.n1316 0.152939
R6473 vdd.n1325 vdd.n1316 0.152939
R6474 vdd.n1325 vdd.n1324 0.152939
R6475 vdd.n1427 vdd.n1426 0.152939
R6476 vdd.n1427 vdd.n1183 0.152939
R6477 vdd.n1442 vdd.n1183 0.152939
R6478 vdd.n1443 vdd.n1442 0.152939
R6479 vdd.n1444 vdd.n1443 0.152939
R6480 vdd.n1444 vdd.n1172 0.152939
R6481 vdd.n1459 vdd.n1172 0.152939
R6482 vdd.n1460 vdd.n1459 0.152939
R6483 vdd.n1462 vdd.n1460 0.152939
R6484 vdd.n1462 vdd.n1461 0.152939
R6485 vdd.n1929 vdd.n1514 0.110256
R6486 vdd.n2836 vdd.n481 0.110256
R6487 vdd.n2708 vdd.n2707 0.110256
R6488 vdd.n1952 vdd.n1951 0.110256
R6489 vdd.n1476 vdd.n1161 0.0695946
R6490 vdd.n3047 vdd.n298 0.0695946
R6491 vdd.n3047 vdd.n3046 0.0695946
R6492 vdd.n1461 vdd.n1161 0.0695946
R6493 vdd.n1929 vdd.n1715 0.0431829
R6494 vdd.n1952 vdd.n854 0.0431829
R6495 vdd.n2836 vdd.n519 0.0431829
R6496 vdd.n2707 vdd.n572 0.0431829
R6497 vdd vdd.n28 0.00833333
R6498 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R6499 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R6500 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R6501 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R6502 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R6503 a_n2848_n452.n1 a_n2848_n452.t40 533.058
R6504 a_n2848_n452.n101 a_n2848_n452.t24 512.366
R6505 a_n2848_n452.n100 a_n2848_n452.t26 512.366
R6506 a_n2848_n452.n69 a_n2848_n452.t36 512.366
R6507 a_n2848_n452.n98 a_n2848_n452.t44 512.366
R6508 a_n2848_n452.n19 a_n2848_n452.t38 539.01
R6509 a_n2848_n452.n78 a_n2848_n452.t28 512.366
R6510 a_n2848_n452.n79 a_n2848_n452.t32 512.366
R6511 a_n2848_n452.n73 a_n2848_n452.t46 512.366
R6512 a_n2848_n452.n80 a_n2848_n452.t34 512.366
R6513 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R6514 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R6515 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R6516 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R6517 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R6518 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R6519 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R6520 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R6521 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R6522 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R6523 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R6524 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R6525 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R6526 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R6527 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R6528 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R6529 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R6530 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R6531 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R6532 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R6533 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R6534 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R6535 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R6536 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R6537 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R6538 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R6539 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R6540 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R6541 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R6542 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R6543 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R6544 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R6545 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R6546 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R6547 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R6548 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R6549 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R6550 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R6551 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R6552 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R6553 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R6554 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R6555 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R6556 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R6557 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R6558 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R6559 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R6560 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R6561 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R6562 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R6563 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R6564 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R6565 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R6566 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R6567 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R6568 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R6569 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R6570 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R6571 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R6572 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R6573 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R6574 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R6575 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R6576 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R6577 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R6578 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R6579 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R6580 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R6581 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R6582 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R6583 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R6584 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R6585 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R6586 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R6587 a_n2848_n452.n27 a_n2848_n452.t31 74.6477
R6588 a_n2848_n452.n24 a_n2848_n452.t39 74.6477
R6589 a_n2848_n452.n26 a_n2848_n452.t41 74.2899
R6590 a_n2848_n452.n25 a_n2848_n452.t43 74.2897
R6591 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R6592 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R6593 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R6594 a_n2848_n452.n104 a_n2848_n452.n27 70.6782
R6595 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R6596 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R6597 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R6598 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R6599 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R6600 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R6601 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R6602 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R6603 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R6604 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R6605 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R6606 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R6607 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R6608 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R6609 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R6610 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R6611 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R6612 a_n2848_n452.n47 a_n2848_n452.t30 533.058
R6613 a_n2848_n452.t42 a_n2848_n452.n37 533.058
R6614 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R6615 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R6616 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R6617 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R6618 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R6619 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R6620 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R6621 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R6622 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R6623 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R6624 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R6625 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R6626 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R6627 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R6628 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R6629 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R6630 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R6631 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R6632 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R6633 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R6634 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R6635 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R6636 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R6637 a_n2848_n452.n103 a_n2848_n452.t37 3.61217
R6638 a_n2848_n452.n103 a_n2848_n452.t45 3.61217
R6639 a_n2848_n452.n72 a_n2848_n452.t47 3.61217
R6640 a_n2848_n452.n72 a_n2848_n452.t35 3.61217
R6641 a_n2848_n452.n71 a_n2848_n452.t29 3.61217
R6642 a_n2848_n452.n71 a_n2848_n452.t33 3.61217
R6643 a_n2848_n452.t25 a_n2848_n452.n104 3.61217
R6644 a_n2848_n452.n104 a_n2848_n452.t27 3.61217
R6645 a_n2848_n452.n65 a_n2848_n452.t0 2.82907
R6646 a_n2848_n452.n65 a_n2848_n452.t21 2.82907
R6647 a_n2848_n452.n66 a_n2848_n452.t8 2.82907
R6648 a_n2848_n452.n66 a_n2848_n452.t9 2.82907
R6649 a_n2848_n452.n68 a_n2848_n452.t3 2.82907
R6650 a_n2848_n452.n68 a_n2848_n452.t4 2.82907
R6651 a_n2848_n452.n64 a_n2848_n452.t23 2.82907
R6652 a_n2848_n452.n64 a_n2848_n452.t19 2.82907
R6653 a_n2848_n452.n62 a_n2848_n452.t16 2.82907
R6654 a_n2848_n452.n62 a_n2848_n452.t13 2.82907
R6655 a_n2848_n452.n60 a_n2848_n452.t2 2.82907
R6656 a_n2848_n452.n60 a_n2848_n452.t15 2.82907
R6657 a_n2848_n452.n56 a_n2848_n452.t11 2.82907
R6658 a_n2848_n452.n56 a_n2848_n452.t6 2.82907
R6659 a_n2848_n452.n57 a_n2848_n452.t7 2.82907
R6660 a_n2848_n452.n57 a_n2848_n452.t12 2.82907
R6661 a_n2848_n452.n59 a_n2848_n452.t17 2.82907
R6662 a_n2848_n452.n59 a_n2848_n452.t14 2.82907
R6663 a_n2848_n452.n55 a_n2848_n452.t20 2.82907
R6664 a_n2848_n452.n55 a_n2848_n452.t22 2.82907
R6665 a_n2848_n452.n53 a_n2848_n452.t1 2.82907
R6666 a_n2848_n452.n53 a_n2848_n452.t5 2.82907
R6667 a_n2848_n452.n52 a_n2848_n452.t18 2.82907
R6668 a_n2848_n452.n52 a_n2848_n452.t10 2.82907
R6669 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R6670 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R6671 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R6672 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R6673 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R6674 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R6675 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R6676 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R6677 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R6678 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R6679 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R6680 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R6681 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R6682 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R6683 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R6684 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R6685 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R6686 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R6687 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R6688 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R6689 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R6690 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R6691 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R6692 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R6693 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R6694 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R6695 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R6696 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R6697 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R6698 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R6699 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R6700 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R6701 a_n1986_8322.n6 a_n1986_8322.t6 74.6477
R6702 a_n1986_8322.n1 a_n1986_8322.t13 74.6477
R6703 a_n1986_8322.t22 a_n1986_8322.n18 74.6476
R6704 a_n1986_8322.n14 a_n1986_8322.t15 74.2899
R6705 a_n1986_8322.n7 a_n1986_8322.t4 74.2899
R6706 a_n1986_8322.n8 a_n1986_8322.t7 74.2899
R6707 a_n1986_8322.n11 a_n1986_8322.t8 74.2899
R6708 a_n1986_8322.n4 a_n1986_8322.t12 74.2899
R6709 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R6710 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R6711 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R6712 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R6713 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R6714 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R6715 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R6716 a_n1986_8322.n13 a_n1986_8322.t0 10.2757
R6717 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R6718 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R6719 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R6720 a_n1986_8322.n17 a_n1986_8322.t20 3.61217
R6721 a_n1986_8322.n17 a_n1986_8322.t17 3.61217
R6722 a_n1986_8322.n15 a_n1986_8322.t14 3.61217
R6723 a_n1986_8322.n15 a_n1986_8322.t23 3.61217
R6724 a_n1986_8322.n5 a_n1986_8322.t10 3.61217
R6725 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R6726 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R6727 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R6728 a_n1986_8322.n0 a_n1986_8322.t21 3.61217
R6729 a_n1986_8322.n0 a_n1986_8322.t16 3.61217
R6730 a_n1986_8322.n2 a_n1986_8322.t19 3.61217
R6731 a_n1986_8322.n2 a_n1986_8322.t18 3.61217
R6732 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R6733 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R6734 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R6735 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R6736 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R6737 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R6738 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R6739 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R6740 a_n1986_8322.t3 a_n1986_8322.t2 0.0788333
R6741 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R6742 a_n1986_8322.t0 a_n1986_8322.t1 0.0471944
R6743 a_n1986_8322.t0 a_n1986_8322.t2 0.0453889
R6744 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R6745 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R6746 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R6747 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R6748 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R6749 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R6750 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R6751 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R6752 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R6753 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R6754 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R6755 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R6756 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R6757 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R6758 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R6759 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R6760 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R6761 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R6762 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R6763 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R6764 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R6765 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R6766 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R6767 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R6768 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R6769 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R6770 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R6771 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R6772 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R6773 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R6774 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R6775 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R6776 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R6777 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R6778 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R6779 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R6780 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R6781 plus.n76 plus.t11 250.337
R6782 plus.n15 plus.t14 250.337
R6783 plus.n124 plus.t2 243.97
R6784 plus.n120 plus.t24 231.093
R6785 plus.n59 plus.t20 231.093
R6786 plus.n124 plus.n123 223.454
R6787 plus.n126 plus.n125 223.454
R6788 plus.n77 plus.t5 187.445
R6789 plus.n74 plus.t22 187.445
R6790 plus.n72 plus.t21 187.445
R6791 plus.n89 plus.t16 187.445
R6792 plus.n95 plus.t17 187.445
R6793 plus.n68 plus.t13 187.445
R6794 plus.n66 plus.t15 187.445
R6795 plus.n107 plus.t10 187.445
R6796 plus.n113 plus.t26 187.445
R6797 plus.n62 plus.t28 187.445
R6798 plus.n1 plus.t23 187.445
R6799 plus.n52 plus.t6 187.445
R6800 plus.n46 plus.t12 187.445
R6801 plus.n5 plus.t8 187.445
R6802 plus.n7 plus.t7 187.445
R6803 plus.n34 plus.t19 187.445
R6804 plus.n28 plus.t18 187.445
R6805 plus.n11 plus.t27 187.445
R6806 plus.n13 plus.t25 187.445
R6807 plus.n16 plus.t9 187.445
R6808 plus.n121 plus.n120 161.3
R6809 plus.n119 plus.n61 161.3
R6810 plus.n118 plus.n117 161.3
R6811 plus.n116 plus.n115 161.3
R6812 plus.n114 plus.n63 161.3
R6813 plus.n112 plus.n111 161.3
R6814 plus.n110 plus.n64 161.3
R6815 plus.n109 plus.n108 161.3
R6816 plus.n106 plus.n65 161.3
R6817 plus.n105 plus.n104 161.3
R6818 plus.n103 plus.n102 161.3
R6819 plus.n101 plus.n67 161.3
R6820 plus.n100 plus.n99 161.3
R6821 plus.n98 plus.n97 161.3
R6822 plus.n96 plus.n69 161.3
R6823 plus.n94 plus.n93 161.3
R6824 plus.n92 plus.n70 161.3
R6825 plus.n91 plus.n90 161.3
R6826 plus.n88 plus.n71 161.3
R6827 plus.n87 plus.n86 161.3
R6828 plus.n85 plus.n84 161.3
R6829 plus.n83 plus.n73 161.3
R6830 plus.n82 plus.n81 161.3
R6831 plus.n80 plus.n79 161.3
R6832 plus.n78 plus.n75 161.3
R6833 plus.n17 plus.n14 161.3
R6834 plus.n19 plus.n18 161.3
R6835 plus.n21 plus.n20 161.3
R6836 plus.n22 plus.n12 161.3
R6837 plus.n24 plus.n23 161.3
R6838 plus.n26 plus.n25 161.3
R6839 plus.n27 plus.n10 161.3
R6840 plus.n30 plus.n29 161.3
R6841 plus.n31 plus.n9 161.3
R6842 plus.n33 plus.n32 161.3
R6843 plus.n35 plus.n8 161.3
R6844 plus.n37 plus.n36 161.3
R6845 plus.n39 plus.n38 161.3
R6846 plus.n40 plus.n6 161.3
R6847 plus.n42 plus.n41 161.3
R6848 plus.n44 plus.n43 161.3
R6849 plus.n45 plus.n4 161.3
R6850 plus.n48 plus.n47 161.3
R6851 plus.n49 plus.n3 161.3
R6852 plus.n51 plus.n50 161.3
R6853 plus.n53 plus.n2 161.3
R6854 plus.n55 plus.n54 161.3
R6855 plus.n57 plus.n56 161.3
R6856 plus.n58 plus.n0 161.3
R6857 plus.n60 plus.n59 161.3
R6858 plus.n88 plus.n87 56.5617
R6859 plus.n97 plus.n96 56.5617
R6860 plus.n106 plus.n105 56.5617
R6861 plus.n45 plus.n44 56.5617
R6862 plus.n36 plus.n35 56.5617
R6863 plus.n27 plus.n26 56.5617
R6864 plus.n79 plus.n78 56.5617
R6865 plus.n115 plus.n114 56.5617
R6866 plus.n54 plus.n53 56.5617
R6867 plus.n18 plus.n17 56.5617
R6868 plus.n119 plus.n118 50.2647
R6869 plus.n58 plus.n57 50.2647
R6870 plus.n84 plus.n83 46.3896
R6871 plus.n108 plus.n64 46.3896
R6872 plus.n47 plus.n3 46.3896
R6873 plus.n23 plus.n22 46.3896
R6874 plus.n76 plus.n75 43.1929
R6875 plus.n15 plus.n14 43.1929
R6876 plus.n94 plus.n70 42.5146
R6877 plus.n101 plus.n100 42.5146
R6878 plus.n40 plus.n39 42.5146
R6879 plus.n33 plus.n9 42.5146
R6880 plus.n77 plus.n76 40.6041
R6881 plus.n16 plus.n15 40.6041
R6882 plus.n90 plus.n70 38.6395
R6883 plus.n102 plus.n101 38.6395
R6884 plus.n41 plus.n40 38.6395
R6885 plus.n29 plus.n9 38.6395
R6886 plus.n122 plus.n121 35.2031
R6887 plus.n83 plus.n82 34.7644
R6888 plus.n112 plus.n64 34.7644
R6889 plus.n51 plus.n3 34.7644
R6890 plus.n22 plus.n21 34.7644
R6891 plus.n79 plus.n74 21.8872
R6892 plus.n114 plus.n113 21.8872
R6893 plus.n53 plus.n52 21.8872
R6894 plus.n18 plus.n13 21.8872
R6895 plus.n89 plus.n88 19.9199
R6896 plus.n105 plus.n66 19.9199
R6897 plus.n44 plus.n5 19.9199
R6898 plus.n28 plus.n27 19.9199
R6899 plus.n123 plus.t4 19.8005
R6900 plus.n123 plus.t0 19.8005
R6901 plus.n125 plus.t3 19.8005
R6902 plus.n125 plus.t1 19.8005
R6903 plus.n96 plus.n95 17.9525
R6904 plus.n97 plus.n68 17.9525
R6905 plus.n36 plus.n7 17.9525
R6906 plus.n35 plus.n34 17.9525
R6907 plus.n87 plus.n72 15.9852
R6908 plus.n107 plus.n106 15.9852
R6909 plus.n46 plus.n45 15.9852
R6910 plus.n26 plus.n11 15.9852
R6911 plus plus.n127 15.3578
R6912 plus.n78 plus.n77 14.0178
R6913 plus.n115 plus.n62 14.0178
R6914 plus.n54 plus.n1 14.0178
R6915 plus.n17 plus.n16 14.0178
R6916 plus.n122 plus.n60 11.9342
R6917 plus.n118 plus.n62 10.575
R6918 plus.n57 plus.n1 10.575
R6919 plus.n120 plus.n119 9.49444
R6920 plus.n59 plus.n58 9.49444
R6921 plus.n84 plus.n72 8.60764
R6922 plus.n108 plus.n107 8.60764
R6923 plus.n47 plus.n46 8.60764
R6924 plus.n23 plus.n11 8.60764
R6925 plus.n95 plus.n94 6.6403
R6926 plus.n100 plus.n68 6.6403
R6927 plus.n39 plus.n7 6.6403
R6928 plus.n34 plus.n33 6.6403
R6929 plus.n127 plus.n126 5.40567
R6930 plus.n90 plus.n89 4.67295
R6931 plus.n102 plus.n66 4.67295
R6932 plus.n41 plus.n5 4.67295
R6933 plus.n29 plus.n28 4.67295
R6934 plus.n82 plus.n74 2.7056
R6935 plus.n113 plus.n112 2.7056
R6936 plus.n52 plus.n51 2.7056
R6937 plus.n21 plus.n13 2.7056
R6938 plus.n127 plus.n122 1.188
R6939 plus.n126 plus.n124 0.716017
R6940 plus.n80 plus.n75 0.189894
R6941 plus.n81 plus.n80 0.189894
R6942 plus.n81 plus.n73 0.189894
R6943 plus.n85 plus.n73 0.189894
R6944 plus.n86 plus.n85 0.189894
R6945 plus.n86 plus.n71 0.189894
R6946 plus.n91 plus.n71 0.189894
R6947 plus.n92 plus.n91 0.189894
R6948 plus.n93 plus.n92 0.189894
R6949 plus.n93 plus.n69 0.189894
R6950 plus.n98 plus.n69 0.189894
R6951 plus.n99 plus.n98 0.189894
R6952 plus.n99 plus.n67 0.189894
R6953 plus.n103 plus.n67 0.189894
R6954 plus.n104 plus.n103 0.189894
R6955 plus.n104 plus.n65 0.189894
R6956 plus.n109 plus.n65 0.189894
R6957 plus.n110 plus.n109 0.189894
R6958 plus.n111 plus.n110 0.189894
R6959 plus.n111 plus.n63 0.189894
R6960 plus.n116 plus.n63 0.189894
R6961 plus.n117 plus.n116 0.189894
R6962 plus.n117 plus.n61 0.189894
R6963 plus.n121 plus.n61 0.189894
R6964 plus.n60 plus.n0 0.189894
R6965 plus.n56 plus.n0 0.189894
R6966 plus.n56 plus.n55 0.189894
R6967 plus.n55 plus.n2 0.189894
R6968 plus.n50 plus.n2 0.189894
R6969 plus.n50 plus.n49 0.189894
R6970 plus.n49 plus.n48 0.189894
R6971 plus.n48 plus.n4 0.189894
R6972 plus.n43 plus.n4 0.189894
R6973 plus.n43 plus.n42 0.189894
R6974 plus.n42 plus.n6 0.189894
R6975 plus.n38 plus.n6 0.189894
R6976 plus.n38 plus.n37 0.189894
R6977 plus.n37 plus.n8 0.189894
R6978 plus.n32 plus.n8 0.189894
R6979 plus.n32 plus.n31 0.189894
R6980 plus.n31 plus.n30 0.189894
R6981 plus.n30 plus.n10 0.189894
R6982 plus.n25 plus.n10 0.189894
R6983 plus.n25 plus.n24 0.189894
R6984 plus.n24 plus.n12 0.189894
R6985 plus.n20 plus.n12 0.189894
R6986 plus.n20 plus.n19 0.189894
R6987 plus.n19 plus.n14 0.189894
R6988 a_n3827_n3924.n22 a_n3827_n3924.t27 214.938
R6989 a_n3827_n3924.n1 a_n3827_n3924.t57 214.409
R6990 a_n3827_n3924.n14 a_n3827_n3924.t26 214.321
R6991 a_n3827_n3924.n15 a_n3827_n3924.t55 214.321
R6992 a_n3827_n3924.n16 a_n3827_n3924.t46 214.321
R6993 a_n3827_n3924.n17 a_n3827_n3924.t56 214.321
R6994 a_n3827_n3924.n18 a_n3827_n3924.t25 214.321
R6995 a_n3827_n3924.n19 a_n3827_n3924.t54 214.321
R6996 a_n3827_n3924.n20 a_n3827_n3924.t24 214.321
R6997 a_n3827_n3924.n21 a_n3827_n3924.t28 214.321
R6998 a_n3827_n3924.n0 a_n3827_n3924.t17 55.8337
R6999 a_n3827_n3924.n2 a_n3827_n3924.t51 55.8337
R7000 a_n3827_n3924.n13 a_n3827_n3924.t31 55.8337
R7001 a_n3827_n3924.n49 a_n3827_n3924.t4 55.8335
R7002 a_n3827_n3924.n47 a_n3827_n3924.t35 55.8335
R7003 a_n3827_n3924.n36 a_n3827_n3924.t48 55.8335
R7004 a_n3827_n3924.n35 a_n3827_n3924.t14 55.8335
R7005 a_n3827_n3924.n24 a_n3827_n3924.t8 55.8335
R7006 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0052
R7007 a_n3827_n3924.n53 a_n3827_n3924.n52 53.0052
R7008 a_n3827_n3924.n55 a_n3827_n3924.n54 53.0052
R7009 a_n3827_n3924.n57 a_n3827_n3924.n56 53.0052
R7010 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R7011 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R7012 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R7013 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R7014 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R7015 a_n3827_n3924.n46 a_n3827_n3924.n45 53.0051
R7016 a_n3827_n3924.n44 a_n3827_n3924.n43 53.0051
R7017 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R7018 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R7019 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0051
R7020 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R7021 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R7022 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R7023 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R7024 a_n3827_n3924.n26 a_n3827_n3924.n25 53.0051
R7025 a_n3827_n3924.n59 a_n3827_n3924.n58 53.0051
R7026 a_n3827_n3924.n23 a_n3827_n3924.n13 12.2417
R7027 a_n3827_n3924.n49 a_n3827_n3924.n48 12.2417
R7028 a_n3827_n3924.n24 a_n3827_n3924.n23 5.16214
R7029 a_n3827_n3924.n48 a_n3827_n3924.n47 5.16214
R7030 a_n3827_n3924.n50 a_n3827_n3924.t2 2.82907
R7031 a_n3827_n3924.n50 a_n3827_n3924.t0 2.82907
R7032 a_n3827_n3924.n52 a_n3827_n3924.t13 2.82907
R7033 a_n3827_n3924.n52 a_n3827_n3924.t18 2.82907
R7034 a_n3827_n3924.n54 a_n3827_n3924.t11 2.82907
R7035 a_n3827_n3924.n54 a_n3827_n3924.t15 2.82907
R7036 a_n3827_n3924.n56 a_n3827_n3924.t7 2.82907
R7037 a_n3827_n3924.n56 a_n3827_n3924.t12 2.82907
R7038 a_n3827_n3924.n3 a_n3827_n3924.t38 2.82907
R7039 a_n3827_n3924.n3 a_n3827_n3924.t29 2.82907
R7040 a_n3827_n3924.n5 a_n3827_n3924.t33 2.82907
R7041 a_n3827_n3924.n5 a_n3827_n3924.t37 2.82907
R7042 a_n3827_n3924.n7 a_n3827_n3924.t49 2.82907
R7043 a_n3827_n3924.n7 a_n3827_n3924.t32 2.82907
R7044 a_n3827_n3924.n9 a_n3827_n3924.t42 2.82907
R7045 a_n3827_n3924.n9 a_n3827_n3924.t53 2.82907
R7046 a_n3827_n3924.n11 a_n3827_n3924.t44 2.82907
R7047 a_n3827_n3924.n11 a_n3827_n3924.t45 2.82907
R7048 a_n3827_n3924.n45 a_n3827_n3924.t41 2.82907
R7049 a_n3827_n3924.n45 a_n3827_n3924.t40 2.82907
R7050 a_n3827_n3924.n43 a_n3827_n3924.t43 2.82907
R7051 a_n3827_n3924.n43 a_n3827_n3924.t36 2.82907
R7052 a_n3827_n3924.n41 a_n3827_n3924.t52 2.82907
R7053 a_n3827_n3924.n41 a_n3827_n3924.t47 2.82907
R7054 a_n3827_n3924.n39 a_n3827_n3924.t34 2.82907
R7055 a_n3827_n3924.n39 a_n3827_n3924.t50 2.82907
R7056 a_n3827_n3924.n37 a_n3827_n3924.t39 2.82907
R7057 a_n3827_n3924.n37 a_n3827_n3924.t30 2.82907
R7058 a_n3827_n3924.n33 a_n3827_n3924.t3 2.82907
R7059 a_n3827_n3924.n33 a_n3827_n3924.t19 2.82907
R7060 a_n3827_n3924.n31 a_n3827_n3924.t10 2.82907
R7061 a_n3827_n3924.n31 a_n3827_n3924.t1 2.82907
R7062 a_n3827_n3924.n29 a_n3827_n3924.t21 2.82907
R7063 a_n3827_n3924.n29 a_n3827_n3924.t9 2.82907
R7064 a_n3827_n3924.n27 a_n3827_n3924.t16 2.82907
R7065 a_n3827_n3924.n27 a_n3827_n3924.t20 2.82907
R7066 a_n3827_n3924.n25 a_n3827_n3924.t5 2.82907
R7067 a_n3827_n3924.n25 a_n3827_n3924.t22 2.82907
R7068 a_n3827_n3924.t23 a_n3827_n3924.n59 2.82907
R7069 a_n3827_n3924.n59 a_n3827_n3924.t6 2.82907
R7070 a_n3827_n3924.n48 a_n3827_n3924.n1 1.95694
R7071 a_n3827_n3924.n23 a_n3827_n3924.n22 1.95694
R7072 a_n3827_n3924.n21 a_n3827_n3924.n20 0.672012
R7073 a_n3827_n3924.n20 a_n3827_n3924.n19 0.672012
R7074 a_n3827_n3924.n19 a_n3827_n3924.n18 0.672012
R7075 a_n3827_n3924.n18 a_n3827_n3924.n17 0.672012
R7076 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R7077 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R7078 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R7079 a_n3827_n3924.n14 a_n3827_n3924.n1 0.585529
R7080 a_n3827_n3924.n26 a_n3827_n3924.n24 0.530672
R7081 a_n3827_n3924.n28 a_n3827_n3924.n26 0.530672
R7082 a_n3827_n3924.n30 a_n3827_n3924.n28 0.530672
R7083 a_n3827_n3924.n32 a_n3827_n3924.n30 0.530672
R7084 a_n3827_n3924.n34 a_n3827_n3924.n32 0.530672
R7085 a_n3827_n3924.n35 a_n3827_n3924.n34 0.530672
R7086 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R7087 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R7088 a_n3827_n3924.n42 a_n3827_n3924.n40 0.530672
R7089 a_n3827_n3924.n44 a_n3827_n3924.n42 0.530672
R7090 a_n3827_n3924.n46 a_n3827_n3924.n44 0.530672
R7091 a_n3827_n3924.n47 a_n3827_n3924.n46 0.530672
R7092 a_n3827_n3924.n13 a_n3827_n3924.n12 0.530672
R7093 a_n3827_n3924.n12 a_n3827_n3924.n10 0.530672
R7094 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R7095 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R7096 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R7097 a_n3827_n3924.n4 a_n3827_n3924.n2 0.530672
R7098 a_n3827_n3924.n58 a_n3827_n3924.n0 0.530672
R7099 a_n3827_n3924.n58 a_n3827_n3924.n57 0.530672
R7100 a_n3827_n3924.n57 a_n3827_n3924.n55 0.530672
R7101 a_n3827_n3924.n55 a_n3827_n3924.n53 0.530672
R7102 a_n3827_n3924.n53 a_n3827_n3924.n51 0.530672
R7103 a_n3827_n3924.n51 a_n3827_n3924.n49 0.530672
R7104 a_n3827_n3924.n36 a_n3827_n3924.n35 0.235414
R7105 a_n3827_n3924.n2 a_n3827_n3924.n0 0.235414
R7106 a_n3827_n3924.n22 a_n3827_n3924.n21 0.0564593
R7107 gnd.n3608 gnd.n2228 766.379
R7108 gnd.n3611 gnd.n3610 766.379
R7109 gnd.n2850 gnd.n2753 766.379
R7110 gnd.n2846 gnd.n2751 766.379
R7111 gnd.n3699 gnd.n2250 756.769
R7112 gnd.n3602 gnd.n3601 756.769
R7113 gnd.n2943 gnd.n2660 756.769
R7114 gnd.n2941 gnd.n2663 756.769
R7115 gnd.n7397 gnd.n129 751.963
R7116 gnd.n7555 gnd.n7554 751.963
R7117 gnd.n7103 gnd.n452 751.963
R7118 gnd.n7156 gnd.n454 751.963
R7119 gnd.n4499 gnd.n1095 751.963
R7120 gnd.n4775 gnd.n4449 751.963
R7121 gnd.n4150 gnd.n3703 751.963
R7122 gnd.n4191 gnd.n3986 751.963
R7123 gnd.n7552 gnd.n131 732.745
R7124 gnd.n199 gnd.n127 732.745
R7125 gnd.n7029 gnd.n451 732.745
R7126 gnd.n7158 gnd.n449 732.745
R7127 gnd.n1959 gnd.n1090 732.745
R7128 gnd.n4790 gnd.n1992 732.745
R7129 gnd.n3842 gnd.n3702 732.745
R7130 gnd.n4193 gnd.n2226 732.745
R7131 gnd.n4763 gnd.n1101 711.122
R7132 gnd.n5900 gnd.n459 711.122
R7133 gnd.n4583 gnd.n4582 711.122
R7134 gnd.n5889 gnd.n1228 711.122
R7135 gnd.n6248 gnd.n922 655.866
R7136 gnd.n6575 gnd.n731 655.866
R7137 gnd.n6788 gnd.n6787 655.866
R7138 gnd.n6081 gnd.n6080 655.866
R7139 gnd.n6576 gnd.n730 636.496
R7140 gnd.n4406 gnd.n4405 585
R7141 gnd.n4406 gnd.n969 585
R7142 gnd.n4408 gnd.n4407 585
R7143 gnd.n4407 gnd.n927 585
R7144 gnd.n4409 gnd.n2012 585
R7145 gnd.n4424 gnd.n2012 585
R7146 gnd.n4410 gnd.n2022 585
R7147 gnd.n2022 gnd.n2010 585
R7148 gnd.n4412 gnd.n4411 585
R7149 gnd.n4413 gnd.n4412 585
R7150 gnd.n2023 gnd.n2021 585
R7151 gnd.n2029 gnd.n2021 585
R7152 gnd.n4394 gnd.n4393 585
R7153 gnd.n4393 gnd.n4392 585
R7154 gnd.n2026 gnd.n2025 585
R7155 gnd.n2038 gnd.n2026 585
R7156 gnd.n4383 gnd.n4382 585
R7157 gnd.n4384 gnd.n4383 585
R7158 gnd.n2040 gnd.n2039 585
R7159 gnd.n2039 gnd.n2035 585
R7160 gnd.n4378 gnd.n4377 585
R7161 gnd.n4377 gnd.n4376 585
R7162 gnd.n2043 gnd.n2042 585
R7163 gnd.n2044 gnd.n2043 585
R7164 gnd.n4367 gnd.n4366 585
R7165 gnd.n4368 gnd.n4367 585
R7166 gnd.n2055 gnd.n2054 585
R7167 gnd.n2061 gnd.n2054 585
R7168 gnd.n4362 gnd.n4361 585
R7169 gnd.n4361 gnd.n4360 585
R7170 gnd.n2058 gnd.n2057 585
R7171 gnd.n2070 gnd.n2058 585
R7172 gnd.n4351 gnd.n4350 585
R7173 gnd.n4352 gnd.n4351 585
R7174 gnd.n2072 gnd.n2071 585
R7175 gnd.n2071 gnd.n2067 585
R7176 gnd.n4346 gnd.n4345 585
R7177 gnd.n4345 gnd.n4344 585
R7178 gnd.n2075 gnd.n2074 585
R7179 gnd.n2076 gnd.n2075 585
R7180 gnd.n4335 gnd.n4334 585
R7181 gnd.n4336 gnd.n4335 585
R7182 gnd.n2087 gnd.n2086 585
R7183 gnd.n2093 gnd.n2086 585
R7184 gnd.n4330 gnd.n4329 585
R7185 gnd.n4329 gnd.n4328 585
R7186 gnd.n2090 gnd.n2089 585
R7187 gnd.n2102 gnd.n2090 585
R7188 gnd.n4319 gnd.n4318 585
R7189 gnd.n4320 gnd.n4319 585
R7190 gnd.n2104 gnd.n2103 585
R7191 gnd.n2103 gnd.n2099 585
R7192 gnd.n4314 gnd.n4313 585
R7193 gnd.n4313 gnd.n4312 585
R7194 gnd.n2108 gnd.n2107 585
R7195 gnd.n2109 gnd.n2108 585
R7196 gnd.n4303 gnd.n4302 585
R7197 gnd.n4304 gnd.n4303 585
R7198 gnd.n2121 gnd.n2120 585
R7199 gnd.n2120 gnd.n2117 585
R7200 gnd.n4298 gnd.n4297 585
R7201 gnd.n4297 gnd.n4296 585
R7202 gnd.n2124 gnd.n2123 585
R7203 gnd.n2135 gnd.n2124 585
R7204 gnd.n4287 gnd.n4286 585
R7205 gnd.n4288 gnd.n4287 585
R7206 gnd.n2137 gnd.n2136 585
R7207 gnd.n2136 gnd.n2132 585
R7208 gnd.n4282 gnd.n4281 585
R7209 gnd.n4281 gnd.n4280 585
R7210 gnd.n2140 gnd.n2139 585
R7211 gnd.n2141 gnd.n2140 585
R7212 gnd.n4271 gnd.n4270 585
R7213 gnd.n4272 gnd.n4271 585
R7214 gnd.n2153 gnd.n2152 585
R7215 gnd.n2152 gnd.n2149 585
R7216 gnd.n4266 gnd.n4265 585
R7217 gnd.n4265 gnd.n4264 585
R7218 gnd.n2156 gnd.n2155 585
R7219 gnd.n2167 gnd.n2156 585
R7220 gnd.n4255 gnd.n4254 585
R7221 gnd.n4256 gnd.n4255 585
R7222 gnd.n2169 gnd.n2168 585
R7223 gnd.n2168 gnd.n2164 585
R7224 gnd.n4250 gnd.n4249 585
R7225 gnd.n4249 gnd.n4248 585
R7226 gnd.n2172 gnd.n2171 585
R7227 gnd.n2173 gnd.n2172 585
R7228 gnd.n4239 gnd.n4238 585
R7229 gnd.n4240 gnd.n4239 585
R7230 gnd.n2185 gnd.n2184 585
R7231 gnd.n2184 gnd.n2181 585
R7232 gnd.n4234 gnd.n4233 585
R7233 gnd.n4233 gnd.n4232 585
R7234 gnd.n2188 gnd.n2187 585
R7235 gnd.n2199 gnd.n2188 585
R7236 gnd.n4223 gnd.n4222 585
R7237 gnd.n4224 gnd.n4223 585
R7238 gnd.n2201 gnd.n2200 585
R7239 gnd.n2200 gnd.n2196 585
R7240 gnd.n4218 gnd.n4217 585
R7241 gnd.n4217 gnd.n4216 585
R7242 gnd.n2204 gnd.n2203 585
R7243 gnd.n2205 gnd.n2204 585
R7244 gnd.n4207 gnd.n4206 585
R7245 gnd.n4208 gnd.n4207 585
R7246 gnd.n2217 gnd.n2216 585
R7247 gnd.n2216 gnd.n2213 585
R7248 gnd.n4202 gnd.n4201 585
R7249 gnd.n4201 gnd.n4200 585
R7250 gnd.n2220 gnd.n2219 585
R7251 gnd.n3985 gnd.n2220 585
R7252 gnd.n4191 gnd.n4190 585
R7253 gnd.n4192 gnd.n4191 585
R7254 gnd.n4187 gnd.n3986 585
R7255 gnd.n4186 gnd.n4185 585
R7256 gnd.n4183 gnd.n3988 585
R7257 gnd.n4181 gnd.n4180 585
R7258 gnd.n4179 gnd.n3989 585
R7259 gnd.n4178 gnd.n4177 585
R7260 gnd.n4175 gnd.n3994 585
R7261 gnd.n4173 gnd.n4172 585
R7262 gnd.n4171 gnd.n3995 585
R7263 gnd.n4170 gnd.n4169 585
R7264 gnd.n4167 gnd.n4000 585
R7265 gnd.n4165 gnd.n4164 585
R7266 gnd.n4163 gnd.n4001 585
R7267 gnd.n4162 gnd.n4161 585
R7268 gnd.n4159 gnd.n4006 585
R7269 gnd.n4157 gnd.n4156 585
R7270 gnd.n4155 gnd.n4007 585
R7271 gnd.n4149 gnd.n4012 585
R7272 gnd.n4151 gnd.n4150 585
R7273 gnd.n4150 gnd.n3701 585
R7274 gnd.n4428 gnd.n4427 585
R7275 gnd.n4427 gnd.n969 585
R7276 gnd.n4426 gnd.n2007 585
R7277 gnd.n4426 gnd.n927 585
R7278 gnd.n4425 gnd.n2009 585
R7279 gnd.n4425 gnd.n4424 585
R7280 gnd.n4064 gnd.n2008 585
R7281 gnd.n2010 gnd.n2008 585
R7282 gnd.n4068 gnd.n2020 585
R7283 gnd.n4413 gnd.n2020 585
R7284 gnd.n4069 gnd.n4063 585
R7285 gnd.n4063 gnd.n2029 585
R7286 gnd.n4070 gnd.n2028 585
R7287 gnd.n4392 gnd.n2028 585
R7288 gnd.n4061 gnd.n4060 585
R7289 gnd.n4060 gnd.n2038 585
R7290 gnd.n4074 gnd.n2037 585
R7291 gnd.n4384 gnd.n2037 585
R7292 gnd.n4075 gnd.n4059 585
R7293 gnd.n4059 gnd.n2035 585
R7294 gnd.n4076 gnd.n2046 585
R7295 gnd.n4376 gnd.n2046 585
R7296 gnd.n4057 gnd.n4056 585
R7297 gnd.n4056 gnd.n2044 585
R7298 gnd.n4080 gnd.n2053 585
R7299 gnd.n4368 gnd.n2053 585
R7300 gnd.n4081 gnd.n4055 585
R7301 gnd.n4055 gnd.n2061 585
R7302 gnd.n4082 gnd.n2060 585
R7303 gnd.n4360 gnd.n2060 585
R7304 gnd.n4053 gnd.n4052 585
R7305 gnd.n4052 gnd.n2070 585
R7306 gnd.n4086 gnd.n2069 585
R7307 gnd.n4352 gnd.n2069 585
R7308 gnd.n4087 gnd.n4051 585
R7309 gnd.n4051 gnd.n2067 585
R7310 gnd.n4088 gnd.n2078 585
R7311 gnd.n4344 gnd.n2078 585
R7312 gnd.n4049 gnd.n4048 585
R7313 gnd.n4048 gnd.n2076 585
R7314 gnd.n4092 gnd.n2085 585
R7315 gnd.n4336 gnd.n2085 585
R7316 gnd.n4093 gnd.n4047 585
R7317 gnd.n4047 gnd.n2093 585
R7318 gnd.n4094 gnd.n2092 585
R7319 gnd.n4328 gnd.n2092 585
R7320 gnd.n4045 gnd.n4044 585
R7321 gnd.n4044 gnd.n2102 585
R7322 gnd.n4098 gnd.n2101 585
R7323 gnd.n4320 gnd.n2101 585
R7324 gnd.n4100 gnd.n4099 585
R7325 gnd.n4099 gnd.n2099 585
R7326 gnd.n4101 gnd.n2111 585
R7327 gnd.n4312 gnd.n2111 585
R7328 gnd.n4103 gnd.n4102 585
R7329 gnd.n4102 gnd.n2109 585
R7330 gnd.n4104 gnd.n2119 585
R7331 gnd.n4304 gnd.n2119 585
R7332 gnd.n4106 gnd.n4105 585
R7333 gnd.n4105 gnd.n2117 585
R7334 gnd.n4107 gnd.n2126 585
R7335 gnd.n4296 gnd.n2126 585
R7336 gnd.n4109 gnd.n4108 585
R7337 gnd.n4108 gnd.n2135 585
R7338 gnd.n4110 gnd.n2134 585
R7339 gnd.n4288 gnd.n2134 585
R7340 gnd.n4112 gnd.n4111 585
R7341 gnd.n4111 gnd.n2132 585
R7342 gnd.n4113 gnd.n2143 585
R7343 gnd.n4280 gnd.n2143 585
R7344 gnd.n4115 gnd.n4114 585
R7345 gnd.n4114 gnd.n2141 585
R7346 gnd.n4116 gnd.n2151 585
R7347 gnd.n4272 gnd.n2151 585
R7348 gnd.n4118 gnd.n4117 585
R7349 gnd.n4117 gnd.n2149 585
R7350 gnd.n4119 gnd.n2158 585
R7351 gnd.n4264 gnd.n2158 585
R7352 gnd.n4121 gnd.n4120 585
R7353 gnd.n4120 gnd.n2167 585
R7354 gnd.n4122 gnd.n2166 585
R7355 gnd.n4256 gnd.n2166 585
R7356 gnd.n4124 gnd.n4123 585
R7357 gnd.n4123 gnd.n2164 585
R7358 gnd.n4125 gnd.n2175 585
R7359 gnd.n4248 gnd.n2175 585
R7360 gnd.n4127 gnd.n4126 585
R7361 gnd.n4126 gnd.n2173 585
R7362 gnd.n4128 gnd.n2183 585
R7363 gnd.n4240 gnd.n2183 585
R7364 gnd.n4130 gnd.n4129 585
R7365 gnd.n4129 gnd.n2181 585
R7366 gnd.n4131 gnd.n2190 585
R7367 gnd.n4232 gnd.n2190 585
R7368 gnd.n4133 gnd.n4132 585
R7369 gnd.n4132 gnd.n2199 585
R7370 gnd.n4134 gnd.n2198 585
R7371 gnd.n4224 gnd.n2198 585
R7372 gnd.n4136 gnd.n4135 585
R7373 gnd.n4135 gnd.n2196 585
R7374 gnd.n4137 gnd.n2207 585
R7375 gnd.n4216 gnd.n2207 585
R7376 gnd.n4139 gnd.n4138 585
R7377 gnd.n4138 gnd.n2205 585
R7378 gnd.n4140 gnd.n2215 585
R7379 gnd.n4208 gnd.n2215 585
R7380 gnd.n4142 gnd.n4141 585
R7381 gnd.n4141 gnd.n2213 585
R7382 gnd.n4143 gnd.n2222 585
R7383 gnd.n4200 gnd.n2222 585
R7384 gnd.n4145 gnd.n4144 585
R7385 gnd.n4144 gnd.n3985 585
R7386 gnd.n4146 gnd.n3703 585
R7387 gnd.n4192 gnd.n3703 585
R7388 gnd.n3608 gnd.n3607 585
R7389 gnd.n3609 gnd.n3608 585
R7390 gnd.n2303 gnd.n2302 585
R7391 gnd.n2309 gnd.n2302 585
R7392 gnd.n3583 gnd.n2321 585
R7393 gnd.n2321 gnd.n2308 585
R7394 gnd.n3585 gnd.n3584 585
R7395 gnd.n3586 gnd.n3585 585
R7396 gnd.n2322 gnd.n2320 585
R7397 gnd.n2320 gnd.n2316 585
R7398 gnd.n3317 gnd.n3316 585
R7399 gnd.n3316 gnd.n3315 585
R7400 gnd.n2327 gnd.n2326 585
R7401 gnd.n3286 gnd.n2327 585
R7402 gnd.n3306 gnd.n3305 585
R7403 gnd.n3305 gnd.n3304 585
R7404 gnd.n2334 gnd.n2333 585
R7405 gnd.n3292 gnd.n2334 585
R7406 gnd.n3262 gnd.n2354 585
R7407 gnd.n2354 gnd.n2353 585
R7408 gnd.n3264 gnd.n3263 585
R7409 gnd.n3265 gnd.n3264 585
R7410 gnd.n2355 gnd.n2352 585
R7411 gnd.n2363 gnd.n2352 585
R7412 gnd.n3240 gnd.n2375 585
R7413 gnd.n2375 gnd.n2362 585
R7414 gnd.n3242 gnd.n3241 585
R7415 gnd.n3243 gnd.n3242 585
R7416 gnd.n2376 gnd.n2374 585
R7417 gnd.n2374 gnd.n2370 585
R7418 gnd.n3228 gnd.n3227 585
R7419 gnd.n3227 gnd.n3226 585
R7420 gnd.n2381 gnd.n2380 585
R7421 gnd.n2391 gnd.n2381 585
R7422 gnd.n3217 gnd.n3216 585
R7423 gnd.n3216 gnd.n3215 585
R7424 gnd.n2388 gnd.n2387 585
R7425 gnd.n3203 gnd.n2388 585
R7426 gnd.n3177 gnd.n2409 585
R7427 gnd.n2409 gnd.n2398 585
R7428 gnd.n3179 gnd.n3178 585
R7429 gnd.n3180 gnd.n3179 585
R7430 gnd.n2410 gnd.n2408 585
R7431 gnd.n2418 gnd.n2408 585
R7432 gnd.n3155 gnd.n2430 585
R7433 gnd.n2430 gnd.n2417 585
R7434 gnd.n3157 gnd.n3156 585
R7435 gnd.n3158 gnd.n3157 585
R7436 gnd.n2431 gnd.n2429 585
R7437 gnd.n2429 gnd.n2425 585
R7438 gnd.n3143 gnd.n3142 585
R7439 gnd.n3142 gnd.n3141 585
R7440 gnd.n2436 gnd.n2435 585
R7441 gnd.n2445 gnd.n2436 585
R7442 gnd.n3132 gnd.n3131 585
R7443 gnd.n3131 gnd.n3130 585
R7444 gnd.n2443 gnd.n2442 585
R7445 gnd.n3118 gnd.n2443 585
R7446 gnd.n2556 gnd.n2555 585
R7447 gnd.n2556 gnd.n2452 585
R7448 gnd.n3075 gnd.n3074 585
R7449 gnd.n3074 gnd.n3073 585
R7450 gnd.n3076 gnd.n2550 585
R7451 gnd.n2561 gnd.n2550 585
R7452 gnd.n3078 gnd.n3077 585
R7453 gnd.n3079 gnd.n3078 585
R7454 gnd.n2551 gnd.n2549 585
R7455 gnd.n2574 gnd.n2549 585
R7456 gnd.n2534 gnd.n2533 585
R7457 gnd.n2537 gnd.n2534 585
R7458 gnd.n3089 gnd.n3088 585
R7459 gnd.n3088 gnd.n3087 585
R7460 gnd.n3090 gnd.n2528 585
R7461 gnd.n3049 gnd.n2528 585
R7462 gnd.n3092 gnd.n3091 585
R7463 gnd.n3093 gnd.n3092 585
R7464 gnd.n2529 gnd.n2527 585
R7465 gnd.n2588 gnd.n2527 585
R7466 gnd.n3041 gnd.n3040 585
R7467 gnd.n3040 gnd.n3039 585
R7468 gnd.n2585 gnd.n2584 585
R7469 gnd.n3023 gnd.n2585 585
R7470 gnd.n3010 gnd.n2604 585
R7471 gnd.n2604 gnd.n2603 585
R7472 gnd.n3012 gnd.n3011 585
R7473 gnd.n3013 gnd.n3012 585
R7474 gnd.n2605 gnd.n2602 585
R7475 gnd.n2611 gnd.n2602 585
R7476 gnd.n2991 gnd.n2990 585
R7477 gnd.n2992 gnd.n2991 585
R7478 gnd.n2622 gnd.n2621 585
R7479 gnd.n2621 gnd.n2617 585
R7480 gnd.n2981 gnd.n2980 585
R7481 gnd.n2982 gnd.n2981 585
R7482 gnd.n2632 gnd.n2631 585
R7483 gnd.n2637 gnd.n2631 585
R7484 gnd.n2959 gnd.n2650 585
R7485 gnd.n2650 gnd.n2636 585
R7486 gnd.n2961 gnd.n2960 585
R7487 gnd.n2962 gnd.n2961 585
R7488 gnd.n2651 gnd.n2649 585
R7489 gnd.n2649 gnd.n2645 585
R7490 gnd.n2950 gnd.n2949 585
R7491 gnd.n2951 gnd.n2950 585
R7492 gnd.n2658 gnd.n2657 585
R7493 gnd.n2662 gnd.n2657 585
R7494 gnd.n2927 gnd.n2679 585
R7495 gnd.n2679 gnd.n2661 585
R7496 gnd.n2929 gnd.n2928 585
R7497 gnd.n2930 gnd.n2929 585
R7498 gnd.n2680 gnd.n2678 585
R7499 gnd.n2678 gnd.n2669 585
R7500 gnd.n2922 gnd.n2921 585
R7501 gnd.n2921 gnd.n2920 585
R7502 gnd.n2727 gnd.n2726 585
R7503 gnd.n2728 gnd.n2727 585
R7504 gnd.n2881 gnd.n2880 585
R7505 gnd.n2882 gnd.n2881 585
R7506 gnd.n2737 gnd.n2736 585
R7507 gnd.n2736 gnd.n2735 585
R7508 gnd.n2876 gnd.n2875 585
R7509 gnd.n2875 gnd.n2874 585
R7510 gnd.n2740 gnd.n2739 585
R7511 gnd.n2741 gnd.n2740 585
R7512 gnd.n2865 gnd.n2864 585
R7513 gnd.n2866 gnd.n2865 585
R7514 gnd.n2748 gnd.n2747 585
R7515 gnd.n2857 gnd.n2747 585
R7516 gnd.n2860 gnd.n2859 585
R7517 gnd.n2859 gnd.n2858 585
R7518 gnd.n2751 gnd.n2750 585
R7519 gnd.n2752 gnd.n2751 585
R7520 gnd.n2846 gnd.n2845 585
R7521 gnd.n2844 gnd.n2770 585
R7522 gnd.n2843 gnd.n2769 585
R7523 gnd.n2848 gnd.n2769 585
R7524 gnd.n2842 gnd.n2841 585
R7525 gnd.n2840 gnd.n2839 585
R7526 gnd.n2838 gnd.n2837 585
R7527 gnd.n2836 gnd.n2835 585
R7528 gnd.n2834 gnd.n2833 585
R7529 gnd.n2832 gnd.n2831 585
R7530 gnd.n2830 gnd.n2829 585
R7531 gnd.n2828 gnd.n2827 585
R7532 gnd.n2826 gnd.n2825 585
R7533 gnd.n2824 gnd.n2823 585
R7534 gnd.n2822 gnd.n2821 585
R7535 gnd.n2820 gnd.n2819 585
R7536 gnd.n2818 gnd.n2817 585
R7537 gnd.n2816 gnd.n2815 585
R7538 gnd.n2814 gnd.n2813 585
R7539 gnd.n2812 gnd.n2811 585
R7540 gnd.n2810 gnd.n2809 585
R7541 gnd.n2808 gnd.n2807 585
R7542 gnd.n2806 gnd.n2805 585
R7543 gnd.n2804 gnd.n2803 585
R7544 gnd.n2802 gnd.n2801 585
R7545 gnd.n2800 gnd.n2799 585
R7546 gnd.n2757 gnd.n2756 585
R7547 gnd.n2851 gnd.n2850 585
R7548 gnd.n3612 gnd.n3611 585
R7549 gnd.n3614 gnd.n3613 585
R7550 gnd.n3616 gnd.n3615 585
R7551 gnd.n3618 gnd.n3617 585
R7552 gnd.n3620 gnd.n3619 585
R7553 gnd.n3622 gnd.n3621 585
R7554 gnd.n3624 gnd.n3623 585
R7555 gnd.n3626 gnd.n3625 585
R7556 gnd.n3628 gnd.n3627 585
R7557 gnd.n3630 gnd.n3629 585
R7558 gnd.n3632 gnd.n3631 585
R7559 gnd.n3634 gnd.n3633 585
R7560 gnd.n3636 gnd.n3635 585
R7561 gnd.n3638 gnd.n3637 585
R7562 gnd.n3640 gnd.n3639 585
R7563 gnd.n3642 gnd.n3641 585
R7564 gnd.n3644 gnd.n3643 585
R7565 gnd.n3646 gnd.n3645 585
R7566 gnd.n3648 gnd.n3647 585
R7567 gnd.n3650 gnd.n3649 585
R7568 gnd.n3652 gnd.n3651 585
R7569 gnd.n3654 gnd.n3653 585
R7570 gnd.n3656 gnd.n3655 585
R7571 gnd.n3658 gnd.n3657 585
R7572 gnd.n3660 gnd.n3659 585
R7573 gnd.n3661 gnd.n2270 585
R7574 gnd.n3662 gnd.n2228 585
R7575 gnd.n3700 gnd.n2228 585
R7576 gnd.n3610 gnd.n2300 585
R7577 gnd.n3610 gnd.n3609 585
R7578 gnd.n3279 gnd.n2299 585
R7579 gnd.n2309 gnd.n2299 585
R7580 gnd.n3281 gnd.n3280 585
R7581 gnd.n3280 gnd.n2308 585
R7582 gnd.n3282 gnd.n2318 585
R7583 gnd.n3586 gnd.n2318 585
R7584 gnd.n3284 gnd.n3283 585
R7585 gnd.n3283 gnd.n2316 585
R7586 gnd.n3285 gnd.n2329 585
R7587 gnd.n3315 gnd.n2329 585
R7588 gnd.n3288 gnd.n3287 585
R7589 gnd.n3287 gnd.n3286 585
R7590 gnd.n3289 gnd.n2336 585
R7591 gnd.n3304 gnd.n2336 585
R7592 gnd.n3291 gnd.n3290 585
R7593 gnd.n3292 gnd.n3291 585
R7594 gnd.n2346 gnd.n2345 585
R7595 gnd.n2353 gnd.n2345 585
R7596 gnd.n3267 gnd.n3266 585
R7597 gnd.n3266 gnd.n3265 585
R7598 gnd.n2349 gnd.n2348 585
R7599 gnd.n2363 gnd.n2349 585
R7600 gnd.n3193 gnd.n3192 585
R7601 gnd.n3192 gnd.n2362 585
R7602 gnd.n3194 gnd.n2372 585
R7603 gnd.n3243 gnd.n2372 585
R7604 gnd.n3196 gnd.n3195 585
R7605 gnd.n3195 gnd.n2370 585
R7606 gnd.n3197 gnd.n2383 585
R7607 gnd.n3226 gnd.n2383 585
R7608 gnd.n3199 gnd.n3198 585
R7609 gnd.n3198 gnd.n2391 585
R7610 gnd.n3200 gnd.n2390 585
R7611 gnd.n3215 gnd.n2390 585
R7612 gnd.n3202 gnd.n3201 585
R7613 gnd.n3203 gnd.n3202 585
R7614 gnd.n2402 gnd.n2401 585
R7615 gnd.n2401 gnd.n2398 585
R7616 gnd.n3182 gnd.n3181 585
R7617 gnd.n3181 gnd.n3180 585
R7618 gnd.n2405 gnd.n2404 585
R7619 gnd.n2418 gnd.n2405 585
R7620 gnd.n3106 gnd.n3105 585
R7621 gnd.n3105 gnd.n2417 585
R7622 gnd.n3107 gnd.n2427 585
R7623 gnd.n3158 gnd.n2427 585
R7624 gnd.n3109 gnd.n3108 585
R7625 gnd.n3108 gnd.n2425 585
R7626 gnd.n3110 gnd.n2438 585
R7627 gnd.n3141 gnd.n2438 585
R7628 gnd.n3112 gnd.n3111 585
R7629 gnd.n3111 gnd.n2445 585
R7630 gnd.n3113 gnd.n2444 585
R7631 gnd.n3130 gnd.n2444 585
R7632 gnd.n3115 gnd.n3114 585
R7633 gnd.n3118 gnd.n3115 585
R7634 gnd.n2455 gnd.n2454 585
R7635 gnd.n2454 gnd.n2452 585
R7636 gnd.n2558 gnd.n2557 585
R7637 gnd.n3073 gnd.n2557 585
R7638 gnd.n2560 gnd.n2559 585
R7639 gnd.n2561 gnd.n2560 585
R7640 gnd.n2571 gnd.n2547 585
R7641 gnd.n3079 gnd.n2547 585
R7642 gnd.n2573 gnd.n2572 585
R7643 gnd.n2574 gnd.n2573 585
R7644 gnd.n2570 gnd.n2569 585
R7645 gnd.n2570 gnd.n2537 585
R7646 gnd.n2568 gnd.n2535 585
R7647 gnd.n3087 gnd.n2535 585
R7648 gnd.n2524 gnd.n2522 585
R7649 gnd.n3049 gnd.n2524 585
R7650 gnd.n3095 gnd.n3094 585
R7651 gnd.n3094 gnd.n3093 585
R7652 gnd.n2523 gnd.n2521 585
R7653 gnd.n2588 gnd.n2523 585
R7654 gnd.n3020 gnd.n2587 585
R7655 gnd.n3039 gnd.n2587 585
R7656 gnd.n3022 gnd.n3021 585
R7657 gnd.n3023 gnd.n3022 585
R7658 gnd.n2597 gnd.n2596 585
R7659 gnd.n2603 gnd.n2596 585
R7660 gnd.n3015 gnd.n3014 585
R7661 gnd.n3014 gnd.n3013 585
R7662 gnd.n2600 gnd.n2599 585
R7663 gnd.n2611 gnd.n2600 585
R7664 gnd.n2900 gnd.n2619 585
R7665 gnd.n2992 gnd.n2619 585
R7666 gnd.n2902 gnd.n2901 585
R7667 gnd.n2901 gnd.n2617 585
R7668 gnd.n2903 gnd.n2630 585
R7669 gnd.n2982 gnd.n2630 585
R7670 gnd.n2905 gnd.n2904 585
R7671 gnd.n2905 gnd.n2637 585
R7672 gnd.n2907 gnd.n2906 585
R7673 gnd.n2906 gnd.n2636 585
R7674 gnd.n2908 gnd.n2647 585
R7675 gnd.n2962 gnd.n2647 585
R7676 gnd.n2910 gnd.n2909 585
R7677 gnd.n2909 gnd.n2645 585
R7678 gnd.n2911 gnd.n2656 585
R7679 gnd.n2951 gnd.n2656 585
R7680 gnd.n2913 gnd.n2912 585
R7681 gnd.n2913 gnd.n2662 585
R7682 gnd.n2915 gnd.n2914 585
R7683 gnd.n2914 gnd.n2661 585
R7684 gnd.n2916 gnd.n2677 585
R7685 gnd.n2930 gnd.n2677 585
R7686 gnd.n2917 gnd.n2730 585
R7687 gnd.n2730 gnd.n2669 585
R7688 gnd.n2919 gnd.n2918 585
R7689 gnd.n2920 gnd.n2919 585
R7690 gnd.n2731 gnd.n2729 585
R7691 gnd.n2729 gnd.n2728 585
R7692 gnd.n2884 gnd.n2883 585
R7693 gnd.n2883 gnd.n2882 585
R7694 gnd.n2734 gnd.n2733 585
R7695 gnd.n2735 gnd.n2734 585
R7696 gnd.n2873 gnd.n2872 585
R7697 gnd.n2874 gnd.n2873 585
R7698 gnd.n2743 gnd.n2742 585
R7699 gnd.n2742 gnd.n2741 585
R7700 gnd.n2868 gnd.n2867 585
R7701 gnd.n2867 gnd.n2866 585
R7702 gnd.n2746 gnd.n2745 585
R7703 gnd.n2857 gnd.n2746 585
R7704 gnd.n2856 gnd.n2855 585
R7705 gnd.n2858 gnd.n2856 585
R7706 gnd.n2754 gnd.n2753 585
R7707 gnd.n2753 gnd.n2752 585
R7708 gnd.n3595 gnd.n2250 585
R7709 gnd.n2250 gnd.n2227 585
R7710 gnd.n3596 gnd.n2311 585
R7711 gnd.n2311 gnd.n2301 585
R7712 gnd.n3598 gnd.n3597 585
R7713 gnd.n3599 gnd.n3598 585
R7714 gnd.n2312 gnd.n2310 585
R7715 gnd.n2319 gnd.n2310 585
R7716 gnd.n3589 gnd.n3588 585
R7717 gnd.n3588 gnd.n3587 585
R7718 gnd.n2315 gnd.n2314 585
R7719 gnd.n3314 gnd.n2315 585
R7720 gnd.n3300 gnd.n2338 585
R7721 gnd.n2338 gnd.n2328 585
R7722 gnd.n3302 gnd.n3301 585
R7723 gnd.n3303 gnd.n3302 585
R7724 gnd.n2339 gnd.n2337 585
R7725 gnd.n2337 gnd.n2335 585
R7726 gnd.n3295 gnd.n3294 585
R7727 gnd.n3294 gnd.n3293 585
R7728 gnd.n2342 gnd.n2341 585
R7729 gnd.n2351 gnd.n2342 585
R7730 gnd.n3251 gnd.n2365 585
R7731 gnd.n2365 gnd.n2350 585
R7732 gnd.n3253 gnd.n3252 585
R7733 gnd.n3254 gnd.n3253 585
R7734 gnd.n2366 gnd.n2364 585
R7735 gnd.n2373 gnd.n2364 585
R7736 gnd.n3246 gnd.n3245 585
R7737 gnd.n3245 gnd.n3244 585
R7738 gnd.n2369 gnd.n2368 585
R7739 gnd.n3225 gnd.n2369 585
R7740 gnd.n3211 gnd.n2393 585
R7741 gnd.n2393 gnd.n2382 585
R7742 gnd.n3213 gnd.n3212 585
R7743 gnd.n3214 gnd.n3213 585
R7744 gnd.n2394 gnd.n2392 585
R7745 gnd.n2392 gnd.n2389 585
R7746 gnd.n3206 gnd.n3205 585
R7747 gnd.n3205 gnd.n3204 585
R7748 gnd.n2397 gnd.n2396 585
R7749 gnd.n2407 gnd.n2397 585
R7750 gnd.n3166 gnd.n2420 585
R7751 gnd.n2420 gnd.n2406 585
R7752 gnd.n3168 gnd.n3167 585
R7753 gnd.n3169 gnd.n3168 585
R7754 gnd.n2421 gnd.n2419 585
R7755 gnd.n2428 gnd.n2419 585
R7756 gnd.n3161 gnd.n3160 585
R7757 gnd.n3160 gnd.n3159 585
R7758 gnd.n2424 gnd.n2423 585
R7759 gnd.n3140 gnd.n2424 585
R7760 gnd.n3126 gnd.n2447 585
R7761 gnd.n2447 gnd.n2437 585
R7762 gnd.n3128 gnd.n3127 585
R7763 gnd.n3129 gnd.n3128 585
R7764 gnd.n2448 gnd.n2446 585
R7765 gnd.n3117 gnd.n2446 585
R7766 gnd.n3121 gnd.n3120 585
R7767 gnd.n3120 gnd.n3119 585
R7768 gnd.n2451 gnd.n2450 585
R7769 gnd.n3072 gnd.n2451 585
R7770 gnd.n2565 gnd.n2564 585
R7771 gnd.n2566 gnd.n2565 585
R7772 gnd.n2545 gnd.n2544 585
R7773 gnd.n2548 gnd.n2545 585
R7774 gnd.n3082 gnd.n3081 585
R7775 gnd.n3081 gnd.n3080 585
R7776 gnd.n3083 gnd.n2539 585
R7777 gnd.n2575 gnd.n2539 585
R7778 gnd.n3085 gnd.n3084 585
R7779 gnd.n3086 gnd.n3085 585
R7780 gnd.n2540 gnd.n2538 585
R7781 gnd.n3050 gnd.n2538 585
R7782 gnd.n3034 gnd.n3033 585
R7783 gnd.n3033 gnd.n2526 585
R7784 gnd.n3035 gnd.n2590 585
R7785 gnd.n2590 gnd.n2525 585
R7786 gnd.n3037 gnd.n3036 585
R7787 gnd.n3038 gnd.n3037 585
R7788 gnd.n2591 gnd.n2589 585
R7789 gnd.n2589 gnd.n2586 585
R7790 gnd.n3026 gnd.n3025 585
R7791 gnd.n3025 gnd.n3024 585
R7792 gnd.n2594 gnd.n2593 585
R7793 gnd.n2601 gnd.n2594 585
R7794 gnd.n3000 gnd.n2999 585
R7795 gnd.n3001 gnd.n3000 585
R7796 gnd.n2613 gnd.n2612 585
R7797 gnd.n2620 gnd.n2612 585
R7798 gnd.n2995 gnd.n2994 585
R7799 gnd.n2994 gnd.n2993 585
R7800 gnd.n2616 gnd.n2615 585
R7801 gnd.n2983 gnd.n2616 585
R7802 gnd.n2970 gnd.n2640 585
R7803 gnd.n2640 gnd.n2639 585
R7804 gnd.n2972 gnd.n2971 585
R7805 gnd.n2973 gnd.n2972 585
R7806 gnd.n2641 gnd.n2638 585
R7807 gnd.n2648 gnd.n2638 585
R7808 gnd.n2965 gnd.n2964 585
R7809 gnd.n2964 gnd.n2963 585
R7810 gnd.n2644 gnd.n2643 585
R7811 gnd.n2952 gnd.n2644 585
R7812 gnd.n2939 gnd.n2665 585
R7813 gnd.n2665 gnd.n2664 585
R7814 gnd.n2941 gnd.n2940 585
R7815 gnd.n2942 gnd.n2941 585
R7816 gnd.n2935 gnd.n2663 585
R7817 gnd.n2934 gnd.n2933 585
R7818 gnd.n2668 gnd.n2667 585
R7819 gnd.n2931 gnd.n2668 585
R7820 gnd.n2690 gnd.n2689 585
R7821 gnd.n2693 gnd.n2692 585
R7822 gnd.n2691 gnd.n2686 585
R7823 gnd.n2698 gnd.n2697 585
R7824 gnd.n2700 gnd.n2699 585
R7825 gnd.n2703 gnd.n2702 585
R7826 gnd.n2701 gnd.n2684 585
R7827 gnd.n2708 gnd.n2707 585
R7828 gnd.n2710 gnd.n2709 585
R7829 gnd.n2713 gnd.n2712 585
R7830 gnd.n2711 gnd.n2682 585
R7831 gnd.n2718 gnd.n2717 585
R7832 gnd.n2722 gnd.n2719 585
R7833 gnd.n2723 gnd.n2660 585
R7834 gnd.n3601 gnd.n2265 585
R7835 gnd.n3668 gnd.n3667 585
R7836 gnd.n3670 gnd.n3669 585
R7837 gnd.n3672 gnd.n3671 585
R7838 gnd.n3674 gnd.n3673 585
R7839 gnd.n3676 gnd.n3675 585
R7840 gnd.n3678 gnd.n3677 585
R7841 gnd.n3680 gnd.n3679 585
R7842 gnd.n3682 gnd.n3681 585
R7843 gnd.n3684 gnd.n3683 585
R7844 gnd.n3686 gnd.n3685 585
R7845 gnd.n3688 gnd.n3687 585
R7846 gnd.n3690 gnd.n3689 585
R7847 gnd.n3693 gnd.n3692 585
R7848 gnd.n3691 gnd.n2253 585
R7849 gnd.n3697 gnd.n2251 585
R7850 gnd.n3699 gnd.n3698 585
R7851 gnd.n3700 gnd.n3699 585
R7852 gnd.n3602 gnd.n2306 585
R7853 gnd.n3602 gnd.n2227 585
R7854 gnd.n3604 gnd.n3603 585
R7855 gnd.n3603 gnd.n2301 585
R7856 gnd.n3600 gnd.n2305 585
R7857 gnd.n3600 gnd.n3599 585
R7858 gnd.n3579 gnd.n2307 585
R7859 gnd.n2319 gnd.n2307 585
R7860 gnd.n3578 gnd.n2317 585
R7861 gnd.n3587 gnd.n2317 585
R7862 gnd.n3313 gnd.n2324 585
R7863 gnd.n3314 gnd.n3313 585
R7864 gnd.n3312 gnd.n3311 585
R7865 gnd.n3312 gnd.n2328 585
R7866 gnd.n3310 gnd.n2330 585
R7867 gnd.n3303 gnd.n2330 585
R7868 gnd.n2343 gnd.n2331 585
R7869 gnd.n2343 gnd.n2335 585
R7870 gnd.n3259 gnd.n2344 585
R7871 gnd.n3293 gnd.n2344 585
R7872 gnd.n3258 gnd.n3257 585
R7873 gnd.n3257 gnd.n2351 585
R7874 gnd.n3256 gnd.n2359 585
R7875 gnd.n3256 gnd.n2350 585
R7876 gnd.n3255 gnd.n2361 585
R7877 gnd.n3255 gnd.n3254 585
R7878 gnd.n3234 gnd.n2360 585
R7879 gnd.n2373 gnd.n2360 585
R7880 gnd.n3233 gnd.n2371 585
R7881 gnd.n3244 gnd.n2371 585
R7882 gnd.n3224 gnd.n2378 585
R7883 gnd.n3225 gnd.n3224 585
R7884 gnd.n3223 gnd.n3222 585
R7885 gnd.n3223 gnd.n2382 585
R7886 gnd.n3221 gnd.n2384 585
R7887 gnd.n3214 gnd.n2384 585
R7888 gnd.n2399 gnd.n2385 585
R7889 gnd.n2399 gnd.n2389 585
R7890 gnd.n3174 gnd.n2400 585
R7891 gnd.n3204 gnd.n2400 585
R7892 gnd.n3173 gnd.n3172 585
R7893 gnd.n3172 gnd.n2407 585
R7894 gnd.n3171 gnd.n2414 585
R7895 gnd.n3171 gnd.n2406 585
R7896 gnd.n3170 gnd.n2416 585
R7897 gnd.n3170 gnd.n3169 585
R7898 gnd.n3149 gnd.n2415 585
R7899 gnd.n2428 gnd.n2415 585
R7900 gnd.n3148 gnd.n2426 585
R7901 gnd.n3159 gnd.n2426 585
R7902 gnd.n3139 gnd.n2433 585
R7903 gnd.n3140 gnd.n3139 585
R7904 gnd.n3138 gnd.n3137 585
R7905 gnd.n3138 gnd.n2437 585
R7906 gnd.n3136 gnd.n2439 585
R7907 gnd.n3129 gnd.n2439 585
R7908 gnd.n3116 gnd.n2440 585
R7909 gnd.n3117 gnd.n3116 585
R7910 gnd.n3069 gnd.n2453 585
R7911 gnd.n3119 gnd.n2453 585
R7912 gnd.n3071 gnd.n3070 585
R7913 gnd.n3072 gnd.n3071 585
R7914 gnd.n3064 gnd.n2567 585
R7915 gnd.n2567 gnd.n2566 585
R7916 gnd.n3062 gnd.n3061 585
R7917 gnd.n3061 gnd.n2548 585
R7918 gnd.n3059 gnd.n2546 585
R7919 gnd.n3080 gnd.n2546 585
R7920 gnd.n2577 gnd.n2576 585
R7921 gnd.n2576 gnd.n2575 585
R7922 gnd.n3053 gnd.n2536 585
R7923 gnd.n3086 gnd.n2536 585
R7924 gnd.n3052 gnd.n3051 585
R7925 gnd.n3051 gnd.n3050 585
R7926 gnd.n3048 gnd.n2579 585
R7927 gnd.n3048 gnd.n2526 585
R7928 gnd.n3047 gnd.n3046 585
R7929 gnd.n3047 gnd.n2525 585
R7930 gnd.n2582 gnd.n2581 585
R7931 gnd.n3038 gnd.n2581 585
R7932 gnd.n3006 gnd.n3005 585
R7933 gnd.n3005 gnd.n2586 585
R7934 gnd.n3007 gnd.n2595 585
R7935 gnd.n3024 gnd.n2595 585
R7936 gnd.n3004 gnd.n3003 585
R7937 gnd.n3003 gnd.n2601 585
R7938 gnd.n3002 gnd.n2609 585
R7939 gnd.n3002 gnd.n3001 585
R7940 gnd.n2987 gnd.n2610 585
R7941 gnd.n2620 gnd.n2610 585
R7942 gnd.n2986 gnd.n2618 585
R7943 gnd.n2993 gnd.n2618 585
R7944 gnd.n2985 gnd.n2984 585
R7945 gnd.n2984 gnd.n2983 585
R7946 gnd.n2629 gnd.n2626 585
R7947 gnd.n2639 gnd.n2629 585
R7948 gnd.n2975 gnd.n2974 585
R7949 gnd.n2974 gnd.n2973 585
R7950 gnd.n2635 gnd.n2634 585
R7951 gnd.n2648 gnd.n2635 585
R7952 gnd.n2955 gnd.n2646 585
R7953 gnd.n2963 gnd.n2646 585
R7954 gnd.n2954 gnd.n2953 585
R7955 gnd.n2953 gnd.n2952 585
R7956 gnd.n2655 gnd.n2653 585
R7957 gnd.n2664 gnd.n2655 585
R7958 gnd.n2944 gnd.n2943 585
R7959 gnd.n2943 gnd.n2942 585
R7960 gnd.n1062 gnd.n1060 585
R7961 gnd.n1060 gnd.n969 585
R7962 gnd.n4421 gnd.n2014 585
R7963 gnd.n2014 gnd.n927 585
R7964 gnd.n4423 gnd.n4422 585
R7965 gnd.n4424 gnd.n4423 585
R7966 gnd.n2015 gnd.n2013 585
R7967 gnd.n2013 gnd.n2010 585
R7968 gnd.n4415 gnd.n4414 585
R7969 gnd.n4414 gnd.n4413 585
R7970 gnd.n2018 gnd.n2017 585
R7971 gnd.n2029 gnd.n2018 585
R7972 gnd.n4391 gnd.n4390 585
R7973 gnd.n4392 gnd.n4391 585
R7974 gnd.n2031 gnd.n2030 585
R7975 gnd.n2038 gnd.n2030 585
R7976 gnd.n4386 gnd.n4385 585
R7977 gnd.n4385 gnd.n4384 585
R7978 gnd.n2034 gnd.n2033 585
R7979 gnd.n2035 gnd.n2034 585
R7980 gnd.n4375 gnd.n4374 585
R7981 gnd.n4376 gnd.n4375 585
R7982 gnd.n2048 gnd.n2047 585
R7983 gnd.n2047 gnd.n2044 585
R7984 gnd.n4370 gnd.n4369 585
R7985 gnd.n4369 gnd.n4368 585
R7986 gnd.n2051 gnd.n2050 585
R7987 gnd.n2061 gnd.n2051 585
R7988 gnd.n4359 gnd.n4358 585
R7989 gnd.n4360 gnd.n4359 585
R7990 gnd.n2063 gnd.n2062 585
R7991 gnd.n2070 gnd.n2062 585
R7992 gnd.n4354 gnd.n4353 585
R7993 gnd.n4353 gnd.n4352 585
R7994 gnd.n2066 gnd.n2065 585
R7995 gnd.n2067 gnd.n2066 585
R7996 gnd.n4343 gnd.n4342 585
R7997 gnd.n4344 gnd.n4343 585
R7998 gnd.n2080 gnd.n2079 585
R7999 gnd.n2079 gnd.n2076 585
R8000 gnd.n4338 gnd.n4337 585
R8001 gnd.n4337 gnd.n4336 585
R8002 gnd.n2083 gnd.n2082 585
R8003 gnd.n2093 gnd.n2083 585
R8004 gnd.n4327 gnd.n4326 585
R8005 gnd.n4328 gnd.n4327 585
R8006 gnd.n2095 gnd.n2094 585
R8007 gnd.n2102 gnd.n2094 585
R8008 gnd.n4322 gnd.n4321 585
R8009 gnd.n4321 gnd.n4320 585
R8010 gnd.n2098 gnd.n2097 585
R8011 gnd.n2099 gnd.n2098 585
R8012 gnd.n4311 gnd.n4310 585
R8013 gnd.n4312 gnd.n4311 585
R8014 gnd.n2113 gnd.n2112 585
R8015 gnd.n2112 gnd.n2109 585
R8016 gnd.n4306 gnd.n4305 585
R8017 gnd.n4305 gnd.n4304 585
R8018 gnd.n2116 gnd.n2115 585
R8019 gnd.n2117 gnd.n2116 585
R8020 gnd.n4295 gnd.n4294 585
R8021 gnd.n4296 gnd.n4295 585
R8022 gnd.n2128 gnd.n2127 585
R8023 gnd.n2135 gnd.n2127 585
R8024 gnd.n4290 gnd.n4289 585
R8025 gnd.n4289 gnd.n4288 585
R8026 gnd.n2131 gnd.n2130 585
R8027 gnd.n2132 gnd.n2131 585
R8028 gnd.n4279 gnd.n4278 585
R8029 gnd.n4280 gnd.n4279 585
R8030 gnd.n2145 gnd.n2144 585
R8031 gnd.n2144 gnd.n2141 585
R8032 gnd.n4274 gnd.n4273 585
R8033 gnd.n4273 gnd.n4272 585
R8034 gnd.n2148 gnd.n2147 585
R8035 gnd.n2149 gnd.n2148 585
R8036 gnd.n4263 gnd.n4262 585
R8037 gnd.n4264 gnd.n4263 585
R8038 gnd.n2160 gnd.n2159 585
R8039 gnd.n2167 gnd.n2159 585
R8040 gnd.n4258 gnd.n4257 585
R8041 gnd.n4257 gnd.n4256 585
R8042 gnd.n2163 gnd.n2162 585
R8043 gnd.n2164 gnd.n2163 585
R8044 gnd.n4247 gnd.n4246 585
R8045 gnd.n4248 gnd.n4247 585
R8046 gnd.n2177 gnd.n2176 585
R8047 gnd.n2176 gnd.n2173 585
R8048 gnd.n4242 gnd.n4241 585
R8049 gnd.n4241 gnd.n4240 585
R8050 gnd.n2180 gnd.n2179 585
R8051 gnd.n2181 gnd.n2180 585
R8052 gnd.n4231 gnd.n4230 585
R8053 gnd.n4232 gnd.n4231 585
R8054 gnd.n2192 gnd.n2191 585
R8055 gnd.n2199 gnd.n2191 585
R8056 gnd.n4226 gnd.n4225 585
R8057 gnd.n4225 gnd.n4224 585
R8058 gnd.n2195 gnd.n2194 585
R8059 gnd.n2196 gnd.n2195 585
R8060 gnd.n4215 gnd.n4214 585
R8061 gnd.n4216 gnd.n4215 585
R8062 gnd.n2209 gnd.n2208 585
R8063 gnd.n2208 gnd.n2205 585
R8064 gnd.n4210 gnd.n4209 585
R8065 gnd.n4209 gnd.n4208 585
R8066 gnd.n2212 gnd.n2211 585
R8067 gnd.n2213 gnd.n2212 585
R8068 gnd.n4199 gnd.n4198 585
R8069 gnd.n4200 gnd.n4199 585
R8070 gnd.n2224 gnd.n2223 585
R8071 gnd.n3985 gnd.n2223 585
R8072 gnd.n4194 gnd.n4193 585
R8073 gnd.n4193 gnd.n4192 585
R8074 gnd.n3748 gnd.n2226 585
R8075 gnd.n3751 gnd.n3750 585
R8076 gnd.n3747 gnd.n3746 585
R8077 gnd.n3746 gnd.n3701 585
R8078 gnd.n3756 gnd.n3755 585
R8079 gnd.n3758 gnd.n3745 585
R8080 gnd.n3761 gnd.n3760 585
R8081 gnd.n3743 gnd.n3742 585
R8082 gnd.n3766 gnd.n3765 585
R8083 gnd.n3768 gnd.n3741 585
R8084 gnd.n3771 gnd.n3770 585
R8085 gnd.n3739 gnd.n3738 585
R8086 gnd.n3776 gnd.n3775 585
R8087 gnd.n3778 gnd.n3737 585
R8088 gnd.n3781 gnd.n3780 585
R8089 gnd.n3735 gnd.n3734 585
R8090 gnd.n3786 gnd.n3785 585
R8091 gnd.n3788 gnd.n3730 585
R8092 gnd.n3791 gnd.n3790 585
R8093 gnd.n3728 gnd.n3727 585
R8094 gnd.n3796 gnd.n3795 585
R8095 gnd.n3798 gnd.n3726 585
R8096 gnd.n3801 gnd.n3800 585
R8097 gnd.n3724 gnd.n3723 585
R8098 gnd.n3806 gnd.n3805 585
R8099 gnd.n3808 gnd.n3722 585
R8100 gnd.n3811 gnd.n3810 585
R8101 gnd.n3720 gnd.n3719 585
R8102 gnd.n3816 gnd.n3815 585
R8103 gnd.n3818 gnd.n3718 585
R8104 gnd.n3821 gnd.n3820 585
R8105 gnd.n3716 gnd.n3715 585
R8106 gnd.n3826 gnd.n3825 585
R8107 gnd.n3828 gnd.n3714 585
R8108 gnd.n3831 gnd.n3830 585
R8109 gnd.n3712 gnd.n3711 585
R8110 gnd.n3837 gnd.n3836 585
R8111 gnd.n3839 gnd.n3710 585
R8112 gnd.n3840 gnd.n3709 585
R8113 gnd.n3843 gnd.n3842 585
R8114 gnd.n3899 gnd.n3898 585
R8115 gnd.n3899 gnd.n969 585
R8116 gnd.n3901 gnd.n3900 585
R8117 gnd.n3900 gnd.n927 585
R8118 gnd.n3902 gnd.n2011 585
R8119 gnd.n4424 gnd.n2011 585
R8120 gnd.n3904 gnd.n3903 585
R8121 gnd.n3903 gnd.n2010 585
R8122 gnd.n3905 gnd.n2019 585
R8123 gnd.n4413 gnd.n2019 585
R8124 gnd.n3907 gnd.n3906 585
R8125 gnd.n3906 gnd.n2029 585
R8126 gnd.n3908 gnd.n2027 585
R8127 gnd.n4392 gnd.n2027 585
R8128 gnd.n3910 gnd.n3909 585
R8129 gnd.n3909 gnd.n2038 585
R8130 gnd.n3911 gnd.n2036 585
R8131 gnd.n4384 gnd.n2036 585
R8132 gnd.n3913 gnd.n3912 585
R8133 gnd.n3912 gnd.n2035 585
R8134 gnd.n3914 gnd.n2045 585
R8135 gnd.n4376 gnd.n2045 585
R8136 gnd.n3916 gnd.n3915 585
R8137 gnd.n3915 gnd.n2044 585
R8138 gnd.n3917 gnd.n2052 585
R8139 gnd.n4368 gnd.n2052 585
R8140 gnd.n3919 gnd.n3918 585
R8141 gnd.n3918 gnd.n2061 585
R8142 gnd.n3920 gnd.n2059 585
R8143 gnd.n4360 gnd.n2059 585
R8144 gnd.n3922 gnd.n3921 585
R8145 gnd.n3921 gnd.n2070 585
R8146 gnd.n3923 gnd.n2068 585
R8147 gnd.n4352 gnd.n2068 585
R8148 gnd.n3925 gnd.n3924 585
R8149 gnd.n3924 gnd.n2067 585
R8150 gnd.n3926 gnd.n2077 585
R8151 gnd.n4344 gnd.n2077 585
R8152 gnd.n3928 gnd.n3927 585
R8153 gnd.n3927 gnd.n2076 585
R8154 gnd.n3929 gnd.n2084 585
R8155 gnd.n4336 gnd.n2084 585
R8156 gnd.n3931 gnd.n3930 585
R8157 gnd.n3930 gnd.n2093 585
R8158 gnd.n3932 gnd.n2091 585
R8159 gnd.n4328 gnd.n2091 585
R8160 gnd.n3934 gnd.n3933 585
R8161 gnd.n3933 gnd.n2102 585
R8162 gnd.n3935 gnd.n2100 585
R8163 gnd.n4320 gnd.n2100 585
R8164 gnd.n3937 gnd.n3936 585
R8165 gnd.n3936 gnd.n2099 585
R8166 gnd.n3938 gnd.n2110 585
R8167 gnd.n4312 gnd.n2110 585
R8168 gnd.n3940 gnd.n3939 585
R8169 gnd.n3939 gnd.n2109 585
R8170 gnd.n3941 gnd.n2118 585
R8171 gnd.n4304 gnd.n2118 585
R8172 gnd.n3943 gnd.n3942 585
R8173 gnd.n3942 gnd.n2117 585
R8174 gnd.n3944 gnd.n2125 585
R8175 gnd.n4296 gnd.n2125 585
R8176 gnd.n3946 gnd.n3945 585
R8177 gnd.n3945 gnd.n2135 585
R8178 gnd.n3947 gnd.n2133 585
R8179 gnd.n4288 gnd.n2133 585
R8180 gnd.n3949 gnd.n3948 585
R8181 gnd.n3948 gnd.n2132 585
R8182 gnd.n3950 gnd.n2142 585
R8183 gnd.n4280 gnd.n2142 585
R8184 gnd.n3952 gnd.n3951 585
R8185 gnd.n3951 gnd.n2141 585
R8186 gnd.n3953 gnd.n2150 585
R8187 gnd.n4272 gnd.n2150 585
R8188 gnd.n3955 gnd.n3954 585
R8189 gnd.n3954 gnd.n2149 585
R8190 gnd.n3956 gnd.n2157 585
R8191 gnd.n4264 gnd.n2157 585
R8192 gnd.n3958 gnd.n3957 585
R8193 gnd.n3957 gnd.n2167 585
R8194 gnd.n3959 gnd.n2165 585
R8195 gnd.n4256 gnd.n2165 585
R8196 gnd.n3961 gnd.n3960 585
R8197 gnd.n3960 gnd.n2164 585
R8198 gnd.n3962 gnd.n2174 585
R8199 gnd.n4248 gnd.n2174 585
R8200 gnd.n3964 gnd.n3963 585
R8201 gnd.n3963 gnd.n2173 585
R8202 gnd.n3965 gnd.n2182 585
R8203 gnd.n4240 gnd.n2182 585
R8204 gnd.n3967 gnd.n3966 585
R8205 gnd.n3966 gnd.n2181 585
R8206 gnd.n3968 gnd.n2189 585
R8207 gnd.n4232 gnd.n2189 585
R8208 gnd.n3970 gnd.n3969 585
R8209 gnd.n3969 gnd.n2199 585
R8210 gnd.n3971 gnd.n2197 585
R8211 gnd.n4224 gnd.n2197 585
R8212 gnd.n3973 gnd.n3972 585
R8213 gnd.n3972 gnd.n2196 585
R8214 gnd.n3974 gnd.n2206 585
R8215 gnd.n4216 gnd.n2206 585
R8216 gnd.n3976 gnd.n3975 585
R8217 gnd.n3975 gnd.n2205 585
R8218 gnd.n3977 gnd.n2214 585
R8219 gnd.n4208 gnd.n2214 585
R8220 gnd.n3979 gnd.n3978 585
R8221 gnd.n3978 gnd.n2213 585
R8222 gnd.n3705 gnd.n2221 585
R8223 gnd.n4200 gnd.n2221 585
R8224 gnd.n3984 gnd.n3983 585
R8225 gnd.n3985 gnd.n3984 585
R8226 gnd.n3704 gnd.n3702 585
R8227 gnd.n4192 gnd.n3702 585
R8228 gnd.n6249 gnd.n6248 585
R8229 gnd.n926 gnd.n925 585
R8230 gnd.n6245 gnd.n6244 585
R8231 gnd.n6246 gnd.n6245 585
R8232 gnd.n6243 gnd.n970 585
R8233 gnd.n6242 gnd.n6241 585
R8234 gnd.n6240 gnd.n6239 585
R8235 gnd.n6238 gnd.n6237 585
R8236 gnd.n6236 gnd.n6235 585
R8237 gnd.n6234 gnd.n6233 585
R8238 gnd.n6232 gnd.n6231 585
R8239 gnd.n6230 gnd.n6229 585
R8240 gnd.n6228 gnd.n6227 585
R8241 gnd.n6226 gnd.n6225 585
R8242 gnd.n6224 gnd.n6223 585
R8243 gnd.n6222 gnd.n6221 585
R8244 gnd.n6220 gnd.n6219 585
R8245 gnd.n6218 gnd.n6217 585
R8246 gnd.n6216 gnd.n6215 585
R8247 gnd.n6214 gnd.n6213 585
R8248 gnd.n6212 gnd.n6211 585
R8249 gnd.n6210 gnd.n6209 585
R8250 gnd.n6208 gnd.n6207 585
R8251 gnd.n6206 gnd.n6205 585
R8252 gnd.n6204 gnd.n6203 585
R8253 gnd.n6202 gnd.n6201 585
R8254 gnd.n6200 gnd.n6199 585
R8255 gnd.n6198 gnd.n6197 585
R8256 gnd.n6196 gnd.n6195 585
R8257 gnd.n6194 gnd.n6193 585
R8258 gnd.n6192 gnd.n6191 585
R8259 gnd.n6190 gnd.n6189 585
R8260 gnd.n6188 gnd.n6187 585
R8261 gnd.n6186 gnd.n6185 585
R8262 gnd.n6184 gnd.n6183 585
R8263 gnd.n6182 gnd.n6181 585
R8264 gnd.n6180 gnd.n6179 585
R8265 gnd.n6178 gnd.n6177 585
R8266 gnd.n6176 gnd.n6175 585
R8267 gnd.n6174 gnd.n6173 585
R8268 gnd.n6172 gnd.n6171 585
R8269 gnd.n6170 gnd.n6169 585
R8270 gnd.n6168 gnd.n6167 585
R8271 gnd.n6166 gnd.n6165 585
R8272 gnd.n6164 gnd.n6163 585
R8273 gnd.n6162 gnd.n6161 585
R8274 gnd.n6160 gnd.n6159 585
R8275 gnd.n6158 gnd.n6157 585
R8276 gnd.n6156 gnd.n6155 585
R8277 gnd.n6154 gnd.n6153 585
R8278 gnd.n6152 gnd.n6151 585
R8279 gnd.n6150 gnd.n6149 585
R8280 gnd.n6148 gnd.n6147 585
R8281 gnd.n6146 gnd.n6145 585
R8282 gnd.n6144 gnd.n6143 585
R8283 gnd.n6142 gnd.n6141 585
R8284 gnd.n6140 gnd.n6139 585
R8285 gnd.n6138 gnd.n6137 585
R8286 gnd.n6136 gnd.n6135 585
R8287 gnd.n6134 gnd.n6133 585
R8288 gnd.n6132 gnd.n6131 585
R8289 gnd.n6130 gnd.n6129 585
R8290 gnd.n6128 gnd.n6127 585
R8291 gnd.n6126 gnd.n6125 585
R8292 gnd.n6124 gnd.n6123 585
R8293 gnd.n6122 gnd.n6121 585
R8294 gnd.n6120 gnd.n6119 585
R8295 gnd.n6118 gnd.n6117 585
R8296 gnd.n6116 gnd.n6115 585
R8297 gnd.n6114 gnd.n6113 585
R8298 gnd.n6112 gnd.n6111 585
R8299 gnd.n6110 gnd.n6109 585
R8300 gnd.n6108 gnd.n6107 585
R8301 gnd.n6106 gnd.n6105 585
R8302 gnd.n6104 gnd.n6103 585
R8303 gnd.n6102 gnd.n6101 585
R8304 gnd.n6100 gnd.n6099 585
R8305 gnd.n6098 gnd.n6097 585
R8306 gnd.n6096 gnd.n6095 585
R8307 gnd.n6094 gnd.n6093 585
R8308 gnd.n6092 gnd.n6091 585
R8309 gnd.n6090 gnd.n6089 585
R8310 gnd.n6088 gnd.n6087 585
R8311 gnd.n6086 gnd.n6085 585
R8312 gnd.n6084 gnd.n6083 585
R8313 gnd.n6082 gnd.n6081 585
R8314 gnd.n923 gnd.n922 585
R8315 gnd.n922 gnd.n921 585
R8316 gnd.n6254 gnd.n6253 585
R8317 gnd.n6255 gnd.n6254 585
R8318 gnd.n920 gnd.n919 585
R8319 gnd.n6256 gnd.n920 585
R8320 gnd.n6259 gnd.n6258 585
R8321 gnd.n6258 gnd.n6257 585
R8322 gnd.n917 gnd.n916 585
R8323 gnd.n916 gnd.n915 585
R8324 gnd.n6264 gnd.n6263 585
R8325 gnd.n6265 gnd.n6264 585
R8326 gnd.n914 gnd.n913 585
R8327 gnd.n6266 gnd.n914 585
R8328 gnd.n6269 gnd.n6268 585
R8329 gnd.n6268 gnd.n6267 585
R8330 gnd.n911 gnd.n910 585
R8331 gnd.n910 gnd.n909 585
R8332 gnd.n6274 gnd.n6273 585
R8333 gnd.n6275 gnd.n6274 585
R8334 gnd.n908 gnd.n907 585
R8335 gnd.n6276 gnd.n908 585
R8336 gnd.n6279 gnd.n6278 585
R8337 gnd.n6278 gnd.n6277 585
R8338 gnd.n905 gnd.n904 585
R8339 gnd.n904 gnd.n903 585
R8340 gnd.n6284 gnd.n6283 585
R8341 gnd.n6285 gnd.n6284 585
R8342 gnd.n902 gnd.n901 585
R8343 gnd.n6286 gnd.n902 585
R8344 gnd.n6289 gnd.n6288 585
R8345 gnd.n6288 gnd.n6287 585
R8346 gnd.n899 gnd.n898 585
R8347 gnd.n898 gnd.n897 585
R8348 gnd.n6294 gnd.n6293 585
R8349 gnd.n6295 gnd.n6294 585
R8350 gnd.n896 gnd.n895 585
R8351 gnd.n6296 gnd.n896 585
R8352 gnd.n6299 gnd.n6298 585
R8353 gnd.n6298 gnd.n6297 585
R8354 gnd.n893 gnd.n892 585
R8355 gnd.n892 gnd.n891 585
R8356 gnd.n6304 gnd.n6303 585
R8357 gnd.n6305 gnd.n6304 585
R8358 gnd.n890 gnd.n889 585
R8359 gnd.n6306 gnd.n890 585
R8360 gnd.n6309 gnd.n6308 585
R8361 gnd.n6308 gnd.n6307 585
R8362 gnd.n887 gnd.n886 585
R8363 gnd.n886 gnd.n885 585
R8364 gnd.n6314 gnd.n6313 585
R8365 gnd.n6315 gnd.n6314 585
R8366 gnd.n884 gnd.n883 585
R8367 gnd.n6316 gnd.n884 585
R8368 gnd.n6319 gnd.n6318 585
R8369 gnd.n6318 gnd.n6317 585
R8370 gnd.n881 gnd.n880 585
R8371 gnd.n880 gnd.n879 585
R8372 gnd.n6324 gnd.n6323 585
R8373 gnd.n6325 gnd.n6324 585
R8374 gnd.n878 gnd.n877 585
R8375 gnd.n6326 gnd.n878 585
R8376 gnd.n6329 gnd.n6328 585
R8377 gnd.n6328 gnd.n6327 585
R8378 gnd.n875 gnd.n874 585
R8379 gnd.n874 gnd.n873 585
R8380 gnd.n6334 gnd.n6333 585
R8381 gnd.n6335 gnd.n6334 585
R8382 gnd.n872 gnd.n871 585
R8383 gnd.n6336 gnd.n872 585
R8384 gnd.n6339 gnd.n6338 585
R8385 gnd.n6338 gnd.n6337 585
R8386 gnd.n869 gnd.n868 585
R8387 gnd.n868 gnd.n867 585
R8388 gnd.n6344 gnd.n6343 585
R8389 gnd.n6345 gnd.n6344 585
R8390 gnd.n866 gnd.n865 585
R8391 gnd.n6346 gnd.n866 585
R8392 gnd.n6349 gnd.n6348 585
R8393 gnd.n6348 gnd.n6347 585
R8394 gnd.n863 gnd.n862 585
R8395 gnd.n862 gnd.n861 585
R8396 gnd.n6354 gnd.n6353 585
R8397 gnd.n6355 gnd.n6354 585
R8398 gnd.n860 gnd.n859 585
R8399 gnd.n6356 gnd.n860 585
R8400 gnd.n6359 gnd.n6358 585
R8401 gnd.n6358 gnd.n6357 585
R8402 gnd.n857 gnd.n856 585
R8403 gnd.n856 gnd.n855 585
R8404 gnd.n6364 gnd.n6363 585
R8405 gnd.n6365 gnd.n6364 585
R8406 gnd.n854 gnd.n853 585
R8407 gnd.n6366 gnd.n854 585
R8408 gnd.n6369 gnd.n6368 585
R8409 gnd.n6368 gnd.n6367 585
R8410 gnd.n851 gnd.n850 585
R8411 gnd.n850 gnd.n849 585
R8412 gnd.n6374 gnd.n6373 585
R8413 gnd.n6375 gnd.n6374 585
R8414 gnd.n848 gnd.n847 585
R8415 gnd.n6376 gnd.n848 585
R8416 gnd.n6379 gnd.n6378 585
R8417 gnd.n6378 gnd.n6377 585
R8418 gnd.n845 gnd.n844 585
R8419 gnd.n844 gnd.n843 585
R8420 gnd.n6384 gnd.n6383 585
R8421 gnd.n6385 gnd.n6384 585
R8422 gnd.n842 gnd.n841 585
R8423 gnd.n6386 gnd.n842 585
R8424 gnd.n6389 gnd.n6388 585
R8425 gnd.n6388 gnd.n6387 585
R8426 gnd.n839 gnd.n838 585
R8427 gnd.n838 gnd.n837 585
R8428 gnd.n6394 gnd.n6393 585
R8429 gnd.n6395 gnd.n6394 585
R8430 gnd.n836 gnd.n835 585
R8431 gnd.n6396 gnd.n836 585
R8432 gnd.n6399 gnd.n6398 585
R8433 gnd.n6398 gnd.n6397 585
R8434 gnd.n833 gnd.n832 585
R8435 gnd.n832 gnd.n831 585
R8436 gnd.n6404 gnd.n6403 585
R8437 gnd.n6405 gnd.n6404 585
R8438 gnd.n830 gnd.n829 585
R8439 gnd.n6406 gnd.n830 585
R8440 gnd.n6409 gnd.n6408 585
R8441 gnd.n6408 gnd.n6407 585
R8442 gnd.n827 gnd.n826 585
R8443 gnd.n826 gnd.n825 585
R8444 gnd.n6414 gnd.n6413 585
R8445 gnd.n6415 gnd.n6414 585
R8446 gnd.n824 gnd.n823 585
R8447 gnd.n6416 gnd.n824 585
R8448 gnd.n6419 gnd.n6418 585
R8449 gnd.n6418 gnd.n6417 585
R8450 gnd.n821 gnd.n820 585
R8451 gnd.n820 gnd.n819 585
R8452 gnd.n6424 gnd.n6423 585
R8453 gnd.n6425 gnd.n6424 585
R8454 gnd.n818 gnd.n817 585
R8455 gnd.n6426 gnd.n818 585
R8456 gnd.n6429 gnd.n6428 585
R8457 gnd.n6428 gnd.n6427 585
R8458 gnd.n815 gnd.n814 585
R8459 gnd.n814 gnd.n813 585
R8460 gnd.n6434 gnd.n6433 585
R8461 gnd.n6435 gnd.n6434 585
R8462 gnd.n812 gnd.n811 585
R8463 gnd.n6436 gnd.n812 585
R8464 gnd.n6439 gnd.n6438 585
R8465 gnd.n6438 gnd.n6437 585
R8466 gnd.n809 gnd.n808 585
R8467 gnd.n808 gnd.n807 585
R8468 gnd.n6444 gnd.n6443 585
R8469 gnd.n6445 gnd.n6444 585
R8470 gnd.n806 gnd.n805 585
R8471 gnd.n6446 gnd.n806 585
R8472 gnd.n6449 gnd.n6448 585
R8473 gnd.n6448 gnd.n6447 585
R8474 gnd.n803 gnd.n802 585
R8475 gnd.n802 gnd.n801 585
R8476 gnd.n6454 gnd.n6453 585
R8477 gnd.n6455 gnd.n6454 585
R8478 gnd.n800 gnd.n799 585
R8479 gnd.n6456 gnd.n800 585
R8480 gnd.n6459 gnd.n6458 585
R8481 gnd.n6458 gnd.n6457 585
R8482 gnd.n797 gnd.n796 585
R8483 gnd.n796 gnd.n795 585
R8484 gnd.n6464 gnd.n6463 585
R8485 gnd.n6465 gnd.n6464 585
R8486 gnd.n794 gnd.n793 585
R8487 gnd.n6466 gnd.n794 585
R8488 gnd.n6469 gnd.n6468 585
R8489 gnd.n6468 gnd.n6467 585
R8490 gnd.n791 gnd.n790 585
R8491 gnd.n790 gnd.n789 585
R8492 gnd.n6474 gnd.n6473 585
R8493 gnd.n6475 gnd.n6474 585
R8494 gnd.n788 gnd.n787 585
R8495 gnd.n6476 gnd.n788 585
R8496 gnd.n6479 gnd.n6478 585
R8497 gnd.n6478 gnd.n6477 585
R8498 gnd.n785 gnd.n784 585
R8499 gnd.n784 gnd.n783 585
R8500 gnd.n6484 gnd.n6483 585
R8501 gnd.n6485 gnd.n6484 585
R8502 gnd.n782 gnd.n781 585
R8503 gnd.n6486 gnd.n782 585
R8504 gnd.n6489 gnd.n6488 585
R8505 gnd.n6488 gnd.n6487 585
R8506 gnd.n779 gnd.n778 585
R8507 gnd.n778 gnd.n777 585
R8508 gnd.n6494 gnd.n6493 585
R8509 gnd.n6495 gnd.n6494 585
R8510 gnd.n776 gnd.n775 585
R8511 gnd.n6496 gnd.n776 585
R8512 gnd.n6499 gnd.n6498 585
R8513 gnd.n6498 gnd.n6497 585
R8514 gnd.n773 gnd.n772 585
R8515 gnd.n772 gnd.n771 585
R8516 gnd.n6504 gnd.n6503 585
R8517 gnd.n6505 gnd.n6504 585
R8518 gnd.n770 gnd.n769 585
R8519 gnd.n6506 gnd.n770 585
R8520 gnd.n6509 gnd.n6508 585
R8521 gnd.n6508 gnd.n6507 585
R8522 gnd.n767 gnd.n766 585
R8523 gnd.n766 gnd.n765 585
R8524 gnd.n6514 gnd.n6513 585
R8525 gnd.n6515 gnd.n6514 585
R8526 gnd.n764 gnd.n763 585
R8527 gnd.n6516 gnd.n764 585
R8528 gnd.n6519 gnd.n6518 585
R8529 gnd.n6518 gnd.n6517 585
R8530 gnd.n761 gnd.n760 585
R8531 gnd.n760 gnd.n759 585
R8532 gnd.n6524 gnd.n6523 585
R8533 gnd.n6525 gnd.n6524 585
R8534 gnd.n758 gnd.n757 585
R8535 gnd.n6526 gnd.n758 585
R8536 gnd.n6529 gnd.n6528 585
R8537 gnd.n6528 gnd.n6527 585
R8538 gnd.n755 gnd.n754 585
R8539 gnd.n754 gnd.n753 585
R8540 gnd.n6534 gnd.n6533 585
R8541 gnd.n6535 gnd.n6534 585
R8542 gnd.n752 gnd.n751 585
R8543 gnd.n6536 gnd.n752 585
R8544 gnd.n6539 gnd.n6538 585
R8545 gnd.n6538 gnd.n6537 585
R8546 gnd.n749 gnd.n748 585
R8547 gnd.n748 gnd.n747 585
R8548 gnd.n6544 gnd.n6543 585
R8549 gnd.n6545 gnd.n6544 585
R8550 gnd.n746 gnd.n745 585
R8551 gnd.n6546 gnd.n746 585
R8552 gnd.n6549 gnd.n6548 585
R8553 gnd.n6548 gnd.n6547 585
R8554 gnd.n743 gnd.n742 585
R8555 gnd.n742 gnd.n741 585
R8556 gnd.n6554 gnd.n6553 585
R8557 gnd.n6555 gnd.n6554 585
R8558 gnd.n740 gnd.n739 585
R8559 gnd.n6556 gnd.n740 585
R8560 gnd.n6559 gnd.n6558 585
R8561 gnd.n6558 gnd.n6557 585
R8562 gnd.n737 gnd.n736 585
R8563 gnd.n736 gnd.n735 585
R8564 gnd.n6565 gnd.n6564 585
R8565 gnd.n6566 gnd.n6565 585
R8566 gnd.n734 gnd.n733 585
R8567 gnd.n6567 gnd.n734 585
R8568 gnd.n6570 gnd.n6569 585
R8569 gnd.n6569 gnd.n6568 585
R8570 gnd.n6571 gnd.n731 585
R8571 gnd.n731 gnd.n730 585
R8572 gnd.n606 gnd.n605 585
R8573 gnd.n6779 gnd.n605 585
R8574 gnd.n6782 gnd.n6781 585
R8575 gnd.n6781 gnd.n6780 585
R8576 gnd.n609 gnd.n608 585
R8577 gnd.n6777 gnd.n609 585
R8578 gnd.n6775 gnd.n6774 585
R8579 gnd.n6776 gnd.n6775 585
R8580 gnd.n612 gnd.n611 585
R8581 gnd.n611 gnd.n610 585
R8582 gnd.n6770 gnd.n6769 585
R8583 gnd.n6769 gnd.n6768 585
R8584 gnd.n615 gnd.n614 585
R8585 gnd.n6767 gnd.n615 585
R8586 gnd.n6765 gnd.n6764 585
R8587 gnd.n6766 gnd.n6765 585
R8588 gnd.n618 gnd.n617 585
R8589 gnd.n617 gnd.n616 585
R8590 gnd.n6760 gnd.n6759 585
R8591 gnd.n6759 gnd.n6758 585
R8592 gnd.n621 gnd.n620 585
R8593 gnd.n6757 gnd.n621 585
R8594 gnd.n6755 gnd.n6754 585
R8595 gnd.n6756 gnd.n6755 585
R8596 gnd.n624 gnd.n623 585
R8597 gnd.n623 gnd.n622 585
R8598 gnd.n6750 gnd.n6749 585
R8599 gnd.n6749 gnd.n6748 585
R8600 gnd.n627 gnd.n626 585
R8601 gnd.n6747 gnd.n627 585
R8602 gnd.n6745 gnd.n6744 585
R8603 gnd.n6746 gnd.n6745 585
R8604 gnd.n630 gnd.n629 585
R8605 gnd.n629 gnd.n628 585
R8606 gnd.n6740 gnd.n6739 585
R8607 gnd.n6739 gnd.n6738 585
R8608 gnd.n633 gnd.n632 585
R8609 gnd.n6737 gnd.n633 585
R8610 gnd.n6735 gnd.n6734 585
R8611 gnd.n6736 gnd.n6735 585
R8612 gnd.n636 gnd.n635 585
R8613 gnd.n635 gnd.n634 585
R8614 gnd.n6730 gnd.n6729 585
R8615 gnd.n6729 gnd.n6728 585
R8616 gnd.n639 gnd.n638 585
R8617 gnd.n6727 gnd.n639 585
R8618 gnd.n6725 gnd.n6724 585
R8619 gnd.n6726 gnd.n6725 585
R8620 gnd.n642 gnd.n641 585
R8621 gnd.n641 gnd.n640 585
R8622 gnd.n6720 gnd.n6719 585
R8623 gnd.n6719 gnd.n6718 585
R8624 gnd.n645 gnd.n644 585
R8625 gnd.n6717 gnd.n645 585
R8626 gnd.n6715 gnd.n6714 585
R8627 gnd.n6716 gnd.n6715 585
R8628 gnd.n648 gnd.n647 585
R8629 gnd.n647 gnd.n646 585
R8630 gnd.n6710 gnd.n6709 585
R8631 gnd.n6709 gnd.n6708 585
R8632 gnd.n651 gnd.n650 585
R8633 gnd.n6707 gnd.n651 585
R8634 gnd.n6705 gnd.n6704 585
R8635 gnd.n6706 gnd.n6705 585
R8636 gnd.n654 gnd.n653 585
R8637 gnd.n653 gnd.n652 585
R8638 gnd.n6700 gnd.n6699 585
R8639 gnd.n6699 gnd.n6698 585
R8640 gnd.n657 gnd.n656 585
R8641 gnd.n6697 gnd.n657 585
R8642 gnd.n6695 gnd.n6694 585
R8643 gnd.n6696 gnd.n6695 585
R8644 gnd.n660 gnd.n659 585
R8645 gnd.n659 gnd.n658 585
R8646 gnd.n6690 gnd.n6689 585
R8647 gnd.n6689 gnd.n6688 585
R8648 gnd.n663 gnd.n662 585
R8649 gnd.n6687 gnd.n663 585
R8650 gnd.n6685 gnd.n6684 585
R8651 gnd.n6686 gnd.n6685 585
R8652 gnd.n666 gnd.n665 585
R8653 gnd.n665 gnd.n664 585
R8654 gnd.n6680 gnd.n6679 585
R8655 gnd.n6679 gnd.n6678 585
R8656 gnd.n669 gnd.n668 585
R8657 gnd.n6677 gnd.n669 585
R8658 gnd.n6675 gnd.n6674 585
R8659 gnd.n6676 gnd.n6675 585
R8660 gnd.n672 gnd.n671 585
R8661 gnd.n671 gnd.n670 585
R8662 gnd.n6670 gnd.n6669 585
R8663 gnd.n6669 gnd.n6668 585
R8664 gnd.n675 gnd.n674 585
R8665 gnd.n6667 gnd.n675 585
R8666 gnd.n6665 gnd.n6664 585
R8667 gnd.n6666 gnd.n6665 585
R8668 gnd.n678 gnd.n677 585
R8669 gnd.n677 gnd.n676 585
R8670 gnd.n6660 gnd.n6659 585
R8671 gnd.n6659 gnd.n6658 585
R8672 gnd.n681 gnd.n680 585
R8673 gnd.n6657 gnd.n681 585
R8674 gnd.n6655 gnd.n6654 585
R8675 gnd.n6656 gnd.n6655 585
R8676 gnd.n684 gnd.n683 585
R8677 gnd.n683 gnd.n682 585
R8678 gnd.n6650 gnd.n6649 585
R8679 gnd.n6649 gnd.n6648 585
R8680 gnd.n687 gnd.n686 585
R8681 gnd.n6647 gnd.n687 585
R8682 gnd.n6645 gnd.n6644 585
R8683 gnd.n6646 gnd.n6645 585
R8684 gnd.n690 gnd.n689 585
R8685 gnd.n689 gnd.n688 585
R8686 gnd.n6640 gnd.n6639 585
R8687 gnd.n6639 gnd.n6638 585
R8688 gnd.n693 gnd.n692 585
R8689 gnd.n6637 gnd.n693 585
R8690 gnd.n6635 gnd.n6634 585
R8691 gnd.n6636 gnd.n6635 585
R8692 gnd.n696 gnd.n695 585
R8693 gnd.n695 gnd.n694 585
R8694 gnd.n6630 gnd.n6629 585
R8695 gnd.n6629 gnd.n6628 585
R8696 gnd.n699 gnd.n698 585
R8697 gnd.n6627 gnd.n699 585
R8698 gnd.n6625 gnd.n6624 585
R8699 gnd.n6626 gnd.n6625 585
R8700 gnd.n702 gnd.n701 585
R8701 gnd.n701 gnd.n700 585
R8702 gnd.n6620 gnd.n6619 585
R8703 gnd.n6619 gnd.n6618 585
R8704 gnd.n705 gnd.n704 585
R8705 gnd.n6617 gnd.n705 585
R8706 gnd.n6615 gnd.n6614 585
R8707 gnd.n6616 gnd.n6615 585
R8708 gnd.n708 gnd.n707 585
R8709 gnd.n707 gnd.n706 585
R8710 gnd.n6610 gnd.n6609 585
R8711 gnd.n6609 gnd.n6608 585
R8712 gnd.n711 gnd.n710 585
R8713 gnd.n6607 gnd.n711 585
R8714 gnd.n6605 gnd.n6604 585
R8715 gnd.n6606 gnd.n6605 585
R8716 gnd.n714 gnd.n713 585
R8717 gnd.n713 gnd.n712 585
R8718 gnd.n6600 gnd.n6599 585
R8719 gnd.n6599 gnd.n6598 585
R8720 gnd.n717 gnd.n716 585
R8721 gnd.n6597 gnd.n717 585
R8722 gnd.n6595 gnd.n6594 585
R8723 gnd.n6596 gnd.n6595 585
R8724 gnd.n720 gnd.n719 585
R8725 gnd.n719 gnd.n718 585
R8726 gnd.n6590 gnd.n6589 585
R8727 gnd.n6589 gnd.n6588 585
R8728 gnd.n723 gnd.n722 585
R8729 gnd.n6587 gnd.n723 585
R8730 gnd.n6585 gnd.n6584 585
R8731 gnd.n6586 gnd.n6585 585
R8732 gnd.n726 gnd.n725 585
R8733 gnd.n725 gnd.n724 585
R8734 gnd.n6580 gnd.n6579 585
R8735 gnd.n6579 gnd.n6578 585
R8736 gnd.n729 gnd.n728 585
R8737 gnd.n6577 gnd.n729 585
R8738 gnd.n6575 gnd.n6574 585
R8739 gnd.n6576 gnd.n6575 585
R8740 gnd.n6057 gnd.n1095 585
R8741 gnd.n4774 gnd.n1095 585
R8742 gnd.n6059 gnd.n6058 585
R8743 gnd.n6060 gnd.n6059 585
R8744 gnd.n1079 gnd.n1078 585
R8745 gnd.n4782 gnd.n1079 585
R8746 gnd.n6068 gnd.n6067 585
R8747 gnd.n6067 gnd.n6066 585
R8748 gnd.n6069 gnd.n1073 585
R8749 gnd.n4443 gnd.n1073 585
R8750 gnd.n6071 gnd.n6070 585
R8751 gnd.n6072 gnd.n6071 585
R8752 gnd.n1074 gnd.n1072 585
R8753 gnd.n4434 gnd.n1072 585
R8754 gnd.n4404 gnd.n1059 585
R8755 gnd.n6078 gnd.n1059 585
R8756 gnd.n4718 gnd.n4449 585
R8757 gnd.n4556 gnd.n4555 585
R8758 gnd.n4725 gnd.n4551 585
R8759 gnd.n4726 gnd.n4549 585
R8760 gnd.n4548 gnd.n4541 585
R8761 gnd.n4733 gnd.n4540 585
R8762 gnd.n4734 gnd.n4539 585
R8763 gnd.n4537 gnd.n4529 585
R8764 gnd.n4741 gnd.n4528 585
R8765 gnd.n4742 gnd.n4526 585
R8766 gnd.n4525 gnd.n4518 585
R8767 gnd.n4749 gnd.n4517 585
R8768 gnd.n4750 gnd.n4516 585
R8769 gnd.n4514 gnd.n4507 585
R8770 gnd.n4757 gnd.n4506 585
R8771 gnd.n4758 gnd.n4504 585
R8772 gnd.n4503 gnd.n4498 585
R8773 gnd.n4501 gnd.n4500 585
R8774 gnd.n4499 gnd.n1098 585
R8775 gnd.n4499 gnd.n1960 585
R8776 gnd.n4776 gnd.n4775 585
R8777 gnd.n4775 gnd.n4774 585
R8778 gnd.n1998 gnd.n1093 585
R8779 gnd.n6060 gnd.n1093 585
R8780 gnd.n4781 gnd.n4780 585
R8781 gnd.n4782 gnd.n4781 585
R8782 gnd.n1997 gnd.n1082 585
R8783 gnd.n6066 gnd.n1082 585
R8784 gnd.n4445 gnd.n4444 585
R8785 gnd.n4444 gnd.n4443 585
R8786 gnd.n2000 gnd.n1070 585
R8787 gnd.n6072 gnd.n1070 585
R8788 gnd.n4433 gnd.n4432 585
R8789 gnd.n4434 gnd.n4433 585
R8790 gnd.n2005 gnd.n1058 585
R8791 gnd.n6078 gnd.n1058 585
R8792 gnd.n7457 gnd.n129 585
R8793 gnd.n7553 gnd.n129 585
R8794 gnd.n7458 gnd.n7395 585
R8795 gnd.n7395 gnd.n126 585
R8796 gnd.n7459 gnd.n207 585
R8797 gnd.n7473 gnd.n207 585
R8798 gnd.n219 gnd.n217 585
R8799 gnd.n217 gnd.n206 585
R8800 gnd.n7464 gnd.n7463 585
R8801 gnd.n7465 gnd.n7464 585
R8802 gnd.n218 gnd.n216 585
R8803 gnd.n216 gnd.n213 585
R8804 gnd.n7391 gnd.n7390 585
R8805 gnd.n7390 gnd.n7389 585
R8806 gnd.n222 gnd.n221 585
R8807 gnd.n232 gnd.n222 585
R8808 gnd.n7380 gnd.n7379 585
R8809 gnd.n7381 gnd.n7380 585
R8810 gnd.n234 gnd.n233 585
R8811 gnd.n233 gnd.n229 585
R8812 gnd.n7375 gnd.n7374 585
R8813 gnd.n7374 gnd.n7373 585
R8814 gnd.n237 gnd.n236 585
R8815 gnd.n238 gnd.n237 585
R8816 gnd.n7364 gnd.n7363 585
R8817 gnd.n7365 gnd.n7364 585
R8818 gnd.n248 gnd.n247 585
R8819 gnd.n253 gnd.n247 585
R8820 gnd.n7359 gnd.n7358 585
R8821 gnd.n7358 gnd.n7357 585
R8822 gnd.n251 gnd.n250 585
R8823 gnd.n262 gnd.n251 585
R8824 gnd.n7348 gnd.n7347 585
R8825 gnd.n7349 gnd.n7348 585
R8826 gnd.n264 gnd.n263 585
R8827 gnd.n263 gnd.n259 585
R8828 gnd.n7343 gnd.n7342 585
R8829 gnd.n7342 gnd.n7341 585
R8830 gnd.n267 gnd.n266 585
R8831 gnd.n268 gnd.n267 585
R8832 gnd.n7332 gnd.n7331 585
R8833 gnd.n7333 gnd.n7332 585
R8834 gnd.n278 gnd.n277 585
R8835 gnd.n283 gnd.n277 585
R8836 gnd.n7327 gnd.n7326 585
R8837 gnd.n7326 gnd.n7325 585
R8838 gnd.n281 gnd.n280 585
R8839 gnd.n292 gnd.n281 585
R8840 gnd.n7316 gnd.n7315 585
R8841 gnd.n7317 gnd.n7316 585
R8842 gnd.n294 gnd.n293 585
R8843 gnd.n293 gnd.n289 585
R8844 gnd.n7311 gnd.n7310 585
R8845 gnd.n7310 gnd.n7309 585
R8846 gnd.n297 gnd.n296 585
R8847 gnd.n298 gnd.n297 585
R8848 gnd.n7300 gnd.n7299 585
R8849 gnd.n7301 gnd.n7300 585
R8850 gnd.n308 gnd.n307 585
R8851 gnd.n313 gnd.n307 585
R8852 gnd.n7295 gnd.n7294 585
R8853 gnd.n7294 gnd.n7293 585
R8854 gnd.n311 gnd.n310 585
R8855 gnd.n322 gnd.n311 585
R8856 gnd.n7284 gnd.n7283 585
R8857 gnd.n7285 gnd.n7284 585
R8858 gnd.n324 gnd.n323 585
R8859 gnd.n323 gnd.n319 585
R8860 gnd.n7279 gnd.n7278 585
R8861 gnd.n7278 gnd.n7277 585
R8862 gnd.n328 gnd.n327 585
R8863 gnd.n329 gnd.n328 585
R8864 gnd.n7268 gnd.n7267 585
R8865 gnd.n7269 gnd.n7268 585
R8866 gnd.n341 gnd.n340 585
R8867 gnd.n340 gnd.n337 585
R8868 gnd.n7263 gnd.n7262 585
R8869 gnd.n7262 gnd.n7261 585
R8870 gnd.n344 gnd.n343 585
R8871 gnd.n355 gnd.n344 585
R8872 gnd.n7252 gnd.n7251 585
R8873 gnd.n7253 gnd.n7252 585
R8874 gnd.n357 gnd.n356 585
R8875 gnd.n356 gnd.n352 585
R8876 gnd.n7247 gnd.n7246 585
R8877 gnd.n7246 gnd.n7245 585
R8878 gnd.n360 gnd.n359 585
R8879 gnd.n361 gnd.n360 585
R8880 gnd.n7236 gnd.n7235 585
R8881 gnd.n7237 gnd.n7236 585
R8882 gnd.n373 gnd.n372 585
R8883 gnd.n372 gnd.n369 585
R8884 gnd.n7231 gnd.n7230 585
R8885 gnd.n7230 gnd.n7229 585
R8886 gnd.n376 gnd.n375 585
R8887 gnd.n387 gnd.n376 585
R8888 gnd.n7220 gnd.n7219 585
R8889 gnd.n7221 gnd.n7220 585
R8890 gnd.n389 gnd.n388 585
R8891 gnd.n388 gnd.n384 585
R8892 gnd.n7215 gnd.n7214 585
R8893 gnd.n7214 gnd.n7213 585
R8894 gnd.n392 gnd.n391 585
R8895 gnd.n393 gnd.n392 585
R8896 gnd.n7204 gnd.n7203 585
R8897 gnd.n7205 gnd.n7204 585
R8898 gnd.n405 gnd.n404 585
R8899 gnd.n404 gnd.n401 585
R8900 gnd.n7199 gnd.n7198 585
R8901 gnd.n7198 gnd.n7197 585
R8902 gnd.n408 gnd.n407 585
R8903 gnd.n6955 gnd.n408 585
R8904 gnd.n7188 gnd.n7187 585
R8905 gnd.n7189 gnd.n7188 585
R8906 gnd.n421 gnd.n420 585
R8907 gnd.n6818 gnd.n420 585
R8908 gnd.n7183 gnd.n7182 585
R8909 gnd.n7182 gnd.n7181 585
R8910 gnd.n424 gnd.n423 585
R8911 gnd.n6814 gnd.n424 585
R8912 gnd.n7172 gnd.n7171 585
R8913 gnd.n7173 gnd.n7172 585
R8914 gnd.n439 gnd.n438 585
R8915 gnd.n7022 gnd.n438 585
R8916 gnd.n7167 gnd.n7166 585
R8917 gnd.n7166 gnd.n7165 585
R8918 gnd.n442 gnd.n441 585
R8919 gnd.n6800 gnd.n442 585
R8920 gnd.n7156 gnd.n7155 585
R8921 gnd.n7157 gnd.n7156 585
R8922 gnd.n7152 gnd.n454 585
R8923 gnd.n7151 gnd.n456 585
R8924 gnd.n526 gnd.n457 585
R8925 gnd.n7144 gnd.n463 585
R8926 gnd.n7143 gnd.n464 585
R8927 gnd.n528 gnd.n465 585
R8928 gnd.n7136 gnd.n471 585
R8929 gnd.n7135 gnd.n472 585
R8930 gnd.n531 gnd.n473 585
R8931 gnd.n7128 gnd.n479 585
R8932 gnd.n7127 gnd.n480 585
R8933 gnd.n533 gnd.n481 585
R8934 gnd.n7120 gnd.n487 585
R8935 gnd.n7119 gnd.n488 585
R8936 gnd.n536 gnd.n489 585
R8937 gnd.n7112 gnd.n495 585
R8938 gnd.n7111 gnd.n496 585
R8939 gnd.n505 gnd.n499 585
R8940 gnd.n7104 gnd.n7103 585
R8941 gnd.n7103 gnd.n7102 585
R8942 gnd.n7556 gnd.n7555 585
R8943 gnd.n7428 gnd.n124 585
R8944 gnd.n7430 gnd.n7429 585
R8945 gnd.n7426 gnd.n7425 585
R8946 gnd.n7434 gnd.n7424 585
R8947 gnd.n7435 gnd.n7422 585
R8948 gnd.n7436 gnd.n7421 585
R8949 gnd.n7419 gnd.n7417 585
R8950 gnd.n7440 gnd.n7416 585
R8951 gnd.n7441 gnd.n7414 585
R8952 gnd.n7442 gnd.n7413 585
R8953 gnd.n7411 gnd.n7409 585
R8954 gnd.n7446 gnd.n7408 585
R8955 gnd.n7447 gnd.n7406 585
R8956 gnd.n7448 gnd.n7405 585
R8957 gnd.n7403 gnd.n7401 585
R8958 gnd.n7452 gnd.n7400 585
R8959 gnd.n7453 gnd.n7398 585
R8960 gnd.n7454 gnd.n7397 585
R8961 gnd.n7397 gnd.n128 585
R8962 gnd.n7554 gnd.n120 585
R8963 gnd.n7554 gnd.n7553 585
R8964 gnd.n7560 gnd.n119 585
R8965 gnd.n126 gnd.n119 585
R8966 gnd.n7561 gnd.n118 585
R8967 gnd.n7473 gnd.n118 585
R8968 gnd.n7562 gnd.n117 585
R8969 gnd.n206 gnd.n117 585
R8970 gnd.n215 gnd.n115 585
R8971 gnd.n7465 gnd.n215 585
R8972 gnd.n7566 gnd.n114 585
R8973 gnd.n213 gnd.n114 585
R8974 gnd.n7567 gnd.n113 585
R8975 gnd.n7389 gnd.n113 585
R8976 gnd.n7568 gnd.n112 585
R8977 gnd.n232 gnd.n112 585
R8978 gnd.n231 gnd.n110 585
R8979 gnd.n7381 gnd.n231 585
R8980 gnd.n7572 gnd.n109 585
R8981 gnd.n229 gnd.n109 585
R8982 gnd.n7573 gnd.n108 585
R8983 gnd.n7373 gnd.n108 585
R8984 gnd.n7574 gnd.n107 585
R8985 gnd.n238 gnd.n107 585
R8986 gnd.n246 gnd.n105 585
R8987 gnd.n7365 gnd.n246 585
R8988 gnd.n7578 gnd.n104 585
R8989 gnd.n253 gnd.n104 585
R8990 gnd.n7579 gnd.n103 585
R8991 gnd.n7357 gnd.n103 585
R8992 gnd.n7580 gnd.n102 585
R8993 gnd.n262 gnd.n102 585
R8994 gnd.n261 gnd.n100 585
R8995 gnd.n7349 gnd.n261 585
R8996 gnd.n7584 gnd.n99 585
R8997 gnd.n259 gnd.n99 585
R8998 gnd.n7585 gnd.n98 585
R8999 gnd.n7341 gnd.n98 585
R9000 gnd.n7586 gnd.n97 585
R9001 gnd.n268 gnd.n97 585
R9002 gnd.n276 gnd.n95 585
R9003 gnd.n7333 gnd.n276 585
R9004 gnd.n7590 gnd.n94 585
R9005 gnd.n283 gnd.n94 585
R9006 gnd.n7591 gnd.n93 585
R9007 gnd.n7325 gnd.n93 585
R9008 gnd.n7592 gnd.n92 585
R9009 gnd.n292 gnd.n92 585
R9010 gnd.n291 gnd.n90 585
R9011 gnd.n7317 gnd.n291 585
R9012 gnd.n7596 gnd.n89 585
R9013 gnd.n289 gnd.n89 585
R9014 gnd.n7597 gnd.n88 585
R9015 gnd.n7309 gnd.n88 585
R9016 gnd.n7598 gnd.n87 585
R9017 gnd.n298 gnd.n87 585
R9018 gnd.n306 gnd.n85 585
R9019 gnd.n7301 gnd.n306 585
R9020 gnd.n7602 gnd.n84 585
R9021 gnd.n313 gnd.n84 585
R9022 gnd.n7603 gnd.n83 585
R9023 gnd.n7293 gnd.n83 585
R9024 gnd.n7604 gnd.n82 585
R9025 gnd.n322 gnd.n82 585
R9026 gnd.n321 gnd.n80 585
R9027 gnd.n7285 gnd.n321 585
R9028 gnd.n6978 gnd.n6977 585
R9029 gnd.n6977 gnd.n319 585
R9030 gnd.n6979 gnd.n331 585
R9031 gnd.n7277 gnd.n331 585
R9032 gnd.n6980 gnd.n6976 585
R9033 gnd.n6976 gnd.n329 585
R9034 gnd.n6974 gnd.n339 585
R9035 gnd.n7269 gnd.n339 585
R9036 gnd.n6984 gnd.n6973 585
R9037 gnd.n6973 gnd.n337 585
R9038 gnd.n6985 gnd.n346 585
R9039 gnd.n7261 gnd.n346 585
R9040 gnd.n6986 gnd.n6972 585
R9041 gnd.n6972 gnd.n355 585
R9042 gnd.n6970 gnd.n354 585
R9043 gnd.n7253 gnd.n354 585
R9044 gnd.n6990 gnd.n6969 585
R9045 gnd.n6969 gnd.n352 585
R9046 gnd.n6991 gnd.n363 585
R9047 gnd.n7245 gnd.n363 585
R9048 gnd.n6992 gnd.n6968 585
R9049 gnd.n6968 gnd.n361 585
R9050 gnd.n6966 gnd.n371 585
R9051 gnd.n7237 gnd.n371 585
R9052 gnd.n6996 gnd.n6965 585
R9053 gnd.n6965 gnd.n369 585
R9054 gnd.n6997 gnd.n378 585
R9055 gnd.n7229 gnd.n378 585
R9056 gnd.n6998 gnd.n6964 585
R9057 gnd.n6964 gnd.n387 585
R9058 gnd.n6962 gnd.n386 585
R9059 gnd.n7221 gnd.n386 585
R9060 gnd.n7002 gnd.n6961 585
R9061 gnd.n6961 gnd.n384 585
R9062 gnd.n7003 gnd.n395 585
R9063 gnd.n7213 gnd.n395 585
R9064 gnd.n7004 gnd.n6960 585
R9065 gnd.n6960 gnd.n393 585
R9066 gnd.n6958 gnd.n403 585
R9067 gnd.n7205 gnd.n403 585
R9068 gnd.n7008 gnd.n6957 585
R9069 gnd.n6957 gnd.n401 585
R9070 gnd.n7009 gnd.n410 585
R9071 gnd.n7197 gnd.n410 585
R9072 gnd.n7010 gnd.n6956 585
R9073 gnd.n6956 gnd.n6955 585
R9074 gnd.n6808 gnd.n418 585
R9075 gnd.n7189 gnd.n418 585
R9076 gnd.n7014 gnd.n6807 585
R9077 gnd.n6818 gnd.n6807 585
R9078 gnd.n7015 gnd.n427 585
R9079 gnd.n7181 gnd.n427 585
R9080 gnd.n7016 gnd.n6806 585
R9081 gnd.n6814 gnd.n6806 585
R9082 gnd.n590 gnd.n436 585
R9083 gnd.n7173 gnd.n436 585
R9084 gnd.n7021 gnd.n7020 585
R9085 gnd.n7022 gnd.n7021 585
R9086 gnd.n589 gnd.n444 585
R9087 gnd.n7165 gnd.n444 585
R9088 gnd.n6802 gnd.n6801 585
R9089 gnd.n6801 gnd.n6800 585
R9090 gnd.n592 gnd.n452 585
R9091 gnd.n7157 gnd.n452 585
R9092 gnd.n1090 gnd.n1089 585
R9093 gnd.n4774 gnd.n1090 585
R9094 gnd.n6062 gnd.n6061 585
R9095 gnd.n6061 gnd.n6060 585
R9096 gnd.n6063 gnd.n1084 585
R9097 gnd.n4782 gnd.n1084 585
R9098 gnd.n6065 gnd.n6064 585
R9099 gnd.n6066 gnd.n6065 585
R9100 gnd.n1067 gnd.n1066 585
R9101 gnd.n4443 gnd.n1067 585
R9102 gnd.n6074 gnd.n6073 585
R9103 gnd.n6073 gnd.n6072 585
R9104 gnd.n6075 gnd.n1061 585
R9105 gnd.n4434 gnd.n1061 585
R9106 gnd.n6077 gnd.n6076 585
R9107 gnd.n6078 gnd.n6077 585
R9108 gnd.n4790 gnd.n4789 585
R9109 gnd.n4792 gnd.n1990 585
R9110 gnd.n4794 gnd.n4793 585
R9111 gnd.n4795 gnd.n1983 585
R9112 gnd.n4797 gnd.n4796 585
R9113 gnd.n4799 gnd.n1981 585
R9114 gnd.n4801 gnd.n4800 585
R9115 gnd.n4802 gnd.n1976 585
R9116 gnd.n4804 gnd.n4803 585
R9117 gnd.n4806 gnd.n1974 585
R9118 gnd.n4808 gnd.n4807 585
R9119 gnd.n4809 gnd.n1969 585
R9120 gnd.n4811 gnd.n4810 585
R9121 gnd.n4813 gnd.n1967 585
R9122 gnd.n4815 gnd.n4814 585
R9123 gnd.n4816 gnd.n1962 585
R9124 gnd.n4818 gnd.n4817 585
R9125 gnd.n4820 gnd.n1961 585
R9126 gnd.n4821 gnd.n1902 585
R9127 gnd.n4824 gnd.n4823 585
R9128 gnd.n1903 gnd.n1895 585
R9129 gnd.n1930 gnd.n1896 585
R9130 gnd.n1932 gnd.n1931 585
R9131 gnd.n1934 gnd.n1933 585
R9132 gnd.n1936 gnd.n1935 585
R9133 gnd.n1938 gnd.n1937 585
R9134 gnd.n1940 gnd.n1939 585
R9135 gnd.n1942 gnd.n1941 585
R9136 gnd.n1944 gnd.n1943 585
R9137 gnd.n1946 gnd.n1945 585
R9138 gnd.n1948 gnd.n1947 585
R9139 gnd.n1950 gnd.n1949 585
R9140 gnd.n1952 gnd.n1951 585
R9141 gnd.n1954 gnd.n1953 585
R9142 gnd.n1956 gnd.n1955 585
R9143 gnd.n1957 gnd.n1913 585
R9144 gnd.n1959 gnd.n1958 585
R9145 gnd.n1960 gnd.n1959 585
R9146 gnd.n4786 gnd.n1992 585
R9147 gnd.n4774 gnd.n1992 585
R9148 gnd.n4785 gnd.n1092 585
R9149 gnd.n6060 gnd.n1092 585
R9150 gnd.n4784 gnd.n4783 585
R9151 gnd.n4783 gnd.n4782 585
R9152 gnd.n1995 gnd.n1081 585
R9153 gnd.n6066 gnd.n1081 585
R9154 gnd.n4442 gnd.n4441 585
R9155 gnd.n4443 gnd.n4442 585
R9156 gnd.n2001 gnd.n1069 585
R9157 gnd.n6072 gnd.n1069 585
R9158 gnd.n4436 gnd.n4435 585
R9159 gnd.n4435 gnd.n4434 585
R9160 gnd.n2003 gnd.n1057 585
R9161 gnd.n6078 gnd.n1057 585
R9162 gnd.n7552 gnd.n7551 585
R9163 gnd.n7553 gnd.n7552 585
R9164 gnd.n132 gnd.n130 585
R9165 gnd.n130 gnd.n126 585
R9166 gnd.n7472 gnd.n7471 585
R9167 gnd.n7473 gnd.n7472 585
R9168 gnd.n209 gnd.n208 585
R9169 gnd.n208 gnd.n206 585
R9170 gnd.n7467 gnd.n7466 585
R9171 gnd.n7466 gnd.n7465 585
R9172 gnd.n212 gnd.n211 585
R9173 gnd.n213 gnd.n212 585
R9174 gnd.n7388 gnd.n7387 585
R9175 gnd.n7389 gnd.n7388 585
R9176 gnd.n225 gnd.n224 585
R9177 gnd.n232 gnd.n224 585
R9178 gnd.n7383 gnd.n7382 585
R9179 gnd.n7382 gnd.n7381 585
R9180 gnd.n228 gnd.n227 585
R9181 gnd.n229 gnd.n228 585
R9182 gnd.n7372 gnd.n7371 585
R9183 gnd.n7373 gnd.n7372 585
R9184 gnd.n241 gnd.n240 585
R9185 gnd.n240 gnd.n238 585
R9186 gnd.n7367 gnd.n7366 585
R9187 gnd.n7366 gnd.n7365 585
R9188 gnd.n244 gnd.n243 585
R9189 gnd.n253 gnd.n244 585
R9190 gnd.n7356 gnd.n7355 585
R9191 gnd.n7357 gnd.n7356 585
R9192 gnd.n255 gnd.n254 585
R9193 gnd.n262 gnd.n254 585
R9194 gnd.n7351 gnd.n7350 585
R9195 gnd.n7350 gnd.n7349 585
R9196 gnd.n258 gnd.n257 585
R9197 gnd.n259 gnd.n258 585
R9198 gnd.n7340 gnd.n7339 585
R9199 gnd.n7341 gnd.n7340 585
R9200 gnd.n271 gnd.n270 585
R9201 gnd.n270 gnd.n268 585
R9202 gnd.n7335 gnd.n7334 585
R9203 gnd.n7334 gnd.n7333 585
R9204 gnd.n274 gnd.n273 585
R9205 gnd.n283 gnd.n274 585
R9206 gnd.n7324 gnd.n7323 585
R9207 gnd.n7325 gnd.n7324 585
R9208 gnd.n285 gnd.n284 585
R9209 gnd.n292 gnd.n284 585
R9210 gnd.n7319 gnd.n7318 585
R9211 gnd.n7318 gnd.n7317 585
R9212 gnd.n288 gnd.n287 585
R9213 gnd.n289 gnd.n288 585
R9214 gnd.n7308 gnd.n7307 585
R9215 gnd.n7309 gnd.n7308 585
R9216 gnd.n301 gnd.n300 585
R9217 gnd.n300 gnd.n298 585
R9218 gnd.n7303 gnd.n7302 585
R9219 gnd.n7302 gnd.n7301 585
R9220 gnd.n304 gnd.n303 585
R9221 gnd.n313 gnd.n304 585
R9222 gnd.n7292 gnd.n7291 585
R9223 gnd.n7293 gnd.n7292 585
R9224 gnd.n315 gnd.n314 585
R9225 gnd.n322 gnd.n314 585
R9226 gnd.n7287 gnd.n7286 585
R9227 gnd.n7286 gnd.n7285 585
R9228 gnd.n318 gnd.n317 585
R9229 gnd.n319 gnd.n318 585
R9230 gnd.n7276 gnd.n7275 585
R9231 gnd.n7277 gnd.n7276 585
R9232 gnd.n333 gnd.n332 585
R9233 gnd.n332 gnd.n329 585
R9234 gnd.n7271 gnd.n7270 585
R9235 gnd.n7270 gnd.n7269 585
R9236 gnd.n336 gnd.n335 585
R9237 gnd.n337 gnd.n336 585
R9238 gnd.n7260 gnd.n7259 585
R9239 gnd.n7261 gnd.n7260 585
R9240 gnd.n348 gnd.n347 585
R9241 gnd.n355 gnd.n347 585
R9242 gnd.n7255 gnd.n7254 585
R9243 gnd.n7254 gnd.n7253 585
R9244 gnd.n351 gnd.n350 585
R9245 gnd.n352 gnd.n351 585
R9246 gnd.n7244 gnd.n7243 585
R9247 gnd.n7245 gnd.n7244 585
R9248 gnd.n365 gnd.n364 585
R9249 gnd.n364 gnd.n361 585
R9250 gnd.n7239 gnd.n7238 585
R9251 gnd.n7238 gnd.n7237 585
R9252 gnd.n368 gnd.n367 585
R9253 gnd.n369 gnd.n368 585
R9254 gnd.n7228 gnd.n7227 585
R9255 gnd.n7229 gnd.n7228 585
R9256 gnd.n380 gnd.n379 585
R9257 gnd.n387 gnd.n379 585
R9258 gnd.n7223 gnd.n7222 585
R9259 gnd.n7222 gnd.n7221 585
R9260 gnd.n383 gnd.n382 585
R9261 gnd.n384 gnd.n383 585
R9262 gnd.n7212 gnd.n7211 585
R9263 gnd.n7213 gnd.n7212 585
R9264 gnd.n397 gnd.n396 585
R9265 gnd.n396 gnd.n393 585
R9266 gnd.n7207 gnd.n7206 585
R9267 gnd.n7206 gnd.n7205 585
R9268 gnd.n400 gnd.n399 585
R9269 gnd.n401 gnd.n400 585
R9270 gnd.n7196 gnd.n7195 585
R9271 gnd.n7197 gnd.n7196 585
R9272 gnd.n412 gnd.n411 585
R9273 gnd.n6955 gnd.n411 585
R9274 gnd.n7191 gnd.n7190 585
R9275 gnd.n7190 gnd.n7189 585
R9276 gnd.n415 gnd.n414 585
R9277 gnd.n6818 gnd.n415 585
R9278 gnd.n7180 gnd.n7179 585
R9279 gnd.n7181 gnd.n7180 585
R9280 gnd.n430 gnd.n429 585
R9281 gnd.n6814 gnd.n429 585
R9282 gnd.n7175 gnd.n7174 585
R9283 gnd.n7174 gnd.n7173 585
R9284 gnd.n433 gnd.n432 585
R9285 gnd.n7022 gnd.n433 585
R9286 gnd.n7164 gnd.n7163 585
R9287 gnd.n7165 gnd.n7164 585
R9288 gnd.n447 gnd.n446 585
R9289 gnd.n6800 gnd.n446 585
R9290 gnd.n7159 gnd.n7158 585
R9291 gnd.n7158 gnd.n7157 585
R9292 gnd.n540 gnd.n449 585
R9293 gnd.n7100 gnd.n7099 585
R9294 gnd.n7098 gnd.n539 585
R9295 gnd.n7102 gnd.n539 585
R9296 gnd.n7097 gnd.n7096 585
R9297 gnd.n7095 gnd.n7094 585
R9298 gnd.n7093 gnd.n7092 585
R9299 gnd.n7091 gnd.n7090 585
R9300 gnd.n7089 gnd.n7088 585
R9301 gnd.n7087 gnd.n7086 585
R9302 gnd.n7085 gnd.n7084 585
R9303 gnd.n7083 gnd.n7082 585
R9304 gnd.n7081 gnd.n7080 585
R9305 gnd.n7079 gnd.n7078 585
R9306 gnd.n7077 gnd.n7076 585
R9307 gnd.n7075 gnd.n7074 585
R9308 gnd.n7073 gnd.n7072 585
R9309 gnd.n7070 gnd.n7069 585
R9310 gnd.n7068 gnd.n7067 585
R9311 gnd.n7066 gnd.n7065 585
R9312 gnd.n7064 gnd.n7063 585
R9313 gnd.n7062 gnd.n7061 585
R9314 gnd.n7060 gnd.n7059 585
R9315 gnd.n7058 gnd.n7057 585
R9316 gnd.n7056 gnd.n7055 585
R9317 gnd.n7054 gnd.n7053 585
R9318 gnd.n7052 gnd.n7051 585
R9319 gnd.n7050 gnd.n7049 585
R9320 gnd.n7048 gnd.n7047 585
R9321 gnd.n7046 gnd.n7045 585
R9322 gnd.n7044 gnd.n7043 585
R9323 gnd.n7042 gnd.n7041 585
R9324 gnd.n7040 gnd.n7039 585
R9325 gnd.n7038 gnd.n7037 585
R9326 gnd.n7036 gnd.n7035 585
R9327 gnd.n7034 gnd.n579 585
R9328 gnd.n583 gnd.n580 585
R9329 gnd.n7030 gnd.n7029 585
R9330 gnd.n200 gnd.n199 585
R9331 gnd.n7481 gnd.n195 585
R9332 gnd.n7483 gnd.n7482 585
R9333 gnd.n7485 gnd.n193 585
R9334 gnd.n7487 gnd.n7486 585
R9335 gnd.n7488 gnd.n188 585
R9336 gnd.n7490 gnd.n7489 585
R9337 gnd.n7492 gnd.n186 585
R9338 gnd.n7494 gnd.n7493 585
R9339 gnd.n7495 gnd.n181 585
R9340 gnd.n7497 gnd.n7496 585
R9341 gnd.n7499 gnd.n179 585
R9342 gnd.n7501 gnd.n7500 585
R9343 gnd.n7502 gnd.n174 585
R9344 gnd.n7504 gnd.n7503 585
R9345 gnd.n7506 gnd.n172 585
R9346 gnd.n7508 gnd.n7507 585
R9347 gnd.n7509 gnd.n167 585
R9348 gnd.n7511 gnd.n7510 585
R9349 gnd.n7513 gnd.n165 585
R9350 gnd.n7515 gnd.n7514 585
R9351 gnd.n7519 gnd.n160 585
R9352 gnd.n7521 gnd.n7520 585
R9353 gnd.n7523 gnd.n158 585
R9354 gnd.n7525 gnd.n7524 585
R9355 gnd.n7526 gnd.n153 585
R9356 gnd.n7528 gnd.n7527 585
R9357 gnd.n7530 gnd.n151 585
R9358 gnd.n7532 gnd.n7531 585
R9359 gnd.n7533 gnd.n146 585
R9360 gnd.n7535 gnd.n7534 585
R9361 gnd.n7537 gnd.n144 585
R9362 gnd.n7539 gnd.n7538 585
R9363 gnd.n7540 gnd.n139 585
R9364 gnd.n7542 gnd.n7541 585
R9365 gnd.n7544 gnd.n137 585
R9366 gnd.n7546 gnd.n7545 585
R9367 gnd.n7547 gnd.n135 585
R9368 gnd.n7548 gnd.n131 585
R9369 gnd.n131 gnd.n128 585
R9370 gnd.n7477 gnd.n127 585
R9371 gnd.n7553 gnd.n127 585
R9372 gnd.n7476 gnd.n7475 585
R9373 gnd.n7475 gnd.n126 585
R9374 gnd.n7474 gnd.n204 585
R9375 gnd.n7474 gnd.n7473 585
R9376 gnd.n6876 gnd.n205 585
R9377 gnd.n206 gnd.n205 585
R9378 gnd.n6877 gnd.n214 585
R9379 gnd.n7465 gnd.n214 585
R9380 gnd.n6879 gnd.n6878 585
R9381 gnd.n6878 gnd.n213 585
R9382 gnd.n6880 gnd.n223 585
R9383 gnd.n7389 gnd.n223 585
R9384 gnd.n6882 gnd.n6881 585
R9385 gnd.n6881 gnd.n232 585
R9386 gnd.n6883 gnd.n230 585
R9387 gnd.n7381 gnd.n230 585
R9388 gnd.n6885 gnd.n6884 585
R9389 gnd.n6884 gnd.n229 585
R9390 gnd.n6886 gnd.n239 585
R9391 gnd.n7373 gnd.n239 585
R9392 gnd.n6888 gnd.n6887 585
R9393 gnd.n6887 gnd.n238 585
R9394 gnd.n6889 gnd.n245 585
R9395 gnd.n7365 gnd.n245 585
R9396 gnd.n6891 gnd.n6890 585
R9397 gnd.n6890 gnd.n253 585
R9398 gnd.n6892 gnd.n252 585
R9399 gnd.n7357 gnd.n252 585
R9400 gnd.n6894 gnd.n6893 585
R9401 gnd.n6893 gnd.n262 585
R9402 gnd.n6895 gnd.n260 585
R9403 gnd.n7349 gnd.n260 585
R9404 gnd.n6897 gnd.n6896 585
R9405 gnd.n6896 gnd.n259 585
R9406 gnd.n6898 gnd.n269 585
R9407 gnd.n7341 gnd.n269 585
R9408 gnd.n6900 gnd.n6899 585
R9409 gnd.n6899 gnd.n268 585
R9410 gnd.n6901 gnd.n275 585
R9411 gnd.n7333 gnd.n275 585
R9412 gnd.n6903 gnd.n6902 585
R9413 gnd.n6902 gnd.n283 585
R9414 gnd.n6904 gnd.n282 585
R9415 gnd.n7325 gnd.n282 585
R9416 gnd.n6906 gnd.n6905 585
R9417 gnd.n6905 gnd.n292 585
R9418 gnd.n6907 gnd.n290 585
R9419 gnd.n7317 gnd.n290 585
R9420 gnd.n6909 gnd.n6908 585
R9421 gnd.n6908 gnd.n289 585
R9422 gnd.n6910 gnd.n299 585
R9423 gnd.n7309 gnd.n299 585
R9424 gnd.n6912 gnd.n6911 585
R9425 gnd.n6911 gnd.n298 585
R9426 gnd.n6913 gnd.n305 585
R9427 gnd.n7301 gnd.n305 585
R9428 gnd.n6915 gnd.n6914 585
R9429 gnd.n6914 gnd.n313 585
R9430 gnd.n6916 gnd.n312 585
R9431 gnd.n7293 gnd.n312 585
R9432 gnd.n6918 gnd.n6917 585
R9433 gnd.n6917 gnd.n322 585
R9434 gnd.n6919 gnd.n320 585
R9435 gnd.n7285 gnd.n320 585
R9436 gnd.n6921 gnd.n6920 585
R9437 gnd.n6920 gnd.n319 585
R9438 gnd.n6922 gnd.n330 585
R9439 gnd.n7277 gnd.n330 585
R9440 gnd.n6924 gnd.n6923 585
R9441 gnd.n6923 gnd.n329 585
R9442 gnd.n6925 gnd.n338 585
R9443 gnd.n7269 gnd.n338 585
R9444 gnd.n6927 gnd.n6926 585
R9445 gnd.n6926 gnd.n337 585
R9446 gnd.n6928 gnd.n345 585
R9447 gnd.n7261 gnd.n345 585
R9448 gnd.n6930 gnd.n6929 585
R9449 gnd.n6929 gnd.n355 585
R9450 gnd.n6931 gnd.n353 585
R9451 gnd.n7253 gnd.n353 585
R9452 gnd.n6933 gnd.n6932 585
R9453 gnd.n6932 gnd.n352 585
R9454 gnd.n6934 gnd.n362 585
R9455 gnd.n7245 gnd.n362 585
R9456 gnd.n6936 gnd.n6935 585
R9457 gnd.n6935 gnd.n361 585
R9458 gnd.n6937 gnd.n370 585
R9459 gnd.n7237 gnd.n370 585
R9460 gnd.n6939 gnd.n6938 585
R9461 gnd.n6938 gnd.n369 585
R9462 gnd.n6940 gnd.n377 585
R9463 gnd.n7229 gnd.n377 585
R9464 gnd.n6942 gnd.n6941 585
R9465 gnd.n6941 gnd.n387 585
R9466 gnd.n6943 gnd.n385 585
R9467 gnd.n7221 gnd.n385 585
R9468 gnd.n6945 gnd.n6944 585
R9469 gnd.n6944 gnd.n384 585
R9470 gnd.n6946 gnd.n394 585
R9471 gnd.n7213 gnd.n394 585
R9472 gnd.n6948 gnd.n6947 585
R9473 gnd.n6947 gnd.n393 585
R9474 gnd.n6949 gnd.n402 585
R9475 gnd.n7205 gnd.n402 585
R9476 gnd.n6951 gnd.n6950 585
R9477 gnd.n6950 gnd.n401 585
R9478 gnd.n6952 gnd.n409 585
R9479 gnd.n7197 gnd.n409 585
R9480 gnd.n6954 gnd.n6953 585
R9481 gnd.n6955 gnd.n6954 585
R9482 gnd.n6810 gnd.n417 585
R9483 gnd.n7189 gnd.n417 585
R9484 gnd.n6820 gnd.n6819 585
R9485 gnd.n6819 gnd.n6818 585
R9486 gnd.n6817 gnd.n426 585
R9487 gnd.n7181 gnd.n426 585
R9488 gnd.n6816 gnd.n6815 585
R9489 gnd.n6815 gnd.n6814 585
R9490 gnd.n588 gnd.n435 585
R9491 gnd.n7173 gnd.n435 585
R9492 gnd.n7024 gnd.n7023 585
R9493 gnd.n7023 gnd.n7022 585
R9494 gnd.n7025 gnd.n443 585
R9495 gnd.n7165 gnd.n443 585
R9496 gnd.n7026 gnd.n585 585
R9497 gnd.n6800 gnd.n585 585
R9498 gnd.n7027 gnd.n451 585
R9499 gnd.n7157 gnd.n451 585
R9500 gnd.n5744 gnd.n1383 585
R9501 gnd.n1383 gnd.n1339 585
R9502 gnd.n5746 gnd.n5745 585
R9503 gnd.n5747 gnd.n5746 585
R9504 gnd.n5655 gnd.n1382 585
R9505 gnd.n1389 gnd.n1382 585
R9506 gnd.n5654 gnd.n5653 585
R9507 gnd.n5653 gnd.n5652 585
R9508 gnd.n1385 gnd.n1384 585
R9509 gnd.n5556 gnd.n1385 585
R9510 gnd.n5627 gnd.n1396 585
R9511 gnd.n5640 gnd.n1396 585
R9512 gnd.n5628 gnd.n1405 585
R9513 gnd.n5553 gnd.n1405 585
R9514 gnd.n5630 gnd.n5629 585
R9515 gnd.n5631 gnd.n5630 585
R9516 gnd.n5626 gnd.n1404 585
R9517 gnd.n5621 gnd.n1404 585
R9518 gnd.n5625 gnd.n5624 585
R9519 gnd.n5624 gnd.n5623 585
R9520 gnd.n1407 gnd.n1406 585
R9521 gnd.n5610 gnd.n1407 585
R9522 gnd.n5600 gnd.n1423 585
R9523 gnd.n1423 gnd.n1416 585
R9524 gnd.n5602 gnd.n5601 585
R9525 gnd.n5603 gnd.n5602 585
R9526 gnd.n5599 gnd.n1422 585
R9527 gnd.n1428 gnd.n1422 585
R9528 gnd.n5598 gnd.n5597 585
R9529 gnd.n5597 gnd.n5596 585
R9530 gnd.n1425 gnd.n1424 585
R9531 gnd.n5463 gnd.n1425 585
R9532 gnd.n5584 gnd.n5583 585
R9533 gnd.n5585 gnd.n5584 585
R9534 gnd.n5582 gnd.n1439 585
R9535 gnd.n1439 gnd.n1436 585
R9536 gnd.n5581 gnd.n5580 585
R9537 gnd.n5580 gnd.n5579 585
R9538 gnd.n1441 gnd.n1440 585
R9539 gnd.n5472 gnd.n1441 585
R9540 gnd.n5538 gnd.n5537 585
R9541 gnd.n5539 gnd.n5538 585
R9542 gnd.n5536 gnd.n1453 585
R9543 gnd.n1453 gnd.n1450 585
R9544 gnd.n5535 gnd.n5534 585
R9545 gnd.n5534 gnd.n5533 585
R9546 gnd.n1455 gnd.n1454 585
R9547 gnd.n5479 gnd.n1455 585
R9548 gnd.n5519 gnd.n5518 585
R9549 gnd.n5520 gnd.n5519 585
R9550 gnd.n5517 gnd.n1465 585
R9551 gnd.n5512 gnd.n1465 585
R9552 gnd.n5516 gnd.n5515 585
R9553 gnd.n5515 gnd.n5514 585
R9554 gnd.n1467 gnd.n1466 585
R9555 gnd.n1479 gnd.n1467 585
R9556 gnd.n5447 gnd.n5446 585
R9557 gnd.n5447 gnd.n1477 585
R9558 gnd.n5452 gnd.n5451 585
R9559 gnd.n5451 gnd.n5450 585
R9560 gnd.n5453 gnd.n1487 585
R9561 gnd.n5492 gnd.n1487 585
R9562 gnd.n5454 gnd.n1496 585
R9563 gnd.n1496 gnd.n1495 585
R9564 gnd.n5456 gnd.n5455 585
R9565 gnd.n5457 gnd.n5456 585
R9566 gnd.n5445 gnd.n1494 585
R9567 gnd.n5440 gnd.n1494 585
R9568 gnd.n5444 gnd.n5443 585
R9569 gnd.n5443 gnd.n5442 585
R9570 gnd.n1498 gnd.n1497 585
R9571 gnd.n5429 gnd.n1498 585
R9572 gnd.n5419 gnd.n1515 585
R9573 gnd.n1515 gnd.n1507 585
R9574 gnd.n5421 gnd.n5420 585
R9575 gnd.n5422 gnd.n5421 585
R9576 gnd.n5418 gnd.n1514 585
R9577 gnd.n1521 gnd.n1514 585
R9578 gnd.n5417 gnd.n5416 585
R9579 gnd.n5416 gnd.n5415 585
R9580 gnd.n1517 gnd.n1516 585
R9581 gnd.n5318 gnd.n1517 585
R9582 gnd.n5403 gnd.n5402 585
R9583 gnd.n5404 gnd.n5403 585
R9584 gnd.n5401 gnd.n1531 585
R9585 gnd.n1531 gnd.n1528 585
R9586 gnd.n5400 gnd.n5399 585
R9587 gnd.n5399 gnd.n5398 585
R9588 gnd.n1533 gnd.n1532 585
R9589 gnd.n5327 gnd.n1533 585
R9590 gnd.n5366 gnd.n5365 585
R9591 gnd.n5367 gnd.n5366 585
R9592 gnd.n5364 gnd.n1544 585
R9593 gnd.n1544 gnd.n1542 585
R9594 gnd.n5363 gnd.n5362 585
R9595 gnd.n5362 gnd.n5361 585
R9596 gnd.n1546 gnd.n1545 585
R9597 gnd.n5334 gnd.n1546 585
R9598 gnd.n5347 gnd.n5346 585
R9599 gnd.n5348 gnd.n5347 585
R9600 gnd.n5345 gnd.n1559 585
R9601 gnd.n5340 gnd.n1559 585
R9602 gnd.n5344 gnd.n5343 585
R9603 gnd.n5343 gnd.n5342 585
R9604 gnd.n1561 gnd.n1560 585
R9605 gnd.n5312 gnd.n1561 585
R9606 gnd.n5286 gnd.n5285 585
R9607 gnd.n5287 gnd.n5286 585
R9608 gnd.n5291 gnd.n5290 585
R9609 gnd.n5290 gnd.n5289 585
R9610 gnd.n5292 gnd.n1573 585
R9611 gnd.n5303 gnd.n1573 585
R9612 gnd.n5293 gnd.n1584 585
R9613 gnd.n1584 gnd.n1583 585
R9614 gnd.n5295 gnd.n5294 585
R9615 gnd.n5296 gnd.n5295 585
R9616 gnd.n5284 gnd.n1582 585
R9617 gnd.n5279 gnd.n1582 585
R9618 gnd.n5283 gnd.n5282 585
R9619 gnd.n5282 gnd.n5281 585
R9620 gnd.n1586 gnd.n1585 585
R9621 gnd.n5267 gnd.n1586 585
R9622 gnd.n5257 gnd.n1602 585
R9623 gnd.n1602 gnd.n1595 585
R9624 gnd.n5259 gnd.n5258 585
R9625 gnd.n5260 gnd.n5259 585
R9626 gnd.n5256 gnd.n1601 585
R9627 gnd.n1608 gnd.n1601 585
R9628 gnd.n5255 gnd.n5254 585
R9629 gnd.n5254 gnd.n5253 585
R9630 gnd.n1604 gnd.n1603 585
R9631 gnd.n5141 gnd.n1604 585
R9632 gnd.n5240 gnd.n5239 585
R9633 gnd.n5241 gnd.n5240 585
R9634 gnd.n5238 gnd.n1618 585
R9635 gnd.n1618 gnd.n1615 585
R9636 gnd.n5237 gnd.n5236 585
R9637 gnd.n5236 gnd.n5235 585
R9638 gnd.n1620 gnd.n1619 585
R9639 gnd.n5149 gnd.n1620 585
R9640 gnd.n5189 gnd.n5188 585
R9641 gnd.n5190 gnd.n5189 585
R9642 gnd.n5187 gnd.n1632 585
R9643 gnd.n1632 gnd.n1629 585
R9644 gnd.n5186 gnd.n5185 585
R9645 gnd.n5185 gnd.n5184 585
R9646 gnd.n1634 gnd.n1633 585
R9647 gnd.n5156 gnd.n1634 585
R9648 gnd.n5169 gnd.n5168 585
R9649 gnd.n5170 gnd.n5169 585
R9650 gnd.n5167 gnd.n1646 585
R9651 gnd.n5162 gnd.n1646 585
R9652 gnd.n5166 gnd.n5165 585
R9653 gnd.n5165 gnd.n5164 585
R9654 gnd.n1648 gnd.n1647 585
R9655 gnd.n5135 gnd.n1648 585
R9656 gnd.n5109 gnd.n5108 585
R9657 gnd.n5110 gnd.n5109 585
R9658 gnd.n5114 gnd.n5113 585
R9659 gnd.n5113 gnd.n5112 585
R9660 gnd.n5115 gnd.n1660 585
R9661 gnd.n5126 gnd.n1660 585
R9662 gnd.n5116 gnd.n1669 585
R9663 gnd.n5025 gnd.n1669 585
R9664 gnd.n5118 gnd.n5117 585
R9665 gnd.n5119 gnd.n5118 585
R9666 gnd.n5107 gnd.n1668 585
R9667 gnd.n5101 gnd.n1668 585
R9668 gnd.n5106 gnd.n5105 585
R9669 gnd.n5105 gnd.n5104 585
R9670 gnd.n1671 gnd.n1670 585
R9671 gnd.n5090 gnd.n1671 585
R9672 gnd.n5080 gnd.n1687 585
R9673 gnd.n1687 gnd.n1680 585
R9674 gnd.n5082 gnd.n5081 585
R9675 gnd.n5083 gnd.n5082 585
R9676 gnd.n5079 gnd.n1686 585
R9677 gnd.n1693 gnd.n1686 585
R9678 gnd.n5078 gnd.n5077 585
R9679 gnd.n5077 gnd.n5076 585
R9680 gnd.n1689 gnd.n1688 585
R9681 gnd.n4937 gnd.n1689 585
R9682 gnd.n5064 gnd.n5063 585
R9683 gnd.n5065 gnd.n5064 585
R9684 gnd.n5062 gnd.n1703 585
R9685 gnd.n1703 gnd.n1700 585
R9686 gnd.n5061 gnd.n5060 585
R9687 gnd.n5060 gnd.n5059 585
R9688 gnd.n1705 gnd.n1704 585
R9689 gnd.n4945 gnd.n1705 585
R9690 gnd.n5010 gnd.n5009 585
R9691 gnd.n5011 gnd.n5010 585
R9692 gnd.n5008 gnd.n1717 585
R9693 gnd.n1717 gnd.n1714 585
R9694 gnd.n5007 gnd.n5006 585
R9695 gnd.n5006 gnd.n5005 585
R9696 gnd.n1719 gnd.n1718 585
R9697 gnd.n4952 gnd.n1719 585
R9698 gnd.n4991 gnd.n4990 585
R9699 gnd.n4992 gnd.n4991 585
R9700 gnd.n4989 gnd.n1730 585
R9701 gnd.n4984 gnd.n1730 585
R9702 gnd.n4988 gnd.n4987 585
R9703 gnd.n4987 gnd.n4986 585
R9704 gnd.n1732 gnd.n1731 585
R9705 gnd.n1745 gnd.n1732 585
R9706 gnd.n4922 gnd.n4921 585
R9707 gnd.n4922 gnd.n1744 585
R9708 gnd.n4926 gnd.n4925 585
R9709 gnd.n4925 gnd.n4924 585
R9710 gnd.n4927 gnd.n1751 585
R9711 gnd.n4965 gnd.n1751 585
R9712 gnd.n4928 gnd.n1761 585
R9713 gnd.n4671 gnd.n1761 585
R9714 gnd.n4930 gnd.n4929 585
R9715 gnd.n4931 gnd.n4930 585
R9716 gnd.n4920 gnd.n1760 585
R9717 gnd.n4915 gnd.n1760 585
R9718 gnd.n4919 gnd.n4918 585
R9719 gnd.n4918 gnd.n4917 585
R9720 gnd.n1763 gnd.n1762 585
R9721 gnd.n4904 gnd.n1763 585
R9722 gnd.n4894 gnd.n4893 585
R9723 gnd.n4892 gnd.n1810 585
R9724 gnd.n4891 gnd.n1809 585
R9725 gnd.n4896 gnd.n1809 585
R9726 gnd.n4890 gnd.n4889 585
R9727 gnd.n4888 gnd.n4887 585
R9728 gnd.n4886 gnd.n4885 585
R9729 gnd.n4884 gnd.n4883 585
R9730 gnd.n4882 gnd.n4881 585
R9731 gnd.n4880 gnd.n4879 585
R9732 gnd.n4878 gnd.n4877 585
R9733 gnd.n4876 gnd.n4875 585
R9734 gnd.n4874 gnd.n4873 585
R9735 gnd.n4872 gnd.n4871 585
R9736 gnd.n4870 gnd.n4869 585
R9737 gnd.n4868 gnd.n4867 585
R9738 gnd.n4866 gnd.n4865 585
R9739 gnd.n4864 gnd.n4863 585
R9740 gnd.n4862 gnd.n4861 585
R9741 gnd.n4860 gnd.n4859 585
R9742 gnd.n4858 gnd.n4857 585
R9743 gnd.n4856 gnd.n4855 585
R9744 gnd.n4854 gnd.n4853 585
R9745 gnd.n4852 gnd.n4851 585
R9746 gnd.n4850 gnd.n4849 585
R9747 gnd.n4848 gnd.n4847 585
R9748 gnd.n4846 gnd.n4845 585
R9749 gnd.n4844 gnd.n4843 585
R9750 gnd.n4842 gnd.n4841 585
R9751 gnd.n4840 gnd.n4839 585
R9752 gnd.n4838 gnd.n4837 585
R9753 gnd.n4836 gnd.n4835 585
R9754 gnd.n4834 gnd.n4833 585
R9755 gnd.n4832 gnd.n4831 585
R9756 gnd.n4830 gnd.n1894 585
R9757 gnd.n1893 gnd.n1892 585
R9758 gnd.n1891 gnd.n1890 585
R9759 gnd.n1888 gnd.n1887 585
R9760 gnd.n1886 gnd.n1885 585
R9761 gnd.n1884 gnd.n1883 585
R9762 gnd.n1882 gnd.n1881 585
R9763 gnd.n1880 gnd.n1879 585
R9764 gnd.n1878 gnd.n1877 585
R9765 gnd.n1876 gnd.n1875 585
R9766 gnd.n1874 gnd.n1873 585
R9767 gnd.n1872 gnd.n1871 585
R9768 gnd.n1870 gnd.n1869 585
R9769 gnd.n1868 gnd.n1867 585
R9770 gnd.n1866 gnd.n1865 585
R9771 gnd.n1864 gnd.n1863 585
R9772 gnd.n1862 gnd.n1861 585
R9773 gnd.n1860 gnd.n1859 585
R9774 gnd.n1858 gnd.n1857 585
R9775 gnd.n1856 gnd.n1855 585
R9776 gnd.n1854 gnd.n1853 585
R9777 gnd.n1852 gnd.n1851 585
R9778 gnd.n1850 gnd.n1849 585
R9779 gnd.n1848 gnd.n1847 585
R9780 gnd.n1846 gnd.n1845 585
R9781 gnd.n1844 gnd.n1843 585
R9782 gnd.n1842 gnd.n1841 585
R9783 gnd.n1840 gnd.n1839 585
R9784 gnd.n1838 gnd.n1837 585
R9785 gnd.n1776 gnd.n1775 585
R9786 gnd.n4899 gnd.n4898 585
R9787 gnd.n4900 gnd.n1774 585
R9788 gnd.n5751 gnd.n5750 585
R9789 gnd.n5753 gnd.n5752 585
R9790 gnd.n5755 gnd.n5754 585
R9791 gnd.n5757 gnd.n5756 585
R9792 gnd.n5759 gnd.n5758 585
R9793 gnd.n5761 gnd.n5760 585
R9794 gnd.n5763 gnd.n5762 585
R9795 gnd.n5765 gnd.n5764 585
R9796 gnd.n5767 gnd.n5766 585
R9797 gnd.n5769 gnd.n5768 585
R9798 gnd.n5771 gnd.n5770 585
R9799 gnd.n5773 gnd.n5772 585
R9800 gnd.n5775 gnd.n5774 585
R9801 gnd.n5777 gnd.n5776 585
R9802 gnd.n5779 gnd.n5778 585
R9803 gnd.n5781 gnd.n5780 585
R9804 gnd.n5783 gnd.n5782 585
R9805 gnd.n5785 gnd.n5784 585
R9806 gnd.n5787 gnd.n5786 585
R9807 gnd.n5789 gnd.n5788 585
R9808 gnd.n5791 gnd.n5790 585
R9809 gnd.n5793 gnd.n5792 585
R9810 gnd.n5795 gnd.n5794 585
R9811 gnd.n5797 gnd.n5796 585
R9812 gnd.n5799 gnd.n5798 585
R9813 gnd.n5801 gnd.n5800 585
R9814 gnd.n5803 gnd.n5802 585
R9815 gnd.n5805 gnd.n5804 585
R9816 gnd.n5807 gnd.n5806 585
R9817 gnd.n5810 gnd.n5809 585
R9818 gnd.n5812 gnd.n5811 585
R9819 gnd.n5814 gnd.n5813 585
R9820 gnd.n5816 gnd.n5815 585
R9821 gnd.n5677 gnd.n556 585
R9822 gnd.n5679 gnd.n5678 585
R9823 gnd.n5681 gnd.n5680 585
R9824 gnd.n5683 gnd.n5682 585
R9825 gnd.n5686 gnd.n5685 585
R9826 gnd.n5688 gnd.n5687 585
R9827 gnd.n5690 gnd.n5689 585
R9828 gnd.n5692 gnd.n5691 585
R9829 gnd.n5694 gnd.n5693 585
R9830 gnd.n5696 gnd.n5695 585
R9831 gnd.n5698 gnd.n5697 585
R9832 gnd.n5700 gnd.n5699 585
R9833 gnd.n5702 gnd.n5701 585
R9834 gnd.n5704 gnd.n5703 585
R9835 gnd.n5706 gnd.n5705 585
R9836 gnd.n5708 gnd.n5707 585
R9837 gnd.n5710 gnd.n5709 585
R9838 gnd.n5712 gnd.n5711 585
R9839 gnd.n5714 gnd.n5713 585
R9840 gnd.n5716 gnd.n5715 585
R9841 gnd.n5718 gnd.n5717 585
R9842 gnd.n5720 gnd.n5719 585
R9843 gnd.n5722 gnd.n5721 585
R9844 gnd.n5724 gnd.n5723 585
R9845 gnd.n5726 gnd.n5725 585
R9846 gnd.n5728 gnd.n5727 585
R9847 gnd.n5730 gnd.n5729 585
R9848 gnd.n5732 gnd.n5731 585
R9849 gnd.n5734 gnd.n5733 585
R9850 gnd.n5736 gnd.n5735 585
R9851 gnd.n5738 gnd.n5737 585
R9852 gnd.n5740 gnd.n5739 585
R9853 gnd.n5742 gnd.n5741 585
R9854 gnd.n5749 gnd.n1376 585
R9855 gnd.n5749 gnd.n1339 585
R9856 gnd.n5748 gnd.n1378 585
R9857 gnd.n5748 gnd.n5747 585
R9858 gnd.n5635 gnd.n1377 585
R9859 gnd.n1389 gnd.n1377 585
R9860 gnd.n5636 gnd.n1387 585
R9861 gnd.n5652 gnd.n1387 585
R9862 gnd.n5637 gnd.n1398 585
R9863 gnd.n5556 gnd.n1398 585
R9864 gnd.n5639 gnd.n5638 585
R9865 gnd.n5640 gnd.n5639 585
R9866 gnd.n5634 gnd.n1397 585
R9867 gnd.n5553 gnd.n1397 585
R9868 gnd.n5633 gnd.n5632 585
R9869 gnd.n5632 gnd.n5631 585
R9870 gnd.n1400 gnd.n1399 585
R9871 gnd.n5621 gnd.n1400 585
R9872 gnd.n5607 gnd.n1409 585
R9873 gnd.n5623 gnd.n1409 585
R9874 gnd.n5609 gnd.n5608 585
R9875 gnd.n5610 gnd.n5609 585
R9876 gnd.n5606 gnd.n1418 585
R9877 gnd.n1418 gnd.n1416 585
R9878 gnd.n5605 gnd.n5604 585
R9879 gnd.n5604 gnd.n5603 585
R9880 gnd.n1420 gnd.n1419 585
R9881 gnd.n1428 gnd.n1420 585
R9882 gnd.n5461 gnd.n1427 585
R9883 gnd.n5596 gnd.n1427 585
R9884 gnd.n5465 gnd.n5464 585
R9885 gnd.n5464 gnd.n5463 585
R9886 gnd.n5466 gnd.n1438 585
R9887 gnd.n5585 gnd.n1438 585
R9888 gnd.n5468 gnd.n5467 585
R9889 gnd.n5467 gnd.n1436 585
R9890 gnd.n5469 gnd.n1443 585
R9891 gnd.n5579 gnd.n1443 585
R9892 gnd.n5474 gnd.n5473 585
R9893 gnd.n5473 gnd.n5472 585
R9894 gnd.n5475 gnd.n1451 585
R9895 gnd.n5539 gnd.n1451 585
R9896 gnd.n5477 gnd.n5476 585
R9897 gnd.n5476 gnd.n1450 585
R9898 gnd.n5478 gnd.n1456 585
R9899 gnd.n5533 gnd.n1456 585
R9900 gnd.n5481 gnd.n5480 585
R9901 gnd.n5480 gnd.n5479 585
R9902 gnd.n5482 gnd.n1463 585
R9903 gnd.n5520 gnd.n1463 585
R9904 gnd.n5483 gnd.n1469 585
R9905 gnd.n5512 gnd.n1469 585
R9906 gnd.n5484 gnd.n1468 585
R9907 gnd.n5514 gnd.n1468 585
R9908 gnd.n5486 gnd.n5485 585
R9909 gnd.n5486 gnd.n1479 585
R9910 gnd.n5488 gnd.n5487 585
R9911 gnd.n5487 gnd.n1477 585
R9912 gnd.n5489 gnd.n1489 585
R9913 gnd.n5450 gnd.n1489 585
R9914 gnd.n5491 gnd.n5490 585
R9915 gnd.n5492 gnd.n5491 585
R9916 gnd.n5460 gnd.n1488 585
R9917 gnd.n1495 gnd.n1488 585
R9918 gnd.n5459 gnd.n5458 585
R9919 gnd.n5458 gnd.n5457 585
R9920 gnd.n1491 gnd.n1490 585
R9921 gnd.n5440 gnd.n1491 585
R9922 gnd.n5426 gnd.n1500 585
R9923 gnd.n5442 gnd.n1500 585
R9924 gnd.n5428 gnd.n5427 585
R9925 gnd.n5429 gnd.n5428 585
R9926 gnd.n5425 gnd.n1509 585
R9927 gnd.n1509 gnd.n1507 585
R9928 gnd.n5424 gnd.n5423 585
R9929 gnd.n5423 gnd.n5422 585
R9930 gnd.n1511 gnd.n1510 585
R9931 gnd.n1521 gnd.n1511 585
R9932 gnd.n5316 gnd.n1519 585
R9933 gnd.n5415 gnd.n1519 585
R9934 gnd.n5320 gnd.n5319 585
R9935 gnd.n5319 gnd.n5318 585
R9936 gnd.n5321 gnd.n1530 585
R9937 gnd.n5404 gnd.n1530 585
R9938 gnd.n5323 gnd.n5322 585
R9939 gnd.n5322 gnd.n1528 585
R9940 gnd.n5324 gnd.n1535 585
R9941 gnd.n5398 gnd.n1535 585
R9942 gnd.n5329 gnd.n5328 585
R9943 gnd.n5328 gnd.n5327 585
R9944 gnd.n5330 gnd.n1543 585
R9945 gnd.n5367 gnd.n1543 585
R9946 gnd.n5332 gnd.n5331 585
R9947 gnd.n5331 gnd.n1542 585
R9948 gnd.n5333 gnd.n1548 585
R9949 gnd.n5361 gnd.n1548 585
R9950 gnd.n5336 gnd.n5335 585
R9951 gnd.n5335 gnd.n5334 585
R9952 gnd.n5337 gnd.n1556 585
R9953 gnd.n5348 gnd.n1556 585
R9954 gnd.n5339 gnd.n5338 585
R9955 gnd.n5340 gnd.n5339 585
R9956 gnd.n5315 gnd.n1563 585
R9957 gnd.n5342 gnd.n1563 585
R9958 gnd.n5314 gnd.n5313 585
R9959 gnd.n5313 gnd.n5312 585
R9960 gnd.n1565 gnd.n1564 585
R9961 gnd.n5287 gnd.n1565 585
R9962 gnd.n5300 gnd.n1577 585
R9963 gnd.n5289 gnd.n1577 585
R9964 gnd.n5302 gnd.n5301 585
R9965 gnd.n5303 gnd.n5302 585
R9966 gnd.n5299 gnd.n1576 585
R9967 gnd.n1583 gnd.n1576 585
R9968 gnd.n5298 gnd.n5297 585
R9969 gnd.n5297 gnd.n5296 585
R9970 gnd.n1579 gnd.n1578 585
R9971 gnd.n5279 gnd.n1579 585
R9972 gnd.n5264 gnd.n1588 585
R9973 gnd.n5281 gnd.n1588 585
R9974 gnd.n5266 gnd.n5265 585
R9975 gnd.n5267 gnd.n5266 585
R9976 gnd.n5263 gnd.n1597 585
R9977 gnd.n1597 gnd.n1595 585
R9978 gnd.n5262 gnd.n5261 585
R9979 gnd.n5261 gnd.n5260 585
R9980 gnd.n1599 gnd.n1598 585
R9981 gnd.n1608 gnd.n1599 585
R9982 gnd.n5139 gnd.n1606 585
R9983 gnd.n5253 gnd.n1606 585
R9984 gnd.n5143 gnd.n5142 585
R9985 gnd.n5142 gnd.n5141 585
R9986 gnd.n5144 gnd.n1617 585
R9987 gnd.n5241 gnd.n1617 585
R9988 gnd.n5146 gnd.n5145 585
R9989 gnd.n5145 gnd.n1615 585
R9990 gnd.n5147 gnd.n1622 585
R9991 gnd.n5235 gnd.n1622 585
R9992 gnd.n5151 gnd.n5150 585
R9993 gnd.n5150 gnd.n5149 585
R9994 gnd.n5152 gnd.n1630 585
R9995 gnd.n5190 gnd.n1630 585
R9996 gnd.n5154 gnd.n5153 585
R9997 gnd.n5153 gnd.n1629 585
R9998 gnd.n5155 gnd.n1636 585
R9999 gnd.n5184 gnd.n1636 585
R10000 gnd.n5158 gnd.n5157 585
R10001 gnd.n5157 gnd.n5156 585
R10002 gnd.n5159 gnd.n1644 585
R10003 gnd.n5170 gnd.n1644 585
R10004 gnd.n5161 gnd.n5160 585
R10005 gnd.n5162 gnd.n5161 585
R10006 gnd.n5138 gnd.n1650 585
R10007 gnd.n5164 gnd.n1650 585
R10008 gnd.n5137 gnd.n5136 585
R10009 gnd.n5136 gnd.n5135 585
R10010 gnd.n1652 gnd.n1651 585
R10011 gnd.n5110 gnd.n1652 585
R10012 gnd.n5123 gnd.n1663 585
R10013 gnd.n5112 gnd.n1663 585
R10014 gnd.n5125 gnd.n5124 585
R10015 gnd.n5126 gnd.n5125 585
R10016 gnd.n5122 gnd.n1662 585
R10017 gnd.n5025 gnd.n1662 585
R10018 gnd.n5121 gnd.n5120 585
R10019 gnd.n5120 gnd.n5119 585
R10020 gnd.n1665 gnd.n1664 585
R10021 gnd.n5101 gnd.n1665 585
R10022 gnd.n5087 gnd.n1673 585
R10023 gnd.n5104 gnd.n1673 585
R10024 gnd.n5089 gnd.n5088 585
R10025 gnd.n5090 gnd.n5089 585
R10026 gnd.n5086 gnd.n1682 585
R10027 gnd.n1682 gnd.n1680 585
R10028 gnd.n5085 gnd.n5084 585
R10029 gnd.n5084 gnd.n5083 585
R10030 gnd.n1684 gnd.n1683 585
R10031 gnd.n1693 gnd.n1684 585
R10032 gnd.n4935 gnd.n1692 585
R10033 gnd.n5076 gnd.n1692 585
R10034 gnd.n4939 gnd.n4938 585
R10035 gnd.n4938 gnd.n4937 585
R10036 gnd.n4940 gnd.n1702 585
R10037 gnd.n5065 gnd.n1702 585
R10038 gnd.n4942 gnd.n4941 585
R10039 gnd.n4941 gnd.n1700 585
R10040 gnd.n4943 gnd.n1707 585
R10041 gnd.n5059 gnd.n1707 585
R10042 gnd.n4947 gnd.n4946 585
R10043 gnd.n4946 gnd.n4945 585
R10044 gnd.n4948 gnd.n1715 585
R10045 gnd.n5011 gnd.n1715 585
R10046 gnd.n4950 gnd.n4949 585
R10047 gnd.n4949 gnd.n1714 585
R10048 gnd.n4951 gnd.n1721 585
R10049 gnd.n5005 gnd.n1721 585
R10050 gnd.n4954 gnd.n4953 585
R10051 gnd.n4953 gnd.n4952 585
R10052 gnd.n4955 gnd.n1728 585
R10053 gnd.n4992 gnd.n1728 585
R10054 gnd.n4956 gnd.n1736 585
R10055 gnd.n4984 gnd.n1736 585
R10056 gnd.n4957 gnd.n1735 585
R10057 gnd.n4986 gnd.n1735 585
R10058 gnd.n4959 gnd.n4958 585
R10059 gnd.n4959 gnd.n1745 585
R10060 gnd.n4961 gnd.n4960 585
R10061 gnd.n4960 gnd.n1744 585
R10062 gnd.n4962 gnd.n1754 585
R10063 gnd.n4924 gnd.n1754 585
R10064 gnd.n4964 gnd.n4963 585
R10065 gnd.n4965 gnd.n4964 585
R10066 gnd.n4934 gnd.n1753 585
R10067 gnd.n4671 gnd.n1753 585
R10068 gnd.n4933 gnd.n4932 585
R10069 gnd.n4932 gnd.n4931 585
R10070 gnd.n1756 gnd.n1755 585
R10071 gnd.n4915 gnd.n1756 585
R10072 gnd.n4901 gnd.n1765 585
R10073 gnd.n4917 gnd.n1765 585
R10074 gnd.n4903 gnd.n4902 585
R10075 gnd.n4904 gnd.n4903 585
R10076 gnd.n6787 gnd.n6786 585
R10077 gnd.n6787 gnd.n419 585
R10078 gnd.n6789 gnd.n6788 585
R10079 gnd.n6788 gnd.n416 585
R10080 gnd.n6790 gnd.n600 585
R10081 gnd.n600 gnd.n428 585
R10082 gnd.n6792 gnd.n6791 585
R10083 gnd.n6792 gnd.n425 585
R10084 gnd.n6793 gnd.n599 585
R10085 gnd.n6793 gnd.n437 585
R10086 gnd.n6795 gnd.n6794 585
R10087 gnd.n6794 gnd.n434 585
R10088 gnd.n6796 gnd.n594 585
R10089 gnd.n594 gnd.n445 585
R10090 gnd.n6798 gnd.n6797 585
R10091 gnd.n6799 gnd.n6798 585
R10092 gnd.n595 gnd.n593 585
R10093 gnd.n593 gnd.n453 585
R10094 gnd.n1242 gnd.n1237 585
R10095 gnd.n1237 gnd.n450 585
R10096 gnd.n1244 gnd.n1243 585
R10097 gnd.n1244 gnd.n506 585
R10098 gnd.n1245 gnd.n1236 585
R10099 gnd.n5891 gnd.n1245 585
R10100 gnd.n5894 gnd.n5893 585
R10101 gnd.n5893 gnd.n5892 585
R10102 gnd.n5895 gnd.n1231 585
R10103 gnd.n1231 gnd.n1229 585
R10104 gnd.n5897 gnd.n5896 585
R10105 gnd.n5898 gnd.n5897 585
R10106 gnd.n1232 gnd.n1230 585
R10107 gnd.n1230 gnd.n1227 585
R10108 gnd.n5880 gnd.n5879 585
R10109 gnd.n5881 gnd.n5880 585
R10110 gnd.n1304 gnd.n1303 585
R10111 gnd.n5870 gnd.n1303 585
R10112 gnd.n5874 gnd.n5873 585
R10113 gnd.n5873 gnd.n5872 585
R10114 gnd.n1307 gnd.n1306 585
R10115 gnd.n5858 gnd.n1307 585
R10116 gnd.n5856 gnd.n5855 585
R10117 gnd.n5857 gnd.n5856 585
R10118 gnd.n1317 gnd.n1316 585
R10119 gnd.n5847 gnd.n1316 585
R10120 gnd.n5851 gnd.n5850 585
R10121 gnd.n5850 gnd.n5849 585
R10122 gnd.n1320 gnd.n1319 585
R10123 gnd.n5838 gnd.n1320 585
R10124 gnd.n5836 gnd.n5835 585
R10125 gnd.n5837 gnd.n5836 585
R10126 gnd.n1330 gnd.n1329 585
R10127 gnd.n5827 gnd.n1329 585
R10128 gnd.n5831 gnd.n5830 585
R10129 gnd.n5830 gnd.n5829 585
R10130 gnd.n1333 gnd.n1332 585
R10131 gnd.n5818 gnd.n1333 585
R10132 gnd.n5647 gnd.n1391 585
R10133 gnd.n1391 gnd.n1381 585
R10134 gnd.n5649 gnd.n5648 585
R10135 gnd.n5650 gnd.n5649 585
R10136 gnd.n1392 gnd.n1390 585
R10137 gnd.n1390 gnd.n1386 585
R10138 gnd.n5642 gnd.n5641 585
R10139 gnd.n5641 gnd.n5640 585
R10140 gnd.n1395 gnd.n1394 585
R10141 gnd.n1403 gnd.n1395 585
R10142 gnd.n5619 gnd.n5618 585
R10143 gnd.n5620 gnd.n5619 585
R10144 gnd.n1412 gnd.n1411 585
R10145 gnd.n1411 gnd.n1408 585
R10146 gnd.n5614 gnd.n5613 585
R10147 gnd.n5613 gnd.n5612 585
R10148 gnd.n1415 gnd.n1414 585
R10149 gnd.n1421 gnd.n1415 585
R10150 gnd.n5594 gnd.n5593 585
R10151 gnd.n5595 gnd.n5594 585
R10152 gnd.n1432 gnd.n1431 585
R10153 gnd.n5462 gnd.n1431 585
R10154 gnd.n5589 gnd.n5588 585
R10155 gnd.n5588 gnd.n5587 585
R10156 gnd.n1435 gnd.n1434 585
R10157 gnd.n1442 gnd.n1435 585
R10158 gnd.n5528 gnd.n1458 585
R10159 gnd.n1458 gnd.n1452 585
R10160 gnd.n5530 gnd.n5529 585
R10161 gnd.n5531 gnd.n5530 585
R10162 gnd.n1459 gnd.n1457 585
R10163 gnd.n1457 gnd.t59 585
R10164 gnd.n5523 gnd.n5522 585
R10165 gnd.n5522 gnd.n5521 585
R10166 gnd.n1462 gnd.n1461 585
R10167 gnd.n5513 gnd.n1462 585
R10168 gnd.n5499 gnd.n5498 585
R10169 gnd.n5500 gnd.n5499 585
R10170 gnd.n1481 gnd.n1480 585
R10171 gnd.n5449 gnd.n1480 585
R10172 gnd.n5494 gnd.n5493 585
R10173 gnd.n5493 gnd.n5492 585
R10174 gnd.n1484 gnd.n1483 585
R10175 gnd.n1493 gnd.n1484 585
R10176 gnd.n5438 gnd.n5437 585
R10177 gnd.n5439 gnd.n5438 585
R10178 gnd.n1503 gnd.n1502 585
R10179 gnd.n1502 gnd.n1499 585
R10180 gnd.n5433 gnd.n5432 585
R10181 gnd.n5432 gnd.n5431 585
R10182 gnd.n1506 gnd.n1505 585
R10183 gnd.n1520 gnd.n1506 585
R10184 gnd.n5413 gnd.n5412 585
R10185 gnd.n5414 gnd.n5413 585
R10186 gnd.n1524 gnd.n1523 585
R10187 gnd.n5317 gnd.n1523 585
R10188 gnd.n5408 gnd.n5407 585
R10189 gnd.n5407 gnd.n5406 585
R10190 gnd.n1527 gnd.n1526 585
R10191 gnd.n1534 gnd.n1527 585
R10192 gnd.n5356 gnd.n1550 585
R10193 gnd.n5325 gnd.n1550 585
R10194 gnd.n5358 gnd.n5357 585
R10195 gnd.n5359 gnd.n5358 585
R10196 gnd.n1551 gnd.n1549 585
R10197 gnd.n1549 gnd.n1547 585
R10198 gnd.n5351 gnd.n5350 585
R10199 gnd.n5350 gnd.n5349 585
R10200 gnd.n1554 gnd.n1553 585
R10201 gnd.n5341 gnd.n1554 585
R10202 gnd.n5310 gnd.n5309 585
R10203 gnd.n5311 gnd.n5310 585
R10204 gnd.n1568 gnd.n1567 585
R10205 gnd.n5288 gnd.n1567 585
R10206 gnd.n5305 gnd.n5304 585
R10207 gnd.n5304 gnd.n5303 585
R10208 gnd.n1571 gnd.n1570 585
R10209 gnd.n1581 gnd.n1571 585
R10210 gnd.n5277 gnd.n5276 585
R10211 gnd.n5278 gnd.n5277 585
R10212 gnd.n1591 gnd.n1590 585
R10213 gnd.n1590 gnd.n1587 585
R10214 gnd.n5272 gnd.n5271 585
R10215 gnd.n5271 gnd.n5270 585
R10216 gnd.n1594 gnd.n1593 585
R10217 gnd.n1607 gnd.n1594 585
R10218 gnd.n5251 gnd.n5250 585
R10219 gnd.n5252 gnd.n5251 585
R10220 gnd.n1611 gnd.n1610 585
R10221 gnd.n5140 gnd.n1610 585
R10222 gnd.n5246 gnd.n5245 585
R10223 gnd.n5245 gnd.n5244 585
R10224 gnd.n1614 gnd.n1613 585
R10225 gnd.n1621 gnd.n1614 585
R10226 gnd.n5178 gnd.n1638 585
R10227 gnd.n1638 gnd.n1631 585
R10228 gnd.n5180 gnd.n5179 585
R10229 gnd.n5181 gnd.n5180 585
R10230 gnd.n1639 gnd.n1637 585
R10231 gnd.n1637 gnd.n1635 585
R10232 gnd.n5173 gnd.n5172 585
R10233 gnd.n5172 gnd.n5171 585
R10234 gnd.n1642 gnd.n1641 585
R10235 gnd.n5163 gnd.n1642 585
R10236 gnd.n5133 gnd.n5132 585
R10237 gnd.n5134 gnd.n5133 585
R10238 gnd.n1656 gnd.n1655 585
R10239 gnd.n5111 gnd.n1655 585
R10240 gnd.n5128 gnd.n5127 585
R10241 gnd.n5127 gnd.n5126 585
R10242 gnd.n1659 gnd.n1658 585
R10243 gnd.n1667 gnd.n1659 585
R10244 gnd.n5099 gnd.n5098 585
R10245 gnd.n5100 gnd.n5099 585
R10246 gnd.n1676 gnd.n1675 585
R10247 gnd.n1675 gnd.n1672 585
R10248 gnd.n5094 gnd.n5093 585
R10249 gnd.n5093 gnd.n5092 585
R10250 gnd.n1679 gnd.n1678 585
R10251 gnd.t57 gnd.n1679 585
R10252 gnd.n5074 gnd.n5073 585
R10253 gnd.n5075 gnd.n5074 585
R10254 gnd.n1696 gnd.n1695 585
R10255 gnd.n4936 gnd.n1695 585
R10256 gnd.n5069 gnd.n5068 585
R10257 gnd.n5068 gnd.n5067 585
R10258 gnd.n1699 gnd.n1698 585
R10259 gnd.n1706 gnd.n1699 585
R10260 gnd.n5000 gnd.n1723 585
R10261 gnd.n1723 gnd.n1716 585
R10262 gnd.n5002 gnd.n5001 585
R10263 gnd.n5003 gnd.n5002 585
R10264 gnd.n1724 gnd.n1722 585
R10265 gnd.n1722 gnd.n1720 585
R10266 gnd.n4995 gnd.n4994 585
R10267 gnd.n4994 gnd.n4993 585
R10268 gnd.n1727 gnd.n1726 585
R10269 gnd.n4985 gnd.n1727 585
R10270 gnd.n4972 gnd.n4971 585
R10271 gnd.n4973 gnd.n4972 585
R10272 gnd.n1747 gnd.n1746 585
R10273 gnd.n4923 gnd.n1746 585
R10274 gnd.n4967 gnd.n4966 585
R10275 gnd.n4966 gnd.n4965 585
R10276 gnd.n1750 gnd.n1749 585
R10277 gnd.n1759 gnd.n1750 585
R10278 gnd.n4913 gnd.n4912 585
R10279 gnd.n4914 gnd.n4913 585
R10280 gnd.n1768 gnd.n1767 585
R10281 gnd.n1767 gnd.n1764 585
R10282 gnd.n4908 gnd.n4907 585
R10283 gnd.n4907 gnd.n4906 585
R10284 gnd.n1771 gnd.n1770 585
R10285 gnd.n1777 gnd.n1771 585
R10286 gnd.n4663 gnd.n4662 585
R10287 gnd.n4664 gnd.n4663 585
R10288 gnd.n4600 gnd.n4599 585
R10289 gnd.n4654 gnd.n4599 585
R10290 gnd.n4658 gnd.n4657 585
R10291 gnd.n4657 gnd.n4656 585
R10292 gnd.n4603 gnd.n4602 585
R10293 gnd.n4652 gnd.n4603 585
R10294 gnd.n4647 gnd.n4646 585
R10295 gnd.n4648 gnd.n4647 585
R10296 gnd.n4606 gnd.n4605 585
R10297 gnd.n4638 gnd.n4605 585
R10298 gnd.n4642 gnd.n4641 585
R10299 gnd.n4641 gnd.n4640 585
R10300 gnd.n4609 gnd.n4608 585
R10301 gnd.n4636 gnd.n4609 585
R10302 gnd.n4631 gnd.n4630 585
R10303 gnd.n4632 gnd.n4631 585
R10304 gnd.n4612 gnd.n4611 585
R10305 gnd.n4622 gnd.n4611 585
R10306 gnd.n4626 gnd.n4625 585
R10307 gnd.n4625 gnd.n4624 585
R10308 gnd.n4619 gnd.n4614 585
R10309 gnd.n4620 gnd.n4619 585
R10310 gnd.n4618 gnd.n4617 585
R10311 gnd.n4618 gnd.n4491 585
R10312 gnd.n4476 gnd.n4475 585
R10313 gnd.n4766 gnd.n4476 585
R10314 gnd.n4769 gnd.n4768 585
R10315 gnd.n4768 gnd.n4767 585
R10316 gnd.n4770 gnd.n4451 585
R10317 gnd.n4477 gnd.n4451 585
R10318 gnd.n4772 gnd.n4771 585
R10319 gnd.n4773 gnd.n4772 585
R10320 gnd.n4452 gnd.n4450 585
R10321 gnd.n4450 gnd.n1094 585
R10322 gnd.n4469 gnd.n4468 585
R10323 gnd.n4468 gnd.n1091 585
R10324 gnd.n4467 gnd.n4454 585
R10325 gnd.n4467 gnd.n1083 585
R10326 gnd.n4466 gnd.n4465 585
R10327 gnd.n4466 gnd.n1080 585
R10328 gnd.n4456 gnd.n4455 585
R10329 gnd.n4455 gnd.n1071 585
R10330 gnd.n4461 gnd.n4460 585
R10331 gnd.n4460 gnd.n1068 585
R10332 gnd.n4459 gnd.n1054 585
R10333 gnd.n2004 gnd.n1054 585
R10334 gnd.n6080 gnd.n1055 585
R10335 gnd.n6080 gnd.n6079 585
R10336 gnd.n5901 gnd.n5900 585
R10337 gnd.n5900 gnd.n5899 585
R10338 gnd.n5902 gnd.n1226 585
R10339 gnd.n5882 gnd.n1226 585
R10340 gnd.n5868 gnd.n1224 585
R10341 gnd.n5869 gnd.n5868 585
R10342 gnd.n5906 gnd.n1223 585
R10343 gnd.n5871 gnd.n1223 585
R10344 gnd.n5907 gnd.n1222 585
R10345 gnd.n1308 gnd.n1222 585
R10346 gnd.n5908 gnd.n1221 585
R10347 gnd.n5859 gnd.n1221 585
R10348 gnd.n1314 gnd.n1219 585
R10349 gnd.n1315 gnd.n1314 585
R10350 gnd.n5912 gnd.n1218 585
R10351 gnd.n5848 gnd.n1218 585
R10352 gnd.n5913 gnd.n1217 585
R10353 gnd.n1321 gnd.n1217 585
R10354 gnd.n5914 gnd.n1216 585
R10355 gnd.n5839 gnd.n1216 585
R10356 gnd.n1327 gnd.n1214 585
R10357 gnd.n1328 gnd.n1327 585
R10358 gnd.n5918 gnd.n1213 585
R10359 gnd.n5828 gnd.n1213 585
R10360 gnd.n5919 gnd.n1212 585
R10361 gnd.n5817 gnd.n1212 585
R10362 gnd.n5920 gnd.n1211 585
R10363 gnd.n5819 gnd.n1211 585
R10364 gnd.n1379 gnd.n1209 585
R10365 gnd.n1380 gnd.n1379 585
R10366 gnd.n5924 gnd.n1208 585
R10367 gnd.n5651 gnd.n1208 585
R10368 gnd.n5925 gnd.n1207 585
R10369 gnd.n5557 gnd.n1207 585
R10370 gnd.n5926 gnd.n1206 585
R10371 gnd.n5554 gnd.n1206 585
R10372 gnd.n1401 gnd.n1204 585
R10373 gnd.n1402 gnd.n1401 585
R10374 gnd.n5930 gnd.n1203 585
R10375 gnd.n5622 gnd.n1203 585
R10376 gnd.n5931 gnd.n1202 585
R10377 gnd.n5611 gnd.n1202 585
R10378 gnd.n5932 gnd.n1201 585
R10379 gnd.n5548 gnd.n1201 585
R10380 gnd.n1429 gnd.n1199 585
R10381 gnd.n1430 gnd.n1429 585
R10382 gnd.n5936 gnd.n1198 585
R10383 gnd.n1426 gnd.n1198 585
R10384 gnd.n5937 gnd.n1197 585
R10385 gnd.n5586 gnd.n1197 585
R10386 gnd.n5938 gnd.n1196 585
R10387 gnd.n5578 gnd.n1196 585
R10388 gnd.n5470 gnd.n1194 585
R10389 gnd.n5471 gnd.n5470 585
R10390 gnd.n5942 gnd.n1193 585
R10391 gnd.n5540 gnd.n1193 585
R10392 gnd.n5943 gnd.n1192 585
R10393 gnd.n5532 gnd.n1192 585
R10394 gnd.n5944 gnd.n1191 585
R10395 gnd.n1464 gnd.n1191 585
R10396 gnd.n5510 gnd.n1189 585
R10397 gnd.n5511 gnd.n5510 585
R10398 gnd.n5948 gnd.n1188 585
R10399 gnd.n1478 gnd.n1188 585
R10400 gnd.n5949 gnd.n1187 585
R10401 gnd.n5501 gnd.n1187 585
R10402 gnd.n5950 gnd.n1186 585
R10403 gnd.n5448 gnd.n1186 585
R10404 gnd.n1485 gnd.n1184 585
R10405 gnd.n1486 gnd.n1485 585
R10406 gnd.n5954 gnd.n1183 585
R10407 gnd.n1492 gnd.n1183 585
R10408 gnd.n5955 gnd.n1182 585
R10409 gnd.n5441 gnd.n1182 585
R10410 gnd.n5956 gnd.n1181 585
R10411 gnd.n5430 gnd.n1181 585
R10412 gnd.n1512 gnd.n1179 585
R10413 gnd.n1513 gnd.n1512 585
R10414 gnd.n5960 gnd.n1178 585
R10415 gnd.n1522 gnd.n1178 585
R10416 gnd.n5961 gnd.n1177 585
R10417 gnd.n1518 gnd.n1177 585
R10418 gnd.n5962 gnd.n1176 585
R10419 gnd.n5405 gnd.n1176 585
R10420 gnd.n5396 gnd.n1174 585
R10421 gnd.n5397 gnd.n5396 585
R10422 gnd.n5966 gnd.n1173 585
R10423 gnd.n5326 gnd.n1173 585
R10424 gnd.n5967 gnd.n1172 585
R10425 gnd.n5368 gnd.n1172 585
R10426 gnd.n5968 gnd.n1171 585
R10427 gnd.n5360 gnd.n1171 585
R10428 gnd.n1557 gnd.n1169 585
R10429 gnd.n1558 gnd.n1557 585
R10430 gnd.n5972 gnd.n1168 585
R10431 gnd.n1555 gnd.n1168 585
R10432 gnd.n5973 gnd.n1167 585
R10433 gnd.n1562 gnd.n1167 585
R10434 gnd.n5974 gnd.n1166 585
R10435 gnd.n1566 gnd.n1166 585
R10436 gnd.n1574 gnd.n1164 585
R10437 gnd.n1575 gnd.n1574 585
R10438 gnd.n5978 gnd.n1163 585
R10439 gnd.n1572 gnd.n1163 585
R10440 gnd.n5979 gnd.n1162 585
R10441 gnd.n1580 gnd.n1162 585
R10442 gnd.n5980 gnd.n1161 585
R10443 gnd.n5280 gnd.n1161 585
R10444 gnd.n5268 gnd.n1159 585
R10445 gnd.n5269 gnd.n5268 585
R10446 gnd.n5984 gnd.n1158 585
R10447 gnd.n1600 gnd.n1158 585
R10448 gnd.n5985 gnd.n1157 585
R10449 gnd.n1609 gnd.n1157 585
R10450 gnd.n5986 gnd.n1156 585
R10451 gnd.n1605 gnd.n1156 585
R10452 gnd.n5242 gnd.n1154 585
R10453 gnd.n5243 gnd.n5242 585
R10454 gnd.n5990 gnd.n1153 585
R10455 gnd.n5234 gnd.n1153 585
R10456 gnd.n5991 gnd.n1152 585
R10457 gnd.n5148 gnd.n1152 585
R10458 gnd.n5992 gnd.n1151 585
R10459 gnd.n5191 gnd.n1151 585
R10460 gnd.n5182 gnd.n1149 585
R10461 gnd.n5183 gnd.n5182 585
R10462 gnd.n5996 gnd.n1148 585
R10463 gnd.n1645 gnd.n1148 585
R10464 gnd.n5997 gnd.n1147 585
R10465 gnd.n1643 gnd.n1147 585
R10466 gnd.n5998 gnd.n1146 585
R10467 gnd.n1649 gnd.n1146 585
R10468 gnd.n1653 gnd.n1144 585
R10469 gnd.n1654 gnd.n1653 585
R10470 gnd.n6002 gnd.n1143 585
R10471 gnd.n1661 gnd.n1143 585
R10472 gnd.n6003 gnd.n1142 585
R10473 gnd.n5026 gnd.n1142 585
R10474 gnd.n6004 gnd.n1141 585
R10475 gnd.n1666 gnd.n1141 585
R10476 gnd.n5102 gnd.n1139 585
R10477 gnd.n5103 gnd.n5102 585
R10478 gnd.n6008 gnd.n1138 585
R10479 gnd.n5091 gnd.n1138 585
R10480 gnd.n6009 gnd.n1137 585
R10481 gnd.n1685 gnd.n1137 585
R10482 gnd.n6010 gnd.n1136 585
R10483 gnd.n1694 gnd.n1136 585
R10484 gnd.n1690 gnd.n1134 585
R10485 gnd.n1691 gnd.n1690 585
R10486 gnd.n6014 gnd.n1133 585
R10487 gnd.n5066 gnd.n1133 585
R10488 gnd.n6015 gnd.n1132 585
R10489 gnd.n5058 gnd.n1132 585
R10490 gnd.n6016 gnd.n1131 585
R10491 gnd.n4944 gnd.n1131 585
R10492 gnd.n5012 gnd.n1129 585
R10493 gnd.n5013 gnd.n5012 585
R10494 gnd.n6020 gnd.n1128 585
R10495 gnd.n5004 gnd.n1128 585
R10496 gnd.n6021 gnd.n1127 585
R10497 gnd.n1729 gnd.n1127 585
R10498 gnd.n6022 gnd.n1126 585
R10499 gnd.n4983 gnd.n1126 585
R10500 gnd.n1733 gnd.n1124 585
R10501 gnd.n1734 gnd.n1733 585
R10502 gnd.n6026 gnd.n1123 585
R10503 gnd.n4974 gnd.n1123 585
R10504 gnd.n6027 gnd.n1122 585
R10505 gnd.n1752 gnd.n1122 585
R10506 gnd.n6028 gnd.n1121 585
R10507 gnd.n4672 gnd.n1121 585
R10508 gnd.n1757 gnd.n1119 585
R10509 gnd.n1758 gnd.n1757 585
R10510 gnd.n6032 gnd.n1118 585
R10511 gnd.n4916 gnd.n1118 585
R10512 gnd.n6033 gnd.n1117 585
R10513 gnd.n4905 gnd.n1117 585
R10514 gnd.n6034 gnd.n1116 585
R10515 gnd.n1772 gnd.n1116 585
R10516 gnd.n4665 gnd.n1114 585
R10517 gnd.n4666 gnd.n4665 585
R10518 gnd.n6038 gnd.n1113 585
R10519 gnd.n4598 gnd.n1113 585
R10520 gnd.n6039 gnd.n1112 585
R10521 gnd.n4655 gnd.n1112 585
R10522 gnd.n6040 gnd.n1111 585
R10523 gnd.n4653 gnd.n1111 585
R10524 gnd.n4650 gnd.n1109 585
R10525 gnd.n4651 gnd.n4650 585
R10526 gnd.n6044 gnd.n1108 585
R10527 gnd.n4604 gnd.n1108 585
R10528 gnd.n6045 gnd.n1107 585
R10529 gnd.n4639 gnd.n1107 585
R10530 gnd.n6046 gnd.n1106 585
R10531 gnd.n4637 gnd.n1106 585
R10532 gnd.n4634 gnd.n1104 585
R10533 gnd.n4635 gnd.n4634 585
R10534 gnd.n6050 gnd.n1103 585
R10535 gnd.n4610 gnd.n1103 585
R10536 gnd.n6051 gnd.n1102 585
R10537 gnd.n4623 gnd.n1102 585
R10538 gnd.n6052 gnd.n1101 585
R10539 gnd.n4621 gnd.n1101 585
R10540 gnd.n4763 gnd.n4762 585
R10541 gnd.n4761 gnd.n4493 585
R10542 gnd.n4495 gnd.n4492 585
R10543 gnd.n4765 gnd.n4492 585
R10544 gnd.n4754 gnd.n4509 585
R10545 gnd.n4753 gnd.n4510 585
R10546 gnd.n4512 gnd.n4511 585
R10547 gnd.n4746 gnd.n4520 585
R10548 gnd.n4745 gnd.n4521 585
R10549 gnd.n4531 gnd.n4522 585
R10550 gnd.n4738 gnd.n4532 585
R10551 gnd.n4737 gnd.n4533 585
R10552 gnd.n4535 gnd.n4534 585
R10553 gnd.n4730 gnd.n4543 585
R10554 gnd.n4729 gnd.n4544 585
R10555 gnd.n4558 gnd.n4545 585
R10556 gnd.n4722 gnd.n4559 585
R10557 gnd.n4721 gnd.n4560 585
R10558 gnd.n4562 gnd.n4561 585
R10559 gnd.n4715 gnd.n4563 585
R10560 gnd.n4714 gnd.n4564 585
R10561 gnd.n4567 gnd.n4565 585
R10562 gnd.n4710 gnd.n4568 585
R10563 gnd.n4709 gnd.n4569 585
R10564 gnd.n4708 gnd.n4570 585
R10565 gnd.n4576 gnd.n4571 585
R10566 gnd.n4704 gnd.n4577 585
R10567 gnd.n4703 gnd.n4578 585
R10568 gnd.n4702 gnd.n4579 585
R10569 gnd.n4582 gnd.n4580 585
R10570 gnd.n5885 gnd.n1228 585
R10571 gnd.n5899 gnd.n1228 585
R10572 gnd.n5884 gnd.n5883 585
R10573 gnd.n5883 gnd.n5882 585
R10574 gnd.n1302 gnd.n1301 585
R10575 gnd.n5869 gnd.n1302 585
R10576 gnd.n5867 gnd.n5866 585
R10577 gnd.n5871 gnd.n5867 585
R10578 gnd.n1310 gnd.n1309 585
R10579 gnd.n1309 gnd.n1308 585
R10580 gnd.n5861 gnd.n5860 585
R10581 gnd.n5860 gnd.n5859 585
R10582 gnd.n1313 gnd.n1312 585
R10583 gnd.n1315 gnd.n1313 585
R10584 gnd.n5846 gnd.n5845 585
R10585 gnd.n5848 gnd.n5846 585
R10586 gnd.n1323 gnd.n1322 585
R10587 gnd.n1322 gnd.n1321 585
R10588 gnd.n5841 gnd.n5840 585
R10589 gnd.n5840 gnd.n5839 585
R10590 gnd.n1326 gnd.n1325 585
R10591 gnd.n1328 gnd.n1326 585
R10592 gnd.n5826 gnd.n5825 585
R10593 gnd.n5828 gnd.n5826 585
R10594 gnd.n1335 gnd.n1334 585
R10595 gnd.n5817 gnd.n1334 585
R10596 gnd.n5821 gnd.n5820 585
R10597 gnd.n5820 gnd.n5819 585
R10598 gnd.n1338 gnd.n1337 585
R10599 gnd.n1380 gnd.n1338 585
R10600 gnd.n5560 gnd.n1388 585
R10601 gnd.n5651 gnd.n1388 585
R10602 gnd.n5559 gnd.n5558 585
R10603 gnd.n5558 gnd.n5557 585
R10604 gnd.n5564 gnd.n5555 585
R10605 gnd.n5555 gnd.n5554 585
R10606 gnd.n5565 gnd.n5552 585
R10607 gnd.n5552 gnd.n1402 585
R10608 gnd.n5566 gnd.n1410 585
R10609 gnd.n5622 gnd.n1410 585
R10610 gnd.n5550 gnd.n1417 585
R10611 gnd.n5611 gnd.n1417 585
R10612 gnd.n5570 gnd.n5549 585
R10613 gnd.n5549 gnd.n5548 585
R10614 gnd.n5571 gnd.n5547 585
R10615 gnd.n5547 gnd.n1430 585
R10616 gnd.n5572 gnd.n5546 585
R10617 gnd.n5546 gnd.n1426 585
R10618 gnd.n1446 gnd.n1437 585
R10619 gnd.n5586 gnd.n1437 585
R10620 gnd.n5577 gnd.n5576 585
R10621 gnd.n5578 gnd.n5577 585
R10622 gnd.n1445 gnd.n1444 585
R10623 gnd.n5471 gnd.n1444 585
R10624 gnd.n5542 gnd.n5541 585
R10625 gnd.n5541 gnd.n5540 585
R10626 gnd.n1449 gnd.n1448 585
R10627 gnd.n5532 gnd.n1449 585
R10628 gnd.n1473 gnd.n1471 585
R10629 gnd.n1471 gnd.n1464 585
R10630 gnd.n5509 gnd.n5508 585
R10631 gnd.n5511 gnd.n5509 585
R10632 gnd.n1472 gnd.n1470 585
R10633 gnd.n1478 gnd.n1470 585
R10634 gnd.n5503 gnd.n5502 585
R10635 gnd.n5502 gnd.n5501 585
R10636 gnd.n1476 gnd.n1475 585
R10637 gnd.n5448 gnd.n1476 585
R10638 gnd.n5382 gnd.n5380 585
R10639 gnd.n5380 gnd.n1486 585
R10640 gnd.n5383 gnd.n5379 585
R10641 gnd.n5379 gnd.n1492 585
R10642 gnd.n5384 gnd.n1501 585
R10643 gnd.n5441 gnd.n1501 585
R10644 gnd.n5377 gnd.n1508 585
R10645 gnd.n5430 gnd.n1508 585
R10646 gnd.n5388 gnd.n5376 585
R10647 gnd.n5376 gnd.n1513 585
R10648 gnd.n5389 gnd.n5375 585
R10649 gnd.n5375 gnd.n1522 585
R10650 gnd.n5390 gnd.n5374 585
R10651 gnd.n5374 gnd.n1518 585
R10652 gnd.n1538 gnd.n1529 585
R10653 gnd.n5405 gnd.n1529 585
R10654 gnd.n5395 gnd.n5394 585
R10655 gnd.n5397 gnd.n5395 585
R10656 gnd.n1537 gnd.n1536 585
R10657 gnd.n5326 gnd.n1536 585
R10658 gnd.n5370 gnd.n5369 585
R10659 gnd.n5369 gnd.n5368 585
R10660 gnd.n1541 gnd.n1540 585
R10661 gnd.n5360 gnd.n1541 585
R10662 gnd.n5211 gnd.n5210 585
R10663 gnd.n5210 gnd.n1558 585
R10664 gnd.n5214 gnd.n5209 585
R10665 gnd.n5209 gnd.n1555 585
R10666 gnd.n5215 gnd.n5208 585
R10667 gnd.n5208 gnd.n1562 585
R10668 gnd.n5216 gnd.n5207 585
R10669 gnd.n5207 gnd.n1566 585
R10670 gnd.n5206 gnd.n5204 585
R10671 gnd.n5206 gnd.n1575 585
R10672 gnd.n5220 gnd.n5203 585
R10673 gnd.n5203 gnd.n1572 585
R10674 gnd.n5221 gnd.n5202 585
R10675 gnd.n5202 gnd.n1580 585
R10676 gnd.n5222 gnd.n1589 585
R10677 gnd.n5280 gnd.n1589 585
R10678 gnd.n5200 gnd.n1596 585
R10679 gnd.n5269 gnd.n1596 585
R10680 gnd.n5226 gnd.n5199 585
R10681 gnd.n5199 gnd.n1600 585
R10682 gnd.n5227 gnd.n5198 585
R10683 gnd.n5198 gnd.n1609 585
R10684 gnd.n5228 gnd.n5197 585
R10685 gnd.n5197 gnd.n1605 585
R10686 gnd.n1625 gnd.n1616 585
R10687 gnd.n5243 gnd.n1616 585
R10688 gnd.n5233 gnd.n5232 585
R10689 gnd.n5234 gnd.n5233 585
R10690 gnd.n1624 gnd.n1623 585
R10691 gnd.n5148 gnd.n1623 585
R10692 gnd.n5193 gnd.n5192 585
R10693 gnd.n5192 gnd.n5191 585
R10694 gnd.n1628 gnd.n1627 585
R10695 gnd.n5183 gnd.n1628 585
R10696 gnd.n5035 gnd.n5034 585
R10697 gnd.n5034 gnd.n1645 585
R10698 gnd.n5038 gnd.n5033 585
R10699 gnd.n5033 gnd.n1643 585
R10700 gnd.n5039 gnd.n5032 585
R10701 gnd.n5032 gnd.n1649 585
R10702 gnd.n5040 gnd.n5031 585
R10703 gnd.n5031 gnd.n1654 585
R10704 gnd.n5030 gnd.n5028 585
R10705 gnd.n5030 gnd.n1661 585
R10706 gnd.n5044 gnd.n5027 585
R10707 gnd.n5027 gnd.n5026 585
R10708 gnd.n5045 gnd.n5024 585
R10709 gnd.n5024 gnd.n1666 585
R10710 gnd.n5046 gnd.n1674 585
R10711 gnd.n5103 gnd.n1674 585
R10712 gnd.n5022 gnd.n1681 585
R10713 gnd.n5091 gnd.n1681 585
R10714 gnd.n5050 gnd.n5021 585
R10715 gnd.n5021 gnd.n1685 585
R10716 gnd.n5051 gnd.n5020 585
R10717 gnd.n5020 gnd.n1694 585
R10718 gnd.n5052 gnd.n5019 585
R10719 gnd.n5019 gnd.n1691 585
R10720 gnd.n1710 gnd.n1701 585
R10721 gnd.n5066 gnd.n1701 585
R10722 gnd.n5057 gnd.n5056 585
R10723 gnd.n5058 gnd.n5057 585
R10724 gnd.n1709 gnd.n1708 585
R10725 gnd.n4944 gnd.n1708 585
R10726 gnd.n5015 gnd.n5014 585
R10727 gnd.n5014 gnd.n5013 585
R10728 gnd.n1713 gnd.n1712 585
R10729 gnd.n5004 gnd.n1713 585
R10730 gnd.n1740 gnd.n1738 585
R10731 gnd.n1738 gnd.n1729 585
R10732 gnd.n4982 gnd.n4981 585
R10733 gnd.n4983 gnd.n4982 585
R10734 gnd.n1739 gnd.n1737 585
R10735 gnd.n1737 gnd.n1734 585
R10736 gnd.n4976 gnd.n4975 585
R10737 gnd.n4975 gnd.n4974 585
R10738 gnd.n1743 gnd.n1742 585
R10739 gnd.n1752 gnd.n1743 585
R10740 gnd.n4674 gnd.n4673 585
R10741 gnd.n4673 gnd.n4672 585
R10742 gnd.n4670 gnd.n4669 585
R10743 gnd.n4670 gnd.n1758 585
R10744 gnd.n4678 gnd.n1766 585
R10745 gnd.n4916 gnd.n1766 585
R10746 gnd.n4679 gnd.n1773 585
R10747 gnd.n4905 gnd.n1773 585
R10748 gnd.n4680 gnd.n4668 585
R10749 gnd.n4668 gnd.n1772 585
R10750 gnd.n4667 gnd.n4596 585
R10751 gnd.n4667 gnd.n4666 585
R10752 gnd.n4684 gnd.n4595 585
R10753 gnd.n4598 gnd.n4595 585
R10754 gnd.n4685 gnd.n4594 585
R10755 gnd.n4655 gnd.n4594 585
R10756 gnd.n4686 gnd.n4593 585
R10757 gnd.n4653 gnd.n4593 585
R10758 gnd.n4649 gnd.n4591 585
R10759 gnd.n4651 gnd.n4649 585
R10760 gnd.n4690 gnd.n4590 585
R10761 gnd.n4604 gnd.n4590 585
R10762 gnd.n4691 gnd.n4589 585
R10763 gnd.n4639 gnd.n4589 585
R10764 gnd.n4692 gnd.n4588 585
R10765 gnd.n4637 gnd.n4588 585
R10766 gnd.n4633 gnd.n4586 585
R10767 gnd.n4635 gnd.n4633 585
R10768 gnd.n4696 gnd.n4585 585
R10769 gnd.n4610 gnd.n4585 585
R10770 gnd.n4697 gnd.n4584 585
R10771 gnd.n4623 gnd.n4584 585
R10772 gnd.n4698 gnd.n4583 585
R10773 gnd.n4621 gnd.n4583 585
R10774 gnd.n5889 gnd.n5888 585
R10775 gnd.n5890 gnd.n5889 585
R10776 gnd.n1266 gnd.n1265 585
R10777 gnd.n1297 gnd.n1296 585
R10778 gnd.n1295 gnd.n1294 585
R10779 gnd.n1292 gnd.n1272 585
R10780 gnd.n1271 gnd.n1270 585
R10781 gnd.n1288 gnd.n1287 585
R10782 gnd.n1286 gnd.n1285 585
R10783 gnd.n1284 gnd.n1276 585
R10784 gnd.n1275 gnd.n1274 585
R10785 gnd.n1279 gnd.n1278 585
R10786 gnd.n1277 gnd.n503 585
R10787 gnd.n7107 gnd.n502 585
R10788 gnd.n7108 gnd.n501 585
R10789 gnd.n1257 gnd.n493 585
R10790 gnd.n7115 gnd.n492 585
R10791 gnd.n7116 gnd.n491 585
R10792 gnd.n1254 gnd.n485 585
R10793 gnd.n7123 gnd.n484 585
R10794 gnd.n7124 gnd.n483 585
R10795 gnd.n1252 gnd.n477 585
R10796 gnd.n7131 gnd.n476 585
R10797 gnd.n7132 gnd.n475 585
R10798 gnd.n1249 gnd.n469 585
R10799 gnd.n7139 gnd.n468 585
R10800 gnd.n7140 gnd.n467 585
R10801 gnd.n1247 gnd.n461 585
R10802 gnd.n7147 gnd.n460 585
R10803 gnd.n7148 gnd.n459 585
R10804 gnd.n3701 gnd.n3700 537.605
R10805 gnd.n5741 gnd.n1383 506.916
R10806 gnd.n5750 gnd.n5749 506.916
R10807 gnd.n4903 gnd.n1774 506.916
R10808 gnd.n4894 gnd.n1763 506.916
R10809 gnd.n1835 gnd.t172 389.64
R10810 gnd.n1374 gnd.t117 389.64
R10811 gnd.n1832 gnd.t124 389.64
R10812 gnd.n5675 gnd.t155 389.64
R10813 gnd.n4573 gnd.t138 371.625
R10814 gnd.n559 gnd.t131 371.625
R10815 gnd.n581 gnd.t113 371.625
R10816 gnd.n201 gnd.t175 371.625
R10817 gnd.n7516 gnd.t89 371.625
R10818 gnd.n122 gnd.t146 371.625
R10819 gnd.n497 gnd.t161 371.625
R10820 gnd.n4552 gnd.t181 371.625
R10821 gnd.n1988 gnd.t184 371.625
R10822 gnd.n1897 gnd.t106 371.625
R10823 gnd.n3731 gnd.t190 371.625
R10824 gnd.n3707 gnd.t168 371.625
R10825 gnd.n4010 gnd.t187 371.625
R10826 gnd.n1268 gnd.t102 371.625
R10827 gnd.n2720 gnd.t193 323.425
R10828 gnd.n2266 gnd.t134 323.425
R10829 gnd.n3568 gnd.n3542 289.615
R10830 gnd.n3536 gnd.n3510 289.615
R10831 gnd.n3504 gnd.n3478 289.615
R10832 gnd.n3473 gnd.n3447 289.615
R10833 gnd.n3441 gnd.n3415 289.615
R10834 gnd.n3409 gnd.n3383 289.615
R10835 gnd.n3377 gnd.n3351 289.615
R10836 gnd.n3346 gnd.n3320 289.615
R10837 gnd.n2794 gnd.t164 279.217
R10838 gnd.n2292 gnd.t142 279.217
R10839 gnd.n1817 gnd.t154 260.649
R10840 gnd.n5667 gnd.t160 260.649
R10841 gnd.n4896 gnd.n4895 256.663
R10842 gnd.n4896 gnd.n1778 256.663
R10843 gnd.n4896 gnd.n1779 256.663
R10844 gnd.n4896 gnd.n1780 256.663
R10845 gnd.n4896 gnd.n1781 256.663
R10846 gnd.n4896 gnd.n1782 256.663
R10847 gnd.n4896 gnd.n1783 256.663
R10848 gnd.n4896 gnd.n1784 256.663
R10849 gnd.n4896 gnd.n1785 256.663
R10850 gnd.n4896 gnd.n1786 256.663
R10851 gnd.n4896 gnd.n1787 256.663
R10852 gnd.n4896 gnd.n1788 256.663
R10853 gnd.n4896 gnd.n1789 256.663
R10854 gnd.n4896 gnd.n1790 256.663
R10855 gnd.n4896 gnd.n1791 256.663
R10856 gnd.n4896 gnd.n1792 256.663
R10857 gnd.n4832 gnd.n4829 256.663
R10858 gnd.n4896 gnd.n1793 256.663
R10859 gnd.n4896 gnd.n1794 256.663
R10860 gnd.n4896 gnd.n1795 256.663
R10861 gnd.n4896 gnd.n1796 256.663
R10862 gnd.n4896 gnd.n1797 256.663
R10863 gnd.n4896 gnd.n1798 256.663
R10864 gnd.n4896 gnd.n1799 256.663
R10865 gnd.n4896 gnd.n1800 256.663
R10866 gnd.n4896 gnd.n1801 256.663
R10867 gnd.n4896 gnd.n1802 256.663
R10868 gnd.n4896 gnd.n1803 256.663
R10869 gnd.n4896 gnd.n1804 256.663
R10870 gnd.n4896 gnd.n1805 256.663
R10871 gnd.n4896 gnd.n1806 256.663
R10872 gnd.n4896 gnd.n1807 256.663
R10873 gnd.n4896 gnd.n1808 256.663
R10874 gnd.n4897 gnd.n4896 256.663
R10875 gnd.n5816 gnd.n1357 256.663
R10876 gnd.n5816 gnd.n1358 256.663
R10877 gnd.n5816 gnd.n1359 256.663
R10878 gnd.n5816 gnd.n1360 256.663
R10879 gnd.n5816 gnd.n1361 256.663
R10880 gnd.n5816 gnd.n1362 256.663
R10881 gnd.n5816 gnd.n1363 256.663
R10882 gnd.n5816 gnd.n1364 256.663
R10883 gnd.n5816 gnd.n1365 256.663
R10884 gnd.n5816 gnd.n1366 256.663
R10885 gnd.n5816 gnd.n1367 256.663
R10886 gnd.n5816 gnd.n1368 256.663
R10887 gnd.n5816 gnd.n1369 256.663
R10888 gnd.n5816 gnd.n1370 256.663
R10889 gnd.n5816 gnd.n1371 256.663
R10890 gnd.n5816 gnd.n1372 256.663
R10891 gnd.n1373 gnd.n556 256.663
R10892 gnd.n5816 gnd.n1356 256.663
R10893 gnd.n5816 gnd.n1355 256.663
R10894 gnd.n5816 gnd.n1354 256.663
R10895 gnd.n5816 gnd.n1353 256.663
R10896 gnd.n5816 gnd.n1352 256.663
R10897 gnd.n5816 gnd.n1351 256.663
R10898 gnd.n5816 gnd.n1350 256.663
R10899 gnd.n5816 gnd.n1349 256.663
R10900 gnd.n5816 gnd.n1348 256.663
R10901 gnd.n5816 gnd.n1347 256.663
R10902 gnd.n5816 gnd.n1346 256.663
R10903 gnd.n5816 gnd.n1345 256.663
R10904 gnd.n5816 gnd.n1344 256.663
R10905 gnd.n5816 gnd.n1343 256.663
R10906 gnd.n5816 gnd.n1342 256.663
R10907 gnd.n5816 gnd.n1341 256.663
R10908 gnd.n5816 gnd.n1340 256.663
R10909 gnd.n4184 gnd.n3701 242.672
R10910 gnd.n4182 gnd.n3701 242.672
R10911 gnd.n4176 gnd.n3701 242.672
R10912 gnd.n4174 gnd.n3701 242.672
R10913 gnd.n4168 gnd.n3701 242.672
R10914 gnd.n4166 gnd.n3701 242.672
R10915 gnd.n4160 gnd.n3701 242.672
R10916 gnd.n4158 gnd.n3701 242.672
R10917 gnd.n4148 gnd.n3701 242.672
R10918 gnd.n2848 gnd.n2847 242.672
R10919 gnd.n2848 gnd.n2758 242.672
R10920 gnd.n2848 gnd.n2759 242.672
R10921 gnd.n2848 gnd.n2760 242.672
R10922 gnd.n2848 gnd.n2761 242.672
R10923 gnd.n2848 gnd.n2762 242.672
R10924 gnd.n2848 gnd.n2763 242.672
R10925 gnd.n2848 gnd.n2764 242.672
R10926 gnd.n2848 gnd.n2765 242.672
R10927 gnd.n2848 gnd.n2766 242.672
R10928 gnd.n2848 gnd.n2767 242.672
R10929 gnd.n2848 gnd.n2768 242.672
R10930 gnd.n2849 gnd.n2848 242.672
R10931 gnd.n3700 gnd.n2241 242.672
R10932 gnd.n3700 gnd.n2240 242.672
R10933 gnd.n3700 gnd.n2239 242.672
R10934 gnd.n3700 gnd.n2238 242.672
R10935 gnd.n3700 gnd.n2237 242.672
R10936 gnd.n3700 gnd.n2236 242.672
R10937 gnd.n3700 gnd.n2235 242.672
R10938 gnd.n3700 gnd.n2234 242.672
R10939 gnd.n3700 gnd.n2233 242.672
R10940 gnd.n3700 gnd.n2232 242.672
R10941 gnd.n3700 gnd.n2231 242.672
R10942 gnd.n3700 gnd.n2230 242.672
R10943 gnd.n3700 gnd.n2229 242.672
R10944 gnd.n2932 gnd.n2931 242.672
R10945 gnd.n2931 gnd.n2670 242.672
R10946 gnd.n2931 gnd.n2671 242.672
R10947 gnd.n2931 gnd.n2672 242.672
R10948 gnd.n2931 gnd.n2673 242.672
R10949 gnd.n2931 gnd.n2674 242.672
R10950 gnd.n2931 gnd.n2675 242.672
R10951 gnd.n2931 gnd.n2676 242.672
R10952 gnd.n3700 gnd.n2242 242.672
R10953 gnd.n3700 gnd.n2243 242.672
R10954 gnd.n3700 gnd.n2244 242.672
R10955 gnd.n3700 gnd.n2245 242.672
R10956 gnd.n3700 gnd.n2246 242.672
R10957 gnd.n3700 gnd.n2247 242.672
R10958 gnd.n3700 gnd.n2248 242.672
R10959 gnd.n3700 gnd.n2249 242.672
R10960 gnd.n3749 gnd.n3701 242.672
R10961 gnd.n3757 gnd.n3701 242.672
R10962 gnd.n3759 gnd.n3701 242.672
R10963 gnd.n3767 gnd.n3701 242.672
R10964 gnd.n3769 gnd.n3701 242.672
R10965 gnd.n3777 gnd.n3701 242.672
R10966 gnd.n3779 gnd.n3701 242.672
R10967 gnd.n3787 gnd.n3701 242.672
R10968 gnd.n3789 gnd.n3701 242.672
R10969 gnd.n3797 gnd.n3701 242.672
R10970 gnd.n3799 gnd.n3701 242.672
R10971 gnd.n3807 gnd.n3701 242.672
R10972 gnd.n3809 gnd.n3701 242.672
R10973 gnd.n3817 gnd.n3701 242.672
R10974 gnd.n3819 gnd.n3701 242.672
R10975 gnd.n3827 gnd.n3701 242.672
R10976 gnd.n3829 gnd.n3701 242.672
R10977 gnd.n3838 gnd.n3701 242.672
R10978 gnd.n3841 gnd.n3701 242.672
R10979 gnd.n6247 gnd.n6246 242.672
R10980 gnd.n6246 gnd.n928 242.672
R10981 gnd.n6246 gnd.n929 242.672
R10982 gnd.n6246 gnd.n930 242.672
R10983 gnd.n6246 gnd.n931 242.672
R10984 gnd.n6246 gnd.n932 242.672
R10985 gnd.n6246 gnd.n933 242.672
R10986 gnd.n6246 gnd.n934 242.672
R10987 gnd.n6246 gnd.n935 242.672
R10988 gnd.n6246 gnd.n936 242.672
R10989 gnd.n6246 gnd.n937 242.672
R10990 gnd.n6246 gnd.n938 242.672
R10991 gnd.n6246 gnd.n939 242.672
R10992 gnd.n6246 gnd.n940 242.672
R10993 gnd.n6246 gnd.n941 242.672
R10994 gnd.n6246 gnd.n942 242.672
R10995 gnd.n6246 gnd.n943 242.672
R10996 gnd.n6246 gnd.n944 242.672
R10997 gnd.n6246 gnd.n945 242.672
R10998 gnd.n6246 gnd.n946 242.672
R10999 gnd.n6246 gnd.n947 242.672
R11000 gnd.n6246 gnd.n948 242.672
R11001 gnd.n6246 gnd.n949 242.672
R11002 gnd.n6246 gnd.n950 242.672
R11003 gnd.n6246 gnd.n951 242.672
R11004 gnd.n6246 gnd.n952 242.672
R11005 gnd.n6246 gnd.n953 242.672
R11006 gnd.n6246 gnd.n954 242.672
R11007 gnd.n6246 gnd.n955 242.672
R11008 gnd.n6246 gnd.n956 242.672
R11009 gnd.n6246 gnd.n957 242.672
R11010 gnd.n6246 gnd.n958 242.672
R11011 gnd.n6246 gnd.n959 242.672
R11012 gnd.n6246 gnd.n960 242.672
R11013 gnd.n6246 gnd.n961 242.672
R11014 gnd.n6246 gnd.n962 242.672
R11015 gnd.n6246 gnd.n963 242.672
R11016 gnd.n6246 gnd.n964 242.672
R11017 gnd.n6246 gnd.n965 242.672
R11018 gnd.n6246 gnd.n966 242.672
R11019 gnd.n6246 gnd.n967 242.672
R11020 gnd.n6246 gnd.n968 242.672
R11021 gnd.n4554 gnd.n1960 242.672
R11022 gnd.n4550 gnd.n1960 242.672
R11023 gnd.n4547 gnd.n1960 242.672
R11024 gnd.n4538 gnd.n1960 242.672
R11025 gnd.n4527 gnd.n1960 242.672
R11026 gnd.n4524 gnd.n1960 242.672
R11027 gnd.n4515 gnd.n1960 242.672
R11028 gnd.n4505 gnd.n1960 242.672
R11029 gnd.n4502 gnd.n1960 242.672
R11030 gnd.n7102 gnd.n525 242.672
R11031 gnd.n7102 gnd.n527 242.672
R11032 gnd.n7102 gnd.n529 242.672
R11033 gnd.n7102 gnd.n530 242.672
R11034 gnd.n7102 gnd.n532 242.672
R11035 gnd.n7102 gnd.n534 242.672
R11036 gnd.n7102 gnd.n535 242.672
R11037 gnd.n7102 gnd.n537 242.672
R11038 gnd.n7102 gnd.n538 242.672
R11039 gnd.n128 gnd.n125 242.672
R11040 gnd.n7427 gnd.n128 242.672
R11041 gnd.n7423 gnd.n128 242.672
R11042 gnd.n7420 gnd.n128 242.672
R11043 gnd.n7415 gnd.n128 242.672
R11044 gnd.n7412 gnd.n128 242.672
R11045 gnd.n7407 gnd.n128 242.672
R11046 gnd.n7404 gnd.n128 242.672
R11047 gnd.n7399 gnd.n128 242.672
R11048 gnd.n4791 gnd.n1960 242.672
R11049 gnd.n1991 gnd.n1960 242.672
R11050 gnd.n4798 gnd.n1960 242.672
R11051 gnd.n1982 gnd.n1960 242.672
R11052 gnd.n4805 gnd.n1960 242.672
R11053 gnd.n1975 gnd.n1960 242.672
R11054 gnd.n4812 gnd.n1960 242.672
R11055 gnd.n1968 gnd.n1960 242.672
R11056 gnd.n4819 gnd.n1960 242.672
R11057 gnd.n4822 gnd.n1960 242.672
R11058 gnd.n1960 gnd.n1904 242.672
R11059 gnd.n4828 gnd.n1899 242.672
R11060 gnd.n1960 gnd.n1905 242.672
R11061 gnd.n1960 gnd.n1906 242.672
R11062 gnd.n1960 gnd.n1907 242.672
R11063 gnd.n1960 gnd.n1908 242.672
R11064 gnd.n1960 gnd.n1909 242.672
R11065 gnd.n1960 gnd.n1910 242.672
R11066 gnd.n1960 gnd.n1911 242.672
R11067 gnd.n1960 gnd.n1912 242.672
R11068 gnd.n7102 gnd.n7101 242.672
R11069 gnd.n7102 gnd.n507 242.672
R11070 gnd.n7102 gnd.n508 242.672
R11071 gnd.n7102 gnd.n509 242.672
R11072 gnd.n7102 gnd.n510 242.672
R11073 gnd.n7102 gnd.n511 242.672
R11074 gnd.n7102 gnd.n512 242.672
R11075 gnd.n7102 gnd.n513 242.672
R11076 gnd.n7071 gnd.n557 242.672
R11077 gnd.n7102 gnd.n514 242.672
R11078 gnd.n7102 gnd.n515 242.672
R11079 gnd.n7102 gnd.n516 242.672
R11080 gnd.n7102 gnd.n517 242.672
R11081 gnd.n7102 gnd.n518 242.672
R11082 gnd.n7102 gnd.n519 242.672
R11083 gnd.n7102 gnd.n520 242.672
R11084 gnd.n7102 gnd.n521 242.672
R11085 gnd.n7102 gnd.n522 242.672
R11086 gnd.n7102 gnd.n523 242.672
R11087 gnd.n7102 gnd.n524 242.672
R11088 gnd.n198 gnd.n128 242.672
R11089 gnd.n7484 gnd.n128 242.672
R11090 gnd.n194 gnd.n128 242.672
R11091 gnd.n7491 gnd.n128 242.672
R11092 gnd.n187 gnd.n128 242.672
R11093 gnd.n7498 gnd.n128 242.672
R11094 gnd.n180 gnd.n128 242.672
R11095 gnd.n7505 gnd.n128 242.672
R11096 gnd.n173 gnd.n128 242.672
R11097 gnd.n7512 gnd.n128 242.672
R11098 gnd.n166 gnd.n128 242.672
R11099 gnd.n7522 gnd.n128 242.672
R11100 gnd.n159 gnd.n128 242.672
R11101 gnd.n7529 gnd.n128 242.672
R11102 gnd.n152 gnd.n128 242.672
R11103 gnd.n7536 gnd.n128 242.672
R11104 gnd.n145 gnd.n128 242.672
R11105 gnd.n7543 gnd.n128 242.672
R11106 gnd.n138 gnd.n128 242.672
R11107 gnd.n4765 gnd.n4764 242.672
R11108 gnd.n4765 gnd.n4478 242.672
R11109 gnd.n4765 gnd.n4479 242.672
R11110 gnd.n4765 gnd.n4480 242.672
R11111 gnd.n4765 gnd.n4481 242.672
R11112 gnd.n4765 gnd.n4482 242.672
R11113 gnd.n4765 gnd.n4483 242.672
R11114 gnd.n4765 gnd.n4484 242.672
R11115 gnd.n4765 gnd.n4485 242.672
R11116 gnd.n4765 gnd.n4486 242.672
R11117 gnd.n4765 gnd.n4487 242.672
R11118 gnd.n4765 gnd.n4488 242.672
R11119 gnd.n4765 gnd.n4489 242.672
R11120 gnd.n4765 gnd.n4490 242.672
R11121 gnd.n5890 gnd.n1264 242.672
R11122 gnd.n5890 gnd.n1263 242.672
R11123 gnd.n5890 gnd.n1262 242.672
R11124 gnd.n5890 gnd.n1261 242.672
R11125 gnd.n5890 gnd.n1260 242.672
R11126 gnd.n5890 gnd.n1259 242.672
R11127 gnd.n5890 gnd.n1258 242.672
R11128 gnd.n5890 gnd.n1256 242.672
R11129 gnd.n5890 gnd.n1255 242.672
R11130 gnd.n5890 gnd.n1253 242.672
R11131 gnd.n5890 gnd.n1251 242.672
R11132 gnd.n5890 gnd.n1250 242.672
R11133 gnd.n5890 gnd.n1248 242.672
R11134 gnd.n5890 gnd.n1246 242.672
R11135 gnd.n135 gnd.n131 240.244
R11136 gnd.n7545 gnd.n7544 240.244
R11137 gnd.n7542 gnd.n139 240.244
R11138 gnd.n7538 gnd.n7537 240.244
R11139 gnd.n7535 gnd.n146 240.244
R11140 gnd.n7531 gnd.n7530 240.244
R11141 gnd.n7528 gnd.n153 240.244
R11142 gnd.n7524 gnd.n7523 240.244
R11143 gnd.n7521 gnd.n160 240.244
R11144 gnd.n7514 gnd.n7513 240.244
R11145 gnd.n7511 gnd.n167 240.244
R11146 gnd.n7507 gnd.n7506 240.244
R11147 gnd.n7504 gnd.n174 240.244
R11148 gnd.n7500 gnd.n7499 240.244
R11149 gnd.n7497 gnd.n181 240.244
R11150 gnd.n7493 gnd.n7492 240.244
R11151 gnd.n7490 gnd.n188 240.244
R11152 gnd.n7486 gnd.n7485 240.244
R11153 gnd.n7483 gnd.n195 240.244
R11154 gnd.n585 gnd.n451 240.244
R11155 gnd.n585 gnd.n443 240.244
R11156 gnd.n7023 gnd.n443 240.244
R11157 gnd.n7023 gnd.n435 240.244
R11158 gnd.n6815 gnd.n435 240.244
R11159 gnd.n6815 gnd.n426 240.244
R11160 gnd.n6819 gnd.n426 240.244
R11161 gnd.n6819 gnd.n417 240.244
R11162 gnd.n6954 gnd.n417 240.244
R11163 gnd.n6954 gnd.n409 240.244
R11164 gnd.n6950 gnd.n409 240.244
R11165 gnd.n6950 gnd.n402 240.244
R11166 gnd.n6947 gnd.n402 240.244
R11167 gnd.n6947 gnd.n394 240.244
R11168 gnd.n6944 gnd.n394 240.244
R11169 gnd.n6944 gnd.n385 240.244
R11170 gnd.n6941 gnd.n385 240.244
R11171 gnd.n6941 gnd.n377 240.244
R11172 gnd.n6938 gnd.n377 240.244
R11173 gnd.n6938 gnd.n370 240.244
R11174 gnd.n6935 gnd.n370 240.244
R11175 gnd.n6935 gnd.n362 240.244
R11176 gnd.n6932 gnd.n362 240.244
R11177 gnd.n6932 gnd.n353 240.244
R11178 gnd.n6929 gnd.n353 240.244
R11179 gnd.n6929 gnd.n345 240.244
R11180 gnd.n6926 gnd.n345 240.244
R11181 gnd.n6926 gnd.n338 240.244
R11182 gnd.n6923 gnd.n338 240.244
R11183 gnd.n6923 gnd.n330 240.244
R11184 gnd.n6920 gnd.n330 240.244
R11185 gnd.n6920 gnd.n320 240.244
R11186 gnd.n6917 gnd.n320 240.244
R11187 gnd.n6917 gnd.n312 240.244
R11188 gnd.n6914 gnd.n312 240.244
R11189 gnd.n6914 gnd.n305 240.244
R11190 gnd.n6911 gnd.n305 240.244
R11191 gnd.n6911 gnd.n299 240.244
R11192 gnd.n6908 gnd.n299 240.244
R11193 gnd.n6908 gnd.n290 240.244
R11194 gnd.n6905 gnd.n290 240.244
R11195 gnd.n6905 gnd.n282 240.244
R11196 gnd.n6902 gnd.n282 240.244
R11197 gnd.n6902 gnd.n275 240.244
R11198 gnd.n6899 gnd.n275 240.244
R11199 gnd.n6899 gnd.n269 240.244
R11200 gnd.n6896 gnd.n269 240.244
R11201 gnd.n6896 gnd.n260 240.244
R11202 gnd.n6893 gnd.n260 240.244
R11203 gnd.n6893 gnd.n252 240.244
R11204 gnd.n6890 gnd.n252 240.244
R11205 gnd.n6890 gnd.n245 240.244
R11206 gnd.n6887 gnd.n245 240.244
R11207 gnd.n6887 gnd.n239 240.244
R11208 gnd.n6884 gnd.n239 240.244
R11209 gnd.n6884 gnd.n230 240.244
R11210 gnd.n6881 gnd.n230 240.244
R11211 gnd.n6881 gnd.n223 240.244
R11212 gnd.n6878 gnd.n223 240.244
R11213 gnd.n6878 gnd.n214 240.244
R11214 gnd.n214 gnd.n205 240.244
R11215 gnd.n7474 gnd.n205 240.244
R11216 gnd.n7475 gnd.n7474 240.244
R11217 gnd.n7475 gnd.n127 240.244
R11218 gnd.n7100 gnd.n539 240.244
R11219 gnd.n7096 gnd.n539 240.244
R11220 gnd.n7094 gnd.n7093 240.244
R11221 gnd.n7090 gnd.n7089 240.244
R11222 gnd.n7086 gnd.n7085 240.244
R11223 gnd.n7082 gnd.n7081 240.244
R11224 gnd.n7078 gnd.n7077 240.244
R11225 gnd.n7074 gnd.n7073 240.244
R11226 gnd.n7069 gnd.n7068 240.244
R11227 gnd.n7065 gnd.n7064 240.244
R11228 gnd.n7061 gnd.n7060 240.244
R11229 gnd.n7057 gnd.n7056 240.244
R11230 gnd.n7053 gnd.n7052 240.244
R11231 gnd.n7049 gnd.n7048 240.244
R11232 gnd.n7045 gnd.n7044 240.244
R11233 gnd.n7041 gnd.n7040 240.244
R11234 gnd.n7037 gnd.n7036 240.244
R11235 gnd.n580 gnd.n579 240.244
R11236 gnd.n7158 gnd.n446 240.244
R11237 gnd.n7164 gnd.n446 240.244
R11238 gnd.n7164 gnd.n433 240.244
R11239 gnd.n7174 gnd.n433 240.244
R11240 gnd.n7174 gnd.n429 240.244
R11241 gnd.n7180 gnd.n429 240.244
R11242 gnd.n7180 gnd.n415 240.244
R11243 gnd.n7190 gnd.n415 240.244
R11244 gnd.n7190 gnd.n411 240.244
R11245 gnd.n7196 gnd.n411 240.244
R11246 gnd.n7196 gnd.n400 240.244
R11247 gnd.n7206 gnd.n400 240.244
R11248 gnd.n7206 gnd.n396 240.244
R11249 gnd.n7212 gnd.n396 240.244
R11250 gnd.n7212 gnd.n383 240.244
R11251 gnd.n7222 gnd.n383 240.244
R11252 gnd.n7222 gnd.n379 240.244
R11253 gnd.n7228 gnd.n379 240.244
R11254 gnd.n7228 gnd.n368 240.244
R11255 gnd.n7238 gnd.n368 240.244
R11256 gnd.n7238 gnd.n364 240.244
R11257 gnd.n7244 gnd.n364 240.244
R11258 gnd.n7244 gnd.n351 240.244
R11259 gnd.n7254 gnd.n351 240.244
R11260 gnd.n7254 gnd.n347 240.244
R11261 gnd.n7260 gnd.n347 240.244
R11262 gnd.n7260 gnd.n336 240.244
R11263 gnd.n7270 gnd.n336 240.244
R11264 gnd.n7270 gnd.n332 240.244
R11265 gnd.n7276 gnd.n332 240.244
R11266 gnd.n7276 gnd.n318 240.244
R11267 gnd.n7286 gnd.n318 240.244
R11268 gnd.n7286 gnd.n314 240.244
R11269 gnd.n7292 gnd.n314 240.244
R11270 gnd.n7292 gnd.n304 240.244
R11271 gnd.n7302 gnd.n304 240.244
R11272 gnd.n7302 gnd.n300 240.244
R11273 gnd.n7308 gnd.n300 240.244
R11274 gnd.n7308 gnd.n288 240.244
R11275 gnd.n7318 gnd.n288 240.244
R11276 gnd.n7318 gnd.n284 240.244
R11277 gnd.n7324 gnd.n284 240.244
R11278 gnd.n7324 gnd.n274 240.244
R11279 gnd.n7334 gnd.n274 240.244
R11280 gnd.n7334 gnd.n270 240.244
R11281 gnd.n7340 gnd.n270 240.244
R11282 gnd.n7340 gnd.n258 240.244
R11283 gnd.n7350 gnd.n258 240.244
R11284 gnd.n7350 gnd.n254 240.244
R11285 gnd.n7356 gnd.n254 240.244
R11286 gnd.n7356 gnd.n244 240.244
R11287 gnd.n7366 gnd.n244 240.244
R11288 gnd.n7366 gnd.n240 240.244
R11289 gnd.n7372 gnd.n240 240.244
R11290 gnd.n7372 gnd.n228 240.244
R11291 gnd.n7382 gnd.n228 240.244
R11292 gnd.n7382 gnd.n224 240.244
R11293 gnd.n7388 gnd.n224 240.244
R11294 gnd.n7388 gnd.n212 240.244
R11295 gnd.n7466 gnd.n212 240.244
R11296 gnd.n7466 gnd.n208 240.244
R11297 gnd.n7472 gnd.n208 240.244
R11298 gnd.n7472 gnd.n130 240.244
R11299 gnd.n7552 gnd.n130 240.244
R11300 gnd.n7398 gnd.n7397 240.244
R11301 gnd.n7403 gnd.n7400 240.244
R11302 gnd.n7406 gnd.n7405 240.244
R11303 gnd.n7411 gnd.n7408 240.244
R11304 gnd.n7414 gnd.n7413 240.244
R11305 gnd.n7419 gnd.n7416 240.244
R11306 gnd.n7422 gnd.n7421 240.244
R11307 gnd.n7426 gnd.n7424 240.244
R11308 gnd.n7429 gnd.n7428 240.244
R11309 gnd.n6801 gnd.n452 240.244
R11310 gnd.n6801 gnd.n444 240.244
R11311 gnd.n7021 gnd.n444 240.244
R11312 gnd.n7021 gnd.n436 240.244
R11313 gnd.n6806 gnd.n436 240.244
R11314 gnd.n6806 gnd.n427 240.244
R11315 gnd.n6807 gnd.n427 240.244
R11316 gnd.n6807 gnd.n418 240.244
R11317 gnd.n6956 gnd.n418 240.244
R11318 gnd.n6956 gnd.n410 240.244
R11319 gnd.n6957 gnd.n410 240.244
R11320 gnd.n6957 gnd.n403 240.244
R11321 gnd.n6960 gnd.n403 240.244
R11322 gnd.n6960 gnd.n395 240.244
R11323 gnd.n6961 gnd.n395 240.244
R11324 gnd.n6961 gnd.n386 240.244
R11325 gnd.n6964 gnd.n386 240.244
R11326 gnd.n6964 gnd.n378 240.244
R11327 gnd.n6965 gnd.n378 240.244
R11328 gnd.n6965 gnd.n371 240.244
R11329 gnd.n6968 gnd.n371 240.244
R11330 gnd.n6968 gnd.n363 240.244
R11331 gnd.n6969 gnd.n363 240.244
R11332 gnd.n6969 gnd.n354 240.244
R11333 gnd.n6972 gnd.n354 240.244
R11334 gnd.n6972 gnd.n346 240.244
R11335 gnd.n6973 gnd.n346 240.244
R11336 gnd.n6973 gnd.n339 240.244
R11337 gnd.n6976 gnd.n339 240.244
R11338 gnd.n6976 gnd.n331 240.244
R11339 gnd.n6977 gnd.n331 240.244
R11340 gnd.n6977 gnd.n321 240.244
R11341 gnd.n321 gnd.n82 240.244
R11342 gnd.n83 gnd.n82 240.244
R11343 gnd.n84 gnd.n83 240.244
R11344 gnd.n306 gnd.n84 240.244
R11345 gnd.n306 gnd.n87 240.244
R11346 gnd.n88 gnd.n87 240.244
R11347 gnd.n89 gnd.n88 240.244
R11348 gnd.n291 gnd.n89 240.244
R11349 gnd.n291 gnd.n92 240.244
R11350 gnd.n93 gnd.n92 240.244
R11351 gnd.n94 gnd.n93 240.244
R11352 gnd.n276 gnd.n94 240.244
R11353 gnd.n276 gnd.n97 240.244
R11354 gnd.n98 gnd.n97 240.244
R11355 gnd.n99 gnd.n98 240.244
R11356 gnd.n261 gnd.n99 240.244
R11357 gnd.n261 gnd.n102 240.244
R11358 gnd.n103 gnd.n102 240.244
R11359 gnd.n104 gnd.n103 240.244
R11360 gnd.n246 gnd.n104 240.244
R11361 gnd.n246 gnd.n107 240.244
R11362 gnd.n108 gnd.n107 240.244
R11363 gnd.n109 gnd.n108 240.244
R11364 gnd.n231 gnd.n109 240.244
R11365 gnd.n231 gnd.n112 240.244
R11366 gnd.n113 gnd.n112 240.244
R11367 gnd.n114 gnd.n113 240.244
R11368 gnd.n215 gnd.n114 240.244
R11369 gnd.n215 gnd.n117 240.244
R11370 gnd.n118 gnd.n117 240.244
R11371 gnd.n119 gnd.n118 240.244
R11372 gnd.n7554 gnd.n119 240.244
R11373 gnd.n526 gnd.n456 240.244
R11374 gnd.n464 gnd.n463 240.244
R11375 gnd.n528 gnd.n471 240.244
R11376 gnd.n531 gnd.n472 240.244
R11377 gnd.n480 gnd.n479 240.244
R11378 gnd.n533 gnd.n487 240.244
R11379 gnd.n536 gnd.n488 240.244
R11380 gnd.n496 gnd.n495 240.244
R11381 gnd.n7103 gnd.n505 240.244
R11382 gnd.n7156 gnd.n442 240.244
R11383 gnd.n7166 gnd.n442 240.244
R11384 gnd.n7166 gnd.n438 240.244
R11385 gnd.n7172 gnd.n438 240.244
R11386 gnd.n7172 gnd.n424 240.244
R11387 gnd.n7182 gnd.n424 240.244
R11388 gnd.n7182 gnd.n420 240.244
R11389 gnd.n7188 gnd.n420 240.244
R11390 gnd.n7188 gnd.n408 240.244
R11391 gnd.n7198 gnd.n408 240.244
R11392 gnd.n7198 gnd.n404 240.244
R11393 gnd.n7204 gnd.n404 240.244
R11394 gnd.n7204 gnd.n392 240.244
R11395 gnd.n7214 gnd.n392 240.244
R11396 gnd.n7214 gnd.n388 240.244
R11397 gnd.n7220 gnd.n388 240.244
R11398 gnd.n7220 gnd.n376 240.244
R11399 gnd.n7230 gnd.n376 240.244
R11400 gnd.n7230 gnd.n372 240.244
R11401 gnd.n7236 gnd.n372 240.244
R11402 gnd.n7236 gnd.n360 240.244
R11403 gnd.n7246 gnd.n360 240.244
R11404 gnd.n7246 gnd.n356 240.244
R11405 gnd.n7252 gnd.n356 240.244
R11406 gnd.n7252 gnd.n344 240.244
R11407 gnd.n7262 gnd.n344 240.244
R11408 gnd.n7262 gnd.n340 240.244
R11409 gnd.n7268 gnd.n340 240.244
R11410 gnd.n7268 gnd.n328 240.244
R11411 gnd.n7278 gnd.n328 240.244
R11412 gnd.n7278 gnd.n323 240.244
R11413 gnd.n7284 gnd.n323 240.244
R11414 gnd.n7284 gnd.n311 240.244
R11415 gnd.n7294 gnd.n311 240.244
R11416 gnd.n7294 gnd.n307 240.244
R11417 gnd.n7300 gnd.n307 240.244
R11418 gnd.n7300 gnd.n297 240.244
R11419 gnd.n7310 gnd.n297 240.244
R11420 gnd.n7310 gnd.n293 240.244
R11421 gnd.n7316 gnd.n293 240.244
R11422 gnd.n7316 gnd.n281 240.244
R11423 gnd.n7326 gnd.n281 240.244
R11424 gnd.n7326 gnd.n277 240.244
R11425 gnd.n7332 gnd.n277 240.244
R11426 gnd.n7332 gnd.n267 240.244
R11427 gnd.n7342 gnd.n267 240.244
R11428 gnd.n7342 gnd.n263 240.244
R11429 gnd.n7348 gnd.n263 240.244
R11430 gnd.n7348 gnd.n251 240.244
R11431 gnd.n7358 gnd.n251 240.244
R11432 gnd.n7358 gnd.n247 240.244
R11433 gnd.n7364 gnd.n247 240.244
R11434 gnd.n7364 gnd.n237 240.244
R11435 gnd.n7374 gnd.n237 240.244
R11436 gnd.n7374 gnd.n233 240.244
R11437 gnd.n7380 gnd.n233 240.244
R11438 gnd.n7380 gnd.n222 240.244
R11439 gnd.n7390 gnd.n222 240.244
R11440 gnd.n7390 gnd.n216 240.244
R11441 gnd.n7464 gnd.n216 240.244
R11442 gnd.n7464 gnd.n217 240.244
R11443 gnd.n217 gnd.n207 240.244
R11444 gnd.n7395 gnd.n207 240.244
R11445 gnd.n7395 gnd.n129 240.244
R11446 gnd.n6254 gnd.n922 240.244
R11447 gnd.n6254 gnd.n920 240.244
R11448 gnd.n6258 gnd.n920 240.244
R11449 gnd.n6258 gnd.n916 240.244
R11450 gnd.n6264 gnd.n916 240.244
R11451 gnd.n6264 gnd.n914 240.244
R11452 gnd.n6268 gnd.n914 240.244
R11453 gnd.n6268 gnd.n910 240.244
R11454 gnd.n6274 gnd.n910 240.244
R11455 gnd.n6274 gnd.n908 240.244
R11456 gnd.n6278 gnd.n908 240.244
R11457 gnd.n6278 gnd.n904 240.244
R11458 gnd.n6284 gnd.n904 240.244
R11459 gnd.n6284 gnd.n902 240.244
R11460 gnd.n6288 gnd.n902 240.244
R11461 gnd.n6288 gnd.n898 240.244
R11462 gnd.n6294 gnd.n898 240.244
R11463 gnd.n6294 gnd.n896 240.244
R11464 gnd.n6298 gnd.n896 240.244
R11465 gnd.n6298 gnd.n892 240.244
R11466 gnd.n6304 gnd.n892 240.244
R11467 gnd.n6304 gnd.n890 240.244
R11468 gnd.n6308 gnd.n890 240.244
R11469 gnd.n6308 gnd.n886 240.244
R11470 gnd.n6314 gnd.n886 240.244
R11471 gnd.n6314 gnd.n884 240.244
R11472 gnd.n6318 gnd.n884 240.244
R11473 gnd.n6318 gnd.n880 240.244
R11474 gnd.n6324 gnd.n880 240.244
R11475 gnd.n6324 gnd.n878 240.244
R11476 gnd.n6328 gnd.n878 240.244
R11477 gnd.n6328 gnd.n874 240.244
R11478 gnd.n6334 gnd.n874 240.244
R11479 gnd.n6334 gnd.n872 240.244
R11480 gnd.n6338 gnd.n872 240.244
R11481 gnd.n6338 gnd.n868 240.244
R11482 gnd.n6344 gnd.n868 240.244
R11483 gnd.n6344 gnd.n866 240.244
R11484 gnd.n6348 gnd.n866 240.244
R11485 gnd.n6348 gnd.n862 240.244
R11486 gnd.n6354 gnd.n862 240.244
R11487 gnd.n6354 gnd.n860 240.244
R11488 gnd.n6358 gnd.n860 240.244
R11489 gnd.n6358 gnd.n856 240.244
R11490 gnd.n6364 gnd.n856 240.244
R11491 gnd.n6364 gnd.n854 240.244
R11492 gnd.n6368 gnd.n854 240.244
R11493 gnd.n6368 gnd.n850 240.244
R11494 gnd.n6374 gnd.n850 240.244
R11495 gnd.n6374 gnd.n848 240.244
R11496 gnd.n6378 gnd.n848 240.244
R11497 gnd.n6378 gnd.n844 240.244
R11498 gnd.n6384 gnd.n844 240.244
R11499 gnd.n6384 gnd.n842 240.244
R11500 gnd.n6388 gnd.n842 240.244
R11501 gnd.n6388 gnd.n838 240.244
R11502 gnd.n6394 gnd.n838 240.244
R11503 gnd.n6394 gnd.n836 240.244
R11504 gnd.n6398 gnd.n836 240.244
R11505 gnd.n6398 gnd.n832 240.244
R11506 gnd.n6404 gnd.n832 240.244
R11507 gnd.n6404 gnd.n830 240.244
R11508 gnd.n6408 gnd.n830 240.244
R11509 gnd.n6408 gnd.n826 240.244
R11510 gnd.n6414 gnd.n826 240.244
R11511 gnd.n6414 gnd.n824 240.244
R11512 gnd.n6418 gnd.n824 240.244
R11513 gnd.n6418 gnd.n820 240.244
R11514 gnd.n6424 gnd.n820 240.244
R11515 gnd.n6424 gnd.n818 240.244
R11516 gnd.n6428 gnd.n818 240.244
R11517 gnd.n6428 gnd.n814 240.244
R11518 gnd.n6434 gnd.n814 240.244
R11519 gnd.n6434 gnd.n812 240.244
R11520 gnd.n6438 gnd.n812 240.244
R11521 gnd.n6438 gnd.n808 240.244
R11522 gnd.n6444 gnd.n808 240.244
R11523 gnd.n6444 gnd.n806 240.244
R11524 gnd.n6448 gnd.n806 240.244
R11525 gnd.n6448 gnd.n802 240.244
R11526 gnd.n6454 gnd.n802 240.244
R11527 gnd.n6454 gnd.n800 240.244
R11528 gnd.n6458 gnd.n800 240.244
R11529 gnd.n6458 gnd.n796 240.244
R11530 gnd.n6464 gnd.n796 240.244
R11531 gnd.n6464 gnd.n794 240.244
R11532 gnd.n6468 gnd.n794 240.244
R11533 gnd.n6468 gnd.n790 240.244
R11534 gnd.n6474 gnd.n790 240.244
R11535 gnd.n6474 gnd.n788 240.244
R11536 gnd.n6478 gnd.n788 240.244
R11537 gnd.n6478 gnd.n784 240.244
R11538 gnd.n6484 gnd.n784 240.244
R11539 gnd.n6484 gnd.n782 240.244
R11540 gnd.n6488 gnd.n782 240.244
R11541 gnd.n6488 gnd.n778 240.244
R11542 gnd.n6494 gnd.n778 240.244
R11543 gnd.n6494 gnd.n776 240.244
R11544 gnd.n6498 gnd.n776 240.244
R11545 gnd.n6498 gnd.n772 240.244
R11546 gnd.n6504 gnd.n772 240.244
R11547 gnd.n6504 gnd.n770 240.244
R11548 gnd.n6508 gnd.n770 240.244
R11549 gnd.n6508 gnd.n766 240.244
R11550 gnd.n6514 gnd.n766 240.244
R11551 gnd.n6514 gnd.n764 240.244
R11552 gnd.n6518 gnd.n764 240.244
R11553 gnd.n6518 gnd.n760 240.244
R11554 gnd.n6524 gnd.n760 240.244
R11555 gnd.n6524 gnd.n758 240.244
R11556 gnd.n6528 gnd.n758 240.244
R11557 gnd.n6528 gnd.n754 240.244
R11558 gnd.n6534 gnd.n754 240.244
R11559 gnd.n6534 gnd.n752 240.244
R11560 gnd.n6538 gnd.n752 240.244
R11561 gnd.n6538 gnd.n748 240.244
R11562 gnd.n6544 gnd.n748 240.244
R11563 gnd.n6544 gnd.n746 240.244
R11564 gnd.n6548 gnd.n746 240.244
R11565 gnd.n6548 gnd.n742 240.244
R11566 gnd.n6554 gnd.n742 240.244
R11567 gnd.n6554 gnd.n740 240.244
R11568 gnd.n6558 gnd.n740 240.244
R11569 gnd.n6558 gnd.n736 240.244
R11570 gnd.n6565 gnd.n736 240.244
R11571 gnd.n6565 gnd.n734 240.244
R11572 gnd.n6569 gnd.n734 240.244
R11573 gnd.n6569 gnd.n731 240.244
R11574 gnd.n6575 gnd.n729 240.244
R11575 gnd.n6579 gnd.n729 240.244
R11576 gnd.n6579 gnd.n725 240.244
R11577 gnd.n6585 gnd.n725 240.244
R11578 gnd.n6585 gnd.n723 240.244
R11579 gnd.n6589 gnd.n723 240.244
R11580 gnd.n6589 gnd.n719 240.244
R11581 gnd.n6595 gnd.n719 240.244
R11582 gnd.n6595 gnd.n717 240.244
R11583 gnd.n6599 gnd.n717 240.244
R11584 gnd.n6599 gnd.n713 240.244
R11585 gnd.n6605 gnd.n713 240.244
R11586 gnd.n6605 gnd.n711 240.244
R11587 gnd.n6609 gnd.n711 240.244
R11588 gnd.n6609 gnd.n707 240.244
R11589 gnd.n6615 gnd.n707 240.244
R11590 gnd.n6615 gnd.n705 240.244
R11591 gnd.n6619 gnd.n705 240.244
R11592 gnd.n6619 gnd.n701 240.244
R11593 gnd.n6625 gnd.n701 240.244
R11594 gnd.n6625 gnd.n699 240.244
R11595 gnd.n6629 gnd.n699 240.244
R11596 gnd.n6629 gnd.n695 240.244
R11597 gnd.n6635 gnd.n695 240.244
R11598 gnd.n6635 gnd.n693 240.244
R11599 gnd.n6639 gnd.n693 240.244
R11600 gnd.n6639 gnd.n689 240.244
R11601 gnd.n6645 gnd.n689 240.244
R11602 gnd.n6645 gnd.n687 240.244
R11603 gnd.n6649 gnd.n687 240.244
R11604 gnd.n6649 gnd.n683 240.244
R11605 gnd.n6655 gnd.n683 240.244
R11606 gnd.n6655 gnd.n681 240.244
R11607 gnd.n6659 gnd.n681 240.244
R11608 gnd.n6659 gnd.n677 240.244
R11609 gnd.n6665 gnd.n677 240.244
R11610 gnd.n6665 gnd.n675 240.244
R11611 gnd.n6669 gnd.n675 240.244
R11612 gnd.n6669 gnd.n671 240.244
R11613 gnd.n6675 gnd.n671 240.244
R11614 gnd.n6675 gnd.n669 240.244
R11615 gnd.n6679 gnd.n669 240.244
R11616 gnd.n6679 gnd.n665 240.244
R11617 gnd.n6685 gnd.n665 240.244
R11618 gnd.n6685 gnd.n663 240.244
R11619 gnd.n6689 gnd.n663 240.244
R11620 gnd.n6689 gnd.n659 240.244
R11621 gnd.n6695 gnd.n659 240.244
R11622 gnd.n6695 gnd.n657 240.244
R11623 gnd.n6699 gnd.n657 240.244
R11624 gnd.n6699 gnd.n653 240.244
R11625 gnd.n6705 gnd.n653 240.244
R11626 gnd.n6705 gnd.n651 240.244
R11627 gnd.n6709 gnd.n651 240.244
R11628 gnd.n6709 gnd.n647 240.244
R11629 gnd.n6715 gnd.n647 240.244
R11630 gnd.n6715 gnd.n645 240.244
R11631 gnd.n6719 gnd.n645 240.244
R11632 gnd.n6719 gnd.n641 240.244
R11633 gnd.n6725 gnd.n641 240.244
R11634 gnd.n6725 gnd.n639 240.244
R11635 gnd.n6729 gnd.n639 240.244
R11636 gnd.n6729 gnd.n635 240.244
R11637 gnd.n6735 gnd.n635 240.244
R11638 gnd.n6735 gnd.n633 240.244
R11639 gnd.n6739 gnd.n633 240.244
R11640 gnd.n6739 gnd.n629 240.244
R11641 gnd.n6745 gnd.n629 240.244
R11642 gnd.n6745 gnd.n627 240.244
R11643 gnd.n6749 gnd.n627 240.244
R11644 gnd.n6749 gnd.n623 240.244
R11645 gnd.n6755 gnd.n623 240.244
R11646 gnd.n6755 gnd.n621 240.244
R11647 gnd.n6759 gnd.n621 240.244
R11648 gnd.n6759 gnd.n617 240.244
R11649 gnd.n6765 gnd.n617 240.244
R11650 gnd.n6765 gnd.n615 240.244
R11651 gnd.n6769 gnd.n615 240.244
R11652 gnd.n6769 gnd.n611 240.244
R11653 gnd.n6775 gnd.n611 240.244
R11654 gnd.n6775 gnd.n609 240.244
R11655 gnd.n6781 gnd.n609 240.244
R11656 gnd.n6781 gnd.n605 240.244
R11657 gnd.n6787 gnd.n605 240.244
R11658 gnd.n6080 gnd.n1054 240.244
R11659 gnd.n4460 gnd.n1054 240.244
R11660 gnd.n4460 gnd.n4455 240.244
R11661 gnd.n4466 gnd.n4455 240.244
R11662 gnd.n4467 gnd.n4466 240.244
R11663 gnd.n4468 gnd.n4467 240.244
R11664 gnd.n4468 gnd.n4450 240.244
R11665 gnd.n4772 gnd.n4450 240.244
R11666 gnd.n4772 gnd.n4451 240.244
R11667 gnd.n4768 gnd.n4451 240.244
R11668 gnd.n4768 gnd.n4476 240.244
R11669 gnd.n4618 gnd.n4476 240.244
R11670 gnd.n4619 gnd.n4618 240.244
R11671 gnd.n4625 gnd.n4619 240.244
R11672 gnd.n4625 gnd.n4611 240.244
R11673 gnd.n4631 gnd.n4611 240.244
R11674 gnd.n4631 gnd.n4609 240.244
R11675 gnd.n4641 gnd.n4609 240.244
R11676 gnd.n4641 gnd.n4605 240.244
R11677 gnd.n4647 gnd.n4605 240.244
R11678 gnd.n4647 gnd.n4603 240.244
R11679 gnd.n4657 gnd.n4603 240.244
R11680 gnd.n4657 gnd.n4599 240.244
R11681 gnd.n4663 gnd.n4599 240.244
R11682 gnd.n4663 gnd.n1771 240.244
R11683 gnd.n4907 gnd.n1771 240.244
R11684 gnd.n4907 gnd.n1767 240.244
R11685 gnd.n4913 gnd.n1767 240.244
R11686 gnd.n4913 gnd.n1750 240.244
R11687 gnd.n4966 gnd.n1750 240.244
R11688 gnd.n4966 gnd.n1746 240.244
R11689 gnd.n4972 gnd.n1746 240.244
R11690 gnd.n4972 gnd.n1727 240.244
R11691 gnd.n4994 gnd.n1727 240.244
R11692 gnd.n4994 gnd.n1722 240.244
R11693 gnd.n5002 gnd.n1722 240.244
R11694 gnd.n5002 gnd.n1723 240.244
R11695 gnd.n1723 gnd.n1699 240.244
R11696 gnd.n5068 gnd.n1699 240.244
R11697 gnd.n5068 gnd.n1695 240.244
R11698 gnd.n5074 gnd.n1695 240.244
R11699 gnd.n5074 gnd.n1679 240.244
R11700 gnd.n5093 gnd.n1679 240.244
R11701 gnd.n5093 gnd.n1675 240.244
R11702 gnd.n5099 gnd.n1675 240.244
R11703 gnd.n5099 gnd.n1659 240.244
R11704 gnd.n5127 gnd.n1659 240.244
R11705 gnd.n5127 gnd.n1655 240.244
R11706 gnd.n5133 gnd.n1655 240.244
R11707 gnd.n5133 gnd.n1642 240.244
R11708 gnd.n5172 gnd.n1642 240.244
R11709 gnd.n5172 gnd.n1637 240.244
R11710 gnd.n5180 gnd.n1637 240.244
R11711 gnd.n5180 gnd.n1638 240.244
R11712 gnd.n1638 gnd.n1614 240.244
R11713 gnd.n5245 gnd.n1614 240.244
R11714 gnd.n5245 gnd.n1610 240.244
R11715 gnd.n5251 gnd.n1610 240.244
R11716 gnd.n5251 gnd.n1594 240.244
R11717 gnd.n5271 gnd.n1594 240.244
R11718 gnd.n5271 gnd.n1590 240.244
R11719 gnd.n5277 gnd.n1590 240.244
R11720 gnd.n5277 gnd.n1571 240.244
R11721 gnd.n5304 gnd.n1571 240.244
R11722 gnd.n5304 gnd.n1567 240.244
R11723 gnd.n5310 gnd.n1567 240.244
R11724 gnd.n5310 gnd.n1554 240.244
R11725 gnd.n5350 gnd.n1554 240.244
R11726 gnd.n5350 gnd.n1549 240.244
R11727 gnd.n5358 gnd.n1549 240.244
R11728 gnd.n5358 gnd.n1550 240.244
R11729 gnd.n1550 gnd.n1527 240.244
R11730 gnd.n5407 gnd.n1527 240.244
R11731 gnd.n5407 gnd.n1523 240.244
R11732 gnd.n5413 gnd.n1523 240.244
R11733 gnd.n5413 gnd.n1506 240.244
R11734 gnd.n5432 gnd.n1506 240.244
R11735 gnd.n5432 gnd.n1502 240.244
R11736 gnd.n5438 gnd.n1502 240.244
R11737 gnd.n5438 gnd.n1484 240.244
R11738 gnd.n5493 gnd.n1484 240.244
R11739 gnd.n5493 gnd.n1480 240.244
R11740 gnd.n5499 gnd.n1480 240.244
R11741 gnd.n5499 gnd.n1462 240.244
R11742 gnd.n5522 gnd.n1462 240.244
R11743 gnd.n5522 gnd.n1457 240.244
R11744 gnd.n5530 gnd.n1457 240.244
R11745 gnd.n5530 gnd.n1458 240.244
R11746 gnd.n1458 gnd.n1435 240.244
R11747 gnd.n5588 gnd.n1435 240.244
R11748 gnd.n5588 gnd.n1431 240.244
R11749 gnd.n5594 gnd.n1431 240.244
R11750 gnd.n5594 gnd.n1415 240.244
R11751 gnd.n5613 gnd.n1415 240.244
R11752 gnd.n5613 gnd.n1411 240.244
R11753 gnd.n5619 gnd.n1411 240.244
R11754 gnd.n5619 gnd.n1395 240.244
R11755 gnd.n5641 gnd.n1395 240.244
R11756 gnd.n5641 gnd.n1390 240.244
R11757 gnd.n5649 gnd.n1390 240.244
R11758 gnd.n5649 gnd.n1391 240.244
R11759 gnd.n1391 gnd.n1333 240.244
R11760 gnd.n5830 gnd.n1333 240.244
R11761 gnd.n5830 gnd.n1329 240.244
R11762 gnd.n5836 gnd.n1329 240.244
R11763 gnd.n5836 gnd.n1320 240.244
R11764 gnd.n5850 gnd.n1320 240.244
R11765 gnd.n5850 gnd.n1316 240.244
R11766 gnd.n5856 gnd.n1316 240.244
R11767 gnd.n5856 gnd.n1307 240.244
R11768 gnd.n5873 gnd.n1307 240.244
R11769 gnd.n5873 gnd.n1303 240.244
R11770 gnd.n5880 gnd.n1303 240.244
R11771 gnd.n5880 gnd.n1230 240.244
R11772 gnd.n5897 gnd.n1230 240.244
R11773 gnd.n5897 gnd.n1231 240.244
R11774 gnd.n5893 gnd.n1231 240.244
R11775 gnd.n5893 gnd.n1245 240.244
R11776 gnd.n1245 gnd.n1244 240.244
R11777 gnd.n1244 gnd.n1237 240.244
R11778 gnd.n1237 gnd.n593 240.244
R11779 gnd.n6798 gnd.n593 240.244
R11780 gnd.n6798 gnd.n594 240.244
R11781 gnd.n6794 gnd.n594 240.244
R11782 gnd.n6794 gnd.n6793 240.244
R11783 gnd.n6793 gnd.n6792 240.244
R11784 gnd.n6792 gnd.n600 240.244
R11785 gnd.n6788 gnd.n600 240.244
R11786 gnd.n6245 gnd.n926 240.244
R11787 gnd.n6245 gnd.n970 240.244
R11788 gnd.n6241 gnd.n6240 240.244
R11789 gnd.n6237 gnd.n6236 240.244
R11790 gnd.n6233 gnd.n6232 240.244
R11791 gnd.n6229 gnd.n6228 240.244
R11792 gnd.n6225 gnd.n6224 240.244
R11793 gnd.n6221 gnd.n6220 240.244
R11794 gnd.n6217 gnd.n6216 240.244
R11795 gnd.n6213 gnd.n6212 240.244
R11796 gnd.n6209 gnd.n6208 240.244
R11797 gnd.n6205 gnd.n6204 240.244
R11798 gnd.n6201 gnd.n6200 240.244
R11799 gnd.n6197 gnd.n6196 240.244
R11800 gnd.n6193 gnd.n6192 240.244
R11801 gnd.n6189 gnd.n6188 240.244
R11802 gnd.n6185 gnd.n6184 240.244
R11803 gnd.n6181 gnd.n6180 240.244
R11804 gnd.n6177 gnd.n6176 240.244
R11805 gnd.n6173 gnd.n6172 240.244
R11806 gnd.n6169 gnd.n6168 240.244
R11807 gnd.n6165 gnd.n6164 240.244
R11808 gnd.n6161 gnd.n6160 240.244
R11809 gnd.n6157 gnd.n6156 240.244
R11810 gnd.n6153 gnd.n6152 240.244
R11811 gnd.n6149 gnd.n6148 240.244
R11812 gnd.n6145 gnd.n6144 240.244
R11813 gnd.n6141 gnd.n6140 240.244
R11814 gnd.n6137 gnd.n6136 240.244
R11815 gnd.n6133 gnd.n6132 240.244
R11816 gnd.n6129 gnd.n6128 240.244
R11817 gnd.n6125 gnd.n6124 240.244
R11818 gnd.n6121 gnd.n6120 240.244
R11819 gnd.n6117 gnd.n6116 240.244
R11820 gnd.n6113 gnd.n6112 240.244
R11821 gnd.n6109 gnd.n6108 240.244
R11822 gnd.n6105 gnd.n6104 240.244
R11823 gnd.n6101 gnd.n6100 240.244
R11824 gnd.n6097 gnd.n6096 240.244
R11825 gnd.n6093 gnd.n6092 240.244
R11826 gnd.n6089 gnd.n6088 240.244
R11827 gnd.n6085 gnd.n6084 240.244
R11828 gnd.n1959 gnd.n1913 240.244
R11829 gnd.n1955 gnd.n1954 240.244
R11830 gnd.n1951 gnd.n1950 240.244
R11831 gnd.n1947 gnd.n1946 240.244
R11832 gnd.n1943 gnd.n1942 240.244
R11833 gnd.n1939 gnd.n1938 240.244
R11834 gnd.n1935 gnd.n1934 240.244
R11835 gnd.n1931 gnd.n1930 240.244
R11836 gnd.n4823 gnd.n1903 240.244
R11837 gnd.n4821 gnd.n4820 240.244
R11838 gnd.n4818 gnd.n1962 240.244
R11839 gnd.n4814 gnd.n4813 240.244
R11840 gnd.n4811 gnd.n1969 240.244
R11841 gnd.n4807 gnd.n4806 240.244
R11842 gnd.n4804 gnd.n1976 240.244
R11843 gnd.n4800 gnd.n4799 240.244
R11844 gnd.n4797 gnd.n1983 240.244
R11845 gnd.n4793 gnd.n4792 240.244
R11846 gnd.n3984 gnd.n3702 240.244
R11847 gnd.n3984 gnd.n2221 240.244
R11848 gnd.n3978 gnd.n2221 240.244
R11849 gnd.n3978 gnd.n2214 240.244
R11850 gnd.n3975 gnd.n2214 240.244
R11851 gnd.n3975 gnd.n2206 240.244
R11852 gnd.n3972 gnd.n2206 240.244
R11853 gnd.n3972 gnd.n2197 240.244
R11854 gnd.n3969 gnd.n2197 240.244
R11855 gnd.n3969 gnd.n2189 240.244
R11856 gnd.n3966 gnd.n2189 240.244
R11857 gnd.n3966 gnd.n2182 240.244
R11858 gnd.n3963 gnd.n2182 240.244
R11859 gnd.n3963 gnd.n2174 240.244
R11860 gnd.n3960 gnd.n2174 240.244
R11861 gnd.n3960 gnd.n2165 240.244
R11862 gnd.n3957 gnd.n2165 240.244
R11863 gnd.n3957 gnd.n2157 240.244
R11864 gnd.n3954 gnd.n2157 240.244
R11865 gnd.n3954 gnd.n2150 240.244
R11866 gnd.n3951 gnd.n2150 240.244
R11867 gnd.n3951 gnd.n2142 240.244
R11868 gnd.n3948 gnd.n2142 240.244
R11869 gnd.n3948 gnd.n2133 240.244
R11870 gnd.n3945 gnd.n2133 240.244
R11871 gnd.n3945 gnd.n2125 240.244
R11872 gnd.n3942 gnd.n2125 240.244
R11873 gnd.n3942 gnd.n2118 240.244
R11874 gnd.n3939 gnd.n2118 240.244
R11875 gnd.n3939 gnd.n2110 240.244
R11876 gnd.n3936 gnd.n2110 240.244
R11877 gnd.n3936 gnd.n2100 240.244
R11878 gnd.n3933 gnd.n2100 240.244
R11879 gnd.n3933 gnd.n2091 240.244
R11880 gnd.n3930 gnd.n2091 240.244
R11881 gnd.n3930 gnd.n2084 240.244
R11882 gnd.n3927 gnd.n2084 240.244
R11883 gnd.n3927 gnd.n2077 240.244
R11884 gnd.n3924 gnd.n2077 240.244
R11885 gnd.n3924 gnd.n2068 240.244
R11886 gnd.n3921 gnd.n2068 240.244
R11887 gnd.n3921 gnd.n2059 240.244
R11888 gnd.n3918 gnd.n2059 240.244
R11889 gnd.n3918 gnd.n2052 240.244
R11890 gnd.n3915 gnd.n2052 240.244
R11891 gnd.n3915 gnd.n2045 240.244
R11892 gnd.n3912 gnd.n2045 240.244
R11893 gnd.n3912 gnd.n2036 240.244
R11894 gnd.n3909 gnd.n2036 240.244
R11895 gnd.n3909 gnd.n2027 240.244
R11896 gnd.n3906 gnd.n2027 240.244
R11897 gnd.n3906 gnd.n2019 240.244
R11898 gnd.n3903 gnd.n2019 240.244
R11899 gnd.n3903 gnd.n2011 240.244
R11900 gnd.n3900 gnd.n2011 240.244
R11901 gnd.n3900 gnd.n3899 240.244
R11902 gnd.n3899 gnd.n1057 240.244
R11903 gnd.n4435 gnd.n1057 240.244
R11904 gnd.n4435 gnd.n1069 240.244
R11905 gnd.n4442 gnd.n1069 240.244
R11906 gnd.n4442 gnd.n1081 240.244
R11907 gnd.n4783 gnd.n1081 240.244
R11908 gnd.n4783 gnd.n1092 240.244
R11909 gnd.n1992 gnd.n1092 240.244
R11910 gnd.n3750 gnd.n3746 240.244
R11911 gnd.n3756 gnd.n3746 240.244
R11912 gnd.n3760 gnd.n3758 240.244
R11913 gnd.n3766 gnd.n3742 240.244
R11914 gnd.n3770 gnd.n3768 240.244
R11915 gnd.n3776 gnd.n3738 240.244
R11916 gnd.n3780 gnd.n3778 240.244
R11917 gnd.n3786 gnd.n3734 240.244
R11918 gnd.n3790 gnd.n3788 240.244
R11919 gnd.n3796 gnd.n3727 240.244
R11920 gnd.n3800 gnd.n3798 240.244
R11921 gnd.n3806 gnd.n3723 240.244
R11922 gnd.n3810 gnd.n3808 240.244
R11923 gnd.n3816 gnd.n3719 240.244
R11924 gnd.n3820 gnd.n3818 240.244
R11925 gnd.n3826 gnd.n3715 240.244
R11926 gnd.n3830 gnd.n3828 240.244
R11927 gnd.n3837 gnd.n3711 240.244
R11928 gnd.n3840 gnd.n3839 240.244
R11929 gnd.n4193 gnd.n2223 240.244
R11930 gnd.n4199 gnd.n2223 240.244
R11931 gnd.n4199 gnd.n2212 240.244
R11932 gnd.n4209 gnd.n2212 240.244
R11933 gnd.n4209 gnd.n2208 240.244
R11934 gnd.n4215 gnd.n2208 240.244
R11935 gnd.n4215 gnd.n2195 240.244
R11936 gnd.n4225 gnd.n2195 240.244
R11937 gnd.n4225 gnd.n2191 240.244
R11938 gnd.n4231 gnd.n2191 240.244
R11939 gnd.n4231 gnd.n2180 240.244
R11940 gnd.n4241 gnd.n2180 240.244
R11941 gnd.n4241 gnd.n2176 240.244
R11942 gnd.n4247 gnd.n2176 240.244
R11943 gnd.n4247 gnd.n2163 240.244
R11944 gnd.n4257 gnd.n2163 240.244
R11945 gnd.n4257 gnd.n2159 240.244
R11946 gnd.n4263 gnd.n2159 240.244
R11947 gnd.n4263 gnd.n2148 240.244
R11948 gnd.n4273 gnd.n2148 240.244
R11949 gnd.n4273 gnd.n2144 240.244
R11950 gnd.n4279 gnd.n2144 240.244
R11951 gnd.n4279 gnd.n2131 240.244
R11952 gnd.n4289 gnd.n2131 240.244
R11953 gnd.n4289 gnd.n2127 240.244
R11954 gnd.n4295 gnd.n2127 240.244
R11955 gnd.n4295 gnd.n2116 240.244
R11956 gnd.n4305 gnd.n2116 240.244
R11957 gnd.n4305 gnd.n2112 240.244
R11958 gnd.n4311 gnd.n2112 240.244
R11959 gnd.n4311 gnd.n2098 240.244
R11960 gnd.n4321 gnd.n2098 240.244
R11961 gnd.n4321 gnd.n2094 240.244
R11962 gnd.n4327 gnd.n2094 240.244
R11963 gnd.n4327 gnd.n2083 240.244
R11964 gnd.n4337 gnd.n2083 240.244
R11965 gnd.n4337 gnd.n2079 240.244
R11966 gnd.n4343 gnd.n2079 240.244
R11967 gnd.n4343 gnd.n2066 240.244
R11968 gnd.n4353 gnd.n2066 240.244
R11969 gnd.n4353 gnd.n2062 240.244
R11970 gnd.n4359 gnd.n2062 240.244
R11971 gnd.n4359 gnd.n2051 240.244
R11972 gnd.n4369 gnd.n2051 240.244
R11973 gnd.n4369 gnd.n2047 240.244
R11974 gnd.n4375 gnd.n2047 240.244
R11975 gnd.n4375 gnd.n2034 240.244
R11976 gnd.n4385 gnd.n2034 240.244
R11977 gnd.n4385 gnd.n2030 240.244
R11978 gnd.n4391 gnd.n2030 240.244
R11979 gnd.n4391 gnd.n2018 240.244
R11980 gnd.n4414 gnd.n2018 240.244
R11981 gnd.n4414 gnd.n2013 240.244
R11982 gnd.n4423 gnd.n2013 240.244
R11983 gnd.n4423 gnd.n2014 240.244
R11984 gnd.n2014 gnd.n1060 240.244
R11985 gnd.n6077 gnd.n1060 240.244
R11986 gnd.n6077 gnd.n1061 240.244
R11987 gnd.n6073 gnd.n1061 240.244
R11988 gnd.n6073 gnd.n1067 240.244
R11989 gnd.n6065 gnd.n1067 240.244
R11990 gnd.n6065 gnd.n1084 240.244
R11991 gnd.n6061 gnd.n1084 240.244
R11992 gnd.n6061 gnd.n1090 240.244
R11993 gnd.n3699 gnd.n2251 240.244
R11994 gnd.n3692 gnd.n3691 240.244
R11995 gnd.n3689 gnd.n3688 240.244
R11996 gnd.n3685 gnd.n3684 240.244
R11997 gnd.n3681 gnd.n3680 240.244
R11998 gnd.n3677 gnd.n3676 240.244
R11999 gnd.n3673 gnd.n3672 240.244
R12000 gnd.n3669 gnd.n3668 240.244
R12001 gnd.n2943 gnd.n2655 240.244
R12002 gnd.n2953 gnd.n2655 240.244
R12003 gnd.n2953 gnd.n2646 240.244
R12004 gnd.n2646 gnd.n2635 240.244
R12005 gnd.n2974 gnd.n2635 240.244
R12006 gnd.n2974 gnd.n2629 240.244
R12007 gnd.n2984 gnd.n2629 240.244
R12008 gnd.n2984 gnd.n2618 240.244
R12009 gnd.n2618 gnd.n2610 240.244
R12010 gnd.n3002 gnd.n2610 240.244
R12011 gnd.n3003 gnd.n3002 240.244
R12012 gnd.n3003 gnd.n2595 240.244
R12013 gnd.n3005 gnd.n2595 240.244
R12014 gnd.n3005 gnd.n2581 240.244
R12015 gnd.n3047 gnd.n2581 240.244
R12016 gnd.n3048 gnd.n3047 240.244
R12017 gnd.n3051 gnd.n3048 240.244
R12018 gnd.n3051 gnd.n2536 240.244
R12019 gnd.n2576 gnd.n2536 240.244
R12020 gnd.n2576 gnd.n2546 240.244
R12021 gnd.n3061 gnd.n2546 240.244
R12022 gnd.n3061 gnd.n2567 240.244
R12023 gnd.n3071 gnd.n2567 240.244
R12024 gnd.n3071 gnd.n2453 240.244
R12025 gnd.n3116 gnd.n2453 240.244
R12026 gnd.n3116 gnd.n2439 240.244
R12027 gnd.n3138 gnd.n2439 240.244
R12028 gnd.n3139 gnd.n3138 240.244
R12029 gnd.n3139 gnd.n2426 240.244
R12030 gnd.n2426 gnd.n2415 240.244
R12031 gnd.n3170 gnd.n2415 240.244
R12032 gnd.n3171 gnd.n3170 240.244
R12033 gnd.n3172 gnd.n3171 240.244
R12034 gnd.n3172 gnd.n2400 240.244
R12035 gnd.n2400 gnd.n2399 240.244
R12036 gnd.n2399 gnd.n2384 240.244
R12037 gnd.n3223 gnd.n2384 240.244
R12038 gnd.n3224 gnd.n3223 240.244
R12039 gnd.n3224 gnd.n2371 240.244
R12040 gnd.n2371 gnd.n2360 240.244
R12041 gnd.n3255 gnd.n2360 240.244
R12042 gnd.n3256 gnd.n3255 240.244
R12043 gnd.n3257 gnd.n3256 240.244
R12044 gnd.n3257 gnd.n2344 240.244
R12045 gnd.n2344 gnd.n2343 240.244
R12046 gnd.n2343 gnd.n2330 240.244
R12047 gnd.n3312 gnd.n2330 240.244
R12048 gnd.n3313 gnd.n3312 240.244
R12049 gnd.n3313 gnd.n2317 240.244
R12050 gnd.n2317 gnd.n2307 240.244
R12051 gnd.n3600 gnd.n2307 240.244
R12052 gnd.n3603 gnd.n3600 240.244
R12053 gnd.n3603 gnd.n3602 240.244
R12054 gnd.n2933 gnd.n2668 240.244
R12055 gnd.n2689 gnd.n2668 240.244
R12056 gnd.n2692 gnd.n2691 240.244
R12057 gnd.n2699 gnd.n2698 240.244
R12058 gnd.n2702 gnd.n2701 240.244
R12059 gnd.n2709 gnd.n2708 240.244
R12060 gnd.n2712 gnd.n2711 240.244
R12061 gnd.n2719 gnd.n2718 240.244
R12062 gnd.n2941 gnd.n2665 240.244
R12063 gnd.n2665 gnd.n2644 240.244
R12064 gnd.n2964 gnd.n2644 240.244
R12065 gnd.n2964 gnd.n2638 240.244
R12066 gnd.n2972 gnd.n2638 240.244
R12067 gnd.n2972 gnd.n2640 240.244
R12068 gnd.n2640 gnd.n2616 240.244
R12069 gnd.n2994 gnd.n2616 240.244
R12070 gnd.n2994 gnd.n2612 240.244
R12071 gnd.n3000 gnd.n2612 240.244
R12072 gnd.n3000 gnd.n2594 240.244
R12073 gnd.n3025 gnd.n2594 240.244
R12074 gnd.n3025 gnd.n2589 240.244
R12075 gnd.n3037 gnd.n2589 240.244
R12076 gnd.n3037 gnd.n2590 240.244
R12077 gnd.n3033 gnd.n2590 240.244
R12078 gnd.n3033 gnd.n2538 240.244
R12079 gnd.n3085 gnd.n2538 240.244
R12080 gnd.n3085 gnd.n2539 240.244
R12081 gnd.n3081 gnd.n2539 240.244
R12082 gnd.n3081 gnd.n2545 240.244
R12083 gnd.n2565 gnd.n2545 240.244
R12084 gnd.n2565 gnd.n2451 240.244
R12085 gnd.n3120 gnd.n2451 240.244
R12086 gnd.n3120 gnd.n2446 240.244
R12087 gnd.n3128 gnd.n2446 240.244
R12088 gnd.n3128 gnd.n2447 240.244
R12089 gnd.n2447 gnd.n2424 240.244
R12090 gnd.n3160 gnd.n2424 240.244
R12091 gnd.n3160 gnd.n2419 240.244
R12092 gnd.n3168 gnd.n2419 240.244
R12093 gnd.n3168 gnd.n2420 240.244
R12094 gnd.n2420 gnd.n2397 240.244
R12095 gnd.n3205 gnd.n2397 240.244
R12096 gnd.n3205 gnd.n2392 240.244
R12097 gnd.n3213 gnd.n2392 240.244
R12098 gnd.n3213 gnd.n2393 240.244
R12099 gnd.n2393 gnd.n2369 240.244
R12100 gnd.n3245 gnd.n2369 240.244
R12101 gnd.n3245 gnd.n2364 240.244
R12102 gnd.n3253 gnd.n2364 240.244
R12103 gnd.n3253 gnd.n2365 240.244
R12104 gnd.n2365 gnd.n2342 240.244
R12105 gnd.n3294 gnd.n2342 240.244
R12106 gnd.n3294 gnd.n2337 240.244
R12107 gnd.n3302 gnd.n2337 240.244
R12108 gnd.n3302 gnd.n2338 240.244
R12109 gnd.n2338 gnd.n2315 240.244
R12110 gnd.n3588 gnd.n2315 240.244
R12111 gnd.n3588 gnd.n2310 240.244
R12112 gnd.n3598 gnd.n2310 240.244
R12113 gnd.n3598 gnd.n2311 240.244
R12114 gnd.n2311 gnd.n2250 240.244
R12115 gnd.n2270 gnd.n2228 240.244
R12116 gnd.n3659 gnd.n3658 240.244
R12117 gnd.n3655 gnd.n3654 240.244
R12118 gnd.n3651 gnd.n3650 240.244
R12119 gnd.n3647 gnd.n3646 240.244
R12120 gnd.n3643 gnd.n3642 240.244
R12121 gnd.n3639 gnd.n3638 240.244
R12122 gnd.n3635 gnd.n3634 240.244
R12123 gnd.n3631 gnd.n3630 240.244
R12124 gnd.n3627 gnd.n3626 240.244
R12125 gnd.n3623 gnd.n3622 240.244
R12126 gnd.n3619 gnd.n3618 240.244
R12127 gnd.n3615 gnd.n3614 240.244
R12128 gnd.n2856 gnd.n2753 240.244
R12129 gnd.n2856 gnd.n2746 240.244
R12130 gnd.n2867 gnd.n2746 240.244
R12131 gnd.n2867 gnd.n2742 240.244
R12132 gnd.n2873 gnd.n2742 240.244
R12133 gnd.n2873 gnd.n2734 240.244
R12134 gnd.n2883 gnd.n2734 240.244
R12135 gnd.n2883 gnd.n2729 240.244
R12136 gnd.n2919 gnd.n2729 240.244
R12137 gnd.n2919 gnd.n2730 240.244
R12138 gnd.n2730 gnd.n2677 240.244
R12139 gnd.n2914 gnd.n2677 240.244
R12140 gnd.n2914 gnd.n2913 240.244
R12141 gnd.n2913 gnd.n2656 240.244
R12142 gnd.n2909 gnd.n2656 240.244
R12143 gnd.n2909 gnd.n2647 240.244
R12144 gnd.n2906 gnd.n2647 240.244
R12145 gnd.n2906 gnd.n2905 240.244
R12146 gnd.n2905 gnd.n2630 240.244
R12147 gnd.n2901 gnd.n2630 240.244
R12148 gnd.n2901 gnd.n2619 240.244
R12149 gnd.n2619 gnd.n2600 240.244
R12150 gnd.n3014 gnd.n2600 240.244
R12151 gnd.n3014 gnd.n2596 240.244
R12152 gnd.n3022 gnd.n2596 240.244
R12153 gnd.n3022 gnd.n2587 240.244
R12154 gnd.n2587 gnd.n2523 240.244
R12155 gnd.n3094 gnd.n2523 240.244
R12156 gnd.n3094 gnd.n2524 240.244
R12157 gnd.n2535 gnd.n2524 240.244
R12158 gnd.n2570 gnd.n2535 240.244
R12159 gnd.n2573 gnd.n2570 240.244
R12160 gnd.n2573 gnd.n2547 240.244
R12161 gnd.n2560 gnd.n2547 240.244
R12162 gnd.n2560 gnd.n2557 240.244
R12163 gnd.n2557 gnd.n2454 240.244
R12164 gnd.n3115 gnd.n2454 240.244
R12165 gnd.n3115 gnd.n2444 240.244
R12166 gnd.n3111 gnd.n2444 240.244
R12167 gnd.n3111 gnd.n2438 240.244
R12168 gnd.n3108 gnd.n2438 240.244
R12169 gnd.n3108 gnd.n2427 240.244
R12170 gnd.n3105 gnd.n2427 240.244
R12171 gnd.n3105 gnd.n2405 240.244
R12172 gnd.n3181 gnd.n2405 240.244
R12173 gnd.n3181 gnd.n2401 240.244
R12174 gnd.n3202 gnd.n2401 240.244
R12175 gnd.n3202 gnd.n2390 240.244
R12176 gnd.n3198 gnd.n2390 240.244
R12177 gnd.n3198 gnd.n2383 240.244
R12178 gnd.n3195 gnd.n2383 240.244
R12179 gnd.n3195 gnd.n2372 240.244
R12180 gnd.n3192 gnd.n2372 240.244
R12181 gnd.n3192 gnd.n2349 240.244
R12182 gnd.n3266 gnd.n2349 240.244
R12183 gnd.n3266 gnd.n2345 240.244
R12184 gnd.n3291 gnd.n2345 240.244
R12185 gnd.n3291 gnd.n2336 240.244
R12186 gnd.n3287 gnd.n2336 240.244
R12187 gnd.n3287 gnd.n2329 240.244
R12188 gnd.n3283 gnd.n2329 240.244
R12189 gnd.n3283 gnd.n2318 240.244
R12190 gnd.n3280 gnd.n2318 240.244
R12191 gnd.n3280 gnd.n2299 240.244
R12192 gnd.n3610 gnd.n2299 240.244
R12193 gnd.n2770 gnd.n2769 240.244
R12194 gnd.n2841 gnd.n2769 240.244
R12195 gnd.n2839 gnd.n2838 240.244
R12196 gnd.n2835 gnd.n2834 240.244
R12197 gnd.n2831 gnd.n2830 240.244
R12198 gnd.n2827 gnd.n2826 240.244
R12199 gnd.n2823 gnd.n2822 240.244
R12200 gnd.n2819 gnd.n2818 240.244
R12201 gnd.n2815 gnd.n2814 240.244
R12202 gnd.n2811 gnd.n2810 240.244
R12203 gnd.n2807 gnd.n2806 240.244
R12204 gnd.n2803 gnd.n2802 240.244
R12205 gnd.n2799 gnd.n2757 240.244
R12206 gnd.n2859 gnd.n2751 240.244
R12207 gnd.n2859 gnd.n2747 240.244
R12208 gnd.n2865 gnd.n2747 240.244
R12209 gnd.n2865 gnd.n2740 240.244
R12210 gnd.n2875 gnd.n2740 240.244
R12211 gnd.n2875 gnd.n2736 240.244
R12212 gnd.n2881 gnd.n2736 240.244
R12213 gnd.n2881 gnd.n2727 240.244
R12214 gnd.n2921 gnd.n2727 240.244
R12215 gnd.n2921 gnd.n2678 240.244
R12216 gnd.n2929 gnd.n2678 240.244
R12217 gnd.n2929 gnd.n2679 240.244
R12218 gnd.n2679 gnd.n2657 240.244
R12219 gnd.n2950 gnd.n2657 240.244
R12220 gnd.n2950 gnd.n2649 240.244
R12221 gnd.n2961 gnd.n2649 240.244
R12222 gnd.n2961 gnd.n2650 240.244
R12223 gnd.n2650 gnd.n2631 240.244
R12224 gnd.n2981 gnd.n2631 240.244
R12225 gnd.n2981 gnd.n2621 240.244
R12226 gnd.n2991 gnd.n2621 240.244
R12227 gnd.n2991 gnd.n2602 240.244
R12228 gnd.n3012 gnd.n2602 240.244
R12229 gnd.n3012 gnd.n2604 240.244
R12230 gnd.n2604 gnd.n2585 240.244
R12231 gnd.n3040 gnd.n2585 240.244
R12232 gnd.n3040 gnd.n2527 240.244
R12233 gnd.n3092 gnd.n2527 240.244
R12234 gnd.n3092 gnd.n2528 240.244
R12235 gnd.n3088 gnd.n2528 240.244
R12236 gnd.n3088 gnd.n2534 240.244
R12237 gnd.n2549 gnd.n2534 240.244
R12238 gnd.n3078 gnd.n2549 240.244
R12239 gnd.n3078 gnd.n2550 240.244
R12240 gnd.n3074 gnd.n2550 240.244
R12241 gnd.n3074 gnd.n2556 240.244
R12242 gnd.n2556 gnd.n2443 240.244
R12243 gnd.n3131 gnd.n2443 240.244
R12244 gnd.n3131 gnd.n2436 240.244
R12245 gnd.n3142 gnd.n2436 240.244
R12246 gnd.n3142 gnd.n2429 240.244
R12247 gnd.n3157 gnd.n2429 240.244
R12248 gnd.n3157 gnd.n2430 240.244
R12249 gnd.n2430 gnd.n2408 240.244
R12250 gnd.n3179 gnd.n2408 240.244
R12251 gnd.n3179 gnd.n2409 240.244
R12252 gnd.n2409 gnd.n2388 240.244
R12253 gnd.n3216 gnd.n2388 240.244
R12254 gnd.n3216 gnd.n2381 240.244
R12255 gnd.n3227 gnd.n2381 240.244
R12256 gnd.n3227 gnd.n2374 240.244
R12257 gnd.n3242 gnd.n2374 240.244
R12258 gnd.n3242 gnd.n2375 240.244
R12259 gnd.n2375 gnd.n2352 240.244
R12260 gnd.n3264 gnd.n2352 240.244
R12261 gnd.n3264 gnd.n2354 240.244
R12262 gnd.n2354 gnd.n2334 240.244
R12263 gnd.n3305 gnd.n2334 240.244
R12264 gnd.n3305 gnd.n2327 240.244
R12265 gnd.n3316 gnd.n2327 240.244
R12266 gnd.n3316 gnd.n2320 240.244
R12267 gnd.n3585 gnd.n2320 240.244
R12268 gnd.n3585 gnd.n2321 240.244
R12269 gnd.n2321 gnd.n2302 240.244
R12270 gnd.n3608 gnd.n2302 240.244
R12271 gnd.n4501 gnd.n4499 240.244
R12272 gnd.n4504 gnd.n4503 240.244
R12273 gnd.n4514 gnd.n4506 240.244
R12274 gnd.n4517 gnd.n4516 240.244
R12275 gnd.n4526 gnd.n4525 240.244
R12276 gnd.n4537 gnd.n4528 240.244
R12277 gnd.n4540 gnd.n4539 240.244
R12278 gnd.n4549 gnd.n4548 240.244
R12279 gnd.n4555 gnd.n4551 240.244
R12280 gnd.n4144 gnd.n3703 240.244
R12281 gnd.n4144 gnd.n2222 240.244
R12282 gnd.n4141 gnd.n2222 240.244
R12283 gnd.n4141 gnd.n2215 240.244
R12284 gnd.n4138 gnd.n2215 240.244
R12285 gnd.n4138 gnd.n2207 240.244
R12286 gnd.n4135 gnd.n2207 240.244
R12287 gnd.n4135 gnd.n2198 240.244
R12288 gnd.n4132 gnd.n2198 240.244
R12289 gnd.n4132 gnd.n2190 240.244
R12290 gnd.n4129 gnd.n2190 240.244
R12291 gnd.n4129 gnd.n2183 240.244
R12292 gnd.n4126 gnd.n2183 240.244
R12293 gnd.n4126 gnd.n2175 240.244
R12294 gnd.n4123 gnd.n2175 240.244
R12295 gnd.n4123 gnd.n2166 240.244
R12296 gnd.n4120 gnd.n2166 240.244
R12297 gnd.n4120 gnd.n2158 240.244
R12298 gnd.n4117 gnd.n2158 240.244
R12299 gnd.n4117 gnd.n2151 240.244
R12300 gnd.n4114 gnd.n2151 240.244
R12301 gnd.n4114 gnd.n2143 240.244
R12302 gnd.n4111 gnd.n2143 240.244
R12303 gnd.n4111 gnd.n2134 240.244
R12304 gnd.n4108 gnd.n2134 240.244
R12305 gnd.n4108 gnd.n2126 240.244
R12306 gnd.n4105 gnd.n2126 240.244
R12307 gnd.n4105 gnd.n2119 240.244
R12308 gnd.n4102 gnd.n2119 240.244
R12309 gnd.n4102 gnd.n2111 240.244
R12310 gnd.n4099 gnd.n2111 240.244
R12311 gnd.n4099 gnd.n2101 240.244
R12312 gnd.n4044 gnd.n2101 240.244
R12313 gnd.n4044 gnd.n2092 240.244
R12314 gnd.n4047 gnd.n2092 240.244
R12315 gnd.n4047 gnd.n2085 240.244
R12316 gnd.n4048 gnd.n2085 240.244
R12317 gnd.n4048 gnd.n2078 240.244
R12318 gnd.n4051 gnd.n2078 240.244
R12319 gnd.n4051 gnd.n2069 240.244
R12320 gnd.n4052 gnd.n2069 240.244
R12321 gnd.n4052 gnd.n2060 240.244
R12322 gnd.n4055 gnd.n2060 240.244
R12323 gnd.n4055 gnd.n2053 240.244
R12324 gnd.n4056 gnd.n2053 240.244
R12325 gnd.n4056 gnd.n2046 240.244
R12326 gnd.n4059 gnd.n2046 240.244
R12327 gnd.n4059 gnd.n2037 240.244
R12328 gnd.n4060 gnd.n2037 240.244
R12329 gnd.n4060 gnd.n2028 240.244
R12330 gnd.n4063 gnd.n2028 240.244
R12331 gnd.n4063 gnd.n2020 240.244
R12332 gnd.n2020 gnd.n2008 240.244
R12333 gnd.n4425 gnd.n2008 240.244
R12334 gnd.n4426 gnd.n4425 240.244
R12335 gnd.n4427 gnd.n4426 240.244
R12336 gnd.n4427 gnd.n1058 240.244
R12337 gnd.n4433 gnd.n1058 240.244
R12338 gnd.n4433 gnd.n1070 240.244
R12339 gnd.n4444 gnd.n1070 240.244
R12340 gnd.n4444 gnd.n1082 240.244
R12341 gnd.n4781 gnd.n1082 240.244
R12342 gnd.n4781 gnd.n1093 240.244
R12343 gnd.n4775 gnd.n1093 240.244
R12344 gnd.n4185 gnd.n4183 240.244
R12345 gnd.n4181 gnd.n3989 240.244
R12346 gnd.n4177 gnd.n4175 240.244
R12347 gnd.n4173 gnd.n3995 240.244
R12348 gnd.n4169 gnd.n4167 240.244
R12349 gnd.n4165 gnd.n4001 240.244
R12350 gnd.n4161 gnd.n4159 240.244
R12351 gnd.n4157 gnd.n4007 240.244
R12352 gnd.n4150 gnd.n4149 240.244
R12353 gnd.n4191 gnd.n2220 240.244
R12354 gnd.n4201 gnd.n2220 240.244
R12355 gnd.n4201 gnd.n2216 240.244
R12356 gnd.n4207 gnd.n2216 240.244
R12357 gnd.n4207 gnd.n2204 240.244
R12358 gnd.n4217 gnd.n2204 240.244
R12359 gnd.n4217 gnd.n2200 240.244
R12360 gnd.n4223 gnd.n2200 240.244
R12361 gnd.n4223 gnd.n2188 240.244
R12362 gnd.n4233 gnd.n2188 240.244
R12363 gnd.n4233 gnd.n2184 240.244
R12364 gnd.n4239 gnd.n2184 240.244
R12365 gnd.n4239 gnd.n2172 240.244
R12366 gnd.n4249 gnd.n2172 240.244
R12367 gnd.n4249 gnd.n2168 240.244
R12368 gnd.n4255 gnd.n2168 240.244
R12369 gnd.n4255 gnd.n2156 240.244
R12370 gnd.n4265 gnd.n2156 240.244
R12371 gnd.n4265 gnd.n2152 240.244
R12372 gnd.n4271 gnd.n2152 240.244
R12373 gnd.n4271 gnd.n2140 240.244
R12374 gnd.n4281 gnd.n2140 240.244
R12375 gnd.n4281 gnd.n2136 240.244
R12376 gnd.n4287 gnd.n2136 240.244
R12377 gnd.n4287 gnd.n2124 240.244
R12378 gnd.n4297 gnd.n2124 240.244
R12379 gnd.n4297 gnd.n2120 240.244
R12380 gnd.n4303 gnd.n2120 240.244
R12381 gnd.n4303 gnd.n2108 240.244
R12382 gnd.n4313 gnd.n2108 240.244
R12383 gnd.n4313 gnd.n2103 240.244
R12384 gnd.n4319 gnd.n2103 240.244
R12385 gnd.n4319 gnd.n2090 240.244
R12386 gnd.n4329 gnd.n2090 240.244
R12387 gnd.n4329 gnd.n2086 240.244
R12388 gnd.n4335 gnd.n2086 240.244
R12389 gnd.n4335 gnd.n2075 240.244
R12390 gnd.n4345 gnd.n2075 240.244
R12391 gnd.n4345 gnd.n2071 240.244
R12392 gnd.n4351 gnd.n2071 240.244
R12393 gnd.n4351 gnd.n2058 240.244
R12394 gnd.n4361 gnd.n2058 240.244
R12395 gnd.n4361 gnd.n2054 240.244
R12396 gnd.n4367 gnd.n2054 240.244
R12397 gnd.n4367 gnd.n2043 240.244
R12398 gnd.n4377 gnd.n2043 240.244
R12399 gnd.n4377 gnd.n2039 240.244
R12400 gnd.n4383 gnd.n2039 240.244
R12401 gnd.n4383 gnd.n2026 240.244
R12402 gnd.n4393 gnd.n2026 240.244
R12403 gnd.n4393 gnd.n2021 240.244
R12404 gnd.n4412 gnd.n2021 240.244
R12405 gnd.n4412 gnd.n2022 240.244
R12406 gnd.n2022 gnd.n2012 240.244
R12407 gnd.n4407 gnd.n2012 240.244
R12408 gnd.n4407 gnd.n4406 240.244
R12409 gnd.n4406 gnd.n1059 240.244
R12410 gnd.n1072 gnd.n1059 240.244
R12411 gnd.n6071 gnd.n1072 240.244
R12412 gnd.n6071 gnd.n1073 240.244
R12413 gnd.n6067 gnd.n1073 240.244
R12414 gnd.n6067 gnd.n1079 240.244
R12415 gnd.n6059 gnd.n1079 240.244
R12416 gnd.n6059 gnd.n1095 240.244
R12417 gnd.n1102 gnd.n1101 240.244
R12418 gnd.n1103 gnd.n1102 240.244
R12419 gnd.n4634 gnd.n1103 240.244
R12420 gnd.n4634 gnd.n1106 240.244
R12421 gnd.n1107 gnd.n1106 240.244
R12422 gnd.n1108 gnd.n1107 240.244
R12423 gnd.n4650 gnd.n1108 240.244
R12424 gnd.n4650 gnd.n1111 240.244
R12425 gnd.n1112 gnd.n1111 240.244
R12426 gnd.n1113 gnd.n1112 240.244
R12427 gnd.n4665 gnd.n1113 240.244
R12428 gnd.n4665 gnd.n1116 240.244
R12429 gnd.n1117 gnd.n1116 240.244
R12430 gnd.n1118 gnd.n1117 240.244
R12431 gnd.n1757 gnd.n1118 240.244
R12432 gnd.n1757 gnd.n1121 240.244
R12433 gnd.n1122 gnd.n1121 240.244
R12434 gnd.n1123 gnd.n1122 240.244
R12435 gnd.n1733 gnd.n1123 240.244
R12436 gnd.n1733 gnd.n1126 240.244
R12437 gnd.n1127 gnd.n1126 240.244
R12438 gnd.n1128 gnd.n1127 240.244
R12439 gnd.n5012 gnd.n1128 240.244
R12440 gnd.n5012 gnd.n1131 240.244
R12441 gnd.n1132 gnd.n1131 240.244
R12442 gnd.n1133 gnd.n1132 240.244
R12443 gnd.n1690 gnd.n1133 240.244
R12444 gnd.n1690 gnd.n1136 240.244
R12445 gnd.n1137 gnd.n1136 240.244
R12446 gnd.n1138 gnd.n1137 240.244
R12447 gnd.n5102 gnd.n1138 240.244
R12448 gnd.n5102 gnd.n1141 240.244
R12449 gnd.n1142 gnd.n1141 240.244
R12450 gnd.n1143 gnd.n1142 240.244
R12451 gnd.n1653 gnd.n1143 240.244
R12452 gnd.n1653 gnd.n1146 240.244
R12453 gnd.n1147 gnd.n1146 240.244
R12454 gnd.n1148 gnd.n1147 240.244
R12455 gnd.n5182 gnd.n1148 240.244
R12456 gnd.n5182 gnd.n1151 240.244
R12457 gnd.n1152 gnd.n1151 240.244
R12458 gnd.n1153 gnd.n1152 240.244
R12459 gnd.n5242 gnd.n1153 240.244
R12460 gnd.n5242 gnd.n1156 240.244
R12461 gnd.n1157 gnd.n1156 240.244
R12462 gnd.n1158 gnd.n1157 240.244
R12463 gnd.n5268 gnd.n1158 240.244
R12464 gnd.n5268 gnd.n1161 240.244
R12465 gnd.n1162 gnd.n1161 240.244
R12466 gnd.n1163 gnd.n1162 240.244
R12467 gnd.n1574 gnd.n1163 240.244
R12468 gnd.n1574 gnd.n1166 240.244
R12469 gnd.n1167 gnd.n1166 240.244
R12470 gnd.n1168 gnd.n1167 240.244
R12471 gnd.n1557 gnd.n1168 240.244
R12472 gnd.n1557 gnd.n1171 240.244
R12473 gnd.n1172 gnd.n1171 240.244
R12474 gnd.n1173 gnd.n1172 240.244
R12475 gnd.n5396 gnd.n1173 240.244
R12476 gnd.n5396 gnd.n1176 240.244
R12477 gnd.n1177 gnd.n1176 240.244
R12478 gnd.n1178 gnd.n1177 240.244
R12479 gnd.n1512 gnd.n1178 240.244
R12480 gnd.n1512 gnd.n1181 240.244
R12481 gnd.n1182 gnd.n1181 240.244
R12482 gnd.n1183 gnd.n1182 240.244
R12483 gnd.n1485 gnd.n1183 240.244
R12484 gnd.n1485 gnd.n1186 240.244
R12485 gnd.n1187 gnd.n1186 240.244
R12486 gnd.n1188 gnd.n1187 240.244
R12487 gnd.n5510 gnd.n1188 240.244
R12488 gnd.n5510 gnd.n1191 240.244
R12489 gnd.n1192 gnd.n1191 240.244
R12490 gnd.n1193 gnd.n1192 240.244
R12491 gnd.n5470 gnd.n1193 240.244
R12492 gnd.n5470 gnd.n1196 240.244
R12493 gnd.n1197 gnd.n1196 240.244
R12494 gnd.n1198 gnd.n1197 240.244
R12495 gnd.n1429 gnd.n1198 240.244
R12496 gnd.n1429 gnd.n1201 240.244
R12497 gnd.n1202 gnd.n1201 240.244
R12498 gnd.n1203 gnd.n1202 240.244
R12499 gnd.n1401 gnd.n1203 240.244
R12500 gnd.n1401 gnd.n1206 240.244
R12501 gnd.n1207 gnd.n1206 240.244
R12502 gnd.n1208 gnd.n1207 240.244
R12503 gnd.n1379 gnd.n1208 240.244
R12504 gnd.n1379 gnd.n1211 240.244
R12505 gnd.n1212 gnd.n1211 240.244
R12506 gnd.n1213 gnd.n1212 240.244
R12507 gnd.n1327 gnd.n1213 240.244
R12508 gnd.n1327 gnd.n1216 240.244
R12509 gnd.n1217 gnd.n1216 240.244
R12510 gnd.n1218 gnd.n1217 240.244
R12511 gnd.n1314 gnd.n1218 240.244
R12512 gnd.n1314 gnd.n1221 240.244
R12513 gnd.n1222 gnd.n1221 240.244
R12514 gnd.n1223 gnd.n1222 240.244
R12515 gnd.n5868 gnd.n1223 240.244
R12516 gnd.n5868 gnd.n1226 240.244
R12517 gnd.n5900 gnd.n1226 240.244
R12518 gnd.n4493 gnd.n4492 240.244
R12519 gnd.n4509 gnd.n4492 240.244
R12520 gnd.n4511 gnd.n4510 240.244
R12521 gnd.n4521 gnd.n4520 240.244
R12522 gnd.n4532 gnd.n4531 240.244
R12523 gnd.n4534 gnd.n4533 240.244
R12524 gnd.n4544 gnd.n4543 240.244
R12525 gnd.n4559 gnd.n4558 240.244
R12526 gnd.n4561 gnd.n4560 240.244
R12527 gnd.n4564 gnd.n4563 240.244
R12528 gnd.n4568 gnd.n4567 240.244
R12529 gnd.n4570 gnd.n4569 240.244
R12530 gnd.n4577 gnd.n4576 240.244
R12531 gnd.n4579 gnd.n4578 240.244
R12532 gnd.n4584 gnd.n4583 240.244
R12533 gnd.n4585 gnd.n4584 240.244
R12534 gnd.n4633 gnd.n4585 240.244
R12535 gnd.n4633 gnd.n4588 240.244
R12536 gnd.n4589 gnd.n4588 240.244
R12537 gnd.n4590 gnd.n4589 240.244
R12538 gnd.n4649 gnd.n4590 240.244
R12539 gnd.n4649 gnd.n4593 240.244
R12540 gnd.n4594 gnd.n4593 240.244
R12541 gnd.n4595 gnd.n4594 240.244
R12542 gnd.n4667 gnd.n4595 240.244
R12543 gnd.n4668 gnd.n4667 240.244
R12544 gnd.n4668 gnd.n1773 240.244
R12545 gnd.n1773 gnd.n1766 240.244
R12546 gnd.n4670 gnd.n1766 240.244
R12547 gnd.n4673 gnd.n4670 240.244
R12548 gnd.n4673 gnd.n1743 240.244
R12549 gnd.n4975 gnd.n1743 240.244
R12550 gnd.n4975 gnd.n1737 240.244
R12551 gnd.n4982 gnd.n1737 240.244
R12552 gnd.n4982 gnd.n1738 240.244
R12553 gnd.n1738 gnd.n1713 240.244
R12554 gnd.n5014 gnd.n1713 240.244
R12555 gnd.n5014 gnd.n1708 240.244
R12556 gnd.n5057 gnd.n1708 240.244
R12557 gnd.n5057 gnd.n1701 240.244
R12558 gnd.n5019 gnd.n1701 240.244
R12559 gnd.n5020 gnd.n5019 240.244
R12560 gnd.n5021 gnd.n5020 240.244
R12561 gnd.n5021 gnd.n1681 240.244
R12562 gnd.n1681 gnd.n1674 240.244
R12563 gnd.n5024 gnd.n1674 240.244
R12564 gnd.n5027 gnd.n5024 240.244
R12565 gnd.n5030 gnd.n5027 240.244
R12566 gnd.n5031 gnd.n5030 240.244
R12567 gnd.n5032 gnd.n5031 240.244
R12568 gnd.n5033 gnd.n5032 240.244
R12569 gnd.n5034 gnd.n5033 240.244
R12570 gnd.n5034 gnd.n1628 240.244
R12571 gnd.n5192 gnd.n1628 240.244
R12572 gnd.n5192 gnd.n1623 240.244
R12573 gnd.n5233 gnd.n1623 240.244
R12574 gnd.n5233 gnd.n1616 240.244
R12575 gnd.n5197 gnd.n1616 240.244
R12576 gnd.n5198 gnd.n5197 240.244
R12577 gnd.n5199 gnd.n5198 240.244
R12578 gnd.n5199 gnd.n1596 240.244
R12579 gnd.n1596 gnd.n1589 240.244
R12580 gnd.n5202 gnd.n1589 240.244
R12581 gnd.n5203 gnd.n5202 240.244
R12582 gnd.n5206 gnd.n5203 240.244
R12583 gnd.n5207 gnd.n5206 240.244
R12584 gnd.n5208 gnd.n5207 240.244
R12585 gnd.n5209 gnd.n5208 240.244
R12586 gnd.n5210 gnd.n5209 240.244
R12587 gnd.n5210 gnd.n1541 240.244
R12588 gnd.n5369 gnd.n1541 240.244
R12589 gnd.n5369 gnd.n1536 240.244
R12590 gnd.n5395 gnd.n1536 240.244
R12591 gnd.n5395 gnd.n1529 240.244
R12592 gnd.n5374 gnd.n1529 240.244
R12593 gnd.n5375 gnd.n5374 240.244
R12594 gnd.n5376 gnd.n5375 240.244
R12595 gnd.n5376 gnd.n1508 240.244
R12596 gnd.n1508 gnd.n1501 240.244
R12597 gnd.n5379 gnd.n1501 240.244
R12598 gnd.n5380 gnd.n5379 240.244
R12599 gnd.n5380 gnd.n1476 240.244
R12600 gnd.n5502 gnd.n1476 240.244
R12601 gnd.n5502 gnd.n1470 240.244
R12602 gnd.n5509 gnd.n1470 240.244
R12603 gnd.n5509 gnd.n1471 240.244
R12604 gnd.n1471 gnd.n1449 240.244
R12605 gnd.n5541 gnd.n1449 240.244
R12606 gnd.n5541 gnd.n1444 240.244
R12607 gnd.n5577 gnd.n1444 240.244
R12608 gnd.n5577 gnd.n1437 240.244
R12609 gnd.n5546 gnd.n1437 240.244
R12610 gnd.n5547 gnd.n5546 240.244
R12611 gnd.n5549 gnd.n5547 240.244
R12612 gnd.n5549 gnd.n1417 240.244
R12613 gnd.n1417 gnd.n1410 240.244
R12614 gnd.n5552 gnd.n1410 240.244
R12615 gnd.n5555 gnd.n5552 240.244
R12616 gnd.n5558 gnd.n5555 240.244
R12617 gnd.n5558 gnd.n1388 240.244
R12618 gnd.n1388 gnd.n1338 240.244
R12619 gnd.n5820 gnd.n1338 240.244
R12620 gnd.n5820 gnd.n1334 240.244
R12621 gnd.n5826 gnd.n1334 240.244
R12622 gnd.n5826 gnd.n1326 240.244
R12623 gnd.n5840 gnd.n1326 240.244
R12624 gnd.n5840 gnd.n1322 240.244
R12625 gnd.n5846 gnd.n1322 240.244
R12626 gnd.n5846 gnd.n1313 240.244
R12627 gnd.n5860 gnd.n1313 240.244
R12628 gnd.n5860 gnd.n1309 240.244
R12629 gnd.n5867 gnd.n1309 240.244
R12630 gnd.n5867 gnd.n1302 240.244
R12631 gnd.n5883 gnd.n1302 240.244
R12632 gnd.n5883 gnd.n1228 240.244
R12633 gnd.n1247 gnd.n460 240.244
R12634 gnd.n468 gnd.n467 240.244
R12635 gnd.n1249 gnd.n475 240.244
R12636 gnd.n1252 gnd.n476 240.244
R12637 gnd.n484 gnd.n483 240.244
R12638 gnd.n1254 gnd.n491 240.244
R12639 gnd.n1257 gnd.n492 240.244
R12640 gnd.n502 gnd.n501 240.244
R12641 gnd.n1278 gnd.n1277 240.244
R12642 gnd.n1276 gnd.n1275 240.244
R12643 gnd.n1287 gnd.n1286 240.244
R12644 gnd.n1272 gnd.n1271 240.244
R12645 gnd.n1296 gnd.n1295 240.244
R12646 gnd.n5889 gnd.n1265 240.244
R12647 gnd.n1817 gnd.n1816 240.132
R12648 gnd.n5667 gnd.n5666 240.132
R12649 gnd.n6255 gnd.n921 225.874
R12650 gnd.n6256 gnd.n6255 225.874
R12651 gnd.n6257 gnd.n6256 225.874
R12652 gnd.n6257 gnd.n915 225.874
R12653 gnd.n6265 gnd.n915 225.874
R12654 gnd.n6266 gnd.n6265 225.874
R12655 gnd.n6267 gnd.n6266 225.874
R12656 gnd.n6267 gnd.n909 225.874
R12657 gnd.n6275 gnd.n909 225.874
R12658 gnd.n6276 gnd.n6275 225.874
R12659 gnd.n6277 gnd.n6276 225.874
R12660 gnd.n6277 gnd.n903 225.874
R12661 gnd.n6285 gnd.n903 225.874
R12662 gnd.n6286 gnd.n6285 225.874
R12663 gnd.n6287 gnd.n6286 225.874
R12664 gnd.n6287 gnd.n897 225.874
R12665 gnd.n6295 gnd.n897 225.874
R12666 gnd.n6296 gnd.n6295 225.874
R12667 gnd.n6297 gnd.n6296 225.874
R12668 gnd.n6297 gnd.n891 225.874
R12669 gnd.n6305 gnd.n891 225.874
R12670 gnd.n6306 gnd.n6305 225.874
R12671 gnd.n6307 gnd.n6306 225.874
R12672 gnd.n6307 gnd.n885 225.874
R12673 gnd.n6315 gnd.n885 225.874
R12674 gnd.n6316 gnd.n6315 225.874
R12675 gnd.n6317 gnd.n6316 225.874
R12676 gnd.n6317 gnd.n879 225.874
R12677 gnd.n6325 gnd.n879 225.874
R12678 gnd.n6326 gnd.n6325 225.874
R12679 gnd.n6327 gnd.n6326 225.874
R12680 gnd.n6327 gnd.n873 225.874
R12681 gnd.n6335 gnd.n873 225.874
R12682 gnd.n6336 gnd.n6335 225.874
R12683 gnd.n6337 gnd.n6336 225.874
R12684 gnd.n6337 gnd.n867 225.874
R12685 gnd.n6345 gnd.n867 225.874
R12686 gnd.n6346 gnd.n6345 225.874
R12687 gnd.n6347 gnd.n6346 225.874
R12688 gnd.n6347 gnd.n861 225.874
R12689 gnd.n6355 gnd.n861 225.874
R12690 gnd.n6356 gnd.n6355 225.874
R12691 gnd.n6357 gnd.n6356 225.874
R12692 gnd.n6357 gnd.n855 225.874
R12693 gnd.n6365 gnd.n855 225.874
R12694 gnd.n6366 gnd.n6365 225.874
R12695 gnd.n6367 gnd.n6366 225.874
R12696 gnd.n6367 gnd.n849 225.874
R12697 gnd.n6375 gnd.n849 225.874
R12698 gnd.n6376 gnd.n6375 225.874
R12699 gnd.n6377 gnd.n6376 225.874
R12700 gnd.n6377 gnd.n843 225.874
R12701 gnd.n6385 gnd.n843 225.874
R12702 gnd.n6386 gnd.n6385 225.874
R12703 gnd.n6387 gnd.n6386 225.874
R12704 gnd.n6387 gnd.n837 225.874
R12705 gnd.n6395 gnd.n837 225.874
R12706 gnd.n6396 gnd.n6395 225.874
R12707 gnd.n6397 gnd.n6396 225.874
R12708 gnd.n6397 gnd.n831 225.874
R12709 gnd.n6405 gnd.n831 225.874
R12710 gnd.n6406 gnd.n6405 225.874
R12711 gnd.n6407 gnd.n6406 225.874
R12712 gnd.n6407 gnd.n825 225.874
R12713 gnd.n6415 gnd.n825 225.874
R12714 gnd.n6416 gnd.n6415 225.874
R12715 gnd.n6417 gnd.n6416 225.874
R12716 gnd.n6417 gnd.n819 225.874
R12717 gnd.n6425 gnd.n819 225.874
R12718 gnd.n6426 gnd.n6425 225.874
R12719 gnd.n6427 gnd.n6426 225.874
R12720 gnd.n6427 gnd.n813 225.874
R12721 gnd.n6435 gnd.n813 225.874
R12722 gnd.n6436 gnd.n6435 225.874
R12723 gnd.n6437 gnd.n6436 225.874
R12724 gnd.n6437 gnd.n807 225.874
R12725 gnd.n6445 gnd.n807 225.874
R12726 gnd.n6446 gnd.n6445 225.874
R12727 gnd.n6447 gnd.n6446 225.874
R12728 gnd.n6447 gnd.n801 225.874
R12729 gnd.n6455 gnd.n801 225.874
R12730 gnd.n6456 gnd.n6455 225.874
R12731 gnd.n6457 gnd.n6456 225.874
R12732 gnd.n6457 gnd.n795 225.874
R12733 gnd.n6465 gnd.n795 225.874
R12734 gnd.n6466 gnd.n6465 225.874
R12735 gnd.n6467 gnd.n6466 225.874
R12736 gnd.n6467 gnd.n789 225.874
R12737 gnd.n6475 gnd.n789 225.874
R12738 gnd.n6476 gnd.n6475 225.874
R12739 gnd.n6477 gnd.n6476 225.874
R12740 gnd.n6477 gnd.n783 225.874
R12741 gnd.n6485 gnd.n783 225.874
R12742 gnd.n6486 gnd.n6485 225.874
R12743 gnd.n6487 gnd.n6486 225.874
R12744 gnd.n6487 gnd.n777 225.874
R12745 gnd.n6495 gnd.n777 225.874
R12746 gnd.n6496 gnd.n6495 225.874
R12747 gnd.n6497 gnd.n6496 225.874
R12748 gnd.n6497 gnd.n771 225.874
R12749 gnd.n6505 gnd.n771 225.874
R12750 gnd.n6506 gnd.n6505 225.874
R12751 gnd.n6507 gnd.n6506 225.874
R12752 gnd.n6507 gnd.n765 225.874
R12753 gnd.n6515 gnd.n765 225.874
R12754 gnd.n6516 gnd.n6515 225.874
R12755 gnd.n6517 gnd.n6516 225.874
R12756 gnd.n6517 gnd.n759 225.874
R12757 gnd.n6525 gnd.n759 225.874
R12758 gnd.n6526 gnd.n6525 225.874
R12759 gnd.n6527 gnd.n6526 225.874
R12760 gnd.n6527 gnd.n753 225.874
R12761 gnd.n6535 gnd.n753 225.874
R12762 gnd.n6536 gnd.n6535 225.874
R12763 gnd.n6537 gnd.n6536 225.874
R12764 gnd.n6537 gnd.n747 225.874
R12765 gnd.n6545 gnd.n747 225.874
R12766 gnd.n6546 gnd.n6545 225.874
R12767 gnd.n6547 gnd.n6546 225.874
R12768 gnd.n6547 gnd.n741 225.874
R12769 gnd.n6555 gnd.n741 225.874
R12770 gnd.n6556 gnd.n6555 225.874
R12771 gnd.n6557 gnd.n6556 225.874
R12772 gnd.n6557 gnd.n735 225.874
R12773 gnd.n6566 gnd.n735 225.874
R12774 gnd.n6567 gnd.n6566 225.874
R12775 gnd.n6568 gnd.n6567 225.874
R12776 gnd.n6568 gnd.n730 225.874
R12777 gnd.n2794 gnd.t167 224.174
R12778 gnd.n2292 gnd.t144 224.174
R12779 gnd.n557 gnd.n513 199.319
R12780 gnd.n557 gnd.n514 199.319
R12781 gnd.n1905 gnd.n1899 199.319
R12782 gnd.n1904 gnd.n1899 199.319
R12783 gnd.n1818 gnd.n1815 186.49
R12784 gnd.n5668 gnd.n5665 186.49
R12785 gnd.n3569 gnd.n3568 185
R12786 gnd.n3567 gnd.n3566 185
R12787 gnd.n3546 gnd.n3545 185
R12788 gnd.n3561 gnd.n3560 185
R12789 gnd.n3559 gnd.n3558 185
R12790 gnd.n3550 gnd.n3549 185
R12791 gnd.n3553 gnd.n3552 185
R12792 gnd.n3537 gnd.n3536 185
R12793 gnd.n3535 gnd.n3534 185
R12794 gnd.n3514 gnd.n3513 185
R12795 gnd.n3529 gnd.n3528 185
R12796 gnd.n3527 gnd.n3526 185
R12797 gnd.n3518 gnd.n3517 185
R12798 gnd.n3521 gnd.n3520 185
R12799 gnd.n3505 gnd.n3504 185
R12800 gnd.n3503 gnd.n3502 185
R12801 gnd.n3482 gnd.n3481 185
R12802 gnd.n3497 gnd.n3496 185
R12803 gnd.n3495 gnd.n3494 185
R12804 gnd.n3486 gnd.n3485 185
R12805 gnd.n3489 gnd.n3488 185
R12806 gnd.n3474 gnd.n3473 185
R12807 gnd.n3472 gnd.n3471 185
R12808 gnd.n3451 gnd.n3450 185
R12809 gnd.n3466 gnd.n3465 185
R12810 gnd.n3464 gnd.n3463 185
R12811 gnd.n3455 gnd.n3454 185
R12812 gnd.n3458 gnd.n3457 185
R12813 gnd.n3442 gnd.n3441 185
R12814 gnd.n3440 gnd.n3439 185
R12815 gnd.n3419 gnd.n3418 185
R12816 gnd.n3434 gnd.n3433 185
R12817 gnd.n3432 gnd.n3431 185
R12818 gnd.n3423 gnd.n3422 185
R12819 gnd.n3426 gnd.n3425 185
R12820 gnd.n3410 gnd.n3409 185
R12821 gnd.n3408 gnd.n3407 185
R12822 gnd.n3387 gnd.n3386 185
R12823 gnd.n3402 gnd.n3401 185
R12824 gnd.n3400 gnd.n3399 185
R12825 gnd.n3391 gnd.n3390 185
R12826 gnd.n3394 gnd.n3393 185
R12827 gnd.n3378 gnd.n3377 185
R12828 gnd.n3376 gnd.n3375 185
R12829 gnd.n3355 gnd.n3354 185
R12830 gnd.n3370 gnd.n3369 185
R12831 gnd.n3368 gnd.n3367 185
R12832 gnd.n3359 gnd.n3358 185
R12833 gnd.n3362 gnd.n3361 185
R12834 gnd.n3347 gnd.n3346 185
R12835 gnd.n3345 gnd.n3344 185
R12836 gnd.n3324 gnd.n3323 185
R12837 gnd.n3339 gnd.n3338 185
R12838 gnd.n3337 gnd.n3336 185
R12839 gnd.n3328 gnd.n3327 185
R12840 gnd.n3331 gnd.n3330 185
R12841 gnd.n2795 gnd.t166 178.987
R12842 gnd.n2293 gnd.t145 178.987
R12843 gnd.n1 gnd.t281 170.774
R12844 gnd.n9 gnd.t361 170.103
R12845 gnd.n8 gnd.t227 170.103
R12846 gnd.n7 gnd.t350 170.103
R12847 gnd.n6 gnd.t316 170.103
R12848 gnd.n5 gnd.t359 170.103
R12849 gnd.n4 gnd.t220 170.103
R12850 gnd.n3 gnd.t346 170.103
R12851 gnd.n2 gnd.t201 170.103
R12852 gnd.n1 gnd.t307 170.103
R12853 gnd.n5739 gnd.n5738 163.367
R12854 gnd.n5735 gnd.n5734 163.367
R12855 gnd.n5731 gnd.n5730 163.367
R12856 gnd.n5727 gnd.n5726 163.367
R12857 gnd.n5723 gnd.n5722 163.367
R12858 gnd.n5719 gnd.n5718 163.367
R12859 gnd.n5715 gnd.n5714 163.367
R12860 gnd.n5711 gnd.n5710 163.367
R12861 gnd.n5707 gnd.n5706 163.367
R12862 gnd.n5703 gnd.n5702 163.367
R12863 gnd.n5699 gnd.n5698 163.367
R12864 gnd.n5695 gnd.n5694 163.367
R12865 gnd.n5691 gnd.n5690 163.367
R12866 gnd.n5687 gnd.n5686 163.367
R12867 gnd.n5682 gnd.n5681 163.367
R12868 gnd.n5678 gnd.n5677 163.367
R12869 gnd.n5815 gnd.n5814 163.367
R12870 gnd.n5811 gnd.n5810 163.367
R12871 gnd.n5806 gnd.n5805 163.367
R12872 gnd.n5802 gnd.n5801 163.367
R12873 gnd.n5798 gnd.n5797 163.367
R12874 gnd.n5794 gnd.n5793 163.367
R12875 gnd.n5790 gnd.n5789 163.367
R12876 gnd.n5786 gnd.n5785 163.367
R12877 gnd.n5782 gnd.n5781 163.367
R12878 gnd.n5778 gnd.n5777 163.367
R12879 gnd.n5774 gnd.n5773 163.367
R12880 gnd.n5770 gnd.n5769 163.367
R12881 gnd.n5766 gnd.n5765 163.367
R12882 gnd.n5762 gnd.n5761 163.367
R12883 gnd.n5758 gnd.n5757 163.367
R12884 gnd.n5754 gnd.n5753 163.367
R12885 gnd.n4903 gnd.n1765 163.367
R12886 gnd.n1765 gnd.n1756 163.367
R12887 gnd.n4932 gnd.n1756 163.367
R12888 gnd.n4932 gnd.n1753 163.367
R12889 gnd.n4964 gnd.n1753 163.367
R12890 gnd.n4964 gnd.n1754 163.367
R12891 gnd.n4960 gnd.n1754 163.367
R12892 gnd.n4960 gnd.n4959 163.367
R12893 gnd.n4959 gnd.n1735 163.367
R12894 gnd.n1736 gnd.n1735 163.367
R12895 gnd.n1736 gnd.n1728 163.367
R12896 gnd.n4953 gnd.n1728 163.367
R12897 gnd.n4953 gnd.n1721 163.367
R12898 gnd.n4949 gnd.n1721 163.367
R12899 gnd.n4949 gnd.n1715 163.367
R12900 gnd.n4946 gnd.n1715 163.367
R12901 gnd.n4946 gnd.n1707 163.367
R12902 gnd.n4941 gnd.n1707 163.367
R12903 gnd.n4941 gnd.n1702 163.367
R12904 gnd.n4938 gnd.n1702 163.367
R12905 gnd.n4938 gnd.n1692 163.367
R12906 gnd.n1692 gnd.n1684 163.367
R12907 gnd.n5084 gnd.n1684 163.367
R12908 gnd.n5084 gnd.n1682 163.367
R12909 gnd.n5089 gnd.n1682 163.367
R12910 gnd.n5089 gnd.n1673 163.367
R12911 gnd.n1673 gnd.n1665 163.367
R12912 gnd.n5120 gnd.n1665 163.367
R12913 gnd.n5120 gnd.n1662 163.367
R12914 gnd.n5125 gnd.n1662 163.367
R12915 gnd.n5125 gnd.n1663 163.367
R12916 gnd.n1663 gnd.n1652 163.367
R12917 gnd.n5136 gnd.n1652 163.367
R12918 gnd.n5136 gnd.n1650 163.367
R12919 gnd.n5161 gnd.n1650 163.367
R12920 gnd.n5161 gnd.n1644 163.367
R12921 gnd.n5157 gnd.n1644 163.367
R12922 gnd.n5157 gnd.n1636 163.367
R12923 gnd.n5153 gnd.n1636 163.367
R12924 gnd.n5153 gnd.n1630 163.367
R12925 gnd.n5150 gnd.n1630 163.367
R12926 gnd.n5150 gnd.n1622 163.367
R12927 gnd.n5145 gnd.n1622 163.367
R12928 gnd.n5145 gnd.n1617 163.367
R12929 gnd.n5142 gnd.n1617 163.367
R12930 gnd.n5142 gnd.n1606 163.367
R12931 gnd.n1606 gnd.n1599 163.367
R12932 gnd.n5261 gnd.n1599 163.367
R12933 gnd.n5261 gnd.n1597 163.367
R12934 gnd.n5266 gnd.n1597 163.367
R12935 gnd.n5266 gnd.n1588 163.367
R12936 gnd.n1588 gnd.n1579 163.367
R12937 gnd.n5297 gnd.n1579 163.367
R12938 gnd.n5297 gnd.n1576 163.367
R12939 gnd.n5302 gnd.n1576 163.367
R12940 gnd.n5302 gnd.n1577 163.367
R12941 gnd.n1577 gnd.n1565 163.367
R12942 gnd.n5313 gnd.n1565 163.367
R12943 gnd.n5313 gnd.n1563 163.367
R12944 gnd.n5339 gnd.n1563 163.367
R12945 gnd.n5339 gnd.n1556 163.367
R12946 gnd.n5335 gnd.n1556 163.367
R12947 gnd.n5335 gnd.n1548 163.367
R12948 gnd.n5331 gnd.n1548 163.367
R12949 gnd.n5331 gnd.n1543 163.367
R12950 gnd.n5328 gnd.n1543 163.367
R12951 gnd.n5328 gnd.n1535 163.367
R12952 gnd.n5322 gnd.n1535 163.367
R12953 gnd.n5322 gnd.n1530 163.367
R12954 gnd.n5319 gnd.n1530 163.367
R12955 gnd.n5319 gnd.n1519 163.367
R12956 gnd.n1519 gnd.n1511 163.367
R12957 gnd.n5423 gnd.n1511 163.367
R12958 gnd.n5423 gnd.n1509 163.367
R12959 gnd.n5428 gnd.n1509 163.367
R12960 gnd.n5428 gnd.n1500 163.367
R12961 gnd.n1500 gnd.n1491 163.367
R12962 gnd.n5458 gnd.n1491 163.367
R12963 gnd.n5458 gnd.n1488 163.367
R12964 gnd.n5491 gnd.n1488 163.367
R12965 gnd.n5491 gnd.n1489 163.367
R12966 gnd.n5487 gnd.n1489 163.367
R12967 gnd.n5487 gnd.n5486 163.367
R12968 gnd.n5486 gnd.n1468 163.367
R12969 gnd.n1469 gnd.n1468 163.367
R12970 gnd.n1469 gnd.n1463 163.367
R12971 gnd.n5480 gnd.n1463 163.367
R12972 gnd.n5480 gnd.n1456 163.367
R12973 gnd.n5476 gnd.n1456 163.367
R12974 gnd.n5476 gnd.n1451 163.367
R12975 gnd.n5473 gnd.n1451 163.367
R12976 gnd.n5473 gnd.n1443 163.367
R12977 gnd.n5467 gnd.n1443 163.367
R12978 gnd.n5467 gnd.n1438 163.367
R12979 gnd.n5464 gnd.n1438 163.367
R12980 gnd.n5464 gnd.n1427 163.367
R12981 gnd.n1427 gnd.n1420 163.367
R12982 gnd.n5604 gnd.n1420 163.367
R12983 gnd.n5604 gnd.n1418 163.367
R12984 gnd.n5609 gnd.n1418 163.367
R12985 gnd.n5609 gnd.n1409 163.367
R12986 gnd.n1409 gnd.n1400 163.367
R12987 gnd.n5632 gnd.n1400 163.367
R12988 gnd.n5632 gnd.n1397 163.367
R12989 gnd.n5639 gnd.n1397 163.367
R12990 gnd.n5639 gnd.n1398 163.367
R12991 gnd.n1398 gnd.n1387 163.367
R12992 gnd.n1387 gnd.n1377 163.367
R12993 gnd.n5748 gnd.n1377 163.367
R12994 gnd.n5749 gnd.n5748 163.367
R12995 gnd.n1810 gnd.n1809 163.367
R12996 gnd.n4889 gnd.n1809 163.367
R12997 gnd.n4887 gnd.n4886 163.367
R12998 gnd.n4883 gnd.n4882 163.367
R12999 gnd.n4879 gnd.n4878 163.367
R13000 gnd.n4875 gnd.n4874 163.367
R13001 gnd.n4871 gnd.n4870 163.367
R13002 gnd.n4867 gnd.n4866 163.367
R13003 gnd.n4863 gnd.n4862 163.367
R13004 gnd.n4859 gnd.n4858 163.367
R13005 gnd.n4855 gnd.n4854 163.367
R13006 gnd.n4851 gnd.n4850 163.367
R13007 gnd.n4847 gnd.n4846 163.367
R13008 gnd.n4843 gnd.n4842 163.367
R13009 gnd.n4839 gnd.n4838 163.367
R13010 gnd.n4835 gnd.n4834 163.367
R13011 gnd.n4831 gnd.n4830 163.367
R13012 gnd.n1892 gnd.n1891 163.367
R13013 gnd.n1887 gnd.n1886 163.367
R13014 gnd.n1883 gnd.n1882 163.367
R13015 gnd.n1879 gnd.n1878 163.367
R13016 gnd.n1875 gnd.n1874 163.367
R13017 gnd.n1871 gnd.n1870 163.367
R13018 gnd.n1867 gnd.n1866 163.367
R13019 gnd.n1863 gnd.n1862 163.367
R13020 gnd.n1859 gnd.n1858 163.367
R13021 gnd.n1855 gnd.n1854 163.367
R13022 gnd.n1851 gnd.n1850 163.367
R13023 gnd.n1847 gnd.n1846 163.367
R13024 gnd.n1843 gnd.n1842 163.367
R13025 gnd.n1839 gnd.n1838 163.367
R13026 gnd.n4898 gnd.n1776 163.367
R13027 gnd.n4918 gnd.n1763 163.367
R13028 gnd.n4918 gnd.n1760 163.367
R13029 gnd.n4930 gnd.n1760 163.367
R13030 gnd.n4930 gnd.n1761 163.367
R13031 gnd.n1761 gnd.n1751 163.367
R13032 gnd.n4925 gnd.n1751 163.367
R13033 gnd.n4925 gnd.n4922 163.367
R13034 gnd.n4922 gnd.n1732 163.367
R13035 gnd.n4987 gnd.n1732 163.367
R13036 gnd.n4987 gnd.n1730 163.367
R13037 gnd.n4991 gnd.n1730 163.367
R13038 gnd.n4991 gnd.n1719 163.367
R13039 gnd.n5006 gnd.n1719 163.367
R13040 gnd.n5006 gnd.n1717 163.367
R13041 gnd.n5010 gnd.n1717 163.367
R13042 gnd.n5010 gnd.n1705 163.367
R13043 gnd.n5060 gnd.n1705 163.367
R13044 gnd.n5060 gnd.n1703 163.367
R13045 gnd.n5064 gnd.n1703 163.367
R13046 gnd.n5064 gnd.n1689 163.367
R13047 gnd.n5077 gnd.n1689 163.367
R13048 gnd.n5077 gnd.n1686 163.367
R13049 gnd.n5082 gnd.n1686 163.367
R13050 gnd.n5082 gnd.n1687 163.367
R13051 gnd.n1687 gnd.n1671 163.367
R13052 gnd.n5105 gnd.n1671 163.367
R13053 gnd.n5105 gnd.n1668 163.367
R13054 gnd.n5118 gnd.n1668 163.367
R13055 gnd.n5118 gnd.n1669 163.367
R13056 gnd.n1669 gnd.n1660 163.367
R13057 gnd.n5113 gnd.n1660 163.367
R13058 gnd.n5113 gnd.n5109 163.367
R13059 gnd.n5109 gnd.n1648 163.367
R13060 gnd.n5165 gnd.n1648 163.367
R13061 gnd.n5165 gnd.n1646 163.367
R13062 gnd.n5169 gnd.n1646 163.367
R13063 gnd.n5169 gnd.n1634 163.367
R13064 gnd.n5185 gnd.n1634 163.367
R13065 gnd.n5185 gnd.n1632 163.367
R13066 gnd.n5189 gnd.n1632 163.367
R13067 gnd.n5189 gnd.n1620 163.367
R13068 gnd.n5236 gnd.n1620 163.367
R13069 gnd.n5236 gnd.n1618 163.367
R13070 gnd.n5240 gnd.n1618 163.367
R13071 gnd.n5240 gnd.n1604 163.367
R13072 gnd.n5254 gnd.n1604 163.367
R13073 gnd.n5254 gnd.n1601 163.367
R13074 gnd.n5259 gnd.n1601 163.367
R13075 gnd.n5259 gnd.n1602 163.367
R13076 gnd.n1602 gnd.n1586 163.367
R13077 gnd.n5282 gnd.n1586 163.367
R13078 gnd.n5282 gnd.n1582 163.367
R13079 gnd.n5295 gnd.n1582 163.367
R13080 gnd.n5295 gnd.n1584 163.367
R13081 gnd.n1584 gnd.n1573 163.367
R13082 gnd.n5290 gnd.n1573 163.367
R13083 gnd.n5290 gnd.n5286 163.367
R13084 gnd.n5286 gnd.n1561 163.367
R13085 gnd.n5343 gnd.n1561 163.367
R13086 gnd.n5343 gnd.n1559 163.367
R13087 gnd.n5347 gnd.n1559 163.367
R13088 gnd.n5347 gnd.n1546 163.367
R13089 gnd.n5362 gnd.n1546 163.367
R13090 gnd.n5362 gnd.n1544 163.367
R13091 gnd.n5366 gnd.n1544 163.367
R13092 gnd.n5366 gnd.n1533 163.367
R13093 gnd.n5399 gnd.n1533 163.367
R13094 gnd.n5399 gnd.n1531 163.367
R13095 gnd.n5403 gnd.n1531 163.367
R13096 gnd.n5403 gnd.n1517 163.367
R13097 gnd.n5416 gnd.n1517 163.367
R13098 gnd.n5416 gnd.n1514 163.367
R13099 gnd.n5421 gnd.n1514 163.367
R13100 gnd.n5421 gnd.n1515 163.367
R13101 gnd.n1515 gnd.n1498 163.367
R13102 gnd.n5443 gnd.n1498 163.367
R13103 gnd.n5443 gnd.n1494 163.367
R13104 gnd.n5456 gnd.n1494 163.367
R13105 gnd.n5456 gnd.n1496 163.367
R13106 gnd.n1496 gnd.n1487 163.367
R13107 gnd.n5451 gnd.n1487 163.367
R13108 gnd.n5451 gnd.n5447 163.367
R13109 gnd.n5447 gnd.n1467 163.367
R13110 gnd.n5515 gnd.n1467 163.367
R13111 gnd.n5515 gnd.n1465 163.367
R13112 gnd.n5519 gnd.n1465 163.367
R13113 gnd.n5519 gnd.n1455 163.367
R13114 gnd.n5534 gnd.n1455 163.367
R13115 gnd.n5534 gnd.n1453 163.367
R13116 gnd.n5538 gnd.n1453 163.367
R13117 gnd.n5538 gnd.n1441 163.367
R13118 gnd.n5580 gnd.n1441 163.367
R13119 gnd.n5580 gnd.n1439 163.367
R13120 gnd.n5584 gnd.n1439 163.367
R13121 gnd.n5584 gnd.n1425 163.367
R13122 gnd.n5597 gnd.n1425 163.367
R13123 gnd.n5597 gnd.n1422 163.367
R13124 gnd.n5602 gnd.n1422 163.367
R13125 gnd.n5602 gnd.n1423 163.367
R13126 gnd.n1423 gnd.n1407 163.367
R13127 gnd.n5624 gnd.n1407 163.367
R13128 gnd.n5624 gnd.n1404 163.367
R13129 gnd.n5630 gnd.n1404 163.367
R13130 gnd.n5630 gnd.n1405 163.367
R13131 gnd.n1405 gnd.n1396 163.367
R13132 gnd.n1396 gnd.n1385 163.367
R13133 gnd.n5653 gnd.n1385 163.367
R13134 gnd.n5653 gnd.n1382 163.367
R13135 gnd.n5746 gnd.n1382 163.367
R13136 gnd.n5746 gnd.n1383 163.367
R13137 gnd.n5674 gnd.n5673 156.462
R13138 gnd.n3509 gnd.n3477 153.042
R13139 gnd.n3573 gnd.n3572 152.079
R13140 gnd.n3541 gnd.n3540 152.079
R13141 gnd.n3509 gnd.n3508 152.079
R13142 gnd.n1823 gnd.n1822 152
R13143 gnd.n1824 gnd.n1813 152
R13144 gnd.n1826 gnd.n1825 152
R13145 gnd.n1828 gnd.n1811 152
R13146 gnd.n1830 gnd.n1829 152
R13147 gnd.n5672 gnd.n5656 152
R13148 gnd.n5664 gnd.n5657 152
R13149 gnd.n5663 gnd.n5662 152
R13150 gnd.n5661 gnd.n5658 152
R13151 gnd.n5659 gnd.t158 150.546
R13152 gnd.t352 gnd.n3551 147.661
R13153 gnd.t330 gnd.n3519 147.661
R13154 gnd.t231 gnd.n3487 147.661
R13155 gnd.t229 gnd.n3456 147.661
R13156 gnd.t1 gnd.n3424 147.661
R13157 gnd.t21 gnd.n3392 147.661
R13158 gnd.t322 gnd.n3360 147.661
R13159 gnd.t3 gnd.n3329 147.661
R13160 gnd.n1373 gnd.n1356 143.351
R13161 gnd.n4829 gnd.n1792 143.351
R13162 gnd.n4829 gnd.n1793 143.351
R13163 gnd.n1820 gnd.t99 130.484
R13164 gnd.n1829 gnd.t152 126.766
R13165 gnd.n1827 gnd.t96 126.766
R13166 gnd.n1813 gnd.t121 126.766
R13167 gnd.n1821 gnd.t178 126.766
R13168 gnd.n5660 gnd.t149 126.766
R13169 gnd.n5662 gnd.t93 126.766
R13170 gnd.n5671 gnd.t128 126.766
R13171 gnd.n5673 gnd.t110 126.766
R13172 gnd.n7071 gnd.n556 104.897
R13173 gnd.n4832 gnd.n4828 104.897
R13174 gnd.n3568 gnd.n3567 104.615
R13175 gnd.n3567 gnd.n3545 104.615
R13176 gnd.n3560 gnd.n3545 104.615
R13177 gnd.n3560 gnd.n3559 104.615
R13178 gnd.n3559 gnd.n3549 104.615
R13179 gnd.n3552 gnd.n3549 104.615
R13180 gnd.n3536 gnd.n3535 104.615
R13181 gnd.n3535 gnd.n3513 104.615
R13182 gnd.n3528 gnd.n3513 104.615
R13183 gnd.n3528 gnd.n3527 104.615
R13184 gnd.n3527 gnd.n3517 104.615
R13185 gnd.n3520 gnd.n3517 104.615
R13186 gnd.n3504 gnd.n3503 104.615
R13187 gnd.n3503 gnd.n3481 104.615
R13188 gnd.n3496 gnd.n3481 104.615
R13189 gnd.n3496 gnd.n3495 104.615
R13190 gnd.n3495 gnd.n3485 104.615
R13191 gnd.n3488 gnd.n3485 104.615
R13192 gnd.n3473 gnd.n3472 104.615
R13193 gnd.n3472 gnd.n3450 104.615
R13194 gnd.n3465 gnd.n3450 104.615
R13195 gnd.n3465 gnd.n3464 104.615
R13196 gnd.n3464 gnd.n3454 104.615
R13197 gnd.n3457 gnd.n3454 104.615
R13198 gnd.n3441 gnd.n3440 104.615
R13199 gnd.n3440 gnd.n3418 104.615
R13200 gnd.n3433 gnd.n3418 104.615
R13201 gnd.n3433 gnd.n3432 104.615
R13202 gnd.n3432 gnd.n3422 104.615
R13203 gnd.n3425 gnd.n3422 104.615
R13204 gnd.n3409 gnd.n3408 104.615
R13205 gnd.n3408 gnd.n3386 104.615
R13206 gnd.n3401 gnd.n3386 104.615
R13207 gnd.n3401 gnd.n3400 104.615
R13208 gnd.n3400 gnd.n3390 104.615
R13209 gnd.n3393 gnd.n3390 104.615
R13210 gnd.n3377 gnd.n3376 104.615
R13211 gnd.n3376 gnd.n3354 104.615
R13212 gnd.n3369 gnd.n3354 104.615
R13213 gnd.n3369 gnd.n3368 104.615
R13214 gnd.n3368 gnd.n3358 104.615
R13215 gnd.n3361 gnd.n3358 104.615
R13216 gnd.n3346 gnd.n3345 104.615
R13217 gnd.n3345 gnd.n3323 104.615
R13218 gnd.n3338 gnd.n3323 104.615
R13219 gnd.n3338 gnd.n3337 104.615
R13220 gnd.n3337 gnd.n3327 104.615
R13221 gnd.n3330 gnd.n3327 104.615
R13222 gnd.n2720 gnd.t196 100.632
R13223 gnd.n2266 gnd.t136 100.632
R13224 gnd.n7545 gnd.n138 99.6594
R13225 gnd.n7543 gnd.n7542 99.6594
R13226 gnd.n7538 gnd.n145 99.6594
R13227 gnd.n7536 gnd.n7535 99.6594
R13228 gnd.n7531 gnd.n152 99.6594
R13229 gnd.n7529 gnd.n7528 99.6594
R13230 gnd.n7524 gnd.n159 99.6594
R13231 gnd.n7522 gnd.n7521 99.6594
R13232 gnd.n7514 gnd.n166 99.6594
R13233 gnd.n7512 gnd.n7511 99.6594
R13234 gnd.n7507 gnd.n173 99.6594
R13235 gnd.n7505 gnd.n7504 99.6594
R13236 gnd.n7500 gnd.n180 99.6594
R13237 gnd.n7498 gnd.n7497 99.6594
R13238 gnd.n7493 gnd.n187 99.6594
R13239 gnd.n7491 gnd.n7490 99.6594
R13240 gnd.n7486 gnd.n194 99.6594
R13241 gnd.n7484 gnd.n7483 99.6594
R13242 gnd.n199 gnd.n198 99.6594
R13243 gnd.n7101 gnd.n449 99.6594
R13244 gnd.n7096 gnd.n507 99.6594
R13245 gnd.n7093 gnd.n508 99.6594
R13246 gnd.n7089 gnd.n509 99.6594
R13247 gnd.n7085 gnd.n510 99.6594
R13248 gnd.n7081 gnd.n511 99.6594
R13249 gnd.n7077 gnd.n512 99.6594
R13250 gnd.n7073 gnd.n513 99.6594
R13251 gnd.n7068 gnd.n515 99.6594
R13252 gnd.n7064 gnd.n516 99.6594
R13253 gnd.n7060 gnd.n517 99.6594
R13254 gnd.n7056 gnd.n518 99.6594
R13255 gnd.n7052 gnd.n519 99.6594
R13256 gnd.n7048 gnd.n520 99.6594
R13257 gnd.n7044 gnd.n521 99.6594
R13258 gnd.n7040 gnd.n522 99.6594
R13259 gnd.n7036 gnd.n523 99.6594
R13260 gnd.n580 gnd.n524 99.6594
R13261 gnd.n7400 gnd.n7399 99.6594
R13262 gnd.n7405 gnd.n7404 99.6594
R13263 gnd.n7408 gnd.n7407 99.6594
R13264 gnd.n7413 gnd.n7412 99.6594
R13265 gnd.n7416 gnd.n7415 99.6594
R13266 gnd.n7421 gnd.n7420 99.6594
R13267 gnd.n7424 gnd.n7423 99.6594
R13268 gnd.n7429 gnd.n7427 99.6594
R13269 gnd.n7555 gnd.n125 99.6594
R13270 gnd.n525 gnd.n454 99.6594
R13271 gnd.n527 gnd.n526 99.6594
R13272 gnd.n529 gnd.n464 99.6594
R13273 gnd.n530 gnd.n471 99.6594
R13274 gnd.n532 gnd.n531 99.6594
R13275 gnd.n534 gnd.n480 99.6594
R13276 gnd.n535 gnd.n487 99.6594
R13277 gnd.n537 gnd.n536 99.6594
R13278 gnd.n538 gnd.n496 99.6594
R13279 gnd.n6248 gnd.n6247 99.6594
R13280 gnd.n970 gnd.n928 99.6594
R13281 gnd.n6240 gnd.n929 99.6594
R13282 gnd.n6236 gnd.n930 99.6594
R13283 gnd.n6232 gnd.n931 99.6594
R13284 gnd.n6228 gnd.n932 99.6594
R13285 gnd.n6224 gnd.n933 99.6594
R13286 gnd.n6220 gnd.n934 99.6594
R13287 gnd.n6216 gnd.n935 99.6594
R13288 gnd.n6212 gnd.n936 99.6594
R13289 gnd.n6208 gnd.n937 99.6594
R13290 gnd.n6204 gnd.n938 99.6594
R13291 gnd.n6200 gnd.n939 99.6594
R13292 gnd.n6196 gnd.n940 99.6594
R13293 gnd.n6192 gnd.n941 99.6594
R13294 gnd.n6188 gnd.n942 99.6594
R13295 gnd.n6184 gnd.n943 99.6594
R13296 gnd.n6180 gnd.n944 99.6594
R13297 gnd.n6176 gnd.n945 99.6594
R13298 gnd.n6172 gnd.n946 99.6594
R13299 gnd.n6168 gnd.n947 99.6594
R13300 gnd.n6164 gnd.n948 99.6594
R13301 gnd.n6160 gnd.n949 99.6594
R13302 gnd.n6156 gnd.n950 99.6594
R13303 gnd.n6152 gnd.n951 99.6594
R13304 gnd.n6148 gnd.n952 99.6594
R13305 gnd.n6144 gnd.n953 99.6594
R13306 gnd.n6140 gnd.n954 99.6594
R13307 gnd.n6136 gnd.n955 99.6594
R13308 gnd.n6132 gnd.n956 99.6594
R13309 gnd.n6128 gnd.n957 99.6594
R13310 gnd.n6124 gnd.n958 99.6594
R13311 gnd.n6120 gnd.n959 99.6594
R13312 gnd.n6116 gnd.n960 99.6594
R13313 gnd.n6112 gnd.n961 99.6594
R13314 gnd.n6108 gnd.n962 99.6594
R13315 gnd.n6104 gnd.n963 99.6594
R13316 gnd.n6100 gnd.n964 99.6594
R13317 gnd.n6096 gnd.n965 99.6594
R13318 gnd.n6092 gnd.n966 99.6594
R13319 gnd.n6088 gnd.n967 99.6594
R13320 gnd.n6084 gnd.n968 99.6594
R13321 gnd.n1955 gnd.n1912 99.6594
R13322 gnd.n1951 gnd.n1911 99.6594
R13323 gnd.n1947 gnd.n1910 99.6594
R13324 gnd.n1943 gnd.n1909 99.6594
R13325 gnd.n1939 gnd.n1908 99.6594
R13326 gnd.n1935 gnd.n1907 99.6594
R13327 gnd.n1931 gnd.n1906 99.6594
R13328 gnd.n1904 gnd.n1903 99.6594
R13329 gnd.n4822 gnd.n4821 99.6594
R13330 gnd.n4819 gnd.n4818 99.6594
R13331 gnd.n4814 gnd.n1968 99.6594
R13332 gnd.n4812 gnd.n4811 99.6594
R13333 gnd.n4807 gnd.n1975 99.6594
R13334 gnd.n4805 gnd.n4804 99.6594
R13335 gnd.n4800 gnd.n1982 99.6594
R13336 gnd.n4798 gnd.n4797 99.6594
R13337 gnd.n4793 gnd.n1991 99.6594
R13338 gnd.n4791 gnd.n4790 99.6594
R13339 gnd.n3749 gnd.n2226 99.6594
R13340 gnd.n3757 gnd.n3756 99.6594
R13341 gnd.n3760 gnd.n3759 99.6594
R13342 gnd.n3767 gnd.n3766 99.6594
R13343 gnd.n3770 gnd.n3769 99.6594
R13344 gnd.n3777 gnd.n3776 99.6594
R13345 gnd.n3780 gnd.n3779 99.6594
R13346 gnd.n3787 gnd.n3786 99.6594
R13347 gnd.n3790 gnd.n3789 99.6594
R13348 gnd.n3797 gnd.n3796 99.6594
R13349 gnd.n3800 gnd.n3799 99.6594
R13350 gnd.n3807 gnd.n3806 99.6594
R13351 gnd.n3810 gnd.n3809 99.6594
R13352 gnd.n3817 gnd.n3816 99.6594
R13353 gnd.n3820 gnd.n3819 99.6594
R13354 gnd.n3827 gnd.n3826 99.6594
R13355 gnd.n3830 gnd.n3829 99.6594
R13356 gnd.n3838 gnd.n3837 99.6594
R13357 gnd.n3841 gnd.n3840 99.6594
R13358 gnd.n3691 gnd.n2249 99.6594
R13359 gnd.n3689 gnd.n2248 99.6594
R13360 gnd.n3685 gnd.n2247 99.6594
R13361 gnd.n3681 gnd.n2246 99.6594
R13362 gnd.n3677 gnd.n2245 99.6594
R13363 gnd.n3673 gnd.n2244 99.6594
R13364 gnd.n3669 gnd.n2243 99.6594
R13365 gnd.n3601 gnd.n2242 99.6594
R13366 gnd.n2932 gnd.n2663 99.6594
R13367 gnd.n2689 gnd.n2670 99.6594
R13368 gnd.n2691 gnd.n2671 99.6594
R13369 gnd.n2699 gnd.n2672 99.6594
R13370 gnd.n2701 gnd.n2673 99.6594
R13371 gnd.n2709 gnd.n2674 99.6594
R13372 gnd.n2711 gnd.n2675 99.6594
R13373 gnd.n2719 gnd.n2676 99.6594
R13374 gnd.n3659 gnd.n2229 99.6594
R13375 gnd.n3655 gnd.n2230 99.6594
R13376 gnd.n3651 gnd.n2231 99.6594
R13377 gnd.n3647 gnd.n2232 99.6594
R13378 gnd.n3643 gnd.n2233 99.6594
R13379 gnd.n3639 gnd.n2234 99.6594
R13380 gnd.n3635 gnd.n2235 99.6594
R13381 gnd.n3631 gnd.n2236 99.6594
R13382 gnd.n3627 gnd.n2237 99.6594
R13383 gnd.n3623 gnd.n2238 99.6594
R13384 gnd.n3619 gnd.n2239 99.6594
R13385 gnd.n3615 gnd.n2240 99.6594
R13386 gnd.n3611 gnd.n2241 99.6594
R13387 gnd.n2847 gnd.n2846 99.6594
R13388 gnd.n2841 gnd.n2758 99.6594
R13389 gnd.n2838 gnd.n2759 99.6594
R13390 gnd.n2834 gnd.n2760 99.6594
R13391 gnd.n2830 gnd.n2761 99.6594
R13392 gnd.n2826 gnd.n2762 99.6594
R13393 gnd.n2822 gnd.n2763 99.6594
R13394 gnd.n2818 gnd.n2764 99.6594
R13395 gnd.n2814 gnd.n2765 99.6594
R13396 gnd.n2810 gnd.n2766 99.6594
R13397 gnd.n2806 gnd.n2767 99.6594
R13398 gnd.n2802 gnd.n2768 99.6594
R13399 gnd.n2849 gnd.n2757 99.6594
R13400 gnd.n4503 gnd.n4502 99.6594
R13401 gnd.n4506 gnd.n4505 99.6594
R13402 gnd.n4516 gnd.n4515 99.6594
R13403 gnd.n4525 gnd.n4524 99.6594
R13404 gnd.n4528 gnd.n4527 99.6594
R13405 gnd.n4539 gnd.n4538 99.6594
R13406 gnd.n4548 gnd.n4547 99.6594
R13407 gnd.n4551 gnd.n4550 99.6594
R13408 gnd.n4554 gnd.n4449 99.6594
R13409 gnd.n4184 gnd.n3986 99.6594
R13410 gnd.n4183 gnd.n4182 99.6594
R13411 gnd.n4176 gnd.n3989 99.6594
R13412 gnd.n4175 gnd.n4174 99.6594
R13413 gnd.n4168 gnd.n3995 99.6594
R13414 gnd.n4167 gnd.n4166 99.6594
R13415 gnd.n4160 gnd.n4001 99.6594
R13416 gnd.n4159 gnd.n4158 99.6594
R13417 gnd.n4148 gnd.n4007 99.6594
R13418 gnd.n4185 gnd.n4184 99.6594
R13419 gnd.n4182 gnd.n4181 99.6594
R13420 gnd.n4177 gnd.n4176 99.6594
R13421 gnd.n4174 gnd.n4173 99.6594
R13422 gnd.n4169 gnd.n4168 99.6594
R13423 gnd.n4166 gnd.n4165 99.6594
R13424 gnd.n4161 gnd.n4160 99.6594
R13425 gnd.n4158 gnd.n4157 99.6594
R13426 gnd.n4149 gnd.n4148 99.6594
R13427 gnd.n2847 gnd.n2770 99.6594
R13428 gnd.n2839 gnd.n2758 99.6594
R13429 gnd.n2835 gnd.n2759 99.6594
R13430 gnd.n2831 gnd.n2760 99.6594
R13431 gnd.n2827 gnd.n2761 99.6594
R13432 gnd.n2823 gnd.n2762 99.6594
R13433 gnd.n2819 gnd.n2763 99.6594
R13434 gnd.n2815 gnd.n2764 99.6594
R13435 gnd.n2811 gnd.n2765 99.6594
R13436 gnd.n2807 gnd.n2766 99.6594
R13437 gnd.n2803 gnd.n2767 99.6594
R13438 gnd.n2799 gnd.n2768 99.6594
R13439 gnd.n2850 gnd.n2849 99.6594
R13440 gnd.n3614 gnd.n2241 99.6594
R13441 gnd.n3618 gnd.n2240 99.6594
R13442 gnd.n3622 gnd.n2239 99.6594
R13443 gnd.n3626 gnd.n2238 99.6594
R13444 gnd.n3630 gnd.n2237 99.6594
R13445 gnd.n3634 gnd.n2236 99.6594
R13446 gnd.n3638 gnd.n2235 99.6594
R13447 gnd.n3642 gnd.n2234 99.6594
R13448 gnd.n3646 gnd.n2233 99.6594
R13449 gnd.n3650 gnd.n2232 99.6594
R13450 gnd.n3654 gnd.n2231 99.6594
R13451 gnd.n3658 gnd.n2230 99.6594
R13452 gnd.n2270 gnd.n2229 99.6594
R13453 gnd.n2933 gnd.n2932 99.6594
R13454 gnd.n2692 gnd.n2670 99.6594
R13455 gnd.n2698 gnd.n2671 99.6594
R13456 gnd.n2702 gnd.n2672 99.6594
R13457 gnd.n2708 gnd.n2673 99.6594
R13458 gnd.n2712 gnd.n2674 99.6594
R13459 gnd.n2718 gnd.n2675 99.6594
R13460 gnd.n2676 gnd.n2660 99.6594
R13461 gnd.n3668 gnd.n2242 99.6594
R13462 gnd.n3672 gnd.n2243 99.6594
R13463 gnd.n3676 gnd.n2244 99.6594
R13464 gnd.n3680 gnd.n2245 99.6594
R13465 gnd.n3684 gnd.n2246 99.6594
R13466 gnd.n3688 gnd.n2247 99.6594
R13467 gnd.n3692 gnd.n2248 99.6594
R13468 gnd.n2251 gnd.n2249 99.6594
R13469 gnd.n3750 gnd.n3749 99.6594
R13470 gnd.n3758 gnd.n3757 99.6594
R13471 gnd.n3759 gnd.n3742 99.6594
R13472 gnd.n3768 gnd.n3767 99.6594
R13473 gnd.n3769 gnd.n3738 99.6594
R13474 gnd.n3778 gnd.n3777 99.6594
R13475 gnd.n3779 gnd.n3734 99.6594
R13476 gnd.n3788 gnd.n3787 99.6594
R13477 gnd.n3789 gnd.n3727 99.6594
R13478 gnd.n3798 gnd.n3797 99.6594
R13479 gnd.n3799 gnd.n3723 99.6594
R13480 gnd.n3808 gnd.n3807 99.6594
R13481 gnd.n3809 gnd.n3719 99.6594
R13482 gnd.n3818 gnd.n3817 99.6594
R13483 gnd.n3819 gnd.n3715 99.6594
R13484 gnd.n3828 gnd.n3827 99.6594
R13485 gnd.n3829 gnd.n3711 99.6594
R13486 gnd.n3839 gnd.n3838 99.6594
R13487 gnd.n3842 gnd.n3841 99.6594
R13488 gnd.n6247 gnd.n926 99.6594
R13489 gnd.n6241 gnd.n928 99.6594
R13490 gnd.n6237 gnd.n929 99.6594
R13491 gnd.n6233 gnd.n930 99.6594
R13492 gnd.n6229 gnd.n931 99.6594
R13493 gnd.n6225 gnd.n932 99.6594
R13494 gnd.n6221 gnd.n933 99.6594
R13495 gnd.n6217 gnd.n934 99.6594
R13496 gnd.n6213 gnd.n935 99.6594
R13497 gnd.n6209 gnd.n936 99.6594
R13498 gnd.n6205 gnd.n937 99.6594
R13499 gnd.n6201 gnd.n938 99.6594
R13500 gnd.n6197 gnd.n939 99.6594
R13501 gnd.n6193 gnd.n940 99.6594
R13502 gnd.n6189 gnd.n941 99.6594
R13503 gnd.n6185 gnd.n942 99.6594
R13504 gnd.n6181 gnd.n943 99.6594
R13505 gnd.n6177 gnd.n944 99.6594
R13506 gnd.n6173 gnd.n945 99.6594
R13507 gnd.n6169 gnd.n946 99.6594
R13508 gnd.n6165 gnd.n947 99.6594
R13509 gnd.n6161 gnd.n948 99.6594
R13510 gnd.n6157 gnd.n949 99.6594
R13511 gnd.n6153 gnd.n950 99.6594
R13512 gnd.n6149 gnd.n951 99.6594
R13513 gnd.n6145 gnd.n952 99.6594
R13514 gnd.n6141 gnd.n953 99.6594
R13515 gnd.n6137 gnd.n954 99.6594
R13516 gnd.n6133 gnd.n955 99.6594
R13517 gnd.n6129 gnd.n956 99.6594
R13518 gnd.n6125 gnd.n957 99.6594
R13519 gnd.n6121 gnd.n958 99.6594
R13520 gnd.n6117 gnd.n959 99.6594
R13521 gnd.n6113 gnd.n960 99.6594
R13522 gnd.n6109 gnd.n961 99.6594
R13523 gnd.n6105 gnd.n962 99.6594
R13524 gnd.n6101 gnd.n963 99.6594
R13525 gnd.n6097 gnd.n964 99.6594
R13526 gnd.n6093 gnd.n965 99.6594
R13527 gnd.n6089 gnd.n966 99.6594
R13528 gnd.n6085 gnd.n967 99.6594
R13529 gnd.n6081 gnd.n968 99.6594
R13530 gnd.n4555 gnd.n4554 99.6594
R13531 gnd.n4550 gnd.n4549 99.6594
R13532 gnd.n4547 gnd.n4540 99.6594
R13533 gnd.n4538 gnd.n4537 99.6594
R13534 gnd.n4527 gnd.n4526 99.6594
R13535 gnd.n4524 gnd.n4517 99.6594
R13536 gnd.n4515 gnd.n4514 99.6594
R13537 gnd.n4505 gnd.n4504 99.6594
R13538 gnd.n4502 gnd.n4501 99.6594
R13539 gnd.n525 gnd.n456 99.6594
R13540 gnd.n527 gnd.n463 99.6594
R13541 gnd.n529 gnd.n528 99.6594
R13542 gnd.n530 gnd.n472 99.6594
R13543 gnd.n532 gnd.n479 99.6594
R13544 gnd.n534 gnd.n533 99.6594
R13545 gnd.n535 gnd.n488 99.6594
R13546 gnd.n537 gnd.n495 99.6594
R13547 gnd.n538 gnd.n505 99.6594
R13548 gnd.n7428 gnd.n125 99.6594
R13549 gnd.n7427 gnd.n7426 99.6594
R13550 gnd.n7423 gnd.n7422 99.6594
R13551 gnd.n7420 gnd.n7419 99.6594
R13552 gnd.n7415 gnd.n7414 99.6594
R13553 gnd.n7412 gnd.n7411 99.6594
R13554 gnd.n7407 gnd.n7406 99.6594
R13555 gnd.n7404 gnd.n7403 99.6594
R13556 gnd.n7399 gnd.n7398 99.6594
R13557 gnd.n4792 gnd.n4791 99.6594
R13558 gnd.n1991 gnd.n1983 99.6594
R13559 gnd.n4799 gnd.n4798 99.6594
R13560 gnd.n1982 gnd.n1976 99.6594
R13561 gnd.n4806 gnd.n4805 99.6594
R13562 gnd.n1975 gnd.n1969 99.6594
R13563 gnd.n4813 gnd.n4812 99.6594
R13564 gnd.n1968 gnd.n1962 99.6594
R13565 gnd.n4820 gnd.n4819 99.6594
R13566 gnd.n4823 gnd.n4822 99.6594
R13567 gnd.n1930 gnd.n1905 99.6594
R13568 gnd.n1934 gnd.n1906 99.6594
R13569 gnd.n1938 gnd.n1907 99.6594
R13570 gnd.n1942 gnd.n1908 99.6594
R13571 gnd.n1946 gnd.n1909 99.6594
R13572 gnd.n1950 gnd.n1910 99.6594
R13573 gnd.n1954 gnd.n1911 99.6594
R13574 gnd.n1913 gnd.n1912 99.6594
R13575 gnd.n7101 gnd.n7100 99.6594
R13576 gnd.n7094 gnd.n507 99.6594
R13577 gnd.n7090 gnd.n508 99.6594
R13578 gnd.n7086 gnd.n509 99.6594
R13579 gnd.n7082 gnd.n510 99.6594
R13580 gnd.n7078 gnd.n511 99.6594
R13581 gnd.n7074 gnd.n512 99.6594
R13582 gnd.n7069 gnd.n514 99.6594
R13583 gnd.n7065 gnd.n515 99.6594
R13584 gnd.n7061 gnd.n516 99.6594
R13585 gnd.n7057 gnd.n517 99.6594
R13586 gnd.n7053 gnd.n518 99.6594
R13587 gnd.n7049 gnd.n519 99.6594
R13588 gnd.n7045 gnd.n520 99.6594
R13589 gnd.n7041 gnd.n521 99.6594
R13590 gnd.n7037 gnd.n522 99.6594
R13591 gnd.n579 gnd.n523 99.6594
R13592 gnd.n7029 gnd.n524 99.6594
R13593 gnd.n198 gnd.n195 99.6594
R13594 gnd.n7485 gnd.n7484 99.6594
R13595 gnd.n194 gnd.n188 99.6594
R13596 gnd.n7492 gnd.n7491 99.6594
R13597 gnd.n187 gnd.n181 99.6594
R13598 gnd.n7499 gnd.n7498 99.6594
R13599 gnd.n180 gnd.n174 99.6594
R13600 gnd.n7506 gnd.n7505 99.6594
R13601 gnd.n173 gnd.n167 99.6594
R13602 gnd.n7513 gnd.n7512 99.6594
R13603 gnd.n166 gnd.n160 99.6594
R13604 gnd.n7523 gnd.n7522 99.6594
R13605 gnd.n159 gnd.n153 99.6594
R13606 gnd.n7530 gnd.n7529 99.6594
R13607 gnd.n152 gnd.n146 99.6594
R13608 gnd.n7537 gnd.n7536 99.6594
R13609 gnd.n145 gnd.n139 99.6594
R13610 gnd.n7544 gnd.n7543 99.6594
R13611 gnd.n138 gnd.n135 99.6594
R13612 gnd.n4764 gnd.n4763 99.6594
R13613 gnd.n4509 gnd.n4478 99.6594
R13614 gnd.n4511 gnd.n4479 99.6594
R13615 gnd.n4521 gnd.n4480 99.6594
R13616 gnd.n4532 gnd.n4481 99.6594
R13617 gnd.n4534 gnd.n4482 99.6594
R13618 gnd.n4544 gnd.n4483 99.6594
R13619 gnd.n4559 gnd.n4484 99.6594
R13620 gnd.n4561 gnd.n4485 99.6594
R13621 gnd.n4564 gnd.n4486 99.6594
R13622 gnd.n4568 gnd.n4487 99.6594
R13623 gnd.n4570 gnd.n4488 99.6594
R13624 gnd.n4577 gnd.n4489 99.6594
R13625 gnd.n4579 gnd.n4490 99.6594
R13626 gnd.n4764 gnd.n4493 99.6594
R13627 gnd.n4510 gnd.n4478 99.6594
R13628 gnd.n4520 gnd.n4479 99.6594
R13629 gnd.n4531 gnd.n4480 99.6594
R13630 gnd.n4533 gnd.n4481 99.6594
R13631 gnd.n4543 gnd.n4482 99.6594
R13632 gnd.n4558 gnd.n4483 99.6594
R13633 gnd.n4560 gnd.n4484 99.6594
R13634 gnd.n4563 gnd.n4485 99.6594
R13635 gnd.n4567 gnd.n4486 99.6594
R13636 gnd.n4569 gnd.n4487 99.6594
R13637 gnd.n4576 gnd.n4488 99.6594
R13638 gnd.n4578 gnd.n4489 99.6594
R13639 gnd.n4582 gnd.n4490 99.6594
R13640 gnd.n1246 gnd.n460 99.6594
R13641 gnd.n1248 gnd.n467 99.6594
R13642 gnd.n1250 gnd.n1249 99.6594
R13643 gnd.n1251 gnd.n476 99.6594
R13644 gnd.n1253 gnd.n483 99.6594
R13645 gnd.n1255 gnd.n1254 99.6594
R13646 gnd.n1256 gnd.n492 99.6594
R13647 gnd.n1258 gnd.n501 99.6594
R13648 gnd.n1277 gnd.n1259 99.6594
R13649 gnd.n1275 gnd.n1260 99.6594
R13650 gnd.n1286 gnd.n1261 99.6594
R13651 gnd.n1271 gnd.n1262 99.6594
R13652 gnd.n1295 gnd.n1263 99.6594
R13653 gnd.n1265 gnd.n1264 99.6594
R13654 gnd.n1296 gnd.n1264 99.6594
R13655 gnd.n1272 gnd.n1263 99.6594
R13656 gnd.n1287 gnd.n1262 99.6594
R13657 gnd.n1276 gnd.n1261 99.6594
R13658 gnd.n1278 gnd.n1260 99.6594
R13659 gnd.n1259 gnd.n502 99.6594
R13660 gnd.n1258 gnd.n1257 99.6594
R13661 gnd.n1256 gnd.n491 99.6594
R13662 gnd.n1255 gnd.n484 99.6594
R13663 gnd.n1253 gnd.n1252 99.6594
R13664 gnd.n1251 gnd.n475 99.6594
R13665 gnd.n1250 gnd.n468 99.6594
R13666 gnd.n1248 gnd.n1247 99.6594
R13667 gnd.n1246 gnd.n459 99.6594
R13668 gnd.n4573 gnd.t141 98.63
R13669 gnd.n559 gnd.t133 98.63
R13670 gnd.n581 gnd.t116 98.63
R13671 gnd.n201 gnd.t176 98.63
R13672 gnd.n7516 gnd.t91 98.63
R13673 gnd.n122 gnd.t147 98.63
R13674 gnd.n497 gnd.t163 98.63
R13675 gnd.n4552 gnd.t182 98.63
R13676 gnd.n1988 gnd.t185 98.63
R13677 gnd.n1897 gnd.t108 98.63
R13678 gnd.n3731 gnd.t192 98.63
R13679 gnd.n3707 gnd.t171 98.63
R13680 gnd.n4010 gnd.t189 98.63
R13681 gnd.n1268 gnd.t104 98.63
R13682 gnd.n1835 gnd.t174 96.6984
R13683 gnd.n1374 gnd.t119 96.6984
R13684 gnd.n1832 gnd.t127 96.6906
R13685 gnd.n5675 gnd.t156 96.6906
R13686 gnd.n1820 gnd.n1819 81.8399
R13687 gnd.n2721 gnd.t195 74.8376
R13688 gnd.n2267 gnd.t137 74.8376
R13689 gnd.n1836 gnd.t173 72.8438
R13690 gnd.n1375 gnd.t120 72.8438
R13691 gnd.n1821 gnd.n1814 72.8411
R13692 gnd.n1827 gnd.n1812 72.8411
R13693 gnd.n5671 gnd.n5670 72.8411
R13694 gnd.n4574 gnd.t140 72.836
R13695 gnd.n1833 gnd.t126 72.836
R13696 gnd.n5676 gnd.t157 72.836
R13697 gnd.n560 gnd.t132 72.836
R13698 gnd.n582 gnd.t115 72.836
R13699 gnd.n202 gnd.t177 72.836
R13700 gnd.n7517 gnd.t92 72.836
R13701 gnd.n123 gnd.t148 72.836
R13702 gnd.n498 gnd.t162 72.836
R13703 gnd.n4553 gnd.t183 72.836
R13704 gnd.n1989 gnd.t186 72.836
R13705 gnd.n1898 gnd.t109 72.836
R13706 gnd.n3732 gnd.t191 72.836
R13707 gnd.n3708 gnd.t170 72.836
R13708 gnd.n4011 gnd.t188 72.836
R13709 gnd.n1269 gnd.t105 72.836
R13710 gnd.n5739 gnd.n1340 71.676
R13711 gnd.n5735 gnd.n1341 71.676
R13712 gnd.n5731 gnd.n1342 71.676
R13713 gnd.n5727 gnd.n1343 71.676
R13714 gnd.n5723 gnd.n1344 71.676
R13715 gnd.n5719 gnd.n1345 71.676
R13716 gnd.n5715 gnd.n1346 71.676
R13717 gnd.n5711 gnd.n1347 71.676
R13718 gnd.n5707 gnd.n1348 71.676
R13719 gnd.n5703 gnd.n1349 71.676
R13720 gnd.n5699 gnd.n1350 71.676
R13721 gnd.n5695 gnd.n1351 71.676
R13722 gnd.n5691 gnd.n1352 71.676
R13723 gnd.n5687 gnd.n1353 71.676
R13724 gnd.n5682 gnd.n1354 71.676
R13725 gnd.n5678 gnd.n1355 71.676
R13726 gnd.n5815 gnd.n1373 71.676
R13727 gnd.n5811 gnd.n1372 71.676
R13728 gnd.n5806 gnd.n1371 71.676
R13729 gnd.n5802 gnd.n1370 71.676
R13730 gnd.n5798 gnd.n1369 71.676
R13731 gnd.n5794 gnd.n1368 71.676
R13732 gnd.n5790 gnd.n1367 71.676
R13733 gnd.n5786 gnd.n1366 71.676
R13734 gnd.n5782 gnd.n1365 71.676
R13735 gnd.n5778 gnd.n1364 71.676
R13736 gnd.n5774 gnd.n1363 71.676
R13737 gnd.n5770 gnd.n1362 71.676
R13738 gnd.n5766 gnd.n1361 71.676
R13739 gnd.n5762 gnd.n1360 71.676
R13740 gnd.n5758 gnd.n1359 71.676
R13741 gnd.n5754 gnd.n1358 71.676
R13742 gnd.n5750 gnd.n1357 71.676
R13743 gnd.n4895 gnd.n4894 71.676
R13744 gnd.n4889 gnd.n1778 71.676
R13745 gnd.n4886 gnd.n1779 71.676
R13746 gnd.n4882 gnd.n1780 71.676
R13747 gnd.n4878 gnd.n1781 71.676
R13748 gnd.n4874 gnd.n1782 71.676
R13749 gnd.n4870 gnd.n1783 71.676
R13750 gnd.n4866 gnd.n1784 71.676
R13751 gnd.n4862 gnd.n1785 71.676
R13752 gnd.n4858 gnd.n1786 71.676
R13753 gnd.n4854 gnd.n1787 71.676
R13754 gnd.n4850 gnd.n1788 71.676
R13755 gnd.n4846 gnd.n1789 71.676
R13756 gnd.n4842 gnd.n1790 71.676
R13757 gnd.n4838 gnd.n1791 71.676
R13758 gnd.n4834 gnd.n1792 71.676
R13759 gnd.n4830 gnd.n1794 71.676
R13760 gnd.n1891 gnd.n1795 71.676
R13761 gnd.n1886 gnd.n1796 71.676
R13762 gnd.n1882 gnd.n1797 71.676
R13763 gnd.n1878 gnd.n1798 71.676
R13764 gnd.n1874 gnd.n1799 71.676
R13765 gnd.n1870 gnd.n1800 71.676
R13766 gnd.n1866 gnd.n1801 71.676
R13767 gnd.n1862 gnd.n1802 71.676
R13768 gnd.n1858 gnd.n1803 71.676
R13769 gnd.n1854 gnd.n1804 71.676
R13770 gnd.n1850 gnd.n1805 71.676
R13771 gnd.n1846 gnd.n1806 71.676
R13772 gnd.n1842 gnd.n1807 71.676
R13773 gnd.n1838 gnd.n1808 71.676
R13774 gnd.n4898 gnd.n4897 71.676
R13775 gnd.n4895 gnd.n1810 71.676
R13776 gnd.n4887 gnd.n1778 71.676
R13777 gnd.n4883 gnd.n1779 71.676
R13778 gnd.n4879 gnd.n1780 71.676
R13779 gnd.n4875 gnd.n1781 71.676
R13780 gnd.n4871 gnd.n1782 71.676
R13781 gnd.n4867 gnd.n1783 71.676
R13782 gnd.n4863 gnd.n1784 71.676
R13783 gnd.n4859 gnd.n1785 71.676
R13784 gnd.n4855 gnd.n1786 71.676
R13785 gnd.n4851 gnd.n1787 71.676
R13786 gnd.n4847 gnd.n1788 71.676
R13787 gnd.n4843 gnd.n1789 71.676
R13788 gnd.n4839 gnd.n1790 71.676
R13789 gnd.n4835 gnd.n1791 71.676
R13790 gnd.n4831 gnd.n1793 71.676
R13791 gnd.n1892 gnd.n1794 71.676
R13792 gnd.n1887 gnd.n1795 71.676
R13793 gnd.n1883 gnd.n1796 71.676
R13794 gnd.n1879 gnd.n1797 71.676
R13795 gnd.n1875 gnd.n1798 71.676
R13796 gnd.n1871 gnd.n1799 71.676
R13797 gnd.n1867 gnd.n1800 71.676
R13798 gnd.n1863 gnd.n1801 71.676
R13799 gnd.n1859 gnd.n1802 71.676
R13800 gnd.n1855 gnd.n1803 71.676
R13801 gnd.n1851 gnd.n1804 71.676
R13802 gnd.n1847 gnd.n1805 71.676
R13803 gnd.n1843 gnd.n1806 71.676
R13804 gnd.n1839 gnd.n1807 71.676
R13805 gnd.n1808 gnd.n1776 71.676
R13806 gnd.n4897 gnd.n1774 71.676
R13807 gnd.n5753 gnd.n1357 71.676
R13808 gnd.n5757 gnd.n1358 71.676
R13809 gnd.n5761 gnd.n1359 71.676
R13810 gnd.n5765 gnd.n1360 71.676
R13811 gnd.n5769 gnd.n1361 71.676
R13812 gnd.n5773 gnd.n1362 71.676
R13813 gnd.n5777 gnd.n1363 71.676
R13814 gnd.n5781 gnd.n1364 71.676
R13815 gnd.n5785 gnd.n1365 71.676
R13816 gnd.n5789 gnd.n1366 71.676
R13817 gnd.n5793 gnd.n1367 71.676
R13818 gnd.n5797 gnd.n1368 71.676
R13819 gnd.n5801 gnd.n1369 71.676
R13820 gnd.n5805 gnd.n1370 71.676
R13821 gnd.n5810 gnd.n1371 71.676
R13822 gnd.n5814 gnd.n1372 71.676
R13823 gnd.n5677 gnd.n1356 71.676
R13824 gnd.n5681 gnd.n1355 71.676
R13825 gnd.n5686 gnd.n1354 71.676
R13826 gnd.n5690 gnd.n1353 71.676
R13827 gnd.n5694 gnd.n1352 71.676
R13828 gnd.n5698 gnd.n1351 71.676
R13829 gnd.n5702 gnd.n1350 71.676
R13830 gnd.n5706 gnd.n1349 71.676
R13831 gnd.n5710 gnd.n1348 71.676
R13832 gnd.n5714 gnd.n1347 71.676
R13833 gnd.n5718 gnd.n1346 71.676
R13834 gnd.n5722 gnd.n1345 71.676
R13835 gnd.n5726 gnd.n1344 71.676
R13836 gnd.n5730 gnd.n1343 71.676
R13837 gnd.n5734 gnd.n1342 71.676
R13838 gnd.n5738 gnd.n1341 71.676
R13839 gnd.n5741 gnd.n1340 71.676
R13840 gnd.n10 gnd.t296 69.1507
R13841 gnd.n18 gnd.t283 68.4792
R13842 gnd.n17 gnd.t320 68.4792
R13843 gnd.n16 gnd.t318 68.4792
R13844 gnd.n15 gnd.t233 68.4792
R13845 gnd.n14 gnd.t348 68.4792
R13846 gnd.n13 gnd.t25 68.4792
R13847 gnd.n12 gnd.t23 68.4792
R13848 gnd.n11 gnd.t235 68.4792
R13849 gnd.n10 gnd.t237 68.4792
R13850 gnd.n6577 gnd.n6576 61.3075
R13851 gnd.n6578 gnd.n6577 61.3075
R13852 gnd.n6578 gnd.n724 61.3075
R13853 gnd.n6586 gnd.n724 61.3075
R13854 gnd.n6587 gnd.n6586 61.3075
R13855 gnd.n6588 gnd.n6587 61.3075
R13856 gnd.n6588 gnd.n718 61.3075
R13857 gnd.n6596 gnd.n718 61.3075
R13858 gnd.n6597 gnd.n6596 61.3075
R13859 gnd.n6598 gnd.n6597 61.3075
R13860 gnd.n6598 gnd.n712 61.3075
R13861 gnd.n6606 gnd.n712 61.3075
R13862 gnd.n6607 gnd.n6606 61.3075
R13863 gnd.n6608 gnd.n6607 61.3075
R13864 gnd.n6608 gnd.n706 61.3075
R13865 gnd.n6616 gnd.n706 61.3075
R13866 gnd.n6617 gnd.n6616 61.3075
R13867 gnd.n6618 gnd.n6617 61.3075
R13868 gnd.n6618 gnd.n700 61.3075
R13869 gnd.n6626 gnd.n700 61.3075
R13870 gnd.n6627 gnd.n6626 61.3075
R13871 gnd.n6628 gnd.n6627 61.3075
R13872 gnd.n6628 gnd.n694 61.3075
R13873 gnd.n6636 gnd.n694 61.3075
R13874 gnd.n6637 gnd.n6636 61.3075
R13875 gnd.n6638 gnd.n6637 61.3075
R13876 gnd.n6638 gnd.n688 61.3075
R13877 gnd.n6646 gnd.n688 61.3075
R13878 gnd.n6647 gnd.n6646 61.3075
R13879 gnd.n6648 gnd.n6647 61.3075
R13880 gnd.n6648 gnd.n682 61.3075
R13881 gnd.n6656 gnd.n682 61.3075
R13882 gnd.n6657 gnd.n6656 61.3075
R13883 gnd.n6658 gnd.n6657 61.3075
R13884 gnd.n6658 gnd.n676 61.3075
R13885 gnd.n6666 gnd.n676 61.3075
R13886 gnd.n6667 gnd.n6666 61.3075
R13887 gnd.n6668 gnd.n6667 61.3075
R13888 gnd.n6668 gnd.n670 61.3075
R13889 gnd.n6676 gnd.n670 61.3075
R13890 gnd.n6677 gnd.n6676 61.3075
R13891 gnd.n6678 gnd.n6677 61.3075
R13892 gnd.n6678 gnd.n664 61.3075
R13893 gnd.n6686 gnd.n664 61.3075
R13894 gnd.n6687 gnd.n6686 61.3075
R13895 gnd.n6688 gnd.n6687 61.3075
R13896 gnd.n6688 gnd.n658 61.3075
R13897 gnd.n6696 gnd.n658 61.3075
R13898 gnd.n6697 gnd.n6696 61.3075
R13899 gnd.n6698 gnd.n6697 61.3075
R13900 gnd.n6698 gnd.n652 61.3075
R13901 gnd.n6706 gnd.n652 61.3075
R13902 gnd.n6707 gnd.n6706 61.3075
R13903 gnd.n6708 gnd.n6707 61.3075
R13904 gnd.n6708 gnd.n646 61.3075
R13905 gnd.n6716 gnd.n646 61.3075
R13906 gnd.n6717 gnd.n6716 61.3075
R13907 gnd.n6718 gnd.n6717 61.3075
R13908 gnd.n6718 gnd.n640 61.3075
R13909 gnd.n6726 gnd.n640 61.3075
R13910 gnd.n6727 gnd.n6726 61.3075
R13911 gnd.n6728 gnd.n6727 61.3075
R13912 gnd.n6728 gnd.n634 61.3075
R13913 gnd.n6736 gnd.n634 61.3075
R13914 gnd.n6737 gnd.n6736 61.3075
R13915 gnd.n6738 gnd.n6737 61.3075
R13916 gnd.n6738 gnd.n628 61.3075
R13917 gnd.n6746 gnd.n628 61.3075
R13918 gnd.n6747 gnd.n6746 61.3075
R13919 gnd.n6748 gnd.n6747 61.3075
R13920 gnd.n6748 gnd.n622 61.3075
R13921 gnd.n6756 gnd.n622 61.3075
R13922 gnd.n6757 gnd.n6756 61.3075
R13923 gnd.n6758 gnd.n6757 61.3075
R13924 gnd.n6758 gnd.n616 61.3075
R13925 gnd.n6766 gnd.n616 61.3075
R13926 gnd.n6767 gnd.n6766 61.3075
R13927 gnd.n6768 gnd.n6767 61.3075
R13928 gnd.n6768 gnd.n610 61.3075
R13929 gnd.n6776 gnd.n610 61.3075
R13930 gnd.n6777 gnd.n6776 61.3075
R13931 gnd.n6780 gnd.n6777 61.3075
R13932 gnd.n6780 gnd.n6779 61.3075
R13933 gnd.n1889 gnd.n1836 59.5399
R13934 gnd.n5808 gnd.n1375 59.5399
R13935 gnd.n1834 gnd.n1833 59.5399
R13936 gnd.n5684 gnd.n5676 59.5399
R13937 gnd.n1831 gnd.n1830 59.1804
R13938 gnd.n2499 gnd.t35 56.607
R13939 gnd.n60 gnd.t225 56.607
R13940 gnd.n2460 gnd.t336 56.407
R13941 gnd.n2479 gnd.t285 56.407
R13942 gnd.n21 gnd.t252 56.407
R13943 gnd.n40 gnd.t343 56.407
R13944 gnd.n2516 gnd.t309 55.8337
R13945 gnd.n2477 gnd.t251 55.8337
R13946 gnd.n2496 gnd.t286 55.8337
R13947 gnd.n77 gnd.t303 55.8337
R13948 gnd.n38 gnd.t254 55.8337
R13949 gnd.n57 gnd.t338 55.8337
R13950 gnd.n1818 gnd.n1817 54.358
R13951 gnd.n5668 gnd.n5667 54.358
R13952 gnd.n2499 gnd.n2498 53.0052
R13953 gnd.n2501 gnd.n2500 53.0052
R13954 gnd.n2503 gnd.n2502 53.0052
R13955 gnd.n2505 gnd.n2504 53.0052
R13956 gnd.n2507 gnd.n2506 53.0052
R13957 gnd.n2509 gnd.n2508 53.0052
R13958 gnd.n2511 gnd.n2510 53.0052
R13959 gnd.n2513 gnd.n2512 53.0052
R13960 gnd.n2515 gnd.n2514 53.0052
R13961 gnd.n2460 gnd.n2459 53.0052
R13962 gnd.n2462 gnd.n2461 53.0052
R13963 gnd.n2464 gnd.n2463 53.0052
R13964 gnd.n2466 gnd.n2465 53.0052
R13965 gnd.n2468 gnd.n2467 53.0052
R13966 gnd.n2470 gnd.n2469 53.0052
R13967 gnd.n2472 gnd.n2471 53.0052
R13968 gnd.n2474 gnd.n2473 53.0052
R13969 gnd.n2476 gnd.n2475 53.0052
R13970 gnd.n2479 gnd.n2478 53.0052
R13971 gnd.n2481 gnd.n2480 53.0052
R13972 gnd.n2483 gnd.n2482 53.0052
R13973 gnd.n2485 gnd.n2484 53.0052
R13974 gnd.n2487 gnd.n2486 53.0052
R13975 gnd.n2489 gnd.n2488 53.0052
R13976 gnd.n2491 gnd.n2490 53.0052
R13977 gnd.n2493 gnd.n2492 53.0052
R13978 gnd.n2495 gnd.n2494 53.0052
R13979 gnd.n76 gnd.n75 53.0052
R13980 gnd.n74 gnd.n73 53.0052
R13981 gnd.n72 gnd.n71 53.0052
R13982 gnd.n70 gnd.n69 53.0052
R13983 gnd.n68 gnd.n67 53.0052
R13984 gnd.n66 gnd.n65 53.0052
R13985 gnd.n64 gnd.n63 53.0052
R13986 gnd.n62 gnd.n61 53.0052
R13987 gnd.n60 gnd.n59 53.0052
R13988 gnd.n37 gnd.n36 53.0052
R13989 gnd.n35 gnd.n34 53.0052
R13990 gnd.n33 gnd.n32 53.0052
R13991 gnd.n31 gnd.n30 53.0052
R13992 gnd.n29 gnd.n28 53.0052
R13993 gnd.n27 gnd.n26 53.0052
R13994 gnd.n25 gnd.n24 53.0052
R13995 gnd.n23 gnd.n22 53.0052
R13996 gnd.n21 gnd.n20 53.0052
R13997 gnd.n56 gnd.n55 53.0052
R13998 gnd.n54 gnd.n53 53.0052
R13999 gnd.n52 gnd.n51 53.0052
R14000 gnd.n50 gnd.n49 53.0052
R14001 gnd.n48 gnd.n47 53.0052
R14002 gnd.n46 gnd.n45 53.0052
R14003 gnd.n44 gnd.n43 53.0052
R14004 gnd.n42 gnd.n41 53.0052
R14005 gnd.n40 gnd.n39 53.0052
R14006 gnd.n5659 gnd.n5658 52.4801
R14007 gnd.n3552 gnd.t352 52.3082
R14008 gnd.n3520 gnd.t330 52.3082
R14009 gnd.n3488 gnd.t231 52.3082
R14010 gnd.n3457 gnd.t229 52.3082
R14011 gnd.n3425 gnd.t1 52.3082
R14012 gnd.n3393 gnd.t21 52.3082
R14013 gnd.n3361 gnd.t322 52.3082
R14014 gnd.n3330 gnd.t3 52.3082
R14015 gnd.n7553 gnd.n128 51.6227
R14016 gnd.n3382 gnd.n3350 51.4173
R14017 gnd.n3446 gnd.n3445 50.455
R14018 gnd.n3414 gnd.n3413 50.455
R14019 gnd.n3382 gnd.n3381 50.455
R14020 gnd.n2795 gnd.n2794 45.1884
R14021 gnd.n2293 gnd.n2292 45.1884
R14022 gnd.n5743 gnd.n5674 44.3322
R14023 gnd.n1821 gnd.n1820 44.3189
R14024 gnd.n4575 gnd.n4574 42.4732
R14025 gnd.n1293 gnd.n1269 42.4732
R14026 gnd.n583 gnd.n582 42.2793
R14027 gnd.n7481 gnd.n202 42.2793
R14028 gnd.n7518 gnd.n7517 42.2793
R14029 gnd.n124 gnd.n123 42.2793
R14030 gnd.n499 gnd.n498 42.2793
R14031 gnd.n4556 gnd.n4553 42.2793
R14032 gnd.n2796 gnd.n2795 42.2793
R14033 gnd.n2294 gnd.n2293 42.2793
R14034 gnd.n2722 gnd.n2721 42.2793
R14035 gnd.n3667 gnd.n2267 42.2793
R14036 gnd.n1990 gnd.n1989 42.2793
R14037 gnd.n3733 gnd.n3732 42.2793
R14038 gnd.n3709 gnd.n3708 42.2793
R14039 gnd.n4012 gnd.n4011 42.2793
R14040 gnd.n1819 gnd.n1818 41.6274
R14041 gnd.n5669 gnd.n5668 41.6274
R14042 gnd.n1828 gnd.n1827 40.8975
R14043 gnd.n5672 gnd.n5671 40.8975
R14044 gnd.n7071 gnd.n560 36.9518
R14045 gnd.n4828 gnd.n1898 36.9518
R14046 gnd.n2848 gnd.n2752 36.8252
R14047 gnd.n6779 gnd.n6778 36.7847
R14048 gnd.n1827 gnd.n1826 35.055
R14049 gnd.n1822 gnd.n1821 35.055
R14050 gnd.n5661 gnd.n5660 35.055
R14051 gnd.n5671 gnd.n5657 35.055
R14052 gnd.n5751 gnd.n1376 32.9371
R14053 gnd.n4902 gnd.n4900 32.9371
R14054 gnd.n3700 gnd.n2227 32.8146
R14055 gnd.n4767 gnd.n4477 31.8661
R14056 gnd.n4767 gnd.n4766 31.8661
R14057 gnd.n4620 gnd.n4491 31.8661
R14058 gnd.n5898 gnd.n1229 31.8661
R14059 gnd.n5892 gnd.n5891 31.8661
R14060 gnd.n5891 gnd.n506 31.8661
R14061 gnd.n7197 gnd.n401 31.8661
R14062 gnd.n7205 gnd.n401 31.8661
R14063 gnd.n7213 gnd.n393 31.8661
R14064 gnd.n7221 gnd.n384 31.8661
R14065 gnd.n7221 gnd.n387 31.8661
R14066 gnd.n7229 gnd.n369 31.8661
R14067 gnd.n7237 gnd.n369 31.8661
R14068 gnd.n7245 gnd.n361 31.8661
R14069 gnd.n7253 gnd.n352 31.8661
R14070 gnd.n7253 gnd.n355 31.8661
R14071 gnd.n7261 gnd.n337 31.8661
R14072 gnd.n7269 gnd.n337 31.8661
R14073 gnd.n7277 gnd.n329 31.8661
R14074 gnd.n7285 gnd.n319 31.8661
R14075 gnd.n7285 gnd.n322 31.8661
R14076 gnd.n7293 gnd.n313 31.8661
R14077 gnd.n7301 gnd.n298 31.8661
R14078 gnd.n7309 gnd.n298 31.8661
R14079 gnd.n7317 gnd.n289 31.8661
R14080 gnd.n7317 gnd.n292 31.8661
R14081 gnd.n7325 gnd.n283 31.8661
R14082 gnd.n7333 gnd.n268 31.8661
R14083 gnd.n7341 gnd.n268 31.8661
R14084 gnd.n7349 gnd.n259 31.8661
R14085 gnd.n7349 gnd.n262 31.8661
R14086 gnd.n7357 gnd.n253 31.8661
R14087 gnd.n7365 gnd.n238 31.8661
R14088 gnd.n7373 gnd.n238 31.8661
R14089 gnd.n7381 gnd.n229 31.8661
R14090 gnd.n7381 gnd.n232 31.8661
R14091 gnd.n7389 gnd.n213 31.8661
R14092 gnd.n7465 gnd.n213 31.8661
R14093 gnd.n7465 gnd.n206 31.8661
R14094 gnd.n7473 gnd.n206 31.8661
R14095 gnd.n7553 gnd.n126 31.8661
R14096 gnd.t214 gnd.n329 31.5474
R14097 gnd.n313 gnd.t210 31.5474
R14098 gnd.t82 gnd.n361 30.9101
R14099 gnd.t12 gnd.n393 30.2728
R14100 gnd.n253 gnd.t14 30.2728
R14101 gnd.n4192 gnd.n3701 29.5331
R14102 gnd.t90 gnd.n126 28.3609
R14103 gnd.n4773 gnd.n1960 28.0422
R14104 gnd.n7102 gnd.n450 28.0422
R14105 gnd.n1056 gnd.n921 27.1052
R14106 gnd.n4574 gnd.n4573 25.7944
R14107 gnd.n560 gnd.n559 25.7944
R14108 gnd.n582 gnd.n581 25.7944
R14109 gnd.n202 gnd.n201 25.7944
R14110 gnd.n7517 gnd.n7516 25.7944
R14111 gnd.n123 gnd.n122 25.7944
R14112 gnd.n498 gnd.n497 25.7944
R14113 gnd.n4553 gnd.n4552 25.7944
R14114 gnd.n2721 gnd.n2720 25.7944
R14115 gnd.n2267 gnd.n2266 25.7944
R14116 gnd.n1989 gnd.n1988 25.7944
R14117 gnd.n1898 gnd.n1897 25.7944
R14118 gnd.n3732 gnd.n3731 25.7944
R14119 gnd.n3708 gnd.n3707 25.7944
R14120 gnd.n4011 gnd.n4010 25.7944
R14121 gnd.n1269 gnd.n1268 25.7944
R14122 gnd.n7189 gnd.n419 25.1743
R14123 gnd.n4766 gnd.n4765 23.8997
R14124 gnd.n5892 gnd.n5890 23.8997
R14125 gnd.n1836 gnd.n1835 23.855
R14126 gnd.n1375 gnd.n1374 23.855
R14127 gnd.n1833 gnd.n1832 23.855
R14128 gnd.n5676 gnd.n5675 23.855
R14129 gnd.n4434 gnd.n1068 23.581
R14130 gnd.n6072 gnd.n1071 23.581
R14131 gnd.n4443 gnd.n1080 23.581
R14132 gnd.n6066 gnd.n1083 23.581
R14133 gnd.n6060 gnd.n1094 23.581
R14134 gnd.n4774 gnd.n4773 23.581
R14135 gnd.n7157 gnd.n450 23.581
R14136 gnd.n6800 gnd.n453 23.581
R14137 gnd.n7022 gnd.n445 23.581
R14138 gnd.n7173 gnd.n434 23.581
R14139 gnd.n6814 gnd.n437 23.581
R14140 gnd.n7181 gnd.n425 23.581
R14141 gnd.n7189 gnd.n416 23.581
R14142 gnd.n7389 gnd.t253 23.2624
R14143 gnd.n7213 gnd.t216 22.6251
R14144 gnd.n7357 gnd.t73 22.6251
R14145 gnd.n6778 gnd.t30 22.3064
R14146 gnd.n7245 gnd.t6 21.9878
R14147 gnd.n7325 gnd.t32 21.9878
R14148 gnd.n7277 gnd.t87 21.3504
R14149 gnd.n7293 gnd.t202 21.3504
R14150 gnd.n1831 gnd.n1762 20.7615
R14151 gnd.n5744 gnd.n5743 20.7615
R14152 gnd.n7261 gnd.t28 20.7131
R14153 gnd.n7309 gnd.t207 20.7131
R14154 gnd.t107 gnd.n1091 20.0758
R14155 gnd.n6799 gnd.t114 20.0758
R14156 gnd.n7229 gnd.t75 20.0758
R14157 gnd.n7341 gnd.t248 20.0758
R14158 gnd.n1815 gnd.t180 19.8005
R14159 gnd.n1815 gnd.t101 19.8005
R14160 gnd.n1816 gnd.t98 19.8005
R14161 gnd.n1816 gnd.t123 19.8005
R14162 gnd.n5665 gnd.t130 19.8005
R14163 gnd.n5665 gnd.t112 19.8005
R14164 gnd.n5666 gnd.t151 19.8005
R14165 gnd.n5666 gnd.t95 19.8005
R14166 gnd.n1812 gnd.n1811 19.5087
R14167 gnd.n1825 gnd.n1812 19.5087
R14168 gnd.n1823 gnd.n1814 19.5087
R14169 gnd.n5670 gnd.n5664 19.5087
R14170 gnd.n7197 gnd.t212 19.4385
R14171 gnd.n7373 gnd.t8 19.4385
R14172 gnd.n4698 gnd.n4697 19.3944
R14173 gnd.n4697 gnd.n4696 19.3944
R14174 gnd.n4696 gnd.n4586 19.3944
R14175 gnd.n4692 gnd.n4586 19.3944
R14176 gnd.n4692 gnd.n4691 19.3944
R14177 gnd.n4691 gnd.n4690 19.3944
R14178 gnd.n4690 gnd.n4591 19.3944
R14179 gnd.n4686 gnd.n4591 19.3944
R14180 gnd.n4686 gnd.n4685 19.3944
R14181 gnd.n4685 gnd.n4684 19.3944
R14182 gnd.n4684 gnd.n4596 19.3944
R14183 gnd.n4680 gnd.n4596 19.3944
R14184 gnd.n4680 gnd.n4679 19.3944
R14185 gnd.n4679 gnd.n4678 19.3944
R14186 gnd.n4678 gnd.n4669 19.3944
R14187 gnd.n4674 gnd.n4669 19.3944
R14188 gnd.n4674 gnd.n1742 19.3944
R14189 gnd.n4976 gnd.n1742 19.3944
R14190 gnd.n4976 gnd.n1739 19.3944
R14191 gnd.n4981 gnd.n1739 19.3944
R14192 gnd.n4981 gnd.n1740 19.3944
R14193 gnd.n1740 gnd.n1712 19.3944
R14194 gnd.n5015 gnd.n1712 19.3944
R14195 gnd.n5015 gnd.n1709 19.3944
R14196 gnd.n5056 gnd.n1709 19.3944
R14197 gnd.n5056 gnd.n1710 19.3944
R14198 gnd.n5052 gnd.n1710 19.3944
R14199 gnd.n5052 gnd.n5051 19.3944
R14200 gnd.n5051 gnd.n5050 19.3944
R14201 gnd.n5050 gnd.n5022 19.3944
R14202 gnd.n5046 gnd.n5022 19.3944
R14203 gnd.n5046 gnd.n5045 19.3944
R14204 gnd.n5045 gnd.n5044 19.3944
R14205 gnd.n5044 gnd.n5028 19.3944
R14206 gnd.n5040 gnd.n5028 19.3944
R14207 gnd.n5040 gnd.n5039 19.3944
R14208 gnd.n5039 gnd.n5038 19.3944
R14209 gnd.n5038 gnd.n5035 19.3944
R14210 gnd.n5035 gnd.n1627 19.3944
R14211 gnd.n5193 gnd.n1627 19.3944
R14212 gnd.n5193 gnd.n1624 19.3944
R14213 gnd.n5232 gnd.n1624 19.3944
R14214 gnd.n5232 gnd.n1625 19.3944
R14215 gnd.n5228 gnd.n1625 19.3944
R14216 gnd.n5228 gnd.n5227 19.3944
R14217 gnd.n5227 gnd.n5226 19.3944
R14218 gnd.n5226 gnd.n5200 19.3944
R14219 gnd.n5222 gnd.n5200 19.3944
R14220 gnd.n5222 gnd.n5221 19.3944
R14221 gnd.n5221 gnd.n5220 19.3944
R14222 gnd.n5220 gnd.n5204 19.3944
R14223 gnd.n5216 gnd.n5204 19.3944
R14224 gnd.n5216 gnd.n5215 19.3944
R14225 gnd.n5215 gnd.n5214 19.3944
R14226 gnd.n5214 gnd.n5211 19.3944
R14227 gnd.n5211 gnd.n1540 19.3944
R14228 gnd.n5370 gnd.n1540 19.3944
R14229 gnd.n5370 gnd.n1537 19.3944
R14230 gnd.n5394 gnd.n1537 19.3944
R14231 gnd.n5394 gnd.n1538 19.3944
R14232 gnd.n5390 gnd.n1538 19.3944
R14233 gnd.n5390 gnd.n5389 19.3944
R14234 gnd.n5389 gnd.n5388 19.3944
R14235 gnd.n5388 gnd.n5377 19.3944
R14236 gnd.n5384 gnd.n5377 19.3944
R14237 gnd.n5384 gnd.n5383 19.3944
R14238 gnd.n5383 gnd.n5382 19.3944
R14239 gnd.n5382 gnd.n1475 19.3944
R14240 gnd.n5503 gnd.n1475 19.3944
R14241 gnd.n5503 gnd.n1472 19.3944
R14242 gnd.n5508 gnd.n1472 19.3944
R14243 gnd.n5508 gnd.n1473 19.3944
R14244 gnd.n1473 gnd.n1448 19.3944
R14245 gnd.n5542 gnd.n1448 19.3944
R14246 gnd.n5542 gnd.n1445 19.3944
R14247 gnd.n5576 gnd.n1445 19.3944
R14248 gnd.n5576 gnd.n1446 19.3944
R14249 gnd.n5572 gnd.n1446 19.3944
R14250 gnd.n5572 gnd.n5571 19.3944
R14251 gnd.n5571 gnd.n5570 19.3944
R14252 gnd.n5570 gnd.n5550 19.3944
R14253 gnd.n5566 gnd.n5550 19.3944
R14254 gnd.n5566 gnd.n5565 19.3944
R14255 gnd.n5565 gnd.n5564 19.3944
R14256 gnd.n5564 gnd.n5559 19.3944
R14257 gnd.n5560 gnd.n5559 19.3944
R14258 gnd.n5560 gnd.n1337 19.3944
R14259 gnd.n5821 gnd.n1337 19.3944
R14260 gnd.n5821 gnd.n1335 19.3944
R14261 gnd.n5825 gnd.n1335 19.3944
R14262 gnd.n5825 gnd.n1325 19.3944
R14263 gnd.n5841 gnd.n1325 19.3944
R14264 gnd.n5841 gnd.n1323 19.3944
R14265 gnd.n5845 gnd.n1323 19.3944
R14266 gnd.n5845 gnd.n1312 19.3944
R14267 gnd.n5861 gnd.n1312 19.3944
R14268 gnd.n5861 gnd.n1310 19.3944
R14269 gnd.n5866 gnd.n1310 19.3944
R14270 gnd.n5866 gnd.n1301 19.3944
R14271 gnd.n5884 gnd.n1301 19.3944
R14272 gnd.n5885 gnd.n5884 19.3944
R14273 gnd.n4704 gnd.n4703 19.3944
R14274 gnd.n4703 gnd.n4702 19.3944
R14275 gnd.n4702 gnd.n4580 19.3944
R14276 gnd.n4762 gnd.n4761 19.3944
R14277 gnd.n4761 gnd.n4495 19.3944
R14278 gnd.n4754 gnd.n4495 19.3944
R14279 gnd.n4754 gnd.n4753 19.3944
R14280 gnd.n4753 gnd.n4512 19.3944
R14281 gnd.n4746 gnd.n4512 19.3944
R14282 gnd.n4746 gnd.n4745 19.3944
R14283 gnd.n4745 gnd.n4522 19.3944
R14284 gnd.n4738 gnd.n4522 19.3944
R14285 gnd.n4738 gnd.n4737 19.3944
R14286 gnd.n4737 gnd.n4535 19.3944
R14287 gnd.n4730 gnd.n4535 19.3944
R14288 gnd.n4730 gnd.n4729 19.3944
R14289 gnd.n4729 gnd.n4545 19.3944
R14290 gnd.n4722 gnd.n4545 19.3944
R14291 gnd.n4722 gnd.n4721 19.3944
R14292 gnd.n4721 gnd.n4562 19.3944
R14293 gnd.n4715 gnd.n4562 19.3944
R14294 gnd.n4715 gnd.n4714 19.3944
R14295 gnd.n4714 gnd.n4565 19.3944
R14296 gnd.n4710 gnd.n4565 19.3944
R14297 gnd.n4710 gnd.n4709 19.3944
R14298 gnd.n4709 gnd.n4708 19.3944
R14299 gnd.n4708 gnd.n4571 19.3944
R14300 gnd.n7099 gnd.n540 19.3944
R14301 gnd.n7099 gnd.n7098 19.3944
R14302 gnd.n7098 gnd.n7097 19.3944
R14303 gnd.n7097 gnd.n7095 19.3944
R14304 gnd.n7095 gnd.n7092 19.3944
R14305 gnd.n7092 gnd.n7091 19.3944
R14306 gnd.n7091 gnd.n7088 19.3944
R14307 gnd.n7088 gnd.n7087 19.3944
R14308 gnd.n7087 gnd.n7084 19.3944
R14309 gnd.n7084 gnd.n7083 19.3944
R14310 gnd.n7083 gnd.n7080 19.3944
R14311 gnd.n7080 gnd.n7079 19.3944
R14312 gnd.n7079 gnd.n7076 19.3944
R14313 gnd.n7076 gnd.n7075 19.3944
R14314 gnd.n7075 gnd.n7072 19.3944
R14315 gnd.n7070 gnd.n7067 19.3944
R14316 gnd.n7067 gnd.n7066 19.3944
R14317 gnd.n7066 gnd.n7063 19.3944
R14318 gnd.n7063 gnd.n7062 19.3944
R14319 gnd.n7062 gnd.n7059 19.3944
R14320 gnd.n7059 gnd.n7058 19.3944
R14321 gnd.n7058 gnd.n7055 19.3944
R14322 gnd.n7055 gnd.n7054 19.3944
R14323 gnd.n7054 gnd.n7051 19.3944
R14324 gnd.n7051 gnd.n7050 19.3944
R14325 gnd.n7050 gnd.n7047 19.3944
R14326 gnd.n7047 gnd.n7046 19.3944
R14327 gnd.n7046 gnd.n7043 19.3944
R14328 gnd.n7043 gnd.n7042 19.3944
R14329 gnd.n7042 gnd.n7039 19.3944
R14330 gnd.n7039 gnd.n7038 19.3944
R14331 gnd.n7038 gnd.n7035 19.3944
R14332 gnd.n7035 gnd.n7034 19.3944
R14333 gnd.n7027 gnd.n7026 19.3944
R14334 gnd.n7026 gnd.n7025 19.3944
R14335 gnd.n7025 gnd.n7024 19.3944
R14336 gnd.n7024 gnd.n588 19.3944
R14337 gnd.n6816 gnd.n588 19.3944
R14338 gnd.n6817 gnd.n6816 19.3944
R14339 gnd.n6820 gnd.n6817 19.3944
R14340 gnd.n6820 gnd.n6810 19.3944
R14341 gnd.n6953 gnd.n6810 19.3944
R14342 gnd.n6953 gnd.n6952 19.3944
R14343 gnd.n6952 gnd.n6951 19.3944
R14344 gnd.n6951 gnd.n6949 19.3944
R14345 gnd.n6949 gnd.n6948 19.3944
R14346 gnd.n6948 gnd.n6946 19.3944
R14347 gnd.n6946 gnd.n6945 19.3944
R14348 gnd.n6945 gnd.n6943 19.3944
R14349 gnd.n6943 gnd.n6942 19.3944
R14350 gnd.n6942 gnd.n6940 19.3944
R14351 gnd.n6940 gnd.n6939 19.3944
R14352 gnd.n6939 gnd.n6937 19.3944
R14353 gnd.n6937 gnd.n6936 19.3944
R14354 gnd.n6936 gnd.n6934 19.3944
R14355 gnd.n6934 gnd.n6933 19.3944
R14356 gnd.n6933 gnd.n6931 19.3944
R14357 gnd.n6931 gnd.n6930 19.3944
R14358 gnd.n6930 gnd.n6928 19.3944
R14359 gnd.n6928 gnd.n6927 19.3944
R14360 gnd.n6927 gnd.n6925 19.3944
R14361 gnd.n6925 gnd.n6924 19.3944
R14362 gnd.n6924 gnd.n6922 19.3944
R14363 gnd.n6922 gnd.n6921 19.3944
R14364 gnd.n6921 gnd.n6919 19.3944
R14365 gnd.n6919 gnd.n6918 19.3944
R14366 gnd.n6918 gnd.n6916 19.3944
R14367 gnd.n6916 gnd.n6915 19.3944
R14368 gnd.n6915 gnd.n6913 19.3944
R14369 gnd.n6913 gnd.n6912 19.3944
R14370 gnd.n6912 gnd.n6910 19.3944
R14371 gnd.n6910 gnd.n6909 19.3944
R14372 gnd.n6909 gnd.n6907 19.3944
R14373 gnd.n6907 gnd.n6906 19.3944
R14374 gnd.n6906 gnd.n6904 19.3944
R14375 gnd.n6904 gnd.n6903 19.3944
R14376 gnd.n6903 gnd.n6901 19.3944
R14377 gnd.n6901 gnd.n6900 19.3944
R14378 gnd.n6900 gnd.n6898 19.3944
R14379 gnd.n6898 gnd.n6897 19.3944
R14380 gnd.n6897 gnd.n6895 19.3944
R14381 gnd.n6895 gnd.n6894 19.3944
R14382 gnd.n6894 gnd.n6892 19.3944
R14383 gnd.n6892 gnd.n6891 19.3944
R14384 gnd.n6891 gnd.n6889 19.3944
R14385 gnd.n6889 gnd.n6888 19.3944
R14386 gnd.n6888 gnd.n6886 19.3944
R14387 gnd.n6886 gnd.n6885 19.3944
R14388 gnd.n6885 gnd.n6883 19.3944
R14389 gnd.n6883 gnd.n6882 19.3944
R14390 gnd.n6882 gnd.n6880 19.3944
R14391 gnd.n6880 gnd.n6879 19.3944
R14392 gnd.n6879 gnd.n6877 19.3944
R14393 gnd.n6877 gnd.n6876 19.3944
R14394 gnd.n6876 gnd.n204 19.3944
R14395 gnd.n7476 gnd.n204 19.3944
R14396 gnd.n7477 gnd.n7476 19.3944
R14397 gnd.n7515 gnd.n165 19.3944
R14398 gnd.n7510 gnd.n165 19.3944
R14399 gnd.n7510 gnd.n7509 19.3944
R14400 gnd.n7509 gnd.n7508 19.3944
R14401 gnd.n7508 gnd.n172 19.3944
R14402 gnd.n7503 gnd.n172 19.3944
R14403 gnd.n7503 gnd.n7502 19.3944
R14404 gnd.n7502 gnd.n7501 19.3944
R14405 gnd.n7501 gnd.n179 19.3944
R14406 gnd.n7496 gnd.n179 19.3944
R14407 gnd.n7496 gnd.n7495 19.3944
R14408 gnd.n7495 gnd.n7494 19.3944
R14409 gnd.n7494 gnd.n186 19.3944
R14410 gnd.n7489 gnd.n186 19.3944
R14411 gnd.n7489 gnd.n7488 19.3944
R14412 gnd.n7488 gnd.n7487 19.3944
R14413 gnd.n7487 gnd.n193 19.3944
R14414 gnd.n7482 gnd.n193 19.3944
R14415 gnd.n7548 gnd.n7547 19.3944
R14416 gnd.n7547 gnd.n7546 19.3944
R14417 gnd.n7546 gnd.n137 19.3944
R14418 gnd.n7541 gnd.n137 19.3944
R14419 gnd.n7541 gnd.n7540 19.3944
R14420 gnd.n7540 gnd.n7539 19.3944
R14421 gnd.n7539 gnd.n144 19.3944
R14422 gnd.n7534 gnd.n144 19.3944
R14423 gnd.n7534 gnd.n7533 19.3944
R14424 gnd.n7533 gnd.n7532 19.3944
R14425 gnd.n7532 gnd.n151 19.3944
R14426 gnd.n7527 gnd.n151 19.3944
R14427 gnd.n7527 gnd.n7526 19.3944
R14428 gnd.n7526 gnd.n7525 19.3944
R14429 gnd.n7525 gnd.n158 19.3944
R14430 gnd.n7520 gnd.n158 19.3944
R14431 gnd.n7520 gnd.n7519 19.3944
R14432 gnd.n7159 gnd.n447 19.3944
R14433 gnd.n7163 gnd.n447 19.3944
R14434 gnd.n7163 gnd.n432 19.3944
R14435 gnd.n7175 gnd.n432 19.3944
R14436 gnd.n7175 gnd.n430 19.3944
R14437 gnd.n7179 gnd.n430 19.3944
R14438 gnd.n7179 gnd.n414 19.3944
R14439 gnd.n7191 gnd.n414 19.3944
R14440 gnd.n7191 gnd.n412 19.3944
R14441 gnd.n7195 gnd.n412 19.3944
R14442 gnd.n7195 gnd.n399 19.3944
R14443 gnd.n7207 gnd.n399 19.3944
R14444 gnd.n7207 gnd.n397 19.3944
R14445 gnd.n7211 gnd.n397 19.3944
R14446 gnd.n7211 gnd.n382 19.3944
R14447 gnd.n7223 gnd.n382 19.3944
R14448 gnd.n7223 gnd.n380 19.3944
R14449 gnd.n7227 gnd.n380 19.3944
R14450 gnd.n7227 gnd.n367 19.3944
R14451 gnd.n7239 gnd.n367 19.3944
R14452 gnd.n7239 gnd.n365 19.3944
R14453 gnd.n7243 gnd.n365 19.3944
R14454 gnd.n7243 gnd.n350 19.3944
R14455 gnd.n7255 gnd.n350 19.3944
R14456 gnd.n7255 gnd.n348 19.3944
R14457 gnd.n7259 gnd.n348 19.3944
R14458 gnd.n7259 gnd.n335 19.3944
R14459 gnd.n7271 gnd.n335 19.3944
R14460 gnd.n7271 gnd.n333 19.3944
R14461 gnd.n7275 gnd.n333 19.3944
R14462 gnd.n7275 gnd.n317 19.3944
R14463 gnd.n7287 gnd.n317 19.3944
R14464 gnd.n7287 gnd.n315 19.3944
R14465 gnd.n7291 gnd.n315 19.3944
R14466 gnd.n7291 gnd.n303 19.3944
R14467 gnd.n7303 gnd.n303 19.3944
R14468 gnd.n7303 gnd.n301 19.3944
R14469 gnd.n7307 gnd.n301 19.3944
R14470 gnd.n7307 gnd.n287 19.3944
R14471 gnd.n7319 gnd.n287 19.3944
R14472 gnd.n7319 gnd.n285 19.3944
R14473 gnd.n7323 gnd.n285 19.3944
R14474 gnd.n7323 gnd.n273 19.3944
R14475 gnd.n7335 gnd.n273 19.3944
R14476 gnd.n7335 gnd.n271 19.3944
R14477 gnd.n7339 gnd.n271 19.3944
R14478 gnd.n7339 gnd.n257 19.3944
R14479 gnd.n7351 gnd.n257 19.3944
R14480 gnd.n7351 gnd.n255 19.3944
R14481 gnd.n7355 gnd.n255 19.3944
R14482 gnd.n7355 gnd.n243 19.3944
R14483 gnd.n7367 gnd.n243 19.3944
R14484 gnd.n7367 gnd.n241 19.3944
R14485 gnd.n7371 gnd.n241 19.3944
R14486 gnd.n7371 gnd.n227 19.3944
R14487 gnd.n7383 gnd.n227 19.3944
R14488 gnd.n7383 gnd.n225 19.3944
R14489 gnd.n7387 gnd.n225 19.3944
R14490 gnd.n7387 gnd.n211 19.3944
R14491 gnd.n7467 gnd.n211 19.3944
R14492 gnd.n7467 gnd.n209 19.3944
R14493 gnd.n7471 gnd.n209 19.3944
R14494 gnd.n7471 gnd.n132 19.3944
R14495 gnd.n7551 gnd.n132 19.3944
R14496 gnd.n6802 gnd.n592 19.3944
R14497 gnd.n6802 gnd.n589 19.3944
R14498 gnd.n7020 gnd.n589 19.3944
R14499 gnd.n7020 gnd.n590 19.3944
R14500 gnd.n7016 gnd.n590 19.3944
R14501 gnd.n7016 gnd.n7015 19.3944
R14502 gnd.n7015 gnd.n7014 19.3944
R14503 gnd.n7014 gnd.n6808 19.3944
R14504 gnd.n7010 gnd.n6808 19.3944
R14505 gnd.n7010 gnd.n7009 19.3944
R14506 gnd.n7009 gnd.n7008 19.3944
R14507 gnd.n7008 gnd.n6958 19.3944
R14508 gnd.n7004 gnd.n6958 19.3944
R14509 gnd.n7004 gnd.n7003 19.3944
R14510 gnd.n7003 gnd.n7002 19.3944
R14511 gnd.n7002 gnd.n6962 19.3944
R14512 gnd.n6998 gnd.n6962 19.3944
R14513 gnd.n6998 gnd.n6997 19.3944
R14514 gnd.n6997 gnd.n6996 19.3944
R14515 gnd.n6996 gnd.n6966 19.3944
R14516 gnd.n6992 gnd.n6966 19.3944
R14517 gnd.n6992 gnd.n6991 19.3944
R14518 gnd.n6991 gnd.n6990 19.3944
R14519 gnd.n6990 gnd.n6970 19.3944
R14520 gnd.n6986 gnd.n6970 19.3944
R14521 gnd.n6986 gnd.n6985 19.3944
R14522 gnd.n6985 gnd.n6984 19.3944
R14523 gnd.n6984 gnd.n6974 19.3944
R14524 gnd.n6980 gnd.n6974 19.3944
R14525 gnd.n6980 gnd.n6979 19.3944
R14526 gnd.n6979 gnd.n6978 19.3944
R14527 gnd.n6978 gnd.n80 19.3944
R14528 gnd.n7604 gnd.n80 19.3944
R14529 gnd.n7604 gnd.n7603 19.3944
R14530 gnd.n7603 gnd.n7602 19.3944
R14531 gnd.n7602 gnd.n85 19.3944
R14532 gnd.n7598 gnd.n85 19.3944
R14533 gnd.n7598 gnd.n7597 19.3944
R14534 gnd.n7597 gnd.n7596 19.3944
R14535 gnd.n7596 gnd.n90 19.3944
R14536 gnd.n7592 gnd.n90 19.3944
R14537 gnd.n7592 gnd.n7591 19.3944
R14538 gnd.n7591 gnd.n7590 19.3944
R14539 gnd.n7590 gnd.n95 19.3944
R14540 gnd.n7586 gnd.n95 19.3944
R14541 gnd.n7586 gnd.n7585 19.3944
R14542 gnd.n7585 gnd.n7584 19.3944
R14543 gnd.n7584 gnd.n100 19.3944
R14544 gnd.n7580 gnd.n100 19.3944
R14545 gnd.n7580 gnd.n7579 19.3944
R14546 gnd.n7579 gnd.n7578 19.3944
R14547 gnd.n7578 gnd.n105 19.3944
R14548 gnd.n7574 gnd.n105 19.3944
R14549 gnd.n7574 gnd.n7573 19.3944
R14550 gnd.n7573 gnd.n7572 19.3944
R14551 gnd.n7572 gnd.n110 19.3944
R14552 gnd.n7568 gnd.n110 19.3944
R14553 gnd.n7568 gnd.n7567 19.3944
R14554 gnd.n7567 gnd.n7566 19.3944
R14555 gnd.n7566 gnd.n115 19.3944
R14556 gnd.n7562 gnd.n115 19.3944
R14557 gnd.n7562 gnd.n7561 19.3944
R14558 gnd.n7561 gnd.n7560 19.3944
R14559 gnd.n7560 gnd.n120 19.3944
R14560 gnd.n7454 gnd.n7453 19.3944
R14561 gnd.n7453 gnd.n7452 19.3944
R14562 gnd.n7452 gnd.n7401 19.3944
R14563 gnd.n7448 gnd.n7401 19.3944
R14564 gnd.n7448 gnd.n7447 19.3944
R14565 gnd.n7447 gnd.n7446 19.3944
R14566 gnd.n7446 gnd.n7409 19.3944
R14567 gnd.n7442 gnd.n7409 19.3944
R14568 gnd.n7442 gnd.n7441 19.3944
R14569 gnd.n7441 gnd.n7440 19.3944
R14570 gnd.n7440 gnd.n7417 19.3944
R14571 gnd.n7436 gnd.n7417 19.3944
R14572 gnd.n7436 gnd.n7435 19.3944
R14573 gnd.n7435 gnd.n7434 19.3944
R14574 gnd.n7434 gnd.n7425 19.3944
R14575 gnd.n7430 gnd.n7425 19.3944
R14576 gnd.n7152 gnd.n7151 19.3944
R14577 gnd.n7151 gnd.n457 19.3944
R14578 gnd.n7144 gnd.n457 19.3944
R14579 gnd.n7144 gnd.n7143 19.3944
R14580 gnd.n7143 gnd.n465 19.3944
R14581 gnd.n7136 gnd.n465 19.3944
R14582 gnd.n7136 gnd.n7135 19.3944
R14583 gnd.n7135 gnd.n473 19.3944
R14584 gnd.n7128 gnd.n473 19.3944
R14585 gnd.n7128 gnd.n7127 19.3944
R14586 gnd.n7127 gnd.n481 19.3944
R14587 gnd.n7120 gnd.n481 19.3944
R14588 gnd.n7120 gnd.n7119 19.3944
R14589 gnd.n7119 gnd.n489 19.3944
R14590 gnd.n7112 gnd.n489 19.3944
R14591 gnd.n7112 gnd.n7111 19.3944
R14592 gnd.n7155 gnd.n441 19.3944
R14593 gnd.n7167 gnd.n441 19.3944
R14594 gnd.n7167 gnd.n439 19.3944
R14595 gnd.n7171 gnd.n439 19.3944
R14596 gnd.n7171 gnd.n423 19.3944
R14597 gnd.n7183 gnd.n423 19.3944
R14598 gnd.n7183 gnd.n421 19.3944
R14599 gnd.n7187 gnd.n421 19.3944
R14600 gnd.n7187 gnd.n407 19.3944
R14601 gnd.n7199 gnd.n407 19.3944
R14602 gnd.n7199 gnd.n405 19.3944
R14603 gnd.n7203 gnd.n405 19.3944
R14604 gnd.n7203 gnd.n391 19.3944
R14605 gnd.n7215 gnd.n391 19.3944
R14606 gnd.n7215 gnd.n389 19.3944
R14607 gnd.n7219 gnd.n389 19.3944
R14608 gnd.n7219 gnd.n375 19.3944
R14609 gnd.n7231 gnd.n375 19.3944
R14610 gnd.n7231 gnd.n373 19.3944
R14611 gnd.n7235 gnd.n373 19.3944
R14612 gnd.n7235 gnd.n359 19.3944
R14613 gnd.n7247 gnd.n359 19.3944
R14614 gnd.n7247 gnd.n357 19.3944
R14615 gnd.n7251 gnd.n357 19.3944
R14616 gnd.n7251 gnd.n343 19.3944
R14617 gnd.n7263 gnd.n343 19.3944
R14618 gnd.n7263 gnd.n341 19.3944
R14619 gnd.n7267 gnd.n341 19.3944
R14620 gnd.n7267 gnd.n327 19.3944
R14621 gnd.n7279 gnd.n327 19.3944
R14622 gnd.n7279 gnd.n324 19.3944
R14623 gnd.n7283 gnd.n324 19.3944
R14624 gnd.n7283 gnd.n310 19.3944
R14625 gnd.n7295 gnd.n310 19.3944
R14626 gnd.n7295 gnd.n308 19.3944
R14627 gnd.n7299 gnd.n308 19.3944
R14628 gnd.n7299 gnd.n296 19.3944
R14629 gnd.n7311 gnd.n296 19.3944
R14630 gnd.n7311 gnd.n294 19.3944
R14631 gnd.n7315 gnd.n294 19.3944
R14632 gnd.n7315 gnd.n280 19.3944
R14633 gnd.n7327 gnd.n280 19.3944
R14634 gnd.n7327 gnd.n278 19.3944
R14635 gnd.n7331 gnd.n278 19.3944
R14636 gnd.n7331 gnd.n266 19.3944
R14637 gnd.n7343 gnd.n266 19.3944
R14638 gnd.n7343 gnd.n264 19.3944
R14639 gnd.n7347 gnd.n264 19.3944
R14640 gnd.n7347 gnd.n250 19.3944
R14641 gnd.n7359 gnd.n250 19.3944
R14642 gnd.n7359 gnd.n248 19.3944
R14643 gnd.n7363 gnd.n248 19.3944
R14644 gnd.n7363 gnd.n236 19.3944
R14645 gnd.n7375 gnd.n236 19.3944
R14646 gnd.n7375 gnd.n234 19.3944
R14647 gnd.n7379 gnd.n234 19.3944
R14648 gnd.n7379 gnd.n221 19.3944
R14649 gnd.n7391 gnd.n221 19.3944
R14650 gnd.n7391 gnd.n218 19.3944
R14651 gnd.n7463 gnd.n218 19.3944
R14652 gnd.n7463 gnd.n219 19.3944
R14653 gnd.n7459 gnd.n219 19.3944
R14654 gnd.n7459 gnd.n7458 19.3944
R14655 gnd.n7458 gnd.n7457 19.3944
R14656 gnd.n4500 gnd.n1098 19.3944
R14657 gnd.n4500 gnd.n4498 19.3944
R14658 gnd.n4758 gnd.n4498 19.3944
R14659 gnd.n4758 gnd.n4757 19.3944
R14660 gnd.n4757 gnd.n4507 19.3944
R14661 gnd.n4750 gnd.n4507 19.3944
R14662 gnd.n4750 gnd.n4749 19.3944
R14663 gnd.n4749 gnd.n4518 19.3944
R14664 gnd.n4742 gnd.n4518 19.3944
R14665 gnd.n4742 gnd.n4741 19.3944
R14666 gnd.n4741 gnd.n4529 19.3944
R14667 gnd.n4734 gnd.n4529 19.3944
R14668 gnd.n4734 gnd.n4733 19.3944
R14669 gnd.n4733 gnd.n4541 19.3944
R14670 gnd.n4726 gnd.n4541 19.3944
R14671 gnd.n4726 gnd.n4725 19.3944
R14672 gnd.n4459 gnd.n1055 19.3944
R14673 gnd.n4461 gnd.n4459 19.3944
R14674 gnd.n4461 gnd.n4456 19.3944
R14675 gnd.n4465 gnd.n4456 19.3944
R14676 gnd.n4465 gnd.n4454 19.3944
R14677 gnd.n4469 gnd.n4454 19.3944
R14678 gnd.n4469 gnd.n4452 19.3944
R14679 gnd.n4771 gnd.n4452 19.3944
R14680 gnd.n4771 gnd.n4770 19.3944
R14681 gnd.n4770 gnd.n4769 19.3944
R14682 gnd.n4769 gnd.n4475 19.3944
R14683 gnd.n4617 gnd.n4475 19.3944
R14684 gnd.n4617 gnd.n4614 19.3944
R14685 gnd.n4626 gnd.n4614 19.3944
R14686 gnd.n4626 gnd.n4612 19.3944
R14687 gnd.n4630 gnd.n4612 19.3944
R14688 gnd.n4630 gnd.n4608 19.3944
R14689 gnd.n4642 gnd.n4608 19.3944
R14690 gnd.n4642 gnd.n4606 19.3944
R14691 gnd.n4646 gnd.n4606 19.3944
R14692 gnd.n4646 gnd.n4602 19.3944
R14693 gnd.n4658 gnd.n4602 19.3944
R14694 gnd.n4658 gnd.n4600 19.3944
R14695 gnd.n4662 gnd.n4600 19.3944
R14696 gnd.n4662 gnd.n1770 19.3944
R14697 gnd.n4908 gnd.n1770 19.3944
R14698 gnd.n4908 gnd.n1768 19.3944
R14699 gnd.n4912 gnd.n1768 19.3944
R14700 gnd.n4912 gnd.n1749 19.3944
R14701 gnd.n4967 gnd.n1749 19.3944
R14702 gnd.n4967 gnd.n1747 19.3944
R14703 gnd.n4971 gnd.n1747 19.3944
R14704 gnd.n4971 gnd.n1726 19.3944
R14705 gnd.n4995 gnd.n1726 19.3944
R14706 gnd.n4995 gnd.n1724 19.3944
R14707 gnd.n5001 gnd.n1724 19.3944
R14708 gnd.n5001 gnd.n5000 19.3944
R14709 gnd.n5000 gnd.n1698 19.3944
R14710 gnd.n5069 gnd.n1698 19.3944
R14711 gnd.n5069 gnd.n1696 19.3944
R14712 gnd.n5073 gnd.n1696 19.3944
R14713 gnd.n5073 gnd.n1678 19.3944
R14714 gnd.n5094 gnd.n1678 19.3944
R14715 gnd.n5094 gnd.n1676 19.3944
R14716 gnd.n5098 gnd.n1676 19.3944
R14717 gnd.n5098 gnd.n1658 19.3944
R14718 gnd.n5128 gnd.n1658 19.3944
R14719 gnd.n5128 gnd.n1656 19.3944
R14720 gnd.n5132 gnd.n1656 19.3944
R14721 gnd.n5132 gnd.n1641 19.3944
R14722 gnd.n5173 gnd.n1641 19.3944
R14723 gnd.n5173 gnd.n1639 19.3944
R14724 gnd.n5179 gnd.n1639 19.3944
R14725 gnd.n5179 gnd.n5178 19.3944
R14726 gnd.n5178 gnd.n1613 19.3944
R14727 gnd.n5246 gnd.n1613 19.3944
R14728 gnd.n5246 gnd.n1611 19.3944
R14729 gnd.n5250 gnd.n1611 19.3944
R14730 gnd.n5250 gnd.n1593 19.3944
R14731 gnd.n5272 gnd.n1593 19.3944
R14732 gnd.n5272 gnd.n1591 19.3944
R14733 gnd.n5276 gnd.n1591 19.3944
R14734 gnd.n5276 gnd.n1570 19.3944
R14735 gnd.n5305 gnd.n1570 19.3944
R14736 gnd.n5305 gnd.n1568 19.3944
R14737 gnd.n5309 gnd.n1568 19.3944
R14738 gnd.n5309 gnd.n1553 19.3944
R14739 gnd.n5351 gnd.n1553 19.3944
R14740 gnd.n5351 gnd.n1551 19.3944
R14741 gnd.n5357 gnd.n1551 19.3944
R14742 gnd.n5357 gnd.n5356 19.3944
R14743 gnd.n5356 gnd.n1526 19.3944
R14744 gnd.n5408 gnd.n1526 19.3944
R14745 gnd.n5408 gnd.n1524 19.3944
R14746 gnd.n5412 gnd.n1524 19.3944
R14747 gnd.n5412 gnd.n1505 19.3944
R14748 gnd.n5433 gnd.n1505 19.3944
R14749 gnd.n5433 gnd.n1503 19.3944
R14750 gnd.n5437 gnd.n1503 19.3944
R14751 gnd.n5437 gnd.n1483 19.3944
R14752 gnd.n5494 gnd.n1483 19.3944
R14753 gnd.n5494 gnd.n1481 19.3944
R14754 gnd.n5498 gnd.n1481 19.3944
R14755 gnd.n5498 gnd.n1461 19.3944
R14756 gnd.n5523 gnd.n1461 19.3944
R14757 gnd.n5523 gnd.n1459 19.3944
R14758 gnd.n5529 gnd.n1459 19.3944
R14759 gnd.n5529 gnd.n5528 19.3944
R14760 gnd.n5528 gnd.n1434 19.3944
R14761 gnd.n5589 gnd.n1434 19.3944
R14762 gnd.n5589 gnd.n1432 19.3944
R14763 gnd.n5593 gnd.n1432 19.3944
R14764 gnd.n5593 gnd.n1414 19.3944
R14765 gnd.n5614 gnd.n1414 19.3944
R14766 gnd.n5614 gnd.n1412 19.3944
R14767 gnd.n5618 gnd.n1412 19.3944
R14768 gnd.n5618 gnd.n1394 19.3944
R14769 gnd.n5642 gnd.n1394 19.3944
R14770 gnd.n5642 gnd.n1392 19.3944
R14771 gnd.n5648 gnd.n1392 19.3944
R14772 gnd.n5648 gnd.n5647 19.3944
R14773 gnd.n5647 gnd.n1332 19.3944
R14774 gnd.n5831 gnd.n1332 19.3944
R14775 gnd.n5831 gnd.n1330 19.3944
R14776 gnd.n5835 gnd.n1330 19.3944
R14777 gnd.n5835 gnd.n1319 19.3944
R14778 gnd.n5851 gnd.n1319 19.3944
R14779 gnd.n5851 gnd.n1317 19.3944
R14780 gnd.n5855 gnd.n1317 19.3944
R14781 gnd.n5855 gnd.n1306 19.3944
R14782 gnd.n5874 gnd.n1306 19.3944
R14783 gnd.n5874 gnd.n1304 19.3944
R14784 gnd.n5879 gnd.n1304 19.3944
R14785 gnd.n5879 gnd.n1232 19.3944
R14786 gnd.n5896 gnd.n1232 19.3944
R14787 gnd.n5896 gnd.n5895 19.3944
R14788 gnd.n5895 gnd.n5894 19.3944
R14789 gnd.n5894 gnd.n1236 19.3944
R14790 gnd.n1243 gnd.n1236 19.3944
R14791 gnd.n1243 gnd.n1242 19.3944
R14792 gnd.n1242 gnd.n595 19.3944
R14793 gnd.n6797 gnd.n595 19.3944
R14794 gnd.n6797 gnd.n6796 19.3944
R14795 gnd.n6796 gnd.n6795 19.3944
R14796 gnd.n6795 gnd.n599 19.3944
R14797 gnd.n6791 gnd.n599 19.3944
R14798 gnd.n6791 gnd.n6790 19.3944
R14799 gnd.n6790 gnd.n6789 19.3944
R14800 gnd.n6574 gnd.n728 19.3944
R14801 gnd.n6580 gnd.n728 19.3944
R14802 gnd.n6580 gnd.n726 19.3944
R14803 gnd.n6584 gnd.n726 19.3944
R14804 gnd.n6584 gnd.n722 19.3944
R14805 gnd.n6590 gnd.n722 19.3944
R14806 gnd.n6590 gnd.n720 19.3944
R14807 gnd.n6594 gnd.n720 19.3944
R14808 gnd.n6594 gnd.n716 19.3944
R14809 gnd.n6600 gnd.n716 19.3944
R14810 gnd.n6600 gnd.n714 19.3944
R14811 gnd.n6604 gnd.n714 19.3944
R14812 gnd.n6604 gnd.n710 19.3944
R14813 gnd.n6610 gnd.n710 19.3944
R14814 gnd.n6610 gnd.n708 19.3944
R14815 gnd.n6614 gnd.n708 19.3944
R14816 gnd.n6614 gnd.n704 19.3944
R14817 gnd.n6620 gnd.n704 19.3944
R14818 gnd.n6620 gnd.n702 19.3944
R14819 gnd.n6624 gnd.n702 19.3944
R14820 gnd.n6624 gnd.n698 19.3944
R14821 gnd.n6630 gnd.n698 19.3944
R14822 gnd.n6630 gnd.n696 19.3944
R14823 gnd.n6634 gnd.n696 19.3944
R14824 gnd.n6634 gnd.n692 19.3944
R14825 gnd.n6640 gnd.n692 19.3944
R14826 gnd.n6640 gnd.n690 19.3944
R14827 gnd.n6644 gnd.n690 19.3944
R14828 gnd.n6644 gnd.n686 19.3944
R14829 gnd.n6650 gnd.n686 19.3944
R14830 gnd.n6650 gnd.n684 19.3944
R14831 gnd.n6654 gnd.n684 19.3944
R14832 gnd.n6654 gnd.n680 19.3944
R14833 gnd.n6660 gnd.n680 19.3944
R14834 gnd.n6660 gnd.n678 19.3944
R14835 gnd.n6664 gnd.n678 19.3944
R14836 gnd.n6664 gnd.n674 19.3944
R14837 gnd.n6670 gnd.n674 19.3944
R14838 gnd.n6670 gnd.n672 19.3944
R14839 gnd.n6674 gnd.n672 19.3944
R14840 gnd.n6674 gnd.n668 19.3944
R14841 gnd.n6680 gnd.n668 19.3944
R14842 gnd.n6680 gnd.n666 19.3944
R14843 gnd.n6684 gnd.n666 19.3944
R14844 gnd.n6684 gnd.n662 19.3944
R14845 gnd.n6690 gnd.n662 19.3944
R14846 gnd.n6690 gnd.n660 19.3944
R14847 gnd.n6694 gnd.n660 19.3944
R14848 gnd.n6694 gnd.n656 19.3944
R14849 gnd.n6700 gnd.n656 19.3944
R14850 gnd.n6700 gnd.n654 19.3944
R14851 gnd.n6704 gnd.n654 19.3944
R14852 gnd.n6704 gnd.n650 19.3944
R14853 gnd.n6710 gnd.n650 19.3944
R14854 gnd.n6710 gnd.n648 19.3944
R14855 gnd.n6714 gnd.n648 19.3944
R14856 gnd.n6714 gnd.n644 19.3944
R14857 gnd.n6720 gnd.n644 19.3944
R14858 gnd.n6720 gnd.n642 19.3944
R14859 gnd.n6724 gnd.n642 19.3944
R14860 gnd.n6724 gnd.n638 19.3944
R14861 gnd.n6730 gnd.n638 19.3944
R14862 gnd.n6730 gnd.n636 19.3944
R14863 gnd.n6734 gnd.n636 19.3944
R14864 gnd.n6734 gnd.n632 19.3944
R14865 gnd.n6740 gnd.n632 19.3944
R14866 gnd.n6740 gnd.n630 19.3944
R14867 gnd.n6744 gnd.n630 19.3944
R14868 gnd.n6744 gnd.n626 19.3944
R14869 gnd.n6750 gnd.n626 19.3944
R14870 gnd.n6750 gnd.n624 19.3944
R14871 gnd.n6754 gnd.n624 19.3944
R14872 gnd.n6754 gnd.n620 19.3944
R14873 gnd.n6760 gnd.n620 19.3944
R14874 gnd.n6760 gnd.n618 19.3944
R14875 gnd.n6764 gnd.n618 19.3944
R14876 gnd.n6764 gnd.n614 19.3944
R14877 gnd.n6770 gnd.n614 19.3944
R14878 gnd.n6770 gnd.n612 19.3944
R14879 gnd.n6774 gnd.n612 19.3944
R14880 gnd.n6774 gnd.n608 19.3944
R14881 gnd.n6782 gnd.n608 19.3944
R14882 gnd.n6782 gnd.n606 19.3944
R14883 gnd.n6786 gnd.n606 19.3944
R14884 gnd.n6253 gnd.n923 19.3944
R14885 gnd.n6253 gnd.n919 19.3944
R14886 gnd.n6259 gnd.n919 19.3944
R14887 gnd.n6259 gnd.n917 19.3944
R14888 gnd.n6263 gnd.n917 19.3944
R14889 gnd.n6263 gnd.n913 19.3944
R14890 gnd.n6269 gnd.n913 19.3944
R14891 gnd.n6269 gnd.n911 19.3944
R14892 gnd.n6273 gnd.n911 19.3944
R14893 gnd.n6273 gnd.n907 19.3944
R14894 gnd.n6279 gnd.n907 19.3944
R14895 gnd.n6279 gnd.n905 19.3944
R14896 gnd.n6283 gnd.n905 19.3944
R14897 gnd.n6283 gnd.n901 19.3944
R14898 gnd.n6289 gnd.n901 19.3944
R14899 gnd.n6289 gnd.n899 19.3944
R14900 gnd.n6293 gnd.n899 19.3944
R14901 gnd.n6293 gnd.n895 19.3944
R14902 gnd.n6299 gnd.n895 19.3944
R14903 gnd.n6299 gnd.n893 19.3944
R14904 gnd.n6303 gnd.n893 19.3944
R14905 gnd.n6303 gnd.n889 19.3944
R14906 gnd.n6309 gnd.n889 19.3944
R14907 gnd.n6309 gnd.n887 19.3944
R14908 gnd.n6313 gnd.n887 19.3944
R14909 gnd.n6313 gnd.n883 19.3944
R14910 gnd.n6319 gnd.n883 19.3944
R14911 gnd.n6319 gnd.n881 19.3944
R14912 gnd.n6323 gnd.n881 19.3944
R14913 gnd.n6323 gnd.n877 19.3944
R14914 gnd.n6329 gnd.n877 19.3944
R14915 gnd.n6329 gnd.n875 19.3944
R14916 gnd.n6333 gnd.n875 19.3944
R14917 gnd.n6333 gnd.n871 19.3944
R14918 gnd.n6339 gnd.n871 19.3944
R14919 gnd.n6339 gnd.n869 19.3944
R14920 gnd.n6343 gnd.n869 19.3944
R14921 gnd.n6343 gnd.n865 19.3944
R14922 gnd.n6349 gnd.n865 19.3944
R14923 gnd.n6349 gnd.n863 19.3944
R14924 gnd.n6353 gnd.n863 19.3944
R14925 gnd.n6353 gnd.n859 19.3944
R14926 gnd.n6359 gnd.n859 19.3944
R14927 gnd.n6359 gnd.n857 19.3944
R14928 gnd.n6363 gnd.n857 19.3944
R14929 gnd.n6363 gnd.n853 19.3944
R14930 gnd.n6369 gnd.n853 19.3944
R14931 gnd.n6369 gnd.n851 19.3944
R14932 gnd.n6373 gnd.n851 19.3944
R14933 gnd.n6373 gnd.n847 19.3944
R14934 gnd.n6379 gnd.n847 19.3944
R14935 gnd.n6379 gnd.n845 19.3944
R14936 gnd.n6383 gnd.n845 19.3944
R14937 gnd.n6383 gnd.n841 19.3944
R14938 gnd.n6389 gnd.n841 19.3944
R14939 gnd.n6389 gnd.n839 19.3944
R14940 gnd.n6393 gnd.n839 19.3944
R14941 gnd.n6393 gnd.n835 19.3944
R14942 gnd.n6399 gnd.n835 19.3944
R14943 gnd.n6399 gnd.n833 19.3944
R14944 gnd.n6403 gnd.n833 19.3944
R14945 gnd.n6403 gnd.n829 19.3944
R14946 gnd.n6409 gnd.n829 19.3944
R14947 gnd.n6409 gnd.n827 19.3944
R14948 gnd.n6413 gnd.n827 19.3944
R14949 gnd.n6413 gnd.n823 19.3944
R14950 gnd.n6419 gnd.n823 19.3944
R14951 gnd.n6419 gnd.n821 19.3944
R14952 gnd.n6423 gnd.n821 19.3944
R14953 gnd.n6423 gnd.n817 19.3944
R14954 gnd.n6429 gnd.n817 19.3944
R14955 gnd.n6429 gnd.n815 19.3944
R14956 gnd.n6433 gnd.n815 19.3944
R14957 gnd.n6433 gnd.n811 19.3944
R14958 gnd.n6439 gnd.n811 19.3944
R14959 gnd.n6439 gnd.n809 19.3944
R14960 gnd.n6443 gnd.n809 19.3944
R14961 gnd.n6443 gnd.n805 19.3944
R14962 gnd.n6449 gnd.n805 19.3944
R14963 gnd.n6449 gnd.n803 19.3944
R14964 gnd.n6453 gnd.n803 19.3944
R14965 gnd.n6453 gnd.n799 19.3944
R14966 gnd.n6459 gnd.n799 19.3944
R14967 gnd.n6459 gnd.n797 19.3944
R14968 gnd.n6463 gnd.n797 19.3944
R14969 gnd.n6463 gnd.n793 19.3944
R14970 gnd.n6469 gnd.n793 19.3944
R14971 gnd.n6469 gnd.n791 19.3944
R14972 gnd.n6473 gnd.n791 19.3944
R14973 gnd.n6473 gnd.n787 19.3944
R14974 gnd.n6479 gnd.n787 19.3944
R14975 gnd.n6479 gnd.n785 19.3944
R14976 gnd.n6483 gnd.n785 19.3944
R14977 gnd.n6483 gnd.n781 19.3944
R14978 gnd.n6489 gnd.n781 19.3944
R14979 gnd.n6489 gnd.n779 19.3944
R14980 gnd.n6493 gnd.n779 19.3944
R14981 gnd.n6493 gnd.n775 19.3944
R14982 gnd.n6499 gnd.n775 19.3944
R14983 gnd.n6499 gnd.n773 19.3944
R14984 gnd.n6503 gnd.n773 19.3944
R14985 gnd.n6503 gnd.n769 19.3944
R14986 gnd.n6509 gnd.n769 19.3944
R14987 gnd.n6509 gnd.n767 19.3944
R14988 gnd.n6513 gnd.n767 19.3944
R14989 gnd.n6513 gnd.n763 19.3944
R14990 gnd.n6519 gnd.n763 19.3944
R14991 gnd.n6519 gnd.n761 19.3944
R14992 gnd.n6523 gnd.n761 19.3944
R14993 gnd.n6523 gnd.n757 19.3944
R14994 gnd.n6529 gnd.n757 19.3944
R14995 gnd.n6529 gnd.n755 19.3944
R14996 gnd.n6533 gnd.n755 19.3944
R14997 gnd.n6533 gnd.n751 19.3944
R14998 gnd.n6539 gnd.n751 19.3944
R14999 gnd.n6539 gnd.n749 19.3944
R15000 gnd.n6543 gnd.n749 19.3944
R15001 gnd.n6543 gnd.n745 19.3944
R15002 gnd.n6549 gnd.n745 19.3944
R15003 gnd.n6549 gnd.n743 19.3944
R15004 gnd.n6553 gnd.n743 19.3944
R15005 gnd.n6553 gnd.n739 19.3944
R15006 gnd.n6559 gnd.n739 19.3944
R15007 gnd.n6559 gnd.n737 19.3944
R15008 gnd.n6564 gnd.n737 19.3944
R15009 gnd.n6564 gnd.n733 19.3944
R15010 gnd.n6570 gnd.n733 19.3944
R15011 gnd.n6571 gnd.n6570 19.3944
R15012 gnd.n6249 gnd.n925 19.3944
R15013 gnd.n6244 gnd.n925 19.3944
R15014 gnd.n6244 gnd.n6243 19.3944
R15015 gnd.n6243 gnd.n6242 19.3944
R15016 gnd.n6242 gnd.n6239 19.3944
R15017 gnd.n6239 gnd.n6238 19.3944
R15018 gnd.n6238 gnd.n6235 19.3944
R15019 gnd.n6235 gnd.n6234 19.3944
R15020 gnd.n6234 gnd.n6231 19.3944
R15021 gnd.n6231 gnd.n6230 19.3944
R15022 gnd.n6230 gnd.n6227 19.3944
R15023 gnd.n6227 gnd.n6226 19.3944
R15024 gnd.n6226 gnd.n6223 19.3944
R15025 gnd.n6223 gnd.n6222 19.3944
R15026 gnd.n6222 gnd.n6219 19.3944
R15027 gnd.n6219 gnd.n6218 19.3944
R15028 gnd.n6218 gnd.n6215 19.3944
R15029 gnd.n6215 gnd.n6214 19.3944
R15030 gnd.n6214 gnd.n6211 19.3944
R15031 gnd.n6211 gnd.n6210 19.3944
R15032 gnd.n6210 gnd.n6207 19.3944
R15033 gnd.n6207 gnd.n6206 19.3944
R15034 gnd.n6206 gnd.n6203 19.3944
R15035 gnd.n6203 gnd.n6202 19.3944
R15036 gnd.n6202 gnd.n6199 19.3944
R15037 gnd.n6199 gnd.n6198 19.3944
R15038 gnd.n6198 gnd.n6195 19.3944
R15039 gnd.n6195 gnd.n6194 19.3944
R15040 gnd.n6194 gnd.n6191 19.3944
R15041 gnd.n6191 gnd.n6190 19.3944
R15042 gnd.n6190 gnd.n6187 19.3944
R15043 gnd.n6187 gnd.n6186 19.3944
R15044 gnd.n6186 gnd.n6183 19.3944
R15045 gnd.n6183 gnd.n6182 19.3944
R15046 gnd.n6182 gnd.n6179 19.3944
R15047 gnd.n6179 gnd.n6178 19.3944
R15048 gnd.n6178 gnd.n6175 19.3944
R15049 gnd.n6175 gnd.n6174 19.3944
R15050 gnd.n6174 gnd.n6171 19.3944
R15051 gnd.n6171 gnd.n6170 19.3944
R15052 gnd.n6170 gnd.n6167 19.3944
R15053 gnd.n6167 gnd.n6166 19.3944
R15054 gnd.n6166 gnd.n6163 19.3944
R15055 gnd.n6163 gnd.n6162 19.3944
R15056 gnd.n6162 gnd.n6159 19.3944
R15057 gnd.n6159 gnd.n6158 19.3944
R15058 gnd.n6158 gnd.n6155 19.3944
R15059 gnd.n6155 gnd.n6154 19.3944
R15060 gnd.n6154 gnd.n6151 19.3944
R15061 gnd.n6151 gnd.n6150 19.3944
R15062 gnd.n6150 gnd.n6147 19.3944
R15063 gnd.n6147 gnd.n6146 19.3944
R15064 gnd.n6146 gnd.n6143 19.3944
R15065 gnd.n6143 gnd.n6142 19.3944
R15066 gnd.n6142 gnd.n6139 19.3944
R15067 gnd.n6139 gnd.n6138 19.3944
R15068 gnd.n6138 gnd.n6135 19.3944
R15069 gnd.n6135 gnd.n6134 19.3944
R15070 gnd.n6134 gnd.n6131 19.3944
R15071 gnd.n6131 gnd.n6130 19.3944
R15072 gnd.n6130 gnd.n6127 19.3944
R15073 gnd.n6127 gnd.n6126 19.3944
R15074 gnd.n6126 gnd.n6123 19.3944
R15075 gnd.n6123 gnd.n6122 19.3944
R15076 gnd.n6122 gnd.n6119 19.3944
R15077 gnd.n6119 gnd.n6118 19.3944
R15078 gnd.n6118 gnd.n6115 19.3944
R15079 gnd.n6115 gnd.n6114 19.3944
R15080 gnd.n6114 gnd.n6111 19.3944
R15081 gnd.n6111 gnd.n6110 19.3944
R15082 gnd.n6110 gnd.n6107 19.3944
R15083 gnd.n6107 gnd.n6106 19.3944
R15084 gnd.n6106 gnd.n6103 19.3944
R15085 gnd.n6103 gnd.n6102 19.3944
R15086 gnd.n6102 gnd.n6099 19.3944
R15087 gnd.n6099 gnd.n6098 19.3944
R15088 gnd.n6098 gnd.n6095 19.3944
R15089 gnd.n6095 gnd.n6094 19.3944
R15090 gnd.n6094 gnd.n6091 19.3944
R15091 gnd.n6091 gnd.n6090 19.3944
R15092 gnd.n6090 gnd.n6087 19.3944
R15093 gnd.n6087 gnd.n6086 19.3944
R15094 gnd.n6086 gnd.n6083 19.3944
R15095 gnd.n6083 gnd.n6082 19.3944
R15096 gnd.n2845 gnd.n2844 19.3944
R15097 gnd.n2844 gnd.n2843 19.3944
R15098 gnd.n2843 gnd.n2842 19.3944
R15099 gnd.n2842 gnd.n2840 19.3944
R15100 gnd.n2840 gnd.n2837 19.3944
R15101 gnd.n2837 gnd.n2836 19.3944
R15102 gnd.n2836 gnd.n2833 19.3944
R15103 gnd.n2833 gnd.n2832 19.3944
R15104 gnd.n2832 gnd.n2829 19.3944
R15105 gnd.n2829 gnd.n2828 19.3944
R15106 gnd.n2828 gnd.n2825 19.3944
R15107 gnd.n2825 gnd.n2824 19.3944
R15108 gnd.n2824 gnd.n2821 19.3944
R15109 gnd.n2821 gnd.n2820 19.3944
R15110 gnd.n2820 gnd.n2817 19.3944
R15111 gnd.n2817 gnd.n2816 19.3944
R15112 gnd.n2816 gnd.n2813 19.3944
R15113 gnd.n2813 gnd.n2812 19.3944
R15114 gnd.n2812 gnd.n2809 19.3944
R15115 gnd.n2809 gnd.n2808 19.3944
R15116 gnd.n2808 gnd.n2805 19.3944
R15117 gnd.n2805 gnd.n2804 19.3944
R15118 gnd.n2801 gnd.n2800 19.3944
R15119 gnd.n2800 gnd.n2756 19.3944
R15120 gnd.n2851 gnd.n2756 19.3944
R15121 gnd.n3617 gnd.n3616 19.3944
R15122 gnd.n3616 gnd.n3613 19.3944
R15123 gnd.n3613 gnd.n3612 19.3944
R15124 gnd.n3662 gnd.n3661 19.3944
R15125 gnd.n3661 gnd.n3660 19.3944
R15126 gnd.n3660 gnd.n3657 19.3944
R15127 gnd.n3657 gnd.n3656 19.3944
R15128 gnd.n3656 gnd.n3653 19.3944
R15129 gnd.n3653 gnd.n3652 19.3944
R15130 gnd.n3652 gnd.n3649 19.3944
R15131 gnd.n3649 gnd.n3648 19.3944
R15132 gnd.n3648 gnd.n3645 19.3944
R15133 gnd.n3645 gnd.n3644 19.3944
R15134 gnd.n3644 gnd.n3641 19.3944
R15135 gnd.n3641 gnd.n3640 19.3944
R15136 gnd.n3640 gnd.n3637 19.3944
R15137 gnd.n3637 gnd.n3636 19.3944
R15138 gnd.n3636 gnd.n3633 19.3944
R15139 gnd.n3633 gnd.n3632 19.3944
R15140 gnd.n3632 gnd.n3629 19.3944
R15141 gnd.n3629 gnd.n3628 19.3944
R15142 gnd.n3628 gnd.n3625 19.3944
R15143 gnd.n3625 gnd.n3624 19.3944
R15144 gnd.n3624 gnd.n3621 19.3944
R15145 gnd.n3621 gnd.n3620 19.3944
R15146 gnd.n2944 gnd.n2653 19.3944
R15147 gnd.n2954 gnd.n2653 19.3944
R15148 gnd.n2955 gnd.n2954 19.3944
R15149 gnd.n2955 gnd.n2634 19.3944
R15150 gnd.n2975 gnd.n2634 19.3944
R15151 gnd.n2975 gnd.n2626 19.3944
R15152 gnd.n2985 gnd.n2626 19.3944
R15153 gnd.n2986 gnd.n2985 19.3944
R15154 gnd.n2987 gnd.n2986 19.3944
R15155 gnd.n2987 gnd.n2609 19.3944
R15156 gnd.n3004 gnd.n2609 19.3944
R15157 gnd.n3007 gnd.n3004 19.3944
R15158 gnd.n3007 gnd.n3006 19.3944
R15159 gnd.n3006 gnd.n2582 19.3944
R15160 gnd.n3046 gnd.n2582 19.3944
R15161 gnd.n3046 gnd.n2579 19.3944
R15162 gnd.n3052 gnd.n2579 19.3944
R15163 gnd.n3053 gnd.n3052 19.3944
R15164 gnd.n3053 gnd.n2577 19.3944
R15165 gnd.n3059 gnd.n2577 19.3944
R15166 gnd.n3062 gnd.n3059 19.3944
R15167 gnd.n3064 gnd.n3062 19.3944
R15168 gnd.n3070 gnd.n3064 19.3944
R15169 gnd.n3070 gnd.n3069 19.3944
R15170 gnd.n3069 gnd.n2440 19.3944
R15171 gnd.n3136 gnd.n2440 19.3944
R15172 gnd.n3137 gnd.n3136 19.3944
R15173 gnd.n3137 gnd.n2433 19.3944
R15174 gnd.n3148 gnd.n2433 19.3944
R15175 gnd.n3149 gnd.n3148 19.3944
R15176 gnd.n3149 gnd.n2416 19.3944
R15177 gnd.n2416 gnd.n2414 19.3944
R15178 gnd.n3173 gnd.n2414 19.3944
R15179 gnd.n3174 gnd.n3173 19.3944
R15180 gnd.n3174 gnd.n2385 19.3944
R15181 gnd.n3221 gnd.n2385 19.3944
R15182 gnd.n3222 gnd.n3221 19.3944
R15183 gnd.n3222 gnd.n2378 19.3944
R15184 gnd.n3233 gnd.n2378 19.3944
R15185 gnd.n3234 gnd.n3233 19.3944
R15186 gnd.n3234 gnd.n2361 19.3944
R15187 gnd.n2361 gnd.n2359 19.3944
R15188 gnd.n3258 gnd.n2359 19.3944
R15189 gnd.n3259 gnd.n3258 19.3944
R15190 gnd.n3259 gnd.n2331 19.3944
R15191 gnd.n3310 gnd.n2331 19.3944
R15192 gnd.n3311 gnd.n3310 19.3944
R15193 gnd.n3311 gnd.n2324 19.3944
R15194 gnd.n3578 gnd.n2324 19.3944
R15195 gnd.n3579 gnd.n3578 19.3944
R15196 gnd.n3579 gnd.n2305 19.3944
R15197 gnd.n3604 gnd.n2305 19.3944
R15198 gnd.n3604 gnd.n2306 19.3944
R15199 gnd.n2935 gnd.n2934 19.3944
R15200 gnd.n2934 gnd.n2667 19.3944
R15201 gnd.n2690 gnd.n2667 19.3944
R15202 gnd.n2693 gnd.n2690 19.3944
R15203 gnd.n2693 gnd.n2686 19.3944
R15204 gnd.n2697 gnd.n2686 19.3944
R15205 gnd.n2700 gnd.n2697 19.3944
R15206 gnd.n2703 gnd.n2700 19.3944
R15207 gnd.n2703 gnd.n2684 19.3944
R15208 gnd.n2707 gnd.n2684 19.3944
R15209 gnd.n2710 gnd.n2707 19.3944
R15210 gnd.n2713 gnd.n2710 19.3944
R15211 gnd.n2713 gnd.n2682 19.3944
R15212 gnd.n2717 gnd.n2682 19.3944
R15213 gnd.n2940 gnd.n2939 19.3944
R15214 gnd.n2939 gnd.n2643 19.3944
R15215 gnd.n2965 gnd.n2643 19.3944
R15216 gnd.n2965 gnd.n2641 19.3944
R15217 gnd.n2971 gnd.n2641 19.3944
R15218 gnd.n2971 gnd.n2970 19.3944
R15219 gnd.n2970 gnd.n2615 19.3944
R15220 gnd.n2995 gnd.n2615 19.3944
R15221 gnd.n2995 gnd.n2613 19.3944
R15222 gnd.n2999 gnd.n2613 19.3944
R15223 gnd.n2999 gnd.n2593 19.3944
R15224 gnd.n3026 gnd.n2593 19.3944
R15225 gnd.n3026 gnd.n2591 19.3944
R15226 gnd.n3036 gnd.n2591 19.3944
R15227 gnd.n3036 gnd.n3035 19.3944
R15228 gnd.n3035 gnd.n3034 19.3944
R15229 gnd.n3034 gnd.n2540 19.3944
R15230 gnd.n3084 gnd.n2540 19.3944
R15231 gnd.n3084 gnd.n3083 19.3944
R15232 gnd.n3083 gnd.n3082 19.3944
R15233 gnd.n3082 gnd.n2544 19.3944
R15234 gnd.n2564 gnd.n2544 19.3944
R15235 gnd.n2564 gnd.n2450 19.3944
R15236 gnd.n3121 gnd.n2450 19.3944
R15237 gnd.n3121 gnd.n2448 19.3944
R15238 gnd.n3127 gnd.n2448 19.3944
R15239 gnd.n3127 gnd.n3126 19.3944
R15240 gnd.n3126 gnd.n2423 19.3944
R15241 gnd.n3161 gnd.n2423 19.3944
R15242 gnd.n3161 gnd.n2421 19.3944
R15243 gnd.n3167 gnd.n2421 19.3944
R15244 gnd.n3167 gnd.n3166 19.3944
R15245 gnd.n3166 gnd.n2396 19.3944
R15246 gnd.n3206 gnd.n2396 19.3944
R15247 gnd.n3206 gnd.n2394 19.3944
R15248 gnd.n3212 gnd.n2394 19.3944
R15249 gnd.n3212 gnd.n3211 19.3944
R15250 gnd.n3211 gnd.n2368 19.3944
R15251 gnd.n3246 gnd.n2368 19.3944
R15252 gnd.n3246 gnd.n2366 19.3944
R15253 gnd.n3252 gnd.n2366 19.3944
R15254 gnd.n3252 gnd.n3251 19.3944
R15255 gnd.n3251 gnd.n2341 19.3944
R15256 gnd.n3295 gnd.n2341 19.3944
R15257 gnd.n3295 gnd.n2339 19.3944
R15258 gnd.n3301 gnd.n2339 19.3944
R15259 gnd.n3301 gnd.n3300 19.3944
R15260 gnd.n3300 gnd.n2314 19.3944
R15261 gnd.n3589 gnd.n2314 19.3944
R15262 gnd.n3589 gnd.n2312 19.3944
R15263 gnd.n3597 gnd.n2312 19.3944
R15264 gnd.n3597 gnd.n3596 19.3944
R15265 gnd.n3596 gnd.n3595 19.3944
R15266 gnd.n3698 gnd.n3697 19.3944
R15267 gnd.n3697 gnd.n2253 19.3944
R15268 gnd.n3693 gnd.n2253 19.3944
R15269 gnd.n3693 gnd.n3690 19.3944
R15270 gnd.n3690 gnd.n3687 19.3944
R15271 gnd.n3687 gnd.n3686 19.3944
R15272 gnd.n3686 gnd.n3683 19.3944
R15273 gnd.n3683 gnd.n3682 19.3944
R15274 gnd.n3682 gnd.n3679 19.3944
R15275 gnd.n3679 gnd.n3678 19.3944
R15276 gnd.n3678 gnd.n3675 19.3944
R15277 gnd.n3675 gnd.n3674 19.3944
R15278 gnd.n3674 gnd.n3671 19.3944
R15279 gnd.n3671 gnd.n3670 19.3944
R15280 gnd.n2855 gnd.n2754 19.3944
R15281 gnd.n2855 gnd.n2745 19.3944
R15282 gnd.n2868 gnd.n2745 19.3944
R15283 gnd.n2868 gnd.n2743 19.3944
R15284 gnd.n2872 gnd.n2743 19.3944
R15285 gnd.n2872 gnd.n2733 19.3944
R15286 gnd.n2884 gnd.n2733 19.3944
R15287 gnd.n2884 gnd.n2731 19.3944
R15288 gnd.n2918 gnd.n2731 19.3944
R15289 gnd.n2918 gnd.n2917 19.3944
R15290 gnd.n2917 gnd.n2916 19.3944
R15291 gnd.n2916 gnd.n2915 19.3944
R15292 gnd.n2915 gnd.n2912 19.3944
R15293 gnd.n2912 gnd.n2911 19.3944
R15294 gnd.n2911 gnd.n2910 19.3944
R15295 gnd.n2910 gnd.n2908 19.3944
R15296 gnd.n2908 gnd.n2907 19.3944
R15297 gnd.n2907 gnd.n2904 19.3944
R15298 gnd.n2904 gnd.n2903 19.3944
R15299 gnd.n2903 gnd.n2902 19.3944
R15300 gnd.n2902 gnd.n2900 19.3944
R15301 gnd.n2900 gnd.n2599 19.3944
R15302 gnd.n3015 gnd.n2599 19.3944
R15303 gnd.n3015 gnd.n2597 19.3944
R15304 gnd.n3021 gnd.n2597 19.3944
R15305 gnd.n3021 gnd.n3020 19.3944
R15306 gnd.n3020 gnd.n2521 19.3944
R15307 gnd.n3095 gnd.n2521 19.3944
R15308 gnd.n3095 gnd.n2522 19.3944
R15309 gnd.n2569 gnd.n2568 19.3944
R15310 gnd.n2572 gnd.n2571 19.3944
R15311 gnd.n2559 gnd.n2558 19.3944
R15312 gnd.n3114 gnd.n2455 19.3944
R15313 gnd.n3114 gnd.n3113 19.3944
R15314 gnd.n3113 gnd.n3112 19.3944
R15315 gnd.n3112 gnd.n3110 19.3944
R15316 gnd.n3110 gnd.n3109 19.3944
R15317 gnd.n3109 gnd.n3107 19.3944
R15318 gnd.n3107 gnd.n3106 19.3944
R15319 gnd.n3106 gnd.n2404 19.3944
R15320 gnd.n3182 gnd.n2404 19.3944
R15321 gnd.n3182 gnd.n2402 19.3944
R15322 gnd.n3201 gnd.n2402 19.3944
R15323 gnd.n3201 gnd.n3200 19.3944
R15324 gnd.n3200 gnd.n3199 19.3944
R15325 gnd.n3199 gnd.n3197 19.3944
R15326 gnd.n3197 gnd.n3196 19.3944
R15327 gnd.n3196 gnd.n3194 19.3944
R15328 gnd.n3194 gnd.n3193 19.3944
R15329 gnd.n3193 gnd.n2348 19.3944
R15330 gnd.n3267 gnd.n2348 19.3944
R15331 gnd.n3267 gnd.n2346 19.3944
R15332 gnd.n3290 gnd.n2346 19.3944
R15333 gnd.n3290 gnd.n3289 19.3944
R15334 gnd.n3289 gnd.n3288 19.3944
R15335 gnd.n3288 gnd.n3285 19.3944
R15336 gnd.n3285 gnd.n3284 19.3944
R15337 gnd.n3284 gnd.n3282 19.3944
R15338 gnd.n3282 gnd.n3281 19.3944
R15339 gnd.n3281 gnd.n3279 19.3944
R15340 gnd.n3279 gnd.n2300 19.3944
R15341 gnd.n2860 gnd.n2750 19.3944
R15342 gnd.n2860 gnd.n2748 19.3944
R15343 gnd.n2864 gnd.n2748 19.3944
R15344 gnd.n2864 gnd.n2739 19.3944
R15345 gnd.n2876 gnd.n2739 19.3944
R15346 gnd.n2876 gnd.n2737 19.3944
R15347 gnd.n2880 gnd.n2737 19.3944
R15348 gnd.n2880 gnd.n2726 19.3944
R15349 gnd.n2922 gnd.n2726 19.3944
R15350 gnd.n2922 gnd.n2680 19.3944
R15351 gnd.n2928 gnd.n2680 19.3944
R15352 gnd.n2928 gnd.n2927 19.3944
R15353 gnd.n2927 gnd.n2658 19.3944
R15354 gnd.n2949 gnd.n2658 19.3944
R15355 gnd.n2949 gnd.n2651 19.3944
R15356 gnd.n2960 gnd.n2651 19.3944
R15357 gnd.n2960 gnd.n2959 19.3944
R15358 gnd.n2959 gnd.n2632 19.3944
R15359 gnd.n2980 gnd.n2632 19.3944
R15360 gnd.n2980 gnd.n2622 19.3944
R15361 gnd.n2990 gnd.n2622 19.3944
R15362 gnd.n2990 gnd.n2605 19.3944
R15363 gnd.n3011 gnd.n2605 19.3944
R15364 gnd.n3011 gnd.n3010 19.3944
R15365 gnd.n3010 gnd.n2584 19.3944
R15366 gnd.n3041 gnd.n2584 19.3944
R15367 gnd.n3041 gnd.n2529 19.3944
R15368 gnd.n3091 gnd.n2529 19.3944
R15369 gnd.n3091 gnd.n3090 19.3944
R15370 gnd.n3090 gnd.n3089 19.3944
R15371 gnd.n3089 gnd.n2533 19.3944
R15372 gnd.n2551 gnd.n2533 19.3944
R15373 gnd.n3077 gnd.n2551 19.3944
R15374 gnd.n3077 gnd.n3076 19.3944
R15375 gnd.n3076 gnd.n3075 19.3944
R15376 gnd.n3075 gnd.n2555 19.3944
R15377 gnd.n2555 gnd.n2442 19.3944
R15378 gnd.n3132 gnd.n2442 19.3944
R15379 gnd.n3132 gnd.n2435 19.3944
R15380 gnd.n3143 gnd.n2435 19.3944
R15381 gnd.n3143 gnd.n2431 19.3944
R15382 gnd.n3156 gnd.n2431 19.3944
R15383 gnd.n3156 gnd.n3155 19.3944
R15384 gnd.n3155 gnd.n2410 19.3944
R15385 gnd.n3178 gnd.n2410 19.3944
R15386 gnd.n3178 gnd.n3177 19.3944
R15387 gnd.n3177 gnd.n2387 19.3944
R15388 gnd.n3217 gnd.n2387 19.3944
R15389 gnd.n3217 gnd.n2380 19.3944
R15390 gnd.n3228 gnd.n2380 19.3944
R15391 gnd.n3228 gnd.n2376 19.3944
R15392 gnd.n3241 gnd.n2376 19.3944
R15393 gnd.n3241 gnd.n3240 19.3944
R15394 gnd.n3240 gnd.n2355 19.3944
R15395 gnd.n3263 gnd.n2355 19.3944
R15396 gnd.n3263 gnd.n3262 19.3944
R15397 gnd.n3262 gnd.n2333 19.3944
R15398 gnd.n3306 gnd.n2333 19.3944
R15399 gnd.n3306 gnd.n2326 19.3944
R15400 gnd.n3317 gnd.n2326 19.3944
R15401 gnd.n3317 gnd.n2322 19.3944
R15402 gnd.n3584 gnd.n2322 19.3944
R15403 gnd.n3584 gnd.n3583 19.3944
R15404 gnd.n3583 gnd.n2303 19.3944
R15405 gnd.n3607 gnd.n2303 19.3944
R15406 gnd.n3983 gnd.n3704 19.3944
R15407 gnd.n3983 gnd.n3705 19.3944
R15408 gnd.n3979 gnd.n3705 19.3944
R15409 gnd.n3979 gnd.n3977 19.3944
R15410 gnd.n3977 gnd.n3976 19.3944
R15411 gnd.n3976 gnd.n3974 19.3944
R15412 gnd.n3974 gnd.n3973 19.3944
R15413 gnd.n3973 gnd.n3971 19.3944
R15414 gnd.n3971 gnd.n3970 19.3944
R15415 gnd.n3970 gnd.n3968 19.3944
R15416 gnd.n3968 gnd.n3967 19.3944
R15417 gnd.n3967 gnd.n3965 19.3944
R15418 gnd.n3965 gnd.n3964 19.3944
R15419 gnd.n3964 gnd.n3962 19.3944
R15420 gnd.n3962 gnd.n3961 19.3944
R15421 gnd.n3961 gnd.n3959 19.3944
R15422 gnd.n3959 gnd.n3958 19.3944
R15423 gnd.n3958 gnd.n3956 19.3944
R15424 gnd.n3956 gnd.n3955 19.3944
R15425 gnd.n3955 gnd.n3953 19.3944
R15426 gnd.n3953 gnd.n3952 19.3944
R15427 gnd.n3952 gnd.n3950 19.3944
R15428 gnd.n3950 gnd.n3949 19.3944
R15429 gnd.n3949 gnd.n3947 19.3944
R15430 gnd.n3947 gnd.n3946 19.3944
R15431 gnd.n3946 gnd.n3944 19.3944
R15432 gnd.n3944 gnd.n3943 19.3944
R15433 gnd.n3943 gnd.n3941 19.3944
R15434 gnd.n3941 gnd.n3940 19.3944
R15435 gnd.n3940 gnd.n3938 19.3944
R15436 gnd.n3938 gnd.n3937 19.3944
R15437 gnd.n3937 gnd.n3935 19.3944
R15438 gnd.n3935 gnd.n3934 19.3944
R15439 gnd.n3934 gnd.n3932 19.3944
R15440 gnd.n3932 gnd.n3931 19.3944
R15441 gnd.n3931 gnd.n3929 19.3944
R15442 gnd.n3929 gnd.n3928 19.3944
R15443 gnd.n3928 gnd.n3926 19.3944
R15444 gnd.n3926 gnd.n3925 19.3944
R15445 gnd.n3925 gnd.n3923 19.3944
R15446 gnd.n3923 gnd.n3922 19.3944
R15447 gnd.n3922 gnd.n3920 19.3944
R15448 gnd.n3920 gnd.n3919 19.3944
R15449 gnd.n3919 gnd.n3917 19.3944
R15450 gnd.n3917 gnd.n3916 19.3944
R15451 gnd.n3916 gnd.n3914 19.3944
R15452 gnd.n3914 gnd.n3913 19.3944
R15453 gnd.n3913 gnd.n3911 19.3944
R15454 gnd.n3911 gnd.n3910 19.3944
R15455 gnd.n3910 gnd.n3908 19.3944
R15456 gnd.n3908 gnd.n3907 19.3944
R15457 gnd.n3907 gnd.n3905 19.3944
R15458 gnd.n3905 gnd.n3904 19.3944
R15459 gnd.n3904 gnd.n3902 19.3944
R15460 gnd.n3902 gnd.n3901 19.3944
R15461 gnd.n3901 gnd.n3898 19.3944
R15462 gnd.n3898 gnd.n2003 19.3944
R15463 gnd.n4436 gnd.n2003 19.3944
R15464 gnd.n4436 gnd.n2001 19.3944
R15465 gnd.n4441 gnd.n2001 19.3944
R15466 gnd.n4441 gnd.n1995 19.3944
R15467 gnd.n4784 gnd.n1995 19.3944
R15468 gnd.n4785 gnd.n4784 19.3944
R15469 gnd.n4786 gnd.n4785 19.3944
R15470 gnd.n4824 gnd.n1895 19.3944
R15471 gnd.n4824 gnd.n1902 19.3944
R15472 gnd.n1961 gnd.n1902 19.3944
R15473 gnd.n4817 gnd.n1961 19.3944
R15474 gnd.n4817 gnd.n4816 19.3944
R15475 gnd.n4816 gnd.n4815 19.3944
R15476 gnd.n4815 gnd.n1967 19.3944
R15477 gnd.n4810 gnd.n1967 19.3944
R15478 gnd.n4810 gnd.n4809 19.3944
R15479 gnd.n4809 gnd.n4808 19.3944
R15480 gnd.n4808 gnd.n1974 19.3944
R15481 gnd.n4803 gnd.n1974 19.3944
R15482 gnd.n4803 gnd.n4802 19.3944
R15483 gnd.n4802 gnd.n4801 19.3944
R15484 gnd.n4801 gnd.n1981 19.3944
R15485 gnd.n4796 gnd.n1981 19.3944
R15486 gnd.n4796 gnd.n4795 19.3944
R15487 gnd.n4795 gnd.n4794 19.3944
R15488 gnd.n1958 gnd.n1957 19.3944
R15489 gnd.n1957 gnd.n1956 19.3944
R15490 gnd.n1956 gnd.n1953 19.3944
R15491 gnd.n1953 gnd.n1952 19.3944
R15492 gnd.n1952 gnd.n1949 19.3944
R15493 gnd.n1949 gnd.n1948 19.3944
R15494 gnd.n1948 gnd.n1945 19.3944
R15495 gnd.n1945 gnd.n1944 19.3944
R15496 gnd.n1944 gnd.n1941 19.3944
R15497 gnd.n1941 gnd.n1940 19.3944
R15498 gnd.n1940 gnd.n1937 19.3944
R15499 gnd.n1937 gnd.n1936 19.3944
R15500 gnd.n1936 gnd.n1933 19.3944
R15501 gnd.n1933 gnd.n1932 19.3944
R15502 gnd.n1932 gnd.n1896 19.3944
R15503 gnd.n4194 gnd.n2224 19.3944
R15504 gnd.n4198 gnd.n2224 19.3944
R15505 gnd.n4198 gnd.n2211 19.3944
R15506 gnd.n4210 gnd.n2211 19.3944
R15507 gnd.n4210 gnd.n2209 19.3944
R15508 gnd.n4214 gnd.n2209 19.3944
R15509 gnd.n4214 gnd.n2194 19.3944
R15510 gnd.n4226 gnd.n2194 19.3944
R15511 gnd.n4226 gnd.n2192 19.3944
R15512 gnd.n4230 gnd.n2192 19.3944
R15513 gnd.n4230 gnd.n2179 19.3944
R15514 gnd.n4242 gnd.n2179 19.3944
R15515 gnd.n4242 gnd.n2177 19.3944
R15516 gnd.n4246 gnd.n2177 19.3944
R15517 gnd.n4246 gnd.n2162 19.3944
R15518 gnd.n4258 gnd.n2162 19.3944
R15519 gnd.n4258 gnd.n2160 19.3944
R15520 gnd.n4262 gnd.n2160 19.3944
R15521 gnd.n4262 gnd.n2147 19.3944
R15522 gnd.n4274 gnd.n2147 19.3944
R15523 gnd.n4274 gnd.n2145 19.3944
R15524 gnd.n4278 gnd.n2145 19.3944
R15525 gnd.n4278 gnd.n2130 19.3944
R15526 gnd.n4290 gnd.n2130 19.3944
R15527 gnd.n4290 gnd.n2128 19.3944
R15528 gnd.n4294 gnd.n2128 19.3944
R15529 gnd.n4294 gnd.n2115 19.3944
R15530 gnd.n4306 gnd.n2115 19.3944
R15531 gnd.n4306 gnd.n2113 19.3944
R15532 gnd.n4310 gnd.n2113 19.3944
R15533 gnd.n4310 gnd.n2097 19.3944
R15534 gnd.n4322 gnd.n2097 19.3944
R15535 gnd.n4322 gnd.n2095 19.3944
R15536 gnd.n4326 gnd.n2095 19.3944
R15537 gnd.n4326 gnd.n2082 19.3944
R15538 gnd.n4338 gnd.n2082 19.3944
R15539 gnd.n4338 gnd.n2080 19.3944
R15540 gnd.n4342 gnd.n2080 19.3944
R15541 gnd.n4342 gnd.n2065 19.3944
R15542 gnd.n4354 gnd.n2065 19.3944
R15543 gnd.n4354 gnd.n2063 19.3944
R15544 gnd.n4358 gnd.n2063 19.3944
R15545 gnd.n4358 gnd.n2050 19.3944
R15546 gnd.n4370 gnd.n2050 19.3944
R15547 gnd.n4370 gnd.n2048 19.3944
R15548 gnd.n4374 gnd.n2048 19.3944
R15549 gnd.n4374 gnd.n2033 19.3944
R15550 gnd.n4386 gnd.n2033 19.3944
R15551 gnd.n4386 gnd.n2031 19.3944
R15552 gnd.n4390 gnd.n2031 19.3944
R15553 gnd.n4390 gnd.n2017 19.3944
R15554 gnd.n4415 gnd.n2017 19.3944
R15555 gnd.n4415 gnd.n2015 19.3944
R15556 gnd.n4422 gnd.n2015 19.3944
R15557 gnd.n4422 gnd.n4421 19.3944
R15558 gnd.n4421 gnd.n1062 19.3944
R15559 gnd.n6076 gnd.n1062 19.3944
R15560 gnd.n6076 gnd.n6075 19.3944
R15561 gnd.n6075 gnd.n6074 19.3944
R15562 gnd.n6074 gnd.n1066 19.3944
R15563 gnd.n6064 gnd.n1066 19.3944
R15564 gnd.n6064 gnd.n6063 19.3944
R15565 gnd.n6063 gnd.n6062 19.3944
R15566 gnd.n6062 gnd.n1089 19.3944
R15567 gnd.n3751 gnd.n3748 19.3944
R15568 gnd.n3751 gnd.n3747 19.3944
R15569 gnd.n3755 gnd.n3747 19.3944
R15570 gnd.n3755 gnd.n3745 19.3944
R15571 gnd.n3761 gnd.n3745 19.3944
R15572 gnd.n3761 gnd.n3743 19.3944
R15573 gnd.n3765 gnd.n3743 19.3944
R15574 gnd.n3765 gnd.n3741 19.3944
R15575 gnd.n3771 gnd.n3741 19.3944
R15576 gnd.n3771 gnd.n3739 19.3944
R15577 gnd.n3775 gnd.n3739 19.3944
R15578 gnd.n3775 gnd.n3737 19.3944
R15579 gnd.n3781 gnd.n3737 19.3944
R15580 gnd.n3781 gnd.n3735 19.3944
R15581 gnd.n3785 gnd.n3735 19.3944
R15582 gnd.n3785 gnd.n3730 19.3944
R15583 gnd.n3791 gnd.n3730 19.3944
R15584 gnd.n3795 gnd.n3728 19.3944
R15585 gnd.n3795 gnd.n3726 19.3944
R15586 gnd.n3801 gnd.n3726 19.3944
R15587 gnd.n3801 gnd.n3724 19.3944
R15588 gnd.n3805 gnd.n3724 19.3944
R15589 gnd.n3805 gnd.n3722 19.3944
R15590 gnd.n3811 gnd.n3722 19.3944
R15591 gnd.n3811 gnd.n3720 19.3944
R15592 gnd.n3815 gnd.n3720 19.3944
R15593 gnd.n3815 gnd.n3718 19.3944
R15594 gnd.n3821 gnd.n3718 19.3944
R15595 gnd.n3821 gnd.n3716 19.3944
R15596 gnd.n3825 gnd.n3716 19.3944
R15597 gnd.n3825 gnd.n3714 19.3944
R15598 gnd.n3831 gnd.n3714 19.3944
R15599 gnd.n3831 gnd.n3712 19.3944
R15600 gnd.n3836 gnd.n3712 19.3944
R15601 gnd.n3836 gnd.n3710 19.3944
R15602 gnd.n4187 gnd.n4186 19.3944
R15603 gnd.n4186 gnd.n3988 19.3944
R15604 gnd.n4180 gnd.n3988 19.3944
R15605 gnd.n4180 gnd.n4179 19.3944
R15606 gnd.n4179 gnd.n4178 19.3944
R15607 gnd.n4178 gnd.n3994 19.3944
R15608 gnd.n4172 gnd.n3994 19.3944
R15609 gnd.n4172 gnd.n4171 19.3944
R15610 gnd.n4171 gnd.n4170 19.3944
R15611 gnd.n4170 gnd.n4000 19.3944
R15612 gnd.n4164 gnd.n4000 19.3944
R15613 gnd.n4164 gnd.n4163 19.3944
R15614 gnd.n4163 gnd.n4162 19.3944
R15615 gnd.n4162 gnd.n4006 19.3944
R15616 gnd.n4156 gnd.n4006 19.3944
R15617 gnd.n4156 gnd.n4155 19.3944
R15618 gnd.n4146 gnd.n4145 19.3944
R15619 gnd.n4145 gnd.n4143 19.3944
R15620 gnd.n4143 gnd.n4142 19.3944
R15621 gnd.n4142 gnd.n4140 19.3944
R15622 gnd.n4140 gnd.n4139 19.3944
R15623 gnd.n4139 gnd.n4137 19.3944
R15624 gnd.n4137 gnd.n4136 19.3944
R15625 gnd.n4136 gnd.n4134 19.3944
R15626 gnd.n4134 gnd.n4133 19.3944
R15627 gnd.n4133 gnd.n4131 19.3944
R15628 gnd.n4131 gnd.n4130 19.3944
R15629 gnd.n4130 gnd.n4128 19.3944
R15630 gnd.n4128 gnd.n4127 19.3944
R15631 gnd.n4127 gnd.n4125 19.3944
R15632 gnd.n4125 gnd.n4124 19.3944
R15633 gnd.n4124 gnd.n4122 19.3944
R15634 gnd.n4122 gnd.n4121 19.3944
R15635 gnd.n4121 gnd.n4119 19.3944
R15636 gnd.n4119 gnd.n4118 19.3944
R15637 gnd.n4118 gnd.n4116 19.3944
R15638 gnd.n4116 gnd.n4115 19.3944
R15639 gnd.n4115 gnd.n4113 19.3944
R15640 gnd.n4113 gnd.n4112 19.3944
R15641 gnd.n4112 gnd.n4110 19.3944
R15642 gnd.n4110 gnd.n4109 19.3944
R15643 gnd.n4109 gnd.n4107 19.3944
R15644 gnd.n4107 gnd.n4106 19.3944
R15645 gnd.n4106 gnd.n4104 19.3944
R15646 gnd.n4104 gnd.n4103 19.3944
R15647 gnd.n4103 gnd.n4101 19.3944
R15648 gnd.n4101 gnd.n4100 19.3944
R15649 gnd.n4100 gnd.n4098 19.3944
R15650 gnd.n4098 gnd.n4045 19.3944
R15651 gnd.n4094 gnd.n4045 19.3944
R15652 gnd.n4094 gnd.n4093 19.3944
R15653 gnd.n4093 gnd.n4092 19.3944
R15654 gnd.n4092 gnd.n4049 19.3944
R15655 gnd.n4088 gnd.n4049 19.3944
R15656 gnd.n4088 gnd.n4087 19.3944
R15657 gnd.n4087 gnd.n4086 19.3944
R15658 gnd.n4086 gnd.n4053 19.3944
R15659 gnd.n4082 gnd.n4053 19.3944
R15660 gnd.n4082 gnd.n4081 19.3944
R15661 gnd.n4081 gnd.n4080 19.3944
R15662 gnd.n4080 gnd.n4057 19.3944
R15663 gnd.n4076 gnd.n4057 19.3944
R15664 gnd.n4076 gnd.n4075 19.3944
R15665 gnd.n4075 gnd.n4074 19.3944
R15666 gnd.n4074 gnd.n4061 19.3944
R15667 gnd.n4070 gnd.n4061 19.3944
R15668 gnd.n4070 gnd.n4069 19.3944
R15669 gnd.n4069 gnd.n4068 19.3944
R15670 gnd.n4068 gnd.n4064 19.3944
R15671 gnd.n4064 gnd.n2009 19.3944
R15672 gnd.n2009 gnd.n2007 19.3944
R15673 gnd.n4428 gnd.n2007 19.3944
R15674 gnd.n4428 gnd.n2005 19.3944
R15675 gnd.n4432 gnd.n2005 19.3944
R15676 gnd.n4432 gnd.n2000 19.3944
R15677 gnd.n4445 gnd.n2000 19.3944
R15678 gnd.n4445 gnd.n1997 19.3944
R15679 gnd.n4780 gnd.n1997 19.3944
R15680 gnd.n4780 gnd.n1998 19.3944
R15681 gnd.n4776 gnd.n1998 19.3944
R15682 gnd.n4190 gnd.n2219 19.3944
R15683 gnd.n4202 gnd.n2219 19.3944
R15684 gnd.n4202 gnd.n2217 19.3944
R15685 gnd.n4206 gnd.n2217 19.3944
R15686 gnd.n4206 gnd.n2203 19.3944
R15687 gnd.n4218 gnd.n2203 19.3944
R15688 gnd.n4218 gnd.n2201 19.3944
R15689 gnd.n4222 gnd.n2201 19.3944
R15690 gnd.n4222 gnd.n2187 19.3944
R15691 gnd.n4234 gnd.n2187 19.3944
R15692 gnd.n4234 gnd.n2185 19.3944
R15693 gnd.n4238 gnd.n2185 19.3944
R15694 gnd.n4238 gnd.n2171 19.3944
R15695 gnd.n4250 gnd.n2171 19.3944
R15696 gnd.n4250 gnd.n2169 19.3944
R15697 gnd.n4254 gnd.n2169 19.3944
R15698 gnd.n4254 gnd.n2155 19.3944
R15699 gnd.n4266 gnd.n2155 19.3944
R15700 gnd.n4266 gnd.n2153 19.3944
R15701 gnd.n4270 gnd.n2153 19.3944
R15702 gnd.n4270 gnd.n2139 19.3944
R15703 gnd.n4282 gnd.n2139 19.3944
R15704 gnd.n4282 gnd.n2137 19.3944
R15705 gnd.n4286 gnd.n2137 19.3944
R15706 gnd.n4286 gnd.n2123 19.3944
R15707 gnd.n4298 gnd.n2123 19.3944
R15708 gnd.n4298 gnd.n2121 19.3944
R15709 gnd.n4302 gnd.n2121 19.3944
R15710 gnd.n4302 gnd.n2107 19.3944
R15711 gnd.n4314 gnd.n2107 19.3944
R15712 gnd.n4314 gnd.n2104 19.3944
R15713 gnd.n4318 gnd.n2104 19.3944
R15714 gnd.n4318 gnd.n2089 19.3944
R15715 gnd.n4330 gnd.n2089 19.3944
R15716 gnd.n4330 gnd.n2087 19.3944
R15717 gnd.n4334 gnd.n2087 19.3944
R15718 gnd.n4334 gnd.n2074 19.3944
R15719 gnd.n4346 gnd.n2074 19.3944
R15720 gnd.n4346 gnd.n2072 19.3944
R15721 gnd.n4350 gnd.n2072 19.3944
R15722 gnd.n4350 gnd.n2057 19.3944
R15723 gnd.n4362 gnd.n2057 19.3944
R15724 gnd.n4362 gnd.n2055 19.3944
R15725 gnd.n4366 gnd.n2055 19.3944
R15726 gnd.n4366 gnd.n2042 19.3944
R15727 gnd.n4378 gnd.n2042 19.3944
R15728 gnd.n4378 gnd.n2040 19.3944
R15729 gnd.n4382 gnd.n2040 19.3944
R15730 gnd.n4382 gnd.n2025 19.3944
R15731 gnd.n4394 gnd.n2025 19.3944
R15732 gnd.n4394 gnd.n2023 19.3944
R15733 gnd.n4411 gnd.n2023 19.3944
R15734 gnd.n4411 gnd.n4410 19.3944
R15735 gnd.n4410 gnd.n4409 19.3944
R15736 gnd.n4409 gnd.n4408 19.3944
R15737 gnd.n4408 gnd.n4405 19.3944
R15738 gnd.n4405 gnd.n4404 19.3944
R15739 gnd.n4404 gnd.n1074 19.3944
R15740 gnd.n6070 gnd.n1074 19.3944
R15741 gnd.n6070 gnd.n6069 19.3944
R15742 gnd.n6069 gnd.n6068 19.3944
R15743 gnd.n6068 gnd.n1078 19.3944
R15744 gnd.n6058 gnd.n1078 19.3944
R15745 gnd.n6058 gnd.n6057 19.3944
R15746 gnd.n6052 gnd.n6051 19.3944
R15747 gnd.n6051 gnd.n6050 19.3944
R15748 gnd.n6050 gnd.n1104 19.3944
R15749 gnd.n6046 gnd.n1104 19.3944
R15750 gnd.n6046 gnd.n6045 19.3944
R15751 gnd.n6045 gnd.n6044 19.3944
R15752 gnd.n6044 gnd.n1109 19.3944
R15753 gnd.n6040 gnd.n1109 19.3944
R15754 gnd.n6040 gnd.n6039 19.3944
R15755 gnd.n6039 gnd.n6038 19.3944
R15756 gnd.n6038 gnd.n1114 19.3944
R15757 gnd.n6034 gnd.n1114 19.3944
R15758 gnd.n6034 gnd.n6033 19.3944
R15759 gnd.n6033 gnd.n6032 19.3944
R15760 gnd.n6032 gnd.n1119 19.3944
R15761 gnd.n6028 gnd.n1119 19.3944
R15762 gnd.n6028 gnd.n6027 19.3944
R15763 gnd.n6027 gnd.n6026 19.3944
R15764 gnd.n6026 gnd.n1124 19.3944
R15765 gnd.n6022 gnd.n1124 19.3944
R15766 gnd.n6022 gnd.n6021 19.3944
R15767 gnd.n6021 gnd.n6020 19.3944
R15768 gnd.n6020 gnd.n1129 19.3944
R15769 gnd.n6016 gnd.n1129 19.3944
R15770 gnd.n6016 gnd.n6015 19.3944
R15771 gnd.n6015 gnd.n6014 19.3944
R15772 gnd.n6014 gnd.n1134 19.3944
R15773 gnd.n6010 gnd.n1134 19.3944
R15774 gnd.n6010 gnd.n6009 19.3944
R15775 gnd.n6009 gnd.n6008 19.3944
R15776 gnd.n6008 gnd.n1139 19.3944
R15777 gnd.n6004 gnd.n1139 19.3944
R15778 gnd.n6004 gnd.n6003 19.3944
R15779 gnd.n6003 gnd.n6002 19.3944
R15780 gnd.n6002 gnd.n1144 19.3944
R15781 gnd.n5998 gnd.n1144 19.3944
R15782 gnd.n5998 gnd.n5997 19.3944
R15783 gnd.n5997 gnd.n5996 19.3944
R15784 gnd.n5996 gnd.n1149 19.3944
R15785 gnd.n5992 gnd.n1149 19.3944
R15786 gnd.n5992 gnd.n5991 19.3944
R15787 gnd.n5991 gnd.n5990 19.3944
R15788 gnd.n5990 gnd.n1154 19.3944
R15789 gnd.n5986 gnd.n1154 19.3944
R15790 gnd.n5986 gnd.n5985 19.3944
R15791 gnd.n5985 gnd.n5984 19.3944
R15792 gnd.n5984 gnd.n1159 19.3944
R15793 gnd.n5980 gnd.n1159 19.3944
R15794 gnd.n5980 gnd.n5979 19.3944
R15795 gnd.n5979 gnd.n5978 19.3944
R15796 gnd.n5978 gnd.n1164 19.3944
R15797 gnd.n5974 gnd.n1164 19.3944
R15798 gnd.n5974 gnd.n5973 19.3944
R15799 gnd.n5973 gnd.n5972 19.3944
R15800 gnd.n5972 gnd.n1169 19.3944
R15801 gnd.n5968 gnd.n1169 19.3944
R15802 gnd.n5968 gnd.n5967 19.3944
R15803 gnd.n5967 gnd.n5966 19.3944
R15804 gnd.n5966 gnd.n1174 19.3944
R15805 gnd.n5962 gnd.n1174 19.3944
R15806 gnd.n5962 gnd.n5961 19.3944
R15807 gnd.n5961 gnd.n5960 19.3944
R15808 gnd.n5960 gnd.n1179 19.3944
R15809 gnd.n5956 gnd.n1179 19.3944
R15810 gnd.n5956 gnd.n5955 19.3944
R15811 gnd.n5955 gnd.n5954 19.3944
R15812 gnd.n5954 gnd.n1184 19.3944
R15813 gnd.n5950 gnd.n1184 19.3944
R15814 gnd.n5950 gnd.n5949 19.3944
R15815 gnd.n5949 gnd.n5948 19.3944
R15816 gnd.n5948 gnd.n1189 19.3944
R15817 gnd.n5944 gnd.n1189 19.3944
R15818 gnd.n5944 gnd.n5943 19.3944
R15819 gnd.n5943 gnd.n5942 19.3944
R15820 gnd.n5942 gnd.n1194 19.3944
R15821 gnd.n5938 gnd.n1194 19.3944
R15822 gnd.n5938 gnd.n5937 19.3944
R15823 gnd.n5937 gnd.n5936 19.3944
R15824 gnd.n5936 gnd.n1199 19.3944
R15825 gnd.n5932 gnd.n1199 19.3944
R15826 gnd.n5932 gnd.n5931 19.3944
R15827 gnd.n5931 gnd.n5930 19.3944
R15828 gnd.n5930 gnd.n1204 19.3944
R15829 gnd.n5926 gnd.n1204 19.3944
R15830 gnd.n5926 gnd.n5925 19.3944
R15831 gnd.n5925 gnd.n5924 19.3944
R15832 gnd.n5924 gnd.n1209 19.3944
R15833 gnd.n5920 gnd.n1209 19.3944
R15834 gnd.n5920 gnd.n5919 19.3944
R15835 gnd.n5919 gnd.n5918 19.3944
R15836 gnd.n5918 gnd.n1214 19.3944
R15837 gnd.n5914 gnd.n1214 19.3944
R15838 gnd.n5914 gnd.n5913 19.3944
R15839 gnd.n5913 gnd.n5912 19.3944
R15840 gnd.n5912 gnd.n1219 19.3944
R15841 gnd.n5908 gnd.n1219 19.3944
R15842 gnd.n5908 gnd.n5907 19.3944
R15843 gnd.n5907 gnd.n5906 19.3944
R15844 gnd.n5906 gnd.n1224 19.3944
R15845 gnd.n5902 gnd.n1224 19.3944
R15846 gnd.n5902 gnd.n5901 19.3944
R15847 gnd.n1297 gnd.n1294 19.3944
R15848 gnd.n1297 gnd.n1266 19.3944
R15849 gnd.n5888 gnd.n1266 19.3944
R15850 gnd.n7148 gnd.n7147 19.3944
R15851 gnd.n7147 gnd.n461 19.3944
R15852 gnd.n7140 gnd.n461 19.3944
R15853 gnd.n7140 gnd.n7139 19.3944
R15854 gnd.n7139 gnd.n469 19.3944
R15855 gnd.n7132 gnd.n469 19.3944
R15856 gnd.n7132 gnd.n7131 19.3944
R15857 gnd.n7131 gnd.n477 19.3944
R15858 gnd.n7124 gnd.n477 19.3944
R15859 gnd.n7124 gnd.n7123 19.3944
R15860 gnd.n7123 gnd.n485 19.3944
R15861 gnd.n7116 gnd.n485 19.3944
R15862 gnd.n7116 gnd.n7115 19.3944
R15863 gnd.n7115 gnd.n493 19.3944
R15864 gnd.n7108 gnd.n493 19.3944
R15865 gnd.n7108 gnd.n7107 19.3944
R15866 gnd.n7107 gnd.n503 19.3944
R15867 gnd.n1279 gnd.n503 19.3944
R15868 gnd.n1279 gnd.n1274 19.3944
R15869 gnd.n1284 gnd.n1274 19.3944
R15870 gnd.n1285 gnd.n1284 19.3944
R15871 gnd.n1288 gnd.n1285 19.3944
R15872 gnd.n1288 gnd.n1270 19.3944
R15873 gnd.n1292 gnd.n1270 19.3944
R15874 gnd.n7072 gnd.n7071 18.4247
R15875 gnd.n4828 gnd.n1896 18.4247
R15876 gnd.n7430 gnd.n124 18.2308
R15877 gnd.n7111 gnd.n499 18.2308
R15878 gnd.n4725 gnd.n4556 18.2308
R15879 gnd.n4155 gnd.n4012 18.2308
R15880 gnd.n2858 gnd.n2752 18.2305
R15881 gnd.n2858 gnd.n2857 18.2305
R15882 gnd.n2866 gnd.n2741 18.2305
R15883 gnd.n2874 gnd.n2741 18.2305
R15884 gnd.n2874 gnd.n2735 18.2305
R15885 gnd.n2882 gnd.n2735 18.2305
R15886 gnd.n2882 gnd.n2728 18.2305
R15887 gnd.n2920 gnd.n2728 18.2305
R15888 gnd.n2930 gnd.n2661 18.2305
R15889 gnd.n4192 gnd.n3985 18.2305
R15890 gnd.n4200 gnd.n2213 18.2305
R15891 gnd.n4208 gnd.n2213 18.2305
R15892 gnd.n4208 gnd.n2205 18.2305
R15893 gnd.n4216 gnd.n2205 18.2305
R15894 gnd.n4224 gnd.n2196 18.2305
R15895 gnd.n4224 gnd.n2199 18.2305
R15896 gnd.n4232 gnd.n2181 18.2305
R15897 gnd.n4240 gnd.n2181 18.2305
R15898 gnd.n4248 gnd.n2173 18.2305
R15899 gnd.n4256 gnd.n2164 18.2305
R15900 gnd.n4256 gnd.n2167 18.2305
R15901 gnd.n4264 gnd.n2149 18.2305
R15902 gnd.n4272 gnd.n2149 18.2305
R15903 gnd.n4280 gnd.n2141 18.2305
R15904 gnd.n4288 gnd.n2132 18.2305
R15905 gnd.n4288 gnd.n2135 18.2305
R15906 gnd.n4296 gnd.n2117 18.2305
R15907 gnd.n4304 gnd.n2117 18.2305
R15908 gnd.n4312 gnd.n2109 18.2305
R15909 gnd.n4320 gnd.n2099 18.2305
R15910 gnd.n4320 gnd.n2102 18.2305
R15911 gnd.n4328 gnd.n2093 18.2305
R15912 gnd.n4336 gnd.n2076 18.2305
R15913 gnd.n4344 gnd.n2076 18.2305
R15914 gnd.n4352 gnd.n2067 18.2305
R15915 gnd.n4352 gnd.n2070 18.2305
R15916 gnd.n4360 gnd.n2061 18.2305
R15917 gnd.n4368 gnd.n2044 18.2305
R15918 gnd.n4376 gnd.n2044 18.2305
R15919 gnd.n4384 gnd.n2035 18.2305
R15920 gnd.n4384 gnd.n2038 18.2305
R15921 gnd.n4392 gnd.n2029 18.2305
R15922 gnd.n4413 gnd.n2010 18.2305
R15923 gnd.n4424 gnd.n2010 18.2305
R15924 gnd.t26 gnd.n2109 18.0482
R15925 gnd.n2093 gnd.t69 18.0482
R15926 gnd.t85 gnd.n2141 17.6836
R15927 gnd.n2061 gnd.t16 17.6836
R15928 gnd.t65 gnd.n2173 17.319
R15929 gnd.n2029 gnd.t36 17.319
R15930 gnd.n3985 gnd.t169 16.2252
R15931 gnd.n4621 gnd.n4620 15.9333
R15932 gnd.n4624 gnd.n4621 15.9333
R15933 gnd.n4624 gnd.n4623 15.9333
R15934 gnd.n4623 gnd.n4622 15.9333
R15935 gnd.n4632 gnd.n4610 15.9333
R15936 gnd.n4635 gnd.n4632 15.9333
R15937 gnd.n4636 gnd.n4635 15.9333
R15938 gnd.n4637 gnd.n4636 15.9333
R15939 gnd.n4640 gnd.n4637 15.9333
R15940 gnd.n4640 gnd.n4639 15.9333
R15941 gnd.n4639 gnd.n4638 15.9333
R15942 gnd.n4638 gnd.n4604 15.9333
R15943 gnd.n4648 gnd.n4604 15.9333
R15944 gnd.n4652 gnd.n4651 15.9333
R15945 gnd.n4653 gnd.n4652 15.9333
R15946 gnd.n4656 gnd.n4653 15.9333
R15947 gnd.n4656 gnd.n4655 15.9333
R15948 gnd.n4655 gnd.n4654 15.9333
R15949 gnd.n4654 gnd.n4598 15.9333
R15950 gnd.n4664 gnd.n4598 15.9333
R15951 gnd.n4666 gnd.n4664 15.9333
R15952 gnd.n4906 gnd.n1772 15.9333
R15953 gnd.n4914 gnd.n1758 15.9333
R15954 gnd.n4965 gnd.n1752 15.9333
R15955 gnd.n4974 gnd.n4973 15.9333
R15956 gnd.n5004 gnd.n5003 15.9333
R15957 gnd.n4944 gnd.n1706 15.9333
R15958 gnd.n5067 gnd.n5066 15.9333
R15959 gnd.n5075 gnd.n1694 15.9333
R15960 gnd.n5100 gnd.n1666 15.9333
R15961 gnd.n5126 gnd.n1661 15.9333
R15962 gnd.n5134 gnd.n1654 15.9333
R15963 gnd.n5171 gnd.n1643 15.9333
R15964 gnd.n5183 gnd.n5181 15.9333
R15965 gnd.n5148 gnd.n1621 15.9333
R15966 gnd.n5244 gnd.n5243 15.9333
R15967 gnd.n5252 gnd.n1609 15.9333
R15968 gnd.n5270 gnd.n5269 15.9333
R15969 gnd.n5278 gnd.n1580 15.9333
R15970 gnd.n5303 gnd.n1572 15.9333
R15971 gnd.n5303 gnd.n1575 15.9333
R15972 gnd.n5311 gnd.n1566 15.9333
R15973 gnd.n5349 gnd.n1555 15.9333
R15974 gnd.n5360 gnd.n5359 15.9333
R15975 gnd.n5326 gnd.n1534 15.9333
R15976 gnd.n5406 gnd.n5405 15.9333
R15977 gnd.n5414 gnd.n1522 15.9333
R15978 gnd.n5431 gnd.n5430 15.9333
R15979 gnd.n5439 gnd.n1492 15.9333
R15980 gnd.n5492 gnd.n1486 15.9333
R15981 gnd.n5501 gnd.n5500 15.9333
R15982 gnd.n5532 gnd.n5531 15.9333
R15983 gnd.n5471 gnd.n1442 15.9333
R15984 gnd.n5587 gnd.n5586 15.9333
R15985 gnd.n5595 gnd.n1430 15.9333
R15986 gnd.n5819 gnd.n5818 15.9333
R15987 gnd.n5818 gnd.n5817 15.9333
R15988 gnd.n5828 gnd.n5827 15.9333
R15989 gnd.n5827 gnd.n1328 15.9333
R15990 gnd.n5837 gnd.n1328 15.9333
R15991 gnd.n5839 gnd.n5837 15.9333
R15992 gnd.n5839 gnd.n5838 15.9333
R15993 gnd.n5838 gnd.n1321 15.9333
R15994 gnd.n5849 gnd.n1321 15.9333
R15995 gnd.n5849 gnd.n5848 15.9333
R15996 gnd.n5847 gnd.n1315 15.9333
R15997 gnd.n5857 gnd.n1315 15.9333
R15998 gnd.n5859 gnd.n5857 15.9333
R15999 gnd.n5859 gnd.n5858 15.9333
R16000 gnd.n5858 gnd.n1308 15.9333
R16001 gnd.n5872 gnd.n1308 15.9333
R16002 gnd.n5872 gnd.n5871 15.9333
R16003 gnd.n5871 gnd.n5870 15.9333
R16004 gnd.n5870 gnd.n5869 15.9333
R16005 gnd.n5882 gnd.n5881 15.9333
R16006 gnd.n5882 gnd.n1227 15.9333
R16007 gnd.n5899 gnd.n1227 15.9333
R16008 gnd.n5899 gnd.n5898 15.9333
R16009 gnd.n3553 gnd.n3551 15.6674
R16010 gnd.n3521 gnd.n3519 15.6674
R16011 gnd.n3489 gnd.n3487 15.6674
R16012 gnd.n3458 gnd.n3456 15.6674
R16013 gnd.n3426 gnd.n3424 15.6674
R16014 gnd.n3394 gnd.n3392 15.6674
R16015 gnd.n3362 gnd.n3360 15.6674
R16016 gnd.n3331 gnd.n3329 15.6674
R16017 gnd.n5557 gnd.t118 15.296
R16018 gnd.n5660 gnd.n5659 15.0827
R16019 gnd.n1819 gnd.n1814 15.0481
R16020 gnd.n5670 gnd.n5669 15.0481
R16021 gnd.n2004 gnd.t34 14.9773
R16022 gnd.n4983 gnd.t236 14.9773
R16023 gnd.t226 gnd.n5611 14.9773
R16024 gnd.t224 gnd.n428 14.9773
R16025 gnd.n1745 gnd.n1734 14.6587
R16026 gnd.n4936 gnd.t63 14.6587
R16027 gnd.n5103 gnd.n5101 14.6587
R16028 gnd.n1479 gnd.n1478 14.6587
R16029 gnd.t43 gnd.n1452 14.6587
R16030 gnd.n5622 gnd.n5621 14.6587
R16031 gnd.n1389 gnd.n1380 14.6587
R16032 gnd.n6246 gnd.n969 14.4022
R16033 gnd.n2942 gnd.n2662 14.2199
R16034 gnd.n2952 gnd.n2645 14.2199
R16035 gnd.n2648 gnd.n2636 14.2199
R16036 gnd.n2973 gnd.n2637 14.2199
R16037 gnd.n2983 gnd.n2617 14.2199
R16038 gnd.n2993 gnd.n2992 14.2199
R16039 gnd.n2603 gnd.n2601 14.2199
R16040 gnd.n3024 gnd.n3023 14.2199
R16041 gnd.n3039 gnd.n2586 14.2199
R16042 gnd.n3093 gnd.n2525 14.2199
R16043 gnd.n3049 gnd.n2526 14.2199
R16044 gnd.n3086 gnd.n2537 14.2199
R16045 gnd.n2575 gnd.n2574 14.2199
R16046 gnd.n3080 gnd.n3079 14.2199
R16047 gnd.n2561 gnd.n2548 14.2199
R16048 gnd.n3119 gnd.n3118 14.2199
R16049 gnd.n3129 gnd.n2445 14.2199
R16050 gnd.n3141 gnd.n2437 14.2199
R16051 gnd.n3140 gnd.n2425 14.2199
R16052 gnd.n3159 gnd.n3158 14.2199
R16053 gnd.n3169 gnd.n2418 14.2199
R16054 gnd.n3180 gnd.n2406 14.2199
R16055 gnd.n3204 gnd.n3203 14.2199
R16056 gnd.n3215 gnd.n2389 14.2199
R16057 gnd.n3214 gnd.n2391 14.2199
R16058 gnd.n3226 gnd.n2382 14.2199
R16059 gnd.n3244 gnd.n3243 14.2199
R16060 gnd.n2373 gnd.n2362 14.2199
R16061 gnd.n3265 gnd.n2350 14.2199
R16062 gnd.n3293 gnd.n3292 14.2199
R16063 gnd.n3304 gnd.n2335 14.2199
R16064 gnd.n3315 gnd.n2328 14.2199
R16065 gnd.n3314 gnd.n2316 14.2199
R16066 gnd.n3587 gnd.n3586 14.2199
R16067 gnd.n3609 gnd.n2301 14.2199
R16068 gnd.n5005 gnd.n1720 14.0214
R16069 gnd.n1693 gnd.t57 14.0214
R16070 gnd.n5184 gnd.n1635 14.0214
R16071 gnd.n1608 gnd.n1607 14.0214
R16072 gnd.n5361 gnd.n1547 14.0214
R16073 gnd.n1521 gnd.n1520 14.0214
R16074 gnd.n5533 gnd.t59 14.0214
R16075 gnd.n1428 gnd.n1421 14.0214
R16076 gnd.t94 gnd.n5650 14.0214
R16077 gnd.n7034 gnd.n583 13.5763
R16078 gnd.n7482 gnd.n7481 13.5763
R16079 gnd.n2723 gnd.n2722 13.5763
R16080 gnd.n3667 gnd.n2265 13.5763
R16081 gnd.n4794 gnd.n1990 13.5763
R16082 gnd.n3710 gnd.n3709 13.5763
R16083 gnd.n4916 gnd.t97 13.384
R16084 gnd.n4992 gnd.n1729 13.384
R16085 gnd.n1685 gnd.n1680 13.384
R16086 gnd.n5026 gnd.t62 13.384
R16087 gnd.n5170 gnd.n1645 13.384
R16088 gnd.n1600 gnd.n1595 13.384
R16089 gnd.n5348 gnd.n1558 13.384
R16090 gnd.n1513 gnd.n1507 13.384
R16091 gnd.n5448 gnd.t56 13.384
R16092 gnd.n5520 gnd.n1464 13.384
R16093 gnd.n5548 gnd.n1416 13.384
R16094 gnd.n2963 gnd.t2 13.3084
R16095 gnd.n4216 gnd.t250 13.3084
R16096 gnd.n1830 gnd.n1811 13.1884
R16097 gnd.n1825 gnd.n1824 13.1884
R16098 gnd.n1824 gnd.n1823 13.1884
R16099 gnd.n5663 gnd.n5658 13.1884
R16100 gnd.n5664 gnd.n5663 13.1884
R16101 gnd.n1826 gnd.n1813 13.146
R16102 gnd.n1822 gnd.n1813 13.146
R16103 gnd.n5662 gnd.n5661 13.146
R16104 gnd.n5662 gnd.n5657 13.146
R16105 gnd.n2664 gnd.t194 12.9438
R16106 gnd.n4248 gnd.t261 12.9438
R16107 gnd.n4392 gnd.t71 12.9438
R16108 gnd.n3554 gnd.n3550 12.8005
R16109 gnd.n3522 gnd.n3518 12.8005
R16110 gnd.n3490 gnd.n3486 12.8005
R16111 gnd.n3459 gnd.n3455 12.8005
R16112 gnd.n3427 gnd.n3423 12.8005
R16113 gnd.n3395 gnd.n3391 12.8005
R16114 gnd.n3363 gnd.n3359 12.8005
R16115 gnd.n3332 gnd.n3328 12.8005
R16116 gnd.n4904 gnd.n1764 12.7467
R16117 gnd.t122 gnd.t125 12.7467
R16118 gnd.n4985 gnd.n4984 12.7467
R16119 gnd.n4945 gnd.t46 12.7467
R16120 gnd.n5090 gnd.n1672 12.7467
R16121 gnd.n5163 gnd.n5162 12.7467
R16122 gnd.n5267 gnd.n1587 12.7467
R16123 gnd.n5341 gnd.n5340 12.7467
R16124 gnd.n5429 gnd.n1499 12.7467
R16125 gnd.n5513 gnd.n5512 12.7467
R16126 gnd.n5585 gnd.t41 12.7467
R16127 gnd.n5610 gnd.n1408 12.7467
R16128 gnd.n5554 gnd.t150 12.7467
R16129 gnd.n4280 gnd.t67 12.5792
R16130 gnd.n4360 gnd.t18 12.5792
R16131 gnd.n4651 gnd.t280 12.4281
R16132 gnd.n5848 gnd.t282 12.4281
R16133 gnd.n6955 gnd.t212 12.4281
R16134 gnd.t8 gnd.n229 12.4281
R16135 gnd.n7030 gnd.n583 12.4126
R16136 gnd.n7481 gnd.n200 12.4126
R16137 gnd.n2722 gnd.n2717 12.4126
R16138 gnd.n3670 gnd.n3667 12.4126
R16139 gnd.n4789 gnd.n1990 12.4126
R16140 gnd.n3843 gnd.n3709 12.4126
R16141 gnd.t228 gnd.n2669 12.2146
R16142 gnd.n4312 gnd.t4 12.2146
R16143 gnd.n4328 gnd.t10 12.2146
R16144 gnd.n4893 gnd.n1831 12.1761
R16145 gnd.n5743 gnd.n5742 12.1761
R16146 gnd.n5013 gnd.n1714 12.1094
R16147 gnd.n5076 gnd.n1691 12.1094
R16148 gnd.n5191 gnd.n1629 12.1094
R16149 gnd.n5253 gnd.n1605 12.1094
R16150 gnd.n5368 gnd.n1542 12.1094
R16151 gnd.n5415 gnd.n1518 12.1094
R16152 gnd.n5540 gnd.n1450 12.1094
R16153 gnd.n5596 gnd.n1426 12.1094
R16154 gnd.n3558 gnd.n3557 12.0247
R16155 gnd.n3526 gnd.n3525 12.0247
R16156 gnd.n3494 gnd.n3493 12.0247
R16157 gnd.n3463 gnd.n3462 12.0247
R16158 gnd.n3431 gnd.n3430 12.0247
R16159 gnd.n3399 gnd.n3398 12.0247
R16160 gnd.n3367 gnd.n3366 12.0247
R16161 gnd.n3336 gnd.n3335 12.0247
R16162 gnd.t265 gnd.n2363 11.85
R16163 gnd.n4296 gnd.t39 11.85
R16164 gnd.n4344 gnd.t292 11.85
R16165 gnd.t34 gnd.n1056 11.85
R16166 gnd.n387 gnd.t75 11.7908
R16167 gnd.t248 gnd.n259 11.7908
R16168 gnd.t267 gnd.n2398 11.4854
R16169 gnd.n4264 gnd.t221 11.4854
R16170 gnd.n4376 gnd.t204 11.4854
R16171 gnd.n4931 gnd.n1759 11.4721
R16172 gnd.n5119 gnd.n1667 11.4721
R16173 gnd.n5111 gnd.n5110 11.4721
R16174 gnd.n5296 gnd.n1581 11.4721
R16175 gnd.n5288 gnd.n5287 11.4721
R16176 gnd.n5457 gnd.n1493 11.4721
R16177 gnd.n5449 gnd.n1477 11.4721
R16178 gnd.n5631 gnd.n1403 11.4721
R16179 gnd.n5652 gnd.n1386 11.4721
R16180 gnd.n1056 gnd.n969 11.3031
R16181 gnd.n3561 gnd.n3548 11.249
R16182 gnd.n3529 gnd.n3516 11.249
R16183 gnd.n3497 gnd.n3484 11.249
R16184 gnd.n3466 gnd.n3453 11.249
R16185 gnd.n3434 gnd.n3421 11.249
R16186 gnd.n3402 gnd.n3389 11.249
R16187 gnd.n3370 gnd.n3357 11.249
R16188 gnd.n3339 gnd.n3326 11.249
R16189 gnd.n355 gnd.t28 11.1535
R16190 gnd.t207 gnd.n289 11.1535
R16191 gnd.n3130 gnd.t273 11.1208
R16192 gnd.n4232 gnd.t255 11.1208
R16193 gnd.n4424 gnd.t77 11.1208
R16194 gnd.n5059 gnd.n5058 10.8348
R16195 gnd.n5135 gnd.t50 10.8348
R16196 gnd.n5235 gnd.n5234 10.8348
R16197 gnd.n5234 gnd.n1615 10.8348
R16198 gnd.n5398 gnd.n5397 10.8348
R16199 gnd.n5397 gnd.n1528 10.8348
R16200 gnd.t52 gnd.n5440 10.8348
R16201 gnd.n5578 gnd.n1436 10.8348
R16202 gnd.n3087 gnd.t279 10.7562
R16203 gnd.n3072 gnd.t329 10.7562
R16204 gnd.n5813 gnd.n5812 10.6151
R16205 gnd.n5812 gnd.n5809 10.6151
R16206 gnd.n5807 gnd.n5804 10.6151
R16207 gnd.n5804 gnd.n5803 10.6151
R16208 gnd.n5803 gnd.n5800 10.6151
R16209 gnd.n5800 gnd.n5799 10.6151
R16210 gnd.n5799 gnd.n5796 10.6151
R16211 gnd.n5796 gnd.n5795 10.6151
R16212 gnd.n5795 gnd.n5792 10.6151
R16213 gnd.n5792 gnd.n5791 10.6151
R16214 gnd.n5791 gnd.n5788 10.6151
R16215 gnd.n5788 gnd.n5787 10.6151
R16216 gnd.n5787 gnd.n5784 10.6151
R16217 gnd.n5784 gnd.n5783 10.6151
R16218 gnd.n5783 gnd.n5780 10.6151
R16219 gnd.n5780 gnd.n5779 10.6151
R16220 gnd.n5779 gnd.n5776 10.6151
R16221 gnd.n5776 gnd.n5775 10.6151
R16222 gnd.n5775 gnd.n5772 10.6151
R16223 gnd.n5772 gnd.n5771 10.6151
R16224 gnd.n5771 gnd.n5768 10.6151
R16225 gnd.n5768 gnd.n5767 10.6151
R16226 gnd.n5767 gnd.n5764 10.6151
R16227 gnd.n5764 gnd.n5763 10.6151
R16228 gnd.n5763 gnd.n5760 10.6151
R16229 gnd.n5760 gnd.n5759 10.6151
R16230 gnd.n5759 gnd.n5756 10.6151
R16231 gnd.n5756 gnd.n5755 10.6151
R16232 gnd.n5755 gnd.n5752 10.6151
R16233 gnd.n5752 gnd.n5751 10.6151
R16234 gnd.n4902 gnd.n4901 10.6151
R16235 gnd.n4901 gnd.n1755 10.6151
R16236 gnd.n4933 gnd.n1755 10.6151
R16237 gnd.n4934 gnd.n4933 10.6151
R16238 gnd.n4963 gnd.n4934 10.6151
R16239 gnd.n4963 gnd.n4962 10.6151
R16240 gnd.n4962 gnd.n4961 10.6151
R16241 gnd.n4961 gnd.n4958 10.6151
R16242 gnd.n4958 gnd.n4957 10.6151
R16243 gnd.n4957 gnd.n4956 10.6151
R16244 gnd.n4956 gnd.n4955 10.6151
R16245 gnd.n4955 gnd.n4954 10.6151
R16246 gnd.n4954 gnd.n4951 10.6151
R16247 gnd.n4951 gnd.n4950 10.6151
R16248 gnd.n4950 gnd.n4948 10.6151
R16249 gnd.n4948 gnd.n4947 10.6151
R16250 gnd.n4947 gnd.n4943 10.6151
R16251 gnd.n4943 gnd.n4942 10.6151
R16252 gnd.n4942 gnd.n4940 10.6151
R16253 gnd.n4940 gnd.n4939 10.6151
R16254 gnd.n4939 gnd.n4935 10.6151
R16255 gnd.n4935 gnd.n1683 10.6151
R16256 gnd.n5085 gnd.n1683 10.6151
R16257 gnd.n5086 gnd.n5085 10.6151
R16258 gnd.n5088 gnd.n5086 10.6151
R16259 gnd.n5088 gnd.n5087 10.6151
R16260 gnd.n5087 gnd.n1664 10.6151
R16261 gnd.n5121 gnd.n1664 10.6151
R16262 gnd.n5122 gnd.n5121 10.6151
R16263 gnd.n5124 gnd.n5122 10.6151
R16264 gnd.n5124 gnd.n5123 10.6151
R16265 gnd.n5123 gnd.n1651 10.6151
R16266 gnd.n5137 gnd.n1651 10.6151
R16267 gnd.n5138 gnd.n5137 10.6151
R16268 gnd.n5160 gnd.n5138 10.6151
R16269 gnd.n5160 gnd.n5159 10.6151
R16270 gnd.n5159 gnd.n5158 10.6151
R16271 gnd.n5158 gnd.n5155 10.6151
R16272 gnd.n5155 gnd.n5154 10.6151
R16273 gnd.n5154 gnd.n5152 10.6151
R16274 gnd.n5152 gnd.n5151 10.6151
R16275 gnd.n5151 gnd.n5147 10.6151
R16276 gnd.n5147 gnd.n5146 10.6151
R16277 gnd.n5146 gnd.n5144 10.6151
R16278 gnd.n5144 gnd.n5143 10.6151
R16279 gnd.n5143 gnd.n5139 10.6151
R16280 gnd.n5139 gnd.n1598 10.6151
R16281 gnd.n5262 gnd.n1598 10.6151
R16282 gnd.n5263 gnd.n5262 10.6151
R16283 gnd.n5265 gnd.n5263 10.6151
R16284 gnd.n5265 gnd.n5264 10.6151
R16285 gnd.n5264 gnd.n1578 10.6151
R16286 gnd.n5298 gnd.n1578 10.6151
R16287 gnd.n5299 gnd.n5298 10.6151
R16288 gnd.n5301 gnd.n5299 10.6151
R16289 gnd.n5301 gnd.n5300 10.6151
R16290 gnd.n5300 gnd.n1564 10.6151
R16291 gnd.n5314 gnd.n1564 10.6151
R16292 gnd.n5315 gnd.n5314 10.6151
R16293 gnd.n5338 gnd.n5315 10.6151
R16294 gnd.n5338 gnd.n5337 10.6151
R16295 gnd.n5337 gnd.n5336 10.6151
R16296 gnd.n5336 gnd.n5333 10.6151
R16297 gnd.n5333 gnd.n5332 10.6151
R16298 gnd.n5332 gnd.n5330 10.6151
R16299 gnd.n5330 gnd.n5329 10.6151
R16300 gnd.n5329 gnd.n5324 10.6151
R16301 gnd.n5324 gnd.n5323 10.6151
R16302 gnd.n5323 gnd.n5321 10.6151
R16303 gnd.n5321 gnd.n5320 10.6151
R16304 gnd.n5320 gnd.n5316 10.6151
R16305 gnd.n5316 gnd.n1510 10.6151
R16306 gnd.n5424 gnd.n1510 10.6151
R16307 gnd.n5425 gnd.n5424 10.6151
R16308 gnd.n5427 gnd.n5425 10.6151
R16309 gnd.n5427 gnd.n5426 10.6151
R16310 gnd.n5426 gnd.n1490 10.6151
R16311 gnd.n5459 gnd.n1490 10.6151
R16312 gnd.n5460 gnd.n5459 10.6151
R16313 gnd.n5490 gnd.n5460 10.6151
R16314 gnd.n5490 gnd.n5489 10.6151
R16315 gnd.n5489 gnd.n5488 10.6151
R16316 gnd.n5488 gnd.n5485 10.6151
R16317 gnd.n5485 gnd.n5484 10.6151
R16318 gnd.n5484 gnd.n5483 10.6151
R16319 gnd.n5483 gnd.n5482 10.6151
R16320 gnd.n5482 gnd.n5481 10.6151
R16321 gnd.n5481 gnd.n5478 10.6151
R16322 gnd.n5478 gnd.n5477 10.6151
R16323 gnd.n5477 gnd.n5475 10.6151
R16324 gnd.n5475 gnd.n5474 10.6151
R16325 gnd.n5474 gnd.n5469 10.6151
R16326 gnd.n5469 gnd.n5468 10.6151
R16327 gnd.n5468 gnd.n5466 10.6151
R16328 gnd.n5466 gnd.n5465 10.6151
R16329 gnd.n5465 gnd.n5461 10.6151
R16330 gnd.n5461 gnd.n1419 10.6151
R16331 gnd.n5605 gnd.n1419 10.6151
R16332 gnd.n5606 gnd.n5605 10.6151
R16333 gnd.n5608 gnd.n5606 10.6151
R16334 gnd.n5608 gnd.n5607 10.6151
R16335 gnd.n5607 gnd.n1399 10.6151
R16336 gnd.n5633 gnd.n1399 10.6151
R16337 gnd.n5634 gnd.n5633 10.6151
R16338 gnd.n5638 gnd.n5634 10.6151
R16339 gnd.n5638 gnd.n5637 10.6151
R16340 gnd.n5637 gnd.n5636 10.6151
R16341 gnd.n5636 gnd.n5635 10.6151
R16342 gnd.n5635 gnd.n1378 10.6151
R16343 gnd.n1378 gnd.n1376 10.6151
R16344 gnd.n1894 gnd.n1893 10.6151
R16345 gnd.n1893 gnd.n1890 10.6151
R16346 gnd.n1888 gnd.n1885 10.6151
R16347 gnd.n1885 gnd.n1884 10.6151
R16348 gnd.n1884 gnd.n1881 10.6151
R16349 gnd.n1881 gnd.n1880 10.6151
R16350 gnd.n1880 gnd.n1877 10.6151
R16351 gnd.n1877 gnd.n1876 10.6151
R16352 gnd.n1876 gnd.n1873 10.6151
R16353 gnd.n1873 gnd.n1872 10.6151
R16354 gnd.n1872 gnd.n1869 10.6151
R16355 gnd.n1869 gnd.n1868 10.6151
R16356 gnd.n1868 gnd.n1865 10.6151
R16357 gnd.n1865 gnd.n1864 10.6151
R16358 gnd.n1864 gnd.n1861 10.6151
R16359 gnd.n1861 gnd.n1860 10.6151
R16360 gnd.n1860 gnd.n1857 10.6151
R16361 gnd.n1857 gnd.n1856 10.6151
R16362 gnd.n1856 gnd.n1853 10.6151
R16363 gnd.n1853 gnd.n1852 10.6151
R16364 gnd.n1852 gnd.n1849 10.6151
R16365 gnd.n1849 gnd.n1848 10.6151
R16366 gnd.n1848 gnd.n1845 10.6151
R16367 gnd.n1845 gnd.n1844 10.6151
R16368 gnd.n1844 gnd.n1841 10.6151
R16369 gnd.n1841 gnd.n1840 10.6151
R16370 gnd.n1840 gnd.n1837 10.6151
R16371 gnd.n1837 gnd.n1775 10.6151
R16372 gnd.n4899 gnd.n1775 10.6151
R16373 gnd.n4900 gnd.n4899 10.6151
R16374 gnd.n4893 gnd.n4892 10.6151
R16375 gnd.n4892 gnd.n4891 10.6151
R16376 gnd.n4891 gnd.n4890 10.6151
R16377 gnd.n4890 gnd.n4888 10.6151
R16378 gnd.n4888 gnd.n4885 10.6151
R16379 gnd.n4885 gnd.n4884 10.6151
R16380 gnd.n4884 gnd.n4881 10.6151
R16381 gnd.n4881 gnd.n4880 10.6151
R16382 gnd.n4880 gnd.n4877 10.6151
R16383 gnd.n4877 gnd.n4876 10.6151
R16384 gnd.n4876 gnd.n4873 10.6151
R16385 gnd.n4873 gnd.n4872 10.6151
R16386 gnd.n4872 gnd.n4869 10.6151
R16387 gnd.n4869 gnd.n4868 10.6151
R16388 gnd.n4868 gnd.n4865 10.6151
R16389 gnd.n4865 gnd.n4864 10.6151
R16390 gnd.n4864 gnd.n4861 10.6151
R16391 gnd.n4861 gnd.n4860 10.6151
R16392 gnd.n4860 gnd.n4857 10.6151
R16393 gnd.n4857 gnd.n4856 10.6151
R16394 gnd.n4856 gnd.n4853 10.6151
R16395 gnd.n4853 gnd.n4852 10.6151
R16396 gnd.n4852 gnd.n4849 10.6151
R16397 gnd.n4849 gnd.n4848 10.6151
R16398 gnd.n4848 gnd.n4845 10.6151
R16399 gnd.n4845 gnd.n4844 10.6151
R16400 gnd.n4844 gnd.n4841 10.6151
R16401 gnd.n4841 gnd.n4840 10.6151
R16402 gnd.n4837 gnd.n4836 10.6151
R16403 gnd.n4836 gnd.n4833 10.6151
R16404 gnd.n5742 gnd.n5740 10.6151
R16405 gnd.n5740 gnd.n5737 10.6151
R16406 gnd.n5737 gnd.n5736 10.6151
R16407 gnd.n5736 gnd.n5733 10.6151
R16408 gnd.n5733 gnd.n5732 10.6151
R16409 gnd.n5732 gnd.n5729 10.6151
R16410 gnd.n5729 gnd.n5728 10.6151
R16411 gnd.n5728 gnd.n5725 10.6151
R16412 gnd.n5725 gnd.n5724 10.6151
R16413 gnd.n5724 gnd.n5721 10.6151
R16414 gnd.n5721 gnd.n5720 10.6151
R16415 gnd.n5720 gnd.n5717 10.6151
R16416 gnd.n5717 gnd.n5716 10.6151
R16417 gnd.n5716 gnd.n5713 10.6151
R16418 gnd.n5713 gnd.n5712 10.6151
R16419 gnd.n5712 gnd.n5709 10.6151
R16420 gnd.n5709 gnd.n5708 10.6151
R16421 gnd.n5708 gnd.n5705 10.6151
R16422 gnd.n5705 gnd.n5704 10.6151
R16423 gnd.n5704 gnd.n5701 10.6151
R16424 gnd.n5701 gnd.n5700 10.6151
R16425 gnd.n5700 gnd.n5697 10.6151
R16426 gnd.n5697 gnd.n5696 10.6151
R16427 gnd.n5696 gnd.n5693 10.6151
R16428 gnd.n5693 gnd.n5692 10.6151
R16429 gnd.n5692 gnd.n5689 10.6151
R16430 gnd.n5689 gnd.n5688 10.6151
R16431 gnd.n5688 gnd.n5685 10.6151
R16432 gnd.n5683 gnd.n5680 10.6151
R16433 gnd.n5680 gnd.n5679 10.6151
R16434 gnd.n4919 gnd.n1762 10.6151
R16435 gnd.n4920 gnd.n4919 10.6151
R16436 gnd.n4929 gnd.n4920 10.6151
R16437 gnd.n4929 gnd.n4928 10.6151
R16438 gnd.n4928 gnd.n4927 10.6151
R16439 gnd.n4927 gnd.n4926 10.6151
R16440 gnd.n4926 gnd.n4921 10.6151
R16441 gnd.n4921 gnd.n1731 10.6151
R16442 gnd.n4988 gnd.n1731 10.6151
R16443 gnd.n4989 gnd.n4988 10.6151
R16444 gnd.n4990 gnd.n4989 10.6151
R16445 gnd.n4990 gnd.n1718 10.6151
R16446 gnd.n5007 gnd.n1718 10.6151
R16447 gnd.n5008 gnd.n5007 10.6151
R16448 gnd.n5009 gnd.n5008 10.6151
R16449 gnd.n5009 gnd.n1704 10.6151
R16450 gnd.n5061 gnd.n1704 10.6151
R16451 gnd.n5062 gnd.n5061 10.6151
R16452 gnd.n5063 gnd.n5062 10.6151
R16453 gnd.n5063 gnd.n1688 10.6151
R16454 gnd.n5078 gnd.n1688 10.6151
R16455 gnd.n5079 gnd.n5078 10.6151
R16456 gnd.n5081 gnd.n5079 10.6151
R16457 gnd.n5081 gnd.n5080 10.6151
R16458 gnd.n5080 gnd.n1670 10.6151
R16459 gnd.n5106 gnd.n1670 10.6151
R16460 gnd.n5107 gnd.n5106 10.6151
R16461 gnd.n5117 gnd.n5107 10.6151
R16462 gnd.n5117 gnd.n5116 10.6151
R16463 gnd.n5116 gnd.n5115 10.6151
R16464 gnd.n5115 gnd.n5114 10.6151
R16465 gnd.n5114 gnd.n5108 10.6151
R16466 gnd.n5108 gnd.n1647 10.6151
R16467 gnd.n5166 gnd.n1647 10.6151
R16468 gnd.n5167 gnd.n5166 10.6151
R16469 gnd.n5168 gnd.n5167 10.6151
R16470 gnd.n5168 gnd.n1633 10.6151
R16471 gnd.n5186 gnd.n1633 10.6151
R16472 gnd.n5187 gnd.n5186 10.6151
R16473 gnd.n5188 gnd.n5187 10.6151
R16474 gnd.n5188 gnd.n1619 10.6151
R16475 gnd.n5237 gnd.n1619 10.6151
R16476 gnd.n5238 gnd.n5237 10.6151
R16477 gnd.n5239 gnd.n5238 10.6151
R16478 gnd.n5239 gnd.n1603 10.6151
R16479 gnd.n5255 gnd.n1603 10.6151
R16480 gnd.n5256 gnd.n5255 10.6151
R16481 gnd.n5258 gnd.n5256 10.6151
R16482 gnd.n5258 gnd.n5257 10.6151
R16483 gnd.n5257 gnd.n1585 10.6151
R16484 gnd.n5283 gnd.n1585 10.6151
R16485 gnd.n5284 gnd.n5283 10.6151
R16486 gnd.n5294 gnd.n5284 10.6151
R16487 gnd.n5294 gnd.n5293 10.6151
R16488 gnd.n5293 gnd.n5292 10.6151
R16489 gnd.n5292 gnd.n5291 10.6151
R16490 gnd.n5291 gnd.n5285 10.6151
R16491 gnd.n5285 gnd.n1560 10.6151
R16492 gnd.n5344 gnd.n1560 10.6151
R16493 gnd.n5345 gnd.n5344 10.6151
R16494 gnd.n5346 gnd.n5345 10.6151
R16495 gnd.n5346 gnd.n1545 10.6151
R16496 gnd.n5363 gnd.n1545 10.6151
R16497 gnd.n5364 gnd.n5363 10.6151
R16498 gnd.n5365 gnd.n5364 10.6151
R16499 gnd.n5365 gnd.n1532 10.6151
R16500 gnd.n5400 gnd.n1532 10.6151
R16501 gnd.n5401 gnd.n5400 10.6151
R16502 gnd.n5402 gnd.n5401 10.6151
R16503 gnd.n5402 gnd.n1516 10.6151
R16504 gnd.n5417 gnd.n1516 10.6151
R16505 gnd.n5418 gnd.n5417 10.6151
R16506 gnd.n5420 gnd.n5418 10.6151
R16507 gnd.n5420 gnd.n5419 10.6151
R16508 gnd.n5419 gnd.n1497 10.6151
R16509 gnd.n5444 gnd.n1497 10.6151
R16510 gnd.n5445 gnd.n5444 10.6151
R16511 gnd.n5455 gnd.n5445 10.6151
R16512 gnd.n5455 gnd.n5454 10.6151
R16513 gnd.n5454 gnd.n5453 10.6151
R16514 gnd.n5453 gnd.n5452 10.6151
R16515 gnd.n5452 gnd.n5446 10.6151
R16516 gnd.n5446 gnd.n1466 10.6151
R16517 gnd.n5516 gnd.n1466 10.6151
R16518 gnd.n5517 gnd.n5516 10.6151
R16519 gnd.n5518 gnd.n5517 10.6151
R16520 gnd.n5518 gnd.n1454 10.6151
R16521 gnd.n5535 gnd.n1454 10.6151
R16522 gnd.n5536 gnd.n5535 10.6151
R16523 gnd.n5537 gnd.n5536 10.6151
R16524 gnd.n5537 gnd.n1440 10.6151
R16525 gnd.n5581 gnd.n1440 10.6151
R16526 gnd.n5582 gnd.n5581 10.6151
R16527 gnd.n5583 gnd.n5582 10.6151
R16528 gnd.n5583 gnd.n1424 10.6151
R16529 gnd.n5598 gnd.n1424 10.6151
R16530 gnd.n5599 gnd.n5598 10.6151
R16531 gnd.n5601 gnd.n5599 10.6151
R16532 gnd.n5601 gnd.n5600 10.6151
R16533 gnd.n5600 gnd.n1406 10.6151
R16534 gnd.n5625 gnd.n1406 10.6151
R16535 gnd.n5626 gnd.n5625 10.6151
R16536 gnd.n5629 gnd.n5626 10.6151
R16537 gnd.n5629 gnd.n5628 10.6151
R16538 gnd.n5628 gnd.n5627 10.6151
R16539 gnd.n5627 gnd.n1384 10.6151
R16540 gnd.n5654 gnd.n1384 10.6151
R16541 gnd.n5655 gnd.n5654 10.6151
R16542 gnd.n5745 gnd.n5655 10.6151
R16543 gnd.n5745 gnd.n5744 10.6151
R16544 gnd.n2931 gnd.n2930 10.5739
R16545 gnd.t87 gnd.n319 10.5161
R16546 gnd.n322 gnd.t202 10.5161
R16547 gnd.n3562 gnd.n3546 10.4732
R16548 gnd.n3530 gnd.n3514 10.4732
R16549 gnd.n3498 gnd.n3482 10.4732
R16550 gnd.n3467 gnd.n3451 10.4732
R16551 gnd.n3435 gnd.n3419 10.4732
R16552 gnd.n3403 gnd.n3387 10.4732
R16553 gnd.n3371 gnd.n3355 10.4732
R16554 gnd.n3340 gnd.n3324 10.4732
R16555 gnd.t264 gnd.n2611 10.3916
R16556 gnd.n4671 gnd.n1759 10.1975
R16557 gnd.n4924 gnd.n4923 10.1975
R16558 gnd.n5025 gnd.n1667 10.1975
R16559 gnd.n1583 gnd.n1581 10.1975
R16560 gnd.n5289 gnd.n5288 10.1975
R16561 gnd.n5450 gnd.n5449 10.1975
R16562 gnd.n5553 gnd.n1403 10.1975
R16563 gnd.n5556 gnd.n1386 10.1975
R16564 gnd.n2639 gnd.t277 10.027
R16565 gnd.t6 gnd.n352 9.87883
R16566 gnd.n292 gnd.t32 9.87883
R16567 gnd.n7607 gnd.n78 9.81789
R16568 gnd.n3566 gnd.n3565 9.69747
R16569 gnd.n3534 gnd.n3533 9.69747
R16570 gnd.n3502 gnd.n3501 9.69747
R16571 gnd.n3471 gnd.n3470 9.69747
R16572 gnd.n3439 gnd.n3438 9.69747
R16573 gnd.n3407 gnd.n3406 9.69747
R16574 gnd.n3375 gnd.n3374 9.69747
R16575 gnd.n3344 gnd.n3343 9.69747
R16576 gnd.n3038 gnd.t272 9.66242
R16577 gnd.n5013 gnd.n5011 9.56018
R16578 gnd.n4937 gnd.n1691 9.56018
R16579 gnd.n5191 gnd.n5190 9.56018
R16580 gnd.t42 gnd.n1631 9.56018
R16581 gnd.n5141 gnd.n1605 9.56018
R16582 gnd.n5368 gnd.n5367 9.56018
R16583 gnd.n5317 gnd.t48 9.56018
R16584 gnd.n5318 gnd.n1518 9.56018
R16585 gnd.n5540 gnd.n5539 9.56018
R16586 gnd.n5463 gnd.n1426 9.56018
R16587 gnd.n6055 gnd.n1098 9.45751
R16588 gnd.n7153 gnd.n7152 9.45599
R16589 gnd.n3572 gnd.n3571 9.45567
R16590 gnd.n3540 gnd.n3539 9.45567
R16591 gnd.n3508 gnd.n3507 9.45567
R16592 gnd.n3477 gnd.n3476 9.45567
R16593 gnd.n3445 gnd.n3444 9.45567
R16594 gnd.n3413 gnd.n3412 9.45567
R16595 gnd.n3381 gnd.n3380 9.45567
R16596 gnd.n3350 gnd.n3349 9.45567
R16597 gnd.n2518 gnd.n2517 9.39724
R16598 gnd.n7547 gnd.n134 9.3005
R16599 gnd.n7546 gnd.n136 9.3005
R16600 gnd.n140 gnd.n137 9.3005
R16601 gnd.n7541 gnd.n141 9.3005
R16602 gnd.n7540 gnd.n142 9.3005
R16603 gnd.n7539 gnd.n143 9.3005
R16604 gnd.n147 gnd.n144 9.3005
R16605 gnd.n7534 gnd.n148 9.3005
R16606 gnd.n7533 gnd.n149 9.3005
R16607 gnd.n7532 gnd.n150 9.3005
R16608 gnd.n154 gnd.n151 9.3005
R16609 gnd.n7527 gnd.n155 9.3005
R16610 gnd.n7526 gnd.n156 9.3005
R16611 gnd.n7525 gnd.n157 9.3005
R16612 gnd.n161 gnd.n158 9.3005
R16613 gnd.n7520 gnd.n162 9.3005
R16614 gnd.n7519 gnd.n163 9.3005
R16615 gnd.n7515 gnd.n164 9.3005
R16616 gnd.n168 gnd.n165 9.3005
R16617 gnd.n7510 gnd.n169 9.3005
R16618 gnd.n7509 gnd.n170 9.3005
R16619 gnd.n7508 gnd.n171 9.3005
R16620 gnd.n175 gnd.n172 9.3005
R16621 gnd.n7503 gnd.n176 9.3005
R16622 gnd.n7502 gnd.n177 9.3005
R16623 gnd.n7501 gnd.n178 9.3005
R16624 gnd.n182 gnd.n179 9.3005
R16625 gnd.n7496 gnd.n183 9.3005
R16626 gnd.n7495 gnd.n184 9.3005
R16627 gnd.n7494 gnd.n185 9.3005
R16628 gnd.n189 gnd.n186 9.3005
R16629 gnd.n7489 gnd.n190 9.3005
R16630 gnd.n7488 gnd.n191 9.3005
R16631 gnd.n7487 gnd.n192 9.3005
R16632 gnd.n196 gnd.n193 9.3005
R16633 gnd.n7482 gnd.n197 9.3005
R16634 gnd.n7481 gnd.n7480 9.3005
R16635 gnd.n7479 gnd.n200 9.3005
R16636 gnd.n7549 gnd.n7548 9.3005
R16637 gnd.n7026 gnd.n584 9.3005
R16638 gnd.n7025 gnd.n586 9.3005
R16639 gnd.n7024 gnd.n587 9.3005
R16640 gnd.n6812 gnd.n588 9.3005
R16641 gnd.n6816 gnd.n6813 9.3005
R16642 gnd.n6817 gnd.n6811 9.3005
R16643 gnd.n6821 gnd.n6820 9.3005
R16644 gnd.n6822 gnd.n6810 9.3005
R16645 gnd.n6953 gnd.n6823 9.3005
R16646 gnd.n6952 gnd.n6824 9.3005
R16647 gnd.n6951 gnd.n6825 9.3005
R16648 gnd.n6949 gnd.n6826 9.3005
R16649 gnd.n6948 gnd.n6827 9.3005
R16650 gnd.n6946 gnd.n6828 9.3005
R16651 gnd.n6945 gnd.n6829 9.3005
R16652 gnd.n6943 gnd.n6830 9.3005
R16653 gnd.n6942 gnd.n6831 9.3005
R16654 gnd.n6940 gnd.n6832 9.3005
R16655 gnd.n6939 gnd.n6833 9.3005
R16656 gnd.n6937 gnd.n6834 9.3005
R16657 gnd.n6936 gnd.n6835 9.3005
R16658 gnd.n6934 gnd.n6836 9.3005
R16659 gnd.n6933 gnd.n6837 9.3005
R16660 gnd.n6931 gnd.n6838 9.3005
R16661 gnd.n6930 gnd.n6839 9.3005
R16662 gnd.n6928 gnd.n6840 9.3005
R16663 gnd.n6927 gnd.n6841 9.3005
R16664 gnd.n6925 gnd.n6842 9.3005
R16665 gnd.n6924 gnd.n6843 9.3005
R16666 gnd.n6922 gnd.n6844 9.3005
R16667 gnd.n6921 gnd.n6845 9.3005
R16668 gnd.n6919 gnd.n325 9.3005
R16669 gnd.n6918 gnd.n6846 9.3005
R16670 gnd.n6916 gnd.n6847 9.3005
R16671 gnd.n6915 gnd.n6848 9.3005
R16672 gnd.n6913 gnd.n6849 9.3005
R16673 gnd.n6912 gnd.n6850 9.3005
R16674 gnd.n6910 gnd.n6851 9.3005
R16675 gnd.n6909 gnd.n6852 9.3005
R16676 gnd.n6907 gnd.n6853 9.3005
R16677 gnd.n6906 gnd.n6854 9.3005
R16678 gnd.n6904 gnd.n6855 9.3005
R16679 gnd.n6903 gnd.n6856 9.3005
R16680 gnd.n6901 gnd.n6857 9.3005
R16681 gnd.n6900 gnd.n6858 9.3005
R16682 gnd.n6898 gnd.n6859 9.3005
R16683 gnd.n6897 gnd.n6860 9.3005
R16684 gnd.n6895 gnd.n6861 9.3005
R16685 gnd.n6894 gnd.n6862 9.3005
R16686 gnd.n6892 gnd.n6863 9.3005
R16687 gnd.n6891 gnd.n6864 9.3005
R16688 gnd.n6889 gnd.n6865 9.3005
R16689 gnd.n6888 gnd.n6866 9.3005
R16690 gnd.n6886 gnd.n6867 9.3005
R16691 gnd.n6885 gnd.n6868 9.3005
R16692 gnd.n6883 gnd.n6869 9.3005
R16693 gnd.n6882 gnd.n6870 9.3005
R16694 gnd.n6880 gnd.n6871 9.3005
R16695 gnd.n6879 gnd.n6872 9.3005
R16696 gnd.n6877 gnd.n6873 9.3005
R16697 gnd.n6876 gnd.n6875 9.3005
R16698 gnd.n6874 gnd.n204 9.3005
R16699 gnd.n7476 gnd.n203 9.3005
R16700 gnd.n7478 gnd.n7477 9.3005
R16701 gnd.n7028 gnd.n7027 9.3005
R16702 gnd.n7034 gnd.n7033 9.3005
R16703 gnd.n7035 gnd.n578 9.3005
R16704 gnd.n7038 gnd.n577 9.3005
R16705 gnd.n7039 gnd.n576 9.3005
R16706 gnd.n7042 gnd.n575 9.3005
R16707 gnd.n7043 gnd.n574 9.3005
R16708 gnd.n7046 gnd.n573 9.3005
R16709 gnd.n7047 gnd.n572 9.3005
R16710 gnd.n7050 gnd.n571 9.3005
R16711 gnd.n7051 gnd.n570 9.3005
R16712 gnd.n7054 gnd.n569 9.3005
R16713 gnd.n7055 gnd.n568 9.3005
R16714 gnd.n7058 gnd.n567 9.3005
R16715 gnd.n7059 gnd.n566 9.3005
R16716 gnd.n7062 gnd.n565 9.3005
R16717 gnd.n7063 gnd.n564 9.3005
R16718 gnd.n7066 gnd.n563 9.3005
R16719 gnd.n7067 gnd.n562 9.3005
R16720 gnd.n7070 gnd.n561 9.3005
R16721 gnd.n7072 gnd.n555 9.3005
R16722 gnd.n7075 gnd.n554 9.3005
R16723 gnd.n7076 gnd.n553 9.3005
R16724 gnd.n7079 gnd.n552 9.3005
R16725 gnd.n7080 gnd.n551 9.3005
R16726 gnd.n7083 gnd.n550 9.3005
R16727 gnd.n7084 gnd.n549 9.3005
R16728 gnd.n7087 gnd.n548 9.3005
R16729 gnd.n7088 gnd.n547 9.3005
R16730 gnd.n7091 gnd.n546 9.3005
R16731 gnd.n7092 gnd.n545 9.3005
R16732 gnd.n7095 gnd.n544 9.3005
R16733 gnd.n7097 gnd.n543 9.3005
R16734 gnd.n7098 gnd.n542 9.3005
R16735 gnd.n7099 gnd.n541 9.3005
R16736 gnd.n540 gnd.n448 9.3005
R16737 gnd.n7032 gnd.n583 9.3005
R16738 gnd.n7031 gnd.n7030 9.3005
R16739 gnd.n7161 gnd.n447 9.3005
R16740 gnd.n7163 gnd.n7162 9.3005
R16741 gnd.n432 gnd.n431 9.3005
R16742 gnd.n7176 gnd.n7175 9.3005
R16743 gnd.n7177 gnd.n430 9.3005
R16744 gnd.n7179 gnd.n7178 9.3005
R16745 gnd.n414 gnd.n413 9.3005
R16746 gnd.n7192 gnd.n7191 9.3005
R16747 gnd.n7193 gnd.n412 9.3005
R16748 gnd.n7195 gnd.n7194 9.3005
R16749 gnd.n399 gnd.n398 9.3005
R16750 gnd.n7208 gnd.n7207 9.3005
R16751 gnd.n7209 gnd.n397 9.3005
R16752 gnd.n7211 gnd.n7210 9.3005
R16753 gnd.n382 gnd.n381 9.3005
R16754 gnd.n7224 gnd.n7223 9.3005
R16755 gnd.n7225 gnd.n380 9.3005
R16756 gnd.n7227 gnd.n7226 9.3005
R16757 gnd.n367 gnd.n366 9.3005
R16758 gnd.n7240 gnd.n7239 9.3005
R16759 gnd.n7241 gnd.n365 9.3005
R16760 gnd.n7243 gnd.n7242 9.3005
R16761 gnd.n350 gnd.n349 9.3005
R16762 gnd.n7256 gnd.n7255 9.3005
R16763 gnd.n7257 gnd.n348 9.3005
R16764 gnd.n7259 gnd.n7258 9.3005
R16765 gnd.n335 gnd.n334 9.3005
R16766 gnd.n7272 gnd.n7271 9.3005
R16767 gnd.n7273 gnd.n333 9.3005
R16768 gnd.n7275 gnd.n7274 9.3005
R16769 gnd.n317 gnd.n316 9.3005
R16770 gnd.n7288 gnd.n7287 9.3005
R16771 gnd.n7289 gnd.n315 9.3005
R16772 gnd.n7291 gnd.n7290 9.3005
R16773 gnd.n303 gnd.n302 9.3005
R16774 gnd.n7304 gnd.n7303 9.3005
R16775 gnd.n7305 gnd.n301 9.3005
R16776 gnd.n7307 gnd.n7306 9.3005
R16777 gnd.n287 gnd.n286 9.3005
R16778 gnd.n7320 gnd.n7319 9.3005
R16779 gnd.n7321 gnd.n285 9.3005
R16780 gnd.n7323 gnd.n7322 9.3005
R16781 gnd.n273 gnd.n272 9.3005
R16782 gnd.n7336 gnd.n7335 9.3005
R16783 gnd.n7337 gnd.n271 9.3005
R16784 gnd.n7339 gnd.n7338 9.3005
R16785 gnd.n257 gnd.n256 9.3005
R16786 gnd.n7352 gnd.n7351 9.3005
R16787 gnd.n7353 gnd.n255 9.3005
R16788 gnd.n7355 gnd.n7354 9.3005
R16789 gnd.n243 gnd.n242 9.3005
R16790 gnd.n7368 gnd.n7367 9.3005
R16791 gnd.n7369 gnd.n241 9.3005
R16792 gnd.n7371 gnd.n7370 9.3005
R16793 gnd.n227 gnd.n226 9.3005
R16794 gnd.n7384 gnd.n7383 9.3005
R16795 gnd.n7385 gnd.n225 9.3005
R16796 gnd.n7387 gnd.n7386 9.3005
R16797 gnd.n211 gnd.n210 9.3005
R16798 gnd.n7468 gnd.n7467 9.3005
R16799 gnd.n7469 gnd.n209 9.3005
R16800 gnd.n7471 gnd.n7470 9.3005
R16801 gnd.n133 gnd.n132 9.3005
R16802 gnd.n7551 gnd.n7550 9.3005
R16803 gnd.n7160 gnd.n7159 9.3005
R16804 gnd.n6251 gnd.n923 9.3005
R16805 gnd.n6253 gnd.n6252 9.3005
R16806 gnd.n919 gnd.n918 9.3005
R16807 gnd.n6260 gnd.n6259 9.3005
R16808 gnd.n6261 gnd.n917 9.3005
R16809 gnd.n6263 gnd.n6262 9.3005
R16810 gnd.n913 gnd.n912 9.3005
R16811 gnd.n6270 gnd.n6269 9.3005
R16812 gnd.n6271 gnd.n911 9.3005
R16813 gnd.n6273 gnd.n6272 9.3005
R16814 gnd.n907 gnd.n906 9.3005
R16815 gnd.n6280 gnd.n6279 9.3005
R16816 gnd.n6281 gnd.n905 9.3005
R16817 gnd.n6283 gnd.n6282 9.3005
R16818 gnd.n901 gnd.n900 9.3005
R16819 gnd.n6290 gnd.n6289 9.3005
R16820 gnd.n6291 gnd.n899 9.3005
R16821 gnd.n6293 gnd.n6292 9.3005
R16822 gnd.n895 gnd.n894 9.3005
R16823 gnd.n6300 gnd.n6299 9.3005
R16824 gnd.n6301 gnd.n893 9.3005
R16825 gnd.n6303 gnd.n6302 9.3005
R16826 gnd.n889 gnd.n888 9.3005
R16827 gnd.n6310 gnd.n6309 9.3005
R16828 gnd.n6311 gnd.n887 9.3005
R16829 gnd.n6313 gnd.n6312 9.3005
R16830 gnd.n883 gnd.n882 9.3005
R16831 gnd.n6320 gnd.n6319 9.3005
R16832 gnd.n6321 gnd.n881 9.3005
R16833 gnd.n6323 gnd.n6322 9.3005
R16834 gnd.n877 gnd.n876 9.3005
R16835 gnd.n6330 gnd.n6329 9.3005
R16836 gnd.n6331 gnd.n875 9.3005
R16837 gnd.n6333 gnd.n6332 9.3005
R16838 gnd.n871 gnd.n870 9.3005
R16839 gnd.n6340 gnd.n6339 9.3005
R16840 gnd.n6341 gnd.n869 9.3005
R16841 gnd.n6343 gnd.n6342 9.3005
R16842 gnd.n865 gnd.n864 9.3005
R16843 gnd.n6350 gnd.n6349 9.3005
R16844 gnd.n6351 gnd.n863 9.3005
R16845 gnd.n6353 gnd.n6352 9.3005
R16846 gnd.n859 gnd.n858 9.3005
R16847 gnd.n6360 gnd.n6359 9.3005
R16848 gnd.n6361 gnd.n857 9.3005
R16849 gnd.n6363 gnd.n6362 9.3005
R16850 gnd.n853 gnd.n852 9.3005
R16851 gnd.n6370 gnd.n6369 9.3005
R16852 gnd.n6371 gnd.n851 9.3005
R16853 gnd.n6373 gnd.n6372 9.3005
R16854 gnd.n847 gnd.n846 9.3005
R16855 gnd.n6380 gnd.n6379 9.3005
R16856 gnd.n6381 gnd.n845 9.3005
R16857 gnd.n6383 gnd.n6382 9.3005
R16858 gnd.n841 gnd.n840 9.3005
R16859 gnd.n6390 gnd.n6389 9.3005
R16860 gnd.n6391 gnd.n839 9.3005
R16861 gnd.n6393 gnd.n6392 9.3005
R16862 gnd.n835 gnd.n834 9.3005
R16863 gnd.n6400 gnd.n6399 9.3005
R16864 gnd.n6401 gnd.n833 9.3005
R16865 gnd.n6403 gnd.n6402 9.3005
R16866 gnd.n829 gnd.n828 9.3005
R16867 gnd.n6410 gnd.n6409 9.3005
R16868 gnd.n6411 gnd.n827 9.3005
R16869 gnd.n6413 gnd.n6412 9.3005
R16870 gnd.n823 gnd.n822 9.3005
R16871 gnd.n6420 gnd.n6419 9.3005
R16872 gnd.n6421 gnd.n821 9.3005
R16873 gnd.n6423 gnd.n6422 9.3005
R16874 gnd.n817 gnd.n816 9.3005
R16875 gnd.n6430 gnd.n6429 9.3005
R16876 gnd.n6431 gnd.n815 9.3005
R16877 gnd.n6433 gnd.n6432 9.3005
R16878 gnd.n811 gnd.n810 9.3005
R16879 gnd.n6440 gnd.n6439 9.3005
R16880 gnd.n6441 gnd.n809 9.3005
R16881 gnd.n6443 gnd.n6442 9.3005
R16882 gnd.n805 gnd.n804 9.3005
R16883 gnd.n6450 gnd.n6449 9.3005
R16884 gnd.n6451 gnd.n803 9.3005
R16885 gnd.n6453 gnd.n6452 9.3005
R16886 gnd.n799 gnd.n798 9.3005
R16887 gnd.n6460 gnd.n6459 9.3005
R16888 gnd.n6461 gnd.n797 9.3005
R16889 gnd.n6463 gnd.n6462 9.3005
R16890 gnd.n793 gnd.n792 9.3005
R16891 gnd.n6470 gnd.n6469 9.3005
R16892 gnd.n6471 gnd.n791 9.3005
R16893 gnd.n6473 gnd.n6472 9.3005
R16894 gnd.n787 gnd.n786 9.3005
R16895 gnd.n6480 gnd.n6479 9.3005
R16896 gnd.n6481 gnd.n785 9.3005
R16897 gnd.n6483 gnd.n6482 9.3005
R16898 gnd.n781 gnd.n780 9.3005
R16899 gnd.n6490 gnd.n6489 9.3005
R16900 gnd.n6491 gnd.n779 9.3005
R16901 gnd.n6493 gnd.n6492 9.3005
R16902 gnd.n775 gnd.n774 9.3005
R16903 gnd.n6500 gnd.n6499 9.3005
R16904 gnd.n6501 gnd.n773 9.3005
R16905 gnd.n6503 gnd.n6502 9.3005
R16906 gnd.n769 gnd.n768 9.3005
R16907 gnd.n6510 gnd.n6509 9.3005
R16908 gnd.n6511 gnd.n767 9.3005
R16909 gnd.n6513 gnd.n6512 9.3005
R16910 gnd.n763 gnd.n762 9.3005
R16911 gnd.n6520 gnd.n6519 9.3005
R16912 gnd.n6521 gnd.n761 9.3005
R16913 gnd.n6523 gnd.n6522 9.3005
R16914 gnd.n757 gnd.n756 9.3005
R16915 gnd.n6530 gnd.n6529 9.3005
R16916 gnd.n6531 gnd.n755 9.3005
R16917 gnd.n6533 gnd.n6532 9.3005
R16918 gnd.n751 gnd.n750 9.3005
R16919 gnd.n6540 gnd.n6539 9.3005
R16920 gnd.n6541 gnd.n749 9.3005
R16921 gnd.n6543 gnd.n6542 9.3005
R16922 gnd.n745 gnd.n744 9.3005
R16923 gnd.n6550 gnd.n6549 9.3005
R16924 gnd.n6551 gnd.n743 9.3005
R16925 gnd.n6553 gnd.n6552 9.3005
R16926 gnd.n739 gnd.n738 9.3005
R16927 gnd.n6560 gnd.n6559 9.3005
R16928 gnd.n6561 gnd.n737 9.3005
R16929 gnd.n6564 gnd.n6563 9.3005
R16930 gnd.n6562 gnd.n733 9.3005
R16931 gnd.n6570 gnd.n732 9.3005
R16932 gnd.n6572 gnd.n6571 9.3005
R16933 gnd.n728 gnd.n727 9.3005
R16934 gnd.n6581 gnd.n6580 9.3005
R16935 gnd.n6582 gnd.n726 9.3005
R16936 gnd.n6584 gnd.n6583 9.3005
R16937 gnd.n722 gnd.n721 9.3005
R16938 gnd.n6591 gnd.n6590 9.3005
R16939 gnd.n6592 gnd.n720 9.3005
R16940 gnd.n6594 gnd.n6593 9.3005
R16941 gnd.n716 gnd.n715 9.3005
R16942 gnd.n6601 gnd.n6600 9.3005
R16943 gnd.n6602 gnd.n714 9.3005
R16944 gnd.n6604 gnd.n6603 9.3005
R16945 gnd.n710 gnd.n709 9.3005
R16946 gnd.n6611 gnd.n6610 9.3005
R16947 gnd.n6612 gnd.n708 9.3005
R16948 gnd.n6614 gnd.n6613 9.3005
R16949 gnd.n704 gnd.n703 9.3005
R16950 gnd.n6621 gnd.n6620 9.3005
R16951 gnd.n6622 gnd.n702 9.3005
R16952 gnd.n6624 gnd.n6623 9.3005
R16953 gnd.n698 gnd.n697 9.3005
R16954 gnd.n6631 gnd.n6630 9.3005
R16955 gnd.n6632 gnd.n696 9.3005
R16956 gnd.n6634 gnd.n6633 9.3005
R16957 gnd.n692 gnd.n691 9.3005
R16958 gnd.n6641 gnd.n6640 9.3005
R16959 gnd.n6642 gnd.n690 9.3005
R16960 gnd.n6644 gnd.n6643 9.3005
R16961 gnd.n686 gnd.n685 9.3005
R16962 gnd.n6651 gnd.n6650 9.3005
R16963 gnd.n6652 gnd.n684 9.3005
R16964 gnd.n6654 gnd.n6653 9.3005
R16965 gnd.n680 gnd.n679 9.3005
R16966 gnd.n6661 gnd.n6660 9.3005
R16967 gnd.n6662 gnd.n678 9.3005
R16968 gnd.n6664 gnd.n6663 9.3005
R16969 gnd.n674 gnd.n673 9.3005
R16970 gnd.n6671 gnd.n6670 9.3005
R16971 gnd.n6672 gnd.n672 9.3005
R16972 gnd.n6674 gnd.n6673 9.3005
R16973 gnd.n668 gnd.n667 9.3005
R16974 gnd.n6681 gnd.n6680 9.3005
R16975 gnd.n6682 gnd.n666 9.3005
R16976 gnd.n6684 gnd.n6683 9.3005
R16977 gnd.n662 gnd.n661 9.3005
R16978 gnd.n6691 gnd.n6690 9.3005
R16979 gnd.n6692 gnd.n660 9.3005
R16980 gnd.n6694 gnd.n6693 9.3005
R16981 gnd.n656 gnd.n655 9.3005
R16982 gnd.n6701 gnd.n6700 9.3005
R16983 gnd.n6702 gnd.n654 9.3005
R16984 gnd.n6704 gnd.n6703 9.3005
R16985 gnd.n650 gnd.n649 9.3005
R16986 gnd.n6711 gnd.n6710 9.3005
R16987 gnd.n6712 gnd.n648 9.3005
R16988 gnd.n6714 gnd.n6713 9.3005
R16989 gnd.n644 gnd.n643 9.3005
R16990 gnd.n6721 gnd.n6720 9.3005
R16991 gnd.n6722 gnd.n642 9.3005
R16992 gnd.n6724 gnd.n6723 9.3005
R16993 gnd.n638 gnd.n637 9.3005
R16994 gnd.n6731 gnd.n6730 9.3005
R16995 gnd.n6732 gnd.n636 9.3005
R16996 gnd.n6734 gnd.n6733 9.3005
R16997 gnd.n632 gnd.n631 9.3005
R16998 gnd.n6741 gnd.n6740 9.3005
R16999 gnd.n6742 gnd.n630 9.3005
R17000 gnd.n6744 gnd.n6743 9.3005
R17001 gnd.n626 gnd.n625 9.3005
R17002 gnd.n6751 gnd.n6750 9.3005
R17003 gnd.n6752 gnd.n624 9.3005
R17004 gnd.n6754 gnd.n6753 9.3005
R17005 gnd.n620 gnd.n619 9.3005
R17006 gnd.n6761 gnd.n6760 9.3005
R17007 gnd.n6762 gnd.n618 9.3005
R17008 gnd.n6764 gnd.n6763 9.3005
R17009 gnd.n614 gnd.n613 9.3005
R17010 gnd.n6771 gnd.n6770 9.3005
R17011 gnd.n6772 gnd.n612 9.3005
R17012 gnd.n6774 gnd.n6773 9.3005
R17013 gnd.n608 gnd.n607 9.3005
R17014 gnd.n6783 gnd.n6782 9.3005
R17015 gnd.n6784 gnd.n606 9.3005
R17016 gnd.n6786 gnd.n6785 9.3005
R17017 gnd.n6574 gnd.n6573 9.3005
R17018 gnd.n4459 gnd.n4458 9.3005
R17019 gnd.n4462 gnd.n4461 9.3005
R17020 gnd.n4463 gnd.n4456 9.3005
R17021 gnd.n4465 gnd.n4464 9.3005
R17022 gnd.n4454 gnd.n4453 9.3005
R17023 gnd.n4470 gnd.n4469 9.3005
R17024 gnd.n4471 gnd.n4452 9.3005
R17025 gnd.n4771 gnd.n4472 9.3005
R17026 gnd.n4770 gnd.n4473 9.3005
R17027 gnd.n4769 gnd.n4474 9.3005
R17028 gnd.n4615 gnd.n4475 9.3005
R17029 gnd.n4617 gnd.n4616 9.3005
R17030 gnd.n4614 gnd.n4613 9.3005
R17031 gnd.n4627 gnd.n4626 9.3005
R17032 gnd.n4628 gnd.n4612 9.3005
R17033 gnd.n4630 gnd.n4629 9.3005
R17034 gnd.n4608 gnd.n4607 9.3005
R17035 gnd.n4643 gnd.n4642 9.3005
R17036 gnd.n4644 gnd.n4606 9.3005
R17037 gnd.n4646 gnd.n4645 9.3005
R17038 gnd.n4602 gnd.n4601 9.3005
R17039 gnd.n4659 gnd.n4658 9.3005
R17040 gnd.n4660 gnd.n4600 9.3005
R17041 gnd.n4662 gnd.n4661 9.3005
R17042 gnd.n1770 gnd.n1769 9.3005
R17043 gnd.n4909 gnd.n4908 9.3005
R17044 gnd.n4910 gnd.n1768 9.3005
R17045 gnd.n4912 gnd.n4911 9.3005
R17046 gnd.n1749 gnd.n1748 9.3005
R17047 gnd.n4968 gnd.n4967 9.3005
R17048 gnd.n4969 gnd.n1747 9.3005
R17049 gnd.n4971 gnd.n4970 9.3005
R17050 gnd.n1726 gnd.n1725 9.3005
R17051 gnd.n4996 gnd.n4995 9.3005
R17052 gnd.n4997 gnd.n1724 9.3005
R17053 gnd.n5001 gnd.n4998 9.3005
R17054 gnd.n5000 gnd.n4999 9.3005
R17055 gnd.n1698 gnd.n1697 9.3005
R17056 gnd.n5070 gnd.n5069 9.3005
R17057 gnd.n5071 gnd.n1696 9.3005
R17058 gnd.n5073 gnd.n5072 9.3005
R17059 gnd.n1678 gnd.n1677 9.3005
R17060 gnd.n5095 gnd.n5094 9.3005
R17061 gnd.n5096 gnd.n1676 9.3005
R17062 gnd.n5098 gnd.n5097 9.3005
R17063 gnd.n1658 gnd.n1657 9.3005
R17064 gnd.n5129 gnd.n5128 9.3005
R17065 gnd.n5130 gnd.n1656 9.3005
R17066 gnd.n5132 gnd.n5131 9.3005
R17067 gnd.n1641 gnd.n1640 9.3005
R17068 gnd.n5174 gnd.n5173 9.3005
R17069 gnd.n5175 gnd.n1639 9.3005
R17070 gnd.n5179 gnd.n5176 9.3005
R17071 gnd.n5178 gnd.n5177 9.3005
R17072 gnd.n1613 gnd.n1612 9.3005
R17073 gnd.n5247 gnd.n5246 9.3005
R17074 gnd.n5248 gnd.n1611 9.3005
R17075 gnd.n5250 gnd.n5249 9.3005
R17076 gnd.n1593 gnd.n1592 9.3005
R17077 gnd.n5273 gnd.n5272 9.3005
R17078 gnd.n5274 gnd.n1591 9.3005
R17079 gnd.n5276 gnd.n5275 9.3005
R17080 gnd.n1570 gnd.n1569 9.3005
R17081 gnd.n5306 gnd.n5305 9.3005
R17082 gnd.n5307 gnd.n1568 9.3005
R17083 gnd.n5309 gnd.n5308 9.3005
R17084 gnd.n1553 gnd.n1552 9.3005
R17085 gnd.n5352 gnd.n5351 9.3005
R17086 gnd.n5353 gnd.n1551 9.3005
R17087 gnd.n5357 gnd.n5354 9.3005
R17088 gnd.n5356 gnd.n5355 9.3005
R17089 gnd.n1526 gnd.n1525 9.3005
R17090 gnd.n5409 gnd.n5408 9.3005
R17091 gnd.n5410 gnd.n1524 9.3005
R17092 gnd.n5412 gnd.n5411 9.3005
R17093 gnd.n1505 gnd.n1504 9.3005
R17094 gnd.n5434 gnd.n5433 9.3005
R17095 gnd.n5435 gnd.n1503 9.3005
R17096 gnd.n5437 gnd.n5436 9.3005
R17097 gnd.n1483 gnd.n1482 9.3005
R17098 gnd.n5495 gnd.n5494 9.3005
R17099 gnd.n5496 gnd.n1481 9.3005
R17100 gnd.n5498 gnd.n5497 9.3005
R17101 gnd.n1461 gnd.n1460 9.3005
R17102 gnd.n5524 gnd.n5523 9.3005
R17103 gnd.n5525 gnd.n1459 9.3005
R17104 gnd.n5529 gnd.n5526 9.3005
R17105 gnd.n5528 gnd.n5527 9.3005
R17106 gnd.n1434 gnd.n1433 9.3005
R17107 gnd.n5590 gnd.n5589 9.3005
R17108 gnd.n5591 gnd.n1432 9.3005
R17109 gnd.n5593 gnd.n5592 9.3005
R17110 gnd.n1414 gnd.n1413 9.3005
R17111 gnd.n5615 gnd.n5614 9.3005
R17112 gnd.n5616 gnd.n1412 9.3005
R17113 gnd.n5618 gnd.n5617 9.3005
R17114 gnd.n1394 gnd.n1393 9.3005
R17115 gnd.n5643 gnd.n5642 9.3005
R17116 gnd.n5644 gnd.n1392 9.3005
R17117 gnd.n5648 gnd.n5645 9.3005
R17118 gnd.n5647 gnd.n5646 9.3005
R17119 gnd.n1332 gnd.n1331 9.3005
R17120 gnd.n5832 gnd.n5831 9.3005
R17121 gnd.n5833 gnd.n1330 9.3005
R17122 gnd.n5835 gnd.n5834 9.3005
R17123 gnd.n1319 gnd.n1318 9.3005
R17124 gnd.n5852 gnd.n5851 9.3005
R17125 gnd.n5853 gnd.n1317 9.3005
R17126 gnd.n5855 gnd.n5854 9.3005
R17127 gnd.n1306 gnd.n1305 9.3005
R17128 gnd.n5875 gnd.n5874 9.3005
R17129 gnd.n5876 gnd.n1304 9.3005
R17130 gnd.n5879 gnd.n5878 9.3005
R17131 gnd.n5877 gnd.n1232 9.3005
R17132 gnd.n5896 gnd.n1233 9.3005
R17133 gnd.n5895 gnd.n1234 9.3005
R17134 gnd.n5894 gnd.n1235 9.3005
R17135 gnd.n1238 gnd.n1236 9.3005
R17136 gnd.n1243 gnd.n1239 9.3005
R17137 gnd.n1242 gnd.n1241 9.3005
R17138 gnd.n1240 gnd.n595 9.3005
R17139 gnd.n6797 gnd.n596 9.3005
R17140 gnd.n6796 gnd.n597 9.3005
R17141 gnd.n6795 gnd.n598 9.3005
R17142 gnd.n601 gnd.n599 9.3005
R17143 gnd.n6791 gnd.n602 9.3005
R17144 gnd.n6790 gnd.n603 9.3005
R17145 gnd.n6789 gnd.n604 9.3005
R17146 gnd.n4457 gnd.n1055 9.3005
R17147 gnd.n6083 gnd.n1052 9.3005
R17148 gnd.n6086 gnd.n1051 9.3005
R17149 gnd.n6087 gnd.n1050 9.3005
R17150 gnd.n6090 gnd.n1049 9.3005
R17151 gnd.n6091 gnd.n1048 9.3005
R17152 gnd.n6094 gnd.n1047 9.3005
R17153 gnd.n6095 gnd.n1046 9.3005
R17154 gnd.n6098 gnd.n1045 9.3005
R17155 gnd.n6099 gnd.n1044 9.3005
R17156 gnd.n6102 gnd.n1043 9.3005
R17157 gnd.n6103 gnd.n1042 9.3005
R17158 gnd.n6106 gnd.n1041 9.3005
R17159 gnd.n6107 gnd.n1040 9.3005
R17160 gnd.n6110 gnd.n1039 9.3005
R17161 gnd.n6111 gnd.n1038 9.3005
R17162 gnd.n6114 gnd.n1037 9.3005
R17163 gnd.n6115 gnd.n1036 9.3005
R17164 gnd.n6118 gnd.n1035 9.3005
R17165 gnd.n6119 gnd.n1034 9.3005
R17166 gnd.n6122 gnd.n1033 9.3005
R17167 gnd.n6123 gnd.n1032 9.3005
R17168 gnd.n6126 gnd.n1031 9.3005
R17169 gnd.n6127 gnd.n1030 9.3005
R17170 gnd.n6130 gnd.n1029 9.3005
R17171 gnd.n6131 gnd.n1028 9.3005
R17172 gnd.n6134 gnd.n1027 9.3005
R17173 gnd.n6135 gnd.n1026 9.3005
R17174 gnd.n6138 gnd.n1025 9.3005
R17175 gnd.n6139 gnd.n1024 9.3005
R17176 gnd.n6142 gnd.n1023 9.3005
R17177 gnd.n6143 gnd.n1022 9.3005
R17178 gnd.n6146 gnd.n1021 9.3005
R17179 gnd.n6147 gnd.n1020 9.3005
R17180 gnd.n6150 gnd.n1019 9.3005
R17181 gnd.n6151 gnd.n1018 9.3005
R17182 gnd.n6154 gnd.n1017 9.3005
R17183 gnd.n6155 gnd.n1016 9.3005
R17184 gnd.n6158 gnd.n1015 9.3005
R17185 gnd.n6159 gnd.n1014 9.3005
R17186 gnd.n6162 gnd.n1013 9.3005
R17187 gnd.n6163 gnd.n1012 9.3005
R17188 gnd.n6166 gnd.n1011 9.3005
R17189 gnd.n6167 gnd.n1010 9.3005
R17190 gnd.n6170 gnd.n1009 9.3005
R17191 gnd.n6171 gnd.n1008 9.3005
R17192 gnd.n6174 gnd.n1007 9.3005
R17193 gnd.n6175 gnd.n1006 9.3005
R17194 gnd.n6178 gnd.n1005 9.3005
R17195 gnd.n6179 gnd.n1004 9.3005
R17196 gnd.n6182 gnd.n1003 9.3005
R17197 gnd.n6183 gnd.n1002 9.3005
R17198 gnd.n6186 gnd.n1001 9.3005
R17199 gnd.n6187 gnd.n1000 9.3005
R17200 gnd.n6190 gnd.n999 9.3005
R17201 gnd.n6191 gnd.n998 9.3005
R17202 gnd.n6194 gnd.n997 9.3005
R17203 gnd.n6195 gnd.n996 9.3005
R17204 gnd.n6198 gnd.n995 9.3005
R17205 gnd.n6199 gnd.n994 9.3005
R17206 gnd.n6202 gnd.n993 9.3005
R17207 gnd.n6203 gnd.n992 9.3005
R17208 gnd.n6206 gnd.n991 9.3005
R17209 gnd.n6207 gnd.n990 9.3005
R17210 gnd.n6210 gnd.n989 9.3005
R17211 gnd.n6211 gnd.n988 9.3005
R17212 gnd.n6214 gnd.n987 9.3005
R17213 gnd.n6215 gnd.n986 9.3005
R17214 gnd.n6218 gnd.n985 9.3005
R17215 gnd.n6219 gnd.n984 9.3005
R17216 gnd.n6222 gnd.n983 9.3005
R17217 gnd.n6223 gnd.n982 9.3005
R17218 gnd.n6226 gnd.n981 9.3005
R17219 gnd.n6227 gnd.n980 9.3005
R17220 gnd.n6230 gnd.n979 9.3005
R17221 gnd.n6231 gnd.n978 9.3005
R17222 gnd.n6234 gnd.n977 9.3005
R17223 gnd.n6235 gnd.n976 9.3005
R17224 gnd.n6238 gnd.n975 9.3005
R17225 gnd.n6239 gnd.n974 9.3005
R17226 gnd.n6242 gnd.n973 9.3005
R17227 gnd.n6243 gnd.n972 9.3005
R17228 gnd.n6244 gnd.n971 9.3005
R17229 gnd.n925 gnd.n924 9.3005
R17230 gnd.n6250 gnd.n6249 9.3005
R17231 gnd.n6082 gnd.n1053 9.3005
R17232 gnd.n3571 gnd.n3570 9.3005
R17233 gnd.n3544 gnd.n3543 9.3005
R17234 gnd.n3565 gnd.n3564 9.3005
R17235 gnd.n3563 gnd.n3562 9.3005
R17236 gnd.n3548 gnd.n3547 9.3005
R17237 gnd.n3557 gnd.n3556 9.3005
R17238 gnd.n3555 gnd.n3554 9.3005
R17239 gnd.n3539 gnd.n3538 9.3005
R17240 gnd.n3512 gnd.n3511 9.3005
R17241 gnd.n3533 gnd.n3532 9.3005
R17242 gnd.n3531 gnd.n3530 9.3005
R17243 gnd.n3516 gnd.n3515 9.3005
R17244 gnd.n3525 gnd.n3524 9.3005
R17245 gnd.n3523 gnd.n3522 9.3005
R17246 gnd.n3507 gnd.n3506 9.3005
R17247 gnd.n3480 gnd.n3479 9.3005
R17248 gnd.n3501 gnd.n3500 9.3005
R17249 gnd.n3499 gnd.n3498 9.3005
R17250 gnd.n3484 gnd.n3483 9.3005
R17251 gnd.n3493 gnd.n3492 9.3005
R17252 gnd.n3491 gnd.n3490 9.3005
R17253 gnd.n3476 gnd.n3475 9.3005
R17254 gnd.n3449 gnd.n3448 9.3005
R17255 gnd.n3470 gnd.n3469 9.3005
R17256 gnd.n3468 gnd.n3467 9.3005
R17257 gnd.n3453 gnd.n3452 9.3005
R17258 gnd.n3462 gnd.n3461 9.3005
R17259 gnd.n3460 gnd.n3459 9.3005
R17260 gnd.n3444 gnd.n3443 9.3005
R17261 gnd.n3417 gnd.n3416 9.3005
R17262 gnd.n3438 gnd.n3437 9.3005
R17263 gnd.n3436 gnd.n3435 9.3005
R17264 gnd.n3421 gnd.n3420 9.3005
R17265 gnd.n3430 gnd.n3429 9.3005
R17266 gnd.n3428 gnd.n3427 9.3005
R17267 gnd.n3412 gnd.n3411 9.3005
R17268 gnd.n3385 gnd.n3384 9.3005
R17269 gnd.n3406 gnd.n3405 9.3005
R17270 gnd.n3404 gnd.n3403 9.3005
R17271 gnd.n3389 gnd.n3388 9.3005
R17272 gnd.n3398 gnd.n3397 9.3005
R17273 gnd.n3396 gnd.n3395 9.3005
R17274 gnd.n3380 gnd.n3379 9.3005
R17275 gnd.n3353 gnd.n3352 9.3005
R17276 gnd.n3374 gnd.n3373 9.3005
R17277 gnd.n3372 gnd.n3371 9.3005
R17278 gnd.n3357 gnd.n3356 9.3005
R17279 gnd.n3366 gnd.n3365 9.3005
R17280 gnd.n3364 gnd.n3363 9.3005
R17281 gnd.n3349 gnd.n3348 9.3005
R17282 gnd.n3322 gnd.n3321 9.3005
R17283 gnd.n3343 gnd.n3342 9.3005
R17284 gnd.n3341 gnd.n3340 9.3005
R17285 gnd.n3326 gnd.n3325 9.3005
R17286 gnd.n3335 gnd.n3334 9.3005
R17287 gnd.n3333 gnd.n3332 9.3005
R17288 gnd.n3697 gnd.n3696 9.3005
R17289 gnd.n3695 gnd.n2253 9.3005
R17290 gnd.n3694 gnd.n3693 9.3005
R17291 gnd.n3690 gnd.n2254 9.3005
R17292 gnd.n3687 gnd.n2255 9.3005
R17293 gnd.n3686 gnd.n2256 9.3005
R17294 gnd.n3683 gnd.n2257 9.3005
R17295 gnd.n3682 gnd.n2258 9.3005
R17296 gnd.n3679 gnd.n2259 9.3005
R17297 gnd.n3678 gnd.n2260 9.3005
R17298 gnd.n3675 gnd.n2261 9.3005
R17299 gnd.n3674 gnd.n2262 9.3005
R17300 gnd.n3671 gnd.n2263 9.3005
R17301 gnd.n3670 gnd.n2264 9.3005
R17302 gnd.n3667 gnd.n3666 9.3005
R17303 gnd.n3665 gnd.n2265 9.3005
R17304 gnd.n3698 gnd.n2252 9.3005
R17305 gnd.n2939 gnd.n2938 9.3005
R17306 gnd.n2643 gnd.n2642 9.3005
R17307 gnd.n2966 gnd.n2965 9.3005
R17308 gnd.n2967 gnd.n2641 9.3005
R17309 gnd.n2971 gnd.n2968 9.3005
R17310 gnd.n2970 gnd.n2969 9.3005
R17311 gnd.n2615 gnd.n2614 9.3005
R17312 gnd.n2996 gnd.n2995 9.3005
R17313 gnd.n2997 gnd.n2613 9.3005
R17314 gnd.n2999 gnd.n2998 9.3005
R17315 gnd.n2593 gnd.n2592 9.3005
R17316 gnd.n3027 gnd.n3026 9.3005
R17317 gnd.n3028 gnd.n2591 9.3005
R17318 gnd.n3036 gnd.n3029 9.3005
R17319 gnd.n3035 gnd.n3030 9.3005
R17320 gnd.n3034 gnd.n3032 9.3005
R17321 gnd.n3031 gnd.n2540 9.3005
R17322 gnd.n3084 gnd.n2541 9.3005
R17323 gnd.n3083 gnd.n2542 9.3005
R17324 gnd.n3082 gnd.n2543 9.3005
R17325 gnd.n2562 gnd.n2544 9.3005
R17326 gnd.n2564 gnd.n2563 9.3005
R17327 gnd.n2450 gnd.n2449 9.3005
R17328 gnd.n3122 gnd.n3121 9.3005
R17329 gnd.n3123 gnd.n2448 9.3005
R17330 gnd.n3127 gnd.n3124 9.3005
R17331 gnd.n3126 gnd.n3125 9.3005
R17332 gnd.n2423 gnd.n2422 9.3005
R17333 gnd.n3162 gnd.n3161 9.3005
R17334 gnd.n3163 gnd.n2421 9.3005
R17335 gnd.n3167 gnd.n3164 9.3005
R17336 gnd.n3166 gnd.n3165 9.3005
R17337 gnd.n2396 gnd.n2395 9.3005
R17338 gnd.n3207 gnd.n3206 9.3005
R17339 gnd.n3208 gnd.n2394 9.3005
R17340 gnd.n3212 gnd.n3209 9.3005
R17341 gnd.n3211 gnd.n3210 9.3005
R17342 gnd.n2368 gnd.n2367 9.3005
R17343 gnd.n3247 gnd.n3246 9.3005
R17344 gnd.n3248 gnd.n2366 9.3005
R17345 gnd.n3252 gnd.n3249 9.3005
R17346 gnd.n3251 gnd.n3250 9.3005
R17347 gnd.n2341 gnd.n2340 9.3005
R17348 gnd.n3296 gnd.n3295 9.3005
R17349 gnd.n3297 gnd.n2339 9.3005
R17350 gnd.n3301 gnd.n3298 9.3005
R17351 gnd.n3300 gnd.n3299 9.3005
R17352 gnd.n2314 gnd.n2313 9.3005
R17353 gnd.n3590 gnd.n3589 9.3005
R17354 gnd.n3591 gnd.n2312 9.3005
R17355 gnd.n3597 gnd.n3592 9.3005
R17356 gnd.n3596 gnd.n3593 9.3005
R17357 gnd.n3595 gnd.n3594 9.3005
R17358 gnd.n2940 gnd.n2937 9.3005
R17359 gnd.n2722 gnd.n2681 9.3005
R17360 gnd.n2717 gnd.n2716 9.3005
R17361 gnd.n2715 gnd.n2682 9.3005
R17362 gnd.n2714 gnd.n2713 9.3005
R17363 gnd.n2710 gnd.n2683 9.3005
R17364 gnd.n2707 gnd.n2706 9.3005
R17365 gnd.n2705 gnd.n2684 9.3005
R17366 gnd.n2704 gnd.n2703 9.3005
R17367 gnd.n2700 gnd.n2685 9.3005
R17368 gnd.n2697 gnd.n2696 9.3005
R17369 gnd.n2695 gnd.n2686 9.3005
R17370 gnd.n2694 gnd.n2693 9.3005
R17371 gnd.n2690 gnd.n2688 9.3005
R17372 gnd.n2687 gnd.n2667 9.3005
R17373 gnd.n2934 gnd.n2666 9.3005
R17374 gnd.n2936 gnd.n2935 9.3005
R17375 gnd.n2724 gnd.n2723 9.3005
R17376 gnd.n2947 gnd.n2653 9.3005
R17377 gnd.n2954 gnd.n2654 9.3005
R17378 gnd.n2956 gnd.n2955 9.3005
R17379 gnd.n2957 gnd.n2634 9.3005
R17380 gnd.n2976 gnd.n2975 9.3005
R17381 gnd.n2978 gnd.n2626 9.3005
R17382 gnd.n2985 gnd.n2628 9.3005
R17383 gnd.n2986 gnd.n2623 9.3005
R17384 gnd.n2988 gnd.n2987 9.3005
R17385 gnd.n2624 gnd.n2609 9.3005
R17386 gnd.n3004 gnd.n2607 9.3005
R17387 gnd.n3008 gnd.n3007 9.3005
R17388 gnd.n3006 gnd.n2583 9.3005
R17389 gnd.n3043 gnd.n2582 9.3005
R17390 gnd.n3046 gnd.n3045 9.3005
R17391 gnd.n2579 gnd.n2578 9.3005
R17392 gnd.n3052 gnd.n2580 9.3005
R17393 gnd.n3054 gnd.n3053 9.3005
R17394 gnd.n3056 gnd.n2577 9.3005
R17395 gnd.n3059 gnd.n3058 9.3005
R17396 gnd.n3062 gnd.n3060 9.3005
R17397 gnd.n3064 gnd.n3063 9.3005
R17398 gnd.n3070 gnd.n3065 9.3005
R17399 gnd.n3069 gnd.n3068 9.3005
R17400 gnd.n2441 gnd.n2440 9.3005
R17401 gnd.n3136 gnd.n3135 9.3005
R17402 gnd.n3137 gnd.n2434 9.3005
R17403 gnd.n3145 gnd.n2433 9.3005
R17404 gnd.n3148 gnd.n3147 9.3005
R17405 gnd.n3150 gnd.n3149 9.3005
R17406 gnd.n3153 gnd.n2416 9.3005
R17407 gnd.n3151 gnd.n2414 9.3005
R17408 gnd.n3173 gnd.n2412 9.3005
R17409 gnd.n3175 gnd.n3174 9.3005
R17410 gnd.n2386 gnd.n2385 9.3005
R17411 gnd.n3221 gnd.n3220 9.3005
R17412 gnd.n3222 gnd.n2379 9.3005
R17413 gnd.n3230 gnd.n2378 9.3005
R17414 gnd.n3233 gnd.n3232 9.3005
R17415 gnd.n3235 gnd.n3234 9.3005
R17416 gnd.n3238 gnd.n2361 9.3005
R17417 gnd.n3236 gnd.n2359 9.3005
R17418 gnd.n3258 gnd.n2357 9.3005
R17419 gnd.n3260 gnd.n3259 9.3005
R17420 gnd.n2332 gnd.n2331 9.3005
R17421 gnd.n3310 gnd.n3309 9.3005
R17422 gnd.n3311 gnd.n2325 9.3005
R17423 gnd.n3319 gnd.n2324 9.3005
R17424 gnd.n3578 gnd.n3577 9.3005
R17425 gnd.n3580 gnd.n3579 9.3005
R17426 gnd.n3581 gnd.n2305 9.3005
R17427 gnd.n3605 gnd.n3604 9.3005
R17428 gnd.n2306 gnd.n2268 9.3005
R17429 gnd.n2945 gnd.n2944 9.3005
R17430 gnd.n3661 gnd.n2269 9.3005
R17431 gnd.n3660 gnd.n2271 9.3005
R17432 gnd.n3657 gnd.n2272 9.3005
R17433 gnd.n3656 gnd.n2273 9.3005
R17434 gnd.n3653 gnd.n2274 9.3005
R17435 gnd.n3652 gnd.n2275 9.3005
R17436 gnd.n3649 gnd.n2276 9.3005
R17437 gnd.n3648 gnd.n2277 9.3005
R17438 gnd.n3645 gnd.n2278 9.3005
R17439 gnd.n3644 gnd.n2279 9.3005
R17440 gnd.n3641 gnd.n2280 9.3005
R17441 gnd.n3640 gnd.n2281 9.3005
R17442 gnd.n3637 gnd.n2282 9.3005
R17443 gnd.n3636 gnd.n2283 9.3005
R17444 gnd.n3633 gnd.n2284 9.3005
R17445 gnd.n3632 gnd.n2285 9.3005
R17446 gnd.n3629 gnd.n2286 9.3005
R17447 gnd.n3628 gnd.n2287 9.3005
R17448 gnd.n3625 gnd.n2288 9.3005
R17449 gnd.n3624 gnd.n2289 9.3005
R17450 gnd.n3621 gnd.n2290 9.3005
R17451 gnd.n3620 gnd.n2291 9.3005
R17452 gnd.n3617 gnd.n2295 9.3005
R17453 gnd.n3616 gnd.n2296 9.3005
R17454 gnd.n3613 gnd.n2297 9.3005
R17455 gnd.n3612 gnd.n2298 9.3005
R17456 gnd.n3663 gnd.n3662 9.3005
R17457 gnd.n3114 gnd.n3098 9.3005
R17458 gnd.n3113 gnd.n3099 9.3005
R17459 gnd.n3112 gnd.n3100 9.3005
R17460 gnd.n3110 gnd.n3101 9.3005
R17461 gnd.n3109 gnd.n3102 9.3005
R17462 gnd.n3107 gnd.n3103 9.3005
R17463 gnd.n3106 gnd.n3104 9.3005
R17464 gnd.n2404 gnd.n2403 9.3005
R17465 gnd.n3183 gnd.n3182 9.3005
R17466 gnd.n3184 gnd.n2402 9.3005
R17467 gnd.n3201 gnd.n3185 9.3005
R17468 gnd.n3200 gnd.n3186 9.3005
R17469 gnd.n3199 gnd.n3187 9.3005
R17470 gnd.n3197 gnd.n3188 9.3005
R17471 gnd.n3196 gnd.n3189 9.3005
R17472 gnd.n3194 gnd.n3190 9.3005
R17473 gnd.n3193 gnd.n3191 9.3005
R17474 gnd.n2348 gnd.n2347 9.3005
R17475 gnd.n3268 gnd.n3267 9.3005
R17476 gnd.n3269 gnd.n2346 9.3005
R17477 gnd.n3290 gnd.n3270 9.3005
R17478 gnd.n3289 gnd.n3271 9.3005
R17479 gnd.n3288 gnd.n3272 9.3005
R17480 gnd.n3285 gnd.n3273 9.3005
R17481 gnd.n3284 gnd.n3274 9.3005
R17482 gnd.n3282 gnd.n3275 9.3005
R17483 gnd.n3281 gnd.n3276 9.3005
R17484 gnd.n3279 gnd.n3278 9.3005
R17485 gnd.n3277 gnd.n2300 9.3005
R17486 gnd.n2855 gnd.n2854 9.3005
R17487 gnd.n2745 gnd.n2744 9.3005
R17488 gnd.n2869 gnd.n2868 9.3005
R17489 gnd.n2870 gnd.n2743 9.3005
R17490 gnd.n2872 gnd.n2871 9.3005
R17491 gnd.n2733 gnd.n2732 9.3005
R17492 gnd.n2885 gnd.n2884 9.3005
R17493 gnd.n2886 gnd.n2731 9.3005
R17494 gnd.n2918 gnd.n2887 9.3005
R17495 gnd.n2917 gnd.n2888 9.3005
R17496 gnd.n2916 gnd.n2889 9.3005
R17497 gnd.n2915 gnd.n2890 9.3005
R17498 gnd.n2912 gnd.n2891 9.3005
R17499 gnd.n2911 gnd.n2892 9.3005
R17500 gnd.n2910 gnd.n2893 9.3005
R17501 gnd.n2908 gnd.n2894 9.3005
R17502 gnd.n2907 gnd.n2895 9.3005
R17503 gnd.n2904 gnd.n2896 9.3005
R17504 gnd.n2903 gnd.n2897 9.3005
R17505 gnd.n2902 gnd.n2898 9.3005
R17506 gnd.n2900 gnd.n2899 9.3005
R17507 gnd.n2599 gnd.n2598 9.3005
R17508 gnd.n3016 gnd.n3015 9.3005
R17509 gnd.n3017 gnd.n2597 9.3005
R17510 gnd.n3021 gnd.n3018 9.3005
R17511 gnd.n3020 gnd.n3019 9.3005
R17512 gnd.n2521 gnd.n2520 9.3005
R17513 gnd.n3096 gnd.n3095 9.3005
R17514 gnd.n2853 gnd.n2754 9.3005
R17515 gnd.n2756 gnd.n2755 9.3005
R17516 gnd.n2800 gnd.n2798 9.3005
R17517 gnd.n2801 gnd.n2797 9.3005
R17518 gnd.n2804 gnd.n2793 9.3005
R17519 gnd.n2805 gnd.n2792 9.3005
R17520 gnd.n2808 gnd.n2791 9.3005
R17521 gnd.n2809 gnd.n2790 9.3005
R17522 gnd.n2812 gnd.n2789 9.3005
R17523 gnd.n2813 gnd.n2788 9.3005
R17524 gnd.n2816 gnd.n2787 9.3005
R17525 gnd.n2817 gnd.n2786 9.3005
R17526 gnd.n2820 gnd.n2785 9.3005
R17527 gnd.n2821 gnd.n2784 9.3005
R17528 gnd.n2824 gnd.n2783 9.3005
R17529 gnd.n2825 gnd.n2782 9.3005
R17530 gnd.n2828 gnd.n2781 9.3005
R17531 gnd.n2829 gnd.n2780 9.3005
R17532 gnd.n2832 gnd.n2779 9.3005
R17533 gnd.n2833 gnd.n2778 9.3005
R17534 gnd.n2836 gnd.n2777 9.3005
R17535 gnd.n2837 gnd.n2776 9.3005
R17536 gnd.n2840 gnd.n2775 9.3005
R17537 gnd.n2842 gnd.n2774 9.3005
R17538 gnd.n2843 gnd.n2773 9.3005
R17539 gnd.n2844 gnd.n2772 9.3005
R17540 gnd.n2845 gnd.n2771 9.3005
R17541 gnd.n2852 gnd.n2851 9.3005
R17542 gnd.n2861 gnd.n2860 9.3005
R17543 gnd.n2862 gnd.n2748 9.3005
R17544 gnd.n2864 gnd.n2863 9.3005
R17545 gnd.n2739 gnd.n2738 9.3005
R17546 gnd.n2877 gnd.n2876 9.3005
R17547 gnd.n2878 gnd.n2737 9.3005
R17548 gnd.n2880 gnd.n2879 9.3005
R17549 gnd.n2726 gnd.n2725 9.3005
R17550 gnd.n2923 gnd.n2922 9.3005
R17551 gnd.n2924 gnd.n2680 9.3005
R17552 gnd.n2928 gnd.n2926 9.3005
R17553 gnd.n2927 gnd.n2659 9.3005
R17554 gnd.n2946 gnd.n2658 9.3005
R17555 gnd.n2949 gnd.n2948 9.3005
R17556 gnd.n2652 gnd.n2651 9.3005
R17557 gnd.n2960 gnd.n2958 9.3005
R17558 gnd.n2959 gnd.n2633 9.3005
R17559 gnd.n2977 gnd.n2632 9.3005
R17560 gnd.n2980 gnd.n2979 9.3005
R17561 gnd.n2627 gnd.n2622 9.3005
R17562 gnd.n2990 gnd.n2989 9.3005
R17563 gnd.n2625 gnd.n2605 9.3005
R17564 gnd.n3011 gnd.n2606 9.3005
R17565 gnd.n3010 gnd.n3009 9.3005
R17566 gnd.n2608 gnd.n2584 9.3005
R17567 gnd.n3042 gnd.n3041 9.3005
R17568 gnd.n3044 gnd.n2529 9.3005
R17569 gnd.n3091 gnd.n2530 9.3005
R17570 gnd.n3090 gnd.n2531 9.3005
R17571 gnd.n3089 gnd.n2532 9.3005
R17572 gnd.n3055 gnd.n2533 9.3005
R17573 gnd.n3057 gnd.n2551 9.3005
R17574 gnd.n3077 gnd.n2552 9.3005
R17575 gnd.n3076 gnd.n2553 9.3005
R17576 gnd.n3075 gnd.n2554 9.3005
R17577 gnd.n3066 gnd.n2555 9.3005
R17578 gnd.n3067 gnd.n2442 9.3005
R17579 gnd.n3133 gnd.n3132 9.3005
R17580 gnd.n3134 gnd.n2435 9.3005
R17581 gnd.n3144 gnd.n3143 9.3005
R17582 gnd.n3146 gnd.n2431 9.3005
R17583 gnd.n3156 gnd.n2432 9.3005
R17584 gnd.n3155 gnd.n3154 9.3005
R17585 gnd.n3152 gnd.n2410 9.3005
R17586 gnd.n3178 gnd.n2411 9.3005
R17587 gnd.n3177 gnd.n3176 9.3005
R17588 gnd.n2413 gnd.n2387 9.3005
R17589 gnd.n3218 gnd.n3217 9.3005
R17590 gnd.n3219 gnd.n2380 9.3005
R17591 gnd.n3229 gnd.n3228 9.3005
R17592 gnd.n3231 gnd.n2376 9.3005
R17593 gnd.n3241 gnd.n2377 9.3005
R17594 gnd.n3240 gnd.n3239 9.3005
R17595 gnd.n3237 gnd.n2355 9.3005
R17596 gnd.n3263 gnd.n2356 9.3005
R17597 gnd.n3262 gnd.n3261 9.3005
R17598 gnd.n2358 gnd.n2333 9.3005
R17599 gnd.n3307 gnd.n3306 9.3005
R17600 gnd.n3308 gnd.n2326 9.3005
R17601 gnd.n3318 gnd.n3317 9.3005
R17602 gnd.n3576 gnd.n2322 9.3005
R17603 gnd.n3584 gnd.n2323 9.3005
R17604 gnd.n3583 gnd.n3582 9.3005
R17605 gnd.n2304 gnd.n2303 9.3005
R17606 gnd.n3607 gnd.n3606 9.3005
R17607 gnd.n2750 gnd.n2749 9.3005
R17608 gnd.n3834 gnd.n3710 9.3005
R17609 gnd.n3836 gnd.n3835 9.3005
R17610 gnd.n3833 gnd.n3712 9.3005
R17611 gnd.n3832 gnd.n3831 9.3005
R17612 gnd.n3714 gnd.n3713 9.3005
R17613 gnd.n3825 gnd.n3824 9.3005
R17614 gnd.n3823 gnd.n3716 9.3005
R17615 gnd.n3822 gnd.n3821 9.3005
R17616 gnd.n3718 gnd.n3717 9.3005
R17617 gnd.n3815 gnd.n3814 9.3005
R17618 gnd.n3813 gnd.n3720 9.3005
R17619 gnd.n3812 gnd.n3811 9.3005
R17620 gnd.n3722 gnd.n3721 9.3005
R17621 gnd.n3805 gnd.n3804 9.3005
R17622 gnd.n3803 gnd.n3724 9.3005
R17623 gnd.n3802 gnd.n3801 9.3005
R17624 gnd.n3726 gnd.n3725 9.3005
R17625 gnd.n3795 gnd.n3794 9.3005
R17626 gnd.n3793 gnd.n3728 9.3005
R17627 gnd.n3792 gnd.n3791 9.3005
R17628 gnd.n3730 gnd.n3729 9.3005
R17629 gnd.n3785 gnd.n3784 9.3005
R17630 gnd.n3783 gnd.n3735 9.3005
R17631 gnd.n3782 gnd.n3781 9.3005
R17632 gnd.n3737 gnd.n3736 9.3005
R17633 gnd.n3775 gnd.n3774 9.3005
R17634 gnd.n3773 gnd.n3739 9.3005
R17635 gnd.n3772 gnd.n3771 9.3005
R17636 gnd.n3741 gnd.n3740 9.3005
R17637 gnd.n3765 gnd.n3764 9.3005
R17638 gnd.n3763 gnd.n3743 9.3005
R17639 gnd.n3762 gnd.n3761 9.3005
R17640 gnd.n3745 gnd.n3744 9.3005
R17641 gnd.n3755 gnd.n3754 9.3005
R17642 gnd.n3753 gnd.n3747 9.3005
R17643 gnd.n3752 gnd.n3751 9.3005
R17644 gnd.n3748 gnd.n2225 9.3005
R17645 gnd.n3709 gnd.n3706 9.3005
R17646 gnd.n3844 gnd.n3843 9.3005
R17647 gnd.n4196 gnd.n2224 9.3005
R17648 gnd.n4198 gnd.n4197 9.3005
R17649 gnd.n2211 gnd.n2210 9.3005
R17650 gnd.n4211 gnd.n4210 9.3005
R17651 gnd.n4212 gnd.n2209 9.3005
R17652 gnd.n4214 gnd.n4213 9.3005
R17653 gnd.n2194 gnd.n2193 9.3005
R17654 gnd.n4227 gnd.n4226 9.3005
R17655 gnd.n4228 gnd.n2192 9.3005
R17656 gnd.n4230 gnd.n4229 9.3005
R17657 gnd.n2179 gnd.n2178 9.3005
R17658 gnd.n4243 gnd.n4242 9.3005
R17659 gnd.n4244 gnd.n2177 9.3005
R17660 gnd.n4246 gnd.n4245 9.3005
R17661 gnd.n2162 gnd.n2161 9.3005
R17662 gnd.n4259 gnd.n4258 9.3005
R17663 gnd.n4260 gnd.n2160 9.3005
R17664 gnd.n4262 gnd.n4261 9.3005
R17665 gnd.n2147 gnd.n2146 9.3005
R17666 gnd.n4275 gnd.n4274 9.3005
R17667 gnd.n4276 gnd.n2145 9.3005
R17668 gnd.n4278 gnd.n4277 9.3005
R17669 gnd.n2130 gnd.n2129 9.3005
R17670 gnd.n4291 gnd.n4290 9.3005
R17671 gnd.n4292 gnd.n2128 9.3005
R17672 gnd.n4294 gnd.n4293 9.3005
R17673 gnd.n2115 gnd.n2114 9.3005
R17674 gnd.n4195 gnd.n4194 9.3005
R17675 gnd.n4307 gnd.n4306 9.3005
R17676 gnd.n4308 gnd.n2113 9.3005
R17677 gnd.n4310 gnd.n4309 9.3005
R17678 gnd.n2097 gnd.n2096 9.3005
R17679 gnd.n4323 gnd.n4322 9.3005
R17680 gnd.n4324 gnd.n2095 9.3005
R17681 gnd.n4326 gnd.n4325 9.3005
R17682 gnd.n2082 gnd.n2081 9.3005
R17683 gnd.n4339 gnd.n4338 9.3005
R17684 gnd.n4340 gnd.n2080 9.3005
R17685 gnd.n4342 gnd.n4341 9.3005
R17686 gnd.n2065 gnd.n2064 9.3005
R17687 gnd.n4355 gnd.n4354 9.3005
R17688 gnd.n4356 gnd.n2063 9.3005
R17689 gnd.n4358 gnd.n4357 9.3005
R17690 gnd.n2050 gnd.n2049 9.3005
R17691 gnd.n4371 gnd.n4370 9.3005
R17692 gnd.n4372 gnd.n2048 9.3005
R17693 gnd.n4374 gnd.n4373 9.3005
R17694 gnd.n2033 gnd.n2032 9.3005
R17695 gnd.n4387 gnd.n4386 9.3005
R17696 gnd.n4388 gnd.n2031 9.3005
R17697 gnd.n4390 gnd.n4389 9.3005
R17698 gnd.n2017 gnd.n2016 9.3005
R17699 gnd.n4416 gnd.n4415 9.3005
R17700 gnd.n4417 gnd.n2015 9.3005
R17701 gnd.n4422 gnd.n4418 9.3005
R17702 gnd.n4421 gnd.n4420 9.3005
R17703 gnd.n4419 gnd.n1062 9.3005
R17704 gnd.n6076 gnd.n1063 9.3005
R17705 gnd.n6075 gnd.n1064 9.3005
R17706 gnd.n6074 gnd.n1065 9.3005
R17707 gnd.n1085 gnd.n1066 9.3005
R17708 gnd.n6064 gnd.n1086 9.3005
R17709 gnd.n6063 gnd.n1087 9.3005
R17710 gnd.n6062 gnd.n1088 9.3005
R17711 gnd.n1914 gnd.n1089 9.3005
R17712 gnd.n1900 gnd.n1896 9.3005
R17713 gnd.n1932 gnd.n1929 9.3005
R17714 gnd.n1933 gnd.n1928 9.3005
R17715 gnd.n1936 gnd.n1927 9.3005
R17716 gnd.n1937 gnd.n1926 9.3005
R17717 gnd.n1940 gnd.n1925 9.3005
R17718 gnd.n1941 gnd.n1924 9.3005
R17719 gnd.n1944 gnd.n1923 9.3005
R17720 gnd.n1945 gnd.n1922 9.3005
R17721 gnd.n1948 gnd.n1921 9.3005
R17722 gnd.n1949 gnd.n1920 9.3005
R17723 gnd.n1952 gnd.n1919 9.3005
R17724 gnd.n1953 gnd.n1918 9.3005
R17725 gnd.n1956 gnd.n1917 9.3005
R17726 gnd.n1957 gnd.n1916 9.3005
R17727 gnd.n1958 gnd.n1915 9.3005
R17728 gnd.n4825 gnd.n4824 9.3005
R17729 gnd.n1902 gnd.n1901 9.3005
R17730 gnd.n1963 gnd.n1961 9.3005
R17731 gnd.n4817 gnd.n1964 9.3005
R17732 gnd.n4816 gnd.n1965 9.3005
R17733 gnd.n4815 gnd.n1966 9.3005
R17734 gnd.n1970 gnd.n1967 9.3005
R17735 gnd.n4810 gnd.n1971 9.3005
R17736 gnd.n4809 gnd.n1972 9.3005
R17737 gnd.n4808 gnd.n1973 9.3005
R17738 gnd.n1977 gnd.n1974 9.3005
R17739 gnd.n4803 gnd.n1978 9.3005
R17740 gnd.n4802 gnd.n1979 9.3005
R17741 gnd.n4801 gnd.n1980 9.3005
R17742 gnd.n1984 gnd.n1981 9.3005
R17743 gnd.n4796 gnd.n1985 9.3005
R17744 gnd.n4795 gnd.n1986 9.3005
R17745 gnd.n4794 gnd.n1987 9.3005
R17746 gnd.n1993 gnd.n1990 9.3005
R17747 gnd.n4789 gnd.n4788 9.3005
R17748 gnd.n4826 gnd.n1895 9.3005
R17749 gnd.n3983 gnd.n3982 9.3005
R17750 gnd.n3981 gnd.n3705 9.3005
R17751 gnd.n3980 gnd.n3979 9.3005
R17752 gnd.n3977 gnd.n3846 9.3005
R17753 gnd.n3976 gnd.n3847 9.3005
R17754 gnd.n3974 gnd.n3848 9.3005
R17755 gnd.n3973 gnd.n3849 9.3005
R17756 gnd.n3971 gnd.n3850 9.3005
R17757 gnd.n3970 gnd.n3851 9.3005
R17758 gnd.n3968 gnd.n3852 9.3005
R17759 gnd.n3967 gnd.n3853 9.3005
R17760 gnd.n3965 gnd.n3854 9.3005
R17761 gnd.n3964 gnd.n3855 9.3005
R17762 gnd.n3962 gnd.n3856 9.3005
R17763 gnd.n3961 gnd.n3857 9.3005
R17764 gnd.n3959 gnd.n3858 9.3005
R17765 gnd.n3958 gnd.n3859 9.3005
R17766 gnd.n3956 gnd.n3860 9.3005
R17767 gnd.n3955 gnd.n3861 9.3005
R17768 gnd.n3953 gnd.n3862 9.3005
R17769 gnd.n3952 gnd.n3863 9.3005
R17770 gnd.n3950 gnd.n3864 9.3005
R17771 gnd.n3949 gnd.n3865 9.3005
R17772 gnd.n3947 gnd.n3866 9.3005
R17773 gnd.n3946 gnd.n3867 9.3005
R17774 gnd.n3944 gnd.n3868 9.3005
R17775 gnd.n3943 gnd.n3869 9.3005
R17776 gnd.n3941 gnd.n3870 9.3005
R17777 gnd.n3940 gnd.n3871 9.3005
R17778 gnd.n3938 gnd.n3872 9.3005
R17779 gnd.n3937 gnd.n3873 9.3005
R17780 gnd.n3935 gnd.n2105 9.3005
R17781 gnd.n3934 gnd.n3874 9.3005
R17782 gnd.n3932 gnd.n3875 9.3005
R17783 gnd.n3931 gnd.n3876 9.3005
R17784 gnd.n3929 gnd.n3877 9.3005
R17785 gnd.n3928 gnd.n3878 9.3005
R17786 gnd.n3926 gnd.n3879 9.3005
R17787 gnd.n3925 gnd.n3880 9.3005
R17788 gnd.n3923 gnd.n3881 9.3005
R17789 gnd.n3922 gnd.n3882 9.3005
R17790 gnd.n3920 gnd.n3883 9.3005
R17791 gnd.n3919 gnd.n3884 9.3005
R17792 gnd.n3917 gnd.n3885 9.3005
R17793 gnd.n3916 gnd.n3886 9.3005
R17794 gnd.n3914 gnd.n3887 9.3005
R17795 gnd.n3913 gnd.n3888 9.3005
R17796 gnd.n3911 gnd.n3889 9.3005
R17797 gnd.n3910 gnd.n3890 9.3005
R17798 gnd.n3908 gnd.n3891 9.3005
R17799 gnd.n3907 gnd.n3892 9.3005
R17800 gnd.n3905 gnd.n3893 9.3005
R17801 gnd.n3904 gnd.n3894 9.3005
R17802 gnd.n3902 gnd.n3895 9.3005
R17803 gnd.n3901 gnd.n3896 9.3005
R17804 gnd.n3898 gnd.n3897 9.3005
R17805 gnd.n2003 gnd.n2002 9.3005
R17806 gnd.n4437 gnd.n4436 9.3005
R17807 gnd.n4438 gnd.n2001 9.3005
R17808 gnd.n4441 gnd.n4440 9.3005
R17809 gnd.n4439 gnd.n1995 9.3005
R17810 gnd.n4784 gnd.n1996 9.3005
R17811 gnd.n4785 gnd.n1994 9.3005
R17812 gnd.n4787 gnd.n4786 9.3005
R17813 gnd.n3845 gnd.n3704 9.3005
R17814 gnd.n4098 gnd.n4097 9.3005
R17815 gnd.n4145 gnd.n4013 9.3005
R17816 gnd.n4143 gnd.n4014 9.3005
R17817 gnd.n4142 gnd.n4015 9.3005
R17818 gnd.n4140 gnd.n4016 9.3005
R17819 gnd.n4139 gnd.n4017 9.3005
R17820 gnd.n4137 gnd.n4018 9.3005
R17821 gnd.n4136 gnd.n4019 9.3005
R17822 gnd.n4134 gnd.n4020 9.3005
R17823 gnd.n4133 gnd.n4021 9.3005
R17824 gnd.n4131 gnd.n4022 9.3005
R17825 gnd.n4130 gnd.n4023 9.3005
R17826 gnd.n4128 gnd.n4024 9.3005
R17827 gnd.n4127 gnd.n4025 9.3005
R17828 gnd.n4125 gnd.n4026 9.3005
R17829 gnd.n4124 gnd.n4027 9.3005
R17830 gnd.n4122 gnd.n4028 9.3005
R17831 gnd.n4121 gnd.n4029 9.3005
R17832 gnd.n4119 gnd.n4030 9.3005
R17833 gnd.n4118 gnd.n4031 9.3005
R17834 gnd.n4116 gnd.n4032 9.3005
R17835 gnd.n4115 gnd.n4033 9.3005
R17836 gnd.n4113 gnd.n4034 9.3005
R17837 gnd.n4112 gnd.n4035 9.3005
R17838 gnd.n4110 gnd.n4036 9.3005
R17839 gnd.n4109 gnd.n4037 9.3005
R17840 gnd.n4107 gnd.n4038 9.3005
R17841 gnd.n4106 gnd.n4039 9.3005
R17842 gnd.n4104 gnd.n4040 9.3005
R17843 gnd.n4103 gnd.n4041 9.3005
R17844 gnd.n4101 gnd.n4042 9.3005
R17845 gnd.n4100 gnd.n4043 9.3005
R17846 gnd.n4147 gnd.n4146 9.3005
R17847 gnd.n4155 gnd.n4154 9.3005
R17848 gnd.n4156 gnd.n4009 9.3005
R17849 gnd.n4008 gnd.n4006 9.3005
R17850 gnd.n4162 gnd.n4005 9.3005
R17851 gnd.n4163 gnd.n4004 9.3005
R17852 gnd.n4164 gnd.n4003 9.3005
R17853 gnd.n4002 gnd.n4000 9.3005
R17854 gnd.n4170 gnd.n3999 9.3005
R17855 gnd.n4171 gnd.n3998 9.3005
R17856 gnd.n4172 gnd.n3997 9.3005
R17857 gnd.n3996 gnd.n3994 9.3005
R17858 gnd.n4178 gnd.n3993 9.3005
R17859 gnd.n4179 gnd.n3992 9.3005
R17860 gnd.n4180 gnd.n3991 9.3005
R17861 gnd.n3990 gnd.n3988 9.3005
R17862 gnd.n4186 gnd.n3987 9.3005
R17863 gnd.n4188 gnd.n4187 9.3005
R17864 gnd.n4153 gnd.n4012 9.3005
R17865 gnd.n4152 gnd.n4151 9.3005
R17866 gnd.n2219 gnd.n2218 9.3005
R17867 gnd.n4203 gnd.n4202 9.3005
R17868 gnd.n4204 gnd.n2217 9.3005
R17869 gnd.n4206 gnd.n4205 9.3005
R17870 gnd.n2203 gnd.n2202 9.3005
R17871 gnd.n4219 gnd.n4218 9.3005
R17872 gnd.n4220 gnd.n2201 9.3005
R17873 gnd.n4222 gnd.n4221 9.3005
R17874 gnd.n2187 gnd.n2186 9.3005
R17875 gnd.n4235 gnd.n4234 9.3005
R17876 gnd.n4236 gnd.n2185 9.3005
R17877 gnd.n4238 gnd.n4237 9.3005
R17878 gnd.n2171 gnd.n2170 9.3005
R17879 gnd.n4251 gnd.n4250 9.3005
R17880 gnd.n4252 gnd.n2169 9.3005
R17881 gnd.n4254 gnd.n4253 9.3005
R17882 gnd.n2155 gnd.n2154 9.3005
R17883 gnd.n4267 gnd.n4266 9.3005
R17884 gnd.n4268 gnd.n2153 9.3005
R17885 gnd.n4270 gnd.n4269 9.3005
R17886 gnd.n2139 gnd.n2138 9.3005
R17887 gnd.n4283 gnd.n4282 9.3005
R17888 gnd.n4284 gnd.n2137 9.3005
R17889 gnd.n4286 gnd.n4285 9.3005
R17890 gnd.n2123 gnd.n2122 9.3005
R17891 gnd.n4299 gnd.n4298 9.3005
R17892 gnd.n4300 gnd.n2121 9.3005
R17893 gnd.n4302 gnd.n4301 9.3005
R17894 gnd.n2107 gnd.n2106 9.3005
R17895 gnd.n4315 gnd.n4314 9.3005
R17896 gnd.n4316 gnd.n2104 9.3005
R17897 gnd.n4318 gnd.n4317 9.3005
R17898 gnd.n2089 gnd.n2088 9.3005
R17899 gnd.n4331 gnd.n4330 9.3005
R17900 gnd.n4332 gnd.n2087 9.3005
R17901 gnd.n4334 gnd.n4333 9.3005
R17902 gnd.n2074 gnd.n2073 9.3005
R17903 gnd.n4347 gnd.n4346 9.3005
R17904 gnd.n4348 gnd.n2072 9.3005
R17905 gnd.n4350 gnd.n4349 9.3005
R17906 gnd.n2057 gnd.n2056 9.3005
R17907 gnd.n4363 gnd.n4362 9.3005
R17908 gnd.n4364 gnd.n2055 9.3005
R17909 gnd.n4366 gnd.n4365 9.3005
R17910 gnd.n2042 gnd.n2041 9.3005
R17911 gnd.n4379 gnd.n4378 9.3005
R17912 gnd.n4380 gnd.n2040 9.3005
R17913 gnd.n4382 gnd.n4381 9.3005
R17914 gnd.n2025 gnd.n2024 9.3005
R17915 gnd.n4395 gnd.n4394 9.3005
R17916 gnd.n4396 gnd.n2023 9.3005
R17917 gnd.n4411 gnd.n4397 9.3005
R17918 gnd.n4410 gnd.n4398 9.3005
R17919 gnd.n4409 gnd.n4399 9.3005
R17920 gnd.n4408 gnd.n4400 9.3005
R17921 gnd.n4405 gnd.n4401 9.3005
R17922 gnd.n4404 gnd.n4403 9.3005
R17923 gnd.n4402 gnd.n1074 9.3005
R17924 gnd.n6070 gnd.n1075 9.3005
R17925 gnd.n6069 gnd.n1076 9.3005
R17926 gnd.n6068 gnd.n1077 9.3005
R17927 gnd.n1096 gnd.n1078 9.3005
R17928 gnd.n6058 gnd.n1097 9.3005
R17929 gnd.n6057 gnd.n6056 9.3005
R17930 gnd.n4190 gnd.n4189 9.3005
R17931 gnd.n7147 gnd.n7146 9.3005
R17932 gnd.n462 gnd.n461 9.3005
R17933 gnd.n7141 gnd.n7140 9.3005
R17934 gnd.n7139 gnd.n7138 9.3005
R17935 gnd.n470 gnd.n469 9.3005
R17936 gnd.n7133 gnd.n7132 9.3005
R17937 gnd.n7131 gnd.n7130 9.3005
R17938 gnd.n478 gnd.n477 9.3005
R17939 gnd.n7125 gnd.n7124 9.3005
R17940 gnd.n7123 gnd.n7122 9.3005
R17941 gnd.n486 gnd.n485 9.3005
R17942 gnd.n7117 gnd.n7116 9.3005
R17943 gnd.n7115 gnd.n7114 9.3005
R17944 gnd.n494 gnd.n493 9.3005
R17945 gnd.n7109 gnd.n7108 9.3005
R17946 gnd.n7107 gnd.n7106 9.3005
R17947 gnd.n504 gnd.n503 9.3005
R17948 gnd.n1280 gnd.n1279 9.3005
R17949 gnd.n7149 gnd.n7148 9.3005
R17950 gnd.n7111 gnd.n7110 9.3005
R17951 gnd.n7113 gnd.n7112 9.3005
R17952 gnd.n490 gnd.n489 9.3005
R17953 gnd.n7119 gnd.n7118 9.3005
R17954 gnd.n7121 gnd.n7120 9.3005
R17955 gnd.n482 gnd.n481 9.3005
R17956 gnd.n7127 gnd.n7126 9.3005
R17957 gnd.n7129 gnd.n7128 9.3005
R17958 gnd.n474 gnd.n473 9.3005
R17959 gnd.n7135 gnd.n7134 9.3005
R17960 gnd.n7137 gnd.n7136 9.3005
R17961 gnd.n466 gnd.n465 9.3005
R17962 gnd.n7143 gnd.n7142 9.3005
R17963 gnd.n7145 gnd.n7144 9.3005
R17964 gnd.n458 gnd.n457 9.3005
R17965 gnd.n7151 gnd.n7150 9.3005
R17966 gnd.n500 gnd.n499 9.3005
R17967 gnd.n7105 gnd.n7104 9.3005
R17968 gnd.n1282 gnd.n1274 9.3005
R17969 gnd.n1284 gnd.n1283 9.3005
R17970 gnd.n1285 gnd.n1273 9.3005
R17971 gnd.n1289 gnd.n1288 9.3005
R17972 gnd.n1290 gnd.n1270 9.3005
R17973 gnd.n1292 gnd.n1291 9.3005
R17974 gnd.n1294 gnd.n1267 9.3005
R17975 gnd.n1298 gnd.n1297 9.3005
R17976 gnd.n1299 gnd.n1266 9.3005
R17977 gnd.n5888 gnd.n5887 9.3005
R17978 gnd.n4697 gnd.n4581 9.3005
R17979 gnd.n4696 gnd.n4695 9.3005
R17980 gnd.n4694 gnd.n4586 9.3005
R17981 gnd.n4693 gnd.n4692 9.3005
R17982 gnd.n4691 gnd.n4587 9.3005
R17983 gnd.n4690 gnd.n4689 9.3005
R17984 gnd.n4688 gnd.n4591 9.3005
R17985 gnd.n4687 gnd.n4686 9.3005
R17986 gnd.n4685 gnd.n4592 9.3005
R17987 gnd.n4684 gnd.n4683 9.3005
R17988 gnd.n4682 gnd.n4596 9.3005
R17989 gnd.n4681 gnd.n4680 9.3005
R17990 gnd.n4679 gnd.n4597 9.3005
R17991 gnd.n4678 gnd.n4677 9.3005
R17992 gnd.n4676 gnd.n4669 9.3005
R17993 gnd.n4675 gnd.n4674 9.3005
R17994 gnd.n1742 gnd.n1741 9.3005
R17995 gnd.n4977 gnd.n4976 9.3005
R17996 gnd.n4978 gnd.n1739 9.3005
R17997 gnd.n4981 gnd.n4980 9.3005
R17998 gnd.n4979 gnd.n1740 9.3005
R17999 gnd.n1712 gnd.n1711 9.3005
R18000 gnd.n5016 gnd.n5015 9.3005
R18001 gnd.n5017 gnd.n1709 9.3005
R18002 gnd.n5056 gnd.n5055 9.3005
R18003 gnd.n5054 gnd.n1710 9.3005
R18004 gnd.n5053 gnd.n5052 9.3005
R18005 gnd.n5051 gnd.n5018 9.3005
R18006 gnd.n5050 gnd.n5049 9.3005
R18007 gnd.n5048 gnd.n5022 9.3005
R18008 gnd.n5047 gnd.n5046 9.3005
R18009 gnd.n5045 gnd.n5023 9.3005
R18010 gnd.n5044 gnd.n5043 9.3005
R18011 gnd.n5042 gnd.n5028 9.3005
R18012 gnd.n5041 gnd.n5040 9.3005
R18013 gnd.n5039 gnd.n5029 9.3005
R18014 gnd.n5038 gnd.n5037 9.3005
R18015 gnd.n5036 gnd.n5035 9.3005
R18016 gnd.n1627 gnd.n1626 9.3005
R18017 gnd.n5194 gnd.n5193 9.3005
R18018 gnd.n5195 gnd.n1624 9.3005
R18019 gnd.n5232 gnd.n5231 9.3005
R18020 gnd.n5230 gnd.n1625 9.3005
R18021 gnd.n5229 gnd.n5228 9.3005
R18022 gnd.n5227 gnd.n5196 9.3005
R18023 gnd.n5226 gnd.n5225 9.3005
R18024 gnd.n5224 gnd.n5200 9.3005
R18025 gnd.n5223 gnd.n5222 9.3005
R18026 gnd.n5221 gnd.n5201 9.3005
R18027 gnd.n5220 gnd.n5219 9.3005
R18028 gnd.n5218 gnd.n5204 9.3005
R18029 gnd.n5217 gnd.n5216 9.3005
R18030 gnd.n5215 gnd.n5205 9.3005
R18031 gnd.n5214 gnd.n5213 9.3005
R18032 gnd.n5212 gnd.n5211 9.3005
R18033 gnd.n1540 gnd.n1539 9.3005
R18034 gnd.n5371 gnd.n5370 9.3005
R18035 gnd.n5372 gnd.n1537 9.3005
R18036 gnd.n5394 gnd.n5393 9.3005
R18037 gnd.n5392 gnd.n1538 9.3005
R18038 gnd.n5391 gnd.n5390 9.3005
R18039 gnd.n5389 gnd.n5373 9.3005
R18040 gnd.n5388 gnd.n5387 9.3005
R18041 gnd.n5386 gnd.n5377 9.3005
R18042 gnd.n5385 gnd.n5384 9.3005
R18043 gnd.n5383 gnd.n5378 9.3005
R18044 gnd.n5382 gnd.n5381 9.3005
R18045 gnd.n1475 gnd.n1474 9.3005
R18046 gnd.n5504 gnd.n5503 9.3005
R18047 gnd.n5505 gnd.n1472 9.3005
R18048 gnd.n5508 gnd.n5507 9.3005
R18049 gnd.n5506 gnd.n1473 9.3005
R18050 gnd.n1448 gnd.n1447 9.3005
R18051 gnd.n5543 gnd.n5542 9.3005
R18052 gnd.n5544 gnd.n1445 9.3005
R18053 gnd.n5576 gnd.n5575 9.3005
R18054 gnd.n5574 gnd.n1446 9.3005
R18055 gnd.n5573 gnd.n5572 9.3005
R18056 gnd.n5571 gnd.n5545 9.3005
R18057 gnd.n5570 gnd.n5569 9.3005
R18058 gnd.n5568 gnd.n5550 9.3005
R18059 gnd.n5567 gnd.n5566 9.3005
R18060 gnd.n5565 gnd.n5551 9.3005
R18061 gnd.n5564 gnd.n5563 9.3005
R18062 gnd.n5562 gnd.n5559 9.3005
R18063 gnd.n5561 gnd.n5560 9.3005
R18064 gnd.n1337 gnd.n1336 9.3005
R18065 gnd.n5822 gnd.n5821 9.3005
R18066 gnd.n5823 gnd.n1335 9.3005
R18067 gnd.n5825 gnd.n5824 9.3005
R18068 gnd.n1325 gnd.n1324 9.3005
R18069 gnd.n5842 gnd.n5841 9.3005
R18070 gnd.n5843 gnd.n1323 9.3005
R18071 gnd.n5845 gnd.n5844 9.3005
R18072 gnd.n1312 gnd.n1311 9.3005
R18073 gnd.n5862 gnd.n5861 9.3005
R18074 gnd.n5863 gnd.n1310 9.3005
R18075 gnd.n5866 gnd.n5865 9.3005
R18076 gnd.n5864 gnd.n1301 9.3005
R18077 gnd.n5884 gnd.n1300 9.3005
R18078 gnd.n5886 gnd.n5885 9.3005
R18079 gnd.n4699 gnd.n4698 9.3005
R18080 gnd.n4702 gnd.n4701 9.3005
R18081 gnd.n4703 gnd.n4572 9.3005
R18082 gnd.n4705 gnd.n4704 9.3005
R18083 gnd.n4706 gnd.n4571 9.3005
R18084 gnd.n4708 gnd.n4707 9.3005
R18085 gnd.n4709 gnd.n4566 9.3005
R18086 gnd.n4711 gnd.n4710 9.3005
R18087 gnd.n4712 gnd.n4565 9.3005
R18088 gnd.n4714 gnd.n4713 9.3005
R18089 gnd.n4700 gnd.n4580 9.3005
R18090 gnd.n4096 gnd.n4045 9.3005
R18091 gnd.n4095 gnd.n4094 9.3005
R18092 gnd.n4093 gnd.n4046 9.3005
R18093 gnd.n4092 gnd.n4091 9.3005
R18094 gnd.n4090 gnd.n4049 9.3005
R18095 gnd.n4089 gnd.n4088 9.3005
R18096 gnd.n4087 gnd.n4050 9.3005
R18097 gnd.n4086 gnd.n4085 9.3005
R18098 gnd.n4084 gnd.n4053 9.3005
R18099 gnd.n4083 gnd.n4082 9.3005
R18100 gnd.n4081 gnd.n4054 9.3005
R18101 gnd.n4080 gnd.n4079 9.3005
R18102 gnd.n4078 gnd.n4057 9.3005
R18103 gnd.n4077 gnd.n4076 9.3005
R18104 gnd.n4075 gnd.n4058 9.3005
R18105 gnd.n4074 gnd.n4073 9.3005
R18106 gnd.n4072 gnd.n4061 9.3005
R18107 gnd.n4071 gnd.n4070 9.3005
R18108 gnd.n4069 gnd.n4062 9.3005
R18109 gnd.n4068 gnd.n4067 9.3005
R18110 gnd.n4066 gnd.n4064 9.3005
R18111 gnd.n4065 gnd.n2009 9.3005
R18112 gnd.n2007 gnd.n2006 9.3005
R18113 gnd.n4429 gnd.n4428 9.3005
R18114 gnd.n4430 gnd.n2005 9.3005
R18115 gnd.n4432 gnd.n4431 9.3005
R18116 gnd.n2000 gnd.n1999 9.3005
R18117 gnd.n4446 gnd.n4445 9.3005
R18118 gnd.n4447 gnd.n1997 9.3005
R18119 gnd.n4780 gnd.n4779 9.3005
R18120 gnd.n4778 gnd.n1998 9.3005
R18121 gnd.n4777 gnd.n4776 9.3005
R18122 gnd.n4716 gnd.n4715 9.3005
R18123 gnd.n4717 gnd.n4562 9.3005
R18124 gnd.n4721 gnd.n4720 9.3005
R18125 gnd.n4723 gnd.n4722 9.3005
R18126 gnd.n4546 gnd.n4545 9.3005
R18127 gnd.n4729 gnd.n4728 9.3005
R18128 gnd.n4731 gnd.n4730 9.3005
R18129 gnd.n4536 gnd.n4535 9.3005
R18130 gnd.n4737 gnd.n4736 9.3005
R18131 gnd.n4739 gnd.n4738 9.3005
R18132 gnd.n4523 gnd.n4522 9.3005
R18133 gnd.n4745 gnd.n4744 9.3005
R18134 gnd.n4747 gnd.n4746 9.3005
R18135 gnd.n4513 gnd.n4512 9.3005
R18136 gnd.n4753 gnd.n4752 9.3005
R18137 gnd.n4755 gnd.n4754 9.3005
R18138 gnd.n4497 gnd.n4495 9.3005
R18139 gnd.n4761 gnd.n4760 9.3005
R18140 gnd.n4762 gnd.n4494 9.3005
R18141 gnd.n4500 gnd.n1099 9.3005
R18142 gnd.n4498 gnd.n4496 9.3005
R18143 gnd.n4759 gnd.n4758 9.3005
R18144 gnd.n4757 gnd.n4756 9.3005
R18145 gnd.n4508 gnd.n4507 9.3005
R18146 gnd.n4751 gnd.n4750 9.3005
R18147 gnd.n4749 gnd.n4748 9.3005
R18148 gnd.n4519 gnd.n4518 9.3005
R18149 gnd.n4743 gnd.n4742 9.3005
R18150 gnd.n4741 gnd.n4740 9.3005
R18151 gnd.n4530 gnd.n4529 9.3005
R18152 gnd.n4735 gnd.n4734 9.3005
R18153 gnd.n4733 gnd.n4732 9.3005
R18154 gnd.n4542 gnd.n4541 9.3005
R18155 gnd.n4727 gnd.n4726 9.3005
R18156 gnd.n4725 gnd.n4724 9.3005
R18157 gnd.n4557 gnd.n4556 9.3005
R18158 gnd.n4719 gnd.n4718 9.3005
R18159 gnd.n6051 gnd.n1100 9.3005
R18160 gnd.n6050 gnd.n6049 9.3005
R18161 gnd.n6048 gnd.n1104 9.3005
R18162 gnd.n6047 gnd.n6046 9.3005
R18163 gnd.n6045 gnd.n1105 9.3005
R18164 gnd.n6044 gnd.n6043 9.3005
R18165 gnd.n6042 gnd.n1109 9.3005
R18166 gnd.n6041 gnd.n6040 9.3005
R18167 gnd.n6039 gnd.n1110 9.3005
R18168 gnd.n6038 gnd.n6037 9.3005
R18169 gnd.n6036 gnd.n1114 9.3005
R18170 gnd.n6035 gnd.n6034 9.3005
R18171 gnd.n6033 gnd.n1115 9.3005
R18172 gnd.n6032 gnd.n6031 9.3005
R18173 gnd.n6030 gnd.n1119 9.3005
R18174 gnd.n6029 gnd.n6028 9.3005
R18175 gnd.n6027 gnd.n1120 9.3005
R18176 gnd.n6026 gnd.n6025 9.3005
R18177 gnd.n6024 gnd.n1124 9.3005
R18178 gnd.n6023 gnd.n6022 9.3005
R18179 gnd.n6021 gnd.n1125 9.3005
R18180 gnd.n6020 gnd.n6019 9.3005
R18181 gnd.n6018 gnd.n1129 9.3005
R18182 gnd.n6017 gnd.n6016 9.3005
R18183 gnd.n6015 gnd.n1130 9.3005
R18184 gnd.n6014 gnd.n6013 9.3005
R18185 gnd.n6012 gnd.n1134 9.3005
R18186 gnd.n6011 gnd.n6010 9.3005
R18187 gnd.n6009 gnd.n1135 9.3005
R18188 gnd.n6008 gnd.n6007 9.3005
R18189 gnd.n6006 gnd.n1139 9.3005
R18190 gnd.n6005 gnd.n6004 9.3005
R18191 gnd.n6003 gnd.n1140 9.3005
R18192 gnd.n6002 gnd.n6001 9.3005
R18193 gnd.n6000 gnd.n1144 9.3005
R18194 gnd.n5999 gnd.n5998 9.3005
R18195 gnd.n5997 gnd.n1145 9.3005
R18196 gnd.n5996 gnd.n5995 9.3005
R18197 gnd.n5994 gnd.n1149 9.3005
R18198 gnd.n5993 gnd.n5992 9.3005
R18199 gnd.n5991 gnd.n1150 9.3005
R18200 gnd.n5990 gnd.n5989 9.3005
R18201 gnd.n5988 gnd.n1154 9.3005
R18202 gnd.n5987 gnd.n5986 9.3005
R18203 gnd.n5985 gnd.n1155 9.3005
R18204 gnd.n5984 gnd.n5983 9.3005
R18205 gnd.n5982 gnd.n1159 9.3005
R18206 gnd.n5981 gnd.n5980 9.3005
R18207 gnd.n5979 gnd.n1160 9.3005
R18208 gnd.n5978 gnd.n5977 9.3005
R18209 gnd.n5976 gnd.n1164 9.3005
R18210 gnd.n5975 gnd.n5974 9.3005
R18211 gnd.n5973 gnd.n1165 9.3005
R18212 gnd.n5972 gnd.n5971 9.3005
R18213 gnd.n5970 gnd.n1169 9.3005
R18214 gnd.n5969 gnd.n5968 9.3005
R18215 gnd.n5967 gnd.n1170 9.3005
R18216 gnd.n5966 gnd.n5965 9.3005
R18217 gnd.n5964 gnd.n1174 9.3005
R18218 gnd.n5963 gnd.n5962 9.3005
R18219 gnd.n5961 gnd.n1175 9.3005
R18220 gnd.n5960 gnd.n5959 9.3005
R18221 gnd.n5958 gnd.n1179 9.3005
R18222 gnd.n5957 gnd.n5956 9.3005
R18223 gnd.n5955 gnd.n1180 9.3005
R18224 gnd.n5954 gnd.n5953 9.3005
R18225 gnd.n5952 gnd.n1184 9.3005
R18226 gnd.n5951 gnd.n5950 9.3005
R18227 gnd.n5949 gnd.n1185 9.3005
R18228 gnd.n5948 gnd.n5947 9.3005
R18229 gnd.n5946 gnd.n1189 9.3005
R18230 gnd.n5945 gnd.n5944 9.3005
R18231 gnd.n5943 gnd.n1190 9.3005
R18232 gnd.n5942 gnd.n5941 9.3005
R18233 gnd.n5940 gnd.n1194 9.3005
R18234 gnd.n5939 gnd.n5938 9.3005
R18235 gnd.n5937 gnd.n1195 9.3005
R18236 gnd.n5936 gnd.n5935 9.3005
R18237 gnd.n5934 gnd.n1199 9.3005
R18238 gnd.n5933 gnd.n5932 9.3005
R18239 gnd.n5931 gnd.n1200 9.3005
R18240 gnd.n5930 gnd.n5929 9.3005
R18241 gnd.n5928 gnd.n1204 9.3005
R18242 gnd.n5927 gnd.n5926 9.3005
R18243 gnd.n5925 gnd.n1205 9.3005
R18244 gnd.n5924 gnd.n5923 9.3005
R18245 gnd.n5922 gnd.n1209 9.3005
R18246 gnd.n5921 gnd.n5920 9.3005
R18247 gnd.n5919 gnd.n1210 9.3005
R18248 gnd.n5918 gnd.n5917 9.3005
R18249 gnd.n5916 gnd.n1214 9.3005
R18250 gnd.n5915 gnd.n5914 9.3005
R18251 gnd.n5913 gnd.n1215 9.3005
R18252 gnd.n5912 gnd.n5911 9.3005
R18253 gnd.n5910 gnd.n1219 9.3005
R18254 gnd.n5909 gnd.n5908 9.3005
R18255 gnd.n5907 gnd.n1220 9.3005
R18256 gnd.n5906 gnd.n5905 9.3005
R18257 gnd.n5904 gnd.n1224 9.3005
R18258 gnd.n5903 gnd.n5902 9.3005
R18259 gnd.n5901 gnd.n1225 9.3005
R18260 gnd.n6053 gnd.n6052 9.3005
R18261 gnd.n441 gnd.n440 9.3005
R18262 gnd.n7168 gnd.n7167 9.3005
R18263 gnd.n7169 gnd.n439 9.3005
R18264 gnd.n7171 gnd.n7170 9.3005
R18265 gnd.n423 gnd.n422 9.3005
R18266 gnd.n7184 gnd.n7183 9.3005
R18267 gnd.n7185 gnd.n421 9.3005
R18268 gnd.n7187 gnd.n7186 9.3005
R18269 gnd.n407 gnd.n406 9.3005
R18270 gnd.n7200 gnd.n7199 9.3005
R18271 gnd.n7201 gnd.n405 9.3005
R18272 gnd.n7203 gnd.n7202 9.3005
R18273 gnd.n391 gnd.n390 9.3005
R18274 gnd.n7216 gnd.n7215 9.3005
R18275 gnd.n7217 gnd.n389 9.3005
R18276 gnd.n7219 gnd.n7218 9.3005
R18277 gnd.n375 gnd.n374 9.3005
R18278 gnd.n7232 gnd.n7231 9.3005
R18279 gnd.n7233 gnd.n373 9.3005
R18280 gnd.n7235 gnd.n7234 9.3005
R18281 gnd.n359 gnd.n358 9.3005
R18282 gnd.n7248 gnd.n7247 9.3005
R18283 gnd.n7249 gnd.n357 9.3005
R18284 gnd.n7251 gnd.n7250 9.3005
R18285 gnd.n343 gnd.n342 9.3005
R18286 gnd.n7264 gnd.n7263 9.3005
R18287 gnd.n7265 gnd.n341 9.3005
R18288 gnd.n7267 gnd.n7266 9.3005
R18289 gnd.n327 gnd.n326 9.3005
R18290 gnd.n7280 gnd.n7279 9.3005
R18291 gnd.n7281 gnd.n324 9.3005
R18292 gnd.n7283 gnd.n7282 9.3005
R18293 gnd.n310 gnd.n309 9.3005
R18294 gnd.n7296 gnd.n7295 9.3005
R18295 gnd.n7297 gnd.n308 9.3005
R18296 gnd.n7299 gnd.n7298 9.3005
R18297 gnd.n296 gnd.n295 9.3005
R18298 gnd.n7312 gnd.n7311 9.3005
R18299 gnd.n7313 gnd.n294 9.3005
R18300 gnd.n7315 gnd.n7314 9.3005
R18301 gnd.n280 gnd.n279 9.3005
R18302 gnd.n7328 gnd.n7327 9.3005
R18303 gnd.n7329 gnd.n278 9.3005
R18304 gnd.n7331 gnd.n7330 9.3005
R18305 gnd.n266 gnd.n265 9.3005
R18306 gnd.n7344 gnd.n7343 9.3005
R18307 gnd.n7345 gnd.n264 9.3005
R18308 gnd.n7347 gnd.n7346 9.3005
R18309 gnd.n250 gnd.n249 9.3005
R18310 gnd.n7360 gnd.n7359 9.3005
R18311 gnd.n7361 gnd.n248 9.3005
R18312 gnd.n7363 gnd.n7362 9.3005
R18313 gnd.n236 gnd.n235 9.3005
R18314 gnd.n7376 gnd.n7375 9.3005
R18315 gnd.n7377 gnd.n234 9.3005
R18316 gnd.n7379 gnd.n7378 9.3005
R18317 gnd.n221 gnd.n220 9.3005
R18318 gnd.n7392 gnd.n7391 9.3005
R18319 gnd.n7393 gnd.n218 9.3005
R18320 gnd.n7463 gnd.n7462 9.3005
R18321 gnd.n7461 gnd.n219 9.3005
R18322 gnd.n7460 gnd.n7459 9.3005
R18323 gnd.n7458 gnd.n7394 9.3005
R18324 gnd.n7457 gnd.n7456 9.3005
R18325 gnd.n7155 gnd.n7154 9.3005
R18326 gnd.n7453 gnd.n7396 9.3005
R18327 gnd.n7452 gnd.n7451 9.3005
R18328 gnd.n7450 gnd.n7401 9.3005
R18329 gnd.n7449 gnd.n7448 9.3005
R18330 gnd.n7447 gnd.n7402 9.3005
R18331 gnd.n7446 gnd.n7445 9.3005
R18332 gnd.n7444 gnd.n7409 9.3005
R18333 gnd.n7443 gnd.n7442 9.3005
R18334 gnd.n7441 gnd.n7410 9.3005
R18335 gnd.n7440 gnd.n7439 9.3005
R18336 gnd.n7438 gnd.n7417 9.3005
R18337 gnd.n7437 gnd.n7436 9.3005
R18338 gnd.n7435 gnd.n7418 9.3005
R18339 gnd.n7434 gnd.n7433 9.3005
R18340 gnd.n7432 gnd.n7425 9.3005
R18341 gnd.n7431 gnd.n7430 9.3005
R18342 gnd.n124 gnd.n121 9.3005
R18343 gnd.n7557 gnd.n7556 9.3005
R18344 gnd.n7455 gnd.n7454 9.3005
R18345 gnd.n6803 gnd.n6802 9.3005
R18346 gnd.n6804 gnd.n589 9.3005
R18347 gnd.n7020 gnd.n7019 9.3005
R18348 gnd.n7018 gnd.n590 9.3005
R18349 gnd.n7017 gnd.n7016 9.3005
R18350 gnd.n7015 gnd.n6805 9.3005
R18351 gnd.n7014 gnd.n7013 9.3005
R18352 gnd.n7012 gnd.n6808 9.3005
R18353 gnd.n7011 gnd.n7010 9.3005
R18354 gnd.n7009 gnd.n6809 9.3005
R18355 gnd.n7008 gnd.n7007 9.3005
R18356 gnd.n7006 gnd.n6958 9.3005
R18357 gnd.n7005 gnd.n7004 9.3005
R18358 gnd.n7003 gnd.n6959 9.3005
R18359 gnd.n7002 gnd.n7001 9.3005
R18360 gnd.n7000 gnd.n6962 9.3005
R18361 gnd.n6999 gnd.n6998 9.3005
R18362 gnd.n6997 gnd.n6963 9.3005
R18363 gnd.n6996 gnd.n6995 9.3005
R18364 gnd.n6994 gnd.n6966 9.3005
R18365 gnd.n6993 gnd.n6992 9.3005
R18366 gnd.n6991 gnd.n6967 9.3005
R18367 gnd.n6990 gnd.n6989 9.3005
R18368 gnd.n6988 gnd.n6970 9.3005
R18369 gnd.n6987 gnd.n6986 9.3005
R18370 gnd.n6985 gnd.n6971 9.3005
R18371 gnd.n6984 gnd.n6983 9.3005
R18372 gnd.n6982 gnd.n6974 9.3005
R18373 gnd.n6981 gnd.n6980 9.3005
R18374 gnd.n6979 gnd.n6975 9.3005
R18375 gnd.n6978 gnd.n79 9.3005
R18376 gnd.n7606 gnd.n80 9.3005
R18377 gnd.n7605 gnd.n7604 9.3005
R18378 gnd.n7603 gnd.n81 9.3005
R18379 gnd.n7602 gnd.n7601 9.3005
R18380 gnd.n7600 gnd.n85 9.3005
R18381 gnd.n7599 gnd.n7598 9.3005
R18382 gnd.n7597 gnd.n86 9.3005
R18383 gnd.n7596 gnd.n7595 9.3005
R18384 gnd.n7594 gnd.n90 9.3005
R18385 gnd.n7593 gnd.n7592 9.3005
R18386 gnd.n7591 gnd.n91 9.3005
R18387 gnd.n7590 gnd.n7589 9.3005
R18388 gnd.n7588 gnd.n95 9.3005
R18389 gnd.n7587 gnd.n7586 9.3005
R18390 gnd.n7585 gnd.n96 9.3005
R18391 gnd.n7584 gnd.n7583 9.3005
R18392 gnd.n7582 gnd.n100 9.3005
R18393 gnd.n7581 gnd.n7580 9.3005
R18394 gnd.n7579 gnd.n101 9.3005
R18395 gnd.n7578 gnd.n7577 9.3005
R18396 gnd.n7576 gnd.n105 9.3005
R18397 gnd.n7575 gnd.n7574 9.3005
R18398 gnd.n7573 gnd.n106 9.3005
R18399 gnd.n7572 gnd.n7571 9.3005
R18400 gnd.n7570 gnd.n110 9.3005
R18401 gnd.n7569 gnd.n7568 9.3005
R18402 gnd.n7567 gnd.n111 9.3005
R18403 gnd.n7566 gnd.n7565 9.3005
R18404 gnd.n7564 gnd.n115 9.3005
R18405 gnd.n7563 gnd.n7562 9.3005
R18406 gnd.n7561 gnd.n116 9.3005
R18407 gnd.n7560 gnd.n7559 9.3005
R18408 gnd.n7558 gnd.n120 9.3005
R18409 gnd.n592 gnd.n591 9.3005
R18410 gnd.n2866 gnd.t165 9.29782
R18411 gnd.n2566 gnd.t271 9.29782
R18412 gnd.t234 gnd.n5091 9.24152
R18413 gnd.n5511 gnd.t349 9.24152
R18414 gnd.t216 gnd.n384 9.24152
R18415 gnd.n262 gnd.t73 9.24152
R18416 gnd.n2857 gnd.t165 8.93321
R18417 gnd.t143 gnd.n2308 8.93321
R18418 gnd.t135 gnd.n2309 8.93321
R18419 gnd.n4917 gnd.n1764 8.92286
R18420 gnd.n5104 gnd.n1672 8.92286
R18421 gnd.n5164 gnd.n5163 8.92286
R18422 gnd.n5281 gnd.n1587 8.92286
R18423 gnd.n5342 gnd.n5341 8.92286
R18424 gnd.n5442 gnd.n1499 8.92286
R18425 gnd.n5514 gnd.n5513 8.92286
R18426 gnd.n5623 gnd.n1408 8.92286
R18427 gnd.n5747 gnd.n1381 8.92286
R18428 gnd.n3569 gnd.n3544 8.92171
R18429 gnd.n3537 gnd.n3512 8.92171
R18430 gnd.n3505 gnd.n3480 8.92171
R18431 gnd.n3474 gnd.n3449 8.92171
R18432 gnd.n3442 gnd.n3417 8.92171
R18433 gnd.n3410 gnd.n3385 8.92171
R18434 gnd.n3378 gnd.n3353 8.92171
R18435 gnd.n3347 gnd.n3322 8.92171
R18436 gnd.n5674 gnd.n5656 8.72777
R18437 gnd.n6078 gnd.t34 8.60421
R18438 gnd.n4622 gnd.t139 8.60421
R18439 gnd.t295 gnd.n1777 8.60421
R18440 gnd.n4896 gnd.n1777 8.60421
R18441 gnd.t24 gnd.n5279 8.60421
R18442 gnd.n5312 gnd.t358 8.60421
R18443 gnd.n5829 gnd.t360 8.60421
R18444 gnd.n5881 gnd.t103 8.60421
R18445 gnd.n6818 gnd.t224 8.60421
R18446 gnd.n6778 gnd.n283 8.60421
R18447 gnd.n232 gnd.t253 8.60421
R18448 gnd.n3225 gnd.t266 8.56861
R18449 gnd.n2497 gnd.n2477 8.43467
R18450 gnd.n58 gnd.n38 8.43467
R18451 gnd.n4097 gnd.n0 8.41456
R18452 gnd.n7607 gnd.n7606 8.41456
R18453 gnd.n6079 gnd.n6078 8.28555
R18454 gnd.n4434 gnd.n2004 8.28555
R18455 gnd.n6072 gnd.n1068 8.28555
R18456 gnd.n4443 gnd.n1071 8.28555
R18457 gnd.n6066 gnd.n1080 8.28555
R18458 gnd.n4782 gnd.n1083 8.28555
R18459 gnd.n6060 gnd.n1091 8.28555
R18460 gnd.n4774 gnd.n1094 8.28555
R18461 gnd.n4906 gnd.t153 8.28555
R18462 gnd.n5083 gnd.n1685 8.28555
R18463 gnd.n5156 gnd.n1645 8.28555
R18464 gnd.n5260 gnd.n1600 8.28555
R18465 gnd.n5334 gnd.n1558 8.28555
R18466 gnd.n5422 gnd.n1513 8.28555
R18467 gnd.n5479 gnd.n1464 8.28555
R18468 gnd.t159 gnd.n1402 8.28555
R18469 gnd.n7157 gnd.n453 8.28555
R18470 gnd.n6800 gnd.n6799 8.28555
R18471 gnd.n7165 gnd.n445 8.28555
R18472 gnd.n7022 gnd.n434 8.28555
R18473 gnd.n7173 gnd.n437 8.28555
R18474 gnd.n6814 gnd.n425 8.28555
R18475 gnd.n7181 gnd.n428 8.28555
R18476 gnd.n6818 gnd.n416 8.28555
R18477 gnd.t0 gnd.n2351 8.20401
R18478 gnd.n3303 gnd.t276 8.20401
R18479 gnd.n3570 gnd.n3542 8.14595
R18480 gnd.n3538 gnd.n3510 8.14595
R18481 gnd.n3506 gnd.n3478 8.14595
R18482 gnd.n3475 gnd.n3447 8.14595
R18483 gnd.n3443 gnd.n3415 8.14595
R18484 gnd.n3411 gnd.n3383 8.14595
R18485 gnd.n3379 gnd.n3351 8.14595
R18486 gnd.n3348 gnd.n3320 8.14595
R18487 gnd.n3575 gnd.n3574 7.97301
R18488 gnd.n4765 gnd.n4491 7.9669
R18489 gnd.t200 gnd.n1700 7.9669
R18490 gnd.n5579 gnd.t317 7.9669
R18491 gnd.n5890 gnd.n1229 7.9669
R18492 gnd.n3013 gnd.t230 7.83941
R18493 gnd.n7556 gnd.n124 7.75808
R18494 gnd.n7104 gnd.n499 7.75808
R18495 gnd.n4718 gnd.n4556 7.75808
R18496 gnd.n4151 gnd.n4012 7.75808
R18497 gnd.n2931 gnd.n2669 7.65711
R18498 gnd.t153 gnd.n4905 7.64824
R18499 gnd.n4923 gnd.t179 7.64824
R18500 gnd.n4952 gnd.n1720 7.64824
R18501 gnd.n5083 gnd.t57 7.64824
R18502 gnd.n5241 gnd.t44 7.64824
R18503 gnd.n5140 gnd.t44 7.64824
R18504 gnd.t47 gnd.n5325 7.64824
R18505 gnd.n5327 gnd.t47 7.64824
R18506 gnd.n5479 gnd.t59 7.64824
R18507 gnd.n5603 gnd.n1421 7.64824
R18508 gnd.n5620 gnd.t159 7.64824
R18509 gnd.t139 gnd.n4610 7.32958
R18510 gnd.n4666 gnd.t295 7.32958
R18511 gnd.n4896 gnd.n1772 7.32958
R18512 gnd.n5817 gnd.n5816 7.32958
R18513 gnd.t360 gnd.n5828 7.32958
R18514 gnd.n5869 gnd.t103 7.32958
R18515 gnd.n1829 gnd.n1828 7.30353
R18516 gnd.n5673 gnd.n5672 7.30353
R18517 gnd.n2199 gnd.t255 7.11021
R18518 gnd.t77 gnd.n927 7.11021
R18519 gnd.n4917 gnd.n4916 7.01093
R18520 gnd.n4986 gnd.n1734 7.01093
R18521 gnd.n5164 gnd.n1649 7.01093
R18522 gnd.n1607 gnd.t60 7.01093
R18523 gnd.n5281 gnd.n5280 7.01093
R18524 gnd.n5342 gnd.n1562 7.01093
R18525 gnd.t64 gnd.n1547 7.01093
R18526 gnd.n5442 gnd.n5441 7.01093
R18527 gnd.n5623 gnd.n5622 7.01093
R18528 gnd.n5747 gnd.n1380 7.01093
R18529 gnd.n1381 gnd.t129 7.01093
R18530 gnd.n2167 gnd.t221 6.74561
R18531 gnd.t204 gnd.n2035 6.74561
R18532 gnd.n5092 gnd.t234 6.69227
R18533 gnd.n5521 gnd.t349 6.69227
R18534 gnd.n6955 gnd.n419 6.69227
R18535 gnd.n5809 gnd.n5808 6.5566
R18536 gnd.n1890 gnd.n1889 6.5566
R18537 gnd.n4837 gnd.n1834 6.5566
R18538 gnd.n5684 gnd.n5683 6.5566
R18539 gnd.n3001 gnd.t230 6.38101
R18540 gnd.n2135 gnd.t39 6.38101
R18541 gnd.t292 gnd.n2067 6.38101
R18542 gnd.n5011 gnd.n1716 6.37362
R18543 gnd.n4937 gnd.n4936 6.37362
R18544 gnd.n5190 gnd.n1631 6.37362
R18545 gnd.n5318 gnd.n5317 6.37362
R18546 gnd.n5539 gnd.n1452 6.37362
R18547 gnd.n5463 gnd.n5462 6.37362
R18548 gnd.n4704 gnd.n4575 6.20656
R18549 gnd.n7518 gnd.n7515 6.20656
R18550 gnd.n3733 gnd.n3728 6.20656
R18551 gnd.n1294 gnd.n1293 6.20656
R18552 gnd.n2920 gnd.t228 6.01641
R18553 gnd.n2353 gnd.t0 6.01641
R18554 gnd.n3286 gnd.t276 6.01641
R18555 gnd.t4 gnd.n2099 6.01641
R18556 gnd.n2102 gnd.t10 6.01641
R18557 gnd.n3572 gnd.n3542 5.81868
R18558 gnd.n3540 gnd.n3510 5.81868
R18559 gnd.n3508 gnd.n3478 5.81868
R18560 gnd.n3477 gnd.n3447 5.81868
R18561 gnd.n3445 gnd.n3415 5.81868
R18562 gnd.n3413 gnd.n3383 5.81868
R18563 gnd.n3381 gnd.n3351 5.81868
R18564 gnd.n3350 gnd.n3320 5.81868
R18565 gnd.n4924 gnd.n1752 5.73631
R18566 gnd.n4986 gnd.t100 5.73631
R18567 gnd.n5104 gnd.t61 5.73631
R18568 gnd.n5026 gnd.n5025 5.73631
R18569 gnd.n5112 gnd.n1661 5.73631
R18570 gnd.n5149 gnd.t42 5.73631
R18571 gnd.n5280 gnd.t55 5.73631
R18572 gnd.n1583 gnd.n1572 5.73631
R18573 gnd.n5289 gnd.n1575 5.73631
R18574 gnd.t58 gnd.n1562 5.73631
R18575 gnd.n5404 gnd.t48 5.73631
R18576 gnd.n1495 gnd.n1486 5.73631
R18577 gnd.n5450 gnd.n5448 5.73631
R18578 gnd.n5514 gnd.t54 5.73631
R18579 gnd.n5554 gnd.n5553 5.73631
R18580 gnd.t129 gnd.n1339 5.73631
R18581 gnd.t266 gnd.n2370 5.65181
R18582 gnd.t67 gnd.n2132 5.65181
R18583 gnd.n2070 gnd.t18 5.65181
R18584 gnd.n5813 gnd.n556 5.62001
R18585 gnd.n4832 gnd.n1894 5.62001
R18586 gnd.n4833 gnd.n4832 5.62001
R18587 gnd.n5679 gnd.n556 5.62001
R18588 gnd.n2801 gnd.n2796 5.4308
R18589 gnd.n3617 gnd.n2294 5.4308
R18590 gnd.t345 gnd.n5111 5.41765
R18591 gnd.t232 gnd.n1493 5.41765
R18592 gnd.t269 gnd.n2417 5.28721
R18593 gnd.n2319 gnd.t143 5.28721
R18594 gnd.n3599 gnd.t135 5.28721
R18595 gnd.t261 gnd.n2164 5.28721
R18596 gnd.n2038 gnd.t71 5.28721
R18597 gnd.t20 gnd.t269 5.10491
R18598 gnd.n5059 gnd.n1706 5.09899
R18599 gnd.n5067 gnd.n1700 5.09899
R18600 gnd.t51 gnd.n1635 5.09899
R18601 gnd.n5235 gnd.n1621 5.09899
R18602 gnd.n5244 gnd.n1615 5.09899
R18603 gnd.n5398 gnd.n1534 5.09899
R18604 gnd.n5406 gnd.n1528 5.09899
R18605 gnd.n1520 gnd.t53 5.09899
R18606 gnd.n5579 gnd.n1442 5.09899
R18607 gnd.n5587 gnd.n1436 5.09899
R18608 gnd.n3570 gnd.n3569 5.04292
R18609 gnd.n3538 gnd.n3537 5.04292
R18610 gnd.n3506 gnd.n3505 5.04292
R18611 gnd.n3475 gnd.n3474 5.04292
R18612 gnd.n3443 gnd.n3442 5.04292
R18613 gnd.n3411 gnd.n3410 5.04292
R18614 gnd.n3379 gnd.n3378 5.04292
R18615 gnd.n3348 gnd.n3347 5.04292
R18616 gnd.n3073 gnd.t271 4.92261
R18617 gnd.t250 gnd.n2196 4.92261
R18618 gnd.n2517 gnd.n2516 4.82753
R18619 gnd.n78 gnd.n77 4.82753
R18620 gnd.n4672 gnd.t306 4.78034
R18621 gnd.n5112 gnd.t345 4.78034
R18622 gnd.n1495 gnd.t232 4.78034
R18623 gnd.n5557 gnd.t319 4.78034
R18624 gnd.n5816 gnd.t111 4.78034
R18625 gnd.n2522 gnd.n2519 4.74817
R18626 gnd.n2572 gnd.n2458 4.74817
R18627 gnd.n2559 gnd.n2457 4.74817
R18628 gnd.n2456 gnd.n2455 4.74817
R18629 gnd.n2568 gnd.n2519 4.74817
R18630 gnd.n2569 gnd.n2458 4.74817
R18631 gnd.n2571 gnd.n2457 4.74817
R18632 gnd.n2558 gnd.n2456 4.74817
R18633 gnd.n2497 gnd.n2496 4.7074
R18634 gnd.n58 gnd.n57 4.7074
R18635 gnd.n2517 gnd.n2497 4.65959
R18636 gnd.n78 gnd.n58 4.65959
R18637 gnd.n7071 gnd.n558 4.6132
R18638 gnd.n4828 gnd.n4827 4.6132
R18639 gnd.t272 gnd.n2588 4.55801
R18640 gnd.n4931 gnd.n1758 4.46168
R18641 gnd.n4974 gnd.n1744 4.46168
R18642 gnd.n4952 gnd.t49 4.46168
R18643 gnd.n5119 gnd.n1666 4.46168
R18644 gnd.n5110 gnd.n1654 4.46168
R18645 gnd.n5296 gnd.n1580 4.46168
R18646 gnd.n5287 gnd.n1566 4.46168
R18647 gnd.n5457 gnd.n1492 4.46168
R18648 gnd.n5501 gnd.n1477 4.46168
R18649 gnd.n5603 gnd.t45 4.46168
R18650 gnd.n5631 gnd.n1402 4.46168
R18651 gnd.n5652 gnd.n5651 4.46168
R18652 gnd.n5669 gnd.n5656 4.46111
R18653 gnd.n3555 gnd.n3551 4.38594
R18654 gnd.n3523 gnd.n3519 4.38594
R18655 gnd.n3491 gnd.n3487 4.38594
R18656 gnd.n3460 gnd.n3456 4.38594
R18657 gnd.n3428 gnd.n3424 4.38594
R18658 gnd.n3396 gnd.n3392 4.38594
R18659 gnd.n3364 gnd.n3360 4.38594
R18660 gnd.n3333 gnd.n3329 4.38594
R18661 gnd.n3566 gnd.n3544 4.26717
R18662 gnd.n3534 gnd.n3512 4.26717
R18663 gnd.n3502 gnd.n3480 4.26717
R18664 gnd.n3471 gnd.n3449 4.26717
R18665 gnd.n3439 gnd.n3417 4.26717
R18666 gnd.n3407 gnd.n3385 4.26717
R18667 gnd.n3375 gnd.n3353 4.26717
R18668 gnd.n3344 gnd.n3322 4.26717
R18669 gnd.n2982 gnd.t277 4.19341
R18670 gnd.n5141 gnd.t219 4.14303
R18671 gnd.n5367 gnd.t347 4.14303
R18672 gnd.n3574 gnd.n3573 4.08274
R18673 gnd.n5808 gnd.n5807 4.05904
R18674 gnd.n1889 gnd.n1888 4.05904
R18675 gnd.n4840 gnd.n1834 4.05904
R18676 gnd.n5685 gnd.n5684 4.05904
R18677 gnd.n2942 gnd.n2661 4.01111
R18678 gnd.n2664 gnd.n2662 4.01111
R18679 gnd.n2952 gnd.n2951 4.01111
R18680 gnd.n2963 gnd.n2645 4.01111
R18681 gnd.n2962 gnd.n2648 4.01111
R18682 gnd.n2973 gnd.n2636 4.01111
R18683 gnd.n2639 gnd.n2637 4.01111
R18684 gnd.n2983 gnd.n2982 4.01111
R18685 gnd.n2993 gnd.n2617 4.01111
R18686 gnd.n2992 gnd.n2620 4.01111
R18687 gnd.n3001 gnd.n2611 4.01111
R18688 gnd.n3013 gnd.n2601 4.01111
R18689 gnd.n3023 gnd.n2586 4.01111
R18690 gnd.n3039 gnd.n3038 4.01111
R18691 gnd.n2588 gnd.n2525 4.01111
R18692 gnd.n3093 gnd.n2526 4.01111
R18693 gnd.n3087 gnd.n3086 4.01111
R18694 gnd.n2575 gnd.n2537 4.01111
R18695 gnd.n3079 gnd.n2548 4.01111
R18696 gnd.n2566 gnd.n2561 4.01111
R18697 gnd.n3073 gnd.n3072 4.01111
R18698 gnd.n3119 gnd.n2452 4.01111
R18699 gnd.n3118 gnd.n3117 4.01111
R18700 gnd.n3130 gnd.n3129 4.01111
R18701 gnd.n2445 gnd.n2437 4.01111
R18702 gnd.n3159 gnd.n2425 4.01111
R18703 gnd.n3158 gnd.n2428 4.01111
R18704 gnd.n3169 gnd.n2417 4.01111
R18705 gnd.n2418 gnd.n2406 4.01111
R18706 gnd.n3180 gnd.n2407 4.01111
R18707 gnd.n3204 gnd.n2398 4.01111
R18708 gnd.n3203 gnd.n2389 4.01111
R18709 gnd.n3226 gnd.n3225 4.01111
R18710 gnd.n3244 gnd.n2370 4.01111
R18711 gnd.n3243 gnd.n2373 4.01111
R18712 gnd.n3254 gnd.n2362 4.01111
R18713 gnd.n2363 gnd.n2350 4.01111
R18714 gnd.n3265 gnd.n2351 4.01111
R18715 gnd.n3292 gnd.n2335 4.01111
R18716 gnd.n3304 gnd.n3303 4.01111
R18717 gnd.n3286 gnd.n2328 4.01111
R18718 gnd.n3315 gnd.n3314 4.01111
R18719 gnd.n3587 gnd.n2316 4.01111
R18720 gnd.n3586 gnd.n2319 4.01111
R18721 gnd.n3599 gnd.n2308 4.01111
R18722 gnd.n2309 gnd.n2301 4.01111
R18723 gnd.n3609 gnd.n2227 4.01111
R18724 gnd.n19 gnd.n9 3.99943
R18725 gnd.n2620 gnd.t264 3.82881
R18726 gnd.n2428 gnd.t20 3.82881
R18727 gnd.n3293 gnd.t270 3.82881
R18728 gnd.n6246 gnd.n927 3.82881
R18729 gnd.n6079 gnd.n1056 3.82437
R18730 gnd.n4477 gnd.n1960 3.82437
R18731 gnd.t179 gnd.n1744 3.82437
R18732 gnd.t49 gnd.n1729 3.82437
R18733 gnd.n5003 gnd.n1714 3.82437
R18734 gnd.n5076 gnd.n5075 3.82437
R18735 gnd.t50 gnd.n1649 3.82437
R18736 gnd.n5181 gnd.n1629 3.82437
R18737 gnd.n5253 gnd.n5252 3.82437
R18738 gnd.n5359 gnd.n1542 3.82437
R18739 gnd.n5415 gnd.n5414 3.82437
R18740 gnd.n5441 gnd.t52 3.82437
R18741 gnd.n5531 gnd.n1450 3.82437
R18742 gnd.n5596 gnd.n5595 3.82437
R18743 gnd.n5548 gnd.t45 3.82437
R18744 gnd.n5829 gnd.t111 3.82437
R18745 gnd.n7102 gnd.n506 3.82437
R18746 gnd.n3574 gnd.n3446 3.70378
R18747 gnd.n3097 gnd.n2518 3.65935
R18748 gnd.n19 gnd.n18 3.60163
R18749 gnd.n4782 gnd.t107 3.50571
R18750 gnd.t280 gnd.n4648 3.50571
R18751 gnd.t282 gnd.n5847 3.50571
R18752 gnd.n7165 gnd.t114 3.50571
R18753 gnd.n7473 gnd.t90 3.50571
R18754 gnd.n3565 gnd.n3546 3.49141
R18755 gnd.n3533 gnd.n3514 3.49141
R18756 gnd.n3501 gnd.n3482 3.49141
R18757 gnd.n3470 gnd.n3451 3.49141
R18758 gnd.n3438 gnd.n3419 3.49141
R18759 gnd.n3406 gnd.n3387 3.49141
R18760 gnd.n3374 gnd.n3355 3.49141
R18761 gnd.n3343 gnd.n3324 3.49141
R18762 gnd.t321 gnd.n3049 3.46421
R18763 gnd.n3050 gnd.t279 3.46421
R18764 gnd.t329 gnd.n2452 3.46421
R18765 gnd.t274 gnd.n3214 3.46421
R18766 gnd.n4905 gnd.n4904 3.18706
R18767 gnd.t100 gnd.n4985 3.18706
R18768 gnd.n4984 gnd.n4983 3.18706
R18769 gnd.n5091 gnd.n5090 3.18706
R18770 gnd.n5162 gnd.n1643 3.18706
R18771 gnd.n5269 gnd.n5267 3.18706
R18772 gnd.n5340 gnd.n1555 3.18706
R18773 gnd.n5430 gnd.n5429 3.18706
R18774 gnd.n5512 gnd.n5511 3.18706
R18775 gnd.n5611 gnd.n5610 3.18706
R18776 gnd.n5640 gnd.t150 3.18706
R18777 gnd.n5819 gnd.n1339 3.18706
R18778 gnd.n3117 gnd.t273 3.0996
R18779 gnd.t275 gnd.n3140 3.0996
R18780 gnd.t351 gnd.n2382 3.0996
R18781 gnd.n5058 gnd.t200 2.8684
R18782 gnd.t317 gnd.n5578 2.8684
R18783 gnd.n2498 gnd.t218 2.82907
R18784 gnd.n2498 gnd.t78 2.82907
R18785 gnd.n2500 gnd.t344 2.82907
R18786 gnd.n2500 gnd.t310 2.82907
R18787 gnd.n2502 gnd.t199 2.82907
R18788 gnd.n2502 gnd.t312 2.82907
R18789 gnd.n2504 gnd.t259 2.82907
R18790 gnd.n2504 gnd.t326 2.82907
R18791 gnd.n2506 gnd.t294 2.82907
R18792 gnd.n2506 gnd.t11 2.82907
R18793 gnd.n2508 gnd.t40 2.82907
R18794 gnd.n2508 gnd.t197 2.82907
R18795 gnd.n2510 gnd.t86 2.82907
R18796 gnd.n2510 gnd.t263 2.82907
R18797 gnd.n2512 gnd.t262 2.82907
R18798 gnd.n2512 gnd.t357 2.82907
R18799 gnd.n2514 gnd.t314 2.82907
R18800 gnd.n2514 gnd.t198 2.82907
R18801 gnd.n2459 gnd.t289 2.82907
R18802 gnd.n2459 gnd.t241 2.82907
R18803 gnd.n2461 gnd.t287 2.82907
R18804 gnd.n2461 gnd.t245 2.82907
R18805 gnd.n2463 gnd.t19 2.82907
R18806 gnd.n2463 gnd.t80 2.82907
R18807 gnd.n2465 gnd.t70 2.82907
R18808 gnd.n2465 gnd.t293 2.82907
R18809 gnd.n2467 gnd.t5 2.82907
R18810 gnd.n2467 gnd.t239 2.82907
R18811 gnd.n2469 gnd.t84 2.82907
R18812 gnd.n2469 gnd.t288 2.82907
R18813 gnd.n2471 gnd.t355 2.82907
R18814 gnd.n2471 gnd.t68 2.82907
R18815 gnd.n2473 gnd.t340 2.82907
R18816 gnd.n2473 gnd.t222 2.82907
R18817 gnd.n2475 gnd.t256 2.82907
R18818 gnd.n2475 gnd.t324 2.82907
R18819 gnd.n2478 gnd.t37 2.82907
R18820 gnd.n2478 gnd.t353 2.82907
R18821 gnd.n2480 gnd.t205 2.82907
R18822 gnd.n2480 gnd.t72 2.82907
R18823 gnd.n2482 gnd.t332 2.82907
R18824 gnd.n2482 gnd.t17 2.82907
R18825 gnd.n2484 gnd.t362 2.82907
R18826 gnd.n2484 gnd.t342 2.82907
R18827 gnd.n2486 gnd.t301 2.82907
R18828 gnd.n2486 gnd.t38 2.82907
R18829 gnd.n2488 gnd.t240 2.82907
R18830 gnd.n2488 gnd.t27 2.82907
R18831 gnd.n2490 gnd.t298 2.82907
R18832 gnd.n2490 gnd.t238 2.82907
R18833 gnd.n2492 gnd.t284 2.82907
R18834 gnd.n2492 gnd.t243 2.82907
R18835 gnd.n2494 gnd.t300 2.82907
R18836 gnd.n2494 gnd.t66 2.82907
R18837 gnd.n75 gnd.t313 2.82907
R18838 gnd.n75 gnd.t328 2.82907
R18839 gnd.n73 gnd.t311 2.82907
R18840 gnd.n73 gnd.t327 2.82907
R18841 gnd.n71 gnd.t33 2.82907
R18842 gnd.n71 gnd.t260 2.82907
R18843 gnd.n69 gnd.t211 2.82907
R18844 gnd.n69 gnd.t208 2.82907
R18845 gnd.n67 gnd.t308 2.82907
R18846 gnd.n67 gnd.t304 2.82907
R18847 gnd.n65 gnd.t209 2.82907
R18848 gnd.n65 gnd.t215 2.82907
R18849 gnd.n63 gnd.t333 2.82907
R18850 gnd.n63 gnd.t79 2.82907
R18851 gnd.n61 gnd.t217 2.82907
R18852 gnd.n61 gnd.t258 2.82907
R18853 gnd.n59 gnd.t213 2.82907
R18854 gnd.n59 gnd.t305 2.82907
R18855 gnd.n36 gnd.t81 2.82907
R18856 gnd.n36 gnd.t9 2.82907
R18857 gnd.n34 gnd.t356 2.82907
R18858 gnd.n34 gnd.t244 2.82907
R18859 gnd.n32 gnd.t337 2.82907
R18860 gnd.n32 gnd.t31 2.82907
R18861 gnd.n30 gnd.t246 2.82907
R18862 gnd.n30 gnd.t299 2.82907
R18863 gnd.n28 gnd.t363 2.82907
R18864 gnd.n28 gnd.t203 2.82907
R18865 gnd.n26 gnd.t302 2.82907
R18866 gnd.n26 gnd.t341 2.82907
R18867 gnd.n24 gnd.t83 2.82907
R18868 gnd.n24 gnd.t7 2.82907
R18869 gnd.n22 gnd.t257 2.82907
R18870 gnd.n22 gnd.t247 2.82907
R18871 gnd.n20 gnd.t339 2.82907
R18872 gnd.n20 gnd.t354 2.82907
R18873 gnd.n55 gnd.t15 2.82907
R18874 gnd.n55 gnd.t223 2.82907
R18875 gnd.n53 gnd.t249 2.82907
R18876 gnd.n53 gnd.t74 2.82907
R18877 gnd.n51 gnd.t290 2.82907
R18878 gnd.n51 gnd.t242 2.82907
R18879 gnd.n49 gnd.t335 2.82907
R18880 gnd.n49 gnd.t334 2.82907
R18881 gnd.n47 gnd.t88 2.82907
R18882 gnd.n47 gnd.t331 2.82907
R18883 gnd.n45 gnd.t29 2.82907
R18884 gnd.n45 gnd.t325 2.82907
R18885 gnd.n43 gnd.t206 2.82907
R18886 gnd.n43 gnd.t291 2.82907
R18887 gnd.n41 gnd.t297 2.82907
R18888 gnd.n41 gnd.t76 2.82907
R18889 gnd.n39 gnd.t323 2.82907
R18890 gnd.n39 gnd.t13 2.82907
R18891 gnd.n3080 gnd.t278 2.735
R18892 gnd.n2407 gnd.t267 2.735
R18893 gnd.n3562 gnd.n3561 2.71565
R18894 gnd.n3530 gnd.n3529 2.71565
R18895 gnd.n3498 gnd.n3497 2.71565
R18896 gnd.n3467 gnd.n3466 2.71565
R18897 gnd.n3435 gnd.n3434 2.71565
R18898 gnd.n3403 gnd.n3402 2.71565
R18899 gnd.n3371 gnd.n3370 2.71565
R18900 gnd.n3340 gnd.n3339 2.71565
R18901 gnd.n4672 gnd.t122 2.54975
R18902 gnd.n4993 gnd.n4992 2.54975
R18903 gnd.t46 gnd.n1716 2.54975
R18904 gnd.n5092 gnd.n1680 2.54975
R18905 gnd.n5126 gnd.t62 2.54975
R18906 gnd.n5171 gnd.n5170 2.54975
R18907 gnd.n5156 gnd.t51 2.54975
R18908 gnd.n5270 gnd.n1595 2.54975
R18909 gnd.n5349 gnd.n5348 2.54975
R18910 gnd.n5422 gnd.t53 2.54975
R18911 gnd.n5431 gnd.n1507 2.54975
R18912 gnd.n5492 gnd.t56 2.54975
R18913 gnd.n5521 gnd.n5520 2.54975
R18914 gnd.n5462 gnd.t41 2.54975
R18915 gnd.n5612 gnd.n1416 2.54975
R18916 gnd.n3024 gnd.t268 2.3704
R18917 gnd.n3254 gnd.t265 2.3704
R18918 gnd.n3097 gnd.n2519 2.27742
R18919 gnd.n3097 gnd.n2458 2.27742
R18920 gnd.n3097 gnd.n2457 2.27742
R18921 gnd.n3097 gnd.n2456 2.27742
R18922 gnd.t219 gnd.n5140 2.23109
R18923 gnd.n5325 gnd.t347 2.23109
R18924 gnd.n4200 gnd.t169 2.0058
R18925 gnd.n3558 gnd.n3548 1.93989
R18926 gnd.n3526 gnd.n3516 1.93989
R18927 gnd.n3494 gnd.n3484 1.93989
R18928 gnd.n3463 gnd.n3453 1.93989
R18929 gnd.n3431 gnd.n3421 1.93989
R18930 gnd.n3399 gnd.n3389 1.93989
R18931 gnd.n3367 gnd.n3357 1.93989
R18932 gnd.n3336 gnd.n3326 1.93989
R18933 gnd.n5005 gnd.n5004 1.91244
R18934 gnd.n1694 gnd.n1693 1.91244
R18935 gnd.n1609 gnd.n1608 1.91244
R18936 gnd.n5361 gnd.n5360 1.91244
R18937 gnd.n5533 gnd.n5532 1.91244
R18938 gnd.n1430 gnd.n1428 1.91244
R18939 gnd.n5651 gnd.t94 1.91244
R18940 gnd.n2603 gnd.t268 1.6412
R18941 gnd.t22 gnd.n5183 1.59378
R18942 gnd.n1522 gnd.t315 1.59378
R18943 gnd.n7205 gnd.t12 1.59378
R18944 gnd.n7365 gnd.t14 1.59378
R18945 gnd.n2951 gnd.t194 1.2766
R18946 gnd.n2574 gnd.t278 1.2766
R18947 gnd.t97 gnd.n4915 1.27512
R18948 gnd.n4915 gnd.n4914 1.27512
R18949 gnd.n4973 gnd.n1745 1.27512
R18950 gnd.t61 gnd.n5103 1.27512
R18951 gnd.n5101 gnd.n5100 1.27512
R18952 gnd.n5135 gnd.n5134 1.27512
R18953 gnd.n5279 gnd.n5278 1.27512
R18954 gnd.n5312 gnd.n5311 1.27512
R18955 gnd.n5440 gnd.n5439 1.27512
R18956 gnd.n5500 gnd.n1479 1.27512
R18957 gnd.n1478 gnd.t54 1.27512
R18958 gnd.n5621 gnd.n5620 1.27512
R18959 gnd.n5650 gnd.n1389 1.27512
R18960 gnd.n2804 gnd.n2796 1.16414
R18961 gnd.n3620 gnd.n2294 1.16414
R18962 gnd.n3557 gnd.n3550 1.16414
R18963 gnd.n3525 gnd.n3518 1.16414
R18964 gnd.n3493 gnd.n3486 1.16414
R18965 gnd.n3462 gnd.n3455 1.16414
R18966 gnd.n3430 gnd.n3423 1.16414
R18967 gnd.n3398 gnd.n3391 1.16414
R18968 gnd.n3366 gnd.n3359 1.16414
R18969 gnd.n3335 gnd.n3328 1.16414
R18970 gnd.n7071 gnd.n7070 0.970197
R18971 gnd.n4828 gnd.n1895 0.970197
R18972 gnd.n3541 gnd.n3509 0.962709
R18973 gnd.n3573 gnd.n3541 0.962709
R18974 gnd.n3414 gnd.n3382 0.962709
R18975 gnd.n3446 gnd.n3414 0.962709
R18976 gnd.t306 gnd.n4671 0.956468
R18977 gnd.n4993 gnd.t236 0.956468
R18978 gnd.n5612 gnd.t226 0.956468
R18979 gnd.t319 gnd.n5556 0.956468
R18980 gnd.n7237 gnd.t82 0.956468
R18981 gnd.n7333 gnd.t30 0.956468
R18982 gnd.t2 gnd.n2962 0.912001
R18983 gnd.n3141 gnd.t275 0.912001
R18984 gnd.n2391 gnd.t351 0.912001
R18985 gnd.n4240 gnd.t65 0.912001
R18986 gnd.n4413 gnd.t36 0.912001
R18987 gnd.n2509 gnd.n2507 0.773756
R18988 gnd.n70 gnd.n68 0.773756
R18989 gnd.n2516 gnd.n2515 0.773756
R18990 gnd.n2515 gnd.n2513 0.773756
R18991 gnd.n2513 gnd.n2511 0.773756
R18992 gnd.n2511 gnd.n2509 0.773756
R18993 gnd.n2507 gnd.n2505 0.773756
R18994 gnd.n2505 gnd.n2503 0.773756
R18995 gnd.n2503 gnd.n2501 0.773756
R18996 gnd.n2501 gnd.n2499 0.773756
R18997 gnd.n62 gnd.n60 0.773756
R18998 gnd.n64 gnd.n62 0.773756
R18999 gnd.n66 gnd.n64 0.773756
R19000 gnd.n68 gnd.n66 0.773756
R19001 gnd.n72 gnd.n70 0.773756
R19002 gnd.n74 gnd.n72 0.773756
R19003 gnd.n76 gnd.n74 0.773756
R19004 gnd.n77 gnd.n76 0.773756
R19005 gnd gnd.n0 0.70738
R19006 gnd.n2 gnd.n1 0.672012
R19007 gnd.n3 gnd.n2 0.672012
R19008 gnd.n4 gnd.n3 0.672012
R19009 gnd.n5 gnd.n4 0.672012
R19010 gnd.n6 gnd.n5 0.672012
R19011 gnd.n7 gnd.n6 0.672012
R19012 gnd.n8 gnd.n7 0.672012
R19013 gnd.n9 gnd.n8 0.672012
R19014 gnd.n11 gnd.n10 0.672012
R19015 gnd.n12 gnd.n11 0.672012
R19016 gnd.n13 gnd.n12 0.672012
R19017 gnd.n14 gnd.n13 0.672012
R19018 gnd.n15 gnd.n14 0.672012
R19019 gnd.n16 gnd.n15 0.672012
R19020 gnd.n17 gnd.n16 0.672012
R19021 gnd.n18 gnd.n17 0.672012
R19022 gnd.n4965 gnd.t125 0.637812
R19023 gnd.n4945 gnd.n4944 0.637812
R19024 gnd.n5066 gnd.n5065 0.637812
R19025 gnd.n5065 gnd.t63 0.637812
R19026 gnd.n5149 gnd.n5148 0.637812
R19027 gnd.n5243 gnd.n5241 0.637812
R19028 gnd.n5260 gnd.t60 0.637812
R19029 gnd.n5334 gnd.t64 0.637812
R19030 gnd.n5327 gnd.n5326 0.637812
R19031 gnd.n5405 gnd.n5404 0.637812
R19032 gnd.n5472 gnd.t43 0.637812
R19033 gnd.n5472 gnd.n5471 0.637812
R19034 gnd.n5586 gnd.n5585 0.637812
R19035 gnd.n5640 gnd.t118 0.637812
R19036 gnd.n7608 gnd.n7607 0.637193
R19037 gnd.n2477 gnd.n2476 0.573776
R19038 gnd.n2476 gnd.n2474 0.573776
R19039 gnd.n2474 gnd.n2472 0.573776
R19040 gnd.n2472 gnd.n2470 0.573776
R19041 gnd.n2470 gnd.n2468 0.573776
R19042 gnd.n2468 gnd.n2466 0.573776
R19043 gnd.n2466 gnd.n2464 0.573776
R19044 gnd.n2464 gnd.n2462 0.573776
R19045 gnd.n2462 gnd.n2460 0.573776
R19046 gnd.n2496 gnd.n2495 0.573776
R19047 gnd.n2495 gnd.n2493 0.573776
R19048 gnd.n2493 gnd.n2491 0.573776
R19049 gnd.n2491 gnd.n2489 0.573776
R19050 gnd.n2489 gnd.n2487 0.573776
R19051 gnd.n2487 gnd.n2485 0.573776
R19052 gnd.n2485 gnd.n2483 0.573776
R19053 gnd.n2483 gnd.n2481 0.573776
R19054 gnd.n2481 gnd.n2479 0.573776
R19055 gnd.n23 gnd.n21 0.573776
R19056 gnd.n25 gnd.n23 0.573776
R19057 gnd.n27 gnd.n25 0.573776
R19058 gnd.n29 gnd.n27 0.573776
R19059 gnd.n31 gnd.n29 0.573776
R19060 gnd.n33 gnd.n31 0.573776
R19061 gnd.n35 gnd.n33 0.573776
R19062 gnd.n37 gnd.n35 0.573776
R19063 gnd.n38 gnd.n37 0.573776
R19064 gnd.n42 gnd.n40 0.573776
R19065 gnd.n44 gnd.n42 0.573776
R19066 gnd.n46 gnd.n44 0.573776
R19067 gnd.n48 gnd.n46 0.573776
R19068 gnd.n50 gnd.n48 0.573776
R19069 gnd.n52 gnd.n50 0.573776
R19070 gnd.n54 gnd.n52 0.573776
R19071 gnd.n56 gnd.n54 0.573776
R19072 gnd.n57 gnd.n56 0.573776
R19073 gnd.n3050 gnd.t321 0.547401
R19074 gnd.n3215 gnd.t274 0.547401
R19075 gnd.n4272 gnd.t85 0.547401
R19076 gnd.n4368 gnd.t16 0.547401
R19077 gnd.n3277 gnd.n2298 0.486781
R19078 gnd.n1225 gnd.n455 0.486781
R19079 gnd.n2853 gnd.n2852 0.48678
R19080 gnd.n6054 gnd.n6053 0.485256
R19081 gnd.n3594 gnd.n2252 0.480683
R19082 gnd.n2937 gnd.n2936 0.480683
R19083 gnd.n4152 gnd.n4147 0.477634
R19084 gnd.n4189 gnd.n4188 0.477634
R19085 gnd.n7456 gnd.n7455 0.477634
R19086 gnd.n7558 gnd.n7557 0.477634
R19087 gnd.n7550 gnd.n7549 0.465439
R19088 gnd.n7479 gnd.n7478 0.465439
R19089 gnd.n7031 gnd.n7028 0.465439
R19090 gnd.n7160 gnd.n448 0.465439
R19091 gnd.n4195 gnd.n2225 0.465439
R19092 gnd.n3845 gnd.n3844 0.465439
R19093 gnd.n1915 gnd.n1914 0.465439
R19094 gnd.n4788 gnd.n4787 0.465439
R19095 gnd.n5887 gnd.n5886 0.451719
R19096 gnd.n4700 gnd.n4699 0.451719
R19097 gnd.n6251 gnd.n6250 0.416659
R19098 gnd.n6573 gnd.n6572 0.416659
R19099 gnd.n6785 gnd.n604 0.416659
R19100 gnd.n4457 gnd.n1053 0.416659
R19101 gnd.n4575 gnd.n4571 0.388379
R19102 gnd.n7519 gnd.n7518 0.388379
R19103 gnd.n3554 gnd.n3553 0.388379
R19104 gnd.n3522 gnd.n3521 0.388379
R19105 gnd.n3490 gnd.n3489 0.388379
R19106 gnd.n3459 gnd.n3458 0.388379
R19107 gnd.n3427 gnd.n3426 0.388379
R19108 gnd.n3395 gnd.n3394 0.388379
R19109 gnd.n3363 gnd.n3362 0.388379
R19110 gnd.n3332 gnd.n3331 0.388379
R19111 gnd.n3791 gnd.n3733 0.388379
R19112 gnd.n1293 gnd.n1292 0.388379
R19113 gnd.n6056 gnd.n6055 0.378829
R19114 gnd.n7154 gnd.n7153 0.377553
R19115 gnd.n7608 gnd.n19 0.374463
R19116 gnd gnd.n7608 0.367492
R19117 gnd.n5184 gnd.t22 0.319156
R19118 gnd.t55 gnd.t24 0.319156
R19119 gnd.t358 gnd.t58 0.319156
R19120 gnd.t315 gnd.n1521 0.319156
R19121 gnd.n7269 gnd.t214 0.319156
R19122 gnd.n7301 gnd.t210 0.319156
R19123 gnd.n2771 gnd.n2749 0.311721
R19124 gnd.n3665 gnd.n3664 0.268793
R19125 gnd.n4777 gnd.n4448 0.247451
R19126 gnd.n1281 gnd.n591 0.247451
R19127 gnd.n3664 gnd.n3663 0.241354
R19128 gnd.n558 gnd.n555 0.229039
R19129 gnd.n561 gnd.n558 0.229039
R19130 gnd.n4827 gnd.n1900 0.229039
R19131 gnd.n4827 gnd.n4826 0.229039
R19132 gnd.n2518 gnd.n0 0.210825
R19133 gnd.n2925 gnd.n2724 0.206293
R19134 gnd.n2353 gnd.t270 0.1828
R19135 gnd.n4304 gnd.t26 0.1828
R19136 gnd.n4336 gnd.t69 0.1828
R19137 gnd.n3571 gnd.n3543 0.155672
R19138 gnd.n3564 gnd.n3543 0.155672
R19139 gnd.n3564 gnd.n3563 0.155672
R19140 gnd.n3563 gnd.n3547 0.155672
R19141 gnd.n3556 gnd.n3547 0.155672
R19142 gnd.n3556 gnd.n3555 0.155672
R19143 gnd.n3539 gnd.n3511 0.155672
R19144 gnd.n3532 gnd.n3511 0.155672
R19145 gnd.n3532 gnd.n3531 0.155672
R19146 gnd.n3531 gnd.n3515 0.155672
R19147 gnd.n3524 gnd.n3515 0.155672
R19148 gnd.n3524 gnd.n3523 0.155672
R19149 gnd.n3507 gnd.n3479 0.155672
R19150 gnd.n3500 gnd.n3479 0.155672
R19151 gnd.n3500 gnd.n3499 0.155672
R19152 gnd.n3499 gnd.n3483 0.155672
R19153 gnd.n3492 gnd.n3483 0.155672
R19154 gnd.n3492 gnd.n3491 0.155672
R19155 gnd.n3476 gnd.n3448 0.155672
R19156 gnd.n3469 gnd.n3448 0.155672
R19157 gnd.n3469 gnd.n3468 0.155672
R19158 gnd.n3468 gnd.n3452 0.155672
R19159 gnd.n3461 gnd.n3452 0.155672
R19160 gnd.n3461 gnd.n3460 0.155672
R19161 gnd.n3444 gnd.n3416 0.155672
R19162 gnd.n3437 gnd.n3416 0.155672
R19163 gnd.n3437 gnd.n3436 0.155672
R19164 gnd.n3436 gnd.n3420 0.155672
R19165 gnd.n3429 gnd.n3420 0.155672
R19166 gnd.n3429 gnd.n3428 0.155672
R19167 gnd.n3412 gnd.n3384 0.155672
R19168 gnd.n3405 gnd.n3384 0.155672
R19169 gnd.n3405 gnd.n3404 0.155672
R19170 gnd.n3404 gnd.n3388 0.155672
R19171 gnd.n3397 gnd.n3388 0.155672
R19172 gnd.n3397 gnd.n3396 0.155672
R19173 gnd.n3380 gnd.n3352 0.155672
R19174 gnd.n3373 gnd.n3352 0.155672
R19175 gnd.n3373 gnd.n3372 0.155672
R19176 gnd.n3372 gnd.n3356 0.155672
R19177 gnd.n3365 gnd.n3356 0.155672
R19178 gnd.n3365 gnd.n3364 0.155672
R19179 gnd.n3349 gnd.n3321 0.155672
R19180 gnd.n3342 gnd.n3321 0.155672
R19181 gnd.n3342 gnd.n3341 0.155672
R19182 gnd.n3341 gnd.n3325 0.155672
R19183 gnd.n3334 gnd.n3325 0.155672
R19184 gnd.n3334 gnd.n3333 0.155672
R19185 gnd.n7306 gnd.n7305 0.152939
R19186 gnd.n7306 gnd.n286 0.152939
R19187 gnd.n7320 gnd.n286 0.152939
R19188 gnd.n7321 gnd.n7320 0.152939
R19189 gnd.n7322 gnd.n7321 0.152939
R19190 gnd.n7322 gnd.n272 0.152939
R19191 gnd.n7336 gnd.n272 0.152939
R19192 gnd.n7337 gnd.n7336 0.152939
R19193 gnd.n7338 gnd.n7337 0.152939
R19194 gnd.n7338 gnd.n256 0.152939
R19195 gnd.n7352 gnd.n256 0.152939
R19196 gnd.n7353 gnd.n7352 0.152939
R19197 gnd.n7354 gnd.n7353 0.152939
R19198 gnd.n7354 gnd.n242 0.152939
R19199 gnd.n7368 gnd.n242 0.152939
R19200 gnd.n7369 gnd.n7368 0.152939
R19201 gnd.n7370 gnd.n7369 0.152939
R19202 gnd.n7370 gnd.n226 0.152939
R19203 gnd.n7384 gnd.n226 0.152939
R19204 gnd.n7385 gnd.n7384 0.152939
R19205 gnd.n7386 gnd.n7385 0.152939
R19206 gnd.n7386 gnd.n210 0.152939
R19207 gnd.n7468 gnd.n210 0.152939
R19208 gnd.n7469 gnd.n7468 0.152939
R19209 gnd.n7470 gnd.n7469 0.152939
R19210 gnd.n7470 gnd.n133 0.152939
R19211 gnd.n7550 gnd.n133 0.152939
R19212 gnd.n7549 gnd.n134 0.152939
R19213 gnd.n136 gnd.n134 0.152939
R19214 gnd.n140 gnd.n136 0.152939
R19215 gnd.n141 gnd.n140 0.152939
R19216 gnd.n142 gnd.n141 0.152939
R19217 gnd.n143 gnd.n142 0.152939
R19218 gnd.n147 gnd.n143 0.152939
R19219 gnd.n148 gnd.n147 0.152939
R19220 gnd.n149 gnd.n148 0.152939
R19221 gnd.n150 gnd.n149 0.152939
R19222 gnd.n154 gnd.n150 0.152939
R19223 gnd.n155 gnd.n154 0.152939
R19224 gnd.n156 gnd.n155 0.152939
R19225 gnd.n157 gnd.n156 0.152939
R19226 gnd.n161 gnd.n157 0.152939
R19227 gnd.n162 gnd.n161 0.152939
R19228 gnd.n163 gnd.n162 0.152939
R19229 gnd.n164 gnd.n163 0.152939
R19230 gnd.n168 gnd.n164 0.152939
R19231 gnd.n169 gnd.n168 0.152939
R19232 gnd.n170 gnd.n169 0.152939
R19233 gnd.n171 gnd.n170 0.152939
R19234 gnd.n175 gnd.n171 0.152939
R19235 gnd.n176 gnd.n175 0.152939
R19236 gnd.n177 gnd.n176 0.152939
R19237 gnd.n178 gnd.n177 0.152939
R19238 gnd.n182 gnd.n178 0.152939
R19239 gnd.n183 gnd.n182 0.152939
R19240 gnd.n184 gnd.n183 0.152939
R19241 gnd.n185 gnd.n184 0.152939
R19242 gnd.n189 gnd.n185 0.152939
R19243 gnd.n190 gnd.n189 0.152939
R19244 gnd.n191 gnd.n190 0.152939
R19245 gnd.n192 gnd.n191 0.152939
R19246 gnd.n196 gnd.n192 0.152939
R19247 gnd.n197 gnd.n196 0.152939
R19248 gnd.n7480 gnd.n197 0.152939
R19249 gnd.n7480 gnd.n7479 0.152939
R19250 gnd.n7028 gnd.n584 0.152939
R19251 gnd.n586 gnd.n584 0.152939
R19252 gnd.n587 gnd.n586 0.152939
R19253 gnd.n6812 gnd.n587 0.152939
R19254 gnd.n6813 gnd.n6812 0.152939
R19255 gnd.n6813 gnd.n6811 0.152939
R19256 gnd.n6821 gnd.n6811 0.152939
R19257 gnd.n6822 gnd.n6821 0.152939
R19258 gnd.n6823 gnd.n6822 0.152939
R19259 gnd.n6824 gnd.n6823 0.152939
R19260 gnd.n6825 gnd.n6824 0.152939
R19261 gnd.n6826 gnd.n6825 0.152939
R19262 gnd.n6827 gnd.n6826 0.152939
R19263 gnd.n6828 gnd.n6827 0.152939
R19264 gnd.n6829 gnd.n6828 0.152939
R19265 gnd.n6830 gnd.n6829 0.152939
R19266 gnd.n6831 gnd.n6830 0.152939
R19267 gnd.n6832 gnd.n6831 0.152939
R19268 gnd.n6833 gnd.n6832 0.152939
R19269 gnd.n6834 gnd.n6833 0.152939
R19270 gnd.n6835 gnd.n6834 0.152939
R19271 gnd.n6836 gnd.n6835 0.152939
R19272 gnd.n6837 gnd.n6836 0.152939
R19273 gnd.n6838 gnd.n6837 0.152939
R19274 gnd.n6839 gnd.n6838 0.152939
R19275 gnd.n6840 gnd.n6839 0.152939
R19276 gnd.n6841 gnd.n6840 0.152939
R19277 gnd.n6842 gnd.n6841 0.152939
R19278 gnd.n6843 gnd.n6842 0.152939
R19279 gnd.n6844 gnd.n6843 0.152939
R19280 gnd.n6845 gnd.n6844 0.152939
R19281 gnd.n6845 gnd.n325 0.152939
R19282 gnd.n6846 gnd.n325 0.152939
R19283 gnd.n6847 gnd.n6846 0.152939
R19284 gnd.n6848 gnd.n6847 0.152939
R19285 gnd.n6849 gnd.n6848 0.152939
R19286 gnd.n6850 gnd.n6849 0.152939
R19287 gnd.n6851 gnd.n6850 0.152939
R19288 gnd.n6852 gnd.n6851 0.152939
R19289 gnd.n6853 gnd.n6852 0.152939
R19290 gnd.n6854 gnd.n6853 0.152939
R19291 gnd.n6855 gnd.n6854 0.152939
R19292 gnd.n6856 gnd.n6855 0.152939
R19293 gnd.n6857 gnd.n6856 0.152939
R19294 gnd.n6858 gnd.n6857 0.152939
R19295 gnd.n6859 gnd.n6858 0.152939
R19296 gnd.n6860 gnd.n6859 0.152939
R19297 gnd.n6861 gnd.n6860 0.152939
R19298 gnd.n6862 gnd.n6861 0.152939
R19299 gnd.n6863 gnd.n6862 0.152939
R19300 gnd.n6864 gnd.n6863 0.152939
R19301 gnd.n6865 gnd.n6864 0.152939
R19302 gnd.n6866 gnd.n6865 0.152939
R19303 gnd.n6867 gnd.n6866 0.152939
R19304 gnd.n6868 gnd.n6867 0.152939
R19305 gnd.n6869 gnd.n6868 0.152939
R19306 gnd.n6870 gnd.n6869 0.152939
R19307 gnd.n6871 gnd.n6870 0.152939
R19308 gnd.n6872 gnd.n6871 0.152939
R19309 gnd.n6873 gnd.n6872 0.152939
R19310 gnd.n6875 gnd.n6873 0.152939
R19311 gnd.n6875 gnd.n6874 0.152939
R19312 gnd.n6874 gnd.n203 0.152939
R19313 gnd.n7478 gnd.n203 0.152939
R19314 gnd.n541 gnd.n448 0.152939
R19315 gnd.n542 gnd.n541 0.152939
R19316 gnd.n543 gnd.n542 0.152939
R19317 gnd.n544 gnd.n543 0.152939
R19318 gnd.n545 gnd.n544 0.152939
R19319 gnd.n546 gnd.n545 0.152939
R19320 gnd.n547 gnd.n546 0.152939
R19321 gnd.n548 gnd.n547 0.152939
R19322 gnd.n549 gnd.n548 0.152939
R19323 gnd.n550 gnd.n549 0.152939
R19324 gnd.n551 gnd.n550 0.152939
R19325 gnd.n552 gnd.n551 0.152939
R19326 gnd.n553 gnd.n552 0.152939
R19327 gnd.n554 gnd.n553 0.152939
R19328 gnd.n555 gnd.n554 0.152939
R19329 gnd.n562 gnd.n561 0.152939
R19330 gnd.n563 gnd.n562 0.152939
R19331 gnd.n564 gnd.n563 0.152939
R19332 gnd.n565 gnd.n564 0.152939
R19333 gnd.n566 gnd.n565 0.152939
R19334 gnd.n567 gnd.n566 0.152939
R19335 gnd.n568 gnd.n567 0.152939
R19336 gnd.n569 gnd.n568 0.152939
R19337 gnd.n570 gnd.n569 0.152939
R19338 gnd.n571 gnd.n570 0.152939
R19339 gnd.n572 gnd.n571 0.152939
R19340 gnd.n573 gnd.n572 0.152939
R19341 gnd.n574 gnd.n573 0.152939
R19342 gnd.n575 gnd.n574 0.152939
R19343 gnd.n576 gnd.n575 0.152939
R19344 gnd.n577 gnd.n576 0.152939
R19345 gnd.n578 gnd.n577 0.152939
R19346 gnd.n7033 gnd.n578 0.152939
R19347 gnd.n7033 gnd.n7032 0.152939
R19348 gnd.n7032 gnd.n7031 0.152939
R19349 gnd.n7161 gnd.n7160 0.152939
R19350 gnd.n7162 gnd.n7161 0.152939
R19351 gnd.n7162 gnd.n431 0.152939
R19352 gnd.n7176 gnd.n431 0.152939
R19353 gnd.n7177 gnd.n7176 0.152939
R19354 gnd.n7178 gnd.n7177 0.152939
R19355 gnd.n7178 gnd.n413 0.152939
R19356 gnd.n7192 gnd.n413 0.152939
R19357 gnd.n7193 gnd.n7192 0.152939
R19358 gnd.n7194 gnd.n7193 0.152939
R19359 gnd.n7194 gnd.n398 0.152939
R19360 gnd.n7208 gnd.n398 0.152939
R19361 gnd.n7209 gnd.n7208 0.152939
R19362 gnd.n7210 gnd.n7209 0.152939
R19363 gnd.n7210 gnd.n381 0.152939
R19364 gnd.n7224 gnd.n381 0.152939
R19365 gnd.n7225 gnd.n7224 0.152939
R19366 gnd.n7226 gnd.n7225 0.152939
R19367 gnd.n7226 gnd.n366 0.152939
R19368 gnd.n7240 gnd.n366 0.152939
R19369 gnd.n7241 gnd.n7240 0.152939
R19370 gnd.n7242 gnd.n7241 0.152939
R19371 gnd.n7242 gnd.n349 0.152939
R19372 gnd.n7256 gnd.n349 0.152939
R19373 gnd.n7257 gnd.n7256 0.152939
R19374 gnd.n7258 gnd.n7257 0.152939
R19375 gnd.n7258 gnd.n334 0.152939
R19376 gnd.n6252 gnd.n6251 0.152939
R19377 gnd.n6252 gnd.n918 0.152939
R19378 gnd.n6260 gnd.n918 0.152939
R19379 gnd.n6261 gnd.n6260 0.152939
R19380 gnd.n6262 gnd.n6261 0.152939
R19381 gnd.n6262 gnd.n912 0.152939
R19382 gnd.n6270 gnd.n912 0.152939
R19383 gnd.n6271 gnd.n6270 0.152939
R19384 gnd.n6272 gnd.n6271 0.152939
R19385 gnd.n6272 gnd.n906 0.152939
R19386 gnd.n6280 gnd.n906 0.152939
R19387 gnd.n6281 gnd.n6280 0.152939
R19388 gnd.n6282 gnd.n6281 0.152939
R19389 gnd.n6282 gnd.n900 0.152939
R19390 gnd.n6290 gnd.n900 0.152939
R19391 gnd.n6291 gnd.n6290 0.152939
R19392 gnd.n6292 gnd.n6291 0.152939
R19393 gnd.n6292 gnd.n894 0.152939
R19394 gnd.n6300 gnd.n894 0.152939
R19395 gnd.n6301 gnd.n6300 0.152939
R19396 gnd.n6302 gnd.n6301 0.152939
R19397 gnd.n6302 gnd.n888 0.152939
R19398 gnd.n6310 gnd.n888 0.152939
R19399 gnd.n6311 gnd.n6310 0.152939
R19400 gnd.n6312 gnd.n6311 0.152939
R19401 gnd.n6312 gnd.n882 0.152939
R19402 gnd.n6320 gnd.n882 0.152939
R19403 gnd.n6321 gnd.n6320 0.152939
R19404 gnd.n6322 gnd.n6321 0.152939
R19405 gnd.n6322 gnd.n876 0.152939
R19406 gnd.n6330 gnd.n876 0.152939
R19407 gnd.n6331 gnd.n6330 0.152939
R19408 gnd.n6332 gnd.n6331 0.152939
R19409 gnd.n6332 gnd.n870 0.152939
R19410 gnd.n6340 gnd.n870 0.152939
R19411 gnd.n6341 gnd.n6340 0.152939
R19412 gnd.n6342 gnd.n6341 0.152939
R19413 gnd.n6342 gnd.n864 0.152939
R19414 gnd.n6350 gnd.n864 0.152939
R19415 gnd.n6351 gnd.n6350 0.152939
R19416 gnd.n6352 gnd.n6351 0.152939
R19417 gnd.n6352 gnd.n858 0.152939
R19418 gnd.n6360 gnd.n858 0.152939
R19419 gnd.n6361 gnd.n6360 0.152939
R19420 gnd.n6362 gnd.n6361 0.152939
R19421 gnd.n6362 gnd.n852 0.152939
R19422 gnd.n6370 gnd.n852 0.152939
R19423 gnd.n6371 gnd.n6370 0.152939
R19424 gnd.n6372 gnd.n6371 0.152939
R19425 gnd.n6372 gnd.n846 0.152939
R19426 gnd.n6380 gnd.n846 0.152939
R19427 gnd.n6381 gnd.n6380 0.152939
R19428 gnd.n6382 gnd.n6381 0.152939
R19429 gnd.n6382 gnd.n840 0.152939
R19430 gnd.n6390 gnd.n840 0.152939
R19431 gnd.n6391 gnd.n6390 0.152939
R19432 gnd.n6392 gnd.n6391 0.152939
R19433 gnd.n6392 gnd.n834 0.152939
R19434 gnd.n6400 gnd.n834 0.152939
R19435 gnd.n6401 gnd.n6400 0.152939
R19436 gnd.n6402 gnd.n6401 0.152939
R19437 gnd.n6402 gnd.n828 0.152939
R19438 gnd.n6410 gnd.n828 0.152939
R19439 gnd.n6411 gnd.n6410 0.152939
R19440 gnd.n6412 gnd.n6411 0.152939
R19441 gnd.n6412 gnd.n822 0.152939
R19442 gnd.n6420 gnd.n822 0.152939
R19443 gnd.n6421 gnd.n6420 0.152939
R19444 gnd.n6422 gnd.n6421 0.152939
R19445 gnd.n6422 gnd.n816 0.152939
R19446 gnd.n6430 gnd.n816 0.152939
R19447 gnd.n6431 gnd.n6430 0.152939
R19448 gnd.n6432 gnd.n6431 0.152939
R19449 gnd.n6432 gnd.n810 0.152939
R19450 gnd.n6440 gnd.n810 0.152939
R19451 gnd.n6441 gnd.n6440 0.152939
R19452 gnd.n6442 gnd.n6441 0.152939
R19453 gnd.n6442 gnd.n804 0.152939
R19454 gnd.n6450 gnd.n804 0.152939
R19455 gnd.n6451 gnd.n6450 0.152939
R19456 gnd.n6452 gnd.n6451 0.152939
R19457 gnd.n6452 gnd.n798 0.152939
R19458 gnd.n6460 gnd.n798 0.152939
R19459 gnd.n6461 gnd.n6460 0.152939
R19460 gnd.n6462 gnd.n6461 0.152939
R19461 gnd.n6462 gnd.n792 0.152939
R19462 gnd.n6470 gnd.n792 0.152939
R19463 gnd.n6471 gnd.n6470 0.152939
R19464 gnd.n6472 gnd.n6471 0.152939
R19465 gnd.n6472 gnd.n786 0.152939
R19466 gnd.n6480 gnd.n786 0.152939
R19467 gnd.n6481 gnd.n6480 0.152939
R19468 gnd.n6482 gnd.n6481 0.152939
R19469 gnd.n6482 gnd.n780 0.152939
R19470 gnd.n6490 gnd.n780 0.152939
R19471 gnd.n6491 gnd.n6490 0.152939
R19472 gnd.n6492 gnd.n6491 0.152939
R19473 gnd.n6492 gnd.n774 0.152939
R19474 gnd.n6500 gnd.n774 0.152939
R19475 gnd.n6501 gnd.n6500 0.152939
R19476 gnd.n6502 gnd.n6501 0.152939
R19477 gnd.n6502 gnd.n768 0.152939
R19478 gnd.n6510 gnd.n768 0.152939
R19479 gnd.n6511 gnd.n6510 0.152939
R19480 gnd.n6512 gnd.n6511 0.152939
R19481 gnd.n6512 gnd.n762 0.152939
R19482 gnd.n6520 gnd.n762 0.152939
R19483 gnd.n6521 gnd.n6520 0.152939
R19484 gnd.n6522 gnd.n6521 0.152939
R19485 gnd.n6522 gnd.n756 0.152939
R19486 gnd.n6530 gnd.n756 0.152939
R19487 gnd.n6531 gnd.n6530 0.152939
R19488 gnd.n6532 gnd.n6531 0.152939
R19489 gnd.n6532 gnd.n750 0.152939
R19490 gnd.n6540 gnd.n750 0.152939
R19491 gnd.n6541 gnd.n6540 0.152939
R19492 gnd.n6542 gnd.n6541 0.152939
R19493 gnd.n6542 gnd.n744 0.152939
R19494 gnd.n6550 gnd.n744 0.152939
R19495 gnd.n6551 gnd.n6550 0.152939
R19496 gnd.n6552 gnd.n6551 0.152939
R19497 gnd.n6552 gnd.n738 0.152939
R19498 gnd.n6560 gnd.n738 0.152939
R19499 gnd.n6561 gnd.n6560 0.152939
R19500 gnd.n6563 gnd.n6561 0.152939
R19501 gnd.n6563 gnd.n6562 0.152939
R19502 gnd.n6562 gnd.n732 0.152939
R19503 gnd.n6572 gnd.n732 0.152939
R19504 gnd.n6573 gnd.n727 0.152939
R19505 gnd.n6581 gnd.n727 0.152939
R19506 gnd.n6582 gnd.n6581 0.152939
R19507 gnd.n6583 gnd.n6582 0.152939
R19508 gnd.n6583 gnd.n721 0.152939
R19509 gnd.n6591 gnd.n721 0.152939
R19510 gnd.n6592 gnd.n6591 0.152939
R19511 gnd.n6593 gnd.n6592 0.152939
R19512 gnd.n6593 gnd.n715 0.152939
R19513 gnd.n6601 gnd.n715 0.152939
R19514 gnd.n6602 gnd.n6601 0.152939
R19515 gnd.n6603 gnd.n6602 0.152939
R19516 gnd.n6603 gnd.n709 0.152939
R19517 gnd.n6611 gnd.n709 0.152939
R19518 gnd.n6612 gnd.n6611 0.152939
R19519 gnd.n6613 gnd.n6612 0.152939
R19520 gnd.n6613 gnd.n703 0.152939
R19521 gnd.n6621 gnd.n703 0.152939
R19522 gnd.n6622 gnd.n6621 0.152939
R19523 gnd.n6623 gnd.n6622 0.152939
R19524 gnd.n6623 gnd.n697 0.152939
R19525 gnd.n6631 gnd.n697 0.152939
R19526 gnd.n6632 gnd.n6631 0.152939
R19527 gnd.n6633 gnd.n6632 0.152939
R19528 gnd.n6633 gnd.n691 0.152939
R19529 gnd.n6641 gnd.n691 0.152939
R19530 gnd.n6642 gnd.n6641 0.152939
R19531 gnd.n6643 gnd.n6642 0.152939
R19532 gnd.n6643 gnd.n685 0.152939
R19533 gnd.n6651 gnd.n685 0.152939
R19534 gnd.n6652 gnd.n6651 0.152939
R19535 gnd.n6653 gnd.n6652 0.152939
R19536 gnd.n6653 gnd.n679 0.152939
R19537 gnd.n6661 gnd.n679 0.152939
R19538 gnd.n6662 gnd.n6661 0.152939
R19539 gnd.n6663 gnd.n6662 0.152939
R19540 gnd.n6663 gnd.n673 0.152939
R19541 gnd.n6671 gnd.n673 0.152939
R19542 gnd.n6672 gnd.n6671 0.152939
R19543 gnd.n6673 gnd.n6672 0.152939
R19544 gnd.n6673 gnd.n667 0.152939
R19545 gnd.n6681 gnd.n667 0.152939
R19546 gnd.n6682 gnd.n6681 0.152939
R19547 gnd.n6683 gnd.n6682 0.152939
R19548 gnd.n6683 gnd.n661 0.152939
R19549 gnd.n6691 gnd.n661 0.152939
R19550 gnd.n6692 gnd.n6691 0.152939
R19551 gnd.n6693 gnd.n6692 0.152939
R19552 gnd.n6693 gnd.n655 0.152939
R19553 gnd.n6701 gnd.n655 0.152939
R19554 gnd.n6702 gnd.n6701 0.152939
R19555 gnd.n6703 gnd.n6702 0.152939
R19556 gnd.n6703 gnd.n649 0.152939
R19557 gnd.n6711 gnd.n649 0.152939
R19558 gnd.n6712 gnd.n6711 0.152939
R19559 gnd.n6713 gnd.n6712 0.152939
R19560 gnd.n6713 gnd.n643 0.152939
R19561 gnd.n6721 gnd.n643 0.152939
R19562 gnd.n6722 gnd.n6721 0.152939
R19563 gnd.n6723 gnd.n6722 0.152939
R19564 gnd.n6723 gnd.n637 0.152939
R19565 gnd.n6731 gnd.n637 0.152939
R19566 gnd.n6732 gnd.n6731 0.152939
R19567 gnd.n6733 gnd.n6732 0.152939
R19568 gnd.n6733 gnd.n631 0.152939
R19569 gnd.n6741 gnd.n631 0.152939
R19570 gnd.n6742 gnd.n6741 0.152939
R19571 gnd.n6743 gnd.n6742 0.152939
R19572 gnd.n6743 gnd.n625 0.152939
R19573 gnd.n6751 gnd.n625 0.152939
R19574 gnd.n6752 gnd.n6751 0.152939
R19575 gnd.n6753 gnd.n6752 0.152939
R19576 gnd.n6753 gnd.n619 0.152939
R19577 gnd.n6761 gnd.n619 0.152939
R19578 gnd.n6762 gnd.n6761 0.152939
R19579 gnd.n6763 gnd.n6762 0.152939
R19580 gnd.n6763 gnd.n613 0.152939
R19581 gnd.n6771 gnd.n613 0.152939
R19582 gnd.n6772 gnd.n6771 0.152939
R19583 gnd.n6773 gnd.n6772 0.152939
R19584 gnd.n6773 gnd.n607 0.152939
R19585 gnd.n6783 gnd.n607 0.152939
R19586 gnd.n6784 gnd.n6783 0.152939
R19587 gnd.n6785 gnd.n6784 0.152939
R19588 gnd.n4458 gnd.n4457 0.152939
R19589 gnd.n4462 gnd.n4458 0.152939
R19590 gnd.n4463 gnd.n4462 0.152939
R19591 gnd.n4464 gnd.n4463 0.152939
R19592 gnd.n4464 gnd.n4453 0.152939
R19593 gnd.n4470 gnd.n4453 0.152939
R19594 gnd.n4471 gnd.n4470 0.152939
R19595 gnd.n4472 gnd.n4471 0.152939
R19596 gnd.n4473 gnd.n4472 0.152939
R19597 gnd.n4474 gnd.n4473 0.152939
R19598 gnd.n4615 gnd.n4474 0.152939
R19599 gnd.n4616 gnd.n4615 0.152939
R19600 gnd.n4616 gnd.n4613 0.152939
R19601 gnd.n4627 gnd.n4613 0.152939
R19602 gnd.n4628 gnd.n4627 0.152939
R19603 gnd.n4629 gnd.n4628 0.152939
R19604 gnd.n4629 gnd.n4607 0.152939
R19605 gnd.n4643 gnd.n4607 0.152939
R19606 gnd.n4644 gnd.n4643 0.152939
R19607 gnd.n4645 gnd.n4644 0.152939
R19608 gnd.n4645 gnd.n4601 0.152939
R19609 gnd.n4659 gnd.n4601 0.152939
R19610 gnd.n4660 gnd.n4659 0.152939
R19611 gnd.n4661 gnd.n4660 0.152939
R19612 gnd.n4661 gnd.n1769 0.152939
R19613 gnd.n4909 gnd.n1769 0.152939
R19614 gnd.n4910 gnd.n4909 0.152939
R19615 gnd.n4911 gnd.n4910 0.152939
R19616 gnd.n4911 gnd.n1748 0.152939
R19617 gnd.n4968 gnd.n1748 0.152939
R19618 gnd.n4969 gnd.n4968 0.152939
R19619 gnd.n4970 gnd.n4969 0.152939
R19620 gnd.n4970 gnd.n1725 0.152939
R19621 gnd.n4996 gnd.n1725 0.152939
R19622 gnd.n4997 gnd.n4996 0.152939
R19623 gnd.n4998 gnd.n4997 0.152939
R19624 gnd.n4999 gnd.n4998 0.152939
R19625 gnd.n4999 gnd.n1697 0.152939
R19626 gnd.n5070 gnd.n1697 0.152939
R19627 gnd.n5071 gnd.n5070 0.152939
R19628 gnd.n5072 gnd.n5071 0.152939
R19629 gnd.n5072 gnd.n1677 0.152939
R19630 gnd.n5095 gnd.n1677 0.152939
R19631 gnd.n5096 gnd.n5095 0.152939
R19632 gnd.n5097 gnd.n5096 0.152939
R19633 gnd.n5097 gnd.n1657 0.152939
R19634 gnd.n5129 gnd.n1657 0.152939
R19635 gnd.n5130 gnd.n5129 0.152939
R19636 gnd.n5131 gnd.n5130 0.152939
R19637 gnd.n5131 gnd.n1640 0.152939
R19638 gnd.n5174 gnd.n1640 0.152939
R19639 gnd.n5175 gnd.n5174 0.152939
R19640 gnd.n5176 gnd.n5175 0.152939
R19641 gnd.n5177 gnd.n5176 0.152939
R19642 gnd.n5177 gnd.n1612 0.152939
R19643 gnd.n5247 gnd.n1612 0.152939
R19644 gnd.n5248 gnd.n5247 0.152939
R19645 gnd.n5249 gnd.n5248 0.152939
R19646 gnd.n5249 gnd.n1592 0.152939
R19647 gnd.n5273 gnd.n1592 0.152939
R19648 gnd.n5274 gnd.n5273 0.152939
R19649 gnd.n5275 gnd.n5274 0.152939
R19650 gnd.n5275 gnd.n1569 0.152939
R19651 gnd.n5306 gnd.n1569 0.152939
R19652 gnd.n5307 gnd.n5306 0.152939
R19653 gnd.n5308 gnd.n5307 0.152939
R19654 gnd.n5308 gnd.n1552 0.152939
R19655 gnd.n5352 gnd.n1552 0.152939
R19656 gnd.n5353 gnd.n5352 0.152939
R19657 gnd.n5354 gnd.n5353 0.152939
R19658 gnd.n5355 gnd.n5354 0.152939
R19659 gnd.n5355 gnd.n1525 0.152939
R19660 gnd.n5409 gnd.n1525 0.152939
R19661 gnd.n5410 gnd.n5409 0.152939
R19662 gnd.n5411 gnd.n5410 0.152939
R19663 gnd.n5411 gnd.n1504 0.152939
R19664 gnd.n5434 gnd.n1504 0.152939
R19665 gnd.n5435 gnd.n5434 0.152939
R19666 gnd.n5436 gnd.n5435 0.152939
R19667 gnd.n5436 gnd.n1482 0.152939
R19668 gnd.n5495 gnd.n1482 0.152939
R19669 gnd.n5496 gnd.n5495 0.152939
R19670 gnd.n5497 gnd.n5496 0.152939
R19671 gnd.n5497 gnd.n1460 0.152939
R19672 gnd.n5524 gnd.n1460 0.152939
R19673 gnd.n5525 gnd.n5524 0.152939
R19674 gnd.n5526 gnd.n5525 0.152939
R19675 gnd.n5527 gnd.n5526 0.152939
R19676 gnd.n5527 gnd.n1433 0.152939
R19677 gnd.n5590 gnd.n1433 0.152939
R19678 gnd.n5591 gnd.n5590 0.152939
R19679 gnd.n5592 gnd.n5591 0.152939
R19680 gnd.n5592 gnd.n1413 0.152939
R19681 gnd.n5615 gnd.n1413 0.152939
R19682 gnd.n5616 gnd.n5615 0.152939
R19683 gnd.n5617 gnd.n5616 0.152939
R19684 gnd.n5617 gnd.n1393 0.152939
R19685 gnd.n5643 gnd.n1393 0.152939
R19686 gnd.n5644 gnd.n5643 0.152939
R19687 gnd.n5645 gnd.n5644 0.152939
R19688 gnd.n5646 gnd.n5645 0.152939
R19689 gnd.n5646 gnd.n1331 0.152939
R19690 gnd.n5832 gnd.n1331 0.152939
R19691 gnd.n5833 gnd.n5832 0.152939
R19692 gnd.n5834 gnd.n5833 0.152939
R19693 gnd.n5834 gnd.n1318 0.152939
R19694 gnd.n5852 gnd.n1318 0.152939
R19695 gnd.n5853 gnd.n5852 0.152939
R19696 gnd.n5854 gnd.n5853 0.152939
R19697 gnd.n5854 gnd.n1305 0.152939
R19698 gnd.n5875 gnd.n1305 0.152939
R19699 gnd.n5876 gnd.n5875 0.152939
R19700 gnd.n5878 gnd.n5876 0.152939
R19701 gnd.n5878 gnd.n5877 0.152939
R19702 gnd.n5877 gnd.n1233 0.152939
R19703 gnd.n1234 gnd.n1233 0.152939
R19704 gnd.n1235 gnd.n1234 0.152939
R19705 gnd.n1238 gnd.n1235 0.152939
R19706 gnd.n1239 gnd.n1238 0.152939
R19707 gnd.n1241 gnd.n1239 0.152939
R19708 gnd.n1241 gnd.n1240 0.152939
R19709 gnd.n1240 gnd.n596 0.152939
R19710 gnd.n597 gnd.n596 0.152939
R19711 gnd.n598 gnd.n597 0.152939
R19712 gnd.n601 gnd.n598 0.152939
R19713 gnd.n602 gnd.n601 0.152939
R19714 gnd.n603 gnd.n602 0.152939
R19715 gnd.n604 gnd.n603 0.152939
R19716 gnd.n6250 gnd.n924 0.152939
R19717 gnd.n971 gnd.n924 0.152939
R19718 gnd.n972 gnd.n971 0.152939
R19719 gnd.n973 gnd.n972 0.152939
R19720 gnd.n974 gnd.n973 0.152939
R19721 gnd.n975 gnd.n974 0.152939
R19722 gnd.n976 gnd.n975 0.152939
R19723 gnd.n977 gnd.n976 0.152939
R19724 gnd.n978 gnd.n977 0.152939
R19725 gnd.n979 gnd.n978 0.152939
R19726 gnd.n980 gnd.n979 0.152939
R19727 gnd.n981 gnd.n980 0.152939
R19728 gnd.n982 gnd.n981 0.152939
R19729 gnd.n983 gnd.n982 0.152939
R19730 gnd.n984 gnd.n983 0.152939
R19731 gnd.n985 gnd.n984 0.152939
R19732 gnd.n986 gnd.n985 0.152939
R19733 gnd.n987 gnd.n986 0.152939
R19734 gnd.n988 gnd.n987 0.152939
R19735 gnd.n989 gnd.n988 0.152939
R19736 gnd.n990 gnd.n989 0.152939
R19737 gnd.n991 gnd.n990 0.152939
R19738 gnd.n992 gnd.n991 0.152939
R19739 gnd.n993 gnd.n992 0.152939
R19740 gnd.n994 gnd.n993 0.152939
R19741 gnd.n995 gnd.n994 0.152939
R19742 gnd.n996 gnd.n995 0.152939
R19743 gnd.n997 gnd.n996 0.152939
R19744 gnd.n998 gnd.n997 0.152939
R19745 gnd.n999 gnd.n998 0.152939
R19746 gnd.n1000 gnd.n999 0.152939
R19747 gnd.n1001 gnd.n1000 0.152939
R19748 gnd.n1002 gnd.n1001 0.152939
R19749 gnd.n1003 gnd.n1002 0.152939
R19750 gnd.n1004 gnd.n1003 0.152939
R19751 gnd.n1005 gnd.n1004 0.152939
R19752 gnd.n1006 gnd.n1005 0.152939
R19753 gnd.n1007 gnd.n1006 0.152939
R19754 gnd.n1008 gnd.n1007 0.152939
R19755 gnd.n1009 gnd.n1008 0.152939
R19756 gnd.n1010 gnd.n1009 0.152939
R19757 gnd.n1011 gnd.n1010 0.152939
R19758 gnd.n1012 gnd.n1011 0.152939
R19759 gnd.n1013 gnd.n1012 0.152939
R19760 gnd.n1014 gnd.n1013 0.152939
R19761 gnd.n1015 gnd.n1014 0.152939
R19762 gnd.n1016 gnd.n1015 0.152939
R19763 gnd.n1017 gnd.n1016 0.152939
R19764 gnd.n1018 gnd.n1017 0.152939
R19765 gnd.n1019 gnd.n1018 0.152939
R19766 gnd.n1020 gnd.n1019 0.152939
R19767 gnd.n1021 gnd.n1020 0.152939
R19768 gnd.n1022 gnd.n1021 0.152939
R19769 gnd.n1023 gnd.n1022 0.152939
R19770 gnd.n1024 gnd.n1023 0.152939
R19771 gnd.n1025 gnd.n1024 0.152939
R19772 gnd.n1026 gnd.n1025 0.152939
R19773 gnd.n1027 gnd.n1026 0.152939
R19774 gnd.n1028 gnd.n1027 0.152939
R19775 gnd.n1029 gnd.n1028 0.152939
R19776 gnd.n1030 gnd.n1029 0.152939
R19777 gnd.n1031 gnd.n1030 0.152939
R19778 gnd.n1032 gnd.n1031 0.152939
R19779 gnd.n1033 gnd.n1032 0.152939
R19780 gnd.n1034 gnd.n1033 0.152939
R19781 gnd.n1035 gnd.n1034 0.152939
R19782 gnd.n1036 gnd.n1035 0.152939
R19783 gnd.n1037 gnd.n1036 0.152939
R19784 gnd.n1038 gnd.n1037 0.152939
R19785 gnd.n1039 gnd.n1038 0.152939
R19786 gnd.n1040 gnd.n1039 0.152939
R19787 gnd.n1041 gnd.n1040 0.152939
R19788 gnd.n1042 gnd.n1041 0.152939
R19789 gnd.n1043 gnd.n1042 0.152939
R19790 gnd.n1044 gnd.n1043 0.152939
R19791 gnd.n1045 gnd.n1044 0.152939
R19792 gnd.n1046 gnd.n1045 0.152939
R19793 gnd.n1047 gnd.n1046 0.152939
R19794 gnd.n1048 gnd.n1047 0.152939
R19795 gnd.n1049 gnd.n1048 0.152939
R19796 gnd.n1050 gnd.n1049 0.152939
R19797 gnd.n1051 gnd.n1050 0.152939
R19798 gnd.n1052 gnd.n1051 0.152939
R19799 gnd.n1053 gnd.n1052 0.152939
R19800 gnd.n3696 gnd.n2252 0.152939
R19801 gnd.n3696 gnd.n3695 0.152939
R19802 gnd.n3695 gnd.n3694 0.152939
R19803 gnd.n3694 gnd.n2254 0.152939
R19804 gnd.n2255 gnd.n2254 0.152939
R19805 gnd.n2256 gnd.n2255 0.152939
R19806 gnd.n2257 gnd.n2256 0.152939
R19807 gnd.n2258 gnd.n2257 0.152939
R19808 gnd.n2259 gnd.n2258 0.152939
R19809 gnd.n2260 gnd.n2259 0.152939
R19810 gnd.n2261 gnd.n2260 0.152939
R19811 gnd.n2262 gnd.n2261 0.152939
R19812 gnd.n2263 gnd.n2262 0.152939
R19813 gnd.n2264 gnd.n2263 0.152939
R19814 gnd.n3666 gnd.n2264 0.152939
R19815 gnd.n3666 gnd.n3665 0.152939
R19816 gnd.n2938 gnd.n2937 0.152939
R19817 gnd.n2938 gnd.n2642 0.152939
R19818 gnd.n2966 gnd.n2642 0.152939
R19819 gnd.n2967 gnd.n2966 0.152939
R19820 gnd.n2968 gnd.n2967 0.152939
R19821 gnd.n2969 gnd.n2968 0.152939
R19822 gnd.n2969 gnd.n2614 0.152939
R19823 gnd.n2996 gnd.n2614 0.152939
R19824 gnd.n2997 gnd.n2996 0.152939
R19825 gnd.n2998 gnd.n2997 0.152939
R19826 gnd.n2998 gnd.n2592 0.152939
R19827 gnd.n3027 gnd.n2592 0.152939
R19828 gnd.n3028 gnd.n3027 0.152939
R19829 gnd.n3029 gnd.n3028 0.152939
R19830 gnd.n3030 gnd.n3029 0.152939
R19831 gnd.n3032 gnd.n3030 0.152939
R19832 gnd.n3032 gnd.n3031 0.152939
R19833 gnd.n3031 gnd.n2541 0.152939
R19834 gnd.n2542 gnd.n2541 0.152939
R19835 gnd.n2543 gnd.n2542 0.152939
R19836 gnd.n2562 gnd.n2543 0.152939
R19837 gnd.n2563 gnd.n2562 0.152939
R19838 gnd.n2563 gnd.n2449 0.152939
R19839 gnd.n3122 gnd.n2449 0.152939
R19840 gnd.n3123 gnd.n3122 0.152939
R19841 gnd.n3124 gnd.n3123 0.152939
R19842 gnd.n3125 gnd.n3124 0.152939
R19843 gnd.n3125 gnd.n2422 0.152939
R19844 gnd.n3162 gnd.n2422 0.152939
R19845 gnd.n3163 gnd.n3162 0.152939
R19846 gnd.n3164 gnd.n3163 0.152939
R19847 gnd.n3165 gnd.n3164 0.152939
R19848 gnd.n3165 gnd.n2395 0.152939
R19849 gnd.n3207 gnd.n2395 0.152939
R19850 gnd.n3208 gnd.n3207 0.152939
R19851 gnd.n3209 gnd.n3208 0.152939
R19852 gnd.n3210 gnd.n3209 0.152939
R19853 gnd.n3210 gnd.n2367 0.152939
R19854 gnd.n3247 gnd.n2367 0.152939
R19855 gnd.n3248 gnd.n3247 0.152939
R19856 gnd.n3249 gnd.n3248 0.152939
R19857 gnd.n3250 gnd.n3249 0.152939
R19858 gnd.n3250 gnd.n2340 0.152939
R19859 gnd.n3296 gnd.n2340 0.152939
R19860 gnd.n3297 gnd.n3296 0.152939
R19861 gnd.n3298 gnd.n3297 0.152939
R19862 gnd.n3299 gnd.n3298 0.152939
R19863 gnd.n3299 gnd.n2313 0.152939
R19864 gnd.n3590 gnd.n2313 0.152939
R19865 gnd.n3591 gnd.n3590 0.152939
R19866 gnd.n3592 gnd.n3591 0.152939
R19867 gnd.n3593 gnd.n3592 0.152939
R19868 gnd.n3594 gnd.n3593 0.152939
R19869 gnd.n2936 gnd.n2666 0.152939
R19870 gnd.n2687 gnd.n2666 0.152939
R19871 gnd.n2688 gnd.n2687 0.152939
R19872 gnd.n2694 gnd.n2688 0.152939
R19873 gnd.n2695 gnd.n2694 0.152939
R19874 gnd.n2696 gnd.n2695 0.152939
R19875 gnd.n2696 gnd.n2685 0.152939
R19876 gnd.n2704 gnd.n2685 0.152939
R19877 gnd.n2705 gnd.n2704 0.152939
R19878 gnd.n2706 gnd.n2705 0.152939
R19879 gnd.n2706 gnd.n2683 0.152939
R19880 gnd.n2714 gnd.n2683 0.152939
R19881 gnd.n2715 gnd.n2714 0.152939
R19882 gnd.n2716 gnd.n2715 0.152939
R19883 gnd.n2716 gnd.n2681 0.152939
R19884 gnd.n2724 gnd.n2681 0.152939
R19885 gnd.n3663 gnd.n2269 0.152939
R19886 gnd.n2271 gnd.n2269 0.152939
R19887 gnd.n2272 gnd.n2271 0.152939
R19888 gnd.n2273 gnd.n2272 0.152939
R19889 gnd.n2274 gnd.n2273 0.152939
R19890 gnd.n2275 gnd.n2274 0.152939
R19891 gnd.n2276 gnd.n2275 0.152939
R19892 gnd.n2277 gnd.n2276 0.152939
R19893 gnd.n2278 gnd.n2277 0.152939
R19894 gnd.n2279 gnd.n2278 0.152939
R19895 gnd.n2280 gnd.n2279 0.152939
R19896 gnd.n2281 gnd.n2280 0.152939
R19897 gnd.n2282 gnd.n2281 0.152939
R19898 gnd.n2283 gnd.n2282 0.152939
R19899 gnd.n2284 gnd.n2283 0.152939
R19900 gnd.n2285 gnd.n2284 0.152939
R19901 gnd.n2286 gnd.n2285 0.152939
R19902 gnd.n2287 gnd.n2286 0.152939
R19903 gnd.n2288 gnd.n2287 0.152939
R19904 gnd.n2289 gnd.n2288 0.152939
R19905 gnd.n2290 gnd.n2289 0.152939
R19906 gnd.n2291 gnd.n2290 0.152939
R19907 gnd.n2295 gnd.n2291 0.152939
R19908 gnd.n2296 gnd.n2295 0.152939
R19909 gnd.n2297 gnd.n2296 0.152939
R19910 gnd.n2298 gnd.n2297 0.152939
R19911 gnd.n3099 gnd.n3098 0.152939
R19912 gnd.n3100 gnd.n3099 0.152939
R19913 gnd.n3101 gnd.n3100 0.152939
R19914 gnd.n3102 gnd.n3101 0.152939
R19915 gnd.n3103 gnd.n3102 0.152939
R19916 gnd.n3104 gnd.n3103 0.152939
R19917 gnd.n3104 gnd.n2403 0.152939
R19918 gnd.n3183 gnd.n2403 0.152939
R19919 gnd.n3184 gnd.n3183 0.152939
R19920 gnd.n3185 gnd.n3184 0.152939
R19921 gnd.n3186 gnd.n3185 0.152939
R19922 gnd.n3187 gnd.n3186 0.152939
R19923 gnd.n3188 gnd.n3187 0.152939
R19924 gnd.n3189 gnd.n3188 0.152939
R19925 gnd.n3190 gnd.n3189 0.152939
R19926 gnd.n3191 gnd.n3190 0.152939
R19927 gnd.n3191 gnd.n2347 0.152939
R19928 gnd.n3268 gnd.n2347 0.152939
R19929 gnd.n3269 gnd.n3268 0.152939
R19930 gnd.n3270 gnd.n3269 0.152939
R19931 gnd.n3271 gnd.n3270 0.152939
R19932 gnd.n3272 gnd.n3271 0.152939
R19933 gnd.n3273 gnd.n3272 0.152939
R19934 gnd.n3274 gnd.n3273 0.152939
R19935 gnd.n3275 gnd.n3274 0.152939
R19936 gnd.n3276 gnd.n3275 0.152939
R19937 gnd.n3278 gnd.n3276 0.152939
R19938 gnd.n3278 gnd.n3277 0.152939
R19939 gnd.n2854 gnd.n2853 0.152939
R19940 gnd.n2854 gnd.n2744 0.152939
R19941 gnd.n2869 gnd.n2744 0.152939
R19942 gnd.n2870 gnd.n2869 0.152939
R19943 gnd.n2871 gnd.n2870 0.152939
R19944 gnd.n2871 gnd.n2732 0.152939
R19945 gnd.n2885 gnd.n2732 0.152939
R19946 gnd.n2886 gnd.n2885 0.152939
R19947 gnd.n2887 gnd.n2886 0.152939
R19948 gnd.n2888 gnd.n2887 0.152939
R19949 gnd.n2889 gnd.n2888 0.152939
R19950 gnd.n2890 gnd.n2889 0.152939
R19951 gnd.n2891 gnd.n2890 0.152939
R19952 gnd.n2892 gnd.n2891 0.152939
R19953 gnd.n2893 gnd.n2892 0.152939
R19954 gnd.n2894 gnd.n2893 0.152939
R19955 gnd.n2895 gnd.n2894 0.152939
R19956 gnd.n2896 gnd.n2895 0.152939
R19957 gnd.n2897 gnd.n2896 0.152939
R19958 gnd.n2898 gnd.n2897 0.152939
R19959 gnd.n2899 gnd.n2898 0.152939
R19960 gnd.n2899 gnd.n2598 0.152939
R19961 gnd.n3016 gnd.n2598 0.152939
R19962 gnd.n3017 gnd.n3016 0.152939
R19963 gnd.n3018 gnd.n3017 0.152939
R19964 gnd.n3019 gnd.n3018 0.152939
R19965 gnd.n3019 gnd.n2520 0.152939
R19966 gnd.n3096 gnd.n2520 0.152939
R19967 gnd.n2772 gnd.n2771 0.152939
R19968 gnd.n2773 gnd.n2772 0.152939
R19969 gnd.n2774 gnd.n2773 0.152939
R19970 gnd.n2775 gnd.n2774 0.152939
R19971 gnd.n2776 gnd.n2775 0.152939
R19972 gnd.n2777 gnd.n2776 0.152939
R19973 gnd.n2778 gnd.n2777 0.152939
R19974 gnd.n2779 gnd.n2778 0.152939
R19975 gnd.n2780 gnd.n2779 0.152939
R19976 gnd.n2781 gnd.n2780 0.152939
R19977 gnd.n2782 gnd.n2781 0.152939
R19978 gnd.n2783 gnd.n2782 0.152939
R19979 gnd.n2784 gnd.n2783 0.152939
R19980 gnd.n2785 gnd.n2784 0.152939
R19981 gnd.n2786 gnd.n2785 0.152939
R19982 gnd.n2787 gnd.n2786 0.152939
R19983 gnd.n2788 gnd.n2787 0.152939
R19984 gnd.n2789 gnd.n2788 0.152939
R19985 gnd.n2790 gnd.n2789 0.152939
R19986 gnd.n2791 gnd.n2790 0.152939
R19987 gnd.n2792 gnd.n2791 0.152939
R19988 gnd.n2793 gnd.n2792 0.152939
R19989 gnd.n2797 gnd.n2793 0.152939
R19990 gnd.n2798 gnd.n2797 0.152939
R19991 gnd.n2798 gnd.n2755 0.152939
R19992 gnd.n2852 gnd.n2755 0.152939
R19993 gnd.n3752 gnd.n2225 0.152939
R19994 gnd.n3753 gnd.n3752 0.152939
R19995 gnd.n3754 gnd.n3753 0.152939
R19996 gnd.n3754 gnd.n3744 0.152939
R19997 gnd.n3762 gnd.n3744 0.152939
R19998 gnd.n3763 gnd.n3762 0.152939
R19999 gnd.n3764 gnd.n3763 0.152939
R20000 gnd.n3764 gnd.n3740 0.152939
R20001 gnd.n3772 gnd.n3740 0.152939
R20002 gnd.n3773 gnd.n3772 0.152939
R20003 gnd.n3774 gnd.n3773 0.152939
R20004 gnd.n3774 gnd.n3736 0.152939
R20005 gnd.n3782 gnd.n3736 0.152939
R20006 gnd.n3783 gnd.n3782 0.152939
R20007 gnd.n3784 gnd.n3783 0.152939
R20008 gnd.n3784 gnd.n3729 0.152939
R20009 gnd.n3792 gnd.n3729 0.152939
R20010 gnd.n3793 gnd.n3792 0.152939
R20011 gnd.n3794 gnd.n3793 0.152939
R20012 gnd.n3794 gnd.n3725 0.152939
R20013 gnd.n3802 gnd.n3725 0.152939
R20014 gnd.n3803 gnd.n3802 0.152939
R20015 gnd.n3804 gnd.n3803 0.152939
R20016 gnd.n3804 gnd.n3721 0.152939
R20017 gnd.n3812 gnd.n3721 0.152939
R20018 gnd.n3813 gnd.n3812 0.152939
R20019 gnd.n3814 gnd.n3813 0.152939
R20020 gnd.n3814 gnd.n3717 0.152939
R20021 gnd.n3822 gnd.n3717 0.152939
R20022 gnd.n3823 gnd.n3822 0.152939
R20023 gnd.n3824 gnd.n3823 0.152939
R20024 gnd.n3824 gnd.n3713 0.152939
R20025 gnd.n3832 gnd.n3713 0.152939
R20026 gnd.n3833 gnd.n3832 0.152939
R20027 gnd.n3835 gnd.n3833 0.152939
R20028 gnd.n3835 gnd.n3834 0.152939
R20029 gnd.n3834 gnd.n3706 0.152939
R20030 gnd.n3844 gnd.n3706 0.152939
R20031 gnd.n4196 gnd.n4195 0.152939
R20032 gnd.n4197 gnd.n4196 0.152939
R20033 gnd.n4197 gnd.n2210 0.152939
R20034 gnd.n4211 gnd.n2210 0.152939
R20035 gnd.n4212 gnd.n4211 0.152939
R20036 gnd.n4213 gnd.n4212 0.152939
R20037 gnd.n4213 gnd.n2193 0.152939
R20038 gnd.n4227 gnd.n2193 0.152939
R20039 gnd.n4228 gnd.n4227 0.152939
R20040 gnd.n4229 gnd.n4228 0.152939
R20041 gnd.n4229 gnd.n2178 0.152939
R20042 gnd.n4243 gnd.n2178 0.152939
R20043 gnd.n4244 gnd.n4243 0.152939
R20044 gnd.n4245 gnd.n4244 0.152939
R20045 gnd.n4245 gnd.n2161 0.152939
R20046 gnd.n4259 gnd.n2161 0.152939
R20047 gnd.n4260 gnd.n4259 0.152939
R20048 gnd.n4261 gnd.n4260 0.152939
R20049 gnd.n4261 gnd.n2146 0.152939
R20050 gnd.n4275 gnd.n2146 0.152939
R20051 gnd.n4276 gnd.n4275 0.152939
R20052 gnd.n4277 gnd.n4276 0.152939
R20053 gnd.n4277 gnd.n2129 0.152939
R20054 gnd.n4291 gnd.n2129 0.152939
R20055 gnd.n4292 gnd.n4291 0.152939
R20056 gnd.n4293 gnd.n4292 0.152939
R20057 gnd.n4293 gnd.n2114 0.152939
R20058 gnd.n4341 gnd.n4340 0.152939
R20059 gnd.n4341 gnd.n2064 0.152939
R20060 gnd.n4355 gnd.n2064 0.152939
R20061 gnd.n4356 gnd.n4355 0.152939
R20062 gnd.n4357 gnd.n4356 0.152939
R20063 gnd.n4357 gnd.n2049 0.152939
R20064 gnd.n4371 gnd.n2049 0.152939
R20065 gnd.n4372 gnd.n4371 0.152939
R20066 gnd.n4373 gnd.n4372 0.152939
R20067 gnd.n4373 gnd.n2032 0.152939
R20068 gnd.n4387 gnd.n2032 0.152939
R20069 gnd.n4388 gnd.n4387 0.152939
R20070 gnd.n4389 gnd.n4388 0.152939
R20071 gnd.n4389 gnd.n2016 0.152939
R20072 gnd.n4416 gnd.n2016 0.152939
R20073 gnd.n4417 gnd.n4416 0.152939
R20074 gnd.n4418 gnd.n4417 0.152939
R20075 gnd.n4420 gnd.n4418 0.152939
R20076 gnd.n4420 gnd.n4419 0.152939
R20077 gnd.n4419 gnd.n1063 0.152939
R20078 gnd.n1064 gnd.n1063 0.152939
R20079 gnd.n1065 gnd.n1064 0.152939
R20080 gnd.n1085 gnd.n1065 0.152939
R20081 gnd.n1086 gnd.n1085 0.152939
R20082 gnd.n1087 gnd.n1086 0.152939
R20083 gnd.n1088 gnd.n1087 0.152939
R20084 gnd.n1914 gnd.n1088 0.152939
R20085 gnd.n1916 gnd.n1915 0.152939
R20086 gnd.n1917 gnd.n1916 0.152939
R20087 gnd.n1918 gnd.n1917 0.152939
R20088 gnd.n1919 gnd.n1918 0.152939
R20089 gnd.n1920 gnd.n1919 0.152939
R20090 gnd.n1921 gnd.n1920 0.152939
R20091 gnd.n1922 gnd.n1921 0.152939
R20092 gnd.n1923 gnd.n1922 0.152939
R20093 gnd.n1924 gnd.n1923 0.152939
R20094 gnd.n1925 gnd.n1924 0.152939
R20095 gnd.n1926 gnd.n1925 0.152939
R20096 gnd.n1927 gnd.n1926 0.152939
R20097 gnd.n1928 gnd.n1927 0.152939
R20098 gnd.n1929 gnd.n1928 0.152939
R20099 gnd.n1929 gnd.n1900 0.152939
R20100 gnd.n4826 gnd.n4825 0.152939
R20101 gnd.n4825 gnd.n1901 0.152939
R20102 gnd.n1963 gnd.n1901 0.152939
R20103 gnd.n1964 gnd.n1963 0.152939
R20104 gnd.n1965 gnd.n1964 0.152939
R20105 gnd.n1966 gnd.n1965 0.152939
R20106 gnd.n1970 gnd.n1966 0.152939
R20107 gnd.n1971 gnd.n1970 0.152939
R20108 gnd.n1972 gnd.n1971 0.152939
R20109 gnd.n1973 gnd.n1972 0.152939
R20110 gnd.n1977 gnd.n1973 0.152939
R20111 gnd.n1978 gnd.n1977 0.152939
R20112 gnd.n1979 gnd.n1978 0.152939
R20113 gnd.n1980 gnd.n1979 0.152939
R20114 gnd.n1984 gnd.n1980 0.152939
R20115 gnd.n1985 gnd.n1984 0.152939
R20116 gnd.n1986 gnd.n1985 0.152939
R20117 gnd.n1987 gnd.n1986 0.152939
R20118 gnd.n1993 gnd.n1987 0.152939
R20119 gnd.n4788 gnd.n1993 0.152939
R20120 gnd.n3982 gnd.n3845 0.152939
R20121 gnd.n3982 gnd.n3981 0.152939
R20122 gnd.n3981 gnd.n3980 0.152939
R20123 gnd.n3980 gnd.n3846 0.152939
R20124 gnd.n3847 gnd.n3846 0.152939
R20125 gnd.n3848 gnd.n3847 0.152939
R20126 gnd.n3849 gnd.n3848 0.152939
R20127 gnd.n3850 gnd.n3849 0.152939
R20128 gnd.n3851 gnd.n3850 0.152939
R20129 gnd.n3852 gnd.n3851 0.152939
R20130 gnd.n3853 gnd.n3852 0.152939
R20131 gnd.n3854 gnd.n3853 0.152939
R20132 gnd.n3855 gnd.n3854 0.152939
R20133 gnd.n3856 gnd.n3855 0.152939
R20134 gnd.n3857 gnd.n3856 0.152939
R20135 gnd.n3858 gnd.n3857 0.152939
R20136 gnd.n3859 gnd.n3858 0.152939
R20137 gnd.n3860 gnd.n3859 0.152939
R20138 gnd.n3861 gnd.n3860 0.152939
R20139 gnd.n3862 gnd.n3861 0.152939
R20140 gnd.n3863 gnd.n3862 0.152939
R20141 gnd.n3864 gnd.n3863 0.152939
R20142 gnd.n3865 gnd.n3864 0.152939
R20143 gnd.n3866 gnd.n3865 0.152939
R20144 gnd.n3867 gnd.n3866 0.152939
R20145 gnd.n3868 gnd.n3867 0.152939
R20146 gnd.n3869 gnd.n3868 0.152939
R20147 gnd.n3870 gnd.n3869 0.152939
R20148 gnd.n3871 gnd.n3870 0.152939
R20149 gnd.n3872 gnd.n3871 0.152939
R20150 gnd.n3873 gnd.n3872 0.152939
R20151 gnd.n3873 gnd.n2105 0.152939
R20152 gnd.n3874 gnd.n2105 0.152939
R20153 gnd.n3875 gnd.n3874 0.152939
R20154 gnd.n3876 gnd.n3875 0.152939
R20155 gnd.n3877 gnd.n3876 0.152939
R20156 gnd.n3878 gnd.n3877 0.152939
R20157 gnd.n3879 gnd.n3878 0.152939
R20158 gnd.n3880 gnd.n3879 0.152939
R20159 gnd.n3881 gnd.n3880 0.152939
R20160 gnd.n3882 gnd.n3881 0.152939
R20161 gnd.n3883 gnd.n3882 0.152939
R20162 gnd.n3884 gnd.n3883 0.152939
R20163 gnd.n3885 gnd.n3884 0.152939
R20164 gnd.n3886 gnd.n3885 0.152939
R20165 gnd.n3887 gnd.n3886 0.152939
R20166 gnd.n3888 gnd.n3887 0.152939
R20167 gnd.n3889 gnd.n3888 0.152939
R20168 gnd.n3890 gnd.n3889 0.152939
R20169 gnd.n3891 gnd.n3890 0.152939
R20170 gnd.n3892 gnd.n3891 0.152939
R20171 gnd.n3893 gnd.n3892 0.152939
R20172 gnd.n3894 gnd.n3893 0.152939
R20173 gnd.n3895 gnd.n3894 0.152939
R20174 gnd.n3896 gnd.n3895 0.152939
R20175 gnd.n3897 gnd.n3896 0.152939
R20176 gnd.n3897 gnd.n2002 0.152939
R20177 gnd.n4437 gnd.n2002 0.152939
R20178 gnd.n4438 gnd.n4437 0.152939
R20179 gnd.n4440 gnd.n4438 0.152939
R20180 gnd.n4440 gnd.n4439 0.152939
R20181 gnd.n4439 gnd.n1996 0.152939
R20182 gnd.n1996 gnd.n1994 0.152939
R20183 gnd.n4787 gnd.n1994 0.152939
R20184 gnd.n4147 gnd.n4013 0.152939
R20185 gnd.n4014 gnd.n4013 0.152939
R20186 gnd.n4015 gnd.n4014 0.152939
R20187 gnd.n4016 gnd.n4015 0.152939
R20188 gnd.n4017 gnd.n4016 0.152939
R20189 gnd.n4018 gnd.n4017 0.152939
R20190 gnd.n4019 gnd.n4018 0.152939
R20191 gnd.n4020 gnd.n4019 0.152939
R20192 gnd.n4021 gnd.n4020 0.152939
R20193 gnd.n4022 gnd.n4021 0.152939
R20194 gnd.n4023 gnd.n4022 0.152939
R20195 gnd.n4024 gnd.n4023 0.152939
R20196 gnd.n4025 gnd.n4024 0.152939
R20197 gnd.n4026 gnd.n4025 0.152939
R20198 gnd.n4027 gnd.n4026 0.152939
R20199 gnd.n4028 gnd.n4027 0.152939
R20200 gnd.n4029 gnd.n4028 0.152939
R20201 gnd.n4030 gnd.n4029 0.152939
R20202 gnd.n4031 gnd.n4030 0.152939
R20203 gnd.n4032 gnd.n4031 0.152939
R20204 gnd.n4033 gnd.n4032 0.152939
R20205 gnd.n4034 gnd.n4033 0.152939
R20206 gnd.n4035 gnd.n4034 0.152939
R20207 gnd.n4036 gnd.n4035 0.152939
R20208 gnd.n4037 gnd.n4036 0.152939
R20209 gnd.n4038 gnd.n4037 0.152939
R20210 gnd.n4039 gnd.n4038 0.152939
R20211 gnd.n4040 gnd.n4039 0.152939
R20212 gnd.n4041 gnd.n4040 0.152939
R20213 gnd.n4042 gnd.n4041 0.152939
R20214 gnd.n4043 gnd.n4042 0.152939
R20215 gnd.n4188 gnd.n3987 0.152939
R20216 gnd.n3990 gnd.n3987 0.152939
R20217 gnd.n3991 gnd.n3990 0.152939
R20218 gnd.n3992 gnd.n3991 0.152939
R20219 gnd.n3993 gnd.n3992 0.152939
R20220 gnd.n3996 gnd.n3993 0.152939
R20221 gnd.n3997 gnd.n3996 0.152939
R20222 gnd.n3998 gnd.n3997 0.152939
R20223 gnd.n3999 gnd.n3998 0.152939
R20224 gnd.n4002 gnd.n3999 0.152939
R20225 gnd.n4003 gnd.n4002 0.152939
R20226 gnd.n4004 gnd.n4003 0.152939
R20227 gnd.n4005 gnd.n4004 0.152939
R20228 gnd.n4008 gnd.n4005 0.152939
R20229 gnd.n4009 gnd.n4008 0.152939
R20230 gnd.n4154 gnd.n4009 0.152939
R20231 gnd.n4154 gnd.n4153 0.152939
R20232 gnd.n4153 gnd.n4152 0.152939
R20233 gnd.n4189 gnd.n2218 0.152939
R20234 gnd.n4203 gnd.n2218 0.152939
R20235 gnd.n4204 gnd.n4203 0.152939
R20236 gnd.n4205 gnd.n4204 0.152939
R20237 gnd.n4205 gnd.n2202 0.152939
R20238 gnd.n4219 gnd.n2202 0.152939
R20239 gnd.n4220 gnd.n4219 0.152939
R20240 gnd.n4221 gnd.n4220 0.152939
R20241 gnd.n4221 gnd.n2186 0.152939
R20242 gnd.n4235 gnd.n2186 0.152939
R20243 gnd.n4236 gnd.n4235 0.152939
R20244 gnd.n4237 gnd.n4236 0.152939
R20245 gnd.n4237 gnd.n2170 0.152939
R20246 gnd.n4251 gnd.n2170 0.152939
R20247 gnd.n4252 gnd.n4251 0.152939
R20248 gnd.n4253 gnd.n4252 0.152939
R20249 gnd.n4253 gnd.n2154 0.152939
R20250 gnd.n4267 gnd.n2154 0.152939
R20251 gnd.n4268 gnd.n4267 0.152939
R20252 gnd.n4269 gnd.n4268 0.152939
R20253 gnd.n4269 gnd.n2138 0.152939
R20254 gnd.n4283 gnd.n2138 0.152939
R20255 gnd.n4284 gnd.n4283 0.152939
R20256 gnd.n4285 gnd.n4284 0.152939
R20257 gnd.n4285 gnd.n2122 0.152939
R20258 gnd.n4299 gnd.n2122 0.152939
R20259 gnd.n4300 gnd.n4299 0.152939
R20260 gnd.n4301 gnd.n4300 0.152939
R20261 gnd.n4301 gnd.n2106 0.152939
R20262 gnd.n4315 gnd.n2106 0.152939
R20263 gnd.n4316 gnd.n4315 0.152939
R20264 gnd.n4317 gnd.n4316 0.152939
R20265 gnd.n4317 gnd.n2088 0.152939
R20266 gnd.n4331 gnd.n2088 0.152939
R20267 gnd.n4332 gnd.n4331 0.152939
R20268 gnd.n4333 gnd.n4332 0.152939
R20269 gnd.n4333 gnd.n2073 0.152939
R20270 gnd.n4347 gnd.n2073 0.152939
R20271 gnd.n4348 gnd.n4347 0.152939
R20272 gnd.n4349 gnd.n4348 0.152939
R20273 gnd.n4349 gnd.n2056 0.152939
R20274 gnd.n4363 gnd.n2056 0.152939
R20275 gnd.n4364 gnd.n4363 0.152939
R20276 gnd.n4365 gnd.n4364 0.152939
R20277 gnd.n4365 gnd.n2041 0.152939
R20278 gnd.n4379 gnd.n2041 0.152939
R20279 gnd.n4380 gnd.n4379 0.152939
R20280 gnd.n4381 gnd.n4380 0.152939
R20281 gnd.n4381 gnd.n2024 0.152939
R20282 gnd.n4395 gnd.n2024 0.152939
R20283 gnd.n4396 gnd.n4395 0.152939
R20284 gnd.n4397 gnd.n4396 0.152939
R20285 gnd.n4398 gnd.n4397 0.152939
R20286 gnd.n4399 gnd.n4398 0.152939
R20287 gnd.n4400 gnd.n4399 0.152939
R20288 gnd.n4401 gnd.n4400 0.152939
R20289 gnd.n4403 gnd.n4401 0.152939
R20290 gnd.n4403 gnd.n4402 0.152939
R20291 gnd.n4402 gnd.n1075 0.152939
R20292 gnd.n1076 gnd.n1075 0.152939
R20293 gnd.n1077 gnd.n1076 0.152939
R20294 gnd.n1096 gnd.n1077 0.152939
R20295 gnd.n1097 gnd.n1096 0.152939
R20296 gnd.n6056 gnd.n1097 0.152939
R20297 gnd.n1283 gnd.n1282 0.152939
R20298 gnd.n1283 gnd.n1273 0.152939
R20299 gnd.n1289 gnd.n1273 0.152939
R20300 gnd.n1290 gnd.n1289 0.152939
R20301 gnd.n1291 gnd.n1290 0.152939
R20302 gnd.n1291 gnd.n1267 0.152939
R20303 gnd.n1298 gnd.n1267 0.152939
R20304 gnd.n1299 gnd.n1298 0.152939
R20305 gnd.n5887 gnd.n1299 0.152939
R20306 gnd.n4699 gnd.n4581 0.152939
R20307 gnd.n4695 gnd.n4581 0.152939
R20308 gnd.n4695 gnd.n4694 0.152939
R20309 gnd.n4694 gnd.n4693 0.152939
R20310 gnd.n4693 gnd.n4587 0.152939
R20311 gnd.n4689 gnd.n4587 0.152939
R20312 gnd.n4689 gnd.n4688 0.152939
R20313 gnd.n4688 gnd.n4687 0.152939
R20314 gnd.n4687 gnd.n4592 0.152939
R20315 gnd.n4683 gnd.n4592 0.152939
R20316 gnd.n4683 gnd.n4682 0.152939
R20317 gnd.n4682 gnd.n4681 0.152939
R20318 gnd.n4681 gnd.n4597 0.152939
R20319 gnd.n4677 gnd.n4597 0.152939
R20320 gnd.n4677 gnd.n4676 0.152939
R20321 gnd.n4676 gnd.n4675 0.152939
R20322 gnd.n4675 gnd.n1741 0.152939
R20323 gnd.n4977 gnd.n1741 0.152939
R20324 gnd.n4978 gnd.n4977 0.152939
R20325 gnd.n4980 gnd.n4978 0.152939
R20326 gnd.n4980 gnd.n4979 0.152939
R20327 gnd.n4979 gnd.n1711 0.152939
R20328 gnd.n5016 gnd.n1711 0.152939
R20329 gnd.n5017 gnd.n5016 0.152939
R20330 gnd.n5055 gnd.n5017 0.152939
R20331 gnd.n5055 gnd.n5054 0.152939
R20332 gnd.n5054 gnd.n5053 0.152939
R20333 gnd.n5053 gnd.n5018 0.152939
R20334 gnd.n5049 gnd.n5018 0.152939
R20335 gnd.n5049 gnd.n5048 0.152939
R20336 gnd.n5048 gnd.n5047 0.152939
R20337 gnd.n5047 gnd.n5023 0.152939
R20338 gnd.n5043 gnd.n5023 0.152939
R20339 gnd.n5043 gnd.n5042 0.152939
R20340 gnd.n5042 gnd.n5041 0.152939
R20341 gnd.n5041 gnd.n5029 0.152939
R20342 gnd.n5037 gnd.n5029 0.152939
R20343 gnd.n5037 gnd.n5036 0.152939
R20344 gnd.n5036 gnd.n1626 0.152939
R20345 gnd.n5194 gnd.n1626 0.152939
R20346 gnd.n5195 gnd.n5194 0.152939
R20347 gnd.n5231 gnd.n5195 0.152939
R20348 gnd.n5231 gnd.n5230 0.152939
R20349 gnd.n5230 gnd.n5229 0.152939
R20350 gnd.n5229 gnd.n5196 0.152939
R20351 gnd.n5225 gnd.n5196 0.152939
R20352 gnd.n5225 gnd.n5224 0.152939
R20353 gnd.n5224 gnd.n5223 0.152939
R20354 gnd.n5223 gnd.n5201 0.152939
R20355 gnd.n5219 gnd.n5201 0.152939
R20356 gnd.n5219 gnd.n5218 0.152939
R20357 gnd.n5218 gnd.n5217 0.152939
R20358 gnd.n5217 gnd.n5205 0.152939
R20359 gnd.n5213 gnd.n5205 0.152939
R20360 gnd.n5213 gnd.n5212 0.152939
R20361 gnd.n5212 gnd.n1539 0.152939
R20362 gnd.n5371 gnd.n1539 0.152939
R20363 gnd.n5372 gnd.n5371 0.152939
R20364 gnd.n5393 gnd.n5372 0.152939
R20365 gnd.n5393 gnd.n5392 0.152939
R20366 gnd.n5392 gnd.n5391 0.152939
R20367 gnd.n5391 gnd.n5373 0.152939
R20368 gnd.n5387 gnd.n5373 0.152939
R20369 gnd.n5387 gnd.n5386 0.152939
R20370 gnd.n5386 gnd.n5385 0.152939
R20371 gnd.n5385 gnd.n5378 0.152939
R20372 gnd.n5381 gnd.n5378 0.152939
R20373 gnd.n5381 gnd.n1474 0.152939
R20374 gnd.n5504 gnd.n1474 0.152939
R20375 gnd.n5505 gnd.n5504 0.152939
R20376 gnd.n5507 gnd.n5505 0.152939
R20377 gnd.n5507 gnd.n5506 0.152939
R20378 gnd.n5506 gnd.n1447 0.152939
R20379 gnd.n5543 gnd.n1447 0.152939
R20380 gnd.n5544 gnd.n5543 0.152939
R20381 gnd.n5575 gnd.n5544 0.152939
R20382 gnd.n5575 gnd.n5574 0.152939
R20383 gnd.n5574 gnd.n5573 0.152939
R20384 gnd.n5573 gnd.n5545 0.152939
R20385 gnd.n5569 gnd.n5545 0.152939
R20386 gnd.n5569 gnd.n5568 0.152939
R20387 gnd.n5568 gnd.n5567 0.152939
R20388 gnd.n5567 gnd.n5551 0.152939
R20389 gnd.n5563 gnd.n5551 0.152939
R20390 gnd.n5563 gnd.n5562 0.152939
R20391 gnd.n5562 gnd.n5561 0.152939
R20392 gnd.n5561 gnd.n1336 0.152939
R20393 gnd.n5822 gnd.n1336 0.152939
R20394 gnd.n5823 gnd.n5822 0.152939
R20395 gnd.n5824 gnd.n5823 0.152939
R20396 gnd.n5824 gnd.n1324 0.152939
R20397 gnd.n5842 gnd.n1324 0.152939
R20398 gnd.n5843 gnd.n5842 0.152939
R20399 gnd.n5844 gnd.n5843 0.152939
R20400 gnd.n5844 gnd.n1311 0.152939
R20401 gnd.n5862 gnd.n1311 0.152939
R20402 gnd.n5863 gnd.n5862 0.152939
R20403 gnd.n5865 gnd.n5863 0.152939
R20404 gnd.n5865 gnd.n5864 0.152939
R20405 gnd.n5864 gnd.n1300 0.152939
R20406 gnd.n5886 gnd.n1300 0.152939
R20407 gnd.n4713 gnd.n4712 0.152939
R20408 gnd.n4712 gnd.n4711 0.152939
R20409 gnd.n4711 gnd.n4566 0.152939
R20410 gnd.n4707 gnd.n4566 0.152939
R20411 gnd.n4707 gnd.n4706 0.152939
R20412 gnd.n4706 gnd.n4705 0.152939
R20413 gnd.n4705 gnd.n4572 0.152939
R20414 gnd.n4701 gnd.n4572 0.152939
R20415 gnd.n4701 gnd.n4700 0.152939
R20416 gnd.n4096 gnd.n4095 0.152939
R20417 gnd.n4095 gnd.n4046 0.152939
R20418 gnd.n4091 gnd.n4046 0.152939
R20419 gnd.n4091 gnd.n4090 0.152939
R20420 gnd.n4090 gnd.n4089 0.152939
R20421 gnd.n4089 gnd.n4050 0.152939
R20422 gnd.n4085 gnd.n4050 0.152939
R20423 gnd.n4085 gnd.n4084 0.152939
R20424 gnd.n4084 gnd.n4083 0.152939
R20425 gnd.n4083 gnd.n4054 0.152939
R20426 gnd.n4079 gnd.n4054 0.152939
R20427 gnd.n4079 gnd.n4078 0.152939
R20428 gnd.n4078 gnd.n4077 0.152939
R20429 gnd.n4077 gnd.n4058 0.152939
R20430 gnd.n4073 gnd.n4058 0.152939
R20431 gnd.n4073 gnd.n4072 0.152939
R20432 gnd.n4072 gnd.n4071 0.152939
R20433 gnd.n4071 gnd.n4062 0.152939
R20434 gnd.n4067 gnd.n4062 0.152939
R20435 gnd.n4067 gnd.n4066 0.152939
R20436 gnd.n4066 gnd.n4065 0.152939
R20437 gnd.n4065 gnd.n2006 0.152939
R20438 gnd.n4429 gnd.n2006 0.152939
R20439 gnd.n4430 gnd.n4429 0.152939
R20440 gnd.n4431 gnd.n4430 0.152939
R20441 gnd.n4431 gnd.n1999 0.152939
R20442 gnd.n4446 gnd.n1999 0.152939
R20443 gnd.n4447 gnd.n4446 0.152939
R20444 gnd.n4779 gnd.n4447 0.152939
R20445 gnd.n4779 gnd.n4778 0.152939
R20446 gnd.n4778 gnd.n4777 0.152939
R20447 gnd.n6053 gnd.n1100 0.152939
R20448 gnd.n6049 gnd.n1100 0.152939
R20449 gnd.n6049 gnd.n6048 0.152939
R20450 gnd.n6048 gnd.n6047 0.152939
R20451 gnd.n6047 gnd.n1105 0.152939
R20452 gnd.n6043 gnd.n1105 0.152939
R20453 gnd.n6043 gnd.n6042 0.152939
R20454 gnd.n6042 gnd.n6041 0.152939
R20455 gnd.n6041 gnd.n1110 0.152939
R20456 gnd.n6037 gnd.n1110 0.152939
R20457 gnd.n6037 gnd.n6036 0.152939
R20458 gnd.n6036 gnd.n6035 0.152939
R20459 gnd.n6035 gnd.n1115 0.152939
R20460 gnd.n6031 gnd.n1115 0.152939
R20461 gnd.n6031 gnd.n6030 0.152939
R20462 gnd.n6030 gnd.n6029 0.152939
R20463 gnd.n6029 gnd.n1120 0.152939
R20464 gnd.n6025 gnd.n1120 0.152939
R20465 gnd.n6025 gnd.n6024 0.152939
R20466 gnd.n6024 gnd.n6023 0.152939
R20467 gnd.n6023 gnd.n1125 0.152939
R20468 gnd.n6019 gnd.n1125 0.152939
R20469 gnd.n6019 gnd.n6018 0.152939
R20470 gnd.n6018 gnd.n6017 0.152939
R20471 gnd.n6017 gnd.n1130 0.152939
R20472 gnd.n6013 gnd.n1130 0.152939
R20473 gnd.n6013 gnd.n6012 0.152939
R20474 gnd.n6012 gnd.n6011 0.152939
R20475 gnd.n6011 gnd.n1135 0.152939
R20476 gnd.n6007 gnd.n1135 0.152939
R20477 gnd.n6007 gnd.n6006 0.152939
R20478 gnd.n6006 gnd.n6005 0.152939
R20479 gnd.n6005 gnd.n1140 0.152939
R20480 gnd.n6001 gnd.n1140 0.152939
R20481 gnd.n6001 gnd.n6000 0.152939
R20482 gnd.n6000 gnd.n5999 0.152939
R20483 gnd.n5999 gnd.n1145 0.152939
R20484 gnd.n5995 gnd.n1145 0.152939
R20485 gnd.n5995 gnd.n5994 0.152939
R20486 gnd.n5994 gnd.n5993 0.152939
R20487 gnd.n5993 gnd.n1150 0.152939
R20488 gnd.n5989 gnd.n1150 0.152939
R20489 gnd.n5989 gnd.n5988 0.152939
R20490 gnd.n5988 gnd.n5987 0.152939
R20491 gnd.n5987 gnd.n1155 0.152939
R20492 gnd.n5983 gnd.n1155 0.152939
R20493 gnd.n5983 gnd.n5982 0.152939
R20494 gnd.n5982 gnd.n5981 0.152939
R20495 gnd.n5981 gnd.n1160 0.152939
R20496 gnd.n5977 gnd.n1160 0.152939
R20497 gnd.n5977 gnd.n5976 0.152939
R20498 gnd.n5976 gnd.n5975 0.152939
R20499 gnd.n5975 gnd.n1165 0.152939
R20500 gnd.n5971 gnd.n1165 0.152939
R20501 gnd.n5971 gnd.n5970 0.152939
R20502 gnd.n5970 gnd.n5969 0.152939
R20503 gnd.n5969 gnd.n1170 0.152939
R20504 gnd.n5965 gnd.n1170 0.152939
R20505 gnd.n5965 gnd.n5964 0.152939
R20506 gnd.n5964 gnd.n5963 0.152939
R20507 gnd.n5963 gnd.n1175 0.152939
R20508 gnd.n5959 gnd.n1175 0.152939
R20509 gnd.n5959 gnd.n5958 0.152939
R20510 gnd.n5958 gnd.n5957 0.152939
R20511 gnd.n5957 gnd.n1180 0.152939
R20512 gnd.n5953 gnd.n1180 0.152939
R20513 gnd.n5953 gnd.n5952 0.152939
R20514 gnd.n5952 gnd.n5951 0.152939
R20515 gnd.n5951 gnd.n1185 0.152939
R20516 gnd.n5947 gnd.n1185 0.152939
R20517 gnd.n5947 gnd.n5946 0.152939
R20518 gnd.n5946 gnd.n5945 0.152939
R20519 gnd.n5945 gnd.n1190 0.152939
R20520 gnd.n5941 gnd.n1190 0.152939
R20521 gnd.n5941 gnd.n5940 0.152939
R20522 gnd.n5940 gnd.n5939 0.152939
R20523 gnd.n5939 gnd.n1195 0.152939
R20524 gnd.n5935 gnd.n1195 0.152939
R20525 gnd.n5935 gnd.n5934 0.152939
R20526 gnd.n5934 gnd.n5933 0.152939
R20527 gnd.n5933 gnd.n1200 0.152939
R20528 gnd.n5929 gnd.n1200 0.152939
R20529 gnd.n5929 gnd.n5928 0.152939
R20530 gnd.n5928 gnd.n5927 0.152939
R20531 gnd.n5927 gnd.n1205 0.152939
R20532 gnd.n5923 gnd.n1205 0.152939
R20533 gnd.n5923 gnd.n5922 0.152939
R20534 gnd.n5922 gnd.n5921 0.152939
R20535 gnd.n5921 gnd.n1210 0.152939
R20536 gnd.n5917 gnd.n1210 0.152939
R20537 gnd.n5917 gnd.n5916 0.152939
R20538 gnd.n5916 gnd.n5915 0.152939
R20539 gnd.n5915 gnd.n1215 0.152939
R20540 gnd.n5911 gnd.n1215 0.152939
R20541 gnd.n5911 gnd.n5910 0.152939
R20542 gnd.n5910 gnd.n5909 0.152939
R20543 gnd.n5909 gnd.n1220 0.152939
R20544 gnd.n5905 gnd.n1220 0.152939
R20545 gnd.n5905 gnd.n5904 0.152939
R20546 gnd.n5904 gnd.n5903 0.152939
R20547 gnd.n5903 gnd.n1225 0.152939
R20548 gnd.n7154 gnd.n440 0.152939
R20549 gnd.n7168 gnd.n440 0.152939
R20550 gnd.n7169 gnd.n7168 0.152939
R20551 gnd.n7170 gnd.n7169 0.152939
R20552 gnd.n7170 gnd.n422 0.152939
R20553 gnd.n7184 gnd.n422 0.152939
R20554 gnd.n7185 gnd.n7184 0.152939
R20555 gnd.n7186 gnd.n7185 0.152939
R20556 gnd.n7186 gnd.n406 0.152939
R20557 gnd.n7200 gnd.n406 0.152939
R20558 gnd.n7201 gnd.n7200 0.152939
R20559 gnd.n7202 gnd.n7201 0.152939
R20560 gnd.n7202 gnd.n390 0.152939
R20561 gnd.n7216 gnd.n390 0.152939
R20562 gnd.n7217 gnd.n7216 0.152939
R20563 gnd.n7218 gnd.n7217 0.152939
R20564 gnd.n7218 gnd.n374 0.152939
R20565 gnd.n7232 gnd.n374 0.152939
R20566 gnd.n7233 gnd.n7232 0.152939
R20567 gnd.n7234 gnd.n7233 0.152939
R20568 gnd.n7234 gnd.n358 0.152939
R20569 gnd.n7248 gnd.n358 0.152939
R20570 gnd.n7249 gnd.n7248 0.152939
R20571 gnd.n7250 gnd.n7249 0.152939
R20572 gnd.n7250 gnd.n342 0.152939
R20573 gnd.n7264 gnd.n342 0.152939
R20574 gnd.n7265 gnd.n7264 0.152939
R20575 gnd.n7266 gnd.n7265 0.152939
R20576 gnd.n7266 gnd.n326 0.152939
R20577 gnd.n7280 gnd.n326 0.152939
R20578 gnd.n7281 gnd.n7280 0.152939
R20579 gnd.n7282 gnd.n7281 0.152939
R20580 gnd.n7282 gnd.n309 0.152939
R20581 gnd.n7296 gnd.n309 0.152939
R20582 gnd.n7297 gnd.n7296 0.152939
R20583 gnd.n7298 gnd.n7297 0.152939
R20584 gnd.n7298 gnd.n295 0.152939
R20585 gnd.n7312 gnd.n295 0.152939
R20586 gnd.n7313 gnd.n7312 0.152939
R20587 gnd.n7314 gnd.n7313 0.152939
R20588 gnd.n7314 gnd.n279 0.152939
R20589 gnd.n7328 gnd.n279 0.152939
R20590 gnd.n7329 gnd.n7328 0.152939
R20591 gnd.n7330 gnd.n7329 0.152939
R20592 gnd.n7330 gnd.n265 0.152939
R20593 gnd.n7344 gnd.n265 0.152939
R20594 gnd.n7345 gnd.n7344 0.152939
R20595 gnd.n7346 gnd.n7345 0.152939
R20596 gnd.n7346 gnd.n249 0.152939
R20597 gnd.n7360 gnd.n249 0.152939
R20598 gnd.n7361 gnd.n7360 0.152939
R20599 gnd.n7362 gnd.n7361 0.152939
R20600 gnd.n7362 gnd.n235 0.152939
R20601 gnd.n7376 gnd.n235 0.152939
R20602 gnd.n7377 gnd.n7376 0.152939
R20603 gnd.n7378 gnd.n7377 0.152939
R20604 gnd.n7378 gnd.n220 0.152939
R20605 gnd.n7392 gnd.n220 0.152939
R20606 gnd.n7393 gnd.n7392 0.152939
R20607 gnd.n7462 gnd.n7393 0.152939
R20608 gnd.n7462 gnd.n7461 0.152939
R20609 gnd.n7461 gnd.n7460 0.152939
R20610 gnd.n7460 gnd.n7394 0.152939
R20611 gnd.n7456 gnd.n7394 0.152939
R20612 gnd.n7455 gnd.n7396 0.152939
R20613 gnd.n7451 gnd.n7396 0.152939
R20614 gnd.n7451 gnd.n7450 0.152939
R20615 gnd.n7450 gnd.n7449 0.152939
R20616 gnd.n7449 gnd.n7402 0.152939
R20617 gnd.n7445 gnd.n7402 0.152939
R20618 gnd.n7445 gnd.n7444 0.152939
R20619 gnd.n7444 gnd.n7443 0.152939
R20620 gnd.n7443 gnd.n7410 0.152939
R20621 gnd.n7439 gnd.n7410 0.152939
R20622 gnd.n7439 gnd.n7438 0.152939
R20623 gnd.n7438 gnd.n7437 0.152939
R20624 gnd.n7437 gnd.n7418 0.152939
R20625 gnd.n7433 gnd.n7418 0.152939
R20626 gnd.n7433 gnd.n7432 0.152939
R20627 gnd.n7432 gnd.n7431 0.152939
R20628 gnd.n7431 gnd.n121 0.152939
R20629 gnd.n7557 gnd.n121 0.152939
R20630 gnd.n6803 gnd.n591 0.152939
R20631 gnd.n6804 gnd.n6803 0.152939
R20632 gnd.n7019 gnd.n6804 0.152939
R20633 gnd.n7019 gnd.n7018 0.152939
R20634 gnd.n7018 gnd.n7017 0.152939
R20635 gnd.n7017 gnd.n6805 0.152939
R20636 gnd.n7013 gnd.n6805 0.152939
R20637 gnd.n7013 gnd.n7012 0.152939
R20638 gnd.n7012 gnd.n7011 0.152939
R20639 gnd.n7011 gnd.n6809 0.152939
R20640 gnd.n7007 gnd.n6809 0.152939
R20641 gnd.n7007 gnd.n7006 0.152939
R20642 gnd.n7006 gnd.n7005 0.152939
R20643 gnd.n7005 gnd.n6959 0.152939
R20644 gnd.n7001 gnd.n6959 0.152939
R20645 gnd.n7001 gnd.n7000 0.152939
R20646 gnd.n7000 gnd.n6999 0.152939
R20647 gnd.n6999 gnd.n6963 0.152939
R20648 gnd.n6995 gnd.n6963 0.152939
R20649 gnd.n6995 gnd.n6994 0.152939
R20650 gnd.n6994 gnd.n6993 0.152939
R20651 gnd.n6993 gnd.n6967 0.152939
R20652 gnd.n6989 gnd.n6967 0.152939
R20653 gnd.n6989 gnd.n6988 0.152939
R20654 gnd.n6988 gnd.n6987 0.152939
R20655 gnd.n6987 gnd.n6971 0.152939
R20656 gnd.n6983 gnd.n6971 0.152939
R20657 gnd.n6983 gnd.n6982 0.152939
R20658 gnd.n6982 gnd.n6981 0.152939
R20659 gnd.n6981 gnd.n6975 0.152939
R20660 gnd.n6975 gnd.n79 0.152939
R20661 gnd.n7606 gnd.n79 0.152939
R20662 gnd.n7606 gnd.n7605 0.152939
R20663 gnd.n7605 gnd.n81 0.152939
R20664 gnd.n7601 gnd.n81 0.152939
R20665 gnd.n7601 gnd.n7600 0.152939
R20666 gnd.n7600 gnd.n7599 0.152939
R20667 gnd.n7599 gnd.n86 0.152939
R20668 gnd.n7595 gnd.n86 0.152939
R20669 gnd.n7595 gnd.n7594 0.152939
R20670 gnd.n7594 gnd.n7593 0.152939
R20671 gnd.n7593 gnd.n91 0.152939
R20672 gnd.n7589 gnd.n91 0.152939
R20673 gnd.n7589 gnd.n7588 0.152939
R20674 gnd.n7588 gnd.n7587 0.152939
R20675 gnd.n7587 gnd.n96 0.152939
R20676 gnd.n7583 gnd.n96 0.152939
R20677 gnd.n7583 gnd.n7582 0.152939
R20678 gnd.n7582 gnd.n7581 0.152939
R20679 gnd.n7581 gnd.n101 0.152939
R20680 gnd.n7577 gnd.n101 0.152939
R20681 gnd.n7577 gnd.n7576 0.152939
R20682 gnd.n7576 gnd.n7575 0.152939
R20683 gnd.n7575 gnd.n106 0.152939
R20684 gnd.n7571 gnd.n106 0.152939
R20685 gnd.n7571 gnd.n7570 0.152939
R20686 gnd.n7570 gnd.n7569 0.152939
R20687 gnd.n7569 gnd.n111 0.152939
R20688 gnd.n7565 gnd.n111 0.152939
R20689 gnd.n7565 gnd.n7564 0.152939
R20690 gnd.n7564 gnd.n7563 0.152939
R20691 gnd.n7563 gnd.n116 0.152939
R20692 gnd.n7559 gnd.n116 0.152939
R20693 gnd.n7559 gnd.n7558 0.152939
R20694 gnd.n1282 gnd.n1281 0.151415
R20695 gnd.n4713 gnd.n4448 0.151415
R20696 gnd.n4097 gnd.n4043 0.145814
R20697 gnd.n4097 gnd.n4096 0.145814
R20698 gnd.n3098 gnd.n3097 0.0767195
R20699 gnd.n3097 gnd.n3096 0.0767195
R20700 gnd.n6055 gnd.n6054 0.063
R20701 gnd.n7153 gnd.n455 0.063
R20702 gnd.n3664 gnd.n2268 0.0477147
R20703 gnd.n2861 gnd.n2749 0.0442063
R20704 gnd.n2862 gnd.n2861 0.0442063
R20705 gnd.n2863 gnd.n2862 0.0442063
R20706 gnd.n2863 gnd.n2738 0.0442063
R20707 gnd.n2877 gnd.n2738 0.0442063
R20708 gnd.n2878 gnd.n2877 0.0442063
R20709 gnd.n2879 gnd.n2878 0.0442063
R20710 gnd.n2879 gnd.n2725 0.0442063
R20711 gnd.n2923 gnd.n2725 0.0442063
R20712 gnd.n2924 gnd.n2923 0.0442063
R20713 gnd.n2926 gnd.n2659 0.0344674
R20714 gnd.n1280 gnd.n504 0.0343753
R20715 gnd.n4717 gnd.n4716 0.0343753
R20716 gnd.n2946 gnd.n2945 0.0269946
R20717 gnd.n2948 gnd.n2947 0.0269946
R20718 gnd.n2654 gnd.n2652 0.0269946
R20719 gnd.n2958 gnd.n2956 0.0269946
R20720 gnd.n2957 gnd.n2633 0.0269946
R20721 gnd.n2977 gnd.n2976 0.0269946
R20722 gnd.n2979 gnd.n2978 0.0269946
R20723 gnd.n2628 gnd.n2627 0.0269946
R20724 gnd.n2989 gnd.n2623 0.0269946
R20725 gnd.n2988 gnd.n2625 0.0269946
R20726 gnd.n2624 gnd.n2606 0.0269946
R20727 gnd.n3009 gnd.n2607 0.0269946
R20728 gnd.n3008 gnd.n2608 0.0269946
R20729 gnd.n3042 gnd.n2583 0.0269946
R20730 gnd.n3044 gnd.n3043 0.0269946
R20731 gnd.n3045 gnd.n2530 0.0269946
R20732 gnd.n2578 gnd.n2531 0.0269946
R20733 gnd.n2580 gnd.n2532 0.0269946
R20734 gnd.n3055 gnd.n3054 0.0269946
R20735 gnd.n3057 gnd.n3056 0.0269946
R20736 gnd.n3058 gnd.n2552 0.0269946
R20737 gnd.n3060 gnd.n2553 0.0269946
R20738 gnd.n3063 gnd.n2554 0.0269946
R20739 gnd.n3066 gnd.n3065 0.0269946
R20740 gnd.n3068 gnd.n3067 0.0269946
R20741 gnd.n3133 gnd.n2441 0.0269946
R20742 gnd.n3135 gnd.n3134 0.0269946
R20743 gnd.n3144 gnd.n2434 0.0269946
R20744 gnd.n3146 gnd.n3145 0.0269946
R20745 gnd.n3147 gnd.n2432 0.0269946
R20746 gnd.n3154 gnd.n3150 0.0269946
R20747 gnd.n3153 gnd.n3152 0.0269946
R20748 gnd.n3151 gnd.n2411 0.0269946
R20749 gnd.n3176 gnd.n2412 0.0269946
R20750 gnd.n3175 gnd.n2413 0.0269946
R20751 gnd.n3218 gnd.n2386 0.0269946
R20752 gnd.n3220 gnd.n3219 0.0269946
R20753 gnd.n3229 gnd.n2379 0.0269946
R20754 gnd.n3231 gnd.n3230 0.0269946
R20755 gnd.n3232 gnd.n2377 0.0269946
R20756 gnd.n3239 gnd.n3235 0.0269946
R20757 gnd.n3238 gnd.n3237 0.0269946
R20758 gnd.n3236 gnd.n2356 0.0269946
R20759 gnd.n3261 gnd.n2357 0.0269946
R20760 gnd.n3260 gnd.n2358 0.0269946
R20761 gnd.n3307 gnd.n2332 0.0269946
R20762 gnd.n3309 gnd.n3308 0.0269946
R20763 gnd.n3318 gnd.n2325 0.0269946
R20764 gnd.n3577 gnd.n2323 0.0269946
R20765 gnd.n3582 gnd.n3580 0.0269946
R20766 gnd.n3581 gnd.n2304 0.0269946
R20767 gnd.n3606 gnd.n3605 0.0269946
R20768 gnd.n7150 gnd.n455 0.0245515
R20769 gnd.n6054 gnd.n1099 0.0245515
R20770 gnd.n2926 gnd.n2925 0.0202011
R20771 gnd.n7150 gnd.n7149 0.0174377
R20772 gnd.n7149 gnd.n458 0.0174377
R20773 gnd.n7146 gnd.n458 0.0174377
R20774 gnd.n7146 gnd.n7145 0.0174377
R20775 gnd.n7145 gnd.n462 0.0174377
R20776 gnd.n7142 gnd.n462 0.0174377
R20777 gnd.n7142 gnd.n7141 0.0174377
R20778 gnd.n7141 gnd.n466 0.0174377
R20779 gnd.n7138 gnd.n466 0.0174377
R20780 gnd.n7138 gnd.n7137 0.0174377
R20781 gnd.n7137 gnd.n470 0.0174377
R20782 gnd.n7134 gnd.n470 0.0174377
R20783 gnd.n7134 gnd.n7133 0.0174377
R20784 gnd.n7133 gnd.n474 0.0174377
R20785 gnd.n7130 gnd.n474 0.0174377
R20786 gnd.n7130 gnd.n7129 0.0174377
R20787 gnd.n7129 gnd.n478 0.0174377
R20788 gnd.n7126 gnd.n478 0.0174377
R20789 gnd.n7126 gnd.n7125 0.0174377
R20790 gnd.n7125 gnd.n482 0.0174377
R20791 gnd.n7122 gnd.n482 0.0174377
R20792 gnd.n7122 gnd.n7121 0.0174377
R20793 gnd.n7121 gnd.n486 0.0174377
R20794 gnd.n7118 gnd.n486 0.0174377
R20795 gnd.n7118 gnd.n7117 0.0174377
R20796 gnd.n7117 gnd.n490 0.0174377
R20797 gnd.n7114 gnd.n490 0.0174377
R20798 gnd.n7114 gnd.n7113 0.0174377
R20799 gnd.n7113 gnd.n494 0.0174377
R20800 gnd.n7110 gnd.n494 0.0174377
R20801 gnd.n7110 gnd.n7109 0.0174377
R20802 gnd.n7109 gnd.n500 0.0174377
R20803 gnd.n7106 gnd.n500 0.0174377
R20804 gnd.n7106 gnd.n7105 0.0174377
R20805 gnd.n7105 gnd.n504 0.0174377
R20806 gnd.n4494 gnd.n1099 0.0174377
R20807 gnd.n4496 gnd.n4494 0.0174377
R20808 gnd.n4760 gnd.n4496 0.0174377
R20809 gnd.n4760 gnd.n4759 0.0174377
R20810 gnd.n4759 gnd.n4497 0.0174377
R20811 gnd.n4756 gnd.n4497 0.0174377
R20812 gnd.n4756 gnd.n4755 0.0174377
R20813 gnd.n4755 gnd.n4508 0.0174377
R20814 gnd.n4752 gnd.n4508 0.0174377
R20815 gnd.n4752 gnd.n4751 0.0174377
R20816 gnd.n4751 gnd.n4513 0.0174377
R20817 gnd.n4748 gnd.n4513 0.0174377
R20818 gnd.n4748 gnd.n4747 0.0174377
R20819 gnd.n4747 gnd.n4519 0.0174377
R20820 gnd.n4744 gnd.n4519 0.0174377
R20821 gnd.n4744 gnd.n4743 0.0174377
R20822 gnd.n4743 gnd.n4523 0.0174377
R20823 gnd.n4740 gnd.n4523 0.0174377
R20824 gnd.n4740 gnd.n4739 0.0174377
R20825 gnd.n4739 gnd.n4530 0.0174377
R20826 gnd.n4736 gnd.n4530 0.0174377
R20827 gnd.n4736 gnd.n4735 0.0174377
R20828 gnd.n4735 gnd.n4536 0.0174377
R20829 gnd.n4732 gnd.n4536 0.0174377
R20830 gnd.n4732 gnd.n4731 0.0174377
R20831 gnd.n4731 gnd.n4542 0.0174377
R20832 gnd.n4728 gnd.n4542 0.0174377
R20833 gnd.n4728 gnd.n4727 0.0174377
R20834 gnd.n4727 gnd.n4546 0.0174377
R20835 gnd.n4724 gnd.n4546 0.0174377
R20836 gnd.n4724 gnd.n4723 0.0174377
R20837 gnd.n4723 gnd.n4557 0.0174377
R20838 gnd.n4720 gnd.n4557 0.0174377
R20839 gnd.n4720 gnd.n4719 0.0174377
R20840 gnd.n4719 gnd.n4717 0.0174377
R20841 gnd.n2925 gnd.n2924 0.0148637
R20842 gnd.n3575 gnd.n3319 0.0144266
R20843 gnd.n3576 gnd.n3575 0.0130679
R20844 gnd.n2945 gnd.n2659 0.00797283
R20845 gnd.n2947 gnd.n2946 0.00797283
R20846 gnd.n2948 gnd.n2654 0.00797283
R20847 gnd.n2956 gnd.n2652 0.00797283
R20848 gnd.n2958 gnd.n2957 0.00797283
R20849 gnd.n2976 gnd.n2633 0.00797283
R20850 gnd.n2978 gnd.n2977 0.00797283
R20851 gnd.n2979 gnd.n2628 0.00797283
R20852 gnd.n2627 gnd.n2623 0.00797283
R20853 gnd.n2989 gnd.n2988 0.00797283
R20854 gnd.n2625 gnd.n2624 0.00797283
R20855 gnd.n2607 gnd.n2606 0.00797283
R20856 gnd.n3009 gnd.n3008 0.00797283
R20857 gnd.n2608 gnd.n2583 0.00797283
R20858 gnd.n3043 gnd.n3042 0.00797283
R20859 gnd.n3045 gnd.n3044 0.00797283
R20860 gnd.n2578 gnd.n2530 0.00797283
R20861 gnd.n2580 gnd.n2531 0.00797283
R20862 gnd.n3054 gnd.n2532 0.00797283
R20863 gnd.n3056 gnd.n3055 0.00797283
R20864 gnd.n3058 gnd.n3057 0.00797283
R20865 gnd.n3060 gnd.n2552 0.00797283
R20866 gnd.n3063 gnd.n2553 0.00797283
R20867 gnd.n3065 gnd.n2554 0.00797283
R20868 gnd.n3068 gnd.n3066 0.00797283
R20869 gnd.n3067 gnd.n2441 0.00797283
R20870 gnd.n3135 gnd.n3133 0.00797283
R20871 gnd.n3134 gnd.n2434 0.00797283
R20872 gnd.n3145 gnd.n3144 0.00797283
R20873 gnd.n3147 gnd.n3146 0.00797283
R20874 gnd.n3150 gnd.n2432 0.00797283
R20875 gnd.n3154 gnd.n3153 0.00797283
R20876 gnd.n3152 gnd.n3151 0.00797283
R20877 gnd.n2412 gnd.n2411 0.00797283
R20878 gnd.n3176 gnd.n3175 0.00797283
R20879 gnd.n2413 gnd.n2386 0.00797283
R20880 gnd.n3220 gnd.n3218 0.00797283
R20881 gnd.n3219 gnd.n2379 0.00797283
R20882 gnd.n3230 gnd.n3229 0.00797283
R20883 gnd.n3232 gnd.n3231 0.00797283
R20884 gnd.n3235 gnd.n2377 0.00797283
R20885 gnd.n3239 gnd.n3238 0.00797283
R20886 gnd.n3237 gnd.n3236 0.00797283
R20887 gnd.n2357 gnd.n2356 0.00797283
R20888 gnd.n3261 gnd.n3260 0.00797283
R20889 gnd.n2358 gnd.n2332 0.00797283
R20890 gnd.n3309 gnd.n3307 0.00797283
R20891 gnd.n3308 gnd.n2325 0.00797283
R20892 gnd.n3319 gnd.n3318 0.00797283
R20893 gnd.n3577 gnd.n3576 0.00797283
R20894 gnd.n3580 gnd.n2323 0.00797283
R20895 gnd.n3582 gnd.n3581 0.00797283
R20896 gnd.n3605 gnd.n2304 0.00797283
R20897 gnd.n3606 gnd.n2268 0.00797283
R20898 gnd.n7282 gnd.n325 0.00433921
R20899 gnd.n4317 gnd.n2105 0.00433921
R20900 gnd.n7272 gnd.n334 0.00335063
R20901 gnd.n7273 gnd.n7272 0.00335063
R20902 gnd.n7274 gnd.n7273 0.00335063
R20903 gnd.n7274 gnd.n316 0.00335063
R20904 gnd.n7288 gnd.n316 0.00335063
R20905 gnd.n7289 gnd.n7288 0.00335063
R20906 gnd.n7290 gnd.n7289 0.00335063
R20907 gnd.n7290 gnd.n302 0.00335063
R20908 gnd.n7304 gnd.n302 0.00335063
R20909 gnd.n7305 gnd.n7304 0.00335063
R20910 gnd.n4307 gnd.n2114 0.00335063
R20911 gnd.n4308 gnd.n4307 0.00335063
R20912 gnd.n4309 gnd.n4308 0.00335063
R20913 gnd.n4309 gnd.n2096 0.00335063
R20914 gnd.n4323 gnd.n2096 0.00335063
R20915 gnd.n4324 gnd.n4323 0.00335063
R20916 gnd.n4325 gnd.n4324 0.00335063
R20917 gnd.n4325 gnd.n2081 0.00335063
R20918 gnd.n4339 gnd.n2081 0.00335063
R20919 gnd.n4340 gnd.n4339 0.00335063
R20920 gnd.n1281 gnd.n1280 0.000838753
R20921 gnd.n4716 gnd.n4448 0.000838753
R20922 outputibias.n27 outputibias.n1 289.615
R20923 outputibias.n58 outputibias.n32 289.615
R20924 outputibias.n90 outputibias.n64 289.615
R20925 outputibias.n122 outputibias.n96 289.615
R20926 outputibias.n28 outputibias.n27 185
R20927 outputibias.n26 outputibias.n25 185
R20928 outputibias.n5 outputibias.n4 185
R20929 outputibias.n20 outputibias.n19 185
R20930 outputibias.n18 outputibias.n17 185
R20931 outputibias.n9 outputibias.n8 185
R20932 outputibias.n12 outputibias.n11 185
R20933 outputibias.n59 outputibias.n58 185
R20934 outputibias.n57 outputibias.n56 185
R20935 outputibias.n36 outputibias.n35 185
R20936 outputibias.n51 outputibias.n50 185
R20937 outputibias.n49 outputibias.n48 185
R20938 outputibias.n40 outputibias.n39 185
R20939 outputibias.n43 outputibias.n42 185
R20940 outputibias.n91 outputibias.n90 185
R20941 outputibias.n89 outputibias.n88 185
R20942 outputibias.n68 outputibias.n67 185
R20943 outputibias.n83 outputibias.n82 185
R20944 outputibias.n81 outputibias.n80 185
R20945 outputibias.n72 outputibias.n71 185
R20946 outputibias.n75 outputibias.n74 185
R20947 outputibias.n123 outputibias.n122 185
R20948 outputibias.n121 outputibias.n120 185
R20949 outputibias.n100 outputibias.n99 185
R20950 outputibias.n115 outputibias.n114 185
R20951 outputibias.n113 outputibias.n112 185
R20952 outputibias.n104 outputibias.n103 185
R20953 outputibias.n107 outputibias.n106 185
R20954 outputibias.n0 outputibias.t8 178.945
R20955 outputibias.n133 outputibias.t9 177.018
R20956 outputibias.n132 outputibias.t11 177.018
R20957 outputibias.n0 outputibias.t10 177.018
R20958 outputibias.t5 outputibias.n10 147.661
R20959 outputibias.t3 outputibias.n41 147.661
R20960 outputibias.t1 outputibias.n73 147.661
R20961 outputibias.t7 outputibias.n105 147.661
R20962 outputibias.n128 outputibias.t4 132.363
R20963 outputibias.n128 outputibias.t2 130.436
R20964 outputibias.n129 outputibias.t0 130.436
R20965 outputibias.n130 outputibias.t6 130.436
R20966 outputibias.n27 outputibias.n26 104.615
R20967 outputibias.n26 outputibias.n4 104.615
R20968 outputibias.n19 outputibias.n4 104.615
R20969 outputibias.n19 outputibias.n18 104.615
R20970 outputibias.n18 outputibias.n8 104.615
R20971 outputibias.n11 outputibias.n8 104.615
R20972 outputibias.n58 outputibias.n57 104.615
R20973 outputibias.n57 outputibias.n35 104.615
R20974 outputibias.n50 outputibias.n35 104.615
R20975 outputibias.n50 outputibias.n49 104.615
R20976 outputibias.n49 outputibias.n39 104.615
R20977 outputibias.n42 outputibias.n39 104.615
R20978 outputibias.n90 outputibias.n89 104.615
R20979 outputibias.n89 outputibias.n67 104.615
R20980 outputibias.n82 outputibias.n67 104.615
R20981 outputibias.n82 outputibias.n81 104.615
R20982 outputibias.n81 outputibias.n71 104.615
R20983 outputibias.n74 outputibias.n71 104.615
R20984 outputibias.n122 outputibias.n121 104.615
R20985 outputibias.n121 outputibias.n99 104.615
R20986 outputibias.n114 outputibias.n99 104.615
R20987 outputibias.n114 outputibias.n113 104.615
R20988 outputibias.n113 outputibias.n103 104.615
R20989 outputibias.n106 outputibias.n103 104.615
R20990 outputibias.n63 outputibias.n31 95.6354
R20991 outputibias.n63 outputibias.n62 94.6732
R20992 outputibias.n95 outputibias.n94 94.6732
R20993 outputibias.n127 outputibias.n126 94.6732
R20994 outputibias.n11 outputibias.t5 52.3082
R20995 outputibias.n42 outputibias.t3 52.3082
R20996 outputibias.n74 outputibias.t1 52.3082
R20997 outputibias.n106 outputibias.t7 52.3082
R20998 outputibias.n12 outputibias.n10 15.6674
R20999 outputibias.n43 outputibias.n41 15.6674
R21000 outputibias.n75 outputibias.n73 15.6674
R21001 outputibias.n107 outputibias.n105 15.6674
R21002 outputibias.n13 outputibias.n9 12.8005
R21003 outputibias.n44 outputibias.n40 12.8005
R21004 outputibias.n76 outputibias.n72 12.8005
R21005 outputibias.n108 outputibias.n104 12.8005
R21006 outputibias.n17 outputibias.n16 12.0247
R21007 outputibias.n48 outputibias.n47 12.0247
R21008 outputibias.n80 outputibias.n79 12.0247
R21009 outputibias.n112 outputibias.n111 12.0247
R21010 outputibias.n20 outputibias.n7 11.249
R21011 outputibias.n51 outputibias.n38 11.249
R21012 outputibias.n83 outputibias.n70 11.249
R21013 outputibias.n115 outputibias.n102 11.249
R21014 outputibias.n21 outputibias.n5 10.4732
R21015 outputibias.n52 outputibias.n36 10.4732
R21016 outputibias.n84 outputibias.n68 10.4732
R21017 outputibias.n116 outputibias.n100 10.4732
R21018 outputibias.n25 outputibias.n24 9.69747
R21019 outputibias.n56 outputibias.n55 9.69747
R21020 outputibias.n88 outputibias.n87 9.69747
R21021 outputibias.n120 outputibias.n119 9.69747
R21022 outputibias.n31 outputibias.n30 9.45567
R21023 outputibias.n62 outputibias.n61 9.45567
R21024 outputibias.n94 outputibias.n93 9.45567
R21025 outputibias.n126 outputibias.n125 9.45567
R21026 outputibias.n30 outputibias.n29 9.3005
R21027 outputibias.n3 outputibias.n2 9.3005
R21028 outputibias.n24 outputibias.n23 9.3005
R21029 outputibias.n22 outputibias.n21 9.3005
R21030 outputibias.n7 outputibias.n6 9.3005
R21031 outputibias.n16 outputibias.n15 9.3005
R21032 outputibias.n14 outputibias.n13 9.3005
R21033 outputibias.n61 outputibias.n60 9.3005
R21034 outputibias.n34 outputibias.n33 9.3005
R21035 outputibias.n55 outputibias.n54 9.3005
R21036 outputibias.n53 outputibias.n52 9.3005
R21037 outputibias.n38 outputibias.n37 9.3005
R21038 outputibias.n47 outputibias.n46 9.3005
R21039 outputibias.n45 outputibias.n44 9.3005
R21040 outputibias.n93 outputibias.n92 9.3005
R21041 outputibias.n66 outputibias.n65 9.3005
R21042 outputibias.n87 outputibias.n86 9.3005
R21043 outputibias.n85 outputibias.n84 9.3005
R21044 outputibias.n70 outputibias.n69 9.3005
R21045 outputibias.n79 outputibias.n78 9.3005
R21046 outputibias.n77 outputibias.n76 9.3005
R21047 outputibias.n125 outputibias.n124 9.3005
R21048 outputibias.n98 outputibias.n97 9.3005
R21049 outputibias.n119 outputibias.n118 9.3005
R21050 outputibias.n117 outputibias.n116 9.3005
R21051 outputibias.n102 outputibias.n101 9.3005
R21052 outputibias.n111 outputibias.n110 9.3005
R21053 outputibias.n109 outputibias.n108 9.3005
R21054 outputibias.n28 outputibias.n3 8.92171
R21055 outputibias.n59 outputibias.n34 8.92171
R21056 outputibias.n91 outputibias.n66 8.92171
R21057 outputibias.n123 outputibias.n98 8.92171
R21058 outputibias.n29 outputibias.n1 8.14595
R21059 outputibias.n60 outputibias.n32 8.14595
R21060 outputibias.n92 outputibias.n64 8.14595
R21061 outputibias.n124 outputibias.n96 8.14595
R21062 outputibias.n31 outputibias.n1 5.81868
R21063 outputibias.n62 outputibias.n32 5.81868
R21064 outputibias.n94 outputibias.n64 5.81868
R21065 outputibias.n126 outputibias.n96 5.81868
R21066 outputibias.n131 outputibias.n130 5.20947
R21067 outputibias.n29 outputibias.n28 5.04292
R21068 outputibias.n60 outputibias.n59 5.04292
R21069 outputibias.n92 outputibias.n91 5.04292
R21070 outputibias.n124 outputibias.n123 5.04292
R21071 outputibias.n131 outputibias.n127 4.42209
R21072 outputibias.n14 outputibias.n10 4.38594
R21073 outputibias.n45 outputibias.n41 4.38594
R21074 outputibias.n77 outputibias.n73 4.38594
R21075 outputibias.n109 outputibias.n105 4.38594
R21076 outputibias.n132 outputibias.n131 4.28454
R21077 outputibias.n25 outputibias.n3 4.26717
R21078 outputibias.n56 outputibias.n34 4.26717
R21079 outputibias.n88 outputibias.n66 4.26717
R21080 outputibias.n120 outputibias.n98 4.26717
R21081 outputibias.n24 outputibias.n5 3.49141
R21082 outputibias.n55 outputibias.n36 3.49141
R21083 outputibias.n87 outputibias.n68 3.49141
R21084 outputibias.n119 outputibias.n100 3.49141
R21085 outputibias.n21 outputibias.n20 2.71565
R21086 outputibias.n52 outputibias.n51 2.71565
R21087 outputibias.n84 outputibias.n83 2.71565
R21088 outputibias.n116 outputibias.n115 2.71565
R21089 outputibias.n17 outputibias.n7 1.93989
R21090 outputibias.n48 outputibias.n38 1.93989
R21091 outputibias.n80 outputibias.n70 1.93989
R21092 outputibias.n112 outputibias.n102 1.93989
R21093 outputibias.n130 outputibias.n129 1.9266
R21094 outputibias.n129 outputibias.n128 1.9266
R21095 outputibias.n133 outputibias.n132 1.92658
R21096 outputibias.n134 outputibias.n133 1.29913
R21097 outputibias.n16 outputibias.n9 1.16414
R21098 outputibias.n47 outputibias.n40 1.16414
R21099 outputibias.n79 outputibias.n72 1.16414
R21100 outputibias.n111 outputibias.n104 1.16414
R21101 outputibias.n127 outputibias.n95 0.962709
R21102 outputibias.n95 outputibias.n63 0.962709
R21103 outputibias.n13 outputibias.n12 0.388379
R21104 outputibias.n44 outputibias.n43 0.388379
R21105 outputibias.n76 outputibias.n75 0.388379
R21106 outputibias.n108 outputibias.n107 0.388379
R21107 outputibias.n134 outputibias.n0 0.337251
R21108 outputibias outputibias.n134 0.302375
R21109 outputibias.n30 outputibias.n2 0.155672
R21110 outputibias.n23 outputibias.n2 0.155672
R21111 outputibias.n23 outputibias.n22 0.155672
R21112 outputibias.n22 outputibias.n6 0.155672
R21113 outputibias.n15 outputibias.n6 0.155672
R21114 outputibias.n15 outputibias.n14 0.155672
R21115 outputibias.n61 outputibias.n33 0.155672
R21116 outputibias.n54 outputibias.n33 0.155672
R21117 outputibias.n54 outputibias.n53 0.155672
R21118 outputibias.n53 outputibias.n37 0.155672
R21119 outputibias.n46 outputibias.n37 0.155672
R21120 outputibias.n46 outputibias.n45 0.155672
R21121 outputibias.n93 outputibias.n65 0.155672
R21122 outputibias.n86 outputibias.n65 0.155672
R21123 outputibias.n86 outputibias.n85 0.155672
R21124 outputibias.n85 outputibias.n69 0.155672
R21125 outputibias.n78 outputibias.n69 0.155672
R21126 outputibias.n78 outputibias.n77 0.155672
R21127 outputibias.n125 outputibias.n97 0.155672
R21128 outputibias.n118 outputibias.n97 0.155672
R21129 outputibias.n118 outputibias.n117 0.155672
R21130 outputibias.n117 outputibias.n101 0.155672
R21131 outputibias.n110 outputibias.n101 0.155672
R21132 outputibias.n110 outputibias.n109 0.155672
R21133 commonsourceibias.n281 commonsourceibias.t101 222.032
R21134 commonsourceibias.n44 commonsourceibias.t78 222.032
R21135 commonsourceibias.n166 commonsourceibias.t118 222.032
R21136 commonsourceibias.n643 commonsourceibias.t107 222.032
R21137 commonsourceibias.n413 commonsourceibias.t30 222.032
R21138 commonsourceibias.n529 commonsourceibias.t123 222.032
R21139 commonsourceibias.n364 commonsourceibias.t100 207.983
R21140 commonsourceibias.n127 commonsourceibias.t74 207.983
R21141 commonsourceibias.n249 commonsourceibias.t115 207.983
R21142 commonsourceibias.n731 commonsourceibias.t122 207.983
R21143 commonsourceibias.n501 commonsourceibias.t12 207.983
R21144 commonsourceibias.n616 commonsourceibias.t140 207.983
R21145 commonsourceibias.n280 commonsourceibias.t87 168.701
R21146 commonsourceibias.n286 commonsourceibias.t129 168.701
R21147 commonsourceibias.n292 commonsourceibias.t110 168.701
R21148 commonsourceibias.n276 commonsourceibias.t93 168.701
R21149 commonsourceibias.n300 commonsourceibias.t95 168.701
R21150 commonsourceibias.n306 commonsourceibias.t121 168.701
R21151 commonsourceibias.n271 commonsourceibias.t102 168.701
R21152 commonsourceibias.n314 commonsourceibias.t108 168.701
R21153 commonsourceibias.n320 commonsourceibias.t159 168.701
R21154 commonsourceibias.n266 commonsourceibias.t138 168.701
R21155 commonsourceibias.n328 commonsourceibias.t117 168.701
R21156 commonsourceibias.n334 commonsourceibias.t83 168.701
R21157 commonsourceibias.n261 commonsourceibias.t86 168.701
R21158 commonsourceibias.n342 commonsourceibias.t127 168.701
R21159 commonsourceibias.n348 commonsourceibias.t109 168.701
R21160 commonsourceibias.n256 commonsourceibias.t91 168.701
R21161 commonsourceibias.n356 commonsourceibias.t137 168.701
R21162 commonsourceibias.n362 commonsourceibias.t119 168.701
R21163 commonsourceibias.n125 commonsourceibias.t20 168.701
R21164 commonsourceibias.n119 commonsourceibias.t50 168.701
R21165 commonsourceibias.n19 commonsourceibias.t8 168.701
R21166 commonsourceibias.n111 commonsourceibias.t36 168.701
R21167 commonsourceibias.n105 commonsourceibias.t76 168.701
R21168 commonsourceibias.n24 commonsourceibias.t24 168.701
R21169 commonsourceibias.n97 commonsourceibias.t34 168.701
R21170 commonsourceibias.n91 commonsourceibias.t10 168.701
R21171 commonsourceibias.n29 commonsourceibias.t40 168.701
R21172 commonsourceibias.n83 commonsourceibias.t56 168.701
R21173 commonsourceibias.n77 commonsourceibias.t26 168.701
R21174 commonsourceibias.n34 commonsourceibias.t38 168.701
R21175 commonsourceibias.n69 commonsourceibias.t70 168.701
R21176 commonsourceibias.n63 commonsourceibias.t18 168.701
R21177 commonsourceibias.n39 commonsourceibias.t22 168.701
R21178 commonsourceibias.n55 commonsourceibias.t52 168.701
R21179 commonsourceibias.n49 commonsourceibias.t4 168.701
R21180 commonsourceibias.n43 commonsourceibias.t46 168.701
R21181 commonsourceibias.n247 commonsourceibias.t136 168.701
R21182 commonsourceibias.n241 commonsourceibias.t151 168.701
R21183 commonsourceibias.n5 commonsourceibias.t104 168.701
R21184 commonsourceibias.n233 commonsourceibias.t126 168.701
R21185 commonsourceibias.n227 commonsourceibias.t144 168.701
R21186 commonsourceibias.n10 commonsourceibias.t96 168.701
R21187 commonsourceibias.n219 commonsourceibias.t94 168.701
R21188 commonsourceibias.n213 commonsourceibias.t134 168.701
R21189 commonsourceibias.n150 commonsourceibias.t152 168.701
R21190 commonsourceibias.n151 commonsourceibias.t88 168.701
R21191 commonsourceibias.n153 commonsourceibias.t124 168.701
R21192 commonsourceibias.n155 commonsourceibias.t120 168.701
R21193 commonsourceibias.n191 commonsourceibias.t139 168.701
R21194 commonsourceibias.n185 commonsourceibias.t112 168.701
R21195 commonsourceibias.n161 commonsourceibias.t106 168.701
R21196 commonsourceibias.n177 commonsourceibias.t128 168.701
R21197 commonsourceibias.n171 commonsourceibias.t145 168.701
R21198 commonsourceibias.n165 commonsourceibias.t99 168.701
R21199 commonsourceibias.n642 commonsourceibias.t90 168.701
R21200 commonsourceibias.n648 commonsourceibias.t135 168.701
R21201 commonsourceibias.n654 commonsourceibias.t116 168.701
R21202 commonsourceibias.n656 commonsourceibias.t98 168.701
R21203 commonsourceibias.n663 commonsourceibias.t92 168.701
R21204 commonsourceibias.n669 commonsourceibias.t146 168.701
R21205 commonsourceibias.n671 commonsourceibias.t125 168.701
R21206 commonsourceibias.n678 commonsourceibias.t132 168.701
R21207 commonsourceibias.n684 commonsourceibias.t153 168.701
R21208 commonsourceibias.n686 commonsourceibias.t157 168.701
R21209 commonsourceibias.n693 commonsourceibias.t142 168.701
R21210 commonsourceibias.n699 commonsourceibias.t97 168.701
R21211 commonsourceibias.n701 commonsourceibias.t81 168.701
R21212 commonsourceibias.n708 commonsourceibias.t149 168.701
R21213 commonsourceibias.n714 commonsourceibias.t131 168.701
R21214 commonsourceibias.n716 commonsourceibias.t111 168.701
R21215 commonsourceibias.n723 commonsourceibias.t156 168.701
R21216 commonsourceibias.n729 commonsourceibias.t141 168.701
R21217 commonsourceibias.n412 commonsourceibias.t2 168.701
R21218 commonsourceibias.n418 commonsourceibias.t48 168.701
R21219 commonsourceibias.n424 commonsourceibias.t14 168.701
R21220 commonsourceibias.n426 commonsourceibias.t68 168.701
R21221 commonsourceibias.n433 commonsourceibias.t66 168.701
R21222 commonsourceibias.n439 commonsourceibias.t6 168.701
R21223 commonsourceibias.n441 commonsourceibias.t62 168.701
R21224 commonsourceibias.n448 commonsourceibias.t54 168.701
R21225 commonsourceibias.n454 commonsourceibias.t72 168.701
R21226 commonsourceibias.n456 commonsourceibias.t64 168.701
R21227 commonsourceibias.n463 commonsourceibias.t32 168.701
R21228 commonsourceibias.n469 commonsourceibias.t58 168.701
R21229 commonsourceibias.n471 commonsourceibias.t44 168.701
R21230 commonsourceibias.n478 commonsourceibias.t16 168.701
R21231 commonsourceibias.n484 commonsourceibias.t60 168.701
R21232 commonsourceibias.n486 commonsourceibias.t28 168.701
R21233 commonsourceibias.n493 commonsourceibias.t0 168.701
R21234 commonsourceibias.n499 commonsourceibias.t42 168.701
R21235 commonsourceibias.n614 commonsourceibias.t154 168.701
R21236 commonsourceibias.n608 commonsourceibias.t84 168.701
R21237 commonsourceibias.n601 commonsourceibias.t130 168.701
R21238 commonsourceibias.n599 commonsourceibias.t147 168.701
R21239 commonsourceibias.n593 commonsourceibias.t80 168.701
R21240 commonsourceibias.n586 commonsourceibias.t89 168.701
R21241 commonsourceibias.n584 commonsourceibias.t114 168.701
R21242 commonsourceibias.n578 commonsourceibias.t155 168.701
R21243 commonsourceibias.n571 commonsourceibias.t85 168.701
R21244 commonsourceibias.n528 commonsourceibias.t103 168.701
R21245 commonsourceibias.n534 commonsourceibias.t150 168.701
R21246 commonsourceibias.n540 commonsourceibias.t133 168.701
R21247 commonsourceibias.n542 commonsourceibias.t113 168.701
R21248 commonsourceibias.n549 commonsourceibias.t105 168.701
R21249 commonsourceibias.n555 commonsourceibias.t158 168.701
R21250 commonsourceibias.n519 commonsourceibias.t143 168.701
R21251 commonsourceibias.n517 commonsourceibias.t148 168.701
R21252 commonsourceibias.n515 commonsourceibias.t82 168.701
R21253 commonsourceibias.n363 commonsourceibias.n251 161.3
R21254 commonsourceibias.n361 commonsourceibias.n360 161.3
R21255 commonsourceibias.n359 commonsourceibias.n252 161.3
R21256 commonsourceibias.n358 commonsourceibias.n357 161.3
R21257 commonsourceibias.n355 commonsourceibias.n253 161.3
R21258 commonsourceibias.n354 commonsourceibias.n353 161.3
R21259 commonsourceibias.n352 commonsourceibias.n254 161.3
R21260 commonsourceibias.n351 commonsourceibias.n350 161.3
R21261 commonsourceibias.n349 commonsourceibias.n255 161.3
R21262 commonsourceibias.n347 commonsourceibias.n346 161.3
R21263 commonsourceibias.n345 commonsourceibias.n257 161.3
R21264 commonsourceibias.n344 commonsourceibias.n343 161.3
R21265 commonsourceibias.n341 commonsourceibias.n258 161.3
R21266 commonsourceibias.n340 commonsourceibias.n339 161.3
R21267 commonsourceibias.n338 commonsourceibias.n259 161.3
R21268 commonsourceibias.n337 commonsourceibias.n336 161.3
R21269 commonsourceibias.n335 commonsourceibias.n260 161.3
R21270 commonsourceibias.n333 commonsourceibias.n332 161.3
R21271 commonsourceibias.n331 commonsourceibias.n262 161.3
R21272 commonsourceibias.n330 commonsourceibias.n329 161.3
R21273 commonsourceibias.n327 commonsourceibias.n263 161.3
R21274 commonsourceibias.n326 commonsourceibias.n325 161.3
R21275 commonsourceibias.n324 commonsourceibias.n264 161.3
R21276 commonsourceibias.n323 commonsourceibias.n322 161.3
R21277 commonsourceibias.n321 commonsourceibias.n265 161.3
R21278 commonsourceibias.n319 commonsourceibias.n318 161.3
R21279 commonsourceibias.n317 commonsourceibias.n267 161.3
R21280 commonsourceibias.n316 commonsourceibias.n315 161.3
R21281 commonsourceibias.n313 commonsourceibias.n268 161.3
R21282 commonsourceibias.n312 commonsourceibias.n311 161.3
R21283 commonsourceibias.n310 commonsourceibias.n269 161.3
R21284 commonsourceibias.n309 commonsourceibias.n308 161.3
R21285 commonsourceibias.n307 commonsourceibias.n270 161.3
R21286 commonsourceibias.n305 commonsourceibias.n304 161.3
R21287 commonsourceibias.n303 commonsourceibias.n272 161.3
R21288 commonsourceibias.n302 commonsourceibias.n301 161.3
R21289 commonsourceibias.n299 commonsourceibias.n273 161.3
R21290 commonsourceibias.n298 commonsourceibias.n297 161.3
R21291 commonsourceibias.n296 commonsourceibias.n274 161.3
R21292 commonsourceibias.n295 commonsourceibias.n294 161.3
R21293 commonsourceibias.n293 commonsourceibias.n275 161.3
R21294 commonsourceibias.n291 commonsourceibias.n290 161.3
R21295 commonsourceibias.n289 commonsourceibias.n277 161.3
R21296 commonsourceibias.n288 commonsourceibias.n287 161.3
R21297 commonsourceibias.n285 commonsourceibias.n278 161.3
R21298 commonsourceibias.n284 commonsourceibias.n283 161.3
R21299 commonsourceibias.n282 commonsourceibias.n279 161.3
R21300 commonsourceibias.n45 commonsourceibias.n42 161.3
R21301 commonsourceibias.n47 commonsourceibias.n46 161.3
R21302 commonsourceibias.n48 commonsourceibias.n41 161.3
R21303 commonsourceibias.n51 commonsourceibias.n50 161.3
R21304 commonsourceibias.n52 commonsourceibias.n40 161.3
R21305 commonsourceibias.n54 commonsourceibias.n53 161.3
R21306 commonsourceibias.n56 commonsourceibias.n38 161.3
R21307 commonsourceibias.n58 commonsourceibias.n57 161.3
R21308 commonsourceibias.n59 commonsourceibias.n37 161.3
R21309 commonsourceibias.n61 commonsourceibias.n60 161.3
R21310 commonsourceibias.n62 commonsourceibias.n36 161.3
R21311 commonsourceibias.n65 commonsourceibias.n64 161.3
R21312 commonsourceibias.n66 commonsourceibias.n35 161.3
R21313 commonsourceibias.n68 commonsourceibias.n67 161.3
R21314 commonsourceibias.n70 commonsourceibias.n33 161.3
R21315 commonsourceibias.n72 commonsourceibias.n71 161.3
R21316 commonsourceibias.n73 commonsourceibias.n32 161.3
R21317 commonsourceibias.n75 commonsourceibias.n74 161.3
R21318 commonsourceibias.n76 commonsourceibias.n31 161.3
R21319 commonsourceibias.n79 commonsourceibias.n78 161.3
R21320 commonsourceibias.n80 commonsourceibias.n30 161.3
R21321 commonsourceibias.n82 commonsourceibias.n81 161.3
R21322 commonsourceibias.n84 commonsourceibias.n28 161.3
R21323 commonsourceibias.n86 commonsourceibias.n85 161.3
R21324 commonsourceibias.n87 commonsourceibias.n27 161.3
R21325 commonsourceibias.n89 commonsourceibias.n88 161.3
R21326 commonsourceibias.n90 commonsourceibias.n26 161.3
R21327 commonsourceibias.n93 commonsourceibias.n92 161.3
R21328 commonsourceibias.n94 commonsourceibias.n25 161.3
R21329 commonsourceibias.n96 commonsourceibias.n95 161.3
R21330 commonsourceibias.n98 commonsourceibias.n23 161.3
R21331 commonsourceibias.n100 commonsourceibias.n99 161.3
R21332 commonsourceibias.n101 commonsourceibias.n22 161.3
R21333 commonsourceibias.n103 commonsourceibias.n102 161.3
R21334 commonsourceibias.n104 commonsourceibias.n21 161.3
R21335 commonsourceibias.n107 commonsourceibias.n106 161.3
R21336 commonsourceibias.n108 commonsourceibias.n20 161.3
R21337 commonsourceibias.n110 commonsourceibias.n109 161.3
R21338 commonsourceibias.n112 commonsourceibias.n18 161.3
R21339 commonsourceibias.n114 commonsourceibias.n113 161.3
R21340 commonsourceibias.n115 commonsourceibias.n17 161.3
R21341 commonsourceibias.n117 commonsourceibias.n116 161.3
R21342 commonsourceibias.n118 commonsourceibias.n16 161.3
R21343 commonsourceibias.n121 commonsourceibias.n120 161.3
R21344 commonsourceibias.n122 commonsourceibias.n15 161.3
R21345 commonsourceibias.n124 commonsourceibias.n123 161.3
R21346 commonsourceibias.n126 commonsourceibias.n14 161.3
R21347 commonsourceibias.n167 commonsourceibias.n164 161.3
R21348 commonsourceibias.n169 commonsourceibias.n168 161.3
R21349 commonsourceibias.n170 commonsourceibias.n163 161.3
R21350 commonsourceibias.n173 commonsourceibias.n172 161.3
R21351 commonsourceibias.n174 commonsourceibias.n162 161.3
R21352 commonsourceibias.n176 commonsourceibias.n175 161.3
R21353 commonsourceibias.n178 commonsourceibias.n160 161.3
R21354 commonsourceibias.n180 commonsourceibias.n179 161.3
R21355 commonsourceibias.n181 commonsourceibias.n159 161.3
R21356 commonsourceibias.n183 commonsourceibias.n182 161.3
R21357 commonsourceibias.n184 commonsourceibias.n158 161.3
R21358 commonsourceibias.n187 commonsourceibias.n186 161.3
R21359 commonsourceibias.n188 commonsourceibias.n157 161.3
R21360 commonsourceibias.n190 commonsourceibias.n189 161.3
R21361 commonsourceibias.n192 commonsourceibias.n156 161.3
R21362 commonsourceibias.n194 commonsourceibias.n193 161.3
R21363 commonsourceibias.n196 commonsourceibias.n195 161.3
R21364 commonsourceibias.n197 commonsourceibias.n154 161.3
R21365 commonsourceibias.n199 commonsourceibias.n198 161.3
R21366 commonsourceibias.n201 commonsourceibias.n200 161.3
R21367 commonsourceibias.n202 commonsourceibias.n152 161.3
R21368 commonsourceibias.n204 commonsourceibias.n203 161.3
R21369 commonsourceibias.n206 commonsourceibias.n205 161.3
R21370 commonsourceibias.n208 commonsourceibias.n207 161.3
R21371 commonsourceibias.n209 commonsourceibias.n13 161.3
R21372 commonsourceibias.n211 commonsourceibias.n210 161.3
R21373 commonsourceibias.n212 commonsourceibias.n12 161.3
R21374 commonsourceibias.n215 commonsourceibias.n214 161.3
R21375 commonsourceibias.n216 commonsourceibias.n11 161.3
R21376 commonsourceibias.n218 commonsourceibias.n217 161.3
R21377 commonsourceibias.n220 commonsourceibias.n9 161.3
R21378 commonsourceibias.n222 commonsourceibias.n221 161.3
R21379 commonsourceibias.n223 commonsourceibias.n8 161.3
R21380 commonsourceibias.n225 commonsourceibias.n224 161.3
R21381 commonsourceibias.n226 commonsourceibias.n7 161.3
R21382 commonsourceibias.n229 commonsourceibias.n228 161.3
R21383 commonsourceibias.n230 commonsourceibias.n6 161.3
R21384 commonsourceibias.n232 commonsourceibias.n231 161.3
R21385 commonsourceibias.n234 commonsourceibias.n4 161.3
R21386 commonsourceibias.n236 commonsourceibias.n235 161.3
R21387 commonsourceibias.n237 commonsourceibias.n3 161.3
R21388 commonsourceibias.n239 commonsourceibias.n238 161.3
R21389 commonsourceibias.n240 commonsourceibias.n2 161.3
R21390 commonsourceibias.n243 commonsourceibias.n242 161.3
R21391 commonsourceibias.n244 commonsourceibias.n1 161.3
R21392 commonsourceibias.n246 commonsourceibias.n245 161.3
R21393 commonsourceibias.n248 commonsourceibias.n0 161.3
R21394 commonsourceibias.n730 commonsourceibias.n618 161.3
R21395 commonsourceibias.n728 commonsourceibias.n727 161.3
R21396 commonsourceibias.n726 commonsourceibias.n619 161.3
R21397 commonsourceibias.n725 commonsourceibias.n724 161.3
R21398 commonsourceibias.n722 commonsourceibias.n620 161.3
R21399 commonsourceibias.n721 commonsourceibias.n720 161.3
R21400 commonsourceibias.n719 commonsourceibias.n621 161.3
R21401 commonsourceibias.n718 commonsourceibias.n717 161.3
R21402 commonsourceibias.n715 commonsourceibias.n622 161.3
R21403 commonsourceibias.n713 commonsourceibias.n712 161.3
R21404 commonsourceibias.n711 commonsourceibias.n623 161.3
R21405 commonsourceibias.n710 commonsourceibias.n709 161.3
R21406 commonsourceibias.n707 commonsourceibias.n624 161.3
R21407 commonsourceibias.n706 commonsourceibias.n705 161.3
R21408 commonsourceibias.n704 commonsourceibias.n625 161.3
R21409 commonsourceibias.n703 commonsourceibias.n702 161.3
R21410 commonsourceibias.n700 commonsourceibias.n626 161.3
R21411 commonsourceibias.n698 commonsourceibias.n697 161.3
R21412 commonsourceibias.n696 commonsourceibias.n627 161.3
R21413 commonsourceibias.n695 commonsourceibias.n694 161.3
R21414 commonsourceibias.n692 commonsourceibias.n628 161.3
R21415 commonsourceibias.n691 commonsourceibias.n690 161.3
R21416 commonsourceibias.n689 commonsourceibias.n629 161.3
R21417 commonsourceibias.n688 commonsourceibias.n687 161.3
R21418 commonsourceibias.n685 commonsourceibias.n630 161.3
R21419 commonsourceibias.n683 commonsourceibias.n682 161.3
R21420 commonsourceibias.n681 commonsourceibias.n631 161.3
R21421 commonsourceibias.n680 commonsourceibias.n679 161.3
R21422 commonsourceibias.n677 commonsourceibias.n632 161.3
R21423 commonsourceibias.n676 commonsourceibias.n675 161.3
R21424 commonsourceibias.n674 commonsourceibias.n633 161.3
R21425 commonsourceibias.n673 commonsourceibias.n672 161.3
R21426 commonsourceibias.n670 commonsourceibias.n634 161.3
R21427 commonsourceibias.n668 commonsourceibias.n667 161.3
R21428 commonsourceibias.n666 commonsourceibias.n635 161.3
R21429 commonsourceibias.n665 commonsourceibias.n664 161.3
R21430 commonsourceibias.n662 commonsourceibias.n636 161.3
R21431 commonsourceibias.n661 commonsourceibias.n660 161.3
R21432 commonsourceibias.n659 commonsourceibias.n637 161.3
R21433 commonsourceibias.n658 commonsourceibias.n657 161.3
R21434 commonsourceibias.n655 commonsourceibias.n638 161.3
R21435 commonsourceibias.n653 commonsourceibias.n652 161.3
R21436 commonsourceibias.n651 commonsourceibias.n639 161.3
R21437 commonsourceibias.n650 commonsourceibias.n649 161.3
R21438 commonsourceibias.n647 commonsourceibias.n640 161.3
R21439 commonsourceibias.n646 commonsourceibias.n645 161.3
R21440 commonsourceibias.n644 commonsourceibias.n641 161.3
R21441 commonsourceibias.n500 commonsourceibias.n388 161.3
R21442 commonsourceibias.n498 commonsourceibias.n497 161.3
R21443 commonsourceibias.n496 commonsourceibias.n389 161.3
R21444 commonsourceibias.n495 commonsourceibias.n494 161.3
R21445 commonsourceibias.n492 commonsourceibias.n390 161.3
R21446 commonsourceibias.n491 commonsourceibias.n490 161.3
R21447 commonsourceibias.n489 commonsourceibias.n391 161.3
R21448 commonsourceibias.n488 commonsourceibias.n487 161.3
R21449 commonsourceibias.n485 commonsourceibias.n392 161.3
R21450 commonsourceibias.n483 commonsourceibias.n482 161.3
R21451 commonsourceibias.n481 commonsourceibias.n393 161.3
R21452 commonsourceibias.n480 commonsourceibias.n479 161.3
R21453 commonsourceibias.n477 commonsourceibias.n394 161.3
R21454 commonsourceibias.n476 commonsourceibias.n475 161.3
R21455 commonsourceibias.n474 commonsourceibias.n395 161.3
R21456 commonsourceibias.n473 commonsourceibias.n472 161.3
R21457 commonsourceibias.n470 commonsourceibias.n396 161.3
R21458 commonsourceibias.n468 commonsourceibias.n467 161.3
R21459 commonsourceibias.n466 commonsourceibias.n397 161.3
R21460 commonsourceibias.n465 commonsourceibias.n464 161.3
R21461 commonsourceibias.n462 commonsourceibias.n398 161.3
R21462 commonsourceibias.n461 commonsourceibias.n460 161.3
R21463 commonsourceibias.n459 commonsourceibias.n399 161.3
R21464 commonsourceibias.n458 commonsourceibias.n457 161.3
R21465 commonsourceibias.n455 commonsourceibias.n400 161.3
R21466 commonsourceibias.n453 commonsourceibias.n452 161.3
R21467 commonsourceibias.n451 commonsourceibias.n401 161.3
R21468 commonsourceibias.n450 commonsourceibias.n449 161.3
R21469 commonsourceibias.n447 commonsourceibias.n402 161.3
R21470 commonsourceibias.n446 commonsourceibias.n445 161.3
R21471 commonsourceibias.n444 commonsourceibias.n403 161.3
R21472 commonsourceibias.n443 commonsourceibias.n442 161.3
R21473 commonsourceibias.n440 commonsourceibias.n404 161.3
R21474 commonsourceibias.n438 commonsourceibias.n437 161.3
R21475 commonsourceibias.n436 commonsourceibias.n405 161.3
R21476 commonsourceibias.n435 commonsourceibias.n434 161.3
R21477 commonsourceibias.n432 commonsourceibias.n406 161.3
R21478 commonsourceibias.n431 commonsourceibias.n430 161.3
R21479 commonsourceibias.n429 commonsourceibias.n407 161.3
R21480 commonsourceibias.n428 commonsourceibias.n427 161.3
R21481 commonsourceibias.n425 commonsourceibias.n408 161.3
R21482 commonsourceibias.n423 commonsourceibias.n422 161.3
R21483 commonsourceibias.n421 commonsourceibias.n409 161.3
R21484 commonsourceibias.n420 commonsourceibias.n419 161.3
R21485 commonsourceibias.n417 commonsourceibias.n410 161.3
R21486 commonsourceibias.n416 commonsourceibias.n415 161.3
R21487 commonsourceibias.n414 commonsourceibias.n411 161.3
R21488 commonsourceibias.n570 commonsourceibias.n569 161.3
R21489 commonsourceibias.n568 commonsourceibias.n567 161.3
R21490 commonsourceibias.n566 commonsourceibias.n516 161.3
R21491 commonsourceibias.n565 commonsourceibias.n564 161.3
R21492 commonsourceibias.n563 commonsourceibias.n562 161.3
R21493 commonsourceibias.n561 commonsourceibias.n518 161.3
R21494 commonsourceibias.n560 commonsourceibias.n559 161.3
R21495 commonsourceibias.n558 commonsourceibias.n557 161.3
R21496 commonsourceibias.n556 commonsourceibias.n520 161.3
R21497 commonsourceibias.n554 commonsourceibias.n553 161.3
R21498 commonsourceibias.n552 commonsourceibias.n521 161.3
R21499 commonsourceibias.n551 commonsourceibias.n550 161.3
R21500 commonsourceibias.n548 commonsourceibias.n522 161.3
R21501 commonsourceibias.n547 commonsourceibias.n546 161.3
R21502 commonsourceibias.n545 commonsourceibias.n523 161.3
R21503 commonsourceibias.n544 commonsourceibias.n543 161.3
R21504 commonsourceibias.n541 commonsourceibias.n524 161.3
R21505 commonsourceibias.n539 commonsourceibias.n538 161.3
R21506 commonsourceibias.n537 commonsourceibias.n525 161.3
R21507 commonsourceibias.n536 commonsourceibias.n535 161.3
R21508 commonsourceibias.n533 commonsourceibias.n526 161.3
R21509 commonsourceibias.n532 commonsourceibias.n531 161.3
R21510 commonsourceibias.n530 commonsourceibias.n527 161.3
R21511 commonsourceibias.n615 commonsourceibias.n367 161.3
R21512 commonsourceibias.n613 commonsourceibias.n612 161.3
R21513 commonsourceibias.n611 commonsourceibias.n368 161.3
R21514 commonsourceibias.n610 commonsourceibias.n609 161.3
R21515 commonsourceibias.n607 commonsourceibias.n369 161.3
R21516 commonsourceibias.n606 commonsourceibias.n605 161.3
R21517 commonsourceibias.n604 commonsourceibias.n370 161.3
R21518 commonsourceibias.n603 commonsourceibias.n602 161.3
R21519 commonsourceibias.n600 commonsourceibias.n371 161.3
R21520 commonsourceibias.n598 commonsourceibias.n597 161.3
R21521 commonsourceibias.n596 commonsourceibias.n372 161.3
R21522 commonsourceibias.n595 commonsourceibias.n594 161.3
R21523 commonsourceibias.n592 commonsourceibias.n373 161.3
R21524 commonsourceibias.n591 commonsourceibias.n590 161.3
R21525 commonsourceibias.n589 commonsourceibias.n374 161.3
R21526 commonsourceibias.n588 commonsourceibias.n587 161.3
R21527 commonsourceibias.n585 commonsourceibias.n375 161.3
R21528 commonsourceibias.n583 commonsourceibias.n582 161.3
R21529 commonsourceibias.n581 commonsourceibias.n376 161.3
R21530 commonsourceibias.n580 commonsourceibias.n579 161.3
R21531 commonsourceibias.n577 commonsourceibias.n377 161.3
R21532 commonsourceibias.n576 commonsourceibias.n575 161.3
R21533 commonsourceibias.n574 commonsourceibias.n378 161.3
R21534 commonsourceibias.n573 commonsourceibias.n572 161.3
R21535 commonsourceibias.n141 commonsourceibias.n139 81.5057
R21536 commonsourceibias.n381 commonsourceibias.n379 81.5057
R21537 commonsourceibias.n141 commonsourceibias.n140 80.9324
R21538 commonsourceibias.n143 commonsourceibias.n142 80.9324
R21539 commonsourceibias.n145 commonsourceibias.n144 80.9324
R21540 commonsourceibias.n147 commonsourceibias.n146 80.9324
R21541 commonsourceibias.n138 commonsourceibias.n137 80.9324
R21542 commonsourceibias.n136 commonsourceibias.n135 80.9324
R21543 commonsourceibias.n134 commonsourceibias.n133 80.9324
R21544 commonsourceibias.n132 commonsourceibias.n131 80.9324
R21545 commonsourceibias.n130 commonsourceibias.n129 80.9324
R21546 commonsourceibias.n504 commonsourceibias.n503 80.9324
R21547 commonsourceibias.n506 commonsourceibias.n505 80.9324
R21548 commonsourceibias.n508 commonsourceibias.n507 80.9324
R21549 commonsourceibias.n510 commonsourceibias.n509 80.9324
R21550 commonsourceibias.n512 commonsourceibias.n511 80.9324
R21551 commonsourceibias.n387 commonsourceibias.n386 80.9324
R21552 commonsourceibias.n385 commonsourceibias.n384 80.9324
R21553 commonsourceibias.n383 commonsourceibias.n382 80.9324
R21554 commonsourceibias.n381 commonsourceibias.n380 80.9324
R21555 commonsourceibias.n365 commonsourceibias.n364 80.6037
R21556 commonsourceibias.n128 commonsourceibias.n127 80.6037
R21557 commonsourceibias.n250 commonsourceibias.n249 80.6037
R21558 commonsourceibias.n732 commonsourceibias.n731 80.6037
R21559 commonsourceibias.n502 commonsourceibias.n501 80.6037
R21560 commonsourceibias.n617 commonsourceibias.n616 80.6037
R21561 commonsourceibias.n322 commonsourceibias.n321 56.5617
R21562 commonsourceibias.n336 commonsourceibias.n335 56.5617
R21563 commonsourceibias.n85 commonsourceibias.n84 56.5617
R21564 commonsourceibias.n71 commonsourceibias.n70 56.5617
R21565 commonsourceibias.n207 commonsourceibias.n206 56.5617
R21566 commonsourceibias.n193 commonsourceibias.n192 56.5617
R21567 commonsourceibias.n687 commonsourceibias.n685 56.5617
R21568 commonsourceibias.n702 commonsourceibias.n700 56.5617
R21569 commonsourceibias.n457 commonsourceibias.n455 56.5617
R21570 commonsourceibias.n472 commonsourceibias.n470 56.5617
R21571 commonsourceibias.n572 commonsourceibias.n570 56.5617
R21572 commonsourceibias.n294 commonsourceibias.n293 56.5617
R21573 commonsourceibias.n308 commonsourceibias.n307 56.5617
R21574 commonsourceibias.n350 commonsourceibias.n349 56.5617
R21575 commonsourceibias.n113 commonsourceibias.n112 56.5617
R21576 commonsourceibias.n99 commonsourceibias.n98 56.5617
R21577 commonsourceibias.n57 commonsourceibias.n56 56.5617
R21578 commonsourceibias.n235 commonsourceibias.n234 56.5617
R21579 commonsourceibias.n221 commonsourceibias.n220 56.5617
R21580 commonsourceibias.n179 commonsourceibias.n178 56.5617
R21581 commonsourceibias.n657 commonsourceibias.n655 56.5617
R21582 commonsourceibias.n672 commonsourceibias.n670 56.5617
R21583 commonsourceibias.n717 commonsourceibias.n715 56.5617
R21584 commonsourceibias.n427 commonsourceibias.n425 56.5617
R21585 commonsourceibias.n442 commonsourceibias.n440 56.5617
R21586 commonsourceibias.n487 commonsourceibias.n485 56.5617
R21587 commonsourceibias.n602 commonsourceibias.n600 56.5617
R21588 commonsourceibias.n587 commonsourceibias.n585 56.5617
R21589 commonsourceibias.n543 commonsourceibias.n541 56.5617
R21590 commonsourceibias.n557 commonsourceibias.n556 56.5617
R21591 commonsourceibias.n285 commonsourceibias.n284 51.2335
R21592 commonsourceibias.n357 commonsourceibias.n252 51.2335
R21593 commonsourceibias.n120 commonsourceibias.n15 51.2335
R21594 commonsourceibias.n48 commonsourceibias.n47 51.2335
R21595 commonsourceibias.n242 commonsourceibias.n1 51.2335
R21596 commonsourceibias.n170 commonsourceibias.n169 51.2335
R21597 commonsourceibias.n647 commonsourceibias.n646 51.2335
R21598 commonsourceibias.n724 commonsourceibias.n619 51.2335
R21599 commonsourceibias.n417 commonsourceibias.n416 51.2335
R21600 commonsourceibias.n494 commonsourceibias.n389 51.2335
R21601 commonsourceibias.n609 commonsourceibias.n368 51.2335
R21602 commonsourceibias.n533 commonsourceibias.n532 51.2335
R21603 commonsourceibias.n364 commonsourceibias.n363 50.9056
R21604 commonsourceibias.n127 commonsourceibias.n126 50.9056
R21605 commonsourceibias.n249 commonsourceibias.n248 50.9056
R21606 commonsourceibias.n731 commonsourceibias.n730 50.9056
R21607 commonsourceibias.n501 commonsourceibias.n500 50.9056
R21608 commonsourceibias.n616 commonsourceibias.n615 50.9056
R21609 commonsourceibias.n299 commonsourceibias.n298 50.2647
R21610 commonsourceibias.n343 commonsourceibias.n257 50.2647
R21611 commonsourceibias.n106 commonsourceibias.n20 50.2647
R21612 commonsourceibias.n62 commonsourceibias.n61 50.2647
R21613 commonsourceibias.n228 commonsourceibias.n6 50.2647
R21614 commonsourceibias.n184 commonsourceibias.n183 50.2647
R21615 commonsourceibias.n662 commonsourceibias.n661 50.2647
R21616 commonsourceibias.n709 commonsourceibias.n623 50.2647
R21617 commonsourceibias.n432 commonsourceibias.n431 50.2647
R21618 commonsourceibias.n479 commonsourceibias.n393 50.2647
R21619 commonsourceibias.n594 commonsourceibias.n372 50.2647
R21620 commonsourceibias.n548 commonsourceibias.n547 50.2647
R21621 commonsourceibias.n281 commonsourceibias.n280 49.9027
R21622 commonsourceibias.n44 commonsourceibias.n43 49.9027
R21623 commonsourceibias.n166 commonsourceibias.n165 49.9027
R21624 commonsourceibias.n643 commonsourceibias.n642 49.9027
R21625 commonsourceibias.n413 commonsourceibias.n412 49.9027
R21626 commonsourceibias.n529 commonsourceibias.n528 49.9027
R21627 commonsourceibias.n313 commonsourceibias.n312 49.296
R21628 commonsourceibias.n329 commonsourceibias.n262 49.296
R21629 commonsourceibias.n92 commonsourceibias.n25 49.296
R21630 commonsourceibias.n76 commonsourceibias.n75 49.296
R21631 commonsourceibias.n214 commonsourceibias.n11 49.296
R21632 commonsourceibias.n198 commonsourceibias.n197 49.296
R21633 commonsourceibias.n677 commonsourceibias.n676 49.296
R21634 commonsourceibias.n694 commonsourceibias.n627 49.296
R21635 commonsourceibias.n447 commonsourceibias.n446 49.296
R21636 commonsourceibias.n464 commonsourceibias.n397 49.296
R21637 commonsourceibias.n579 commonsourceibias.n376 49.296
R21638 commonsourceibias.n562 commonsourceibias.n561 49.296
R21639 commonsourceibias.n315 commonsourceibias.n267 48.3272
R21640 commonsourceibias.n327 commonsourceibias.n326 48.3272
R21641 commonsourceibias.n90 commonsourceibias.n89 48.3272
R21642 commonsourceibias.n78 commonsourceibias.n30 48.3272
R21643 commonsourceibias.n212 commonsourceibias.n211 48.3272
R21644 commonsourceibias.n202 commonsourceibias.n201 48.3272
R21645 commonsourceibias.n679 commonsourceibias.n631 48.3272
R21646 commonsourceibias.n692 commonsourceibias.n691 48.3272
R21647 commonsourceibias.n449 commonsourceibias.n401 48.3272
R21648 commonsourceibias.n462 commonsourceibias.n461 48.3272
R21649 commonsourceibias.n577 commonsourceibias.n576 48.3272
R21650 commonsourceibias.n566 commonsourceibias.n565 48.3272
R21651 commonsourceibias.n301 commonsourceibias.n272 47.3584
R21652 commonsourceibias.n341 commonsourceibias.n340 47.3584
R21653 commonsourceibias.n104 commonsourceibias.n103 47.3584
R21654 commonsourceibias.n64 commonsourceibias.n35 47.3584
R21655 commonsourceibias.n226 commonsourceibias.n225 47.3584
R21656 commonsourceibias.n186 commonsourceibias.n157 47.3584
R21657 commonsourceibias.n664 commonsourceibias.n635 47.3584
R21658 commonsourceibias.n707 commonsourceibias.n706 47.3584
R21659 commonsourceibias.n434 commonsourceibias.n405 47.3584
R21660 commonsourceibias.n477 commonsourceibias.n476 47.3584
R21661 commonsourceibias.n592 commonsourceibias.n591 47.3584
R21662 commonsourceibias.n550 commonsourceibias.n521 47.3584
R21663 commonsourceibias.n287 commonsourceibias.n277 46.3896
R21664 commonsourceibias.n355 commonsourceibias.n354 46.3896
R21665 commonsourceibias.n118 commonsourceibias.n117 46.3896
R21666 commonsourceibias.n50 commonsourceibias.n40 46.3896
R21667 commonsourceibias.n240 commonsourceibias.n239 46.3896
R21668 commonsourceibias.n172 commonsourceibias.n162 46.3896
R21669 commonsourceibias.n649 commonsourceibias.n639 46.3896
R21670 commonsourceibias.n722 commonsourceibias.n721 46.3896
R21671 commonsourceibias.n419 commonsourceibias.n409 46.3896
R21672 commonsourceibias.n492 commonsourceibias.n491 46.3896
R21673 commonsourceibias.n607 commonsourceibias.n606 46.3896
R21674 commonsourceibias.n535 commonsourceibias.n525 46.3896
R21675 commonsourceibias.n282 commonsourceibias.n281 44.7059
R21676 commonsourceibias.n644 commonsourceibias.n643 44.7059
R21677 commonsourceibias.n414 commonsourceibias.n413 44.7059
R21678 commonsourceibias.n530 commonsourceibias.n529 44.7059
R21679 commonsourceibias.n45 commonsourceibias.n44 44.7059
R21680 commonsourceibias.n167 commonsourceibias.n166 44.7059
R21681 commonsourceibias.n291 commonsourceibias.n277 34.7644
R21682 commonsourceibias.n354 commonsourceibias.n254 34.7644
R21683 commonsourceibias.n117 commonsourceibias.n17 34.7644
R21684 commonsourceibias.n54 commonsourceibias.n40 34.7644
R21685 commonsourceibias.n239 commonsourceibias.n3 34.7644
R21686 commonsourceibias.n176 commonsourceibias.n162 34.7644
R21687 commonsourceibias.n653 commonsourceibias.n639 34.7644
R21688 commonsourceibias.n721 commonsourceibias.n621 34.7644
R21689 commonsourceibias.n423 commonsourceibias.n409 34.7644
R21690 commonsourceibias.n491 commonsourceibias.n391 34.7644
R21691 commonsourceibias.n606 commonsourceibias.n370 34.7644
R21692 commonsourceibias.n539 commonsourceibias.n525 34.7644
R21693 commonsourceibias.n305 commonsourceibias.n272 33.7956
R21694 commonsourceibias.n340 commonsourceibias.n259 33.7956
R21695 commonsourceibias.n103 commonsourceibias.n22 33.7956
R21696 commonsourceibias.n68 commonsourceibias.n35 33.7956
R21697 commonsourceibias.n225 commonsourceibias.n8 33.7956
R21698 commonsourceibias.n190 commonsourceibias.n157 33.7956
R21699 commonsourceibias.n668 commonsourceibias.n635 33.7956
R21700 commonsourceibias.n706 commonsourceibias.n625 33.7956
R21701 commonsourceibias.n438 commonsourceibias.n405 33.7956
R21702 commonsourceibias.n476 commonsourceibias.n395 33.7956
R21703 commonsourceibias.n591 commonsourceibias.n374 33.7956
R21704 commonsourceibias.n554 commonsourceibias.n521 33.7956
R21705 commonsourceibias.n319 commonsourceibias.n267 32.8269
R21706 commonsourceibias.n326 commonsourceibias.n264 32.8269
R21707 commonsourceibias.n89 commonsourceibias.n27 32.8269
R21708 commonsourceibias.n82 commonsourceibias.n30 32.8269
R21709 commonsourceibias.n211 commonsourceibias.n13 32.8269
R21710 commonsourceibias.n203 commonsourceibias.n202 32.8269
R21711 commonsourceibias.n683 commonsourceibias.n631 32.8269
R21712 commonsourceibias.n691 commonsourceibias.n629 32.8269
R21713 commonsourceibias.n453 commonsourceibias.n401 32.8269
R21714 commonsourceibias.n461 commonsourceibias.n399 32.8269
R21715 commonsourceibias.n576 commonsourceibias.n378 32.8269
R21716 commonsourceibias.n567 commonsourceibias.n566 32.8269
R21717 commonsourceibias.n312 commonsourceibias.n269 31.8581
R21718 commonsourceibias.n333 commonsourceibias.n262 31.8581
R21719 commonsourceibias.n96 commonsourceibias.n25 31.8581
R21720 commonsourceibias.n75 commonsourceibias.n32 31.8581
R21721 commonsourceibias.n218 commonsourceibias.n11 31.8581
R21722 commonsourceibias.n197 commonsourceibias.n196 31.8581
R21723 commonsourceibias.n676 commonsourceibias.n633 31.8581
R21724 commonsourceibias.n698 commonsourceibias.n627 31.8581
R21725 commonsourceibias.n446 commonsourceibias.n403 31.8581
R21726 commonsourceibias.n468 commonsourceibias.n397 31.8581
R21727 commonsourceibias.n583 commonsourceibias.n376 31.8581
R21728 commonsourceibias.n561 commonsourceibias.n560 31.8581
R21729 commonsourceibias.n298 commonsourceibias.n274 30.8893
R21730 commonsourceibias.n347 commonsourceibias.n257 30.8893
R21731 commonsourceibias.n110 commonsourceibias.n20 30.8893
R21732 commonsourceibias.n61 commonsourceibias.n37 30.8893
R21733 commonsourceibias.n232 commonsourceibias.n6 30.8893
R21734 commonsourceibias.n183 commonsourceibias.n159 30.8893
R21735 commonsourceibias.n661 commonsourceibias.n637 30.8893
R21736 commonsourceibias.n713 commonsourceibias.n623 30.8893
R21737 commonsourceibias.n431 commonsourceibias.n407 30.8893
R21738 commonsourceibias.n483 commonsourceibias.n393 30.8893
R21739 commonsourceibias.n598 commonsourceibias.n372 30.8893
R21740 commonsourceibias.n547 commonsourceibias.n523 30.8893
R21741 commonsourceibias.n284 commonsourceibias.n279 29.9206
R21742 commonsourceibias.n361 commonsourceibias.n252 29.9206
R21743 commonsourceibias.n124 commonsourceibias.n15 29.9206
R21744 commonsourceibias.n47 commonsourceibias.n42 29.9206
R21745 commonsourceibias.n246 commonsourceibias.n1 29.9206
R21746 commonsourceibias.n169 commonsourceibias.n164 29.9206
R21747 commonsourceibias.n646 commonsourceibias.n641 29.9206
R21748 commonsourceibias.n728 commonsourceibias.n619 29.9206
R21749 commonsourceibias.n416 commonsourceibias.n411 29.9206
R21750 commonsourceibias.n498 commonsourceibias.n389 29.9206
R21751 commonsourceibias.n613 commonsourceibias.n368 29.9206
R21752 commonsourceibias.n532 commonsourceibias.n527 29.9206
R21753 commonsourceibias.n363 commonsourceibias.n362 21.8872
R21754 commonsourceibias.n126 commonsourceibias.n125 21.8872
R21755 commonsourceibias.n248 commonsourceibias.n247 21.8872
R21756 commonsourceibias.n730 commonsourceibias.n729 21.8872
R21757 commonsourceibias.n500 commonsourceibias.n499 21.8872
R21758 commonsourceibias.n615 commonsourceibias.n614 21.8872
R21759 commonsourceibias.n294 commonsourceibias.n276 21.3954
R21760 commonsourceibias.n349 commonsourceibias.n348 21.3954
R21761 commonsourceibias.n112 commonsourceibias.n111 21.3954
R21762 commonsourceibias.n57 commonsourceibias.n39 21.3954
R21763 commonsourceibias.n234 commonsourceibias.n233 21.3954
R21764 commonsourceibias.n179 commonsourceibias.n161 21.3954
R21765 commonsourceibias.n657 commonsourceibias.n656 21.3954
R21766 commonsourceibias.n715 commonsourceibias.n714 21.3954
R21767 commonsourceibias.n427 commonsourceibias.n426 21.3954
R21768 commonsourceibias.n485 commonsourceibias.n484 21.3954
R21769 commonsourceibias.n600 commonsourceibias.n599 21.3954
R21770 commonsourceibias.n543 commonsourceibias.n542 21.3954
R21771 commonsourceibias.n308 commonsourceibias.n271 20.9036
R21772 commonsourceibias.n335 commonsourceibias.n334 20.9036
R21773 commonsourceibias.n98 commonsourceibias.n97 20.9036
R21774 commonsourceibias.n71 commonsourceibias.n34 20.9036
R21775 commonsourceibias.n220 commonsourceibias.n219 20.9036
R21776 commonsourceibias.n193 commonsourceibias.n155 20.9036
R21777 commonsourceibias.n672 commonsourceibias.n671 20.9036
R21778 commonsourceibias.n700 commonsourceibias.n699 20.9036
R21779 commonsourceibias.n442 commonsourceibias.n441 20.9036
R21780 commonsourceibias.n470 commonsourceibias.n469 20.9036
R21781 commonsourceibias.n585 commonsourceibias.n584 20.9036
R21782 commonsourceibias.n557 commonsourceibias.n519 20.9036
R21783 commonsourceibias.n321 commonsourceibias.n320 20.4117
R21784 commonsourceibias.n322 commonsourceibias.n266 20.4117
R21785 commonsourceibias.n85 commonsourceibias.n29 20.4117
R21786 commonsourceibias.n84 commonsourceibias.n83 20.4117
R21787 commonsourceibias.n207 commonsourceibias.n150 20.4117
R21788 commonsourceibias.n206 commonsourceibias.n151 20.4117
R21789 commonsourceibias.n685 commonsourceibias.n684 20.4117
R21790 commonsourceibias.n687 commonsourceibias.n686 20.4117
R21791 commonsourceibias.n455 commonsourceibias.n454 20.4117
R21792 commonsourceibias.n457 commonsourceibias.n456 20.4117
R21793 commonsourceibias.n572 commonsourceibias.n571 20.4117
R21794 commonsourceibias.n570 commonsourceibias.n515 20.4117
R21795 commonsourceibias.n307 commonsourceibias.n306 19.9199
R21796 commonsourceibias.n336 commonsourceibias.n261 19.9199
R21797 commonsourceibias.n99 commonsourceibias.n24 19.9199
R21798 commonsourceibias.n70 commonsourceibias.n69 19.9199
R21799 commonsourceibias.n221 commonsourceibias.n10 19.9199
R21800 commonsourceibias.n192 commonsourceibias.n191 19.9199
R21801 commonsourceibias.n670 commonsourceibias.n669 19.9199
R21802 commonsourceibias.n702 commonsourceibias.n701 19.9199
R21803 commonsourceibias.n440 commonsourceibias.n439 19.9199
R21804 commonsourceibias.n472 commonsourceibias.n471 19.9199
R21805 commonsourceibias.n587 commonsourceibias.n586 19.9199
R21806 commonsourceibias.n556 commonsourceibias.n555 19.9199
R21807 commonsourceibias.n293 commonsourceibias.n292 19.4281
R21808 commonsourceibias.n350 commonsourceibias.n256 19.4281
R21809 commonsourceibias.n113 commonsourceibias.n19 19.4281
R21810 commonsourceibias.n56 commonsourceibias.n55 19.4281
R21811 commonsourceibias.n235 commonsourceibias.n5 19.4281
R21812 commonsourceibias.n178 commonsourceibias.n177 19.4281
R21813 commonsourceibias.n655 commonsourceibias.n654 19.4281
R21814 commonsourceibias.n717 commonsourceibias.n716 19.4281
R21815 commonsourceibias.n425 commonsourceibias.n424 19.4281
R21816 commonsourceibias.n487 commonsourceibias.n486 19.4281
R21817 commonsourceibias.n602 commonsourceibias.n601 19.4281
R21818 commonsourceibias.n541 commonsourceibias.n540 19.4281
R21819 commonsourceibias.n286 commonsourceibias.n285 13.526
R21820 commonsourceibias.n357 commonsourceibias.n356 13.526
R21821 commonsourceibias.n120 commonsourceibias.n119 13.526
R21822 commonsourceibias.n49 commonsourceibias.n48 13.526
R21823 commonsourceibias.n242 commonsourceibias.n241 13.526
R21824 commonsourceibias.n171 commonsourceibias.n170 13.526
R21825 commonsourceibias.n648 commonsourceibias.n647 13.526
R21826 commonsourceibias.n724 commonsourceibias.n723 13.526
R21827 commonsourceibias.n418 commonsourceibias.n417 13.526
R21828 commonsourceibias.n494 commonsourceibias.n493 13.526
R21829 commonsourceibias.n609 commonsourceibias.n608 13.526
R21830 commonsourceibias.n534 commonsourceibias.n533 13.526
R21831 commonsourceibias.n130 commonsourceibias.n128 13.2322
R21832 commonsourceibias.n504 commonsourceibias.n502 13.2322
R21833 commonsourceibias.n300 commonsourceibias.n299 13.0342
R21834 commonsourceibias.n343 commonsourceibias.n342 13.0342
R21835 commonsourceibias.n106 commonsourceibias.n105 13.0342
R21836 commonsourceibias.n63 commonsourceibias.n62 13.0342
R21837 commonsourceibias.n228 commonsourceibias.n227 13.0342
R21838 commonsourceibias.n185 commonsourceibias.n184 13.0342
R21839 commonsourceibias.n663 commonsourceibias.n662 13.0342
R21840 commonsourceibias.n709 commonsourceibias.n708 13.0342
R21841 commonsourceibias.n433 commonsourceibias.n432 13.0342
R21842 commonsourceibias.n479 commonsourceibias.n478 13.0342
R21843 commonsourceibias.n594 commonsourceibias.n593 13.0342
R21844 commonsourceibias.n549 commonsourceibias.n548 13.0342
R21845 commonsourceibias.n314 commonsourceibias.n313 12.5423
R21846 commonsourceibias.n329 commonsourceibias.n328 12.5423
R21847 commonsourceibias.n92 commonsourceibias.n91 12.5423
R21848 commonsourceibias.n77 commonsourceibias.n76 12.5423
R21849 commonsourceibias.n214 commonsourceibias.n213 12.5423
R21850 commonsourceibias.n198 commonsourceibias.n153 12.5423
R21851 commonsourceibias.n678 commonsourceibias.n677 12.5423
R21852 commonsourceibias.n694 commonsourceibias.n693 12.5423
R21853 commonsourceibias.n448 commonsourceibias.n447 12.5423
R21854 commonsourceibias.n464 commonsourceibias.n463 12.5423
R21855 commonsourceibias.n579 commonsourceibias.n578 12.5423
R21856 commonsourceibias.n562 commonsourceibias.n517 12.5423
R21857 commonsourceibias.n734 commonsourceibias.n366 12.2777
R21858 commonsourceibias.n315 commonsourceibias.n314 12.0505
R21859 commonsourceibias.n328 commonsourceibias.n327 12.0505
R21860 commonsourceibias.n91 commonsourceibias.n90 12.0505
R21861 commonsourceibias.n78 commonsourceibias.n77 12.0505
R21862 commonsourceibias.n213 commonsourceibias.n212 12.0505
R21863 commonsourceibias.n201 commonsourceibias.n153 12.0505
R21864 commonsourceibias.n679 commonsourceibias.n678 12.0505
R21865 commonsourceibias.n693 commonsourceibias.n692 12.0505
R21866 commonsourceibias.n449 commonsourceibias.n448 12.0505
R21867 commonsourceibias.n463 commonsourceibias.n462 12.0505
R21868 commonsourceibias.n578 commonsourceibias.n577 12.0505
R21869 commonsourceibias.n565 commonsourceibias.n517 12.0505
R21870 commonsourceibias.n301 commonsourceibias.n300 11.5587
R21871 commonsourceibias.n342 commonsourceibias.n341 11.5587
R21872 commonsourceibias.n105 commonsourceibias.n104 11.5587
R21873 commonsourceibias.n64 commonsourceibias.n63 11.5587
R21874 commonsourceibias.n227 commonsourceibias.n226 11.5587
R21875 commonsourceibias.n186 commonsourceibias.n185 11.5587
R21876 commonsourceibias.n664 commonsourceibias.n663 11.5587
R21877 commonsourceibias.n708 commonsourceibias.n707 11.5587
R21878 commonsourceibias.n434 commonsourceibias.n433 11.5587
R21879 commonsourceibias.n478 commonsourceibias.n477 11.5587
R21880 commonsourceibias.n593 commonsourceibias.n592 11.5587
R21881 commonsourceibias.n550 commonsourceibias.n549 11.5587
R21882 commonsourceibias.n287 commonsourceibias.n286 11.0668
R21883 commonsourceibias.n356 commonsourceibias.n355 11.0668
R21884 commonsourceibias.n119 commonsourceibias.n118 11.0668
R21885 commonsourceibias.n50 commonsourceibias.n49 11.0668
R21886 commonsourceibias.n241 commonsourceibias.n240 11.0668
R21887 commonsourceibias.n172 commonsourceibias.n171 11.0668
R21888 commonsourceibias.n649 commonsourceibias.n648 11.0668
R21889 commonsourceibias.n723 commonsourceibias.n722 11.0668
R21890 commonsourceibias.n419 commonsourceibias.n418 11.0668
R21891 commonsourceibias.n493 commonsourceibias.n492 11.0668
R21892 commonsourceibias.n608 commonsourceibias.n607 11.0668
R21893 commonsourceibias.n535 commonsourceibias.n534 11.0668
R21894 commonsourceibias.n734 commonsourceibias.n733 10.3347
R21895 commonsourceibias.n149 commonsourceibias.n148 9.50363
R21896 commonsourceibias.n514 commonsourceibias.n513 9.50363
R21897 commonsourceibias.n366 commonsourceibias.n250 8.75852
R21898 commonsourceibias.n733 commonsourceibias.n617 8.75852
R21899 commonsourceibias.n292 commonsourceibias.n291 5.16479
R21900 commonsourceibias.n256 commonsourceibias.n254 5.16479
R21901 commonsourceibias.n19 commonsourceibias.n17 5.16479
R21902 commonsourceibias.n55 commonsourceibias.n54 5.16479
R21903 commonsourceibias.n5 commonsourceibias.n3 5.16479
R21904 commonsourceibias.n177 commonsourceibias.n176 5.16479
R21905 commonsourceibias.n654 commonsourceibias.n653 5.16479
R21906 commonsourceibias.n716 commonsourceibias.n621 5.16479
R21907 commonsourceibias.n424 commonsourceibias.n423 5.16479
R21908 commonsourceibias.n486 commonsourceibias.n391 5.16479
R21909 commonsourceibias.n601 commonsourceibias.n370 5.16479
R21910 commonsourceibias.n540 commonsourceibias.n539 5.16479
R21911 commonsourceibias.n366 commonsourceibias.n365 5.03125
R21912 commonsourceibias.n733 commonsourceibias.n732 5.03125
R21913 commonsourceibias.n306 commonsourceibias.n305 4.67295
R21914 commonsourceibias.n261 commonsourceibias.n259 4.67295
R21915 commonsourceibias.n24 commonsourceibias.n22 4.67295
R21916 commonsourceibias.n69 commonsourceibias.n68 4.67295
R21917 commonsourceibias.n10 commonsourceibias.n8 4.67295
R21918 commonsourceibias.n191 commonsourceibias.n190 4.67295
R21919 commonsourceibias.n669 commonsourceibias.n668 4.67295
R21920 commonsourceibias.n701 commonsourceibias.n625 4.67295
R21921 commonsourceibias.n439 commonsourceibias.n438 4.67295
R21922 commonsourceibias.n471 commonsourceibias.n395 4.67295
R21923 commonsourceibias.n586 commonsourceibias.n374 4.67295
R21924 commonsourceibias.n555 commonsourceibias.n554 4.67295
R21925 commonsourceibias commonsourceibias.n734 4.20978
R21926 commonsourceibias.n320 commonsourceibias.n319 4.18111
R21927 commonsourceibias.n266 commonsourceibias.n264 4.18111
R21928 commonsourceibias.n29 commonsourceibias.n27 4.18111
R21929 commonsourceibias.n83 commonsourceibias.n82 4.18111
R21930 commonsourceibias.n150 commonsourceibias.n13 4.18111
R21931 commonsourceibias.n203 commonsourceibias.n151 4.18111
R21932 commonsourceibias.n684 commonsourceibias.n683 4.18111
R21933 commonsourceibias.n686 commonsourceibias.n629 4.18111
R21934 commonsourceibias.n454 commonsourceibias.n453 4.18111
R21935 commonsourceibias.n456 commonsourceibias.n399 4.18111
R21936 commonsourceibias.n571 commonsourceibias.n378 4.18111
R21937 commonsourceibias.n567 commonsourceibias.n515 4.18111
R21938 commonsourceibias.n271 commonsourceibias.n269 3.68928
R21939 commonsourceibias.n334 commonsourceibias.n333 3.68928
R21940 commonsourceibias.n97 commonsourceibias.n96 3.68928
R21941 commonsourceibias.n34 commonsourceibias.n32 3.68928
R21942 commonsourceibias.n219 commonsourceibias.n218 3.68928
R21943 commonsourceibias.n196 commonsourceibias.n155 3.68928
R21944 commonsourceibias.n671 commonsourceibias.n633 3.68928
R21945 commonsourceibias.n699 commonsourceibias.n698 3.68928
R21946 commonsourceibias.n441 commonsourceibias.n403 3.68928
R21947 commonsourceibias.n469 commonsourceibias.n468 3.68928
R21948 commonsourceibias.n584 commonsourceibias.n583 3.68928
R21949 commonsourceibias.n560 commonsourceibias.n519 3.68928
R21950 commonsourceibias.n276 commonsourceibias.n274 3.19744
R21951 commonsourceibias.n348 commonsourceibias.n347 3.19744
R21952 commonsourceibias.n111 commonsourceibias.n110 3.19744
R21953 commonsourceibias.n39 commonsourceibias.n37 3.19744
R21954 commonsourceibias.n233 commonsourceibias.n232 3.19744
R21955 commonsourceibias.n161 commonsourceibias.n159 3.19744
R21956 commonsourceibias.n656 commonsourceibias.n637 3.19744
R21957 commonsourceibias.n714 commonsourceibias.n713 3.19744
R21958 commonsourceibias.n426 commonsourceibias.n407 3.19744
R21959 commonsourceibias.n484 commonsourceibias.n483 3.19744
R21960 commonsourceibias.n599 commonsourceibias.n598 3.19744
R21961 commonsourceibias.n542 commonsourceibias.n523 3.19744
R21962 commonsourceibias.n139 commonsourceibias.t47 2.82907
R21963 commonsourceibias.n139 commonsourceibias.t79 2.82907
R21964 commonsourceibias.n140 commonsourceibias.t53 2.82907
R21965 commonsourceibias.n140 commonsourceibias.t5 2.82907
R21966 commonsourceibias.n142 commonsourceibias.t19 2.82907
R21967 commonsourceibias.n142 commonsourceibias.t23 2.82907
R21968 commonsourceibias.n144 commonsourceibias.t39 2.82907
R21969 commonsourceibias.n144 commonsourceibias.t71 2.82907
R21970 commonsourceibias.n146 commonsourceibias.t57 2.82907
R21971 commonsourceibias.n146 commonsourceibias.t27 2.82907
R21972 commonsourceibias.n137 commonsourceibias.t11 2.82907
R21973 commonsourceibias.n137 commonsourceibias.t41 2.82907
R21974 commonsourceibias.n135 commonsourceibias.t25 2.82907
R21975 commonsourceibias.n135 commonsourceibias.t35 2.82907
R21976 commonsourceibias.n133 commonsourceibias.t37 2.82907
R21977 commonsourceibias.n133 commonsourceibias.t77 2.82907
R21978 commonsourceibias.n131 commonsourceibias.t51 2.82907
R21979 commonsourceibias.n131 commonsourceibias.t9 2.82907
R21980 commonsourceibias.n129 commonsourceibias.t75 2.82907
R21981 commonsourceibias.n129 commonsourceibias.t21 2.82907
R21982 commonsourceibias.n503 commonsourceibias.t43 2.82907
R21983 commonsourceibias.n503 commonsourceibias.t13 2.82907
R21984 commonsourceibias.n505 commonsourceibias.t29 2.82907
R21985 commonsourceibias.n505 commonsourceibias.t1 2.82907
R21986 commonsourceibias.n507 commonsourceibias.t17 2.82907
R21987 commonsourceibias.n507 commonsourceibias.t61 2.82907
R21988 commonsourceibias.n509 commonsourceibias.t59 2.82907
R21989 commonsourceibias.n509 commonsourceibias.t45 2.82907
R21990 commonsourceibias.n511 commonsourceibias.t65 2.82907
R21991 commonsourceibias.n511 commonsourceibias.t33 2.82907
R21992 commonsourceibias.n386 commonsourceibias.t55 2.82907
R21993 commonsourceibias.n386 commonsourceibias.t73 2.82907
R21994 commonsourceibias.n384 commonsourceibias.t7 2.82907
R21995 commonsourceibias.n384 commonsourceibias.t63 2.82907
R21996 commonsourceibias.n382 commonsourceibias.t69 2.82907
R21997 commonsourceibias.n382 commonsourceibias.t67 2.82907
R21998 commonsourceibias.n380 commonsourceibias.t49 2.82907
R21999 commonsourceibias.n380 commonsourceibias.t15 2.82907
R22000 commonsourceibias.n379 commonsourceibias.t31 2.82907
R22001 commonsourceibias.n379 commonsourceibias.t3 2.82907
R22002 commonsourceibias.n280 commonsourceibias.n279 2.7056
R22003 commonsourceibias.n362 commonsourceibias.n361 2.7056
R22004 commonsourceibias.n125 commonsourceibias.n124 2.7056
R22005 commonsourceibias.n43 commonsourceibias.n42 2.7056
R22006 commonsourceibias.n247 commonsourceibias.n246 2.7056
R22007 commonsourceibias.n165 commonsourceibias.n164 2.7056
R22008 commonsourceibias.n642 commonsourceibias.n641 2.7056
R22009 commonsourceibias.n729 commonsourceibias.n728 2.7056
R22010 commonsourceibias.n412 commonsourceibias.n411 2.7056
R22011 commonsourceibias.n499 commonsourceibias.n498 2.7056
R22012 commonsourceibias.n614 commonsourceibias.n613 2.7056
R22013 commonsourceibias.n528 commonsourceibias.n527 2.7056
R22014 commonsourceibias.n132 commonsourceibias.n130 0.573776
R22015 commonsourceibias.n134 commonsourceibias.n132 0.573776
R22016 commonsourceibias.n136 commonsourceibias.n134 0.573776
R22017 commonsourceibias.n138 commonsourceibias.n136 0.573776
R22018 commonsourceibias.n147 commonsourceibias.n145 0.573776
R22019 commonsourceibias.n145 commonsourceibias.n143 0.573776
R22020 commonsourceibias.n143 commonsourceibias.n141 0.573776
R22021 commonsourceibias.n383 commonsourceibias.n381 0.573776
R22022 commonsourceibias.n385 commonsourceibias.n383 0.573776
R22023 commonsourceibias.n387 commonsourceibias.n385 0.573776
R22024 commonsourceibias.n512 commonsourceibias.n510 0.573776
R22025 commonsourceibias.n510 commonsourceibias.n508 0.573776
R22026 commonsourceibias.n508 commonsourceibias.n506 0.573776
R22027 commonsourceibias.n506 commonsourceibias.n504 0.573776
R22028 commonsourceibias.n148 commonsourceibias.n138 0.287138
R22029 commonsourceibias.n148 commonsourceibias.n147 0.287138
R22030 commonsourceibias.n513 commonsourceibias.n387 0.287138
R22031 commonsourceibias.n513 commonsourceibias.n512 0.287138
R22032 commonsourceibias.n365 commonsourceibias.n251 0.285035
R22033 commonsourceibias.n128 commonsourceibias.n14 0.285035
R22034 commonsourceibias.n250 commonsourceibias.n0 0.285035
R22035 commonsourceibias.n732 commonsourceibias.n618 0.285035
R22036 commonsourceibias.n502 commonsourceibias.n388 0.285035
R22037 commonsourceibias.n617 commonsourceibias.n367 0.285035
R22038 commonsourceibias.n360 commonsourceibias.n251 0.189894
R22039 commonsourceibias.n360 commonsourceibias.n359 0.189894
R22040 commonsourceibias.n359 commonsourceibias.n358 0.189894
R22041 commonsourceibias.n358 commonsourceibias.n253 0.189894
R22042 commonsourceibias.n353 commonsourceibias.n253 0.189894
R22043 commonsourceibias.n353 commonsourceibias.n352 0.189894
R22044 commonsourceibias.n352 commonsourceibias.n351 0.189894
R22045 commonsourceibias.n351 commonsourceibias.n255 0.189894
R22046 commonsourceibias.n346 commonsourceibias.n255 0.189894
R22047 commonsourceibias.n346 commonsourceibias.n345 0.189894
R22048 commonsourceibias.n345 commonsourceibias.n344 0.189894
R22049 commonsourceibias.n344 commonsourceibias.n258 0.189894
R22050 commonsourceibias.n339 commonsourceibias.n258 0.189894
R22051 commonsourceibias.n339 commonsourceibias.n338 0.189894
R22052 commonsourceibias.n338 commonsourceibias.n337 0.189894
R22053 commonsourceibias.n337 commonsourceibias.n260 0.189894
R22054 commonsourceibias.n332 commonsourceibias.n260 0.189894
R22055 commonsourceibias.n332 commonsourceibias.n331 0.189894
R22056 commonsourceibias.n331 commonsourceibias.n330 0.189894
R22057 commonsourceibias.n330 commonsourceibias.n263 0.189894
R22058 commonsourceibias.n325 commonsourceibias.n263 0.189894
R22059 commonsourceibias.n325 commonsourceibias.n324 0.189894
R22060 commonsourceibias.n324 commonsourceibias.n323 0.189894
R22061 commonsourceibias.n323 commonsourceibias.n265 0.189894
R22062 commonsourceibias.n318 commonsourceibias.n265 0.189894
R22063 commonsourceibias.n318 commonsourceibias.n317 0.189894
R22064 commonsourceibias.n317 commonsourceibias.n316 0.189894
R22065 commonsourceibias.n316 commonsourceibias.n268 0.189894
R22066 commonsourceibias.n311 commonsourceibias.n268 0.189894
R22067 commonsourceibias.n311 commonsourceibias.n310 0.189894
R22068 commonsourceibias.n310 commonsourceibias.n309 0.189894
R22069 commonsourceibias.n309 commonsourceibias.n270 0.189894
R22070 commonsourceibias.n304 commonsourceibias.n270 0.189894
R22071 commonsourceibias.n304 commonsourceibias.n303 0.189894
R22072 commonsourceibias.n303 commonsourceibias.n302 0.189894
R22073 commonsourceibias.n302 commonsourceibias.n273 0.189894
R22074 commonsourceibias.n297 commonsourceibias.n273 0.189894
R22075 commonsourceibias.n297 commonsourceibias.n296 0.189894
R22076 commonsourceibias.n296 commonsourceibias.n295 0.189894
R22077 commonsourceibias.n295 commonsourceibias.n275 0.189894
R22078 commonsourceibias.n290 commonsourceibias.n275 0.189894
R22079 commonsourceibias.n290 commonsourceibias.n289 0.189894
R22080 commonsourceibias.n289 commonsourceibias.n288 0.189894
R22081 commonsourceibias.n288 commonsourceibias.n278 0.189894
R22082 commonsourceibias.n283 commonsourceibias.n278 0.189894
R22083 commonsourceibias.n283 commonsourceibias.n282 0.189894
R22084 commonsourceibias.n123 commonsourceibias.n14 0.189894
R22085 commonsourceibias.n123 commonsourceibias.n122 0.189894
R22086 commonsourceibias.n122 commonsourceibias.n121 0.189894
R22087 commonsourceibias.n121 commonsourceibias.n16 0.189894
R22088 commonsourceibias.n116 commonsourceibias.n16 0.189894
R22089 commonsourceibias.n116 commonsourceibias.n115 0.189894
R22090 commonsourceibias.n115 commonsourceibias.n114 0.189894
R22091 commonsourceibias.n114 commonsourceibias.n18 0.189894
R22092 commonsourceibias.n109 commonsourceibias.n18 0.189894
R22093 commonsourceibias.n109 commonsourceibias.n108 0.189894
R22094 commonsourceibias.n108 commonsourceibias.n107 0.189894
R22095 commonsourceibias.n107 commonsourceibias.n21 0.189894
R22096 commonsourceibias.n102 commonsourceibias.n21 0.189894
R22097 commonsourceibias.n102 commonsourceibias.n101 0.189894
R22098 commonsourceibias.n101 commonsourceibias.n100 0.189894
R22099 commonsourceibias.n100 commonsourceibias.n23 0.189894
R22100 commonsourceibias.n95 commonsourceibias.n23 0.189894
R22101 commonsourceibias.n95 commonsourceibias.n94 0.189894
R22102 commonsourceibias.n94 commonsourceibias.n93 0.189894
R22103 commonsourceibias.n93 commonsourceibias.n26 0.189894
R22104 commonsourceibias.n88 commonsourceibias.n26 0.189894
R22105 commonsourceibias.n88 commonsourceibias.n87 0.189894
R22106 commonsourceibias.n87 commonsourceibias.n86 0.189894
R22107 commonsourceibias.n86 commonsourceibias.n28 0.189894
R22108 commonsourceibias.n81 commonsourceibias.n28 0.189894
R22109 commonsourceibias.n81 commonsourceibias.n80 0.189894
R22110 commonsourceibias.n80 commonsourceibias.n79 0.189894
R22111 commonsourceibias.n79 commonsourceibias.n31 0.189894
R22112 commonsourceibias.n74 commonsourceibias.n31 0.189894
R22113 commonsourceibias.n74 commonsourceibias.n73 0.189894
R22114 commonsourceibias.n73 commonsourceibias.n72 0.189894
R22115 commonsourceibias.n72 commonsourceibias.n33 0.189894
R22116 commonsourceibias.n67 commonsourceibias.n33 0.189894
R22117 commonsourceibias.n67 commonsourceibias.n66 0.189894
R22118 commonsourceibias.n66 commonsourceibias.n65 0.189894
R22119 commonsourceibias.n65 commonsourceibias.n36 0.189894
R22120 commonsourceibias.n60 commonsourceibias.n36 0.189894
R22121 commonsourceibias.n60 commonsourceibias.n59 0.189894
R22122 commonsourceibias.n59 commonsourceibias.n58 0.189894
R22123 commonsourceibias.n58 commonsourceibias.n38 0.189894
R22124 commonsourceibias.n53 commonsourceibias.n38 0.189894
R22125 commonsourceibias.n53 commonsourceibias.n52 0.189894
R22126 commonsourceibias.n52 commonsourceibias.n51 0.189894
R22127 commonsourceibias.n51 commonsourceibias.n41 0.189894
R22128 commonsourceibias.n46 commonsourceibias.n41 0.189894
R22129 commonsourceibias.n46 commonsourceibias.n45 0.189894
R22130 commonsourceibias.n205 commonsourceibias.n204 0.189894
R22131 commonsourceibias.n204 commonsourceibias.n152 0.189894
R22132 commonsourceibias.n200 commonsourceibias.n152 0.189894
R22133 commonsourceibias.n200 commonsourceibias.n199 0.189894
R22134 commonsourceibias.n199 commonsourceibias.n154 0.189894
R22135 commonsourceibias.n195 commonsourceibias.n154 0.189894
R22136 commonsourceibias.n195 commonsourceibias.n194 0.189894
R22137 commonsourceibias.n194 commonsourceibias.n156 0.189894
R22138 commonsourceibias.n189 commonsourceibias.n156 0.189894
R22139 commonsourceibias.n189 commonsourceibias.n188 0.189894
R22140 commonsourceibias.n188 commonsourceibias.n187 0.189894
R22141 commonsourceibias.n187 commonsourceibias.n158 0.189894
R22142 commonsourceibias.n182 commonsourceibias.n158 0.189894
R22143 commonsourceibias.n182 commonsourceibias.n181 0.189894
R22144 commonsourceibias.n181 commonsourceibias.n180 0.189894
R22145 commonsourceibias.n180 commonsourceibias.n160 0.189894
R22146 commonsourceibias.n175 commonsourceibias.n160 0.189894
R22147 commonsourceibias.n175 commonsourceibias.n174 0.189894
R22148 commonsourceibias.n174 commonsourceibias.n173 0.189894
R22149 commonsourceibias.n173 commonsourceibias.n163 0.189894
R22150 commonsourceibias.n168 commonsourceibias.n163 0.189894
R22151 commonsourceibias.n168 commonsourceibias.n167 0.189894
R22152 commonsourceibias.n245 commonsourceibias.n0 0.189894
R22153 commonsourceibias.n245 commonsourceibias.n244 0.189894
R22154 commonsourceibias.n244 commonsourceibias.n243 0.189894
R22155 commonsourceibias.n243 commonsourceibias.n2 0.189894
R22156 commonsourceibias.n238 commonsourceibias.n2 0.189894
R22157 commonsourceibias.n238 commonsourceibias.n237 0.189894
R22158 commonsourceibias.n237 commonsourceibias.n236 0.189894
R22159 commonsourceibias.n236 commonsourceibias.n4 0.189894
R22160 commonsourceibias.n231 commonsourceibias.n4 0.189894
R22161 commonsourceibias.n231 commonsourceibias.n230 0.189894
R22162 commonsourceibias.n230 commonsourceibias.n229 0.189894
R22163 commonsourceibias.n229 commonsourceibias.n7 0.189894
R22164 commonsourceibias.n224 commonsourceibias.n7 0.189894
R22165 commonsourceibias.n224 commonsourceibias.n223 0.189894
R22166 commonsourceibias.n223 commonsourceibias.n222 0.189894
R22167 commonsourceibias.n222 commonsourceibias.n9 0.189894
R22168 commonsourceibias.n217 commonsourceibias.n9 0.189894
R22169 commonsourceibias.n217 commonsourceibias.n216 0.189894
R22170 commonsourceibias.n216 commonsourceibias.n215 0.189894
R22171 commonsourceibias.n215 commonsourceibias.n12 0.189894
R22172 commonsourceibias.n210 commonsourceibias.n12 0.189894
R22173 commonsourceibias.n210 commonsourceibias.n209 0.189894
R22174 commonsourceibias.n209 commonsourceibias.n208 0.189894
R22175 commonsourceibias.n645 commonsourceibias.n644 0.189894
R22176 commonsourceibias.n645 commonsourceibias.n640 0.189894
R22177 commonsourceibias.n650 commonsourceibias.n640 0.189894
R22178 commonsourceibias.n651 commonsourceibias.n650 0.189894
R22179 commonsourceibias.n652 commonsourceibias.n651 0.189894
R22180 commonsourceibias.n652 commonsourceibias.n638 0.189894
R22181 commonsourceibias.n658 commonsourceibias.n638 0.189894
R22182 commonsourceibias.n659 commonsourceibias.n658 0.189894
R22183 commonsourceibias.n660 commonsourceibias.n659 0.189894
R22184 commonsourceibias.n660 commonsourceibias.n636 0.189894
R22185 commonsourceibias.n665 commonsourceibias.n636 0.189894
R22186 commonsourceibias.n666 commonsourceibias.n665 0.189894
R22187 commonsourceibias.n667 commonsourceibias.n666 0.189894
R22188 commonsourceibias.n667 commonsourceibias.n634 0.189894
R22189 commonsourceibias.n673 commonsourceibias.n634 0.189894
R22190 commonsourceibias.n674 commonsourceibias.n673 0.189894
R22191 commonsourceibias.n675 commonsourceibias.n674 0.189894
R22192 commonsourceibias.n675 commonsourceibias.n632 0.189894
R22193 commonsourceibias.n680 commonsourceibias.n632 0.189894
R22194 commonsourceibias.n681 commonsourceibias.n680 0.189894
R22195 commonsourceibias.n682 commonsourceibias.n681 0.189894
R22196 commonsourceibias.n682 commonsourceibias.n630 0.189894
R22197 commonsourceibias.n688 commonsourceibias.n630 0.189894
R22198 commonsourceibias.n689 commonsourceibias.n688 0.189894
R22199 commonsourceibias.n690 commonsourceibias.n689 0.189894
R22200 commonsourceibias.n690 commonsourceibias.n628 0.189894
R22201 commonsourceibias.n695 commonsourceibias.n628 0.189894
R22202 commonsourceibias.n696 commonsourceibias.n695 0.189894
R22203 commonsourceibias.n697 commonsourceibias.n696 0.189894
R22204 commonsourceibias.n697 commonsourceibias.n626 0.189894
R22205 commonsourceibias.n703 commonsourceibias.n626 0.189894
R22206 commonsourceibias.n704 commonsourceibias.n703 0.189894
R22207 commonsourceibias.n705 commonsourceibias.n704 0.189894
R22208 commonsourceibias.n705 commonsourceibias.n624 0.189894
R22209 commonsourceibias.n710 commonsourceibias.n624 0.189894
R22210 commonsourceibias.n711 commonsourceibias.n710 0.189894
R22211 commonsourceibias.n712 commonsourceibias.n711 0.189894
R22212 commonsourceibias.n712 commonsourceibias.n622 0.189894
R22213 commonsourceibias.n718 commonsourceibias.n622 0.189894
R22214 commonsourceibias.n719 commonsourceibias.n718 0.189894
R22215 commonsourceibias.n720 commonsourceibias.n719 0.189894
R22216 commonsourceibias.n720 commonsourceibias.n620 0.189894
R22217 commonsourceibias.n725 commonsourceibias.n620 0.189894
R22218 commonsourceibias.n726 commonsourceibias.n725 0.189894
R22219 commonsourceibias.n727 commonsourceibias.n726 0.189894
R22220 commonsourceibias.n727 commonsourceibias.n618 0.189894
R22221 commonsourceibias.n415 commonsourceibias.n414 0.189894
R22222 commonsourceibias.n415 commonsourceibias.n410 0.189894
R22223 commonsourceibias.n420 commonsourceibias.n410 0.189894
R22224 commonsourceibias.n421 commonsourceibias.n420 0.189894
R22225 commonsourceibias.n422 commonsourceibias.n421 0.189894
R22226 commonsourceibias.n422 commonsourceibias.n408 0.189894
R22227 commonsourceibias.n428 commonsourceibias.n408 0.189894
R22228 commonsourceibias.n429 commonsourceibias.n428 0.189894
R22229 commonsourceibias.n430 commonsourceibias.n429 0.189894
R22230 commonsourceibias.n430 commonsourceibias.n406 0.189894
R22231 commonsourceibias.n435 commonsourceibias.n406 0.189894
R22232 commonsourceibias.n436 commonsourceibias.n435 0.189894
R22233 commonsourceibias.n437 commonsourceibias.n436 0.189894
R22234 commonsourceibias.n437 commonsourceibias.n404 0.189894
R22235 commonsourceibias.n443 commonsourceibias.n404 0.189894
R22236 commonsourceibias.n444 commonsourceibias.n443 0.189894
R22237 commonsourceibias.n445 commonsourceibias.n444 0.189894
R22238 commonsourceibias.n445 commonsourceibias.n402 0.189894
R22239 commonsourceibias.n450 commonsourceibias.n402 0.189894
R22240 commonsourceibias.n451 commonsourceibias.n450 0.189894
R22241 commonsourceibias.n452 commonsourceibias.n451 0.189894
R22242 commonsourceibias.n452 commonsourceibias.n400 0.189894
R22243 commonsourceibias.n458 commonsourceibias.n400 0.189894
R22244 commonsourceibias.n459 commonsourceibias.n458 0.189894
R22245 commonsourceibias.n460 commonsourceibias.n459 0.189894
R22246 commonsourceibias.n460 commonsourceibias.n398 0.189894
R22247 commonsourceibias.n465 commonsourceibias.n398 0.189894
R22248 commonsourceibias.n466 commonsourceibias.n465 0.189894
R22249 commonsourceibias.n467 commonsourceibias.n466 0.189894
R22250 commonsourceibias.n467 commonsourceibias.n396 0.189894
R22251 commonsourceibias.n473 commonsourceibias.n396 0.189894
R22252 commonsourceibias.n474 commonsourceibias.n473 0.189894
R22253 commonsourceibias.n475 commonsourceibias.n474 0.189894
R22254 commonsourceibias.n475 commonsourceibias.n394 0.189894
R22255 commonsourceibias.n480 commonsourceibias.n394 0.189894
R22256 commonsourceibias.n481 commonsourceibias.n480 0.189894
R22257 commonsourceibias.n482 commonsourceibias.n481 0.189894
R22258 commonsourceibias.n482 commonsourceibias.n392 0.189894
R22259 commonsourceibias.n488 commonsourceibias.n392 0.189894
R22260 commonsourceibias.n489 commonsourceibias.n488 0.189894
R22261 commonsourceibias.n490 commonsourceibias.n489 0.189894
R22262 commonsourceibias.n490 commonsourceibias.n390 0.189894
R22263 commonsourceibias.n495 commonsourceibias.n390 0.189894
R22264 commonsourceibias.n496 commonsourceibias.n495 0.189894
R22265 commonsourceibias.n497 commonsourceibias.n496 0.189894
R22266 commonsourceibias.n497 commonsourceibias.n388 0.189894
R22267 commonsourceibias.n531 commonsourceibias.n530 0.189894
R22268 commonsourceibias.n531 commonsourceibias.n526 0.189894
R22269 commonsourceibias.n536 commonsourceibias.n526 0.189894
R22270 commonsourceibias.n537 commonsourceibias.n536 0.189894
R22271 commonsourceibias.n538 commonsourceibias.n537 0.189894
R22272 commonsourceibias.n538 commonsourceibias.n524 0.189894
R22273 commonsourceibias.n544 commonsourceibias.n524 0.189894
R22274 commonsourceibias.n545 commonsourceibias.n544 0.189894
R22275 commonsourceibias.n546 commonsourceibias.n545 0.189894
R22276 commonsourceibias.n546 commonsourceibias.n522 0.189894
R22277 commonsourceibias.n551 commonsourceibias.n522 0.189894
R22278 commonsourceibias.n552 commonsourceibias.n551 0.189894
R22279 commonsourceibias.n553 commonsourceibias.n552 0.189894
R22280 commonsourceibias.n553 commonsourceibias.n520 0.189894
R22281 commonsourceibias.n558 commonsourceibias.n520 0.189894
R22282 commonsourceibias.n559 commonsourceibias.n558 0.189894
R22283 commonsourceibias.n559 commonsourceibias.n518 0.189894
R22284 commonsourceibias.n563 commonsourceibias.n518 0.189894
R22285 commonsourceibias.n564 commonsourceibias.n563 0.189894
R22286 commonsourceibias.n564 commonsourceibias.n516 0.189894
R22287 commonsourceibias.n568 commonsourceibias.n516 0.189894
R22288 commonsourceibias.n569 commonsourceibias.n568 0.189894
R22289 commonsourceibias.n574 commonsourceibias.n573 0.189894
R22290 commonsourceibias.n575 commonsourceibias.n574 0.189894
R22291 commonsourceibias.n575 commonsourceibias.n377 0.189894
R22292 commonsourceibias.n580 commonsourceibias.n377 0.189894
R22293 commonsourceibias.n581 commonsourceibias.n580 0.189894
R22294 commonsourceibias.n582 commonsourceibias.n581 0.189894
R22295 commonsourceibias.n582 commonsourceibias.n375 0.189894
R22296 commonsourceibias.n588 commonsourceibias.n375 0.189894
R22297 commonsourceibias.n589 commonsourceibias.n588 0.189894
R22298 commonsourceibias.n590 commonsourceibias.n589 0.189894
R22299 commonsourceibias.n590 commonsourceibias.n373 0.189894
R22300 commonsourceibias.n595 commonsourceibias.n373 0.189894
R22301 commonsourceibias.n596 commonsourceibias.n595 0.189894
R22302 commonsourceibias.n597 commonsourceibias.n596 0.189894
R22303 commonsourceibias.n597 commonsourceibias.n371 0.189894
R22304 commonsourceibias.n603 commonsourceibias.n371 0.189894
R22305 commonsourceibias.n604 commonsourceibias.n603 0.189894
R22306 commonsourceibias.n605 commonsourceibias.n604 0.189894
R22307 commonsourceibias.n605 commonsourceibias.n369 0.189894
R22308 commonsourceibias.n610 commonsourceibias.n369 0.189894
R22309 commonsourceibias.n611 commonsourceibias.n610 0.189894
R22310 commonsourceibias.n612 commonsourceibias.n611 0.189894
R22311 commonsourceibias.n612 commonsourceibias.n367 0.189894
R22312 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R22313 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R22314 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R22315 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R22316 diffpairibias.n0 diffpairibias.t27 436.822
R22317 diffpairibias.n27 diffpairibias.t24 435.479
R22318 diffpairibias.n26 diffpairibias.t21 435.479
R22319 diffpairibias.n25 diffpairibias.t22 435.479
R22320 diffpairibias.n24 diffpairibias.t26 435.479
R22321 diffpairibias.n23 diffpairibias.t20 435.479
R22322 diffpairibias.n0 diffpairibias.t23 435.479
R22323 diffpairibias.n1 diffpairibias.t28 435.479
R22324 diffpairibias.n2 diffpairibias.t25 435.479
R22325 diffpairibias.n3 diffpairibias.t29 435.479
R22326 diffpairibias.n13 diffpairibias.t14 377.536
R22327 diffpairibias.n13 diffpairibias.t0 376.193
R22328 diffpairibias.n14 diffpairibias.t10 376.193
R22329 diffpairibias.n15 diffpairibias.t12 376.193
R22330 diffpairibias.n16 diffpairibias.t6 376.193
R22331 diffpairibias.n17 diffpairibias.t2 376.193
R22332 diffpairibias.n18 diffpairibias.t16 376.193
R22333 diffpairibias.n19 diffpairibias.t4 376.193
R22334 diffpairibias.n20 diffpairibias.t18 376.193
R22335 diffpairibias.n21 diffpairibias.t8 376.193
R22336 diffpairibias.n4 diffpairibias.t15 113.368
R22337 diffpairibias.n4 diffpairibias.t1 112.698
R22338 diffpairibias.n5 diffpairibias.t11 112.698
R22339 diffpairibias.n6 diffpairibias.t13 112.698
R22340 diffpairibias.n7 diffpairibias.t7 112.698
R22341 diffpairibias.n8 diffpairibias.t3 112.698
R22342 diffpairibias.n9 diffpairibias.t17 112.698
R22343 diffpairibias.n10 diffpairibias.t5 112.698
R22344 diffpairibias.n11 diffpairibias.t19 112.698
R22345 diffpairibias.n12 diffpairibias.t9 112.698
R22346 diffpairibias.n22 diffpairibias.n21 4.77242
R22347 diffpairibias.n22 diffpairibias.n12 4.30807
R22348 diffpairibias.n23 diffpairibias.n22 4.13945
R22349 diffpairibias.n21 diffpairibias.n20 1.34352
R22350 diffpairibias.n20 diffpairibias.n19 1.34352
R22351 diffpairibias.n19 diffpairibias.n18 1.34352
R22352 diffpairibias.n18 diffpairibias.n17 1.34352
R22353 diffpairibias.n17 diffpairibias.n16 1.34352
R22354 diffpairibias.n16 diffpairibias.n15 1.34352
R22355 diffpairibias.n15 diffpairibias.n14 1.34352
R22356 diffpairibias.n14 diffpairibias.n13 1.34352
R22357 diffpairibias.n3 diffpairibias.n2 1.34352
R22358 diffpairibias.n2 diffpairibias.n1 1.34352
R22359 diffpairibias.n1 diffpairibias.n0 1.34352
R22360 diffpairibias.n24 diffpairibias.n23 1.34352
R22361 diffpairibias.n25 diffpairibias.n24 1.34352
R22362 diffpairibias.n26 diffpairibias.n25 1.34352
R22363 diffpairibias.n27 diffpairibias.n26 1.34352
R22364 diffpairibias.n28 diffpairibias.n27 0.862419
R22365 diffpairibias diffpairibias.n28 0.684875
R22366 diffpairibias.n12 diffpairibias.n11 0.672012
R22367 diffpairibias.n11 diffpairibias.n10 0.672012
R22368 diffpairibias.n10 diffpairibias.n9 0.672012
R22369 diffpairibias.n9 diffpairibias.n8 0.672012
R22370 diffpairibias.n8 diffpairibias.n7 0.672012
R22371 diffpairibias.n7 diffpairibias.n6 0.672012
R22372 diffpairibias.n6 diffpairibias.n5 0.672012
R22373 diffpairibias.n5 diffpairibias.n4 0.672012
R22374 diffpairibias.n28 diffpairibias.n3 0.190907
R22375 minus.n76 minus.t28 250.337
R22376 minus.n15 minus.t20 250.337
R22377 minus.n126 minus.t1 243.255
R22378 minus.n120 minus.t8 231.093
R22379 minus.n59 minus.t10 231.093
R22380 minus.n125 minus.n123 224.169
R22381 minus.n125 minus.n124 223.454
R22382 minus.n62 minus.t12 187.445
R22383 minus.n113 minus.t18 187.445
R22384 minus.n107 minus.t25 187.445
R22385 minus.n66 minus.t22 187.445
R22386 minus.n68 minus.t19 187.445
R22387 minus.n95 minus.t7 187.445
R22388 minus.n89 minus.t6 187.445
R22389 minus.n72 minus.t16 187.445
R22390 minus.n74 minus.t15 187.445
R22391 minus.n77 minus.t23 187.445
R22392 minus.n16 minus.t14 187.445
R22393 minus.n13 minus.t9 187.445
R22394 minus.n11 minus.t5 187.445
R22395 minus.n28 minus.t26 187.445
R22396 minus.n34 minus.t27 187.445
R22397 minus.n7 minus.t21 187.445
R22398 minus.n5 minus.t24 187.445
R22399 minus.n46 minus.t17 187.445
R22400 minus.n52 minus.t11 187.445
R22401 minus.n1 minus.t13 187.445
R22402 minus.n78 minus.n75 161.3
R22403 minus.n80 minus.n79 161.3
R22404 minus.n82 minus.n81 161.3
R22405 minus.n83 minus.n73 161.3
R22406 minus.n85 minus.n84 161.3
R22407 minus.n87 minus.n86 161.3
R22408 minus.n88 minus.n71 161.3
R22409 minus.n91 minus.n90 161.3
R22410 minus.n92 minus.n70 161.3
R22411 minus.n94 minus.n93 161.3
R22412 minus.n96 minus.n69 161.3
R22413 minus.n98 minus.n97 161.3
R22414 minus.n100 minus.n99 161.3
R22415 minus.n101 minus.n67 161.3
R22416 minus.n103 minus.n102 161.3
R22417 minus.n105 minus.n104 161.3
R22418 minus.n106 minus.n65 161.3
R22419 minus.n109 minus.n108 161.3
R22420 minus.n110 minus.n64 161.3
R22421 minus.n112 minus.n111 161.3
R22422 minus.n114 minus.n63 161.3
R22423 minus.n116 minus.n115 161.3
R22424 minus.n118 minus.n117 161.3
R22425 minus.n119 minus.n61 161.3
R22426 minus.n121 minus.n120 161.3
R22427 minus.n60 minus.n59 161.3
R22428 minus.n58 minus.n0 161.3
R22429 minus.n57 minus.n56 161.3
R22430 minus.n55 minus.n54 161.3
R22431 minus.n53 minus.n2 161.3
R22432 minus.n51 minus.n50 161.3
R22433 minus.n49 minus.n3 161.3
R22434 minus.n48 minus.n47 161.3
R22435 minus.n45 minus.n4 161.3
R22436 minus.n44 minus.n43 161.3
R22437 minus.n42 minus.n41 161.3
R22438 minus.n40 minus.n6 161.3
R22439 minus.n39 minus.n38 161.3
R22440 minus.n37 minus.n36 161.3
R22441 minus.n35 minus.n8 161.3
R22442 minus.n33 minus.n32 161.3
R22443 minus.n31 minus.n9 161.3
R22444 minus.n30 minus.n29 161.3
R22445 minus.n27 minus.n10 161.3
R22446 minus.n26 minus.n25 161.3
R22447 minus.n24 minus.n23 161.3
R22448 minus.n22 minus.n12 161.3
R22449 minus.n21 minus.n20 161.3
R22450 minus.n19 minus.n18 161.3
R22451 minus.n17 minus.n14 161.3
R22452 minus.n106 minus.n105 56.5617
R22453 minus.n97 minus.n96 56.5617
R22454 minus.n88 minus.n87 56.5617
R22455 minus.n27 minus.n26 56.5617
R22456 minus.n36 minus.n35 56.5617
R22457 minus.n45 minus.n44 56.5617
R22458 minus.n115 minus.n114 56.5617
R22459 minus.n79 minus.n78 56.5617
R22460 minus.n18 minus.n17 56.5617
R22461 minus.n54 minus.n53 56.5617
R22462 minus.n119 minus.n118 50.2647
R22463 minus.n58 minus.n57 50.2647
R22464 minus.n108 minus.n64 46.3896
R22465 minus.n84 minus.n83 46.3896
R22466 minus.n23 minus.n22 46.3896
R22467 minus.n47 minus.n3 46.3896
R22468 minus.n76 minus.n75 43.1929
R22469 minus.n15 minus.n14 43.1929
R22470 minus.n101 minus.n100 42.5146
R22471 minus.n94 minus.n70 42.5146
R22472 minus.n33 minus.n9 42.5146
R22473 minus.n40 minus.n39 42.5146
R22474 minus.n77 minus.n76 40.6041
R22475 minus.n16 minus.n15 40.6041
R22476 minus.n102 minus.n101 38.6395
R22477 minus.n90 minus.n70 38.6395
R22478 minus.n29 minus.n9 38.6395
R22479 minus.n41 minus.n40 38.6395
R22480 minus.n122 minus.n121 35.4191
R22481 minus.n112 minus.n64 34.7644
R22482 minus.n83 minus.n82 34.7644
R22483 minus.n22 minus.n21 34.7644
R22484 minus.n51 minus.n3 34.7644
R22485 minus.n114 minus.n113 21.8872
R22486 minus.n79 minus.n74 21.8872
R22487 minus.n18 minus.n13 21.8872
R22488 minus.n53 minus.n52 21.8872
R22489 minus.n105 minus.n66 19.9199
R22490 minus.n89 minus.n88 19.9199
R22491 minus.n28 minus.n27 19.9199
R22492 minus.n44 minus.n5 19.9199
R22493 minus.n124 minus.t0 19.8005
R22494 minus.n124 minus.t2 19.8005
R22495 minus.n123 minus.t4 19.8005
R22496 minus.n123 minus.t3 19.8005
R22497 minus.n97 minus.n68 17.9525
R22498 minus.n96 minus.n95 17.9525
R22499 minus.n35 minus.n34 17.9525
R22500 minus.n36 minus.n7 17.9525
R22501 minus.n107 minus.n106 15.9852
R22502 minus.n87 minus.n72 15.9852
R22503 minus.n26 minus.n11 15.9852
R22504 minus.n46 minus.n45 15.9852
R22505 minus.n115 minus.n62 14.0178
R22506 minus.n78 minus.n77 14.0178
R22507 minus.n17 minus.n16 14.0178
R22508 minus.n54 minus.n1 14.0178
R22509 minus.n122 minus.n60 12.1501
R22510 minus minus.n127 11.8706
R22511 minus.n118 minus.n62 10.575
R22512 minus.n57 minus.n1 10.575
R22513 minus.n120 minus.n119 9.49444
R22514 minus.n59 minus.n58 9.49444
R22515 minus.n108 minus.n107 8.60764
R22516 minus.n84 minus.n72 8.60764
R22517 minus.n23 minus.n11 8.60764
R22518 minus.n47 minus.n46 8.60764
R22519 minus.n100 minus.n68 6.6403
R22520 minus.n95 minus.n94 6.6403
R22521 minus.n34 minus.n33 6.6403
R22522 minus.n39 minus.n7 6.6403
R22523 minus.n127 minus.n126 4.80222
R22524 minus.n102 minus.n66 4.67295
R22525 minus.n90 minus.n89 4.67295
R22526 minus.n29 minus.n28 4.67295
R22527 minus.n41 minus.n5 4.67295
R22528 minus.n113 minus.n112 2.7056
R22529 minus.n82 minus.n74 2.7056
R22530 minus.n21 minus.n13 2.7056
R22531 minus.n52 minus.n51 2.7056
R22532 minus.n127 minus.n122 0.972091
R22533 minus.n126 minus.n125 0.716017
R22534 minus.n121 minus.n61 0.189894
R22535 minus.n117 minus.n61 0.189894
R22536 minus.n117 minus.n116 0.189894
R22537 minus.n116 minus.n63 0.189894
R22538 minus.n111 minus.n63 0.189894
R22539 minus.n111 minus.n110 0.189894
R22540 minus.n110 minus.n109 0.189894
R22541 minus.n109 minus.n65 0.189894
R22542 minus.n104 minus.n65 0.189894
R22543 minus.n104 minus.n103 0.189894
R22544 minus.n103 minus.n67 0.189894
R22545 minus.n99 minus.n67 0.189894
R22546 minus.n99 minus.n98 0.189894
R22547 minus.n98 minus.n69 0.189894
R22548 minus.n93 minus.n69 0.189894
R22549 minus.n93 minus.n92 0.189894
R22550 minus.n92 minus.n91 0.189894
R22551 minus.n91 minus.n71 0.189894
R22552 minus.n86 minus.n71 0.189894
R22553 minus.n86 minus.n85 0.189894
R22554 minus.n85 minus.n73 0.189894
R22555 minus.n81 minus.n73 0.189894
R22556 minus.n81 minus.n80 0.189894
R22557 minus.n80 minus.n75 0.189894
R22558 minus.n19 minus.n14 0.189894
R22559 minus.n20 minus.n19 0.189894
R22560 minus.n20 minus.n12 0.189894
R22561 minus.n24 minus.n12 0.189894
R22562 minus.n25 minus.n24 0.189894
R22563 minus.n25 minus.n10 0.189894
R22564 minus.n30 minus.n10 0.189894
R22565 minus.n31 minus.n30 0.189894
R22566 minus.n32 minus.n31 0.189894
R22567 minus.n32 minus.n8 0.189894
R22568 minus.n37 minus.n8 0.189894
R22569 minus.n38 minus.n37 0.189894
R22570 minus.n38 minus.n6 0.189894
R22571 minus.n42 minus.n6 0.189894
R22572 minus.n43 minus.n42 0.189894
R22573 minus.n43 minus.n4 0.189894
R22574 minus.n48 minus.n4 0.189894
R22575 minus.n49 minus.n48 0.189894
R22576 minus.n50 minus.n49 0.189894
R22577 minus.n50 minus.n2 0.189894
R22578 minus.n55 minus.n2 0.189894
R22579 minus.n56 minus.n55 0.189894
R22580 minus.n56 minus.n0 0.189894
R22581 minus.n60 minus.n0 0.189894
R22582 output.n41 output.n15 289.615
R22583 output.n72 output.n46 289.615
R22584 output.n104 output.n78 289.615
R22585 output.n136 output.n110 289.615
R22586 output.n77 output.n45 197.26
R22587 output.n77 output.n76 196.298
R22588 output.n109 output.n108 196.298
R22589 output.n141 output.n140 196.298
R22590 output.n42 output.n41 185
R22591 output.n40 output.n39 185
R22592 output.n19 output.n18 185
R22593 output.n34 output.n33 185
R22594 output.n32 output.n31 185
R22595 output.n23 output.n22 185
R22596 output.n26 output.n25 185
R22597 output.n73 output.n72 185
R22598 output.n71 output.n70 185
R22599 output.n50 output.n49 185
R22600 output.n65 output.n64 185
R22601 output.n63 output.n62 185
R22602 output.n54 output.n53 185
R22603 output.n57 output.n56 185
R22604 output.n105 output.n104 185
R22605 output.n103 output.n102 185
R22606 output.n82 output.n81 185
R22607 output.n97 output.n96 185
R22608 output.n95 output.n94 185
R22609 output.n86 output.n85 185
R22610 output.n89 output.n88 185
R22611 output.n137 output.n136 185
R22612 output.n135 output.n134 185
R22613 output.n114 output.n113 185
R22614 output.n129 output.n128 185
R22615 output.n127 output.n126 185
R22616 output.n118 output.n117 185
R22617 output.n121 output.n120 185
R22618 output.t3 output.n24 147.661
R22619 output.t1 output.n55 147.661
R22620 output.t2 output.n87 147.661
R22621 output.t0 output.n119 147.661
R22622 output.n41 output.n40 104.615
R22623 output.n40 output.n18 104.615
R22624 output.n33 output.n18 104.615
R22625 output.n33 output.n32 104.615
R22626 output.n32 output.n22 104.615
R22627 output.n25 output.n22 104.615
R22628 output.n72 output.n71 104.615
R22629 output.n71 output.n49 104.615
R22630 output.n64 output.n49 104.615
R22631 output.n64 output.n63 104.615
R22632 output.n63 output.n53 104.615
R22633 output.n56 output.n53 104.615
R22634 output.n104 output.n103 104.615
R22635 output.n103 output.n81 104.615
R22636 output.n96 output.n81 104.615
R22637 output.n96 output.n95 104.615
R22638 output.n95 output.n85 104.615
R22639 output.n88 output.n85 104.615
R22640 output.n136 output.n135 104.615
R22641 output.n135 output.n113 104.615
R22642 output.n128 output.n113 104.615
R22643 output.n128 output.n127 104.615
R22644 output.n127 output.n117 104.615
R22645 output.n120 output.n117 104.615
R22646 output.n1 output.t16 77.056
R22647 output.n14 output.t17 76.6694
R22648 output.n1 output.n0 72.7095
R22649 output.n3 output.n2 72.7095
R22650 output.n5 output.n4 72.7095
R22651 output.n7 output.n6 72.7095
R22652 output.n9 output.n8 72.7095
R22653 output.n11 output.n10 72.7095
R22654 output.n13 output.n12 72.7095
R22655 output.n25 output.t3 52.3082
R22656 output.n56 output.t1 52.3082
R22657 output.n88 output.t2 52.3082
R22658 output.n120 output.t0 52.3082
R22659 output.n26 output.n24 15.6674
R22660 output.n57 output.n55 15.6674
R22661 output.n89 output.n87 15.6674
R22662 output.n121 output.n119 15.6674
R22663 output.n27 output.n23 12.8005
R22664 output.n58 output.n54 12.8005
R22665 output.n90 output.n86 12.8005
R22666 output.n122 output.n118 12.8005
R22667 output.n31 output.n30 12.0247
R22668 output.n62 output.n61 12.0247
R22669 output.n94 output.n93 12.0247
R22670 output.n126 output.n125 12.0247
R22671 output.n34 output.n21 11.249
R22672 output.n65 output.n52 11.249
R22673 output.n97 output.n84 11.249
R22674 output.n129 output.n116 11.249
R22675 output.n35 output.n19 10.4732
R22676 output.n66 output.n50 10.4732
R22677 output.n98 output.n82 10.4732
R22678 output.n130 output.n114 10.4732
R22679 output.n39 output.n38 9.69747
R22680 output.n70 output.n69 9.69747
R22681 output.n102 output.n101 9.69747
R22682 output.n134 output.n133 9.69747
R22683 output.n45 output.n44 9.45567
R22684 output.n76 output.n75 9.45567
R22685 output.n108 output.n107 9.45567
R22686 output.n140 output.n139 9.45567
R22687 output.n44 output.n43 9.3005
R22688 output.n17 output.n16 9.3005
R22689 output.n38 output.n37 9.3005
R22690 output.n36 output.n35 9.3005
R22691 output.n21 output.n20 9.3005
R22692 output.n30 output.n29 9.3005
R22693 output.n28 output.n27 9.3005
R22694 output.n75 output.n74 9.3005
R22695 output.n48 output.n47 9.3005
R22696 output.n69 output.n68 9.3005
R22697 output.n67 output.n66 9.3005
R22698 output.n52 output.n51 9.3005
R22699 output.n61 output.n60 9.3005
R22700 output.n59 output.n58 9.3005
R22701 output.n107 output.n106 9.3005
R22702 output.n80 output.n79 9.3005
R22703 output.n101 output.n100 9.3005
R22704 output.n99 output.n98 9.3005
R22705 output.n84 output.n83 9.3005
R22706 output.n93 output.n92 9.3005
R22707 output.n91 output.n90 9.3005
R22708 output.n139 output.n138 9.3005
R22709 output.n112 output.n111 9.3005
R22710 output.n133 output.n132 9.3005
R22711 output.n131 output.n130 9.3005
R22712 output.n116 output.n115 9.3005
R22713 output.n125 output.n124 9.3005
R22714 output.n123 output.n122 9.3005
R22715 output.n42 output.n17 8.92171
R22716 output.n73 output.n48 8.92171
R22717 output.n105 output.n80 8.92171
R22718 output.n137 output.n112 8.92171
R22719 output output.n141 8.15037
R22720 output.n43 output.n15 8.14595
R22721 output.n74 output.n46 8.14595
R22722 output.n106 output.n78 8.14595
R22723 output.n138 output.n110 8.14595
R22724 output.n45 output.n15 5.81868
R22725 output.n76 output.n46 5.81868
R22726 output.n108 output.n78 5.81868
R22727 output.n140 output.n110 5.81868
R22728 output.n43 output.n42 5.04292
R22729 output.n74 output.n73 5.04292
R22730 output.n106 output.n105 5.04292
R22731 output.n138 output.n137 5.04292
R22732 output.n28 output.n24 4.38594
R22733 output.n59 output.n55 4.38594
R22734 output.n91 output.n87 4.38594
R22735 output.n123 output.n119 4.38594
R22736 output.n39 output.n17 4.26717
R22737 output.n70 output.n48 4.26717
R22738 output.n102 output.n80 4.26717
R22739 output.n134 output.n112 4.26717
R22740 output.n0 output.t5 3.9605
R22741 output.n0 output.t10 3.9605
R22742 output.n2 output.t14 3.9605
R22743 output.n2 output.t6 3.9605
R22744 output.n4 output.t9 3.9605
R22745 output.n4 output.t7 3.9605
R22746 output.n6 output.t13 3.9605
R22747 output.n6 output.t15 3.9605
R22748 output.n8 output.t18 3.9605
R22749 output.n8 output.t11 3.9605
R22750 output.n10 output.t12 3.9605
R22751 output.n10 output.t19 3.9605
R22752 output.n12 output.t4 3.9605
R22753 output.n12 output.t8 3.9605
R22754 output.n38 output.n19 3.49141
R22755 output.n69 output.n50 3.49141
R22756 output.n101 output.n82 3.49141
R22757 output.n133 output.n114 3.49141
R22758 output.n35 output.n34 2.71565
R22759 output.n66 output.n65 2.71565
R22760 output.n98 output.n97 2.71565
R22761 output.n130 output.n129 2.71565
R22762 output.n31 output.n21 1.93989
R22763 output.n62 output.n52 1.93989
R22764 output.n94 output.n84 1.93989
R22765 output.n126 output.n116 1.93989
R22766 output.n30 output.n23 1.16414
R22767 output.n61 output.n54 1.16414
R22768 output.n93 output.n86 1.16414
R22769 output.n125 output.n118 1.16414
R22770 output.n141 output.n109 0.962709
R22771 output.n109 output.n77 0.962709
R22772 output.n27 output.n26 0.388379
R22773 output.n58 output.n57 0.388379
R22774 output.n90 output.n89 0.388379
R22775 output.n122 output.n121 0.388379
R22776 output.n14 output.n13 0.387128
R22777 output.n13 output.n11 0.387128
R22778 output.n11 output.n9 0.387128
R22779 output.n9 output.n7 0.387128
R22780 output.n7 output.n5 0.387128
R22781 output.n5 output.n3 0.387128
R22782 output.n3 output.n1 0.387128
R22783 output.n44 output.n16 0.155672
R22784 output.n37 output.n16 0.155672
R22785 output.n37 output.n36 0.155672
R22786 output.n36 output.n20 0.155672
R22787 output.n29 output.n20 0.155672
R22788 output.n29 output.n28 0.155672
R22789 output.n75 output.n47 0.155672
R22790 output.n68 output.n47 0.155672
R22791 output.n68 output.n67 0.155672
R22792 output.n67 output.n51 0.155672
R22793 output.n60 output.n51 0.155672
R22794 output.n60 output.n59 0.155672
R22795 output.n107 output.n79 0.155672
R22796 output.n100 output.n79 0.155672
R22797 output.n100 output.n99 0.155672
R22798 output.n99 output.n83 0.155672
R22799 output.n92 output.n83 0.155672
R22800 output.n92 output.n91 0.155672
R22801 output.n139 output.n111 0.155672
R22802 output.n132 output.n111 0.155672
R22803 output.n132 output.n131 0.155672
R22804 output.n131 output.n115 0.155672
R22805 output.n124 output.n115 0.155672
R22806 output.n124 output.n123 0.155672
R22807 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 67.66129f
C5 minus diffpairibias 5.39e-19
C6 commonsourceibias output 0.006808f
C7 CSoutput minus 3.03921f
C8 vdd plus 0.072837f
C9 plus diffpairibias 4.4e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.931998f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 45.462303f
C15 minus plus 10.7649f
C16 minus commonsourceibias 0.343793f
C17 plus commonsourceibias 0.290384f
C18 diffpairibias gnd 59.991528f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.181983p
C22 plus gnd 40.3801f
C23 minus gnd 32.59889f
C24 CSoutput gnd 0.11623p
C25 vdd gnd 0.346521p
C26 output.t16 gnd 0.464308f
C27 output.t5 gnd 0.044422f
C28 output.t10 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t14 gnd 0.044422f
C32 output.t6 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t9 gnd 0.044422f
C36 output.t7 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t13 gnd 0.044422f
C40 output.t15 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t18 gnd 0.044422f
C44 output.t11 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t12 gnd 0.044422f
C48 output.t19 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t4 gnd 0.044422f
C52 output.t8 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t17 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t3 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t1 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t2 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t0 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 minus.n0 gnd 0.030269f
C189 minus.t13 gnd 0.508973f
C190 minus.n1 gnd 0.205851f
C191 minus.n2 gnd 0.030269f
C192 minus.t11 gnd 0.508973f
C193 minus.n3 gnd 0.025866f
C194 minus.n4 gnd 0.030269f
C195 minus.t17 gnd 0.508973f
C196 minus.t24 gnd 0.508973f
C197 minus.n5 gnd 0.205851f
C198 minus.n6 gnd 0.030269f
C199 minus.t21 gnd 0.508973f
C200 minus.n7 gnd 0.205851f
C201 minus.n8 gnd 0.030269f
C202 minus.t27 gnd 0.508973f
C203 minus.n9 gnd 0.024602f
C204 minus.n10 gnd 0.030269f
C205 minus.t26 gnd 0.508973f
C206 minus.t5 gnd 0.508973f
C207 minus.n11 gnd 0.205851f
C208 minus.n12 gnd 0.030269f
C209 minus.t9 gnd 0.508973f
C210 minus.n13 gnd 0.205851f
C211 minus.n14 gnd 0.128459f
C212 minus.t14 gnd 0.508973f
C213 minus.t20 gnd 0.569378f
C214 minus.n15 gnd 0.240661f
C215 minus.n16 gnd 0.235738f
C216 minus.n17 gnd 0.038785f
C217 minus.n18 gnd 0.034253f
C218 minus.n19 gnd 0.030269f
C219 minus.n20 gnd 0.030269f
C220 minus.n21 gnd 0.036172f
C221 minus.n22 gnd 0.025866f
C222 minus.n23 gnd 0.039422f
C223 minus.n24 gnd 0.030269f
C224 minus.n25 gnd 0.030269f
C225 minus.n26 gnd 0.037652f
C226 minus.n27 gnd 0.035386f
C227 minus.n28 gnd 0.205851f
C228 minus.n29 gnd 0.037917f
C229 minus.n30 gnd 0.030269f
C230 minus.n31 gnd 0.030269f
C231 minus.n32 gnd 0.030269f
C232 minus.n33 gnd 0.03894f
C233 minus.n34 gnd 0.205851f
C234 minus.n35 gnd 0.036519f
C235 minus.n36 gnd 0.036519f
C236 minus.n37 gnd 0.030269f
C237 minus.n38 gnd 0.030269f
C238 minus.n39 gnd 0.03894f
C239 minus.n40 gnd 0.024602f
C240 minus.n41 gnd 0.037917f
C241 minus.n42 gnd 0.030269f
C242 minus.n43 gnd 0.030269f
C243 minus.n44 gnd 0.035386f
C244 minus.n45 gnd 0.037652f
C245 minus.n46 gnd 0.205851f
C246 minus.n47 gnd 0.039422f
C247 minus.n48 gnd 0.030269f
C248 minus.n49 gnd 0.030269f
C249 minus.n50 gnd 0.030269f
C250 minus.n51 gnd 0.036172f
C251 minus.n52 gnd 0.205851f
C252 minus.n53 gnd 0.034253f
C253 minus.n54 gnd 0.038785f
C254 minus.n55 gnd 0.030269f
C255 minus.n56 gnd 0.030269f
C256 minus.n57 gnd 0.039487f
C257 minus.n58 gnd 0.011001f
C258 minus.t10 gnd 0.550454f
C259 minus.n59 gnd 0.238341f
C260 minus.n60 gnd 0.354592f
C261 minus.n61 gnd 0.030269f
C262 minus.t8 gnd 0.550454f
C263 minus.t12 gnd 0.508973f
C264 minus.n62 gnd 0.205851f
C265 minus.n63 gnd 0.030269f
C266 minus.t18 gnd 0.508973f
C267 minus.n64 gnd 0.025866f
C268 minus.n65 gnd 0.030269f
C269 minus.t25 gnd 0.508973f
C270 minus.t22 gnd 0.508973f
C271 minus.n66 gnd 0.205851f
C272 minus.n67 gnd 0.030269f
C273 minus.t19 gnd 0.508973f
C274 minus.n68 gnd 0.205851f
C275 minus.n69 gnd 0.030269f
C276 minus.t7 gnd 0.508973f
C277 minus.n70 gnd 0.024602f
C278 minus.n71 gnd 0.030269f
C279 minus.t6 gnd 0.508973f
C280 minus.t16 gnd 0.508973f
C281 minus.n72 gnd 0.205851f
C282 minus.n73 gnd 0.030269f
C283 minus.t15 gnd 0.508973f
C284 minus.n74 gnd 0.205851f
C285 minus.n75 gnd 0.128459f
C286 minus.t23 gnd 0.508973f
C287 minus.t28 gnd 0.569378f
C288 minus.n76 gnd 0.240661f
C289 minus.n77 gnd 0.235738f
C290 minus.n78 gnd 0.038785f
C291 minus.n79 gnd 0.034253f
C292 minus.n80 gnd 0.030269f
C293 minus.n81 gnd 0.030269f
C294 minus.n82 gnd 0.036172f
C295 minus.n83 gnd 0.025866f
C296 minus.n84 gnd 0.039422f
C297 minus.n85 gnd 0.030269f
C298 minus.n86 gnd 0.030269f
C299 minus.n87 gnd 0.037652f
C300 minus.n88 gnd 0.035386f
C301 minus.n89 gnd 0.205851f
C302 minus.n90 gnd 0.037917f
C303 minus.n91 gnd 0.030269f
C304 minus.n92 gnd 0.030269f
C305 minus.n93 gnd 0.030269f
C306 minus.n94 gnd 0.03894f
C307 minus.n95 gnd 0.205851f
C308 minus.n96 gnd 0.036519f
C309 minus.n97 gnd 0.036519f
C310 minus.n98 gnd 0.030269f
C311 minus.n99 gnd 0.030269f
C312 minus.n100 gnd 0.03894f
C313 minus.n101 gnd 0.024602f
C314 minus.n102 gnd 0.037917f
C315 minus.n103 gnd 0.030269f
C316 minus.n104 gnd 0.030269f
C317 minus.n105 gnd 0.035386f
C318 minus.n106 gnd 0.037652f
C319 minus.n107 gnd 0.205851f
C320 minus.n108 gnd 0.039422f
C321 minus.n109 gnd 0.030269f
C322 minus.n110 gnd 0.030269f
C323 minus.n111 gnd 0.030269f
C324 minus.n112 gnd 0.036172f
C325 minus.n113 gnd 0.205851f
C326 minus.n114 gnd 0.034253f
C327 minus.n115 gnd 0.038785f
C328 minus.n116 gnd 0.030269f
C329 minus.n117 gnd 0.030269f
C330 minus.n118 gnd 0.039487f
C331 minus.n119 gnd 0.011001f
C332 minus.n120 gnd 0.238341f
C333 minus.n121 gnd 1.10421f
C334 minus.n122 gnd 1.622f
C335 minus.t4 gnd 0.009331f
C336 minus.t3 gnd 0.009331f
C337 minus.n123 gnd 0.030683f
C338 minus.t0 gnd 0.009331f
C339 minus.t2 gnd 0.009331f
C340 minus.n124 gnd 0.030263f
C341 minus.n125 gnd 0.258277f
C342 minus.t1 gnd 0.051936f
C343 minus.n126 gnd 0.140939f
C344 minus.n127 gnd 2.12621f
C345 diffpairibias.t27 gnd 0.090128f
C346 diffpairibias.t23 gnd 0.08996f
C347 diffpairibias.n0 gnd 0.105991f
C348 diffpairibias.t28 gnd 0.08996f
C349 diffpairibias.n1 gnd 0.051736f
C350 diffpairibias.t25 gnd 0.08996f
C351 diffpairibias.n2 gnd 0.051736f
C352 diffpairibias.t29 gnd 0.08996f
C353 diffpairibias.n3 gnd 0.041084f
C354 diffpairibias.t15 gnd 0.086371f
C355 diffpairibias.t1 gnd 0.085993f
C356 diffpairibias.n4 gnd 0.13579f
C357 diffpairibias.t11 gnd 0.085993f
C358 diffpairibias.n5 gnd 0.072463f
C359 diffpairibias.t13 gnd 0.085993f
C360 diffpairibias.n6 gnd 0.072463f
C361 diffpairibias.t7 gnd 0.085993f
C362 diffpairibias.n7 gnd 0.072463f
C363 diffpairibias.t3 gnd 0.085993f
C364 diffpairibias.n8 gnd 0.072463f
C365 diffpairibias.t17 gnd 0.085993f
C366 diffpairibias.n9 gnd 0.072463f
C367 diffpairibias.t5 gnd 0.085993f
C368 diffpairibias.n10 gnd 0.072463f
C369 diffpairibias.t19 gnd 0.085993f
C370 diffpairibias.n11 gnd 0.072463f
C371 diffpairibias.t9 gnd 0.085993f
C372 diffpairibias.n12 gnd 0.102883f
C373 diffpairibias.t14 gnd 0.086899f
C374 diffpairibias.t0 gnd 0.086748f
C375 diffpairibias.n13 gnd 0.094648f
C376 diffpairibias.t10 gnd 0.086748f
C377 diffpairibias.n14 gnd 0.052262f
C378 diffpairibias.t12 gnd 0.086748f
C379 diffpairibias.n15 gnd 0.052262f
C380 diffpairibias.t6 gnd 0.086748f
C381 diffpairibias.n16 gnd 0.052262f
C382 diffpairibias.t2 gnd 0.086748f
C383 diffpairibias.n17 gnd 0.052262f
C384 diffpairibias.t16 gnd 0.086748f
C385 diffpairibias.n18 gnd 0.052262f
C386 diffpairibias.t4 gnd 0.086748f
C387 diffpairibias.n19 gnd 0.052262f
C388 diffpairibias.t18 gnd 0.086748f
C389 diffpairibias.n20 gnd 0.052262f
C390 diffpairibias.t8 gnd 0.086748f
C391 diffpairibias.n21 gnd 0.061849f
C392 diffpairibias.n22 gnd 0.233513f
C393 diffpairibias.t20 gnd 0.08996f
C394 diffpairibias.n23 gnd 0.051747f
C395 diffpairibias.t26 gnd 0.08996f
C396 diffpairibias.n24 gnd 0.051736f
C397 diffpairibias.t22 gnd 0.08996f
C398 diffpairibias.n25 gnd 0.051736f
C399 diffpairibias.t21 gnd 0.08996f
C400 diffpairibias.n26 gnd 0.051736f
C401 diffpairibias.t24 gnd 0.08996f
C402 diffpairibias.n27 gnd 0.04729f
C403 diffpairibias.n28 gnd 0.047711f
C404 commonsourceibias.n0 gnd 0.010724f
C405 commonsourceibias.t115 gnd 0.162395f
C406 commonsourceibias.t136 gnd 0.150157f
C407 commonsourceibias.n1 gnd 0.007823f
C408 commonsourceibias.n2 gnd 0.008037f
C409 commonsourceibias.t151 gnd 0.150157f
C410 commonsourceibias.n3 gnd 0.01034f
C411 commonsourceibias.n4 gnd 0.008037f
C412 commonsourceibias.t104 gnd 0.150157f
C413 commonsourceibias.n5 gnd 0.059912f
C414 commonsourceibias.t126 gnd 0.150157f
C415 commonsourceibias.n6 gnd 0.007578f
C416 commonsourceibias.n7 gnd 0.008037f
C417 commonsourceibias.t144 gnd 0.150157f
C418 commonsourceibias.n8 gnd 0.010186f
C419 commonsourceibias.n9 gnd 0.008037f
C420 commonsourceibias.t96 gnd 0.150157f
C421 commonsourceibias.n10 gnd 0.059912f
C422 commonsourceibias.t94 gnd 0.150157f
C423 commonsourceibias.n11 gnd 0.007361f
C424 commonsourceibias.n12 gnd 0.008037f
C425 commonsourceibias.t134 gnd 0.150157f
C426 commonsourceibias.n13 gnd 0.010015f
C427 commonsourceibias.n14 gnd 0.010724f
C428 commonsourceibias.t74 gnd 0.162395f
C429 commonsourceibias.t20 gnd 0.150157f
C430 commonsourceibias.n15 gnd 0.007823f
C431 commonsourceibias.n16 gnd 0.008037f
C432 commonsourceibias.t50 gnd 0.150157f
C433 commonsourceibias.n17 gnd 0.01034f
C434 commonsourceibias.n18 gnd 0.008037f
C435 commonsourceibias.t8 gnd 0.150157f
C436 commonsourceibias.n19 gnd 0.059912f
C437 commonsourceibias.t36 gnd 0.150157f
C438 commonsourceibias.n20 gnd 0.007578f
C439 commonsourceibias.n21 gnd 0.008037f
C440 commonsourceibias.t76 gnd 0.150157f
C441 commonsourceibias.n22 gnd 0.010186f
C442 commonsourceibias.n23 gnd 0.008037f
C443 commonsourceibias.t24 gnd 0.150157f
C444 commonsourceibias.n24 gnd 0.059912f
C445 commonsourceibias.t34 gnd 0.150157f
C446 commonsourceibias.n25 gnd 0.007361f
C447 commonsourceibias.n26 gnd 0.008037f
C448 commonsourceibias.t10 gnd 0.150157f
C449 commonsourceibias.n27 gnd 0.010015f
C450 commonsourceibias.n28 gnd 0.008037f
C451 commonsourceibias.t40 gnd 0.150157f
C452 commonsourceibias.n29 gnd 0.059912f
C453 commonsourceibias.t56 gnd 0.150157f
C454 commonsourceibias.n30 gnd 0.007172f
C455 commonsourceibias.n31 gnd 0.008037f
C456 commonsourceibias.t26 gnd 0.150157f
C457 commonsourceibias.n32 gnd 0.009825f
C458 commonsourceibias.n33 gnd 0.008037f
C459 commonsourceibias.t38 gnd 0.150157f
C460 commonsourceibias.n34 gnd 0.059912f
C461 commonsourceibias.t70 gnd 0.150157f
C462 commonsourceibias.n35 gnd 0.007008f
C463 commonsourceibias.n36 gnd 0.008037f
C464 commonsourceibias.t18 gnd 0.150157f
C465 commonsourceibias.n37 gnd 0.009613f
C466 commonsourceibias.n38 gnd 0.008037f
C467 commonsourceibias.t22 gnd 0.150157f
C468 commonsourceibias.n39 gnd 0.059912f
C469 commonsourceibias.t52 gnd 0.150157f
C470 commonsourceibias.n40 gnd 0.006868f
C471 commonsourceibias.n41 gnd 0.008037f
C472 commonsourceibias.t4 gnd 0.150157f
C473 commonsourceibias.n42 gnd 0.009378f
C474 commonsourceibias.t78 gnd 0.166947f
C475 commonsourceibias.t46 gnd 0.150157f
C476 commonsourceibias.n43 gnd 0.065449f
C477 commonsourceibias.n44 gnd 0.071822f
C478 commonsourceibias.n45 gnd 0.033327f
C479 commonsourceibias.n46 gnd 0.008037f
C480 commonsourceibias.n47 gnd 0.007823f
C481 commonsourceibias.n48 gnd 0.01121f
C482 commonsourceibias.n49 gnd 0.059912f
C483 commonsourceibias.n50 gnd 0.011203f
C484 commonsourceibias.n51 gnd 0.008037f
C485 commonsourceibias.n52 gnd 0.008037f
C486 commonsourceibias.n53 gnd 0.008037f
C487 commonsourceibias.n54 gnd 0.01034f
C488 commonsourceibias.n55 gnd 0.059912f
C489 commonsourceibias.n56 gnd 0.010583f
C490 commonsourceibias.n57 gnd 0.010282f
C491 commonsourceibias.n58 gnd 0.008037f
C492 commonsourceibias.n59 gnd 0.008037f
C493 commonsourceibias.n60 gnd 0.008037f
C494 commonsourceibias.n61 gnd 0.007578f
C495 commonsourceibias.n62 gnd 0.01122f
C496 commonsourceibias.n63 gnd 0.059912f
C497 commonsourceibias.n64 gnd 0.011217f
C498 commonsourceibias.n65 gnd 0.008037f
C499 commonsourceibias.n66 gnd 0.008037f
C500 commonsourceibias.n67 gnd 0.008037f
C501 commonsourceibias.n68 gnd 0.010186f
C502 commonsourceibias.n69 gnd 0.059912f
C503 commonsourceibias.n70 gnd 0.010507f
C504 commonsourceibias.n71 gnd 0.010357f
C505 commonsourceibias.n72 gnd 0.008037f
C506 commonsourceibias.n73 gnd 0.008037f
C507 commonsourceibias.n74 gnd 0.008037f
C508 commonsourceibias.n75 gnd 0.007361f
C509 commonsourceibias.n76 gnd 0.011225f
C510 commonsourceibias.n77 gnd 0.059912f
C511 commonsourceibias.n78 gnd 0.011224f
C512 commonsourceibias.n79 gnd 0.008037f
C513 commonsourceibias.n80 gnd 0.008037f
C514 commonsourceibias.n81 gnd 0.008037f
C515 commonsourceibias.n82 gnd 0.010015f
C516 commonsourceibias.n83 gnd 0.059912f
C517 commonsourceibias.n84 gnd 0.010432f
C518 commonsourceibias.n85 gnd 0.010432f
C519 commonsourceibias.n86 gnd 0.008037f
C520 commonsourceibias.n87 gnd 0.008037f
C521 commonsourceibias.n88 gnd 0.008037f
C522 commonsourceibias.n89 gnd 0.007172f
C523 commonsourceibias.n90 gnd 0.011224f
C524 commonsourceibias.n91 gnd 0.059912f
C525 commonsourceibias.n92 gnd 0.011225f
C526 commonsourceibias.n93 gnd 0.008037f
C527 commonsourceibias.n94 gnd 0.008037f
C528 commonsourceibias.n95 gnd 0.008037f
C529 commonsourceibias.n96 gnd 0.009825f
C530 commonsourceibias.n97 gnd 0.059912f
C531 commonsourceibias.n98 gnd 0.010357f
C532 commonsourceibias.n99 gnd 0.010507f
C533 commonsourceibias.n100 gnd 0.008037f
C534 commonsourceibias.n101 gnd 0.008037f
C535 commonsourceibias.n102 gnd 0.008037f
C536 commonsourceibias.n103 gnd 0.007008f
C537 commonsourceibias.n104 gnd 0.011217f
C538 commonsourceibias.n105 gnd 0.059912f
C539 commonsourceibias.n106 gnd 0.01122f
C540 commonsourceibias.n107 gnd 0.008037f
C541 commonsourceibias.n108 gnd 0.008037f
C542 commonsourceibias.n109 gnd 0.008037f
C543 commonsourceibias.n110 gnd 0.009613f
C544 commonsourceibias.n111 gnd 0.059912f
C545 commonsourceibias.n112 gnd 0.010282f
C546 commonsourceibias.n113 gnd 0.010583f
C547 commonsourceibias.n114 gnd 0.008037f
C548 commonsourceibias.n115 gnd 0.008037f
C549 commonsourceibias.n116 gnd 0.008037f
C550 commonsourceibias.n117 gnd 0.006868f
C551 commonsourceibias.n118 gnd 0.011203f
C552 commonsourceibias.n119 gnd 0.059912f
C553 commonsourceibias.n120 gnd 0.01121f
C554 commonsourceibias.n121 gnd 0.008037f
C555 commonsourceibias.n122 gnd 0.008037f
C556 commonsourceibias.n123 gnd 0.008037f
C557 commonsourceibias.n124 gnd 0.009378f
C558 commonsourceibias.n125 gnd 0.059912f
C559 commonsourceibias.n126 gnd 0.009861f
C560 commonsourceibias.n127 gnd 0.07189f
C561 commonsourceibias.n128 gnd 0.080075f
C562 commonsourceibias.t75 gnd 0.017343f
C563 commonsourceibias.t21 gnd 0.017343f
C564 commonsourceibias.n129 gnd 0.15325f
C565 commonsourceibias.n130 gnd 0.132562f
C566 commonsourceibias.t51 gnd 0.017343f
C567 commonsourceibias.t9 gnd 0.017343f
C568 commonsourceibias.n131 gnd 0.15325f
C569 commonsourceibias.n132 gnd 0.070394f
C570 commonsourceibias.t37 gnd 0.017343f
C571 commonsourceibias.t77 gnd 0.017343f
C572 commonsourceibias.n133 gnd 0.15325f
C573 commonsourceibias.n134 gnd 0.070394f
C574 commonsourceibias.t25 gnd 0.017343f
C575 commonsourceibias.t35 gnd 0.017343f
C576 commonsourceibias.n135 gnd 0.15325f
C577 commonsourceibias.n136 gnd 0.070394f
C578 commonsourceibias.t11 gnd 0.017343f
C579 commonsourceibias.t41 gnd 0.017343f
C580 commonsourceibias.n137 gnd 0.15325f
C581 commonsourceibias.n138 gnd 0.058811f
C582 commonsourceibias.t47 gnd 0.017343f
C583 commonsourceibias.t79 gnd 0.017343f
C584 commonsourceibias.n139 gnd 0.153763f
C585 commonsourceibias.t53 gnd 0.017343f
C586 commonsourceibias.t5 gnd 0.017343f
C587 commonsourceibias.n140 gnd 0.15325f
C588 commonsourceibias.n141 gnd 0.1428f
C589 commonsourceibias.t19 gnd 0.017343f
C590 commonsourceibias.t23 gnd 0.017343f
C591 commonsourceibias.n142 gnd 0.15325f
C592 commonsourceibias.n143 gnd 0.070394f
C593 commonsourceibias.t39 gnd 0.017343f
C594 commonsourceibias.t71 gnd 0.017343f
C595 commonsourceibias.n144 gnd 0.15325f
C596 commonsourceibias.n145 gnd 0.070394f
C597 commonsourceibias.t57 gnd 0.017343f
C598 commonsourceibias.t27 gnd 0.017343f
C599 commonsourceibias.n146 gnd 0.15325f
C600 commonsourceibias.n147 gnd 0.058811f
C601 commonsourceibias.n148 gnd 0.071213f
C602 commonsourceibias.n149 gnd 0.052016f
C603 commonsourceibias.t152 gnd 0.150157f
C604 commonsourceibias.n150 gnd 0.059912f
C605 commonsourceibias.t88 gnd 0.150157f
C606 commonsourceibias.n151 gnd 0.059912f
C607 commonsourceibias.n152 gnd 0.008037f
C608 commonsourceibias.t124 gnd 0.150157f
C609 commonsourceibias.n153 gnd 0.059912f
C610 commonsourceibias.n154 gnd 0.008037f
C611 commonsourceibias.t120 gnd 0.150157f
C612 commonsourceibias.n155 gnd 0.059912f
C613 commonsourceibias.n156 gnd 0.008037f
C614 commonsourceibias.t139 gnd 0.150157f
C615 commonsourceibias.n157 gnd 0.007008f
C616 commonsourceibias.n158 gnd 0.008037f
C617 commonsourceibias.t112 gnd 0.150157f
C618 commonsourceibias.n159 gnd 0.009613f
C619 commonsourceibias.n160 gnd 0.008037f
C620 commonsourceibias.t106 gnd 0.150157f
C621 commonsourceibias.n161 gnd 0.059912f
C622 commonsourceibias.t128 gnd 0.150157f
C623 commonsourceibias.n162 gnd 0.006868f
C624 commonsourceibias.n163 gnd 0.008037f
C625 commonsourceibias.t145 gnd 0.150157f
C626 commonsourceibias.n164 gnd 0.009378f
C627 commonsourceibias.t118 gnd 0.166947f
C628 commonsourceibias.t99 gnd 0.150157f
C629 commonsourceibias.n165 gnd 0.065449f
C630 commonsourceibias.n166 gnd 0.071822f
C631 commonsourceibias.n167 gnd 0.033327f
C632 commonsourceibias.n168 gnd 0.008037f
C633 commonsourceibias.n169 gnd 0.007823f
C634 commonsourceibias.n170 gnd 0.01121f
C635 commonsourceibias.n171 gnd 0.059912f
C636 commonsourceibias.n172 gnd 0.011203f
C637 commonsourceibias.n173 gnd 0.008037f
C638 commonsourceibias.n174 gnd 0.008037f
C639 commonsourceibias.n175 gnd 0.008037f
C640 commonsourceibias.n176 gnd 0.01034f
C641 commonsourceibias.n177 gnd 0.059912f
C642 commonsourceibias.n178 gnd 0.010583f
C643 commonsourceibias.n179 gnd 0.010282f
C644 commonsourceibias.n180 gnd 0.008037f
C645 commonsourceibias.n181 gnd 0.008037f
C646 commonsourceibias.n182 gnd 0.008037f
C647 commonsourceibias.n183 gnd 0.007578f
C648 commonsourceibias.n184 gnd 0.01122f
C649 commonsourceibias.n185 gnd 0.059912f
C650 commonsourceibias.n186 gnd 0.011217f
C651 commonsourceibias.n187 gnd 0.008037f
C652 commonsourceibias.n188 gnd 0.008037f
C653 commonsourceibias.n189 gnd 0.008037f
C654 commonsourceibias.n190 gnd 0.010186f
C655 commonsourceibias.n191 gnd 0.059912f
C656 commonsourceibias.n192 gnd 0.010507f
C657 commonsourceibias.n193 gnd 0.010357f
C658 commonsourceibias.n194 gnd 0.008037f
C659 commonsourceibias.n195 gnd 0.008037f
C660 commonsourceibias.n196 gnd 0.009825f
C661 commonsourceibias.n197 gnd 0.007361f
C662 commonsourceibias.n198 gnd 0.011225f
C663 commonsourceibias.n199 gnd 0.008037f
C664 commonsourceibias.n200 gnd 0.008037f
C665 commonsourceibias.n201 gnd 0.011224f
C666 commonsourceibias.n202 gnd 0.007172f
C667 commonsourceibias.n203 gnd 0.010015f
C668 commonsourceibias.n204 gnd 0.008037f
C669 commonsourceibias.n205 gnd 0.007021f
C670 commonsourceibias.n206 gnd 0.010432f
C671 commonsourceibias.n207 gnd 0.010432f
C672 commonsourceibias.n208 gnd 0.007021f
C673 commonsourceibias.n209 gnd 0.008037f
C674 commonsourceibias.n210 gnd 0.008037f
C675 commonsourceibias.n211 gnd 0.007172f
C676 commonsourceibias.n212 gnd 0.011224f
C677 commonsourceibias.n213 gnd 0.059912f
C678 commonsourceibias.n214 gnd 0.011225f
C679 commonsourceibias.n215 gnd 0.008037f
C680 commonsourceibias.n216 gnd 0.008037f
C681 commonsourceibias.n217 gnd 0.008037f
C682 commonsourceibias.n218 gnd 0.009825f
C683 commonsourceibias.n219 gnd 0.059912f
C684 commonsourceibias.n220 gnd 0.010357f
C685 commonsourceibias.n221 gnd 0.010507f
C686 commonsourceibias.n222 gnd 0.008037f
C687 commonsourceibias.n223 gnd 0.008037f
C688 commonsourceibias.n224 gnd 0.008037f
C689 commonsourceibias.n225 gnd 0.007008f
C690 commonsourceibias.n226 gnd 0.011217f
C691 commonsourceibias.n227 gnd 0.059912f
C692 commonsourceibias.n228 gnd 0.01122f
C693 commonsourceibias.n229 gnd 0.008037f
C694 commonsourceibias.n230 gnd 0.008037f
C695 commonsourceibias.n231 gnd 0.008037f
C696 commonsourceibias.n232 gnd 0.009613f
C697 commonsourceibias.n233 gnd 0.059912f
C698 commonsourceibias.n234 gnd 0.010282f
C699 commonsourceibias.n235 gnd 0.010583f
C700 commonsourceibias.n236 gnd 0.008037f
C701 commonsourceibias.n237 gnd 0.008037f
C702 commonsourceibias.n238 gnd 0.008037f
C703 commonsourceibias.n239 gnd 0.006868f
C704 commonsourceibias.n240 gnd 0.011203f
C705 commonsourceibias.n241 gnd 0.059912f
C706 commonsourceibias.n242 gnd 0.01121f
C707 commonsourceibias.n243 gnd 0.008037f
C708 commonsourceibias.n244 gnd 0.008037f
C709 commonsourceibias.n245 gnd 0.008037f
C710 commonsourceibias.n246 gnd 0.009378f
C711 commonsourceibias.n247 gnd 0.059912f
C712 commonsourceibias.n248 gnd 0.009861f
C713 commonsourceibias.n249 gnd 0.07189f
C714 commonsourceibias.n250 gnd 0.04697f
C715 commonsourceibias.n251 gnd 0.010724f
C716 commonsourceibias.t119 gnd 0.150157f
C717 commonsourceibias.n252 gnd 0.007823f
C718 commonsourceibias.n253 gnd 0.008037f
C719 commonsourceibias.t137 gnd 0.150157f
C720 commonsourceibias.n254 gnd 0.01034f
C721 commonsourceibias.n255 gnd 0.008037f
C722 commonsourceibias.t91 gnd 0.150157f
C723 commonsourceibias.n256 gnd 0.059912f
C724 commonsourceibias.t109 gnd 0.150157f
C725 commonsourceibias.n257 gnd 0.007578f
C726 commonsourceibias.n258 gnd 0.008037f
C727 commonsourceibias.t127 gnd 0.150157f
C728 commonsourceibias.n259 gnd 0.010186f
C729 commonsourceibias.n260 gnd 0.008037f
C730 commonsourceibias.t86 gnd 0.150157f
C731 commonsourceibias.n261 gnd 0.059912f
C732 commonsourceibias.t83 gnd 0.150157f
C733 commonsourceibias.n262 gnd 0.007361f
C734 commonsourceibias.n263 gnd 0.008037f
C735 commonsourceibias.t117 gnd 0.150157f
C736 commonsourceibias.n264 gnd 0.010015f
C737 commonsourceibias.n265 gnd 0.008037f
C738 commonsourceibias.t138 gnd 0.150157f
C739 commonsourceibias.n266 gnd 0.059912f
C740 commonsourceibias.t159 gnd 0.150157f
C741 commonsourceibias.n267 gnd 0.007172f
C742 commonsourceibias.n268 gnd 0.008037f
C743 commonsourceibias.t108 gnd 0.150157f
C744 commonsourceibias.n269 gnd 0.009825f
C745 commonsourceibias.n270 gnd 0.008037f
C746 commonsourceibias.t102 gnd 0.150157f
C747 commonsourceibias.n271 gnd 0.059912f
C748 commonsourceibias.t121 gnd 0.150157f
C749 commonsourceibias.n272 gnd 0.007008f
C750 commonsourceibias.n273 gnd 0.008037f
C751 commonsourceibias.t95 gnd 0.150157f
C752 commonsourceibias.n274 gnd 0.009613f
C753 commonsourceibias.n275 gnd 0.008037f
C754 commonsourceibias.t93 gnd 0.150157f
C755 commonsourceibias.n276 gnd 0.059912f
C756 commonsourceibias.t110 gnd 0.150157f
C757 commonsourceibias.n277 gnd 0.006868f
C758 commonsourceibias.n278 gnd 0.008037f
C759 commonsourceibias.t129 gnd 0.150157f
C760 commonsourceibias.n279 gnd 0.009378f
C761 commonsourceibias.t101 gnd 0.166947f
C762 commonsourceibias.t87 gnd 0.150157f
C763 commonsourceibias.n280 gnd 0.065449f
C764 commonsourceibias.n281 gnd 0.071822f
C765 commonsourceibias.n282 gnd 0.033327f
C766 commonsourceibias.n283 gnd 0.008037f
C767 commonsourceibias.n284 gnd 0.007823f
C768 commonsourceibias.n285 gnd 0.01121f
C769 commonsourceibias.n286 gnd 0.059912f
C770 commonsourceibias.n287 gnd 0.011203f
C771 commonsourceibias.n288 gnd 0.008037f
C772 commonsourceibias.n289 gnd 0.008037f
C773 commonsourceibias.n290 gnd 0.008037f
C774 commonsourceibias.n291 gnd 0.01034f
C775 commonsourceibias.n292 gnd 0.059912f
C776 commonsourceibias.n293 gnd 0.010583f
C777 commonsourceibias.n294 gnd 0.010282f
C778 commonsourceibias.n295 gnd 0.008037f
C779 commonsourceibias.n296 gnd 0.008037f
C780 commonsourceibias.n297 gnd 0.008037f
C781 commonsourceibias.n298 gnd 0.007578f
C782 commonsourceibias.n299 gnd 0.01122f
C783 commonsourceibias.n300 gnd 0.059912f
C784 commonsourceibias.n301 gnd 0.011217f
C785 commonsourceibias.n302 gnd 0.008037f
C786 commonsourceibias.n303 gnd 0.008037f
C787 commonsourceibias.n304 gnd 0.008037f
C788 commonsourceibias.n305 gnd 0.010186f
C789 commonsourceibias.n306 gnd 0.059912f
C790 commonsourceibias.n307 gnd 0.010507f
C791 commonsourceibias.n308 gnd 0.010357f
C792 commonsourceibias.n309 gnd 0.008037f
C793 commonsourceibias.n310 gnd 0.008037f
C794 commonsourceibias.n311 gnd 0.008037f
C795 commonsourceibias.n312 gnd 0.007361f
C796 commonsourceibias.n313 gnd 0.011225f
C797 commonsourceibias.n314 gnd 0.059912f
C798 commonsourceibias.n315 gnd 0.011224f
C799 commonsourceibias.n316 gnd 0.008037f
C800 commonsourceibias.n317 gnd 0.008037f
C801 commonsourceibias.n318 gnd 0.008037f
C802 commonsourceibias.n319 gnd 0.010015f
C803 commonsourceibias.n320 gnd 0.059912f
C804 commonsourceibias.n321 gnd 0.010432f
C805 commonsourceibias.n322 gnd 0.010432f
C806 commonsourceibias.n323 gnd 0.008037f
C807 commonsourceibias.n324 gnd 0.008037f
C808 commonsourceibias.n325 gnd 0.008037f
C809 commonsourceibias.n326 gnd 0.007172f
C810 commonsourceibias.n327 gnd 0.011224f
C811 commonsourceibias.n328 gnd 0.059912f
C812 commonsourceibias.n329 gnd 0.011225f
C813 commonsourceibias.n330 gnd 0.008037f
C814 commonsourceibias.n331 gnd 0.008037f
C815 commonsourceibias.n332 gnd 0.008037f
C816 commonsourceibias.n333 gnd 0.009825f
C817 commonsourceibias.n334 gnd 0.059912f
C818 commonsourceibias.n335 gnd 0.010357f
C819 commonsourceibias.n336 gnd 0.010507f
C820 commonsourceibias.n337 gnd 0.008037f
C821 commonsourceibias.n338 gnd 0.008037f
C822 commonsourceibias.n339 gnd 0.008037f
C823 commonsourceibias.n340 gnd 0.007008f
C824 commonsourceibias.n341 gnd 0.011217f
C825 commonsourceibias.n342 gnd 0.059912f
C826 commonsourceibias.n343 gnd 0.01122f
C827 commonsourceibias.n344 gnd 0.008037f
C828 commonsourceibias.n345 gnd 0.008037f
C829 commonsourceibias.n346 gnd 0.008037f
C830 commonsourceibias.n347 gnd 0.009613f
C831 commonsourceibias.n348 gnd 0.059912f
C832 commonsourceibias.n349 gnd 0.010282f
C833 commonsourceibias.n350 gnd 0.010583f
C834 commonsourceibias.n351 gnd 0.008037f
C835 commonsourceibias.n352 gnd 0.008037f
C836 commonsourceibias.n353 gnd 0.008037f
C837 commonsourceibias.n354 gnd 0.006868f
C838 commonsourceibias.n355 gnd 0.011203f
C839 commonsourceibias.n356 gnd 0.059912f
C840 commonsourceibias.n357 gnd 0.01121f
C841 commonsourceibias.n358 gnd 0.008037f
C842 commonsourceibias.n359 gnd 0.008037f
C843 commonsourceibias.n360 gnd 0.008037f
C844 commonsourceibias.n361 gnd 0.009378f
C845 commonsourceibias.n362 gnd 0.059912f
C846 commonsourceibias.n363 gnd 0.009861f
C847 commonsourceibias.t100 gnd 0.162395f
C848 commonsourceibias.n364 gnd 0.07189f
C849 commonsourceibias.n365 gnd 0.025003f
C850 commonsourceibias.n366 gnd 0.464917f
C851 commonsourceibias.n367 gnd 0.010724f
C852 commonsourceibias.t140 gnd 0.162395f
C853 commonsourceibias.t154 gnd 0.150157f
C854 commonsourceibias.n368 gnd 0.007823f
C855 commonsourceibias.n369 gnd 0.008037f
C856 commonsourceibias.t84 gnd 0.150157f
C857 commonsourceibias.n370 gnd 0.01034f
C858 commonsourceibias.n371 gnd 0.008037f
C859 commonsourceibias.t147 gnd 0.150157f
C860 commonsourceibias.n372 gnd 0.007578f
C861 commonsourceibias.n373 gnd 0.008037f
C862 commonsourceibias.t80 gnd 0.150157f
C863 commonsourceibias.n374 gnd 0.010186f
C864 commonsourceibias.n375 gnd 0.008037f
C865 commonsourceibias.t114 gnd 0.150157f
C866 commonsourceibias.n376 gnd 0.007361f
C867 commonsourceibias.n377 gnd 0.008037f
C868 commonsourceibias.t155 gnd 0.150157f
C869 commonsourceibias.n378 gnd 0.010015f
C870 commonsourceibias.t31 gnd 0.017343f
C871 commonsourceibias.t3 gnd 0.017343f
C872 commonsourceibias.n379 gnd 0.153763f
C873 commonsourceibias.t49 gnd 0.017343f
C874 commonsourceibias.t15 gnd 0.017343f
C875 commonsourceibias.n380 gnd 0.15325f
C876 commonsourceibias.n381 gnd 0.1428f
C877 commonsourceibias.t69 gnd 0.017343f
C878 commonsourceibias.t67 gnd 0.017343f
C879 commonsourceibias.n382 gnd 0.15325f
C880 commonsourceibias.n383 gnd 0.070394f
C881 commonsourceibias.t7 gnd 0.017343f
C882 commonsourceibias.t63 gnd 0.017343f
C883 commonsourceibias.n384 gnd 0.15325f
C884 commonsourceibias.n385 gnd 0.070394f
C885 commonsourceibias.t55 gnd 0.017343f
C886 commonsourceibias.t73 gnd 0.017343f
C887 commonsourceibias.n386 gnd 0.15325f
C888 commonsourceibias.n387 gnd 0.058811f
C889 commonsourceibias.n388 gnd 0.010724f
C890 commonsourceibias.t42 gnd 0.150157f
C891 commonsourceibias.n389 gnd 0.007823f
C892 commonsourceibias.n390 gnd 0.008037f
C893 commonsourceibias.t0 gnd 0.150157f
C894 commonsourceibias.n391 gnd 0.01034f
C895 commonsourceibias.n392 gnd 0.008037f
C896 commonsourceibias.t60 gnd 0.150157f
C897 commonsourceibias.n393 gnd 0.007578f
C898 commonsourceibias.n394 gnd 0.008037f
C899 commonsourceibias.t16 gnd 0.150157f
C900 commonsourceibias.n395 gnd 0.010186f
C901 commonsourceibias.n396 gnd 0.008037f
C902 commonsourceibias.t58 gnd 0.150157f
C903 commonsourceibias.n397 gnd 0.007361f
C904 commonsourceibias.n398 gnd 0.008037f
C905 commonsourceibias.t32 gnd 0.150157f
C906 commonsourceibias.n399 gnd 0.010015f
C907 commonsourceibias.n400 gnd 0.008037f
C908 commonsourceibias.t72 gnd 0.150157f
C909 commonsourceibias.n401 gnd 0.007172f
C910 commonsourceibias.n402 gnd 0.008037f
C911 commonsourceibias.t54 gnd 0.150157f
C912 commonsourceibias.n403 gnd 0.009825f
C913 commonsourceibias.n404 gnd 0.008037f
C914 commonsourceibias.t6 gnd 0.150157f
C915 commonsourceibias.n405 gnd 0.007008f
C916 commonsourceibias.n406 gnd 0.008037f
C917 commonsourceibias.t66 gnd 0.150157f
C918 commonsourceibias.n407 gnd 0.009613f
C919 commonsourceibias.n408 gnd 0.008037f
C920 commonsourceibias.t14 gnd 0.150157f
C921 commonsourceibias.n409 gnd 0.006868f
C922 commonsourceibias.n410 gnd 0.008037f
C923 commonsourceibias.t48 gnd 0.150157f
C924 commonsourceibias.n411 gnd 0.009378f
C925 commonsourceibias.t30 gnd 0.166947f
C926 commonsourceibias.t2 gnd 0.150157f
C927 commonsourceibias.n412 gnd 0.065449f
C928 commonsourceibias.n413 gnd 0.071822f
C929 commonsourceibias.n414 gnd 0.033327f
C930 commonsourceibias.n415 gnd 0.008037f
C931 commonsourceibias.n416 gnd 0.007823f
C932 commonsourceibias.n417 gnd 0.01121f
C933 commonsourceibias.n418 gnd 0.059912f
C934 commonsourceibias.n419 gnd 0.011203f
C935 commonsourceibias.n420 gnd 0.008037f
C936 commonsourceibias.n421 gnd 0.008037f
C937 commonsourceibias.n422 gnd 0.008037f
C938 commonsourceibias.n423 gnd 0.01034f
C939 commonsourceibias.n424 gnd 0.059912f
C940 commonsourceibias.n425 gnd 0.010583f
C941 commonsourceibias.t68 gnd 0.150157f
C942 commonsourceibias.n426 gnd 0.059912f
C943 commonsourceibias.n427 gnd 0.010282f
C944 commonsourceibias.n428 gnd 0.008037f
C945 commonsourceibias.n429 gnd 0.008037f
C946 commonsourceibias.n430 gnd 0.008037f
C947 commonsourceibias.n431 gnd 0.007578f
C948 commonsourceibias.n432 gnd 0.01122f
C949 commonsourceibias.n433 gnd 0.059912f
C950 commonsourceibias.n434 gnd 0.011217f
C951 commonsourceibias.n435 gnd 0.008037f
C952 commonsourceibias.n436 gnd 0.008037f
C953 commonsourceibias.n437 gnd 0.008037f
C954 commonsourceibias.n438 gnd 0.010186f
C955 commonsourceibias.n439 gnd 0.059912f
C956 commonsourceibias.n440 gnd 0.010507f
C957 commonsourceibias.t62 gnd 0.150157f
C958 commonsourceibias.n441 gnd 0.059912f
C959 commonsourceibias.n442 gnd 0.010357f
C960 commonsourceibias.n443 gnd 0.008037f
C961 commonsourceibias.n444 gnd 0.008037f
C962 commonsourceibias.n445 gnd 0.008037f
C963 commonsourceibias.n446 gnd 0.007361f
C964 commonsourceibias.n447 gnd 0.011225f
C965 commonsourceibias.n448 gnd 0.059912f
C966 commonsourceibias.n449 gnd 0.011224f
C967 commonsourceibias.n450 gnd 0.008037f
C968 commonsourceibias.n451 gnd 0.008037f
C969 commonsourceibias.n452 gnd 0.008037f
C970 commonsourceibias.n453 gnd 0.010015f
C971 commonsourceibias.n454 gnd 0.059912f
C972 commonsourceibias.n455 gnd 0.010432f
C973 commonsourceibias.t64 gnd 0.150157f
C974 commonsourceibias.n456 gnd 0.059912f
C975 commonsourceibias.n457 gnd 0.010432f
C976 commonsourceibias.n458 gnd 0.008037f
C977 commonsourceibias.n459 gnd 0.008037f
C978 commonsourceibias.n460 gnd 0.008037f
C979 commonsourceibias.n461 gnd 0.007172f
C980 commonsourceibias.n462 gnd 0.011224f
C981 commonsourceibias.n463 gnd 0.059912f
C982 commonsourceibias.n464 gnd 0.011225f
C983 commonsourceibias.n465 gnd 0.008037f
C984 commonsourceibias.n466 gnd 0.008037f
C985 commonsourceibias.n467 gnd 0.008037f
C986 commonsourceibias.n468 gnd 0.009825f
C987 commonsourceibias.n469 gnd 0.059912f
C988 commonsourceibias.n470 gnd 0.010357f
C989 commonsourceibias.t44 gnd 0.150157f
C990 commonsourceibias.n471 gnd 0.059912f
C991 commonsourceibias.n472 gnd 0.010507f
C992 commonsourceibias.n473 gnd 0.008037f
C993 commonsourceibias.n474 gnd 0.008037f
C994 commonsourceibias.n475 gnd 0.008037f
C995 commonsourceibias.n476 gnd 0.007008f
C996 commonsourceibias.n477 gnd 0.011217f
C997 commonsourceibias.n478 gnd 0.059912f
C998 commonsourceibias.n479 gnd 0.01122f
C999 commonsourceibias.n480 gnd 0.008037f
C1000 commonsourceibias.n481 gnd 0.008037f
C1001 commonsourceibias.n482 gnd 0.008037f
C1002 commonsourceibias.n483 gnd 0.009613f
C1003 commonsourceibias.n484 gnd 0.059912f
C1004 commonsourceibias.n485 gnd 0.010282f
C1005 commonsourceibias.t28 gnd 0.150157f
C1006 commonsourceibias.n486 gnd 0.059912f
C1007 commonsourceibias.n487 gnd 0.010583f
C1008 commonsourceibias.n488 gnd 0.008037f
C1009 commonsourceibias.n489 gnd 0.008037f
C1010 commonsourceibias.n490 gnd 0.008037f
C1011 commonsourceibias.n491 gnd 0.006868f
C1012 commonsourceibias.n492 gnd 0.011203f
C1013 commonsourceibias.n493 gnd 0.059912f
C1014 commonsourceibias.n494 gnd 0.01121f
C1015 commonsourceibias.n495 gnd 0.008037f
C1016 commonsourceibias.n496 gnd 0.008037f
C1017 commonsourceibias.n497 gnd 0.008037f
C1018 commonsourceibias.n498 gnd 0.009378f
C1019 commonsourceibias.n499 gnd 0.059912f
C1020 commonsourceibias.n500 gnd 0.009861f
C1021 commonsourceibias.t12 gnd 0.162395f
C1022 commonsourceibias.n501 gnd 0.07189f
C1023 commonsourceibias.n502 gnd 0.080075f
C1024 commonsourceibias.t43 gnd 0.017343f
C1025 commonsourceibias.t13 gnd 0.017343f
C1026 commonsourceibias.n503 gnd 0.15325f
C1027 commonsourceibias.n504 gnd 0.132562f
C1028 commonsourceibias.t29 gnd 0.017343f
C1029 commonsourceibias.t1 gnd 0.017343f
C1030 commonsourceibias.n505 gnd 0.15325f
C1031 commonsourceibias.n506 gnd 0.070394f
C1032 commonsourceibias.t17 gnd 0.017343f
C1033 commonsourceibias.t61 gnd 0.017343f
C1034 commonsourceibias.n507 gnd 0.15325f
C1035 commonsourceibias.n508 gnd 0.070394f
C1036 commonsourceibias.t59 gnd 0.017343f
C1037 commonsourceibias.t45 gnd 0.017343f
C1038 commonsourceibias.n509 gnd 0.15325f
C1039 commonsourceibias.n510 gnd 0.070394f
C1040 commonsourceibias.t65 gnd 0.017343f
C1041 commonsourceibias.t33 gnd 0.017343f
C1042 commonsourceibias.n511 gnd 0.15325f
C1043 commonsourceibias.n512 gnd 0.058811f
C1044 commonsourceibias.n513 gnd 0.071213f
C1045 commonsourceibias.n514 gnd 0.052016f
C1046 commonsourceibias.t82 gnd 0.150157f
C1047 commonsourceibias.n515 gnd 0.059912f
C1048 commonsourceibias.n516 gnd 0.008037f
C1049 commonsourceibias.t148 gnd 0.150157f
C1050 commonsourceibias.n517 gnd 0.059912f
C1051 commonsourceibias.n518 gnd 0.008037f
C1052 commonsourceibias.t143 gnd 0.150157f
C1053 commonsourceibias.n519 gnd 0.059912f
C1054 commonsourceibias.n520 gnd 0.008037f
C1055 commonsourceibias.t158 gnd 0.150157f
C1056 commonsourceibias.n521 gnd 0.007008f
C1057 commonsourceibias.n522 gnd 0.008037f
C1058 commonsourceibias.t105 gnd 0.150157f
C1059 commonsourceibias.n523 gnd 0.009613f
C1060 commonsourceibias.n524 gnd 0.008037f
C1061 commonsourceibias.t133 gnd 0.150157f
C1062 commonsourceibias.n525 gnd 0.006868f
C1063 commonsourceibias.n526 gnd 0.008037f
C1064 commonsourceibias.t150 gnd 0.150157f
C1065 commonsourceibias.n527 gnd 0.009378f
C1066 commonsourceibias.t123 gnd 0.166947f
C1067 commonsourceibias.t103 gnd 0.150157f
C1068 commonsourceibias.n528 gnd 0.065449f
C1069 commonsourceibias.n529 gnd 0.071822f
C1070 commonsourceibias.n530 gnd 0.033327f
C1071 commonsourceibias.n531 gnd 0.008037f
C1072 commonsourceibias.n532 gnd 0.007823f
C1073 commonsourceibias.n533 gnd 0.01121f
C1074 commonsourceibias.n534 gnd 0.059912f
C1075 commonsourceibias.n535 gnd 0.011203f
C1076 commonsourceibias.n536 gnd 0.008037f
C1077 commonsourceibias.n537 gnd 0.008037f
C1078 commonsourceibias.n538 gnd 0.008037f
C1079 commonsourceibias.n539 gnd 0.01034f
C1080 commonsourceibias.n540 gnd 0.059912f
C1081 commonsourceibias.n541 gnd 0.010583f
C1082 commonsourceibias.t113 gnd 0.150157f
C1083 commonsourceibias.n542 gnd 0.059912f
C1084 commonsourceibias.n543 gnd 0.010282f
C1085 commonsourceibias.n544 gnd 0.008037f
C1086 commonsourceibias.n545 gnd 0.008037f
C1087 commonsourceibias.n546 gnd 0.008037f
C1088 commonsourceibias.n547 gnd 0.007578f
C1089 commonsourceibias.n548 gnd 0.01122f
C1090 commonsourceibias.n549 gnd 0.059912f
C1091 commonsourceibias.n550 gnd 0.011217f
C1092 commonsourceibias.n551 gnd 0.008037f
C1093 commonsourceibias.n552 gnd 0.008037f
C1094 commonsourceibias.n553 gnd 0.008037f
C1095 commonsourceibias.n554 gnd 0.010186f
C1096 commonsourceibias.n555 gnd 0.059912f
C1097 commonsourceibias.n556 gnd 0.010507f
C1098 commonsourceibias.n557 gnd 0.010357f
C1099 commonsourceibias.n558 gnd 0.008037f
C1100 commonsourceibias.n559 gnd 0.008037f
C1101 commonsourceibias.n560 gnd 0.009825f
C1102 commonsourceibias.n561 gnd 0.007361f
C1103 commonsourceibias.n562 gnd 0.011225f
C1104 commonsourceibias.n563 gnd 0.008037f
C1105 commonsourceibias.n564 gnd 0.008037f
C1106 commonsourceibias.n565 gnd 0.011224f
C1107 commonsourceibias.n566 gnd 0.007172f
C1108 commonsourceibias.n567 gnd 0.010015f
C1109 commonsourceibias.n568 gnd 0.008037f
C1110 commonsourceibias.n569 gnd 0.007021f
C1111 commonsourceibias.n570 gnd 0.010432f
C1112 commonsourceibias.t85 gnd 0.150157f
C1113 commonsourceibias.n571 gnd 0.059912f
C1114 commonsourceibias.n572 gnd 0.010432f
C1115 commonsourceibias.n573 gnd 0.007021f
C1116 commonsourceibias.n574 gnd 0.008037f
C1117 commonsourceibias.n575 gnd 0.008037f
C1118 commonsourceibias.n576 gnd 0.007172f
C1119 commonsourceibias.n577 gnd 0.011224f
C1120 commonsourceibias.n578 gnd 0.059912f
C1121 commonsourceibias.n579 gnd 0.011225f
C1122 commonsourceibias.n580 gnd 0.008037f
C1123 commonsourceibias.n581 gnd 0.008037f
C1124 commonsourceibias.n582 gnd 0.008037f
C1125 commonsourceibias.n583 gnd 0.009825f
C1126 commonsourceibias.n584 gnd 0.059912f
C1127 commonsourceibias.n585 gnd 0.010357f
C1128 commonsourceibias.t89 gnd 0.150157f
C1129 commonsourceibias.n586 gnd 0.059912f
C1130 commonsourceibias.n587 gnd 0.010507f
C1131 commonsourceibias.n588 gnd 0.008037f
C1132 commonsourceibias.n589 gnd 0.008037f
C1133 commonsourceibias.n590 gnd 0.008037f
C1134 commonsourceibias.n591 gnd 0.007008f
C1135 commonsourceibias.n592 gnd 0.011217f
C1136 commonsourceibias.n593 gnd 0.059912f
C1137 commonsourceibias.n594 gnd 0.01122f
C1138 commonsourceibias.n595 gnd 0.008037f
C1139 commonsourceibias.n596 gnd 0.008037f
C1140 commonsourceibias.n597 gnd 0.008037f
C1141 commonsourceibias.n598 gnd 0.009613f
C1142 commonsourceibias.n599 gnd 0.059912f
C1143 commonsourceibias.n600 gnd 0.010282f
C1144 commonsourceibias.t130 gnd 0.150157f
C1145 commonsourceibias.n601 gnd 0.059912f
C1146 commonsourceibias.n602 gnd 0.010583f
C1147 commonsourceibias.n603 gnd 0.008037f
C1148 commonsourceibias.n604 gnd 0.008037f
C1149 commonsourceibias.n605 gnd 0.008037f
C1150 commonsourceibias.n606 gnd 0.006868f
C1151 commonsourceibias.n607 gnd 0.011203f
C1152 commonsourceibias.n608 gnd 0.059912f
C1153 commonsourceibias.n609 gnd 0.01121f
C1154 commonsourceibias.n610 gnd 0.008037f
C1155 commonsourceibias.n611 gnd 0.008037f
C1156 commonsourceibias.n612 gnd 0.008037f
C1157 commonsourceibias.n613 gnd 0.009378f
C1158 commonsourceibias.n614 gnd 0.059912f
C1159 commonsourceibias.n615 gnd 0.009861f
C1160 commonsourceibias.n616 gnd 0.07189f
C1161 commonsourceibias.n617 gnd 0.04697f
C1162 commonsourceibias.n618 gnd 0.010724f
C1163 commonsourceibias.t141 gnd 0.150157f
C1164 commonsourceibias.n619 gnd 0.007823f
C1165 commonsourceibias.n620 gnd 0.008037f
C1166 commonsourceibias.t156 gnd 0.150157f
C1167 commonsourceibias.n621 gnd 0.01034f
C1168 commonsourceibias.n622 gnd 0.008037f
C1169 commonsourceibias.t131 gnd 0.150157f
C1170 commonsourceibias.n623 gnd 0.007578f
C1171 commonsourceibias.n624 gnd 0.008037f
C1172 commonsourceibias.t149 gnd 0.150157f
C1173 commonsourceibias.n625 gnd 0.010186f
C1174 commonsourceibias.n626 gnd 0.008037f
C1175 commonsourceibias.t97 gnd 0.150157f
C1176 commonsourceibias.n627 gnd 0.007361f
C1177 commonsourceibias.n628 gnd 0.008037f
C1178 commonsourceibias.t142 gnd 0.150157f
C1179 commonsourceibias.n629 gnd 0.010015f
C1180 commonsourceibias.n630 gnd 0.008037f
C1181 commonsourceibias.t153 gnd 0.150157f
C1182 commonsourceibias.n631 gnd 0.007172f
C1183 commonsourceibias.n632 gnd 0.008037f
C1184 commonsourceibias.t132 gnd 0.150157f
C1185 commonsourceibias.n633 gnd 0.009825f
C1186 commonsourceibias.n634 gnd 0.008037f
C1187 commonsourceibias.t146 gnd 0.150157f
C1188 commonsourceibias.n635 gnd 0.007008f
C1189 commonsourceibias.n636 gnd 0.008037f
C1190 commonsourceibias.t92 gnd 0.150157f
C1191 commonsourceibias.n637 gnd 0.009613f
C1192 commonsourceibias.n638 gnd 0.008037f
C1193 commonsourceibias.t116 gnd 0.150157f
C1194 commonsourceibias.n639 gnd 0.006868f
C1195 commonsourceibias.n640 gnd 0.008037f
C1196 commonsourceibias.t135 gnd 0.150157f
C1197 commonsourceibias.n641 gnd 0.009378f
C1198 commonsourceibias.t107 gnd 0.166947f
C1199 commonsourceibias.t90 gnd 0.150157f
C1200 commonsourceibias.n642 gnd 0.065449f
C1201 commonsourceibias.n643 gnd 0.071822f
C1202 commonsourceibias.n644 gnd 0.033327f
C1203 commonsourceibias.n645 gnd 0.008037f
C1204 commonsourceibias.n646 gnd 0.007823f
C1205 commonsourceibias.n647 gnd 0.01121f
C1206 commonsourceibias.n648 gnd 0.059912f
C1207 commonsourceibias.n649 gnd 0.011203f
C1208 commonsourceibias.n650 gnd 0.008037f
C1209 commonsourceibias.n651 gnd 0.008037f
C1210 commonsourceibias.n652 gnd 0.008037f
C1211 commonsourceibias.n653 gnd 0.01034f
C1212 commonsourceibias.n654 gnd 0.059912f
C1213 commonsourceibias.n655 gnd 0.010583f
C1214 commonsourceibias.t98 gnd 0.150157f
C1215 commonsourceibias.n656 gnd 0.059912f
C1216 commonsourceibias.n657 gnd 0.010282f
C1217 commonsourceibias.n658 gnd 0.008037f
C1218 commonsourceibias.n659 gnd 0.008037f
C1219 commonsourceibias.n660 gnd 0.008037f
C1220 commonsourceibias.n661 gnd 0.007578f
C1221 commonsourceibias.n662 gnd 0.01122f
C1222 commonsourceibias.n663 gnd 0.059912f
C1223 commonsourceibias.n664 gnd 0.011217f
C1224 commonsourceibias.n665 gnd 0.008037f
C1225 commonsourceibias.n666 gnd 0.008037f
C1226 commonsourceibias.n667 gnd 0.008037f
C1227 commonsourceibias.n668 gnd 0.010186f
C1228 commonsourceibias.n669 gnd 0.059912f
C1229 commonsourceibias.n670 gnd 0.010507f
C1230 commonsourceibias.t125 gnd 0.150157f
C1231 commonsourceibias.n671 gnd 0.059912f
C1232 commonsourceibias.n672 gnd 0.010357f
C1233 commonsourceibias.n673 gnd 0.008037f
C1234 commonsourceibias.n674 gnd 0.008037f
C1235 commonsourceibias.n675 gnd 0.008037f
C1236 commonsourceibias.n676 gnd 0.007361f
C1237 commonsourceibias.n677 gnd 0.011225f
C1238 commonsourceibias.n678 gnd 0.059912f
C1239 commonsourceibias.n679 gnd 0.011224f
C1240 commonsourceibias.n680 gnd 0.008037f
C1241 commonsourceibias.n681 gnd 0.008037f
C1242 commonsourceibias.n682 gnd 0.008037f
C1243 commonsourceibias.n683 gnd 0.010015f
C1244 commonsourceibias.n684 gnd 0.059912f
C1245 commonsourceibias.n685 gnd 0.010432f
C1246 commonsourceibias.t157 gnd 0.150157f
C1247 commonsourceibias.n686 gnd 0.059912f
C1248 commonsourceibias.n687 gnd 0.010432f
C1249 commonsourceibias.n688 gnd 0.008037f
C1250 commonsourceibias.n689 gnd 0.008037f
C1251 commonsourceibias.n690 gnd 0.008037f
C1252 commonsourceibias.n691 gnd 0.007172f
C1253 commonsourceibias.n692 gnd 0.011224f
C1254 commonsourceibias.n693 gnd 0.059912f
C1255 commonsourceibias.n694 gnd 0.011225f
C1256 commonsourceibias.n695 gnd 0.008037f
C1257 commonsourceibias.n696 gnd 0.008037f
C1258 commonsourceibias.n697 gnd 0.008037f
C1259 commonsourceibias.n698 gnd 0.009825f
C1260 commonsourceibias.n699 gnd 0.059912f
C1261 commonsourceibias.n700 gnd 0.010357f
C1262 commonsourceibias.t81 gnd 0.150157f
C1263 commonsourceibias.n701 gnd 0.059912f
C1264 commonsourceibias.n702 gnd 0.010507f
C1265 commonsourceibias.n703 gnd 0.008037f
C1266 commonsourceibias.n704 gnd 0.008037f
C1267 commonsourceibias.n705 gnd 0.008037f
C1268 commonsourceibias.n706 gnd 0.007008f
C1269 commonsourceibias.n707 gnd 0.011217f
C1270 commonsourceibias.n708 gnd 0.059912f
C1271 commonsourceibias.n709 gnd 0.01122f
C1272 commonsourceibias.n710 gnd 0.008037f
C1273 commonsourceibias.n711 gnd 0.008037f
C1274 commonsourceibias.n712 gnd 0.008037f
C1275 commonsourceibias.n713 gnd 0.009613f
C1276 commonsourceibias.n714 gnd 0.059912f
C1277 commonsourceibias.n715 gnd 0.010282f
C1278 commonsourceibias.t111 gnd 0.150157f
C1279 commonsourceibias.n716 gnd 0.059912f
C1280 commonsourceibias.n717 gnd 0.010583f
C1281 commonsourceibias.n718 gnd 0.008037f
C1282 commonsourceibias.n719 gnd 0.008037f
C1283 commonsourceibias.n720 gnd 0.008037f
C1284 commonsourceibias.n721 gnd 0.006868f
C1285 commonsourceibias.n722 gnd 0.011203f
C1286 commonsourceibias.n723 gnd 0.059912f
C1287 commonsourceibias.n724 gnd 0.01121f
C1288 commonsourceibias.n725 gnd 0.008037f
C1289 commonsourceibias.n726 gnd 0.008037f
C1290 commonsourceibias.n727 gnd 0.008037f
C1291 commonsourceibias.n728 gnd 0.009378f
C1292 commonsourceibias.n729 gnd 0.059912f
C1293 commonsourceibias.n730 gnd 0.009861f
C1294 commonsourceibias.t122 gnd 0.162395f
C1295 commonsourceibias.n731 gnd 0.07189f
C1296 commonsourceibias.n732 gnd 0.025003f
C1297 commonsourceibias.n733 gnd 0.221951f
C1298 commonsourceibias.n734 gnd 4.85761f
C1299 outputibias.t10 gnd 0.11477f
C1300 outputibias.t8 gnd 0.115567f
C1301 outputibias.n0 gnd 0.130108f
C1302 outputibias.n1 gnd 0.001372f
C1303 outputibias.n2 gnd 9.76e-19
C1304 outputibias.n3 gnd 5.24e-19
C1305 outputibias.n4 gnd 0.001239f
C1306 outputibias.n5 gnd 5.55e-19
C1307 outputibias.n6 gnd 9.76e-19
C1308 outputibias.n7 gnd 5.24e-19
C1309 outputibias.n8 gnd 0.001239f
C1310 outputibias.n9 gnd 5.55e-19
C1311 outputibias.n10 gnd 0.004176f
C1312 outputibias.t5 gnd 0.00202f
C1313 outputibias.n11 gnd 9.3e-19
C1314 outputibias.n12 gnd 7.32e-19
C1315 outputibias.n13 gnd 5.24e-19
C1316 outputibias.n14 gnd 0.02322f
C1317 outputibias.n15 gnd 9.76e-19
C1318 outputibias.n16 gnd 5.24e-19
C1319 outputibias.n17 gnd 5.55e-19
C1320 outputibias.n18 gnd 0.001239f
C1321 outputibias.n19 gnd 0.001239f
C1322 outputibias.n20 gnd 5.55e-19
C1323 outputibias.n21 gnd 5.24e-19
C1324 outputibias.n22 gnd 9.76e-19
C1325 outputibias.n23 gnd 9.76e-19
C1326 outputibias.n24 gnd 5.24e-19
C1327 outputibias.n25 gnd 5.55e-19
C1328 outputibias.n26 gnd 0.001239f
C1329 outputibias.n27 gnd 0.002683f
C1330 outputibias.n28 gnd 5.55e-19
C1331 outputibias.n29 gnd 5.24e-19
C1332 outputibias.n30 gnd 0.002256f
C1333 outputibias.n31 gnd 0.005781f
C1334 outputibias.n32 gnd 0.001372f
C1335 outputibias.n33 gnd 9.76e-19
C1336 outputibias.n34 gnd 5.24e-19
C1337 outputibias.n35 gnd 0.001239f
C1338 outputibias.n36 gnd 5.55e-19
C1339 outputibias.n37 gnd 9.76e-19
C1340 outputibias.n38 gnd 5.24e-19
C1341 outputibias.n39 gnd 0.001239f
C1342 outputibias.n40 gnd 5.55e-19
C1343 outputibias.n41 gnd 0.004176f
C1344 outputibias.t3 gnd 0.00202f
C1345 outputibias.n42 gnd 9.3e-19
C1346 outputibias.n43 gnd 7.32e-19
C1347 outputibias.n44 gnd 5.24e-19
C1348 outputibias.n45 gnd 0.02322f
C1349 outputibias.n46 gnd 9.76e-19
C1350 outputibias.n47 gnd 5.24e-19
C1351 outputibias.n48 gnd 5.55e-19
C1352 outputibias.n49 gnd 0.001239f
C1353 outputibias.n50 gnd 0.001239f
C1354 outputibias.n51 gnd 5.55e-19
C1355 outputibias.n52 gnd 5.24e-19
C1356 outputibias.n53 gnd 9.76e-19
C1357 outputibias.n54 gnd 9.76e-19
C1358 outputibias.n55 gnd 5.24e-19
C1359 outputibias.n56 gnd 5.55e-19
C1360 outputibias.n57 gnd 0.001239f
C1361 outputibias.n58 gnd 0.002683f
C1362 outputibias.n59 gnd 5.55e-19
C1363 outputibias.n60 gnd 5.24e-19
C1364 outputibias.n61 gnd 0.002256f
C1365 outputibias.n62 gnd 0.005197f
C1366 outputibias.n63 gnd 0.121892f
C1367 outputibias.n64 gnd 0.001372f
C1368 outputibias.n65 gnd 9.76e-19
C1369 outputibias.n66 gnd 5.24e-19
C1370 outputibias.n67 gnd 0.001239f
C1371 outputibias.n68 gnd 5.55e-19
C1372 outputibias.n69 gnd 9.76e-19
C1373 outputibias.n70 gnd 5.24e-19
C1374 outputibias.n71 gnd 0.001239f
C1375 outputibias.n72 gnd 5.55e-19
C1376 outputibias.n73 gnd 0.004176f
C1377 outputibias.t1 gnd 0.00202f
C1378 outputibias.n74 gnd 9.3e-19
C1379 outputibias.n75 gnd 7.32e-19
C1380 outputibias.n76 gnd 5.24e-19
C1381 outputibias.n77 gnd 0.02322f
C1382 outputibias.n78 gnd 9.76e-19
C1383 outputibias.n79 gnd 5.24e-19
C1384 outputibias.n80 gnd 5.55e-19
C1385 outputibias.n81 gnd 0.001239f
C1386 outputibias.n82 gnd 0.001239f
C1387 outputibias.n83 gnd 5.55e-19
C1388 outputibias.n84 gnd 5.24e-19
C1389 outputibias.n85 gnd 9.76e-19
C1390 outputibias.n86 gnd 9.76e-19
C1391 outputibias.n87 gnd 5.24e-19
C1392 outputibias.n88 gnd 5.55e-19
C1393 outputibias.n89 gnd 0.001239f
C1394 outputibias.n90 gnd 0.002683f
C1395 outputibias.n91 gnd 5.55e-19
C1396 outputibias.n92 gnd 5.24e-19
C1397 outputibias.n93 gnd 0.002256f
C1398 outputibias.n94 gnd 0.005197f
C1399 outputibias.n95 gnd 0.064513f
C1400 outputibias.n96 gnd 0.001372f
C1401 outputibias.n97 gnd 9.76e-19
C1402 outputibias.n98 gnd 5.24e-19
C1403 outputibias.n99 gnd 0.001239f
C1404 outputibias.n100 gnd 5.55e-19
C1405 outputibias.n101 gnd 9.76e-19
C1406 outputibias.n102 gnd 5.24e-19
C1407 outputibias.n103 gnd 0.001239f
C1408 outputibias.n104 gnd 5.55e-19
C1409 outputibias.n105 gnd 0.004176f
C1410 outputibias.t7 gnd 0.00202f
C1411 outputibias.n106 gnd 9.3e-19
C1412 outputibias.n107 gnd 7.32e-19
C1413 outputibias.n108 gnd 5.24e-19
C1414 outputibias.n109 gnd 0.02322f
C1415 outputibias.n110 gnd 9.76e-19
C1416 outputibias.n111 gnd 5.24e-19
C1417 outputibias.n112 gnd 5.55e-19
C1418 outputibias.n113 gnd 0.001239f
C1419 outputibias.n114 gnd 0.001239f
C1420 outputibias.n115 gnd 5.55e-19
C1421 outputibias.n116 gnd 5.24e-19
C1422 outputibias.n117 gnd 9.76e-19
C1423 outputibias.n118 gnd 9.76e-19
C1424 outputibias.n119 gnd 5.24e-19
C1425 outputibias.n120 gnd 5.55e-19
C1426 outputibias.n121 gnd 0.001239f
C1427 outputibias.n122 gnd 0.002683f
C1428 outputibias.n123 gnd 5.55e-19
C1429 outputibias.n124 gnd 5.24e-19
C1430 outputibias.n125 gnd 0.002256f
C1431 outputibias.n126 gnd 0.005197f
C1432 outputibias.n127 gnd 0.084814f
C1433 outputibias.t6 gnd 0.108319f
C1434 outputibias.t0 gnd 0.108319f
C1435 outputibias.t2 gnd 0.108319f
C1436 outputibias.t4 gnd 0.109238f
C1437 outputibias.n128 gnd 0.134674f
C1438 outputibias.n129 gnd 0.07244f
C1439 outputibias.n130 gnd 0.079818f
C1440 outputibias.n131 gnd 0.164901f
C1441 outputibias.t11 gnd 0.11477f
C1442 outputibias.n132 gnd 0.067481f
C1443 outputibias.t9 gnd 0.11477f
C1444 outputibias.n133 gnd 0.065115f
C1445 outputibias.n134 gnd 0.029159f
C1446 a_n3827_n3924.t6 gnd 0.095164f
C1447 a_n3827_n3924.t17 gnd 0.989057f
C1448 a_n3827_n3924.n0 gnd 0.373908f
C1449 a_n3827_n3924.t57 gnd 1.2292f
C1450 a_n3827_n3924.n1 gnd 1.25966f
C1451 a_n3827_n3924.t51 gnd 0.989057f
C1452 a_n3827_n3924.n2 gnd 0.373908f
C1453 a_n3827_n3924.t38 gnd 0.095164f
C1454 a_n3827_n3924.t29 gnd 0.095164f
C1455 a_n3827_n3924.n3 gnd 0.777221f
C1456 a_n3827_n3924.n4 gnd 0.391675f
C1457 a_n3827_n3924.t33 gnd 0.095164f
C1458 a_n3827_n3924.t37 gnd 0.095164f
C1459 a_n3827_n3924.n5 gnd 0.777221f
C1460 a_n3827_n3924.n6 gnd 0.391675f
C1461 a_n3827_n3924.t49 gnd 0.095164f
C1462 a_n3827_n3924.t32 gnd 0.095164f
C1463 a_n3827_n3924.n7 gnd 0.777221f
C1464 a_n3827_n3924.n8 gnd 0.391675f
C1465 a_n3827_n3924.t42 gnd 0.095164f
C1466 a_n3827_n3924.t53 gnd 0.095164f
C1467 a_n3827_n3924.n9 gnd 0.777221f
C1468 a_n3827_n3924.n10 gnd 0.391675f
C1469 a_n3827_n3924.t44 gnd 0.095164f
C1470 a_n3827_n3924.t45 gnd 0.095164f
C1471 a_n3827_n3924.n11 gnd 0.777221f
C1472 a_n3827_n3924.n12 gnd 0.391675f
C1473 a_n3827_n3924.t31 gnd 0.989057f
C1474 a_n3827_n3924.n13 gnd 0.925833f
C1475 a_n3827_n3924.t27 gnd 1.23041f
C1476 a_n3827_n3924.t26 gnd 1.22888f
C1477 a_n3827_n3924.n14 gnd 0.823361f
C1478 a_n3827_n3924.t55 gnd 1.22888f
C1479 a_n3827_n3924.n15 gnd 0.865521f
C1480 a_n3827_n3924.t46 gnd 1.22888f
C1481 a_n3827_n3924.n16 gnd 0.865521f
C1482 a_n3827_n3924.t56 gnd 1.22888f
C1483 a_n3827_n3924.n17 gnd 0.865521f
C1484 a_n3827_n3924.t25 gnd 1.22888f
C1485 a_n3827_n3924.n18 gnd 0.865521f
C1486 a_n3827_n3924.t54 gnd 1.22888f
C1487 a_n3827_n3924.n19 gnd 0.865521f
C1488 a_n3827_n3924.t24 gnd 1.22888f
C1489 a_n3827_n3924.n20 gnd 0.865521f
C1490 a_n3827_n3924.t28 gnd 1.22888f
C1491 a_n3827_n3924.n21 gnd 0.565437f
C1492 a_n3827_n3924.n22 gnd 1.00053f
C1493 a_n3827_n3924.n23 gnd 0.897154f
C1494 a_n3827_n3924.t8 gnd 0.989054f
C1495 a_n3827_n3924.n24 gnd 0.61435f
C1496 a_n3827_n3924.t5 gnd 0.095164f
C1497 a_n3827_n3924.t22 gnd 0.095164f
C1498 a_n3827_n3924.n25 gnd 0.777219f
C1499 a_n3827_n3924.n26 gnd 0.391677f
C1500 a_n3827_n3924.t16 gnd 0.095164f
C1501 a_n3827_n3924.t20 gnd 0.095164f
C1502 a_n3827_n3924.n27 gnd 0.777219f
C1503 a_n3827_n3924.n28 gnd 0.391677f
C1504 a_n3827_n3924.t21 gnd 0.095164f
C1505 a_n3827_n3924.t9 gnd 0.095164f
C1506 a_n3827_n3924.n29 gnd 0.777219f
C1507 a_n3827_n3924.n30 gnd 0.391677f
C1508 a_n3827_n3924.t10 gnd 0.095164f
C1509 a_n3827_n3924.t1 gnd 0.095164f
C1510 a_n3827_n3924.n31 gnd 0.777219f
C1511 a_n3827_n3924.n32 gnd 0.391677f
C1512 a_n3827_n3924.t3 gnd 0.095164f
C1513 a_n3827_n3924.t19 gnd 0.095164f
C1514 a_n3827_n3924.n33 gnd 0.777219f
C1515 a_n3827_n3924.n34 gnd 0.391677f
C1516 a_n3827_n3924.t14 gnd 0.989054f
C1517 a_n3827_n3924.n35 gnd 0.373911f
C1518 a_n3827_n3924.t48 gnd 0.989054f
C1519 a_n3827_n3924.n36 gnd 0.373911f
C1520 a_n3827_n3924.t39 gnd 0.095164f
C1521 a_n3827_n3924.t30 gnd 0.095164f
C1522 a_n3827_n3924.n37 gnd 0.777219f
C1523 a_n3827_n3924.n38 gnd 0.391677f
C1524 a_n3827_n3924.t34 gnd 0.095164f
C1525 a_n3827_n3924.t50 gnd 0.095164f
C1526 a_n3827_n3924.n39 gnd 0.777219f
C1527 a_n3827_n3924.n40 gnd 0.391677f
C1528 a_n3827_n3924.t52 gnd 0.095164f
C1529 a_n3827_n3924.t47 gnd 0.095164f
C1530 a_n3827_n3924.n41 gnd 0.777219f
C1531 a_n3827_n3924.n42 gnd 0.391677f
C1532 a_n3827_n3924.t43 gnd 0.095164f
C1533 a_n3827_n3924.t36 gnd 0.095164f
C1534 a_n3827_n3924.n43 gnd 0.777219f
C1535 a_n3827_n3924.n44 gnd 0.391677f
C1536 a_n3827_n3924.t41 gnd 0.095164f
C1537 a_n3827_n3924.t40 gnd 0.095164f
C1538 a_n3827_n3924.n45 gnd 0.777219f
C1539 a_n3827_n3924.n46 gnd 0.391677f
C1540 a_n3827_n3924.t35 gnd 0.989054f
C1541 a_n3827_n3924.n47 gnd 0.61435f
C1542 a_n3827_n3924.n48 gnd 0.897154f
C1543 a_n3827_n3924.t4 gnd 0.989053f
C1544 a_n3827_n3924.n49 gnd 0.925837f
C1545 a_n3827_n3924.t2 gnd 0.095164f
C1546 a_n3827_n3924.t0 gnd 0.095164f
C1547 a_n3827_n3924.n50 gnd 0.777221f
C1548 a_n3827_n3924.n51 gnd 0.391675f
C1549 a_n3827_n3924.t13 gnd 0.095164f
C1550 a_n3827_n3924.t18 gnd 0.095164f
C1551 a_n3827_n3924.n52 gnd 0.777221f
C1552 a_n3827_n3924.n53 gnd 0.391675f
C1553 a_n3827_n3924.t11 gnd 0.095164f
C1554 a_n3827_n3924.t15 gnd 0.095164f
C1555 a_n3827_n3924.n54 gnd 0.777221f
C1556 a_n3827_n3924.n55 gnd 0.391675f
C1557 a_n3827_n3924.t7 gnd 0.095164f
C1558 a_n3827_n3924.t12 gnd 0.095164f
C1559 a_n3827_n3924.n56 gnd 0.777221f
C1560 a_n3827_n3924.n57 gnd 0.391675f
C1561 a_n3827_n3924.n58 gnd 0.391674f
C1562 a_n3827_n3924.n59 gnd 0.777222f
C1563 a_n3827_n3924.t23 gnd 0.095164f
C1564 plus.n0 gnd 0.022575f
C1565 plus.t20 gnd 0.410529f
C1566 plus.t23 gnd 0.379592f
C1567 plus.n1 gnd 0.153524f
C1568 plus.n2 gnd 0.022575f
C1569 plus.t6 gnd 0.379592f
C1570 plus.n3 gnd 0.019291f
C1571 plus.n4 gnd 0.022575f
C1572 plus.t12 gnd 0.379592f
C1573 plus.t8 gnd 0.379592f
C1574 plus.n5 gnd 0.153524f
C1575 plus.n6 gnd 0.022575f
C1576 plus.t7 gnd 0.379592f
C1577 plus.n7 gnd 0.153524f
C1578 plus.n8 gnd 0.022575f
C1579 plus.t19 gnd 0.379592f
C1580 plus.n9 gnd 0.018348f
C1581 plus.n10 gnd 0.022575f
C1582 plus.t18 gnd 0.379592f
C1583 plus.t27 gnd 0.379592f
C1584 plus.n11 gnd 0.153524f
C1585 plus.n12 gnd 0.022575f
C1586 plus.t25 gnd 0.379592f
C1587 plus.n13 gnd 0.153524f
C1588 plus.n14 gnd 0.095805f
C1589 plus.t9 gnd 0.379592f
C1590 plus.t14 gnd 0.424642f
C1591 plus.n15 gnd 0.179485f
C1592 plus.n16 gnd 0.175814f
C1593 plus.n17 gnd 0.028926f
C1594 plus.n18 gnd 0.025546f
C1595 plus.n19 gnd 0.022575f
C1596 plus.n20 gnd 0.022575f
C1597 plus.n21 gnd 0.026977f
C1598 plus.n22 gnd 0.019291f
C1599 plus.n23 gnd 0.029401f
C1600 plus.n24 gnd 0.022575f
C1601 plus.n25 gnd 0.022575f
C1602 plus.n26 gnd 0.028081f
C1603 plus.n27 gnd 0.026391f
C1604 plus.n28 gnd 0.153524f
C1605 plus.n29 gnd 0.028279f
C1606 plus.n30 gnd 0.022575f
C1607 plus.n31 gnd 0.022575f
C1608 plus.n32 gnd 0.022575f
C1609 plus.n33 gnd 0.029042f
C1610 plus.n34 gnd 0.153524f
C1611 plus.n35 gnd 0.027236f
C1612 plus.n36 gnd 0.027236f
C1613 plus.n37 gnd 0.022575f
C1614 plus.n38 gnd 0.022575f
C1615 plus.n39 gnd 0.029042f
C1616 plus.n40 gnd 0.018348f
C1617 plus.n41 gnd 0.028279f
C1618 plus.n42 gnd 0.022575f
C1619 plus.n43 gnd 0.022575f
C1620 plus.n44 gnd 0.026391f
C1621 plus.n45 gnd 0.028081f
C1622 plus.n46 gnd 0.153524f
C1623 plus.n47 gnd 0.029401f
C1624 plus.n48 gnd 0.022575f
C1625 plus.n49 gnd 0.022575f
C1626 plus.n50 gnd 0.022575f
C1627 plus.n51 gnd 0.026977f
C1628 plus.n52 gnd 0.153524f
C1629 plus.n53 gnd 0.025546f
C1630 plus.n54 gnd 0.028926f
C1631 plus.n55 gnd 0.022575f
C1632 plus.n56 gnd 0.022575f
C1633 plus.n57 gnd 0.02945f
C1634 plus.n58 gnd 0.008204f
C1635 plus.n59 gnd 0.177755f
C1636 plus.n60 gnd 0.258648f
C1637 plus.n61 gnd 0.022575f
C1638 plus.t28 gnd 0.379592f
C1639 plus.n62 gnd 0.153524f
C1640 plus.n63 gnd 0.022575f
C1641 plus.t26 gnd 0.379592f
C1642 plus.n64 gnd 0.019291f
C1643 plus.n65 gnd 0.022575f
C1644 plus.t10 gnd 0.379592f
C1645 plus.t15 gnd 0.379592f
C1646 plus.n66 gnd 0.153524f
C1647 plus.n67 gnd 0.022575f
C1648 plus.t13 gnd 0.379592f
C1649 plus.n68 gnd 0.153524f
C1650 plus.n69 gnd 0.022575f
C1651 plus.t17 gnd 0.379592f
C1652 plus.n70 gnd 0.018348f
C1653 plus.n71 gnd 0.022575f
C1654 plus.t16 gnd 0.379592f
C1655 plus.t21 gnd 0.379592f
C1656 plus.n72 gnd 0.153524f
C1657 plus.n73 gnd 0.022575f
C1658 plus.t22 gnd 0.379592f
C1659 plus.n74 gnd 0.153524f
C1660 plus.n75 gnd 0.095805f
C1661 plus.t5 gnd 0.379592f
C1662 plus.t11 gnd 0.424642f
C1663 plus.n76 gnd 0.179485f
C1664 plus.n77 gnd 0.175814f
C1665 plus.n78 gnd 0.028926f
C1666 plus.n79 gnd 0.025546f
C1667 plus.n80 gnd 0.022575f
C1668 plus.n81 gnd 0.022575f
C1669 plus.n82 gnd 0.026977f
C1670 plus.n83 gnd 0.019291f
C1671 plus.n84 gnd 0.029401f
C1672 plus.n85 gnd 0.022575f
C1673 plus.n86 gnd 0.022575f
C1674 plus.n87 gnd 0.028081f
C1675 plus.n88 gnd 0.026391f
C1676 plus.n89 gnd 0.153524f
C1677 plus.n90 gnd 0.028279f
C1678 plus.n91 gnd 0.022575f
C1679 plus.n92 gnd 0.022575f
C1680 plus.n93 gnd 0.022575f
C1681 plus.n94 gnd 0.029042f
C1682 plus.n95 gnd 0.153524f
C1683 plus.n96 gnd 0.027236f
C1684 plus.n97 gnd 0.027236f
C1685 plus.n98 gnd 0.022575f
C1686 plus.n99 gnd 0.022575f
C1687 plus.n100 gnd 0.029042f
C1688 plus.n101 gnd 0.018348f
C1689 plus.n102 gnd 0.028279f
C1690 plus.n103 gnd 0.022575f
C1691 plus.n104 gnd 0.022575f
C1692 plus.n105 gnd 0.026391f
C1693 plus.n106 gnd 0.028081f
C1694 plus.n107 gnd 0.153524f
C1695 plus.n108 gnd 0.029401f
C1696 plus.n109 gnd 0.022575f
C1697 plus.n110 gnd 0.022575f
C1698 plus.n111 gnd 0.022575f
C1699 plus.n112 gnd 0.026977f
C1700 plus.n113 gnd 0.153524f
C1701 plus.n114 gnd 0.025546f
C1702 plus.n115 gnd 0.028926f
C1703 plus.n116 gnd 0.022575f
C1704 plus.n117 gnd 0.022575f
C1705 plus.n118 gnd 0.02945f
C1706 plus.n119 gnd 0.008204f
C1707 plus.t24 gnd 0.410529f
C1708 plus.n120 gnd 0.177755f
C1709 plus.n121 gnd 0.814491f
C1710 plus.n122 gnd 1.20072f
C1711 plus.t2 gnd 0.038971f
C1712 plus.t4 gnd 0.006959f
C1713 plus.t0 gnd 0.006959f
C1714 plus.n123 gnd 0.02257f
C1715 plus.n124 gnd 0.175211f
C1716 plus.t3 gnd 0.006959f
C1717 plus.t1 gnd 0.006959f
C1718 plus.n125 gnd 0.02257f
C1719 plus.n126 gnd 0.131517f
C1720 plus.n127 gnd 3.2133f
C1721 a_n1808_13878.t11 gnd 0.185683f
C1722 a_n1808_13878.t13 gnd 0.185683f
C1723 a_n1808_13878.t17 gnd 0.185683f
C1724 a_n1808_13878.n0 gnd 1.46451f
C1725 a_n1808_13878.t8 gnd 0.185683f
C1726 a_n1808_13878.t10 gnd 0.185683f
C1727 a_n1808_13878.n1 gnd 1.46364f
C1728 a_n1808_13878.t14 gnd 0.185683f
C1729 a_n1808_13878.t9 gnd 0.185683f
C1730 a_n1808_13878.n2 gnd 1.46209f
C1731 a_n1808_13878.n3 gnd 2.04299f
C1732 a_n1808_13878.t12 gnd 0.185683f
C1733 a_n1808_13878.t19 gnd 0.185683f
C1734 a_n1808_13878.n4 gnd 1.46209f
C1735 a_n1808_13878.n5 gnd 3.70273f
C1736 a_n1808_13878.t1 gnd 1.73864f
C1737 a_n1808_13878.t4 gnd 0.185683f
C1738 a_n1808_13878.t5 gnd 0.185683f
C1739 a_n1808_13878.n6 gnd 1.30795f
C1740 a_n1808_13878.n7 gnd 1.46144f
C1741 a_n1808_13878.t0 gnd 1.73518f
C1742 a_n1808_13878.n8 gnd 0.735417f
C1743 a_n1808_13878.t3 gnd 1.73518f
C1744 a_n1808_13878.n9 gnd 0.735417f
C1745 a_n1808_13878.t6 gnd 0.185683f
C1746 a_n1808_13878.t7 gnd 0.185683f
C1747 a_n1808_13878.n10 gnd 1.30795f
C1748 a_n1808_13878.n11 gnd 0.742539f
C1749 a_n1808_13878.t2 gnd 1.73518f
C1750 a_n1808_13878.n12 gnd 1.73174f
C1751 a_n1808_13878.n13 gnd 2.52099f
C1752 a_n1808_13878.t15 gnd 0.185683f
C1753 a_n1808_13878.t16 gnd 0.185683f
C1754 a_n1808_13878.n14 gnd 1.46209f
C1755 a_n1808_13878.n15 gnd 1.80499f
C1756 a_n1808_13878.n16 gnd 1.31424f
C1757 a_n1808_13878.n17 gnd 1.46209f
C1758 a_n1808_13878.t18 gnd 0.185683f
C1759 a_n1986_8322.t2 gnd 38.6505f
C1760 a_n1986_8322.t0 gnd 29.5428f
C1761 a_n1986_8322.t3 gnd 19.257301f
C1762 a_n1986_8322.t1 gnd 38.6505f
C1763 a_n1986_8322.t13 gnd 0.875297f
C1764 a_n1986_8322.t21 gnd 0.09348f
C1765 a_n1986_8322.t16 gnd 0.09348f
C1766 a_n1986_8322.n0 gnd 0.658471f
C1767 a_n1986_8322.n1 gnd 0.735745f
C1768 a_n1986_8322.t19 gnd 0.09348f
C1769 a_n1986_8322.t18 gnd 0.09348f
C1770 a_n1986_8322.n2 gnd 0.658471f
C1771 a_n1986_8322.n3 gnd 0.373822f
C1772 a_n1986_8322.t12 gnd 0.873554f
C1773 a_n1986_8322.n4 gnd 1.39817f
C1774 a_n1986_8322.t6 gnd 0.875297f
C1775 a_n1986_8322.t10 gnd 0.09348f
C1776 a_n1986_8322.t9 gnd 0.09348f
C1777 a_n1986_8322.n5 gnd 0.658471f
C1778 a_n1986_8322.n6 gnd 0.735745f
C1779 a_n1986_8322.t4 gnd 0.873554f
C1780 a_n1986_8322.n7 gnd 0.370237f
C1781 a_n1986_8322.t7 gnd 0.873554f
C1782 a_n1986_8322.n8 gnd 0.370237f
C1783 a_n1986_8322.t5 gnd 0.09348f
C1784 a_n1986_8322.t11 gnd 0.09348f
C1785 a_n1986_8322.n9 gnd 0.658471f
C1786 a_n1986_8322.n10 gnd 0.373822f
C1787 a_n1986_8322.t8 gnd 0.873554f
C1788 a_n1986_8322.n11 gnd 0.871824f
C1789 a_n1986_8322.n12 gnd 1.58981f
C1790 a_n1986_8322.n13 gnd 4.0376f
C1791 a_n1986_8322.t15 gnd 0.873554f
C1792 a_n1986_8322.n14 gnd 0.766087f
C1793 a_n1986_8322.t14 gnd 0.09348f
C1794 a_n1986_8322.t23 gnd 0.09348f
C1795 a_n1986_8322.n15 gnd 0.658471f
C1796 a_n1986_8322.n16 gnd 0.373822f
C1797 a_n1986_8322.t20 gnd 0.09348f
C1798 a_n1986_8322.t17 gnd 0.09348f
C1799 a_n1986_8322.n17 gnd 0.658471f
C1800 a_n1986_8322.n18 gnd 0.735743f
C1801 a_n1986_8322.t22 gnd 0.875299f
C1802 a_n2848_n452.n0 gnd 3.415f
C1803 a_n2848_n452.n1 gnd 0.285666f
C1804 a_n2848_n452.n2 gnd 0.492471f
C1805 a_n2848_n452.n3 gnd 0.664435f
C1806 a_n2848_n452.n4 gnd 0.215942f
C1807 a_n2848_n452.n5 gnd 0.282512f
C1808 a_n2848_n452.n6 gnd 0.546457f
C1809 a_n2848_n452.n7 gnd 0.526038f
C1810 a_n2848_n452.n8 gnd 0.204894f
C1811 a_n2848_n452.n9 gnd 0.150908f
C1812 a_n2848_n452.n10 gnd 0.23718f
C1813 a_n2848_n452.n11 gnd 0.183194f
C1814 a_n2848_n452.n12 gnd 0.204894f
C1815 a_n2848_n452.n13 gnd 1.0063f
C1816 a_n2848_n452.n14 gnd 0.150908f
C1817 a_n2848_n452.n15 gnd 0.580023f
C1818 a_n2848_n452.n16 gnd 0.432289f
C1819 a_n2848_n452.n17 gnd 0.215942f
C1820 a_n2848_n452.n18 gnd 0.492471f
C1821 a_n2848_n452.n19 gnd 0.282512f
C1822 a_n2848_n452.n20 gnd 0.438486f
C1823 a_n2848_n452.n21 gnd 0.215942f
C1824 a_n2848_n452.n22 gnd 0.731535f
C1825 a_n2848_n452.n23 gnd 0.282512f
C1826 a_n2848_n452.n24 gnd 1.17886f
C1827 a_n2848_n452.n25 gnd 1.91568f
C1828 a_n2848_n452.n26 gnd 1.14458f
C1829 a_n2848_n452.n27 gnd 1.77783f
C1830 a_n2848_n452.n28 gnd 0.377489f
C1831 a_n2848_n452.n29 gnd 3.11576f
C1832 a_n2848_n452.n30 gnd 0.377488f
C1833 a_n2848_n452.n31 gnd 3.20158f
C1834 a_n2848_n452.n32 gnd 0.008361f
C1835 a_n2848_n452.n34 gnd 0.285666f
C1836 a_n2848_n452.n35 gnd 0.008361f
C1837 a_n2848_n452.n37 gnd 0.285666f
C1838 a_n2848_n452.n38 gnd 0.008361f
C1839 a_n2848_n452.n39 gnd 0.28526f
C1840 a_n2848_n452.n40 gnd 0.008361f
C1841 a_n2848_n452.n41 gnd 0.28526f
C1842 a_n2848_n452.n42 gnd 0.008361f
C1843 a_n2848_n452.n43 gnd 0.28526f
C1844 a_n2848_n452.n44 gnd 0.008361f
C1845 a_n2848_n452.n45 gnd 0.28526f
C1846 a_n2848_n452.n47 gnd 0.285666f
C1847 a_n2848_n452.n48 gnd 0.008361f
C1848 a_n2848_n452.n50 gnd 0.285666f
C1849 a_n2848_n452.t27 gnd 0.14978f
C1850 a_n2848_n452.t40 gnd 0.708223f
C1851 a_n2848_n452.t24 gnd 0.696704f
C1852 a_n2848_n452.t26 gnd 0.696704f
C1853 a_n2848_n452.t18 gnd 0.116496f
C1854 a_n2848_n452.t10 gnd 0.116496f
C1855 a_n2848_n452.n52 gnd 1.03243f
C1856 a_n2848_n452.t1 gnd 0.116496f
C1857 a_n2848_n452.t5 gnd 0.116496f
C1858 a_n2848_n452.n53 gnd 1.0294f
C1859 a_n2848_n452.n54 gnd 0.912817f
C1860 a_n2848_n452.t20 gnd 0.116496f
C1861 a_n2848_n452.t22 gnd 0.116496f
C1862 a_n2848_n452.n55 gnd 1.0294f
C1863 a_n2848_n452.t11 gnd 0.116496f
C1864 a_n2848_n452.t6 gnd 0.116496f
C1865 a_n2848_n452.n56 gnd 1.03243f
C1866 a_n2848_n452.t7 gnd 0.116496f
C1867 a_n2848_n452.t12 gnd 0.116496f
C1868 a_n2848_n452.n57 gnd 1.0294f
C1869 a_n2848_n452.n58 gnd 0.912817f
C1870 a_n2848_n452.t17 gnd 0.116496f
C1871 a_n2848_n452.t14 gnd 0.116496f
C1872 a_n2848_n452.n59 gnd 1.0294f
C1873 a_n2848_n452.t2 gnd 0.116496f
C1874 a_n2848_n452.t15 gnd 0.116496f
C1875 a_n2848_n452.n60 gnd 1.0294f
C1876 a_n2848_n452.n61 gnd 3.15028f
C1877 a_n2848_n452.t16 gnd 0.116496f
C1878 a_n2848_n452.t13 gnd 0.116496f
C1879 a_n2848_n452.n62 gnd 1.0294f
C1880 a_n2848_n452.n63 gnd 0.449443f
C1881 a_n2848_n452.t23 gnd 0.116496f
C1882 a_n2848_n452.t19 gnd 0.116496f
C1883 a_n2848_n452.n64 gnd 1.0294f
C1884 a_n2848_n452.t0 gnd 0.116496f
C1885 a_n2848_n452.t21 gnd 0.116496f
C1886 a_n2848_n452.n65 gnd 1.03243f
C1887 a_n2848_n452.t8 gnd 0.116496f
C1888 a_n2848_n452.t9 gnd 0.116496f
C1889 a_n2848_n452.n66 gnd 1.0294f
C1890 a_n2848_n452.n67 gnd 0.912814f
C1891 a_n2848_n452.t3 gnd 0.116496f
C1892 a_n2848_n452.t4 gnd 0.116496f
C1893 a_n2848_n452.n68 gnd 1.0294f
C1894 a_n2848_n452.t36 gnd 0.696704f
C1895 a_n2848_n452.n69 gnd 0.302425f
C1896 a_n2848_n452.t44 gnd 0.696704f
C1897 a_n2848_n452.t30 gnd 0.708223f
C1898 a_n2848_n452.t75 gnd 0.711378f
C1899 a_n2848_n452.t58 gnd 0.696704f
C1900 a_n2848_n452.t62 gnd 0.696704f
C1901 a_n2848_n452.t52 gnd 0.696704f
C1902 a_n2848_n452.n70 gnd 0.306315f
C1903 a_n2848_n452.t67 gnd 0.696704f
C1904 a_n2848_n452.t73 gnd 0.708223f
C1905 a_n2848_n452.t39 gnd 1.40246f
C1906 a_n2848_n452.t29 gnd 0.14978f
C1907 a_n2848_n452.t33 gnd 0.14978f
C1908 a_n2848_n452.n71 gnd 1.05505f
C1909 a_n2848_n452.t47 gnd 0.14978f
C1910 a_n2848_n452.t35 gnd 0.14978f
C1911 a_n2848_n452.n72 gnd 1.05505f
C1912 a_n2848_n452.t43 gnd 1.39967f
C1913 a_n2848_n452.t46 gnd 0.696704f
C1914 a_n2848_n452.n73 gnd 0.306315f
C1915 a_n2848_n452.t34 gnd 0.696704f
C1916 a_n2848_n452.t28 gnd 0.696704f
C1917 a_n2848_n452.t56 gnd 0.696704f
C1918 a_n2848_n452.n74 gnd 0.306315f
C1919 a_n2848_n452.t65 gnd 0.696704f
C1920 a_n2848_n452.t71 gnd 0.696704f
C1921 a_n2848_n452.t70 gnd 0.711378f
C1922 a_n2848_n452.n75 gnd 0.308932f
C1923 a_n2848_n452.t50 gnd 0.696704f
C1924 a_n2848_n452.n76 gnd 0.302425f
C1925 a_n2848_n452.n77 gnd 0.308933f
C1926 a_n2848_n452.t51 gnd 0.708223f
C1927 a_n2848_n452.t38 gnd 0.711378f
C1928 a_n2848_n452.n78 gnd 0.308932f
C1929 a_n2848_n452.t32 gnd 0.696704f
C1930 a_n2848_n452.n79 gnd 0.302425f
C1931 a_n2848_n452.n80 gnd 0.308933f
C1932 a_n2848_n452.t42 gnd 0.708223f
C1933 a_n2848_n452.n81 gnd 1.13204f
C1934 a_n2848_n452.t55 gnd 0.696704f
C1935 a_n2848_n452.n82 gnd 0.302425f
C1936 a_n2848_n452.t61 gnd 0.696704f
C1937 a_n2848_n452.n83 gnd 0.302425f
C1938 a_n2848_n452.t53 gnd 0.696704f
C1939 a_n2848_n452.n84 gnd 0.302425f
C1940 a_n2848_n452.t66 gnd 0.696704f
C1941 a_n2848_n452.n85 gnd 0.302425f
C1942 a_n2848_n452.t57 gnd 0.696704f
C1943 a_n2848_n452.n86 gnd 0.296933f
C1944 a_n2848_n452.t48 gnd 0.696704f
C1945 a_n2848_n452.n87 gnd 0.306315f
C1946 a_n2848_n452.t59 gnd 0.708378f
C1947 a_n2848_n452.t68 gnd 0.696704f
C1948 a_n2848_n452.n88 gnd 0.296933f
C1949 a_n2848_n452.t54 gnd 0.696704f
C1950 a_n2848_n452.n89 gnd 0.306315f
C1951 a_n2848_n452.t63 gnd 0.708378f
C1952 a_n2848_n452.t72 gnd 0.696704f
C1953 a_n2848_n452.n90 gnd 0.296933f
C1954 a_n2848_n452.t60 gnd 0.696704f
C1955 a_n2848_n452.n91 gnd 0.306315f
C1956 a_n2848_n452.t74 gnd 0.708378f
C1957 a_n2848_n452.t64 gnd 0.696704f
C1958 a_n2848_n452.n92 gnd 0.296933f
C1959 a_n2848_n452.t49 gnd 0.696704f
C1960 a_n2848_n452.n93 gnd 0.306315f
C1961 a_n2848_n452.t69 gnd 0.708378f
C1962 a_n2848_n452.n94 gnd 1.33845f
C1963 a_n2848_n452.n95 gnd 0.308933f
C1964 a_n2848_n452.n96 gnd 0.302425f
C1965 a_n2848_n452.n97 gnd 0.308932f
C1966 a_n2848_n452.n98 gnd 0.308933f
C1967 a_n2848_n452.n99 gnd 0.01225f
C1968 a_n2848_n452.n100 gnd 0.302425f
C1969 a_n2848_n452.n101 gnd 0.308933f
C1970 a_n2848_n452.n102 gnd 0.786935f
C1971 a_n2848_n452.t41 gnd 1.39967f
C1972 a_n2848_n452.t31 gnd 1.40246f
C1973 a_n2848_n452.t37 gnd 0.14978f
C1974 a_n2848_n452.t45 gnd 0.14978f
C1975 a_n2848_n452.n103 gnd 1.05505f
C1976 a_n2848_n452.n104 gnd 1.05505f
C1977 a_n2848_n452.t25 gnd 0.14978f
C1978 vdd.t191 gnd 0.032819f
C1979 vdd.t195 gnd 0.032819f
C1980 vdd.n0 gnd 0.258853f
C1981 vdd.t28 gnd 0.032819f
C1982 vdd.t113 gnd 0.032819f
C1983 vdd.n1 gnd 0.258425f
C1984 vdd.n2 gnd 0.238317f
C1985 vdd.t197 gnd 0.032819f
C1986 vdd.t185 gnd 0.032819f
C1987 vdd.n3 gnd 0.258425f
C1988 vdd.n4 gnd 0.120526f
C1989 vdd.t115 gnd 0.032819f
C1990 vdd.t119 gnd 0.032819f
C1991 vdd.n5 gnd 0.258425f
C1992 vdd.n6 gnd 0.113091f
C1993 vdd.t30 gnd 0.032819f
C1994 vdd.t199 gnd 0.032819f
C1995 vdd.n7 gnd 0.258853f
C1996 vdd.t193 gnd 0.032819f
C1997 vdd.t117 gnd 0.032819f
C1998 vdd.n8 gnd 0.258425f
C1999 vdd.n9 gnd 0.238317f
C2000 vdd.t187 gnd 0.032819f
C2001 vdd.t20 gnd 0.032819f
C2002 vdd.n10 gnd 0.258425f
C2003 vdd.n11 gnd 0.120526f
C2004 vdd.t23 gnd 0.032819f
C2005 vdd.t189 gnd 0.032819f
C2006 vdd.n12 gnd 0.258425f
C2007 vdd.n13 gnd 0.113091f
C2008 vdd.n14 gnd 0.079954f
C2009 vdd.t14 gnd 0.018233f
C2010 vdd.t18 gnd 0.018233f
C2011 vdd.n15 gnd 0.167828f
C2012 vdd.t6 gnd 0.018233f
C2013 vdd.t17 gnd 0.018233f
C2014 vdd.n16 gnd 0.167337f
C2015 vdd.n17 gnd 0.291218f
C2016 vdd.t7 gnd 0.018233f
C2017 vdd.t13 gnd 0.018233f
C2018 vdd.n18 gnd 0.167337f
C2019 vdd.n19 gnd 0.120481f
C2020 vdd.t10 gnd 0.018233f
C2021 vdd.t11 gnd 0.018233f
C2022 vdd.n20 gnd 0.167828f
C2023 vdd.t8 gnd 0.018233f
C2024 vdd.t5 gnd 0.018233f
C2025 vdd.n21 gnd 0.167337f
C2026 vdd.n22 gnd 0.291218f
C2027 vdd.t16 gnd 0.018233f
C2028 vdd.t15 gnd 0.018233f
C2029 vdd.n23 gnd 0.167337f
C2030 vdd.n24 gnd 0.120481f
C2031 vdd.t3 gnd 0.018233f
C2032 vdd.t4 gnd 0.018233f
C2033 vdd.n25 gnd 0.167337f
C2034 vdd.t12 gnd 0.018233f
C2035 vdd.t9 gnd 0.018233f
C2036 vdd.n26 gnd 0.167337f
C2037 vdd.n27 gnd 19.652802f
C2038 vdd.n28 gnd 7.29364f
C2039 vdd.n29 gnd 0.004973f
C2040 vdd.n30 gnd 0.004615f
C2041 vdd.n31 gnd 0.002553f
C2042 vdd.n32 gnd 0.005861f
C2043 vdd.n33 gnd 0.00248f
C2044 vdd.n34 gnd 0.002626f
C2045 vdd.n35 gnd 0.004615f
C2046 vdd.n36 gnd 0.00248f
C2047 vdd.n37 gnd 0.005861f
C2048 vdd.n38 gnd 0.002626f
C2049 vdd.n39 gnd 0.004615f
C2050 vdd.n40 gnd 0.00248f
C2051 vdd.n41 gnd 0.004396f
C2052 vdd.n42 gnd 0.004409f
C2053 vdd.t123 gnd 0.012592f
C2054 vdd.n43 gnd 0.028017f
C2055 vdd.n44 gnd 0.145808f
C2056 vdd.n45 gnd 0.00248f
C2057 vdd.n46 gnd 0.002626f
C2058 vdd.n47 gnd 0.005861f
C2059 vdd.n48 gnd 0.005861f
C2060 vdd.n49 gnd 0.002626f
C2061 vdd.n50 gnd 0.00248f
C2062 vdd.n51 gnd 0.004615f
C2063 vdd.n52 gnd 0.004615f
C2064 vdd.n53 gnd 0.00248f
C2065 vdd.n54 gnd 0.002626f
C2066 vdd.n55 gnd 0.005861f
C2067 vdd.n56 gnd 0.005861f
C2068 vdd.n57 gnd 0.002626f
C2069 vdd.n58 gnd 0.00248f
C2070 vdd.n59 gnd 0.004615f
C2071 vdd.n60 gnd 0.004615f
C2072 vdd.n61 gnd 0.00248f
C2073 vdd.n62 gnd 0.002626f
C2074 vdd.n63 gnd 0.005861f
C2075 vdd.n64 gnd 0.005861f
C2076 vdd.n65 gnd 0.013857f
C2077 vdd.n66 gnd 0.002553f
C2078 vdd.n67 gnd 0.00248f
C2079 vdd.n68 gnd 0.011927f
C2080 vdd.n69 gnd 0.008327f
C2081 vdd.t175 gnd 0.029173f
C2082 vdd.t149 gnd 0.029173f
C2083 vdd.n70 gnd 0.200496f
C2084 vdd.n71 gnd 0.15766f
C2085 vdd.t182 gnd 0.029173f
C2086 vdd.t138 gnd 0.029173f
C2087 vdd.n72 gnd 0.200496f
C2088 vdd.n73 gnd 0.12723f
C2089 vdd.t168 gnd 0.029173f
C2090 vdd.t143 gnd 0.029173f
C2091 vdd.n74 gnd 0.200496f
C2092 vdd.n75 gnd 0.12723f
C2093 vdd.n76 gnd 0.004973f
C2094 vdd.n77 gnd 0.004615f
C2095 vdd.n78 gnd 0.002553f
C2096 vdd.n79 gnd 0.005861f
C2097 vdd.n80 gnd 0.00248f
C2098 vdd.n81 gnd 0.002626f
C2099 vdd.n82 gnd 0.004615f
C2100 vdd.n83 gnd 0.00248f
C2101 vdd.n84 gnd 0.005861f
C2102 vdd.n85 gnd 0.002626f
C2103 vdd.n86 gnd 0.004615f
C2104 vdd.n87 gnd 0.00248f
C2105 vdd.n88 gnd 0.004396f
C2106 vdd.n89 gnd 0.004409f
C2107 vdd.t181 gnd 0.012592f
C2108 vdd.n90 gnd 0.028017f
C2109 vdd.n91 gnd 0.145808f
C2110 vdd.n92 gnd 0.00248f
C2111 vdd.n93 gnd 0.002626f
C2112 vdd.n94 gnd 0.005861f
C2113 vdd.n95 gnd 0.005861f
C2114 vdd.n96 gnd 0.002626f
C2115 vdd.n97 gnd 0.00248f
C2116 vdd.n98 gnd 0.004615f
C2117 vdd.n99 gnd 0.004615f
C2118 vdd.n100 gnd 0.00248f
C2119 vdd.n101 gnd 0.002626f
C2120 vdd.n102 gnd 0.005861f
C2121 vdd.n103 gnd 0.005861f
C2122 vdd.n104 gnd 0.002626f
C2123 vdd.n105 gnd 0.00248f
C2124 vdd.n106 gnd 0.004615f
C2125 vdd.n107 gnd 0.004615f
C2126 vdd.n108 gnd 0.00248f
C2127 vdd.n109 gnd 0.002626f
C2128 vdd.n110 gnd 0.005861f
C2129 vdd.n111 gnd 0.005861f
C2130 vdd.n112 gnd 0.013857f
C2131 vdd.n113 gnd 0.002553f
C2132 vdd.n114 gnd 0.00248f
C2133 vdd.n115 gnd 0.011927f
C2134 vdd.n116 gnd 0.008066f
C2135 vdd.n117 gnd 0.09466f
C2136 vdd.n118 gnd 0.004973f
C2137 vdd.n119 gnd 0.004615f
C2138 vdd.n120 gnd 0.002553f
C2139 vdd.n121 gnd 0.005861f
C2140 vdd.n122 gnd 0.00248f
C2141 vdd.n123 gnd 0.002626f
C2142 vdd.n124 gnd 0.004615f
C2143 vdd.n125 gnd 0.00248f
C2144 vdd.n126 gnd 0.005861f
C2145 vdd.n127 gnd 0.002626f
C2146 vdd.n128 gnd 0.004615f
C2147 vdd.n129 gnd 0.00248f
C2148 vdd.n130 gnd 0.004396f
C2149 vdd.n131 gnd 0.004409f
C2150 vdd.t150 gnd 0.012592f
C2151 vdd.n132 gnd 0.028017f
C2152 vdd.n133 gnd 0.145808f
C2153 vdd.n134 gnd 0.00248f
C2154 vdd.n135 gnd 0.002626f
C2155 vdd.n136 gnd 0.005861f
C2156 vdd.n137 gnd 0.005861f
C2157 vdd.n138 gnd 0.002626f
C2158 vdd.n139 gnd 0.00248f
C2159 vdd.n140 gnd 0.004615f
C2160 vdd.n141 gnd 0.004615f
C2161 vdd.n142 gnd 0.00248f
C2162 vdd.n143 gnd 0.002626f
C2163 vdd.n144 gnd 0.005861f
C2164 vdd.n145 gnd 0.005861f
C2165 vdd.n146 gnd 0.002626f
C2166 vdd.n147 gnd 0.00248f
C2167 vdd.n148 gnd 0.004615f
C2168 vdd.n149 gnd 0.004615f
C2169 vdd.n150 gnd 0.00248f
C2170 vdd.n151 gnd 0.002626f
C2171 vdd.n152 gnd 0.005861f
C2172 vdd.n153 gnd 0.005861f
C2173 vdd.n154 gnd 0.013857f
C2174 vdd.n155 gnd 0.002553f
C2175 vdd.n156 gnd 0.00248f
C2176 vdd.n157 gnd 0.011927f
C2177 vdd.n158 gnd 0.008327f
C2178 vdd.t152 gnd 0.029173f
C2179 vdd.t163 gnd 0.029173f
C2180 vdd.n159 gnd 0.200496f
C2181 vdd.n160 gnd 0.15766f
C2182 vdd.t127 gnd 0.029173f
C2183 vdd.t146 gnd 0.029173f
C2184 vdd.n161 gnd 0.200496f
C2185 vdd.n162 gnd 0.12723f
C2186 vdd.t162 gnd 0.029173f
C2187 vdd.t183 gnd 0.029173f
C2188 vdd.n163 gnd 0.200496f
C2189 vdd.n164 gnd 0.12723f
C2190 vdd.n165 gnd 0.004973f
C2191 vdd.n166 gnd 0.004615f
C2192 vdd.n167 gnd 0.002553f
C2193 vdd.n168 gnd 0.005861f
C2194 vdd.n169 gnd 0.00248f
C2195 vdd.n170 gnd 0.002626f
C2196 vdd.n171 gnd 0.004615f
C2197 vdd.n172 gnd 0.00248f
C2198 vdd.n173 gnd 0.005861f
C2199 vdd.n174 gnd 0.002626f
C2200 vdd.n175 gnd 0.004615f
C2201 vdd.n176 gnd 0.00248f
C2202 vdd.n177 gnd 0.004396f
C2203 vdd.n178 gnd 0.004409f
C2204 vdd.t140 gnd 0.012592f
C2205 vdd.n179 gnd 0.028017f
C2206 vdd.n180 gnd 0.145808f
C2207 vdd.n181 gnd 0.00248f
C2208 vdd.n182 gnd 0.002626f
C2209 vdd.n183 gnd 0.005861f
C2210 vdd.n184 gnd 0.005861f
C2211 vdd.n185 gnd 0.002626f
C2212 vdd.n186 gnd 0.00248f
C2213 vdd.n187 gnd 0.004615f
C2214 vdd.n188 gnd 0.004615f
C2215 vdd.n189 gnd 0.00248f
C2216 vdd.n190 gnd 0.002626f
C2217 vdd.n191 gnd 0.005861f
C2218 vdd.n192 gnd 0.005861f
C2219 vdd.n193 gnd 0.002626f
C2220 vdd.n194 gnd 0.00248f
C2221 vdd.n195 gnd 0.004615f
C2222 vdd.n196 gnd 0.004615f
C2223 vdd.n197 gnd 0.00248f
C2224 vdd.n198 gnd 0.002626f
C2225 vdd.n199 gnd 0.005861f
C2226 vdd.n200 gnd 0.005861f
C2227 vdd.n201 gnd 0.013857f
C2228 vdd.n202 gnd 0.002553f
C2229 vdd.n203 gnd 0.00248f
C2230 vdd.n204 gnd 0.011927f
C2231 vdd.n205 gnd 0.008066f
C2232 vdd.n206 gnd 0.056313f
C2233 vdd.n207 gnd 0.202911f
C2234 vdd.n208 gnd 0.004973f
C2235 vdd.n209 gnd 0.004615f
C2236 vdd.n210 gnd 0.002553f
C2237 vdd.n211 gnd 0.005861f
C2238 vdd.n212 gnd 0.00248f
C2239 vdd.n213 gnd 0.002626f
C2240 vdd.n214 gnd 0.004615f
C2241 vdd.n215 gnd 0.00248f
C2242 vdd.n216 gnd 0.005861f
C2243 vdd.n217 gnd 0.002626f
C2244 vdd.n218 gnd 0.004615f
C2245 vdd.n219 gnd 0.00248f
C2246 vdd.n220 gnd 0.004396f
C2247 vdd.n221 gnd 0.004409f
C2248 vdd.t155 gnd 0.012592f
C2249 vdd.n222 gnd 0.028017f
C2250 vdd.n223 gnd 0.145808f
C2251 vdd.n224 gnd 0.00248f
C2252 vdd.n225 gnd 0.002626f
C2253 vdd.n226 gnd 0.005861f
C2254 vdd.n227 gnd 0.005861f
C2255 vdd.n228 gnd 0.002626f
C2256 vdd.n229 gnd 0.00248f
C2257 vdd.n230 gnd 0.004615f
C2258 vdd.n231 gnd 0.004615f
C2259 vdd.n232 gnd 0.00248f
C2260 vdd.n233 gnd 0.002626f
C2261 vdd.n234 gnd 0.005861f
C2262 vdd.n235 gnd 0.005861f
C2263 vdd.n236 gnd 0.002626f
C2264 vdd.n237 gnd 0.00248f
C2265 vdd.n238 gnd 0.004615f
C2266 vdd.n239 gnd 0.004615f
C2267 vdd.n240 gnd 0.00248f
C2268 vdd.n241 gnd 0.002626f
C2269 vdd.n242 gnd 0.005861f
C2270 vdd.n243 gnd 0.005861f
C2271 vdd.n244 gnd 0.013857f
C2272 vdd.n245 gnd 0.002553f
C2273 vdd.n246 gnd 0.00248f
C2274 vdd.n247 gnd 0.011927f
C2275 vdd.n248 gnd 0.008327f
C2276 vdd.t156 gnd 0.029173f
C2277 vdd.t172 gnd 0.029173f
C2278 vdd.n249 gnd 0.200496f
C2279 vdd.n250 gnd 0.15766f
C2280 vdd.t133 gnd 0.029173f
C2281 vdd.t154 gnd 0.029173f
C2282 vdd.n251 gnd 0.200496f
C2283 vdd.n252 gnd 0.12723f
C2284 vdd.t167 gnd 0.029173f
C2285 vdd.t131 gnd 0.029173f
C2286 vdd.n253 gnd 0.200496f
C2287 vdd.n254 gnd 0.12723f
C2288 vdd.n255 gnd 0.004973f
C2289 vdd.n256 gnd 0.004615f
C2290 vdd.n257 gnd 0.002553f
C2291 vdd.n258 gnd 0.005861f
C2292 vdd.n259 gnd 0.00248f
C2293 vdd.n260 gnd 0.002626f
C2294 vdd.n261 gnd 0.004615f
C2295 vdd.n262 gnd 0.00248f
C2296 vdd.n263 gnd 0.005861f
C2297 vdd.n264 gnd 0.002626f
C2298 vdd.n265 gnd 0.004615f
C2299 vdd.n266 gnd 0.00248f
C2300 vdd.n267 gnd 0.004396f
C2301 vdd.n268 gnd 0.004409f
C2302 vdd.t144 gnd 0.012592f
C2303 vdd.n269 gnd 0.028017f
C2304 vdd.n270 gnd 0.145808f
C2305 vdd.n271 gnd 0.00248f
C2306 vdd.n272 gnd 0.002626f
C2307 vdd.n273 gnd 0.005861f
C2308 vdd.n274 gnd 0.005861f
C2309 vdd.n275 gnd 0.002626f
C2310 vdd.n276 gnd 0.00248f
C2311 vdd.n277 gnd 0.004615f
C2312 vdd.n278 gnd 0.004615f
C2313 vdd.n279 gnd 0.00248f
C2314 vdd.n280 gnd 0.002626f
C2315 vdd.n281 gnd 0.005861f
C2316 vdd.n282 gnd 0.005861f
C2317 vdd.n283 gnd 0.002626f
C2318 vdd.n284 gnd 0.00248f
C2319 vdd.n285 gnd 0.004615f
C2320 vdd.n286 gnd 0.004615f
C2321 vdd.n287 gnd 0.00248f
C2322 vdd.n288 gnd 0.002626f
C2323 vdd.n289 gnd 0.005861f
C2324 vdd.n290 gnd 0.005861f
C2325 vdd.n291 gnd 0.013857f
C2326 vdd.n292 gnd 0.002553f
C2327 vdd.n293 gnd 0.00248f
C2328 vdd.n294 gnd 0.011927f
C2329 vdd.n295 gnd 0.008066f
C2330 vdd.n296 gnd 0.056313f
C2331 vdd.n297 gnd 0.219627f
C2332 vdd.n298 gnd 0.006964f
C2333 vdd.n299 gnd 0.009061f
C2334 vdd.n300 gnd 0.007293f
C2335 vdd.n301 gnd 0.007293f
C2336 vdd.n302 gnd 0.009061f
C2337 vdd.n303 gnd 0.009061f
C2338 vdd.n304 gnd 0.662103f
C2339 vdd.n305 gnd 0.009061f
C2340 vdd.n306 gnd 0.009061f
C2341 vdd.n307 gnd 0.009061f
C2342 vdd.n308 gnd 0.717664f
C2343 vdd.n309 gnd 0.009061f
C2344 vdd.n310 gnd 0.009061f
C2345 vdd.n311 gnd 0.009061f
C2346 vdd.n312 gnd 0.009061f
C2347 vdd.n313 gnd 0.007293f
C2348 vdd.n314 gnd 0.009061f
C2349 vdd.t130 gnd 0.463009f
C2350 vdd.n315 gnd 0.009061f
C2351 vdd.n316 gnd 0.009061f
C2352 vdd.n317 gnd 0.009061f
C2353 vdd.n318 gnd 0.926018f
C2354 vdd.n319 gnd 0.009061f
C2355 vdd.n320 gnd 0.009061f
C2356 vdd.n321 gnd 0.009061f
C2357 vdd.n322 gnd 0.009061f
C2358 vdd.n323 gnd 0.009061f
C2359 vdd.n324 gnd 0.007293f
C2360 vdd.n325 gnd 0.009061f
C2361 vdd.n326 gnd 0.009061f
C2362 vdd.n327 gnd 0.009061f
C2363 vdd.n328 gnd 0.022083f
C2364 vdd.n329 gnd 2.21318f
C2365 vdd.n330 gnd 0.022589f
C2366 vdd.n331 gnd 0.009061f
C2367 vdd.n332 gnd 0.009061f
C2368 vdd.n334 gnd 0.009061f
C2369 vdd.n335 gnd 0.009061f
C2370 vdd.n336 gnd 0.007293f
C2371 vdd.n337 gnd 0.007293f
C2372 vdd.n338 gnd 0.009061f
C2373 vdd.n339 gnd 0.009061f
C2374 vdd.n340 gnd 0.009061f
C2375 vdd.n341 gnd 0.009061f
C2376 vdd.n342 gnd 0.009061f
C2377 vdd.n343 gnd 0.009061f
C2378 vdd.n344 gnd 0.007293f
C2379 vdd.n346 gnd 0.009061f
C2380 vdd.n347 gnd 0.009061f
C2381 vdd.n348 gnd 0.009061f
C2382 vdd.n349 gnd 0.009061f
C2383 vdd.n350 gnd 0.009061f
C2384 vdd.n351 gnd 0.007293f
C2385 vdd.n353 gnd 0.009061f
C2386 vdd.n354 gnd 0.009061f
C2387 vdd.n355 gnd 0.009061f
C2388 vdd.n356 gnd 0.009061f
C2389 vdd.n357 gnd 0.009061f
C2390 vdd.n358 gnd 0.007293f
C2391 vdd.n360 gnd 0.009061f
C2392 vdd.n361 gnd 0.009061f
C2393 vdd.n362 gnd 0.009061f
C2394 vdd.n363 gnd 0.009061f
C2395 vdd.n364 gnd 0.00609f
C2396 vdd.t63 gnd 0.111477f
C2397 vdd.t62 gnd 0.119139f
C2398 vdd.t61 gnd 0.145588f
C2399 vdd.n365 gnd 0.186623f
C2400 vdd.n366 gnd 0.157527f
C2401 vdd.n368 gnd 0.009061f
C2402 vdd.n369 gnd 0.009061f
C2403 vdd.n370 gnd 0.007293f
C2404 vdd.n371 gnd 0.009061f
C2405 vdd.n373 gnd 0.009061f
C2406 vdd.n374 gnd 0.009061f
C2407 vdd.n375 gnd 0.009061f
C2408 vdd.n376 gnd 0.009061f
C2409 vdd.n377 gnd 0.007293f
C2410 vdd.n379 gnd 0.009061f
C2411 vdd.n380 gnd 0.009061f
C2412 vdd.n381 gnd 0.009061f
C2413 vdd.n382 gnd 0.009061f
C2414 vdd.n383 gnd 0.009061f
C2415 vdd.n384 gnd 0.007293f
C2416 vdd.n386 gnd 0.009061f
C2417 vdd.n387 gnd 0.009061f
C2418 vdd.n388 gnd 0.009061f
C2419 vdd.n389 gnd 0.009061f
C2420 vdd.n390 gnd 0.009061f
C2421 vdd.n391 gnd 0.007293f
C2422 vdd.n393 gnd 0.009061f
C2423 vdd.n394 gnd 0.009061f
C2424 vdd.n395 gnd 0.009061f
C2425 vdd.n396 gnd 0.009061f
C2426 vdd.n397 gnd 0.009061f
C2427 vdd.n398 gnd 0.007293f
C2428 vdd.n400 gnd 0.009061f
C2429 vdd.n401 gnd 0.009061f
C2430 vdd.n402 gnd 0.009061f
C2431 vdd.n403 gnd 0.009061f
C2432 vdd.n404 gnd 0.00722f
C2433 vdd.t57 gnd 0.111477f
C2434 vdd.t56 gnd 0.119139f
C2435 vdd.t54 gnd 0.145588f
C2436 vdd.n405 gnd 0.186623f
C2437 vdd.n406 gnd 0.157527f
C2438 vdd.n408 gnd 0.009061f
C2439 vdd.n409 gnd 0.009061f
C2440 vdd.n410 gnd 0.007293f
C2441 vdd.n411 gnd 0.009061f
C2442 vdd.n413 gnd 0.009061f
C2443 vdd.n414 gnd 0.009061f
C2444 vdd.n415 gnd 0.009061f
C2445 vdd.n416 gnd 0.009061f
C2446 vdd.n417 gnd 0.007293f
C2447 vdd.n419 gnd 0.009061f
C2448 vdd.n420 gnd 0.009061f
C2449 vdd.n421 gnd 0.009061f
C2450 vdd.n422 gnd 0.009061f
C2451 vdd.n423 gnd 0.009061f
C2452 vdd.n424 gnd 0.007293f
C2453 vdd.n426 gnd 0.009061f
C2454 vdd.n427 gnd 0.009061f
C2455 vdd.n428 gnd 0.009061f
C2456 vdd.n429 gnd 0.009061f
C2457 vdd.n430 gnd 0.009061f
C2458 vdd.n431 gnd 0.007293f
C2459 vdd.n433 gnd 0.009061f
C2460 vdd.n434 gnd 0.009061f
C2461 vdd.n435 gnd 0.009061f
C2462 vdd.n436 gnd 0.009061f
C2463 vdd.n437 gnd 0.009061f
C2464 vdd.n438 gnd 0.007293f
C2465 vdd.n440 gnd 0.009061f
C2466 vdd.n441 gnd 0.009061f
C2467 vdd.n442 gnd 0.009061f
C2468 vdd.n443 gnd 0.009061f
C2469 vdd.n444 gnd 0.009061f
C2470 vdd.n445 gnd 0.009061f
C2471 vdd.n446 gnd 0.007293f
C2472 vdd.n447 gnd 0.009061f
C2473 vdd.n448 gnd 0.009061f
C2474 vdd.n449 gnd 0.007293f
C2475 vdd.n450 gnd 0.009061f
C2476 vdd.n451 gnd 0.007293f
C2477 vdd.n452 gnd 0.009061f
C2478 vdd.n453 gnd 0.007293f
C2479 vdd.n454 gnd 0.009061f
C2480 vdd.n455 gnd 0.009061f
C2481 vdd.n456 gnd 0.50468f
C2482 vdd.t126 gnd 0.463009f
C2483 vdd.n457 gnd 0.009061f
C2484 vdd.n458 gnd 0.007293f
C2485 vdd.n459 gnd 0.009061f
C2486 vdd.n460 gnd 0.007293f
C2487 vdd.n461 gnd 0.009061f
C2488 vdd.t151 gnd 0.463009f
C2489 vdd.n462 gnd 0.009061f
C2490 vdd.n463 gnd 0.007293f
C2491 vdd.n464 gnd 0.009061f
C2492 vdd.n465 gnd 0.007293f
C2493 vdd.n466 gnd 0.009061f
C2494 vdd.t122 gnd 0.463009f
C2495 vdd.n467 gnd 0.578761f
C2496 vdd.n468 gnd 0.009061f
C2497 vdd.n469 gnd 0.007293f
C2498 vdd.n470 gnd 0.009061f
C2499 vdd.n471 gnd 0.007293f
C2500 vdd.n472 gnd 0.009061f
C2501 vdd.n473 gnd 0.926018f
C2502 vdd.n474 gnd 0.009061f
C2503 vdd.n475 gnd 0.007293f
C2504 vdd.n476 gnd 0.022083f
C2505 vdd.n477 gnd 0.006053f
C2506 vdd.n478 gnd 0.022083f
C2507 vdd.t33 gnd 0.463009f
C2508 vdd.n479 gnd 0.022083f
C2509 vdd.n480 gnd 0.006053f
C2510 vdd.n481 gnd 0.007793f
C2511 vdd.n482 gnd 0.007293f
C2512 vdd.n483 gnd 0.009061f
C2513 vdd.n484 gnd 6.38027f
C2514 vdd.n515 gnd 0.022589f
C2515 vdd.n516 gnd 1.27328f
C2516 vdd.n517 gnd 0.009061f
C2517 vdd.n518 gnd 0.007293f
C2518 vdd.n519 gnd 0.005799f
C2519 vdd.n520 gnd 0.014807f
C2520 vdd.n521 gnd 0.007293f
C2521 vdd.n522 gnd 0.009061f
C2522 vdd.n523 gnd 0.009061f
C2523 vdd.n524 gnd 0.009061f
C2524 vdd.n525 gnd 0.009061f
C2525 vdd.n526 gnd 0.009061f
C2526 vdd.n527 gnd 0.009061f
C2527 vdd.n528 gnd 0.009061f
C2528 vdd.n529 gnd 0.009061f
C2529 vdd.n530 gnd 0.009061f
C2530 vdd.n531 gnd 0.009061f
C2531 vdd.n532 gnd 0.009061f
C2532 vdd.n533 gnd 0.009061f
C2533 vdd.n534 gnd 0.009061f
C2534 vdd.n535 gnd 0.009061f
C2535 vdd.n536 gnd 0.00609f
C2536 vdd.n537 gnd 0.009061f
C2537 vdd.n538 gnd 0.009061f
C2538 vdd.n539 gnd 0.009061f
C2539 vdd.n540 gnd 0.009061f
C2540 vdd.n541 gnd 0.009061f
C2541 vdd.n542 gnd 0.009061f
C2542 vdd.n543 gnd 0.009061f
C2543 vdd.n544 gnd 0.009061f
C2544 vdd.n545 gnd 0.009061f
C2545 vdd.n546 gnd 0.009061f
C2546 vdd.n547 gnd 0.009061f
C2547 vdd.n548 gnd 0.009061f
C2548 vdd.n549 gnd 0.009061f
C2549 vdd.n550 gnd 0.009061f
C2550 vdd.n551 gnd 0.009061f
C2551 vdd.n552 gnd 0.009061f
C2552 vdd.n553 gnd 0.009061f
C2553 vdd.n554 gnd 0.009061f
C2554 vdd.n555 gnd 0.009061f
C2555 vdd.n556 gnd 0.00722f
C2556 vdd.t34 gnd 0.111477f
C2557 vdd.t35 gnd 0.119139f
C2558 vdd.t32 gnd 0.145588f
C2559 vdd.n557 gnd 0.186623f
C2560 vdd.n558 gnd 0.156797f
C2561 vdd.n559 gnd 0.009061f
C2562 vdd.n560 gnd 0.009061f
C2563 vdd.n561 gnd 0.009061f
C2564 vdd.n562 gnd 0.009061f
C2565 vdd.n563 gnd 0.009061f
C2566 vdd.n564 gnd 0.009061f
C2567 vdd.n565 gnd 0.009061f
C2568 vdd.n566 gnd 0.009061f
C2569 vdd.n567 gnd 0.009061f
C2570 vdd.n568 gnd 0.009061f
C2571 vdd.n569 gnd 0.009061f
C2572 vdd.n570 gnd 0.009061f
C2573 vdd.n571 gnd 0.009061f
C2574 vdd.n572 gnd 0.005799f
C2575 vdd.n575 gnd 0.006162f
C2576 vdd.n576 gnd 0.006162f
C2577 vdd.n577 gnd 0.006162f
C2578 vdd.n578 gnd 0.006162f
C2579 vdd.n579 gnd 0.006162f
C2580 vdd.n580 gnd 0.006162f
C2581 vdd.n582 gnd 0.006162f
C2582 vdd.n583 gnd 0.006162f
C2583 vdd.n585 gnd 0.006162f
C2584 vdd.n586 gnd 0.004485f
C2585 vdd.n588 gnd 0.006162f
C2586 vdd.t78 gnd 0.248992f
C2587 vdd.t77 gnd 0.254874f
C2588 vdd.t76 gnd 0.162551f
C2589 vdd.n589 gnd 0.08785f
C2590 vdd.n590 gnd 0.049831f
C2591 vdd.n591 gnd 0.008806f
C2592 vdd.n592 gnd 0.014401f
C2593 vdd.n594 gnd 0.006162f
C2594 vdd.n595 gnd 0.629692f
C2595 vdd.n596 gnd 0.013651f
C2596 vdd.n597 gnd 0.013651f
C2597 vdd.n598 gnd 0.006162f
C2598 vdd.n599 gnd 0.014621f
C2599 vdd.n600 gnd 0.006162f
C2600 vdd.n601 gnd 0.006162f
C2601 vdd.n602 gnd 0.006162f
C2602 vdd.n603 gnd 0.006162f
C2603 vdd.n604 gnd 0.006162f
C2604 vdd.n606 gnd 0.006162f
C2605 vdd.n607 gnd 0.006162f
C2606 vdd.n609 gnd 0.006162f
C2607 vdd.n610 gnd 0.006162f
C2608 vdd.n612 gnd 0.006162f
C2609 vdd.n613 gnd 0.006162f
C2610 vdd.n615 gnd 0.006162f
C2611 vdd.n616 gnd 0.006162f
C2612 vdd.n618 gnd 0.006162f
C2613 vdd.n619 gnd 0.006162f
C2614 vdd.n621 gnd 0.006162f
C2615 vdd.t71 gnd 0.248992f
C2616 vdd.t70 gnd 0.254874f
C2617 vdd.t68 gnd 0.162551f
C2618 vdd.n622 gnd 0.08785f
C2619 vdd.n623 gnd 0.049831f
C2620 vdd.n624 gnd 0.006162f
C2621 vdd.n626 gnd 0.006162f
C2622 vdd.n627 gnd 0.006162f
C2623 vdd.t69 gnd 0.314846f
C2624 vdd.n628 gnd 0.006162f
C2625 vdd.n629 gnd 0.006162f
C2626 vdd.n630 gnd 0.006162f
C2627 vdd.n631 gnd 0.006162f
C2628 vdd.n632 gnd 0.006162f
C2629 vdd.n633 gnd 0.629692f
C2630 vdd.n634 gnd 0.006162f
C2631 vdd.n635 gnd 0.006162f
C2632 vdd.n636 gnd 0.550981f
C2633 vdd.n637 gnd 0.006162f
C2634 vdd.n638 gnd 0.006162f
C2635 vdd.n639 gnd 0.005437f
C2636 vdd.n640 gnd 0.006162f
C2637 vdd.n641 gnd 0.555611f
C2638 vdd.n642 gnd 0.006162f
C2639 vdd.n643 gnd 0.006162f
C2640 vdd.n644 gnd 0.006162f
C2641 vdd.n645 gnd 0.006162f
C2642 vdd.n646 gnd 0.006162f
C2643 vdd.n647 gnd 0.629692f
C2644 vdd.n648 gnd 0.006162f
C2645 vdd.n649 gnd 0.006162f
C2646 vdd.t48 gnd 0.282436f
C2647 vdd.t24 gnd 0.074081f
C2648 vdd.n650 gnd 0.006162f
C2649 vdd.n651 gnd 0.006162f
C2650 vdd.n652 gnd 0.006162f
C2651 vdd.t2 gnd 0.314846f
C2652 vdd.n653 gnd 0.006162f
C2653 vdd.n654 gnd 0.006162f
C2654 vdd.n655 gnd 0.006162f
C2655 vdd.n656 gnd 0.006162f
C2656 vdd.n657 gnd 0.006162f
C2657 vdd.t26 gnd 0.314846f
C2658 vdd.n658 gnd 0.006162f
C2659 vdd.n659 gnd 0.006162f
C2660 vdd.n660 gnd 0.5232f
C2661 vdd.n661 gnd 0.006162f
C2662 vdd.n662 gnd 0.006162f
C2663 vdd.n663 gnd 0.006162f
C2664 vdd.n664 gnd 0.384298f
C2665 vdd.n665 gnd 0.006162f
C2666 vdd.n666 gnd 0.006162f
C2667 vdd.t198 gnd 0.314846f
C2668 vdd.n667 gnd 0.006162f
C2669 vdd.n668 gnd 0.006162f
C2670 vdd.n669 gnd 0.006162f
C2671 vdd.n670 gnd 0.5232f
C2672 vdd.n671 gnd 0.006162f
C2673 vdd.n672 gnd 0.006162f
C2674 vdd.t108 gnd 0.268545f
C2675 vdd.t29 gnd 0.245395f
C2676 vdd.n673 gnd 0.006162f
C2677 vdd.n674 gnd 0.006162f
C2678 vdd.n675 gnd 0.006162f
C2679 vdd.t116 gnd 0.314846f
C2680 vdd.n676 gnd 0.006162f
C2681 vdd.n677 gnd 0.006162f
C2682 vdd.t1 gnd 0.314846f
C2683 vdd.n678 gnd 0.006162f
C2684 vdd.n679 gnd 0.006162f
C2685 vdd.n680 gnd 0.006162f
C2686 vdd.t21 gnd 0.231505f
C2687 vdd.n681 gnd 0.006162f
C2688 vdd.n682 gnd 0.006162f
C2689 vdd.n683 gnd 0.537091f
C2690 vdd.n684 gnd 0.006162f
C2691 vdd.n685 gnd 0.006162f
C2692 vdd.n686 gnd 0.006162f
C2693 vdd.n687 gnd 0.629692f
C2694 vdd.n688 gnd 0.006162f
C2695 vdd.n689 gnd 0.006162f
C2696 vdd.t192 gnd 0.282436f
C2697 vdd.n690 gnd 0.398188f
C2698 vdd.n691 gnd 0.006162f
C2699 vdd.n692 gnd 0.006162f
C2700 vdd.n693 gnd 0.006162f
C2701 vdd.t19 gnd 0.314846f
C2702 vdd.n694 gnd 0.006162f
C2703 vdd.n695 gnd 0.006162f
C2704 vdd.n696 gnd 0.006162f
C2705 vdd.n697 gnd 0.006162f
C2706 vdd.n698 gnd 0.006162f
C2707 vdd.t186 gnd 0.629692f
C2708 vdd.n699 gnd 0.006162f
C2709 vdd.n700 gnd 0.006162f
C2710 vdd.t73 gnd 0.314846f
C2711 vdd.n701 gnd 0.006162f
C2712 vdd.n702 gnd 0.014621f
C2713 vdd.n703 gnd 0.014621f
C2714 vdd.t188 gnd 0.592652f
C2715 vdd.n704 gnd 0.013651f
C2716 vdd.n705 gnd 0.013651f
C2717 vdd.n706 gnd 0.014621f
C2718 vdd.n707 gnd 0.006162f
C2719 vdd.n708 gnd 0.006162f
C2720 vdd.t114 gnd 0.592652f
C2721 vdd.n726 gnd 0.014621f
C2722 vdd.n744 gnd 0.013651f
C2723 vdd.n745 gnd 0.006162f
C2724 vdd.n746 gnd 0.013651f
C2725 vdd.t98 gnd 0.248992f
C2726 vdd.t97 gnd 0.254874f
C2727 vdd.t96 gnd 0.162551f
C2728 vdd.n747 gnd 0.08785f
C2729 vdd.n748 gnd 0.049831f
C2730 vdd.n749 gnd 0.014401f
C2731 vdd.n750 gnd 0.006162f
C2732 vdd.t184 gnd 0.629692f
C2733 vdd.n751 gnd 0.013651f
C2734 vdd.n752 gnd 0.006162f
C2735 vdd.n753 gnd 0.014621f
C2736 vdd.n754 gnd 0.006162f
C2737 vdd.t67 gnd 0.248992f
C2738 vdd.t66 gnd 0.254874f
C2739 vdd.t64 gnd 0.162551f
C2740 vdd.n755 gnd 0.08785f
C2741 vdd.n756 gnd 0.049831f
C2742 vdd.n757 gnd 0.008806f
C2743 vdd.n758 gnd 0.006162f
C2744 vdd.n759 gnd 0.006162f
C2745 vdd.t65 gnd 0.314846f
C2746 vdd.n760 gnd 0.006162f
C2747 vdd.n761 gnd 0.006162f
C2748 vdd.n762 gnd 0.006162f
C2749 vdd.n763 gnd 0.006162f
C2750 vdd.n764 gnd 0.006162f
C2751 vdd.n765 gnd 0.006162f
C2752 vdd.n766 gnd 0.629692f
C2753 vdd.n767 gnd 0.006162f
C2754 vdd.n768 gnd 0.006162f
C2755 vdd.t196 gnd 0.314846f
C2756 vdd.n769 gnd 0.006162f
C2757 vdd.n770 gnd 0.006162f
C2758 vdd.n771 gnd 0.006162f
C2759 vdd.n772 gnd 0.006162f
C2760 vdd.n773 gnd 0.398188f
C2761 vdd.n774 gnd 0.006162f
C2762 vdd.n775 gnd 0.006162f
C2763 vdd.n776 gnd 0.006162f
C2764 vdd.n777 gnd 0.006162f
C2765 vdd.n778 gnd 0.006162f
C2766 vdd.n779 gnd 0.537091f
C2767 vdd.n780 gnd 0.006162f
C2768 vdd.n781 gnd 0.006162f
C2769 vdd.t112 gnd 0.282436f
C2770 vdd.t111 gnd 0.231505f
C2771 vdd.n782 gnd 0.006162f
C2772 vdd.n783 gnd 0.006162f
C2773 vdd.n784 gnd 0.006162f
C2774 vdd.t25 gnd 0.314846f
C2775 vdd.n785 gnd 0.006162f
C2776 vdd.n786 gnd 0.006162f
C2777 vdd.t27 gnd 0.314846f
C2778 vdd.n787 gnd 0.006162f
C2779 vdd.n788 gnd 0.006162f
C2780 vdd.n789 gnd 0.006162f
C2781 vdd.t194 gnd 0.245395f
C2782 vdd.n790 gnd 0.006162f
C2783 vdd.n791 gnd 0.006162f
C2784 vdd.n792 gnd 0.5232f
C2785 vdd.n793 gnd 0.006162f
C2786 vdd.n794 gnd 0.006162f
C2787 vdd.n795 gnd 0.006162f
C2788 vdd.t190 gnd 0.314846f
C2789 vdd.n796 gnd 0.006162f
C2790 vdd.n797 gnd 0.006162f
C2791 vdd.t31 gnd 0.268545f
C2792 vdd.n798 gnd 0.384298f
C2793 vdd.n799 gnd 0.006162f
C2794 vdd.n800 gnd 0.006162f
C2795 vdd.n801 gnd 0.006162f
C2796 vdd.n802 gnd 0.5232f
C2797 vdd.n803 gnd 0.006162f
C2798 vdd.n804 gnd 0.006162f
C2799 vdd.t0 gnd 0.314846f
C2800 vdd.n805 gnd 0.006162f
C2801 vdd.n806 gnd 0.006162f
C2802 vdd.n807 gnd 0.006162f
C2803 vdd.n808 gnd 0.629692f
C2804 vdd.n809 gnd 0.006162f
C2805 vdd.n810 gnd 0.006162f
C2806 vdd.t110 gnd 0.314846f
C2807 vdd.n811 gnd 0.006162f
C2808 vdd.n812 gnd 0.006162f
C2809 vdd.n813 gnd 0.006162f
C2810 vdd.t109 gnd 0.074081f
C2811 vdd.n814 gnd 0.006162f
C2812 vdd.n815 gnd 0.006162f
C2813 vdd.n816 gnd 0.006162f
C2814 vdd.t85 gnd 0.254874f
C2815 vdd.t83 gnd 0.162551f
C2816 vdd.t86 gnd 0.254874f
C2817 vdd.n817 gnd 0.14325f
C2818 vdd.n818 gnd 0.006162f
C2819 vdd.n819 gnd 0.006162f
C2820 vdd.n820 gnd 0.629692f
C2821 vdd.n821 gnd 0.006162f
C2822 vdd.n822 gnd 0.006162f
C2823 vdd.t84 gnd 0.282436f
C2824 vdd.n823 gnd 0.555611f
C2825 vdd.n824 gnd 0.006162f
C2826 vdd.n825 gnd 0.006162f
C2827 vdd.n826 gnd 0.006162f
C2828 vdd.n827 gnd 0.550981f
C2829 vdd.n828 gnd 0.006162f
C2830 vdd.n829 gnd 0.006162f
C2831 vdd.n830 gnd 0.006162f
C2832 vdd.n831 gnd 0.006162f
C2833 vdd.n832 gnd 0.006162f
C2834 vdd.n833 gnd 0.629692f
C2835 vdd.n834 gnd 0.006162f
C2836 vdd.n835 gnd 0.006162f
C2837 vdd.t80 gnd 0.314846f
C2838 vdd.n836 gnd 0.006162f
C2839 vdd.n837 gnd 0.014621f
C2840 vdd.n838 gnd 0.014621f
C2841 vdd.n839 gnd 6.38027f
C2842 vdd.n840 gnd 0.013651f
C2843 vdd.n841 gnd 0.013651f
C2844 vdd.n842 gnd 0.014621f
C2845 vdd.n843 gnd 0.006162f
C2846 vdd.n844 gnd 0.006162f
C2847 vdd.n845 gnd 0.006162f
C2848 vdd.n846 gnd 0.006162f
C2849 vdd.n847 gnd 0.006162f
C2850 vdd.n848 gnd 0.006162f
C2851 vdd.n849 gnd 0.006162f
C2852 vdd.n850 gnd 0.006162f
C2853 vdd.n852 gnd 0.006162f
C2854 vdd.n853 gnd 0.006162f
C2855 vdd.n854 gnd 0.005799f
C2856 vdd.n857 gnd 0.022589f
C2857 vdd.n858 gnd 0.007293f
C2858 vdd.n859 gnd 0.009061f
C2859 vdd.n861 gnd 0.009061f
C2860 vdd.n862 gnd 0.006053f
C2861 vdd.t40 gnd 0.463009f
C2862 vdd.n863 gnd 6.71363f
C2863 vdd.n864 gnd 0.009061f
C2864 vdd.n865 gnd 0.022589f
C2865 vdd.n866 gnd 0.007293f
C2866 vdd.n867 gnd 0.009061f
C2867 vdd.n868 gnd 0.007293f
C2868 vdd.n869 gnd 0.009061f
C2869 vdd.n870 gnd 0.926018f
C2870 vdd.n871 gnd 0.009061f
C2871 vdd.n872 gnd 0.007293f
C2872 vdd.n873 gnd 0.007293f
C2873 vdd.n874 gnd 0.009061f
C2874 vdd.n875 gnd 0.007293f
C2875 vdd.n876 gnd 0.009061f
C2876 vdd.t120 gnd 0.463009f
C2877 vdd.n877 gnd 0.009061f
C2878 vdd.n878 gnd 0.007293f
C2879 vdd.n879 gnd 0.009061f
C2880 vdd.n880 gnd 0.007293f
C2881 vdd.n881 gnd 0.009061f
C2882 vdd.t173 gnd 0.463009f
C2883 vdd.n882 gnd 0.009061f
C2884 vdd.n883 gnd 0.007293f
C2885 vdd.n884 gnd 0.009061f
C2886 vdd.n885 gnd 0.007293f
C2887 vdd.n886 gnd 0.009061f
C2888 vdd.n887 gnd 0.726924f
C2889 vdd.n888 gnd 0.768595f
C2890 vdd.t128 gnd 0.463009f
C2891 vdd.n889 gnd 0.009061f
C2892 vdd.n890 gnd 0.007293f
C2893 vdd.n891 gnd 0.004973f
C2894 vdd.n892 gnd 0.004615f
C2895 vdd.n893 gnd 0.002553f
C2896 vdd.n894 gnd 0.005861f
C2897 vdd.n895 gnd 0.00248f
C2898 vdd.n896 gnd 0.002626f
C2899 vdd.n897 gnd 0.004615f
C2900 vdd.n898 gnd 0.00248f
C2901 vdd.n899 gnd 0.005861f
C2902 vdd.n900 gnd 0.002626f
C2903 vdd.n901 gnd 0.004615f
C2904 vdd.n902 gnd 0.00248f
C2905 vdd.n903 gnd 0.004396f
C2906 vdd.n904 gnd 0.004409f
C2907 vdd.t121 gnd 0.012592f
C2908 vdd.n905 gnd 0.028017f
C2909 vdd.n906 gnd 0.145808f
C2910 vdd.n907 gnd 0.00248f
C2911 vdd.n908 gnd 0.002626f
C2912 vdd.n909 gnd 0.005861f
C2913 vdd.n910 gnd 0.005861f
C2914 vdd.n911 gnd 0.002626f
C2915 vdd.n912 gnd 0.00248f
C2916 vdd.n913 gnd 0.004615f
C2917 vdd.n914 gnd 0.004615f
C2918 vdd.n915 gnd 0.00248f
C2919 vdd.n916 gnd 0.002626f
C2920 vdd.n917 gnd 0.005861f
C2921 vdd.n918 gnd 0.005861f
C2922 vdd.n919 gnd 0.002626f
C2923 vdd.n920 gnd 0.00248f
C2924 vdd.n921 gnd 0.004615f
C2925 vdd.n922 gnd 0.004615f
C2926 vdd.n923 gnd 0.00248f
C2927 vdd.n924 gnd 0.002626f
C2928 vdd.n925 gnd 0.005861f
C2929 vdd.n926 gnd 0.005861f
C2930 vdd.n927 gnd 0.013857f
C2931 vdd.n928 gnd 0.002553f
C2932 vdd.n929 gnd 0.00248f
C2933 vdd.n930 gnd 0.011927f
C2934 vdd.n931 gnd 0.008327f
C2935 vdd.t147 gnd 0.029173f
C2936 vdd.t176 gnd 0.029173f
C2937 vdd.n932 gnd 0.200496f
C2938 vdd.n933 gnd 0.15766f
C2939 vdd.t136 gnd 0.029173f
C2940 vdd.t164 gnd 0.029173f
C2941 vdd.n934 gnd 0.200496f
C2942 vdd.n935 gnd 0.12723f
C2943 vdd.t142 gnd 0.029173f
C2944 vdd.t170 gnd 0.029173f
C2945 vdd.n936 gnd 0.200496f
C2946 vdd.n937 gnd 0.12723f
C2947 vdd.n938 gnd 0.004973f
C2948 vdd.n939 gnd 0.004615f
C2949 vdd.n940 gnd 0.002553f
C2950 vdd.n941 gnd 0.005861f
C2951 vdd.n942 gnd 0.00248f
C2952 vdd.n943 gnd 0.002626f
C2953 vdd.n944 gnd 0.004615f
C2954 vdd.n945 gnd 0.00248f
C2955 vdd.n946 gnd 0.005861f
C2956 vdd.n947 gnd 0.002626f
C2957 vdd.n948 gnd 0.004615f
C2958 vdd.n949 gnd 0.00248f
C2959 vdd.n950 gnd 0.004396f
C2960 vdd.n951 gnd 0.004409f
C2961 vdd.t180 gnd 0.012592f
C2962 vdd.n952 gnd 0.028017f
C2963 vdd.n953 gnd 0.145808f
C2964 vdd.n954 gnd 0.00248f
C2965 vdd.n955 gnd 0.002626f
C2966 vdd.n956 gnd 0.005861f
C2967 vdd.n957 gnd 0.005861f
C2968 vdd.n958 gnd 0.002626f
C2969 vdd.n959 gnd 0.00248f
C2970 vdd.n960 gnd 0.004615f
C2971 vdd.n961 gnd 0.004615f
C2972 vdd.n962 gnd 0.00248f
C2973 vdd.n963 gnd 0.002626f
C2974 vdd.n964 gnd 0.005861f
C2975 vdd.n965 gnd 0.005861f
C2976 vdd.n966 gnd 0.002626f
C2977 vdd.n967 gnd 0.00248f
C2978 vdd.n968 gnd 0.004615f
C2979 vdd.n969 gnd 0.004615f
C2980 vdd.n970 gnd 0.00248f
C2981 vdd.n971 gnd 0.002626f
C2982 vdd.n972 gnd 0.005861f
C2983 vdd.n973 gnd 0.005861f
C2984 vdd.n974 gnd 0.013857f
C2985 vdd.n975 gnd 0.002553f
C2986 vdd.n976 gnd 0.00248f
C2987 vdd.n977 gnd 0.011927f
C2988 vdd.n978 gnd 0.008066f
C2989 vdd.n979 gnd 0.09466f
C2990 vdd.n980 gnd 0.004973f
C2991 vdd.n981 gnd 0.004615f
C2992 vdd.n982 gnd 0.002553f
C2993 vdd.n983 gnd 0.005861f
C2994 vdd.n984 gnd 0.00248f
C2995 vdd.n985 gnd 0.002626f
C2996 vdd.n986 gnd 0.004615f
C2997 vdd.n987 gnd 0.00248f
C2998 vdd.n988 gnd 0.005861f
C2999 vdd.n989 gnd 0.002626f
C3000 vdd.n990 gnd 0.004615f
C3001 vdd.n991 gnd 0.00248f
C3002 vdd.n992 gnd 0.004396f
C3003 vdd.n993 gnd 0.004409f
C3004 vdd.t171 gnd 0.012592f
C3005 vdd.n994 gnd 0.028017f
C3006 vdd.n995 gnd 0.145808f
C3007 vdd.n996 gnd 0.00248f
C3008 vdd.n997 gnd 0.002626f
C3009 vdd.n998 gnd 0.005861f
C3010 vdd.n999 gnd 0.005861f
C3011 vdd.n1000 gnd 0.002626f
C3012 vdd.n1001 gnd 0.00248f
C3013 vdd.n1002 gnd 0.004615f
C3014 vdd.n1003 gnd 0.004615f
C3015 vdd.n1004 gnd 0.00248f
C3016 vdd.n1005 gnd 0.002626f
C3017 vdd.n1006 gnd 0.005861f
C3018 vdd.n1007 gnd 0.005861f
C3019 vdd.n1008 gnd 0.002626f
C3020 vdd.n1009 gnd 0.00248f
C3021 vdd.n1010 gnd 0.004615f
C3022 vdd.n1011 gnd 0.004615f
C3023 vdd.n1012 gnd 0.00248f
C3024 vdd.n1013 gnd 0.002626f
C3025 vdd.n1014 gnd 0.005861f
C3026 vdd.n1015 gnd 0.005861f
C3027 vdd.n1016 gnd 0.013857f
C3028 vdd.n1017 gnd 0.002553f
C3029 vdd.n1018 gnd 0.00248f
C3030 vdd.n1019 gnd 0.011927f
C3031 vdd.n1020 gnd 0.008327f
C3032 vdd.t129 gnd 0.029173f
C3033 vdd.t174 gnd 0.029173f
C3034 vdd.n1021 gnd 0.200496f
C3035 vdd.n1022 gnd 0.15766f
C3036 vdd.t169 gnd 0.029173f
C3037 vdd.t160 gnd 0.029173f
C3038 vdd.n1023 gnd 0.200496f
C3039 vdd.n1024 gnd 0.12723f
C3040 vdd.t145 gnd 0.029173f
C3041 vdd.t125 gnd 0.029173f
C3042 vdd.n1025 gnd 0.200496f
C3043 vdd.n1026 gnd 0.12723f
C3044 vdd.n1027 gnd 0.004973f
C3045 vdd.n1028 gnd 0.004615f
C3046 vdd.n1029 gnd 0.002553f
C3047 vdd.n1030 gnd 0.005861f
C3048 vdd.n1031 gnd 0.00248f
C3049 vdd.n1032 gnd 0.002626f
C3050 vdd.n1033 gnd 0.004615f
C3051 vdd.n1034 gnd 0.00248f
C3052 vdd.n1035 gnd 0.005861f
C3053 vdd.n1036 gnd 0.002626f
C3054 vdd.n1037 gnd 0.004615f
C3055 vdd.n1038 gnd 0.00248f
C3056 vdd.n1039 gnd 0.004396f
C3057 vdd.n1040 gnd 0.004409f
C3058 vdd.t158 gnd 0.012592f
C3059 vdd.n1041 gnd 0.028017f
C3060 vdd.n1042 gnd 0.145808f
C3061 vdd.n1043 gnd 0.00248f
C3062 vdd.n1044 gnd 0.002626f
C3063 vdd.n1045 gnd 0.005861f
C3064 vdd.n1046 gnd 0.005861f
C3065 vdd.n1047 gnd 0.002626f
C3066 vdd.n1048 gnd 0.00248f
C3067 vdd.n1049 gnd 0.004615f
C3068 vdd.n1050 gnd 0.004615f
C3069 vdd.n1051 gnd 0.00248f
C3070 vdd.n1052 gnd 0.002626f
C3071 vdd.n1053 gnd 0.005861f
C3072 vdd.n1054 gnd 0.005861f
C3073 vdd.n1055 gnd 0.002626f
C3074 vdd.n1056 gnd 0.00248f
C3075 vdd.n1057 gnd 0.004615f
C3076 vdd.n1058 gnd 0.004615f
C3077 vdd.n1059 gnd 0.00248f
C3078 vdd.n1060 gnd 0.002626f
C3079 vdd.n1061 gnd 0.005861f
C3080 vdd.n1062 gnd 0.005861f
C3081 vdd.n1063 gnd 0.013857f
C3082 vdd.n1064 gnd 0.002553f
C3083 vdd.n1065 gnd 0.00248f
C3084 vdd.n1066 gnd 0.011927f
C3085 vdd.n1067 gnd 0.008066f
C3086 vdd.n1068 gnd 0.056313f
C3087 vdd.n1069 gnd 0.202911f
C3088 vdd.n1070 gnd 0.004973f
C3089 vdd.n1071 gnd 0.004615f
C3090 vdd.n1072 gnd 0.002553f
C3091 vdd.n1073 gnd 0.005861f
C3092 vdd.n1074 gnd 0.00248f
C3093 vdd.n1075 gnd 0.002626f
C3094 vdd.n1076 gnd 0.004615f
C3095 vdd.n1077 gnd 0.00248f
C3096 vdd.n1078 gnd 0.005861f
C3097 vdd.n1079 gnd 0.002626f
C3098 vdd.n1080 gnd 0.004615f
C3099 vdd.n1081 gnd 0.00248f
C3100 vdd.n1082 gnd 0.004396f
C3101 vdd.n1083 gnd 0.004409f
C3102 vdd.t179 gnd 0.012592f
C3103 vdd.n1084 gnd 0.028017f
C3104 vdd.n1085 gnd 0.145808f
C3105 vdd.n1086 gnd 0.00248f
C3106 vdd.n1087 gnd 0.002626f
C3107 vdd.n1088 gnd 0.005861f
C3108 vdd.n1089 gnd 0.005861f
C3109 vdd.n1090 gnd 0.002626f
C3110 vdd.n1091 gnd 0.00248f
C3111 vdd.n1092 gnd 0.004615f
C3112 vdd.n1093 gnd 0.004615f
C3113 vdd.n1094 gnd 0.00248f
C3114 vdd.n1095 gnd 0.002626f
C3115 vdd.n1096 gnd 0.005861f
C3116 vdd.n1097 gnd 0.005861f
C3117 vdd.n1098 gnd 0.002626f
C3118 vdd.n1099 gnd 0.00248f
C3119 vdd.n1100 gnd 0.004615f
C3120 vdd.n1101 gnd 0.004615f
C3121 vdd.n1102 gnd 0.00248f
C3122 vdd.n1103 gnd 0.002626f
C3123 vdd.n1104 gnd 0.005861f
C3124 vdd.n1105 gnd 0.005861f
C3125 vdd.n1106 gnd 0.013857f
C3126 vdd.n1107 gnd 0.002553f
C3127 vdd.n1108 gnd 0.00248f
C3128 vdd.n1109 gnd 0.011927f
C3129 vdd.n1110 gnd 0.008327f
C3130 vdd.t134 gnd 0.029173f
C3131 vdd.t178 gnd 0.029173f
C3132 vdd.n1111 gnd 0.200496f
C3133 vdd.n1112 gnd 0.15766f
C3134 vdd.t177 gnd 0.029173f
C3135 vdd.t166 gnd 0.029173f
C3136 vdd.n1113 gnd 0.200496f
C3137 vdd.n1114 gnd 0.12723f
C3138 vdd.t153 gnd 0.029173f
C3139 vdd.t132 gnd 0.029173f
C3140 vdd.n1115 gnd 0.200496f
C3141 vdd.n1116 gnd 0.12723f
C3142 vdd.n1117 gnd 0.004973f
C3143 vdd.n1118 gnd 0.004615f
C3144 vdd.n1119 gnd 0.002553f
C3145 vdd.n1120 gnd 0.005861f
C3146 vdd.n1121 gnd 0.00248f
C3147 vdd.n1122 gnd 0.002626f
C3148 vdd.n1123 gnd 0.004615f
C3149 vdd.n1124 gnd 0.00248f
C3150 vdd.n1125 gnd 0.005861f
C3151 vdd.n1126 gnd 0.002626f
C3152 vdd.n1127 gnd 0.004615f
C3153 vdd.n1128 gnd 0.00248f
C3154 vdd.n1129 gnd 0.004396f
C3155 vdd.n1130 gnd 0.004409f
C3156 vdd.t165 gnd 0.012592f
C3157 vdd.n1131 gnd 0.028017f
C3158 vdd.n1132 gnd 0.145808f
C3159 vdd.n1133 gnd 0.00248f
C3160 vdd.n1134 gnd 0.002626f
C3161 vdd.n1135 gnd 0.005861f
C3162 vdd.n1136 gnd 0.005861f
C3163 vdd.n1137 gnd 0.002626f
C3164 vdd.n1138 gnd 0.00248f
C3165 vdd.n1139 gnd 0.004615f
C3166 vdd.n1140 gnd 0.004615f
C3167 vdd.n1141 gnd 0.00248f
C3168 vdd.n1142 gnd 0.002626f
C3169 vdd.n1143 gnd 0.005861f
C3170 vdd.n1144 gnd 0.005861f
C3171 vdd.n1145 gnd 0.002626f
C3172 vdd.n1146 gnd 0.00248f
C3173 vdd.n1147 gnd 0.004615f
C3174 vdd.n1148 gnd 0.004615f
C3175 vdd.n1149 gnd 0.00248f
C3176 vdd.n1150 gnd 0.002626f
C3177 vdd.n1151 gnd 0.005861f
C3178 vdd.n1152 gnd 0.005861f
C3179 vdd.n1153 gnd 0.013857f
C3180 vdd.n1154 gnd 0.002553f
C3181 vdd.n1155 gnd 0.00248f
C3182 vdd.n1156 gnd 0.011927f
C3183 vdd.n1157 gnd 0.008066f
C3184 vdd.n1158 gnd 0.056313f
C3185 vdd.n1159 gnd 0.219627f
C3186 vdd.n1160 gnd 1.8458f
C3187 vdd.n1161 gnd 0.534468f
C3188 vdd.n1162 gnd 0.007293f
C3189 vdd.n1163 gnd 0.009061f
C3190 vdd.n1164 gnd 0.569501f
C3191 vdd.n1165 gnd 0.009061f
C3192 vdd.n1166 gnd 0.007293f
C3193 vdd.n1167 gnd 0.009061f
C3194 vdd.n1168 gnd 0.007293f
C3195 vdd.n1169 gnd 0.009061f
C3196 vdd.t124 gnd 0.463009f
C3197 vdd.t135 gnd 0.463009f
C3198 vdd.n1170 gnd 0.009061f
C3199 vdd.n1171 gnd 0.007293f
C3200 vdd.n1172 gnd 0.009061f
C3201 vdd.n1173 gnd 0.007293f
C3202 vdd.n1174 gnd 0.009061f
C3203 vdd.t141 gnd 0.463009f
C3204 vdd.n1175 gnd 0.009061f
C3205 vdd.n1176 gnd 0.007293f
C3206 vdd.n1177 gnd 0.009061f
C3207 vdd.n1178 gnd 0.007293f
C3208 vdd.n1179 gnd 0.009061f
C3209 vdd.t157 gnd 0.463009f
C3210 vdd.n1180 gnd 0.671363f
C3211 vdd.n1181 gnd 0.009061f
C3212 vdd.n1182 gnd 0.007293f
C3213 vdd.n1183 gnd 0.009061f
C3214 vdd.n1184 gnd 0.007293f
C3215 vdd.n1185 gnd 0.009061f
C3216 vdd.n1186 gnd 0.926018f
C3217 vdd.n1187 gnd 0.009061f
C3218 vdd.n1188 gnd 0.007293f
C3219 vdd.n1189 gnd 0.022083f
C3220 vdd.n1190 gnd 0.006053f
C3221 vdd.n1191 gnd 0.022083f
C3222 vdd.t44 gnd 0.463009f
C3223 vdd.n1192 gnd 0.022083f
C3224 vdd.n1193 gnd 0.006053f
C3225 vdd.n1194 gnd 0.009061f
C3226 vdd.n1195 gnd 0.007293f
C3227 vdd.n1196 gnd 0.009061f
C3228 vdd.n1227 gnd 0.022589f
C3229 vdd.n1228 gnd 1.36588f
C3230 vdd.n1229 gnd 0.009061f
C3231 vdd.n1230 gnd 0.007293f
C3232 vdd.n1231 gnd 0.009061f
C3233 vdd.n1232 gnd 0.009061f
C3234 vdd.n1233 gnd 0.009061f
C3235 vdd.n1234 gnd 0.009061f
C3236 vdd.n1235 gnd 0.009061f
C3237 vdd.n1236 gnd 0.007293f
C3238 vdd.n1237 gnd 0.009061f
C3239 vdd.n1238 gnd 0.009061f
C3240 vdd.n1239 gnd 0.009061f
C3241 vdd.n1240 gnd 0.009061f
C3242 vdd.n1241 gnd 0.009061f
C3243 vdd.n1242 gnd 0.007293f
C3244 vdd.n1243 gnd 0.009061f
C3245 vdd.n1244 gnd 0.009061f
C3246 vdd.n1245 gnd 0.009061f
C3247 vdd.n1246 gnd 0.009061f
C3248 vdd.n1247 gnd 0.009061f
C3249 vdd.n1248 gnd 0.007293f
C3250 vdd.n1249 gnd 0.009061f
C3251 vdd.n1250 gnd 0.009061f
C3252 vdd.n1251 gnd 0.009061f
C3253 vdd.n1252 gnd 0.009061f
C3254 vdd.n1253 gnd 0.009061f
C3255 vdd.t94 gnd 0.111477f
C3256 vdd.t95 gnd 0.119139f
C3257 vdd.t93 gnd 0.145588f
C3258 vdd.n1254 gnd 0.186623f
C3259 vdd.n1255 gnd 0.157527f
C3260 vdd.n1256 gnd 0.015608f
C3261 vdd.n1257 gnd 0.009061f
C3262 vdd.n1258 gnd 0.009061f
C3263 vdd.n1259 gnd 0.009061f
C3264 vdd.n1260 gnd 0.009061f
C3265 vdd.n1261 gnd 0.009061f
C3266 vdd.n1262 gnd 0.007293f
C3267 vdd.n1263 gnd 0.009061f
C3268 vdd.n1264 gnd 0.009061f
C3269 vdd.n1265 gnd 0.009061f
C3270 vdd.n1266 gnd 0.009061f
C3271 vdd.n1267 gnd 0.009061f
C3272 vdd.n1268 gnd 0.007293f
C3273 vdd.n1269 gnd 0.009061f
C3274 vdd.n1270 gnd 0.009061f
C3275 vdd.n1271 gnd 0.009061f
C3276 vdd.n1272 gnd 0.009061f
C3277 vdd.n1273 gnd 0.009061f
C3278 vdd.n1274 gnd 0.007293f
C3279 vdd.n1275 gnd 0.009061f
C3280 vdd.n1276 gnd 0.009061f
C3281 vdd.n1277 gnd 0.009061f
C3282 vdd.n1278 gnd 0.009061f
C3283 vdd.n1279 gnd 0.009061f
C3284 vdd.n1280 gnd 0.007293f
C3285 vdd.n1281 gnd 0.009061f
C3286 vdd.n1282 gnd 0.009061f
C3287 vdd.n1283 gnd 0.009061f
C3288 vdd.n1284 gnd 0.009061f
C3289 vdd.n1285 gnd 0.009061f
C3290 vdd.n1286 gnd 0.007293f
C3291 vdd.n1287 gnd 0.009061f
C3292 vdd.n1288 gnd 0.009061f
C3293 vdd.n1289 gnd 0.009061f
C3294 vdd.n1290 gnd 0.009061f
C3295 vdd.n1291 gnd 0.007293f
C3296 vdd.n1292 gnd 0.009061f
C3297 vdd.n1293 gnd 0.009061f
C3298 vdd.n1294 gnd 0.009061f
C3299 vdd.n1295 gnd 0.009061f
C3300 vdd.n1296 gnd 0.009061f
C3301 vdd.n1297 gnd 0.007293f
C3302 vdd.n1298 gnd 0.009061f
C3303 vdd.n1299 gnd 0.009061f
C3304 vdd.n1300 gnd 0.009061f
C3305 vdd.n1301 gnd 0.009061f
C3306 vdd.n1302 gnd 0.009061f
C3307 vdd.n1303 gnd 0.007293f
C3308 vdd.n1304 gnd 0.009061f
C3309 vdd.n1305 gnd 0.009061f
C3310 vdd.n1306 gnd 0.009061f
C3311 vdd.n1307 gnd 0.009061f
C3312 vdd.n1308 gnd 0.009061f
C3313 vdd.n1309 gnd 0.007293f
C3314 vdd.n1310 gnd 0.009061f
C3315 vdd.n1311 gnd 0.009061f
C3316 vdd.n1312 gnd 0.009061f
C3317 vdd.n1313 gnd 0.009061f
C3318 vdd.n1314 gnd 0.009061f
C3319 vdd.n1315 gnd 0.007293f
C3320 vdd.n1316 gnd 0.009061f
C3321 vdd.n1317 gnd 0.009061f
C3322 vdd.n1318 gnd 0.009061f
C3323 vdd.n1319 gnd 0.009061f
C3324 vdd.t45 gnd 0.111477f
C3325 vdd.t46 gnd 0.119139f
C3326 vdd.t43 gnd 0.145588f
C3327 vdd.n1320 gnd 0.186623f
C3328 vdd.n1321 gnd 0.157527f
C3329 vdd.n1322 gnd 0.011961f
C3330 vdd.n1323 gnd 0.003464f
C3331 vdd.n1324 gnd 0.022589f
C3332 vdd.n1325 gnd 0.009061f
C3333 vdd.n1326 gnd 0.003829f
C3334 vdd.n1327 gnd 0.007293f
C3335 vdd.n1328 gnd 0.007293f
C3336 vdd.n1329 gnd 0.009061f
C3337 vdd.n1330 gnd 0.009061f
C3338 vdd.n1331 gnd 0.009061f
C3339 vdd.n1332 gnd 0.007293f
C3340 vdd.n1333 gnd 0.007293f
C3341 vdd.n1334 gnd 0.007293f
C3342 vdd.n1335 gnd 0.009061f
C3343 vdd.n1336 gnd 0.009061f
C3344 vdd.n1337 gnd 0.009061f
C3345 vdd.n1338 gnd 0.007293f
C3346 vdd.n1339 gnd 0.007293f
C3347 vdd.n1340 gnd 0.007293f
C3348 vdd.n1341 gnd 0.009061f
C3349 vdd.n1342 gnd 0.009061f
C3350 vdd.n1343 gnd 0.009061f
C3351 vdd.n1344 gnd 0.007293f
C3352 vdd.n1345 gnd 0.007293f
C3353 vdd.n1346 gnd 0.007293f
C3354 vdd.n1347 gnd 0.009061f
C3355 vdd.n1348 gnd 0.009061f
C3356 vdd.n1349 gnd 0.009061f
C3357 vdd.n1350 gnd 0.007293f
C3358 vdd.n1351 gnd 0.007293f
C3359 vdd.n1352 gnd 0.007293f
C3360 vdd.n1353 gnd 0.009061f
C3361 vdd.n1354 gnd 0.009061f
C3362 vdd.n1355 gnd 0.009061f
C3363 vdd.n1356 gnd 0.00722f
C3364 vdd.n1357 gnd 0.009061f
C3365 vdd.t91 gnd 0.111477f
C3366 vdd.t92 gnd 0.119139f
C3367 vdd.t90 gnd 0.145588f
C3368 vdd.n1358 gnd 0.186623f
C3369 vdd.n1359 gnd 0.157527f
C3370 vdd.n1360 gnd 0.015608f
C3371 vdd.n1361 gnd 0.004959f
C3372 vdd.n1362 gnd 0.009061f
C3373 vdd.n1363 gnd 0.009061f
C3374 vdd.n1364 gnd 0.009061f
C3375 vdd.n1365 gnd 0.007293f
C3376 vdd.n1366 gnd 0.007293f
C3377 vdd.n1367 gnd 0.007293f
C3378 vdd.n1368 gnd 0.009061f
C3379 vdd.n1369 gnd 0.009061f
C3380 vdd.n1370 gnd 0.009061f
C3381 vdd.n1371 gnd 0.007293f
C3382 vdd.n1372 gnd 0.007293f
C3383 vdd.n1373 gnd 0.007293f
C3384 vdd.n1374 gnd 0.009061f
C3385 vdd.n1375 gnd 0.009061f
C3386 vdd.n1376 gnd 0.009061f
C3387 vdd.n1377 gnd 0.007293f
C3388 vdd.n1378 gnd 0.007293f
C3389 vdd.n1379 gnd 0.007293f
C3390 vdd.n1380 gnd 0.009061f
C3391 vdd.n1381 gnd 0.009061f
C3392 vdd.n1382 gnd 0.009061f
C3393 vdd.n1383 gnd 0.007293f
C3394 vdd.n1384 gnd 0.007293f
C3395 vdd.n1385 gnd 0.007293f
C3396 vdd.n1386 gnd 0.009061f
C3397 vdd.n1387 gnd 0.009061f
C3398 vdd.n1388 gnd 0.009061f
C3399 vdd.n1389 gnd 0.007293f
C3400 vdd.n1390 gnd 0.007293f
C3401 vdd.n1391 gnd 0.00609f
C3402 vdd.n1392 gnd 0.009061f
C3403 vdd.n1393 gnd 0.009061f
C3404 vdd.n1394 gnd 0.009061f
C3405 vdd.n1395 gnd 0.00609f
C3406 vdd.n1396 gnd 0.007293f
C3407 vdd.n1397 gnd 0.007293f
C3408 vdd.n1398 gnd 0.009061f
C3409 vdd.n1399 gnd 0.009061f
C3410 vdd.n1400 gnd 0.009061f
C3411 vdd.n1401 gnd 0.007293f
C3412 vdd.n1402 gnd 0.007293f
C3413 vdd.n1403 gnd 0.007293f
C3414 vdd.n1404 gnd 0.009061f
C3415 vdd.n1405 gnd 0.009061f
C3416 vdd.n1406 gnd 0.009061f
C3417 vdd.n1407 gnd 0.007293f
C3418 vdd.n1408 gnd 0.007293f
C3419 vdd.n1409 gnd 0.007293f
C3420 vdd.n1410 gnd 0.009061f
C3421 vdd.n1411 gnd 0.009061f
C3422 vdd.n1412 gnd 0.009061f
C3423 vdd.n1413 gnd 0.007293f
C3424 vdd.n1414 gnd 0.007293f
C3425 vdd.n1415 gnd 0.007293f
C3426 vdd.n1416 gnd 0.009061f
C3427 vdd.n1417 gnd 0.009061f
C3428 vdd.n1418 gnd 0.009061f
C3429 vdd.n1419 gnd 0.007293f
C3430 vdd.n1420 gnd 0.009061f
C3431 vdd.n1421 gnd 2.21318f
C3432 vdd.n1423 gnd 0.022589f
C3433 vdd.n1424 gnd 0.006053f
C3434 vdd.n1425 gnd 0.022589f
C3435 vdd.n1426 gnd 0.022083f
C3436 vdd.n1427 gnd 0.009061f
C3437 vdd.n1428 gnd 0.007293f
C3438 vdd.n1429 gnd 0.009061f
C3439 vdd.n1430 gnd 0.48616f
C3440 vdd.n1431 gnd 0.009061f
C3441 vdd.n1432 gnd 0.007293f
C3442 vdd.n1433 gnd 0.009061f
C3443 vdd.n1434 gnd 0.009061f
C3444 vdd.n1435 gnd 0.009061f
C3445 vdd.n1436 gnd 0.007293f
C3446 vdd.n1437 gnd 0.009061f
C3447 vdd.n1438 gnd 0.828786f
C3448 vdd.n1439 gnd 0.926018f
C3449 vdd.n1440 gnd 0.009061f
C3450 vdd.n1441 gnd 0.007293f
C3451 vdd.n1442 gnd 0.009061f
C3452 vdd.n1443 gnd 0.009061f
C3453 vdd.n1444 gnd 0.009061f
C3454 vdd.n1445 gnd 0.007293f
C3455 vdd.n1446 gnd 0.009061f
C3456 vdd.n1447 gnd 0.560241f
C3457 vdd.n1448 gnd 0.009061f
C3458 vdd.n1449 gnd 0.007293f
C3459 vdd.n1450 gnd 0.009061f
C3460 vdd.n1451 gnd 0.009061f
C3461 vdd.n1452 gnd 0.009061f
C3462 vdd.n1453 gnd 0.007293f
C3463 vdd.n1454 gnd 0.009061f
C3464 vdd.n1455 gnd 0.51394f
C3465 vdd.n1456 gnd 0.717664f
C3466 vdd.n1457 gnd 0.009061f
C3467 vdd.n1458 gnd 0.007293f
C3468 vdd.n1459 gnd 0.009061f
C3469 vdd.n1460 gnd 0.009061f
C3470 vdd.n1461 gnd 0.006964f
C3471 vdd.n1462 gnd 0.009061f
C3472 vdd.n1463 gnd 0.007293f
C3473 vdd.n1464 gnd 0.009061f
C3474 vdd.n1465 gnd 0.768595f
C3475 vdd.n1466 gnd 0.009061f
C3476 vdd.n1467 gnd 0.007293f
C3477 vdd.n1468 gnd 0.009061f
C3478 vdd.n1469 gnd 0.009061f
C3479 vdd.n1470 gnd 0.009061f
C3480 vdd.n1471 gnd 0.007293f
C3481 vdd.n1472 gnd 0.009061f
C3482 vdd.t159 gnd 0.463009f
C3483 vdd.n1473 gnd 0.662103f
C3484 vdd.n1474 gnd 0.009061f
C3485 vdd.n1475 gnd 0.007293f
C3486 vdd.n1476 gnd 0.006964f
C3487 vdd.n1477 gnd 0.009061f
C3488 vdd.n1478 gnd 0.009061f
C3489 vdd.n1479 gnd 0.007293f
C3490 vdd.n1480 gnd 0.009061f
C3491 vdd.n1481 gnd 0.50468f
C3492 vdd.n1482 gnd 0.009061f
C3493 vdd.n1483 gnd 0.007293f
C3494 vdd.n1484 gnd 0.009061f
C3495 vdd.n1485 gnd 0.009061f
C3496 vdd.n1486 gnd 0.009061f
C3497 vdd.n1487 gnd 0.007293f
C3498 vdd.n1488 gnd 0.009061f
C3499 vdd.n1489 gnd 0.652843f
C3500 vdd.n1490 gnd 0.578761f
C3501 vdd.n1491 gnd 0.009061f
C3502 vdd.n1492 gnd 0.007293f
C3503 vdd.n1493 gnd 0.009061f
C3504 vdd.n1494 gnd 0.009061f
C3505 vdd.n1495 gnd 0.009061f
C3506 vdd.n1496 gnd 0.007293f
C3507 vdd.n1497 gnd 0.009061f
C3508 vdd.n1498 gnd 0.736185f
C3509 vdd.n1499 gnd 0.009061f
C3510 vdd.n1500 gnd 0.007293f
C3511 vdd.n1501 gnd 0.009061f
C3512 vdd.n1502 gnd 0.009061f
C3513 vdd.n1503 gnd 0.022083f
C3514 vdd.n1504 gnd 0.009061f
C3515 vdd.n1505 gnd 0.009061f
C3516 vdd.n1506 gnd 0.007293f
C3517 vdd.n1507 gnd 0.009061f
C3518 vdd.n1508 gnd 0.578761f
C3519 vdd.n1509 gnd 0.926018f
C3520 vdd.n1510 gnd 0.009061f
C3521 vdd.n1511 gnd 0.007293f
C3522 vdd.n1512 gnd 0.009061f
C3523 vdd.n1513 gnd 0.009061f
C3524 vdd.n1514 gnd 0.007793f
C3525 vdd.n1515 gnd 0.007293f
C3526 vdd.n1517 gnd 0.009061f
C3527 vdd.n1519 gnd 0.007293f
C3528 vdd.n1520 gnd 0.009061f
C3529 vdd.n1521 gnd 0.007293f
C3530 vdd.n1523 gnd 0.009061f
C3531 vdd.n1524 gnd 0.007293f
C3532 vdd.n1525 gnd 0.009061f
C3533 vdd.n1526 gnd 0.009061f
C3534 vdd.n1527 gnd 0.009061f
C3535 vdd.n1528 gnd 0.009061f
C3536 vdd.n1529 gnd 0.009061f
C3537 vdd.n1530 gnd 0.007293f
C3538 vdd.n1532 gnd 0.009061f
C3539 vdd.n1533 gnd 0.009061f
C3540 vdd.n1534 gnd 0.009061f
C3541 vdd.n1535 gnd 0.009061f
C3542 vdd.n1536 gnd 0.009061f
C3543 vdd.n1537 gnd 0.007293f
C3544 vdd.n1539 gnd 0.009061f
C3545 vdd.n1540 gnd 0.009061f
C3546 vdd.n1541 gnd 0.009061f
C3547 vdd.n1542 gnd 0.009061f
C3548 vdd.n1543 gnd 0.00609f
C3549 vdd.t60 gnd 0.111477f
C3550 vdd.t59 gnd 0.119139f
C3551 vdd.t58 gnd 0.145588f
C3552 vdd.n1544 gnd 0.186623f
C3553 vdd.n1545 gnd 0.156797f
C3554 vdd.n1547 gnd 0.009061f
C3555 vdd.n1548 gnd 0.009061f
C3556 vdd.n1549 gnd 0.007293f
C3557 vdd.n1550 gnd 0.009061f
C3558 vdd.n1552 gnd 0.009061f
C3559 vdd.n1553 gnd 0.009061f
C3560 vdd.n1554 gnd 0.009061f
C3561 vdd.n1555 gnd 0.009061f
C3562 vdd.n1556 gnd 0.007293f
C3563 vdd.n1558 gnd 0.009061f
C3564 vdd.n1559 gnd 0.009061f
C3565 vdd.n1560 gnd 0.009061f
C3566 vdd.n1561 gnd 0.009061f
C3567 vdd.n1562 gnd 0.009061f
C3568 vdd.n1563 gnd 0.007293f
C3569 vdd.n1565 gnd 0.009061f
C3570 vdd.n1566 gnd 0.009061f
C3571 vdd.n1567 gnd 0.009061f
C3572 vdd.n1568 gnd 0.009061f
C3573 vdd.n1569 gnd 0.009061f
C3574 vdd.n1570 gnd 0.007293f
C3575 vdd.n1572 gnd 0.009061f
C3576 vdd.n1573 gnd 0.009061f
C3577 vdd.n1574 gnd 0.009061f
C3578 vdd.n1575 gnd 0.009061f
C3579 vdd.n1576 gnd 0.009061f
C3580 vdd.n1577 gnd 0.007293f
C3581 vdd.n1579 gnd 0.009061f
C3582 vdd.n1580 gnd 0.009061f
C3583 vdd.n1581 gnd 0.009061f
C3584 vdd.n1582 gnd 0.009061f
C3585 vdd.n1583 gnd 0.00722f
C3586 vdd.t53 gnd 0.111477f
C3587 vdd.t52 gnd 0.119139f
C3588 vdd.t51 gnd 0.145588f
C3589 vdd.n1584 gnd 0.186623f
C3590 vdd.n1585 gnd 0.156797f
C3591 vdd.n1587 gnd 0.009061f
C3592 vdd.n1588 gnd 0.009061f
C3593 vdd.n1589 gnd 0.007293f
C3594 vdd.n1590 gnd 0.009061f
C3595 vdd.n1592 gnd 0.009061f
C3596 vdd.n1593 gnd 0.009061f
C3597 vdd.n1594 gnd 0.009061f
C3598 vdd.n1595 gnd 0.009061f
C3599 vdd.n1596 gnd 0.007293f
C3600 vdd.n1598 gnd 0.009061f
C3601 vdd.n1599 gnd 0.009061f
C3602 vdd.n1600 gnd 0.009061f
C3603 vdd.n1601 gnd 0.009061f
C3604 vdd.n1602 gnd 0.009061f
C3605 vdd.n1603 gnd 0.007293f
C3606 vdd.n1605 gnd 0.009061f
C3607 vdd.n1606 gnd 0.009061f
C3608 vdd.n1607 gnd 0.009061f
C3609 vdd.n1608 gnd 0.009061f
C3610 vdd.n1609 gnd 0.009061f
C3611 vdd.n1610 gnd 0.009061f
C3612 vdd.n1611 gnd 0.007293f
C3613 vdd.n1613 gnd 0.009061f
C3614 vdd.n1615 gnd 0.009061f
C3615 vdd.n1616 gnd 0.007293f
C3616 vdd.n1617 gnd 0.007293f
C3617 vdd.n1618 gnd 0.009061f
C3618 vdd.n1620 gnd 0.009061f
C3619 vdd.n1621 gnd 0.007293f
C3620 vdd.n1622 gnd 0.007293f
C3621 vdd.n1623 gnd 0.009061f
C3622 vdd.n1625 gnd 0.009061f
C3623 vdd.n1626 gnd 0.009061f
C3624 vdd.n1627 gnd 0.007293f
C3625 vdd.n1628 gnd 0.007293f
C3626 vdd.n1629 gnd 0.007293f
C3627 vdd.n1630 gnd 0.009061f
C3628 vdd.n1632 gnd 0.009061f
C3629 vdd.n1633 gnd 0.009061f
C3630 vdd.n1634 gnd 0.007293f
C3631 vdd.n1635 gnd 0.007293f
C3632 vdd.n1636 gnd 0.007293f
C3633 vdd.n1637 gnd 0.009061f
C3634 vdd.n1639 gnd 0.009061f
C3635 vdd.n1640 gnd 0.009061f
C3636 vdd.n1641 gnd 0.007293f
C3637 vdd.n1642 gnd 0.007293f
C3638 vdd.n1643 gnd 0.007293f
C3639 vdd.n1644 gnd 0.009061f
C3640 vdd.n1646 gnd 0.009061f
C3641 vdd.n1647 gnd 0.009061f
C3642 vdd.n1648 gnd 0.007293f
C3643 vdd.n1649 gnd 0.009061f
C3644 vdd.n1650 gnd 0.009061f
C3645 vdd.n1651 gnd 0.009061f
C3646 vdd.n1652 gnd 0.014878f
C3647 vdd.n1653 gnd 0.004959f
C3648 vdd.n1654 gnd 0.007293f
C3649 vdd.n1655 gnd 0.009061f
C3650 vdd.n1657 gnd 0.009061f
C3651 vdd.n1658 gnd 0.009061f
C3652 vdd.n1659 gnd 0.007293f
C3653 vdd.n1660 gnd 0.007293f
C3654 vdd.n1661 gnd 0.007293f
C3655 vdd.n1662 gnd 0.009061f
C3656 vdd.n1664 gnd 0.009061f
C3657 vdd.n1665 gnd 0.009061f
C3658 vdd.n1666 gnd 0.007293f
C3659 vdd.n1667 gnd 0.007293f
C3660 vdd.n1668 gnd 0.007293f
C3661 vdd.n1669 gnd 0.009061f
C3662 vdd.n1671 gnd 0.009061f
C3663 vdd.n1672 gnd 0.009061f
C3664 vdd.n1673 gnd 0.007293f
C3665 vdd.n1674 gnd 0.007293f
C3666 vdd.n1675 gnd 0.007293f
C3667 vdd.n1676 gnd 0.009061f
C3668 vdd.n1678 gnd 0.009061f
C3669 vdd.n1679 gnd 0.009061f
C3670 vdd.n1680 gnd 0.007293f
C3671 vdd.n1681 gnd 0.007293f
C3672 vdd.n1682 gnd 0.007293f
C3673 vdd.n1683 gnd 0.009061f
C3674 vdd.n1685 gnd 0.009061f
C3675 vdd.n1686 gnd 0.009061f
C3676 vdd.n1687 gnd 0.007293f
C3677 vdd.n1688 gnd 0.009061f
C3678 vdd.n1689 gnd 0.009061f
C3679 vdd.n1690 gnd 0.009061f
C3680 vdd.n1691 gnd 0.014878f
C3681 vdd.n1692 gnd 0.00609f
C3682 vdd.n1693 gnd 0.007293f
C3683 vdd.n1694 gnd 0.009061f
C3684 vdd.n1696 gnd 0.009061f
C3685 vdd.n1697 gnd 0.009061f
C3686 vdd.n1698 gnd 0.007293f
C3687 vdd.n1699 gnd 0.007293f
C3688 vdd.n1700 gnd 0.007293f
C3689 vdd.n1701 gnd 0.009061f
C3690 vdd.n1703 gnd 0.009061f
C3691 vdd.n1704 gnd 0.009061f
C3692 vdd.n1705 gnd 0.007293f
C3693 vdd.n1706 gnd 0.007293f
C3694 vdd.n1707 gnd 0.007293f
C3695 vdd.n1708 gnd 0.009061f
C3696 vdd.n1710 gnd 0.009061f
C3697 vdd.n1711 gnd 0.009061f
C3698 vdd.n1713 gnd 0.009061f
C3699 vdd.n1714 gnd 0.007293f
C3700 vdd.n1715 gnd 0.005799f
C3701 vdd.n1716 gnd 0.006162f
C3702 vdd.n1717 gnd 0.006162f
C3703 vdd.n1718 gnd 0.006162f
C3704 vdd.n1719 gnd 0.006162f
C3705 vdd.n1720 gnd 0.006162f
C3706 vdd.n1721 gnd 0.006162f
C3707 vdd.n1722 gnd 0.006162f
C3708 vdd.n1723 gnd 0.006162f
C3709 vdd.n1725 gnd 0.006162f
C3710 vdd.n1726 gnd 0.006162f
C3711 vdd.n1727 gnd 0.006162f
C3712 vdd.n1728 gnd 0.006162f
C3713 vdd.n1729 gnd 0.006162f
C3714 vdd.n1731 gnd 0.006162f
C3715 vdd.n1733 gnd 0.006162f
C3716 vdd.n1734 gnd 0.006162f
C3717 vdd.n1735 gnd 0.006162f
C3718 vdd.n1736 gnd 0.006162f
C3719 vdd.n1737 gnd 0.006162f
C3720 vdd.n1739 gnd 0.006162f
C3721 vdd.n1741 gnd 0.006162f
C3722 vdd.n1742 gnd 0.006162f
C3723 vdd.n1743 gnd 0.006162f
C3724 vdd.n1744 gnd 0.006162f
C3725 vdd.n1745 gnd 0.006162f
C3726 vdd.n1747 gnd 0.006162f
C3727 vdd.n1749 gnd 0.006162f
C3728 vdd.n1750 gnd 0.006162f
C3729 vdd.n1751 gnd 0.006162f
C3730 vdd.n1752 gnd 0.006162f
C3731 vdd.n1753 gnd 0.006162f
C3732 vdd.n1755 gnd 0.006162f
C3733 vdd.n1756 gnd 0.006162f
C3734 vdd.n1757 gnd 0.006162f
C3735 vdd.n1758 gnd 0.006162f
C3736 vdd.n1759 gnd 0.006162f
C3737 vdd.n1760 gnd 0.006162f
C3738 vdd.n1761 gnd 0.006162f
C3739 vdd.n1762 gnd 0.006162f
C3740 vdd.n1763 gnd 0.004485f
C3741 vdd.n1764 gnd 0.006162f
C3742 vdd.t106 gnd 0.248992f
C3743 vdd.t107 gnd 0.254874f
C3744 vdd.t105 gnd 0.162551f
C3745 vdd.n1765 gnd 0.08785f
C3746 vdd.n1766 gnd 0.049831f
C3747 vdd.n1767 gnd 0.008806f
C3748 vdd.n1768 gnd 0.006162f
C3749 vdd.n1769 gnd 0.006162f
C3750 vdd.n1770 gnd 0.375037f
C3751 vdd.n1771 gnd 0.006162f
C3752 vdd.n1772 gnd 0.006162f
C3753 vdd.n1773 gnd 0.006162f
C3754 vdd.n1774 gnd 0.006162f
C3755 vdd.n1775 gnd 0.006162f
C3756 vdd.n1776 gnd 0.006162f
C3757 vdd.n1777 gnd 0.006162f
C3758 vdd.n1778 gnd 0.006162f
C3759 vdd.n1779 gnd 0.006162f
C3760 vdd.n1780 gnd 0.006162f
C3761 vdd.n1781 gnd 0.006162f
C3762 vdd.n1782 gnd 0.006162f
C3763 vdd.n1783 gnd 0.006162f
C3764 vdd.n1784 gnd 0.006162f
C3765 vdd.n1785 gnd 0.006162f
C3766 vdd.n1786 gnd 0.006162f
C3767 vdd.n1787 gnd 0.006162f
C3768 vdd.n1788 gnd 0.006162f
C3769 vdd.n1789 gnd 0.006162f
C3770 vdd.n1790 gnd 0.006162f
C3771 vdd.t81 gnd 0.248992f
C3772 vdd.t82 gnd 0.254874f
C3773 vdd.t79 gnd 0.162551f
C3774 vdd.n1791 gnd 0.08785f
C3775 vdd.n1792 gnd 0.049831f
C3776 vdd.n1793 gnd 0.006162f
C3777 vdd.n1794 gnd 0.006162f
C3778 vdd.n1795 gnd 0.006162f
C3779 vdd.n1796 gnd 0.006162f
C3780 vdd.n1797 gnd 0.006162f
C3781 vdd.n1798 gnd 0.006162f
C3782 vdd.n1800 gnd 0.006162f
C3783 vdd.n1801 gnd 0.006162f
C3784 vdd.n1802 gnd 0.006162f
C3785 vdd.n1803 gnd 0.006162f
C3786 vdd.n1805 gnd 0.006162f
C3787 vdd.n1807 gnd 0.006162f
C3788 vdd.n1808 gnd 0.006162f
C3789 vdd.n1809 gnd 0.006162f
C3790 vdd.n1810 gnd 0.006162f
C3791 vdd.n1811 gnd 0.006162f
C3792 vdd.n1813 gnd 0.006162f
C3793 vdd.n1815 gnd 0.006162f
C3794 vdd.n1816 gnd 0.006162f
C3795 vdd.n1817 gnd 0.006162f
C3796 vdd.n1818 gnd 0.006162f
C3797 vdd.n1819 gnd 0.006162f
C3798 vdd.n1821 gnd 0.006162f
C3799 vdd.n1823 gnd 0.006162f
C3800 vdd.n1824 gnd 0.006162f
C3801 vdd.n1825 gnd 0.004485f
C3802 vdd.n1826 gnd 0.008806f
C3803 vdd.n1827 gnd 0.004757f
C3804 vdd.n1828 gnd 0.006162f
C3805 vdd.n1830 gnd 0.006162f
C3806 vdd.n1831 gnd 0.014621f
C3807 vdd.n1832 gnd 0.014621f
C3808 vdd.n1833 gnd 0.013651f
C3809 vdd.n1834 gnd 0.006162f
C3810 vdd.n1835 gnd 0.006162f
C3811 vdd.n1836 gnd 0.006162f
C3812 vdd.n1837 gnd 0.006162f
C3813 vdd.n1838 gnd 0.006162f
C3814 vdd.n1839 gnd 0.006162f
C3815 vdd.n1840 gnd 0.006162f
C3816 vdd.n1841 gnd 0.006162f
C3817 vdd.n1842 gnd 0.006162f
C3818 vdd.n1843 gnd 0.006162f
C3819 vdd.n1844 gnd 0.006162f
C3820 vdd.n1845 gnd 0.006162f
C3821 vdd.n1846 gnd 0.006162f
C3822 vdd.n1847 gnd 0.006162f
C3823 vdd.n1848 gnd 0.006162f
C3824 vdd.n1849 gnd 0.006162f
C3825 vdd.n1850 gnd 0.006162f
C3826 vdd.n1851 gnd 0.006162f
C3827 vdd.n1852 gnd 0.006162f
C3828 vdd.n1853 gnd 0.006162f
C3829 vdd.n1854 gnd 0.006162f
C3830 vdd.n1855 gnd 0.006162f
C3831 vdd.n1856 gnd 0.006162f
C3832 vdd.n1857 gnd 0.006162f
C3833 vdd.n1858 gnd 0.006162f
C3834 vdd.n1859 gnd 0.006162f
C3835 vdd.n1860 gnd 0.006162f
C3836 vdd.n1861 gnd 0.006162f
C3837 vdd.n1862 gnd 0.006162f
C3838 vdd.n1863 gnd 0.006162f
C3839 vdd.n1864 gnd 0.006162f
C3840 vdd.n1865 gnd 0.006162f
C3841 vdd.n1866 gnd 0.006162f
C3842 vdd.n1867 gnd 0.006162f
C3843 vdd.n1868 gnd 0.006162f
C3844 vdd.n1869 gnd 0.006162f
C3845 vdd.n1870 gnd 0.006162f
C3846 vdd.n1871 gnd 0.199094f
C3847 vdd.n1872 gnd 0.006162f
C3848 vdd.n1873 gnd 0.006162f
C3849 vdd.n1874 gnd 0.006162f
C3850 vdd.n1875 gnd 0.006162f
C3851 vdd.n1876 gnd 0.006162f
C3852 vdd.n1877 gnd 0.006162f
C3853 vdd.n1878 gnd 0.006162f
C3854 vdd.n1879 gnd 0.006162f
C3855 vdd.n1880 gnd 0.006162f
C3856 vdd.n1881 gnd 0.006162f
C3857 vdd.n1882 gnd 0.006162f
C3858 vdd.n1883 gnd 0.006162f
C3859 vdd.n1884 gnd 0.006162f
C3860 vdd.n1885 gnd 0.006162f
C3861 vdd.n1886 gnd 0.006162f
C3862 vdd.n1887 gnd 0.006162f
C3863 vdd.n1888 gnd 0.006162f
C3864 vdd.n1889 gnd 0.006162f
C3865 vdd.n1890 gnd 0.006162f
C3866 vdd.n1891 gnd 0.006162f
C3867 vdd.n1892 gnd 0.013651f
C3868 vdd.n1894 gnd 0.014621f
C3869 vdd.n1895 gnd 0.014621f
C3870 vdd.n1896 gnd 0.006162f
C3871 vdd.n1897 gnd 0.004757f
C3872 vdd.n1898 gnd 0.006162f
C3873 vdd.n1900 gnd 0.006162f
C3874 vdd.n1902 gnd 0.006162f
C3875 vdd.n1903 gnd 0.006162f
C3876 vdd.n1904 gnd 0.006162f
C3877 vdd.n1905 gnd 0.006162f
C3878 vdd.n1906 gnd 0.006162f
C3879 vdd.n1908 gnd 0.006162f
C3880 vdd.n1910 gnd 0.006162f
C3881 vdd.n1911 gnd 0.006162f
C3882 vdd.n1912 gnd 0.006162f
C3883 vdd.n1913 gnd 0.006162f
C3884 vdd.n1914 gnd 0.006162f
C3885 vdd.n1916 gnd 0.006162f
C3886 vdd.n1918 gnd 0.006162f
C3887 vdd.n1919 gnd 0.006162f
C3888 vdd.n1920 gnd 0.006162f
C3889 vdd.n1921 gnd 0.006162f
C3890 vdd.n1922 gnd 0.006162f
C3891 vdd.n1924 gnd 0.006162f
C3892 vdd.n1926 gnd 0.006162f
C3893 vdd.n1927 gnd 0.006162f
C3894 vdd.n1928 gnd 0.018379f
C3895 vdd.n1929 gnd 0.54483f
C3896 vdd.n1931 gnd 0.007293f
C3897 vdd.n1932 gnd 0.007293f
C3898 vdd.n1933 gnd 0.009061f
C3899 vdd.n1935 gnd 0.009061f
C3900 vdd.n1936 gnd 0.009061f
C3901 vdd.n1937 gnd 0.007293f
C3902 vdd.n1938 gnd 0.006053f
C3903 vdd.n1939 gnd 0.022589f
C3904 vdd.n1940 gnd 0.022083f
C3905 vdd.n1941 gnd 0.006053f
C3906 vdd.n1942 gnd 0.022083f
C3907 vdd.n1943 gnd 1.27328f
C3908 vdd.n1944 gnd 0.022083f
C3909 vdd.n1945 gnd 0.022589f
C3910 vdd.n1946 gnd 0.003464f
C3911 vdd.t42 gnd 0.111477f
C3912 vdd.t41 gnd 0.119139f
C3913 vdd.t39 gnd 0.145588f
C3914 vdd.n1947 gnd 0.186623f
C3915 vdd.n1948 gnd 0.156797f
C3916 vdd.n1949 gnd 0.011232f
C3917 vdd.n1950 gnd 0.003829f
C3918 vdd.n1951 gnd 0.007793f
C3919 vdd.n1952 gnd 0.54483f
C3920 vdd.n1953 gnd 0.018379f
C3921 vdd.n1954 gnd 0.006162f
C3922 vdd.n1955 gnd 0.006162f
C3923 vdd.n1956 gnd 0.006162f
C3924 vdd.n1958 gnd 0.006162f
C3925 vdd.n1960 gnd 0.006162f
C3926 vdd.n1961 gnd 0.006162f
C3927 vdd.n1962 gnd 0.006162f
C3928 vdd.n1963 gnd 0.006162f
C3929 vdd.n1964 gnd 0.006162f
C3930 vdd.n1966 gnd 0.006162f
C3931 vdd.n1968 gnd 0.006162f
C3932 vdd.n1969 gnd 0.006162f
C3933 vdd.n1970 gnd 0.006162f
C3934 vdd.n1971 gnd 0.006162f
C3935 vdd.n1972 gnd 0.006162f
C3936 vdd.n1974 gnd 0.006162f
C3937 vdd.n1976 gnd 0.006162f
C3938 vdd.n1977 gnd 0.006162f
C3939 vdd.n1978 gnd 0.006162f
C3940 vdd.n1979 gnd 0.006162f
C3941 vdd.n1980 gnd 0.006162f
C3942 vdd.n1982 gnd 0.006162f
C3943 vdd.n1984 gnd 0.006162f
C3944 vdd.n1985 gnd 0.006162f
C3945 vdd.n1986 gnd 0.014621f
C3946 vdd.n1987 gnd 0.013651f
C3947 vdd.n1988 gnd 0.013651f
C3948 vdd.n1989 gnd 0.907498f
C3949 vdd.n1990 gnd 0.013651f
C3950 vdd.n1991 gnd 0.013651f
C3951 vdd.n1992 gnd 0.006162f
C3952 vdd.n1993 gnd 0.006162f
C3953 vdd.n1994 gnd 0.006162f
C3954 vdd.n1995 gnd 0.393558f
C3955 vdd.n1996 gnd 0.006162f
C3956 vdd.n1997 gnd 0.006162f
C3957 vdd.n1998 gnd 0.006162f
C3958 vdd.n1999 gnd 0.006162f
C3959 vdd.n2000 gnd 0.006162f
C3960 vdd.n2001 gnd 0.629692f
C3961 vdd.n2002 gnd 0.006162f
C3962 vdd.n2003 gnd 0.006162f
C3963 vdd.n2004 gnd 0.006162f
C3964 vdd.n2005 gnd 0.006162f
C3965 vdd.n2006 gnd 0.006162f
C3966 vdd.n2007 gnd 0.629692f
C3967 vdd.n2008 gnd 0.006162f
C3968 vdd.n2009 gnd 0.006162f
C3969 vdd.n2010 gnd 0.005437f
C3970 vdd.n2011 gnd 0.01785f
C3971 vdd.n2012 gnd 0.003806f
C3972 vdd.n2013 gnd 0.006162f
C3973 vdd.n2014 gnd 0.347257f
C3974 vdd.n2015 gnd 0.006162f
C3975 vdd.n2016 gnd 0.006162f
C3976 vdd.n2017 gnd 0.006162f
C3977 vdd.n2018 gnd 0.006162f
C3978 vdd.n2019 gnd 0.006162f
C3979 vdd.n2020 gnd 0.421338f
C3980 vdd.n2021 gnd 0.006162f
C3981 vdd.n2022 gnd 0.006162f
C3982 vdd.n2023 gnd 0.006162f
C3983 vdd.n2024 gnd 0.006162f
C3984 vdd.n2025 gnd 0.006162f
C3985 vdd.n2026 gnd 0.560241f
C3986 vdd.n2027 gnd 0.006162f
C3987 vdd.n2028 gnd 0.006162f
C3988 vdd.n2029 gnd 0.006162f
C3989 vdd.n2030 gnd 0.006162f
C3990 vdd.n2031 gnd 0.006162f
C3991 vdd.n2032 gnd 0.50005f
C3992 vdd.n2033 gnd 0.006162f
C3993 vdd.n2034 gnd 0.006162f
C3994 vdd.n2035 gnd 0.006162f
C3995 vdd.n2036 gnd 0.006162f
C3996 vdd.n2037 gnd 0.006162f
C3997 vdd.n2038 gnd 0.361147f
C3998 vdd.n2039 gnd 0.006162f
C3999 vdd.n2040 gnd 0.006162f
C4000 vdd.n2041 gnd 0.006162f
C4001 vdd.n2042 gnd 0.006162f
C4002 vdd.n2043 gnd 0.006162f
C4003 vdd.n2044 gnd 0.199094f
C4004 vdd.n2045 gnd 0.006162f
C4005 vdd.n2046 gnd 0.006162f
C4006 vdd.n2047 gnd 0.006162f
C4007 vdd.n2048 gnd 0.006162f
C4008 vdd.n2049 gnd 0.006162f
C4009 vdd.n2050 gnd 0.347257f
C4010 vdd.n2051 gnd 0.006162f
C4011 vdd.n2052 gnd 0.006162f
C4012 vdd.n2053 gnd 0.006162f
C4013 vdd.n2054 gnd 0.006162f
C4014 vdd.n2055 gnd 0.006162f
C4015 vdd.n2056 gnd 0.629692f
C4016 vdd.n2057 gnd 0.006162f
C4017 vdd.n2058 gnd 0.006162f
C4018 vdd.n2059 gnd 0.006162f
C4019 vdd.n2060 gnd 0.006162f
C4020 vdd.n2061 gnd 0.006162f
C4021 vdd.n2062 gnd 0.006162f
C4022 vdd.n2063 gnd 0.006162f
C4023 vdd.n2064 gnd 0.49079f
C4024 vdd.n2065 gnd 0.006162f
C4025 vdd.n2066 gnd 0.006162f
C4026 vdd.n2067 gnd 0.006162f
C4027 vdd.n2068 gnd 0.006162f
C4028 vdd.n2069 gnd 0.006162f
C4029 vdd.n2070 gnd 0.006162f
C4030 vdd.n2071 gnd 0.393558f
C4031 vdd.n2072 gnd 0.006162f
C4032 vdd.n2073 gnd 0.006162f
C4033 vdd.n2074 gnd 0.006162f
C4034 vdd.n2075 gnd 0.014401f
C4035 vdd.n2076 gnd 0.01387f
C4036 vdd.n2077 gnd 0.006162f
C4037 vdd.n2078 gnd 0.006162f
C4038 vdd.n2079 gnd 0.004757f
C4039 vdd.n2080 gnd 0.006162f
C4040 vdd.n2081 gnd 0.006162f
C4041 vdd.n2082 gnd 0.004485f
C4042 vdd.n2083 gnd 0.006162f
C4043 vdd.n2084 gnd 0.006162f
C4044 vdd.n2085 gnd 0.006162f
C4045 vdd.n2086 gnd 0.006162f
C4046 vdd.n2087 gnd 0.006162f
C4047 vdd.n2088 gnd 0.006162f
C4048 vdd.n2089 gnd 0.006162f
C4049 vdd.n2090 gnd 0.006162f
C4050 vdd.n2091 gnd 0.006162f
C4051 vdd.n2092 gnd 0.006162f
C4052 vdd.n2093 gnd 0.006162f
C4053 vdd.n2094 gnd 0.006162f
C4054 vdd.n2095 gnd 0.006162f
C4055 vdd.n2096 gnd 0.006162f
C4056 vdd.n2097 gnd 0.006162f
C4057 vdd.n2098 gnd 0.006162f
C4058 vdd.n2099 gnd 0.006162f
C4059 vdd.n2100 gnd 0.006162f
C4060 vdd.n2101 gnd 0.006162f
C4061 vdd.n2102 gnd 0.006162f
C4062 vdd.n2103 gnd 0.006162f
C4063 vdd.n2104 gnd 0.006162f
C4064 vdd.n2105 gnd 0.006162f
C4065 vdd.n2106 gnd 0.006162f
C4066 vdd.n2107 gnd 0.006162f
C4067 vdd.n2108 gnd 0.006162f
C4068 vdd.n2109 gnd 0.006162f
C4069 vdd.n2110 gnd 0.006162f
C4070 vdd.n2111 gnd 0.006162f
C4071 vdd.n2112 gnd 0.006162f
C4072 vdd.n2113 gnd 0.006162f
C4073 vdd.n2114 gnd 0.006162f
C4074 vdd.n2115 gnd 0.006162f
C4075 vdd.n2116 gnd 0.006162f
C4076 vdd.n2117 gnd 0.006162f
C4077 vdd.n2118 gnd 0.006162f
C4078 vdd.n2119 gnd 0.006162f
C4079 vdd.n2120 gnd 0.006162f
C4080 vdd.n2121 gnd 0.006162f
C4081 vdd.n2122 gnd 0.006162f
C4082 vdd.n2123 gnd 0.006162f
C4083 vdd.n2124 gnd 0.006162f
C4084 vdd.n2125 gnd 0.006162f
C4085 vdd.n2126 gnd 0.006162f
C4086 vdd.n2127 gnd 0.006162f
C4087 vdd.n2128 gnd 0.006162f
C4088 vdd.n2129 gnd 0.006162f
C4089 vdd.n2130 gnd 0.006162f
C4090 vdd.n2131 gnd 0.006162f
C4091 vdd.n2132 gnd 0.006162f
C4092 vdd.n2133 gnd 0.006162f
C4093 vdd.n2134 gnd 0.006162f
C4094 vdd.n2135 gnd 0.006162f
C4095 vdd.n2136 gnd 0.006162f
C4096 vdd.n2137 gnd 0.006162f
C4097 vdd.n2138 gnd 0.006162f
C4098 vdd.n2139 gnd 0.006162f
C4099 vdd.n2140 gnd 0.006162f
C4100 vdd.n2141 gnd 0.006162f
C4101 vdd.n2142 gnd 0.006162f
C4102 vdd.n2143 gnd 0.014621f
C4103 vdd.n2144 gnd 0.013651f
C4104 vdd.n2145 gnd 0.013651f
C4105 vdd.n2146 gnd 0.768595f
C4106 vdd.n2147 gnd 0.013651f
C4107 vdd.n2148 gnd 0.014621f
C4108 vdd.n2149 gnd 0.01387f
C4109 vdd.n2150 gnd 0.006162f
C4110 vdd.n2151 gnd 0.006162f
C4111 vdd.n2152 gnd 0.006162f
C4112 vdd.n2153 gnd 0.004757f
C4113 vdd.n2154 gnd 0.008806f
C4114 vdd.n2155 gnd 0.004485f
C4115 vdd.n2156 gnd 0.006162f
C4116 vdd.n2157 gnd 0.006162f
C4117 vdd.n2158 gnd 0.006162f
C4118 vdd.n2159 gnd 0.006162f
C4119 vdd.n2160 gnd 0.006162f
C4120 vdd.n2161 gnd 0.006162f
C4121 vdd.n2162 gnd 0.006162f
C4122 vdd.n2163 gnd 0.006162f
C4123 vdd.n2164 gnd 0.006162f
C4124 vdd.n2165 gnd 0.006162f
C4125 vdd.n2166 gnd 0.006162f
C4126 vdd.n2167 gnd 0.006162f
C4127 vdd.n2168 gnd 0.006162f
C4128 vdd.n2169 gnd 0.006162f
C4129 vdd.n2170 gnd 0.006162f
C4130 vdd.n2171 gnd 0.006162f
C4131 vdd.n2172 gnd 0.006162f
C4132 vdd.n2173 gnd 0.006162f
C4133 vdd.n2174 gnd 0.006162f
C4134 vdd.n2175 gnd 0.006162f
C4135 vdd.n2176 gnd 0.006162f
C4136 vdd.n2177 gnd 0.006162f
C4137 vdd.n2178 gnd 0.006162f
C4138 vdd.n2179 gnd 0.006162f
C4139 vdd.n2180 gnd 0.006162f
C4140 vdd.n2181 gnd 0.006162f
C4141 vdd.n2182 gnd 0.006162f
C4142 vdd.n2183 gnd 0.006162f
C4143 vdd.n2184 gnd 0.006162f
C4144 vdd.n2185 gnd 0.006162f
C4145 vdd.n2186 gnd 0.006162f
C4146 vdd.n2187 gnd 0.006162f
C4147 vdd.n2188 gnd 0.006162f
C4148 vdd.n2189 gnd 0.006162f
C4149 vdd.n2190 gnd 0.006162f
C4150 vdd.n2191 gnd 0.006162f
C4151 vdd.n2192 gnd 0.006162f
C4152 vdd.n2193 gnd 0.006162f
C4153 vdd.n2194 gnd 0.006162f
C4154 vdd.n2195 gnd 0.006162f
C4155 vdd.n2196 gnd 0.006162f
C4156 vdd.n2197 gnd 0.006162f
C4157 vdd.n2198 gnd 0.006162f
C4158 vdd.n2199 gnd 0.006162f
C4159 vdd.n2200 gnd 0.006162f
C4160 vdd.n2201 gnd 0.006162f
C4161 vdd.n2202 gnd 0.006162f
C4162 vdd.n2203 gnd 0.006162f
C4163 vdd.n2204 gnd 0.006162f
C4164 vdd.n2205 gnd 0.006162f
C4165 vdd.n2206 gnd 0.006162f
C4166 vdd.n2207 gnd 0.006162f
C4167 vdd.n2208 gnd 0.006162f
C4168 vdd.n2209 gnd 0.006162f
C4169 vdd.n2210 gnd 0.006162f
C4170 vdd.n2211 gnd 0.006162f
C4171 vdd.n2212 gnd 0.006162f
C4172 vdd.n2213 gnd 0.006162f
C4173 vdd.n2214 gnd 0.006162f
C4174 vdd.n2215 gnd 0.006162f
C4175 vdd.n2216 gnd 0.014621f
C4176 vdd.n2217 gnd 0.014621f
C4177 vdd.n2218 gnd 0.768595f
C4178 vdd.t118 gnd 2.73175f
C4179 vdd.t22 gnd 2.73175f
C4180 vdd.n2251 gnd 0.014621f
C4181 vdd.n2252 gnd 0.006162f
C4182 vdd.t74 gnd 0.248992f
C4183 vdd.t75 gnd 0.254874f
C4184 vdd.t72 gnd 0.162551f
C4185 vdd.n2253 gnd 0.08785f
C4186 vdd.n2254 gnd 0.049831f
C4187 vdd.n2255 gnd 0.006162f
C4188 vdd.t88 gnd 0.248992f
C4189 vdd.t89 gnd 0.254874f
C4190 vdd.t87 gnd 0.162551f
C4191 vdd.n2256 gnd 0.08785f
C4192 vdd.n2257 gnd 0.049831f
C4193 vdd.n2258 gnd 0.008806f
C4194 vdd.n2259 gnd 0.006162f
C4195 vdd.n2260 gnd 0.006162f
C4196 vdd.n2261 gnd 0.006162f
C4197 vdd.n2262 gnd 0.006162f
C4198 vdd.n2263 gnd 0.006162f
C4199 vdd.n2264 gnd 0.006162f
C4200 vdd.n2265 gnd 0.006162f
C4201 vdd.n2266 gnd 0.006162f
C4202 vdd.n2267 gnd 0.006162f
C4203 vdd.n2268 gnd 0.006162f
C4204 vdd.n2269 gnd 0.006162f
C4205 vdd.n2270 gnd 0.006162f
C4206 vdd.n2271 gnd 0.006162f
C4207 vdd.n2272 gnd 0.006162f
C4208 vdd.n2273 gnd 0.006162f
C4209 vdd.n2274 gnd 0.006162f
C4210 vdd.n2275 gnd 0.006162f
C4211 vdd.n2276 gnd 0.006162f
C4212 vdd.n2277 gnd 0.006162f
C4213 vdd.n2278 gnd 0.006162f
C4214 vdd.n2279 gnd 0.006162f
C4215 vdd.n2280 gnd 0.006162f
C4216 vdd.n2281 gnd 0.006162f
C4217 vdd.n2282 gnd 0.006162f
C4218 vdd.n2283 gnd 0.006162f
C4219 vdd.n2284 gnd 0.006162f
C4220 vdd.n2285 gnd 0.006162f
C4221 vdd.n2286 gnd 0.006162f
C4222 vdd.n2287 gnd 0.006162f
C4223 vdd.n2288 gnd 0.006162f
C4224 vdd.n2289 gnd 0.006162f
C4225 vdd.n2290 gnd 0.006162f
C4226 vdd.n2291 gnd 0.006162f
C4227 vdd.n2292 gnd 0.006162f
C4228 vdd.n2293 gnd 0.006162f
C4229 vdd.n2294 gnd 0.006162f
C4230 vdd.n2295 gnd 0.006162f
C4231 vdd.n2296 gnd 0.006162f
C4232 vdd.n2297 gnd 0.006162f
C4233 vdd.n2298 gnd 0.006162f
C4234 vdd.n2299 gnd 0.006162f
C4235 vdd.n2300 gnd 0.006162f
C4236 vdd.n2301 gnd 0.006162f
C4237 vdd.n2302 gnd 0.006162f
C4238 vdd.n2303 gnd 0.006162f
C4239 vdd.n2304 gnd 0.006162f
C4240 vdd.n2305 gnd 0.006162f
C4241 vdd.n2306 gnd 0.006162f
C4242 vdd.n2307 gnd 0.006162f
C4243 vdd.n2308 gnd 0.006162f
C4244 vdd.n2309 gnd 0.006162f
C4245 vdd.n2310 gnd 0.006162f
C4246 vdd.n2311 gnd 0.006162f
C4247 vdd.n2312 gnd 0.006162f
C4248 vdd.n2313 gnd 0.006162f
C4249 vdd.n2314 gnd 0.006162f
C4250 vdd.n2315 gnd 0.004485f
C4251 vdd.n2316 gnd 0.006162f
C4252 vdd.n2317 gnd 0.006162f
C4253 vdd.n2318 gnd 0.004757f
C4254 vdd.n2319 gnd 0.006162f
C4255 vdd.n2320 gnd 0.006162f
C4256 vdd.n2321 gnd 0.014621f
C4257 vdd.n2322 gnd 0.013651f
C4258 vdd.n2323 gnd 0.006162f
C4259 vdd.n2324 gnd 0.006162f
C4260 vdd.n2325 gnd 0.006162f
C4261 vdd.n2326 gnd 0.006162f
C4262 vdd.n2327 gnd 0.006162f
C4263 vdd.n2328 gnd 0.006162f
C4264 vdd.n2329 gnd 0.006162f
C4265 vdd.n2330 gnd 0.006162f
C4266 vdd.n2331 gnd 0.006162f
C4267 vdd.n2332 gnd 0.006162f
C4268 vdd.n2333 gnd 0.006162f
C4269 vdd.n2334 gnd 0.006162f
C4270 vdd.n2335 gnd 0.006162f
C4271 vdd.n2336 gnd 0.006162f
C4272 vdd.n2337 gnd 0.006162f
C4273 vdd.n2338 gnd 0.006162f
C4274 vdd.n2339 gnd 0.006162f
C4275 vdd.n2340 gnd 0.006162f
C4276 vdd.n2341 gnd 0.006162f
C4277 vdd.n2342 gnd 0.006162f
C4278 vdd.n2343 gnd 0.006162f
C4279 vdd.n2344 gnd 0.006162f
C4280 vdd.n2345 gnd 0.006162f
C4281 vdd.n2346 gnd 0.006162f
C4282 vdd.n2347 gnd 0.006162f
C4283 vdd.n2348 gnd 0.006162f
C4284 vdd.n2349 gnd 0.006162f
C4285 vdd.n2350 gnd 0.006162f
C4286 vdd.n2351 gnd 0.006162f
C4287 vdd.n2352 gnd 0.006162f
C4288 vdd.n2353 gnd 0.006162f
C4289 vdd.n2354 gnd 0.006162f
C4290 vdd.n2355 gnd 0.006162f
C4291 vdd.n2356 gnd 0.006162f
C4292 vdd.n2357 gnd 0.006162f
C4293 vdd.n2358 gnd 0.006162f
C4294 vdd.n2359 gnd 0.006162f
C4295 vdd.n2360 gnd 0.006162f
C4296 vdd.n2361 gnd 0.006162f
C4297 vdd.n2362 gnd 0.006162f
C4298 vdd.n2363 gnd 0.006162f
C4299 vdd.n2364 gnd 0.006162f
C4300 vdd.n2365 gnd 0.006162f
C4301 vdd.n2366 gnd 0.006162f
C4302 vdd.n2367 gnd 0.006162f
C4303 vdd.n2368 gnd 0.006162f
C4304 vdd.n2369 gnd 0.006162f
C4305 vdd.n2370 gnd 0.006162f
C4306 vdd.n2371 gnd 0.006162f
C4307 vdd.n2372 gnd 0.006162f
C4308 vdd.n2373 gnd 0.006162f
C4309 vdd.n2374 gnd 0.199094f
C4310 vdd.n2375 gnd 0.006162f
C4311 vdd.n2376 gnd 0.006162f
C4312 vdd.n2377 gnd 0.006162f
C4313 vdd.n2378 gnd 0.006162f
C4314 vdd.n2379 gnd 0.006162f
C4315 vdd.n2380 gnd 0.006162f
C4316 vdd.n2381 gnd 0.006162f
C4317 vdd.n2382 gnd 0.006162f
C4318 vdd.n2383 gnd 0.006162f
C4319 vdd.n2384 gnd 0.006162f
C4320 vdd.n2385 gnd 0.006162f
C4321 vdd.n2386 gnd 0.006162f
C4322 vdd.n2387 gnd 0.006162f
C4323 vdd.n2388 gnd 0.006162f
C4324 vdd.n2389 gnd 0.006162f
C4325 vdd.n2390 gnd 0.006162f
C4326 vdd.n2391 gnd 0.006162f
C4327 vdd.n2392 gnd 0.006162f
C4328 vdd.n2393 gnd 0.006162f
C4329 vdd.n2394 gnd 0.006162f
C4330 vdd.n2395 gnd 0.375037f
C4331 vdd.n2396 gnd 0.006162f
C4332 vdd.n2397 gnd 0.006162f
C4333 vdd.n2398 gnd 0.006162f
C4334 vdd.n2399 gnd 0.006162f
C4335 vdd.n2400 gnd 0.006162f
C4336 vdd.n2401 gnd 0.013651f
C4337 vdd.n2402 gnd 0.014621f
C4338 vdd.n2403 gnd 0.014621f
C4339 vdd.n2404 gnd 0.006162f
C4340 vdd.n2405 gnd 0.006162f
C4341 vdd.n2406 gnd 0.006162f
C4342 vdd.n2407 gnd 0.004757f
C4343 vdd.n2408 gnd 0.008806f
C4344 vdd.n2409 gnd 0.004485f
C4345 vdd.n2410 gnd 0.006162f
C4346 vdd.n2411 gnd 0.006162f
C4347 vdd.n2412 gnd 0.006162f
C4348 vdd.n2413 gnd 0.006162f
C4349 vdd.n2414 gnd 0.006162f
C4350 vdd.n2415 gnd 0.006162f
C4351 vdd.n2416 gnd 0.006162f
C4352 vdd.n2417 gnd 0.006162f
C4353 vdd.n2418 gnd 0.006162f
C4354 vdd.n2419 gnd 0.006162f
C4355 vdd.n2420 gnd 0.006162f
C4356 vdd.n2421 gnd 0.006162f
C4357 vdd.n2422 gnd 0.006162f
C4358 vdd.n2423 gnd 0.006162f
C4359 vdd.n2424 gnd 0.006162f
C4360 vdd.n2425 gnd 0.006162f
C4361 vdd.n2426 gnd 0.006162f
C4362 vdd.n2427 gnd 0.006162f
C4363 vdd.n2428 gnd 0.006162f
C4364 vdd.n2429 gnd 0.006162f
C4365 vdd.n2430 gnd 0.006162f
C4366 vdd.n2431 gnd 0.006162f
C4367 vdd.n2432 gnd 0.006162f
C4368 vdd.n2433 gnd 0.006162f
C4369 vdd.n2434 gnd 0.006162f
C4370 vdd.n2435 gnd 0.006162f
C4371 vdd.n2436 gnd 0.006162f
C4372 vdd.n2437 gnd 0.006162f
C4373 vdd.n2438 gnd 0.006162f
C4374 vdd.n2439 gnd 0.006162f
C4375 vdd.n2440 gnd 0.006162f
C4376 vdd.n2441 gnd 0.006162f
C4377 vdd.n2442 gnd 0.006162f
C4378 vdd.n2443 gnd 0.006162f
C4379 vdd.n2444 gnd 0.006162f
C4380 vdd.n2445 gnd 0.006162f
C4381 vdd.n2446 gnd 0.006162f
C4382 vdd.n2447 gnd 0.006162f
C4383 vdd.n2448 gnd 0.006162f
C4384 vdd.n2449 gnd 0.006162f
C4385 vdd.n2450 gnd 0.006162f
C4386 vdd.n2451 gnd 0.006162f
C4387 vdd.n2452 gnd 0.006162f
C4388 vdd.n2453 gnd 0.006162f
C4389 vdd.n2454 gnd 0.006162f
C4390 vdd.n2455 gnd 0.006162f
C4391 vdd.n2456 gnd 0.006162f
C4392 vdd.n2457 gnd 0.006162f
C4393 vdd.n2458 gnd 0.006162f
C4394 vdd.n2459 gnd 0.006162f
C4395 vdd.n2460 gnd 0.006162f
C4396 vdd.n2461 gnd 0.006162f
C4397 vdd.n2462 gnd 0.006162f
C4398 vdd.n2463 gnd 0.006162f
C4399 vdd.n2464 gnd 0.006162f
C4400 vdd.n2465 gnd 0.006162f
C4401 vdd.n2466 gnd 0.006162f
C4402 vdd.n2467 gnd 0.006162f
C4403 vdd.n2468 gnd 0.006162f
C4404 vdd.n2469 gnd 0.006162f
C4405 vdd.n2471 gnd 0.768595f
C4406 vdd.n2473 gnd 0.006162f
C4407 vdd.n2474 gnd 0.006162f
C4408 vdd.n2475 gnd 0.014621f
C4409 vdd.n2476 gnd 0.013651f
C4410 vdd.n2477 gnd 0.013651f
C4411 vdd.n2478 gnd 0.768595f
C4412 vdd.n2479 gnd 0.013651f
C4413 vdd.n2480 gnd 0.013651f
C4414 vdd.n2481 gnd 0.006162f
C4415 vdd.n2482 gnd 0.006162f
C4416 vdd.n2483 gnd 0.006162f
C4417 vdd.n2484 gnd 0.393558f
C4418 vdd.n2485 gnd 0.006162f
C4419 vdd.n2486 gnd 0.006162f
C4420 vdd.n2487 gnd 0.006162f
C4421 vdd.n2488 gnd 0.006162f
C4422 vdd.n2489 gnd 0.006162f
C4423 vdd.n2490 gnd 0.49079f
C4424 vdd.n2491 gnd 0.006162f
C4425 vdd.n2492 gnd 0.006162f
C4426 vdd.n2493 gnd 0.006162f
C4427 vdd.n2494 gnd 0.006162f
C4428 vdd.n2495 gnd 0.006162f
C4429 vdd.n2496 gnd 0.629692f
C4430 vdd.n2497 gnd 0.006162f
C4431 vdd.n2498 gnd 0.006162f
C4432 vdd.n2499 gnd 0.006162f
C4433 vdd.n2500 gnd 0.006162f
C4434 vdd.n2501 gnd 0.006162f
C4435 vdd.n2502 gnd 0.347257f
C4436 vdd.n2503 gnd 0.006162f
C4437 vdd.n2504 gnd 0.006162f
C4438 vdd.n2505 gnd 0.006162f
C4439 vdd.n2506 gnd 0.006162f
C4440 vdd.n2507 gnd 0.006162f
C4441 vdd.n2508 gnd 0.199094f
C4442 vdd.n2509 gnd 0.006162f
C4443 vdd.n2510 gnd 0.006162f
C4444 vdd.n2511 gnd 0.006162f
C4445 vdd.n2512 gnd 0.006162f
C4446 vdd.n2513 gnd 0.006162f
C4447 vdd.n2514 gnd 0.361147f
C4448 vdd.n2515 gnd 0.006162f
C4449 vdd.n2516 gnd 0.006162f
C4450 vdd.n2517 gnd 0.006162f
C4451 vdd.n2518 gnd 0.006162f
C4452 vdd.n2519 gnd 0.006162f
C4453 vdd.n2520 gnd 0.50005f
C4454 vdd.n2521 gnd 0.006162f
C4455 vdd.n2522 gnd 0.006162f
C4456 vdd.n2523 gnd 0.006162f
C4457 vdd.n2524 gnd 0.006162f
C4458 vdd.n2525 gnd 0.006162f
C4459 vdd.n2526 gnd 0.560241f
C4460 vdd.n2527 gnd 0.006162f
C4461 vdd.n2528 gnd 0.006162f
C4462 vdd.n2529 gnd 0.006162f
C4463 vdd.n2530 gnd 0.006162f
C4464 vdd.n2531 gnd 0.006162f
C4465 vdd.n2532 gnd 0.421338f
C4466 vdd.n2533 gnd 0.006162f
C4467 vdd.n2534 gnd 0.006162f
C4468 vdd.n2535 gnd 0.006162f
C4469 vdd.t49 gnd 0.254874f
C4470 vdd.t47 gnd 0.162551f
C4471 vdd.t50 gnd 0.254874f
C4472 vdd.n2536 gnd 0.14325f
C4473 vdd.n2537 gnd 0.01785f
C4474 vdd.n2538 gnd 0.003806f
C4475 vdd.n2539 gnd 0.006162f
C4476 vdd.n2540 gnd 0.347257f
C4477 vdd.n2541 gnd 0.006162f
C4478 vdd.n2542 gnd 0.006162f
C4479 vdd.n2543 gnd 0.006162f
C4480 vdd.n2544 gnd 0.006162f
C4481 vdd.n2545 gnd 0.006162f
C4482 vdd.n2546 gnd 0.629692f
C4483 vdd.n2547 gnd 0.006162f
C4484 vdd.n2548 gnd 0.006162f
C4485 vdd.n2549 gnd 0.006162f
C4486 vdd.n2550 gnd 0.006162f
C4487 vdd.n2551 gnd 0.006162f
C4488 vdd.n2552 gnd 0.006162f
C4489 vdd.n2554 gnd 0.006162f
C4490 vdd.n2555 gnd 0.006162f
C4491 vdd.n2557 gnd 0.006162f
C4492 vdd.n2558 gnd 0.006162f
C4493 vdd.n2561 gnd 0.006162f
C4494 vdd.n2562 gnd 0.006162f
C4495 vdd.n2563 gnd 0.006162f
C4496 vdd.n2564 gnd 0.006162f
C4497 vdd.n2566 gnd 0.006162f
C4498 vdd.n2567 gnd 0.006162f
C4499 vdd.n2568 gnd 0.006162f
C4500 vdd.n2569 gnd 0.006162f
C4501 vdd.n2570 gnd 0.006162f
C4502 vdd.n2571 gnd 0.006162f
C4503 vdd.n2573 gnd 0.006162f
C4504 vdd.n2574 gnd 0.006162f
C4505 vdd.n2575 gnd 0.006162f
C4506 vdd.n2576 gnd 0.006162f
C4507 vdd.n2577 gnd 0.006162f
C4508 vdd.n2578 gnd 0.006162f
C4509 vdd.n2580 gnd 0.006162f
C4510 vdd.n2581 gnd 0.006162f
C4511 vdd.n2582 gnd 0.006162f
C4512 vdd.n2583 gnd 0.006162f
C4513 vdd.n2584 gnd 0.006162f
C4514 vdd.n2585 gnd 0.006162f
C4515 vdd.n2587 gnd 0.006162f
C4516 vdd.n2588 gnd 0.014621f
C4517 vdd.n2589 gnd 0.014621f
C4518 vdd.n2590 gnd 0.013651f
C4519 vdd.n2591 gnd 0.006162f
C4520 vdd.n2592 gnd 0.006162f
C4521 vdd.n2593 gnd 0.006162f
C4522 vdd.n2594 gnd 0.006162f
C4523 vdd.n2595 gnd 0.006162f
C4524 vdd.n2596 gnd 0.006162f
C4525 vdd.n2597 gnd 0.629692f
C4526 vdd.n2598 gnd 0.006162f
C4527 vdd.n2599 gnd 0.006162f
C4528 vdd.n2600 gnd 0.006162f
C4529 vdd.n2601 gnd 0.006162f
C4530 vdd.n2602 gnd 0.006162f
C4531 vdd.n2603 gnd 0.393558f
C4532 vdd.n2604 gnd 0.006162f
C4533 vdd.n2605 gnd 0.006162f
C4534 vdd.n2606 gnd 0.006162f
C4535 vdd.n2607 gnd 0.014401f
C4536 vdd.n2608 gnd 0.01387f
C4537 vdd.n2609 gnd 0.014621f
C4538 vdd.n2611 gnd 0.006162f
C4539 vdd.n2612 gnd 0.006162f
C4540 vdd.n2613 gnd 0.004757f
C4541 vdd.n2614 gnd 0.008806f
C4542 vdd.n2615 gnd 0.004485f
C4543 vdd.n2616 gnd 0.006162f
C4544 vdd.n2617 gnd 0.006162f
C4545 vdd.n2619 gnd 0.006162f
C4546 vdd.n2620 gnd 0.006162f
C4547 vdd.n2621 gnd 0.006162f
C4548 vdd.n2622 gnd 0.006162f
C4549 vdd.n2623 gnd 0.006162f
C4550 vdd.n2624 gnd 0.006162f
C4551 vdd.n2626 gnd 0.006162f
C4552 vdd.n2627 gnd 0.006162f
C4553 vdd.n2628 gnd 0.006162f
C4554 vdd.n2629 gnd 0.006162f
C4555 vdd.n2630 gnd 0.006162f
C4556 vdd.n2631 gnd 0.006162f
C4557 vdd.n2633 gnd 0.006162f
C4558 vdd.n2634 gnd 0.006162f
C4559 vdd.n2635 gnd 0.006162f
C4560 vdd.n2636 gnd 0.006162f
C4561 vdd.n2637 gnd 0.006162f
C4562 vdd.n2638 gnd 0.006162f
C4563 vdd.n2640 gnd 0.006162f
C4564 vdd.n2641 gnd 0.006162f
C4565 vdd.n2642 gnd 0.006162f
C4566 vdd.n2644 gnd 0.006162f
C4567 vdd.n2645 gnd 0.006162f
C4568 vdd.n2646 gnd 0.006162f
C4569 vdd.n2647 gnd 0.006162f
C4570 vdd.n2648 gnd 0.006162f
C4571 vdd.n2649 gnd 0.006162f
C4572 vdd.n2651 gnd 0.006162f
C4573 vdd.n2652 gnd 0.006162f
C4574 vdd.n2653 gnd 0.006162f
C4575 vdd.n2654 gnd 0.006162f
C4576 vdd.n2655 gnd 0.006162f
C4577 vdd.n2656 gnd 0.006162f
C4578 vdd.n2658 gnd 0.006162f
C4579 vdd.n2659 gnd 0.006162f
C4580 vdd.n2660 gnd 0.006162f
C4581 vdd.n2661 gnd 0.006162f
C4582 vdd.n2662 gnd 0.006162f
C4583 vdd.n2663 gnd 0.006162f
C4584 vdd.n2665 gnd 0.006162f
C4585 vdd.n2666 gnd 0.006162f
C4586 vdd.n2668 gnd 0.006162f
C4587 vdd.n2669 gnd 0.006162f
C4588 vdd.n2670 gnd 0.014621f
C4589 vdd.n2671 gnd 0.013651f
C4590 vdd.n2672 gnd 0.013651f
C4591 vdd.n2673 gnd 0.907498f
C4592 vdd.n2674 gnd 0.013651f
C4593 vdd.n2675 gnd 0.014621f
C4594 vdd.n2676 gnd 0.01387f
C4595 vdd.n2677 gnd 0.006162f
C4596 vdd.n2678 gnd 0.004757f
C4597 vdd.n2679 gnd 0.006162f
C4598 vdd.n2681 gnd 0.006162f
C4599 vdd.n2682 gnd 0.006162f
C4600 vdd.n2683 gnd 0.006162f
C4601 vdd.n2684 gnd 0.006162f
C4602 vdd.n2685 gnd 0.006162f
C4603 vdd.n2686 gnd 0.006162f
C4604 vdd.n2688 gnd 0.006162f
C4605 vdd.n2689 gnd 0.006162f
C4606 vdd.n2690 gnd 0.006162f
C4607 vdd.n2691 gnd 0.006162f
C4608 vdd.n2692 gnd 0.006162f
C4609 vdd.n2693 gnd 0.006162f
C4610 vdd.n2695 gnd 0.006162f
C4611 vdd.n2696 gnd 0.006162f
C4612 vdd.n2697 gnd 0.006162f
C4613 vdd.n2698 gnd 0.006162f
C4614 vdd.n2699 gnd 0.006162f
C4615 vdd.n2700 gnd 0.006162f
C4616 vdd.n2702 gnd 0.006162f
C4617 vdd.n2703 gnd 0.006162f
C4618 vdd.n2705 gnd 0.006162f
C4619 vdd.n2706 gnd 0.014807f
C4620 vdd.n2707 gnd 0.548403f
C4621 vdd.n2708 gnd 0.007793f
C4622 vdd.n2709 gnd 0.022589f
C4623 vdd.n2710 gnd 0.003464f
C4624 vdd.t100 gnd 0.111477f
C4625 vdd.t101 gnd 0.119139f
C4626 vdd.t99 gnd 0.145588f
C4627 vdd.n2711 gnd 0.186623f
C4628 vdd.n2712 gnd 0.156797f
C4629 vdd.n2713 gnd 0.011232f
C4630 vdd.n2714 gnd 0.009061f
C4631 vdd.n2715 gnd 0.003829f
C4632 vdd.n2716 gnd 0.007293f
C4633 vdd.n2717 gnd 0.009061f
C4634 vdd.n2718 gnd 0.009061f
C4635 vdd.n2719 gnd 0.007293f
C4636 vdd.n2720 gnd 0.007293f
C4637 vdd.n2721 gnd 0.009061f
C4638 vdd.n2722 gnd 0.009061f
C4639 vdd.n2723 gnd 0.007293f
C4640 vdd.n2724 gnd 0.007293f
C4641 vdd.n2725 gnd 0.009061f
C4642 vdd.n2726 gnd 0.009061f
C4643 vdd.n2727 gnd 0.007293f
C4644 vdd.n2728 gnd 0.007293f
C4645 vdd.n2729 gnd 0.009061f
C4646 vdd.n2730 gnd 0.009061f
C4647 vdd.n2731 gnd 0.007293f
C4648 vdd.n2732 gnd 0.007293f
C4649 vdd.n2733 gnd 0.009061f
C4650 vdd.n2734 gnd 0.009061f
C4651 vdd.n2735 gnd 0.007293f
C4652 vdd.n2736 gnd 0.007293f
C4653 vdd.n2737 gnd 0.009061f
C4654 vdd.n2738 gnd 0.009061f
C4655 vdd.n2739 gnd 0.007293f
C4656 vdd.n2740 gnd 0.007293f
C4657 vdd.n2741 gnd 0.009061f
C4658 vdd.n2742 gnd 0.009061f
C4659 vdd.n2743 gnd 0.007293f
C4660 vdd.n2744 gnd 0.007293f
C4661 vdd.n2745 gnd 0.009061f
C4662 vdd.n2746 gnd 0.009061f
C4663 vdd.n2747 gnd 0.007293f
C4664 vdd.n2748 gnd 0.007293f
C4665 vdd.n2749 gnd 0.009061f
C4666 vdd.n2750 gnd 0.009061f
C4667 vdd.n2751 gnd 0.007293f
C4668 vdd.n2752 gnd 0.009061f
C4669 vdd.n2753 gnd 0.009061f
C4670 vdd.n2754 gnd 0.007293f
C4671 vdd.n2755 gnd 0.009061f
C4672 vdd.n2756 gnd 0.009061f
C4673 vdd.n2757 gnd 0.009061f
C4674 vdd.n2758 gnd 0.014878f
C4675 vdd.n2759 gnd 0.009061f
C4676 vdd.n2760 gnd 0.009061f
C4677 vdd.n2761 gnd 0.004959f
C4678 vdd.n2762 gnd 0.007293f
C4679 vdd.n2763 gnd 0.009061f
C4680 vdd.n2764 gnd 0.009061f
C4681 vdd.n2765 gnd 0.007293f
C4682 vdd.n2766 gnd 0.007293f
C4683 vdd.n2767 gnd 0.009061f
C4684 vdd.n2768 gnd 0.009061f
C4685 vdd.n2769 gnd 0.007293f
C4686 vdd.n2770 gnd 0.007293f
C4687 vdd.n2771 gnd 0.009061f
C4688 vdd.n2772 gnd 0.009061f
C4689 vdd.n2773 gnd 0.007293f
C4690 vdd.n2774 gnd 0.007293f
C4691 vdd.n2775 gnd 0.009061f
C4692 vdd.n2776 gnd 0.009061f
C4693 vdd.n2777 gnd 0.007293f
C4694 vdd.n2778 gnd 0.007293f
C4695 vdd.n2779 gnd 0.009061f
C4696 vdd.n2780 gnd 0.009061f
C4697 vdd.n2781 gnd 0.007293f
C4698 vdd.n2782 gnd 0.007293f
C4699 vdd.n2783 gnd 0.009061f
C4700 vdd.n2784 gnd 0.009061f
C4701 vdd.n2785 gnd 0.007293f
C4702 vdd.n2786 gnd 0.007293f
C4703 vdd.n2787 gnd 0.009061f
C4704 vdd.n2788 gnd 0.009061f
C4705 vdd.n2789 gnd 0.007293f
C4706 vdd.n2790 gnd 0.007293f
C4707 vdd.n2791 gnd 0.009061f
C4708 vdd.n2792 gnd 0.009061f
C4709 vdd.n2793 gnd 0.007293f
C4710 vdd.n2794 gnd 0.007293f
C4711 vdd.n2795 gnd 0.009061f
C4712 vdd.n2796 gnd 0.009061f
C4713 vdd.n2797 gnd 0.007293f
C4714 vdd.n2798 gnd 0.009061f
C4715 vdd.n2799 gnd 0.009061f
C4716 vdd.n2800 gnd 0.007293f
C4717 vdd.n2801 gnd 0.009061f
C4718 vdd.n2802 gnd 0.009061f
C4719 vdd.n2803 gnd 0.009061f
C4720 vdd.t37 gnd 0.111477f
C4721 vdd.t38 gnd 0.119139f
C4722 vdd.t36 gnd 0.145588f
C4723 vdd.n2804 gnd 0.186623f
C4724 vdd.n2805 gnd 0.156797f
C4725 vdd.n2806 gnd 0.014878f
C4726 vdd.n2807 gnd 0.009061f
C4727 vdd.n2808 gnd 0.009061f
C4728 vdd.n2809 gnd 0.00609f
C4729 vdd.n2810 gnd 0.007293f
C4730 vdd.n2811 gnd 0.009061f
C4731 vdd.n2812 gnd 0.009061f
C4732 vdd.n2813 gnd 0.007293f
C4733 vdd.n2814 gnd 0.007293f
C4734 vdd.n2815 gnd 0.009061f
C4735 vdd.n2816 gnd 0.009061f
C4736 vdd.n2817 gnd 0.007293f
C4737 vdd.n2818 gnd 0.007293f
C4738 vdd.n2819 gnd 0.009061f
C4739 vdd.n2820 gnd 0.009061f
C4740 vdd.n2821 gnd 0.007293f
C4741 vdd.n2822 gnd 0.007293f
C4742 vdd.n2823 gnd 0.009061f
C4743 vdd.n2824 gnd 0.009061f
C4744 vdd.n2825 gnd 0.007293f
C4745 vdd.n2826 gnd 0.007293f
C4746 vdd.n2827 gnd 0.009061f
C4747 vdd.n2828 gnd 0.009061f
C4748 vdd.n2829 gnd 0.007293f
C4749 vdd.n2830 gnd 0.007293f
C4750 vdd.n2831 gnd 0.009061f
C4751 vdd.n2832 gnd 0.009061f
C4752 vdd.n2833 gnd 0.007293f
C4753 vdd.n2834 gnd 0.007293f
C4754 vdd.n2836 gnd 0.548403f
C4755 vdd.n2838 gnd 0.007293f
C4756 vdd.n2839 gnd 0.009061f
C4757 vdd.n2840 gnd 6.71363f
C4758 vdd.n2842 gnd 0.022589f
C4759 vdd.n2843 gnd 0.006053f
C4760 vdd.n2844 gnd 0.022589f
C4761 vdd.n2845 gnd 0.022083f
C4762 vdd.n2846 gnd 0.009061f
C4763 vdd.n2847 gnd 0.007293f
C4764 vdd.n2848 gnd 0.009061f
C4765 vdd.n2849 gnd 0.578761f
C4766 vdd.n2850 gnd 0.009061f
C4767 vdd.n2851 gnd 0.007293f
C4768 vdd.n2852 gnd 0.009061f
C4769 vdd.n2853 gnd 0.009061f
C4770 vdd.n2854 gnd 0.009061f
C4771 vdd.n2855 gnd 0.007293f
C4772 vdd.n2856 gnd 0.009061f
C4773 vdd.n2857 gnd 0.736185f
C4774 vdd.n2858 gnd 0.926018f
C4775 vdd.n2859 gnd 0.009061f
C4776 vdd.n2860 gnd 0.007293f
C4777 vdd.n2861 gnd 0.009061f
C4778 vdd.n2862 gnd 0.009061f
C4779 vdd.n2863 gnd 0.009061f
C4780 vdd.n2864 gnd 0.007293f
C4781 vdd.n2865 gnd 0.009061f
C4782 vdd.n2866 gnd 0.652843f
C4783 vdd.n2867 gnd 0.009061f
C4784 vdd.n2868 gnd 0.007293f
C4785 vdd.n2869 gnd 0.009061f
C4786 vdd.n2870 gnd 0.009061f
C4787 vdd.n2871 gnd 0.009061f
C4788 vdd.n2872 gnd 0.007293f
C4789 vdd.n2873 gnd 0.009061f
C4790 vdd.t148 gnd 0.463009f
C4791 vdd.n2874 gnd 0.768595f
C4792 vdd.n2875 gnd 0.009061f
C4793 vdd.n2876 gnd 0.007293f
C4794 vdd.n2877 gnd 0.009061f
C4795 vdd.n2878 gnd 0.009061f
C4796 vdd.n2879 gnd 0.009061f
C4797 vdd.n2880 gnd 0.007293f
C4798 vdd.n2881 gnd 0.009061f
C4799 vdd.n2882 gnd 0.726924f
C4800 vdd.n2883 gnd 0.009061f
C4801 vdd.n2884 gnd 0.007293f
C4802 vdd.n2885 gnd 0.009061f
C4803 vdd.n2886 gnd 0.009061f
C4804 vdd.n2887 gnd 0.009061f
C4805 vdd.n2888 gnd 0.007293f
C4806 vdd.n2889 gnd 0.007293f
C4807 vdd.n2890 gnd 0.007293f
C4808 vdd.n2891 gnd 0.009061f
C4809 vdd.n2892 gnd 0.009061f
C4810 vdd.n2893 gnd 0.009061f
C4811 vdd.n2894 gnd 0.007293f
C4812 vdd.n2895 gnd 0.007293f
C4813 vdd.n2896 gnd 0.007293f
C4814 vdd.n2897 gnd 0.009061f
C4815 vdd.n2898 gnd 0.009061f
C4816 vdd.n2899 gnd 0.009061f
C4817 vdd.n2900 gnd 0.007293f
C4818 vdd.n2901 gnd 0.007293f
C4819 vdd.n2902 gnd 0.006053f
C4820 vdd.n2903 gnd 0.022083f
C4821 vdd.n2904 gnd 0.022589f
C4822 vdd.n2906 gnd 0.022589f
C4823 vdd.n2907 gnd 0.003464f
C4824 vdd.t104 gnd 0.111477f
C4825 vdd.t103 gnd 0.119139f
C4826 vdd.t102 gnd 0.145588f
C4827 vdd.n2908 gnd 0.186623f
C4828 vdd.n2909 gnd 0.157527f
C4829 vdd.n2910 gnd 0.011961f
C4830 vdd.n2911 gnd 0.003829f
C4831 vdd.n2912 gnd 0.007293f
C4832 vdd.n2913 gnd 0.009061f
C4833 vdd.n2915 gnd 0.009061f
C4834 vdd.n2916 gnd 0.009061f
C4835 vdd.n2917 gnd 0.007293f
C4836 vdd.n2918 gnd 0.007293f
C4837 vdd.n2919 gnd 0.007293f
C4838 vdd.n2920 gnd 0.009061f
C4839 vdd.n2922 gnd 0.009061f
C4840 vdd.n2923 gnd 0.009061f
C4841 vdd.n2924 gnd 0.007293f
C4842 vdd.n2925 gnd 0.007293f
C4843 vdd.n2926 gnd 0.007293f
C4844 vdd.n2927 gnd 0.009061f
C4845 vdd.n2929 gnd 0.009061f
C4846 vdd.n2930 gnd 0.009061f
C4847 vdd.n2931 gnd 0.007293f
C4848 vdd.n2932 gnd 0.007293f
C4849 vdd.n2933 gnd 0.007293f
C4850 vdd.n2934 gnd 0.009061f
C4851 vdd.n2936 gnd 0.009061f
C4852 vdd.n2937 gnd 0.009061f
C4853 vdd.n2938 gnd 0.007293f
C4854 vdd.n2939 gnd 0.007293f
C4855 vdd.n2940 gnd 0.007293f
C4856 vdd.n2941 gnd 0.009061f
C4857 vdd.n2943 gnd 0.009061f
C4858 vdd.n2944 gnd 0.009061f
C4859 vdd.n2945 gnd 0.007293f
C4860 vdd.n2946 gnd 0.009061f
C4861 vdd.n2947 gnd 0.009061f
C4862 vdd.n2948 gnd 0.009061f
C4863 vdd.n2949 gnd 0.015608f
C4864 vdd.n2950 gnd 0.004959f
C4865 vdd.n2951 gnd 0.007293f
C4866 vdd.n2952 gnd 0.009061f
C4867 vdd.n2954 gnd 0.009061f
C4868 vdd.n2955 gnd 0.009061f
C4869 vdd.n2956 gnd 0.007293f
C4870 vdd.n2957 gnd 0.007293f
C4871 vdd.n2958 gnd 0.007293f
C4872 vdd.n2959 gnd 0.009061f
C4873 vdd.n2961 gnd 0.009061f
C4874 vdd.n2962 gnd 0.009061f
C4875 vdd.n2963 gnd 0.007293f
C4876 vdd.n2964 gnd 0.007293f
C4877 vdd.n2965 gnd 0.007293f
C4878 vdd.n2966 gnd 0.009061f
C4879 vdd.n2968 gnd 0.009061f
C4880 vdd.n2969 gnd 0.009061f
C4881 vdd.n2970 gnd 0.007293f
C4882 vdd.n2971 gnd 0.007293f
C4883 vdd.n2972 gnd 0.007293f
C4884 vdd.n2973 gnd 0.009061f
C4885 vdd.n2975 gnd 0.009061f
C4886 vdd.n2976 gnd 0.009061f
C4887 vdd.n2977 gnd 0.007293f
C4888 vdd.n2978 gnd 0.007293f
C4889 vdd.n2979 gnd 0.007293f
C4890 vdd.n2980 gnd 0.009061f
C4891 vdd.n2982 gnd 0.009061f
C4892 vdd.n2983 gnd 0.009061f
C4893 vdd.n2984 gnd 0.007293f
C4894 vdd.n2985 gnd 0.009061f
C4895 vdd.n2986 gnd 0.009061f
C4896 vdd.n2987 gnd 0.009061f
C4897 vdd.n2988 gnd 0.015608f
C4898 vdd.n2989 gnd 0.00609f
C4899 vdd.n2990 gnd 0.007293f
C4900 vdd.n2991 gnd 0.009061f
C4901 vdd.n2993 gnd 0.009061f
C4902 vdd.n2994 gnd 0.009061f
C4903 vdd.n2995 gnd 0.007293f
C4904 vdd.n2996 gnd 0.007293f
C4905 vdd.n2997 gnd 0.007293f
C4906 vdd.n2998 gnd 0.009061f
C4907 vdd.n3000 gnd 0.009061f
C4908 vdd.n3001 gnd 0.009061f
C4909 vdd.n3002 gnd 0.007293f
C4910 vdd.n3003 gnd 0.007293f
C4911 vdd.n3004 gnd 0.007293f
C4912 vdd.n3005 gnd 0.009061f
C4913 vdd.n3007 gnd 0.009061f
C4914 vdd.n3008 gnd 0.009061f
C4915 vdd.n3009 gnd 0.007293f
C4916 vdd.n3010 gnd 0.007293f
C4917 vdd.n3011 gnd 0.007293f
C4918 vdd.n3012 gnd 0.009061f
C4919 vdd.n3014 gnd 0.009061f
C4920 vdd.n3015 gnd 0.009061f
C4921 vdd.n3017 gnd 0.009061f
C4922 vdd.n3018 gnd 0.007293f
C4923 vdd.n3019 gnd 0.007293f
C4924 vdd.n3020 gnd 0.006053f
C4925 vdd.n3021 gnd 0.022589f
C4926 vdd.n3022 gnd 0.022083f
C4927 vdd.n3023 gnd 0.006053f
C4928 vdd.n3024 gnd 0.022083f
C4929 vdd.n3025 gnd 1.36588f
C4930 vdd.t55 gnd 0.463009f
C4931 vdd.n3026 gnd 0.48616f
C4932 vdd.n3027 gnd 0.926018f
C4933 vdd.n3028 gnd 0.009061f
C4934 vdd.n3029 gnd 0.007293f
C4935 vdd.n3030 gnd 0.007293f
C4936 vdd.n3031 gnd 0.007293f
C4937 vdd.n3032 gnd 0.009061f
C4938 vdd.n3033 gnd 0.828786f
C4939 vdd.t139 gnd 0.463009f
C4940 vdd.n3034 gnd 0.560241f
C4941 vdd.n3035 gnd 0.671363f
C4942 vdd.n3036 gnd 0.009061f
C4943 vdd.n3037 gnd 0.007293f
C4944 vdd.n3038 gnd 0.007293f
C4945 vdd.n3039 gnd 0.007293f
C4946 vdd.n3040 gnd 0.009061f
C4947 vdd.n3041 gnd 0.51394f
C4948 vdd.t161 gnd 0.463009f
C4949 vdd.n3042 gnd 0.768595f
C4950 vdd.t137 gnd 0.463009f
C4951 vdd.n3043 gnd 0.569501f
C4952 vdd.n3044 gnd 0.009061f
C4953 vdd.n3045 gnd 0.007293f
C4954 vdd.n3046 gnd 0.006964f
C4955 vdd.n3047 gnd 0.534468f
C4956 vdd.n3048 gnd 1.83522f
C4957 CSoutput.n0 gnd 0.036693f
C4958 CSoutput.t142 gnd 0.242719f
C4959 CSoutput.n1 gnd 0.1096f
C4960 CSoutput.n2 gnd 0.036693f
C4961 CSoutput.t148 gnd 0.242719f
C4962 CSoutput.n3 gnd 0.029082f
C4963 CSoutput.n4 gnd 0.036693f
C4964 CSoutput.t134 gnd 0.242719f
C4965 CSoutput.n5 gnd 0.025078f
C4966 CSoutput.n6 gnd 0.036693f
C4967 CSoutput.t146 gnd 0.242719f
C4968 CSoutput.t143 gnd 0.242719f
C4969 CSoutput.n7 gnd 0.108405f
C4970 CSoutput.n8 gnd 0.036693f
C4971 CSoutput.t132 gnd 0.242719f
C4972 CSoutput.n9 gnd 0.023911f
C4973 CSoutput.n10 gnd 0.036693f
C4974 CSoutput.t136 gnd 0.242719f
C4975 CSoutput.t140 gnd 0.242719f
C4976 CSoutput.n11 gnd 0.108405f
C4977 CSoutput.n12 gnd 0.036693f
C4978 CSoutput.t129 gnd 0.242719f
C4979 CSoutput.n13 gnd 0.025078f
C4980 CSoutput.n14 gnd 0.036693f
C4981 CSoutput.t128 gnd 0.242719f
C4982 CSoutput.t139 gnd 0.242719f
C4983 CSoutput.n15 gnd 0.108405f
C4984 CSoutput.n16 gnd 0.036693f
C4985 CSoutput.t144 gnd 0.242719f
C4986 CSoutput.n17 gnd 0.026785f
C4987 CSoutput.t130 gnd 0.290056f
C4988 CSoutput.t149 gnd 0.242719f
C4989 CSoutput.n18 gnd 0.138391f
C4990 CSoutput.n19 gnd 0.134288f
C4991 CSoutput.n20 gnd 0.15579f
C4992 CSoutput.n21 gnd 0.036693f
C4993 CSoutput.n22 gnd 0.030625f
C4994 CSoutput.n23 gnd 0.108405f
C4995 CSoutput.n24 gnd 0.029521f
C4996 CSoutput.n25 gnd 0.029082f
C4997 CSoutput.n26 gnd 0.036693f
C4998 CSoutput.n27 gnd 0.036693f
C4999 CSoutput.n28 gnd 0.030389f
C5000 CSoutput.n29 gnd 0.025801f
C5001 CSoutput.n30 gnd 0.110819f
C5002 CSoutput.n31 gnd 0.026157f
C5003 CSoutput.n32 gnd 0.036693f
C5004 CSoutput.n33 gnd 0.036693f
C5005 CSoutput.n34 gnd 0.036693f
C5006 CSoutput.n35 gnd 0.030066f
C5007 CSoutput.n36 gnd 0.108405f
C5008 CSoutput.n37 gnd 0.028753f
C5009 CSoutput.n38 gnd 0.02985f
C5010 CSoutput.n39 gnd 0.036693f
C5011 CSoutput.n40 gnd 0.036693f
C5012 CSoutput.n41 gnd 0.030618f
C5013 CSoutput.n42 gnd 0.027985f
C5014 CSoutput.n43 gnd 0.108405f
C5015 CSoutput.n44 gnd 0.028695f
C5016 CSoutput.n45 gnd 0.036693f
C5017 CSoutput.n46 gnd 0.036693f
C5018 CSoutput.n47 gnd 0.036693f
C5019 CSoutput.n48 gnd 0.028695f
C5020 CSoutput.n49 gnd 0.108405f
C5021 CSoutput.n50 gnd 0.027985f
C5022 CSoutput.n51 gnd 0.030618f
C5023 CSoutput.n52 gnd 0.036693f
C5024 CSoutput.n53 gnd 0.036693f
C5025 CSoutput.n54 gnd 0.02985f
C5026 CSoutput.n55 gnd 0.028753f
C5027 CSoutput.n56 gnd 0.108405f
C5028 CSoutput.n57 gnd 0.030066f
C5029 CSoutput.n58 gnd 0.036693f
C5030 CSoutput.n59 gnd 0.036693f
C5031 CSoutput.n60 gnd 0.036693f
C5032 CSoutput.n61 gnd 0.026157f
C5033 CSoutput.n62 gnd 0.110819f
C5034 CSoutput.n63 gnd 0.025801f
C5035 CSoutput.t147 gnd 0.242719f
C5036 CSoutput.n64 gnd 0.108405f
C5037 CSoutput.n65 gnd 0.030389f
C5038 CSoutput.n66 gnd 0.036693f
C5039 CSoutput.n67 gnd 0.036693f
C5040 CSoutput.n68 gnd 0.036693f
C5041 CSoutput.n69 gnd 0.029521f
C5042 CSoutput.n70 gnd 0.108405f
C5043 CSoutput.n71 gnd 0.030625f
C5044 CSoutput.n72 gnd 0.026785f
C5045 CSoutput.n73 gnd 0.036693f
C5046 CSoutput.n74 gnd 0.036693f
C5047 CSoutput.n75 gnd 0.027778f
C5048 CSoutput.n76 gnd 0.016497f
C5049 CSoutput.t131 gnd 0.272712f
C5050 CSoutput.n77 gnd 0.135473f
C5051 CSoutput.n78 gnd 0.579675f
C5052 CSoutput.t85 gnd 0.04577f
C5053 CSoutput.t72 gnd 0.04577f
C5054 CSoutput.n79 gnd 0.354366f
C5055 CSoutput.t74 gnd 0.04577f
C5056 CSoutput.t82 gnd 0.04577f
C5057 CSoutput.n80 gnd 0.353734f
C5058 CSoutput.n81 gnd 0.359039f
C5059 CSoutput.t94 gnd 0.04577f
C5060 CSoutput.t105 gnd 0.04577f
C5061 CSoutput.n82 gnd 0.353734f
C5062 CSoutput.n83 gnd 0.17692f
C5063 CSoutput.t66 gnd 0.04577f
C5064 CSoutput.t71 gnd 0.04577f
C5065 CSoutput.n84 gnd 0.353734f
C5066 CSoutput.n85 gnd 0.32443f
C5067 CSoutput.t83 gnd 0.04577f
C5068 CSoutput.t95 gnd 0.04577f
C5069 CSoutput.n86 gnd 0.354366f
C5070 CSoutput.t98 gnd 0.04577f
C5071 CSoutput.t106 gnd 0.04577f
C5072 CSoutput.n87 gnd 0.353734f
C5073 CSoutput.n88 gnd 0.359039f
C5074 CSoutput.t110 gnd 0.04577f
C5075 CSoutput.t93 gnd 0.04577f
C5076 CSoutput.n89 gnd 0.353734f
C5077 CSoutput.n90 gnd 0.17692f
C5078 CSoutput.t97 gnd 0.04577f
C5079 CSoutput.t80 gnd 0.04577f
C5080 CSoutput.n91 gnd 0.353734f
C5081 CSoutput.n92 gnd 0.263831f
C5082 CSoutput.n93 gnd 0.33269f
C5083 CSoutput.t64 gnd 0.04577f
C5084 CSoutput.t65 gnd 0.04577f
C5085 CSoutput.n94 gnd 0.354366f
C5086 CSoutput.t76 gnd 0.04577f
C5087 CSoutput.t104 gnd 0.04577f
C5088 CSoutput.n95 gnd 0.353734f
C5089 CSoutput.n96 gnd 0.359039f
C5090 CSoutput.t108 gnd 0.04577f
C5091 CSoutput.t86 gnd 0.04577f
C5092 CSoutput.n97 gnd 0.353734f
C5093 CSoutput.n98 gnd 0.17692f
C5094 CSoutput.t75 gnd 0.04577f
C5095 CSoutput.t87 gnd 0.04577f
C5096 CSoutput.n99 gnd 0.353734f
C5097 CSoutput.n100 gnd 0.263831f
C5098 CSoutput.n101 gnd 0.371862f
C5099 CSoutput.n102 gnd 7.5385f
C5100 CSoutput.n104 gnd 0.649101f
C5101 CSoutput.n105 gnd 0.486825f
C5102 CSoutput.n106 gnd 0.649101f
C5103 CSoutput.n107 gnd 0.649101f
C5104 CSoutput.n108 gnd 1.74758f
C5105 CSoutput.n109 gnd 0.649101f
C5106 CSoutput.n110 gnd 0.649101f
C5107 CSoutput.t138 gnd 0.811376f
C5108 CSoutput.n111 gnd 0.649101f
C5109 CSoutput.n112 gnd 0.649101f
C5110 CSoutput.n116 gnd 0.649101f
C5111 CSoutput.n120 gnd 0.649101f
C5112 CSoutput.n121 gnd 0.649101f
C5113 CSoutput.n123 gnd 0.649101f
C5114 CSoutput.n128 gnd 0.649101f
C5115 CSoutput.n130 gnd 0.649101f
C5116 CSoutput.n131 gnd 0.649101f
C5117 CSoutput.n133 gnd 0.649101f
C5118 CSoutput.n134 gnd 0.649101f
C5119 CSoutput.n136 gnd 0.649101f
C5120 CSoutput.t133 gnd 10.8464f
C5121 CSoutput.n138 gnd 0.649101f
C5122 CSoutput.n139 gnd 0.486825f
C5123 CSoutput.n140 gnd 0.649101f
C5124 CSoutput.n141 gnd 0.649101f
C5125 CSoutput.n142 gnd 1.74758f
C5126 CSoutput.n143 gnd 0.649101f
C5127 CSoutput.n144 gnd 0.649101f
C5128 CSoutput.t135 gnd 0.811376f
C5129 CSoutput.n145 gnd 0.649101f
C5130 CSoutput.n146 gnd 0.649101f
C5131 CSoutput.n150 gnd 0.649101f
C5132 CSoutput.n154 gnd 0.649101f
C5133 CSoutput.n155 gnd 0.649101f
C5134 CSoutput.n157 gnd 0.649101f
C5135 CSoutput.n162 gnd 0.649101f
C5136 CSoutput.n164 gnd 0.649101f
C5137 CSoutput.n165 gnd 0.649101f
C5138 CSoutput.n167 gnd 0.649101f
C5139 CSoutput.n168 gnd 0.649101f
C5140 CSoutput.n170 gnd 0.649101f
C5141 CSoutput.n171 gnd 0.486825f
C5142 CSoutput.n173 gnd 0.649101f
C5143 CSoutput.n174 gnd 0.486825f
C5144 CSoutput.n175 gnd 0.649101f
C5145 CSoutput.n176 gnd 0.649101f
C5146 CSoutput.n177 gnd 1.74758f
C5147 CSoutput.n178 gnd 0.649101f
C5148 CSoutput.n179 gnd 0.649101f
C5149 CSoutput.t137 gnd 0.811376f
C5150 CSoutput.n180 gnd 0.649101f
C5151 CSoutput.n181 gnd 1.74758f
C5152 CSoutput.n183 gnd 0.649101f
C5153 CSoutput.n184 gnd 0.649101f
C5154 CSoutput.n186 gnd 0.649101f
C5155 CSoutput.n187 gnd 0.649101f
C5156 CSoutput.t145 gnd 10.6696f
C5157 CSoutput.t141 gnd 10.8464f
C5158 CSoutput.n193 gnd 2.03632f
C5159 CSoutput.n194 gnd 8.29524f
C5160 CSoutput.n195 gnd 8.64235f
C5161 CSoutput.n200 gnd 2.20589f
C5162 CSoutput.n206 gnd 0.649101f
C5163 CSoutput.n208 gnd 0.649101f
C5164 CSoutput.n210 gnd 0.649101f
C5165 CSoutput.n212 gnd 0.649101f
C5166 CSoutput.n214 gnd 0.649101f
C5167 CSoutput.n220 gnd 0.649101f
C5168 CSoutput.n227 gnd 1.19085f
C5169 CSoutput.n228 gnd 1.19085f
C5170 CSoutput.n229 gnd 0.649101f
C5171 CSoutput.n230 gnd 0.649101f
C5172 CSoutput.n232 gnd 0.486825f
C5173 CSoutput.n233 gnd 0.416922f
C5174 CSoutput.n235 gnd 0.486825f
C5175 CSoutput.n236 gnd 0.416922f
C5176 CSoutput.n237 gnd 0.486825f
C5177 CSoutput.n239 gnd 0.649101f
C5178 CSoutput.n241 gnd 1.74758f
C5179 CSoutput.n242 gnd 2.03632f
C5180 CSoutput.n243 gnd 7.62949f
C5181 CSoutput.n245 gnd 0.486825f
C5182 CSoutput.n246 gnd 1.25263f
C5183 CSoutput.n247 gnd 0.486825f
C5184 CSoutput.n249 gnd 0.649101f
C5185 CSoutput.n251 gnd 1.74758f
C5186 CSoutput.n252 gnd 3.80651f
C5187 CSoutput.t109 gnd 0.04577f
C5188 CSoutput.t84 gnd 0.04577f
C5189 CSoutput.n253 gnd 0.354366f
C5190 CSoutput.t100 gnd 0.04577f
C5191 CSoutput.t68 gnd 0.04577f
C5192 CSoutput.n254 gnd 0.353734f
C5193 CSoutput.n255 gnd 0.359039f
C5194 CSoutput.t69 gnd 0.04577f
C5195 CSoutput.t92 gnd 0.04577f
C5196 CSoutput.n256 gnd 0.353734f
C5197 CSoutput.n257 gnd 0.17692f
C5198 CSoutput.t78 gnd 0.04577f
C5199 CSoutput.t67 gnd 0.04577f
C5200 CSoutput.n258 gnd 0.353734f
C5201 CSoutput.n259 gnd 0.32443f
C5202 CSoutput.t101 gnd 0.04577f
C5203 CSoutput.t102 gnd 0.04577f
C5204 CSoutput.n260 gnd 0.354366f
C5205 CSoutput.t73 gnd 0.04577f
C5206 CSoutput.t111 gnd 0.04577f
C5207 CSoutput.n261 gnd 0.353734f
C5208 CSoutput.n262 gnd 0.359039f
C5209 CSoutput.t81 gnd 0.04577f
C5210 CSoutput.t99 gnd 0.04577f
C5211 CSoutput.n263 gnd 0.353734f
C5212 CSoutput.n264 gnd 0.17692f
C5213 CSoutput.t91 gnd 0.04577f
C5214 CSoutput.t70 gnd 0.04577f
C5215 CSoutput.n265 gnd 0.353734f
C5216 CSoutput.n266 gnd 0.263831f
C5217 CSoutput.n267 gnd 0.33269f
C5218 CSoutput.t89 gnd 0.04577f
C5219 CSoutput.t90 gnd 0.04577f
C5220 CSoutput.n268 gnd 0.354366f
C5221 CSoutput.t96 gnd 0.04577f
C5222 CSoutput.t103 gnd 0.04577f
C5223 CSoutput.n269 gnd 0.353734f
C5224 CSoutput.n270 gnd 0.359039f
C5225 CSoutput.t88 gnd 0.04577f
C5226 CSoutput.t77 gnd 0.04577f
C5227 CSoutput.n271 gnd 0.353734f
C5228 CSoutput.n272 gnd 0.17692f
C5229 CSoutput.t107 gnd 0.04577f
C5230 CSoutput.t79 gnd 0.04577f
C5231 CSoutput.n273 gnd 0.353733f
C5232 CSoutput.n274 gnd 0.263833f
C5233 CSoutput.n275 gnd 0.371862f
C5234 CSoutput.n276 gnd 10.4353f
C5235 CSoutput.t121 gnd 0.040049f
C5236 CSoutput.t59 gnd 0.040049f
C5237 CSoutput.n277 gnd 0.355068f
C5238 CSoutput.t3 gnd 0.040049f
C5239 CSoutput.t53 gnd 0.040049f
C5240 CSoutput.n278 gnd 0.353884f
C5241 CSoutput.n279 gnd 0.329754f
C5242 CSoutput.t17 gnd 0.040049f
C5243 CSoutput.t25 gnd 0.040049f
C5244 CSoutput.n280 gnd 0.353884f
C5245 CSoutput.n281 gnd 0.162553f
C5246 CSoutput.t51 gnd 0.040049f
C5247 CSoutput.t8 gnd 0.040049f
C5248 CSoutput.n282 gnd 0.353884f
C5249 CSoutput.n283 gnd 0.162553f
C5250 CSoutput.t61 gnd 0.040049f
C5251 CSoutput.t22 gnd 0.040049f
C5252 CSoutput.n284 gnd 0.353884f
C5253 CSoutput.n285 gnd 0.162553f
C5254 CSoutput.t62 gnd 0.040049f
C5255 CSoutput.t113 gnd 0.040049f
C5256 CSoutput.n286 gnd 0.353884f
C5257 CSoutput.n287 gnd 0.162553f
C5258 CSoutput.t112 gnd 0.040049f
C5259 CSoutput.t50 gnd 0.040049f
C5260 CSoutput.n288 gnd 0.353884f
C5261 CSoutput.n289 gnd 0.162553f
C5262 CSoutput.t32 gnd 0.040049f
C5263 CSoutput.t38 gnd 0.040049f
C5264 CSoutput.n290 gnd 0.353884f
C5265 CSoutput.n291 gnd 0.162553f
C5266 CSoutput.t16 gnd 0.040049f
C5267 CSoutput.t4 gnd 0.040049f
C5268 CSoutput.n292 gnd 0.353884f
C5269 CSoutput.n293 gnd 0.162553f
C5270 CSoutput.t27 gnd 0.040049f
C5271 CSoutput.t116 gnd 0.040049f
C5272 CSoutput.n294 gnd 0.353884f
C5273 CSoutput.n295 gnd 0.299781f
C5274 CSoutput.t40 gnd 0.040049f
C5275 CSoutput.t117 gnd 0.040049f
C5276 CSoutput.n296 gnd 0.355068f
C5277 CSoutput.t123 gnd 0.040049f
C5278 CSoutput.t43 gnd 0.040049f
C5279 CSoutput.n297 gnd 0.353884f
C5280 CSoutput.n298 gnd 0.329754f
C5281 CSoutput.t37 gnd 0.040049f
C5282 CSoutput.t20 gnd 0.040049f
C5283 CSoutput.n299 gnd 0.353884f
C5284 CSoutput.n300 gnd 0.162553f
C5285 CSoutput.t1 gnd 0.040049f
C5286 CSoutput.t58 gnd 0.040049f
C5287 CSoutput.n301 gnd 0.353884f
C5288 CSoutput.n302 gnd 0.162553f
C5289 CSoutput.t119 gnd 0.040049f
C5290 CSoutput.t127 gnd 0.040049f
C5291 CSoutput.n303 gnd 0.353884f
C5292 CSoutput.n304 gnd 0.162553f
C5293 CSoutput.t23 gnd 0.040049f
C5294 CSoutput.t36 gnd 0.040049f
C5295 CSoutput.n305 gnd 0.353884f
C5296 CSoutput.n306 gnd 0.162553f
C5297 CSoutput.t55 gnd 0.040049f
C5298 CSoutput.t115 gnd 0.040049f
C5299 CSoutput.n307 gnd 0.353884f
C5300 CSoutput.n308 gnd 0.162553f
C5301 CSoutput.t9 gnd 0.040049f
C5302 CSoutput.t125 gnd 0.040049f
C5303 CSoutput.n309 gnd 0.353884f
C5304 CSoutput.n310 gnd 0.162553f
C5305 CSoutput.t34 gnd 0.040049f
C5306 CSoutput.t19 gnd 0.040049f
C5307 CSoutput.n311 gnd 0.353884f
C5308 CSoutput.n312 gnd 0.162553f
C5309 CSoutput.t2 gnd 0.040049f
C5310 CSoutput.t41 gnd 0.040049f
C5311 CSoutput.n313 gnd 0.353884f
C5312 CSoutput.n314 gnd 0.24679f
C5313 CSoutput.n315 gnd 0.458555f
C5314 CSoutput.n316 gnd 11.6175f
C5315 CSoutput.t122 gnd 0.040049f
C5316 CSoutput.t45 gnd 0.040049f
C5317 CSoutput.n317 gnd 0.355068f
C5318 CSoutput.t15 gnd 0.040049f
C5319 CSoutput.t10 gnd 0.040049f
C5320 CSoutput.n318 gnd 0.353884f
C5321 CSoutput.n319 gnd 0.329754f
C5322 CSoutput.t5 gnd 0.040049f
C5323 CSoutput.t24 gnd 0.040049f
C5324 CSoutput.n320 gnd 0.353884f
C5325 CSoutput.n321 gnd 0.162553f
C5326 CSoutput.t120 gnd 0.040049f
C5327 CSoutput.t63 gnd 0.040049f
C5328 CSoutput.n322 gnd 0.353884f
C5329 CSoutput.n323 gnd 0.162553f
C5330 CSoutput.t11 gnd 0.040049f
C5331 CSoutput.t126 gnd 0.040049f
C5332 CSoutput.n324 gnd 0.353884f
C5333 CSoutput.n325 gnd 0.162553f
C5334 CSoutput.t7 gnd 0.040049f
C5335 CSoutput.t57 gnd 0.040049f
C5336 CSoutput.n326 gnd 0.353884f
C5337 CSoutput.n327 gnd 0.162553f
C5338 CSoutput.t28 gnd 0.040049f
C5339 CSoutput.t30 gnd 0.040049f
C5340 CSoutput.n328 gnd 0.353884f
C5341 CSoutput.n329 gnd 0.162553f
C5342 CSoutput.t33 gnd 0.040049f
C5343 CSoutput.t54 gnd 0.040049f
C5344 CSoutput.n330 gnd 0.353884f
C5345 CSoutput.n331 gnd 0.162553f
C5346 CSoutput.t12 gnd 0.040049f
C5347 CSoutput.t44 gnd 0.040049f
C5348 CSoutput.n332 gnd 0.353884f
C5349 CSoutput.n333 gnd 0.162553f
C5350 CSoutput.t46 gnd 0.040049f
C5351 CSoutput.t56 gnd 0.040049f
C5352 CSoutput.n334 gnd 0.353884f
C5353 CSoutput.n335 gnd 0.299781f
C5354 CSoutput.t31 gnd 0.040049f
C5355 CSoutput.t114 gnd 0.040049f
C5356 CSoutput.n336 gnd 0.355068f
C5357 CSoutput.t35 gnd 0.040049f
C5358 CSoutput.t49 gnd 0.040049f
C5359 CSoutput.n337 gnd 0.353884f
C5360 CSoutput.n338 gnd 0.329754f
C5361 CSoutput.t18 gnd 0.040049f
C5362 CSoutput.t47 gnd 0.040049f
C5363 CSoutput.n339 gnd 0.353884f
C5364 CSoutput.n340 gnd 0.162553f
C5365 CSoutput.t52 gnd 0.040049f
C5366 CSoutput.t6 gnd 0.040049f
C5367 CSoutput.n341 gnd 0.353884f
C5368 CSoutput.n342 gnd 0.162553f
C5369 CSoutput.t29 gnd 0.040049f
C5370 CSoutput.t14 gnd 0.040049f
C5371 CSoutput.n343 gnd 0.353884f
C5372 CSoutput.n344 gnd 0.162553f
C5373 CSoutput.t48 gnd 0.040049f
C5374 CSoutput.t0 gnd 0.040049f
C5375 CSoutput.n345 gnd 0.353884f
C5376 CSoutput.n346 gnd 0.162553f
C5377 CSoutput.t13 gnd 0.040049f
C5378 CSoutput.t21 gnd 0.040049f
C5379 CSoutput.n347 gnd 0.353884f
C5380 CSoutput.n348 gnd 0.162553f
C5381 CSoutput.t26 gnd 0.040049f
C5382 CSoutput.t124 gnd 0.040049f
C5383 CSoutput.n349 gnd 0.353884f
C5384 CSoutput.n350 gnd 0.162553f
C5385 CSoutput.t60 gnd 0.040049f
C5386 CSoutput.t118 gnd 0.040049f
C5387 CSoutput.n351 gnd 0.353884f
C5388 CSoutput.n352 gnd 0.162553f
C5389 CSoutput.t39 gnd 0.040049f
C5390 CSoutput.t42 gnd 0.040049f
C5391 CSoutput.n353 gnd 0.353884f
C5392 CSoutput.n354 gnd 0.24679f
C5393 CSoutput.n355 gnd 0.458555f
C5394 CSoutput.n356 gnd 6.92896f
C5395 CSoutput.n357 gnd 12.168099f
C5396 a_n5644_8799.n0 gnd 0.207688f
C5397 a_n5644_8799.n1 gnd 0.286319f
C5398 a_n5644_8799.n2 gnd 0.217233f
C5399 a_n5644_8799.n3 gnd 0.207688f
C5400 a_n5644_8799.n4 gnd 0.286319f
C5401 a_n5644_8799.n5 gnd 0.217233f
C5402 a_n5644_8799.n6 gnd 0.207688f
C5403 a_n5644_8799.n7 gnd 0.451214f
C5404 a_n5644_8799.n8 gnd 0.217233f
C5405 a_n5644_8799.n9 gnd 0.207688f
C5406 a_n5644_8799.n10 gnd 0.321077f
C5407 a_n5644_8799.n11 gnd 0.182475f
C5408 a_n5644_8799.n12 gnd 0.207688f
C5409 a_n5644_8799.n13 gnd 0.321077f
C5410 a_n5644_8799.n14 gnd 0.182475f
C5411 a_n5644_8799.n15 gnd 0.207688f
C5412 a_n5644_8799.n16 gnd 0.321077f
C5413 a_n5644_8799.n17 gnd 0.34737f
C5414 a_n5644_8799.n18 gnd 4.02716f
C5415 a_n5644_8799.n19 gnd 2.78963f
C5416 a_n5644_8799.n20 gnd 0.363059f
C5417 a_n5644_8799.n21 gnd 3.04277f
C5418 a_n5644_8799.n22 gnd 0.363058f
C5419 a_n5644_8799.n23 gnd 0.855698f
C5420 a_n5644_8799.n24 gnd 0.250037f
C5421 a_n5644_8799.n25 gnd 0.004668f
C5422 a_n5644_8799.n26 gnd 0.010096f
C5423 a_n5644_8799.n27 gnd 0.010096f
C5424 a_n5644_8799.n28 gnd 0.004668f
C5425 a_n5644_8799.n29 gnd 0.250037f
C5426 a_n5644_8799.n30 gnd 0.004668f
C5427 a_n5644_8799.n31 gnd 0.010096f
C5428 a_n5644_8799.n32 gnd 0.010096f
C5429 a_n5644_8799.n33 gnd 0.004668f
C5430 a_n5644_8799.n34 gnd 0.250037f
C5431 a_n5644_8799.n35 gnd 0.004668f
C5432 a_n5644_8799.n36 gnd 0.010096f
C5433 a_n5644_8799.n37 gnd 0.010096f
C5434 a_n5644_8799.n38 gnd 0.004668f
C5435 a_n5644_8799.n39 gnd 0.004668f
C5436 a_n5644_8799.n40 gnd 0.010096f
C5437 a_n5644_8799.n41 gnd 0.010096f
C5438 a_n5644_8799.n42 gnd 0.004668f
C5439 a_n5644_8799.n43 gnd 0.250037f
C5440 a_n5644_8799.n44 gnd 0.004668f
C5441 a_n5644_8799.n45 gnd 0.010096f
C5442 a_n5644_8799.n46 gnd 0.010096f
C5443 a_n5644_8799.n47 gnd 0.004668f
C5444 a_n5644_8799.n48 gnd 0.250037f
C5445 a_n5644_8799.n49 gnd 0.004668f
C5446 a_n5644_8799.n50 gnd 0.010096f
C5447 a_n5644_8799.n51 gnd 0.010096f
C5448 a_n5644_8799.n52 gnd 0.004668f
C5449 a_n5644_8799.n53 gnd 0.250037f
C5450 a_n5644_8799.t27 gnd 0.144055f
C5451 a_n5644_8799.t32 gnd 0.144055f
C5452 a_n5644_8799.t23 gnd 0.144055f
C5453 a_n5644_8799.n54 gnd 1.13618f
C5454 a_n5644_8799.t22 gnd 0.144055f
C5455 a_n5644_8799.t31 gnd 0.144055f
C5456 a_n5644_8799.n55 gnd 1.13431f
C5457 a_n5644_8799.t34 gnd 0.144055f
C5458 a_n5644_8799.t35 gnd 0.144055f
C5459 a_n5644_8799.n56 gnd 1.13431f
C5460 a_n5644_8799.t16 gnd 0.112043f
C5461 a_n5644_8799.t19 gnd 0.112043f
C5462 a_n5644_8799.n57 gnd 0.992966f
C5463 a_n5644_8799.t3 gnd 0.112043f
C5464 a_n5644_8799.t24 gnd 0.112043f
C5465 a_n5644_8799.n58 gnd 0.990047f
C5466 a_n5644_8799.n59 gnd 0.877922f
C5467 a_n5644_8799.t4 gnd 0.112043f
C5468 a_n5644_8799.t2 gnd 0.112043f
C5469 a_n5644_8799.n60 gnd 0.990047f
C5470 a_n5644_8799.t25 gnd 0.112043f
C5471 a_n5644_8799.t15 gnd 0.112043f
C5472 a_n5644_8799.n61 gnd 0.992966f
C5473 a_n5644_8799.t6 gnd 0.112043f
C5474 a_n5644_8799.t21 gnd 0.112043f
C5475 a_n5644_8799.n62 gnd 0.990046f
C5476 a_n5644_8799.n63 gnd 0.877924f
C5477 a_n5644_8799.t14 gnd 0.112043f
C5478 a_n5644_8799.t5 gnd 0.112043f
C5479 a_n5644_8799.n64 gnd 0.990046f
C5480 a_n5644_8799.t13 gnd 0.112043f
C5481 a_n5644_8799.t1 gnd 0.112043f
C5482 a_n5644_8799.n65 gnd 0.992966f
C5483 a_n5644_8799.t8 gnd 0.112043f
C5484 a_n5644_8799.t9 gnd 0.112043f
C5485 a_n5644_8799.n66 gnd 0.990046f
C5486 a_n5644_8799.n67 gnd 0.877924f
C5487 a_n5644_8799.t11 gnd 0.112043f
C5488 a_n5644_8799.t17 gnd 0.112043f
C5489 a_n5644_8799.n68 gnd 0.990046f
C5490 a_n5644_8799.t18 gnd 0.112043f
C5491 a_n5644_8799.t7 gnd 0.112043f
C5492 a_n5644_8799.n69 gnd 0.990047f
C5493 a_n5644_8799.n70 gnd 3.08844f
C5494 a_n5644_8799.t26 gnd 0.112043f
C5495 a_n5644_8799.t20 gnd 0.112043f
C5496 a_n5644_8799.n71 gnd 0.990047f
C5497 a_n5644_8799.n72 gnd 0.432262f
C5498 a_n5644_8799.t29 gnd 0.112043f
C5499 a_n5644_8799.t0 gnd 0.112043f
C5500 a_n5644_8799.n73 gnd 0.990047f
C5501 a_n5644_8799.t75 gnd 0.597318f
C5502 a_n5644_8799.n74 gnd 0.26846f
C5503 a_n5644_8799.t42 gnd 0.597318f
C5504 a_n5644_8799.t62 gnd 0.597318f
C5505 a_n5644_8799.t53 gnd 0.608623f
C5506 a_n5644_8799.n75 gnd 0.250405f
C5507 a_n5644_8799.n76 gnd 0.270847f
C5508 a_n5644_8799.t77 gnd 0.597318f
C5509 a_n5644_8799.n77 gnd 0.26846f
C5510 a_n5644_8799.n78 gnd 0.264052f
C5511 a_n5644_8799.t52 gnd 0.597318f
C5512 a_n5644_8799.n79 gnd 0.264052f
C5513 a_n5644_8799.t41 gnd 0.597318f
C5514 a_n5644_8799.n80 gnd 0.270847f
C5515 a_n5644_8799.t40 gnd 0.608613f
C5516 a_n5644_8799.t79 gnd 0.597318f
C5517 a_n5644_8799.n81 gnd 0.26846f
C5518 a_n5644_8799.t49 gnd 0.597318f
C5519 a_n5644_8799.t68 gnd 0.597318f
C5520 a_n5644_8799.t58 gnd 0.608623f
C5521 a_n5644_8799.n82 gnd 0.250405f
C5522 a_n5644_8799.n83 gnd 0.270847f
C5523 a_n5644_8799.t81 gnd 0.597318f
C5524 a_n5644_8799.n84 gnd 0.26846f
C5525 a_n5644_8799.n85 gnd 0.264052f
C5526 a_n5644_8799.t57 gnd 0.597318f
C5527 a_n5644_8799.n86 gnd 0.264052f
C5528 a_n5644_8799.t45 gnd 0.597318f
C5529 a_n5644_8799.n87 gnd 0.270847f
C5530 a_n5644_8799.t47 gnd 0.608613f
C5531 a_n5644_8799.n88 gnd 0.898345f
C5532 a_n5644_8799.t66 gnd 0.597318f
C5533 a_n5644_8799.n89 gnd 0.26846f
C5534 a_n5644_8799.t74 gnd 0.597318f
C5535 a_n5644_8799.t71 gnd 0.597318f
C5536 a_n5644_8799.t39 gnd 0.608623f
C5537 a_n5644_8799.n90 gnd 0.250405f
C5538 a_n5644_8799.n91 gnd 0.270847f
C5539 a_n5644_8799.t48 gnd 0.597318f
C5540 a_n5644_8799.n92 gnd 0.26846f
C5541 a_n5644_8799.n93 gnd 0.264052f
C5542 a_n5644_8799.t54 gnd 0.597318f
C5543 a_n5644_8799.n94 gnd 0.264052f
C5544 a_n5644_8799.t43 gnd 0.597318f
C5545 a_n5644_8799.n95 gnd 0.270847f
C5546 a_n5644_8799.t83 gnd 0.608613f
C5547 a_n5644_8799.n96 gnd 1.53813f
C5548 a_n5644_8799.t60 gnd 0.608613f
C5549 a_n5644_8799.t59 gnd 0.597318f
C5550 a_n5644_8799.t46 gnd 0.597318f
C5551 a_n5644_8799.n97 gnd 0.26846f
C5552 a_n5644_8799.t76 gnd 0.597318f
C5553 a_n5644_8799.t61 gnd 0.597318f
C5554 a_n5644_8799.t51 gnd 0.597318f
C5555 a_n5644_8799.n98 gnd 0.26846f
C5556 a_n5644_8799.t69 gnd 0.608623f
C5557 a_n5644_8799.n99 gnd 0.250405f
C5558 a_n5644_8799.t78 gnd 0.597318f
C5559 a_n5644_8799.n100 gnd 0.270847f
C5560 a_n5644_8799.n101 gnd 0.264052f
C5561 a_n5644_8799.n102 gnd 0.264052f
C5562 a_n5644_8799.n103 gnd 0.270847f
C5563 a_n5644_8799.t64 gnd 0.608613f
C5564 a_n5644_8799.t63 gnd 0.597318f
C5565 a_n5644_8799.t55 gnd 0.597318f
C5566 a_n5644_8799.n104 gnd 0.26846f
C5567 a_n5644_8799.t80 gnd 0.597318f
C5568 a_n5644_8799.t67 gnd 0.597318f
C5569 a_n5644_8799.t56 gnd 0.597318f
C5570 a_n5644_8799.n105 gnd 0.26846f
C5571 a_n5644_8799.t72 gnd 0.608623f
C5572 a_n5644_8799.n106 gnd 0.250405f
C5573 a_n5644_8799.t36 gnd 0.597318f
C5574 a_n5644_8799.n107 gnd 0.270847f
C5575 a_n5644_8799.n108 gnd 0.264052f
C5576 a_n5644_8799.n109 gnd 0.264052f
C5577 a_n5644_8799.n110 gnd 0.270847f
C5578 a_n5644_8799.n111 gnd 0.898345f
C5579 a_n5644_8799.t82 gnd 0.608613f
C5580 a_n5644_8799.t44 gnd 0.597318f
C5581 a_n5644_8799.t65 gnd 0.597318f
C5582 a_n5644_8799.n112 gnd 0.26846f
C5583 a_n5644_8799.t37 gnd 0.597318f
C5584 a_n5644_8799.t73 gnd 0.597318f
C5585 a_n5644_8799.t50 gnd 0.597318f
C5586 a_n5644_8799.n113 gnd 0.26846f
C5587 a_n5644_8799.t38 gnd 0.608623f
C5588 a_n5644_8799.n114 gnd 0.250405f
C5589 a_n5644_8799.t70 gnd 0.597318f
C5590 a_n5644_8799.n115 gnd 0.270847f
C5591 a_n5644_8799.n116 gnd 0.264052f
C5592 a_n5644_8799.n117 gnd 0.264052f
C5593 a_n5644_8799.n118 gnd 0.270847f
C5594 a_n5644_8799.n119 gnd 1.08536f
C5595 a_n5644_8799.n120 gnd 12.2f
C5596 a_n5644_8799.n121 gnd 4.3715f
C5597 a_n5644_8799.n122 gnd 5.67176f
C5598 a_n5644_8799.t33 gnd 0.144055f
C5599 a_n5644_8799.t12 gnd 0.144055f
C5600 a_n5644_8799.n123 gnd 1.13431f
C5601 a_n5644_8799.t28 gnd 0.144055f
C5602 a_n5644_8799.t30 gnd 0.144055f
C5603 a_n5644_8799.n124 gnd 1.13431f
C5604 a_n5644_8799.n125 gnd 1.13618f
C5605 a_n5644_8799.t10 gnd 0.144055f
.ends

