* NGSPICE file created from opamp606.ext - technology: sky130A

.subckt opamp606 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2804_13878.t31 a_n2982_13878.t37 a_n2982_13878.t38 vdd.t265 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t163 commonsourceibias.t48 gnd.t311 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t1 a_n2982_13878.t72 vdd.t278 vdd.t277 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t296 a_n9628_8799.t48 CSoutput.t180 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t310 commonsourceibias.t49 CSoutput.t162 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 a_n9628_8799.t5 plus.t5 a_n3106_n452.t55 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X6 CSoutput.t161 commonsourceibias.t50 gnd.t309 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t160 commonsourceibias.t51 gnd.t308 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t181 a_n9628_8799.t49 vdd.t297 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 a_n3106_n452.t54 plus.t6 a_n9628_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X10 vdd.t302 a_n9628_8799.t50 CSoutput.t186 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 a_n2982_8322.t37 a_n2982_13878.t73 a_n9628_8799.t43 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 CSoutput.t187 a_n9628_8799.t51 vdd.t303 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 vdd.t80 a_n9628_8799.t52 CSoutput.t46 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 output.t16 CSoutput.t192 vdd.t4 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X15 CSoutput.t47 a_n9628_8799.t53 vdd.t81 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 gnd.t307 commonsourceibias.t52 CSoutput.t159 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X17 vdd.t5 CSoutput.t193 output.t15 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 CSoutput.t158 commonsourceibias.t53 gnd.t306 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t305 commonsourceibias.t54 CSoutput.t157 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X20 vdd.t92 a_n9628_8799.t54 CSoutput.t52 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t93 a_n9628_8799.t55 CSoutput.t53 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X22 CSoutput.t156 commonsourceibias.t55 gnd.t304 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t155 commonsourceibias.t56 gnd.t303 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t166 a_n9628_8799.t56 vdd.t282 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 a_n2982_13878.t71 minus.t5 a_n3106_n452.t31 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 CSoutput.t154 commonsourceibias.t57 gnd.t302 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n9628_8799.t15 plus.t7 a_n3106_n452.t53 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n9628_8799.t42 a_n2982_13878.t74 a_n2982_8322.t36 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 a_n2982_13878.t5 minus.t6 a_n3106_n452.t7 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X30 plus.t4 gnd.t154 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 vdd.t283 a_n9628_8799.t57 CSoutput.t167 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 vdd.t18 a_n9628_8799.t58 CSoutput.t8 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 CSoutput.t9 a_n9628_8799.t59 vdd.t19 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 a_n9628_8799.t41 a_n2982_13878.t75 a_n2982_8322.t35 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 CSoutput.t153 commonsourceibias.t58 gnd.t301 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t300 commonsourceibias.t59 CSoutput.t152 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd.t153 gnd.t151 gnd.t152 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 CSoutput.t151 commonsourceibias.t60 gnd.t299 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 CSoutput.t150 commonsourceibias.t61 gnd.t298 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n3106_n452.t52 plus.t8 a_n9628_8799.t8 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X41 vdd.t99 CSoutput.t194 output.t14 gnd.t172 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X42 CSoutput.t24 a_n9628_8799.t60 vdd.t48 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 a_n3106_n452.t2 diffpairibias.t16 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 a_n3106_n452.t23 minus.t7 a_n2982_13878.t19 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 CSoutput.t25 a_n9628_8799.t61 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 vdd.t118 a_n9628_8799.t62 CSoutput.t66 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 gnd.t297 commonsourceibias.t62 CSoutput.t149 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 vdd.t120 a_n9628_8799.t63 CSoutput.t67 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 CSoutput.t148 commonsourceibias.t63 gnd.t296 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X50 output.t17 outputibias.t8 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X51 gnd.t295 commonsourceibias.t0 commonsourceibias.t1 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t147 commonsourceibias.t64 gnd.t294 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 CSoutput.t195 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X54 vdd.t222 vdd.t220 vdd.t221 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X55 vdd.t113 a_n9628_8799.t64 CSoutput.t62 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 vdd.t100 CSoutput.t196 output.t13 gnd.t173 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X57 a_n2804_13878.t30 a_n2982_13878.t59 a_n2982_13878.t60 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 CSoutput.t146 commonsourceibias.t65 gnd.t293 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 output.t12 CSoutput.t197 vdd.t101 gnd.t174 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X60 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t29 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 vdd.t219 vdd.t217 vdd.t218 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X62 gnd.t150 gnd.t148 gnd.t149 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X63 gnd.t292 commonsourceibias.t66 CSoutput.t145 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 CSoutput.t63 a_n9628_8799.t65 vdd.t114 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 vdd.t216 vdd.t214 vdd.t215 vdd.t193 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X66 gnd.t291 commonsourceibias.t32 commonsourceibias.t33 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t144 commonsourceibias.t67 gnd.t290 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 a_n3106_n452.t51 plus.t9 a_n9628_8799.t4 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X69 vdd.t145 a_n9628_8799.t66 CSoutput.t90 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X70 vdd.t146 a_n9628_8799.t67 CSoutput.t91 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 gnd.t147 gnd.t145 gnd.t146 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X72 gnd.t144 gnd.t141 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X73 gnd.t140 gnd.t138 gnd.t139 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X74 CSoutput.t143 commonsourceibias.t68 gnd.t289 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 diffpairibias.t15 diffpairibias.t14 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 a_n3106_n452.t50 plus.t10 a_n9628_8799.t13 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X77 CSoutput.t70 a_n9628_8799.t68 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 a_n3106_n452.t29 minus.t8 a_n2982_13878.t70 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X79 a_n2982_13878.t52 a_n2982_13878.t51 a_n2804_13878.t28 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X80 CSoutput.t142 commonsourceibias.t69 gnd.t288 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X81 CSoutput.t71 a_n9628_8799.t69 vdd.t125 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t141 commonsourceibias.t70 gnd.t287 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X83 a_n9628_8799.t36 a_n2982_13878.t76 a_n2982_8322.t34 vdd.t255 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X84 gnd.t286 commonsourceibias.t71 CSoutput.t140 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 vdd.t14 a_n9628_8799.t70 CSoutput.t6 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 CSoutput.t7 a_n9628_8799.t71 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 gnd.t281 commonsourceibias.t72 CSoutput.t139 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t198 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X89 a_n2982_13878.t50 a_n2982_13878.t49 a_n2804_13878.t27 vdd.t276 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 vdd.t121 a_n9628_8799.t72 CSoutput.t68 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 vdd.t122 a_n9628_8799.t73 CSoutput.t69 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 a_n9628_8799.t35 a_n2982_13878.t77 a_n2982_8322.t33 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X93 CSoutput.t0 a_n9628_8799.t74 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 CSoutput.t138 commonsourceibias.t73 gnd.t285 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X95 diffpairibias.t13 diffpairibias.t12 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X96 CSoutput.t1 a_n9628_8799.t75 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 gnd.t284 commonsourceibias.t30 commonsourceibias.t31 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 a_n9628_8799.t38 a_n2982_13878.t78 a_n2982_8322.t32 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 CSoutput.t137 commonsourceibias.t74 gnd.t283 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 gnd.t282 commonsourceibias.t75 CSoutput.t136 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 CSoutput.t135 commonsourceibias.t76 gnd.t280 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 a_n2982_8322.t31 a_n2982_13878.t79 a_n9628_8799.t37 vdd.t276 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X103 gnd.t279 commonsourceibias.t77 CSoutput.t134 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 CSoutput.t164 a_n9628_8799.t76 vdd.t280 vdd.t279 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 a_n3106_n452.t19 minus.t9 a_n2982_13878.t15 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X106 a_n3106_n452.t49 plus.t11 a_n9628_8799.t19 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X107 output.t11 CSoutput.t199 vdd.t94 gnd.t165 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X108 vdd.t95 CSoutput.t200 output.t10 gnd.t166 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X109 a_n9628_8799.t17 plus.t12 a_n3106_n452.t48 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X110 vdd.t213 vdd.t210 vdd.t212 vdd.t211 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X111 gnd.t278 commonsourceibias.t78 CSoutput.t133 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 a_n3106_n452.t15 diffpairibias.t17 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X113 CSoutput.t165 a_n9628_8799.t77 vdd.t281 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 vdd.t45 a_n9628_8799.t78 CSoutput.t22 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 gnd.t137 gnd.t135 gnd.t136 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X116 vdd.t47 a_n9628_8799.t79 CSoutput.t23 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 a_n2982_13878.t58 a_n2982_13878.t57 a_n2804_13878.t26 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 a_n3106_n452.t47 plus.t13 a_n9628_8799.t14 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X119 vdd.t115 a_n9628_8799.t80 CSoutput.t64 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 gnd.t277 commonsourceibias.t79 CSoutput.t132 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 a_n9628_8799.t40 a_n2982_13878.t80 a_n2982_8322.t30 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 a_n2982_13878.t64 a_n2982_13878.t63 a_n2804_13878.t25 vdd.t227 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t134 gnd.t132 gnd.t133 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X124 vdd.t96 CSoutput.t201 output.t9 gnd.t167 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t116 a_n9628_8799.t81 CSoutput.t65 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X126 CSoutput.t88 a_n9628_8799.t82 vdd.t143 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 gnd.t276 commonsourceibias.t80 CSoutput.t131 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 a_n2982_13878.t18 minus.t10 a_n3106_n452.t22 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X129 CSoutput.t89 a_n9628_8799.t83 vdd.t144 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X130 vdd.t209 vdd.t207 vdd.t208 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 gnd.t275 commonsourceibias.t24 commonsourceibias.t25 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X132 output.t8 CSoutput.t202 vdd.t26 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X133 gnd.t274 commonsourceibias.t81 CSoutput.t130 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 CSoutput.t178 a_n9628_8799.t84 vdd.t294 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 vdd.t206 vdd.t203 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 a_n2804_13878.t24 a_n2982_13878.t23 a_n2982_13878.t24 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X137 CSoutput.t179 a_n9628_8799.t85 vdd.t295 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 vdd.t306 a_n9628_8799.t86 CSoutput.t190 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X139 vdd.t274 a_n2982_13878.t81 a_n2982_8322.t13 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X140 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t23 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 a_n2982_8322.t12 a_n2982_13878.t82 vdd.t272 vdd.t271 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 a_n3106_n452.t24 diffpairibias.t18 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 CSoutput.t191 a_n9628_8799.t87 vdd.t307 vdd.t279 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 output.t7 CSoutput.t203 vdd.t27 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X145 CSoutput.t129 commonsourceibias.t82 gnd.t273 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 gnd.t131 gnd.t129 gnd.t130 gnd.t76 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X147 CSoutput.t128 commonsourceibias.t83 gnd.t272 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 gnd.t128 gnd.t126 gnd.t127 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X149 gnd.t125 gnd.t123 minus.t4 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X150 vdd.t270 a_n2982_13878.t83 a_n2804_13878.t0 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 vdd.t202 vdd.t199 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X152 gnd.t122 gnd.t120 gnd.t121 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X153 a_n2804_13878.t22 a_n2982_13878.t21 a_n2982_13878.t22 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 vdd.t111 a_n9628_8799.t88 CSoutput.t60 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 vdd.t112 a_n9628_8799.t89 CSoutput.t61 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n2982_8322.t29 a_n2982_13878.t84 a_n9628_8799.t39 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 gnd.t111 gnd.t109 plus.t3 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X158 a_n9628_8799.t10 plus.t14 a_n3106_n452.t46 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X159 vdd.t198 vdd.t196 vdd.t197 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X160 a_n2982_13878.t20 minus.t11 a_n3106_n452.t25 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X161 vdd.t195 vdd.t192 vdd.t194 vdd.t193 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X162 a_n2982_8322.t11 a_n2982_13878.t85 vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X163 a_n9628_8799.t23 a_n2982_13878.t86 a_n2982_8322.t28 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 a_n9628_8799.t1 plus.t15 a_n3106_n452.t45 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X165 CSoutput.t44 a_n9628_8799.t90 vdd.t77 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 diffpairibias.t11 diffpairibias.t10 gnd.t325 gnd.t324 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X167 a_n2982_13878.t1 minus.t12 a_n3106_n452.t3 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X168 vdd.t78 a_n9628_8799.t91 CSoutput.t45 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X169 a_n2982_13878.t42 a_n2982_13878.t41 a_n2804_13878.t21 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X170 CSoutput.t127 commonsourceibias.t84 gnd.t271 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n9628_8799.t22 a_n2982_13878.t87 a_n2982_8322.t27 vdd.t265 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X172 CSoutput.t20 a_n9628_8799.t92 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 CSoutput.t21 a_n9628_8799.t93 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 commonsourceibias.t29 commonsourceibias.t28 gnd.t270 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t269 commonsourceibias.t85 CSoutput.t126 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 a_n2804_13878.t20 a_n2982_13878.t45 a_n2982_13878.t46 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 gnd.t119 gnd.t116 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X178 a_n3106_n452.t10 minus.t13 a_n2982_13878.t8 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 vdd.t191 vdd.t189 vdd.t190 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X180 outputibias.t7 outputibias.t6 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X181 vdd.t28 CSoutput.t204 output.t6 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X182 CSoutput.t12 a_n9628_8799.t94 vdd.t23 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 CSoutput.t125 commonsourceibias.t86 gnd.t268 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 vdd.t263 a_n2982_13878.t88 a_n2982_8322.t10 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X185 a_n2804_13878.t19 a_n2982_13878.t67 a_n2982_13878.t68 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X186 vdd.t25 a_n9628_8799.t95 CSoutput.t13 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 vdd.t65 a_n9628_8799.t96 CSoutput.t36 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 a_n2982_13878.t7 minus.t14 a_n3106_n452.t9 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X189 a_n3106_n452.t44 plus.t16 a_n9628_8799.t16 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X190 a_n2982_13878.t48 a_n2982_13878.t47 a_n2804_13878.t18 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X191 gnd.t267 commonsourceibias.t87 CSoutput.t124 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t266 commonsourceibias.t88 CSoutput.t123 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 commonsourceibias.t27 commonsourceibias.t26 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 outputibias.t5 outputibias.t4 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X195 gnd.t263 commonsourceibias.t89 CSoutput.t122 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X196 vdd.t67 a_n9628_8799.t97 CSoutput.t37 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X197 vdd.t59 a_n9628_8799.t98 CSoutput.t32 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 CSoutput.t121 commonsourceibias.t90 gnd.t262 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 CSoutput.t33 a_n9628_8799.t99 vdd.t60 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 a_n3106_n452.t27 diffpairibias.t19 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X201 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X202 vdd.t188 vdd.t186 vdd.t187 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X203 a_n3106_n452.t17 diffpairibias.t20 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X204 commonsourceibias.t7 commonsourceibias.t6 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 a_n9628_8799.t7 plus.t17 a_n3106_n452.t43 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X206 vdd.t54 a_n9628_8799.t100 CSoutput.t28 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 vdd.t55 a_n9628_8799.t101 CSoutput.t29 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 CSoutput.t42 a_n9628_8799.t102 vdd.t75 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd.t108 gnd.t106 gnd.t107 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X210 vdd.t185 vdd.t183 vdd.t184 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X211 CSoutput.t120 commonsourceibias.t91 gnd.t259 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 a_n9628_8799.t44 plus.t18 a_n3106_n452.t42 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X213 CSoutput.t119 commonsourceibias.t92 gnd.t258 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 a_n2804_13878.t17 a_n2982_13878.t25 a_n2982_13878.t26 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X215 gnd.t105 gnd.t103 gnd.t104 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X216 a_n2982_8322.t26 a_n2982_13878.t89 a_n9628_8799.t25 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 CSoutput.t43 a_n9628_8799.t103 vdd.t76 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 CSoutput.t176 a_n9628_8799.t104 vdd.t292 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 commonsourceibias.t5 commonsourceibias.t4 gnd.t257 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 minus.t3 gnd.t100 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X221 CSoutput.t205 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X222 diffpairibias.t9 diffpairibias.t8 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X223 a_n2804_13878.t6 a_n2982_13878.t90 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 a_n2982_13878.t10 minus.t15 a_n3106_n452.t12 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X225 vdd.t257 a_n2982_13878.t91 a_n2804_13878.t5 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X226 CSoutput.t118 commonsourceibias.t93 gnd.t256 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 CSoutput.t117 commonsourceibias.t94 gnd.t255 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 CSoutput.t177 a_n9628_8799.t105 vdd.t293 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t206 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X230 gnd.t254 commonsourceibias.t42 commonsourceibias.t43 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 a_n3106_n452.t41 plus.t19 a_n9628_8799.t6 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X232 vdd.t300 a_n9628_8799.t106 CSoutput.t184 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 vdd.t301 a_n9628_8799.t107 CSoutput.t185 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 vdd.t90 a_n9628_8799.t108 CSoutput.t50 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X235 commonsourceibias.t41 commonsourceibias.t40 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 CSoutput.t51 a_n9628_8799.t109 vdd.t91 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n2804_13878.t16 a_n2982_13878.t29 a_n2982_13878.t30 vdd.t255 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X238 gnd.t250 commonsourceibias.t95 CSoutput.t116 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 commonsourceibias.t39 commonsourceibias.t38 gnd.t249 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X240 vdd.t286 a_n9628_8799.t110 CSoutput.t170 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X241 vdd.t287 a_n9628_8799.t111 CSoutput.t171 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 output.t19 outputibias.t9 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X243 CSoutput.t4 a_n9628_8799.t112 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 gnd.t248 commonsourceibias.t36 commonsourceibias.t37 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 a_n3106_n452.t18 minus.t16 a_n2982_13878.t14 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X246 a_n2982_8322.t25 a_n2982_13878.t92 a_n9628_8799.t24 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X247 a_n2982_13878.t34 a_n2982_13878.t33 a_n2804_13878.t15 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 CSoutput.t5 a_n9628_8799.t113 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X249 diffpairibias.t7 diffpairibias.t6 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X250 gnd.t99 gnd.t97 gnd.t98 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 vdd.t38 a_n9628_8799.t114 CSoutput.t18 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X252 a_n2804_13878.t14 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X253 commonsourceibias.t35 commonsourceibias.t34 gnd.t247 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X254 vdd.t252 a_n2982_13878.t93 a_n2982_8322.t9 vdd.t251 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X255 vdd.t97 CSoutput.t207 output.t5 gnd.t170 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X256 vdd.t40 a_n9628_8799.t115 CSoutput.t19 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 a_n3106_n452.t1 minus.t17 a_n2982_13878.t0 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X258 a_n3106_n452.t40 plus.t20 a_n9628_8799.t12 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X259 gnd.t246 commonsourceibias.t96 CSoutput.t115 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 a_n3106_n452.t20 minus.t18 a_n2982_13878.t16 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X261 CSoutput.t58 a_n9628_8799.t116 vdd.t108 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 gnd.t245 commonsourceibias.t12 commonsourceibias.t13 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 a_n2804_13878.t7 a_n2982_13878.t94 vdd.t250 vdd.t249 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X264 vdd.t110 a_n9628_8799.t117 CSoutput.t59 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 CSoutput.t86 a_n9628_8799.t118 vdd.t141 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 CSoutput.t87 a_n9628_8799.t119 vdd.t142 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 gnd.t96 gnd.t93 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X268 vdd.t182 vdd.t180 vdd.t181 vdd.t156 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X269 vdd.t132 a_n9628_8799.t120 CSoutput.t78 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X270 a_n3106_n452.t0 diffpairibias.t21 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 minus.t2 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X272 a_n2982_8322.t24 a_n2982_13878.t95 a_n9628_8799.t27 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X273 vdd.t247 a_n2982_13878.t96 a_n2982_8322.t8 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X274 gnd.t243 commonsourceibias.t10 commonsourceibias.t11 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n9628_8799.t18 plus.t21 a_n3106_n452.t39 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X276 a_n2982_13878.t2 minus.t19 a_n3106_n452.t4 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X277 vdd.t133 a_n9628_8799.t121 CSoutput.t79 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 a_n3106_n452.t5 minus.t20 a_n2982_13878.t3 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X279 gnd.t242 commonsourceibias.t8 commonsourceibias.t9 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t179 vdd.t176 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X281 vdd.t139 a_n9628_8799.t122 CSoutput.t84 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 a_n3106_n452.t13 minus.t21 a_n2982_13878.t11 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X283 vdd.t140 a_n9628_8799.t123 CSoutput.t85 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 output.t4 CSoutput.t208 vdd.t98 gnd.t171 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X285 vdd.t130 a_n9628_8799.t124 CSoutput.t76 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 CSoutput.t77 a_n9628_8799.t125 vdd.t131 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 CSoutput.t174 a_n9628_8799.t126 vdd.t290 vdd.t279 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t114 commonsourceibias.t97 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 a_n3106_n452.t11 minus.t22 a_n2982_13878.t9 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X290 a_n2804_13878.t13 a_n2982_13878.t43 a_n2982_13878.t44 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X291 CSoutput.t175 a_n9628_8799.t127 vdd.t291 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t188 a_n9628_8799.t128 vdd.t304 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X293 a_n2982_8322.t23 a_n2982_13878.t97 a_n9628_8799.t26 vdd.t245 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X294 diffpairibias.t5 diffpairibias.t4 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X295 gnd.t89 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X296 CSoutput.t189 a_n9628_8799.t129 vdd.t305 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 CSoutput.t56 a_n9628_8799.t130 vdd.t105 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t175 vdd.t172 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X299 CSoutput.t113 commonsourceibias.t98 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X300 vdd.t107 a_n9628_8799.t131 CSoutput.t57 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t209 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X302 gnd.t85 gnd.t82 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X303 a_n2982_8322.t7 a_n2982_13878.t98 vdd.t244 vdd.t243 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X304 CSoutput.t40 a_n9628_8799.t132 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 outputibias.t3 outputibias.t2 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X306 a_n3106_n452.t16 minus.t23 a_n2982_13878.t13 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X307 vdd.t74 a_n9628_8799.t133 CSoutput.t41 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 gnd.t81 gnd.t79 gnd.t80 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X309 gnd.t237 commonsourceibias.t99 CSoutput.t112 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 CSoutput.t16 a_n9628_8799.t134 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 output.t0 outputibias.t10 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X312 vdd.t242 a_n2982_13878.t99 a_n2804_13878.t4 vdd.t241 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X313 vdd.t36 a_n9628_8799.t135 CSoutput.t17 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X314 CSoutput.t10 a_n9628_8799.t136 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 gnd.t78 gnd.t75 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X316 vdd.t22 a_n9628_8799.t137 CSoutput.t11 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 gnd.t74 gnd.t72 plus.t2 gnd.t73 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X318 gnd.t236 commonsourceibias.t100 CSoutput.t111 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 output.t18 outputibias.t11 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X320 gnd.t235 commonsourceibias.t101 CSoutput.t110 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 a_n2982_8322.t22 a_n2982_13878.t100 a_n9628_8799.t33 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X322 gnd.t71 gnd.t69 gnd.t70 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X323 commonsourceibias.t17 commonsourceibias.t16 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 a_n9628_8799.t32 a_n2982_13878.t101 a_n2982_8322.t21 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X325 a_n2804_13878.t3 a_n2982_13878.t102 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X326 gnd.t232 commonsourceibias.t102 CSoutput.t109 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 vdd.t62 a_n9628_8799.t138 CSoutput.t34 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 vdd.t171 vdd.t169 vdd.t170 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X329 vdd.t168 vdd.t166 vdd.t167 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X330 vdd.t63 a_n9628_8799.t139 CSoutput.t35 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 CSoutput.t30 a_n9628_8799.t140 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t31 a_n9628_8799.t141 vdd.t58 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X333 CSoutput.t26 a_n9628_8799.t142 vdd.t51 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 a_n2982_13878.t66 a_n2982_13878.t65 a_n2804_13878.t12 vdd.t228 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 a_n9628_8799.t21 a_n2982_13878.t103 a_n2982_8322.t20 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X336 a_n3106_n452.t38 plus.t22 a_n9628_8799.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X337 a_n9628_8799.t20 a_n2982_13878.t104 a_n2982_8322.t19 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X338 a_n2982_13878.t4 minus.t24 a_n3106_n452.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X339 a_n9628_8799.t2 plus.t23 a_n3106_n452.t37 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X340 gnd.t231 commonsourceibias.t103 CSoutput.t108 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 gnd.t68 gnd.t66 minus.t1 gnd.t67 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X342 a_n2982_8322.t18 a_n2982_13878.t105 a_n9628_8799.t31 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X343 commonsourceibias.t15 commonsourceibias.t14 gnd.t230 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t228 commonsourceibias.t104 CSoutput.t107 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 a_n2982_13878.t69 minus.t25 a_n3106_n452.t28 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 vdd.t53 a_n9628_8799.t143 CSoutput.t27 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 gnd.t226 commonsourceibias.t22 commonsourceibias.t23 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 CSoutput.t38 a_n9628_8799.t144 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 CSoutput.t39 a_n9628_8799.t145 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X350 CSoutput.t172 a_n9628_8799.t146 vdd.t288 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 CSoutput.t173 a_n9628_8799.t147 vdd.t289 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 a_n2804_13878.t11 a_n2982_13878.t39 a_n2982_13878.t40 vdd.t234 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 vdd.t298 a_n9628_8799.t148 CSoutput.t182 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 vdd.t299 a_n9628_8799.t149 CSoutput.t183 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 vdd.t86 a_n9628_8799.t150 CSoutput.t48 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X356 gnd.t224 commonsourceibias.t20 commonsourceibias.t21 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X357 commonsourceibias.t19 commonsourceibias.t18 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 a_n3106_n452.t8 minus.t26 a_n2982_13878.t6 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X359 gnd.t221 commonsourceibias.t105 CSoutput.t106 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 a_n3106_n452.t26 diffpairibias.t22 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X361 CSoutput.t105 commonsourceibias.t106 gnd.t219 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 output.t3 CSoutput.t210 vdd.t82 gnd.t157 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X363 vdd.t88 a_n9628_8799.t151 CSoutput.t49 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 gnd.t218 commonsourceibias.t107 CSoutput.t104 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 CSoutput.t168 a_n9628_8799.t152 vdd.t284 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 a_n2982_13878.t62 a_n2982_13878.t61 a_n2804_13878.t10 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X367 gnd.t65 gnd.t62 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X368 a_n9628_8799.t30 a_n2982_13878.t106 a_n2982_8322.t17 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 a_n9628_8799.t11 plus.t24 a_n3106_n452.t36 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X370 gnd.t61 gnd.t58 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X371 vdd.t285 a_n9628_8799.t153 CSoutput.t169 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 CSoutput.t211 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X373 CSoutput.t2 a_n9628_8799.t154 vdd.t6 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 vdd.t165 vdd.t163 vdd.t164 vdd.t156 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X375 CSoutput.t103 commonsourceibias.t108 gnd.t216 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 gnd.t215 commonsourceibias.t109 CSoutput.t102 gnd.t214 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X377 commonsourceibias.t47 commonsourceibias.t46 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 diffpairibias.t3 diffpairibias.t2 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X379 gnd.t57 gnd.t54 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X380 CSoutput.t3 a_n9628_8799.t155 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 outputibias.t1 outputibias.t0 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X382 a_n2982_8322.t16 a_n2982_13878.t107 a_n9628_8799.t29 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X383 gnd.t211 commonsourceibias.t110 CSoutput.t101 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 a_n2982_13878.t12 minus.t27 a_n3106_n452.t14 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X385 gnd.t53 gnd.t51 plus.t1 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X386 vdd.t30 a_n9628_8799.t156 CSoutput.t14 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 vdd.t162 vdd.t159 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X388 gnd.t50 gnd.t47 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X389 CSoutput.t15 a_n9628_8799.t157 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X390 CSoutput.t54 a_n9628_8799.t158 vdd.t102 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 diffpairibias.t1 diffpairibias.t0 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X392 commonsourceibias.t45 commonsourceibias.t44 gnd.t209 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 gnd.t210 commonsourceibias.t111 CSoutput.t100 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X394 CSoutput.t99 commonsourceibias.t112 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X395 vdd.t230 a_n2982_13878.t108 a_n2804_13878.t2 vdd.t229 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X396 CSoutput.t55 a_n9628_8799.t159 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 CSoutput.t82 a_n9628_8799.t160 vdd.t137 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X398 vdd.t138 a_n9628_8799.t161 CSoutput.t83 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 plus.t0 gnd.t44 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X400 vdd.t128 a_n9628_8799.t162 CSoutput.t74 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 gnd.t206 commonsourceibias.t2 commonsourceibias.t3 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 a_n9628_8799.t46 plus.t25 a_n3106_n452.t35 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X403 gnd.t43 gnd.t41 minus.t0 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X404 vdd.t83 CSoutput.t212 output.t2 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X405 a_n2982_8322.t15 a_n2982_13878.t109 a_n9628_8799.t28 vdd.t228 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X406 a_n2982_13878.t17 minus.t28 a_n3106_n452.t21 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X407 output.t1 CSoutput.t213 vdd.t84 gnd.t159 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X408 gnd.t204 commonsourceibias.t113 CSoutput.t98 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X409 a_n9628_8799.t45 plus.t26 a_n3106_n452.t34 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X410 gnd.t202 commonsourceibias.t114 CSoutput.t97 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 gnd.t40 gnd.t37 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X412 a_n2982_8322.t14 a_n2982_13878.t110 a_n9628_8799.t34 vdd.t227 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X413 vdd.t129 a_n9628_8799.t163 CSoutput.t75 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 vdd.t134 a_n9628_8799.t164 CSoutput.t80 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 CSoutput.t81 a_n9628_8799.t165 vdd.t136 vdd.t135 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 gnd.t200 commonsourceibias.t115 CSoutput.t96 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X417 vdd.t158 vdd.t155 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X418 a_n2982_8322.t6 a_n2982_13878.t111 vdd.t226 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X419 gnd.t199 commonsourceibias.t116 CSoutput.t95 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X420 a_n2804_13878.t9 a_n2982_13878.t53 a_n2982_13878.t54 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X421 gnd.t197 commonsourceibias.t117 CSoutput.t94 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X422 CSoutput.t93 commonsourceibias.t118 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 CSoutput.t92 commonsourceibias.t119 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 vdd.t154 vdd.t151 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X425 a_n3106_n452.t33 plus.t27 a_n9628_8799.t47 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X426 a_n3106_n452.t30 diffpairibias.t23 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X427 vdd.t150 vdd.t147 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X428 vdd.t126 a_n9628_8799.t166 CSoutput.t72 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X429 CSoutput.t73 a_n9628_8799.t167 vdd.t127 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X430 a_n2982_13878.t32 a_n2982_13878.t31 a_n2804_13878.t8 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X431 a_n3106_n452.t32 plus.t28 a_n9628_8799.t9 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
R0 a_n2982_13878.n15 a_n2982_13878.t110 538.698
R1 a_n2982_13878.n146 a_n2982_13878.t87 512.366
R2 a_n2982_13878.n145 a_n2982_13878.t92 512.366
R3 a_n2982_13878.n98 a_n2982_13878.t80 512.366
R4 a_n2982_13878.n144 a_n2982_13878.t97 512.366
R5 a_n2982_13878.n143 a_n2982_13878.t106 512.366
R6 a_n2982_13878.n99 a_n2982_13878.t107 512.366
R7 a_n2982_13878.n142 a_n2982_13878.t74 512.366
R8 a_n2982_13878.n141 a_n2982_13878.t89 512.366
R9 a_n2982_13878.n100 a_n2982_13878.t77 512.366
R10 a_n2982_13878.n140 a_n2982_13878.t84 512.366
R11 a_n2982_13878.n9 a_n2982_13878.t65 538.698
R12 a_n2982_13878.n154 a_n2982_13878.t21 512.366
R13 a_n2982_13878.n153 a_n2982_13878.t49 512.366
R14 a_n2982_13878.n83 a_n2982_13878.t25 512.366
R15 a_n2982_13878.n152 a_n2982_13878.t35 512.366
R16 a_n2982_13878.n151 a_n2982_13878.t29 512.366
R17 a_n2982_13878.n84 a_n2982_13878.t61 512.366
R18 a_n2982_13878.n150 a_n2982_13878.t43 512.366
R19 a_n2982_13878.n149 a_n2982_13878.t57 512.366
R20 a_n2982_13878.n97 a_n2982_13878.t39 512.366
R21 a_n2982_13878.n147 a_n2982_13878.t41 512.366
R22 a_n2982_13878.n31 a_n2982_13878.t63 538.698
R23 a_n2982_13878.n120 a_n2982_13878.t37 512.366
R24 a_n2982_13878.n109 a_n2982_13878.t31 512.366
R25 a_n2982_13878.n121 a_n2982_13878.t45 512.366
R26 a_n2982_13878.n108 a_n2982_13878.t27 512.366
R27 a_n2982_13878.n122 a_n2982_13878.t59 512.366
R28 a_n2982_13878.n123 a_n2982_13878.t47 512.366
R29 a_n2982_13878.n107 a_n2982_13878.t67 512.366
R30 a_n2982_13878.n124 a_n2982_13878.t51 512.366
R31 a_n2982_13878.n106 a_n2982_13878.t55 512.366
R32 a_n2982_13878.n125 a_n2982_13878.t33 512.366
R33 a_n2982_13878.n37 a_n2982_13878.t109 538.698
R34 a_n2982_13878.n114 a_n2982_13878.t78 512.366
R35 a_n2982_13878.n113 a_n2982_13878.t79 512.366
R36 a_n2982_13878.n115 a_n2982_13878.t104 512.366
R37 a_n2982_13878.n112 a_n2982_13878.t105 512.366
R38 a_n2982_13878.n116 a_n2982_13878.t76 512.366
R39 a_n2982_13878.n117 a_n2982_13878.t100 512.366
R40 a_n2982_13878.n111 a_n2982_13878.t101 512.366
R41 a_n2982_13878.n118 a_n2982_13878.t73 512.366
R42 a_n2982_13878.n110 a_n2982_13878.t86 512.366
R43 a_n2982_13878.n119 a_n2982_13878.t95 512.366
R44 a_n2982_13878.n137 a_n2982_13878.t94 512.366
R45 a_n2982_13878.n127 a_n2982_13878.t83 512.366
R46 a_n2982_13878.n138 a_n2982_13878.t72 512.366
R47 a_n2982_13878.n135 a_n2982_13878.t102 512.366
R48 a_n2982_13878.n128 a_n2982_13878.t91 512.366
R49 a_n2982_13878.n136 a_n2982_13878.t90 512.366
R50 a_n2982_13878.n133 a_n2982_13878.t98 512.366
R51 a_n2982_13878.n129 a_n2982_13878.t81 512.366
R52 a_n2982_13878.n134 a_n2982_13878.t82 512.366
R53 a_n2982_13878.n131 a_n2982_13878.t85 512.366
R54 a_n2982_13878.n130 a_n2982_13878.t96 512.366
R55 a_n2982_13878.n132 a_n2982_13878.t111 512.366
R56 a_n2982_13878.n77 a_n2982_13878.n10 70.5844
R57 a_n2982_13878.n69 a_n2982_13878.n16 70.5844
R58 a_n2982_13878.n27 a_n2982_13878.n59 70.5844
R59 a_n2982_13878.n33 a_n2982_13878.n51 70.5844
R60 a_n2982_13878.n50 a_n2982_13878.n33 70.1674
R61 a_n2982_13878.n50 a_n2982_13878.n110 20.9683
R62 a_n2982_13878.n32 a_n2982_13878.n49 74.73
R63 a_n2982_13878.n118 a_n2982_13878.n49 11.843
R64 a_n2982_13878.n48 a_n2982_13878.n32 80.4688
R65 a_n2982_13878.n48 a_n2982_13878.n111 0.365327
R66 a_n2982_13878.n34 a_n2982_13878.n47 75.0448
R67 a_n2982_13878.n46 a_n2982_13878.n34 70.1674
R68 a_n2982_13878.n46 a_n2982_13878.n112 20.9683
R69 a_n2982_13878.n35 a_n2982_13878.n45 70.3058
R70 a_n2982_13878.n115 a_n2982_13878.n45 20.6913
R71 a_n2982_13878.n44 a_n2982_13878.n35 75.3623
R72 a_n2982_13878.n44 a_n2982_13878.n113 10.5784
R73 a_n2982_13878.n37 a_n2982_13878.n36 44.7878
R74 a_n2982_13878.n58 a_n2982_13878.n27 70.1674
R75 a_n2982_13878.n58 a_n2982_13878.n106 20.9683
R76 a_n2982_13878.n26 a_n2982_13878.n57 74.73
R77 a_n2982_13878.n124 a_n2982_13878.n57 11.843
R78 a_n2982_13878.n56 a_n2982_13878.n26 80.4688
R79 a_n2982_13878.n56 a_n2982_13878.n107 0.365327
R80 a_n2982_13878.n28 a_n2982_13878.n55 75.0448
R81 a_n2982_13878.n54 a_n2982_13878.n28 70.1674
R82 a_n2982_13878.n54 a_n2982_13878.n108 20.9683
R83 a_n2982_13878.n29 a_n2982_13878.n53 70.3058
R84 a_n2982_13878.n121 a_n2982_13878.n53 20.6913
R85 a_n2982_13878.n52 a_n2982_13878.n29 75.3623
R86 a_n2982_13878.n52 a_n2982_13878.n109 10.5784
R87 a_n2982_13878.n31 a_n2982_13878.n30 44.7878
R88 a_n2982_13878.n17 a_n2982_13878.n67 70.1674
R89 a_n2982_13878.n19 a_n2982_13878.n65 70.1674
R90 a_n2982_13878.n21 a_n2982_13878.n63 70.1674
R91 a_n2982_13878.n24 a_n2982_13878.n61 70.1674
R92 a_n2982_13878.n132 a_n2982_13878.n61 20.9683
R93 a_n2982_13878.n60 a_n2982_13878.n25 75.0448
R94 a_n2982_13878.n60 a_n2982_13878.n130 11.2134
R95 a_n2982_13878.n25 a_n2982_13878.n131 161.3
R96 a_n2982_13878.n134 a_n2982_13878.n63 20.9683
R97 a_n2982_13878.n62 a_n2982_13878.n22 75.0448
R98 a_n2982_13878.n62 a_n2982_13878.n129 11.2134
R99 a_n2982_13878.n22 a_n2982_13878.n133 161.3
R100 a_n2982_13878.n136 a_n2982_13878.n65 20.9683
R101 a_n2982_13878.n64 a_n2982_13878.n20 75.0448
R102 a_n2982_13878.n64 a_n2982_13878.n128 11.2134
R103 a_n2982_13878.n20 a_n2982_13878.n135 161.3
R104 a_n2982_13878.n138 a_n2982_13878.n67 20.9683
R105 a_n2982_13878.n66 a_n2982_13878.n18 75.0448
R106 a_n2982_13878.n66 a_n2982_13878.n127 11.2134
R107 a_n2982_13878.n18 a_n2982_13878.n137 161.3
R108 a_n2982_13878.n16 a_n2982_13878.n68 70.1674
R109 a_n2982_13878.n68 a_n2982_13878.n97 20.9683
R110 a_n2982_13878.n148 a_n2982_13878.n5 161.3
R111 a_n2982_13878.n10 a_n2982_13878.n76 70.1674
R112 a_n2982_13878.n76 a_n2982_13878.n100 20.9683
R113 a_n2982_13878.n75 a_n2982_13878.n11 74.73
R114 a_n2982_13878.n141 a_n2982_13878.n75 11.843
R115 a_n2982_13878.n74 a_n2982_13878.n11 80.4688
R116 a_n2982_13878.n74 a_n2982_13878.n142 0.365327
R117 a_n2982_13878.n12 a_n2982_13878.n73 75.0448
R118 a_n2982_13878.n72 a_n2982_13878.n12 70.1674
R119 a_n2982_13878.n144 a_n2982_13878.n72 20.9683
R120 a_n2982_13878.n14 a_n2982_13878.n71 70.3058
R121 a_n2982_13878.n71 a_n2982_13878.n98 20.6913
R122 a_n2982_13878.n70 a_n2982_13878.n14 75.3623
R123 a_n2982_13878.n145 a_n2982_13878.n70 10.5784
R124 a_n2982_13878.n13 a_n2982_13878.n15 44.7878
R125 a_n2982_13878.n82 a_n2982_13878.n5 44.8194
R126 a_n2982_13878.n82 a_n2982_13878.n150 13.6566
R127 a_n2982_13878.n6 a_n2982_13878.n81 75.0448
R128 a_n2982_13878.n80 a_n2982_13878.n6 70.1674
R129 a_n2982_13878.n152 a_n2982_13878.n80 20.9683
R130 a_n2982_13878.n8 a_n2982_13878.n79 70.3058
R131 a_n2982_13878.n79 a_n2982_13878.n83 20.6913
R132 a_n2982_13878.n78 a_n2982_13878.n8 75.3623
R133 a_n2982_13878.n153 a_n2982_13878.n78 10.5784
R134 a_n2982_13878.n7 a_n2982_13878.n9 44.7878
R135 a_n2982_13878.n3 a_n2982_13878.n94 81.4626
R136 a_n2982_13878.n4 a_n2982_13878.n88 81.4626
R137 a_n2982_13878.n0 a_n2982_13878.n85 81.4626
R138 a_n2982_13878.n3 a_n2982_13878.n95 80.9324
R139 a_n2982_13878.n2 a_n2982_13878.n96 80.9324
R140 a_n2982_13878.n2 a_n2982_13878.n93 80.9324
R141 a_n2982_13878.n2 a_n2982_13878.n92 80.9324
R142 a_n2982_13878.n1 a_n2982_13878.n91 80.9324
R143 a_n2982_13878.n4 a_n2982_13878.n89 80.9324
R144 a_n2982_13878.n0 a_n2982_13878.n90 80.9324
R145 a_n2982_13878.n0 a_n2982_13878.n87 80.9324
R146 a_n2982_13878.n0 a_n2982_13878.n86 80.9324
R147 a_n2982_13878.n43 a_n2982_13878.t54 74.6477
R148 a_n2982_13878.n38 a_n2982_13878.t64 74.6477
R149 a_n2982_13878.n42 a_n2982_13878.t66 74.2899
R150 a_n2982_13878.n40 a_n2982_13878.t24 74.2897
R151 a_n2982_13878.n43 a_n2982_13878.n156 70.6783
R152 a_n2982_13878.n43 a_n2982_13878.n157 70.6783
R153 a_n2982_13878.n41 a_n2982_13878.n158 70.6783
R154 a_n2982_13878.n41 a_n2982_13878.n159 70.6783
R155 a_n2982_13878.n40 a_n2982_13878.n105 70.6783
R156 a_n2982_13878.n39 a_n2982_13878.n104 70.6783
R157 a_n2982_13878.n39 a_n2982_13878.n103 70.6783
R158 a_n2982_13878.n38 a_n2982_13878.n102 70.6783
R159 a_n2982_13878.n38 a_n2982_13878.n101 70.6783
R160 a_n2982_13878.n160 a_n2982_13878.n42 70.6782
R161 a_n2982_13878.n146 a_n2982_13878.n145 48.2005
R162 a_n2982_13878.n72 a_n2982_13878.n143 20.9683
R163 a_n2982_13878.n142 a_n2982_13878.n99 48.2005
R164 a_n2982_13878.n140 a_n2982_13878.n76 20.9683
R165 a_n2982_13878.n154 a_n2982_13878.n153 48.2005
R166 a_n2982_13878.n80 a_n2982_13878.n151 20.9683
R167 a_n2982_13878.n150 a_n2982_13878.n84 48.2005
R168 a_n2982_13878.n147 a_n2982_13878.n68 20.9683
R169 a_n2982_13878.n120 a_n2982_13878.n109 48.2005
R170 a_n2982_13878.n122 a_n2982_13878.n54 20.9683
R171 a_n2982_13878.n123 a_n2982_13878.n107 48.2005
R172 a_n2982_13878.n125 a_n2982_13878.n58 20.9683
R173 a_n2982_13878.n114 a_n2982_13878.n113 48.2005
R174 a_n2982_13878.n116 a_n2982_13878.n46 20.9683
R175 a_n2982_13878.n117 a_n2982_13878.n111 48.2005
R176 a_n2982_13878.n119 a_n2982_13878.n50 20.9683
R177 a_n2982_13878.n137 a_n2982_13878.n127 48.2005
R178 a_n2982_13878.t99 a_n2982_13878.n67 533.335
R179 a_n2982_13878.n135 a_n2982_13878.n128 48.2005
R180 a_n2982_13878.t108 a_n2982_13878.n65 533.335
R181 a_n2982_13878.n133 a_n2982_13878.n129 48.2005
R182 a_n2982_13878.t93 a_n2982_13878.n63 533.335
R183 a_n2982_13878.n131 a_n2982_13878.n130 48.2005
R184 a_n2982_13878.t88 a_n2982_13878.n61 533.335
R185 a_n2982_13878.n144 a_n2982_13878.n71 21.4216
R186 a_n2982_13878.n152 a_n2982_13878.n79 21.4216
R187 a_n2982_13878.n108 a_n2982_13878.n53 21.4216
R188 a_n2982_13878.n112 a_n2982_13878.n45 21.4216
R189 a_n2982_13878.n77 a_n2982_13878.t103 532.5
R190 a_n2982_13878.n69 a_n2982_13878.t53 532.5
R191 a_n2982_13878.t23 a_n2982_13878.n59 532.5
R192 a_n2982_13878.t75 a_n2982_13878.n51 532.5
R193 a_n2982_13878.n1 a_n2982_13878.n0 33.585
R194 a_n2982_13878.n75 a_n2982_13878.n100 34.4824
R195 a_n2982_13878.n149 a_n2982_13878.n148 25.5611
R196 a_n2982_13878.n106 a_n2982_13878.n57 34.4824
R197 a_n2982_13878.n110 a_n2982_13878.n49 34.4824
R198 a_n2982_13878.n143 a_n2982_13878.n73 35.3134
R199 a_n2982_13878.n73 a_n2982_13878.n99 11.2134
R200 a_n2982_13878.n151 a_n2982_13878.n81 35.3134
R201 a_n2982_13878.n81 a_n2982_13878.n84 11.2134
R202 a_n2982_13878.n55 a_n2982_13878.n122 35.3134
R203 a_n2982_13878.n123 a_n2982_13878.n55 11.2134
R204 a_n2982_13878.n47 a_n2982_13878.n116 35.3134
R205 a_n2982_13878.n117 a_n2982_13878.n47 11.2134
R206 a_n2982_13878.n138 a_n2982_13878.n66 35.3134
R207 a_n2982_13878.n136 a_n2982_13878.n64 35.3134
R208 a_n2982_13878.n134 a_n2982_13878.n62 35.3134
R209 a_n2982_13878.n132 a_n2982_13878.n60 35.3134
R210 a_n2982_13878.n5 a_n2982_13878.n2 23.891
R211 a_n2982_13878.n70 a_n2982_13878.n98 36.139
R212 a_n2982_13878.n78 a_n2982_13878.n83 36.139
R213 a_n2982_13878.n148 a_n2982_13878.n97 22.6399
R214 a_n2982_13878.n121 a_n2982_13878.n52 36.139
R215 a_n2982_13878.n115 a_n2982_13878.n44 36.139
R216 a_n2982_13878.n36 a_n2982_13878.n23 13.9285
R217 a_n2982_13878.n10 a_n2982_13878.n139 13.724
R218 a_n2982_13878.n155 a_n2982_13878.n7 12.4191
R219 a_n2982_13878.n25 a_n2982_13878.n23 11.2486
R220 a_n2982_13878.n139 a_n2982_13878.n17 11.2486
R221 a_n2982_13878.n126 a_n2982_13878.n40 10.5745
R222 a_n2982_13878.n126 a_n2982_13878.n27 8.58383
R223 a_n2982_13878.n42 a_n2982_13878.n155 6.7311
R224 a_n2982_13878.n139 a_n2982_13878.n126 5.3452
R225 a_n2982_13878.n30 a_n2982_13878.n33 3.94368
R226 a_n2982_13878.n16 a_n2982_13878.n13 3.94368
R227 a_n2982_13878.n156 a_n2982_13878.t40 3.61217
R228 a_n2982_13878.n156 a_n2982_13878.t42 3.61217
R229 a_n2982_13878.n157 a_n2982_13878.t44 3.61217
R230 a_n2982_13878.n157 a_n2982_13878.t58 3.61217
R231 a_n2982_13878.n158 a_n2982_13878.t30 3.61217
R232 a_n2982_13878.n158 a_n2982_13878.t62 3.61217
R233 a_n2982_13878.n159 a_n2982_13878.t26 3.61217
R234 a_n2982_13878.n159 a_n2982_13878.t36 3.61217
R235 a_n2982_13878.n105 a_n2982_13878.t56 3.61217
R236 a_n2982_13878.n105 a_n2982_13878.t34 3.61217
R237 a_n2982_13878.n104 a_n2982_13878.t68 3.61217
R238 a_n2982_13878.n104 a_n2982_13878.t52 3.61217
R239 a_n2982_13878.n103 a_n2982_13878.t60 3.61217
R240 a_n2982_13878.n103 a_n2982_13878.t48 3.61217
R241 a_n2982_13878.n102 a_n2982_13878.t46 3.61217
R242 a_n2982_13878.n102 a_n2982_13878.t28 3.61217
R243 a_n2982_13878.n101 a_n2982_13878.t38 3.61217
R244 a_n2982_13878.n101 a_n2982_13878.t32 3.61217
R245 a_n2982_13878.t22 a_n2982_13878.n160 3.61217
R246 a_n2982_13878.n160 a_n2982_13878.t50 3.61217
R247 a_n2982_13878.n94 a_n2982_13878.t13 2.82907
R248 a_n2982_13878.n94 a_n2982_13878.t17 2.82907
R249 a_n2982_13878.n95 a_n2982_13878.t14 2.82907
R250 a_n2982_13878.n95 a_n2982_13878.t10 2.82907
R251 a_n2982_13878.n96 a_n2982_13878.t19 2.82907
R252 a_n2982_13878.n96 a_n2982_13878.t5 2.82907
R253 a_n2982_13878.n93 a_n2982_13878.t9 2.82907
R254 a_n2982_13878.n93 a_n2982_13878.t2 2.82907
R255 a_n2982_13878.n92 a_n2982_13878.t16 2.82907
R256 a_n2982_13878.n92 a_n2982_13878.t69 2.82907
R257 a_n2982_13878.n91 a_n2982_13878.t70 2.82907
R258 a_n2982_13878.n91 a_n2982_13878.t1 2.82907
R259 a_n2982_13878.n88 a_n2982_13878.t8 2.82907
R260 a_n2982_13878.n88 a_n2982_13878.t18 2.82907
R261 a_n2982_13878.n89 a_n2982_13878.t0 2.82907
R262 a_n2982_13878.n89 a_n2982_13878.t20 2.82907
R263 a_n2982_13878.n90 a_n2982_13878.t11 2.82907
R264 a_n2982_13878.n90 a_n2982_13878.t4 2.82907
R265 a_n2982_13878.n87 a_n2982_13878.t6 2.82907
R266 a_n2982_13878.n87 a_n2982_13878.t12 2.82907
R267 a_n2982_13878.n86 a_n2982_13878.t15 2.82907
R268 a_n2982_13878.n86 a_n2982_13878.t71 2.82907
R269 a_n2982_13878.n85 a_n2982_13878.t3 2.82907
R270 a_n2982_13878.n85 a_n2982_13878.t7 2.82907
R271 a_n2982_13878.n15 a_n2982_13878.n146 14.1668
R272 a_n2982_13878.n140 a_n2982_13878.n77 22.3251
R273 a_n2982_13878.n9 a_n2982_13878.n154 14.1668
R274 a_n2982_13878.n147 a_n2982_13878.n69 22.3251
R275 a_n2982_13878.n120 a_n2982_13878.n31 14.1668
R276 a_n2982_13878.n59 a_n2982_13878.n125 22.3251
R277 a_n2982_13878.n114 a_n2982_13878.n37 14.1668
R278 a_n2982_13878.n51 a_n2982_13878.n119 22.3251
R279 a_n2982_13878.n155 a_n2982_13878.n23 1.30542
R280 a_n2982_13878.n20 a_n2982_13878.n21 1.04595
R281 a_n2982_13878.n74 a_n2982_13878.n141 47.835
R282 a_n2982_13878.n82 a_n2982_13878.n149 26.6438
R283 a_n2982_13878.n124 a_n2982_13878.n56 47.835
R284 a_n2982_13878.n118 a_n2982_13878.n48 47.835
R285 a_n2982_13878.n0 a_n2982_13878.n4 1.59102
R286 a_n2982_13878.n33 a_n2982_13878.n32 1.13686
R287 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R288 a_n2982_13878.n11 a_n2982_13878.n10 1.13686
R289 a_n2982_13878.n5 a_n2982_13878.n16 1.09898
R290 a_n2982_13878.n42 a_n2982_13878.n41 1.07378
R291 a_n2982_13878.n39 a_n2982_13878.n38 1.07378
R292 a_n2982_13878.n2 a_n2982_13878.n3 1.06084
R293 a_n2982_13878.n2 a_n2982_13878.n1 1.06084
R294 a_n2982_13878.n35 a_n2982_13878.n36 0.758076
R295 a_n2982_13878.n34 a_n2982_13878.n35 0.758076
R296 a_n2982_13878.n32 a_n2982_13878.n34 0.758076
R297 a_n2982_13878.n29 a_n2982_13878.n30 0.758076
R298 a_n2982_13878.n28 a_n2982_13878.n29 0.758076
R299 a_n2982_13878.n26 a_n2982_13878.n28 0.758076
R300 a_n2982_13878.n25 a_n2982_13878.n24 0.758076
R301 a_n2982_13878.n22 a_n2982_13878.n21 0.758076
R302 a_n2982_13878.n20 a_n2982_13878.n19 0.758076
R303 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R304 a_n2982_13878.n14 a_n2982_13878.n13 0.758076
R305 a_n2982_13878.n14 a_n2982_13878.n12 0.758076
R306 a_n2982_13878.n12 a_n2982_13878.n11 0.758076
R307 a_n2982_13878.n8 a_n2982_13878.n7 0.758076
R308 a_n2982_13878.n8 a_n2982_13878.n6 0.758076
R309 a_n2982_13878.n6 a_n2982_13878.n5 0.758076
R310 a_n2982_13878.n41 a_n2982_13878.n43 0.716017
R311 a_n2982_13878.n40 a_n2982_13878.n39 0.716017
R312 a_n2982_13878.n22 a_n2982_13878.n24 0.67853
R313 a_n2982_13878.n18 a_n2982_13878.n19 0.67853
R314 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R315 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R316 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R317 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R318 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R319 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R320 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R321 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R322 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R323 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R324 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R325 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R326 a_n2804_13878.n15 a_n2804_13878.t3 74.6477
R327 a_n2804_13878.n20 a_n2804_13878.t4 74.2899
R328 a_n2804_13878.n17 a_n2804_13878.t7 74.2899
R329 a_n2804_13878.n16 a_n2804_13878.t2 74.2899
R330 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R331 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R332 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R333 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R334 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R335 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R336 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R337 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R338 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R339 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R340 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R341 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R342 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R343 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R344 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R345 a_n2804_13878.n18 a_n2804_13878.t0 3.61217
R346 a_n2804_13878.n18 a_n2804_13878.t1 3.61217
R347 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R348 a_n2804_13878.n14 a_n2804_13878.t6 3.61217
R349 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R350 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R351 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R352 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R353 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R354 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R355 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R356 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R357 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R358 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R359 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R360 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R361 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R362 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R363 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R364 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R365 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R366 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R367 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R368 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R369 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R370 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R371 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R372 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R373 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R374 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R375 vdd.n327 vdd.n291 756.745
R376 vdd.n268 vdd.n232 756.745
R377 vdd.n225 vdd.n189 756.745
R378 vdd.n166 vdd.n130 756.745
R379 vdd.n124 vdd.n88 756.745
R380 vdd.n65 vdd.n29 756.745
R381 vdd.n2201 vdd.n2165 756.745
R382 vdd.n2260 vdd.n2224 756.745
R383 vdd.n2099 vdd.n2063 756.745
R384 vdd.n2158 vdd.n2122 756.745
R385 vdd.n1998 vdd.n1962 756.745
R386 vdd.n2057 vdd.n2021 756.745
R387 vdd.n1315 vdd.t151 640.208
R388 vdd.n1010 vdd.t192 640.208
R389 vdd.n1319 vdd.t189 640.208
R390 vdd.n1001 vdd.t214 640.208
R391 vdd.n896 vdd.t176 640.208
R392 vdd.n2823 vdd.t207 640.208
R393 vdd.n832 vdd.t169 640.208
R394 vdd.n2820 vdd.t199 640.208
R395 vdd.n799 vdd.t147 640.208
R396 vdd.n1071 vdd.t203 640.208
R397 vdd.n1772 vdd.t217 592.009
R398 vdd.n1810 vdd.t210 592.009
R399 vdd.n1706 vdd.t220 592.009
R400 vdd.n2362 vdd.t180 592.009
R401 vdd.n1248 vdd.t155 592.009
R402 vdd.n1208 vdd.t163 592.009
R403 vdd.n426 vdd.t186 592.009
R404 vdd.n440 vdd.t159 592.009
R405 vdd.n452 vdd.t166 592.009
R406 vdd.n768 vdd.t183 592.009
R407 vdd.n3456 vdd.t196 592.009
R408 vdd.n688 vdd.t172 592.009
R409 vdd.n328 vdd.n327 585
R410 vdd.n326 vdd.n293 585
R411 vdd.n325 vdd.n324 585
R412 vdd.n296 vdd.n294 585
R413 vdd.n319 vdd.n318 585
R414 vdd.n317 vdd.n316 585
R415 vdd.n300 vdd.n299 585
R416 vdd.n311 vdd.n310 585
R417 vdd.n309 vdd.n308 585
R418 vdd.n304 vdd.n303 585
R419 vdd.n269 vdd.n268 585
R420 vdd.n267 vdd.n234 585
R421 vdd.n266 vdd.n265 585
R422 vdd.n237 vdd.n235 585
R423 vdd.n260 vdd.n259 585
R424 vdd.n258 vdd.n257 585
R425 vdd.n241 vdd.n240 585
R426 vdd.n252 vdd.n251 585
R427 vdd.n250 vdd.n249 585
R428 vdd.n245 vdd.n244 585
R429 vdd.n226 vdd.n225 585
R430 vdd.n224 vdd.n191 585
R431 vdd.n223 vdd.n222 585
R432 vdd.n194 vdd.n192 585
R433 vdd.n217 vdd.n216 585
R434 vdd.n215 vdd.n214 585
R435 vdd.n198 vdd.n197 585
R436 vdd.n209 vdd.n208 585
R437 vdd.n207 vdd.n206 585
R438 vdd.n202 vdd.n201 585
R439 vdd.n167 vdd.n166 585
R440 vdd.n165 vdd.n132 585
R441 vdd.n164 vdd.n163 585
R442 vdd.n135 vdd.n133 585
R443 vdd.n158 vdd.n157 585
R444 vdd.n156 vdd.n155 585
R445 vdd.n139 vdd.n138 585
R446 vdd.n150 vdd.n149 585
R447 vdd.n148 vdd.n147 585
R448 vdd.n143 vdd.n142 585
R449 vdd.n125 vdd.n124 585
R450 vdd.n123 vdd.n90 585
R451 vdd.n122 vdd.n121 585
R452 vdd.n93 vdd.n91 585
R453 vdd.n116 vdd.n115 585
R454 vdd.n114 vdd.n113 585
R455 vdd.n97 vdd.n96 585
R456 vdd.n108 vdd.n107 585
R457 vdd.n106 vdd.n105 585
R458 vdd.n101 vdd.n100 585
R459 vdd.n66 vdd.n65 585
R460 vdd.n64 vdd.n31 585
R461 vdd.n63 vdd.n62 585
R462 vdd.n34 vdd.n32 585
R463 vdd.n57 vdd.n56 585
R464 vdd.n55 vdd.n54 585
R465 vdd.n38 vdd.n37 585
R466 vdd.n49 vdd.n48 585
R467 vdd.n47 vdd.n46 585
R468 vdd.n42 vdd.n41 585
R469 vdd.n2202 vdd.n2201 585
R470 vdd.n2200 vdd.n2167 585
R471 vdd.n2199 vdd.n2198 585
R472 vdd.n2170 vdd.n2168 585
R473 vdd.n2193 vdd.n2192 585
R474 vdd.n2191 vdd.n2190 585
R475 vdd.n2174 vdd.n2173 585
R476 vdd.n2185 vdd.n2184 585
R477 vdd.n2183 vdd.n2182 585
R478 vdd.n2178 vdd.n2177 585
R479 vdd.n2261 vdd.n2260 585
R480 vdd.n2259 vdd.n2226 585
R481 vdd.n2258 vdd.n2257 585
R482 vdd.n2229 vdd.n2227 585
R483 vdd.n2252 vdd.n2251 585
R484 vdd.n2250 vdd.n2249 585
R485 vdd.n2233 vdd.n2232 585
R486 vdd.n2244 vdd.n2243 585
R487 vdd.n2242 vdd.n2241 585
R488 vdd.n2237 vdd.n2236 585
R489 vdd.n2100 vdd.n2099 585
R490 vdd.n2098 vdd.n2065 585
R491 vdd.n2097 vdd.n2096 585
R492 vdd.n2068 vdd.n2066 585
R493 vdd.n2091 vdd.n2090 585
R494 vdd.n2089 vdd.n2088 585
R495 vdd.n2072 vdd.n2071 585
R496 vdd.n2083 vdd.n2082 585
R497 vdd.n2081 vdd.n2080 585
R498 vdd.n2076 vdd.n2075 585
R499 vdd.n2159 vdd.n2158 585
R500 vdd.n2157 vdd.n2124 585
R501 vdd.n2156 vdd.n2155 585
R502 vdd.n2127 vdd.n2125 585
R503 vdd.n2150 vdd.n2149 585
R504 vdd.n2148 vdd.n2147 585
R505 vdd.n2131 vdd.n2130 585
R506 vdd.n2142 vdd.n2141 585
R507 vdd.n2140 vdd.n2139 585
R508 vdd.n2135 vdd.n2134 585
R509 vdd.n1999 vdd.n1998 585
R510 vdd.n1997 vdd.n1964 585
R511 vdd.n1996 vdd.n1995 585
R512 vdd.n1967 vdd.n1965 585
R513 vdd.n1990 vdd.n1989 585
R514 vdd.n1988 vdd.n1987 585
R515 vdd.n1971 vdd.n1970 585
R516 vdd.n1982 vdd.n1981 585
R517 vdd.n1980 vdd.n1979 585
R518 vdd.n1975 vdd.n1974 585
R519 vdd.n2058 vdd.n2057 585
R520 vdd.n2056 vdd.n2023 585
R521 vdd.n2055 vdd.n2054 585
R522 vdd.n2026 vdd.n2024 585
R523 vdd.n2049 vdd.n2048 585
R524 vdd.n2047 vdd.n2046 585
R525 vdd.n2030 vdd.n2029 585
R526 vdd.n2041 vdd.n2040 585
R527 vdd.n2039 vdd.n2038 585
R528 vdd.n2034 vdd.n2033 585
R529 vdd.n3628 vdd.n392 509.269
R530 vdd.n3624 vdd.n393 509.269
R531 vdd.n3496 vdd.n685 509.269
R532 vdd.n3493 vdd.n684 509.269
R533 vdd.n2357 vdd.n1530 509.269
R534 vdd.n2360 vdd.n2359 509.269
R535 vdd.n1679 vdd.n1643 509.269
R536 vdd.n1875 vdd.n1644 509.269
R537 vdd.n305 vdd.t71 329.043
R538 vdd.n246 vdd.t93 329.043
R539 vdd.n203 vdd.t137 329.043
R540 vdd.n144 vdd.t145 329.043
R541 vdd.n102 vdd.t144 329.043
R542 vdd.n43 vdd.t38 329.043
R543 vdd.n2179 vdd.t304 329.043
R544 vdd.n2238 vdd.t67 329.043
R545 vdd.n2077 vdd.t58 329.043
R546 vdd.n2136 vdd.t286 329.043
R547 vdd.n1976 vdd.t12 329.043
R548 vdd.n2035 vdd.t116 329.043
R549 vdd.n1772 vdd.t219 319.788
R550 vdd.n1810 vdd.t213 319.788
R551 vdd.n1706 vdd.t222 319.788
R552 vdd.n2362 vdd.t181 319.788
R553 vdd.n1248 vdd.t157 319.788
R554 vdd.n1208 vdd.t164 319.788
R555 vdd.n426 vdd.t187 319.788
R556 vdd.n440 vdd.t161 319.788
R557 vdd.n452 vdd.t167 319.788
R558 vdd.n768 vdd.t185 319.788
R559 vdd.n3456 vdd.t198 319.788
R560 vdd.n688 vdd.t175 319.788
R561 vdd.n1773 vdd.t218 303.69
R562 vdd.n1811 vdd.t212 303.69
R563 vdd.n1707 vdd.t221 303.69
R564 vdd.n2363 vdd.t182 303.69
R565 vdd.n1249 vdd.t158 303.69
R566 vdd.n1209 vdd.t165 303.69
R567 vdd.n427 vdd.t188 303.69
R568 vdd.n441 vdd.t162 303.69
R569 vdd.n453 vdd.t168 303.69
R570 vdd.n769 vdd.t184 303.69
R571 vdd.n3457 vdd.t197 303.69
R572 vdd.n689 vdd.t174 303.69
R573 vdd.n3090 vdd.n960 279.512
R574 vdd.n3330 vdd.n809 279.512
R575 vdd.n3267 vdd.n806 279.512
R576 vdd.n3022 vdd.n3021 279.512
R577 vdd.n2783 vdd.n998 279.512
R578 vdd.n2714 vdd.n2713 279.512
R579 vdd.n1355 vdd.n1354 279.512
R580 vdd.n2508 vdd.n1138 279.512
R581 vdd.n3246 vdd.n807 279.512
R582 vdd.n3333 vdd.n3332 279.512
R583 vdd.n2895 vdd.n2818 279.512
R584 vdd.n2826 vdd.n956 279.512
R585 vdd.n2711 vdd.n1008 279.512
R586 vdd.n1006 vdd.n980 279.512
R587 vdd.n1480 vdd.n1175 279.512
R588 vdd.n1280 vdd.n1133 279.512
R589 vdd.n2506 vdd.n1141 254.619
R590 vdd.n3495 vdd.n692 254.619
R591 vdd.n3248 vdd.n807 185
R592 vdd.n3331 vdd.n807 185
R593 vdd.n3250 vdd.n3249 185
R594 vdd.n3249 vdd.n805 185
R595 vdd.n3251 vdd.n839 185
R596 vdd.n3261 vdd.n839 185
R597 vdd.n3252 vdd.n848 185
R598 vdd.n848 vdd.n846 185
R599 vdd.n3254 vdd.n3253 185
R600 vdd.n3255 vdd.n3254 185
R601 vdd.n3207 vdd.n847 185
R602 vdd.n847 vdd.n843 185
R603 vdd.n3206 vdd.n3205 185
R604 vdd.n3205 vdd.n3204 185
R605 vdd.n850 vdd.n849 185
R606 vdd.n851 vdd.n850 185
R607 vdd.n3197 vdd.n3196 185
R608 vdd.n3198 vdd.n3197 185
R609 vdd.n3195 vdd.n859 185
R610 vdd.n864 vdd.n859 185
R611 vdd.n3194 vdd.n3193 185
R612 vdd.n3193 vdd.n3192 185
R613 vdd.n861 vdd.n860 185
R614 vdd.n870 vdd.n861 185
R615 vdd.n3185 vdd.n3184 185
R616 vdd.n3186 vdd.n3185 185
R617 vdd.n3183 vdd.n871 185
R618 vdd.n877 vdd.n871 185
R619 vdd.n3182 vdd.n3181 185
R620 vdd.n3181 vdd.n3180 185
R621 vdd.n873 vdd.n872 185
R622 vdd.n874 vdd.n873 185
R623 vdd.n3173 vdd.n3172 185
R624 vdd.n3174 vdd.n3173 185
R625 vdd.n3171 vdd.n884 185
R626 vdd.n884 vdd.n881 185
R627 vdd.n3170 vdd.n3169 185
R628 vdd.n3169 vdd.n3168 185
R629 vdd.n886 vdd.n885 185
R630 vdd.n887 vdd.n886 185
R631 vdd.n3161 vdd.n3160 185
R632 vdd.n3162 vdd.n3161 185
R633 vdd.n3159 vdd.n895 185
R634 vdd.n901 vdd.n895 185
R635 vdd.n3158 vdd.n3157 185
R636 vdd.n3157 vdd.n3156 185
R637 vdd.n3147 vdd.n898 185
R638 vdd.n908 vdd.n898 185
R639 vdd.n3149 vdd.n3148 185
R640 vdd.n3150 vdd.n3149 185
R641 vdd.n3146 vdd.n909 185
R642 vdd.n909 vdd.n905 185
R643 vdd.n3145 vdd.n3144 185
R644 vdd.n3144 vdd.n3143 185
R645 vdd.n911 vdd.n910 185
R646 vdd.n912 vdd.n911 185
R647 vdd.n3136 vdd.n3135 185
R648 vdd.n3137 vdd.n3136 185
R649 vdd.n3134 vdd.n920 185
R650 vdd.n925 vdd.n920 185
R651 vdd.n3133 vdd.n3132 185
R652 vdd.n3132 vdd.n3131 185
R653 vdd.n922 vdd.n921 185
R654 vdd.n931 vdd.n922 185
R655 vdd.n3124 vdd.n3123 185
R656 vdd.n3125 vdd.n3124 185
R657 vdd.n3122 vdd.n932 185
R658 vdd.n2998 vdd.n932 185
R659 vdd.n3121 vdd.n3120 185
R660 vdd.n3120 vdd.n3119 185
R661 vdd.n934 vdd.n933 185
R662 vdd.n3004 vdd.n934 185
R663 vdd.n3112 vdd.n3111 185
R664 vdd.n3113 vdd.n3112 185
R665 vdd.n3110 vdd.n943 185
R666 vdd.n943 vdd.n940 185
R667 vdd.n3109 vdd.n3108 185
R668 vdd.n3108 vdd.n3107 185
R669 vdd.n945 vdd.n944 185
R670 vdd.n946 vdd.n945 185
R671 vdd.n3100 vdd.n3099 185
R672 vdd.n3101 vdd.n3100 185
R673 vdd.n3098 vdd.n954 185
R674 vdd.n3016 vdd.n954 185
R675 vdd.n3097 vdd.n3096 185
R676 vdd.n3096 vdd.n3095 185
R677 vdd.n956 vdd.n955 185
R678 vdd.n957 vdd.n956 185
R679 vdd.n2827 vdd.n2826 185
R680 vdd.n2829 vdd.n2828 185
R681 vdd.n2831 vdd.n2830 185
R682 vdd.n2833 vdd.n2832 185
R683 vdd.n2835 vdd.n2834 185
R684 vdd.n2837 vdd.n2836 185
R685 vdd.n2839 vdd.n2838 185
R686 vdd.n2841 vdd.n2840 185
R687 vdd.n2843 vdd.n2842 185
R688 vdd.n2845 vdd.n2844 185
R689 vdd.n2847 vdd.n2846 185
R690 vdd.n2849 vdd.n2848 185
R691 vdd.n2851 vdd.n2850 185
R692 vdd.n2853 vdd.n2852 185
R693 vdd.n2855 vdd.n2854 185
R694 vdd.n2857 vdd.n2856 185
R695 vdd.n2859 vdd.n2858 185
R696 vdd.n2861 vdd.n2860 185
R697 vdd.n2863 vdd.n2862 185
R698 vdd.n2865 vdd.n2864 185
R699 vdd.n2867 vdd.n2866 185
R700 vdd.n2869 vdd.n2868 185
R701 vdd.n2871 vdd.n2870 185
R702 vdd.n2873 vdd.n2872 185
R703 vdd.n2875 vdd.n2874 185
R704 vdd.n2877 vdd.n2876 185
R705 vdd.n2879 vdd.n2878 185
R706 vdd.n2881 vdd.n2880 185
R707 vdd.n2883 vdd.n2882 185
R708 vdd.n2885 vdd.n2884 185
R709 vdd.n2887 vdd.n2886 185
R710 vdd.n2889 vdd.n2888 185
R711 vdd.n2891 vdd.n2890 185
R712 vdd.n2893 vdd.n2892 185
R713 vdd.n2894 vdd.n2818 185
R714 vdd.n3088 vdd.n2818 185
R715 vdd.n3334 vdd.n3333 185
R716 vdd.n3335 vdd.n798 185
R717 vdd.n3337 vdd.n3336 185
R718 vdd.n3339 vdd.n796 185
R719 vdd.n3341 vdd.n3340 185
R720 vdd.n3342 vdd.n795 185
R721 vdd.n3344 vdd.n3343 185
R722 vdd.n3346 vdd.n793 185
R723 vdd.n3348 vdd.n3347 185
R724 vdd.n3349 vdd.n792 185
R725 vdd.n3351 vdd.n3350 185
R726 vdd.n3353 vdd.n790 185
R727 vdd.n3355 vdd.n3354 185
R728 vdd.n3356 vdd.n789 185
R729 vdd.n3358 vdd.n3357 185
R730 vdd.n3360 vdd.n788 185
R731 vdd.n3361 vdd.n786 185
R732 vdd.n3364 vdd.n3363 185
R733 vdd.n787 vdd.n785 185
R734 vdd.n3220 vdd.n3219 185
R735 vdd.n3222 vdd.n3221 185
R736 vdd.n3224 vdd.n3216 185
R737 vdd.n3226 vdd.n3225 185
R738 vdd.n3227 vdd.n3215 185
R739 vdd.n3229 vdd.n3228 185
R740 vdd.n3231 vdd.n3213 185
R741 vdd.n3233 vdd.n3232 185
R742 vdd.n3234 vdd.n3212 185
R743 vdd.n3236 vdd.n3235 185
R744 vdd.n3238 vdd.n3210 185
R745 vdd.n3240 vdd.n3239 185
R746 vdd.n3241 vdd.n3209 185
R747 vdd.n3243 vdd.n3242 185
R748 vdd.n3245 vdd.n3208 185
R749 vdd.n3247 vdd.n3246 185
R750 vdd.n3246 vdd.n692 185
R751 vdd.n3332 vdd.n802 185
R752 vdd.n3332 vdd.n3331 185
R753 vdd.n2949 vdd.n804 185
R754 vdd.n805 vdd.n804 185
R755 vdd.n2950 vdd.n838 185
R756 vdd.n3261 vdd.n838 185
R757 vdd.n2952 vdd.n2951 185
R758 vdd.n2951 vdd.n846 185
R759 vdd.n2953 vdd.n845 185
R760 vdd.n3255 vdd.n845 185
R761 vdd.n2955 vdd.n2954 185
R762 vdd.n2954 vdd.n843 185
R763 vdd.n2956 vdd.n853 185
R764 vdd.n3204 vdd.n853 185
R765 vdd.n2958 vdd.n2957 185
R766 vdd.n2957 vdd.n851 185
R767 vdd.n2959 vdd.n858 185
R768 vdd.n3198 vdd.n858 185
R769 vdd.n2961 vdd.n2960 185
R770 vdd.n2960 vdd.n864 185
R771 vdd.n2962 vdd.n863 185
R772 vdd.n3192 vdd.n863 185
R773 vdd.n2964 vdd.n2963 185
R774 vdd.n2963 vdd.n870 185
R775 vdd.n2965 vdd.n869 185
R776 vdd.n3186 vdd.n869 185
R777 vdd.n2967 vdd.n2966 185
R778 vdd.n2966 vdd.n877 185
R779 vdd.n2968 vdd.n876 185
R780 vdd.n3180 vdd.n876 185
R781 vdd.n2970 vdd.n2969 185
R782 vdd.n2969 vdd.n874 185
R783 vdd.n2971 vdd.n883 185
R784 vdd.n3174 vdd.n883 185
R785 vdd.n2973 vdd.n2972 185
R786 vdd.n2972 vdd.n881 185
R787 vdd.n2974 vdd.n889 185
R788 vdd.n3168 vdd.n889 185
R789 vdd.n2976 vdd.n2975 185
R790 vdd.n2975 vdd.n887 185
R791 vdd.n2977 vdd.n894 185
R792 vdd.n3162 vdd.n894 185
R793 vdd.n2979 vdd.n2978 185
R794 vdd.n2978 vdd.n901 185
R795 vdd.n2980 vdd.n900 185
R796 vdd.n3156 vdd.n900 185
R797 vdd.n2982 vdd.n2981 185
R798 vdd.n2981 vdd.n908 185
R799 vdd.n2983 vdd.n907 185
R800 vdd.n3150 vdd.n907 185
R801 vdd.n2985 vdd.n2984 185
R802 vdd.n2984 vdd.n905 185
R803 vdd.n2986 vdd.n914 185
R804 vdd.n3143 vdd.n914 185
R805 vdd.n2988 vdd.n2987 185
R806 vdd.n2987 vdd.n912 185
R807 vdd.n2989 vdd.n919 185
R808 vdd.n3137 vdd.n919 185
R809 vdd.n2991 vdd.n2990 185
R810 vdd.n2990 vdd.n925 185
R811 vdd.n2992 vdd.n924 185
R812 vdd.n3131 vdd.n924 185
R813 vdd.n2994 vdd.n2993 185
R814 vdd.n2993 vdd.n931 185
R815 vdd.n2995 vdd.n930 185
R816 vdd.n3125 vdd.n930 185
R817 vdd.n2997 vdd.n2996 185
R818 vdd.n2998 vdd.n2997 185
R819 vdd.n2898 vdd.n936 185
R820 vdd.n3119 vdd.n936 185
R821 vdd.n3006 vdd.n3005 185
R822 vdd.n3005 vdd.n3004 185
R823 vdd.n3007 vdd.n942 185
R824 vdd.n3113 vdd.n942 185
R825 vdd.n3009 vdd.n3008 185
R826 vdd.n3008 vdd.n940 185
R827 vdd.n3010 vdd.n948 185
R828 vdd.n3107 vdd.n948 185
R829 vdd.n3012 vdd.n3011 185
R830 vdd.n3011 vdd.n946 185
R831 vdd.n3013 vdd.n953 185
R832 vdd.n3101 vdd.n953 185
R833 vdd.n3015 vdd.n3014 185
R834 vdd.n3016 vdd.n3015 185
R835 vdd.n2897 vdd.n959 185
R836 vdd.n3095 vdd.n959 185
R837 vdd.n2896 vdd.n2895 185
R838 vdd.n2895 vdd.n957 185
R839 vdd.n2357 vdd.n2356 185
R840 vdd.n2358 vdd.n2357 185
R841 vdd.n1531 vdd.n1529 185
R842 vdd.n2349 vdd.n1529 185
R843 vdd.n2352 vdd.n2351 185
R844 vdd.n2351 vdd.n2350 185
R845 vdd.n1534 vdd.n1533 185
R846 vdd.n1535 vdd.n1534 185
R847 vdd.n2338 vdd.n2337 185
R848 vdd.n2339 vdd.n2338 185
R849 vdd.n1543 vdd.n1542 185
R850 vdd.n2330 vdd.n1542 185
R851 vdd.n2333 vdd.n2332 185
R852 vdd.n2332 vdd.n2331 185
R853 vdd.n1546 vdd.n1545 185
R854 vdd.n1553 vdd.n1546 185
R855 vdd.n2321 vdd.n2320 185
R856 vdd.n2322 vdd.n2321 185
R857 vdd.n1555 vdd.n1554 185
R858 vdd.n1554 vdd.n1552 185
R859 vdd.n2316 vdd.n2315 185
R860 vdd.n2315 vdd.n2314 185
R861 vdd.n1558 vdd.n1557 185
R862 vdd.n1559 vdd.n1558 185
R863 vdd.n2305 vdd.n2304 185
R864 vdd.n2306 vdd.n2305 185
R865 vdd.n1566 vdd.n1565 185
R866 vdd.n2297 vdd.n1565 185
R867 vdd.n2300 vdd.n2299 185
R868 vdd.n2299 vdd.n2298 185
R869 vdd.n1569 vdd.n1568 185
R870 vdd.n1575 vdd.n1569 185
R871 vdd.n2288 vdd.n2287 185
R872 vdd.n2289 vdd.n2288 185
R873 vdd.n1577 vdd.n1576 185
R874 vdd.n2280 vdd.n1576 185
R875 vdd.n2283 vdd.n2282 185
R876 vdd.n2282 vdd.n2281 185
R877 vdd.n1580 vdd.n1579 185
R878 vdd.n1581 vdd.n1580 185
R879 vdd.n2271 vdd.n2270 185
R880 vdd.n2272 vdd.n2271 185
R881 vdd.n1589 vdd.n1588 185
R882 vdd.n1588 vdd.n1587 185
R883 vdd.n1959 vdd.n1958 185
R884 vdd.n1958 vdd.n1957 185
R885 vdd.n1592 vdd.n1591 185
R886 vdd.n1598 vdd.n1592 185
R887 vdd.n1948 vdd.n1947 185
R888 vdd.n1949 vdd.n1948 185
R889 vdd.n1600 vdd.n1599 185
R890 vdd.n1940 vdd.n1599 185
R891 vdd.n1943 vdd.n1942 185
R892 vdd.n1942 vdd.n1941 185
R893 vdd.n1603 vdd.n1602 185
R894 vdd.n1610 vdd.n1603 185
R895 vdd.n1931 vdd.n1930 185
R896 vdd.n1932 vdd.n1931 185
R897 vdd.n1612 vdd.n1611 185
R898 vdd.n1611 vdd.n1609 185
R899 vdd.n1926 vdd.n1925 185
R900 vdd.n1925 vdd.n1924 185
R901 vdd.n1615 vdd.n1614 185
R902 vdd.n1616 vdd.n1615 185
R903 vdd.n1915 vdd.n1914 185
R904 vdd.n1916 vdd.n1915 185
R905 vdd.n1623 vdd.n1622 185
R906 vdd.n1907 vdd.n1622 185
R907 vdd.n1910 vdd.n1909 185
R908 vdd.n1909 vdd.n1908 185
R909 vdd.n1626 vdd.n1625 185
R910 vdd.n1632 vdd.n1626 185
R911 vdd.n1898 vdd.n1897 185
R912 vdd.n1899 vdd.n1898 185
R913 vdd.n1634 vdd.n1633 185
R914 vdd.n1890 vdd.n1633 185
R915 vdd.n1893 vdd.n1892 185
R916 vdd.n1892 vdd.n1891 185
R917 vdd.n1637 vdd.n1636 185
R918 vdd.n1638 vdd.n1637 185
R919 vdd.n1881 vdd.n1880 185
R920 vdd.n1882 vdd.n1881 185
R921 vdd.n1645 vdd.n1644 185
R922 vdd.n1680 vdd.n1644 185
R923 vdd.n1876 vdd.n1875 185
R924 vdd.n1648 vdd.n1647 185
R925 vdd.n1872 vdd.n1871 185
R926 vdd.n1873 vdd.n1872 185
R927 vdd.n1682 vdd.n1681 185
R928 vdd.n1867 vdd.n1684 185
R929 vdd.n1866 vdd.n1685 185
R930 vdd.n1865 vdd.n1686 185
R931 vdd.n1688 vdd.n1687 185
R932 vdd.n1861 vdd.n1690 185
R933 vdd.n1860 vdd.n1691 185
R934 vdd.n1859 vdd.n1692 185
R935 vdd.n1694 vdd.n1693 185
R936 vdd.n1855 vdd.n1696 185
R937 vdd.n1854 vdd.n1697 185
R938 vdd.n1853 vdd.n1698 185
R939 vdd.n1700 vdd.n1699 185
R940 vdd.n1849 vdd.n1702 185
R941 vdd.n1848 vdd.n1703 185
R942 vdd.n1847 vdd.n1704 185
R943 vdd.n1708 vdd.n1705 185
R944 vdd.n1843 vdd.n1710 185
R945 vdd.n1842 vdd.n1711 185
R946 vdd.n1841 vdd.n1712 185
R947 vdd.n1714 vdd.n1713 185
R948 vdd.n1837 vdd.n1716 185
R949 vdd.n1836 vdd.n1717 185
R950 vdd.n1835 vdd.n1718 185
R951 vdd.n1720 vdd.n1719 185
R952 vdd.n1831 vdd.n1722 185
R953 vdd.n1830 vdd.n1723 185
R954 vdd.n1829 vdd.n1724 185
R955 vdd.n1726 vdd.n1725 185
R956 vdd.n1825 vdd.n1728 185
R957 vdd.n1824 vdd.n1729 185
R958 vdd.n1823 vdd.n1730 185
R959 vdd.n1732 vdd.n1731 185
R960 vdd.n1819 vdd.n1734 185
R961 vdd.n1818 vdd.n1735 185
R962 vdd.n1817 vdd.n1736 185
R963 vdd.n1738 vdd.n1737 185
R964 vdd.n1813 vdd.n1740 185
R965 vdd.n1812 vdd.n1809 185
R966 vdd.n1808 vdd.n1741 185
R967 vdd.n1743 vdd.n1742 185
R968 vdd.n1804 vdd.n1745 185
R969 vdd.n1803 vdd.n1746 185
R970 vdd.n1802 vdd.n1747 185
R971 vdd.n1749 vdd.n1748 185
R972 vdd.n1798 vdd.n1751 185
R973 vdd.n1797 vdd.n1752 185
R974 vdd.n1796 vdd.n1753 185
R975 vdd.n1755 vdd.n1754 185
R976 vdd.n1792 vdd.n1757 185
R977 vdd.n1791 vdd.n1758 185
R978 vdd.n1790 vdd.n1759 185
R979 vdd.n1761 vdd.n1760 185
R980 vdd.n1786 vdd.n1763 185
R981 vdd.n1785 vdd.n1764 185
R982 vdd.n1784 vdd.n1765 185
R983 vdd.n1767 vdd.n1766 185
R984 vdd.n1780 vdd.n1769 185
R985 vdd.n1779 vdd.n1770 185
R986 vdd.n1778 vdd.n1771 185
R987 vdd.n1775 vdd.n1679 185
R988 vdd.n1873 vdd.n1679 185
R989 vdd.n2361 vdd.n2360 185
R990 vdd.n2365 vdd.n1525 185
R991 vdd.n1524 vdd.n1518 185
R992 vdd.n1522 vdd.n1521 185
R993 vdd.n1520 vdd.n1279 185
R994 vdd.n2369 vdd.n1276 185
R995 vdd.n2371 vdd.n2370 185
R996 vdd.n2373 vdd.n1274 185
R997 vdd.n2375 vdd.n2374 185
R998 vdd.n2376 vdd.n1269 185
R999 vdd.n2378 vdd.n2377 185
R1000 vdd.n2380 vdd.n1267 185
R1001 vdd.n2382 vdd.n2381 185
R1002 vdd.n2383 vdd.n1262 185
R1003 vdd.n2385 vdd.n2384 185
R1004 vdd.n2387 vdd.n1260 185
R1005 vdd.n2389 vdd.n2388 185
R1006 vdd.n2390 vdd.n1256 185
R1007 vdd.n2392 vdd.n2391 185
R1008 vdd.n2394 vdd.n1253 185
R1009 vdd.n2396 vdd.n2395 185
R1010 vdd.n1254 vdd.n1247 185
R1011 vdd.n2400 vdd.n1251 185
R1012 vdd.n2401 vdd.n1243 185
R1013 vdd.n2403 vdd.n2402 185
R1014 vdd.n2405 vdd.n1241 185
R1015 vdd.n2407 vdd.n2406 185
R1016 vdd.n2408 vdd.n1236 185
R1017 vdd.n2410 vdd.n2409 185
R1018 vdd.n2412 vdd.n1234 185
R1019 vdd.n2414 vdd.n2413 185
R1020 vdd.n2415 vdd.n1229 185
R1021 vdd.n2417 vdd.n2416 185
R1022 vdd.n2419 vdd.n1227 185
R1023 vdd.n2421 vdd.n2420 185
R1024 vdd.n2422 vdd.n1222 185
R1025 vdd.n2424 vdd.n2423 185
R1026 vdd.n2426 vdd.n1220 185
R1027 vdd.n2428 vdd.n2427 185
R1028 vdd.n2429 vdd.n1216 185
R1029 vdd.n2431 vdd.n2430 185
R1030 vdd.n2433 vdd.n1213 185
R1031 vdd.n2435 vdd.n2434 185
R1032 vdd.n1214 vdd.n1207 185
R1033 vdd.n2439 vdd.n1211 185
R1034 vdd.n2440 vdd.n1203 185
R1035 vdd.n2442 vdd.n2441 185
R1036 vdd.n2444 vdd.n1201 185
R1037 vdd.n2446 vdd.n2445 185
R1038 vdd.n2447 vdd.n1196 185
R1039 vdd.n2449 vdd.n2448 185
R1040 vdd.n2451 vdd.n1194 185
R1041 vdd.n2453 vdd.n2452 185
R1042 vdd.n2454 vdd.n1189 185
R1043 vdd.n2456 vdd.n2455 185
R1044 vdd.n2458 vdd.n1187 185
R1045 vdd.n2460 vdd.n2459 185
R1046 vdd.n2461 vdd.n1185 185
R1047 vdd.n2463 vdd.n2462 185
R1048 vdd.n2466 vdd.n2465 185
R1049 vdd.n2468 vdd.n2467 185
R1050 vdd.n2470 vdd.n1183 185
R1051 vdd.n2472 vdd.n2471 185
R1052 vdd.n1530 vdd.n1182 185
R1053 vdd.n2359 vdd.n1528 185
R1054 vdd.n2359 vdd.n2358 185
R1055 vdd.n1538 vdd.n1527 185
R1056 vdd.n2349 vdd.n1527 185
R1057 vdd.n2348 vdd.n2347 185
R1058 vdd.n2350 vdd.n2348 185
R1059 vdd.n1537 vdd.n1536 185
R1060 vdd.n1536 vdd.n1535 185
R1061 vdd.n2341 vdd.n2340 185
R1062 vdd.n2340 vdd.n2339 185
R1063 vdd.n1541 vdd.n1540 185
R1064 vdd.n2330 vdd.n1541 185
R1065 vdd.n2329 vdd.n2328 185
R1066 vdd.n2331 vdd.n2329 185
R1067 vdd.n1548 vdd.n1547 185
R1068 vdd.n1553 vdd.n1547 185
R1069 vdd.n2324 vdd.n2323 185
R1070 vdd.n2323 vdd.n2322 185
R1071 vdd.n1551 vdd.n1550 185
R1072 vdd.n1552 vdd.n1551 185
R1073 vdd.n2313 vdd.n2312 185
R1074 vdd.n2314 vdd.n2313 185
R1075 vdd.n1561 vdd.n1560 185
R1076 vdd.n1560 vdd.n1559 185
R1077 vdd.n2308 vdd.n2307 185
R1078 vdd.n2307 vdd.n2306 185
R1079 vdd.n1564 vdd.n1563 185
R1080 vdd.n2297 vdd.n1564 185
R1081 vdd.n2296 vdd.n2295 185
R1082 vdd.n2298 vdd.n2296 185
R1083 vdd.n1571 vdd.n1570 185
R1084 vdd.n1575 vdd.n1570 185
R1085 vdd.n2291 vdd.n2290 185
R1086 vdd.n2290 vdd.n2289 185
R1087 vdd.n1574 vdd.n1573 185
R1088 vdd.n2280 vdd.n1574 185
R1089 vdd.n2279 vdd.n2278 185
R1090 vdd.n2281 vdd.n2279 185
R1091 vdd.n1583 vdd.n1582 185
R1092 vdd.n1582 vdd.n1581 185
R1093 vdd.n2274 vdd.n2273 185
R1094 vdd.n2273 vdd.n2272 185
R1095 vdd.n1586 vdd.n1585 185
R1096 vdd.n1587 vdd.n1586 185
R1097 vdd.n1956 vdd.n1955 185
R1098 vdd.n1957 vdd.n1956 185
R1099 vdd.n1594 vdd.n1593 185
R1100 vdd.n1598 vdd.n1593 185
R1101 vdd.n1951 vdd.n1950 185
R1102 vdd.n1950 vdd.n1949 185
R1103 vdd.n1597 vdd.n1596 185
R1104 vdd.n1940 vdd.n1597 185
R1105 vdd.n1939 vdd.n1938 185
R1106 vdd.n1941 vdd.n1939 185
R1107 vdd.n1605 vdd.n1604 185
R1108 vdd.n1610 vdd.n1604 185
R1109 vdd.n1934 vdd.n1933 185
R1110 vdd.n1933 vdd.n1932 185
R1111 vdd.n1608 vdd.n1607 185
R1112 vdd.n1609 vdd.n1608 185
R1113 vdd.n1923 vdd.n1922 185
R1114 vdd.n1924 vdd.n1923 185
R1115 vdd.n1618 vdd.n1617 185
R1116 vdd.n1617 vdd.n1616 185
R1117 vdd.n1918 vdd.n1917 185
R1118 vdd.n1917 vdd.n1916 185
R1119 vdd.n1621 vdd.n1620 185
R1120 vdd.n1907 vdd.n1621 185
R1121 vdd.n1906 vdd.n1905 185
R1122 vdd.n1908 vdd.n1906 185
R1123 vdd.n1628 vdd.n1627 185
R1124 vdd.n1632 vdd.n1627 185
R1125 vdd.n1901 vdd.n1900 185
R1126 vdd.n1900 vdd.n1899 185
R1127 vdd.n1631 vdd.n1630 185
R1128 vdd.n1890 vdd.n1631 185
R1129 vdd.n1889 vdd.n1888 185
R1130 vdd.n1891 vdd.n1889 185
R1131 vdd.n1640 vdd.n1639 185
R1132 vdd.n1639 vdd.n1638 185
R1133 vdd.n1884 vdd.n1883 185
R1134 vdd.n1883 vdd.n1882 185
R1135 vdd.n1643 vdd.n1642 185
R1136 vdd.n1680 vdd.n1643 185
R1137 vdd.n1000 vdd.n998 185
R1138 vdd.n2712 vdd.n998 185
R1139 vdd.n2634 vdd.n1018 185
R1140 vdd.n1018 vdd.n1005 185
R1141 vdd.n2636 vdd.n2635 185
R1142 vdd.n2637 vdd.n2636 185
R1143 vdd.n2633 vdd.n1017 185
R1144 vdd.n1399 vdd.n1017 185
R1145 vdd.n2632 vdd.n2631 185
R1146 vdd.n2631 vdd.n2630 185
R1147 vdd.n1020 vdd.n1019 185
R1148 vdd.n1021 vdd.n1020 185
R1149 vdd.n2621 vdd.n2620 185
R1150 vdd.n2622 vdd.n2621 185
R1151 vdd.n2619 vdd.n1031 185
R1152 vdd.n1031 vdd.n1028 185
R1153 vdd.n2618 vdd.n2617 185
R1154 vdd.n2617 vdd.n2616 185
R1155 vdd.n1033 vdd.n1032 185
R1156 vdd.n1425 vdd.n1033 185
R1157 vdd.n2609 vdd.n2608 185
R1158 vdd.n2610 vdd.n2609 185
R1159 vdd.n2607 vdd.n1041 185
R1160 vdd.n1046 vdd.n1041 185
R1161 vdd.n2606 vdd.n2605 185
R1162 vdd.n2605 vdd.n2604 185
R1163 vdd.n1043 vdd.n1042 185
R1164 vdd.n1052 vdd.n1043 185
R1165 vdd.n2597 vdd.n2596 185
R1166 vdd.n2598 vdd.n2597 185
R1167 vdd.n2595 vdd.n1053 185
R1168 vdd.n1437 vdd.n1053 185
R1169 vdd.n2594 vdd.n2593 185
R1170 vdd.n2593 vdd.n2592 185
R1171 vdd.n1055 vdd.n1054 185
R1172 vdd.n1056 vdd.n1055 185
R1173 vdd.n2585 vdd.n2584 185
R1174 vdd.n2586 vdd.n2585 185
R1175 vdd.n2583 vdd.n1065 185
R1176 vdd.n1065 vdd.n1062 185
R1177 vdd.n2582 vdd.n2581 185
R1178 vdd.n2581 vdd.n2580 185
R1179 vdd.n1067 vdd.n1066 185
R1180 vdd.n1076 vdd.n1067 185
R1181 vdd.n2572 vdd.n2571 185
R1182 vdd.n2573 vdd.n2572 185
R1183 vdd.n2570 vdd.n1077 185
R1184 vdd.n1083 vdd.n1077 185
R1185 vdd.n2569 vdd.n2568 185
R1186 vdd.n2568 vdd.n2567 185
R1187 vdd.n1079 vdd.n1078 185
R1188 vdd.n1080 vdd.n1079 185
R1189 vdd.n2560 vdd.n2559 185
R1190 vdd.n2561 vdd.n2560 185
R1191 vdd.n2558 vdd.n1090 185
R1192 vdd.n1090 vdd.n1087 185
R1193 vdd.n2557 vdd.n2556 185
R1194 vdd.n2556 vdd.n2555 185
R1195 vdd.n1092 vdd.n1091 185
R1196 vdd.n1093 vdd.n1092 185
R1197 vdd.n2548 vdd.n2547 185
R1198 vdd.n2549 vdd.n2548 185
R1199 vdd.n2546 vdd.n1101 185
R1200 vdd.n1106 vdd.n1101 185
R1201 vdd.n2545 vdd.n2544 185
R1202 vdd.n2544 vdd.n2543 185
R1203 vdd.n1103 vdd.n1102 185
R1204 vdd.n1112 vdd.n1103 185
R1205 vdd.n2536 vdd.n2535 185
R1206 vdd.n2537 vdd.n2536 185
R1207 vdd.n2534 vdd.n1113 185
R1208 vdd.n1119 vdd.n1113 185
R1209 vdd.n2533 vdd.n2532 185
R1210 vdd.n2532 vdd.n2531 185
R1211 vdd.n1115 vdd.n1114 185
R1212 vdd.n1116 vdd.n1115 185
R1213 vdd.n2524 vdd.n2523 185
R1214 vdd.n2525 vdd.n2524 185
R1215 vdd.n2522 vdd.n1126 185
R1216 vdd.n1126 vdd.n1123 185
R1217 vdd.n2521 vdd.n2520 185
R1218 vdd.n2520 vdd.n2519 185
R1219 vdd.n1128 vdd.n1127 185
R1220 vdd.n1137 vdd.n1128 185
R1221 vdd.n2512 vdd.n2511 185
R1222 vdd.n2513 vdd.n2512 185
R1223 vdd.n2510 vdd.n1138 185
R1224 vdd.n1138 vdd.n1134 185
R1225 vdd.n2509 vdd.n2508 185
R1226 vdd.n1140 vdd.n1139 185
R1227 vdd.n2505 vdd.n2504 185
R1228 vdd.n2506 vdd.n2505 185
R1229 vdd.n2503 vdd.n1176 185
R1230 vdd.n2502 vdd.n2501 185
R1231 vdd.n2500 vdd.n2499 185
R1232 vdd.n2498 vdd.n2497 185
R1233 vdd.n2496 vdd.n2495 185
R1234 vdd.n2494 vdd.n2493 185
R1235 vdd.n2492 vdd.n2491 185
R1236 vdd.n2490 vdd.n2489 185
R1237 vdd.n2488 vdd.n2487 185
R1238 vdd.n2486 vdd.n2485 185
R1239 vdd.n2484 vdd.n2483 185
R1240 vdd.n2482 vdd.n2481 185
R1241 vdd.n2480 vdd.n2479 185
R1242 vdd.n2478 vdd.n2477 185
R1243 vdd.n2476 vdd.n2475 185
R1244 vdd.n1321 vdd.n1177 185
R1245 vdd.n1323 vdd.n1322 185
R1246 vdd.n1325 vdd.n1324 185
R1247 vdd.n1327 vdd.n1326 185
R1248 vdd.n1329 vdd.n1328 185
R1249 vdd.n1331 vdd.n1330 185
R1250 vdd.n1333 vdd.n1332 185
R1251 vdd.n1335 vdd.n1334 185
R1252 vdd.n1337 vdd.n1336 185
R1253 vdd.n1339 vdd.n1338 185
R1254 vdd.n1341 vdd.n1340 185
R1255 vdd.n1343 vdd.n1342 185
R1256 vdd.n1345 vdd.n1344 185
R1257 vdd.n1347 vdd.n1346 185
R1258 vdd.n1350 vdd.n1349 185
R1259 vdd.n1352 vdd.n1351 185
R1260 vdd.n1354 vdd.n1353 185
R1261 vdd.n2715 vdd.n2714 185
R1262 vdd.n2717 vdd.n2716 185
R1263 vdd.n2719 vdd.n2718 185
R1264 vdd.n2722 vdd.n2721 185
R1265 vdd.n2724 vdd.n2723 185
R1266 vdd.n2726 vdd.n2725 185
R1267 vdd.n2728 vdd.n2727 185
R1268 vdd.n2730 vdd.n2729 185
R1269 vdd.n2732 vdd.n2731 185
R1270 vdd.n2734 vdd.n2733 185
R1271 vdd.n2736 vdd.n2735 185
R1272 vdd.n2738 vdd.n2737 185
R1273 vdd.n2740 vdd.n2739 185
R1274 vdd.n2742 vdd.n2741 185
R1275 vdd.n2744 vdd.n2743 185
R1276 vdd.n2746 vdd.n2745 185
R1277 vdd.n2748 vdd.n2747 185
R1278 vdd.n2750 vdd.n2749 185
R1279 vdd.n2752 vdd.n2751 185
R1280 vdd.n2754 vdd.n2753 185
R1281 vdd.n2756 vdd.n2755 185
R1282 vdd.n2758 vdd.n2757 185
R1283 vdd.n2760 vdd.n2759 185
R1284 vdd.n2762 vdd.n2761 185
R1285 vdd.n2764 vdd.n2763 185
R1286 vdd.n2766 vdd.n2765 185
R1287 vdd.n2768 vdd.n2767 185
R1288 vdd.n2770 vdd.n2769 185
R1289 vdd.n2772 vdd.n2771 185
R1290 vdd.n2774 vdd.n2773 185
R1291 vdd.n2776 vdd.n2775 185
R1292 vdd.n2778 vdd.n2777 185
R1293 vdd.n2780 vdd.n2779 185
R1294 vdd.n2781 vdd.n999 185
R1295 vdd.n2783 vdd.n2782 185
R1296 vdd.n2784 vdd.n2783 185
R1297 vdd.n2713 vdd.n1003 185
R1298 vdd.n2713 vdd.n2712 185
R1299 vdd.n1397 vdd.n1004 185
R1300 vdd.n1005 vdd.n1004 185
R1301 vdd.n1398 vdd.n1015 185
R1302 vdd.n2637 vdd.n1015 185
R1303 vdd.n1401 vdd.n1400 185
R1304 vdd.n1400 vdd.n1399 185
R1305 vdd.n1402 vdd.n1022 185
R1306 vdd.n2630 vdd.n1022 185
R1307 vdd.n1404 vdd.n1403 185
R1308 vdd.n1403 vdd.n1021 185
R1309 vdd.n1405 vdd.n1029 185
R1310 vdd.n2622 vdd.n1029 185
R1311 vdd.n1407 vdd.n1406 185
R1312 vdd.n1406 vdd.n1028 185
R1313 vdd.n1408 vdd.n1034 185
R1314 vdd.n2616 vdd.n1034 185
R1315 vdd.n1427 vdd.n1426 185
R1316 vdd.n1426 vdd.n1425 185
R1317 vdd.n1428 vdd.n1039 185
R1318 vdd.n2610 vdd.n1039 185
R1319 vdd.n1430 vdd.n1429 185
R1320 vdd.n1429 vdd.n1046 185
R1321 vdd.n1431 vdd.n1044 185
R1322 vdd.n2604 vdd.n1044 185
R1323 vdd.n1433 vdd.n1432 185
R1324 vdd.n1432 vdd.n1052 185
R1325 vdd.n1434 vdd.n1050 185
R1326 vdd.n2598 vdd.n1050 185
R1327 vdd.n1436 vdd.n1435 185
R1328 vdd.n1437 vdd.n1436 185
R1329 vdd.n1396 vdd.n1057 185
R1330 vdd.n2592 vdd.n1057 185
R1331 vdd.n1395 vdd.n1394 185
R1332 vdd.n1394 vdd.n1056 185
R1333 vdd.n1393 vdd.n1063 185
R1334 vdd.n2586 vdd.n1063 185
R1335 vdd.n1392 vdd.n1391 185
R1336 vdd.n1391 vdd.n1062 185
R1337 vdd.n1390 vdd.n1068 185
R1338 vdd.n2580 vdd.n1068 185
R1339 vdd.n1389 vdd.n1388 185
R1340 vdd.n1388 vdd.n1076 185
R1341 vdd.n1387 vdd.n1074 185
R1342 vdd.n2573 vdd.n1074 185
R1343 vdd.n1386 vdd.n1385 185
R1344 vdd.n1385 vdd.n1083 185
R1345 vdd.n1384 vdd.n1081 185
R1346 vdd.n2567 vdd.n1081 185
R1347 vdd.n1383 vdd.n1382 185
R1348 vdd.n1382 vdd.n1080 185
R1349 vdd.n1381 vdd.n1088 185
R1350 vdd.n2561 vdd.n1088 185
R1351 vdd.n1380 vdd.n1379 185
R1352 vdd.n1379 vdd.n1087 185
R1353 vdd.n1378 vdd.n1094 185
R1354 vdd.n2555 vdd.n1094 185
R1355 vdd.n1377 vdd.n1376 185
R1356 vdd.n1376 vdd.n1093 185
R1357 vdd.n1375 vdd.n1099 185
R1358 vdd.n2549 vdd.n1099 185
R1359 vdd.n1374 vdd.n1373 185
R1360 vdd.n1373 vdd.n1106 185
R1361 vdd.n1372 vdd.n1104 185
R1362 vdd.n2543 vdd.n1104 185
R1363 vdd.n1371 vdd.n1370 185
R1364 vdd.n1370 vdd.n1112 185
R1365 vdd.n1369 vdd.n1110 185
R1366 vdd.n2537 vdd.n1110 185
R1367 vdd.n1368 vdd.n1367 185
R1368 vdd.n1367 vdd.n1119 185
R1369 vdd.n1366 vdd.n1117 185
R1370 vdd.n2531 vdd.n1117 185
R1371 vdd.n1365 vdd.n1364 185
R1372 vdd.n1364 vdd.n1116 185
R1373 vdd.n1363 vdd.n1124 185
R1374 vdd.n2525 vdd.n1124 185
R1375 vdd.n1362 vdd.n1361 185
R1376 vdd.n1361 vdd.n1123 185
R1377 vdd.n1360 vdd.n1129 185
R1378 vdd.n2519 vdd.n1129 185
R1379 vdd.n1359 vdd.n1358 185
R1380 vdd.n1358 vdd.n1137 185
R1381 vdd.n1357 vdd.n1135 185
R1382 vdd.n2513 vdd.n1135 185
R1383 vdd.n1356 vdd.n1355 185
R1384 vdd.n1355 vdd.n1134 185
R1385 vdd.n3629 vdd.n3628 185
R1386 vdd.n3628 vdd.n3627 185
R1387 vdd.n3630 vdd.n387 185
R1388 vdd.n387 vdd.n386 185
R1389 vdd.n3632 vdd.n3631 185
R1390 vdd.n3633 vdd.n3632 185
R1391 vdd.n382 vdd.n381 185
R1392 vdd.n3634 vdd.n382 185
R1393 vdd.n3637 vdd.n3636 185
R1394 vdd.n3636 vdd.n3635 185
R1395 vdd.n3638 vdd.n376 185
R1396 vdd.n376 vdd.n375 185
R1397 vdd.n3640 vdd.n3639 185
R1398 vdd.n3641 vdd.n3640 185
R1399 vdd.n371 vdd.n370 185
R1400 vdd.n3642 vdd.n371 185
R1401 vdd.n3645 vdd.n3644 185
R1402 vdd.n3644 vdd.n3643 185
R1403 vdd.n3646 vdd.n365 185
R1404 vdd.n3603 vdd.n365 185
R1405 vdd.n3648 vdd.n3647 185
R1406 vdd.n3649 vdd.n3648 185
R1407 vdd.n360 vdd.n359 185
R1408 vdd.n3650 vdd.n360 185
R1409 vdd.n3653 vdd.n3652 185
R1410 vdd.n3652 vdd.n3651 185
R1411 vdd.n3654 vdd.n354 185
R1412 vdd.n361 vdd.n354 185
R1413 vdd.n3656 vdd.n3655 185
R1414 vdd.n3657 vdd.n3656 185
R1415 vdd.n350 vdd.n349 185
R1416 vdd.n3658 vdd.n350 185
R1417 vdd.n3661 vdd.n3660 185
R1418 vdd.n3660 vdd.n3659 185
R1419 vdd.n3662 vdd.n345 185
R1420 vdd.n345 vdd.n344 185
R1421 vdd.n3664 vdd.n3663 185
R1422 vdd.n3665 vdd.n3664 185
R1423 vdd.n339 vdd.n337 185
R1424 vdd.n3666 vdd.n339 185
R1425 vdd.n3669 vdd.n3668 185
R1426 vdd.n3668 vdd.n3667 185
R1427 vdd.n338 vdd.n336 185
R1428 vdd.n340 vdd.n338 185
R1429 vdd.n3579 vdd.n3578 185
R1430 vdd.n3580 vdd.n3579 185
R1431 vdd.n635 vdd.n634 185
R1432 vdd.n634 vdd.n633 185
R1433 vdd.n3574 vdd.n3573 185
R1434 vdd.n3573 vdd.n3572 185
R1435 vdd.n638 vdd.n637 185
R1436 vdd.n644 vdd.n638 185
R1437 vdd.n3560 vdd.n3559 185
R1438 vdd.n3561 vdd.n3560 185
R1439 vdd.n646 vdd.n645 185
R1440 vdd.n3552 vdd.n645 185
R1441 vdd.n3555 vdd.n3554 185
R1442 vdd.n3554 vdd.n3553 185
R1443 vdd.n649 vdd.n648 185
R1444 vdd.n656 vdd.n649 185
R1445 vdd.n3543 vdd.n3542 185
R1446 vdd.n3544 vdd.n3543 185
R1447 vdd.n658 vdd.n657 185
R1448 vdd.n657 vdd.n655 185
R1449 vdd.n3538 vdd.n3537 185
R1450 vdd.n3537 vdd.n3536 185
R1451 vdd.n661 vdd.n660 185
R1452 vdd.n662 vdd.n661 185
R1453 vdd.n3527 vdd.n3526 185
R1454 vdd.n3528 vdd.n3527 185
R1455 vdd.n669 vdd.n668 185
R1456 vdd.n3519 vdd.n668 185
R1457 vdd.n3522 vdd.n3521 185
R1458 vdd.n3521 vdd.n3520 185
R1459 vdd.n672 vdd.n671 185
R1460 vdd.n679 vdd.n672 185
R1461 vdd.n3510 vdd.n3509 185
R1462 vdd.n3511 vdd.n3510 185
R1463 vdd.n681 vdd.n680 185
R1464 vdd.n680 vdd.n678 185
R1465 vdd.n3505 vdd.n3504 185
R1466 vdd.n3504 vdd.n3503 185
R1467 vdd.n684 vdd.n683 185
R1468 vdd.n723 vdd.n684 185
R1469 vdd.n3493 vdd.n3492 185
R1470 vdd.n3491 vdd.n725 185
R1471 vdd.n3490 vdd.n724 185
R1472 vdd.n3495 vdd.n724 185
R1473 vdd.n729 vdd.n728 185
R1474 vdd.n733 vdd.n732 185
R1475 vdd.n3486 vdd.n734 185
R1476 vdd.n3485 vdd.n3484 185
R1477 vdd.n3483 vdd.n3482 185
R1478 vdd.n3481 vdd.n3480 185
R1479 vdd.n3479 vdd.n3478 185
R1480 vdd.n3477 vdd.n3476 185
R1481 vdd.n3475 vdd.n3474 185
R1482 vdd.n3473 vdd.n3472 185
R1483 vdd.n3471 vdd.n3470 185
R1484 vdd.n3469 vdd.n3468 185
R1485 vdd.n3467 vdd.n3466 185
R1486 vdd.n3465 vdd.n3464 185
R1487 vdd.n3463 vdd.n3462 185
R1488 vdd.n3461 vdd.n3460 185
R1489 vdd.n3459 vdd.n3458 185
R1490 vdd.n3450 vdd.n747 185
R1491 vdd.n3452 vdd.n3451 185
R1492 vdd.n3449 vdd.n3448 185
R1493 vdd.n3447 vdd.n3446 185
R1494 vdd.n3445 vdd.n3444 185
R1495 vdd.n3443 vdd.n3442 185
R1496 vdd.n3441 vdd.n3440 185
R1497 vdd.n3439 vdd.n3438 185
R1498 vdd.n3437 vdd.n3436 185
R1499 vdd.n3435 vdd.n3434 185
R1500 vdd.n3433 vdd.n3432 185
R1501 vdd.n3431 vdd.n3430 185
R1502 vdd.n3429 vdd.n3428 185
R1503 vdd.n3427 vdd.n3426 185
R1504 vdd.n3425 vdd.n3424 185
R1505 vdd.n3423 vdd.n3422 185
R1506 vdd.n3421 vdd.n3420 185
R1507 vdd.n3419 vdd.n3418 185
R1508 vdd.n3417 vdd.n3416 185
R1509 vdd.n3415 vdd.n3414 185
R1510 vdd.n3413 vdd.n3412 185
R1511 vdd.n3411 vdd.n3410 185
R1512 vdd.n3404 vdd.n767 185
R1513 vdd.n3406 vdd.n3405 185
R1514 vdd.n3403 vdd.n3402 185
R1515 vdd.n3401 vdd.n3400 185
R1516 vdd.n3399 vdd.n3398 185
R1517 vdd.n3397 vdd.n3396 185
R1518 vdd.n3395 vdd.n3394 185
R1519 vdd.n3393 vdd.n3392 185
R1520 vdd.n3391 vdd.n3390 185
R1521 vdd.n3389 vdd.n3388 185
R1522 vdd.n3387 vdd.n3386 185
R1523 vdd.n3385 vdd.n3384 185
R1524 vdd.n3383 vdd.n3382 185
R1525 vdd.n3381 vdd.n3380 185
R1526 vdd.n3379 vdd.n3378 185
R1527 vdd.n3377 vdd.n3376 185
R1528 vdd.n3375 vdd.n3374 185
R1529 vdd.n3373 vdd.n3372 185
R1530 vdd.n3371 vdd.n3370 185
R1531 vdd.n3369 vdd.n3368 185
R1532 vdd.n3367 vdd.n691 185
R1533 vdd.n3497 vdd.n3496 185
R1534 vdd.n3496 vdd.n3495 185
R1535 vdd.n3624 vdd.n3623 185
R1536 vdd.n618 vdd.n425 185
R1537 vdd.n617 vdd.n616 185
R1538 vdd.n615 vdd.n614 185
R1539 vdd.n613 vdd.n430 185
R1540 vdd.n609 vdd.n608 185
R1541 vdd.n607 vdd.n606 185
R1542 vdd.n605 vdd.n604 185
R1543 vdd.n603 vdd.n432 185
R1544 vdd.n599 vdd.n598 185
R1545 vdd.n597 vdd.n596 185
R1546 vdd.n595 vdd.n594 185
R1547 vdd.n593 vdd.n434 185
R1548 vdd.n589 vdd.n588 185
R1549 vdd.n587 vdd.n586 185
R1550 vdd.n585 vdd.n584 185
R1551 vdd.n583 vdd.n436 185
R1552 vdd.n579 vdd.n578 185
R1553 vdd.n577 vdd.n576 185
R1554 vdd.n575 vdd.n574 185
R1555 vdd.n573 vdd.n438 185
R1556 vdd.n569 vdd.n568 185
R1557 vdd.n567 vdd.n566 185
R1558 vdd.n565 vdd.n564 185
R1559 vdd.n563 vdd.n442 185
R1560 vdd.n559 vdd.n558 185
R1561 vdd.n557 vdd.n556 185
R1562 vdd.n555 vdd.n554 185
R1563 vdd.n553 vdd.n444 185
R1564 vdd.n549 vdd.n548 185
R1565 vdd.n547 vdd.n546 185
R1566 vdd.n545 vdd.n544 185
R1567 vdd.n543 vdd.n446 185
R1568 vdd.n539 vdd.n538 185
R1569 vdd.n537 vdd.n536 185
R1570 vdd.n535 vdd.n534 185
R1571 vdd.n533 vdd.n448 185
R1572 vdd.n529 vdd.n528 185
R1573 vdd.n527 vdd.n526 185
R1574 vdd.n525 vdd.n524 185
R1575 vdd.n523 vdd.n450 185
R1576 vdd.n519 vdd.n518 185
R1577 vdd.n517 vdd.n516 185
R1578 vdd.n515 vdd.n514 185
R1579 vdd.n513 vdd.n454 185
R1580 vdd.n509 vdd.n508 185
R1581 vdd.n507 vdd.n506 185
R1582 vdd.n505 vdd.n504 185
R1583 vdd.n503 vdd.n456 185
R1584 vdd.n499 vdd.n498 185
R1585 vdd.n497 vdd.n496 185
R1586 vdd.n495 vdd.n494 185
R1587 vdd.n493 vdd.n458 185
R1588 vdd.n489 vdd.n488 185
R1589 vdd.n487 vdd.n486 185
R1590 vdd.n485 vdd.n484 185
R1591 vdd.n483 vdd.n460 185
R1592 vdd.n479 vdd.n478 185
R1593 vdd.n477 vdd.n476 185
R1594 vdd.n475 vdd.n474 185
R1595 vdd.n473 vdd.n462 185
R1596 vdd.n469 vdd.n468 185
R1597 vdd.n467 vdd.n466 185
R1598 vdd.n465 vdd.n392 185
R1599 vdd.n3620 vdd.n393 185
R1600 vdd.n3627 vdd.n393 185
R1601 vdd.n3619 vdd.n3618 185
R1602 vdd.n3618 vdd.n386 185
R1603 vdd.n3617 vdd.n385 185
R1604 vdd.n3633 vdd.n385 185
R1605 vdd.n621 vdd.n384 185
R1606 vdd.n3634 vdd.n384 185
R1607 vdd.n3613 vdd.n383 185
R1608 vdd.n3635 vdd.n383 185
R1609 vdd.n3612 vdd.n3611 185
R1610 vdd.n3611 vdd.n375 185
R1611 vdd.n3610 vdd.n374 185
R1612 vdd.n3641 vdd.n374 185
R1613 vdd.n623 vdd.n373 185
R1614 vdd.n3642 vdd.n373 185
R1615 vdd.n3606 vdd.n372 185
R1616 vdd.n3643 vdd.n372 185
R1617 vdd.n3605 vdd.n3604 185
R1618 vdd.n3604 vdd.n3603 185
R1619 vdd.n3602 vdd.n364 185
R1620 vdd.n3649 vdd.n364 185
R1621 vdd.n625 vdd.n363 185
R1622 vdd.n3650 vdd.n363 185
R1623 vdd.n3598 vdd.n362 185
R1624 vdd.n3651 vdd.n362 185
R1625 vdd.n3597 vdd.n3596 185
R1626 vdd.n3596 vdd.n361 185
R1627 vdd.n3595 vdd.n353 185
R1628 vdd.n3657 vdd.n353 185
R1629 vdd.n627 vdd.n352 185
R1630 vdd.n3658 vdd.n352 185
R1631 vdd.n3591 vdd.n351 185
R1632 vdd.n3659 vdd.n351 185
R1633 vdd.n3590 vdd.n3589 185
R1634 vdd.n3589 vdd.n344 185
R1635 vdd.n3588 vdd.n343 185
R1636 vdd.n3665 vdd.n343 185
R1637 vdd.n629 vdd.n342 185
R1638 vdd.n3666 vdd.n342 185
R1639 vdd.n3584 vdd.n341 185
R1640 vdd.n3667 vdd.n341 185
R1641 vdd.n3583 vdd.n3582 185
R1642 vdd.n3582 vdd.n340 185
R1643 vdd.n3581 vdd.n631 185
R1644 vdd.n3581 vdd.n3580 185
R1645 vdd.n3569 vdd.n632 185
R1646 vdd.n633 vdd.n632 185
R1647 vdd.n3571 vdd.n3570 185
R1648 vdd.n3572 vdd.n3571 185
R1649 vdd.n640 vdd.n639 185
R1650 vdd.n644 vdd.n639 185
R1651 vdd.n3563 vdd.n3562 185
R1652 vdd.n3562 vdd.n3561 185
R1653 vdd.n643 vdd.n642 185
R1654 vdd.n3552 vdd.n643 185
R1655 vdd.n3551 vdd.n3550 185
R1656 vdd.n3553 vdd.n3551 185
R1657 vdd.n651 vdd.n650 185
R1658 vdd.n656 vdd.n650 185
R1659 vdd.n3546 vdd.n3545 185
R1660 vdd.n3545 vdd.n3544 185
R1661 vdd.n654 vdd.n653 185
R1662 vdd.n655 vdd.n654 185
R1663 vdd.n3535 vdd.n3534 185
R1664 vdd.n3536 vdd.n3535 185
R1665 vdd.n664 vdd.n663 185
R1666 vdd.n663 vdd.n662 185
R1667 vdd.n3530 vdd.n3529 185
R1668 vdd.n3529 vdd.n3528 185
R1669 vdd.n667 vdd.n666 185
R1670 vdd.n3519 vdd.n667 185
R1671 vdd.n3518 vdd.n3517 185
R1672 vdd.n3520 vdd.n3518 185
R1673 vdd.n674 vdd.n673 185
R1674 vdd.n679 vdd.n673 185
R1675 vdd.n3513 vdd.n3512 185
R1676 vdd.n3512 vdd.n3511 185
R1677 vdd.n677 vdd.n676 185
R1678 vdd.n678 vdd.n677 185
R1679 vdd.n3502 vdd.n3501 185
R1680 vdd.n3503 vdd.n3502 185
R1681 vdd.n686 vdd.n685 185
R1682 vdd.n723 vdd.n685 185
R1683 vdd.n3091 vdd.n3090 185
R1684 vdd.n962 vdd.n961 185
R1685 vdd.n3087 vdd.n3086 185
R1686 vdd.n3088 vdd.n3087 185
R1687 vdd.n3085 vdd.n2819 185
R1688 vdd.n3084 vdd.n3083 185
R1689 vdd.n3082 vdd.n3081 185
R1690 vdd.n3080 vdd.n3079 185
R1691 vdd.n3078 vdd.n3077 185
R1692 vdd.n3076 vdd.n3075 185
R1693 vdd.n3074 vdd.n3073 185
R1694 vdd.n3072 vdd.n3071 185
R1695 vdd.n3070 vdd.n3069 185
R1696 vdd.n3068 vdd.n3067 185
R1697 vdd.n3066 vdd.n3065 185
R1698 vdd.n3064 vdd.n3063 185
R1699 vdd.n3062 vdd.n3061 185
R1700 vdd.n3060 vdd.n3059 185
R1701 vdd.n3058 vdd.n3057 185
R1702 vdd.n3056 vdd.n3055 185
R1703 vdd.n3054 vdd.n3053 185
R1704 vdd.n3052 vdd.n3051 185
R1705 vdd.n3050 vdd.n3049 185
R1706 vdd.n3048 vdd.n3047 185
R1707 vdd.n3046 vdd.n3045 185
R1708 vdd.n3044 vdd.n3043 185
R1709 vdd.n3042 vdd.n3041 185
R1710 vdd.n3040 vdd.n3039 185
R1711 vdd.n3038 vdd.n3037 185
R1712 vdd.n3036 vdd.n3035 185
R1713 vdd.n3034 vdd.n3033 185
R1714 vdd.n3032 vdd.n3031 185
R1715 vdd.n3030 vdd.n3029 185
R1716 vdd.n3027 vdd.n3026 185
R1717 vdd.n3025 vdd.n3024 185
R1718 vdd.n3023 vdd.n3022 185
R1719 vdd.n3267 vdd.n3266 185
R1720 vdd.n3269 vdd.n834 185
R1721 vdd.n3271 vdd.n3270 185
R1722 vdd.n3273 vdd.n831 185
R1723 vdd.n3275 vdd.n3274 185
R1724 vdd.n3277 vdd.n829 185
R1725 vdd.n3279 vdd.n3278 185
R1726 vdd.n3280 vdd.n828 185
R1727 vdd.n3282 vdd.n3281 185
R1728 vdd.n3284 vdd.n826 185
R1729 vdd.n3286 vdd.n3285 185
R1730 vdd.n3287 vdd.n825 185
R1731 vdd.n3289 vdd.n3288 185
R1732 vdd.n3291 vdd.n823 185
R1733 vdd.n3293 vdd.n3292 185
R1734 vdd.n3294 vdd.n822 185
R1735 vdd.n3296 vdd.n3295 185
R1736 vdd.n3298 vdd.n731 185
R1737 vdd.n3300 vdd.n3299 185
R1738 vdd.n3302 vdd.n820 185
R1739 vdd.n3304 vdd.n3303 185
R1740 vdd.n3305 vdd.n819 185
R1741 vdd.n3307 vdd.n3306 185
R1742 vdd.n3309 vdd.n817 185
R1743 vdd.n3311 vdd.n3310 185
R1744 vdd.n3312 vdd.n816 185
R1745 vdd.n3314 vdd.n3313 185
R1746 vdd.n3316 vdd.n814 185
R1747 vdd.n3318 vdd.n3317 185
R1748 vdd.n3319 vdd.n813 185
R1749 vdd.n3321 vdd.n3320 185
R1750 vdd.n3323 vdd.n812 185
R1751 vdd.n3324 vdd.n811 185
R1752 vdd.n3327 vdd.n3326 185
R1753 vdd.n3328 vdd.n809 185
R1754 vdd.n809 vdd.n692 185
R1755 vdd.n3265 vdd.n806 185
R1756 vdd.n3331 vdd.n806 185
R1757 vdd.n3264 vdd.n3263 185
R1758 vdd.n3263 vdd.n805 185
R1759 vdd.n3262 vdd.n836 185
R1760 vdd.n3262 vdd.n3261 185
R1761 vdd.n2905 vdd.n837 185
R1762 vdd.n846 vdd.n837 185
R1763 vdd.n2906 vdd.n844 185
R1764 vdd.n3255 vdd.n844 185
R1765 vdd.n2908 vdd.n2907 185
R1766 vdd.n2907 vdd.n843 185
R1767 vdd.n2909 vdd.n852 185
R1768 vdd.n3204 vdd.n852 185
R1769 vdd.n2911 vdd.n2910 185
R1770 vdd.n2910 vdd.n851 185
R1771 vdd.n2912 vdd.n857 185
R1772 vdd.n3198 vdd.n857 185
R1773 vdd.n2914 vdd.n2913 185
R1774 vdd.n2913 vdd.n864 185
R1775 vdd.n2915 vdd.n862 185
R1776 vdd.n3192 vdd.n862 185
R1777 vdd.n2917 vdd.n2916 185
R1778 vdd.n2916 vdd.n870 185
R1779 vdd.n2918 vdd.n868 185
R1780 vdd.n3186 vdd.n868 185
R1781 vdd.n2920 vdd.n2919 185
R1782 vdd.n2919 vdd.n877 185
R1783 vdd.n2921 vdd.n875 185
R1784 vdd.n3180 vdd.n875 185
R1785 vdd.n2923 vdd.n2922 185
R1786 vdd.n2922 vdd.n874 185
R1787 vdd.n2924 vdd.n882 185
R1788 vdd.n3174 vdd.n882 185
R1789 vdd.n2926 vdd.n2925 185
R1790 vdd.n2925 vdd.n881 185
R1791 vdd.n2927 vdd.n888 185
R1792 vdd.n3168 vdd.n888 185
R1793 vdd.n2929 vdd.n2928 185
R1794 vdd.n2928 vdd.n887 185
R1795 vdd.n2930 vdd.n893 185
R1796 vdd.n3162 vdd.n893 185
R1797 vdd.n2932 vdd.n2931 185
R1798 vdd.n2931 vdd.n901 185
R1799 vdd.n2933 vdd.n899 185
R1800 vdd.n3156 vdd.n899 185
R1801 vdd.n2935 vdd.n2934 185
R1802 vdd.n2934 vdd.n908 185
R1803 vdd.n2936 vdd.n906 185
R1804 vdd.n3150 vdd.n906 185
R1805 vdd.n2938 vdd.n2937 185
R1806 vdd.n2937 vdd.n905 185
R1807 vdd.n2939 vdd.n913 185
R1808 vdd.n3143 vdd.n913 185
R1809 vdd.n2941 vdd.n2940 185
R1810 vdd.n2940 vdd.n912 185
R1811 vdd.n2942 vdd.n918 185
R1812 vdd.n3137 vdd.n918 185
R1813 vdd.n2944 vdd.n2943 185
R1814 vdd.n2943 vdd.n925 185
R1815 vdd.n2945 vdd.n923 185
R1816 vdd.n3131 vdd.n923 185
R1817 vdd.n2947 vdd.n2946 185
R1818 vdd.n2946 vdd.n931 185
R1819 vdd.n2948 vdd.n929 185
R1820 vdd.n3125 vdd.n929 185
R1821 vdd.n3000 vdd.n2999 185
R1822 vdd.n2999 vdd.n2998 185
R1823 vdd.n3001 vdd.n935 185
R1824 vdd.n3119 vdd.n935 185
R1825 vdd.n3003 vdd.n3002 185
R1826 vdd.n3004 vdd.n3003 185
R1827 vdd.n2904 vdd.n941 185
R1828 vdd.n3113 vdd.n941 185
R1829 vdd.n2903 vdd.n2902 185
R1830 vdd.n2902 vdd.n940 185
R1831 vdd.n2901 vdd.n947 185
R1832 vdd.n3107 vdd.n947 185
R1833 vdd.n2900 vdd.n2899 185
R1834 vdd.n2899 vdd.n946 185
R1835 vdd.n2822 vdd.n952 185
R1836 vdd.n3101 vdd.n952 185
R1837 vdd.n3018 vdd.n3017 185
R1838 vdd.n3017 vdd.n3016 185
R1839 vdd.n3019 vdd.n958 185
R1840 vdd.n3095 vdd.n958 185
R1841 vdd.n3021 vdd.n3020 185
R1842 vdd.n3021 vdd.n957 185
R1843 vdd.n3092 vdd.n960 185
R1844 vdd.n960 vdd.n957 185
R1845 vdd.n3094 vdd.n3093 185
R1846 vdd.n3095 vdd.n3094 185
R1847 vdd.n951 vdd.n950 185
R1848 vdd.n3016 vdd.n951 185
R1849 vdd.n3103 vdd.n3102 185
R1850 vdd.n3102 vdd.n3101 185
R1851 vdd.n3104 vdd.n949 185
R1852 vdd.n949 vdd.n946 185
R1853 vdd.n3106 vdd.n3105 185
R1854 vdd.n3107 vdd.n3106 185
R1855 vdd.n939 vdd.n938 185
R1856 vdd.n940 vdd.n939 185
R1857 vdd.n3115 vdd.n3114 185
R1858 vdd.n3114 vdd.n3113 185
R1859 vdd.n3116 vdd.n937 185
R1860 vdd.n3004 vdd.n937 185
R1861 vdd.n3118 vdd.n3117 185
R1862 vdd.n3119 vdd.n3118 185
R1863 vdd.n928 vdd.n927 185
R1864 vdd.n2998 vdd.n928 185
R1865 vdd.n3127 vdd.n3126 185
R1866 vdd.n3126 vdd.n3125 185
R1867 vdd.n3128 vdd.n926 185
R1868 vdd.n931 vdd.n926 185
R1869 vdd.n3130 vdd.n3129 185
R1870 vdd.n3131 vdd.n3130 185
R1871 vdd.n917 vdd.n916 185
R1872 vdd.n925 vdd.n917 185
R1873 vdd.n3139 vdd.n3138 185
R1874 vdd.n3138 vdd.n3137 185
R1875 vdd.n3140 vdd.n915 185
R1876 vdd.n915 vdd.n912 185
R1877 vdd.n3142 vdd.n3141 185
R1878 vdd.n3143 vdd.n3142 185
R1879 vdd.n904 vdd.n903 185
R1880 vdd.n905 vdd.n904 185
R1881 vdd.n3152 vdd.n3151 185
R1882 vdd.n3151 vdd.n3150 185
R1883 vdd.n3153 vdd.n902 185
R1884 vdd.n908 vdd.n902 185
R1885 vdd.n3155 vdd.n3154 185
R1886 vdd.n3156 vdd.n3155 185
R1887 vdd.n892 vdd.n891 185
R1888 vdd.n901 vdd.n892 185
R1889 vdd.n3164 vdd.n3163 185
R1890 vdd.n3163 vdd.n3162 185
R1891 vdd.n3165 vdd.n890 185
R1892 vdd.n890 vdd.n887 185
R1893 vdd.n3167 vdd.n3166 185
R1894 vdd.n3168 vdd.n3167 185
R1895 vdd.n880 vdd.n879 185
R1896 vdd.n881 vdd.n880 185
R1897 vdd.n3176 vdd.n3175 185
R1898 vdd.n3175 vdd.n3174 185
R1899 vdd.n3177 vdd.n878 185
R1900 vdd.n878 vdd.n874 185
R1901 vdd.n3179 vdd.n3178 185
R1902 vdd.n3180 vdd.n3179 185
R1903 vdd.n867 vdd.n866 185
R1904 vdd.n877 vdd.n867 185
R1905 vdd.n3188 vdd.n3187 185
R1906 vdd.n3187 vdd.n3186 185
R1907 vdd.n3189 vdd.n865 185
R1908 vdd.n870 vdd.n865 185
R1909 vdd.n3191 vdd.n3190 185
R1910 vdd.n3192 vdd.n3191 185
R1911 vdd.n856 vdd.n855 185
R1912 vdd.n864 vdd.n856 185
R1913 vdd.n3200 vdd.n3199 185
R1914 vdd.n3199 vdd.n3198 185
R1915 vdd.n3201 vdd.n854 185
R1916 vdd.n854 vdd.n851 185
R1917 vdd.n3203 vdd.n3202 185
R1918 vdd.n3204 vdd.n3203 185
R1919 vdd.n842 vdd.n841 185
R1920 vdd.n843 vdd.n842 185
R1921 vdd.n3257 vdd.n3256 185
R1922 vdd.n3256 vdd.n3255 185
R1923 vdd.n3258 vdd.n840 185
R1924 vdd.n846 vdd.n840 185
R1925 vdd.n3260 vdd.n3259 185
R1926 vdd.n3261 vdd.n3260 185
R1927 vdd.n810 vdd.n808 185
R1928 vdd.n808 vdd.n805 185
R1929 vdd.n3330 vdd.n3329 185
R1930 vdd.n3331 vdd.n3330 185
R1931 vdd.n2711 vdd.n2710 185
R1932 vdd.n2712 vdd.n2711 185
R1933 vdd.n1009 vdd.n1007 185
R1934 vdd.n1007 vdd.n1005 185
R1935 vdd.n2626 vdd.n1016 185
R1936 vdd.n2637 vdd.n1016 185
R1937 vdd.n2627 vdd.n1025 185
R1938 vdd.n1399 vdd.n1025 185
R1939 vdd.n2629 vdd.n2628 185
R1940 vdd.n2630 vdd.n2629 185
R1941 vdd.n2625 vdd.n1024 185
R1942 vdd.n1024 vdd.n1021 185
R1943 vdd.n2624 vdd.n2623 185
R1944 vdd.n2623 vdd.n2622 185
R1945 vdd.n1027 vdd.n1026 185
R1946 vdd.n1028 vdd.n1027 185
R1947 vdd.n2615 vdd.n2614 185
R1948 vdd.n2616 vdd.n2615 185
R1949 vdd.n2613 vdd.n1036 185
R1950 vdd.n1425 vdd.n1036 185
R1951 vdd.n2612 vdd.n2611 185
R1952 vdd.n2611 vdd.n2610 185
R1953 vdd.n1038 vdd.n1037 185
R1954 vdd.n1046 vdd.n1038 185
R1955 vdd.n2603 vdd.n2602 185
R1956 vdd.n2604 vdd.n2603 185
R1957 vdd.n2601 vdd.n1047 185
R1958 vdd.n1052 vdd.n1047 185
R1959 vdd.n2600 vdd.n2599 185
R1960 vdd.n2599 vdd.n2598 185
R1961 vdd.n1049 vdd.n1048 185
R1962 vdd.n1437 vdd.n1049 185
R1963 vdd.n2591 vdd.n2590 185
R1964 vdd.n2592 vdd.n2591 185
R1965 vdd.n2589 vdd.n1059 185
R1966 vdd.n1059 vdd.n1056 185
R1967 vdd.n2588 vdd.n2587 185
R1968 vdd.n2587 vdd.n2586 185
R1969 vdd.n1061 vdd.n1060 185
R1970 vdd.n1062 vdd.n1061 185
R1971 vdd.n2579 vdd.n2578 185
R1972 vdd.n2580 vdd.n2579 185
R1973 vdd.n2576 vdd.n1070 185
R1974 vdd.n1076 vdd.n1070 185
R1975 vdd.n2575 vdd.n2574 185
R1976 vdd.n2574 vdd.n2573 185
R1977 vdd.n1073 vdd.n1072 185
R1978 vdd.n1083 vdd.n1073 185
R1979 vdd.n2566 vdd.n2565 185
R1980 vdd.n2567 vdd.n2566 185
R1981 vdd.n2564 vdd.n1084 185
R1982 vdd.n1084 vdd.n1080 185
R1983 vdd.n2563 vdd.n2562 185
R1984 vdd.n2562 vdd.n2561 185
R1985 vdd.n1086 vdd.n1085 185
R1986 vdd.n1087 vdd.n1086 185
R1987 vdd.n2554 vdd.n2553 185
R1988 vdd.n2555 vdd.n2554 185
R1989 vdd.n2552 vdd.n1096 185
R1990 vdd.n1096 vdd.n1093 185
R1991 vdd.n2551 vdd.n2550 185
R1992 vdd.n2550 vdd.n2549 185
R1993 vdd.n1098 vdd.n1097 185
R1994 vdd.n1106 vdd.n1098 185
R1995 vdd.n2542 vdd.n2541 185
R1996 vdd.n2543 vdd.n2542 185
R1997 vdd.n2540 vdd.n1107 185
R1998 vdd.n1112 vdd.n1107 185
R1999 vdd.n2539 vdd.n2538 185
R2000 vdd.n2538 vdd.n2537 185
R2001 vdd.n1109 vdd.n1108 185
R2002 vdd.n1119 vdd.n1109 185
R2003 vdd.n2530 vdd.n2529 185
R2004 vdd.n2531 vdd.n2530 185
R2005 vdd.n2528 vdd.n1120 185
R2006 vdd.n1120 vdd.n1116 185
R2007 vdd.n2527 vdd.n2526 185
R2008 vdd.n2526 vdd.n2525 185
R2009 vdd.n1122 vdd.n1121 185
R2010 vdd.n1123 vdd.n1122 185
R2011 vdd.n2518 vdd.n2517 185
R2012 vdd.n2519 vdd.n2518 185
R2013 vdd.n2516 vdd.n1131 185
R2014 vdd.n1137 vdd.n1131 185
R2015 vdd.n2515 vdd.n2514 185
R2016 vdd.n2514 vdd.n2513 185
R2017 vdd.n1133 vdd.n1132 185
R2018 vdd.n1134 vdd.n1133 185
R2019 vdd.n2642 vdd.n980 185
R2020 vdd.n2784 vdd.n980 185
R2021 vdd.n2644 vdd.n2643 185
R2022 vdd.n2646 vdd.n2645 185
R2023 vdd.n2648 vdd.n2647 185
R2024 vdd.n2650 vdd.n2649 185
R2025 vdd.n2652 vdd.n2651 185
R2026 vdd.n2654 vdd.n2653 185
R2027 vdd.n2656 vdd.n2655 185
R2028 vdd.n2658 vdd.n2657 185
R2029 vdd.n2660 vdd.n2659 185
R2030 vdd.n2662 vdd.n2661 185
R2031 vdd.n2664 vdd.n2663 185
R2032 vdd.n2666 vdd.n2665 185
R2033 vdd.n2668 vdd.n2667 185
R2034 vdd.n2670 vdd.n2669 185
R2035 vdd.n2672 vdd.n2671 185
R2036 vdd.n2674 vdd.n2673 185
R2037 vdd.n2676 vdd.n2675 185
R2038 vdd.n2678 vdd.n2677 185
R2039 vdd.n2680 vdd.n2679 185
R2040 vdd.n2682 vdd.n2681 185
R2041 vdd.n2684 vdd.n2683 185
R2042 vdd.n2686 vdd.n2685 185
R2043 vdd.n2688 vdd.n2687 185
R2044 vdd.n2690 vdd.n2689 185
R2045 vdd.n2692 vdd.n2691 185
R2046 vdd.n2694 vdd.n2693 185
R2047 vdd.n2696 vdd.n2695 185
R2048 vdd.n2698 vdd.n2697 185
R2049 vdd.n2700 vdd.n2699 185
R2050 vdd.n2702 vdd.n2701 185
R2051 vdd.n2704 vdd.n2703 185
R2052 vdd.n2706 vdd.n2705 185
R2053 vdd.n2708 vdd.n2707 185
R2054 vdd.n2709 vdd.n1008 185
R2055 vdd.n2641 vdd.n1006 185
R2056 vdd.n2712 vdd.n1006 185
R2057 vdd.n2640 vdd.n2639 185
R2058 vdd.n2639 vdd.n1005 185
R2059 vdd.n2638 vdd.n1013 185
R2060 vdd.n2638 vdd.n2637 185
R2061 vdd.n1415 vdd.n1014 185
R2062 vdd.n1399 vdd.n1014 185
R2063 vdd.n1416 vdd.n1023 185
R2064 vdd.n2630 vdd.n1023 185
R2065 vdd.n1418 vdd.n1417 185
R2066 vdd.n1417 vdd.n1021 185
R2067 vdd.n1419 vdd.n1030 185
R2068 vdd.n2622 vdd.n1030 185
R2069 vdd.n1421 vdd.n1420 185
R2070 vdd.n1420 vdd.n1028 185
R2071 vdd.n1422 vdd.n1035 185
R2072 vdd.n2616 vdd.n1035 185
R2073 vdd.n1424 vdd.n1423 185
R2074 vdd.n1425 vdd.n1424 185
R2075 vdd.n1414 vdd.n1040 185
R2076 vdd.n2610 vdd.n1040 185
R2077 vdd.n1413 vdd.n1412 185
R2078 vdd.n1412 vdd.n1046 185
R2079 vdd.n1411 vdd.n1045 185
R2080 vdd.n2604 vdd.n1045 185
R2081 vdd.n1410 vdd.n1409 185
R2082 vdd.n1409 vdd.n1052 185
R2083 vdd.n1318 vdd.n1051 185
R2084 vdd.n2598 vdd.n1051 185
R2085 vdd.n1439 vdd.n1438 185
R2086 vdd.n1438 vdd.n1437 185
R2087 vdd.n1440 vdd.n1058 185
R2088 vdd.n2592 vdd.n1058 185
R2089 vdd.n1442 vdd.n1441 185
R2090 vdd.n1441 vdd.n1056 185
R2091 vdd.n1443 vdd.n1064 185
R2092 vdd.n2586 vdd.n1064 185
R2093 vdd.n1445 vdd.n1444 185
R2094 vdd.n1444 vdd.n1062 185
R2095 vdd.n1446 vdd.n1069 185
R2096 vdd.n2580 vdd.n1069 185
R2097 vdd.n1448 vdd.n1447 185
R2098 vdd.n1447 vdd.n1076 185
R2099 vdd.n1449 vdd.n1075 185
R2100 vdd.n2573 vdd.n1075 185
R2101 vdd.n1451 vdd.n1450 185
R2102 vdd.n1450 vdd.n1083 185
R2103 vdd.n1452 vdd.n1082 185
R2104 vdd.n2567 vdd.n1082 185
R2105 vdd.n1454 vdd.n1453 185
R2106 vdd.n1453 vdd.n1080 185
R2107 vdd.n1455 vdd.n1089 185
R2108 vdd.n2561 vdd.n1089 185
R2109 vdd.n1457 vdd.n1456 185
R2110 vdd.n1456 vdd.n1087 185
R2111 vdd.n1458 vdd.n1095 185
R2112 vdd.n2555 vdd.n1095 185
R2113 vdd.n1460 vdd.n1459 185
R2114 vdd.n1459 vdd.n1093 185
R2115 vdd.n1461 vdd.n1100 185
R2116 vdd.n2549 vdd.n1100 185
R2117 vdd.n1463 vdd.n1462 185
R2118 vdd.n1462 vdd.n1106 185
R2119 vdd.n1464 vdd.n1105 185
R2120 vdd.n2543 vdd.n1105 185
R2121 vdd.n1466 vdd.n1465 185
R2122 vdd.n1465 vdd.n1112 185
R2123 vdd.n1467 vdd.n1111 185
R2124 vdd.n2537 vdd.n1111 185
R2125 vdd.n1469 vdd.n1468 185
R2126 vdd.n1468 vdd.n1119 185
R2127 vdd.n1470 vdd.n1118 185
R2128 vdd.n2531 vdd.n1118 185
R2129 vdd.n1472 vdd.n1471 185
R2130 vdd.n1471 vdd.n1116 185
R2131 vdd.n1473 vdd.n1125 185
R2132 vdd.n2525 vdd.n1125 185
R2133 vdd.n1475 vdd.n1474 185
R2134 vdd.n1474 vdd.n1123 185
R2135 vdd.n1476 vdd.n1130 185
R2136 vdd.n2519 vdd.n1130 185
R2137 vdd.n1478 vdd.n1477 185
R2138 vdd.n1477 vdd.n1137 185
R2139 vdd.n1479 vdd.n1136 185
R2140 vdd.n2513 vdd.n1136 185
R2141 vdd.n1481 vdd.n1480 185
R2142 vdd.n1480 vdd.n1134 185
R2143 vdd.n1281 vdd.n1280 185
R2144 vdd.n1283 vdd.n1282 185
R2145 vdd.n1285 vdd.n1284 185
R2146 vdd.n1287 vdd.n1286 185
R2147 vdd.n1289 vdd.n1288 185
R2148 vdd.n1291 vdd.n1290 185
R2149 vdd.n1293 vdd.n1292 185
R2150 vdd.n1295 vdd.n1294 185
R2151 vdd.n1297 vdd.n1296 185
R2152 vdd.n1299 vdd.n1298 185
R2153 vdd.n1301 vdd.n1300 185
R2154 vdd.n1303 vdd.n1302 185
R2155 vdd.n1305 vdd.n1304 185
R2156 vdd.n1307 vdd.n1306 185
R2157 vdd.n1309 vdd.n1308 185
R2158 vdd.n1311 vdd.n1310 185
R2159 vdd.n1313 vdd.n1312 185
R2160 vdd.n1515 vdd.n1314 185
R2161 vdd.n1514 vdd.n1513 185
R2162 vdd.n1512 vdd.n1511 185
R2163 vdd.n1510 vdd.n1509 185
R2164 vdd.n1508 vdd.n1507 185
R2165 vdd.n1506 vdd.n1505 185
R2166 vdd.n1504 vdd.n1503 185
R2167 vdd.n1502 vdd.n1501 185
R2168 vdd.n1500 vdd.n1499 185
R2169 vdd.n1498 vdd.n1497 185
R2170 vdd.n1496 vdd.n1495 185
R2171 vdd.n1494 vdd.n1493 185
R2172 vdd.n1492 vdd.n1491 185
R2173 vdd.n1490 vdd.n1489 185
R2174 vdd.n1488 vdd.n1487 185
R2175 vdd.n1486 vdd.n1485 185
R2176 vdd.n1484 vdd.n1483 185
R2177 vdd.n1482 vdd.n1175 185
R2178 vdd.n2506 vdd.n1175 185
R2179 vdd.n327 vdd.n326 171.744
R2180 vdd.n326 vdd.n325 171.744
R2181 vdd.n325 vdd.n294 171.744
R2182 vdd.n318 vdd.n294 171.744
R2183 vdd.n318 vdd.n317 171.744
R2184 vdd.n317 vdd.n299 171.744
R2185 vdd.n310 vdd.n299 171.744
R2186 vdd.n310 vdd.n309 171.744
R2187 vdd.n309 vdd.n303 171.744
R2188 vdd.n268 vdd.n267 171.744
R2189 vdd.n267 vdd.n266 171.744
R2190 vdd.n266 vdd.n235 171.744
R2191 vdd.n259 vdd.n235 171.744
R2192 vdd.n259 vdd.n258 171.744
R2193 vdd.n258 vdd.n240 171.744
R2194 vdd.n251 vdd.n240 171.744
R2195 vdd.n251 vdd.n250 171.744
R2196 vdd.n250 vdd.n244 171.744
R2197 vdd.n225 vdd.n224 171.744
R2198 vdd.n224 vdd.n223 171.744
R2199 vdd.n223 vdd.n192 171.744
R2200 vdd.n216 vdd.n192 171.744
R2201 vdd.n216 vdd.n215 171.744
R2202 vdd.n215 vdd.n197 171.744
R2203 vdd.n208 vdd.n197 171.744
R2204 vdd.n208 vdd.n207 171.744
R2205 vdd.n207 vdd.n201 171.744
R2206 vdd.n166 vdd.n165 171.744
R2207 vdd.n165 vdd.n164 171.744
R2208 vdd.n164 vdd.n133 171.744
R2209 vdd.n157 vdd.n133 171.744
R2210 vdd.n157 vdd.n156 171.744
R2211 vdd.n156 vdd.n138 171.744
R2212 vdd.n149 vdd.n138 171.744
R2213 vdd.n149 vdd.n148 171.744
R2214 vdd.n148 vdd.n142 171.744
R2215 vdd.n124 vdd.n123 171.744
R2216 vdd.n123 vdd.n122 171.744
R2217 vdd.n122 vdd.n91 171.744
R2218 vdd.n115 vdd.n91 171.744
R2219 vdd.n115 vdd.n114 171.744
R2220 vdd.n114 vdd.n96 171.744
R2221 vdd.n107 vdd.n96 171.744
R2222 vdd.n107 vdd.n106 171.744
R2223 vdd.n106 vdd.n100 171.744
R2224 vdd.n65 vdd.n64 171.744
R2225 vdd.n64 vdd.n63 171.744
R2226 vdd.n63 vdd.n32 171.744
R2227 vdd.n56 vdd.n32 171.744
R2228 vdd.n56 vdd.n55 171.744
R2229 vdd.n55 vdd.n37 171.744
R2230 vdd.n48 vdd.n37 171.744
R2231 vdd.n48 vdd.n47 171.744
R2232 vdd.n47 vdd.n41 171.744
R2233 vdd.n2201 vdd.n2200 171.744
R2234 vdd.n2200 vdd.n2199 171.744
R2235 vdd.n2199 vdd.n2168 171.744
R2236 vdd.n2192 vdd.n2168 171.744
R2237 vdd.n2192 vdd.n2191 171.744
R2238 vdd.n2191 vdd.n2173 171.744
R2239 vdd.n2184 vdd.n2173 171.744
R2240 vdd.n2184 vdd.n2183 171.744
R2241 vdd.n2183 vdd.n2177 171.744
R2242 vdd.n2260 vdd.n2259 171.744
R2243 vdd.n2259 vdd.n2258 171.744
R2244 vdd.n2258 vdd.n2227 171.744
R2245 vdd.n2251 vdd.n2227 171.744
R2246 vdd.n2251 vdd.n2250 171.744
R2247 vdd.n2250 vdd.n2232 171.744
R2248 vdd.n2243 vdd.n2232 171.744
R2249 vdd.n2243 vdd.n2242 171.744
R2250 vdd.n2242 vdd.n2236 171.744
R2251 vdd.n2099 vdd.n2098 171.744
R2252 vdd.n2098 vdd.n2097 171.744
R2253 vdd.n2097 vdd.n2066 171.744
R2254 vdd.n2090 vdd.n2066 171.744
R2255 vdd.n2090 vdd.n2089 171.744
R2256 vdd.n2089 vdd.n2071 171.744
R2257 vdd.n2082 vdd.n2071 171.744
R2258 vdd.n2082 vdd.n2081 171.744
R2259 vdd.n2081 vdd.n2075 171.744
R2260 vdd.n2158 vdd.n2157 171.744
R2261 vdd.n2157 vdd.n2156 171.744
R2262 vdd.n2156 vdd.n2125 171.744
R2263 vdd.n2149 vdd.n2125 171.744
R2264 vdd.n2149 vdd.n2148 171.744
R2265 vdd.n2148 vdd.n2130 171.744
R2266 vdd.n2141 vdd.n2130 171.744
R2267 vdd.n2141 vdd.n2140 171.744
R2268 vdd.n2140 vdd.n2134 171.744
R2269 vdd.n1998 vdd.n1997 171.744
R2270 vdd.n1997 vdd.n1996 171.744
R2271 vdd.n1996 vdd.n1965 171.744
R2272 vdd.n1989 vdd.n1965 171.744
R2273 vdd.n1989 vdd.n1988 171.744
R2274 vdd.n1988 vdd.n1970 171.744
R2275 vdd.n1981 vdd.n1970 171.744
R2276 vdd.n1981 vdd.n1980 171.744
R2277 vdd.n1980 vdd.n1974 171.744
R2278 vdd.n2057 vdd.n2056 171.744
R2279 vdd.n2056 vdd.n2055 171.744
R2280 vdd.n2055 vdd.n2024 171.744
R2281 vdd.n2048 vdd.n2024 171.744
R2282 vdd.n2048 vdd.n2047 171.744
R2283 vdd.n2047 vdd.n2029 171.744
R2284 vdd.n2040 vdd.n2029 171.744
R2285 vdd.n2040 vdd.n2039 171.744
R2286 vdd.n2039 vdd.n2033 171.744
R2287 vdd.n468 vdd.n467 146.341
R2288 vdd.n474 vdd.n473 146.341
R2289 vdd.n478 vdd.n477 146.341
R2290 vdd.n484 vdd.n483 146.341
R2291 vdd.n488 vdd.n487 146.341
R2292 vdd.n494 vdd.n493 146.341
R2293 vdd.n498 vdd.n497 146.341
R2294 vdd.n504 vdd.n503 146.341
R2295 vdd.n508 vdd.n507 146.341
R2296 vdd.n514 vdd.n513 146.341
R2297 vdd.n518 vdd.n517 146.341
R2298 vdd.n524 vdd.n523 146.341
R2299 vdd.n528 vdd.n527 146.341
R2300 vdd.n534 vdd.n533 146.341
R2301 vdd.n538 vdd.n537 146.341
R2302 vdd.n544 vdd.n543 146.341
R2303 vdd.n548 vdd.n547 146.341
R2304 vdd.n554 vdd.n553 146.341
R2305 vdd.n558 vdd.n557 146.341
R2306 vdd.n564 vdd.n563 146.341
R2307 vdd.n568 vdd.n567 146.341
R2308 vdd.n574 vdd.n573 146.341
R2309 vdd.n578 vdd.n577 146.341
R2310 vdd.n584 vdd.n583 146.341
R2311 vdd.n588 vdd.n587 146.341
R2312 vdd.n594 vdd.n593 146.341
R2313 vdd.n598 vdd.n597 146.341
R2314 vdd.n604 vdd.n603 146.341
R2315 vdd.n608 vdd.n607 146.341
R2316 vdd.n614 vdd.n613 146.341
R2317 vdd.n616 vdd.n425 146.341
R2318 vdd.n3502 vdd.n685 146.341
R2319 vdd.n3502 vdd.n677 146.341
R2320 vdd.n3512 vdd.n677 146.341
R2321 vdd.n3512 vdd.n673 146.341
R2322 vdd.n3518 vdd.n673 146.341
R2323 vdd.n3518 vdd.n667 146.341
R2324 vdd.n3529 vdd.n667 146.341
R2325 vdd.n3529 vdd.n663 146.341
R2326 vdd.n3535 vdd.n663 146.341
R2327 vdd.n3535 vdd.n654 146.341
R2328 vdd.n3545 vdd.n654 146.341
R2329 vdd.n3545 vdd.n650 146.341
R2330 vdd.n3551 vdd.n650 146.341
R2331 vdd.n3551 vdd.n643 146.341
R2332 vdd.n3562 vdd.n643 146.341
R2333 vdd.n3562 vdd.n639 146.341
R2334 vdd.n3571 vdd.n639 146.341
R2335 vdd.n3571 vdd.n632 146.341
R2336 vdd.n3581 vdd.n632 146.341
R2337 vdd.n3582 vdd.n3581 146.341
R2338 vdd.n3582 vdd.n341 146.341
R2339 vdd.n342 vdd.n341 146.341
R2340 vdd.n343 vdd.n342 146.341
R2341 vdd.n3589 vdd.n343 146.341
R2342 vdd.n3589 vdd.n351 146.341
R2343 vdd.n352 vdd.n351 146.341
R2344 vdd.n353 vdd.n352 146.341
R2345 vdd.n3596 vdd.n353 146.341
R2346 vdd.n3596 vdd.n362 146.341
R2347 vdd.n363 vdd.n362 146.341
R2348 vdd.n364 vdd.n363 146.341
R2349 vdd.n3604 vdd.n364 146.341
R2350 vdd.n3604 vdd.n372 146.341
R2351 vdd.n373 vdd.n372 146.341
R2352 vdd.n374 vdd.n373 146.341
R2353 vdd.n3611 vdd.n374 146.341
R2354 vdd.n3611 vdd.n383 146.341
R2355 vdd.n384 vdd.n383 146.341
R2356 vdd.n385 vdd.n384 146.341
R2357 vdd.n3618 vdd.n385 146.341
R2358 vdd.n3618 vdd.n393 146.341
R2359 vdd.n725 vdd.n724 146.341
R2360 vdd.n728 vdd.n724 146.341
R2361 vdd.n734 vdd.n733 146.341
R2362 vdd.n3484 vdd.n3483 146.341
R2363 vdd.n3480 vdd.n3479 146.341
R2364 vdd.n3476 vdd.n3475 146.341
R2365 vdd.n3472 vdd.n3471 146.341
R2366 vdd.n3468 vdd.n3467 146.341
R2367 vdd.n3464 vdd.n3463 146.341
R2368 vdd.n3460 vdd.n3459 146.341
R2369 vdd.n3451 vdd.n3450 146.341
R2370 vdd.n3448 vdd.n3447 146.341
R2371 vdd.n3444 vdd.n3443 146.341
R2372 vdd.n3440 vdd.n3439 146.341
R2373 vdd.n3436 vdd.n3435 146.341
R2374 vdd.n3432 vdd.n3431 146.341
R2375 vdd.n3428 vdd.n3427 146.341
R2376 vdd.n3424 vdd.n3423 146.341
R2377 vdd.n3420 vdd.n3419 146.341
R2378 vdd.n3416 vdd.n3415 146.341
R2379 vdd.n3412 vdd.n3411 146.341
R2380 vdd.n3405 vdd.n3404 146.341
R2381 vdd.n3402 vdd.n3401 146.341
R2382 vdd.n3398 vdd.n3397 146.341
R2383 vdd.n3394 vdd.n3393 146.341
R2384 vdd.n3390 vdd.n3389 146.341
R2385 vdd.n3386 vdd.n3385 146.341
R2386 vdd.n3382 vdd.n3381 146.341
R2387 vdd.n3378 vdd.n3377 146.341
R2388 vdd.n3374 vdd.n3373 146.341
R2389 vdd.n3370 vdd.n3369 146.341
R2390 vdd.n3496 vdd.n691 146.341
R2391 vdd.n3504 vdd.n684 146.341
R2392 vdd.n3504 vdd.n680 146.341
R2393 vdd.n3510 vdd.n680 146.341
R2394 vdd.n3510 vdd.n672 146.341
R2395 vdd.n3521 vdd.n672 146.341
R2396 vdd.n3521 vdd.n668 146.341
R2397 vdd.n3527 vdd.n668 146.341
R2398 vdd.n3527 vdd.n661 146.341
R2399 vdd.n3537 vdd.n661 146.341
R2400 vdd.n3537 vdd.n657 146.341
R2401 vdd.n3543 vdd.n657 146.341
R2402 vdd.n3543 vdd.n649 146.341
R2403 vdd.n3554 vdd.n649 146.341
R2404 vdd.n3554 vdd.n645 146.341
R2405 vdd.n3560 vdd.n645 146.341
R2406 vdd.n3560 vdd.n638 146.341
R2407 vdd.n3573 vdd.n638 146.341
R2408 vdd.n3573 vdd.n634 146.341
R2409 vdd.n3579 vdd.n634 146.341
R2410 vdd.n3579 vdd.n338 146.341
R2411 vdd.n3668 vdd.n338 146.341
R2412 vdd.n3668 vdd.n339 146.341
R2413 vdd.n3664 vdd.n339 146.341
R2414 vdd.n3664 vdd.n345 146.341
R2415 vdd.n3660 vdd.n345 146.341
R2416 vdd.n3660 vdd.n350 146.341
R2417 vdd.n3656 vdd.n350 146.341
R2418 vdd.n3656 vdd.n354 146.341
R2419 vdd.n3652 vdd.n354 146.341
R2420 vdd.n3652 vdd.n360 146.341
R2421 vdd.n3648 vdd.n360 146.341
R2422 vdd.n3648 vdd.n365 146.341
R2423 vdd.n3644 vdd.n365 146.341
R2424 vdd.n3644 vdd.n371 146.341
R2425 vdd.n3640 vdd.n371 146.341
R2426 vdd.n3640 vdd.n376 146.341
R2427 vdd.n3636 vdd.n376 146.341
R2428 vdd.n3636 vdd.n382 146.341
R2429 vdd.n3632 vdd.n382 146.341
R2430 vdd.n3632 vdd.n387 146.341
R2431 vdd.n3628 vdd.n387 146.341
R2432 vdd.n2471 vdd.n2470 146.341
R2433 vdd.n2468 vdd.n2465 146.341
R2434 vdd.n2463 vdd.n1185 146.341
R2435 vdd.n2459 vdd.n2458 146.341
R2436 vdd.n2456 vdd.n1189 146.341
R2437 vdd.n2452 vdd.n2451 146.341
R2438 vdd.n2449 vdd.n1196 146.341
R2439 vdd.n2445 vdd.n2444 146.341
R2440 vdd.n2442 vdd.n1203 146.341
R2441 vdd.n1214 vdd.n1211 146.341
R2442 vdd.n2434 vdd.n2433 146.341
R2443 vdd.n2431 vdd.n1216 146.341
R2444 vdd.n2427 vdd.n2426 146.341
R2445 vdd.n2424 vdd.n1222 146.341
R2446 vdd.n2420 vdd.n2419 146.341
R2447 vdd.n2417 vdd.n1229 146.341
R2448 vdd.n2413 vdd.n2412 146.341
R2449 vdd.n2410 vdd.n1236 146.341
R2450 vdd.n2406 vdd.n2405 146.341
R2451 vdd.n2403 vdd.n1243 146.341
R2452 vdd.n1254 vdd.n1251 146.341
R2453 vdd.n2395 vdd.n2394 146.341
R2454 vdd.n2392 vdd.n1256 146.341
R2455 vdd.n2388 vdd.n2387 146.341
R2456 vdd.n2385 vdd.n1262 146.341
R2457 vdd.n2381 vdd.n2380 146.341
R2458 vdd.n2378 vdd.n1269 146.341
R2459 vdd.n2374 vdd.n2373 146.341
R2460 vdd.n2371 vdd.n1276 146.341
R2461 vdd.n1522 vdd.n1520 146.341
R2462 vdd.n1525 vdd.n1524 146.341
R2463 vdd.n1883 vdd.n1643 146.341
R2464 vdd.n1883 vdd.n1639 146.341
R2465 vdd.n1889 vdd.n1639 146.341
R2466 vdd.n1889 vdd.n1631 146.341
R2467 vdd.n1900 vdd.n1631 146.341
R2468 vdd.n1900 vdd.n1627 146.341
R2469 vdd.n1906 vdd.n1627 146.341
R2470 vdd.n1906 vdd.n1621 146.341
R2471 vdd.n1917 vdd.n1621 146.341
R2472 vdd.n1917 vdd.n1617 146.341
R2473 vdd.n1923 vdd.n1617 146.341
R2474 vdd.n1923 vdd.n1608 146.341
R2475 vdd.n1933 vdd.n1608 146.341
R2476 vdd.n1933 vdd.n1604 146.341
R2477 vdd.n1939 vdd.n1604 146.341
R2478 vdd.n1939 vdd.n1597 146.341
R2479 vdd.n1950 vdd.n1597 146.341
R2480 vdd.n1950 vdd.n1593 146.341
R2481 vdd.n1956 vdd.n1593 146.341
R2482 vdd.n1956 vdd.n1586 146.341
R2483 vdd.n2273 vdd.n1586 146.341
R2484 vdd.n2273 vdd.n1582 146.341
R2485 vdd.n2279 vdd.n1582 146.341
R2486 vdd.n2279 vdd.n1574 146.341
R2487 vdd.n2290 vdd.n1574 146.341
R2488 vdd.n2290 vdd.n1570 146.341
R2489 vdd.n2296 vdd.n1570 146.341
R2490 vdd.n2296 vdd.n1564 146.341
R2491 vdd.n2307 vdd.n1564 146.341
R2492 vdd.n2307 vdd.n1560 146.341
R2493 vdd.n2313 vdd.n1560 146.341
R2494 vdd.n2313 vdd.n1551 146.341
R2495 vdd.n2323 vdd.n1551 146.341
R2496 vdd.n2323 vdd.n1547 146.341
R2497 vdd.n2329 vdd.n1547 146.341
R2498 vdd.n2329 vdd.n1541 146.341
R2499 vdd.n2340 vdd.n1541 146.341
R2500 vdd.n2340 vdd.n1536 146.341
R2501 vdd.n2348 vdd.n1536 146.341
R2502 vdd.n2348 vdd.n1527 146.341
R2503 vdd.n2359 vdd.n1527 146.341
R2504 vdd.n1872 vdd.n1648 146.341
R2505 vdd.n1872 vdd.n1681 146.341
R2506 vdd.n1685 vdd.n1684 146.341
R2507 vdd.n1687 vdd.n1686 146.341
R2508 vdd.n1691 vdd.n1690 146.341
R2509 vdd.n1693 vdd.n1692 146.341
R2510 vdd.n1697 vdd.n1696 146.341
R2511 vdd.n1699 vdd.n1698 146.341
R2512 vdd.n1703 vdd.n1702 146.341
R2513 vdd.n1705 vdd.n1704 146.341
R2514 vdd.n1711 vdd.n1710 146.341
R2515 vdd.n1713 vdd.n1712 146.341
R2516 vdd.n1717 vdd.n1716 146.341
R2517 vdd.n1719 vdd.n1718 146.341
R2518 vdd.n1723 vdd.n1722 146.341
R2519 vdd.n1725 vdd.n1724 146.341
R2520 vdd.n1729 vdd.n1728 146.341
R2521 vdd.n1731 vdd.n1730 146.341
R2522 vdd.n1735 vdd.n1734 146.341
R2523 vdd.n1737 vdd.n1736 146.341
R2524 vdd.n1809 vdd.n1740 146.341
R2525 vdd.n1742 vdd.n1741 146.341
R2526 vdd.n1746 vdd.n1745 146.341
R2527 vdd.n1748 vdd.n1747 146.341
R2528 vdd.n1752 vdd.n1751 146.341
R2529 vdd.n1754 vdd.n1753 146.341
R2530 vdd.n1758 vdd.n1757 146.341
R2531 vdd.n1760 vdd.n1759 146.341
R2532 vdd.n1764 vdd.n1763 146.341
R2533 vdd.n1766 vdd.n1765 146.341
R2534 vdd.n1770 vdd.n1769 146.341
R2535 vdd.n1771 vdd.n1679 146.341
R2536 vdd.n1881 vdd.n1644 146.341
R2537 vdd.n1881 vdd.n1637 146.341
R2538 vdd.n1892 vdd.n1637 146.341
R2539 vdd.n1892 vdd.n1633 146.341
R2540 vdd.n1898 vdd.n1633 146.341
R2541 vdd.n1898 vdd.n1626 146.341
R2542 vdd.n1909 vdd.n1626 146.341
R2543 vdd.n1909 vdd.n1622 146.341
R2544 vdd.n1915 vdd.n1622 146.341
R2545 vdd.n1915 vdd.n1615 146.341
R2546 vdd.n1925 vdd.n1615 146.341
R2547 vdd.n1925 vdd.n1611 146.341
R2548 vdd.n1931 vdd.n1611 146.341
R2549 vdd.n1931 vdd.n1603 146.341
R2550 vdd.n1942 vdd.n1603 146.341
R2551 vdd.n1942 vdd.n1599 146.341
R2552 vdd.n1948 vdd.n1599 146.341
R2553 vdd.n1948 vdd.n1592 146.341
R2554 vdd.n1958 vdd.n1592 146.341
R2555 vdd.n1958 vdd.n1588 146.341
R2556 vdd.n2271 vdd.n1588 146.341
R2557 vdd.n2271 vdd.n1580 146.341
R2558 vdd.n2282 vdd.n1580 146.341
R2559 vdd.n2282 vdd.n1576 146.341
R2560 vdd.n2288 vdd.n1576 146.341
R2561 vdd.n2288 vdd.n1569 146.341
R2562 vdd.n2299 vdd.n1569 146.341
R2563 vdd.n2299 vdd.n1565 146.341
R2564 vdd.n2305 vdd.n1565 146.341
R2565 vdd.n2305 vdd.n1558 146.341
R2566 vdd.n2315 vdd.n1558 146.341
R2567 vdd.n2315 vdd.n1554 146.341
R2568 vdd.n2321 vdd.n1554 146.341
R2569 vdd.n2321 vdd.n1546 146.341
R2570 vdd.n2332 vdd.n1546 146.341
R2571 vdd.n2332 vdd.n1542 146.341
R2572 vdd.n2338 vdd.n1542 146.341
R2573 vdd.n2338 vdd.n1534 146.341
R2574 vdd.n2351 vdd.n1534 146.341
R2575 vdd.n2351 vdd.n1529 146.341
R2576 vdd.n2357 vdd.n1529 146.341
R2577 vdd.n1315 vdd.t154 127.284
R2578 vdd.n1010 vdd.t194 127.284
R2579 vdd.n1319 vdd.t191 127.284
R2580 vdd.n1001 vdd.t215 127.284
R2581 vdd.n896 vdd.t178 127.284
R2582 vdd.n896 vdd.t179 127.284
R2583 vdd.n2823 vdd.t209 127.284
R2584 vdd.n832 vdd.t170 127.284
R2585 vdd.n2820 vdd.t202 127.284
R2586 vdd.n799 vdd.t149 127.284
R2587 vdd.n1071 vdd.t205 127.284
R2588 vdd.n1071 vdd.t206 127.284
R2589 vdd.n22 vdd.n20 117.314
R2590 vdd.n17 vdd.n15 117.314
R2591 vdd.n27 vdd.n26 116.927
R2592 vdd.n24 vdd.n23 116.927
R2593 vdd.n22 vdd.n21 116.927
R2594 vdd.n17 vdd.n16 116.927
R2595 vdd.n19 vdd.n18 116.927
R2596 vdd.n27 vdd.n25 116.927
R2597 vdd.n1316 vdd.t153 111.188
R2598 vdd.n1011 vdd.t195 111.188
R2599 vdd.n1320 vdd.t190 111.188
R2600 vdd.n1002 vdd.t216 111.188
R2601 vdd.n2824 vdd.t208 111.188
R2602 vdd.n833 vdd.t171 111.188
R2603 vdd.n2821 vdd.t201 111.188
R2604 vdd.n800 vdd.t150 111.188
R2605 vdd.n3094 vdd.n960 99.5127
R2606 vdd.n3094 vdd.n951 99.5127
R2607 vdd.n3102 vdd.n951 99.5127
R2608 vdd.n3102 vdd.n949 99.5127
R2609 vdd.n3106 vdd.n949 99.5127
R2610 vdd.n3106 vdd.n939 99.5127
R2611 vdd.n3114 vdd.n939 99.5127
R2612 vdd.n3114 vdd.n937 99.5127
R2613 vdd.n3118 vdd.n937 99.5127
R2614 vdd.n3118 vdd.n928 99.5127
R2615 vdd.n3126 vdd.n928 99.5127
R2616 vdd.n3126 vdd.n926 99.5127
R2617 vdd.n3130 vdd.n926 99.5127
R2618 vdd.n3130 vdd.n917 99.5127
R2619 vdd.n3138 vdd.n917 99.5127
R2620 vdd.n3138 vdd.n915 99.5127
R2621 vdd.n3142 vdd.n915 99.5127
R2622 vdd.n3142 vdd.n904 99.5127
R2623 vdd.n3151 vdd.n904 99.5127
R2624 vdd.n3151 vdd.n902 99.5127
R2625 vdd.n3155 vdd.n902 99.5127
R2626 vdd.n3155 vdd.n892 99.5127
R2627 vdd.n3163 vdd.n892 99.5127
R2628 vdd.n3163 vdd.n890 99.5127
R2629 vdd.n3167 vdd.n890 99.5127
R2630 vdd.n3167 vdd.n880 99.5127
R2631 vdd.n3175 vdd.n880 99.5127
R2632 vdd.n3175 vdd.n878 99.5127
R2633 vdd.n3179 vdd.n878 99.5127
R2634 vdd.n3179 vdd.n867 99.5127
R2635 vdd.n3187 vdd.n867 99.5127
R2636 vdd.n3187 vdd.n865 99.5127
R2637 vdd.n3191 vdd.n865 99.5127
R2638 vdd.n3191 vdd.n856 99.5127
R2639 vdd.n3199 vdd.n856 99.5127
R2640 vdd.n3199 vdd.n854 99.5127
R2641 vdd.n3203 vdd.n854 99.5127
R2642 vdd.n3203 vdd.n842 99.5127
R2643 vdd.n3256 vdd.n842 99.5127
R2644 vdd.n3256 vdd.n840 99.5127
R2645 vdd.n3260 vdd.n840 99.5127
R2646 vdd.n3260 vdd.n808 99.5127
R2647 vdd.n3330 vdd.n808 99.5127
R2648 vdd.n3326 vdd.n809 99.5127
R2649 vdd.n3324 vdd.n3323 99.5127
R2650 vdd.n3321 vdd.n813 99.5127
R2651 vdd.n3317 vdd.n3316 99.5127
R2652 vdd.n3314 vdd.n816 99.5127
R2653 vdd.n3310 vdd.n3309 99.5127
R2654 vdd.n3307 vdd.n819 99.5127
R2655 vdd.n3303 vdd.n3302 99.5127
R2656 vdd.n3300 vdd.n3298 99.5127
R2657 vdd.n3296 vdd.n822 99.5127
R2658 vdd.n3292 vdd.n3291 99.5127
R2659 vdd.n3289 vdd.n825 99.5127
R2660 vdd.n3285 vdd.n3284 99.5127
R2661 vdd.n3282 vdd.n828 99.5127
R2662 vdd.n3278 vdd.n3277 99.5127
R2663 vdd.n3275 vdd.n831 99.5127
R2664 vdd.n3270 vdd.n3269 99.5127
R2665 vdd.n3021 vdd.n958 99.5127
R2666 vdd.n3017 vdd.n958 99.5127
R2667 vdd.n3017 vdd.n952 99.5127
R2668 vdd.n2899 vdd.n952 99.5127
R2669 vdd.n2899 vdd.n947 99.5127
R2670 vdd.n2902 vdd.n947 99.5127
R2671 vdd.n2902 vdd.n941 99.5127
R2672 vdd.n3003 vdd.n941 99.5127
R2673 vdd.n3003 vdd.n935 99.5127
R2674 vdd.n2999 vdd.n935 99.5127
R2675 vdd.n2999 vdd.n929 99.5127
R2676 vdd.n2946 vdd.n929 99.5127
R2677 vdd.n2946 vdd.n923 99.5127
R2678 vdd.n2943 vdd.n923 99.5127
R2679 vdd.n2943 vdd.n918 99.5127
R2680 vdd.n2940 vdd.n918 99.5127
R2681 vdd.n2940 vdd.n913 99.5127
R2682 vdd.n2937 vdd.n913 99.5127
R2683 vdd.n2937 vdd.n906 99.5127
R2684 vdd.n2934 vdd.n906 99.5127
R2685 vdd.n2934 vdd.n899 99.5127
R2686 vdd.n2931 vdd.n899 99.5127
R2687 vdd.n2931 vdd.n893 99.5127
R2688 vdd.n2928 vdd.n893 99.5127
R2689 vdd.n2928 vdd.n888 99.5127
R2690 vdd.n2925 vdd.n888 99.5127
R2691 vdd.n2925 vdd.n882 99.5127
R2692 vdd.n2922 vdd.n882 99.5127
R2693 vdd.n2922 vdd.n875 99.5127
R2694 vdd.n2919 vdd.n875 99.5127
R2695 vdd.n2919 vdd.n868 99.5127
R2696 vdd.n2916 vdd.n868 99.5127
R2697 vdd.n2916 vdd.n862 99.5127
R2698 vdd.n2913 vdd.n862 99.5127
R2699 vdd.n2913 vdd.n857 99.5127
R2700 vdd.n2910 vdd.n857 99.5127
R2701 vdd.n2910 vdd.n852 99.5127
R2702 vdd.n2907 vdd.n852 99.5127
R2703 vdd.n2907 vdd.n844 99.5127
R2704 vdd.n844 vdd.n837 99.5127
R2705 vdd.n3262 vdd.n837 99.5127
R2706 vdd.n3263 vdd.n3262 99.5127
R2707 vdd.n3263 vdd.n806 99.5127
R2708 vdd.n3087 vdd.n962 99.5127
R2709 vdd.n3087 vdd.n2819 99.5127
R2710 vdd.n3083 vdd.n3082 99.5127
R2711 vdd.n3079 vdd.n3078 99.5127
R2712 vdd.n3075 vdd.n3074 99.5127
R2713 vdd.n3071 vdd.n3070 99.5127
R2714 vdd.n3067 vdd.n3066 99.5127
R2715 vdd.n3063 vdd.n3062 99.5127
R2716 vdd.n3059 vdd.n3058 99.5127
R2717 vdd.n3055 vdd.n3054 99.5127
R2718 vdd.n3051 vdd.n3050 99.5127
R2719 vdd.n3047 vdd.n3046 99.5127
R2720 vdd.n3043 vdd.n3042 99.5127
R2721 vdd.n3039 vdd.n3038 99.5127
R2722 vdd.n3035 vdd.n3034 99.5127
R2723 vdd.n3031 vdd.n3030 99.5127
R2724 vdd.n3026 vdd.n3025 99.5127
R2725 vdd.n2783 vdd.n999 99.5127
R2726 vdd.n2779 vdd.n2778 99.5127
R2727 vdd.n2775 vdd.n2774 99.5127
R2728 vdd.n2771 vdd.n2770 99.5127
R2729 vdd.n2767 vdd.n2766 99.5127
R2730 vdd.n2763 vdd.n2762 99.5127
R2731 vdd.n2759 vdd.n2758 99.5127
R2732 vdd.n2755 vdd.n2754 99.5127
R2733 vdd.n2751 vdd.n2750 99.5127
R2734 vdd.n2747 vdd.n2746 99.5127
R2735 vdd.n2743 vdd.n2742 99.5127
R2736 vdd.n2739 vdd.n2738 99.5127
R2737 vdd.n2735 vdd.n2734 99.5127
R2738 vdd.n2731 vdd.n2730 99.5127
R2739 vdd.n2727 vdd.n2726 99.5127
R2740 vdd.n2723 vdd.n2722 99.5127
R2741 vdd.n2718 vdd.n2717 99.5127
R2742 vdd.n1355 vdd.n1135 99.5127
R2743 vdd.n1358 vdd.n1135 99.5127
R2744 vdd.n1358 vdd.n1129 99.5127
R2745 vdd.n1361 vdd.n1129 99.5127
R2746 vdd.n1361 vdd.n1124 99.5127
R2747 vdd.n1364 vdd.n1124 99.5127
R2748 vdd.n1364 vdd.n1117 99.5127
R2749 vdd.n1367 vdd.n1117 99.5127
R2750 vdd.n1367 vdd.n1110 99.5127
R2751 vdd.n1370 vdd.n1110 99.5127
R2752 vdd.n1370 vdd.n1104 99.5127
R2753 vdd.n1373 vdd.n1104 99.5127
R2754 vdd.n1373 vdd.n1099 99.5127
R2755 vdd.n1376 vdd.n1099 99.5127
R2756 vdd.n1376 vdd.n1094 99.5127
R2757 vdd.n1379 vdd.n1094 99.5127
R2758 vdd.n1379 vdd.n1088 99.5127
R2759 vdd.n1382 vdd.n1088 99.5127
R2760 vdd.n1382 vdd.n1081 99.5127
R2761 vdd.n1385 vdd.n1081 99.5127
R2762 vdd.n1385 vdd.n1074 99.5127
R2763 vdd.n1388 vdd.n1074 99.5127
R2764 vdd.n1388 vdd.n1068 99.5127
R2765 vdd.n1391 vdd.n1068 99.5127
R2766 vdd.n1391 vdd.n1063 99.5127
R2767 vdd.n1394 vdd.n1063 99.5127
R2768 vdd.n1394 vdd.n1057 99.5127
R2769 vdd.n1436 vdd.n1057 99.5127
R2770 vdd.n1436 vdd.n1050 99.5127
R2771 vdd.n1432 vdd.n1050 99.5127
R2772 vdd.n1432 vdd.n1044 99.5127
R2773 vdd.n1429 vdd.n1044 99.5127
R2774 vdd.n1429 vdd.n1039 99.5127
R2775 vdd.n1426 vdd.n1039 99.5127
R2776 vdd.n1426 vdd.n1034 99.5127
R2777 vdd.n1406 vdd.n1034 99.5127
R2778 vdd.n1406 vdd.n1029 99.5127
R2779 vdd.n1403 vdd.n1029 99.5127
R2780 vdd.n1403 vdd.n1022 99.5127
R2781 vdd.n1400 vdd.n1022 99.5127
R2782 vdd.n1400 vdd.n1015 99.5127
R2783 vdd.n1015 vdd.n1004 99.5127
R2784 vdd.n2713 vdd.n1004 99.5127
R2785 vdd.n2505 vdd.n1140 99.5127
R2786 vdd.n2505 vdd.n1176 99.5127
R2787 vdd.n2501 vdd.n2500 99.5127
R2788 vdd.n2497 vdd.n2496 99.5127
R2789 vdd.n2493 vdd.n2492 99.5127
R2790 vdd.n2489 vdd.n2488 99.5127
R2791 vdd.n2485 vdd.n2484 99.5127
R2792 vdd.n2481 vdd.n2480 99.5127
R2793 vdd.n2477 vdd.n2476 99.5127
R2794 vdd.n1322 vdd.n1321 99.5127
R2795 vdd.n1326 vdd.n1325 99.5127
R2796 vdd.n1330 vdd.n1329 99.5127
R2797 vdd.n1334 vdd.n1333 99.5127
R2798 vdd.n1338 vdd.n1337 99.5127
R2799 vdd.n1342 vdd.n1341 99.5127
R2800 vdd.n1346 vdd.n1345 99.5127
R2801 vdd.n1351 vdd.n1350 99.5127
R2802 vdd.n2512 vdd.n1138 99.5127
R2803 vdd.n2512 vdd.n1128 99.5127
R2804 vdd.n2520 vdd.n1128 99.5127
R2805 vdd.n2520 vdd.n1126 99.5127
R2806 vdd.n2524 vdd.n1126 99.5127
R2807 vdd.n2524 vdd.n1115 99.5127
R2808 vdd.n2532 vdd.n1115 99.5127
R2809 vdd.n2532 vdd.n1113 99.5127
R2810 vdd.n2536 vdd.n1113 99.5127
R2811 vdd.n2536 vdd.n1103 99.5127
R2812 vdd.n2544 vdd.n1103 99.5127
R2813 vdd.n2544 vdd.n1101 99.5127
R2814 vdd.n2548 vdd.n1101 99.5127
R2815 vdd.n2548 vdd.n1092 99.5127
R2816 vdd.n2556 vdd.n1092 99.5127
R2817 vdd.n2556 vdd.n1090 99.5127
R2818 vdd.n2560 vdd.n1090 99.5127
R2819 vdd.n2560 vdd.n1079 99.5127
R2820 vdd.n2568 vdd.n1079 99.5127
R2821 vdd.n2568 vdd.n1077 99.5127
R2822 vdd.n2572 vdd.n1077 99.5127
R2823 vdd.n2572 vdd.n1067 99.5127
R2824 vdd.n2581 vdd.n1067 99.5127
R2825 vdd.n2581 vdd.n1065 99.5127
R2826 vdd.n2585 vdd.n1065 99.5127
R2827 vdd.n2585 vdd.n1055 99.5127
R2828 vdd.n2593 vdd.n1055 99.5127
R2829 vdd.n2593 vdd.n1053 99.5127
R2830 vdd.n2597 vdd.n1053 99.5127
R2831 vdd.n2597 vdd.n1043 99.5127
R2832 vdd.n2605 vdd.n1043 99.5127
R2833 vdd.n2605 vdd.n1041 99.5127
R2834 vdd.n2609 vdd.n1041 99.5127
R2835 vdd.n2609 vdd.n1033 99.5127
R2836 vdd.n2617 vdd.n1033 99.5127
R2837 vdd.n2617 vdd.n1031 99.5127
R2838 vdd.n2621 vdd.n1031 99.5127
R2839 vdd.n2621 vdd.n1020 99.5127
R2840 vdd.n2631 vdd.n1020 99.5127
R2841 vdd.n2631 vdd.n1017 99.5127
R2842 vdd.n2636 vdd.n1017 99.5127
R2843 vdd.n2636 vdd.n1018 99.5127
R2844 vdd.n1018 vdd.n998 99.5127
R2845 vdd.n3246 vdd.n3245 99.5127
R2846 vdd.n3243 vdd.n3209 99.5127
R2847 vdd.n3239 vdd.n3238 99.5127
R2848 vdd.n3236 vdd.n3212 99.5127
R2849 vdd.n3232 vdd.n3231 99.5127
R2850 vdd.n3229 vdd.n3215 99.5127
R2851 vdd.n3225 vdd.n3224 99.5127
R2852 vdd.n3222 vdd.n3219 99.5127
R2853 vdd.n3363 vdd.n787 99.5127
R2854 vdd.n3361 vdd.n3360 99.5127
R2855 vdd.n3358 vdd.n789 99.5127
R2856 vdd.n3354 vdd.n3353 99.5127
R2857 vdd.n3351 vdd.n792 99.5127
R2858 vdd.n3347 vdd.n3346 99.5127
R2859 vdd.n3344 vdd.n795 99.5127
R2860 vdd.n3340 vdd.n3339 99.5127
R2861 vdd.n3337 vdd.n798 99.5127
R2862 vdd.n2895 vdd.n959 99.5127
R2863 vdd.n3015 vdd.n959 99.5127
R2864 vdd.n3015 vdd.n953 99.5127
R2865 vdd.n3011 vdd.n953 99.5127
R2866 vdd.n3011 vdd.n948 99.5127
R2867 vdd.n3008 vdd.n948 99.5127
R2868 vdd.n3008 vdd.n942 99.5127
R2869 vdd.n3005 vdd.n942 99.5127
R2870 vdd.n3005 vdd.n936 99.5127
R2871 vdd.n2997 vdd.n936 99.5127
R2872 vdd.n2997 vdd.n930 99.5127
R2873 vdd.n2993 vdd.n930 99.5127
R2874 vdd.n2993 vdd.n924 99.5127
R2875 vdd.n2990 vdd.n924 99.5127
R2876 vdd.n2990 vdd.n919 99.5127
R2877 vdd.n2987 vdd.n919 99.5127
R2878 vdd.n2987 vdd.n914 99.5127
R2879 vdd.n2984 vdd.n914 99.5127
R2880 vdd.n2984 vdd.n907 99.5127
R2881 vdd.n2981 vdd.n907 99.5127
R2882 vdd.n2981 vdd.n900 99.5127
R2883 vdd.n2978 vdd.n900 99.5127
R2884 vdd.n2978 vdd.n894 99.5127
R2885 vdd.n2975 vdd.n894 99.5127
R2886 vdd.n2975 vdd.n889 99.5127
R2887 vdd.n2972 vdd.n889 99.5127
R2888 vdd.n2972 vdd.n883 99.5127
R2889 vdd.n2969 vdd.n883 99.5127
R2890 vdd.n2969 vdd.n876 99.5127
R2891 vdd.n2966 vdd.n876 99.5127
R2892 vdd.n2966 vdd.n869 99.5127
R2893 vdd.n2963 vdd.n869 99.5127
R2894 vdd.n2963 vdd.n863 99.5127
R2895 vdd.n2960 vdd.n863 99.5127
R2896 vdd.n2960 vdd.n858 99.5127
R2897 vdd.n2957 vdd.n858 99.5127
R2898 vdd.n2957 vdd.n853 99.5127
R2899 vdd.n2954 vdd.n853 99.5127
R2900 vdd.n2954 vdd.n845 99.5127
R2901 vdd.n2951 vdd.n845 99.5127
R2902 vdd.n2951 vdd.n838 99.5127
R2903 vdd.n838 vdd.n804 99.5127
R2904 vdd.n3332 vdd.n804 99.5127
R2905 vdd.n2830 vdd.n2829 99.5127
R2906 vdd.n2834 vdd.n2833 99.5127
R2907 vdd.n2838 vdd.n2837 99.5127
R2908 vdd.n2842 vdd.n2841 99.5127
R2909 vdd.n2846 vdd.n2845 99.5127
R2910 vdd.n2850 vdd.n2849 99.5127
R2911 vdd.n2854 vdd.n2853 99.5127
R2912 vdd.n2858 vdd.n2857 99.5127
R2913 vdd.n2862 vdd.n2861 99.5127
R2914 vdd.n2866 vdd.n2865 99.5127
R2915 vdd.n2870 vdd.n2869 99.5127
R2916 vdd.n2874 vdd.n2873 99.5127
R2917 vdd.n2878 vdd.n2877 99.5127
R2918 vdd.n2882 vdd.n2881 99.5127
R2919 vdd.n2886 vdd.n2885 99.5127
R2920 vdd.n2890 vdd.n2889 99.5127
R2921 vdd.n2892 vdd.n2818 99.5127
R2922 vdd.n3096 vdd.n956 99.5127
R2923 vdd.n3096 vdd.n954 99.5127
R2924 vdd.n3100 vdd.n954 99.5127
R2925 vdd.n3100 vdd.n945 99.5127
R2926 vdd.n3108 vdd.n945 99.5127
R2927 vdd.n3108 vdd.n943 99.5127
R2928 vdd.n3112 vdd.n943 99.5127
R2929 vdd.n3112 vdd.n934 99.5127
R2930 vdd.n3120 vdd.n934 99.5127
R2931 vdd.n3120 vdd.n932 99.5127
R2932 vdd.n3124 vdd.n932 99.5127
R2933 vdd.n3124 vdd.n922 99.5127
R2934 vdd.n3132 vdd.n922 99.5127
R2935 vdd.n3132 vdd.n920 99.5127
R2936 vdd.n3136 vdd.n920 99.5127
R2937 vdd.n3136 vdd.n911 99.5127
R2938 vdd.n3144 vdd.n911 99.5127
R2939 vdd.n3144 vdd.n909 99.5127
R2940 vdd.n3149 vdd.n909 99.5127
R2941 vdd.n3149 vdd.n898 99.5127
R2942 vdd.n3157 vdd.n898 99.5127
R2943 vdd.n3157 vdd.n895 99.5127
R2944 vdd.n3161 vdd.n895 99.5127
R2945 vdd.n3161 vdd.n886 99.5127
R2946 vdd.n3169 vdd.n886 99.5127
R2947 vdd.n3169 vdd.n884 99.5127
R2948 vdd.n3173 vdd.n884 99.5127
R2949 vdd.n3173 vdd.n873 99.5127
R2950 vdd.n3181 vdd.n873 99.5127
R2951 vdd.n3181 vdd.n871 99.5127
R2952 vdd.n3185 vdd.n871 99.5127
R2953 vdd.n3185 vdd.n861 99.5127
R2954 vdd.n3193 vdd.n861 99.5127
R2955 vdd.n3193 vdd.n859 99.5127
R2956 vdd.n3197 vdd.n859 99.5127
R2957 vdd.n3197 vdd.n850 99.5127
R2958 vdd.n3205 vdd.n850 99.5127
R2959 vdd.n3205 vdd.n847 99.5127
R2960 vdd.n3254 vdd.n847 99.5127
R2961 vdd.n3254 vdd.n848 99.5127
R2962 vdd.n848 vdd.n839 99.5127
R2963 vdd.n3249 vdd.n839 99.5127
R2964 vdd.n3249 vdd.n807 99.5127
R2965 vdd.n2707 vdd.n2706 99.5127
R2966 vdd.n2703 vdd.n2702 99.5127
R2967 vdd.n2699 vdd.n2698 99.5127
R2968 vdd.n2695 vdd.n2694 99.5127
R2969 vdd.n2691 vdd.n2690 99.5127
R2970 vdd.n2687 vdd.n2686 99.5127
R2971 vdd.n2683 vdd.n2682 99.5127
R2972 vdd.n2679 vdd.n2678 99.5127
R2973 vdd.n2675 vdd.n2674 99.5127
R2974 vdd.n2671 vdd.n2670 99.5127
R2975 vdd.n2667 vdd.n2666 99.5127
R2976 vdd.n2663 vdd.n2662 99.5127
R2977 vdd.n2659 vdd.n2658 99.5127
R2978 vdd.n2655 vdd.n2654 99.5127
R2979 vdd.n2651 vdd.n2650 99.5127
R2980 vdd.n2647 vdd.n2646 99.5127
R2981 vdd.n2643 vdd.n980 99.5127
R2982 vdd.n1480 vdd.n1136 99.5127
R2983 vdd.n1477 vdd.n1136 99.5127
R2984 vdd.n1477 vdd.n1130 99.5127
R2985 vdd.n1474 vdd.n1130 99.5127
R2986 vdd.n1474 vdd.n1125 99.5127
R2987 vdd.n1471 vdd.n1125 99.5127
R2988 vdd.n1471 vdd.n1118 99.5127
R2989 vdd.n1468 vdd.n1118 99.5127
R2990 vdd.n1468 vdd.n1111 99.5127
R2991 vdd.n1465 vdd.n1111 99.5127
R2992 vdd.n1465 vdd.n1105 99.5127
R2993 vdd.n1462 vdd.n1105 99.5127
R2994 vdd.n1462 vdd.n1100 99.5127
R2995 vdd.n1459 vdd.n1100 99.5127
R2996 vdd.n1459 vdd.n1095 99.5127
R2997 vdd.n1456 vdd.n1095 99.5127
R2998 vdd.n1456 vdd.n1089 99.5127
R2999 vdd.n1453 vdd.n1089 99.5127
R3000 vdd.n1453 vdd.n1082 99.5127
R3001 vdd.n1450 vdd.n1082 99.5127
R3002 vdd.n1450 vdd.n1075 99.5127
R3003 vdd.n1447 vdd.n1075 99.5127
R3004 vdd.n1447 vdd.n1069 99.5127
R3005 vdd.n1444 vdd.n1069 99.5127
R3006 vdd.n1444 vdd.n1064 99.5127
R3007 vdd.n1441 vdd.n1064 99.5127
R3008 vdd.n1441 vdd.n1058 99.5127
R3009 vdd.n1438 vdd.n1058 99.5127
R3010 vdd.n1438 vdd.n1051 99.5127
R3011 vdd.n1409 vdd.n1051 99.5127
R3012 vdd.n1409 vdd.n1045 99.5127
R3013 vdd.n1412 vdd.n1045 99.5127
R3014 vdd.n1412 vdd.n1040 99.5127
R3015 vdd.n1424 vdd.n1040 99.5127
R3016 vdd.n1424 vdd.n1035 99.5127
R3017 vdd.n1420 vdd.n1035 99.5127
R3018 vdd.n1420 vdd.n1030 99.5127
R3019 vdd.n1417 vdd.n1030 99.5127
R3020 vdd.n1417 vdd.n1023 99.5127
R3021 vdd.n1023 vdd.n1014 99.5127
R3022 vdd.n2638 vdd.n1014 99.5127
R3023 vdd.n2639 vdd.n2638 99.5127
R3024 vdd.n2639 vdd.n1006 99.5127
R3025 vdd.n1284 vdd.n1283 99.5127
R3026 vdd.n1288 vdd.n1287 99.5127
R3027 vdd.n1292 vdd.n1291 99.5127
R3028 vdd.n1296 vdd.n1295 99.5127
R3029 vdd.n1300 vdd.n1299 99.5127
R3030 vdd.n1304 vdd.n1303 99.5127
R3031 vdd.n1308 vdd.n1307 99.5127
R3032 vdd.n1312 vdd.n1311 99.5127
R3033 vdd.n1513 vdd.n1314 99.5127
R3034 vdd.n1511 vdd.n1510 99.5127
R3035 vdd.n1507 vdd.n1506 99.5127
R3036 vdd.n1503 vdd.n1502 99.5127
R3037 vdd.n1499 vdd.n1498 99.5127
R3038 vdd.n1495 vdd.n1494 99.5127
R3039 vdd.n1491 vdd.n1490 99.5127
R3040 vdd.n1487 vdd.n1486 99.5127
R3041 vdd.n1483 vdd.n1175 99.5127
R3042 vdd.n2514 vdd.n1133 99.5127
R3043 vdd.n2514 vdd.n1131 99.5127
R3044 vdd.n2518 vdd.n1131 99.5127
R3045 vdd.n2518 vdd.n1122 99.5127
R3046 vdd.n2526 vdd.n1122 99.5127
R3047 vdd.n2526 vdd.n1120 99.5127
R3048 vdd.n2530 vdd.n1120 99.5127
R3049 vdd.n2530 vdd.n1109 99.5127
R3050 vdd.n2538 vdd.n1109 99.5127
R3051 vdd.n2538 vdd.n1107 99.5127
R3052 vdd.n2542 vdd.n1107 99.5127
R3053 vdd.n2542 vdd.n1098 99.5127
R3054 vdd.n2550 vdd.n1098 99.5127
R3055 vdd.n2550 vdd.n1096 99.5127
R3056 vdd.n2554 vdd.n1096 99.5127
R3057 vdd.n2554 vdd.n1086 99.5127
R3058 vdd.n2562 vdd.n1086 99.5127
R3059 vdd.n2562 vdd.n1084 99.5127
R3060 vdd.n2566 vdd.n1084 99.5127
R3061 vdd.n2566 vdd.n1073 99.5127
R3062 vdd.n2574 vdd.n1073 99.5127
R3063 vdd.n2574 vdd.n1070 99.5127
R3064 vdd.n2579 vdd.n1070 99.5127
R3065 vdd.n2579 vdd.n1061 99.5127
R3066 vdd.n2587 vdd.n1061 99.5127
R3067 vdd.n2587 vdd.n1059 99.5127
R3068 vdd.n2591 vdd.n1059 99.5127
R3069 vdd.n2591 vdd.n1049 99.5127
R3070 vdd.n2599 vdd.n1049 99.5127
R3071 vdd.n2599 vdd.n1047 99.5127
R3072 vdd.n2603 vdd.n1047 99.5127
R3073 vdd.n2603 vdd.n1038 99.5127
R3074 vdd.n2611 vdd.n1038 99.5127
R3075 vdd.n2611 vdd.n1036 99.5127
R3076 vdd.n2615 vdd.n1036 99.5127
R3077 vdd.n2615 vdd.n1027 99.5127
R3078 vdd.n2623 vdd.n1027 99.5127
R3079 vdd.n2623 vdd.n1024 99.5127
R3080 vdd.n2629 vdd.n1024 99.5127
R3081 vdd.n2629 vdd.n1025 99.5127
R3082 vdd.n1025 vdd.n1016 99.5127
R3083 vdd.n1016 vdd.n1007 99.5127
R3084 vdd.n2711 vdd.n1007 99.5127
R3085 vdd.n9 vdd.n7 98.9633
R3086 vdd.n2 vdd.n0 98.9633
R3087 vdd.n9 vdd.n8 98.6055
R3088 vdd.n11 vdd.n10 98.6055
R3089 vdd.n13 vdd.n12 98.6055
R3090 vdd.n6 vdd.n5 98.6055
R3091 vdd.n4 vdd.n3 98.6055
R3092 vdd.n2 vdd.n1 98.6055
R3093 vdd.t71 vdd.n303 85.8723
R3094 vdd.t93 vdd.n244 85.8723
R3095 vdd.t137 vdd.n201 85.8723
R3096 vdd.t145 vdd.n142 85.8723
R3097 vdd.t144 vdd.n100 85.8723
R3098 vdd.t38 vdd.n41 85.8723
R3099 vdd.t304 vdd.n2177 85.8723
R3100 vdd.t67 vdd.n2236 85.8723
R3101 vdd.t58 vdd.n2075 85.8723
R3102 vdd.t286 vdd.n2134 85.8723
R3103 vdd.t12 vdd.n1974 85.8723
R3104 vdd.t116 vdd.n2033 85.8723
R3105 vdd.n897 vdd.n896 78.546
R3106 vdd.n2577 vdd.n1071 78.546
R3107 vdd.n290 vdd.n289 75.1835
R3108 vdd.n288 vdd.n287 75.1835
R3109 vdd.n286 vdd.n285 75.1835
R3110 vdd.n284 vdd.n283 75.1835
R3111 vdd.n282 vdd.n281 75.1835
R3112 vdd.n280 vdd.n279 75.1835
R3113 vdd.n278 vdd.n277 75.1835
R3114 vdd.n276 vdd.n275 75.1835
R3115 vdd.n274 vdd.n273 75.1835
R3116 vdd.n188 vdd.n187 75.1835
R3117 vdd.n186 vdd.n185 75.1835
R3118 vdd.n184 vdd.n183 75.1835
R3119 vdd.n182 vdd.n181 75.1835
R3120 vdd.n180 vdd.n179 75.1835
R3121 vdd.n178 vdd.n177 75.1835
R3122 vdd.n176 vdd.n175 75.1835
R3123 vdd.n174 vdd.n173 75.1835
R3124 vdd.n172 vdd.n171 75.1835
R3125 vdd.n87 vdd.n86 75.1835
R3126 vdd.n85 vdd.n84 75.1835
R3127 vdd.n83 vdd.n82 75.1835
R3128 vdd.n81 vdd.n80 75.1835
R3129 vdd.n79 vdd.n78 75.1835
R3130 vdd.n77 vdd.n76 75.1835
R3131 vdd.n75 vdd.n74 75.1835
R3132 vdd.n73 vdd.n72 75.1835
R3133 vdd.n71 vdd.n70 75.1835
R3134 vdd.n2207 vdd.n2206 75.1835
R3135 vdd.n2209 vdd.n2208 75.1835
R3136 vdd.n2211 vdd.n2210 75.1835
R3137 vdd.n2213 vdd.n2212 75.1835
R3138 vdd.n2215 vdd.n2214 75.1835
R3139 vdd.n2217 vdd.n2216 75.1835
R3140 vdd.n2219 vdd.n2218 75.1835
R3141 vdd.n2221 vdd.n2220 75.1835
R3142 vdd.n2223 vdd.n2222 75.1835
R3143 vdd.n2105 vdd.n2104 75.1835
R3144 vdd.n2107 vdd.n2106 75.1835
R3145 vdd.n2109 vdd.n2108 75.1835
R3146 vdd.n2111 vdd.n2110 75.1835
R3147 vdd.n2113 vdd.n2112 75.1835
R3148 vdd.n2115 vdd.n2114 75.1835
R3149 vdd.n2117 vdd.n2116 75.1835
R3150 vdd.n2119 vdd.n2118 75.1835
R3151 vdd.n2121 vdd.n2120 75.1835
R3152 vdd.n2004 vdd.n2003 75.1835
R3153 vdd.n2006 vdd.n2005 75.1835
R3154 vdd.n2008 vdd.n2007 75.1835
R3155 vdd.n2010 vdd.n2009 75.1835
R3156 vdd.n2012 vdd.n2011 75.1835
R3157 vdd.n2014 vdd.n2013 75.1835
R3158 vdd.n2016 vdd.n2015 75.1835
R3159 vdd.n2018 vdd.n2017 75.1835
R3160 vdd.n2020 vdd.n2019 75.1835
R3161 vdd.n3088 vdd.n2801 72.8958
R3162 vdd.n3088 vdd.n2802 72.8958
R3163 vdd.n3088 vdd.n2803 72.8958
R3164 vdd.n3088 vdd.n2804 72.8958
R3165 vdd.n3088 vdd.n2805 72.8958
R3166 vdd.n3088 vdd.n2806 72.8958
R3167 vdd.n3088 vdd.n2807 72.8958
R3168 vdd.n3088 vdd.n2808 72.8958
R3169 vdd.n3088 vdd.n2809 72.8958
R3170 vdd.n3088 vdd.n2810 72.8958
R3171 vdd.n3088 vdd.n2811 72.8958
R3172 vdd.n3088 vdd.n2812 72.8958
R3173 vdd.n3088 vdd.n2813 72.8958
R3174 vdd.n3088 vdd.n2814 72.8958
R3175 vdd.n3088 vdd.n2815 72.8958
R3176 vdd.n3088 vdd.n2816 72.8958
R3177 vdd.n3088 vdd.n2817 72.8958
R3178 vdd.n803 vdd.n692 72.8958
R3179 vdd.n3338 vdd.n692 72.8958
R3180 vdd.n797 vdd.n692 72.8958
R3181 vdd.n3345 vdd.n692 72.8958
R3182 vdd.n794 vdd.n692 72.8958
R3183 vdd.n3352 vdd.n692 72.8958
R3184 vdd.n791 vdd.n692 72.8958
R3185 vdd.n3359 vdd.n692 72.8958
R3186 vdd.n3362 vdd.n692 72.8958
R3187 vdd.n3218 vdd.n692 72.8958
R3188 vdd.n3223 vdd.n692 72.8958
R3189 vdd.n3217 vdd.n692 72.8958
R3190 vdd.n3230 vdd.n692 72.8958
R3191 vdd.n3214 vdd.n692 72.8958
R3192 vdd.n3237 vdd.n692 72.8958
R3193 vdd.n3211 vdd.n692 72.8958
R3194 vdd.n3244 vdd.n692 72.8958
R3195 vdd.n2507 vdd.n2506 72.8958
R3196 vdd.n2506 vdd.n1142 72.8958
R3197 vdd.n2506 vdd.n1143 72.8958
R3198 vdd.n2506 vdd.n1144 72.8958
R3199 vdd.n2506 vdd.n1145 72.8958
R3200 vdd.n2506 vdd.n1146 72.8958
R3201 vdd.n2506 vdd.n1147 72.8958
R3202 vdd.n2506 vdd.n1148 72.8958
R3203 vdd.n2506 vdd.n1149 72.8958
R3204 vdd.n2506 vdd.n1150 72.8958
R3205 vdd.n2506 vdd.n1151 72.8958
R3206 vdd.n2506 vdd.n1152 72.8958
R3207 vdd.n2506 vdd.n1153 72.8958
R3208 vdd.n2506 vdd.n1154 72.8958
R3209 vdd.n2506 vdd.n1155 72.8958
R3210 vdd.n2506 vdd.n1156 72.8958
R3211 vdd.n2506 vdd.n1157 72.8958
R3212 vdd.n2784 vdd.n981 72.8958
R3213 vdd.n2784 vdd.n982 72.8958
R3214 vdd.n2784 vdd.n983 72.8958
R3215 vdd.n2784 vdd.n984 72.8958
R3216 vdd.n2784 vdd.n985 72.8958
R3217 vdd.n2784 vdd.n986 72.8958
R3218 vdd.n2784 vdd.n987 72.8958
R3219 vdd.n2784 vdd.n988 72.8958
R3220 vdd.n2784 vdd.n989 72.8958
R3221 vdd.n2784 vdd.n990 72.8958
R3222 vdd.n2784 vdd.n991 72.8958
R3223 vdd.n2784 vdd.n992 72.8958
R3224 vdd.n2784 vdd.n993 72.8958
R3225 vdd.n2784 vdd.n994 72.8958
R3226 vdd.n2784 vdd.n995 72.8958
R3227 vdd.n2784 vdd.n996 72.8958
R3228 vdd.n2784 vdd.n997 72.8958
R3229 vdd.n3089 vdd.n3088 72.8958
R3230 vdd.n3088 vdd.n2785 72.8958
R3231 vdd.n3088 vdd.n2786 72.8958
R3232 vdd.n3088 vdd.n2787 72.8958
R3233 vdd.n3088 vdd.n2788 72.8958
R3234 vdd.n3088 vdd.n2789 72.8958
R3235 vdd.n3088 vdd.n2790 72.8958
R3236 vdd.n3088 vdd.n2791 72.8958
R3237 vdd.n3088 vdd.n2792 72.8958
R3238 vdd.n3088 vdd.n2793 72.8958
R3239 vdd.n3088 vdd.n2794 72.8958
R3240 vdd.n3088 vdd.n2795 72.8958
R3241 vdd.n3088 vdd.n2796 72.8958
R3242 vdd.n3088 vdd.n2797 72.8958
R3243 vdd.n3088 vdd.n2798 72.8958
R3244 vdd.n3088 vdd.n2799 72.8958
R3245 vdd.n3088 vdd.n2800 72.8958
R3246 vdd.n3268 vdd.n692 72.8958
R3247 vdd.n835 vdd.n692 72.8958
R3248 vdd.n3276 vdd.n692 72.8958
R3249 vdd.n830 vdd.n692 72.8958
R3250 vdd.n3283 vdd.n692 72.8958
R3251 vdd.n827 vdd.n692 72.8958
R3252 vdd.n3290 vdd.n692 72.8958
R3253 vdd.n824 vdd.n692 72.8958
R3254 vdd.n3297 vdd.n692 72.8958
R3255 vdd.n3301 vdd.n692 72.8958
R3256 vdd.n821 vdd.n692 72.8958
R3257 vdd.n3308 vdd.n692 72.8958
R3258 vdd.n818 vdd.n692 72.8958
R3259 vdd.n3315 vdd.n692 72.8958
R3260 vdd.n815 vdd.n692 72.8958
R3261 vdd.n3322 vdd.n692 72.8958
R3262 vdd.n3325 vdd.n692 72.8958
R3263 vdd.n2784 vdd.n979 72.8958
R3264 vdd.n2784 vdd.n978 72.8958
R3265 vdd.n2784 vdd.n977 72.8958
R3266 vdd.n2784 vdd.n976 72.8958
R3267 vdd.n2784 vdd.n975 72.8958
R3268 vdd.n2784 vdd.n974 72.8958
R3269 vdd.n2784 vdd.n973 72.8958
R3270 vdd.n2784 vdd.n972 72.8958
R3271 vdd.n2784 vdd.n971 72.8958
R3272 vdd.n2784 vdd.n970 72.8958
R3273 vdd.n2784 vdd.n969 72.8958
R3274 vdd.n2784 vdd.n968 72.8958
R3275 vdd.n2784 vdd.n967 72.8958
R3276 vdd.n2784 vdd.n966 72.8958
R3277 vdd.n2784 vdd.n965 72.8958
R3278 vdd.n2784 vdd.n964 72.8958
R3279 vdd.n2784 vdd.n963 72.8958
R3280 vdd.n2506 vdd.n1158 72.8958
R3281 vdd.n2506 vdd.n1159 72.8958
R3282 vdd.n2506 vdd.n1160 72.8958
R3283 vdd.n2506 vdd.n1161 72.8958
R3284 vdd.n2506 vdd.n1162 72.8958
R3285 vdd.n2506 vdd.n1163 72.8958
R3286 vdd.n2506 vdd.n1164 72.8958
R3287 vdd.n2506 vdd.n1165 72.8958
R3288 vdd.n2506 vdd.n1166 72.8958
R3289 vdd.n2506 vdd.n1167 72.8958
R3290 vdd.n2506 vdd.n1168 72.8958
R3291 vdd.n2506 vdd.n1169 72.8958
R3292 vdd.n2506 vdd.n1170 72.8958
R3293 vdd.n2506 vdd.n1171 72.8958
R3294 vdd.n2506 vdd.n1172 72.8958
R3295 vdd.n2506 vdd.n1173 72.8958
R3296 vdd.n2506 vdd.n1174 72.8958
R3297 vdd.n1874 vdd.n1873 66.2847
R3298 vdd.n1873 vdd.n1649 66.2847
R3299 vdd.n1873 vdd.n1650 66.2847
R3300 vdd.n1873 vdd.n1651 66.2847
R3301 vdd.n1873 vdd.n1652 66.2847
R3302 vdd.n1873 vdd.n1653 66.2847
R3303 vdd.n1873 vdd.n1654 66.2847
R3304 vdd.n1873 vdd.n1655 66.2847
R3305 vdd.n1873 vdd.n1656 66.2847
R3306 vdd.n1873 vdd.n1657 66.2847
R3307 vdd.n1873 vdd.n1658 66.2847
R3308 vdd.n1873 vdd.n1659 66.2847
R3309 vdd.n1873 vdd.n1660 66.2847
R3310 vdd.n1873 vdd.n1661 66.2847
R3311 vdd.n1873 vdd.n1662 66.2847
R3312 vdd.n1873 vdd.n1663 66.2847
R3313 vdd.n1873 vdd.n1664 66.2847
R3314 vdd.n1873 vdd.n1665 66.2847
R3315 vdd.n1873 vdd.n1666 66.2847
R3316 vdd.n1873 vdd.n1667 66.2847
R3317 vdd.n1873 vdd.n1668 66.2847
R3318 vdd.n1873 vdd.n1669 66.2847
R3319 vdd.n1873 vdd.n1670 66.2847
R3320 vdd.n1873 vdd.n1671 66.2847
R3321 vdd.n1873 vdd.n1672 66.2847
R3322 vdd.n1873 vdd.n1673 66.2847
R3323 vdd.n1873 vdd.n1674 66.2847
R3324 vdd.n1873 vdd.n1675 66.2847
R3325 vdd.n1873 vdd.n1676 66.2847
R3326 vdd.n1873 vdd.n1677 66.2847
R3327 vdd.n1873 vdd.n1678 66.2847
R3328 vdd.n1526 vdd.n1141 66.2847
R3329 vdd.n1523 vdd.n1141 66.2847
R3330 vdd.n1519 vdd.n1141 66.2847
R3331 vdd.n2372 vdd.n1141 66.2847
R3332 vdd.n1275 vdd.n1141 66.2847
R3333 vdd.n2379 vdd.n1141 66.2847
R3334 vdd.n1268 vdd.n1141 66.2847
R3335 vdd.n2386 vdd.n1141 66.2847
R3336 vdd.n1261 vdd.n1141 66.2847
R3337 vdd.n2393 vdd.n1141 66.2847
R3338 vdd.n1255 vdd.n1141 66.2847
R3339 vdd.n1250 vdd.n1141 66.2847
R3340 vdd.n2404 vdd.n1141 66.2847
R3341 vdd.n1242 vdd.n1141 66.2847
R3342 vdd.n2411 vdd.n1141 66.2847
R3343 vdd.n1235 vdd.n1141 66.2847
R3344 vdd.n2418 vdd.n1141 66.2847
R3345 vdd.n1228 vdd.n1141 66.2847
R3346 vdd.n2425 vdd.n1141 66.2847
R3347 vdd.n1221 vdd.n1141 66.2847
R3348 vdd.n2432 vdd.n1141 66.2847
R3349 vdd.n1215 vdd.n1141 66.2847
R3350 vdd.n1210 vdd.n1141 66.2847
R3351 vdd.n2443 vdd.n1141 66.2847
R3352 vdd.n1202 vdd.n1141 66.2847
R3353 vdd.n2450 vdd.n1141 66.2847
R3354 vdd.n1195 vdd.n1141 66.2847
R3355 vdd.n2457 vdd.n1141 66.2847
R3356 vdd.n1188 vdd.n1141 66.2847
R3357 vdd.n2464 vdd.n1141 66.2847
R3358 vdd.n2469 vdd.n1141 66.2847
R3359 vdd.n1184 vdd.n1141 66.2847
R3360 vdd.n3495 vdd.n3494 66.2847
R3361 vdd.n3495 vdd.n693 66.2847
R3362 vdd.n3495 vdd.n694 66.2847
R3363 vdd.n3495 vdd.n695 66.2847
R3364 vdd.n3495 vdd.n696 66.2847
R3365 vdd.n3495 vdd.n697 66.2847
R3366 vdd.n3495 vdd.n698 66.2847
R3367 vdd.n3495 vdd.n699 66.2847
R3368 vdd.n3495 vdd.n700 66.2847
R3369 vdd.n3495 vdd.n701 66.2847
R3370 vdd.n3495 vdd.n702 66.2847
R3371 vdd.n3495 vdd.n703 66.2847
R3372 vdd.n3495 vdd.n704 66.2847
R3373 vdd.n3495 vdd.n705 66.2847
R3374 vdd.n3495 vdd.n706 66.2847
R3375 vdd.n3495 vdd.n707 66.2847
R3376 vdd.n3495 vdd.n708 66.2847
R3377 vdd.n3495 vdd.n709 66.2847
R3378 vdd.n3495 vdd.n710 66.2847
R3379 vdd.n3495 vdd.n711 66.2847
R3380 vdd.n3495 vdd.n712 66.2847
R3381 vdd.n3495 vdd.n713 66.2847
R3382 vdd.n3495 vdd.n714 66.2847
R3383 vdd.n3495 vdd.n715 66.2847
R3384 vdd.n3495 vdd.n716 66.2847
R3385 vdd.n3495 vdd.n717 66.2847
R3386 vdd.n3495 vdd.n718 66.2847
R3387 vdd.n3495 vdd.n719 66.2847
R3388 vdd.n3495 vdd.n720 66.2847
R3389 vdd.n3495 vdd.n721 66.2847
R3390 vdd.n3495 vdd.n722 66.2847
R3391 vdd.n3626 vdd.n3625 66.2847
R3392 vdd.n3626 vdd.n424 66.2847
R3393 vdd.n3626 vdd.n423 66.2847
R3394 vdd.n3626 vdd.n422 66.2847
R3395 vdd.n3626 vdd.n421 66.2847
R3396 vdd.n3626 vdd.n420 66.2847
R3397 vdd.n3626 vdd.n419 66.2847
R3398 vdd.n3626 vdd.n418 66.2847
R3399 vdd.n3626 vdd.n417 66.2847
R3400 vdd.n3626 vdd.n416 66.2847
R3401 vdd.n3626 vdd.n415 66.2847
R3402 vdd.n3626 vdd.n414 66.2847
R3403 vdd.n3626 vdd.n413 66.2847
R3404 vdd.n3626 vdd.n412 66.2847
R3405 vdd.n3626 vdd.n411 66.2847
R3406 vdd.n3626 vdd.n410 66.2847
R3407 vdd.n3626 vdd.n409 66.2847
R3408 vdd.n3626 vdd.n408 66.2847
R3409 vdd.n3626 vdd.n407 66.2847
R3410 vdd.n3626 vdd.n406 66.2847
R3411 vdd.n3626 vdd.n405 66.2847
R3412 vdd.n3626 vdd.n404 66.2847
R3413 vdd.n3626 vdd.n403 66.2847
R3414 vdd.n3626 vdd.n402 66.2847
R3415 vdd.n3626 vdd.n401 66.2847
R3416 vdd.n3626 vdd.n400 66.2847
R3417 vdd.n3626 vdd.n399 66.2847
R3418 vdd.n3626 vdd.n398 66.2847
R3419 vdd.n3626 vdd.n397 66.2847
R3420 vdd.n3626 vdd.n396 66.2847
R3421 vdd.n3626 vdd.n395 66.2847
R3422 vdd.n3626 vdd.n394 66.2847
R3423 vdd.n467 vdd.n394 52.4337
R3424 vdd.n473 vdd.n395 52.4337
R3425 vdd.n477 vdd.n396 52.4337
R3426 vdd.n483 vdd.n397 52.4337
R3427 vdd.n487 vdd.n398 52.4337
R3428 vdd.n493 vdd.n399 52.4337
R3429 vdd.n497 vdd.n400 52.4337
R3430 vdd.n503 vdd.n401 52.4337
R3431 vdd.n507 vdd.n402 52.4337
R3432 vdd.n513 vdd.n403 52.4337
R3433 vdd.n517 vdd.n404 52.4337
R3434 vdd.n523 vdd.n405 52.4337
R3435 vdd.n527 vdd.n406 52.4337
R3436 vdd.n533 vdd.n407 52.4337
R3437 vdd.n537 vdd.n408 52.4337
R3438 vdd.n543 vdd.n409 52.4337
R3439 vdd.n547 vdd.n410 52.4337
R3440 vdd.n553 vdd.n411 52.4337
R3441 vdd.n557 vdd.n412 52.4337
R3442 vdd.n563 vdd.n413 52.4337
R3443 vdd.n567 vdd.n414 52.4337
R3444 vdd.n573 vdd.n415 52.4337
R3445 vdd.n577 vdd.n416 52.4337
R3446 vdd.n583 vdd.n417 52.4337
R3447 vdd.n587 vdd.n418 52.4337
R3448 vdd.n593 vdd.n419 52.4337
R3449 vdd.n597 vdd.n420 52.4337
R3450 vdd.n603 vdd.n421 52.4337
R3451 vdd.n607 vdd.n422 52.4337
R3452 vdd.n613 vdd.n423 52.4337
R3453 vdd.n616 vdd.n424 52.4337
R3454 vdd.n3625 vdd.n3624 52.4337
R3455 vdd.n3494 vdd.n3493 52.4337
R3456 vdd.n728 vdd.n693 52.4337
R3457 vdd.n734 vdd.n694 52.4337
R3458 vdd.n3483 vdd.n695 52.4337
R3459 vdd.n3479 vdd.n696 52.4337
R3460 vdd.n3475 vdd.n697 52.4337
R3461 vdd.n3471 vdd.n698 52.4337
R3462 vdd.n3467 vdd.n699 52.4337
R3463 vdd.n3463 vdd.n700 52.4337
R3464 vdd.n3459 vdd.n701 52.4337
R3465 vdd.n3451 vdd.n702 52.4337
R3466 vdd.n3447 vdd.n703 52.4337
R3467 vdd.n3443 vdd.n704 52.4337
R3468 vdd.n3439 vdd.n705 52.4337
R3469 vdd.n3435 vdd.n706 52.4337
R3470 vdd.n3431 vdd.n707 52.4337
R3471 vdd.n3427 vdd.n708 52.4337
R3472 vdd.n3423 vdd.n709 52.4337
R3473 vdd.n3419 vdd.n710 52.4337
R3474 vdd.n3415 vdd.n711 52.4337
R3475 vdd.n3411 vdd.n712 52.4337
R3476 vdd.n3405 vdd.n713 52.4337
R3477 vdd.n3401 vdd.n714 52.4337
R3478 vdd.n3397 vdd.n715 52.4337
R3479 vdd.n3393 vdd.n716 52.4337
R3480 vdd.n3389 vdd.n717 52.4337
R3481 vdd.n3385 vdd.n718 52.4337
R3482 vdd.n3381 vdd.n719 52.4337
R3483 vdd.n3377 vdd.n720 52.4337
R3484 vdd.n3373 vdd.n721 52.4337
R3485 vdd.n3369 vdd.n722 52.4337
R3486 vdd.n2471 vdd.n1184 52.4337
R3487 vdd.n2469 vdd.n2468 52.4337
R3488 vdd.n2464 vdd.n2463 52.4337
R3489 vdd.n2459 vdd.n1188 52.4337
R3490 vdd.n2457 vdd.n2456 52.4337
R3491 vdd.n2452 vdd.n1195 52.4337
R3492 vdd.n2450 vdd.n2449 52.4337
R3493 vdd.n2445 vdd.n1202 52.4337
R3494 vdd.n2443 vdd.n2442 52.4337
R3495 vdd.n1211 vdd.n1210 52.4337
R3496 vdd.n2434 vdd.n1215 52.4337
R3497 vdd.n2432 vdd.n2431 52.4337
R3498 vdd.n2427 vdd.n1221 52.4337
R3499 vdd.n2425 vdd.n2424 52.4337
R3500 vdd.n2420 vdd.n1228 52.4337
R3501 vdd.n2418 vdd.n2417 52.4337
R3502 vdd.n2413 vdd.n1235 52.4337
R3503 vdd.n2411 vdd.n2410 52.4337
R3504 vdd.n2406 vdd.n1242 52.4337
R3505 vdd.n2404 vdd.n2403 52.4337
R3506 vdd.n1251 vdd.n1250 52.4337
R3507 vdd.n2395 vdd.n1255 52.4337
R3508 vdd.n2393 vdd.n2392 52.4337
R3509 vdd.n2388 vdd.n1261 52.4337
R3510 vdd.n2386 vdd.n2385 52.4337
R3511 vdd.n2381 vdd.n1268 52.4337
R3512 vdd.n2379 vdd.n2378 52.4337
R3513 vdd.n2374 vdd.n1275 52.4337
R3514 vdd.n2372 vdd.n2371 52.4337
R3515 vdd.n1520 vdd.n1519 52.4337
R3516 vdd.n1524 vdd.n1523 52.4337
R3517 vdd.n2360 vdd.n1526 52.4337
R3518 vdd.n1875 vdd.n1874 52.4337
R3519 vdd.n1681 vdd.n1649 52.4337
R3520 vdd.n1685 vdd.n1650 52.4337
R3521 vdd.n1687 vdd.n1651 52.4337
R3522 vdd.n1691 vdd.n1652 52.4337
R3523 vdd.n1693 vdd.n1653 52.4337
R3524 vdd.n1697 vdd.n1654 52.4337
R3525 vdd.n1699 vdd.n1655 52.4337
R3526 vdd.n1703 vdd.n1656 52.4337
R3527 vdd.n1705 vdd.n1657 52.4337
R3528 vdd.n1711 vdd.n1658 52.4337
R3529 vdd.n1713 vdd.n1659 52.4337
R3530 vdd.n1717 vdd.n1660 52.4337
R3531 vdd.n1719 vdd.n1661 52.4337
R3532 vdd.n1723 vdd.n1662 52.4337
R3533 vdd.n1725 vdd.n1663 52.4337
R3534 vdd.n1729 vdd.n1664 52.4337
R3535 vdd.n1731 vdd.n1665 52.4337
R3536 vdd.n1735 vdd.n1666 52.4337
R3537 vdd.n1737 vdd.n1667 52.4337
R3538 vdd.n1809 vdd.n1668 52.4337
R3539 vdd.n1742 vdd.n1669 52.4337
R3540 vdd.n1746 vdd.n1670 52.4337
R3541 vdd.n1748 vdd.n1671 52.4337
R3542 vdd.n1752 vdd.n1672 52.4337
R3543 vdd.n1754 vdd.n1673 52.4337
R3544 vdd.n1758 vdd.n1674 52.4337
R3545 vdd.n1760 vdd.n1675 52.4337
R3546 vdd.n1764 vdd.n1676 52.4337
R3547 vdd.n1766 vdd.n1677 52.4337
R3548 vdd.n1770 vdd.n1678 52.4337
R3549 vdd.n1874 vdd.n1648 52.4337
R3550 vdd.n1684 vdd.n1649 52.4337
R3551 vdd.n1686 vdd.n1650 52.4337
R3552 vdd.n1690 vdd.n1651 52.4337
R3553 vdd.n1692 vdd.n1652 52.4337
R3554 vdd.n1696 vdd.n1653 52.4337
R3555 vdd.n1698 vdd.n1654 52.4337
R3556 vdd.n1702 vdd.n1655 52.4337
R3557 vdd.n1704 vdd.n1656 52.4337
R3558 vdd.n1710 vdd.n1657 52.4337
R3559 vdd.n1712 vdd.n1658 52.4337
R3560 vdd.n1716 vdd.n1659 52.4337
R3561 vdd.n1718 vdd.n1660 52.4337
R3562 vdd.n1722 vdd.n1661 52.4337
R3563 vdd.n1724 vdd.n1662 52.4337
R3564 vdd.n1728 vdd.n1663 52.4337
R3565 vdd.n1730 vdd.n1664 52.4337
R3566 vdd.n1734 vdd.n1665 52.4337
R3567 vdd.n1736 vdd.n1666 52.4337
R3568 vdd.n1740 vdd.n1667 52.4337
R3569 vdd.n1741 vdd.n1668 52.4337
R3570 vdd.n1745 vdd.n1669 52.4337
R3571 vdd.n1747 vdd.n1670 52.4337
R3572 vdd.n1751 vdd.n1671 52.4337
R3573 vdd.n1753 vdd.n1672 52.4337
R3574 vdd.n1757 vdd.n1673 52.4337
R3575 vdd.n1759 vdd.n1674 52.4337
R3576 vdd.n1763 vdd.n1675 52.4337
R3577 vdd.n1765 vdd.n1676 52.4337
R3578 vdd.n1769 vdd.n1677 52.4337
R3579 vdd.n1771 vdd.n1678 52.4337
R3580 vdd.n1526 vdd.n1525 52.4337
R3581 vdd.n1523 vdd.n1522 52.4337
R3582 vdd.n1519 vdd.n1276 52.4337
R3583 vdd.n2373 vdd.n2372 52.4337
R3584 vdd.n1275 vdd.n1269 52.4337
R3585 vdd.n2380 vdd.n2379 52.4337
R3586 vdd.n1268 vdd.n1262 52.4337
R3587 vdd.n2387 vdd.n2386 52.4337
R3588 vdd.n1261 vdd.n1256 52.4337
R3589 vdd.n2394 vdd.n2393 52.4337
R3590 vdd.n1255 vdd.n1254 52.4337
R3591 vdd.n1250 vdd.n1243 52.4337
R3592 vdd.n2405 vdd.n2404 52.4337
R3593 vdd.n1242 vdd.n1236 52.4337
R3594 vdd.n2412 vdd.n2411 52.4337
R3595 vdd.n1235 vdd.n1229 52.4337
R3596 vdd.n2419 vdd.n2418 52.4337
R3597 vdd.n1228 vdd.n1222 52.4337
R3598 vdd.n2426 vdd.n2425 52.4337
R3599 vdd.n1221 vdd.n1216 52.4337
R3600 vdd.n2433 vdd.n2432 52.4337
R3601 vdd.n1215 vdd.n1214 52.4337
R3602 vdd.n1210 vdd.n1203 52.4337
R3603 vdd.n2444 vdd.n2443 52.4337
R3604 vdd.n1202 vdd.n1196 52.4337
R3605 vdd.n2451 vdd.n2450 52.4337
R3606 vdd.n1195 vdd.n1189 52.4337
R3607 vdd.n2458 vdd.n2457 52.4337
R3608 vdd.n1188 vdd.n1185 52.4337
R3609 vdd.n2465 vdd.n2464 52.4337
R3610 vdd.n2470 vdd.n2469 52.4337
R3611 vdd.n1530 vdd.n1184 52.4337
R3612 vdd.n3494 vdd.n725 52.4337
R3613 vdd.n733 vdd.n693 52.4337
R3614 vdd.n3484 vdd.n694 52.4337
R3615 vdd.n3480 vdd.n695 52.4337
R3616 vdd.n3476 vdd.n696 52.4337
R3617 vdd.n3472 vdd.n697 52.4337
R3618 vdd.n3468 vdd.n698 52.4337
R3619 vdd.n3464 vdd.n699 52.4337
R3620 vdd.n3460 vdd.n700 52.4337
R3621 vdd.n3450 vdd.n701 52.4337
R3622 vdd.n3448 vdd.n702 52.4337
R3623 vdd.n3444 vdd.n703 52.4337
R3624 vdd.n3440 vdd.n704 52.4337
R3625 vdd.n3436 vdd.n705 52.4337
R3626 vdd.n3432 vdd.n706 52.4337
R3627 vdd.n3428 vdd.n707 52.4337
R3628 vdd.n3424 vdd.n708 52.4337
R3629 vdd.n3420 vdd.n709 52.4337
R3630 vdd.n3416 vdd.n710 52.4337
R3631 vdd.n3412 vdd.n711 52.4337
R3632 vdd.n3404 vdd.n712 52.4337
R3633 vdd.n3402 vdd.n713 52.4337
R3634 vdd.n3398 vdd.n714 52.4337
R3635 vdd.n3394 vdd.n715 52.4337
R3636 vdd.n3390 vdd.n716 52.4337
R3637 vdd.n3386 vdd.n717 52.4337
R3638 vdd.n3382 vdd.n718 52.4337
R3639 vdd.n3378 vdd.n719 52.4337
R3640 vdd.n3374 vdd.n720 52.4337
R3641 vdd.n3370 vdd.n721 52.4337
R3642 vdd.n722 vdd.n691 52.4337
R3643 vdd.n3625 vdd.n425 52.4337
R3644 vdd.n614 vdd.n424 52.4337
R3645 vdd.n608 vdd.n423 52.4337
R3646 vdd.n604 vdd.n422 52.4337
R3647 vdd.n598 vdd.n421 52.4337
R3648 vdd.n594 vdd.n420 52.4337
R3649 vdd.n588 vdd.n419 52.4337
R3650 vdd.n584 vdd.n418 52.4337
R3651 vdd.n578 vdd.n417 52.4337
R3652 vdd.n574 vdd.n416 52.4337
R3653 vdd.n568 vdd.n415 52.4337
R3654 vdd.n564 vdd.n414 52.4337
R3655 vdd.n558 vdd.n413 52.4337
R3656 vdd.n554 vdd.n412 52.4337
R3657 vdd.n548 vdd.n411 52.4337
R3658 vdd.n544 vdd.n410 52.4337
R3659 vdd.n538 vdd.n409 52.4337
R3660 vdd.n534 vdd.n408 52.4337
R3661 vdd.n528 vdd.n407 52.4337
R3662 vdd.n524 vdd.n406 52.4337
R3663 vdd.n518 vdd.n405 52.4337
R3664 vdd.n514 vdd.n404 52.4337
R3665 vdd.n508 vdd.n403 52.4337
R3666 vdd.n504 vdd.n402 52.4337
R3667 vdd.n498 vdd.n401 52.4337
R3668 vdd.n494 vdd.n400 52.4337
R3669 vdd.n488 vdd.n399 52.4337
R3670 vdd.n484 vdd.n398 52.4337
R3671 vdd.n478 vdd.n397 52.4337
R3672 vdd.n474 vdd.n396 52.4337
R3673 vdd.n468 vdd.n395 52.4337
R3674 vdd.n394 vdd.n392 52.4337
R3675 vdd.t238 vdd.t251 51.4683
R3676 vdd.n274 vdd.n272 42.0461
R3677 vdd.n172 vdd.n170 42.0461
R3678 vdd.n71 vdd.n69 42.0461
R3679 vdd.n2207 vdd.n2205 42.0461
R3680 vdd.n2105 vdd.n2103 42.0461
R3681 vdd.n2004 vdd.n2002 42.0461
R3682 vdd.n332 vdd.n331 41.6884
R3683 vdd.n230 vdd.n229 41.6884
R3684 vdd.n129 vdd.n128 41.6884
R3685 vdd.n2265 vdd.n2264 41.6884
R3686 vdd.n2163 vdd.n2162 41.6884
R3687 vdd.n2062 vdd.n2061 41.6884
R3688 vdd.n1774 vdd.n1773 41.1157
R3689 vdd.n1812 vdd.n1811 41.1157
R3690 vdd.n1708 vdd.n1707 41.1157
R3691 vdd.n428 vdd.n427 41.1157
R3692 vdd.n566 vdd.n441 41.1157
R3693 vdd.n454 vdd.n453 41.1157
R3694 vdd.n3325 vdd.n3324 39.2114
R3695 vdd.n3322 vdd.n3321 39.2114
R3696 vdd.n3317 vdd.n815 39.2114
R3697 vdd.n3315 vdd.n3314 39.2114
R3698 vdd.n3310 vdd.n818 39.2114
R3699 vdd.n3308 vdd.n3307 39.2114
R3700 vdd.n3303 vdd.n821 39.2114
R3701 vdd.n3301 vdd.n3300 39.2114
R3702 vdd.n3297 vdd.n3296 39.2114
R3703 vdd.n3292 vdd.n824 39.2114
R3704 vdd.n3290 vdd.n3289 39.2114
R3705 vdd.n3285 vdd.n827 39.2114
R3706 vdd.n3283 vdd.n3282 39.2114
R3707 vdd.n3278 vdd.n830 39.2114
R3708 vdd.n3276 vdd.n3275 39.2114
R3709 vdd.n3270 vdd.n835 39.2114
R3710 vdd.n3268 vdd.n3267 39.2114
R3711 vdd.n3090 vdd.n3089 39.2114
R3712 vdd.n2819 vdd.n2785 39.2114
R3713 vdd.n3082 vdd.n2786 39.2114
R3714 vdd.n3078 vdd.n2787 39.2114
R3715 vdd.n3074 vdd.n2788 39.2114
R3716 vdd.n3070 vdd.n2789 39.2114
R3717 vdd.n3066 vdd.n2790 39.2114
R3718 vdd.n3062 vdd.n2791 39.2114
R3719 vdd.n3058 vdd.n2792 39.2114
R3720 vdd.n3054 vdd.n2793 39.2114
R3721 vdd.n3050 vdd.n2794 39.2114
R3722 vdd.n3046 vdd.n2795 39.2114
R3723 vdd.n3042 vdd.n2796 39.2114
R3724 vdd.n3038 vdd.n2797 39.2114
R3725 vdd.n3034 vdd.n2798 39.2114
R3726 vdd.n3030 vdd.n2799 39.2114
R3727 vdd.n3025 vdd.n2800 39.2114
R3728 vdd.n2779 vdd.n997 39.2114
R3729 vdd.n2775 vdd.n996 39.2114
R3730 vdd.n2771 vdd.n995 39.2114
R3731 vdd.n2767 vdd.n994 39.2114
R3732 vdd.n2763 vdd.n993 39.2114
R3733 vdd.n2759 vdd.n992 39.2114
R3734 vdd.n2755 vdd.n991 39.2114
R3735 vdd.n2751 vdd.n990 39.2114
R3736 vdd.n2747 vdd.n989 39.2114
R3737 vdd.n2743 vdd.n988 39.2114
R3738 vdd.n2739 vdd.n987 39.2114
R3739 vdd.n2735 vdd.n986 39.2114
R3740 vdd.n2731 vdd.n985 39.2114
R3741 vdd.n2727 vdd.n984 39.2114
R3742 vdd.n2723 vdd.n983 39.2114
R3743 vdd.n2718 vdd.n982 39.2114
R3744 vdd.n2714 vdd.n981 39.2114
R3745 vdd.n2508 vdd.n2507 39.2114
R3746 vdd.n1176 vdd.n1142 39.2114
R3747 vdd.n2500 vdd.n1143 39.2114
R3748 vdd.n2496 vdd.n1144 39.2114
R3749 vdd.n2492 vdd.n1145 39.2114
R3750 vdd.n2488 vdd.n1146 39.2114
R3751 vdd.n2484 vdd.n1147 39.2114
R3752 vdd.n2480 vdd.n1148 39.2114
R3753 vdd.n2476 vdd.n1149 39.2114
R3754 vdd.n1322 vdd.n1150 39.2114
R3755 vdd.n1326 vdd.n1151 39.2114
R3756 vdd.n1330 vdd.n1152 39.2114
R3757 vdd.n1334 vdd.n1153 39.2114
R3758 vdd.n1338 vdd.n1154 39.2114
R3759 vdd.n1342 vdd.n1155 39.2114
R3760 vdd.n1346 vdd.n1156 39.2114
R3761 vdd.n1351 vdd.n1157 39.2114
R3762 vdd.n3244 vdd.n3243 39.2114
R3763 vdd.n3239 vdd.n3211 39.2114
R3764 vdd.n3237 vdd.n3236 39.2114
R3765 vdd.n3232 vdd.n3214 39.2114
R3766 vdd.n3230 vdd.n3229 39.2114
R3767 vdd.n3225 vdd.n3217 39.2114
R3768 vdd.n3223 vdd.n3222 39.2114
R3769 vdd.n3218 vdd.n787 39.2114
R3770 vdd.n3362 vdd.n3361 39.2114
R3771 vdd.n3359 vdd.n3358 39.2114
R3772 vdd.n3354 vdd.n791 39.2114
R3773 vdd.n3352 vdd.n3351 39.2114
R3774 vdd.n3347 vdd.n794 39.2114
R3775 vdd.n3345 vdd.n3344 39.2114
R3776 vdd.n3340 vdd.n797 39.2114
R3777 vdd.n3338 vdd.n3337 39.2114
R3778 vdd.n3333 vdd.n803 39.2114
R3779 vdd.n2826 vdd.n2801 39.2114
R3780 vdd.n2830 vdd.n2802 39.2114
R3781 vdd.n2834 vdd.n2803 39.2114
R3782 vdd.n2838 vdd.n2804 39.2114
R3783 vdd.n2842 vdd.n2805 39.2114
R3784 vdd.n2846 vdd.n2806 39.2114
R3785 vdd.n2850 vdd.n2807 39.2114
R3786 vdd.n2854 vdd.n2808 39.2114
R3787 vdd.n2858 vdd.n2809 39.2114
R3788 vdd.n2862 vdd.n2810 39.2114
R3789 vdd.n2866 vdd.n2811 39.2114
R3790 vdd.n2870 vdd.n2812 39.2114
R3791 vdd.n2874 vdd.n2813 39.2114
R3792 vdd.n2878 vdd.n2814 39.2114
R3793 vdd.n2882 vdd.n2815 39.2114
R3794 vdd.n2886 vdd.n2816 39.2114
R3795 vdd.n2890 vdd.n2817 39.2114
R3796 vdd.n2829 vdd.n2801 39.2114
R3797 vdd.n2833 vdd.n2802 39.2114
R3798 vdd.n2837 vdd.n2803 39.2114
R3799 vdd.n2841 vdd.n2804 39.2114
R3800 vdd.n2845 vdd.n2805 39.2114
R3801 vdd.n2849 vdd.n2806 39.2114
R3802 vdd.n2853 vdd.n2807 39.2114
R3803 vdd.n2857 vdd.n2808 39.2114
R3804 vdd.n2861 vdd.n2809 39.2114
R3805 vdd.n2865 vdd.n2810 39.2114
R3806 vdd.n2869 vdd.n2811 39.2114
R3807 vdd.n2873 vdd.n2812 39.2114
R3808 vdd.n2877 vdd.n2813 39.2114
R3809 vdd.n2881 vdd.n2814 39.2114
R3810 vdd.n2885 vdd.n2815 39.2114
R3811 vdd.n2889 vdd.n2816 39.2114
R3812 vdd.n2892 vdd.n2817 39.2114
R3813 vdd.n803 vdd.n798 39.2114
R3814 vdd.n3339 vdd.n3338 39.2114
R3815 vdd.n797 vdd.n795 39.2114
R3816 vdd.n3346 vdd.n3345 39.2114
R3817 vdd.n794 vdd.n792 39.2114
R3818 vdd.n3353 vdd.n3352 39.2114
R3819 vdd.n791 vdd.n789 39.2114
R3820 vdd.n3360 vdd.n3359 39.2114
R3821 vdd.n3363 vdd.n3362 39.2114
R3822 vdd.n3219 vdd.n3218 39.2114
R3823 vdd.n3224 vdd.n3223 39.2114
R3824 vdd.n3217 vdd.n3215 39.2114
R3825 vdd.n3231 vdd.n3230 39.2114
R3826 vdd.n3214 vdd.n3212 39.2114
R3827 vdd.n3238 vdd.n3237 39.2114
R3828 vdd.n3211 vdd.n3209 39.2114
R3829 vdd.n3245 vdd.n3244 39.2114
R3830 vdd.n2507 vdd.n1140 39.2114
R3831 vdd.n2501 vdd.n1142 39.2114
R3832 vdd.n2497 vdd.n1143 39.2114
R3833 vdd.n2493 vdd.n1144 39.2114
R3834 vdd.n2489 vdd.n1145 39.2114
R3835 vdd.n2485 vdd.n1146 39.2114
R3836 vdd.n2481 vdd.n1147 39.2114
R3837 vdd.n2477 vdd.n1148 39.2114
R3838 vdd.n1321 vdd.n1149 39.2114
R3839 vdd.n1325 vdd.n1150 39.2114
R3840 vdd.n1329 vdd.n1151 39.2114
R3841 vdd.n1333 vdd.n1152 39.2114
R3842 vdd.n1337 vdd.n1153 39.2114
R3843 vdd.n1341 vdd.n1154 39.2114
R3844 vdd.n1345 vdd.n1155 39.2114
R3845 vdd.n1350 vdd.n1156 39.2114
R3846 vdd.n1354 vdd.n1157 39.2114
R3847 vdd.n2717 vdd.n981 39.2114
R3848 vdd.n2722 vdd.n982 39.2114
R3849 vdd.n2726 vdd.n983 39.2114
R3850 vdd.n2730 vdd.n984 39.2114
R3851 vdd.n2734 vdd.n985 39.2114
R3852 vdd.n2738 vdd.n986 39.2114
R3853 vdd.n2742 vdd.n987 39.2114
R3854 vdd.n2746 vdd.n988 39.2114
R3855 vdd.n2750 vdd.n989 39.2114
R3856 vdd.n2754 vdd.n990 39.2114
R3857 vdd.n2758 vdd.n991 39.2114
R3858 vdd.n2762 vdd.n992 39.2114
R3859 vdd.n2766 vdd.n993 39.2114
R3860 vdd.n2770 vdd.n994 39.2114
R3861 vdd.n2774 vdd.n995 39.2114
R3862 vdd.n2778 vdd.n996 39.2114
R3863 vdd.n999 vdd.n997 39.2114
R3864 vdd.n3089 vdd.n962 39.2114
R3865 vdd.n3083 vdd.n2785 39.2114
R3866 vdd.n3079 vdd.n2786 39.2114
R3867 vdd.n3075 vdd.n2787 39.2114
R3868 vdd.n3071 vdd.n2788 39.2114
R3869 vdd.n3067 vdd.n2789 39.2114
R3870 vdd.n3063 vdd.n2790 39.2114
R3871 vdd.n3059 vdd.n2791 39.2114
R3872 vdd.n3055 vdd.n2792 39.2114
R3873 vdd.n3051 vdd.n2793 39.2114
R3874 vdd.n3047 vdd.n2794 39.2114
R3875 vdd.n3043 vdd.n2795 39.2114
R3876 vdd.n3039 vdd.n2796 39.2114
R3877 vdd.n3035 vdd.n2797 39.2114
R3878 vdd.n3031 vdd.n2798 39.2114
R3879 vdd.n3026 vdd.n2799 39.2114
R3880 vdd.n3022 vdd.n2800 39.2114
R3881 vdd.n3269 vdd.n3268 39.2114
R3882 vdd.n835 vdd.n831 39.2114
R3883 vdd.n3277 vdd.n3276 39.2114
R3884 vdd.n830 vdd.n828 39.2114
R3885 vdd.n3284 vdd.n3283 39.2114
R3886 vdd.n827 vdd.n825 39.2114
R3887 vdd.n3291 vdd.n3290 39.2114
R3888 vdd.n824 vdd.n822 39.2114
R3889 vdd.n3298 vdd.n3297 39.2114
R3890 vdd.n3302 vdd.n3301 39.2114
R3891 vdd.n821 vdd.n819 39.2114
R3892 vdd.n3309 vdd.n3308 39.2114
R3893 vdd.n818 vdd.n816 39.2114
R3894 vdd.n3316 vdd.n3315 39.2114
R3895 vdd.n815 vdd.n813 39.2114
R3896 vdd.n3323 vdd.n3322 39.2114
R3897 vdd.n3326 vdd.n3325 39.2114
R3898 vdd.n1008 vdd.n963 39.2114
R3899 vdd.n2706 vdd.n964 39.2114
R3900 vdd.n2702 vdd.n965 39.2114
R3901 vdd.n2698 vdd.n966 39.2114
R3902 vdd.n2694 vdd.n967 39.2114
R3903 vdd.n2690 vdd.n968 39.2114
R3904 vdd.n2686 vdd.n969 39.2114
R3905 vdd.n2682 vdd.n970 39.2114
R3906 vdd.n2678 vdd.n971 39.2114
R3907 vdd.n2674 vdd.n972 39.2114
R3908 vdd.n2670 vdd.n973 39.2114
R3909 vdd.n2666 vdd.n974 39.2114
R3910 vdd.n2662 vdd.n975 39.2114
R3911 vdd.n2658 vdd.n976 39.2114
R3912 vdd.n2654 vdd.n977 39.2114
R3913 vdd.n2650 vdd.n978 39.2114
R3914 vdd.n2646 vdd.n979 39.2114
R3915 vdd.n1280 vdd.n1158 39.2114
R3916 vdd.n1284 vdd.n1159 39.2114
R3917 vdd.n1288 vdd.n1160 39.2114
R3918 vdd.n1292 vdd.n1161 39.2114
R3919 vdd.n1296 vdd.n1162 39.2114
R3920 vdd.n1300 vdd.n1163 39.2114
R3921 vdd.n1304 vdd.n1164 39.2114
R3922 vdd.n1308 vdd.n1165 39.2114
R3923 vdd.n1312 vdd.n1166 39.2114
R3924 vdd.n1513 vdd.n1167 39.2114
R3925 vdd.n1510 vdd.n1168 39.2114
R3926 vdd.n1506 vdd.n1169 39.2114
R3927 vdd.n1502 vdd.n1170 39.2114
R3928 vdd.n1498 vdd.n1171 39.2114
R3929 vdd.n1494 vdd.n1172 39.2114
R3930 vdd.n1490 vdd.n1173 39.2114
R3931 vdd.n1486 vdd.n1174 39.2114
R3932 vdd.n2643 vdd.n979 39.2114
R3933 vdd.n2647 vdd.n978 39.2114
R3934 vdd.n2651 vdd.n977 39.2114
R3935 vdd.n2655 vdd.n976 39.2114
R3936 vdd.n2659 vdd.n975 39.2114
R3937 vdd.n2663 vdd.n974 39.2114
R3938 vdd.n2667 vdd.n973 39.2114
R3939 vdd.n2671 vdd.n972 39.2114
R3940 vdd.n2675 vdd.n971 39.2114
R3941 vdd.n2679 vdd.n970 39.2114
R3942 vdd.n2683 vdd.n969 39.2114
R3943 vdd.n2687 vdd.n968 39.2114
R3944 vdd.n2691 vdd.n967 39.2114
R3945 vdd.n2695 vdd.n966 39.2114
R3946 vdd.n2699 vdd.n965 39.2114
R3947 vdd.n2703 vdd.n964 39.2114
R3948 vdd.n2707 vdd.n963 39.2114
R3949 vdd.n1283 vdd.n1158 39.2114
R3950 vdd.n1287 vdd.n1159 39.2114
R3951 vdd.n1291 vdd.n1160 39.2114
R3952 vdd.n1295 vdd.n1161 39.2114
R3953 vdd.n1299 vdd.n1162 39.2114
R3954 vdd.n1303 vdd.n1163 39.2114
R3955 vdd.n1307 vdd.n1164 39.2114
R3956 vdd.n1311 vdd.n1165 39.2114
R3957 vdd.n1314 vdd.n1166 39.2114
R3958 vdd.n1511 vdd.n1167 39.2114
R3959 vdd.n1507 vdd.n1168 39.2114
R3960 vdd.n1503 vdd.n1169 39.2114
R3961 vdd.n1499 vdd.n1170 39.2114
R3962 vdd.n1495 vdd.n1171 39.2114
R3963 vdd.n1491 vdd.n1172 39.2114
R3964 vdd.n1487 vdd.n1173 39.2114
R3965 vdd.n1483 vdd.n1174 39.2114
R3966 vdd.n2364 vdd.n2363 37.2369
R3967 vdd.n2400 vdd.n1249 37.2369
R3968 vdd.n2439 vdd.n1209 37.2369
R3969 vdd.n3410 vdd.n769 37.2369
R3970 vdd.n3458 vdd.n3457 37.2369
R3971 vdd.n690 vdd.n689 37.2369
R3972 vdd.n1317 vdd.n1316 30.449
R3973 vdd.n1012 vdd.n1011 30.449
R3974 vdd.n1348 vdd.n1320 30.449
R3975 vdd.n2720 vdd.n1002 30.449
R3976 vdd.n2825 vdd.n2824 30.449
R3977 vdd.n3272 vdd.n833 30.449
R3978 vdd.n3028 vdd.n2821 30.449
R3979 vdd.n801 vdd.n800 30.449
R3980 vdd.n2510 vdd.n2509 29.8151
R3981 vdd.n2782 vdd.n1000 29.8151
R3982 vdd.n2715 vdd.n1003 29.8151
R3983 vdd.n1356 vdd.n1353 29.8151
R3984 vdd.n3023 vdd.n3020 29.8151
R3985 vdd.n3266 vdd.n3265 29.8151
R3986 vdd.n3092 vdd.n3091 29.8151
R3987 vdd.n3329 vdd.n3328 29.8151
R3988 vdd.n3248 vdd.n3247 29.8151
R3989 vdd.n3334 vdd.n802 29.8151
R3990 vdd.n2896 vdd.n2894 29.8151
R3991 vdd.n2827 vdd.n955 29.8151
R3992 vdd.n1281 vdd.n1132 29.8151
R3993 vdd.n2710 vdd.n2709 29.8151
R3994 vdd.n2642 vdd.n2641 29.8151
R3995 vdd.n1482 vdd.n1481 29.8151
R3996 vdd.n1873 vdd.n1680 22.2201
R3997 vdd.n2358 vdd.n1141 22.2201
R3998 vdd.n3495 vdd.n723 22.2201
R3999 vdd.n3627 vdd.n3626 22.2201
R4000 vdd.n1884 vdd.n1642 19.3944
R4001 vdd.n1884 vdd.n1640 19.3944
R4002 vdd.n1888 vdd.n1640 19.3944
R4003 vdd.n1888 vdd.n1630 19.3944
R4004 vdd.n1901 vdd.n1630 19.3944
R4005 vdd.n1901 vdd.n1628 19.3944
R4006 vdd.n1905 vdd.n1628 19.3944
R4007 vdd.n1905 vdd.n1620 19.3944
R4008 vdd.n1918 vdd.n1620 19.3944
R4009 vdd.n1918 vdd.n1618 19.3944
R4010 vdd.n1922 vdd.n1618 19.3944
R4011 vdd.n1922 vdd.n1607 19.3944
R4012 vdd.n1934 vdd.n1607 19.3944
R4013 vdd.n1934 vdd.n1605 19.3944
R4014 vdd.n1938 vdd.n1605 19.3944
R4015 vdd.n1938 vdd.n1596 19.3944
R4016 vdd.n1951 vdd.n1596 19.3944
R4017 vdd.n1951 vdd.n1594 19.3944
R4018 vdd.n1955 vdd.n1594 19.3944
R4019 vdd.n1955 vdd.n1585 19.3944
R4020 vdd.n2274 vdd.n1585 19.3944
R4021 vdd.n2274 vdd.n1583 19.3944
R4022 vdd.n2278 vdd.n1583 19.3944
R4023 vdd.n2278 vdd.n1573 19.3944
R4024 vdd.n2291 vdd.n1573 19.3944
R4025 vdd.n2291 vdd.n1571 19.3944
R4026 vdd.n2295 vdd.n1571 19.3944
R4027 vdd.n2295 vdd.n1563 19.3944
R4028 vdd.n2308 vdd.n1563 19.3944
R4029 vdd.n2308 vdd.n1561 19.3944
R4030 vdd.n2312 vdd.n1561 19.3944
R4031 vdd.n2312 vdd.n1550 19.3944
R4032 vdd.n2324 vdd.n1550 19.3944
R4033 vdd.n2324 vdd.n1548 19.3944
R4034 vdd.n2328 vdd.n1548 19.3944
R4035 vdd.n2328 vdd.n1540 19.3944
R4036 vdd.n2341 vdd.n1540 19.3944
R4037 vdd.n2341 vdd.n1537 19.3944
R4038 vdd.n2347 vdd.n1537 19.3944
R4039 vdd.n2347 vdd.n1538 19.3944
R4040 vdd.n1538 vdd.n1528 19.3944
R4041 vdd.n1808 vdd.n1743 19.3944
R4042 vdd.n1804 vdd.n1743 19.3944
R4043 vdd.n1804 vdd.n1803 19.3944
R4044 vdd.n1803 vdd.n1802 19.3944
R4045 vdd.n1802 vdd.n1749 19.3944
R4046 vdd.n1798 vdd.n1749 19.3944
R4047 vdd.n1798 vdd.n1797 19.3944
R4048 vdd.n1797 vdd.n1796 19.3944
R4049 vdd.n1796 vdd.n1755 19.3944
R4050 vdd.n1792 vdd.n1755 19.3944
R4051 vdd.n1792 vdd.n1791 19.3944
R4052 vdd.n1791 vdd.n1790 19.3944
R4053 vdd.n1790 vdd.n1761 19.3944
R4054 vdd.n1786 vdd.n1761 19.3944
R4055 vdd.n1786 vdd.n1785 19.3944
R4056 vdd.n1785 vdd.n1784 19.3944
R4057 vdd.n1784 vdd.n1767 19.3944
R4058 vdd.n1780 vdd.n1767 19.3944
R4059 vdd.n1780 vdd.n1779 19.3944
R4060 vdd.n1779 vdd.n1778 19.3944
R4061 vdd.n1843 vdd.n1842 19.3944
R4062 vdd.n1842 vdd.n1841 19.3944
R4063 vdd.n1841 vdd.n1714 19.3944
R4064 vdd.n1837 vdd.n1714 19.3944
R4065 vdd.n1837 vdd.n1836 19.3944
R4066 vdd.n1836 vdd.n1835 19.3944
R4067 vdd.n1835 vdd.n1720 19.3944
R4068 vdd.n1831 vdd.n1720 19.3944
R4069 vdd.n1831 vdd.n1830 19.3944
R4070 vdd.n1830 vdd.n1829 19.3944
R4071 vdd.n1829 vdd.n1726 19.3944
R4072 vdd.n1825 vdd.n1726 19.3944
R4073 vdd.n1825 vdd.n1824 19.3944
R4074 vdd.n1824 vdd.n1823 19.3944
R4075 vdd.n1823 vdd.n1732 19.3944
R4076 vdd.n1819 vdd.n1732 19.3944
R4077 vdd.n1819 vdd.n1818 19.3944
R4078 vdd.n1818 vdd.n1817 19.3944
R4079 vdd.n1817 vdd.n1738 19.3944
R4080 vdd.n1813 vdd.n1738 19.3944
R4081 vdd.n1876 vdd.n1647 19.3944
R4082 vdd.n1871 vdd.n1647 19.3944
R4083 vdd.n1871 vdd.n1682 19.3944
R4084 vdd.n1867 vdd.n1682 19.3944
R4085 vdd.n1867 vdd.n1866 19.3944
R4086 vdd.n1866 vdd.n1865 19.3944
R4087 vdd.n1865 vdd.n1688 19.3944
R4088 vdd.n1861 vdd.n1688 19.3944
R4089 vdd.n1861 vdd.n1860 19.3944
R4090 vdd.n1860 vdd.n1859 19.3944
R4091 vdd.n1859 vdd.n1694 19.3944
R4092 vdd.n1855 vdd.n1694 19.3944
R4093 vdd.n1855 vdd.n1854 19.3944
R4094 vdd.n1854 vdd.n1853 19.3944
R4095 vdd.n1853 vdd.n1700 19.3944
R4096 vdd.n1849 vdd.n1700 19.3944
R4097 vdd.n1849 vdd.n1848 19.3944
R4098 vdd.n1848 vdd.n1847 19.3944
R4099 vdd.n2396 vdd.n1247 19.3944
R4100 vdd.n2396 vdd.n1253 19.3944
R4101 vdd.n2391 vdd.n1253 19.3944
R4102 vdd.n2391 vdd.n2390 19.3944
R4103 vdd.n2390 vdd.n2389 19.3944
R4104 vdd.n2389 vdd.n1260 19.3944
R4105 vdd.n2384 vdd.n1260 19.3944
R4106 vdd.n2384 vdd.n2383 19.3944
R4107 vdd.n2383 vdd.n2382 19.3944
R4108 vdd.n2382 vdd.n1267 19.3944
R4109 vdd.n2377 vdd.n1267 19.3944
R4110 vdd.n2377 vdd.n2376 19.3944
R4111 vdd.n2376 vdd.n2375 19.3944
R4112 vdd.n2375 vdd.n1274 19.3944
R4113 vdd.n2370 vdd.n1274 19.3944
R4114 vdd.n2370 vdd.n2369 19.3944
R4115 vdd.n1521 vdd.n1279 19.3944
R4116 vdd.n2365 vdd.n1518 19.3944
R4117 vdd.n2435 vdd.n1207 19.3944
R4118 vdd.n2435 vdd.n1213 19.3944
R4119 vdd.n2430 vdd.n1213 19.3944
R4120 vdd.n2430 vdd.n2429 19.3944
R4121 vdd.n2429 vdd.n2428 19.3944
R4122 vdd.n2428 vdd.n1220 19.3944
R4123 vdd.n2423 vdd.n1220 19.3944
R4124 vdd.n2423 vdd.n2422 19.3944
R4125 vdd.n2422 vdd.n2421 19.3944
R4126 vdd.n2421 vdd.n1227 19.3944
R4127 vdd.n2416 vdd.n1227 19.3944
R4128 vdd.n2416 vdd.n2415 19.3944
R4129 vdd.n2415 vdd.n2414 19.3944
R4130 vdd.n2414 vdd.n1234 19.3944
R4131 vdd.n2409 vdd.n1234 19.3944
R4132 vdd.n2409 vdd.n2408 19.3944
R4133 vdd.n2408 vdd.n2407 19.3944
R4134 vdd.n2407 vdd.n1241 19.3944
R4135 vdd.n2402 vdd.n1241 19.3944
R4136 vdd.n2402 vdd.n2401 19.3944
R4137 vdd.n2472 vdd.n1182 19.3944
R4138 vdd.n2472 vdd.n1183 19.3944
R4139 vdd.n2467 vdd.n2466 19.3944
R4140 vdd.n2462 vdd.n2461 19.3944
R4141 vdd.n2461 vdd.n2460 19.3944
R4142 vdd.n2460 vdd.n1187 19.3944
R4143 vdd.n2455 vdd.n1187 19.3944
R4144 vdd.n2455 vdd.n2454 19.3944
R4145 vdd.n2454 vdd.n2453 19.3944
R4146 vdd.n2453 vdd.n1194 19.3944
R4147 vdd.n2448 vdd.n1194 19.3944
R4148 vdd.n2448 vdd.n2447 19.3944
R4149 vdd.n2447 vdd.n2446 19.3944
R4150 vdd.n2446 vdd.n1201 19.3944
R4151 vdd.n2441 vdd.n1201 19.3944
R4152 vdd.n2441 vdd.n2440 19.3944
R4153 vdd.n1880 vdd.n1645 19.3944
R4154 vdd.n1880 vdd.n1636 19.3944
R4155 vdd.n1893 vdd.n1636 19.3944
R4156 vdd.n1893 vdd.n1634 19.3944
R4157 vdd.n1897 vdd.n1634 19.3944
R4158 vdd.n1897 vdd.n1625 19.3944
R4159 vdd.n1910 vdd.n1625 19.3944
R4160 vdd.n1910 vdd.n1623 19.3944
R4161 vdd.n1914 vdd.n1623 19.3944
R4162 vdd.n1914 vdd.n1614 19.3944
R4163 vdd.n1926 vdd.n1614 19.3944
R4164 vdd.n1926 vdd.n1612 19.3944
R4165 vdd.n1930 vdd.n1612 19.3944
R4166 vdd.n1930 vdd.n1602 19.3944
R4167 vdd.n1943 vdd.n1602 19.3944
R4168 vdd.n1943 vdd.n1600 19.3944
R4169 vdd.n1947 vdd.n1600 19.3944
R4170 vdd.n1947 vdd.n1591 19.3944
R4171 vdd.n1959 vdd.n1591 19.3944
R4172 vdd.n1959 vdd.n1589 19.3944
R4173 vdd.n2270 vdd.n1589 19.3944
R4174 vdd.n2270 vdd.n1579 19.3944
R4175 vdd.n2283 vdd.n1579 19.3944
R4176 vdd.n2283 vdd.n1577 19.3944
R4177 vdd.n2287 vdd.n1577 19.3944
R4178 vdd.n2287 vdd.n1568 19.3944
R4179 vdd.n2300 vdd.n1568 19.3944
R4180 vdd.n2300 vdd.n1566 19.3944
R4181 vdd.n2304 vdd.n1566 19.3944
R4182 vdd.n2304 vdd.n1557 19.3944
R4183 vdd.n2316 vdd.n1557 19.3944
R4184 vdd.n2316 vdd.n1555 19.3944
R4185 vdd.n2320 vdd.n1555 19.3944
R4186 vdd.n2320 vdd.n1545 19.3944
R4187 vdd.n2333 vdd.n1545 19.3944
R4188 vdd.n2333 vdd.n1543 19.3944
R4189 vdd.n2337 vdd.n1543 19.3944
R4190 vdd.n2337 vdd.n1533 19.3944
R4191 vdd.n2352 vdd.n1533 19.3944
R4192 vdd.n2352 vdd.n1531 19.3944
R4193 vdd.n2356 vdd.n1531 19.3944
R4194 vdd.n3501 vdd.n686 19.3944
R4195 vdd.n3501 vdd.n676 19.3944
R4196 vdd.n3513 vdd.n676 19.3944
R4197 vdd.n3513 vdd.n674 19.3944
R4198 vdd.n3517 vdd.n674 19.3944
R4199 vdd.n3517 vdd.n666 19.3944
R4200 vdd.n3530 vdd.n666 19.3944
R4201 vdd.n3530 vdd.n664 19.3944
R4202 vdd.n3534 vdd.n664 19.3944
R4203 vdd.n3534 vdd.n653 19.3944
R4204 vdd.n3546 vdd.n653 19.3944
R4205 vdd.n3546 vdd.n651 19.3944
R4206 vdd.n3550 vdd.n651 19.3944
R4207 vdd.n3550 vdd.n642 19.3944
R4208 vdd.n3563 vdd.n642 19.3944
R4209 vdd.n3563 vdd.n640 19.3944
R4210 vdd.n3570 vdd.n640 19.3944
R4211 vdd.n3570 vdd.n3569 19.3944
R4212 vdd.n3569 vdd.n631 19.3944
R4213 vdd.n3583 vdd.n631 19.3944
R4214 vdd.n3584 vdd.n3583 19.3944
R4215 vdd.n3584 vdd.n629 19.3944
R4216 vdd.n3588 vdd.n629 19.3944
R4217 vdd.n3590 vdd.n3588 19.3944
R4218 vdd.n3591 vdd.n3590 19.3944
R4219 vdd.n3591 vdd.n627 19.3944
R4220 vdd.n3595 vdd.n627 19.3944
R4221 vdd.n3597 vdd.n3595 19.3944
R4222 vdd.n3598 vdd.n3597 19.3944
R4223 vdd.n3598 vdd.n625 19.3944
R4224 vdd.n3602 vdd.n625 19.3944
R4225 vdd.n3605 vdd.n3602 19.3944
R4226 vdd.n3606 vdd.n3605 19.3944
R4227 vdd.n3606 vdd.n623 19.3944
R4228 vdd.n3610 vdd.n623 19.3944
R4229 vdd.n3612 vdd.n3610 19.3944
R4230 vdd.n3613 vdd.n3612 19.3944
R4231 vdd.n3613 vdd.n621 19.3944
R4232 vdd.n3617 vdd.n621 19.3944
R4233 vdd.n3619 vdd.n3617 19.3944
R4234 vdd.n3620 vdd.n3619 19.3944
R4235 vdd.n569 vdd.n438 19.3944
R4236 vdd.n575 vdd.n438 19.3944
R4237 vdd.n576 vdd.n575 19.3944
R4238 vdd.n579 vdd.n576 19.3944
R4239 vdd.n579 vdd.n436 19.3944
R4240 vdd.n585 vdd.n436 19.3944
R4241 vdd.n586 vdd.n585 19.3944
R4242 vdd.n589 vdd.n586 19.3944
R4243 vdd.n589 vdd.n434 19.3944
R4244 vdd.n595 vdd.n434 19.3944
R4245 vdd.n596 vdd.n595 19.3944
R4246 vdd.n599 vdd.n596 19.3944
R4247 vdd.n599 vdd.n432 19.3944
R4248 vdd.n605 vdd.n432 19.3944
R4249 vdd.n606 vdd.n605 19.3944
R4250 vdd.n609 vdd.n606 19.3944
R4251 vdd.n609 vdd.n430 19.3944
R4252 vdd.n615 vdd.n430 19.3944
R4253 vdd.n617 vdd.n615 19.3944
R4254 vdd.n618 vdd.n617 19.3944
R4255 vdd.n516 vdd.n515 19.3944
R4256 vdd.n519 vdd.n516 19.3944
R4257 vdd.n519 vdd.n450 19.3944
R4258 vdd.n525 vdd.n450 19.3944
R4259 vdd.n526 vdd.n525 19.3944
R4260 vdd.n529 vdd.n526 19.3944
R4261 vdd.n529 vdd.n448 19.3944
R4262 vdd.n535 vdd.n448 19.3944
R4263 vdd.n536 vdd.n535 19.3944
R4264 vdd.n539 vdd.n536 19.3944
R4265 vdd.n539 vdd.n446 19.3944
R4266 vdd.n545 vdd.n446 19.3944
R4267 vdd.n546 vdd.n545 19.3944
R4268 vdd.n549 vdd.n546 19.3944
R4269 vdd.n549 vdd.n444 19.3944
R4270 vdd.n555 vdd.n444 19.3944
R4271 vdd.n556 vdd.n555 19.3944
R4272 vdd.n559 vdd.n556 19.3944
R4273 vdd.n559 vdd.n442 19.3944
R4274 vdd.n565 vdd.n442 19.3944
R4275 vdd.n466 vdd.n465 19.3944
R4276 vdd.n469 vdd.n466 19.3944
R4277 vdd.n469 vdd.n462 19.3944
R4278 vdd.n475 vdd.n462 19.3944
R4279 vdd.n476 vdd.n475 19.3944
R4280 vdd.n479 vdd.n476 19.3944
R4281 vdd.n479 vdd.n460 19.3944
R4282 vdd.n485 vdd.n460 19.3944
R4283 vdd.n486 vdd.n485 19.3944
R4284 vdd.n489 vdd.n486 19.3944
R4285 vdd.n489 vdd.n458 19.3944
R4286 vdd.n495 vdd.n458 19.3944
R4287 vdd.n496 vdd.n495 19.3944
R4288 vdd.n499 vdd.n496 19.3944
R4289 vdd.n499 vdd.n456 19.3944
R4290 vdd.n505 vdd.n456 19.3944
R4291 vdd.n506 vdd.n505 19.3944
R4292 vdd.n509 vdd.n506 19.3944
R4293 vdd.n3505 vdd.n683 19.3944
R4294 vdd.n3505 vdd.n681 19.3944
R4295 vdd.n3509 vdd.n681 19.3944
R4296 vdd.n3509 vdd.n671 19.3944
R4297 vdd.n3522 vdd.n671 19.3944
R4298 vdd.n3522 vdd.n669 19.3944
R4299 vdd.n3526 vdd.n669 19.3944
R4300 vdd.n3526 vdd.n660 19.3944
R4301 vdd.n3538 vdd.n660 19.3944
R4302 vdd.n3538 vdd.n658 19.3944
R4303 vdd.n3542 vdd.n658 19.3944
R4304 vdd.n3542 vdd.n648 19.3944
R4305 vdd.n3555 vdd.n648 19.3944
R4306 vdd.n3555 vdd.n646 19.3944
R4307 vdd.n3559 vdd.n646 19.3944
R4308 vdd.n3559 vdd.n637 19.3944
R4309 vdd.n3574 vdd.n637 19.3944
R4310 vdd.n3574 vdd.n635 19.3944
R4311 vdd.n3578 vdd.n635 19.3944
R4312 vdd.n3578 vdd.n336 19.3944
R4313 vdd.n3669 vdd.n336 19.3944
R4314 vdd.n3669 vdd.n337 19.3944
R4315 vdd.n3663 vdd.n337 19.3944
R4316 vdd.n3663 vdd.n3662 19.3944
R4317 vdd.n3662 vdd.n3661 19.3944
R4318 vdd.n3661 vdd.n349 19.3944
R4319 vdd.n3655 vdd.n349 19.3944
R4320 vdd.n3655 vdd.n3654 19.3944
R4321 vdd.n3654 vdd.n3653 19.3944
R4322 vdd.n3653 vdd.n359 19.3944
R4323 vdd.n3647 vdd.n359 19.3944
R4324 vdd.n3647 vdd.n3646 19.3944
R4325 vdd.n3646 vdd.n3645 19.3944
R4326 vdd.n3645 vdd.n370 19.3944
R4327 vdd.n3639 vdd.n370 19.3944
R4328 vdd.n3639 vdd.n3638 19.3944
R4329 vdd.n3638 vdd.n3637 19.3944
R4330 vdd.n3637 vdd.n381 19.3944
R4331 vdd.n3631 vdd.n381 19.3944
R4332 vdd.n3631 vdd.n3630 19.3944
R4333 vdd.n3630 vdd.n3629 19.3944
R4334 vdd.n3452 vdd.n747 19.3944
R4335 vdd.n3452 vdd.n3449 19.3944
R4336 vdd.n3449 vdd.n3446 19.3944
R4337 vdd.n3446 vdd.n3445 19.3944
R4338 vdd.n3445 vdd.n3442 19.3944
R4339 vdd.n3442 vdd.n3441 19.3944
R4340 vdd.n3441 vdd.n3438 19.3944
R4341 vdd.n3438 vdd.n3437 19.3944
R4342 vdd.n3437 vdd.n3434 19.3944
R4343 vdd.n3434 vdd.n3433 19.3944
R4344 vdd.n3433 vdd.n3430 19.3944
R4345 vdd.n3430 vdd.n3429 19.3944
R4346 vdd.n3429 vdd.n3426 19.3944
R4347 vdd.n3426 vdd.n3425 19.3944
R4348 vdd.n3425 vdd.n3422 19.3944
R4349 vdd.n3422 vdd.n3421 19.3944
R4350 vdd.n3421 vdd.n3418 19.3944
R4351 vdd.n3418 vdd.n3417 19.3944
R4352 vdd.n3417 vdd.n3414 19.3944
R4353 vdd.n3414 vdd.n3413 19.3944
R4354 vdd.n3492 vdd.n3491 19.3944
R4355 vdd.n3491 vdd.n3490 19.3944
R4356 vdd.n732 vdd.n729 19.3944
R4357 vdd.n3486 vdd.n3485 19.3944
R4358 vdd.n3485 vdd.n3482 19.3944
R4359 vdd.n3482 vdd.n3481 19.3944
R4360 vdd.n3481 vdd.n3478 19.3944
R4361 vdd.n3478 vdd.n3477 19.3944
R4362 vdd.n3477 vdd.n3474 19.3944
R4363 vdd.n3474 vdd.n3473 19.3944
R4364 vdd.n3473 vdd.n3470 19.3944
R4365 vdd.n3470 vdd.n3469 19.3944
R4366 vdd.n3469 vdd.n3466 19.3944
R4367 vdd.n3466 vdd.n3465 19.3944
R4368 vdd.n3465 vdd.n3462 19.3944
R4369 vdd.n3462 vdd.n3461 19.3944
R4370 vdd.n3406 vdd.n767 19.3944
R4371 vdd.n3406 vdd.n3403 19.3944
R4372 vdd.n3403 vdd.n3400 19.3944
R4373 vdd.n3400 vdd.n3399 19.3944
R4374 vdd.n3399 vdd.n3396 19.3944
R4375 vdd.n3396 vdd.n3395 19.3944
R4376 vdd.n3395 vdd.n3392 19.3944
R4377 vdd.n3392 vdd.n3391 19.3944
R4378 vdd.n3391 vdd.n3388 19.3944
R4379 vdd.n3388 vdd.n3387 19.3944
R4380 vdd.n3387 vdd.n3384 19.3944
R4381 vdd.n3384 vdd.n3383 19.3944
R4382 vdd.n3383 vdd.n3380 19.3944
R4383 vdd.n3380 vdd.n3379 19.3944
R4384 vdd.n3379 vdd.n3376 19.3944
R4385 vdd.n3376 vdd.n3375 19.3944
R4386 vdd.n3372 vdd.n3371 19.3944
R4387 vdd.n3368 vdd.n3367 19.3944
R4388 vdd.n1812 vdd.n1808 19.0066
R4389 vdd.n2400 vdd.n1247 19.0066
R4390 vdd.n569 vdd.n566 19.0066
R4391 vdd.n3410 vdd.n767 19.0066
R4392 vdd.n1316 vdd.n1315 16.0975
R4393 vdd.n1011 vdd.n1010 16.0975
R4394 vdd.n1773 vdd.n1772 16.0975
R4395 vdd.n1811 vdd.n1810 16.0975
R4396 vdd.n1707 vdd.n1706 16.0975
R4397 vdd.n2363 vdd.n2362 16.0975
R4398 vdd.n1249 vdd.n1248 16.0975
R4399 vdd.n1209 vdd.n1208 16.0975
R4400 vdd.n1320 vdd.n1319 16.0975
R4401 vdd.n1002 vdd.n1001 16.0975
R4402 vdd.n2824 vdd.n2823 16.0975
R4403 vdd.n427 vdd.n426 16.0975
R4404 vdd.n441 vdd.n440 16.0975
R4405 vdd.n453 vdd.n452 16.0975
R4406 vdd.n769 vdd.n768 16.0975
R4407 vdd.n3457 vdd.n3456 16.0975
R4408 vdd.n833 vdd.n832 16.0975
R4409 vdd.n2821 vdd.n2820 16.0975
R4410 vdd.n689 vdd.n688 16.0975
R4411 vdd.n800 vdd.n799 16.0975
R4412 vdd.t251 vdd.n2784 15.4182
R4413 vdd.n3088 vdd.t238 15.4182
R4414 vdd.n28 vdd.n27 14.6072
R4415 vdd.n328 vdd.n293 13.1884
R4416 vdd.n269 vdd.n234 13.1884
R4417 vdd.n226 vdd.n191 13.1884
R4418 vdd.n167 vdd.n132 13.1884
R4419 vdd.n125 vdd.n90 13.1884
R4420 vdd.n66 vdd.n31 13.1884
R4421 vdd.n2202 vdd.n2167 13.1884
R4422 vdd.n2261 vdd.n2226 13.1884
R4423 vdd.n2100 vdd.n2065 13.1884
R4424 vdd.n2159 vdd.n2124 13.1884
R4425 vdd.n1999 vdd.n1964 13.1884
R4426 vdd.n2058 vdd.n2023 13.1884
R4427 vdd.n2506 vdd.n1134 13.1509
R4428 vdd.n3331 vdd.n692 13.1509
R4429 vdd.n1843 vdd.n1708 12.9944
R4430 vdd.n1847 vdd.n1708 12.9944
R4431 vdd.n2439 vdd.n1207 12.9944
R4432 vdd.n2440 vdd.n2439 12.9944
R4433 vdd.n515 vdd.n454 12.9944
R4434 vdd.n509 vdd.n454 12.9944
R4435 vdd.n3458 vdd.n747 12.9944
R4436 vdd.n3461 vdd.n3458 12.9944
R4437 vdd.n329 vdd.n291 12.8005
R4438 vdd.n324 vdd.n295 12.8005
R4439 vdd.n270 vdd.n232 12.8005
R4440 vdd.n265 vdd.n236 12.8005
R4441 vdd.n227 vdd.n189 12.8005
R4442 vdd.n222 vdd.n193 12.8005
R4443 vdd.n168 vdd.n130 12.8005
R4444 vdd.n163 vdd.n134 12.8005
R4445 vdd.n126 vdd.n88 12.8005
R4446 vdd.n121 vdd.n92 12.8005
R4447 vdd.n67 vdd.n29 12.8005
R4448 vdd.n62 vdd.n33 12.8005
R4449 vdd.n2203 vdd.n2165 12.8005
R4450 vdd.n2198 vdd.n2169 12.8005
R4451 vdd.n2262 vdd.n2224 12.8005
R4452 vdd.n2257 vdd.n2228 12.8005
R4453 vdd.n2101 vdd.n2063 12.8005
R4454 vdd.n2096 vdd.n2067 12.8005
R4455 vdd.n2160 vdd.n2122 12.8005
R4456 vdd.n2155 vdd.n2126 12.8005
R4457 vdd.n2000 vdd.n1962 12.8005
R4458 vdd.n1995 vdd.n1966 12.8005
R4459 vdd.n2059 vdd.n2021 12.8005
R4460 vdd.n2054 vdd.n2025 12.8005
R4461 vdd.n323 vdd.n296 12.0247
R4462 vdd.n264 vdd.n237 12.0247
R4463 vdd.n221 vdd.n194 12.0247
R4464 vdd.n162 vdd.n135 12.0247
R4465 vdd.n120 vdd.n93 12.0247
R4466 vdd.n61 vdd.n34 12.0247
R4467 vdd.n2197 vdd.n2170 12.0247
R4468 vdd.n2256 vdd.n2229 12.0247
R4469 vdd.n2095 vdd.n2068 12.0247
R4470 vdd.n2154 vdd.n2127 12.0247
R4471 vdd.n1994 vdd.n1967 12.0247
R4472 vdd.n2053 vdd.n2026 12.0247
R4473 vdd.n1882 vdd.n1638 11.337
R4474 vdd.n1891 vdd.n1638 11.337
R4475 vdd.n1891 vdd.n1890 11.337
R4476 vdd.n1899 vdd.n1632 11.337
R4477 vdd.n1908 vdd.n1907 11.337
R4478 vdd.n1924 vdd.n1616 11.337
R4479 vdd.n1932 vdd.n1609 11.337
R4480 vdd.n1941 vdd.n1940 11.337
R4481 vdd.n1949 vdd.n1598 11.337
R4482 vdd.n2272 vdd.n1587 11.337
R4483 vdd.n2281 vdd.n1581 11.337
R4484 vdd.n2289 vdd.n1575 11.337
R4485 vdd.n2298 vdd.n2297 11.337
R4486 vdd.n2314 vdd.n1559 11.337
R4487 vdd.n2322 vdd.n1552 11.337
R4488 vdd.n2331 vdd.n2330 11.337
R4489 vdd.n2339 vdd.n1535 11.337
R4490 vdd.n2350 vdd.n1535 11.337
R4491 vdd.n2350 vdd.n2349 11.337
R4492 vdd.n3503 vdd.n678 11.337
R4493 vdd.n3511 vdd.n678 11.337
R4494 vdd.n3511 vdd.n679 11.337
R4495 vdd.n3520 vdd.n3519 11.337
R4496 vdd.n3536 vdd.n662 11.337
R4497 vdd.n3544 vdd.n655 11.337
R4498 vdd.n3553 vdd.n3552 11.337
R4499 vdd.n3561 vdd.n644 11.337
R4500 vdd.n3580 vdd.n633 11.337
R4501 vdd.n3667 vdd.n340 11.337
R4502 vdd.n3665 vdd.n344 11.337
R4503 vdd.n3659 vdd.n3658 11.337
R4504 vdd.n3651 vdd.n361 11.337
R4505 vdd.n3650 vdd.n3649 11.337
R4506 vdd.n3643 vdd.n3642 11.337
R4507 vdd.n3641 vdd.n375 11.337
R4508 vdd.n3635 vdd.n3634 11.337
R4509 vdd.n3634 vdd.n3633 11.337
R4510 vdd.n3633 vdd.n386 11.337
R4511 vdd.n320 vdd.n319 11.249
R4512 vdd.n261 vdd.n260 11.249
R4513 vdd.n218 vdd.n217 11.249
R4514 vdd.n159 vdd.n158 11.249
R4515 vdd.n117 vdd.n116 11.249
R4516 vdd.n58 vdd.n57 11.249
R4517 vdd.n2194 vdd.n2193 11.249
R4518 vdd.n2253 vdd.n2252 11.249
R4519 vdd.n2092 vdd.n2091 11.249
R4520 vdd.n2151 vdd.n2150 11.249
R4521 vdd.n1991 vdd.n1990 11.249
R4522 vdd.n2050 vdd.n2049 11.249
R4523 vdd.n1680 vdd.t211 11.2237
R4524 vdd.n3627 vdd.t160 11.2237
R4525 vdd.t15 vdd.n1553 10.7702
R4526 vdd.n3528 vdd.t29 10.7702
R4527 vdd.n305 vdd.n304 10.7238
R4528 vdd.n246 vdd.n245 10.7238
R4529 vdd.n203 vdd.n202 10.7238
R4530 vdd.n144 vdd.n143 10.7238
R4531 vdd.n102 vdd.n101 10.7238
R4532 vdd.n43 vdd.n42 10.7238
R4533 vdd.n2179 vdd.n2178 10.7238
R4534 vdd.n2238 vdd.n2237 10.7238
R4535 vdd.n2077 vdd.n2076 10.7238
R4536 vdd.n2136 vdd.n2135 10.7238
R4537 vdd.n1976 vdd.n1975 10.7238
R4538 vdd.n2035 vdd.n2034 10.7238
R4539 vdd.n2511 vdd.n2510 10.6151
R4540 vdd.n2511 vdd.n1127 10.6151
R4541 vdd.n2521 vdd.n1127 10.6151
R4542 vdd.n2522 vdd.n2521 10.6151
R4543 vdd.n2523 vdd.n2522 10.6151
R4544 vdd.n2523 vdd.n1114 10.6151
R4545 vdd.n2533 vdd.n1114 10.6151
R4546 vdd.n2534 vdd.n2533 10.6151
R4547 vdd.n2535 vdd.n2534 10.6151
R4548 vdd.n2535 vdd.n1102 10.6151
R4549 vdd.n2545 vdd.n1102 10.6151
R4550 vdd.n2546 vdd.n2545 10.6151
R4551 vdd.n2547 vdd.n2546 10.6151
R4552 vdd.n2547 vdd.n1091 10.6151
R4553 vdd.n2557 vdd.n1091 10.6151
R4554 vdd.n2558 vdd.n2557 10.6151
R4555 vdd.n2559 vdd.n2558 10.6151
R4556 vdd.n2559 vdd.n1078 10.6151
R4557 vdd.n2569 vdd.n1078 10.6151
R4558 vdd.n2570 vdd.n2569 10.6151
R4559 vdd.n2571 vdd.n2570 10.6151
R4560 vdd.n2571 vdd.n1066 10.6151
R4561 vdd.n2582 vdd.n1066 10.6151
R4562 vdd.n2583 vdd.n2582 10.6151
R4563 vdd.n2584 vdd.n2583 10.6151
R4564 vdd.n2584 vdd.n1054 10.6151
R4565 vdd.n2594 vdd.n1054 10.6151
R4566 vdd.n2595 vdd.n2594 10.6151
R4567 vdd.n2596 vdd.n2595 10.6151
R4568 vdd.n2596 vdd.n1042 10.6151
R4569 vdd.n2606 vdd.n1042 10.6151
R4570 vdd.n2607 vdd.n2606 10.6151
R4571 vdd.n2608 vdd.n2607 10.6151
R4572 vdd.n2608 vdd.n1032 10.6151
R4573 vdd.n2618 vdd.n1032 10.6151
R4574 vdd.n2619 vdd.n2618 10.6151
R4575 vdd.n2620 vdd.n2619 10.6151
R4576 vdd.n2620 vdd.n1019 10.6151
R4577 vdd.n2632 vdd.n1019 10.6151
R4578 vdd.n2633 vdd.n2632 10.6151
R4579 vdd.n2635 vdd.n2633 10.6151
R4580 vdd.n2635 vdd.n2634 10.6151
R4581 vdd.n2634 vdd.n1000 10.6151
R4582 vdd.n2782 vdd.n2781 10.6151
R4583 vdd.n2781 vdd.n2780 10.6151
R4584 vdd.n2780 vdd.n2777 10.6151
R4585 vdd.n2777 vdd.n2776 10.6151
R4586 vdd.n2776 vdd.n2773 10.6151
R4587 vdd.n2773 vdd.n2772 10.6151
R4588 vdd.n2772 vdd.n2769 10.6151
R4589 vdd.n2769 vdd.n2768 10.6151
R4590 vdd.n2768 vdd.n2765 10.6151
R4591 vdd.n2765 vdd.n2764 10.6151
R4592 vdd.n2764 vdd.n2761 10.6151
R4593 vdd.n2761 vdd.n2760 10.6151
R4594 vdd.n2760 vdd.n2757 10.6151
R4595 vdd.n2757 vdd.n2756 10.6151
R4596 vdd.n2756 vdd.n2753 10.6151
R4597 vdd.n2753 vdd.n2752 10.6151
R4598 vdd.n2752 vdd.n2749 10.6151
R4599 vdd.n2749 vdd.n2748 10.6151
R4600 vdd.n2748 vdd.n2745 10.6151
R4601 vdd.n2745 vdd.n2744 10.6151
R4602 vdd.n2744 vdd.n2741 10.6151
R4603 vdd.n2741 vdd.n2740 10.6151
R4604 vdd.n2740 vdd.n2737 10.6151
R4605 vdd.n2737 vdd.n2736 10.6151
R4606 vdd.n2736 vdd.n2733 10.6151
R4607 vdd.n2733 vdd.n2732 10.6151
R4608 vdd.n2732 vdd.n2729 10.6151
R4609 vdd.n2729 vdd.n2728 10.6151
R4610 vdd.n2728 vdd.n2725 10.6151
R4611 vdd.n2725 vdd.n2724 10.6151
R4612 vdd.n2724 vdd.n2721 10.6151
R4613 vdd.n2719 vdd.n2716 10.6151
R4614 vdd.n2716 vdd.n2715 10.6151
R4615 vdd.n1357 vdd.n1356 10.6151
R4616 vdd.n1359 vdd.n1357 10.6151
R4617 vdd.n1360 vdd.n1359 10.6151
R4618 vdd.n1362 vdd.n1360 10.6151
R4619 vdd.n1363 vdd.n1362 10.6151
R4620 vdd.n1365 vdd.n1363 10.6151
R4621 vdd.n1366 vdd.n1365 10.6151
R4622 vdd.n1368 vdd.n1366 10.6151
R4623 vdd.n1369 vdd.n1368 10.6151
R4624 vdd.n1371 vdd.n1369 10.6151
R4625 vdd.n1372 vdd.n1371 10.6151
R4626 vdd.n1374 vdd.n1372 10.6151
R4627 vdd.n1375 vdd.n1374 10.6151
R4628 vdd.n1377 vdd.n1375 10.6151
R4629 vdd.n1378 vdd.n1377 10.6151
R4630 vdd.n1380 vdd.n1378 10.6151
R4631 vdd.n1381 vdd.n1380 10.6151
R4632 vdd.n1383 vdd.n1381 10.6151
R4633 vdd.n1384 vdd.n1383 10.6151
R4634 vdd.n1386 vdd.n1384 10.6151
R4635 vdd.n1387 vdd.n1386 10.6151
R4636 vdd.n1389 vdd.n1387 10.6151
R4637 vdd.n1390 vdd.n1389 10.6151
R4638 vdd.n1392 vdd.n1390 10.6151
R4639 vdd.n1393 vdd.n1392 10.6151
R4640 vdd.n1395 vdd.n1393 10.6151
R4641 vdd.n1396 vdd.n1395 10.6151
R4642 vdd.n1435 vdd.n1396 10.6151
R4643 vdd.n1435 vdd.n1434 10.6151
R4644 vdd.n1434 vdd.n1433 10.6151
R4645 vdd.n1433 vdd.n1431 10.6151
R4646 vdd.n1431 vdd.n1430 10.6151
R4647 vdd.n1430 vdd.n1428 10.6151
R4648 vdd.n1428 vdd.n1427 10.6151
R4649 vdd.n1427 vdd.n1408 10.6151
R4650 vdd.n1408 vdd.n1407 10.6151
R4651 vdd.n1407 vdd.n1405 10.6151
R4652 vdd.n1405 vdd.n1404 10.6151
R4653 vdd.n1404 vdd.n1402 10.6151
R4654 vdd.n1402 vdd.n1401 10.6151
R4655 vdd.n1401 vdd.n1398 10.6151
R4656 vdd.n1398 vdd.n1397 10.6151
R4657 vdd.n1397 vdd.n1003 10.6151
R4658 vdd.n2509 vdd.n1139 10.6151
R4659 vdd.n2504 vdd.n1139 10.6151
R4660 vdd.n2504 vdd.n2503 10.6151
R4661 vdd.n2503 vdd.n2502 10.6151
R4662 vdd.n2502 vdd.n2499 10.6151
R4663 vdd.n2499 vdd.n2498 10.6151
R4664 vdd.n2498 vdd.n2495 10.6151
R4665 vdd.n2495 vdd.n2494 10.6151
R4666 vdd.n2494 vdd.n2491 10.6151
R4667 vdd.n2491 vdd.n2490 10.6151
R4668 vdd.n2490 vdd.n2487 10.6151
R4669 vdd.n2487 vdd.n2486 10.6151
R4670 vdd.n2486 vdd.n2483 10.6151
R4671 vdd.n2483 vdd.n2482 10.6151
R4672 vdd.n2482 vdd.n2479 10.6151
R4673 vdd.n2479 vdd.n2478 10.6151
R4674 vdd.n2478 vdd.n2475 10.6151
R4675 vdd.n2475 vdd.n1177 10.6151
R4676 vdd.n1323 vdd.n1177 10.6151
R4677 vdd.n1324 vdd.n1323 10.6151
R4678 vdd.n1327 vdd.n1324 10.6151
R4679 vdd.n1328 vdd.n1327 10.6151
R4680 vdd.n1331 vdd.n1328 10.6151
R4681 vdd.n1332 vdd.n1331 10.6151
R4682 vdd.n1335 vdd.n1332 10.6151
R4683 vdd.n1336 vdd.n1335 10.6151
R4684 vdd.n1339 vdd.n1336 10.6151
R4685 vdd.n1340 vdd.n1339 10.6151
R4686 vdd.n1343 vdd.n1340 10.6151
R4687 vdd.n1344 vdd.n1343 10.6151
R4688 vdd.n1347 vdd.n1344 10.6151
R4689 vdd.n1352 vdd.n1349 10.6151
R4690 vdd.n1353 vdd.n1352 10.6151
R4691 vdd.n3020 vdd.n3019 10.6151
R4692 vdd.n3019 vdd.n3018 10.6151
R4693 vdd.n3018 vdd.n2822 10.6151
R4694 vdd.n2900 vdd.n2822 10.6151
R4695 vdd.n2901 vdd.n2900 10.6151
R4696 vdd.n2903 vdd.n2901 10.6151
R4697 vdd.n2904 vdd.n2903 10.6151
R4698 vdd.n3002 vdd.n2904 10.6151
R4699 vdd.n3002 vdd.n3001 10.6151
R4700 vdd.n3001 vdd.n3000 10.6151
R4701 vdd.n3000 vdd.n2948 10.6151
R4702 vdd.n2948 vdd.n2947 10.6151
R4703 vdd.n2947 vdd.n2945 10.6151
R4704 vdd.n2945 vdd.n2944 10.6151
R4705 vdd.n2944 vdd.n2942 10.6151
R4706 vdd.n2942 vdd.n2941 10.6151
R4707 vdd.n2941 vdd.n2939 10.6151
R4708 vdd.n2939 vdd.n2938 10.6151
R4709 vdd.n2938 vdd.n2936 10.6151
R4710 vdd.n2936 vdd.n2935 10.6151
R4711 vdd.n2935 vdd.n2933 10.6151
R4712 vdd.n2933 vdd.n2932 10.6151
R4713 vdd.n2932 vdd.n2930 10.6151
R4714 vdd.n2930 vdd.n2929 10.6151
R4715 vdd.n2929 vdd.n2927 10.6151
R4716 vdd.n2927 vdd.n2926 10.6151
R4717 vdd.n2926 vdd.n2924 10.6151
R4718 vdd.n2924 vdd.n2923 10.6151
R4719 vdd.n2923 vdd.n2921 10.6151
R4720 vdd.n2921 vdd.n2920 10.6151
R4721 vdd.n2920 vdd.n2918 10.6151
R4722 vdd.n2918 vdd.n2917 10.6151
R4723 vdd.n2917 vdd.n2915 10.6151
R4724 vdd.n2915 vdd.n2914 10.6151
R4725 vdd.n2914 vdd.n2912 10.6151
R4726 vdd.n2912 vdd.n2911 10.6151
R4727 vdd.n2911 vdd.n2909 10.6151
R4728 vdd.n2909 vdd.n2908 10.6151
R4729 vdd.n2908 vdd.n2906 10.6151
R4730 vdd.n2906 vdd.n2905 10.6151
R4731 vdd.n2905 vdd.n836 10.6151
R4732 vdd.n3264 vdd.n836 10.6151
R4733 vdd.n3265 vdd.n3264 10.6151
R4734 vdd.n3091 vdd.n961 10.6151
R4735 vdd.n3086 vdd.n961 10.6151
R4736 vdd.n3086 vdd.n3085 10.6151
R4737 vdd.n3085 vdd.n3084 10.6151
R4738 vdd.n3084 vdd.n3081 10.6151
R4739 vdd.n3081 vdd.n3080 10.6151
R4740 vdd.n3080 vdd.n3077 10.6151
R4741 vdd.n3077 vdd.n3076 10.6151
R4742 vdd.n3076 vdd.n3073 10.6151
R4743 vdd.n3073 vdd.n3072 10.6151
R4744 vdd.n3072 vdd.n3069 10.6151
R4745 vdd.n3069 vdd.n3068 10.6151
R4746 vdd.n3068 vdd.n3065 10.6151
R4747 vdd.n3065 vdd.n3064 10.6151
R4748 vdd.n3064 vdd.n3061 10.6151
R4749 vdd.n3061 vdd.n3060 10.6151
R4750 vdd.n3060 vdd.n3057 10.6151
R4751 vdd.n3057 vdd.n3056 10.6151
R4752 vdd.n3056 vdd.n3053 10.6151
R4753 vdd.n3053 vdd.n3052 10.6151
R4754 vdd.n3052 vdd.n3049 10.6151
R4755 vdd.n3049 vdd.n3048 10.6151
R4756 vdd.n3048 vdd.n3045 10.6151
R4757 vdd.n3045 vdd.n3044 10.6151
R4758 vdd.n3044 vdd.n3041 10.6151
R4759 vdd.n3041 vdd.n3040 10.6151
R4760 vdd.n3040 vdd.n3037 10.6151
R4761 vdd.n3037 vdd.n3036 10.6151
R4762 vdd.n3036 vdd.n3033 10.6151
R4763 vdd.n3033 vdd.n3032 10.6151
R4764 vdd.n3032 vdd.n3029 10.6151
R4765 vdd.n3027 vdd.n3024 10.6151
R4766 vdd.n3024 vdd.n3023 10.6151
R4767 vdd.n3093 vdd.n3092 10.6151
R4768 vdd.n3093 vdd.n950 10.6151
R4769 vdd.n3103 vdd.n950 10.6151
R4770 vdd.n3104 vdd.n3103 10.6151
R4771 vdd.n3105 vdd.n3104 10.6151
R4772 vdd.n3105 vdd.n938 10.6151
R4773 vdd.n3115 vdd.n938 10.6151
R4774 vdd.n3116 vdd.n3115 10.6151
R4775 vdd.n3117 vdd.n3116 10.6151
R4776 vdd.n3117 vdd.n927 10.6151
R4777 vdd.n3127 vdd.n927 10.6151
R4778 vdd.n3128 vdd.n3127 10.6151
R4779 vdd.n3129 vdd.n3128 10.6151
R4780 vdd.n3129 vdd.n916 10.6151
R4781 vdd.n3139 vdd.n916 10.6151
R4782 vdd.n3140 vdd.n3139 10.6151
R4783 vdd.n3141 vdd.n3140 10.6151
R4784 vdd.n3141 vdd.n903 10.6151
R4785 vdd.n3152 vdd.n903 10.6151
R4786 vdd.n3153 vdd.n3152 10.6151
R4787 vdd.n3154 vdd.n3153 10.6151
R4788 vdd.n3154 vdd.n891 10.6151
R4789 vdd.n3164 vdd.n891 10.6151
R4790 vdd.n3165 vdd.n3164 10.6151
R4791 vdd.n3166 vdd.n3165 10.6151
R4792 vdd.n3166 vdd.n879 10.6151
R4793 vdd.n3176 vdd.n879 10.6151
R4794 vdd.n3177 vdd.n3176 10.6151
R4795 vdd.n3178 vdd.n3177 10.6151
R4796 vdd.n3178 vdd.n866 10.6151
R4797 vdd.n3188 vdd.n866 10.6151
R4798 vdd.n3189 vdd.n3188 10.6151
R4799 vdd.n3190 vdd.n3189 10.6151
R4800 vdd.n3190 vdd.n855 10.6151
R4801 vdd.n3200 vdd.n855 10.6151
R4802 vdd.n3201 vdd.n3200 10.6151
R4803 vdd.n3202 vdd.n3201 10.6151
R4804 vdd.n3202 vdd.n841 10.6151
R4805 vdd.n3257 vdd.n841 10.6151
R4806 vdd.n3258 vdd.n3257 10.6151
R4807 vdd.n3259 vdd.n3258 10.6151
R4808 vdd.n3259 vdd.n810 10.6151
R4809 vdd.n3329 vdd.n810 10.6151
R4810 vdd.n3328 vdd.n3327 10.6151
R4811 vdd.n3327 vdd.n811 10.6151
R4812 vdd.n812 vdd.n811 10.6151
R4813 vdd.n3320 vdd.n812 10.6151
R4814 vdd.n3320 vdd.n3319 10.6151
R4815 vdd.n3319 vdd.n3318 10.6151
R4816 vdd.n3318 vdd.n814 10.6151
R4817 vdd.n3313 vdd.n814 10.6151
R4818 vdd.n3313 vdd.n3312 10.6151
R4819 vdd.n3312 vdd.n3311 10.6151
R4820 vdd.n3311 vdd.n817 10.6151
R4821 vdd.n3306 vdd.n817 10.6151
R4822 vdd.n3306 vdd.n3305 10.6151
R4823 vdd.n3305 vdd.n3304 10.6151
R4824 vdd.n3304 vdd.n820 10.6151
R4825 vdd.n3299 vdd.n820 10.6151
R4826 vdd.n3299 vdd.n731 10.6151
R4827 vdd.n3295 vdd.n731 10.6151
R4828 vdd.n3295 vdd.n3294 10.6151
R4829 vdd.n3294 vdd.n3293 10.6151
R4830 vdd.n3293 vdd.n823 10.6151
R4831 vdd.n3288 vdd.n823 10.6151
R4832 vdd.n3288 vdd.n3287 10.6151
R4833 vdd.n3287 vdd.n3286 10.6151
R4834 vdd.n3286 vdd.n826 10.6151
R4835 vdd.n3281 vdd.n826 10.6151
R4836 vdd.n3281 vdd.n3280 10.6151
R4837 vdd.n3280 vdd.n3279 10.6151
R4838 vdd.n3279 vdd.n829 10.6151
R4839 vdd.n3274 vdd.n829 10.6151
R4840 vdd.n3274 vdd.n3273 10.6151
R4841 vdd.n3271 vdd.n834 10.6151
R4842 vdd.n3266 vdd.n834 10.6151
R4843 vdd.n3247 vdd.n3208 10.6151
R4844 vdd.n3242 vdd.n3208 10.6151
R4845 vdd.n3242 vdd.n3241 10.6151
R4846 vdd.n3241 vdd.n3240 10.6151
R4847 vdd.n3240 vdd.n3210 10.6151
R4848 vdd.n3235 vdd.n3210 10.6151
R4849 vdd.n3235 vdd.n3234 10.6151
R4850 vdd.n3234 vdd.n3233 10.6151
R4851 vdd.n3233 vdd.n3213 10.6151
R4852 vdd.n3228 vdd.n3213 10.6151
R4853 vdd.n3228 vdd.n3227 10.6151
R4854 vdd.n3227 vdd.n3226 10.6151
R4855 vdd.n3226 vdd.n3216 10.6151
R4856 vdd.n3221 vdd.n3216 10.6151
R4857 vdd.n3221 vdd.n3220 10.6151
R4858 vdd.n3220 vdd.n785 10.6151
R4859 vdd.n3364 vdd.n785 10.6151
R4860 vdd.n3364 vdd.n786 10.6151
R4861 vdd.n788 vdd.n786 10.6151
R4862 vdd.n3357 vdd.n788 10.6151
R4863 vdd.n3357 vdd.n3356 10.6151
R4864 vdd.n3356 vdd.n3355 10.6151
R4865 vdd.n3355 vdd.n790 10.6151
R4866 vdd.n3350 vdd.n790 10.6151
R4867 vdd.n3350 vdd.n3349 10.6151
R4868 vdd.n3349 vdd.n3348 10.6151
R4869 vdd.n3348 vdd.n793 10.6151
R4870 vdd.n3343 vdd.n793 10.6151
R4871 vdd.n3343 vdd.n3342 10.6151
R4872 vdd.n3342 vdd.n3341 10.6151
R4873 vdd.n3341 vdd.n796 10.6151
R4874 vdd.n3336 vdd.n3335 10.6151
R4875 vdd.n3335 vdd.n3334 10.6151
R4876 vdd.n2897 vdd.n2896 10.6151
R4877 vdd.n3014 vdd.n2897 10.6151
R4878 vdd.n3014 vdd.n3013 10.6151
R4879 vdd.n3013 vdd.n3012 10.6151
R4880 vdd.n3012 vdd.n3010 10.6151
R4881 vdd.n3010 vdd.n3009 10.6151
R4882 vdd.n3009 vdd.n3007 10.6151
R4883 vdd.n3007 vdd.n3006 10.6151
R4884 vdd.n3006 vdd.n2898 10.6151
R4885 vdd.n2996 vdd.n2898 10.6151
R4886 vdd.n2996 vdd.n2995 10.6151
R4887 vdd.n2995 vdd.n2994 10.6151
R4888 vdd.n2994 vdd.n2992 10.6151
R4889 vdd.n2992 vdd.n2991 10.6151
R4890 vdd.n2991 vdd.n2989 10.6151
R4891 vdd.n2989 vdd.n2988 10.6151
R4892 vdd.n2988 vdd.n2986 10.6151
R4893 vdd.n2986 vdd.n2985 10.6151
R4894 vdd.n2985 vdd.n2983 10.6151
R4895 vdd.n2983 vdd.n2982 10.6151
R4896 vdd.n2982 vdd.n2980 10.6151
R4897 vdd.n2980 vdd.n2979 10.6151
R4898 vdd.n2979 vdd.n2977 10.6151
R4899 vdd.n2977 vdd.n2976 10.6151
R4900 vdd.n2976 vdd.n2974 10.6151
R4901 vdd.n2974 vdd.n2973 10.6151
R4902 vdd.n2973 vdd.n2971 10.6151
R4903 vdd.n2971 vdd.n2970 10.6151
R4904 vdd.n2970 vdd.n2968 10.6151
R4905 vdd.n2968 vdd.n2967 10.6151
R4906 vdd.n2967 vdd.n2965 10.6151
R4907 vdd.n2965 vdd.n2964 10.6151
R4908 vdd.n2964 vdd.n2962 10.6151
R4909 vdd.n2962 vdd.n2961 10.6151
R4910 vdd.n2961 vdd.n2959 10.6151
R4911 vdd.n2959 vdd.n2958 10.6151
R4912 vdd.n2958 vdd.n2956 10.6151
R4913 vdd.n2956 vdd.n2955 10.6151
R4914 vdd.n2955 vdd.n2953 10.6151
R4915 vdd.n2953 vdd.n2952 10.6151
R4916 vdd.n2952 vdd.n2950 10.6151
R4917 vdd.n2950 vdd.n2949 10.6151
R4918 vdd.n2949 vdd.n802 10.6151
R4919 vdd.n2828 vdd.n2827 10.6151
R4920 vdd.n2831 vdd.n2828 10.6151
R4921 vdd.n2832 vdd.n2831 10.6151
R4922 vdd.n2835 vdd.n2832 10.6151
R4923 vdd.n2836 vdd.n2835 10.6151
R4924 vdd.n2839 vdd.n2836 10.6151
R4925 vdd.n2840 vdd.n2839 10.6151
R4926 vdd.n2843 vdd.n2840 10.6151
R4927 vdd.n2844 vdd.n2843 10.6151
R4928 vdd.n2847 vdd.n2844 10.6151
R4929 vdd.n2848 vdd.n2847 10.6151
R4930 vdd.n2851 vdd.n2848 10.6151
R4931 vdd.n2852 vdd.n2851 10.6151
R4932 vdd.n2855 vdd.n2852 10.6151
R4933 vdd.n2856 vdd.n2855 10.6151
R4934 vdd.n2859 vdd.n2856 10.6151
R4935 vdd.n2860 vdd.n2859 10.6151
R4936 vdd.n2863 vdd.n2860 10.6151
R4937 vdd.n2864 vdd.n2863 10.6151
R4938 vdd.n2867 vdd.n2864 10.6151
R4939 vdd.n2868 vdd.n2867 10.6151
R4940 vdd.n2871 vdd.n2868 10.6151
R4941 vdd.n2872 vdd.n2871 10.6151
R4942 vdd.n2875 vdd.n2872 10.6151
R4943 vdd.n2876 vdd.n2875 10.6151
R4944 vdd.n2879 vdd.n2876 10.6151
R4945 vdd.n2880 vdd.n2879 10.6151
R4946 vdd.n2883 vdd.n2880 10.6151
R4947 vdd.n2884 vdd.n2883 10.6151
R4948 vdd.n2887 vdd.n2884 10.6151
R4949 vdd.n2888 vdd.n2887 10.6151
R4950 vdd.n2893 vdd.n2891 10.6151
R4951 vdd.n2894 vdd.n2893 10.6151
R4952 vdd.n3097 vdd.n955 10.6151
R4953 vdd.n3098 vdd.n3097 10.6151
R4954 vdd.n3099 vdd.n3098 10.6151
R4955 vdd.n3099 vdd.n944 10.6151
R4956 vdd.n3109 vdd.n944 10.6151
R4957 vdd.n3110 vdd.n3109 10.6151
R4958 vdd.n3111 vdd.n3110 10.6151
R4959 vdd.n3111 vdd.n933 10.6151
R4960 vdd.n3121 vdd.n933 10.6151
R4961 vdd.n3122 vdd.n3121 10.6151
R4962 vdd.n3123 vdd.n3122 10.6151
R4963 vdd.n3123 vdd.n921 10.6151
R4964 vdd.n3133 vdd.n921 10.6151
R4965 vdd.n3134 vdd.n3133 10.6151
R4966 vdd.n3135 vdd.n3134 10.6151
R4967 vdd.n3135 vdd.n910 10.6151
R4968 vdd.n3145 vdd.n910 10.6151
R4969 vdd.n3146 vdd.n3145 10.6151
R4970 vdd.n3148 vdd.n3146 10.6151
R4971 vdd.n3148 vdd.n3147 10.6151
R4972 vdd.n3159 vdd.n3158 10.6151
R4973 vdd.n3160 vdd.n3159 10.6151
R4974 vdd.n3160 vdd.n885 10.6151
R4975 vdd.n3170 vdd.n885 10.6151
R4976 vdd.n3171 vdd.n3170 10.6151
R4977 vdd.n3172 vdd.n3171 10.6151
R4978 vdd.n3172 vdd.n872 10.6151
R4979 vdd.n3182 vdd.n872 10.6151
R4980 vdd.n3183 vdd.n3182 10.6151
R4981 vdd.n3184 vdd.n3183 10.6151
R4982 vdd.n3184 vdd.n860 10.6151
R4983 vdd.n3194 vdd.n860 10.6151
R4984 vdd.n3195 vdd.n3194 10.6151
R4985 vdd.n3196 vdd.n3195 10.6151
R4986 vdd.n3196 vdd.n849 10.6151
R4987 vdd.n3206 vdd.n849 10.6151
R4988 vdd.n3207 vdd.n3206 10.6151
R4989 vdd.n3253 vdd.n3207 10.6151
R4990 vdd.n3253 vdd.n3252 10.6151
R4991 vdd.n3252 vdd.n3251 10.6151
R4992 vdd.n3251 vdd.n3250 10.6151
R4993 vdd.n3250 vdd.n3248 10.6151
R4994 vdd.n2515 vdd.n1132 10.6151
R4995 vdd.n2516 vdd.n2515 10.6151
R4996 vdd.n2517 vdd.n2516 10.6151
R4997 vdd.n2517 vdd.n1121 10.6151
R4998 vdd.n2527 vdd.n1121 10.6151
R4999 vdd.n2528 vdd.n2527 10.6151
R5000 vdd.n2529 vdd.n2528 10.6151
R5001 vdd.n2529 vdd.n1108 10.6151
R5002 vdd.n2539 vdd.n1108 10.6151
R5003 vdd.n2540 vdd.n2539 10.6151
R5004 vdd.n2541 vdd.n2540 10.6151
R5005 vdd.n2541 vdd.n1097 10.6151
R5006 vdd.n2551 vdd.n1097 10.6151
R5007 vdd.n2552 vdd.n2551 10.6151
R5008 vdd.n2553 vdd.n2552 10.6151
R5009 vdd.n2553 vdd.n1085 10.6151
R5010 vdd.n2563 vdd.n1085 10.6151
R5011 vdd.n2564 vdd.n2563 10.6151
R5012 vdd.n2565 vdd.n2564 10.6151
R5013 vdd.n2565 vdd.n1072 10.6151
R5014 vdd.n2575 vdd.n1072 10.6151
R5015 vdd.n2576 vdd.n2575 10.6151
R5016 vdd.n2578 vdd.n1060 10.6151
R5017 vdd.n2588 vdd.n1060 10.6151
R5018 vdd.n2589 vdd.n2588 10.6151
R5019 vdd.n2590 vdd.n2589 10.6151
R5020 vdd.n2590 vdd.n1048 10.6151
R5021 vdd.n2600 vdd.n1048 10.6151
R5022 vdd.n2601 vdd.n2600 10.6151
R5023 vdd.n2602 vdd.n2601 10.6151
R5024 vdd.n2602 vdd.n1037 10.6151
R5025 vdd.n2612 vdd.n1037 10.6151
R5026 vdd.n2613 vdd.n2612 10.6151
R5027 vdd.n2614 vdd.n2613 10.6151
R5028 vdd.n2614 vdd.n1026 10.6151
R5029 vdd.n2624 vdd.n1026 10.6151
R5030 vdd.n2625 vdd.n2624 10.6151
R5031 vdd.n2628 vdd.n2625 10.6151
R5032 vdd.n2628 vdd.n2627 10.6151
R5033 vdd.n2627 vdd.n2626 10.6151
R5034 vdd.n2626 vdd.n1009 10.6151
R5035 vdd.n2710 vdd.n1009 10.6151
R5036 vdd.n2709 vdd.n2708 10.6151
R5037 vdd.n2708 vdd.n2705 10.6151
R5038 vdd.n2705 vdd.n2704 10.6151
R5039 vdd.n2704 vdd.n2701 10.6151
R5040 vdd.n2701 vdd.n2700 10.6151
R5041 vdd.n2700 vdd.n2697 10.6151
R5042 vdd.n2697 vdd.n2696 10.6151
R5043 vdd.n2696 vdd.n2693 10.6151
R5044 vdd.n2693 vdd.n2692 10.6151
R5045 vdd.n2692 vdd.n2689 10.6151
R5046 vdd.n2689 vdd.n2688 10.6151
R5047 vdd.n2688 vdd.n2685 10.6151
R5048 vdd.n2685 vdd.n2684 10.6151
R5049 vdd.n2684 vdd.n2681 10.6151
R5050 vdd.n2681 vdd.n2680 10.6151
R5051 vdd.n2680 vdd.n2677 10.6151
R5052 vdd.n2677 vdd.n2676 10.6151
R5053 vdd.n2676 vdd.n2673 10.6151
R5054 vdd.n2673 vdd.n2672 10.6151
R5055 vdd.n2672 vdd.n2669 10.6151
R5056 vdd.n2669 vdd.n2668 10.6151
R5057 vdd.n2668 vdd.n2665 10.6151
R5058 vdd.n2665 vdd.n2664 10.6151
R5059 vdd.n2664 vdd.n2661 10.6151
R5060 vdd.n2661 vdd.n2660 10.6151
R5061 vdd.n2660 vdd.n2657 10.6151
R5062 vdd.n2657 vdd.n2656 10.6151
R5063 vdd.n2656 vdd.n2653 10.6151
R5064 vdd.n2653 vdd.n2652 10.6151
R5065 vdd.n2652 vdd.n2649 10.6151
R5066 vdd.n2649 vdd.n2648 10.6151
R5067 vdd.n2645 vdd.n2644 10.6151
R5068 vdd.n2644 vdd.n2642 10.6151
R5069 vdd.n1481 vdd.n1479 10.6151
R5070 vdd.n1479 vdd.n1478 10.6151
R5071 vdd.n1478 vdd.n1476 10.6151
R5072 vdd.n1476 vdd.n1475 10.6151
R5073 vdd.n1475 vdd.n1473 10.6151
R5074 vdd.n1473 vdd.n1472 10.6151
R5075 vdd.n1472 vdd.n1470 10.6151
R5076 vdd.n1470 vdd.n1469 10.6151
R5077 vdd.n1469 vdd.n1467 10.6151
R5078 vdd.n1467 vdd.n1466 10.6151
R5079 vdd.n1466 vdd.n1464 10.6151
R5080 vdd.n1464 vdd.n1463 10.6151
R5081 vdd.n1463 vdd.n1461 10.6151
R5082 vdd.n1461 vdd.n1460 10.6151
R5083 vdd.n1460 vdd.n1458 10.6151
R5084 vdd.n1458 vdd.n1457 10.6151
R5085 vdd.n1457 vdd.n1455 10.6151
R5086 vdd.n1455 vdd.n1454 10.6151
R5087 vdd.n1454 vdd.n1452 10.6151
R5088 vdd.n1452 vdd.n1451 10.6151
R5089 vdd.n1451 vdd.n1449 10.6151
R5090 vdd.n1449 vdd.n1448 10.6151
R5091 vdd.n1448 vdd.n1446 10.6151
R5092 vdd.n1446 vdd.n1445 10.6151
R5093 vdd.n1445 vdd.n1443 10.6151
R5094 vdd.n1443 vdd.n1442 10.6151
R5095 vdd.n1442 vdd.n1440 10.6151
R5096 vdd.n1440 vdd.n1439 10.6151
R5097 vdd.n1439 vdd.n1318 10.6151
R5098 vdd.n1410 vdd.n1318 10.6151
R5099 vdd.n1411 vdd.n1410 10.6151
R5100 vdd.n1413 vdd.n1411 10.6151
R5101 vdd.n1414 vdd.n1413 10.6151
R5102 vdd.n1423 vdd.n1414 10.6151
R5103 vdd.n1423 vdd.n1422 10.6151
R5104 vdd.n1422 vdd.n1421 10.6151
R5105 vdd.n1421 vdd.n1419 10.6151
R5106 vdd.n1419 vdd.n1418 10.6151
R5107 vdd.n1418 vdd.n1416 10.6151
R5108 vdd.n1416 vdd.n1415 10.6151
R5109 vdd.n1415 vdd.n1013 10.6151
R5110 vdd.n2640 vdd.n1013 10.6151
R5111 vdd.n2641 vdd.n2640 10.6151
R5112 vdd.n1282 vdd.n1281 10.6151
R5113 vdd.n1285 vdd.n1282 10.6151
R5114 vdd.n1286 vdd.n1285 10.6151
R5115 vdd.n1289 vdd.n1286 10.6151
R5116 vdd.n1290 vdd.n1289 10.6151
R5117 vdd.n1293 vdd.n1290 10.6151
R5118 vdd.n1294 vdd.n1293 10.6151
R5119 vdd.n1297 vdd.n1294 10.6151
R5120 vdd.n1298 vdd.n1297 10.6151
R5121 vdd.n1301 vdd.n1298 10.6151
R5122 vdd.n1302 vdd.n1301 10.6151
R5123 vdd.n1305 vdd.n1302 10.6151
R5124 vdd.n1306 vdd.n1305 10.6151
R5125 vdd.n1309 vdd.n1306 10.6151
R5126 vdd.n1310 vdd.n1309 10.6151
R5127 vdd.n1313 vdd.n1310 10.6151
R5128 vdd.n1515 vdd.n1313 10.6151
R5129 vdd.n1515 vdd.n1514 10.6151
R5130 vdd.n1514 vdd.n1512 10.6151
R5131 vdd.n1512 vdd.n1509 10.6151
R5132 vdd.n1509 vdd.n1508 10.6151
R5133 vdd.n1508 vdd.n1505 10.6151
R5134 vdd.n1505 vdd.n1504 10.6151
R5135 vdd.n1504 vdd.n1501 10.6151
R5136 vdd.n1501 vdd.n1500 10.6151
R5137 vdd.n1500 vdd.n1497 10.6151
R5138 vdd.n1497 vdd.n1496 10.6151
R5139 vdd.n1496 vdd.n1493 10.6151
R5140 vdd.n1493 vdd.n1492 10.6151
R5141 vdd.n1492 vdd.n1489 10.6151
R5142 vdd.n1489 vdd.n1488 10.6151
R5143 vdd.n1485 vdd.n1484 10.6151
R5144 vdd.n1484 vdd.n1482 10.6151
R5145 vdd.n2306 vdd.t52 10.5435
R5146 vdd.n656 vdd.t103 10.5435
R5147 vdd.n316 vdd.n298 10.4732
R5148 vdd.n257 vdd.n239 10.4732
R5149 vdd.n214 vdd.n196 10.4732
R5150 vdd.n155 vdd.n137 10.4732
R5151 vdd.n113 vdd.n95 10.4732
R5152 vdd.n54 vdd.n36 10.4732
R5153 vdd.n2190 vdd.n2172 10.4732
R5154 vdd.n2249 vdd.n2231 10.4732
R5155 vdd.n2088 vdd.n2070 10.4732
R5156 vdd.n2147 vdd.n2129 10.4732
R5157 vdd.n1987 vdd.n1969 10.4732
R5158 vdd.n2046 vdd.n2028 10.4732
R5159 vdd.t49 vdd.n2280 10.3167
R5160 vdd.n3572 vdd.t119 10.3167
R5161 vdd.n1957 vdd.t35 10.09
R5162 vdd.n3666 vdd.t33 10.09
R5163 vdd.n2475 vdd.n2474 9.98956
R5164 vdd.n3488 vdd.n731 9.98956
R5165 vdd.n3365 vdd.n3364 9.98956
R5166 vdd.n2367 vdd.n1515 9.98956
R5167 vdd.t56 vdd.n1610 9.86327
R5168 vdd.n3657 vdd.t79 9.86327
R5169 vdd.n2712 vdd.t271 9.7499
R5170 vdd.t256 vdd.n957 9.7499
R5171 vdd.n315 vdd.n300 9.69747
R5172 vdd.n256 vdd.n241 9.69747
R5173 vdd.n213 vdd.n198 9.69747
R5174 vdd.n154 vdd.n139 9.69747
R5175 vdd.n112 vdd.n97 9.69747
R5176 vdd.n53 vdd.n38 9.69747
R5177 vdd.n2189 vdd.n2174 9.69747
R5178 vdd.n2248 vdd.n2233 9.69747
R5179 vdd.n2087 vdd.n2072 9.69747
R5180 vdd.n2146 vdd.n2131 9.69747
R5181 vdd.n1986 vdd.n1971 9.69747
R5182 vdd.n2045 vdd.n2030 9.69747
R5183 vdd.n1916 vdd.t106 9.63654
R5184 vdd.n3603 vdd.t0 9.63654
R5185 vdd.n331 vdd.n330 9.45567
R5186 vdd.n272 vdd.n271 9.45567
R5187 vdd.n229 vdd.n228 9.45567
R5188 vdd.n170 vdd.n169 9.45567
R5189 vdd.n128 vdd.n127 9.45567
R5190 vdd.n69 vdd.n68 9.45567
R5191 vdd.n2205 vdd.n2204 9.45567
R5192 vdd.n2264 vdd.n2263 9.45567
R5193 vdd.n2103 vdd.n2102 9.45567
R5194 vdd.n2162 vdd.n2161 9.45567
R5195 vdd.n2002 vdd.n2001 9.45567
R5196 vdd.n2061 vdd.n2060 9.45567
R5197 vdd.n1890 vdd.t66 9.40981
R5198 vdd.n3635 vdd.t70 9.40981
R5199 vdd.n2437 vdd.n1207 9.3005
R5200 vdd.n2436 vdd.n2435 9.3005
R5201 vdd.n1213 vdd.n1212 9.3005
R5202 vdd.n2430 vdd.n1217 9.3005
R5203 vdd.n2429 vdd.n1218 9.3005
R5204 vdd.n2428 vdd.n1219 9.3005
R5205 vdd.n1223 vdd.n1220 9.3005
R5206 vdd.n2423 vdd.n1224 9.3005
R5207 vdd.n2422 vdd.n1225 9.3005
R5208 vdd.n2421 vdd.n1226 9.3005
R5209 vdd.n1230 vdd.n1227 9.3005
R5210 vdd.n2416 vdd.n1231 9.3005
R5211 vdd.n2415 vdd.n1232 9.3005
R5212 vdd.n2414 vdd.n1233 9.3005
R5213 vdd.n1237 vdd.n1234 9.3005
R5214 vdd.n2409 vdd.n1238 9.3005
R5215 vdd.n2408 vdd.n1239 9.3005
R5216 vdd.n2407 vdd.n1240 9.3005
R5217 vdd.n1244 vdd.n1241 9.3005
R5218 vdd.n2402 vdd.n1245 9.3005
R5219 vdd.n2401 vdd.n1246 9.3005
R5220 vdd.n2400 vdd.n2399 9.3005
R5221 vdd.n2398 vdd.n1247 9.3005
R5222 vdd.n2397 vdd.n2396 9.3005
R5223 vdd.n1253 vdd.n1252 9.3005
R5224 vdd.n2391 vdd.n1257 9.3005
R5225 vdd.n2390 vdd.n1258 9.3005
R5226 vdd.n2389 vdd.n1259 9.3005
R5227 vdd.n1263 vdd.n1260 9.3005
R5228 vdd.n2384 vdd.n1264 9.3005
R5229 vdd.n2383 vdd.n1265 9.3005
R5230 vdd.n2382 vdd.n1266 9.3005
R5231 vdd.n1270 vdd.n1267 9.3005
R5232 vdd.n2377 vdd.n1271 9.3005
R5233 vdd.n2376 vdd.n1272 9.3005
R5234 vdd.n2375 vdd.n1273 9.3005
R5235 vdd.n1277 vdd.n1274 9.3005
R5236 vdd.n2370 vdd.n1278 9.3005
R5237 vdd.n2439 vdd.n2438 9.3005
R5238 vdd.n2461 vdd.n1178 9.3005
R5239 vdd.n2460 vdd.n1186 9.3005
R5240 vdd.n1190 vdd.n1187 9.3005
R5241 vdd.n2455 vdd.n1191 9.3005
R5242 vdd.n2454 vdd.n1192 9.3005
R5243 vdd.n2453 vdd.n1193 9.3005
R5244 vdd.n1197 vdd.n1194 9.3005
R5245 vdd.n2448 vdd.n1198 9.3005
R5246 vdd.n2447 vdd.n1199 9.3005
R5247 vdd.n2446 vdd.n1200 9.3005
R5248 vdd.n1204 vdd.n1201 9.3005
R5249 vdd.n2441 vdd.n1205 9.3005
R5250 vdd.n2440 vdd.n1206 9.3005
R5251 vdd.n2473 vdd.n2472 9.3005
R5252 vdd.n1182 vdd.n1181 9.3005
R5253 vdd.n2270 vdd.n2269 9.3005
R5254 vdd.n1579 vdd.n1578 9.3005
R5255 vdd.n2284 vdd.n2283 9.3005
R5256 vdd.n2285 vdd.n1577 9.3005
R5257 vdd.n2287 vdd.n2286 9.3005
R5258 vdd.n1568 vdd.n1567 9.3005
R5259 vdd.n2301 vdd.n2300 9.3005
R5260 vdd.n2302 vdd.n1566 9.3005
R5261 vdd.n2304 vdd.n2303 9.3005
R5262 vdd.n1557 vdd.n1556 9.3005
R5263 vdd.n2317 vdd.n2316 9.3005
R5264 vdd.n2318 vdd.n1555 9.3005
R5265 vdd.n2320 vdd.n2319 9.3005
R5266 vdd.n1545 vdd.n1544 9.3005
R5267 vdd.n2334 vdd.n2333 9.3005
R5268 vdd.n2335 vdd.n1543 9.3005
R5269 vdd.n2337 vdd.n2336 9.3005
R5270 vdd.n1533 vdd.n1532 9.3005
R5271 vdd.n2353 vdd.n2352 9.3005
R5272 vdd.n2354 vdd.n1531 9.3005
R5273 vdd.n2356 vdd.n2355 9.3005
R5274 vdd.n307 vdd.n306 9.3005
R5275 vdd.n302 vdd.n301 9.3005
R5276 vdd.n313 vdd.n312 9.3005
R5277 vdd.n315 vdd.n314 9.3005
R5278 vdd.n298 vdd.n297 9.3005
R5279 vdd.n321 vdd.n320 9.3005
R5280 vdd.n323 vdd.n322 9.3005
R5281 vdd.n295 vdd.n292 9.3005
R5282 vdd.n330 vdd.n329 9.3005
R5283 vdd.n248 vdd.n247 9.3005
R5284 vdd.n243 vdd.n242 9.3005
R5285 vdd.n254 vdd.n253 9.3005
R5286 vdd.n256 vdd.n255 9.3005
R5287 vdd.n239 vdd.n238 9.3005
R5288 vdd.n262 vdd.n261 9.3005
R5289 vdd.n264 vdd.n263 9.3005
R5290 vdd.n236 vdd.n233 9.3005
R5291 vdd.n271 vdd.n270 9.3005
R5292 vdd.n205 vdd.n204 9.3005
R5293 vdd.n200 vdd.n199 9.3005
R5294 vdd.n211 vdd.n210 9.3005
R5295 vdd.n213 vdd.n212 9.3005
R5296 vdd.n196 vdd.n195 9.3005
R5297 vdd.n219 vdd.n218 9.3005
R5298 vdd.n221 vdd.n220 9.3005
R5299 vdd.n193 vdd.n190 9.3005
R5300 vdd.n228 vdd.n227 9.3005
R5301 vdd.n146 vdd.n145 9.3005
R5302 vdd.n141 vdd.n140 9.3005
R5303 vdd.n152 vdd.n151 9.3005
R5304 vdd.n154 vdd.n153 9.3005
R5305 vdd.n137 vdd.n136 9.3005
R5306 vdd.n160 vdd.n159 9.3005
R5307 vdd.n162 vdd.n161 9.3005
R5308 vdd.n134 vdd.n131 9.3005
R5309 vdd.n169 vdd.n168 9.3005
R5310 vdd.n104 vdd.n103 9.3005
R5311 vdd.n99 vdd.n98 9.3005
R5312 vdd.n110 vdd.n109 9.3005
R5313 vdd.n112 vdd.n111 9.3005
R5314 vdd.n95 vdd.n94 9.3005
R5315 vdd.n118 vdd.n117 9.3005
R5316 vdd.n120 vdd.n119 9.3005
R5317 vdd.n92 vdd.n89 9.3005
R5318 vdd.n127 vdd.n126 9.3005
R5319 vdd.n45 vdd.n44 9.3005
R5320 vdd.n40 vdd.n39 9.3005
R5321 vdd.n51 vdd.n50 9.3005
R5322 vdd.n53 vdd.n52 9.3005
R5323 vdd.n36 vdd.n35 9.3005
R5324 vdd.n59 vdd.n58 9.3005
R5325 vdd.n61 vdd.n60 9.3005
R5326 vdd.n33 vdd.n30 9.3005
R5327 vdd.n68 vdd.n67 9.3005
R5328 vdd.n3410 vdd.n3409 9.3005
R5329 vdd.n3413 vdd.n766 9.3005
R5330 vdd.n3414 vdd.n765 9.3005
R5331 vdd.n3417 vdd.n764 9.3005
R5332 vdd.n3418 vdd.n763 9.3005
R5333 vdd.n3421 vdd.n762 9.3005
R5334 vdd.n3422 vdd.n761 9.3005
R5335 vdd.n3425 vdd.n760 9.3005
R5336 vdd.n3426 vdd.n759 9.3005
R5337 vdd.n3429 vdd.n758 9.3005
R5338 vdd.n3430 vdd.n757 9.3005
R5339 vdd.n3433 vdd.n756 9.3005
R5340 vdd.n3434 vdd.n755 9.3005
R5341 vdd.n3437 vdd.n754 9.3005
R5342 vdd.n3438 vdd.n753 9.3005
R5343 vdd.n3441 vdd.n752 9.3005
R5344 vdd.n3442 vdd.n751 9.3005
R5345 vdd.n3445 vdd.n750 9.3005
R5346 vdd.n3446 vdd.n749 9.3005
R5347 vdd.n3449 vdd.n748 9.3005
R5348 vdd.n3453 vdd.n3452 9.3005
R5349 vdd.n3454 vdd.n747 9.3005
R5350 vdd.n3458 vdd.n3455 9.3005
R5351 vdd.n3461 vdd.n746 9.3005
R5352 vdd.n3462 vdd.n745 9.3005
R5353 vdd.n3465 vdd.n744 9.3005
R5354 vdd.n3466 vdd.n743 9.3005
R5355 vdd.n3469 vdd.n742 9.3005
R5356 vdd.n3470 vdd.n741 9.3005
R5357 vdd.n3473 vdd.n740 9.3005
R5358 vdd.n3474 vdd.n739 9.3005
R5359 vdd.n3477 vdd.n738 9.3005
R5360 vdd.n3478 vdd.n737 9.3005
R5361 vdd.n3481 vdd.n736 9.3005
R5362 vdd.n3482 vdd.n735 9.3005
R5363 vdd.n3485 vdd.n730 9.3005
R5364 vdd.n3491 vdd.n727 9.3005
R5365 vdd.n3492 vdd.n726 9.3005
R5366 vdd.n3506 vdd.n3505 9.3005
R5367 vdd.n3507 vdd.n681 9.3005
R5368 vdd.n3509 vdd.n3508 9.3005
R5369 vdd.n671 vdd.n670 9.3005
R5370 vdd.n3523 vdd.n3522 9.3005
R5371 vdd.n3524 vdd.n669 9.3005
R5372 vdd.n3526 vdd.n3525 9.3005
R5373 vdd.n660 vdd.n659 9.3005
R5374 vdd.n3539 vdd.n3538 9.3005
R5375 vdd.n3540 vdd.n658 9.3005
R5376 vdd.n3542 vdd.n3541 9.3005
R5377 vdd.n648 vdd.n647 9.3005
R5378 vdd.n3556 vdd.n3555 9.3005
R5379 vdd.n3557 vdd.n646 9.3005
R5380 vdd.n3559 vdd.n3558 9.3005
R5381 vdd.n637 vdd.n636 9.3005
R5382 vdd.n3575 vdd.n3574 9.3005
R5383 vdd.n3576 vdd.n635 9.3005
R5384 vdd.n3578 vdd.n3577 9.3005
R5385 vdd.n336 vdd.n334 9.3005
R5386 vdd.n683 vdd.n682 9.3005
R5387 vdd.n3670 vdd.n3669 9.3005
R5388 vdd.n337 vdd.n335 9.3005
R5389 vdd.n3663 vdd.n346 9.3005
R5390 vdd.n3662 vdd.n347 9.3005
R5391 vdd.n3661 vdd.n348 9.3005
R5392 vdd.n355 vdd.n349 9.3005
R5393 vdd.n3655 vdd.n356 9.3005
R5394 vdd.n3654 vdd.n357 9.3005
R5395 vdd.n3653 vdd.n358 9.3005
R5396 vdd.n366 vdd.n359 9.3005
R5397 vdd.n3647 vdd.n367 9.3005
R5398 vdd.n3646 vdd.n368 9.3005
R5399 vdd.n3645 vdd.n369 9.3005
R5400 vdd.n377 vdd.n370 9.3005
R5401 vdd.n3639 vdd.n378 9.3005
R5402 vdd.n3638 vdd.n379 9.3005
R5403 vdd.n3637 vdd.n380 9.3005
R5404 vdd.n388 vdd.n381 9.3005
R5405 vdd.n3631 vdd.n389 9.3005
R5406 vdd.n3630 vdd.n390 9.3005
R5407 vdd.n3629 vdd.n391 9.3005
R5408 vdd.n466 vdd.n463 9.3005
R5409 vdd.n470 vdd.n469 9.3005
R5410 vdd.n471 vdd.n462 9.3005
R5411 vdd.n475 vdd.n472 9.3005
R5412 vdd.n476 vdd.n461 9.3005
R5413 vdd.n480 vdd.n479 9.3005
R5414 vdd.n481 vdd.n460 9.3005
R5415 vdd.n485 vdd.n482 9.3005
R5416 vdd.n486 vdd.n459 9.3005
R5417 vdd.n490 vdd.n489 9.3005
R5418 vdd.n491 vdd.n458 9.3005
R5419 vdd.n495 vdd.n492 9.3005
R5420 vdd.n496 vdd.n457 9.3005
R5421 vdd.n500 vdd.n499 9.3005
R5422 vdd.n501 vdd.n456 9.3005
R5423 vdd.n505 vdd.n502 9.3005
R5424 vdd.n506 vdd.n455 9.3005
R5425 vdd.n510 vdd.n509 9.3005
R5426 vdd.n511 vdd.n454 9.3005
R5427 vdd.n515 vdd.n512 9.3005
R5428 vdd.n516 vdd.n451 9.3005
R5429 vdd.n520 vdd.n519 9.3005
R5430 vdd.n521 vdd.n450 9.3005
R5431 vdd.n525 vdd.n522 9.3005
R5432 vdd.n526 vdd.n449 9.3005
R5433 vdd.n530 vdd.n529 9.3005
R5434 vdd.n531 vdd.n448 9.3005
R5435 vdd.n535 vdd.n532 9.3005
R5436 vdd.n536 vdd.n447 9.3005
R5437 vdd.n540 vdd.n539 9.3005
R5438 vdd.n541 vdd.n446 9.3005
R5439 vdd.n545 vdd.n542 9.3005
R5440 vdd.n546 vdd.n445 9.3005
R5441 vdd.n550 vdd.n549 9.3005
R5442 vdd.n551 vdd.n444 9.3005
R5443 vdd.n555 vdd.n552 9.3005
R5444 vdd.n556 vdd.n443 9.3005
R5445 vdd.n560 vdd.n559 9.3005
R5446 vdd.n561 vdd.n442 9.3005
R5447 vdd.n565 vdd.n562 9.3005
R5448 vdd.n566 vdd.n439 9.3005
R5449 vdd.n570 vdd.n569 9.3005
R5450 vdd.n571 vdd.n438 9.3005
R5451 vdd.n575 vdd.n572 9.3005
R5452 vdd.n576 vdd.n437 9.3005
R5453 vdd.n580 vdd.n579 9.3005
R5454 vdd.n581 vdd.n436 9.3005
R5455 vdd.n585 vdd.n582 9.3005
R5456 vdd.n586 vdd.n435 9.3005
R5457 vdd.n590 vdd.n589 9.3005
R5458 vdd.n591 vdd.n434 9.3005
R5459 vdd.n595 vdd.n592 9.3005
R5460 vdd.n596 vdd.n433 9.3005
R5461 vdd.n600 vdd.n599 9.3005
R5462 vdd.n601 vdd.n432 9.3005
R5463 vdd.n605 vdd.n602 9.3005
R5464 vdd.n606 vdd.n431 9.3005
R5465 vdd.n610 vdd.n609 9.3005
R5466 vdd.n611 vdd.n430 9.3005
R5467 vdd.n615 vdd.n612 9.3005
R5468 vdd.n617 vdd.n429 9.3005
R5469 vdd.n619 vdd.n618 9.3005
R5470 vdd.n3623 vdd.n3622 9.3005
R5471 vdd.n465 vdd.n464 9.3005
R5472 vdd.n3501 vdd.n3500 9.3005
R5473 vdd.n676 vdd.n675 9.3005
R5474 vdd.n3514 vdd.n3513 9.3005
R5475 vdd.n3515 vdd.n674 9.3005
R5476 vdd.n3517 vdd.n3516 9.3005
R5477 vdd.n666 vdd.n665 9.3005
R5478 vdd.n3531 vdd.n3530 9.3005
R5479 vdd.n3532 vdd.n664 9.3005
R5480 vdd.n3534 vdd.n3533 9.3005
R5481 vdd.n653 vdd.n652 9.3005
R5482 vdd.n3547 vdd.n3546 9.3005
R5483 vdd.n3548 vdd.n651 9.3005
R5484 vdd.n3550 vdd.n3549 9.3005
R5485 vdd.n642 vdd.n641 9.3005
R5486 vdd.n3564 vdd.n3563 9.3005
R5487 vdd.n3565 vdd.n640 9.3005
R5488 vdd.n3570 vdd.n3566 9.3005
R5489 vdd.n3569 vdd.n3568 9.3005
R5490 vdd.n3567 vdd.n631 9.3005
R5491 vdd.n3583 vdd.n630 9.3005
R5492 vdd.n3585 vdd.n3584 9.3005
R5493 vdd.n3586 vdd.n629 9.3005
R5494 vdd.n3588 vdd.n3587 9.3005
R5495 vdd.n3590 vdd.n628 9.3005
R5496 vdd.n3592 vdd.n3591 9.3005
R5497 vdd.n3593 vdd.n627 9.3005
R5498 vdd.n3595 vdd.n3594 9.3005
R5499 vdd.n3597 vdd.n626 9.3005
R5500 vdd.n3599 vdd.n3598 9.3005
R5501 vdd.n3600 vdd.n625 9.3005
R5502 vdd.n3602 vdd.n3601 9.3005
R5503 vdd.n3605 vdd.n624 9.3005
R5504 vdd.n3607 vdd.n3606 9.3005
R5505 vdd.n3608 vdd.n623 9.3005
R5506 vdd.n3610 vdd.n3609 9.3005
R5507 vdd.n3612 vdd.n622 9.3005
R5508 vdd.n3614 vdd.n3613 9.3005
R5509 vdd.n3615 vdd.n621 9.3005
R5510 vdd.n3617 vdd.n3616 9.3005
R5511 vdd.n3619 vdd.n620 9.3005
R5512 vdd.n3621 vdd.n3620 9.3005
R5513 vdd.n3499 vdd.n686 9.3005
R5514 vdd.n3498 vdd.n3497 9.3005
R5515 vdd.n3367 vdd.n687 9.3005
R5516 vdd.n3376 vdd.n783 9.3005
R5517 vdd.n3379 vdd.n782 9.3005
R5518 vdd.n3380 vdd.n781 9.3005
R5519 vdd.n3383 vdd.n780 9.3005
R5520 vdd.n3384 vdd.n779 9.3005
R5521 vdd.n3387 vdd.n778 9.3005
R5522 vdd.n3388 vdd.n777 9.3005
R5523 vdd.n3391 vdd.n776 9.3005
R5524 vdd.n3392 vdd.n775 9.3005
R5525 vdd.n3395 vdd.n774 9.3005
R5526 vdd.n3396 vdd.n773 9.3005
R5527 vdd.n3399 vdd.n772 9.3005
R5528 vdd.n3400 vdd.n771 9.3005
R5529 vdd.n3403 vdd.n770 9.3005
R5530 vdd.n3407 vdd.n3406 9.3005
R5531 vdd.n3408 vdd.n767 9.3005
R5532 vdd.n2366 vdd.n2365 9.3005
R5533 vdd.n2361 vdd.n1517 9.3005
R5534 vdd.n1885 vdd.n1884 9.3005
R5535 vdd.n1886 vdd.n1640 9.3005
R5536 vdd.n1888 vdd.n1887 9.3005
R5537 vdd.n1630 vdd.n1629 9.3005
R5538 vdd.n1902 vdd.n1901 9.3005
R5539 vdd.n1903 vdd.n1628 9.3005
R5540 vdd.n1905 vdd.n1904 9.3005
R5541 vdd.n1620 vdd.n1619 9.3005
R5542 vdd.n1919 vdd.n1918 9.3005
R5543 vdd.n1920 vdd.n1618 9.3005
R5544 vdd.n1922 vdd.n1921 9.3005
R5545 vdd.n1607 vdd.n1606 9.3005
R5546 vdd.n1935 vdd.n1934 9.3005
R5547 vdd.n1936 vdd.n1605 9.3005
R5548 vdd.n1938 vdd.n1937 9.3005
R5549 vdd.n1596 vdd.n1595 9.3005
R5550 vdd.n1952 vdd.n1951 9.3005
R5551 vdd.n1953 vdd.n1594 9.3005
R5552 vdd.n1955 vdd.n1954 9.3005
R5553 vdd.n1585 vdd.n1584 9.3005
R5554 vdd.n2275 vdd.n2274 9.3005
R5555 vdd.n2276 vdd.n1583 9.3005
R5556 vdd.n2278 vdd.n2277 9.3005
R5557 vdd.n1573 vdd.n1572 9.3005
R5558 vdd.n2292 vdd.n2291 9.3005
R5559 vdd.n2293 vdd.n1571 9.3005
R5560 vdd.n2295 vdd.n2294 9.3005
R5561 vdd.n1563 vdd.n1562 9.3005
R5562 vdd.n2309 vdd.n2308 9.3005
R5563 vdd.n2310 vdd.n1561 9.3005
R5564 vdd.n2312 vdd.n2311 9.3005
R5565 vdd.n1550 vdd.n1549 9.3005
R5566 vdd.n2325 vdd.n2324 9.3005
R5567 vdd.n2326 vdd.n1548 9.3005
R5568 vdd.n2328 vdd.n2327 9.3005
R5569 vdd.n1540 vdd.n1539 9.3005
R5570 vdd.n2342 vdd.n2341 9.3005
R5571 vdd.n2343 vdd.n1537 9.3005
R5572 vdd.n2347 vdd.n2346 9.3005
R5573 vdd.n2345 vdd.n1538 9.3005
R5574 vdd.n2344 vdd.n1528 9.3005
R5575 vdd.n1642 vdd.n1641 9.3005
R5576 vdd.n1778 vdd.n1777 9.3005
R5577 vdd.n1779 vdd.n1768 9.3005
R5578 vdd.n1781 vdd.n1780 9.3005
R5579 vdd.n1782 vdd.n1767 9.3005
R5580 vdd.n1784 vdd.n1783 9.3005
R5581 vdd.n1785 vdd.n1762 9.3005
R5582 vdd.n1787 vdd.n1786 9.3005
R5583 vdd.n1788 vdd.n1761 9.3005
R5584 vdd.n1790 vdd.n1789 9.3005
R5585 vdd.n1791 vdd.n1756 9.3005
R5586 vdd.n1793 vdd.n1792 9.3005
R5587 vdd.n1794 vdd.n1755 9.3005
R5588 vdd.n1796 vdd.n1795 9.3005
R5589 vdd.n1797 vdd.n1750 9.3005
R5590 vdd.n1799 vdd.n1798 9.3005
R5591 vdd.n1800 vdd.n1749 9.3005
R5592 vdd.n1802 vdd.n1801 9.3005
R5593 vdd.n1803 vdd.n1744 9.3005
R5594 vdd.n1805 vdd.n1804 9.3005
R5595 vdd.n1806 vdd.n1743 9.3005
R5596 vdd.n1808 vdd.n1807 9.3005
R5597 vdd.n1812 vdd.n1739 9.3005
R5598 vdd.n1814 vdd.n1813 9.3005
R5599 vdd.n1815 vdd.n1738 9.3005
R5600 vdd.n1817 vdd.n1816 9.3005
R5601 vdd.n1818 vdd.n1733 9.3005
R5602 vdd.n1820 vdd.n1819 9.3005
R5603 vdd.n1821 vdd.n1732 9.3005
R5604 vdd.n1823 vdd.n1822 9.3005
R5605 vdd.n1824 vdd.n1727 9.3005
R5606 vdd.n1826 vdd.n1825 9.3005
R5607 vdd.n1827 vdd.n1726 9.3005
R5608 vdd.n1829 vdd.n1828 9.3005
R5609 vdd.n1830 vdd.n1721 9.3005
R5610 vdd.n1832 vdd.n1831 9.3005
R5611 vdd.n1833 vdd.n1720 9.3005
R5612 vdd.n1835 vdd.n1834 9.3005
R5613 vdd.n1836 vdd.n1715 9.3005
R5614 vdd.n1838 vdd.n1837 9.3005
R5615 vdd.n1839 vdd.n1714 9.3005
R5616 vdd.n1841 vdd.n1840 9.3005
R5617 vdd.n1842 vdd.n1709 9.3005
R5618 vdd.n1844 vdd.n1843 9.3005
R5619 vdd.n1845 vdd.n1708 9.3005
R5620 vdd.n1847 vdd.n1846 9.3005
R5621 vdd.n1848 vdd.n1701 9.3005
R5622 vdd.n1850 vdd.n1849 9.3005
R5623 vdd.n1851 vdd.n1700 9.3005
R5624 vdd.n1853 vdd.n1852 9.3005
R5625 vdd.n1854 vdd.n1695 9.3005
R5626 vdd.n1856 vdd.n1855 9.3005
R5627 vdd.n1857 vdd.n1694 9.3005
R5628 vdd.n1859 vdd.n1858 9.3005
R5629 vdd.n1860 vdd.n1689 9.3005
R5630 vdd.n1862 vdd.n1861 9.3005
R5631 vdd.n1863 vdd.n1688 9.3005
R5632 vdd.n1865 vdd.n1864 9.3005
R5633 vdd.n1866 vdd.n1683 9.3005
R5634 vdd.n1868 vdd.n1867 9.3005
R5635 vdd.n1869 vdd.n1682 9.3005
R5636 vdd.n1871 vdd.n1870 9.3005
R5637 vdd.n1647 vdd.n1646 9.3005
R5638 vdd.n1877 vdd.n1876 9.3005
R5639 vdd.n1776 vdd.n1775 9.3005
R5640 vdd.n1880 vdd.n1879 9.3005
R5641 vdd.n1636 vdd.n1635 9.3005
R5642 vdd.n1894 vdd.n1893 9.3005
R5643 vdd.n1895 vdd.n1634 9.3005
R5644 vdd.n1897 vdd.n1896 9.3005
R5645 vdd.n1625 vdd.n1624 9.3005
R5646 vdd.n1911 vdd.n1910 9.3005
R5647 vdd.n1912 vdd.n1623 9.3005
R5648 vdd.n1914 vdd.n1913 9.3005
R5649 vdd.n1614 vdd.n1613 9.3005
R5650 vdd.n1927 vdd.n1926 9.3005
R5651 vdd.n1928 vdd.n1612 9.3005
R5652 vdd.n1930 vdd.n1929 9.3005
R5653 vdd.n1602 vdd.n1601 9.3005
R5654 vdd.n1944 vdd.n1943 9.3005
R5655 vdd.n1945 vdd.n1600 9.3005
R5656 vdd.n1947 vdd.n1946 9.3005
R5657 vdd.n1591 vdd.n1590 9.3005
R5658 vdd.n1960 vdd.n1959 9.3005
R5659 vdd.n1961 vdd.n1589 9.3005
R5660 vdd.n1878 vdd.n1645 9.3005
R5661 vdd.n2181 vdd.n2180 9.3005
R5662 vdd.n2176 vdd.n2175 9.3005
R5663 vdd.n2187 vdd.n2186 9.3005
R5664 vdd.n2189 vdd.n2188 9.3005
R5665 vdd.n2172 vdd.n2171 9.3005
R5666 vdd.n2195 vdd.n2194 9.3005
R5667 vdd.n2197 vdd.n2196 9.3005
R5668 vdd.n2169 vdd.n2166 9.3005
R5669 vdd.n2204 vdd.n2203 9.3005
R5670 vdd.n2240 vdd.n2239 9.3005
R5671 vdd.n2235 vdd.n2234 9.3005
R5672 vdd.n2246 vdd.n2245 9.3005
R5673 vdd.n2248 vdd.n2247 9.3005
R5674 vdd.n2231 vdd.n2230 9.3005
R5675 vdd.n2254 vdd.n2253 9.3005
R5676 vdd.n2256 vdd.n2255 9.3005
R5677 vdd.n2228 vdd.n2225 9.3005
R5678 vdd.n2263 vdd.n2262 9.3005
R5679 vdd.n2079 vdd.n2078 9.3005
R5680 vdd.n2074 vdd.n2073 9.3005
R5681 vdd.n2085 vdd.n2084 9.3005
R5682 vdd.n2087 vdd.n2086 9.3005
R5683 vdd.n2070 vdd.n2069 9.3005
R5684 vdd.n2093 vdd.n2092 9.3005
R5685 vdd.n2095 vdd.n2094 9.3005
R5686 vdd.n2067 vdd.n2064 9.3005
R5687 vdd.n2102 vdd.n2101 9.3005
R5688 vdd.n2138 vdd.n2137 9.3005
R5689 vdd.n2133 vdd.n2132 9.3005
R5690 vdd.n2144 vdd.n2143 9.3005
R5691 vdd.n2146 vdd.n2145 9.3005
R5692 vdd.n2129 vdd.n2128 9.3005
R5693 vdd.n2152 vdd.n2151 9.3005
R5694 vdd.n2154 vdd.n2153 9.3005
R5695 vdd.n2126 vdd.n2123 9.3005
R5696 vdd.n2161 vdd.n2160 9.3005
R5697 vdd.n1978 vdd.n1977 9.3005
R5698 vdd.n1973 vdd.n1972 9.3005
R5699 vdd.n1984 vdd.n1983 9.3005
R5700 vdd.n1986 vdd.n1985 9.3005
R5701 vdd.n1969 vdd.n1968 9.3005
R5702 vdd.n1992 vdd.n1991 9.3005
R5703 vdd.n1994 vdd.n1993 9.3005
R5704 vdd.n1966 vdd.n1963 9.3005
R5705 vdd.n2001 vdd.n2000 9.3005
R5706 vdd.n2037 vdd.n2036 9.3005
R5707 vdd.n2032 vdd.n2031 9.3005
R5708 vdd.n2043 vdd.n2042 9.3005
R5709 vdd.n2045 vdd.n2044 9.3005
R5710 vdd.n2028 vdd.n2027 9.3005
R5711 vdd.n2051 vdd.n2050 9.3005
R5712 vdd.n2053 vdd.n2052 9.3005
R5713 vdd.n2025 vdd.n2022 9.3005
R5714 vdd.n2060 vdd.n2059 9.3005
R5715 vdd.n1916 vdd.t123 9.18308
R5716 vdd.n3603 vdd.t61 9.18308
R5717 vdd.n1610 vdd.t109 8.95635
R5718 vdd.n2358 vdd.t156 8.95635
R5719 vdd.n723 vdd.t173 8.95635
R5720 vdd.t43 vdd.n3657 8.95635
R5721 vdd.n312 vdd.n311 8.92171
R5722 vdd.n253 vdd.n252 8.92171
R5723 vdd.n210 vdd.n209 8.92171
R5724 vdd.n151 vdd.n150 8.92171
R5725 vdd.n109 vdd.n108 8.92171
R5726 vdd.n50 vdd.n49 8.92171
R5727 vdd.n2186 vdd.n2185 8.92171
R5728 vdd.n2245 vdd.n2244 8.92171
R5729 vdd.n2084 vdd.n2083 8.92171
R5730 vdd.n2143 vdd.n2142 8.92171
R5731 vdd.n1983 vdd.n1982 8.92171
R5732 vdd.n2042 vdd.n2041 8.92171
R5733 vdd.n231 vdd.n129 8.81535
R5734 vdd.n2164 vdd.n2062 8.81535
R5735 vdd.n1957 vdd.t7 8.72962
R5736 vdd.t46 vdd.n3666 8.72962
R5737 vdd.n2280 vdd.t87 8.50289
R5738 vdd.n3572 vdd.t279 8.50289
R5739 vdd.n28 vdd.n14 8.42249
R5740 vdd.n2306 vdd.t68 8.27616
R5741 vdd.t17 vdd.n656 8.27616
R5742 vdd.n3672 vdd.n3671 8.16225
R5743 vdd.n2268 vdd.n2267 8.16225
R5744 vdd.n308 vdd.n302 8.14595
R5745 vdd.n249 vdd.n243 8.14595
R5746 vdd.n206 vdd.n200 8.14595
R5747 vdd.n147 vdd.n141 8.14595
R5748 vdd.n105 vdd.n99 8.14595
R5749 vdd.n46 vdd.n40 8.14595
R5750 vdd.n2182 vdd.n2176 8.14595
R5751 vdd.n2241 vdd.n2235 8.14595
R5752 vdd.n2080 vdd.n2074 8.14595
R5753 vdd.n2139 vdd.n2133 8.14595
R5754 vdd.n1979 vdd.n1973 8.14595
R5755 vdd.n2038 vdd.n2032 8.14595
R5756 vdd.n1553 vdd.t64 8.04943
R5757 vdd.n3528 vdd.t20 8.04943
R5758 vdd.n2513 vdd.n1134 7.70933
R5759 vdd.n2513 vdd.n1137 7.70933
R5760 vdd.n2519 vdd.n1123 7.70933
R5761 vdd.n2525 vdd.n1123 7.70933
R5762 vdd.n2525 vdd.n1116 7.70933
R5763 vdd.n2531 vdd.n1116 7.70933
R5764 vdd.n2531 vdd.n1119 7.70933
R5765 vdd.n2537 vdd.n1112 7.70933
R5766 vdd.n2543 vdd.n1106 7.70933
R5767 vdd.n2549 vdd.n1093 7.70933
R5768 vdd.n2555 vdd.n1093 7.70933
R5769 vdd.n2561 vdd.n1087 7.70933
R5770 vdd.n2567 vdd.n1080 7.70933
R5771 vdd.n2567 vdd.n1083 7.70933
R5772 vdd.n2573 vdd.n1076 7.70933
R5773 vdd.n2580 vdd.n1062 7.70933
R5774 vdd.n2586 vdd.n1062 7.70933
R5775 vdd.n2592 vdd.n1056 7.70933
R5776 vdd.n2598 vdd.n1052 7.70933
R5777 vdd.n2604 vdd.n1046 7.70933
R5778 vdd.n2622 vdd.n1028 7.70933
R5779 vdd.n2622 vdd.n1021 7.70933
R5780 vdd.n2630 vdd.n1021 7.70933
R5781 vdd.n2712 vdd.n1005 7.70933
R5782 vdd.n3095 vdd.n957 7.70933
R5783 vdd.n3107 vdd.n946 7.70933
R5784 vdd.n3107 vdd.n940 7.70933
R5785 vdd.n3113 vdd.n940 7.70933
R5786 vdd.n3125 vdd.n931 7.70933
R5787 vdd.n3131 vdd.n925 7.70933
R5788 vdd.n3143 vdd.n912 7.70933
R5789 vdd.n3150 vdd.n905 7.70933
R5790 vdd.n3150 vdd.n908 7.70933
R5791 vdd.n3156 vdd.n901 7.70933
R5792 vdd.n3162 vdd.n887 7.70933
R5793 vdd.n3168 vdd.n887 7.70933
R5794 vdd.n3174 vdd.n881 7.70933
R5795 vdd.n3180 vdd.n874 7.70933
R5796 vdd.n3180 vdd.n877 7.70933
R5797 vdd.n3186 vdd.n870 7.70933
R5798 vdd.n3192 vdd.n864 7.70933
R5799 vdd.n3198 vdd.n851 7.70933
R5800 vdd.n3204 vdd.n851 7.70933
R5801 vdd.n3204 vdd.n843 7.70933
R5802 vdd.n3255 vdd.n843 7.70933
R5803 vdd.n3255 vdd.n846 7.70933
R5804 vdd.n3261 vdd.n805 7.70933
R5805 vdd.n3331 vdd.n805 7.70933
R5806 vdd.n307 vdd.n304 7.3702
R5807 vdd.n248 vdd.n245 7.3702
R5808 vdd.n205 vdd.n202 7.3702
R5809 vdd.n146 vdd.n143 7.3702
R5810 vdd.n104 vdd.n101 7.3702
R5811 vdd.n45 vdd.n42 7.3702
R5812 vdd.n2181 vdd.n2178 7.3702
R5813 vdd.n2240 vdd.n2237 7.3702
R5814 vdd.n2079 vdd.n2076 7.3702
R5815 vdd.n2138 vdd.n2135 7.3702
R5816 vdd.n1978 vdd.n1975 7.3702
R5817 vdd.n2037 vdd.n2034 7.3702
R5818 vdd.n1106 vdd.t276 7.36923
R5819 vdd.n3186 vdd.t253 7.36923
R5820 vdd.n2339 vdd.t11 7.1425
R5821 vdd.n2537 vdd.t228 7.1425
R5822 vdd.n1425 vdd.t224 7.1425
R5823 vdd.n3119 vdd.t227 7.1425
R5824 vdd.n864 vdd.t237 7.1425
R5825 vdd.n679 vdd.t37 7.1425
R5826 vdd.n1813 vdd.n1812 6.98232
R5827 vdd.n2401 vdd.n2400 6.98232
R5828 vdd.n566 vdd.n565 6.98232
R5829 vdd.n3413 vdd.n3410 6.98232
R5830 vdd.t85 vdd.n1552 6.91577
R5831 vdd.n3536 vdd.t2 6.91577
R5832 vdd.n1425 vdd.t225 6.80241
R5833 vdd.n3119 vdd.t269 6.80241
R5834 vdd.n2298 vdd.t135 6.68904
R5835 vdd.n3552 vdd.t39 6.68904
R5836 vdd.t89 vdd.n1581 6.46231
R5837 vdd.n2561 vdd.t235 6.46231
R5838 vdd.t240 vdd.n1056 6.46231
R5839 vdd.n3143 vdd.t245 6.46231
R5840 vdd.t261 vdd.n881 6.46231
R5841 vdd.n3580 vdd.t72 6.46231
R5842 vdd.n3672 vdd.n333 6.38151
R5843 vdd.n2267 vdd.n2266 6.38151
R5844 vdd.n2637 vdd.t273 6.34895
R5845 vdd.n3016 vdd.t258 6.34895
R5846 vdd.n3158 vdd.n897 6.2444
R5847 vdd.n2577 vdd.n2576 6.2444
R5848 vdd.n1949 vdd.t41 6.23558
R5849 vdd.t13 vdd.n344 6.23558
R5850 vdd.t24 vdd.n1609 6.00885
R5851 vdd.n3651 vdd.t31 6.00885
R5852 vdd.n2598 vdd.t266 5.89549
R5853 vdd.n925 vdd.t241 5.89549
R5854 vdd.n308 vdd.n307 5.81868
R5855 vdd.n249 vdd.n248 5.81868
R5856 vdd.n206 vdd.n205 5.81868
R5857 vdd.n147 vdd.n146 5.81868
R5858 vdd.n105 vdd.n104 5.81868
R5859 vdd.n46 vdd.n45 5.81868
R5860 vdd.n2182 vdd.n2181 5.81868
R5861 vdd.n2241 vdd.n2240 5.81868
R5862 vdd.n2080 vdd.n2079 5.81868
R5863 vdd.n2139 vdd.n2138 5.81868
R5864 vdd.n1979 vdd.n1978 5.81868
R5865 vdd.n2038 vdd.n2037 5.81868
R5866 vdd.n1908 vdd.t9 5.78212
R5867 vdd.n3642 vdd.t117 5.78212
R5868 vdd.n2720 vdd.n2719 5.77611
R5869 vdd.n1349 vdd.n1348 5.77611
R5870 vdd.n3028 vdd.n3027 5.77611
R5871 vdd.n3272 vdd.n3271 5.77611
R5872 vdd.n3336 vdd.n801 5.77611
R5873 vdd.n2891 vdd.n2825 5.77611
R5874 vdd.n2645 vdd.n1012 5.77611
R5875 vdd.n1485 vdd.n1317 5.77611
R5876 vdd.n1775 vdd.n1774 5.62474
R5877 vdd.n2364 vdd.n2361 5.62474
R5878 vdd.n3623 vdd.n428 5.62474
R5879 vdd.n3497 vdd.n690 5.62474
R5880 vdd.n1632 vdd.t9 5.55539
R5881 vdd.n2573 vdd.t255 5.55539
R5882 vdd.n901 vdd.t231 5.55539
R5883 vdd.t117 vdd.n3641 5.55539
R5884 vdd.n1924 vdd.t24 5.32866
R5885 vdd.t31 vdd.n3650 5.32866
R5886 vdd.n1940 vdd.t41 5.10193
R5887 vdd.n3659 vdd.t13 5.10193
R5888 vdd.n311 vdd.n302 5.04292
R5889 vdd.n252 vdd.n243 5.04292
R5890 vdd.n209 vdd.n200 5.04292
R5891 vdd.n150 vdd.n141 5.04292
R5892 vdd.n108 vdd.n99 5.04292
R5893 vdd.n49 vdd.n40 5.04292
R5894 vdd.n2185 vdd.n2176 5.04292
R5895 vdd.n2244 vdd.n2235 5.04292
R5896 vdd.n2083 vdd.n2074 5.04292
R5897 vdd.n2142 vdd.n2133 5.04292
R5898 vdd.n1982 vdd.n1973 5.04292
R5899 vdd.n2041 vdd.n2032 5.04292
R5900 vdd.n2272 vdd.t89 4.8752
R5901 vdd.t234 vdd.t246 4.8752
R5902 vdd.t277 vdd.t223 4.8752
R5903 vdd.t72 vdd.n340 4.8752
R5904 vdd.n2721 vdd.n2720 4.83952
R5905 vdd.n1348 vdd.n1347 4.83952
R5906 vdd.n3029 vdd.n3028 4.83952
R5907 vdd.n3273 vdd.n3272 4.83952
R5908 vdd.n801 vdd.n796 4.83952
R5909 vdd.n2888 vdd.n2825 4.83952
R5910 vdd.n2648 vdd.n1012 4.83952
R5911 vdd.n1488 vdd.n1317 4.83952
R5912 vdd.n1399 vdd.t243 4.76184
R5913 vdd.n3101 vdd.t229 4.76184
R5914 vdd.n2369 vdd.n2368 4.74817
R5915 vdd.n1521 vdd.n1516 4.74817
R5916 vdd.n1183 vdd.n1180 4.74817
R5917 vdd.n2462 vdd.n1179 4.74817
R5918 vdd.n2467 vdd.n1180 4.74817
R5919 vdd.n2466 vdd.n1179 4.74817
R5920 vdd.n3490 vdd.n3489 4.74817
R5921 vdd.n3487 vdd.n3486 4.74817
R5922 vdd.n3487 vdd.n732 4.74817
R5923 vdd.n3489 vdd.n729 4.74817
R5924 vdd.n3372 vdd.n784 4.74817
R5925 vdd.n3368 vdd.n3366 4.74817
R5926 vdd.n3371 vdd.n3366 4.74817
R5927 vdd.n3375 vdd.n784 4.74817
R5928 vdd.n2368 vdd.n1279 4.74817
R5929 vdd.n1518 vdd.n1516 4.74817
R5930 vdd.n333 vdd.n332 4.7074
R5931 vdd.n231 vdd.n230 4.7074
R5932 vdd.n2266 vdd.n2265 4.7074
R5933 vdd.n2164 vdd.n2163 4.7074
R5934 vdd.n1575 vdd.t135 4.64847
R5935 vdd.t236 vdd.n1087 4.64847
R5936 vdd.n2592 vdd.t275 4.64847
R5937 vdd.t264 vdd.n912 4.64847
R5938 vdd.n3174 vdd.t260 4.64847
R5939 vdd.n3561 vdd.t39 4.64847
R5940 vdd.n1076 vdd.t204 4.53511
R5941 vdd.n3156 vdd.t177 4.53511
R5942 vdd.n2314 vdd.t85 4.42174
R5943 vdd.n2519 vdd.t152 4.42174
R5944 vdd.n1399 vdd.t193 4.42174
R5945 vdd.n3101 vdd.t200 4.42174
R5946 vdd.n846 vdd.t148 4.42174
R5947 vdd.t2 vdd.n655 4.42174
R5948 vdd.n3147 vdd.n897 4.37123
R5949 vdd.n2578 vdd.n2577 4.37123
R5950 vdd.n2616 vdd.t262 4.30838
R5951 vdd.n3004 vdd.t249 4.30838
R5952 vdd.n312 vdd.n300 4.26717
R5953 vdd.n253 vdd.n241 4.26717
R5954 vdd.n210 vdd.n198 4.26717
R5955 vdd.n151 vdd.n139 4.26717
R5956 vdd.n109 vdd.n97 4.26717
R5957 vdd.n50 vdd.n38 4.26717
R5958 vdd.n2186 vdd.n2174 4.26717
R5959 vdd.n2245 vdd.n2233 4.26717
R5960 vdd.n2084 vdd.n2072 4.26717
R5961 vdd.n2143 vdd.n2131 4.26717
R5962 vdd.n1983 vdd.n1971 4.26717
R5963 vdd.n2042 vdd.n2030 4.26717
R5964 vdd.n2330 vdd.t11 4.19501
R5965 vdd.n3520 vdd.t37 4.19501
R5966 vdd.n333 vdd.n231 4.10845
R5967 vdd.n2266 vdd.n2164 4.10845
R5968 vdd.n289 vdd.t19 4.06363
R5969 vdd.n289 vdd.t299 4.06363
R5970 vdd.n287 vdd.t51 4.06363
R5971 vdd.n287 vdd.t140 4.06363
R5972 vdd.n285 vdd.t44 4.06363
R5973 vdd.n285 vdd.t92 4.06363
R5974 vdd.n283 vdd.t102 4.06363
R5975 vdd.n283 vdd.t133 4.06363
R5976 vdd.n281 vdd.t142 4.06363
R5977 vdd.n281 vdd.t47 4.06363
R5978 vdd.n279 vdd.t280 4.06363
R5979 vdd.n279 vdd.t134 4.06363
R5980 vdd.n277 vdd.t288 4.06363
R5981 vdd.n277 vdd.t55 4.06363
R5982 vdd.n275 vdd.t3 4.06363
R5983 vdd.n275 vdd.t18 4.06363
R5984 vdd.n273 vdd.t81 4.06363
R5985 vdd.n273 vdd.t63 4.06363
R5986 vdd.n187 vdd.t1 4.06363
R5987 vdd.n187 vdd.t138 4.06363
R5988 vdd.n185 vdd.t32 4.06363
R5989 vdd.n185 vdd.t62 4.06363
R5990 vdd.n183 vdd.t76 4.06363
R5991 vdd.n183 vdd.t146 4.06363
R5992 vdd.n181 vdd.t297 4.06363
R5993 vdd.n181 vdd.t22 4.06363
R5994 vdd.n179 vdd.t73 4.06363
R5995 vdd.n179 vdd.t111 4.06363
R5996 vdd.n177 vdd.t307 4.06363
R5997 vdd.n177 vdd.t283 4.06363
R5998 vdd.n175 vdd.t104 4.06363
R5999 vdd.n175 vdd.t40 4.06363
R6000 vdd.n173 vdd.t294 4.06363
R6001 vdd.n173 vdd.t122 4.06363
R6002 vdd.n171 vdd.t114 4.06363
R6003 vdd.n171 vdd.t30 4.06363
R6004 vdd.n86 vdd.t131 4.06363
R6005 vdd.n86 vdd.t118 4.06363
R6006 vdd.n84 vdd.t75 4.06363
R6007 vdd.n84 vdd.t126 4.06363
R6008 vdd.n82 vdd.t141 4.06363
R6009 vdd.n82 vdd.t80 4.06363
R6010 vdd.n80 vdd.t34 4.06363
R6011 vdd.n80 vdd.t14 4.06363
R6012 vdd.n78 vdd.t91 4.06363
R6013 vdd.n78 vdd.t306 4.06363
R6014 vdd.n76 vdd.t290 4.06363
R6015 vdd.n76 vdd.t120 4.06363
R6016 vdd.n74 vdd.t289 4.06363
R6017 vdd.n74 vdd.t45 4.06363
R6018 vdd.n72 vdd.t6 4.06363
R6019 vdd.n72 vdd.t78 4.06363
R6020 vdd.n70 vdd.t21 4.06363
R6021 vdd.n70 vdd.t121 4.06363
R6022 vdd.n2206 vdd.t23 4.06363
R6023 vdd.n2206 vdd.t65 4.06363
R6024 vdd.n2208 vdd.t105 4.06363
R6025 vdd.n2208 vdd.t86 4.06363
R6026 vdd.n2210 vdd.t284 4.06363
R6027 vdd.n2210 vdd.t59 4.06363
R6028 vdd.n2212 vdd.t108 4.06363
R6029 vdd.n2212 vdd.t88 4.06363
R6030 vdd.n2214 vdd.t8 4.06363
R6031 vdd.n2214 vdd.t115 4.06363
R6032 vdd.n2216 vdd.t143 4.06363
R6033 vdd.n2216 vdd.t132 4.06363
R6034 vdd.n2218 vdd.t291 4.06363
R6035 vdd.n2218 vdd.t302 4.06363
R6036 vdd.n2220 vdd.t282 4.06363
R6037 vdd.n2220 vdd.t25 4.06363
R6038 vdd.n2222 vdd.t60 4.06363
R6039 vdd.n2222 vdd.t107 4.06363
R6040 vdd.n2104 vdd.t293 4.06363
R6041 vdd.n2104 vdd.t301 4.06363
R6042 vdd.n2106 vdd.t69 4.06363
R6043 vdd.n2106 vdd.t128 4.06363
R6044 vdd.n2108 vdd.t136 4.06363
R6045 vdd.n2108 vdd.t287 4.06363
R6046 vdd.n2110 vdd.t305 4.06363
R6047 vdd.n2110 vdd.t129 4.06363
R6048 vdd.n2112 vdd.t127 4.06363
R6049 vdd.n2112 vdd.t112 4.06363
R6050 vdd.n2114 vdd.t42 4.06363
R6051 vdd.n2114 vdd.t74 4.06363
R6052 vdd.n2116 vdd.t57 4.06363
R6053 vdd.n2116 vdd.t113 4.06363
R6054 vdd.n2118 vdd.t124 4.06363
R6055 vdd.n2118 vdd.t300 4.06363
R6056 vdd.n2120 vdd.t10 4.06363
R6057 vdd.n2120 vdd.t298 4.06363
R6058 vdd.n2003 vdd.t16 4.06363
R6059 vdd.n2003 vdd.t296 4.06363
R6060 vdd.n2005 vdd.t77 4.06363
R6061 vdd.n2005 vdd.t285 4.06363
R6062 vdd.n2007 vdd.t292 4.06363
R6063 vdd.n2007 vdd.t53 4.06363
R6064 vdd.n2009 vdd.t50 4.06363
R6065 vdd.n2009 vdd.t130 4.06363
R6066 vdd.n2011 vdd.t295 4.06363
R6067 vdd.n2011 vdd.t90 4.06363
R6068 vdd.n2013 vdd.t125 4.06363
R6069 vdd.n2013 vdd.t36 4.06363
R6070 vdd.n2015 vdd.t303 4.06363
R6071 vdd.n2015 vdd.t110 4.06363
R6072 vdd.n2017 vdd.t281 4.06363
R6073 vdd.n2017 vdd.t54 4.06363
R6074 vdd.n2019 vdd.t48 4.06363
R6075 vdd.n2019 vdd.t139 4.06363
R6076 vdd.n1112 vdd.t268 3.96828
R6077 vdd.n2610 vdd.t248 3.96828
R6078 vdd.n2998 vdd.t265 3.96828
R6079 vdd.n3192 vdd.t254 3.96828
R6080 vdd.n26 vdd.t82 3.9605
R6081 vdd.n26 vdd.t97 3.9605
R6082 vdd.n23 vdd.t84 3.9605
R6083 vdd.n23 vdd.t28 3.9605
R6084 vdd.n21 vdd.t27 3.9605
R6085 vdd.n21 vdd.t100 3.9605
R6086 vdd.n20 vdd.t4 3.9605
R6087 vdd.n20 vdd.t96 3.9605
R6088 vdd.n15 vdd.t26 3.9605
R6089 vdd.n15 vdd.t99 3.9605
R6090 vdd.n16 vdd.t98 3.9605
R6091 vdd.n16 vdd.t95 3.9605
R6092 vdd.n18 vdd.t101 3.9605
R6093 vdd.n18 vdd.t83 3.9605
R6094 vdd.n25 vdd.t94 3.9605
R6095 vdd.n25 vdd.t5 3.9605
R6096 vdd.n2543 vdd.t268 3.74155
R6097 vdd.n1046 vdd.t248 3.74155
R6098 vdd.n3125 vdd.t265 3.74155
R6099 vdd.n870 vdd.t254 3.74155
R6100 vdd.n7 vdd.t278 3.61217
R6101 vdd.n7 vdd.t242 3.61217
R6102 vdd.n8 vdd.t250 3.61217
R6103 vdd.n8 vdd.t270 3.61217
R6104 vdd.n10 vdd.t259 3.61217
R6105 vdd.n10 vdd.t230 3.61217
R6106 vdd.n12 vdd.t239 3.61217
R6107 vdd.n12 vdd.t257 3.61217
R6108 vdd.n5 vdd.t272 3.61217
R6109 vdd.n5 vdd.t252 3.61217
R6110 vdd.n3 vdd.t244 3.61217
R6111 vdd.n3 vdd.t274 3.61217
R6112 vdd.n1 vdd.t226 3.61217
R6113 vdd.n1 vdd.t263 3.61217
R6114 vdd.n0 vdd.t267 3.61217
R6115 vdd.n0 vdd.t247 3.61217
R6116 vdd.n316 vdd.n315 3.49141
R6117 vdd.n257 vdd.n256 3.49141
R6118 vdd.n214 vdd.n213 3.49141
R6119 vdd.n155 vdd.n154 3.49141
R6120 vdd.n113 vdd.n112 3.49141
R6121 vdd.n54 vdd.n53 3.49141
R6122 vdd.n2190 vdd.n2189 3.49141
R6123 vdd.n2249 vdd.n2248 3.49141
R6124 vdd.n2088 vdd.n2087 3.49141
R6125 vdd.n2147 vdd.n2146 3.49141
R6126 vdd.n1987 vdd.n1986 3.49141
R6127 vdd.n2046 vdd.n2045 3.49141
R6128 vdd.t262 vdd.n1028 3.40145
R6129 vdd.n2784 vdd.t271 3.40145
R6130 vdd.n3088 vdd.t256 3.40145
R6131 vdd.n3113 vdd.t249 3.40145
R6132 vdd.n2331 vdd.t64 3.28809
R6133 vdd.n1137 vdd.t152 3.28809
R6134 vdd.n2637 vdd.t193 3.28809
R6135 vdd.n3016 vdd.t200 3.28809
R6136 vdd.n3261 vdd.t148 3.28809
R6137 vdd.n3519 vdd.t20 3.28809
R6138 vdd.t68 vdd.n1559 3.06136
R6139 vdd.n2555 vdd.t236 3.06136
R6140 vdd.n1437 vdd.t275 3.06136
R6141 vdd.n3137 vdd.t264 3.06136
R6142 vdd.t260 vdd.n874 3.06136
R6143 vdd.n3544 vdd.t17 3.06136
R6144 vdd.n2630 vdd.t243 2.94799
R6145 vdd.t229 vdd.n946 2.94799
R6146 vdd.n2289 vdd.t87 2.83463
R6147 vdd.n644 vdd.t279 2.83463
R6148 vdd.n319 vdd.n298 2.71565
R6149 vdd.n260 vdd.n239 2.71565
R6150 vdd.n217 vdd.n196 2.71565
R6151 vdd.n158 vdd.n137 2.71565
R6152 vdd.n116 vdd.n95 2.71565
R6153 vdd.n57 vdd.n36 2.71565
R6154 vdd.n2193 vdd.n2172 2.71565
R6155 vdd.n2252 vdd.n2231 2.71565
R6156 vdd.n2091 vdd.n2070 2.71565
R6157 vdd.n2150 vdd.n2129 2.71565
R6158 vdd.n1990 vdd.n1969 2.71565
R6159 vdd.n2049 vdd.n2028 2.71565
R6160 vdd.t7 vdd.n1587 2.6079
R6161 vdd.n3667 vdd.t46 2.6079
R6162 vdd.n2604 vdd.t246 2.49453
R6163 vdd.n931 vdd.t277 2.49453
R6164 vdd.n306 vdd.n305 2.4129
R6165 vdd.n247 vdd.n246 2.4129
R6166 vdd.n204 vdd.n203 2.4129
R6167 vdd.n145 vdd.n144 2.4129
R6168 vdd.n103 vdd.n102 2.4129
R6169 vdd.n44 vdd.n43 2.4129
R6170 vdd.n2180 vdd.n2179 2.4129
R6171 vdd.n2239 vdd.n2238 2.4129
R6172 vdd.n2078 vdd.n2077 2.4129
R6173 vdd.n2137 vdd.n2136 2.4129
R6174 vdd.n1977 vdd.n1976 2.4129
R6175 vdd.n2036 vdd.n2035 2.4129
R6176 vdd.n1941 vdd.t109 2.38117
R6177 vdd.n2349 vdd.t156 2.38117
R6178 vdd.n3503 vdd.t173 2.38117
R6179 vdd.n3658 vdd.t43 2.38117
R6180 vdd.n2474 vdd.n1180 2.27742
R6181 vdd.n2474 vdd.n1179 2.27742
R6182 vdd.n3488 vdd.n3487 2.27742
R6183 vdd.n3489 vdd.n3488 2.27742
R6184 vdd.n3366 vdd.n3365 2.27742
R6185 vdd.n3365 vdd.n784 2.27742
R6186 vdd.n2368 vdd.n2367 2.27742
R6187 vdd.n2367 vdd.n1516 2.27742
R6188 vdd.t123 vdd.n1616 2.15444
R6189 vdd.n1083 vdd.t255 2.15444
R6190 vdd.n2580 vdd.t233 2.15444
R6191 vdd.n908 vdd.t232 2.15444
R6192 vdd.n3162 vdd.t231 2.15444
R6193 vdd.n3649 vdd.t61 2.15444
R6194 vdd.n320 vdd.n296 1.93989
R6195 vdd.n261 vdd.n237 1.93989
R6196 vdd.n218 vdd.n194 1.93989
R6197 vdd.n159 vdd.n135 1.93989
R6198 vdd.n117 vdd.n93 1.93989
R6199 vdd.n58 vdd.n34 1.93989
R6200 vdd.n2194 vdd.n2170 1.93989
R6201 vdd.n2253 vdd.n2229 1.93989
R6202 vdd.n2092 vdd.n2068 1.93989
R6203 vdd.n2151 vdd.n2127 1.93989
R6204 vdd.n1991 vdd.n1967 1.93989
R6205 vdd.n2050 vdd.n2026 1.93989
R6206 vdd.n1899 vdd.t66 1.92771
R6207 vdd.t70 vdd.n375 1.92771
R6208 vdd.n1437 vdd.t266 1.81434
R6209 vdd.n3137 vdd.t241 1.81434
R6210 vdd.n1907 vdd.t106 1.70098
R6211 vdd.n3643 vdd.t0 1.70098
R6212 vdd.n1932 vdd.t56 1.47425
R6213 vdd.n361 vdd.t79 1.47425
R6214 vdd.t273 vdd.n1005 1.36088
R6215 vdd.n3095 vdd.t258 1.36088
R6216 vdd.n1598 vdd.t35 1.24752
R6217 vdd.t235 vdd.n1080 1.24752
R6218 vdd.n2586 vdd.t240 1.24752
R6219 vdd.t245 vdd.n905 1.24752
R6220 vdd.n3168 vdd.t261 1.24752
R6221 vdd.t33 vdd.n3665 1.24752
R6222 vdd.n2267 vdd.n28 1.21639
R6223 vdd vdd.n3672 1.20856
R6224 vdd.n331 vdd.n291 1.16414
R6225 vdd.n324 vdd.n323 1.16414
R6226 vdd.n272 vdd.n232 1.16414
R6227 vdd.n265 vdd.n264 1.16414
R6228 vdd.n229 vdd.n189 1.16414
R6229 vdd.n222 vdd.n221 1.16414
R6230 vdd.n170 vdd.n130 1.16414
R6231 vdd.n163 vdd.n162 1.16414
R6232 vdd.n128 vdd.n88 1.16414
R6233 vdd.n121 vdd.n120 1.16414
R6234 vdd.n69 vdd.n29 1.16414
R6235 vdd.n62 vdd.n61 1.16414
R6236 vdd.n2205 vdd.n2165 1.16414
R6237 vdd.n2198 vdd.n2197 1.16414
R6238 vdd.n2264 vdd.n2224 1.16414
R6239 vdd.n2257 vdd.n2256 1.16414
R6240 vdd.n2103 vdd.n2063 1.16414
R6241 vdd.n2096 vdd.n2095 1.16414
R6242 vdd.n2162 vdd.n2122 1.16414
R6243 vdd.n2155 vdd.n2154 1.16414
R6244 vdd.n2002 vdd.n1962 1.16414
R6245 vdd.n1995 vdd.n1994 1.16414
R6246 vdd.n2061 vdd.n2021 1.16414
R6247 vdd.n2054 vdd.n2053 1.16414
R6248 vdd.n2281 vdd.t49 1.02079
R6249 vdd.t204 vdd.t233 1.02079
R6250 vdd.t232 vdd.t177 1.02079
R6251 vdd.t119 vdd.n633 1.02079
R6252 vdd.n1778 vdd.n1774 0.970197
R6253 vdd.n2365 vdd.n2364 0.970197
R6254 vdd.n618 vdd.n428 0.970197
R6255 vdd.n3367 vdd.n690 0.970197
R6256 vdd.n2610 vdd.t225 0.907421
R6257 vdd.n2998 vdd.t269 0.907421
R6258 vdd.n2297 vdd.t52 0.794056
R6259 vdd.n3553 vdd.t103 0.794056
R6260 vdd.n2322 vdd.t15 0.567326
R6261 vdd.n1119 vdd.t228 0.567326
R6262 vdd.n2616 vdd.t224 0.567326
R6263 vdd.n3004 vdd.t227 0.567326
R6264 vdd.n3198 vdd.t237 0.567326
R6265 vdd.t29 vdd.n662 0.567326
R6266 vdd.n2355 vdd.n1181 0.530988
R6267 vdd.n726 vdd.n682 0.530988
R6268 vdd.n464 vdd.n391 0.530988
R6269 vdd.n3622 vdd.n3621 0.530988
R6270 vdd.n3499 vdd.n3498 0.530988
R6271 vdd.n2344 vdd.n1517 0.530988
R6272 vdd.n1776 vdd.n1641 0.530988
R6273 vdd.n1878 vdd.n1877 0.530988
R6274 vdd.n4 vdd.n2 0.459552
R6275 vdd.n11 vdd.n9 0.459552
R6276 vdd.n329 vdd.n328 0.388379
R6277 vdd.n295 vdd.n293 0.388379
R6278 vdd.n270 vdd.n269 0.388379
R6279 vdd.n236 vdd.n234 0.388379
R6280 vdd.n227 vdd.n226 0.388379
R6281 vdd.n193 vdd.n191 0.388379
R6282 vdd.n168 vdd.n167 0.388379
R6283 vdd.n134 vdd.n132 0.388379
R6284 vdd.n126 vdd.n125 0.388379
R6285 vdd.n92 vdd.n90 0.388379
R6286 vdd.n67 vdd.n66 0.388379
R6287 vdd.n33 vdd.n31 0.388379
R6288 vdd.n2203 vdd.n2202 0.388379
R6289 vdd.n2169 vdd.n2167 0.388379
R6290 vdd.n2262 vdd.n2261 0.388379
R6291 vdd.n2228 vdd.n2226 0.388379
R6292 vdd.n2101 vdd.n2100 0.388379
R6293 vdd.n2067 vdd.n2065 0.388379
R6294 vdd.n2160 vdd.n2159 0.388379
R6295 vdd.n2126 vdd.n2124 0.388379
R6296 vdd.n2000 vdd.n1999 0.388379
R6297 vdd.n1966 vdd.n1964 0.388379
R6298 vdd.n2059 vdd.n2058 0.388379
R6299 vdd.n2025 vdd.n2023 0.388379
R6300 vdd.n19 vdd.n17 0.387128
R6301 vdd.n24 vdd.n22 0.387128
R6302 vdd.n6 vdd.n4 0.358259
R6303 vdd.n13 vdd.n11 0.358259
R6304 vdd.n276 vdd.n274 0.358259
R6305 vdd.n278 vdd.n276 0.358259
R6306 vdd.n280 vdd.n278 0.358259
R6307 vdd.n282 vdd.n280 0.358259
R6308 vdd.n284 vdd.n282 0.358259
R6309 vdd.n286 vdd.n284 0.358259
R6310 vdd.n288 vdd.n286 0.358259
R6311 vdd.n290 vdd.n288 0.358259
R6312 vdd.n332 vdd.n290 0.358259
R6313 vdd.n174 vdd.n172 0.358259
R6314 vdd.n176 vdd.n174 0.358259
R6315 vdd.n178 vdd.n176 0.358259
R6316 vdd.n180 vdd.n178 0.358259
R6317 vdd.n182 vdd.n180 0.358259
R6318 vdd.n184 vdd.n182 0.358259
R6319 vdd.n186 vdd.n184 0.358259
R6320 vdd.n188 vdd.n186 0.358259
R6321 vdd.n230 vdd.n188 0.358259
R6322 vdd.n73 vdd.n71 0.358259
R6323 vdd.n75 vdd.n73 0.358259
R6324 vdd.n77 vdd.n75 0.358259
R6325 vdd.n79 vdd.n77 0.358259
R6326 vdd.n81 vdd.n79 0.358259
R6327 vdd.n83 vdd.n81 0.358259
R6328 vdd.n85 vdd.n83 0.358259
R6329 vdd.n87 vdd.n85 0.358259
R6330 vdd.n129 vdd.n87 0.358259
R6331 vdd.n2265 vdd.n2223 0.358259
R6332 vdd.n2223 vdd.n2221 0.358259
R6333 vdd.n2221 vdd.n2219 0.358259
R6334 vdd.n2219 vdd.n2217 0.358259
R6335 vdd.n2217 vdd.n2215 0.358259
R6336 vdd.n2215 vdd.n2213 0.358259
R6337 vdd.n2213 vdd.n2211 0.358259
R6338 vdd.n2211 vdd.n2209 0.358259
R6339 vdd.n2209 vdd.n2207 0.358259
R6340 vdd.n2163 vdd.n2121 0.358259
R6341 vdd.n2121 vdd.n2119 0.358259
R6342 vdd.n2119 vdd.n2117 0.358259
R6343 vdd.n2117 vdd.n2115 0.358259
R6344 vdd.n2115 vdd.n2113 0.358259
R6345 vdd.n2113 vdd.n2111 0.358259
R6346 vdd.n2111 vdd.n2109 0.358259
R6347 vdd.n2109 vdd.n2107 0.358259
R6348 vdd.n2107 vdd.n2105 0.358259
R6349 vdd.n2062 vdd.n2020 0.358259
R6350 vdd.n2020 vdd.n2018 0.358259
R6351 vdd.n2018 vdd.n2016 0.358259
R6352 vdd.n2016 vdd.n2014 0.358259
R6353 vdd.n2014 vdd.n2012 0.358259
R6354 vdd.n2012 vdd.n2010 0.358259
R6355 vdd.n2010 vdd.n2008 0.358259
R6356 vdd.n2008 vdd.n2006 0.358259
R6357 vdd.n2006 vdd.n2004 0.358259
R6358 vdd.n2549 vdd.t276 0.340595
R6359 vdd.n1052 vdd.t234 0.340595
R6360 vdd.n3131 vdd.t223 0.340595
R6361 vdd.n877 vdd.t253 0.340595
R6362 vdd.n14 vdd.n6 0.334552
R6363 vdd.n14 vdd.n13 0.334552
R6364 vdd.n27 vdd.n19 0.21707
R6365 vdd.n27 vdd.n24 0.21707
R6366 vdd.n330 vdd.n292 0.155672
R6367 vdd.n322 vdd.n292 0.155672
R6368 vdd.n322 vdd.n321 0.155672
R6369 vdd.n321 vdd.n297 0.155672
R6370 vdd.n314 vdd.n297 0.155672
R6371 vdd.n314 vdd.n313 0.155672
R6372 vdd.n313 vdd.n301 0.155672
R6373 vdd.n306 vdd.n301 0.155672
R6374 vdd.n271 vdd.n233 0.155672
R6375 vdd.n263 vdd.n233 0.155672
R6376 vdd.n263 vdd.n262 0.155672
R6377 vdd.n262 vdd.n238 0.155672
R6378 vdd.n255 vdd.n238 0.155672
R6379 vdd.n255 vdd.n254 0.155672
R6380 vdd.n254 vdd.n242 0.155672
R6381 vdd.n247 vdd.n242 0.155672
R6382 vdd.n228 vdd.n190 0.155672
R6383 vdd.n220 vdd.n190 0.155672
R6384 vdd.n220 vdd.n219 0.155672
R6385 vdd.n219 vdd.n195 0.155672
R6386 vdd.n212 vdd.n195 0.155672
R6387 vdd.n212 vdd.n211 0.155672
R6388 vdd.n211 vdd.n199 0.155672
R6389 vdd.n204 vdd.n199 0.155672
R6390 vdd.n169 vdd.n131 0.155672
R6391 vdd.n161 vdd.n131 0.155672
R6392 vdd.n161 vdd.n160 0.155672
R6393 vdd.n160 vdd.n136 0.155672
R6394 vdd.n153 vdd.n136 0.155672
R6395 vdd.n153 vdd.n152 0.155672
R6396 vdd.n152 vdd.n140 0.155672
R6397 vdd.n145 vdd.n140 0.155672
R6398 vdd.n127 vdd.n89 0.155672
R6399 vdd.n119 vdd.n89 0.155672
R6400 vdd.n119 vdd.n118 0.155672
R6401 vdd.n118 vdd.n94 0.155672
R6402 vdd.n111 vdd.n94 0.155672
R6403 vdd.n111 vdd.n110 0.155672
R6404 vdd.n110 vdd.n98 0.155672
R6405 vdd.n103 vdd.n98 0.155672
R6406 vdd.n68 vdd.n30 0.155672
R6407 vdd.n60 vdd.n30 0.155672
R6408 vdd.n60 vdd.n59 0.155672
R6409 vdd.n59 vdd.n35 0.155672
R6410 vdd.n52 vdd.n35 0.155672
R6411 vdd.n52 vdd.n51 0.155672
R6412 vdd.n51 vdd.n39 0.155672
R6413 vdd.n44 vdd.n39 0.155672
R6414 vdd.n2204 vdd.n2166 0.155672
R6415 vdd.n2196 vdd.n2166 0.155672
R6416 vdd.n2196 vdd.n2195 0.155672
R6417 vdd.n2195 vdd.n2171 0.155672
R6418 vdd.n2188 vdd.n2171 0.155672
R6419 vdd.n2188 vdd.n2187 0.155672
R6420 vdd.n2187 vdd.n2175 0.155672
R6421 vdd.n2180 vdd.n2175 0.155672
R6422 vdd.n2263 vdd.n2225 0.155672
R6423 vdd.n2255 vdd.n2225 0.155672
R6424 vdd.n2255 vdd.n2254 0.155672
R6425 vdd.n2254 vdd.n2230 0.155672
R6426 vdd.n2247 vdd.n2230 0.155672
R6427 vdd.n2247 vdd.n2246 0.155672
R6428 vdd.n2246 vdd.n2234 0.155672
R6429 vdd.n2239 vdd.n2234 0.155672
R6430 vdd.n2102 vdd.n2064 0.155672
R6431 vdd.n2094 vdd.n2064 0.155672
R6432 vdd.n2094 vdd.n2093 0.155672
R6433 vdd.n2093 vdd.n2069 0.155672
R6434 vdd.n2086 vdd.n2069 0.155672
R6435 vdd.n2086 vdd.n2085 0.155672
R6436 vdd.n2085 vdd.n2073 0.155672
R6437 vdd.n2078 vdd.n2073 0.155672
R6438 vdd.n2161 vdd.n2123 0.155672
R6439 vdd.n2153 vdd.n2123 0.155672
R6440 vdd.n2153 vdd.n2152 0.155672
R6441 vdd.n2152 vdd.n2128 0.155672
R6442 vdd.n2145 vdd.n2128 0.155672
R6443 vdd.n2145 vdd.n2144 0.155672
R6444 vdd.n2144 vdd.n2132 0.155672
R6445 vdd.n2137 vdd.n2132 0.155672
R6446 vdd.n2001 vdd.n1963 0.155672
R6447 vdd.n1993 vdd.n1963 0.155672
R6448 vdd.n1993 vdd.n1992 0.155672
R6449 vdd.n1992 vdd.n1968 0.155672
R6450 vdd.n1985 vdd.n1968 0.155672
R6451 vdd.n1985 vdd.n1984 0.155672
R6452 vdd.n1984 vdd.n1972 0.155672
R6453 vdd.n1977 vdd.n1972 0.155672
R6454 vdd.n2060 vdd.n2022 0.155672
R6455 vdd.n2052 vdd.n2022 0.155672
R6456 vdd.n2052 vdd.n2051 0.155672
R6457 vdd.n2051 vdd.n2027 0.155672
R6458 vdd.n2044 vdd.n2027 0.155672
R6459 vdd.n2044 vdd.n2043 0.155672
R6460 vdd.n2043 vdd.n2031 0.155672
R6461 vdd.n2036 vdd.n2031 0.155672
R6462 vdd.n1186 vdd.n1178 0.152939
R6463 vdd.n1190 vdd.n1186 0.152939
R6464 vdd.n1191 vdd.n1190 0.152939
R6465 vdd.n1192 vdd.n1191 0.152939
R6466 vdd.n1193 vdd.n1192 0.152939
R6467 vdd.n1197 vdd.n1193 0.152939
R6468 vdd.n1198 vdd.n1197 0.152939
R6469 vdd.n1199 vdd.n1198 0.152939
R6470 vdd.n1200 vdd.n1199 0.152939
R6471 vdd.n1204 vdd.n1200 0.152939
R6472 vdd.n1205 vdd.n1204 0.152939
R6473 vdd.n1206 vdd.n1205 0.152939
R6474 vdd.n2438 vdd.n1206 0.152939
R6475 vdd.n2438 vdd.n2437 0.152939
R6476 vdd.n2437 vdd.n2436 0.152939
R6477 vdd.n2436 vdd.n1212 0.152939
R6478 vdd.n1217 vdd.n1212 0.152939
R6479 vdd.n1218 vdd.n1217 0.152939
R6480 vdd.n1219 vdd.n1218 0.152939
R6481 vdd.n1223 vdd.n1219 0.152939
R6482 vdd.n1224 vdd.n1223 0.152939
R6483 vdd.n1225 vdd.n1224 0.152939
R6484 vdd.n1226 vdd.n1225 0.152939
R6485 vdd.n1230 vdd.n1226 0.152939
R6486 vdd.n1231 vdd.n1230 0.152939
R6487 vdd.n1232 vdd.n1231 0.152939
R6488 vdd.n1233 vdd.n1232 0.152939
R6489 vdd.n1237 vdd.n1233 0.152939
R6490 vdd.n1238 vdd.n1237 0.152939
R6491 vdd.n1239 vdd.n1238 0.152939
R6492 vdd.n1240 vdd.n1239 0.152939
R6493 vdd.n1244 vdd.n1240 0.152939
R6494 vdd.n1245 vdd.n1244 0.152939
R6495 vdd.n1246 vdd.n1245 0.152939
R6496 vdd.n2399 vdd.n1246 0.152939
R6497 vdd.n2399 vdd.n2398 0.152939
R6498 vdd.n2398 vdd.n2397 0.152939
R6499 vdd.n2397 vdd.n1252 0.152939
R6500 vdd.n1257 vdd.n1252 0.152939
R6501 vdd.n1258 vdd.n1257 0.152939
R6502 vdd.n1259 vdd.n1258 0.152939
R6503 vdd.n1263 vdd.n1259 0.152939
R6504 vdd.n1264 vdd.n1263 0.152939
R6505 vdd.n1265 vdd.n1264 0.152939
R6506 vdd.n1266 vdd.n1265 0.152939
R6507 vdd.n1270 vdd.n1266 0.152939
R6508 vdd.n1271 vdd.n1270 0.152939
R6509 vdd.n1272 vdd.n1271 0.152939
R6510 vdd.n1273 vdd.n1272 0.152939
R6511 vdd.n1277 vdd.n1273 0.152939
R6512 vdd.n1278 vdd.n1277 0.152939
R6513 vdd.n2473 vdd.n1181 0.152939
R6514 vdd.n2269 vdd.n1578 0.152939
R6515 vdd.n2284 vdd.n1578 0.152939
R6516 vdd.n2285 vdd.n2284 0.152939
R6517 vdd.n2286 vdd.n2285 0.152939
R6518 vdd.n2286 vdd.n1567 0.152939
R6519 vdd.n2301 vdd.n1567 0.152939
R6520 vdd.n2302 vdd.n2301 0.152939
R6521 vdd.n2303 vdd.n2302 0.152939
R6522 vdd.n2303 vdd.n1556 0.152939
R6523 vdd.n2317 vdd.n1556 0.152939
R6524 vdd.n2318 vdd.n2317 0.152939
R6525 vdd.n2319 vdd.n2318 0.152939
R6526 vdd.n2319 vdd.n1544 0.152939
R6527 vdd.n2334 vdd.n1544 0.152939
R6528 vdd.n2335 vdd.n2334 0.152939
R6529 vdd.n2336 vdd.n2335 0.152939
R6530 vdd.n2336 vdd.n1532 0.152939
R6531 vdd.n2353 vdd.n1532 0.152939
R6532 vdd.n2354 vdd.n2353 0.152939
R6533 vdd.n2355 vdd.n2354 0.152939
R6534 vdd.n735 vdd.n730 0.152939
R6535 vdd.n736 vdd.n735 0.152939
R6536 vdd.n737 vdd.n736 0.152939
R6537 vdd.n738 vdd.n737 0.152939
R6538 vdd.n739 vdd.n738 0.152939
R6539 vdd.n740 vdd.n739 0.152939
R6540 vdd.n741 vdd.n740 0.152939
R6541 vdd.n742 vdd.n741 0.152939
R6542 vdd.n743 vdd.n742 0.152939
R6543 vdd.n744 vdd.n743 0.152939
R6544 vdd.n745 vdd.n744 0.152939
R6545 vdd.n746 vdd.n745 0.152939
R6546 vdd.n3455 vdd.n746 0.152939
R6547 vdd.n3455 vdd.n3454 0.152939
R6548 vdd.n3454 vdd.n3453 0.152939
R6549 vdd.n3453 vdd.n748 0.152939
R6550 vdd.n749 vdd.n748 0.152939
R6551 vdd.n750 vdd.n749 0.152939
R6552 vdd.n751 vdd.n750 0.152939
R6553 vdd.n752 vdd.n751 0.152939
R6554 vdd.n753 vdd.n752 0.152939
R6555 vdd.n754 vdd.n753 0.152939
R6556 vdd.n755 vdd.n754 0.152939
R6557 vdd.n756 vdd.n755 0.152939
R6558 vdd.n757 vdd.n756 0.152939
R6559 vdd.n758 vdd.n757 0.152939
R6560 vdd.n759 vdd.n758 0.152939
R6561 vdd.n760 vdd.n759 0.152939
R6562 vdd.n761 vdd.n760 0.152939
R6563 vdd.n762 vdd.n761 0.152939
R6564 vdd.n763 vdd.n762 0.152939
R6565 vdd.n764 vdd.n763 0.152939
R6566 vdd.n765 vdd.n764 0.152939
R6567 vdd.n766 vdd.n765 0.152939
R6568 vdd.n3409 vdd.n766 0.152939
R6569 vdd.n3409 vdd.n3408 0.152939
R6570 vdd.n3408 vdd.n3407 0.152939
R6571 vdd.n3407 vdd.n770 0.152939
R6572 vdd.n771 vdd.n770 0.152939
R6573 vdd.n772 vdd.n771 0.152939
R6574 vdd.n773 vdd.n772 0.152939
R6575 vdd.n774 vdd.n773 0.152939
R6576 vdd.n775 vdd.n774 0.152939
R6577 vdd.n776 vdd.n775 0.152939
R6578 vdd.n777 vdd.n776 0.152939
R6579 vdd.n778 vdd.n777 0.152939
R6580 vdd.n779 vdd.n778 0.152939
R6581 vdd.n780 vdd.n779 0.152939
R6582 vdd.n781 vdd.n780 0.152939
R6583 vdd.n782 vdd.n781 0.152939
R6584 vdd.n783 vdd.n782 0.152939
R6585 vdd.n727 vdd.n726 0.152939
R6586 vdd.n3506 vdd.n682 0.152939
R6587 vdd.n3507 vdd.n3506 0.152939
R6588 vdd.n3508 vdd.n3507 0.152939
R6589 vdd.n3508 vdd.n670 0.152939
R6590 vdd.n3523 vdd.n670 0.152939
R6591 vdd.n3524 vdd.n3523 0.152939
R6592 vdd.n3525 vdd.n3524 0.152939
R6593 vdd.n3525 vdd.n659 0.152939
R6594 vdd.n3539 vdd.n659 0.152939
R6595 vdd.n3540 vdd.n3539 0.152939
R6596 vdd.n3541 vdd.n3540 0.152939
R6597 vdd.n3541 vdd.n647 0.152939
R6598 vdd.n3556 vdd.n647 0.152939
R6599 vdd.n3557 vdd.n3556 0.152939
R6600 vdd.n3558 vdd.n3557 0.152939
R6601 vdd.n3558 vdd.n636 0.152939
R6602 vdd.n3575 vdd.n636 0.152939
R6603 vdd.n3576 vdd.n3575 0.152939
R6604 vdd.n3577 vdd.n3576 0.152939
R6605 vdd.n3577 vdd.n334 0.152939
R6606 vdd.n3670 vdd.n335 0.152939
R6607 vdd.n346 vdd.n335 0.152939
R6608 vdd.n347 vdd.n346 0.152939
R6609 vdd.n348 vdd.n347 0.152939
R6610 vdd.n355 vdd.n348 0.152939
R6611 vdd.n356 vdd.n355 0.152939
R6612 vdd.n357 vdd.n356 0.152939
R6613 vdd.n358 vdd.n357 0.152939
R6614 vdd.n366 vdd.n358 0.152939
R6615 vdd.n367 vdd.n366 0.152939
R6616 vdd.n368 vdd.n367 0.152939
R6617 vdd.n369 vdd.n368 0.152939
R6618 vdd.n377 vdd.n369 0.152939
R6619 vdd.n378 vdd.n377 0.152939
R6620 vdd.n379 vdd.n378 0.152939
R6621 vdd.n380 vdd.n379 0.152939
R6622 vdd.n388 vdd.n380 0.152939
R6623 vdd.n389 vdd.n388 0.152939
R6624 vdd.n390 vdd.n389 0.152939
R6625 vdd.n391 vdd.n390 0.152939
R6626 vdd.n464 vdd.n463 0.152939
R6627 vdd.n470 vdd.n463 0.152939
R6628 vdd.n471 vdd.n470 0.152939
R6629 vdd.n472 vdd.n471 0.152939
R6630 vdd.n472 vdd.n461 0.152939
R6631 vdd.n480 vdd.n461 0.152939
R6632 vdd.n481 vdd.n480 0.152939
R6633 vdd.n482 vdd.n481 0.152939
R6634 vdd.n482 vdd.n459 0.152939
R6635 vdd.n490 vdd.n459 0.152939
R6636 vdd.n491 vdd.n490 0.152939
R6637 vdd.n492 vdd.n491 0.152939
R6638 vdd.n492 vdd.n457 0.152939
R6639 vdd.n500 vdd.n457 0.152939
R6640 vdd.n501 vdd.n500 0.152939
R6641 vdd.n502 vdd.n501 0.152939
R6642 vdd.n502 vdd.n455 0.152939
R6643 vdd.n510 vdd.n455 0.152939
R6644 vdd.n511 vdd.n510 0.152939
R6645 vdd.n512 vdd.n511 0.152939
R6646 vdd.n512 vdd.n451 0.152939
R6647 vdd.n520 vdd.n451 0.152939
R6648 vdd.n521 vdd.n520 0.152939
R6649 vdd.n522 vdd.n521 0.152939
R6650 vdd.n522 vdd.n449 0.152939
R6651 vdd.n530 vdd.n449 0.152939
R6652 vdd.n531 vdd.n530 0.152939
R6653 vdd.n532 vdd.n531 0.152939
R6654 vdd.n532 vdd.n447 0.152939
R6655 vdd.n540 vdd.n447 0.152939
R6656 vdd.n541 vdd.n540 0.152939
R6657 vdd.n542 vdd.n541 0.152939
R6658 vdd.n542 vdd.n445 0.152939
R6659 vdd.n550 vdd.n445 0.152939
R6660 vdd.n551 vdd.n550 0.152939
R6661 vdd.n552 vdd.n551 0.152939
R6662 vdd.n552 vdd.n443 0.152939
R6663 vdd.n560 vdd.n443 0.152939
R6664 vdd.n561 vdd.n560 0.152939
R6665 vdd.n562 vdd.n561 0.152939
R6666 vdd.n562 vdd.n439 0.152939
R6667 vdd.n570 vdd.n439 0.152939
R6668 vdd.n571 vdd.n570 0.152939
R6669 vdd.n572 vdd.n571 0.152939
R6670 vdd.n572 vdd.n437 0.152939
R6671 vdd.n580 vdd.n437 0.152939
R6672 vdd.n581 vdd.n580 0.152939
R6673 vdd.n582 vdd.n581 0.152939
R6674 vdd.n582 vdd.n435 0.152939
R6675 vdd.n590 vdd.n435 0.152939
R6676 vdd.n591 vdd.n590 0.152939
R6677 vdd.n592 vdd.n591 0.152939
R6678 vdd.n592 vdd.n433 0.152939
R6679 vdd.n600 vdd.n433 0.152939
R6680 vdd.n601 vdd.n600 0.152939
R6681 vdd.n602 vdd.n601 0.152939
R6682 vdd.n602 vdd.n431 0.152939
R6683 vdd.n610 vdd.n431 0.152939
R6684 vdd.n611 vdd.n610 0.152939
R6685 vdd.n612 vdd.n611 0.152939
R6686 vdd.n612 vdd.n429 0.152939
R6687 vdd.n619 vdd.n429 0.152939
R6688 vdd.n3622 vdd.n619 0.152939
R6689 vdd.n3500 vdd.n3499 0.152939
R6690 vdd.n3500 vdd.n675 0.152939
R6691 vdd.n3514 vdd.n675 0.152939
R6692 vdd.n3515 vdd.n3514 0.152939
R6693 vdd.n3516 vdd.n3515 0.152939
R6694 vdd.n3516 vdd.n665 0.152939
R6695 vdd.n3531 vdd.n665 0.152939
R6696 vdd.n3532 vdd.n3531 0.152939
R6697 vdd.n3533 vdd.n3532 0.152939
R6698 vdd.n3533 vdd.n652 0.152939
R6699 vdd.n3547 vdd.n652 0.152939
R6700 vdd.n3548 vdd.n3547 0.152939
R6701 vdd.n3549 vdd.n3548 0.152939
R6702 vdd.n3549 vdd.n641 0.152939
R6703 vdd.n3564 vdd.n641 0.152939
R6704 vdd.n3565 vdd.n3564 0.152939
R6705 vdd.n3566 vdd.n3565 0.152939
R6706 vdd.n3568 vdd.n3566 0.152939
R6707 vdd.n3568 vdd.n3567 0.152939
R6708 vdd.n3567 vdd.n630 0.152939
R6709 vdd.n3585 vdd.n630 0.152939
R6710 vdd.n3586 vdd.n3585 0.152939
R6711 vdd.n3587 vdd.n3586 0.152939
R6712 vdd.n3587 vdd.n628 0.152939
R6713 vdd.n3592 vdd.n628 0.152939
R6714 vdd.n3593 vdd.n3592 0.152939
R6715 vdd.n3594 vdd.n3593 0.152939
R6716 vdd.n3594 vdd.n626 0.152939
R6717 vdd.n3599 vdd.n626 0.152939
R6718 vdd.n3600 vdd.n3599 0.152939
R6719 vdd.n3601 vdd.n3600 0.152939
R6720 vdd.n3601 vdd.n624 0.152939
R6721 vdd.n3607 vdd.n624 0.152939
R6722 vdd.n3608 vdd.n3607 0.152939
R6723 vdd.n3609 vdd.n3608 0.152939
R6724 vdd.n3609 vdd.n622 0.152939
R6725 vdd.n3614 vdd.n622 0.152939
R6726 vdd.n3615 vdd.n3614 0.152939
R6727 vdd.n3616 vdd.n3615 0.152939
R6728 vdd.n3616 vdd.n620 0.152939
R6729 vdd.n3621 vdd.n620 0.152939
R6730 vdd.n3498 vdd.n687 0.152939
R6731 vdd.n2366 vdd.n1517 0.152939
R6732 vdd.n1885 vdd.n1641 0.152939
R6733 vdd.n1886 vdd.n1885 0.152939
R6734 vdd.n1887 vdd.n1886 0.152939
R6735 vdd.n1887 vdd.n1629 0.152939
R6736 vdd.n1902 vdd.n1629 0.152939
R6737 vdd.n1903 vdd.n1902 0.152939
R6738 vdd.n1904 vdd.n1903 0.152939
R6739 vdd.n1904 vdd.n1619 0.152939
R6740 vdd.n1919 vdd.n1619 0.152939
R6741 vdd.n1920 vdd.n1919 0.152939
R6742 vdd.n1921 vdd.n1920 0.152939
R6743 vdd.n1921 vdd.n1606 0.152939
R6744 vdd.n1935 vdd.n1606 0.152939
R6745 vdd.n1936 vdd.n1935 0.152939
R6746 vdd.n1937 vdd.n1936 0.152939
R6747 vdd.n1937 vdd.n1595 0.152939
R6748 vdd.n1952 vdd.n1595 0.152939
R6749 vdd.n1953 vdd.n1952 0.152939
R6750 vdd.n1954 vdd.n1953 0.152939
R6751 vdd.n1954 vdd.n1584 0.152939
R6752 vdd.n2275 vdd.n1584 0.152939
R6753 vdd.n2276 vdd.n2275 0.152939
R6754 vdd.n2277 vdd.n2276 0.152939
R6755 vdd.n2277 vdd.n1572 0.152939
R6756 vdd.n2292 vdd.n1572 0.152939
R6757 vdd.n2293 vdd.n2292 0.152939
R6758 vdd.n2294 vdd.n2293 0.152939
R6759 vdd.n2294 vdd.n1562 0.152939
R6760 vdd.n2309 vdd.n1562 0.152939
R6761 vdd.n2310 vdd.n2309 0.152939
R6762 vdd.n2311 vdd.n2310 0.152939
R6763 vdd.n2311 vdd.n1549 0.152939
R6764 vdd.n2325 vdd.n1549 0.152939
R6765 vdd.n2326 vdd.n2325 0.152939
R6766 vdd.n2327 vdd.n2326 0.152939
R6767 vdd.n2327 vdd.n1539 0.152939
R6768 vdd.n2342 vdd.n1539 0.152939
R6769 vdd.n2343 vdd.n2342 0.152939
R6770 vdd.n2346 vdd.n2343 0.152939
R6771 vdd.n2346 vdd.n2345 0.152939
R6772 vdd.n2345 vdd.n2344 0.152939
R6773 vdd.n1877 vdd.n1646 0.152939
R6774 vdd.n1870 vdd.n1646 0.152939
R6775 vdd.n1870 vdd.n1869 0.152939
R6776 vdd.n1869 vdd.n1868 0.152939
R6777 vdd.n1868 vdd.n1683 0.152939
R6778 vdd.n1864 vdd.n1683 0.152939
R6779 vdd.n1864 vdd.n1863 0.152939
R6780 vdd.n1863 vdd.n1862 0.152939
R6781 vdd.n1862 vdd.n1689 0.152939
R6782 vdd.n1858 vdd.n1689 0.152939
R6783 vdd.n1858 vdd.n1857 0.152939
R6784 vdd.n1857 vdd.n1856 0.152939
R6785 vdd.n1856 vdd.n1695 0.152939
R6786 vdd.n1852 vdd.n1695 0.152939
R6787 vdd.n1852 vdd.n1851 0.152939
R6788 vdd.n1851 vdd.n1850 0.152939
R6789 vdd.n1850 vdd.n1701 0.152939
R6790 vdd.n1846 vdd.n1701 0.152939
R6791 vdd.n1846 vdd.n1845 0.152939
R6792 vdd.n1845 vdd.n1844 0.152939
R6793 vdd.n1844 vdd.n1709 0.152939
R6794 vdd.n1840 vdd.n1709 0.152939
R6795 vdd.n1840 vdd.n1839 0.152939
R6796 vdd.n1839 vdd.n1838 0.152939
R6797 vdd.n1838 vdd.n1715 0.152939
R6798 vdd.n1834 vdd.n1715 0.152939
R6799 vdd.n1834 vdd.n1833 0.152939
R6800 vdd.n1833 vdd.n1832 0.152939
R6801 vdd.n1832 vdd.n1721 0.152939
R6802 vdd.n1828 vdd.n1721 0.152939
R6803 vdd.n1828 vdd.n1827 0.152939
R6804 vdd.n1827 vdd.n1826 0.152939
R6805 vdd.n1826 vdd.n1727 0.152939
R6806 vdd.n1822 vdd.n1727 0.152939
R6807 vdd.n1822 vdd.n1821 0.152939
R6808 vdd.n1821 vdd.n1820 0.152939
R6809 vdd.n1820 vdd.n1733 0.152939
R6810 vdd.n1816 vdd.n1733 0.152939
R6811 vdd.n1816 vdd.n1815 0.152939
R6812 vdd.n1815 vdd.n1814 0.152939
R6813 vdd.n1814 vdd.n1739 0.152939
R6814 vdd.n1807 vdd.n1739 0.152939
R6815 vdd.n1807 vdd.n1806 0.152939
R6816 vdd.n1806 vdd.n1805 0.152939
R6817 vdd.n1805 vdd.n1744 0.152939
R6818 vdd.n1801 vdd.n1744 0.152939
R6819 vdd.n1801 vdd.n1800 0.152939
R6820 vdd.n1800 vdd.n1799 0.152939
R6821 vdd.n1799 vdd.n1750 0.152939
R6822 vdd.n1795 vdd.n1750 0.152939
R6823 vdd.n1795 vdd.n1794 0.152939
R6824 vdd.n1794 vdd.n1793 0.152939
R6825 vdd.n1793 vdd.n1756 0.152939
R6826 vdd.n1789 vdd.n1756 0.152939
R6827 vdd.n1789 vdd.n1788 0.152939
R6828 vdd.n1788 vdd.n1787 0.152939
R6829 vdd.n1787 vdd.n1762 0.152939
R6830 vdd.n1783 vdd.n1762 0.152939
R6831 vdd.n1783 vdd.n1782 0.152939
R6832 vdd.n1782 vdd.n1781 0.152939
R6833 vdd.n1781 vdd.n1768 0.152939
R6834 vdd.n1777 vdd.n1768 0.152939
R6835 vdd.n1777 vdd.n1776 0.152939
R6836 vdd.n1879 vdd.n1878 0.152939
R6837 vdd.n1879 vdd.n1635 0.152939
R6838 vdd.n1894 vdd.n1635 0.152939
R6839 vdd.n1895 vdd.n1894 0.152939
R6840 vdd.n1896 vdd.n1895 0.152939
R6841 vdd.n1896 vdd.n1624 0.152939
R6842 vdd.n1911 vdd.n1624 0.152939
R6843 vdd.n1912 vdd.n1911 0.152939
R6844 vdd.n1913 vdd.n1912 0.152939
R6845 vdd.n1913 vdd.n1613 0.152939
R6846 vdd.n1927 vdd.n1613 0.152939
R6847 vdd.n1928 vdd.n1927 0.152939
R6848 vdd.n1929 vdd.n1928 0.152939
R6849 vdd.n1929 vdd.n1601 0.152939
R6850 vdd.n1944 vdd.n1601 0.152939
R6851 vdd.n1945 vdd.n1944 0.152939
R6852 vdd.n1946 vdd.n1945 0.152939
R6853 vdd.n1946 vdd.n1590 0.152939
R6854 vdd.n1960 vdd.n1590 0.152939
R6855 vdd.n1961 vdd.n1960 0.152939
R6856 vdd.n1882 vdd.t211 0.113865
R6857 vdd.t160 vdd.n386 0.113865
R6858 vdd.n2474 vdd.n2473 0.110256
R6859 vdd.n3488 vdd.n727 0.110256
R6860 vdd.n3365 vdd.n687 0.110256
R6861 vdd.n2367 vdd.n2366 0.110256
R6862 vdd.n2269 vdd.n2268 0.0695946
R6863 vdd.n3671 vdd.n334 0.0695946
R6864 vdd.n3671 vdd.n3670 0.0695946
R6865 vdd.n2268 vdd.n1961 0.0695946
R6866 vdd.n2474 vdd.n1178 0.0431829
R6867 vdd.n2367 vdd.n1278 0.0431829
R6868 vdd.n3488 vdd.n730 0.0431829
R6869 vdd.n3365 vdd.n783 0.0431829
R6870 vdd vdd.n28 0.00833333
R6871 commonsourceibias.n25 commonsourceibias.t34 230.006
R6872 commonsourceibias.n91 commonsourceibias.t73 230.006
R6873 commonsourceibias.n218 commonsourceibias.t98 230.006
R6874 commonsourceibias.n154 commonsourceibias.t70 230.006
R6875 commonsourceibias.n322 commonsourceibias.t24 230.006
R6876 commonsourceibias.n281 commonsourceibias.t111 230.006
R6877 commonsourceibias.n483 commonsourceibias.t113 230.006
R6878 commonsourceibias.n419 commonsourceibias.t52 230.006
R6879 commonsourceibias.n70 commonsourceibias.t20 207.983
R6880 commonsourceibias.n136 commonsourceibias.t89 207.983
R6881 commonsourceibias.n263 commonsourceibias.t109 207.983
R6882 commonsourceibias.n199 commonsourceibias.t54 207.983
R6883 commonsourceibias.n368 commonsourceibias.t38 207.983
R6884 commonsourceibias.n402 commonsourceibias.t69 207.983
R6885 commonsourceibias.n529 commonsourceibias.t63 207.983
R6886 commonsourceibias.n465 commonsourceibias.t112 207.983
R6887 commonsourceibias.n10 commonsourceibias.t28 168.701
R6888 commonsourceibias.n63 commonsourceibias.t2 168.701
R6889 commonsourceibias.n57 commonsourceibias.t18 168.701
R6890 commonsourceibias.n16 commonsourceibias.t32 168.701
R6891 commonsourceibias.n49 commonsourceibias.t14 168.701
R6892 commonsourceibias.n43 commonsourceibias.t12 168.701
R6893 commonsourceibias.n19 commonsourceibias.t44 168.701
R6894 commonsourceibias.n21 commonsourceibias.t22 168.701
R6895 commonsourceibias.n23 commonsourceibias.t6 168.701
R6896 commonsourceibias.n26 commonsourceibias.t8 168.701
R6897 commonsourceibias.n1 commonsourceibias.t51 168.701
R6898 commonsourceibias.n129 commonsourceibias.t95 168.701
R6899 commonsourceibias.n123 commonsourceibias.t90 168.701
R6900 commonsourceibias.n7 commonsourceibias.t101 168.701
R6901 commonsourceibias.n115 commonsourceibias.t86 168.701
R6902 commonsourceibias.n109 commonsourceibias.t77 168.701
R6903 commonsourceibias.n85 commonsourceibias.t94 168.701
R6904 commonsourceibias.n87 commonsourceibias.t87 168.701
R6905 commonsourceibias.n89 commonsourceibias.t58 168.701
R6906 commonsourceibias.n92 commonsourceibias.t80 168.701
R6907 commonsourceibias.n219 commonsourceibias.t102 168.701
R6908 commonsourceibias.n216 commonsourceibias.t48 168.701
R6909 commonsourceibias.n214 commonsourceibias.t103 168.701
R6910 commonsourceibias.n212 commonsourceibias.t108 168.701
R6911 commonsourceibias.n236 commonsourceibias.t88 168.701
R6912 commonsourceibias.n242 commonsourceibias.t68 168.701
R6913 commonsourceibias.n209 commonsourceibias.t115 168.701
R6914 commonsourceibias.n250 commonsourceibias.t93 168.701
R6915 commonsourceibias.n256 commonsourceibias.t96 168.701
R6916 commonsourceibias.n203 commonsourceibias.t57 168.701
R6917 commonsourceibias.n139 commonsourceibias.t119 168.701
R6918 commonsourceibias.n192 commonsourceibias.t110 168.701
R6919 commonsourceibias.n186 commonsourceibias.t60 168.701
R6920 commonsourceibias.n145 commonsourceibias.t117 168.701
R6921 commonsourceibias.n178 commonsourceibias.t65 168.701
R6922 commonsourceibias.n172 commonsourceibias.t59 168.701
R6923 commonsourceibias.n148 commonsourceibias.t118 168.701
R6924 commonsourceibias.n150 commonsourceibias.t71 168.701
R6925 commonsourceibias.n152 commonsourceibias.t83 168.701
R6926 commonsourceibias.n155 commonsourceibias.t116 168.701
R6927 commonsourceibias.n323 commonsourceibias.t4 168.701
R6928 commonsourceibias.n320 commonsourceibias.t30 168.701
R6929 commonsourceibias.n318 commonsourceibias.t40 168.701
R6930 commonsourceibias.n316 commonsourceibias.t10 168.701
R6931 commonsourceibias.n340 commonsourceibias.t26 168.701
R6932 commonsourceibias.n346 commonsourceibias.t42 168.701
R6933 commonsourceibias.n348 commonsourceibias.t46 168.701
R6934 commonsourceibias.n355 commonsourceibias.t36 168.701
R6935 commonsourceibias.n361 commonsourceibias.t16 168.701
R6936 commonsourceibias.n308 commonsourceibias.t0 168.701
R6937 commonsourceibias.n267 commonsourceibias.t99 168.701
R6938 commonsourceibias.n395 commonsourceibias.t84 168.701
R6939 commonsourceibias.n389 commonsourceibias.t72 168.701
R6940 commonsourceibias.n382 commonsourceibias.t92 168.701
R6941 commonsourceibias.n380 commonsourceibias.t66 168.701
R6942 commonsourceibias.n282 commonsourceibias.t64 168.701
R6943 commonsourceibias.n279 commonsourceibias.t104 168.701
R6944 commonsourceibias.n277 commonsourceibias.t67 168.701
R6945 commonsourceibias.n275 commonsourceibias.t79 168.701
R6946 commonsourceibias.n299 commonsourceibias.t56 168.701
R6947 commonsourceibias.n484 commonsourceibias.t97 168.701
R6948 commonsourceibias.n481 commonsourceibias.t78 168.701
R6949 commonsourceibias.n479 commonsourceibias.t53 168.701
R6950 commonsourceibias.n477 commonsourceibias.t62 168.701
R6951 commonsourceibias.n501 commonsourceibias.t82 168.701
R6952 commonsourceibias.n507 commonsourceibias.t85 168.701
R6953 commonsourceibias.n509 commonsourceibias.t76 168.701
R6954 commonsourceibias.n516 commonsourceibias.t100 168.701
R6955 commonsourceibias.n522 commonsourceibias.t91 168.701
R6956 commonsourceibias.n469 commonsourceibias.t81 168.701
R6957 commonsourceibias.n420 commonsourceibias.t61 168.701
R6958 commonsourceibias.n417 commonsourceibias.t75 168.701
R6959 commonsourceibias.n415 commonsourceibias.t55 168.701
R6960 commonsourceibias.n413 commonsourceibias.t105 168.701
R6961 commonsourceibias.n437 commonsourceibias.t74 168.701
R6962 commonsourceibias.n443 commonsourceibias.t49 168.701
R6963 commonsourceibias.n445 commonsourceibias.t106 168.701
R6964 commonsourceibias.n452 commonsourceibias.t114 168.701
R6965 commonsourceibias.n458 commonsourceibias.t50 168.701
R6966 commonsourceibias.n405 commonsourceibias.t107 168.701
R6967 commonsourceibias.n27 commonsourceibias.n24 161.3
R6968 commonsourceibias.n29 commonsourceibias.n28 161.3
R6969 commonsourceibias.n31 commonsourceibias.n30 161.3
R6970 commonsourceibias.n32 commonsourceibias.n22 161.3
R6971 commonsourceibias.n34 commonsourceibias.n33 161.3
R6972 commonsourceibias.n36 commonsourceibias.n35 161.3
R6973 commonsourceibias.n37 commonsourceibias.n20 161.3
R6974 commonsourceibias.n39 commonsourceibias.n38 161.3
R6975 commonsourceibias.n41 commonsourceibias.n40 161.3
R6976 commonsourceibias.n42 commonsourceibias.n18 161.3
R6977 commonsourceibias.n45 commonsourceibias.n44 161.3
R6978 commonsourceibias.n46 commonsourceibias.n17 161.3
R6979 commonsourceibias.n48 commonsourceibias.n47 161.3
R6980 commonsourceibias.n50 commonsourceibias.n15 161.3
R6981 commonsourceibias.n52 commonsourceibias.n51 161.3
R6982 commonsourceibias.n53 commonsourceibias.n14 161.3
R6983 commonsourceibias.n55 commonsourceibias.n54 161.3
R6984 commonsourceibias.n56 commonsourceibias.n13 161.3
R6985 commonsourceibias.n59 commonsourceibias.n58 161.3
R6986 commonsourceibias.n60 commonsourceibias.n12 161.3
R6987 commonsourceibias.n62 commonsourceibias.n61 161.3
R6988 commonsourceibias.n64 commonsourceibias.n11 161.3
R6989 commonsourceibias.n66 commonsourceibias.n65 161.3
R6990 commonsourceibias.n68 commonsourceibias.n67 161.3
R6991 commonsourceibias.n69 commonsourceibias.n9 161.3
R6992 commonsourceibias.n93 commonsourceibias.n90 161.3
R6993 commonsourceibias.n95 commonsourceibias.n94 161.3
R6994 commonsourceibias.n97 commonsourceibias.n96 161.3
R6995 commonsourceibias.n98 commonsourceibias.n88 161.3
R6996 commonsourceibias.n100 commonsourceibias.n99 161.3
R6997 commonsourceibias.n102 commonsourceibias.n101 161.3
R6998 commonsourceibias.n103 commonsourceibias.n86 161.3
R6999 commonsourceibias.n105 commonsourceibias.n104 161.3
R7000 commonsourceibias.n107 commonsourceibias.n106 161.3
R7001 commonsourceibias.n108 commonsourceibias.n84 161.3
R7002 commonsourceibias.n111 commonsourceibias.n110 161.3
R7003 commonsourceibias.n112 commonsourceibias.n8 161.3
R7004 commonsourceibias.n114 commonsourceibias.n113 161.3
R7005 commonsourceibias.n116 commonsourceibias.n6 161.3
R7006 commonsourceibias.n118 commonsourceibias.n117 161.3
R7007 commonsourceibias.n119 commonsourceibias.n5 161.3
R7008 commonsourceibias.n121 commonsourceibias.n120 161.3
R7009 commonsourceibias.n122 commonsourceibias.n4 161.3
R7010 commonsourceibias.n125 commonsourceibias.n124 161.3
R7011 commonsourceibias.n126 commonsourceibias.n3 161.3
R7012 commonsourceibias.n128 commonsourceibias.n127 161.3
R7013 commonsourceibias.n130 commonsourceibias.n2 161.3
R7014 commonsourceibias.n132 commonsourceibias.n131 161.3
R7015 commonsourceibias.n134 commonsourceibias.n133 161.3
R7016 commonsourceibias.n135 commonsourceibias.n0 161.3
R7017 commonsourceibias.n262 commonsourceibias.n202 161.3
R7018 commonsourceibias.n261 commonsourceibias.n260 161.3
R7019 commonsourceibias.n259 commonsourceibias.n258 161.3
R7020 commonsourceibias.n257 commonsourceibias.n204 161.3
R7021 commonsourceibias.n255 commonsourceibias.n254 161.3
R7022 commonsourceibias.n253 commonsourceibias.n205 161.3
R7023 commonsourceibias.n252 commonsourceibias.n251 161.3
R7024 commonsourceibias.n249 commonsourceibias.n206 161.3
R7025 commonsourceibias.n248 commonsourceibias.n247 161.3
R7026 commonsourceibias.n246 commonsourceibias.n207 161.3
R7027 commonsourceibias.n245 commonsourceibias.n244 161.3
R7028 commonsourceibias.n243 commonsourceibias.n208 161.3
R7029 commonsourceibias.n241 commonsourceibias.n240 161.3
R7030 commonsourceibias.n239 commonsourceibias.n210 161.3
R7031 commonsourceibias.n238 commonsourceibias.n237 161.3
R7032 commonsourceibias.n235 commonsourceibias.n211 161.3
R7033 commonsourceibias.n234 commonsourceibias.n233 161.3
R7034 commonsourceibias.n232 commonsourceibias.n231 161.3
R7035 commonsourceibias.n230 commonsourceibias.n213 161.3
R7036 commonsourceibias.n229 commonsourceibias.n228 161.3
R7037 commonsourceibias.n227 commonsourceibias.n226 161.3
R7038 commonsourceibias.n225 commonsourceibias.n215 161.3
R7039 commonsourceibias.n224 commonsourceibias.n223 161.3
R7040 commonsourceibias.n222 commonsourceibias.n221 161.3
R7041 commonsourceibias.n220 commonsourceibias.n217 161.3
R7042 commonsourceibias.n156 commonsourceibias.n153 161.3
R7043 commonsourceibias.n158 commonsourceibias.n157 161.3
R7044 commonsourceibias.n160 commonsourceibias.n159 161.3
R7045 commonsourceibias.n161 commonsourceibias.n151 161.3
R7046 commonsourceibias.n163 commonsourceibias.n162 161.3
R7047 commonsourceibias.n165 commonsourceibias.n164 161.3
R7048 commonsourceibias.n166 commonsourceibias.n149 161.3
R7049 commonsourceibias.n168 commonsourceibias.n167 161.3
R7050 commonsourceibias.n170 commonsourceibias.n169 161.3
R7051 commonsourceibias.n171 commonsourceibias.n147 161.3
R7052 commonsourceibias.n174 commonsourceibias.n173 161.3
R7053 commonsourceibias.n175 commonsourceibias.n146 161.3
R7054 commonsourceibias.n177 commonsourceibias.n176 161.3
R7055 commonsourceibias.n179 commonsourceibias.n144 161.3
R7056 commonsourceibias.n181 commonsourceibias.n180 161.3
R7057 commonsourceibias.n182 commonsourceibias.n143 161.3
R7058 commonsourceibias.n184 commonsourceibias.n183 161.3
R7059 commonsourceibias.n185 commonsourceibias.n142 161.3
R7060 commonsourceibias.n188 commonsourceibias.n187 161.3
R7061 commonsourceibias.n189 commonsourceibias.n141 161.3
R7062 commonsourceibias.n191 commonsourceibias.n190 161.3
R7063 commonsourceibias.n193 commonsourceibias.n140 161.3
R7064 commonsourceibias.n195 commonsourceibias.n194 161.3
R7065 commonsourceibias.n197 commonsourceibias.n196 161.3
R7066 commonsourceibias.n198 commonsourceibias.n138 161.3
R7067 commonsourceibias.n367 commonsourceibias.n307 161.3
R7068 commonsourceibias.n366 commonsourceibias.n365 161.3
R7069 commonsourceibias.n364 commonsourceibias.n363 161.3
R7070 commonsourceibias.n362 commonsourceibias.n309 161.3
R7071 commonsourceibias.n360 commonsourceibias.n359 161.3
R7072 commonsourceibias.n358 commonsourceibias.n310 161.3
R7073 commonsourceibias.n357 commonsourceibias.n356 161.3
R7074 commonsourceibias.n354 commonsourceibias.n311 161.3
R7075 commonsourceibias.n353 commonsourceibias.n352 161.3
R7076 commonsourceibias.n351 commonsourceibias.n312 161.3
R7077 commonsourceibias.n350 commonsourceibias.n349 161.3
R7078 commonsourceibias.n347 commonsourceibias.n313 161.3
R7079 commonsourceibias.n345 commonsourceibias.n344 161.3
R7080 commonsourceibias.n343 commonsourceibias.n314 161.3
R7081 commonsourceibias.n342 commonsourceibias.n341 161.3
R7082 commonsourceibias.n339 commonsourceibias.n315 161.3
R7083 commonsourceibias.n338 commonsourceibias.n337 161.3
R7084 commonsourceibias.n336 commonsourceibias.n335 161.3
R7085 commonsourceibias.n334 commonsourceibias.n317 161.3
R7086 commonsourceibias.n333 commonsourceibias.n332 161.3
R7087 commonsourceibias.n331 commonsourceibias.n330 161.3
R7088 commonsourceibias.n329 commonsourceibias.n319 161.3
R7089 commonsourceibias.n328 commonsourceibias.n327 161.3
R7090 commonsourceibias.n326 commonsourceibias.n325 161.3
R7091 commonsourceibias.n324 commonsourceibias.n321 161.3
R7092 commonsourceibias.n301 commonsourceibias.n300 161.3
R7093 commonsourceibias.n298 commonsourceibias.n274 161.3
R7094 commonsourceibias.n297 commonsourceibias.n296 161.3
R7095 commonsourceibias.n295 commonsourceibias.n294 161.3
R7096 commonsourceibias.n293 commonsourceibias.n276 161.3
R7097 commonsourceibias.n292 commonsourceibias.n291 161.3
R7098 commonsourceibias.n290 commonsourceibias.n289 161.3
R7099 commonsourceibias.n288 commonsourceibias.n278 161.3
R7100 commonsourceibias.n287 commonsourceibias.n286 161.3
R7101 commonsourceibias.n285 commonsourceibias.n284 161.3
R7102 commonsourceibias.n283 commonsourceibias.n280 161.3
R7103 commonsourceibias.n377 commonsourceibias.n273 161.3
R7104 commonsourceibias.n401 commonsourceibias.n266 161.3
R7105 commonsourceibias.n400 commonsourceibias.n399 161.3
R7106 commonsourceibias.n398 commonsourceibias.n397 161.3
R7107 commonsourceibias.n396 commonsourceibias.n268 161.3
R7108 commonsourceibias.n394 commonsourceibias.n393 161.3
R7109 commonsourceibias.n392 commonsourceibias.n269 161.3
R7110 commonsourceibias.n391 commonsourceibias.n390 161.3
R7111 commonsourceibias.n388 commonsourceibias.n270 161.3
R7112 commonsourceibias.n387 commonsourceibias.n386 161.3
R7113 commonsourceibias.n385 commonsourceibias.n271 161.3
R7114 commonsourceibias.n384 commonsourceibias.n383 161.3
R7115 commonsourceibias.n381 commonsourceibias.n272 161.3
R7116 commonsourceibias.n379 commonsourceibias.n378 161.3
R7117 commonsourceibias.n528 commonsourceibias.n468 161.3
R7118 commonsourceibias.n527 commonsourceibias.n526 161.3
R7119 commonsourceibias.n525 commonsourceibias.n524 161.3
R7120 commonsourceibias.n523 commonsourceibias.n470 161.3
R7121 commonsourceibias.n521 commonsourceibias.n520 161.3
R7122 commonsourceibias.n519 commonsourceibias.n471 161.3
R7123 commonsourceibias.n518 commonsourceibias.n517 161.3
R7124 commonsourceibias.n515 commonsourceibias.n472 161.3
R7125 commonsourceibias.n514 commonsourceibias.n513 161.3
R7126 commonsourceibias.n512 commonsourceibias.n473 161.3
R7127 commonsourceibias.n511 commonsourceibias.n510 161.3
R7128 commonsourceibias.n508 commonsourceibias.n474 161.3
R7129 commonsourceibias.n506 commonsourceibias.n505 161.3
R7130 commonsourceibias.n504 commonsourceibias.n475 161.3
R7131 commonsourceibias.n503 commonsourceibias.n502 161.3
R7132 commonsourceibias.n500 commonsourceibias.n476 161.3
R7133 commonsourceibias.n499 commonsourceibias.n498 161.3
R7134 commonsourceibias.n497 commonsourceibias.n496 161.3
R7135 commonsourceibias.n495 commonsourceibias.n478 161.3
R7136 commonsourceibias.n494 commonsourceibias.n493 161.3
R7137 commonsourceibias.n492 commonsourceibias.n491 161.3
R7138 commonsourceibias.n490 commonsourceibias.n480 161.3
R7139 commonsourceibias.n489 commonsourceibias.n488 161.3
R7140 commonsourceibias.n487 commonsourceibias.n486 161.3
R7141 commonsourceibias.n485 commonsourceibias.n482 161.3
R7142 commonsourceibias.n464 commonsourceibias.n404 161.3
R7143 commonsourceibias.n463 commonsourceibias.n462 161.3
R7144 commonsourceibias.n461 commonsourceibias.n460 161.3
R7145 commonsourceibias.n459 commonsourceibias.n406 161.3
R7146 commonsourceibias.n457 commonsourceibias.n456 161.3
R7147 commonsourceibias.n455 commonsourceibias.n407 161.3
R7148 commonsourceibias.n454 commonsourceibias.n453 161.3
R7149 commonsourceibias.n451 commonsourceibias.n408 161.3
R7150 commonsourceibias.n450 commonsourceibias.n449 161.3
R7151 commonsourceibias.n448 commonsourceibias.n409 161.3
R7152 commonsourceibias.n447 commonsourceibias.n446 161.3
R7153 commonsourceibias.n444 commonsourceibias.n410 161.3
R7154 commonsourceibias.n442 commonsourceibias.n441 161.3
R7155 commonsourceibias.n440 commonsourceibias.n411 161.3
R7156 commonsourceibias.n439 commonsourceibias.n438 161.3
R7157 commonsourceibias.n436 commonsourceibias.n412 161.3
R7158 commonsourceibias.n435 commonsourceibias.n434 161.3
R7159 commonsourceibias.n433 commonsourceibias.n432 161.3
R7160 commonsourceibias.n431 commonsourceibias.n414 161.3
R7161 commonsourceibias.n430 commonsourceibias.n429 161.3
R7162 commonsourceibias.n428 commonsourceibias.n427 161.3
R7163 commonsourceibias.n426 commonsourceibias.n416 161.3
R7164 commonsourceibias.n425 commonsourceibias.n424 161.3
R7165 commonsourceibias.n423 commonsourceibias.n422 161.3
R7166 commonsourceibias.n421 commonsourceibias.n418 161.3
R7167 commonsourceibias.n80 commonsourceibias.n78 81.5057
R7168 commonsourceibias.n304 commonsourceibias.n302 81.5057
R7169 commonsourceibias.n80 commonsourceibias.n79 80.9324
R7170 commonsourceibias.n82 commonsourceibias.n81 80.9324
R7171 commonsourceibias.n77 commonsourceibias.n76 80.9324
R7172 commonsourceibias.n75 commonsourceibias.n74 80.9324
R7173 commonsourceibias.n73 commonsourceibias.n72 80.9324
R7174 commonsourceibias.n371 commonsourceibias.n370 80.9324
R7175 commonsourceibias.n373 commonsourceibias.n372 80.9324
R7176 commonsourceibias.n375 commonsourceibias.n374 80.9324
R7177 commonsourceibias.n306 commonsourceibias.n305 80.9324
R7178 commonsourceibias.n304 commonsourceibias.n303 80.9324
R7179 commonsourceibias.n71 commonsourceibias.n70 80.6037
R7180 commonsourceibias.n137 commonsourceibias.n136 80.6037
R7181 commonsourceibias.n264 commonsourceibias.n263 80.6037
R7182 commonsourceibias.n200 commonsourceibias.n199 80.6037
R7183 commonsourceibias.n369 commonsourceibias.n368 80.6037
R7184 commonsourceibias.n403 commonsourceibias.n402 80.6037
R7185 commonsourceibias.n530 commonsourceibias.n529 80.6037
R7186 commonsourceibias.n466 commonsourceibias.n465 80.6037
R7187 commonsourceibias.n65 commonsourceibias.n64 56.5617
R7188 commonsourceibias.n51 commonsourceibias.n50 56.5617
R7189 commonsourceibias.n42 commonsourceibias.n41 56.5617
R7190 commonsourceibias.n28 commonsourceibias.n27 56.5617
R7191 commonsourceibias.n131 commonsourceibias.n130 56.5617
R7192 commonsourceibias.n117 commonsourceibias.n116 56.5617
R7193 commonsourceibias.n108 commonsourceibias.n107 56.5617
R7194 commonsourceibias.n94 commonsourceibias.n93 56.5617
R7195 commonsourceibias.n221 commonsourceibias.n220 56.5617
R7196 commonsourceibias.n235 commonsourceibias.n234 56.5617
R7197 commonsourceibias.n244 commonsourceibias.n243 56.5617
R7198 commonsourceibias.n258 commonsourceibias.n257 56.5617
R7199 commonsourceibias.n194 commonsourceibias.n193 56.5617
R7200 commonsourceibias.n180 commonsourceibias.n179 56.5617
R7201 commonsourceibias.n171 commonsourceibias.n170 56.5617
R7202 commonsourceibias.n157 commonsourceibias.n156 56.5617
R7203 commonsourceibias.n325 commonsourceibias.n324 56.5617
R7204 commonsourceibias.n339 commonsourceibias.n338 56.5617
R7205 commonsourceibias.n349 commonsourceibias.n347 56.5617
R7206 commonsourceibias.n363 commonsourceibias.n362 56.5617
R7207 commonsourceibias.n397 commonsourceibias.n396 56.5617
R7208 commonsourceibias.n383 commonsourceibias.n381 56.5617
R7209 commonsourceibias.n284 commonsourceibias.n283 56.5617
R7210 commonsourceibias.n298 commonsourceibias.n297 56.5617
R7211 commonsourceibias.n486 commonsourceibias.n485 56.5617
R7212 commonsourceibias.n500 commonsourceibias.n499 56.5617
R7213 commonsourceibias.n510 commonsourceibias.n508 56.5617
R7214 commonsourceibias.n524 commonsourceibias.n523 56.5617
R7215 commonsourceibias.n422 commonsourceibias.n421 56.5617
R7216 commonsourceibias.n436 commonsourceibias.n435 56.5617
R7217 commonsourceibias.n446 commonsourceibias.n444 56.5617
R7218 commonsourceibias.n460 commonsourceibias.n459 56.5617
R7219 commonsourceibias.n56 commonsourceibias.n55 56.0773
R7220 commonsourceibias.n37 commonsourceibias.n36 56.0773
R7221 commonsourceibias.n122 commonsourceibias.n121 56.0773
R7222 commonsourceibias.n103 commonsourceibias.n102 56.0773
R7223 commonsourceibias.n230 commonsourceibias.n229 56.0773
R7224 commonsourceibias.n249 commonsourceibias.n248 56.0773
R7225 commonsourceibias.n185 commonsourceibias.n184 56.0773
R7226 commonsourceibias.n166 commonsourceibias.n165 56.0773
R7227 commonsourceibias.n334 commonsourceibias.n333 56.0773
R7228 commonsourceibias.n354 commonsourceibias.n353 56.0773
R7229 commonsourceibias.n388 commonsourceibias.n387 56.0773
R7230 commonsourceibias.n293 commonsourceibias.n292 56.0773
R7231 commonsourceibias.n495 commonsourceibias.n494 56.0773
R7232 commonsourceibias.n515 commonsourceibias.n514 56.0773
R7233 commonsourceibias.n431 commonsourceibias.n430 56.0773
R7234 commonsourceibias.n451 commonsourceibias.n450 56.0773
R7235 commonsourceibias.n70 commonsourceibias.n69 46.0096
R7236 commonsourceibias.n136 commonsourceibias.n135 46.0096
R7237 commonsourceibias.n263 commonsourceibias.n262 46.0096
R7238 commonsourceibias.n199 commonsourceibias.n198 46.0096
R7239 commonsourceibias.n368 commonsourceibias.n367 46.0096
R7240 commonsourceibias.n402 commonsourceibias.n401 46.0096
R7241 commonsourceibias.n529 commonsourceibias.n528 46.0096
R7242 commonsourceibias.n465 commonsourceibias.n464 46.0096
R7243 commonsourceibias.n58 commonsourceibias.n12 41.5458
R7244 commonsourceibias.n33 commonsourceibias.n32 41.5458
R7245 commonsourceibias.n124 commonsourceibias.n3 41.5458
R7246 commonsourceibias.n99 commonsourceibias.n98 41.5458
R7247 commonsourceibias.n226 commonsourceibias.n225 41.5458
R7248 commonsourceibias.n251 commonsourceibias.n205 41.5458
R7249 commonsourceibias.n187 commonsourceibias.n141 41.5458
R7250 commonsourceibias.n162 commonsourceibias.n161 41.5458
R7251 commonsourceibias.n330 commonsourceibias.n329 41.5458
R7252 commonsourceibias.n356 commonsourceibias.n310 41.5458
R7253 commonsourceibias.n390 commonsourceibias.n269 41.5458
R7254 commonsourceibias.n289 commonsourceibias.n288 41.5458
R7255 commonsourceibias.n491 commonsourceibias.n490 41.5458
R7256 commonsourceibias.n517 commonsourceibias.n471 41.5458
R7257 commonsourceibias.n427 commonsourceibias.n426 41.5458
R7258 commonsourceibias.n453 commonsourceibias.n407 41.5458
R7259 commonsourceibias.n48 commonsourceibias.n17 40.577
R7260 commonsourceibias.n44 commonsourceibias.n17 40.577
R7261 commonsourceibias.n114 commonsourceibias.n8 40.577
R7262 commonsourceibias.n110 commonsourceibias.n8 40.577
R7263 commonsourceibias.n237 commonsourceibias.n210 40.577
R7264 commonsourceibias.n241 commonsourceibias.n210 40.577
R7265 commonsourceibias.n177 commonsourceibias.n146 40.577
R7266 commonsourceibias.n173 commonsourceibias.n146 40.577
R7267 commonsourceibias.n341 commonsourceibias.n314 40.577
R7268 commonsourceibias.n345 commonsourceibias.n314 40.577
R7269 commonsourceibias.n379 commonsourceibias.n273 40.577
R7270 commonsourceibias.n300 commonsourceibias.n273 40.577
R7271 commonsourceibias.n502 commonsourceibias.n475 40.577
R7272 commonsourceibias.n506 commonsourceibias.n475 40.577
R7273 commonsourceibias.n438 commonsourceibias.n411 40.577
R7274 commonsourceibias.n442 commonsourceibias.n411 40.577
R7275 commonsourceibias.n62 commonsourceibias.n12 39.6083
R7276 commonsourceibias.n32 commonsourceibias.n31 39.6083
R7277 commonsourceibias.n128 commonsourceibias.n3 39.6083
R7278 commonsourceibias.n98 commonsourceibias.n97 39.6083
R7279 commonsourceibias.n225 commonsourceibias.n224 39.6083
R7280 commonsourceibias.n255 commonsourceibias.n205 39.6083
R7281 commonsourceibias.n191 commonsourceibias.n141 39.6083
R7282 commonsourceibias.n161 commonsourceibias.n160 39.6083
R7283 commonsourceibias.n329 commonsourceibias.n328 39.6083
R7284 commonsourceibias.n360 commonsourceibias.n310 39.6083
R7285 commonsourceibias.n394 commonsourceibias.n269 39.6083
R7286 commonsourceibias.n288 commonsourceibias.n287 39.6083
R7287 commonsourceibias.n490 commonsourceibias.n489 39.6083
R7288 commonsourceibias.n521 commonsourceibias.n471 39.6083
R7289 commonsourceibias.n426 commonsourceibias.n425 39.6083
R7290 commonsourceibias.n457 commonsourceibias.n407 39.6083
R7291 commonsourceibias.n26 commonsourceibias.n25 33.0515
R7292 commonsourceibias.n92 commonsourceibias.n91 33.0515
R7293 commonsourceibias.n155 commonsourceibias.n154 33.0515
R7294 commonsourceibias.n219 commonsourceibias.n218 33.0515
R7295 commonsourceibias.n323 commonsourceibias.n322 33.0515
R7296 commonsourceibias.n282 commonsourceibias.n281 33.0515
R7297 commonsourceibias.n484 commonsourceibias.n483 33.0515
R7298 commonsourceibias.n420 commonsourceibias.n419 33.0515
R7299 commonsourceibias.n25 commonsourceibias.n24 28.5514
R7300 commonsourceibias.n91 commonsourceibias.n90 28.5514
R7301 commonsourceibias.n218 commonsourceibias.n217 28.5514
R7302 commonsourceibias.n154 commonsourceibias.n153 28.5514
R7303 commonsourceibias.n322 commonsourceibias.n321 28.5514
R7304 commonsourceibias.n281 commonsourceibias.n280 28.5514
R7305 commonsourceibias.n483 commonsourceibias.n482 28.5514
R7306 commonsourceibias.n419 commonsourceibias.n418 28.5514
R7307 commonsourceibias.n69 commonsourceibias.n68 26.0455
R7308 commonsourceibias.n135 commonsourceibias.n134 26.0455
R7309 commonsourceibias.n262 commonsourceibias.n261 26.0455
R7310 commonsourceibias.n198 commonsourceibias.n197 26.0455
R7311 commonsourceibias.n367 commonsourceibias.n366 26.0455
R7312 commonsourceibias.n401 commonsourceibias.n400 26.0455
R7313 commonsourceibias.n528 commonsourceibias.n527 26.0455
R7314 commonsourceibias.n464 commonsourceibias.n463 26.0455
R7315 commonsourceibias.n55 commonsourceibias.n14 25.0767
R7316 commonsourceibias.n38 commonsourceibias.n37 25.0767
R7317 commonsourceibias.n121 commonsourceibias.n5 25.0767
R7318 commonsourceibias.n104 commonsourceibias.n103 25.0767
R7319 commonsourceibias.n231 commonsourceibias.n230 25.0767
R7320 commonsourceibias.n248 commonsourceibias.n207 25.0767
R7321 commonsourceibias.n184 commonsourceibias.n143 25.0767
R7322 commonsourceibias.n167 commonsourceibias.n166 25.0767
R7323 commonsourceibias.n335 commonsourceibias.n334 25.0767
R7324 commonsourceibias.n353 commonsourceibias.n312 25.0767
R7325 commonsourceibias.n387 commonsourceibias.n271 25.0767
R7326 commonsourceibias.n294 commonsourceibias.n293 25.0767
R7327 commonsourceibias.n496 commonsourceibias.n495 25.0767
R7328 commonsourceibias.n514 commonsourceibias.n473 25.0767
R7329 commonsourceibias.n432 commonsourceibias.n431 25.0767
R7330 commonsourceibias.n450 commonsourceibias.n409 25.0767
R7331 commonsourceibias.n51 commonsourceibias.n16 24.3464
R7332 commonsourceibias.n41 commonsourceibias.n19 24.3464
R7333 commonsourceibias.n117 commonsourceibias.n7 24.3464
R7334 commonsourceibias.n107 commonsourceibias.n85 24.3464
R7335 commonsourceibias.n234 commonsourceibias.n212 24.3464
R7336 commonsourceibias.n244 commonsourceibias.n209 24.3464
R7337 commonsourceibias.n180 commonsourceibias.n145 24.3464
R7338 commonsourceibias.n170 commonsourceibias.n148 24.3464
R7339 commonsourceibias.n338 commonsourceibias.n316 24.3464
R7340 commonsourceibias.n349 commonsourceibias.n348 24.3464
R7341 commonsourceibias.n383 commonsourceibias.n382 24.3464
R7342 commonsourceibias.n297 commonsourceibias.n275 24.3464
R7343 commonsourceibias.n499 commonsourceibias.n477 24.3464
R7344 commonsourceibias.n510 commonsourceibias.n509 24.3464
R7345 commonsourceibias.n435 commonsourceibias.n413 24.3464
R7346 commonsourceibias.n446 commonsourceibias.n445 24.3464
R7347 commonsourceibias.n65 commonsourceibias.n10 23.8546
R7348 commonsourceibias.n27 commonsourceibias.n26 23.8546
R7349 commonsourceibias.n131 commonsourceibias.n1 23.8546
R7350 commonsourceibias.n93 commonsourceibias.n92 23.8546
R7351 commonsourceibias.n220 commonsourceibias.n219 23.8546
R7352 commonsourceibias.n258 commonsourceibias.n203 23.8546
R7353 commonsourceibias.n194 commonsourceibias.n139 23.8546
R7354 commonsourceibias.n156 commonsourceibias.n155 23.8546
R7355 commonsourceibias.n324 commonsourceibias.n323 23.8546
R7356 commonsourceibias.n363 commonsourceibias.n308 23.8546
R7357 commonsourceibias.n397 commonsourceibias.n267 23.8546
R7358 commonsourceibias.n283 commonsourceibias.n282 23.8546
R7359 commonsourceibias.n485 commonsourceibias.n484 23.8546
R7360 commonsourceibias.n524 commonsourceibias.n469 23.8546
R7361 commonsourceibias.n421 commonsourceibias.n420 23.8546
R7362 commonsourceibias.n460 commonsourceibias.n405 23.8546
R7363 commonsourceibias.n64 commonsourceibias.n63 16.9689
R7364 commonsourceibias.n28 commonsourceibias.n23 16.9689
R7365 commonsourceibias.n130 commonsourceibias.n129 16.9689
R7366 commonsourceibias.n94 commonsourceibias.n89 16.9689
R7367 commonsourceibias.n221 commonsourceibias.n216 16.9689
R7368 commonsourceibias.n257 commonsourceibias.n256 16.9689
R7369 commonsourceibias.n193 commonsourceibias.n192 16.9689
R7370 commonsourceibias.n157 commonsourceibias.n152 16.9689
R7371 commonsourceibias.n325 commonsourceibias.n320 16.9689
R7372 commonsourceibias.n362 commonsourceibias.n361 16.9689
R7373 commonsourceibias.n396 commonsourceibias.n395 16.9689
R7374 commonsourceibias.n284 commonsourceibias.n279 16.9689
R7375 commonsourceibias.n486 commonsourceibias.n481 16.9689
R7376 commonsourceibias.n523 commonsourceibias.n522 16.9689
R7377 commonsourceibias.n422 commonsourceibias.n417 16.9689
R7378 commonsourceibias.n459 commonsourceibias.n458 16.9689
R7379 commonsourceibias.n50 commonsourceibias.n49 16.477
R7380 commonsourceibias.n43 commonsourceibias.n42 16.477
R7381 commonsourceibias.n116 commonsourceibias.n115 16.477
R7382 commonsourceibias.n109 commonsourceibias.n108 16.477
R7383 commonsourceibias.n236 commonsourceibias.n235 16.477
R7384 commonsourceibias.n243 commonsourceibias.n242 16.477
R7385 commonsourceibias.n179 commonsourceibias.n178 16.477
R7386 commonsourceibias.n172 commonsourceibias.n171 16.477
R7387 commonsourceibias.n340 commonsourceibias.n339 16.477
R7388 commonsourceibias.n347 commonsourceibias.n346 16.477
R7389 commonsourceibias.n381 commonsourceibias.n380 16.477
R7390 commonsourceibias.n299 commonsourceibias.n298 16.477
R7391 commonsourceibias.n501 commonsourceibias.n500 16.477
R7392 commonsourceibias.n508 commonsourceibias.n507 16.477
R7393 commonsourceibias.n437 commonsourceibias.n436 16.477
R7394 commonsourceibias.n444 commonsourceibias.n443 16.477
R7395 commonsourceibias.n57 commonsourceibias.n56 15.9852
R7396 commonsourceibias.n36 commonsourceibias.n21 15.9852
R7397 commonsourceibias.n123 commonsourceibias.n122 15.9852
R7398 commonsourceibias.n102 commonsourceibias.n87 15.9852
R7399 commonsourceibias.n229 commonsourceibias.n214 15.9852
R7400 commonsourceibias.n250 commonsourceibias.n249 15.9852
R7401 commonsourceibias.n186 commonsourceibias.n185 15.9852
R7402 commonsourceibias.n165 commonsourceibias.n150 15.9852
R7403 commonsourceibias.n333 commonsourceibias.n318 15.9852
R7404 commonsourceibias.n355 commonsourceibias.n354 15.9852
R7405 commonsourceibias.n389 commonsourceibias.n388 15.9852
R7406 commonsourceibias.n292 commonsourceibias.n277 15.9852
R7407 commonsourceibias.n494 commonsourceibias.n479 15.9852
R7408 commonsourceibias.n516 commonsourceibias.n515 15.9852
R7409 commonsourceibias.n430 commonsourceibias.n415 15.9852
R7410 commonsourceibias.n452 commonsourceibias.n451 15.9852
R7411 commonsourceibias.n73 commonsourceibias.n71 13.2057
R7412 commonsourceibias.n371 commonsourceibias.n369 13.2057
R7413 commonsourceibias.n532 commonsourceibias.n265 10.122
R7414 commonsourceibias.n112 commonsourceibias.n83 9.50363
R7415 commonsourceibias.n377 commonsourceibias.n376 9.50363
R7416 commonsourceibias.n201 commonsourceibias.n137 8.7339
R7417 commonsourceibias.n467 commonsourceibias.n403 8.7339
R7418 commonsourceibias.n58 commonsourceibias.n57 8.60764
R7419 commonsourceibias.n33 commonsourceibias.n21 8.60764
R7420 commonsourceibias.n124 commonsourceibias.n123 8.60764
R7421 commonsourceibias.n99 commonsourceibias.n87 8.60764
R7422 commonsourceibias.n226 commonsourceibias.n214 8.60764
R7423 commonsourceibias.n251 commonsourceibias.n250 8.60764
R7424 commonsourceibias.n187 commonsourceibias.n186 8.60764
R7425 commonsourceibias.n162 commonsourceibias.n150 8.60764
R7426 commonsourceibias.n330 commonsourceibias.n318 8.60764
R7427 commonsourceibias.n356 commonsourceibias.n355 8.60764
R7428 commonsourceibias.n390 commonsourceibias.n389 8.60764
R7429 commonsourceibias.n289 commonsourceibias.n277 8.60764
R7430 commonsourceibias.n491 commonsourceibias.n479 8.60764
R7431 commonsourceibias.n517 commonsourceibias.n516 8.60764
R7432 commonsourceibias.n427 commonsourceibias.n415 8.60764
R7433 commonsourceibias.n453 commonsourceibias.n452 8.60764
R7434 commonsourceibias.n532 commonsourceibias.n531 8.46921
R7435 commonsourceibias.n49 commonsourceibias.n48 8.11581
R7436 commonsourceibias.n44 commonsourceibias.n43 8.11581
R7437 commonsourceibias.n115 commonsourceibias.n114 8.11581
R7438 commonsourceibias.n110 commonsourceibias.n109 8.11581
R7439 commonsourceibias.n237 commonsourceibias.n236 8.11581
R7440 commonsourceibias.n242 commonsourceibias.n241 8.11581
R7441 commonsourceibias.n178 commonsourceibias.n177 8.11581
R7442 commonsourceibias.n173 commonsourceibias.n172 8.11581
R7443 commonsourceibias.n341 commonsourceibias.n340 8.11581
R7444 commonsourceibias.n346 commonsourceibias.n345 8.11581
R7445 commonsourceibias.n380 commonsourceibias.n379 8.11581
R7446 commonsourceibias.n300 commonsourceibias.n299 8.11581
R7447 commonsourceibias.n502 commonsourceibias.n501 8.11581
R7448 commonsourceibias.n507 commonsourceibias.n506 8.11581
R7449 commonsourceibias.n438 commonsourceibias.n437 8.11581
R7450 commonsourceibias.n443 commonsourceibias.n442 8.11581
R7451 commonsourceibias.n63 commonsourceibias.n62 7.62397
R7452 commonsourceibias.n31 commonsourceibias.n23 7.62397
R7453 commonsourceibias.n129 commonsourceibias.n128 7.62397
R7454 commonsourceibias.n97 commonsourceibias.n89 7.62397
R7455 commonsourceibias.n224 commonsourceibias.n216 7.62397
R7456 commonsourceibias.n256 commonsourceibias.n255 7.62397
R7457 commonsourceibias.n192 commonsourceibias.n191 7.62397
R7458 commonsourceibias.n160 commonsourceibias.n152 7.62397
R7459 commonsourceibias.n328 commonsourceibias.n320 7.62397
R7460 commonsourceibias.n361 commonsourceibias.n360 7.62397
R7461 commonsourceibias.n395 commonsourceibias.n394 7.62397
R7462 commonsourceibias.n287 commonsourceibias.n279 7.62397
R7463 commonsourceibias.n489 commonsourceibias.n481 7.62397
R7464 commonsourceibias.n522 commonsourceibias.n521 7.62397
R7465 commonsourceibias.n425 commonsourceibias.n417 7.62397
R7466 commonsourceibias.n458 commonsourceibias.n457 7.62397
R7467 commonsourceibias.n265 commonsourceibias.n264 5.00473
R7468 commonsourceibias.n201 commonsourceibias.n200 5.00473
R7469 commonsourceibias.n531 commonsourceibias.n530 5.00473
R7470 commonsourceibias.n467 commonsourceibias.n466 5.00473
R7471 commonsourceibias commonsourceibias.n532 4.08303
R7472 commonsourceibias.n265 commonsourceibias.n201 3.72967
R7473 commonsourceibias.n531 commonsourceibias.n467 3.72967
R7474 commonsourceibias.n78 commonsourceibias.t9 2.82907
R7475 commonsourceibias.n78 commonsourceibias.t35 2.82907
R7476 commonsourceibias.n79 commonsourceibias.t23 2.82907
R7477 commonsourceibias.n79 commonsourceibias.t7 2.82907
R7478 commonsourceibias.n81 commonsourceibias.t13 2.82907
R7479 commonsourceibias.n81 commonsourceibias.t45 2.82907
R7480 commonsourceibias.n76 commonsourceibias.t33 2.82907
R7481 commonsourceibias.n76 commonsourceibias.t15 2.82907
R7482 commonsourceibias.n74 commonsourceibias.t3 2.82907
R7483 commonsourceibias.n74 commonsourceibias.t19 2.82907
R7484 commonsourceibias.n72 commonsourceibias.t21 2.82907
R7485 commonsourceibias.n72 commonsourceibias.t29 2.82907
R7486 commonsourceibias.n370 commonsourceibias.t1 2.82907
R7487 commonsourceibias.n370 commonsourceibias.t39 2.82907
R7488 commonsourceibias.n372 commonsourceibias.t37 2.82907
R7489 commonsourceibias.n372 commonsourceibias.t17 2.82907
R7490 commonsourceibias.n374 commonsourceibias.t43 2.82907
R7491 commonsourceibias.n374 commonsourceibias.t47 2.82907
R7492 commonsourceibias.n305 commonsourceibias.t11 2.82907
R7493 commonsourceibias.n305 commonsourceibias.t27 2.82907
R7494 commonsourceibias.n303 commonsourceibias.t31 2.82907
R7495 commonsourceibias.n303 commonsourceibias.t41 2.82907
R7496 commonsourceibias.n302 commonsourceibias.t25 2.82907
R7497 commonsourceibias.n302 commonsourceibias.t5 2.82907
R7498 commonsourceibias.n68 commonsourceibias.n10 0.738255
R7499 commonsourceibias.n134 commonsourceibias.n1 0.738255
R7500 commonsourceibias.n261 commonsourceibias.n203 0.738255
R7501 commonsourceibias.n197 commonsourceibias.n139 0.738255
R7502 commonsourceibias.n366 commonsourceibias.n308 0.738255
R7503 commonsourceibias.n400 commonsourceibias.n267 0.738255
R7504 commonsourceibias.n527 commonsourceibias.n469 0.738255
R7505 commonsourceibias.n463 commonsourceibias.n405 0.738255
R7506 commonsourceibias.n75 commonsourceibias.n73 0.573776
R7507 commonsourceibias.n77 commonsourceibias.n75 0.573776
R7508 commonsourceibias.n82 commonsourceibias.n80 0.573776
R7509 commonsourceibias.n306 commonsourceibias.n304 0.573776
R7510 commonsourceibias.n375 commonsourceibias.n373 0.573776
R7511 commonsourceibias.n373 commonsourceibias.n371 0.573776
R7512 commonsourceibias.n83 commonsourceibias.n77 0.287138
R7513 commonsourceibias.n83 commonsourceibias.n82 0.287138
R7514 commonsourceibias.n376 commonsourceibias.n306 0.287138
R7515 commonsourceibias.n376 commonsourceibias.n375 0.287138
R7516 commonsourceibias.n71 commonsourceibias.n9 0.285035
R7517 commonsourceibias.n137 commonsourceibias.n0 0.285035
R7518 commonsourceibias.n264 commonsourceibias.n202 0.285035
R7519 commonsourceibias.n200 commonsourceibias.n138 0.285035
R7520 commonsourceibias.n369 commonsourceibias.n307 0.285035
R7521 commonsourceibias.n403 commonsourceibias.n266 0.285035
R7522 commonsourceibias.n530 commonsourceibias.n468 0.285035
R7523 commonsourceibias.n466 commonsourceibias.n404 0.285035
R7524 commonsourceibias.n16 commonsourceibias.n14 0.246418
R7525 commonsourceibias.n38 commonsourceibias.n19 0.246418
R7526 commonsourceibias.n7 commonsourceibias.n5 0.246418
R7527 commonsourceibias.n104 commonsourceibias.n85 0.246418
R7528 commonsourceibias.n231 commonsourceibias.n212 0.246418
R7529 commonsourceibias.n209 commonsourceibias.n207 0.246418
R7530 commonsourceibias.n145 commonsourceibias.n143 0.246418
R7531 commonsourceibias.n167 commonsourceibias.n148 0.246418
R7532 commonsourceibias.n335 commonsourceibias.n316 0.246418
R7533 commonsourceibias.n348 commonsourceibias.n312 0.246418
R7534 commonsourceibias.n382 commonsourceibias.n271 0.246418
R7535 commonsourceibias.n294 commonsourceibias.n275 0.246418
R7536 commonsourceibias.n496 commonsourceibias.n477 0.246418
R7537 commonsourceibias.n509 commonsourceibias.n473 0.246418
R7538 commonsourceibias.n432 commonsourceibias.n413 0.246418
R7539 commonsourceibias.n445 commonsourceibias.n409 0.246418
R7540 commonsourceibias.n67 commonsourceibias.n9 0.189894
R7541 commonsourceibias.n67 commonsourceibias.n66 0.189894
R7542 commonsourceibias.n66 commonsourceibias.n11 0.189894
R7543 commonsourceibias.n61 commonsourceibias.n11 0.189894
R7544 commonsourceibias.n61 commonsourceibias.n60 0.189894
R7545 commonsourceibias.n60 commonsourceibias.n59 0.189894
R7546 commonsourceibias.n59 commonsourceibias.n13 0.189894
R7547 commonsourceibias.n54 commonsourceibias.n13 0.189894
R7548 commonsourceibias.n54 commonsourceibias.n53 0.189894
R7549 commonsourceibias.n53 commonsourceibias.n52 0.189894
R7550 commonsourceibias.n52 commonsourceibias.n15 0.189894
R7551 commonsourceibias.n47 commonsourceibias.n15 0.189894
R7552 commonsourceibias.n47 commonsourceibias.n46 0.189894
R7553 commonsourceibias.n46 commonsourceibias.n45 0.189894
R7554 commonsourceibias.n45 commonsourceibias.n18 0.189894
R7555 commonsourceibias.n40 commonsourceibias.n18 0.189894
R7556 commonsourceibias.n40 commonsourceibias.n39 0.189894
R7557 commonsourceibias.n39 commonsourceibias.n20 0.189894
R7558 commonsourceibias.n35 commonsourceibias.n20 0.189894
R7559 commonsourceibias.n35 commonsourceibias.n34 0.189894
R7560 commonsourceibias.n34 commonsourceibias.n22 0.189894
R7561 commonsourceibias.n30 commonsourceibias.n22 0.189894
R7562 commonsourceibias.n30 commonsourceibias.n29 0.189894
R7563 commonsourceibias.n29 commonsourceibias.n24 0.189894
R7564 commonsourceibias.n111 commonsourceibias.n84 0.189894
R7565 commonsourceibias.n106 commonsourceibias.n84 0.189894
R7566 commonsourceibias.n106 commonsourceibias.n105 0.189894
R7567 commonsourceibias.n105 commonsourceibias.n86 0.189894
R7568 commonsourceibias.n101 commonsourceibias.n86 0.189894
R7569 commonsourceibias.n101 commonsourceibias.n100 0.189894
R7570 commonsourceibias.n100 commonsourceibias.n88 0.189894
R7571 commonsourceibias.n96 commonsourceibias.n88 0.189894
R7572 commonsourceibias.n96 commonsourceibias.n95 0.189894
R7573 commonsourceibias.n95 commonsourceibias.n90 0.189894
R7574 commonsourceibias.n133 commonsourceibias.n0 0.189894
R7575 commonsourceibias.n133 commonsourceibias.n132 0.189894
R7576 commonsourceibias.n132 commonsourceibias.n2 0.189894
R7577 commonsourceibias.n127 commonsourceibias.n2 0.189894
R7578 commonsourceibias.n127 commonsourceibias.n126 0.189894
R7579 commonsourceibias.n126 commonsourceibias.n125 0.189894
R7580 commonsourceibias.n125 commonsourceibias.n4 0.189894
R7581 commonsourceibias.n120 commonsourceibias.n4 0.189894
R7582 commonsourceibias.n120 commonsourceibias.n119 0.189894
R7583 commonsourceibias.n119 commonsourceibias.n118 0.189894
R7584 commonsourceibias.n118 commonsourceibias.n6 0.189894
R7585 commonsourceibias.n113 commonsourceibias.n6 0.189894
R7586 commonsourceibias.n260 commonsourceibias.n202 0.189894
R7587 commonsourceibias.n260 commonsourceibias.n259 0.189894
R7588 commonsourceibias.n259 commonsourceibias.n204 0.189894
R7589 commonsourceibias.n254 commonsourceibias.n204 0.189894
R7590 commonsourceibias.n254 commonsourceibias.n253 0.189894
R7591 commonsourceibias.n253 commonsourceibias.n252 0.189894
R7592 commonsourceibias.n252 commonsourceibias.n206 0.189894
R7593 commonsourceibias.n247 commonsourceibias.n206 0.189894
R7594 commonsourceibias.n247 commonsourceibias.n246 0.189894
R7595 commonsourceibias.n246 commonsourceibias.n245 0.189894
R7596 commonsourceibias.n245 commonsourceibias.n208 0.189894
R7597 commonsourceibias.n240 commonsourceibias.n208 0.189894
R7598 commonsourceibias.n240 commonsourceibias.n239 0.189894
R7599 commonsourceibias.n239 commonsourceibias.n238 0.189894
R7600 commonsourceibias.n238 commonsourceibias.n211 0.189894
R7601 commonsourceibias.n233 commonsourceibias.n211 0.189894
R7602 commonsourceibias.n233 commonsourceibias.n232 0.189894
R7603 commonsourceibias.n232 commonsourceibias.n213 0.189894
R7604 commonsourceibias.n228 commonsourceibias.n213 0.189894
R7605 commonsourceibias.n228 commonsourceibias.n227 0.189894
R7606 commonsourceibias.n227 commonsourceibias.n215 0.189894
R7607 commonsourceibias.n223 commonsourceibias.n215 0.189894
R7608 commonsourceibias.n223 commonsourceibias.n222 0.189894
R7609 commonsourceibias.n222 commonsourceibias.n217 0.189894
R7610 commonsourceibias.n196 commonsourceibias.n138 0.189894
R7611 commonsourceibias.n196 commonsourceibias.n195 0.189894
R7612 commonsourceibias.n195 commonsourceibias.n140 0.189894
R7613 commonsourceibias.n190 commonsourceibias.n140 0.189894
R7614 commonsourceibias.n190 commonsourceibias.n189 0.189894
R7615 commonsourceibias.n189 commonsourceibias.n188 0.189894
R7616 commonsourceibias.n188 commonsourceibias.n142 0.189894
R7617 commonsourceibias.n183 commonsourceibias.n142 0.189894
R7618 commonsourceibias.n183 commonsourceibias.n182 0.189894
R7619 commonsourceibias.n182 commonsourceibias.n181 0.189894
R7620 commonsourceibias.n181 commonsourceibias.n144 0.189894
R7621 commonsourceibias.n176 commonsourceibias.n144 0.189894
R7622 commonsourceibias.n176 commonsourceibias.n175 0.189894
R7623 commonsourceibias.n175 commonsourceibias.n174 0.189894
R7624 commonsourceibias.n174 commonsourceibias.n147 0.189894
R7625 commonsourceibias.n169 commonsourceibias.n147 0.189894
R7626 commonsourceibias.n169 commonsourceibias.n168 0.189894
R7627 commonsourceibias.n168 commonsourceibias.n149 0.189894
R7628 commonsourceibias.n164 commonsourceibias.n149 0.189894
R7629 commonsourceibias.n164 commonsourceibias.n163 0.189894
R7630 commonsourceibias.n163 commonsourceibias.n151 0.189894
R7631 commonsourceibias.n159 commonsourceibias.n151 0.189894
R7632 commonsourceibias.n159 commonsourceibias.n158 0.189894
R7633 commonsourceibias.n158 commonsourceibias.n153 0.189894
R7634 commonsourceibias.n326 commonsourceibias.n321 0.189894
R7635 commonsourceibias.n327 commonsourceibias.n326 0.189894
R7636 commonsourceibias.n327 commonsourceibias.n319 0.189894
R7637 commonsourceibias.n331 commonsourceibias.n319 0.189894
R7638 commonsourceibias.n332 commonsourceibias.n331 0.189894
R7639 commonsourceibias.n332 commonsourceibias.n317 0.189894
R7640 commonsourceibias.n336 commonsourceibias.n317 0.189894
R7641 commonsourceibias.n337 commonsourceibias.n336 0.189894
R7642 commonsourceibias.n337 commonsourceibias.n315 0.189894
R7643 commonsourceibias.n342 commonsourceibias.n315 0.189894
R7644 commonsourceibias.n343 commonsourceibias.n342 0.189894
R7645 commonsourceibias.n344 commonsourceibias.n343 0.189894
R7646 commonsourceibias.n344 commonsourceibias.n313 0.189894
R7647 commonsourceibias.n350 commonsourceibias.n313 0.189894
R7648 commonsourceibias.n351 commonsourceibias.n350 0.189894
R7649 commonsourceibias.n352 commonsourceibias.n351 0.189894
R7650 commonsourceibias.n352 commonsourceibias.n311 0.189894
R7651 commonsourceibias.n357 commonsourceibias.n311 0.189894
R7652 commonsourceibias.n358 commonsourceibias.n357 0.189894
R7653 commonsourceibias.n359 commonsourceibias.n358 0.189894
R7654 commonsourceibias.n359 commonsourceibias.n309 0.189894
R7655 commonsourceibias.n364 commonsourceibias.n309 0.189894
R7656 commonsourceibias.n365 commonsourceibias.n364 0.189894
R7657 commonsourceibias.n365 commonsourceibias.n307 0.189894
R7658 commonsourceibias.n285 commonsourceibias.n280 0.189894
R7659 commonsourceibias.n286 commonsourceibias.n285 0.189894
R7660 commonsourceibias.n286 commonsourceibias.n278 0.189894
R7661 commonsourceibias.n290 commonsourceibias.n278 0.189894
R7662 commonsourceibias.n291 commonsourceibias.n290 0.189894
R7663 commonsourceibias.n291 commonsourceibias.n276 0.189894
R7664 commonsourceibias.n295 commonsourceibias.n276 0.189894
R7665 commonsourceibias.n296 commonsourceibias.n295 0.189894
R7666 commonsourceibias.n296 commonsourceibias.n274 0.189894
R7667 commonsourceibias.n301 commonsourceibias.n274 0.189894
R7668 commonsourceibias.n378 commonsourceibias.n272 0.189894
R7669 commonsourceibias.n384 commonsourceibias.n272 0.189894
R7670 commonsourceibias.n385 commonsourceibias.n384 0.189894
R7671 commonsourceibias.n386 commonsourceibias.n385 0.189894
R7672 commonsourceibias.n386 commonsourceibias.n270 0.189894
R7673 commonsourceibias.n391 commonsourceibias.n270 0.189894
R7674 commonsourceibias.n392 commonsourceibias.n391 0.189894
R7675 commonsourceibias.n393 commonsourceibias.n392 0.189894
R7676 commonsourceibias.n393 commonsourceibias.n268 0.189894
R7677 commonsourceibias.n398 commonsourceibias.n268 0.189894
R7678 commonsourceibias.n399 commonsourceibias.n398 0.189894
R7679 commonsourceibias.n399 commonsourceibias.n266 0.189894
R7680 commonsourceibias.n487 commonsourceibias.n482 0.189894
R7681 commonsourceibias.n488 commonsourceibias.n487 0.189894
R7682 commonsourceibias.n488 commonsourceibias.n480 0.189894
R7683 commonsourceibias.n492 commonsourceibias.n480 0.189894
R7684 commonsourceibias.n493 commonsourceibias.n492 0.189894
R7685 commonsourceibias.n493 commonsourceibias.n478 0.189894
R7686 commonsourceibias.n497 commonsourceibias.n478 0.189894
R7687 commonsourceibias.n498 commonsourceibias.n497 0.189894
R7688 commonsourceibias.n498 commonsourceibias.n476 0.189894
R7689 commonsourceibias.n503 commonsourceibias.n476 0.189894
R7690 commonsourceibias.n504 commonsourceibias.n503 0.189894
R7691 commonsourceibias.n505 commonsourceibias.n504 0.189894
R7692 commonsourceibias.n505 commonsourceibias.n474 0.189894
R7693 commonsourceibias.n511 commonsourceibias.n474 0.189894
R7694 commonsourceibias.n512 commonsourceibias.n511 0.189894
R7695 commonsourceibias.n513 commonsourceibias.n512 0.189894
R7696 commonsourceibias.n513 commonsourceibias.n472 0.189894
R7697 commonsourceibias.n518 commonsourceibias.n472 0.189894
R7698 commonsourceibias.n519 commonsourceibias.n518 0.189894
R7699 commonsourceibias.n520 commonsourceibias.n519 0.189894
R7700 commonsourceibias.n520 commonsourceibias.n470 0.189894
R7701 commonsourceibias.n525 commonsourceibias.n470 0.189894
R7702 commonsourceibias.n526 commonsourceibias.n525 0.189894
R7703 commonsourceibias.n526 commonsourceibias.n468 0.189894
R7704 commonsourceibias.n423 commonsourceibias.n418 0.189894
R7705 commonsourceibias.n424 commonsourceibias.n423 0.189894
R7706 commonsourceibias.n424 commonsourceibias.n416 0.189894
R7707 commonsourceibias.n428 commonsourceibias.n416 0.189894
R7708 commonsourceibias.n429 commonsourceibias.n428 0.189894
R7709 commonsourceibias.n429 commonsourceibias.n414 0.189894
R7710 commonsourceibias.n433 commonsourceibias.n414 0.189894
R7711 commonsourceibias.n434 commonsourceibias.n433 0.189894
R7712 commonsourceibias.n434 commonsourceibias.n412 0.189894
R7713 commonsourceibias.n439 commonsourceibias.n412 0.189894
R7714 commonsourceibias.n440 commonsourceibias.n439 0.189894
R7715 commonsourceibias.n441 commonsourceibias.n440 0.189894
R7716 commonsourceibias.n441 commonsourceibias.n410 0.189894
R7717 commonsourceibias.n447 commonsourceibias.n410 0.189894
R7718 commonsourceibias.n448 commonsourceibias.n447 0.189894
R7719 commonsourceibias.n449 commonsourceibias.n448 0.189894
R7720 commonsourceibias.n449 commonsourceibias.n408 0.189894
R7721 commonsourceibias.n454 commonsourceibias.n408 0.189894
R7722 commonsourceibias.n455 commonsourceibias.n454 0.189894
R7723 commonsourceibias.n456 commonsourceibias.n455 0.189894
R7724 commonsourceibias.n456 commonsourceibias.n406 0.189894
R7725 commonsourceibias.n461 commonsourceibias.n406 0.189894
R7726 commonsourceibias.n462 commonsourceibias.n461 0.189894
R7727 commonsourceibias.n462 commonsourceibias.n404 0.189894
R7728 commonsourceibias.n112 commonsourceibias.n111 0.170955
R7729 commonsourceibias.n113 commonsourceibias.n112 0.170955
R7730 commonsourceibias.n377 commonsourceibias.n301 0.170955
R7731 commonsourceibias.n378 commonsourceibias.n377 0.170955
R7732 gnd.n7211 gnd.n394 1810.87
R7733 gnd.n2339 gnd.n2338 927.927
R7734 gnd.n7674 gnd.n172 838.452
R7735 gnd.n7661 gnd.n170 838.452
R7736 gnd.n5212 gnd.n3058 838.452
R7737 gnd.n5281 gnd.n3060 838.452
R7738 gnd.n6356 gnd.n2575 838.452
R7739 gnd.n6276 gnd.n2573 838.452
R7740 gnd.n3955 gnd.n2365 838.452
R7741 gnd.n3997 gnd.n2367 838.452
R7742 gnd.n7676 gnd.n167 783.196
R7743 gnd.n7536 gnd.n169 783.196
R7744 gnd.n5719 gnd.n3057 783.196
R7745 gnd.n6000 gnd.n3061 783.196
R7746 gnd.n6358 gnd.n2570 783.196
R7747 gnd.n2780 gnd.n2572 783.196
R7748 gnd.n4209 gnd.n2364 783.196
R7749 gnd.n6485 gnd.n2368 783.196
R7750 gnd.n6337 gnd.n2604 771.183
R7751 gnd.n6018 gnd.n3035 771.183
R7752 gnd.n6341 gnd.n2586 771.183
R7753 gnd.n5369 gnd.n3037 771.183
R7754 gnd.n2246 gnd.n878 766.379
R7755 gnd.n2249 gnd.n2248 766.379
R7756 gnd.n1486 gnd.n1389 766.379
R7757 gnd.n1482 gnd.n1387 766.379
R7758 gnd.n2337 gnd.n900 756.769
R7759 gnd.n2240 gnd.n2239 756.769
R7760 gnd.n1579 gnd.n1296 756.769
R7761 gnd.n1577 gnd.n1299 756.769
R7762 gnd.n6689 gnd.n706 737.549
R7763 gnd.n7210 gnd.n395 737.549
R7764 gnd.n7421 gnd.n267 737.549
R7765 gnd.n6513 gnd.n871 737.549
R7766 gnd.n6685 gnd.n706 585
R7767 gnd.n706 gnd.n705 585
R7768 gnd.n6684 gnd.n6683 585
R7769 gnd.n6683 gnd.n6682 585
R7770 gnd.n709 gnd.n708 585
R7771 gnd.n6681 gnd.n709 585
R7772 gnd.n6679 gnd.n6678 585
R7773 gnd.n6680 gnd.n6679 585
R7774 gnd.n6677 gnd.n711 585
R7775 gnd.n711 gnd.n710 585
R7776 gnd.n6676 gnd.n6675 585
R7777 gnd.n6675 gnd.n6674 585
R7778 gnd.n717 gnd.n716 585
R7779 gnd.n6673 gnd.n717 585
R7780 gnd.n6671 gnd.n6670 585
R7781 gnd.n6672 gnd.n6671 585
R7782 gnd.n6669 gnd.n719 585
R7783 gnd.n719 gnd.n718 585
R7784 gnd.n6668 gnd.n6667 585
R7785 gnd.n6667 gnd.n6666 585
R7786 gnd.n725 gnd.n724 585
R7787 gnd.n6665 gnd.n725 585
R7788 gnd.n6663 gnd.n6662 585
R7789 gnd.n6664 gnd.n6663 585
R7790 gnd.n6661 gnd.n727 585
R7791 gnd.n727 gnd.n726 585
R7792 gnd.n6660 gnd.n6659 585
R7793 gnd.n6659 gnd.n6658 585
R7794 gnd.n733 gnd.n732 585
R7795 gnd.n6657 gnd.n733 585
R7796 gnd.n6655 gnd.n6654 585
R7797 gnd.n6656 gnd.n6655 585
R7798 gnd.n6653 gnd.n735 585
R7799 gnd.n735 gnd.n734 585
R7800 gnd.n6652 gnd.n6651 585
R7801 gnd.n6651 gnd.n6650 585
R7802 gnd.n741 gnd.n740 585
R7803 gnd.n6649 gnd.n741 585
R7804 gnd.n6647 gnd.n6646 585
R7805 gnd.n6648 gnd.n6647 585
R7806 gnd.n6645 gnd.n743 585
R7807 gnd.n743 gnd.n742 585
R7808 gnd.n6644 gnd.n6643 585
R7809 gnd.n6643 gnd.n6642 585
R7810 gnd.n749 gnd.n748 585
R7811 gnd.n6641 gnd.n749 585
R7812 gnd.n6639 gnd.n6638 585
R7813 gnd.n6640 gnd.n6639 585
R7814 gnd.n6637 gnd.n751 585
R7815 gnd.n751 gnd.n750 585
R7816 gnd.n6636 gnd.n6635 585
R7817 gnd.n6635 gnd.n6634 585
R7818 gnd.n757 gnd.n756 585
R7819 gnd.n6633 gnd.n757 585
R7820 gnd.n6631 gnd.n6630 585
R7821 gnd.n6632 gnd.n6631 585
R7822 gnd.n6629 gnd.n759 585
R7823 gnd.n759 gnd.n758 585
R7824 gnd.n6628 gnd.n6627 585
R7825 gnd.n6627 gnd.n6626 585
R7826 gnd.n765 gnd.n764 585
R7827 gnd.n6625 gnd.n765 585
R7828 gnd.n6623 gnd.n6622 585
R7829 gnd.n6624 gnd.n6623 585
R7830 gnd.n6621 gnd.n767 585
R7831 gnd.n767 gnd.n766 585
R7832 gnd.n6620 gnd.n6619 585
R7833 gnd.n6619 gnd.n6618 585
R7834 gnd.n773 gnd.n772 585
R7835 gnd.n6617 gnd.n773 585
R7836 gnd.n6615 gnd.n6614 585
R7837 gnd.n6616 gnd.n6615 585
R7838 gnd.n6613 gnd.n775 585
R7839 gnd.n775 gnd.n774 585
R7840 gnd.n6612 gnd.n6611 585
R7841 gnd.n6611 gnd.n6610 585
R7842 gnd.n781 gnd.n780 585
R7843 gnd.n6609 gnd.n781 585
R7844 gnd.n6607 gnd.n6606 585
R7845 gnd.n6608 gnd.n6607 585
R7846 gnd.n6605 gnd.n783 585
R7847 gnd.n783 gnd.n782 585
R7848 gnd.n6604 gnd.n6603 585
R7849 gnd.n6603 gnd.n6602 585
R7850 gnd.n789 gnd.n788 585
R7851 gnd.n6601 gnd.n789 585
R7852 gnd.n6599 gnd.n6598 585
R7853 gnd.n6600 gnd.n6599 585
R7854 gnd.n6597 gnd.n791 585
R7855 gnd.n791 gnd.n790 585
R7856 gnd.n6596 gnd.n6595 585
R7857 gnd.n6595 gnd.n6594 585
R7858 gnd.n797 gnd.n796 585
R7859 gnd.n6593 gnd.n797 585
R7860 gnd.n6591 gnd.n6590 585
R7861 gnd.n6592 gnd.n6591 585
R7862 gnd.n6589 gnd.n799 585
R7863 gnd.n799 gnd.n798 585
R7864 gnd.n6588 gnd.n6587 585
R7865 gnd.n6587 gnd.n6586 585
R7866 gnd.n805 gnd.n804 585
R7867 gnd.n6585 gnd.n805 585
R7868 gnd.n6583 gnd.n6582 585
R7869 gnd.n6584 gnd.n6583 585
R7870 gnd.n6581 gnd.n807 585
R7871 gnd.n807 gnd.n806 585
R7872 gnd.n6580 gnd.n6579 585
R7873 gnd.n6579 gnd.n6578 585
R7874 gnd.n813 gnd.n812 585
R7875 gnd.n6577 gnd.n813 585
R7876 gnd.n6575 gnd.n6574 585
R7877 gnd.n6576 gnd.n6575 585
R7878 gnd.n6573 gnd.n815 585
R7879 gnd.n815 gnd.n814 585
R7880 gnd.n6572 gnd.n6571 585
R7881 gnd.n6571 gnd.n6570 585
R7882 gnd.n821 gnd.n820 585
R7883 gnd.n6569 gnd.n821 585
R7884 gnd.n6567 gnd.n6566 585
R7885 gnd.n6568 gnd.n6567 585
R7886 gnd.n6565 gnd.n823 585
R7887 gnd.n823 gnd.n822 585
R7888 gnd.n6564 gnd.n6563 585
R7889 gnd.n6563 gnd.n6562 585
R7890 gnd.n829 gnd.n828 585
R7891 gnd.n6561 gnd.n829 585
R7892 gnd.n6559 gnd.n6558 585
R7893 gnd.n6560 gnd.n6559 585
R7894 gnd.n6557 gnd.n831 585
R7895 gnd.n831 gnd.n830 585
R7896 gnd.n6556 gnd.n6555 585
R7897 gnd.n6555 gnd.n6554 585
R7898 gnd.n837 gnd.n836 585
R7899 gnd.n6553 gnd.n837 585
R7900 gnd.n6551 gnd.n6550 585
R7901 gnd.n6552 gnd.n6551 585
R7902 gnd.n6549 gnd.n839 585
R7903 gnd.n839 gnd.n838 585
R7904 gnd.n6548 gnd.n6547 585
R7905 gnd.n6547 gnd.n6546 585
R7906 gnd.n845 gnd.n844 585
R7907 gnd.n6545 gnd.n845 585
R7908 gnd.n6543 gnd.n6542 585
R7909 gnd.n6544 gnd.n6543 585
R7910 gnd.n6541 gnd.n847 585
R7911 gnd.n847 gnd.n846 585
R7912 gnd.n6540 gnd.n6539 585
R7913 gnd.n6539 gnd.n6538 585
R7914 gnd.n853 gnd.n852 585
R7915 gnd.n6537 gnd.n853 585
R7916 gnd.n6535 gnd.n6534 585
R7917 gnd.n6536 gnd.n6535 585
R7918 gnd.n6533 gnd.n855 585
R7919 gnd.n855 gnd.n854 585
R7920 gnd.n6532 gnd.n6531 585
R7921 gnd.n6531 gnd.n6530 585
R7922 gnd.n861 gnd.n860 585
R7923 gnd.n6529 gnd.n861 585
R7924 gnd.n6527 gnd.n6526 585
R7925 gnd.n6528 gnd.n6527 585
R7926 gnd.n6525 gnd.n863 585
R7927 gnd.n863 gnd.n862 585
R7928 gnd.n6524 gnd.n6523 585
R7929 gnd.n6523 gnd.n6522 585
R7930 gnd.n869 gnd.n868 585
R7931 gnd.n6521 gnd.n869 585
R7932 gnd.n6519 gnd.n6518 585
R7933 gnd.n6520 gnd.n6519 585
R7934 gnd.n6689 gnd.n6688 585
R7935 gnd.n6690 gnd.n6689 585
R7936 gnd.n704 gnd.n703 585
R7937 gnd.n6691 gnd.n704 585
R7938 gnd.n6694 gnd.n6693 585
R7939 gnd.n6693 gnd.n6692 585
R7940 gnd.n701 gnd.n700 585
R7941 gnd.n700 gnd.n699 585
R7942 gnd.n6699 gnd.n6698 585
R7943 gnd.n6700 gnd.n6699 585
R7944 gnd.n698 gnd.n697 585
R7945 gnd.n6701 gnd.n698 585
R7946 gnd.n6704 gnd.n6703 585
R7947 gnd.n6703 gnd.n6702 585
R7948 gnd.n695 gnd.n694 585
R7949 gnd.n694 gnd.n693 585
R7950 gnd.n6709 gnd.n6708 585
R7951 gnd.n6710 gnd.n6709 585
R7952 gnd.n692 gnd.n691 585
R7953 gnd.n6711 gnd.n692 585
R7954 gnd.n6714 gnd.n6713 585
R7955 gnd.n6713 gnd.n6712 585
R7956 gnd.n689 gnd.n688 585
R7957 gnd.n688 gnd.n687 585
R7958 gnd.n6719 gnd.n6718 585
R7959 gnd.n6720 gnd.n6719 585
R7960 gnd.n686 gnd.n685 585
R7961 gnd.n6721 gnd.n686 585
R7962 gnd.n6724 gnd.n6723 585
R7963 gnd.n6723 gnd.n6722 585
R7964 gnd.n683 gnd.n682 585
R7965 gnd.n682 gnd.n681 585
R7966 gnd.n6729 gnd.n6728 585
R7967 gnd.n6730 gnd.n6729 585
R7968 gnd.n680 gnd.n679 585
R7969 gnd.n6731 gnd.n680 585
R7970 gnd.n6734 gnd.n6733 585
R7971 gnd.n6733 gnd.n6732 585
R7972 gnd.n677 gnd.n676 585
R7973 gnd.n676 gnd.n675 585
R7974 gnd.n6739 gnd.n6738 585
R7975 gnd.n6740 gnd.n6739 585
R7976 gnd.n674 gnd.n673 585
R7977 gnd.n6741 gnd.n674 585
R7978 gnd.n6744 gnd.n6743 585
R7979 gnd.n6743 gnd.n6742 585
R7980 gnd.n671 gnd.n670 585
R7981 gnd.n670 gnd.n669 585
R7982 gnd.n6749 gnd.n6748 585
R7983 gnd.n6750 gnd.n6749 585
R7984 gnd.n668 gnd.n667 585
R7985 gnd.n6751 gnd.n668 585
R7986 gnd.n6754 gnd.n6753 585
R7987 gnd.n6753 gnd.n6752 585
R7988 gnd.n665 gnd.n664 585
R7989 gnd.n664 gnd.n663 585
R7990 gnd.n6759 gnd.n6758 585
R7991 gnd.n6760 gnd.n6759 585
R7992 gnd.n662 gnd.n661 585
R7993 gnd.n6761 gnd.n662 585
R7994 gnd.n6764 gnd.n6763 585
R7995 gnd.n6763 gnd.n6762 585
R7996 gnd.n659 gnd.n658 585
R7997 gnd.n658 gnd.n657 585
R7998 gnd.n6769 gnd.n6768 585
R7999 gnd.n6770 gnd.n6769 585
R8000 gnd.n656 gnd.n655 585
R8001 gnd.n6771 gnd.n656 585
R8002 gnd.n6774 gnd.n6773 585
R8003 gnd.n6773 gnd.n6772 585
R8004 gnd.n653 gnd.n652 585
R8005 gnd.n652 gnd.n651 585
R8006 gnd.n6779 gnd.n6778 585
R8007 gnd.n6780 gnd.n6779 585
R8008 gnd.n650 gnd.n649 585
R8009 gnd.n6781 gnd.n650 585
R8010 gnd.n6784 gnd.n6783 585
R8011 gnd.n6783 gnd.n6782 585
R8012 gnd.n647 gnd.n646 585
R8013 gnd.n646 gnd.n645 585
R8014 gnd.n6789 gnd.n6788 585
R8015 gnd.n6790 gnd.n6789 585
R8016 gnd.n644 gnd.n643 585
R8017 gnd.n6791 gnd.n644 585
R8018 gnd.n6794 gnd.n6793 585
R8019 gnd.n6793 gnd.n6792 585
R8020 gnd.n641 gnd.n640 585
R8021 gnd.n640 gnd.n639 585
R8022 gnd.n6799 gnd.n6798 585
R8023 gnd.n6800 gnd.n6799 585
R8024 gnd.n638 gnd.n637 585
R8025 gnd.n6801 gnd.n638 585
R8026 gnd.n6804 gnd.n6803 585
R8027 gnd.n6803 gnd.n6802 585
R8028 gnd.n635 gnd.n634 585
R8029 gnd.n634 gnd.n633 585
R8030 gnd.n6809 gnd.n6808 585
R8031 gnd.n6810 gnd.n6809 585
R8032 gnd.n632 gnd.n631 585
R8033 gnd.n6811 gnd.n632 585
R8034 gnd.n6814 gnd.n6813 585
R8035 gnd.n6813 gnd.n6812 585
R8036 gnd.n629 gnd.n628 585
R8037 gnd.n628 gnd.n627 585
R8038 gnd.n6819 gnd.n6818 585
R8039 gnd.n6820 gnd.n6819 585
R8040 gnd.n626 gnd.n625 585
R8041 gnd.n6821 gnd.n626 585
R8042 gnd.n6824 gnd.n6823 585
R8043 gnd.n6823 gnd.n6822 585
R8044 gnd.n623 gnd.n622 585
R8045 gnd.n622 gnd.n621 585
R8046 gnd.n6829 gnd.n6828 585
R8047 gnd.n6830 gnd.n6829 585
R8048 gnd.n620 gnd.n619 585
R8049 gnd.n6831 gnd.n620 585
R8050 gnd.n6834 gnd.n6833 585
R8051 gnd.n6833 gnd.n6832 585
R8052 gnd.n617 gnd.n616 585
R8053 gnd.n616 gnd.n615 585
R8054 gnd.n6839 gnd.n6838 585
R8055 gnd.n6840 gnd.n6839 585
R8056 gnd.n614 gnd.n613 585
R8057 gnd.n6841 gnd.n614 585
R8058 gnd.n6844 gnd.n6843 585
R8059 gnd.n6843 gnd.n6842 585
R8060 gnd.n611 gnd.n610 585
R8061 gnd.n610 gnd.n609 585
R8062 gnd.n6849 gnd.n6848 585
R8063 gnd.n6850 gnd.n6849 585
R8064 gnd.n608 gnd.n607 585
R8065 gnd.n6851 gnd.n608 585
R8066 gnd.n6854 gnd.n6853 585
R8067 gnd.n6853 gnd.n6852 585
R8068 gnd.n605 gnd.n604 585
R8069 gnd.n604 gnd.n603 585
R8070 gnd.n6859 gnd.n6858 585
R8071 gnd.n6860 gnd.n6859 585
R8072 gnd.n602 gnd.n601 585
R8073 gnd.n6861 gnd.n602 585
R8074 gnd.n6864 gnd.n6863 585
R8075 gnd.n6863 gnd.n6862 585
R8076 gnd.n599 gnd.n598 585
R8077 gnd.n598 gnd.n597 585
R8078 gnd.n6869 gnd.n6868 585
R8079 gnd.n6870 gnd.n6869 585
R8080 gnd.n596 gnd.n595 585
R8081 gnd.n6871 gnd.n596 585
R8082 gnd.n6874 gnd.n6873 585
R8083 gnd.n6873 gnd.n6872 585
R8084 gnd.n593 gnd.n592 585
R8085 gnd.n592 gnd.n591 585
R8086 gnd.n6879 gnd.n6878 585
R8087 gnd.n6880 gnd.n6879 585
R8088 gnd.n590 gnd.n589 585
R8089 gnd.n6881 gnd.n590 585
R8090 gnd.n6884 gnd.n6883 585
R8091 gnd.n6883 gnd.n6882 585
R8092 gnd.n587 gnd.n586 585
R8093 gnd.n586 gnd.n585 585
R8094 gnd.n6889 gnd.n6888 585
R8095 gnd.n6890 gnd.n6889 585
R8096 gnd.n584 gnd.n583 585
R8097 gnd.n6891 gnd.n584 585
R8098 gnd.n6894 gnd.n6893 585
R8099 gnd.n6893 gnd.n6892 585
R8100 gnd.n581 gnd.n580 585
R8101 gnd.n580 gnd.n579 585
R8102 gnd.n6899 gnd.n6898 585
R8103 gnd.n6900 gnd.n6899 585
R8104 gnd.n578 gnd.n577 585
R8105 gnd.n6901 gnd.n578 585
R8106 gnd.n6904 gnd.n6903 585
R8107 gnd.n6903 gnd.n6902 585
R8108 gnd.n575 gnd.n574 585
R8109 gnd.n574 gnd.n573 585
R8110 gnd.n6909 gnd.n6908 585
R8111 gnd.n6910 gnd.n6909 585
R8112 gnd.n572 gnd.n571 585
R8113 gnd.n6911 gnd.n572 585
R8114 gnd.n6914 gnd.n6913 585
R8115 gnd.n6913 gnd.n6912 585
R8116 gnd.n569 gnd.n568 585
R8117 gnd.n568 gnd.n567 585
R8118 gnd.n6919 gnd.n6918 585
R8119 gnd.n6920 gnd.n6919 585
R8120 gnd.n566 gnd.n565 585
R8121 gnd.n6921 gnd.n566 585
R8122 gnd.n6924 gnd.n6923 585
R8123 gnd.n6923 gnd.n6922 585
R8124 gnd.n563 gnd.n562 585
R8125 gnd.n562 gnd.n561 585
R8126 gnd.n6929 gnd.n6928 585
R8127 gnd.n6930 gnd.n6929 585
R8128 gnd.n560 gnd.n559 585
R8129 gnd.n6931 gnd.n560 585
R8130 gnd.n6934 gnd.n6933 585
R8131 gnd.n6933 gnd.n6932 585
R8132 gnd.n557 gnd.n556 585
R8133 gnd.n556 gnd.n555 585
R8134 gnd.n6939 gnd.n6938 585
R8135 gnd.n6940 gnd.n6939 585
R8136 gnd.n554 gnd.n553 585
R8137 gnd.n6941 gnd.n554 585
R8138 gnd.n6944 gnd.n6943 585
R8139 gnd.n6943 gnd.n6942 585
R8140 gnd.n551 gnd.n550 585
R8141 gnd.n550 gnd.n549 585
R8142 gnd.n6949 gnd.n6948 585
R8143 gnd.n6950 gnd.n6949 585
R8144 gnd.n548 gnd.n547 585
R8145 gnd.n6951 gnd.n548 585
R8146 gnd.n6954 gnd.n6953 585
R8147 gnd.n6953 gnd.n6952 585
R8148 gnd.n545 gnd.n544 585
R8149 gnd.n544 gnd.n543 585
R8150 gnd.n6959 gnd.n6958 585
R8151 gnd.n6960 gnd.n6959 585
R8152 gnd.n542 gnd.n541 585
R8153 gnd.n6961 gnd.n542 585
R8154 gnd.n6964 gnd.n6963 585
R8155 gnd.n6963 gnd.n6962 585
R8156 gnd.n539 gnd.n538 585
R8157 gnd.n538 gnd.n537 585
R8158 gnd.n6969 gnd.n6968 585
R8159 gnd.n6970 gnd.n6969 585
R8160 gnd.n536 gnd.n535 585
R8161 gnd.n6971 gnd.n536 585
R8162 gnd.n6974 gnd.n6973 585
R8163 gnd.n6973 gnd.n6972 585
R8164 gnd.n533 gnd.n532 585
R8165 gnd.n532 gnd.n531 585
R8166 gnd.n6979 gnd.n6978 585
R8167 gnd.n6980 gnd.n6979 585
R8168 gnd.n530 gnd.n529 585
R8169 gnd.n6981 gnd.n530 585
R8170 gnd.n6984 gnd.n6983 585
R8171 gnd.n6983 gnd.n6982 585
R8172 gnd.n527 gnd.n526 585
R8173 gnd.n526 gnd.n525 585
R8174 gnd.n6989 gnd.n6988 585
R8175 gnd.n6990 gnd.n6989 585
R8176 gnd.n524 gnd.n523 585
R8177 gnd.n6991 gnd.n524 585
R8178 gnd.n6994 gnd.n6993 585
R8179 gnd.n6993 gnd.n6992 585
R8180 gnd.n521 gnd.n520 585
R8181 gnd.n520 gnd.n519 585
R8182 gnd.n6999 gnd.n6998 585
R8183 gnd.n7000 gnd.n6999 585
R8184 gnd.n518 gnd.n517 585
R8185 gnd.n7001 gnd.n518 585
R8186 gnd.n7004 gnd.n7003 585
R8187 gnd.n7003 gnd.n7002 585
R8188 gnd.n515 gnd.n514 585
R8189 gnd.n514 gnd.n513 585
R8190 gnd.n7009 gnd.n7008 585
R8191 gnd.n7010 gnd.n7009 585
R8192 gnd.n512 gnd.n511 585
R8193 gnd.n7011 gnd.n512 585
R8194 gnd.n7014 gnd.n7013 585
R8195 gnd.n7013 gnd.n7012 585
R8196 gnd.n509 gnd.n508 585
R8197 gnd.n508 gnd.n507 585
R8198 gnd.n7019 gnd.n7018 585
R8199 gnd.n7020 gnd.n7019 585
R8200 gnd.n506 gnd.n505 585
R8201 gnd.n7021 gnd.n506 585
R8202 gnd.n7024 gnd.n7023 585
R8203 gnd.n7023 gnd.n7022 585
R8204 gnd.n503 gnd.n502 585
R8205 gnd.n502 gnd.n501 585
R8206 gnd.n7029 gnd.n7028 585
R8207 gnd.n7030 gnd.n7029 585
R8208 gnd.n500 gnd.n499 585
R8209 gnd.n7031 gnd.n500 585
R8210 gnd.n7034 gnd.n7033 585
R8211 gnd.n7033 gnd.n7032 585
R8212 gnd.n497 gnd.n496 585
R8213 gnd.n496 gnd.n495 585
R8214 gnd.n7039 gnd.n7038 585
R8215 gnd.n7040 gnd.n7039 585
R8216 gnd.n494 gnd.n493 585
R8217 gnd.n7041 gnd.n494 585
R8218 gnd.n7044 gnd.n7043 585
R8219 gnd.n7043 gnd.n7042 585
R8220 gnd.n491 gnd.n490 585
R8221 gnd.n490 gnd.n489 585
R8222 gnd.n7049 gnd.n7048 585
R8223 gnd.n7050 gnd.n7049 585
R8224 gnd.n488 gnd.n487 585
R8225 gnd.n7051 gnd.n488 585
R8226 gnd.n7054 gnd.n7053 585
R8227 gnd.n7053 gnd.n7052 585
R8228 gnd.n485 gnd.n484 585
R8229 gnd.n484 gnd.n483 585
R8230 gnd.n7059 gnd.n7058 585
R8231 gnd.n7060 gnd.n7059 585
R8232 gnd.n482 gnd.n481 585
R8233 gnd.n7061 gnd.n482 585
R8234 gnd.n7064 gnd.n7063 585
R8235 gnd.n7063 gnd.n7062 585
R8236 gnd.n479 gnd.n478 585
R8237 gnd.n478 gnd.n477 585
R8238 gnd.n7069 gnd.n7068 585
R8239 gnd.n7070 gnd.n7069 585
R8240 gnd.n476 gnd.n475 585
R8241 gnd.n7071 gnd.n476 585
R8242 gnd.n7074 gnd.n7073 585
R8243 gnd.n7073 gnd.n7072 585
R8244 gnd.n473 gnd.n472 585
R8245 gnd.n472 gnd.n471 585
R8246 gnd.n7079 gnd.n7078 585
R8247 gnd.n7080 gnd.n7079 585
R8248 gnd.n470 gnd.n469 585
R8249 gnd.n7081 gnd.n470 585
R8250 gnd.n7084 gnd.n7083 585
R8251 gnd.n7083 gnd.n7082 585
R8252 gnd.n467 gnd.n466 585
R8253 gnd.n466 gnd.n465 585
R8254 gnd.n7089 gnd.n7088 585
R8255 gnd.n7090 gnd.n7089 585
R8256 gnd.n464 gnd.n463 585
R8257 gnd.n7091 gnd.n464 585
R8258 gnd.n7094 gnd.n7093 585
R8259 gnd.n7093 gnd.n7092 585
R8260 gnd.n461 gnd.n460 585
R8261 gnd.n460 gnd.n459 585
R8262 gnd.n7099 gnd.n7098 585
R8263 gnd.n7100 gnd.n7099 585
R8264 gnd.n458 gnd.n457 585
R8265 gnd.n7101 gnd.n458 585
R8266 gnd.n7104 gnd.n7103 585
R8267 gnd.n7103 gnd.n7102 585
R8268 gnd.n455 gnd.n454 585
R8269 gnd.n454 gnd.n453 585
R8270 gnd.n7109 gnd.n7108 585
R8271 gnd.n7110 gnd.n7109 585
R8272 gnd.n452 gnd.n451 585
R8273 gnd.n7111 gnd.n452 585
R8274 gnd.n7114 gnd.n7113 585
R8275 gnd.n7113 gnd.n7112 585
R8276 gnd.n449 gnd.n448 585
R8277 gnd.n448 gnd.n447 585
R8278 gnd.n7119 gnd.n7118 585
R8279 gnd.n7120 gnd.n7119 585
R8280 gnd.n446 gnd.n445 585
R8281 gnd.n7121 gnd.n446 585
R8282 gnd.n7124 gnd.n7123 585
R8283 gnd.n7123 gnd.n7122 585
R8284 gnd.n443 gnd.n442 585
R8285 gnd.n442 gnd.n441 585
R8286 gnd.n7129 gnd.n7128 585
R8287 gnd.n7130 gnd.n7129 585
R8288 gnd.n440 gnd.n439 585
R8289 gnd.n7131 gnd.n440 585
R8290 gnd.n7134 gnd.n7133 585
R8291 gnd.n7133 gnd.n7132 585
R8292 gnd.n437 gnd.n436 585
R8293 gnd.n436 gnd.n435 585
R8294 gnd.n7139 gnd.n7138 585
R8295 gnd.n7140 gnd.n7139 585
R8296 gnd.n434 gnd.n433 585
R8297 gnd.n7141 gnd.n434 585
R8298 gnd.n7144 gnd.n7143 585
R8299 gnd.n7143 gnd.n7142 585
R8300 gnd.n431 gnd.n430 585
R8301 gnd.n430 gnd.n429 585
R8302 gnd.n7149 gnd.n7148 585
R8303 gnd.n7150 gnd.n7149 585
R8304 gnd.n428 gnd.n427 585
R8305 gnd.n7151 gnd.n428 585
R8306 gnd.n7154 gnd.n7153 585
R8307 gnd.n7153 gnd.n7152 585
R8308 gnd.n425 gnd.n424 585
R8309 gnd.n424 gnd.n423 585
R8310 gnd.n7159 gnd.n7158 585
R8311 gnd.n7160 gnd.n7159 585
R8312 gnd.n422 gnd.n421 585
R8313 gnd.n7161 gnd.n422 585
R8314 gnd.n7164 gnd.n7163 585
R8315 gnd.n7163 gnd.n7162 585
R8316 gnd.n419 gnd.n418 585
R8317 gnd.n418 gnd.n417 585
R8318 gnd.n7169 gnd.n7168 585
R8319 gnd.n7170 gnd.n7169 585
R8320 gnd.n416 gnd.n415 585
R8321 gnd.n7171 gnd.n416 585
R8322 gnd.n7174 gnd.n7173 585
R8323 gnd.n7173 gnd.n7172 585
R8324 gnd.n413 gnd.n412 585
R8325 gnd.n412 gnd.n411 585
R8326 gnd.n7179 gnd.n7178 585
R8327 gnd.n7180 gnd.n7179 585
R8328 gnd.n410 gnd.n409 585
R8329 gnd.n7181 gnd.n410 585
R8330 gnd.n7184 gnd.n7183 585
R8331 gnd.n7183 gnd.n7182 585
R8332 gnd.n407 gnd.n406 585
R8333 gnd.n406 gnd.n405 585
R8334 gnd.n7189 gnd.n7188 585
R8335 gnd.n7190 gnd.n7189 585
R8336 gnd.n404 gnd.n403 585
R8337 gnd.n7191 gnd.n404 585
R8338 gnd.n7194 gnd.n7193 585
R8339 gnd.n7193 gnd.n7192 585
R8340 gnd.n401 gnd.n400 585
R8341 gnd.n400 gnd.n399 585
R8342 gnd.n7200 gnd.n7199 585
R8343 gnd.n7201 gnd.n7200 585
R8344 gnd.n398 gnd.n397 585
R8345 gnd.n7202 gnd.n398 585
R8346 gnd.n7205 gnd.n7204 585
R8347 gnd.n7204 gnd.n7203 585
R8348 gnd.n7206 gnd.n395 585
R8349 gnd.n395 gnd.n394 585
R8350 gnd.n270 gnd.n269 585
R8351 gnd.n269 gnd.n268 585
R8352 gnd.n7415 gnd.n7414 585
R8353 gnd.n7414 gnd.n7413 585
R8354 gnd.n273 gnd.n272 585
R8355 gnd.n7412 gnd.n273 585
R8356 gnd.n7410 gnd.n7409 585
R8357 gnd.n7411 gnd.n7410 585
R8358 gnd.n276 gnd.n275 585
R8359 gnd.n275 gnd.n274 585
R8360 gnd.n7405 gnd.n7404 585
R8361 gnd.n7404 gnd.n7403 585
R8362 gnd.n279 gnd.n278 585
R8363 gnd.n7402 gnd.n279 585
R8364 gnd.n7400 gnd.n7399 585
R8365 gnd.n7401 gnd.n7400 585
R8366 gnd.n282 gnd.n281 585
R8367 gnd.n281 gnd.n280 585
R8368 gnd.n7395 gnd.n7394 585
R8369 gnd.n7394 gnd.n7393 585
R8370 gnd.n285 gnd.n284 585
R8371 gnd.n7392 gnd.n285 585
R8372 gnd.n7390 gnd.n7389 585
R8373 gnd.n7391 gnd.n7390 585
R8374 gnd.n288 gnd.n287 585
R8375 gnd.n287 gnd.n286 585
R8376 gnd.n7385 gnd.n7384 585
R8377 gnd.n7384 gnd.n7383 585
R8378 gnd.n291 gnd.n290 585
R8379 gnd.n7382 gnd.n291 585
R8380 gnd.n7380 gnd.n7379 585
R8381 gnd.n7381 gnd.n7380 585
R8382 gnd.n294 gnd.n293 585
R8383 gnd.n293 gnd.n292 585
R8384 gnd.n7375 gnd.n7374 585
R8385 gnd.n7374 gnd.n7373 585
R8386 gnd.n297 gnd.n296 585
R8387 gnd.n7372 gnd.n297 585
R8388 gnd.n7370 gnd.n7369 585
R8389 gnd.n7371 gnd.n7370 585
R8390 gnd.n300 gnd.n299 585
R8391 gnd.n299 gnd.n298 585
R8392 gnd.n7365 gnd.n7364 585
R8393 gnd.n7364 gnd.n7363 585
R8394 gnd.n303 gnd.n302 585
R8395 gnd.n7362 gnd.n303 585
R8396 gnd.n7360 gnd.n7359 585
R8397 gnd.n7361 gnd.n7360 585
R8398 gnd.n306 gnd.n305 585
R8399 gnd.n305 gnd.n304 585
R8400 gnd.n7355 gnd.n7354 585
R8401 gnd.n7354 gnd.n7353 585
R8402 gnd.n309 gnd.n308 585
R8403 gnd.n7352 gnd.n309 585
R8404 gnd.n7350 gnd.n7349 585
R8405 gnd.n7351 gnd.n7350 585
R8406 gnd.n312 gnd.n311 585
R8407 gnd.n311 gnd.n310 585
R8408 gnd.n7345 gnd.n7344 585
R8409 gnd.n7344 gnd.n7343 585
R8410 gnd.n315 gnd.n314 585
R8411 gnd.n7342 gnd.n315 585
R8412 gnd.n7340 gnd.n7339 585
R8413 gnd.n7341 gnd.n7340 585
R8414 gnd.n318 gnd.n317 585
R8415 gnd.n317 gnd.n316 585
R8416 gnd.n7335 gnd.n7334 585
R8417 gnd.n7334 gnd.n7333 585
R8418 gnd.n321 gnd.n320 585
R8419 gnd.n7332 gnd.n321 585
R8420 gnd.n7330 gnd.n7329 585
R8421 gnd.n7331 gnd.n7330 585
R8422 gnd.n324 gnd.n323 585
R8423 gnd.n323 gnd.n322 585
R8424 gnd.n7325 gnd.n7324 585
R8425 gnd.n7324 gnd.n7323 585
R8426 gnd.n327 gnd.n326 585
R8427 gnd.n7322 gnd.n327 585
R8428 gnd.n7320 gnd.n7319 585
R8429 gnd.n7321 gnd.n7320 585
R8430 gnd.n330 gnd.n329 585
R8431 gnd.n329 gnd.n328 585
R8432 gnd.n7315 gnd.n7314 585
R8433 gnd.n7314 gnd.n7313 585
R8434 gnd.n333 gnd.n332 585
R8435 gnd.n7312 gnd.n333 585
R8436 gnd.n7310 gnd.n7309 585
R8437 gnd.n7311 gnd.n7310 585
R8438 gnd.n336 gnd.n335 585
R8439 gnd.n335 gnd.n334 585
R8440 gnd.n7305 gnd.n7304 585
R8441 gnd.n7304 gnd.n7303 585
R8442 gnd.n339 gnd.n338 585
R8443 gnd.n7302 gnd.n339 585
R8444 gnd.n7300 gnd.n7299 585
R8445 gnd.n7301 gnd.n7300 585
R8446 gnd.n342 gnd.n341 585
R8447 gnd.n341 gnd.n340 585
R8448 gnd.n7295 gnd.n7294 585
R8449 gnd.n7294 gnd.n7293 585
R8450 gnd.n345 gnd.n344 585
R8451 gnd.n7292 gnd.n345 585
R8452 gnd.n7290 gnd.n7289 585
R8453 gnd.n7291 gnd.n7290 585
R8454 gnd.n348 gnd.n347 585
R8455 gnd.n347 gnd.n346 585
R8456 gnd.n7285 gnd.n7284 585
R8457 gnd.n7284 gnd.n7283 585
R8458 gnd.n351 gnd.n350 585
R8459 gnd.n7282 gnd.n351 585
R8460 gnd.n7280 gnd.n7279 585
R8461 gnd.n7281 gnd.n7280 585
R8462 gnd.n354 gnd.n353 585
R8463 gnd.n353 gnd.n352 585
R8464 gnd.n7275 gnd.n7274 585
R8465 gnd.n7274 gnd.n7273 585
R8466 gnd.n357 gnd.n356 585
R8467 gnd.n7272 gnd.n357 585
R8468 gnd.n7270 gnd.n7269 585
R8469 gnd.n7271 gnd.n7270 585
R8470 gnd.n360 gnd.n359 585
R8471 gnd.n359 gnd.n358 585
R8472 gnd.n7265 gnd.n7264 585
R8473 gnd.n7264 gnd.n7263 585
R8474 gnd.n363 gnd.n362 585
R8475 gnd.n7262 gnd.n363 585
R8476 gnd.n7260 gnd.n7259 585
R8477 gnd.n7261 gnd.n7260 585
R8478 gnd.n366 gnd.n365 585
R8479 gnd.n365 gnd.n364 585
R8480 gnd.n7255 gnd.n7254 585
R8481 gnd.n7254 gnd.n7253 585
R8482 gnd.n369 gnd.n368 585
R8483 gnd.n7252 gnd.n369 585
R8484 gnd.n7250 gnd.n7249 585
R8485 gnd.n7251 gnd.n7250 585
R8486 gnd.n372 gnd.n371 585
R8487 gnd.n371 gnd.n370 585
R8488 gnd.n7245 gnd.n7244 585
R8489 gnd.n7244 gnd.n7243 585
R8490 gnd.n375 gnd.n374 585
R8491 gnd.n7242 gnd.n375 585
R8492 gnd.n7240 gnd.n7239 585
R8493 gnd.n7241 gnd.n7240 585
R8494 gnd.n378 gnd.n377 585
R8495 gnd.n377 gnd.n376 585
R8496 gnd.n7235 gnd.n7234 585
R8497 gnd.n7234 gnd.n7233 585
R8498 gnd.n381 gnd.n380 585
R8499 gnd.n7232 gnd.n381 585
R8500 gnd.n7230 gnd.n7229 585
R8501 gnd.n7231 gnd.n7230 585
R8502 gnd.n384 gnd.n383 585
R8503 gnd.n383 gnd.n382 585
R8504 gnd.n7225 gnd.n7224 585
R8505 gnd.n7224 gnd.n7223 585
R8506 gnd.n387 gnd.n386 585
R8507 gnd.n7222 gnd.n387 585
R8508 gnd.n7220 gnd.n7219 585
R8509 gnd.n7221 gnd.n7220 585
R8510 gnd.n390 gnd.n389 585
R8511 gnd.n389 gnd.n388 585
R8512 gnd.n7215 gnd.n7214 585
R8513 gnd.n7214 gnd.n7213 585
R8514 gnd.n393 gnd.n392 585
R8515 gnd.n7212 gnd.n393 585
R8516 gnd.n7210 gnd.n7209 585
R8517 gnd.n7211 gnd.n7210 585
R8518 gnd.n6356 gnd.n6355 585
R8519 gnd.n6357 gnd.n6356 585
R8520 gnd.n2560 gnd.n2559 585
R8521 gnd.n6350 gnd.n2560 585
R8522 gnd.n6365 gnd.n6364 585
R8523 gnd.n6364 gnd.n6363 585
R8524 gnd.n6366 gnd.n2555 585
R8525 gnd.n4425 gnd.n2555 585
R8526 gnd.n6368 gnd.n6367 585
R8527 gnd.n6369 gnd.n6368 585
R8528 gnd.n2540 gnd.n2539 585
R8529 gnd.n4419 gnd.n2540 585
R8530 gnd.n6377 gnd.n6376 585
R8531 gnd.n6376 gnd.n6375 585
R8532 gnd.n6378 gnd.n2535 585
R8533 gnd.n4436 gnd.n2535 585
R8534 gnd.n6380 gnd.n6379 585
R8535 gnd.n6381 gnd.n6380 585
R8536 gnd.n2519 gnd.n2518 585
R8537 gnd.n4412 gnd.n2519 585
R8538 gnd.n6389 gnd.n6388 585
R8539 gnd.n6388 gnd.n6387 585
R8540 gnd.n6390 gnd.n2514 585
R8541 gnd.n4404 gnd.n2514 585
R8542 gnd.n6392 gnd.n6391 585
R8543 gnd.n6393 gnd.n6392 585
R8544 gnd.n2500 gnd.n2499 585
R8545 gnd.n4398 gnd.n2500 585
R8546 gnd.n6401 gnd.n6400 585
R8547 gnd.n6400 gnd.n6399 585
R8548 gnd.n6402 gnd.n2495 585
R8549 gnd.n4390 gnd.n2495 585
R8550 gnd.n6404 gnd.n6403 585
R8551 gnd.n6405 gnd.n6404 585
R8552 gnd.n2482 gnd.n2481 585
R8553 gnd.n4341 gnd.n2482 585
R8554 gnd.n6414 gnd.n6413 585
R8555 gnd.n6413 gnd.n6412 585
R8556 gnd.n6415 gnd.n2477 585
R8557 gnd.n4332 gnd.n2477 585
R8558 gnd.n6417 gnd.n6416 585
R8559 gnd.n6418 gnd.n6417 585
R8560 gnd.n2466 gnd.n2465 585
R8561 gnd.n4317 gnd.n2466 585
R8562 gnd.n6427 gnd.n6426 585
R8563 gnd.n6426 gnd.n6425 585
R8564 gnd.n6428 gnd.n2461 585
R8565 gnd.n4354 gnd.n2461 585
R8566 gnd.n6430 gnd.n6429 585
R8567 gnd.n6431 gnd.n6430 585
R8568 gnd.n2447 gnd.n2446 585
R8569 gnd.n4310 gnd.n2447 585
R8570 gnd.n6440 gnd.n6439 585
R8571 gnd.n6439 gnd.n6438 585
R8572 gnd.n6441 gnd.n2442 585
R8573 gnd.n4301 gnd.n2442 585
R8574 gnd.n6443 gnd.n6442 585
R8575 gnd.n6444 gnd.n6443 585
R8576 gnd.n2427 gnd.n2426 585
R8577 gnd.n4295 gnd.n2427 585
R8578 gnd.n6452 gnd.n6451 585
R8579 gnd.n6451 gnd.n6450 585
R8580 gnd.n6453 gnd.n2422 585
R8581 gnd.n4287 gnd.n2422 585
R8582 gnd.n6455 gnd.n6454 585
R8583 gnd.n6456 gnd.n6455 585
R8584 gnd.n2406 gnd.n2405 585
R8585 gnd.n4232 gnd.n2406 585
R8586 gnd.n6464 gnd.n6463 585
R8587 gnd.n6463 gnd.n6462 585
R8588 gnd.n6465 gnd.n2401 585
R8589 gnd.n4238 gnd.n2401 585
R8590 gnd.n6467 gnd.n6466 585
R8591 gnd.n6468 gnd.n6467 585
R8592 gnd.n2385 gnd.n2384 585
R8593 gnd.n4244 gnd.n2385 585
R8594 gnd.n6476 gnd.n6475 585
R8595 gnd.n6475 gnd.n6474 585
R8596 gnd.n6477 gnd.n2379 585
R8597 gnd.n4250 gnd.n2379 585
R8598 gnd.n6479 gnd.n6478 585
R8599 gnd.n6480 gnd.n6479 585
R8600 gnd.n2380 gnd.n2378 585
R8601 gnd.n4256 gnd.n2378 585
R8602 gnd.n4213 gnd.n2367 585
R8603 gnd.n6486 gnd.n2367 585
R8604 gnd.n3998 gnd.n3997 585
R8605 gnd.n3995 gnd.n3932 585
R8606 gnd.n3994 gnd.n3993 585
R8607 gnd.n3992 gnd.n3991 585
R8608 gnd.n3990 gnd.n3936 585
R8609 gnd.n3988 gnd.n3987 585
R8610 gnd.n3986 gnd.n3937 585
R8611 gnd.n3985 gnd.n3984 585
R8612 gnd.n3982 gnd.n3942 585
R8613 gnd.n3980 gnd.n3979 585
R8614 gnd.n3978 gnd.n3943 585
R8615 gnd.n3977 gnd.n3976 585
R8616 gnd.n3974 gnd.n3948 585
R8617 gnd.n3972 gnd.n3971 585
R8618 gnd.n3970 gnd.n3949 585
R8619 gnd.n3969 gnd.n3968 585
R8620 gnd.n3966 gnd.n3954 585
R8621 gnd.n3964 gnd.n3963 585
R8622 gnd.n3956 gnd.n3955 585
R8623 gnd.n3955 gnd.n2363 585
R8624 gnd.n6277 gnd.n6276 585
R8625 gnd.n6278 gnd.n2675 585
R8626 gnd.n6279 gnd.n2670 585
R8627 gnd.n2688 gnd.n2659 585
R8628 gnd.n6286 gnd.n2658 585
R8629 gnd.n6287 gnd.n2657 585
R8630 gnd.n2685 gnd.n2651 585
R8631 gnd.n6294 gnd.n2650 585
R8632 gnd.n6295 gnd.n2649 585
R8633 gnd.n2683 gnd.n2641 585
R8634 gnd.n6302 gnd.n2640 585
R8635 gnd.n6303 gnd.n2639 585
R8636 gnd.n2680 gnd.n2633 585
R8637 gnd.n6310 gnd.n2632 585
R8638 gnd.n6311 gnd.n2631 585
R8639 gnd.n2678 gnd.n2623 585
R8640 gnd.n6318 gnd.n2622 585
R8641 gnd.n6319 gnd.n2621 585
R8642 gnd.n2620 gnd.n2575 585
R8643 gnd.n6274 gnd.n2575 585
R8644 gnd.n2580 gnd.n2573 585
R8645 gnd.n6357 gnd.n2573 585
R8646 gnd.n6349 gnd.n6348 585
R8647 gnd.n6350 gnd.n6349 585
R8648 gnd.n2579 gnd.n2563 585
R8649 gnd.n6363 gnd.n2563 585
R8650 gnd.n4428 gnd.n4426 585
R8651 gnd.n4426 gnd.n4425 585
R8652 gnd.n4429 gnd.n2553 585
R8653 gnd.n6369 gnd.n2553 585
R8654 gnd.n4430 gnd.n3862 585
R8655 gnd.n4419 gnd.n3862 585
R8656 gnd.n3859 gnd.n2542 585
R8657 gnd.n6375 gnd.n2542 585
R8658 gnd.n4435 gnd.n4434 585
R8659 gnd.n4436 gnd.n4435 585
R8660 gnd.n3858 gnd.n2533 585
R8661 gnd.n6381 gnd.n2533 585
R8662 gnd.n4411 gnd.n4410 585
R8663 gnd.n4412 gnd.n4411 585
R8664 gnd.n3865 gnd.n2522 585
R8665 gnd.n6387 gnd.n2522 585
R8666 gnd.n4406 gnd.n4405 585
R8667 gnd.n4405 gnd.n4404 585
R8668 gnd.n3867 gnd.n2513 585
R8669 gnd.n6393 gnd.n2513 585
R8670 gnd.n4397 gnd.n4396 585
R8671 gnd.n4398 gnd.n4397 585
R8672 gnd.n3871 gnd.n2502 585
R8673 gnd.n6399 gnd.n2502 585
R8674 gnd.n4392 gnd.n4391 585
R8675 gnd.n4391 gnd.n4390 585
R8676 gnd.n3873 gnd.n2493 585
R8677 gnd.n6405 gnd.n2493 585
R8678 gnd.n4344 gnd.n4342 585
R8679 gnd.n4342 gnd.n4341 585
R8680 gnd.n4345 gnd.n2485 585
R8681 gnd.n6412 gnd.n2485 585
R8682 gnd.n4346 gnd.n3897 585
R8683 gnd.n4332 gnd.n3897 585
R8684 gnd.n3895 gnd.n2476 585
R8685 gnd.n6418 gnd.n2476 585
R8686 gnd.n4350 gnd.n3894 585
R8687 gnd.n4317 gnd.n3894 585
R8688 gnd.n4351 gnd.n2468 585
R8689 gnd.n6425 gnd.n2468 585
R8690 gnd.n4353 gnd.n4352 585
R8691 gnd.n4354 gnd.n4353 585
R8692 gnd.n3891 gnd.n2459 585
R8693 gnd.n6431 gnd.n2459 585
R8694 gnd.n4309 gnd.n4308 585
R8695 gnd.n4310 gnd.n4309 585
R8696 gnd.n3900 gnd.n2450 585
R8697 gnd.n6438 gnd.n2450 585
R8698 gnd.n4303 gnd.n4302 585
R8699 gnd.n4302 gnd.n4301 585
R8700 gnd.n3902 gnd.n2440 585
R8701 gnd.n6444 gnd.n2440 585
R8702 gnd.n4294 gnd.n4293 585
R8703 gnd.n4295 gnd.n4294 585
R8704 gnd.n3905 gnd.n2429 585
R8705 gnd.n6450 gnd.n2429 585
R8706 gnd.n4289 gnd.n4288 585
R8707 gnd.n4288 gnd.n4287 585
R8708 gnd.n3907 gnd.n2420 585
R8709 gnd.n6456 gnd.n2420 585
R8710 gnd.n4231 gnd.n4230 585
R8711 gnd.n4232 gnd.n4231 585
R8712 gnd.n4224 gnd.n2409 585
R8713 gnd.n6462 gnd.n2409 585
R8714 gnd.n4240 gnd.n4239 585
R8715 gnd.n4239 gnd.n4238 585
R8716 gnd.n4241 gnd.n2399 585
R8717 gnd.n6468 gnd.n2399 585
R8718 gnd.n4243 gnd.n4242 585
R8719 gnd.n4244 gnd.n4243 585
R8720 gnd.n3929 gnd.n2388 585
R8721 gnd.n6474 gnd.n2388 585
R8722 gnd.n4252 gnd.n4251 585
R8723 gnd.n4251 gnd.n4250 585
R8724 gnd.n4253 gnd.n2376 585
R8725 gnd.n6480 gnd.n2376 585
R8726 gnd.n4255 gnd.n4254 585
R8727 gnd.n4256 gnd.n4255 585
R8728 gnd.n3925 gnd.n2365 585
R8729 gnd.n6486 gnd.n2365 585
R8730 gnd.n2246 gnd.n2245 585
R8731 gnd.n2247 gnd.n2246 585
R8732 gnd.n953 gnd.n952 585
R8733 gnd.n959 gnd.n952 585
R8734 gnd.n2221 gnd.n971 585
R8735 gnd.n971 gnd.n958 585
R8736 gnd.n2223 gnd.n2222 585
R8737 gnd.n2224 gnd.n2223 585
R8738 gnd.n972 gnd.n970 585
R8739 gnd.n970 gnd.n966 585
R8740 gnd.n1955 gnd.n1954 585
R8741 gnd.n1954 gnd.n1953 585
R8742 gnd.n977 gnd.n976 585
R8743 gnd.n1924 gnd.n977 585
R8744 gnd.n1944 gnd.n1943 585
R8745 gnd.n1943 gnd.n1942 585
R8746 gnd.n984 gnd.n983 585
R8747 gnd.n1930 gnd.n984 585
R8748 gnd.n1900 gnd.n1004 585
R8749 gnd.n1004 gnd.n1003 585
R8750 gnd.n1902 gnd.n1901 585
R8751 gnd.n1903 gnd.n1902 585
R8752 gnd.n1005 gnd.n1002 585
R8753 gnd.n1013 gnd.n1002 585
R8754 gnd.n1878 gnd.n1025 585
R8755 gnd.n1025 gnd.n1012 585
R8756 gnd.n1880 gnd.n1879 585
R8757 gnd.n1881 gnd.n1880 585
R8758 gnd.n1026 gnd.n1024 585
R8759 gnd.n1024 gnd.n1020 585
R8760 gnd.n1866 gnd.n1865 585
R8761 gnd.n1865 gnd.n1864 585
R8762 gnd.n1031 gnd.n1030 585
R8763 gnd.n1040 gnd.n1031 585
R8764 gnd.n1855 gnd.n1854 585
R8765 gnd.n1854 gnd.n1853 585
R8766 gnd.n1038 gnd.n1037 585
R8767 gnd.n1841 gnd.n1038 585
R8768 gnd.n1813 gnd.n1057 585
R8769 gnd.n1057 gnd.n1047 585
R8770 gnd.n1815 gnd.n1814 585
R8771 gnd.n1816 gnd.n1815 585
R8772 gnd.n1058 gnd.n1056 585
R8773 gnd.n1066 gnd.n1056 585
R8774 gnd.n1791 gnd.n1078 585
R8775 gnd.n1078 gnd.n1065 585
R8776 gnd.n1793 gnd.n1792 585
R8777 gnd.n1794 gnd.n1793 585
R8778 gnd.n1079 gnd.n1077 585
R8779 gnd.n1077 gnd.n1073 585
R8780 gnd.n1779 gnd.n1778 585
R8781 gnd.n1778 gnd.n1777 585
R8782 gnd.n1084 gnd.n1083 585
R8783 gnd.n1093 gnd.n1084 585
R8784 gnd.n1768 gnd.n1767 585
R8785 gnd.n1767 gnd.n1766 585
R8786 gnd.n1091 gnd.n1090 585
R8787 gnd.n1754 gnd.n1091 585
R8788 gnd.n1192 gnd.n1191 585
R8789 gnd.n1192 gnd.n1100 585
R8790 gnd.n1711 gnd.n1710 585
R8791 gnd.n1710 gnd.n1709 585
R8792 gnd.n1712 gnd.n1186 585
R8793 gnd.n1197 gnd.n1186 585
R8794 gnd.n1714 gnd.n1713 585
R8795 gnd.n1715 gnd.n1714 585
R8796 gnd.n1187 gnd.n1185 585
R8797 gnd.n1210 gnd.n1185 585
R8798 gnd.n1170 gnd.n1169 585
R8799 gnd.n1173 gnd.n1170 585
R8800 gnd.n1725 gnd.n1724 585
R8801 gnd.n1724 gnd.n1723 585
R8802 gnd.n1726 gnd.n1164 585
R8803 gnd.n1685 gnd.n1164 585
R8804 gnd.n1728 gnd.n1727 585
R8805 gnd.n1729 gnd.n1728 585
R8806 gnd.n1165 gnd.n1163 585
R8807 gnd.n1224 gnd.n1163 585
R8808 gnd.n1677 gnd.n1676 585
R8809 gnd.n1676 gnd.n1675 585
R8810 gnd.n1221 gnd.n1220 585
R8811 gnd.n1659 gnd.n1221 585
R8812 gnd.n1646 gnd.n1240 585
R8813 gnd.n1240 gnd.n1239 585
R8814 gnd.n1648 gnd.n1647 585
R8815 gnd.n1649 gnd.n1648 585
R8816 gnd.n1241 gnd.n1238 585
R8817 gnd.n1247 gnd.n1238 585
R8818 gnd.n1627 gnd.n1626 585
R8819 gnd.n1628 gnd.n1627 585
R8820 gnd.n1258 gnd.n1257 585
R8821 gnd.n1257 gnd.n1253 585
R8822 gnd.n1617 gnd.n1616 585
R8823 gnd.n1618 gnd.n1617 585
R8824 gnd.n1268 gnd.n1267 585
R8825 gnd.n1273 gnd.n1267 585
R8826 gnd.n1595 gnd.n1286 585
R8827 gnd.n1286 gnd.n1272 585
R8828 gnd.n1597 gnd.n1596 585
R8829 gnd.n1598 gnd.n1597 585
R8830 gnd.n1287 gnd.n1285 585
R8831 gnd.n1285 gnd.n1281 585
R8832 gnd.n1586 gnd.n1585 585
R8833 gnd.n1587 gnd.n1586 585
R8834 gnd.n1294 gnd.n1293 585
R8835 gnd.n1298 gnd.n1293 585
R8836 gnd.n1563 gnd.n1315 585
R8837 gnd.n1315 gnd.n1297 585
R8838 gnd.n1565 gnd.n1564 585
R8839 gnd.n1566 gnd.n1565 585
R8840 gnd.n1316 gnd.n1314 585
R8841 gnd.n1314 gnd.n1305 585
R8842 gnd.n1558 gnd.n1557 585
R8843 gnd.n1557 gnd.n1556 585
R8844 gnd.n1363 gnd.n1362 585
R8845 gnd.n1364 gnd.n1363 585
R8846 gnd.n1517 gnd.n1516 585
R8847 gnd.n1518 gnd.n1517 585
R8848 gnd.n1373 gnd.n1372 585
R8849 gnd.n1372 gnd.n1371 585
R8850 gnd.n1512 gnd.n1511 585
R8851 gnd.n1511 gnd.n1510 585
R8852 gnd.n1376 gnd.n1375 585
R8853 gnd.n1377 gnd.n1376 585
R8854 gnd.n1501 gnd.n1500 585
R8855 gnd.n1502 gnd.n1501 585
R8856 gnd.n1384 gnd.n1383 585
R8857 gnd.n1493 gnd.n1383 585
R8858 gnd.n1496 gnd.n1495 585
R8859 gnd.n1495 gnd.n1494 585
R8860 gnd.n1387 gnd.n1386 585
R8861 gnd.n1388 gnd.n1387 585
R8862 gnd.n1482 gnd.n1481 585
R8863 gnd.n1480 gnd.n1406 585
R8864 gnd.n1479 gnd.n1405 585
R8865 gnd.n1484 gnd.n1405 585
R8866 gnd.n1478 gnd.n1477 585
R8867 gnd.n1476 gnd.n1475 585
R8868 gnd.n1474 gnd.n1473 585
R8869 gnd.n1472 gnd.n1471 585
R8870 gnd.n1470 gnd.n1469 585
R8871 gnd.n1468 gnd.n1467 585
R8872 gnd.n1466 gnd.n1465 585
R8873 gnd.n1464 gnd.n1463 585
R8874 gnd.n1462 gnd.n1461 585
R8875 gnd.n1460 gnd.n1459 585
R8876 gnd.n1458 gnd.n1457 585
R8877 gnd.n1456 gnd.n1455 585
R8878 gnd.n1454 gnd.n1453 585
R8879 gnd.n1452 gnd.n1451 585
R8880 gnd.n1450 gnd.n1449 585
R8881 gnd.n1448 gnd.n1447 585
R8882 gnd.n1446 gnd.n1445 585
R8883 gnd.n1444 gnd.n1443 585
R8884 gnd.n1442 gnd.n1441 585
R8885 gnd.n1440 gnd.n1439 585
R8886 gnd.n1438 gnd.n1437 585
R8887 gnd.n1436 gnd.n1435 585
R8888 gnd.n1393 gnd.n1392 585
R8889 gnd.n1487 gnd.n1486 585
R8890 gnd.n2250 gnd.n2249 585
R8891 gnd.n2252 gnd.n2251 585
R8892 gnd.n2254 gnd.n2253 585
R8893 gnd.n2256 gnd.n2255 585
R8894 gnd.n2258 gnd.n2257 585
R8895 gnd.n2260 gnd.n2259 585
R8896 gnd.n2262 gnd.n2261 585
R8897 gnd.n2264 gnd.n2263 585
R8898 gnd.n2266 gnd.n2265 585
R8899 gnd.n2268 gnd.n2267 585
R8900 gnd.n2270 gnd.n2269 585
R8901 gnd.n2272 gnd.n2271 585
R8902 gnd.n2274 gnd.n2273 585
R8903 gnd.n2276 gnd.n2275 585
R8904 gnd.n2278 gnd.n2277 585
R8905 gnd.n2280 gnd.n2279 585
R8906 gnd.n2282 gnd.n2281 585
R8907 gnd.n2284 gnd.n2283 585
R8908 gnd.n2286 gnd.n2285 585
R8909 gnd.n2288 gnd.n2287 585
R8910 gnd.n2290 gnd.n2289 585
R8911 gnd.n2292 gnd.n2291 585
R8912 gnd.n2294 gnd.n2293 585
R8913 gnd.n2296 gnd.n2295 585
R8914 gnd.n2298 gnd.n2297 585
R8915 gnd.n2299 gnd.n920 585
R8916 gnd.n2300 gnd.n878 585
R8917 gnd.n2338 gnd.n878 585
R8918 gnd.n2248 gnd.n950 585
R8919 gnd.n2248 gnd.n2247 585
R8920 gnd.n1917 gnd.n949 585
R8921 gnd.n959 gnd.n949 585
R8922 gnd.n1919 gnd.n1918 585
R8923 gnd.n1918 gnd.n958 585
R8924 gnd.n1920 gnd.n968 585
R8925 gnd.n2224 gnd.n968 585
R8926 gnd.n1922 gnd.n1921 585
R8927 gnd.n1921 gnd.n966 585
R8928 gnd.n1923 gnd.n979 585
R8929 gnd.n1953 gnd.n979 585
R8930 gnd.n1926 gnd.n1925 585
R8931 gnd.n1925 gnd.n1924 585
R8932 gnd.n1927 gnd.n986 585
R8933 gnd.n1942 gnd.n986 585
R8934 gnd.n1929 gnd.n1928 585
R8935 gnd.n1930 gnd.n1929 585
R8936 gnd.n996 gnd.n995 585
R8937 gnd.n1003 gnd.n995 585
R8938 gnd.n1905 gnd.n1904 585
R8939 gnd.n1904 gnd.n1903 585
R8940 gnd.n999 gnd.n998 585
R8941 gnd.n1013 gnd.n999 585
R8942 gnd.n1829 gnd.n1828 585
R8943 gnd.n1828 gnd.n1012 585
R8944 gnd.n1830 gnd.n1022 585
R8945 gnd.n1881 gnd.n1022 585
R8946 gnd.n1832 gnd.n1831 585
R8947 gnd.n1831 gnd.n1020 585
R8948 gnd.n1833 gnd.n1033 585
R8949 gnd.n1864 gnd.n1033 585
R8950 gnd.n1835 gnd.n1834 585
R8951 gnd.n1834 gnd.n1040 585
R8952 gnd.n1836 gnd.n1039 585
R8953 gnd.n1853 gnd.n1039 585
R8954 gnd.n1838 gnd.n1837 585
R8955 gnd.n1841 gnd.n1838 585
R8956 gnd.n1050 gnd.n1049 585
R8957 gnd.n1049 gnd.n1047 585
R8958 gnd.n1818 gnd.n1817 585
R8959 gnd.n1817 gnd.n1816 585
R8960 gnd.n1053 gnd.n1052 585
R8961 gnd.n1066 gnd.n1053 585
R8962 gnd.n1742 gnd.n1741 585
R8963 gnd.n1741 gnd.n1065 585
R8964 gnd.n1743 gnd.n1075 585
R8965 gnd.n1794 gnd.n1075 585
R8966 gnd.n1745 gnd.n1744 585
R8967 gnd.n1744 gnd.n1073 585
R8968 gnd.n1746 gnd.n1086 585
R8969 gnd.n1777 gnd.n1086 585
R8970 gnd.n1748 gnd.n1747 585
R8971 gnd.n1747 gnd.n1093 585
R8972 gnd.n1749 gnd.n1092 585
R8973 gnd.n1766 gnd.n1092 585
R8974 gnd.n1751 gnd.n1750 585
R8975 gnd.n1754 gnd.n1751 585
R8976 gnd.n1103 gnd.n1102 585
R8977 gnd.n1102 gnd.n1100 585
R8978 gnd.n1194 gnd.n1193 585
R8979 gnd.n1709 gnd.n1193 585
R8980 gnd.n1196 gnd.n1195 585
R8981 gnd.n1197 gnd.n1196 585
R8982 gnd.n1207 gnd.n1183 585
R8983 gnd.n1715 gnd.n1183 585
R8984 gnd.n1209 gnd.n1208 585
R8985 gnd.n1210 gnd.n1209 585
R8986 gnd.n1206 gnd.n1205 585
R8987 gnd.n1206 gnd.n1173 585
R8988 gnd.n1204 gnd.n1171 585
R8989 gnd.n1723 gnd.n1171 585
R8990 gnd.n1160 gnd.n1158 585
R8991 gnd.n1685 gnd.n1160 585
R8992 gnd.n1731 gnd.n1730 585
R8993 gnd.n1730 gnd.n1729 585
R8994 gnd.n1159 gnd.n1157 585
R8995 gnd.n1224 gnd.n1159 585
R8996 gnd.n1656 gnd.n1223 585
R8997 gnd.n1675 gnd.n1223 585
R8998 gnd.n1658 gnd.n1657 585
R8999 gnd.n1659 gnd.n1658 585
R9000 gnd.n1233 gnd.n1232 585
R9001 gnd.n1239 gnd.n1232 585
R9002 gnd.n1651 gnd.n1650 585
R9003 gnd.n1650 gnd.n1649 585
R9004 gnd.n1236 gnd.n1235 585
R9005 gnd.n1247 gnd.n1236 585
R9006 gnd.n1536 gnd.n1255 585
R9007 gnd.n1628 gnd.n1255 585
R9008 gnd.n1538 gnd.n1537 585
R9009 gnd.n1537 gnd.n1253 585
R9010 gnd.n1539 gnd.n1266 585
R9011 gnd.n1618 gnd.n1266 585
R9012 gnd.n1541 gnd.n1540 585
R9013 gnd.n1541 gnd.n1273 585
R9014 gnd.n1543 gnd.n1542 585
R9015 gnd.n1542 gnd.n1272 585
R9016 gnd.n1544 gnd.n1283 585
R9017 gnd.n1598 gnd.n1283 585
R9018 gnd.n1546 gnd.n1545 585
R9019 gnd.n1545 gnd.n1281 585
R9020 gnd.n1547 gnd.n1292 585
R9021 gnd.n1587 gnd.n1292 585
R9022 gnd.n1549 gnd.n1548 585
R9023 gnd.n1549 gnd.n1298 585
R9024 gnd.n1551 gnd.n1550 585
R9025 gnd.n1550 gnd.n1297 585
R9026 gnd.n1552 gnd.n1313 585
R9027 gnd.n1566 gnd.n1313 585
R9028 gnd.n1553 gnd.n1366 585
R9029 gnd.n1366 gnd.n1305 585
R9030 gnd.n1555 gnd.n1554 585
R9031 gnd.n1556 gnd.n1555 585
R9032 gnd.n1367 gnd.n1365 585
R9033 gnd.n1365 gnd.n1364 585
R9034 gnd.n1520 gnd.n1519 585
R9035 gnd.n1519 gnd.n1518 585
R9036 gnd.n1370 gnd.n1369 585
R9037 gnd.n1371 gnd.n1370 585
R9038 gnd.n1509 gnd.n1508 585
R9039 gnd.n1510 gnd.n1509 585
R9040 gnd.n1379 gnd.n1378 585
R9041 gnd.n1378 gnd.n1377 585
R9042 gnd.n1504 gnd.n1503 585
R9043 gnd.n1503 gnd.n1502 585
R9044 gnd.n1382 gnd.n1381 585
R9045 gnd.n1493 gnd.n1382 585
R9046 gnd.n1492 gnd.n1491 585
R9047 gnd.n1494 gnd.n1492 585
R9048 gnd.n1390 gnd.n1389 585
R9049 gnd.n1389 gnd.n1388 585
R9050 gnd.n7674 gnd.n7673 585
R9051 gnd.n7675 gnd.n7674 585
R9052 gnd.n158 gnd.n157 585
R9053 gnd.n7668 gnd.n158 585
R9054 gnd.n7683 gnd.n7682 585
R9055 gnd.n7682 gnd.n7681 585
R9056 gnd.n7684 gnd.n153 585
R9057 gnd.n5889 gnd.n153 585
R9058 gnd.n7686 gnd.n7685 585
R9059 gnd.n7687 gnd.n7686 585
R9060 gnd.n137 gnd.n136 585
R9061 gnd.n5895 gnd.n137 585
R9062 gnd.n7695 gnd.n7694 585
R9063 gnd.n7694 gnd.n7693 585
R9064 gnd.n7696 gnd.n132 585
R9065 gnd.n5901 gnd.n132 585
R9066 gnd.n7698 gnd.n7697 585
R9067 gnd.n7699 gnd.n7698 585
R9068 gnd.n116 gnd.n115 585
R9069 gnd.n5907 gnd.n116 585
R9070 gnd.n7707 gnd.n7706 585
R9071 gnd.n7706 gnd.n7705 585
R9072 gnd.n7708 gnd.n111 585
R9073 gnd.n5913 gnd.n111 585
R9074 gnd.n7710 gnd.n7709 585
R9075 gnd.n7711 gnd.n7710 585
R9076 gnd.n97 gnd.n96 585
R9077 gnd.n5870 gnd.n97 585
R9078 gnd.n7719 gnd.n7718 585
R9079 gnd.n7718 gnd.n7717 585
R9080 gnd.n7720 gnd.n91 585
R9081 gnd.n5861 gnd.n91 585
R9082 gnd.n7722 gnd.n7721 585
R9083 gnd.n7723 gnd.n7722 585
R9084 gnd.n92 gnd.n90 585
R9085 gnd.n5855 gnd.n90 585
R9086 gnd.n5930 gnd.n5929 585
R9087 gnd.n5929 gnd.n5928 585
R9088 gnd.n5931 gnd.n72 585
R9089 gnd.n7731 gnd.n72 585
R9090 gnd.n5932 gnd.n3167 585
R9091 gnd.n5845 gnd.n3167 585
R9092 gnd.n5934 gnd.n5933 585
R9093 gnd.n5935 gnd.n5934 585
R9094 gnd.n3168 gnd.n3160 585
R9095 gnd.n5940 gnd.n3160 585
R9096 gnd.n5840 gnd.n5839 585
R9097 gnd.n5839 gnd.n3156 585
R9098 gnd.n5838 gnd.n5837 585
R9099 gnd.n5838 gnd.n3149 585
R9100 gnd.n3139 gnd.n3138 585
R9101 gnd.n5949 gnd.n3139 585
R9102 gnd.n5955 gnd.n5954 585
R9103 gnd.n5954 gnd.n5953 585
R9104 gnd.n5956 gnd.n3134 585
R9105 gnd.n5828 gnd.n3134 585
R9106 gnd.n5958 gnd.n5957 585
R9107 gnd.n5959 gnd.n5958 585
R9108 gnd.n3120 gnd.n3119 585
R9109 gnd.n5810 gnd.n3120 585
R9110 gnd.n5967 gnd.n5966 585
R9111 gnd.n5966 gnd.n5965 585
R9112 gnd.n5968 gnd.n3115 585
R9113 gnd.n5803 gnd.n3115 585
R9114 gnd.n5970 gnd.n5969 585
R9115 gnd.n5971 gnd.n5970 585
R9116 gnd.n3099 gnd.n3098 585
R9117 gnd.n5747 gnd.n3099 585
R9118 gnd.n5979 gnd.n5978 585
R9119 gnd.n5978 gnd.n5977 585
R9120 gnd.n5980 gnd.n3094 585
R9121 gnd.n5758 gnd.n3094 585
R9122 gnd.n5982 gnd.n5981 585
R9123 gnd.n5983 gnd.n5982 585
R9124 gnd.n3079 gnd.n3078 585
R9125 gnd.n5738 gnd.n3079 585
R9126 gnd.n5991 gnd.n5990 585
R9127 gnd.n5990 gnd.n5989 585
R9128 gnd.n5992 gnd.n3073 585
R9129 gnd.n5730 gnd.n3073 585
R9130 gnd.n5994 gnd.n5993 585
R9131 gnd.n5995 gnd.n5994 585
R9132 gnd.n3074 gnd.n3072 585
R9133 gnd.n5195 gnd.n3072 585
R9134 gnd.n5723 gnd.n3060 585
R9135 gnd.n6001 gnd.n3060 585
R9136 gnd.n5282 gnd.n5281 585
R9137 gnd.n5245 gnd.n5244 585
R9138 gnd.n5296 gnd.n5295 585
R9139 gnd.n5298 gnd.n5243 585
R9140 gnd.n5301 gnd.n5300 585
R9141 gnd.n5236 gnd.n5235 585
R9142 gnd.n5315 gnd.n5314 585
R9143 gnd.n5317 gnd.n5234 585
R9144 gnd.n5320 gnd.n5319 585
R9145 gnd.n5227 gnd.n5226 585
R9146 gnd.n5334 gnd.n5333 585
R9147 gnd.n5336 gnd.n5225 585
R9148 gnd.n5339 gnd.n5338 585
R9149 gnd.n5218 gnd.n5217 585
R9150 gnd.n5354 gnd.n5353 585
R9151 gnd.n5356 gnd.n5216 585
R9152 gnd.n5359 gnd.n5358 585
R9153 gnd.n5360 gnd.n5213 585
R9154 gnd.n5212 gnd.n5211 585
R9155 gnd.n5212 gnd.n3048 585
R9156 gnd.n7662 gnd.n7661 585
R9157 gnd.n183 gnd.n182 585
R9158 gnd.n241 gnd.n240 585
R9159 gnd.n193 gnd.n192 585
R9160 gnd.n236 gnd.n235 585
R9161 gnd.n234 gnd.n233 585
R9162 gnd.n232 gnd.n231 585
R9163 gnd.n225 gnd.n195 585
R9164 gnd.n227 gnd.n226 585
R9165 gnd.n224 gnd.n223 585
R9166 gnd.n222 gnd.n221 585
R9167 gnd.n215 gnd.n197 585
R9168 gnd.n217 gnd.n216 585
R9169 gnd.n214 gnd.n213 585
R9170 gnd.n212 gnd.n211 585
R9171 gnd.n205 gnd.n199 585
R9172 gnd.n207 gnd.n206 585
R9173 gnd.n204 gnd.n203 585
R9174 gnd.n202 gnd.n172 585
R9175 gnd.n7659 gnd.n172 585
R9176 gnd.n7665 gnd.n170 585
R9177 gnd.n7675 gnd.n170 585
R9178 gnd.n7667 gnd.n7666 585
R9179 gnd.n7668 gnd.n7667 585
R9180 gnd.n177 gnd.n161 585
R9181 gnd.n7681 gnd.n161 585
R9182 gnd.n5888 gnd.n5887 585
R9183 gnd.n5889 gnd.n5888 585
R9184 gnd.n5882 gnd.n151 585
R9185 gnd.n7687 gnd.n151 585
R9186 gnd.n5897 gnd.n5896 585
R9187 gnd.n5896 gnd.n5895 585
R9188 gnd.n5898 gnd.n140 585
R9189 gnd.n7693 gnd.n140 585
R9190 gnd.n5900 gnd.n5899 585
R9191 gnd.n5901 gnd.n5900 585
R9192 gnd.n3232 gnd.n130 585
R9193 gnd.n7699 gnd.n130 585
R9194 gnd.n5909 gnd.n5908 585
R9195 gnd.n5908 gnd.n5907 585
R9196 gnd.n5910 gnd.n119 585
R9197 gnd.n7705 gnd.n119 585
R9198 gnd.n5912 gnd.n5911 585
R9199 gnd.n5913 gnd.n5912 585
R9200 gnd.n3228 gnd.n110 585
R9201 gnd.n7711 gnd.n110 585
R9202 gnd.n5869 gnd.n5868 585
R9203 gnd.n5870 gnd.n5869 585
R9204 gnd.n3235 gnd.n100 585
R9205 gnd.n7717 gnd.n100 585
R9206 gnd.n5863 gnd.n5862 585
R9207 gnd.n5862 gnd.n5861 585
R9208 gnd.n3237 gnd.n88 585
R9209 gnd.n7723 gnd.n88 585
R9210 gnd.n5854 gnd.n5853 585
R9211 gnd.n5855 gnd.n5854 585
R9212 gnd.n68 gnd.n67 585
R9213 gnd.n5928 gnd.n68 585
R9214 gnd.n7733 gnd.n7732 585
R9215 gnd.n7732 gnd.n7731 585
R9216 gnd.n7734 gnd.n66 585
R9217 gnd.n5845 gnd.n66 585
R9218 gnd.n3165 gnd.n64 585
R9219 gnd.n5935 gnd.n3165 585
R9220 gnd.n5818 gnd.n3158 585
R9221 gnd.n5940 gnd.n3158 585
R9222 gnd.n5820 gnd.n5817 585
R9223 gnd.n5817 gnd.n3156 585
R9224 gnd.n5821 gnd.n5816 585
R9225 gnd.n5816 gnd.n3149 585
R9226 gnd.n5822 gnd.n3148 585
R9227 gnd.n5949 gnd.n3148 585
R9228 gnd.n3243 gnd.n3142 585
R9229 gnd.n5953 gnd.n3142 585
R9230 gnd.n5827 gnd.n5826 585
R9231 gnd.n5828 gnd.n5827 585
R9232 gnd.n3242 gnd.n3133 585
R9233 gnd.n5959 gnd.n3133 585
R9234 gnd.n5812 gnd.n5811 585
R9235 gnd.n5811 gnd.n5810 585
R9236 gnd.n3245 gnd.n3122 585
R9237 gnd.n5965 gnd.n3122 585
R9238 gnd.n5750 gnd.n3247 585
R9239 gnd.n5803 gnd.n3247 585
R9240 gnd.n5751 gnd.n3113 585
R9241 gnd.n5971 gnd.n3113 585
R9242 gnd.n5752 gnd.n5748 585
R9243 gnd.n5748 gnd.n5747 585
R9244 gnd.n3255 gnd.n3102 585
R9245 gnd.n5977 gnd.n3102 585
R9246 gnd.n5757 gnd.n5756 585
R9247 gnd.n5758 gnd.n5757 585
R9248 gnd.n3254 gnd.n3093 585
R9249 gnd.n5983 gnd.n3093 585
R9250 gnd.n5737 gnd.n5736 585
R9251 gnd.n5738 gnd.n5737 585
R9252 gnd.n3260 gnd.n3082 585
R9253 gnd.n5989 gnd.n3082 585
R9254 gnd.n5732 gnd.n5731 585
R9255 gnd.n5731 gnd.n5730 585
R9256 gnd.n3262 gnd.n3070 585
R9257 gnd.n5995 gnd.n3070 585
R9258 gnd.n5197 gnd.n5196 585
R9259 gnd.n5196 gnd.n5195 585
R9260 gnd.n5198 gnd.n3058 585
R9261 gnd.n6001 gnd.n3058 585
R9262 gnd.n2233 gnd.n900 585
R9263 gnd.n900 gnd.n877 585
R9264 gnd.n2234 gnd.n961 585
R9265 gnd.n961 gnd.n951 585
R9266 gnd.n2236 gnd.n2235 585
R9267 gnd.n2237 gnd.n2236 585
R9268 gnd.n962 gnd.n960 585
R9269 gnd.n969 gnd.n960 585
R9270 gnd.n2227 gnd.n2226 585
R9271 gnd.n2226 gnd.n2225 585
R9272 gnd.n965 gnd.n964 585
R9273 gnd.n1952 gnd.n965 585
R9274 gnd.n1938 gnd.n988 585
R9275 gnd.n988 gnd.n978 585
R9276 gnd.n1940 gnd.n1939 585
R9277 gnd.n1941 gnd.n1940 585
R9278 gnd.n989 gnd.n987 585
R9279 gnd.n987 gnd.n985 585
R9280 gnd.n1933 gnd.n1932 585
R9281 gnd.n1932 gnd.n1931 585
R9282 gnd.n992 gnd.n991 585
R9283 gnd.n1001 gnd.n992 585
R9284 gnd.n1889 gnd.n1015 585
R9285 gnd.n1015 gnd.n1000 585
R9286 gnd.n1891 gnd.n1890 585
R9287 gnd.n1892 gnd.n1891 585
R9288 gnd.n1016 gnd.n1014 585
R9289 gnd.n1023 gnd.n1014 585
R9290 gnd.n1884 gnd.n1883 585
R9291 gnd.n1883 gnd.n1882 585
R9292 gnd.n1019 gnd.n1018 585
R9293 gnd.n1863 gnd.n1019 585
R9294 gnd.n1849 gnd.n1042 585
R9295 gnd.n1042 gnd.n1032 585
R9296 gnd.n1851 gnd.n1850 585
R9297 gnd.n1852 gnd.n1851 585
R9298 gnd.n1043 gnd.n1041 585
R9299 gnd.n1840 gnd.n1041 585
R9300 gnd.n1844 gnd.n1843 585
R9301 gnd.n1843 gnd.n1842 585
R9302 gnd.n1046 gnd.n1045 585
R9303 gnd.n1055 gnd.n1046 585
R9304 gnd.n1802 gnd.n1068 585
R9305 gnd.n1068 gnd.n1054 585
R9306 gnd.n1804 gnd.n1803 585
R9307 gnd.n1805 gnd.n1804 585
R9308 gnd.n1069 gnd.n1067 585
R9309 gnd.n1076 gnd.n1067 585
R9310 gnd.n1797 gnd.n1796 585
R9311 gnd.n1796 gnd.n1795 585
R9312 gnd.n1072 gnd.n1071 585
R9313 gnd.n1776 gnd.n1072 585
R9314 gnd.n1762 gnd.n1095 585
R9315 gnd.n1095 gnd.n1085 585
R9316 gnd.n1764 gnd.n1763 585
R9317 gnd.n1765 gnd.n1764 585
R9318 gnd.n1096 gnd.n1094 585
R9319 gnd.n1753 gnd.n1094 585
R9320 gnd.n1757 gnd.n1756 585
R9321 gnd.n1756 gnd.n1755 585
R9322 gnd.n1099 gnd.n1098 585
R9323 gnd.n1708 gnd.n1099 585
R9324 gnd.n1201 gnd.n1200 585
R9325 gnd.n1202 gnd.n1201 585
R9326 gnd.n1181 gnd.n1180 585
R9327 gnd.n1184 gnd.n1181 585
R9328 gnd.n1718 gnd.n1717 585
R9329 gnd.n1717 gnd.n1716 585
R9330 gnd.n1719 gnd.n1175 585
R9331 gnd.n1211 gnd.n1175 585
R9332 gnd.n1721 gnd.n1720 585
R9333 gnd.n1722 gnd.n1721 585
R9334 gnd.n1176 gnd.n1174 585
R9335 gnd.n1686 gnd.n1174 585
R9336 gnd.n1670 gnd.n1669 585
R9337 gnd.n1669 gnd.n1162 585
R9338 gnd.n1671 gnd.n1226 585
R9339 gnd.n1226 gnd.n1161 585
R9340 gnd.n1673 gnd.n1672 585
R9341 gnd.n1674 gnd.n1673 585
R9342 gnd.n1227 gnd.n1225 585
R9343 gnd.n1225 gnd.n1222 585
R9344 gnd.n1662 gnd.n1661 585
R9345 gnd.n1661 gnd.n1660 585
R9346 gnd.n1230 gnd.n1229 585
R9347 gnd.n1237 gnd.n1230 585
R9348 gnd.n1636 gnd.n1635 585
R9349 gnd.n1637 gnd.n1636 585
R9350 gnd.n1249 gnd.n1248 585
R9351 gnd.n1256 gnd.n1248 585
R9352 gnd.n1631 gnd.n1630 585
R9353 gnd.n1630 gnd.n1629 585
R9354 gnd.n1252 gnd.n1251 585
R9355 gnd.n1619 gnd.n1252 585
R9356 gnd.n1606 gnd.n1276 585
R9357 gnd.n1276 gnd.n1275 585
R9358 gnd.n1608 gnd.n1607 585
R9359 gnd.n1609 gnd.n1608 585
R9360 gnd.n1277 gnd.n1274 585
R9361 gnd.n1284 gnd.n1274 585
R9362 gnd.n1601 gnd.n1600 585
R9363 gnd.n1600 gnd.n1599 585
R9364 gnd.n1280 gnd.n1279 585
R9365 gnd.n1588 gnd.n1280 585
R9366 gnd.n1575 gnd.n1301 585
R9367 gnd.n1301 gnd.n1300 585
R9368 gnd.n1577 gnd.n1576 585
R9369 gnd.n1578 gnd.n1577 585
R9370 gnd.n1571 gnd.n1299 585
R9371 gnd.n1570 gnd.n1569 585
R9372 gnd.n1304 gnd.n1303 585
R9373 gnd.n1567 gnd.n1304 585
R9374 gnd.n1326 gnd.n1325 585
R9375 gnd.n1329 gnd.n1328 585
R9376 gnd.n1327 gnd.n1322 585
R9377 gnd.n1334 gnd.n1333 585
R9378 gnd.n1336 gnd.n1335 585
R9379 gnd.n1339 gnd.n1338 585
R9380 gnd.n1337 gnd.n1320 585
R9381 gnd.n1344 gnd.n1343 585
R9382 gnd.n1346 gnd.n1345 585
R9383 gnd.n1349 gnd.n1348 585
R9384 gnd.n1347 gnd.n1318 585
R9385 gnd.n1354 gnd.n1353 585
R9386 gnd.n1358 gnd.n1355 585
R9387 gnd.n1359 gnd.n1296 585
R9388 gnd.n2239 gnd.n915 585
R9389 gnd.n2306 gnd.n2305 585
R9390 gnd.n2308 gnd.n2307 585
R9391 gnd.n2310 gnd.n2309 585
R9392 gnd.n2312 gnd.n2311 585
R9393 gnd.n2314 gnd.n2313 585
R9394 gnd.n2316 gnd.n2315 585
R9395 gnd.n2318 gnd.n2317 585
R9396 gnd.n2320 gnd.n2319 585
R9397 gnd.n2322 gnd.n2321 585
R9398 gnd.n2324 gnd.n2323 585
R9399 gnd.n2326 gnd.n2325 585
R9400 gnd.n2328 gnd.n2327 585
R9401 gnd.n2331 gnd.n2330 585
R9402 gnd.n2329 gnd.n903 585
R9403 gnd.n2335 gnd.n901 585
R9404 gnd.n2337 gnd.n2336 585
R9405 gnd.n2338 gnd.n2337 585
R9406 gnd.n2240 gnd.n956 585
R9407 gnd.n2240 gnd.n877 585
R9408 gnd.n2242 gnd.n2241 585
R9409 gnd.n2241 gnd.n951 585
R9410 gnd.n2238 gnd.n955 585
R9411 gnd.n2238 gnd.n2237 585
R9412 gnd.n2217 gnd.n957 585
R9413 gnd.n969 gnd.n957 585
R9414 gnd.n2216 gnd.n967 585
R9415 gnd.n2225 gnd.n967 585
R9416 gnd.n1951 gnd.n974 585
R9417 gnd.n1952 gnd.n1951 585
R9418 gnd.n1950 gnd.n1949 585
R9419 gnd.n1950 gnd.n978 585
R9420 gnd.n1948 gnd.n980 585
R9421 gnd.n1941 gnd.n980 585
R9422 gnd.n993 gnd.n981 585
R9423 gnd.n993 gnd.n985 585
R9424 gnd.n1897 gnd.n994 585
R9425 gnd.n1931 gnd.n994 585
R9426 gnd.n1896 gnd.n1895 585
R9427 gnd.n1895 gnd.n1001 585
R9428 gnd.n1894 gnd.n1009 585
R9429 gnd.n1894 gnd.n1000 585
R9430 gnd.n1893 gnd.n1011 585
R9431 gnd.n1893 gnd.n1892 585
R9432 gnd.n1872 gnd.n1010 585
R9433 gnd.n1023 gnd.n1010 585
R9434 gnd.n1871 gnd.n1021 585
R9435 gnd.n1882 gnd.n1021 585
R9436 gnd.n1862 gnd.n1028 585
R9437 gnd.n1863 gnd.n1862 585
R9438 gnd.n1861 gnd.n1860 585
R9439 gnd.n1861 gnd.n1032 585
R9440 gnd.n1859 gnd.n1034 585
R9441 gnd.n1852 gnd.n1034 585
R9442 gnd.n1839 gnd.n1035 585
R9443 gnd.n1840 gnd.n1839 585
R9444 gnd.n1810 gnd.n1048 585
R9445 gnd.n1842 gnd.n1048 585
R9446 gnd.n1809 gnd.n1808 585
R9447 gnd.n1808 gnd.n1055 585
R9448 gnd.n1807 gnd.n1062 585
R9449 gnd.n1807 gnd.n1054 585
R9450 gnd.n1806 gnd.n1064 585
R9451 gnd.n1806 gnd.n1805 585
R9452 gnd.n1785 gnd.n1063 585
R9453 gnd.n1076 gnd.n1063 585
R9454 gnd.n1784 gnd.n1074 585
R9455 gnd.n1795 gnd.n1074 585
R9456 gnd.n1775 gnd.n1081 585
R9457 gnd.n1776 gnd.n1775 585
R9458 gnd.n1774 gnd.n1773 585
R9459 gnd.n1774 gnd.n1085 585
R9460 gnd.n1772 gnd.n1087 585
R9461 gnd.n1765 gnd.n1087 585
R9462 gnd.n1752 gnd.n1088 585
R9463 gnd.n1753 gnd.n1752 585
R9464 gnd.n1705 gnd.n1101 585
R9465 gnd.n1755 gnd.n1101 585
R9466 gnd.n1707 gnd.n1706 585
R9467 gnd.n1708 gnd.n1707 585
R9468 gnd.n1700 gnd.n1203 585
R9469 gnd.n1203 gnd.n1202 585
R9470 gnd.n1698 gnd.n1697 585
R9471 gnd.n1697 gnd.n1184 585
R9472 gnd.n1695 gnd.n1182 585
R9473 gnd.n1716 gnd.n1182 585
R9474 gnd.n1213 gnd.n1212 585
R9475 gnd.n1212 gnd.n1211 585
R9476 gnd.n1689 gnd.n1172 585
R9477 gnd.n1722 gnd.n1172 585
R9478 gnd.n1688 gnd.n1687 585
R9479 gnd.n1687 gnd.n1686 585
R9480 gnd.n1684 gnd.n1215 585
R9481 gnd.n1684 gnd.n1162 585
R9482 gnd.n1683 gnd.n1682 585
R9483 gnd.n1683 gnd.n1161 585
R9484 gnd.n1218 gnd.n1217 585
R9485 gnd.n1674 gnd.n1217 585
R9486 gnd.n1642 gnd.n1641 585
R9487 gnd.n1641 gnd.n1222 585
R9488 gnd.n1643 gnd.n1231 585
R9489 gnd.n1660 gnd.n1231 585
R9490 gnd.n1640 gnd.n1639 585
R9491 gnd.n1639 gnd.n1237 585
R9492 gnd.n1638 gnd.n1245 585
R9493 gnd.n1638 gnd.n1637 585
R9494 gnd.n1623 gnd.n1246 585
R9495 gnd.n1256 gnd.n1246 585
R9496 gnd.n1622 gnd.n1254 585
R9497 gnd.n1629 gnd.n1254 585
R9498 gnd.n1621 gnd.n1620 585
R9499 gnd.n1620 gnd.n1619 585
R9500 gnd.n1265 gnd.n1262 585
R9501 gnd.n1275 gnd.n1265 585
R9502 gnd.n1611 gnd.n1610 585
R9503 gnd.n1610 gnd.n1609 585
R9504 gnd.n1271 gnd.n1270 585
R9505 gnd.n1284 gnd.n1271 585
R9506 gnd.n1591 gnd.n1282 585
R9507 gnd.n1599 gnd.n1282 585
R9508 gnd.n1590 gnd.n1589 585
R9509 gnd.n1589 gnd.n1588 585
R9510 gnd.n1291 gnd.n1289 585
R9511 gnd.n1300 gnd.n1291 585
R9512 gnd.n1580 gnd.n1579 585
R9513 gnd.n1579 gnd.n1578 585
R9514 gnd.n5474 gnd.n5473 585
R9515 gnd.n5475 gnd.n5474 585
R9516 gnd.n5388 gnd.n3341 585
R9517 gnd.n3347 gnd.n3341 585
R9518 gnd.n5387 gnd.n5386 585
R9519 gnd.n5386 gnd.n5385 585
R9520 gnd.n3344 gnd.n3343 585
R9521 gnd.n3434 gnd.n3344 585
R9522 gnd.n5176 gnd.n3371 585
R9523 gnd.n3437 gnd.n3371 585
R9524 gnd.n5178 gnd.n5177 585
R9525 gnd.n5179 gnd.n5178 585
R9526 gnd.n5175 gnd.n3370 585
R9527 gnd.n5170 gnd.n3370 585
R9528 gnd.n5174 gnd.n5173 585
R9529 gnd.n5173 gnd.n5172 585
R9530 gnd.n3373 gnd.n3372 585
R9531 gnd.n5157 gnd.n3373 585
R9532 gnd.n5143 gnd.n3395 585
R9533 gnd.n3395 gnd.n3383 585
R9534 gnd.n5145 gnd.n5144 585
R9535 gnd.n5146 gnd.n5145 585
R9536 gnd.n5142 gnd.n3394 585
R9537 gnd.n3394 gnd.n3390 585
R9538 gnd.n5141 gnd.n5140 585
R9539 gnd.n5140 gnd.n5139 585
R9540 gnd.n3397 gnd.n3396 585
R9541 gnd.n3451 gnd.n3397 585
R9542 gnd.n5128 gnd.n5127 585
R9543 gnd.n5129 gnd.n5128 585
R9544 gnd.n5126 gnd.n3408 585
R9545 gnd.n3408 gnd.n3405 585
R9546 gnd.n5125 gnd.n5124 585
R9547 gnd.n5124 gnd.n5123 585
R9548 gnd.n3410 gnd.n3409 585
R9549 gnd.n5097 gnd.n3410 585
R9550 gnd.n5110 gnd.n5109 585
R9551 gnd.n5111 gnd.n5110 585
R9552 gnd.n5108 gnd.n3422 585
R9553 gnd.n5103 gnd.n3422 585
R9554 gnd.n5107 gnd.n5106 585
R9555 gnd.n5106 gnd.n5105 585
R9556 gnd.n3424 gnd.n3423 585
R9557 gnd.n5083 gnd.n3424 585
R9558 gnd.n5074 gnd.n3470 585
R9559 gnd.n3470 gnd.n3463 585
R9560 gnd.n5076 gnd.n5075 585
R9561 gnd.n5077 gnd.n5076 585
R9562 gnd.n5073 gnd.n3469 585
R9563 gnd.n5034 gnd.n3469 585
R9564 gnd.n5072 gnd.n5071 585
R9565 gnd.n5071 gnd.n5070 585
R9566 gnd.n3472 gnd.n3471 585
R9567 gnd.n4977 gnd.n3472 585
R9568 gnd.n5055 gnd.n5054 585
R9569 gnd.n5056 gnd.n5055 585
R9570 gnd.n5053 gnd.n3484 585
R9571 gnd.n3484 gnd.n3480 585
R9572 gnd.n5052 gnd.n5051 585
R9573 gnd.n5051 gnd.n5050 585
R9574 gnd.n3486 gnd.n3485 585
R9575 gnd.n4984 gnd.n3486 585
R9576 gnd.n5025 gnd.n5024 585
R9577 gnd.n5026 gnd.n5025 585
R9578 gnd.n5023 gnd.n3498 585
R9579 gnd.n3498 gnd.n3495 585
R9580 gnd.n5022 gnd.n5021 585
R9581 gnd.n5021 gnd.n5020 585
R9582 gnd.n3500 gnd.n3499 585
R9583 gnd.n4992 gnd.n3500 585
R9584 gnd.n5005 gnd.n5004 585
R9585 gnd.n5006 gnd.n5005 585
R9586 gnd.n5003 gnd.n3511 585
R9587 gnd.n4998 gnd.n3511 585
R9588 gnd.n5002 gnd.n5001 585
R9589 gnd.n5001 gnd.n5000 585
R9590 gnd.n3513 gnd.n3512 585
R9591 gnd.n4972 gnd.n3513 585
R9592 gnd.n4955 gnd.n3527 585
R9593 gnd.n4940 gnd.n3527 585
R9594 gnd.n4957 gnd.n4956 585
R9595 gnd.n4958 gnd.n4957 585
R9596 gnd.n4954 gnd.n3526 585
R9597 gnd.n3532 gnd.n3526 585
R9598 gnd.n4953 gnd.n4952 585
R9599 gnd.n4952 gnd.n4951 585
R9600 gnd.n3529 gnd.n3528 585
R9601 gnd.n4930 gnd.n3529 585
R9602 gnd.n4917 gnd.n3546 585
R9603 gnd.n3546 gnd.n3539 585
R9604 gnd.n4919 gnd.n4918 585
R9605 gnd.n4920 gnd.n4919 585
R9606 gnd.n4916 gnd.n3545 585
R9607 gnd.n3551 gnd.n3545 585
R9608 gnd.n4915 gnd.n4914 585
R9609 gnd.n4914 gnd.n4913 585
R9610 gnd.n3548 gnd.n3547 585
R9611 gnd.n4824 gnd.n3548 585
R9612 gnd.n4901 gnd.n4900 585
R9613 gnd.n4902 gnd.n4901 585
R9614 gnd.n4899 gnd.n3562 585
R9615 gnd.n3562 gnd.n3558 585
R9616 gnd.n4898 gnd.n4897 585
R9617 gnd.n4897 gnd.n4896 585
R9618 gnd.n3564 gnd.n3563 585
R9619 gnd.n4832 gnd.n3564 585
R9620 gnd.n4870 gnd.n4869 585
R9621 gnd.n4871 gnd.n4870 585
R9622 gnd.n4868 gnd.n3576 585
R9623 gnd.n3576 gnd.n3573 585
R9624 gnd.n4867 gnd.n4866 585
R9625 gnd.n4866 gnd.n4865 585
R9626 gnd.n3578 gnd.n3577 585
R9627 gnd.n4839 gnd.n3578 585
R9628 gnd.n4852 gnd.n4851 585
R9629 gnd.n4853 gnd.n4852 585
R9630 gnd.n4850 gnd.n3591 585
R9631 gnd.n4845 gnd.n3591 585
R9632 gnd.n4849 gnd.n4848 585
R9633 gnd.n4848 gnd.n4847 585
R9634 gnd.n3593 gnd.n3592 585
R9635 gnd.n4819 gnd.n3593 585
R9636 gnd.n4805 gnd.n4804 585
R9637 gnd.n4804 gnd.n4803 585
R9638 gnd.n4806 gnd.n3609 585
R9639 gnd.n4801 gnd.n3609 585
R9640 gnd.n4808 gnd.n4807 585
R9641 gnd.n4809 gnd.n4808 585
R9642 gnd.n3610 gnd.n3608 585
R9643 gnd.n4795 gnd.n3608 585
R9644 gnd.n4792 gnd.n4791 585
R9645 gnd.n4793 gnd.n4792 585
R9646 gnd.n4790 gnd.n3613 585
R9647 gnd.n3619 gnd.n3613 585
R9648 gnd.n4789 gnd.n4788 585
R9649 gnd.n4788 gnd.n4787 585
R9650 gnd.n3615 gnd.n3614 585
R9651 gnd.n4774 gnd.n3615 585
R9652 gnd.n4762 gnd.n3633 585
R9653 gnd.n3633 gnd.n3625 585
R9654 gnd.n4764 gnd.n4763 585
R9655 gnd.n4765 gnd.n4764 585
R9656 gnd.n4761 gnd.n3632 585
R9657 gnd.n3638 gnd.n3632 585
R9658 gnd.n4760 gnd.n4759 585
R9659 gnd.n4759 gnd.n4758 585
R9660 gnd.n3635 gnd.n3634 585
R9661 gnd.n4645 gnd.n3635 585
R9662 gnd.n4745 gnd.n4744 585
R9663 gnd.n4746 gnd.n4745 585
R9664 gnd.n4743 gnd.n3649 585
R9665 gnd.n3649 gnd.n3645 585
R9666 gnd.n4742 gnd.n4741 585
R9667 gnd.n4741 gnd.n4740 585
R9668 gnd.n3651 gnd.n3650 585
R9669 gnd.n4653 gnd.n3651 585
R9670 gnd.n4693 gnd.n4692 585
R9671 gnd.n4694 gnd.n4693 585
R9672 gnd.n4691 gnd.n3662 585
R9673 gnd.n3666 gnd.n3662 585
R9674 gnd.n4690 gnd.n4689 585
R9675 gnd.n4689 gnd.n4688 585
R9676 gnd.n3664 gnd.n3663 585
R9677 gnd.n4661 gnd.n3664 585
R9678 gnd.n4674 gnd.n4673 585
R9679 gnd.n4675 gnd.n4674 585
R9680 gnd.n4672 gnd.n3676 585
R9681 gnd.n4667 gnd.n3676 585
R9682 gnd.n4671 gnd.n4670 585
R9683 gnd.n4670 gnd.n4669 585
R9684 gnd.n3678 gnd.n3677 585
R9685 gnd.n4640 gnd.n3678 585
R9686 gnd.n4626 gnd.n4625 585
R9687 gnd.n4625 gnd.n4624 585
R9688 gnd.n4627 gnd.n3691 585
R9689 gnd.n4572 gnd.n3691 585
R9690 gnd.n4629 gnd.n4628 585
R9691 gnd.n4630 gnd.n4629 585
R9692 gnd.n3692 gnd.n3690 585
R9693 gnd.n4576 gnd.n3690 585
R9694 gnd.n4604 gnd.n4603 585
R9695 gnd.n4605 gnd.n4604 585
R9696 gnd.n4602 gnd.n3703 585
R9697 gnd.n3707 gnd.n3703 585
R9698 gnd.n4601 gnd.n4600 585
R9699 gnd.n4600 gnd.n4599 585
R9700 gnd.n3705 gnd.n3704 585
R9701 gnd.n4586 gnd.n3705 585
R9702 gnd.n4565 gnd.n3721 585
R9703 gnd.n3721 gnd.n3713 585
R9704 gnd.n4567 gnd.n4566 585
R9705 gnd.n4568 gnd.n4567 585
R9706 gnd.n4564 gnd.n3720 585
R9707 gnd.n4554 gnd.n3720 585
R9708 gnd.n4563 gnd.n4562 585
R9709 gnd.n4562 gnd.n4561 585
R9710 gnd.n3723 gnd.n3722 585
R9711 gnd.n4526 gnd.n3723 585
R9712 gnd.n4535 gnd.n4534 585
R9713 gnd.n4534 gnd.n2942 585
R9714 gnd.n4536 gnd.n4533 585
R9715 gnd.n4533 gnd.n2940 585
R9716 gnd.n4538 gnd.n4537 585
R9717 gnd.n4539 gnd.n4538 585
R9718 gnd.n2930 gnd.n2929 585
R9719 gnd.n3734 gnd.n2930 585
R9720 gnd.n6138 gnd.n6137 585
R9721 gnd.n6137 gnd.n6136 585
R9722 gnd.n6139 gnd.n2927 585
R9723 gnd.n4518 gnd.n2927 585
R9724 gnd.n6141 gnd.n6140 585
R9725 gnd.n6142 gnd.n6141 585
R9726 gnd.n2928 gnd.n2926 585
R9727 gnd.n4507 gnd.n2926 585
R9728 gnd.n3746 gnd.n3745 585
R9729 gnd.n3747 gnd.n3746 585
R9730 gnd.n2911 gnd.n2910 585
R9731 gnd.n4501 gnd.n2911 585
R9732 gnd.n6152 gnd.n6151 585
R9733 gnd.n6151 gnd.n6150 585
R9734 gnd.n6153 gnd.n2889 585
R9735 gnd.n3824 gnd.n2889 585
R9736 gnd.n6218 gnd.n6217 585
R9737 gnd.n6216 gnd.n2888 585
R9738 gnd.n6215 gnd.n2887 585
R9739 gnd.n6220 gnd.n2887 585
R9740 gnd.n6214 gnd.n6213 585
R9741 gnd.n6212 gnd.n6211 585
R9742 gnd.n6210 gnd.n6209 585
R9743 gnd.n6208 gnd.n6207 585
R9744 gnd.n6206 gnd.n6205 585
R9745 gnd.n6204 gnd.n6203 585
R9746 gnd.n6202 gnd.n6201 585
R9747 gnd.n6200 gnd.n6199 585
R9748 gnd.n6198 gnd.n6197 585
R9749 gnd.n6196 gnd.n6195 585
R9750 gnd.n6194 gnd.n6193 585
R9751 gnd.n6192 gnd.n6191 585
R9752 gnd.n6190 gnd.n6189 585
R9753 gnd.n6188 gnd.n6187 585
R9754 gnd.n6186 gnd.n6185 585
R9755 gnd.n6184 gnd.n6183 585
R9756 gnd.n6182 gnd.n6181 585
R9757 gnd.n6180 gnd.n6179 585
R9758 gnd.n6178 gnd.n6177 585
R9759 gnd.n6176 gnd.n6175 585
R9760 gnd.n6174 gnd.n6173 585
R9761 gnd.n6172 gnd.n6171 585
R9762 gnd.n6170 gnd.n6169 585
R9763 gnd.n6168 gnd.n6167 585
R9764 gnd.n6166 gnd.n6165 585
R9765 gnd.n6164 gnd.n6163 585
R9766 gnd.n6162 gnd.n6161 585
R9767 gnd.n6160 gnd.n6159 585
R9768 gnd.n6158 gnd.n2851 585
R9769 gnd.n6223 gnd.n6222 585
R9770 gnd.n2853 gnd.n2850 585
R9771 gnd.n3761 gnd.n3760 585
R9772 gnd.n3763 gnd.n3762 585
R9773 gnd.n3766 gnd.n3765 585
R9774 gnd.n3768 gnd.n3767 585
R9775 gnd.n3770 gnd.n3769 585
R9776 gnd.n3772 gnd.n3771 585
R9777 gnd.n3774 gnd.n3773 585
R9778 gnd.n3776 gnd.n3775 585
R9779 gnd.n3778 gnd.n3777 585
R9780 gnd.n3780 gnd.n3779 585
R9781 gnd.n3782 gnd.n3781 585
R9782 gnd.n3784 gnd.n3783 585
R9783 gnd.n3786 gnd.n3785 585
R9784 gnd.n3788 gnd.n3787 585
R9785 gnd.n3790 gnd.n3789 585
R9786 gnd.n3792 gnd.n3791 585
R9787 gnd.n3794 gnd.n3793 585
R9788 gnd.n3796 gnd.n3795 585
R9789 gnd.n3798 gnd.n3797 585
R9790 gnd.n3800 gnd.n3799 585
R9791 gnd.n3802 gnd.n3801 585
R9792 gnd.n3804 gnd.n3803 585
R9793 gnd.n3806 gnd.n3805 585
R9794 gnd.n3808 gnd.n3807 585
R9795 gnd.n3810 gnd.n3809 585
R9796 gnd.n3812 gnd.n3811 585
R9797 gnd.n3814 gnd.n3813 585
R9798 gnd.n3816 gnd.n3815 585
R9799 gnd.n3818 gnd.n3817 585
R9800 gnd.n3820 gnd.n3819 585
R9801 gnd.n3821 gnd.n3757 585
R9802 gnd.n5478 gnd.n5477 585
R9803 gnd.n5480 gnd.n5479 585
R9804 gnd.n5482 gnd.n5481 585
R9805 gnd.n5484 gnd.n5483 585
R9806 gnd.n5486 gnd.n5485 585
R9807 gnd.n5488 gnd.n5487 585
R9808 gnd.n5490 gnd.n5489 585
R9809 gnd.n5492 gnd.n5491 585
R9810 gnd.n5494 gnd.n5493 585
R9811 gnd.n5496 gnd.n5495 585
R9812 gnd.n5498 gnd.n5497 585
R9813 gnd.n5500 gnd.n5499 585
R9814 gnd.n5502 gnd.n5501 585
R9815 gnd.n5504 gnd.n5503 585
R9816 gnd.n5506 gnd.n5505 585
R9817 gnd.n5508 gnd.n5507 585
R9818 gnd.n5510 gnd.n5509 585
R9819 gnd.n5512 gnd.n5511 585
R9820 gnd.n5514 gnd.n5513 585
R9821 gnd.n5516 gnd.n5515 585
R9822 gnd.n5518 gnd.n5517 585
R9823 gnd.n5520 gnd.n5519 585
R9824 gnd.n5522 gnd.n5521 585
R9825 gnd.n5524 gnd.n5523 585
R9826 gnd.n5526 gnd.n5525 585
R9827 gnd.n5528 gnd.n5527 585
R9828 gnd.n5530 gnd.n5529 585
R9829 gnd.n5532 gnd.n5531 585
R9830 gnd.n5534 gnd.n5533 585
R9831 gnd.n5536 gnd.n3335 585
R9832 gnd.n5538 gnd.n5537 585
R9833 gnd.n5540 gnd.n3299 585
R9834 gnd.n5542 gnd.n5541 585
R9835 gnd.n5545 gnd.n5544 585
R9836 gnd.n3302 gnd.n3300 585
R9837 gnd.n5411 gnd.n5410 585
R9838 gnd.n5413 gnd.n5412 585
R9839 gnd.n5416 gnd.n5415 585
R9840 gnd.n5418 gnd.n5417 585
R9841 gnd.n5420 gnd.n5419 585
R9842 gnd.n5422 gnd.n5421 585
R9843 gnd.n5424 gnd.n5423 585
R9844 gnd.n5426 gnd.n5425 585
R9845 gnd.n5428 gnd.n5427 585
R9846 gnd.n5430 gnd.n5429 585
R9847 gnd.n5432 gnd.n5431 585
R9848 gnd.n5434 gnd.n5433 585
R9849 gnd.n5436 gnd.n5435 585
R9850 gnd.n5438 gnd.n5437 585
R9851 gnd.n5440 gnd.n5439 585
R9852 gnd.n5442 gnd.n5441 585
R9853 gnd.n5444 gnd.n5443 585
R9854 gnd.n5446 gnd.n5445 585
R9855 gnd.n5448 gnd.n5447 585
R9856 gnd.n5450 gnd.n5449 585
R9857 gnd.n5452 gnd.n5451 585
R9858 gnd.n5454 gnd.n5453 585
R9859 gnd.n5456 gnd.n5455 585
R9860 gnd.n5458 gnd.n5457 585
R9861 gnd.n5460 gnd.n5459 585
R9862 gnd.n5462 gnd.n5461 585
R9863 gnd.n5464 gnd.n5463 585
R9864 gnd.n5466 gnd.n5465 585
R9865 gnd.n5468 gnd.n5467 585
R9866 gnd.n5470 gnd.n5469 585
R9867 gnd.n5471 gnd.n3342 585
R9868 gnd.n5476 gnd.n3338 585
R9869 gnd.n5476 gnd.n5475 585
R9870 gnd.n3428 gnd.n3339 585
R9871 gnd.n3347 gnd.n3339 585
R9872 gnd.n3429 gnd.n3346 585
R9873 gnd.n5385 gnd.n3346 585
R9874 gnd.n3431 gnd.n3430 585
R9875 gnd.n3434 gnd.n3431 585
R9876 gnd.n3439 gnd.n3438 585
R9877 gnd.n3438 gnd.n3437 585
R9878 gnd.n3440 gnd.n3369 585
R9879 gnd.n5179 gnd.n3369 585
R9880 gnd.n3441 gnd.n3376 585
R9881 gnd.n5170 gnd.n3376 585
R9882 gnd.n3442 gnd.n3375 585
R9883 gnd.n5172 gnd.n3375 585
R9884 gnd.n3443 gnd.n3384 585
R9885 gnd.n5157 gnd.n3384 585
R9886 gnd.n3445 gnd.n3444 585
R9887 gnd.n3444 gnd.n3383 585
R9888 gnd.n3446 gnd.n3391 585
R9889 gnd.n5146 gnd.n3391 585
R9890 gnd.n3448 gnd.n3447 585
R9891 gnd.n3447 gnd.n3390 585
R9892 gnd.n3449 gnd.n3399 585
R9893 gnd.n5139 gnd.n3399 585
R9894 gnd.n3453 gnd.n3452 585
R9895 gnd.n3452 gnd.n3451 585
R9896 gnd.n3454 gnd.n3406 585
R9897 gnd.n5129 gnd.n3406 585
R9898 gnd.n3456 gnd.n3455 585
R9899 gnd.n3455 gnd.n3405 585
R9900 gnd.n3457 gnd.n3412 585
R9901 gnd.n5123 gnd.n3412 585
R9902 gnd.n5099 gnd.n5098 585
R9903 gnd.n5098 gnd.n5097 585
R9904 gnd.n5100 gnd.n3421 585
R9905 gnd.n5111 gnd.n3421 585
R9906 gnd.n5102 gnd.n5101 585
R9907 gnd.n5103 gnd.n5102 585
R9908 gnd.n3427 gnd.n3426 585
R9909 gnd.n5105 gnd.n3426 585
R9910 gnd.n5082 gnd.n5081 585
R9911 gnd.n5083 gnd.n5082 585
R9912 gnd.n5080 gnd.n3465 585
R9913 gnd.n3465 gnd.n3463 585
R9914 gnd.n5079 gnd.n5078 585
R9915 gnd.n5078 gnd.n5077 585
R9916 gnd.n3467 gnd.n3466 585
R9917 gnd.n5034 gnd.n3467 585
R9918 gnd.n4976 gnd.n3474 585
R9919 gnd.n5070 gnd.n3474 585
R9920 gnd.n4979 gnd.n4978 585
R9921 gnd.n4978 gnd.n4977 585
R9922 gnd.n4980 gnd.n3482 585
R9923 gnd.n5056 gnd.n3482 585
R9924 gnd.n4982 gnd.n4981 585
R9925 gnd.n4981 gnd.n3480 585
R9926 gnd.n4983 gnd.n3488 585
R9927 gnd.n5050 gnd.n3488 585
R9928 gnd.n4986 gnd.n4985 585
R9929 gnd.n4985 gnd.n4984 585
R9930 gnd.n4987 gnd.n3496 585
R9931 gnd.n5026 gnd.n3496 585
R9932 gnd.n4989 gnd.n4988 585
R9933 gnd.n4988 gnd.n3495 585
R9934 gnd.n4990 gnd.n3501 585
R9935 gnd.n5020 gnd.n3501 585
R9936 gnd.n4994 gnd.n4993 585
R9937 gnd.n4993 gnd.n4992 585
R9938 gnd.n4995 gnd.n3509 585
R9939 gnd.n5006 gnd.n3509 585
R9940 gnd.n4997 gnd.n4996 585
R9941 gnd.n4998 gnd.n4997 585
R9942 gnd.n4975 gnd.n3514 585
R9943 gnd.n5000 gnd.n3514 585
R9944 gnd.n4974 gnd.n4973 585
R9945 gnd.n4973 gnd.n4972 585
R9946 gnd.n3516 gnd.n3515 585
R9947 gnd.n4940 gnd.n3516 585
R9948 gnd.n4924 gnd.n3524 585
R9949 gnd.n4958 gnd.n3524 585
R9950 gnd.n4926 gnd.n4925 585
R9951 gnd.n4925 gnd.n3532 585
R9952 gnd.n4927 gnd.n3531 585
R9953 gnd.n4951 gnd.n3531 585
R9954 gnd.n4929 gnd.n4928 585
R9955 gnd.n4930 gnd.n4929 585
R9956 gnd.n4923 gnd.n3541 585
R9957 gnd.n3541 gnd.n3539 585
R9958 gnd.n4922 gnd.n4921 585
R9959 gnd.n4921 gnd.n4920 585
R9960 gnd.n3543 gnd.n3542 585
R9961 gnd.n3551 gnd.n3543 585
R9962 gnd.n4823 gnd.n3550 585
R9963 gnd.n4913 gnd.n3550 585
R9964 gnd.n4826 gnd.n4825 585
R9965 gnd.n4825 gnd.n4824 585
R9966 gnd.n4827 gnd.n3560 585
R9967 gnd.n4902 gnd.n3560 585
R9968 gnd.n4829 gnd.n4828 585
R9969 gnd.n4828 gnd.n3558 585
R9970 gnd.n4830 gnd.n3566 585
R9971 gnd.n4896 gnd.n3566 585
R9972 gnd.n4834 gnd.n4833 585
R9973 gnd.n4833 gnd.n4832 585
R9974 gnd.n4835 gnd.n3574 585
R9975 gnd.n4871 gnd.n3574 585
R9976 gnd.n4837 gnd.n4836 585
R9977 gnd.n4836 gnd.n3573 585
R9978 gnd.n4838 gnd.n3580 585
R9979 gnd.n4865 gnd.n3580 585
R9980 gnd.n4841 gnd.n4840 585
R9981 gnd.n4840 gnd.n4839 585
R9982 gnd.n4842 gnd.n3588 585
R9983 gnd.n4853 gnd.n3588 585
R9984 gnd.n4844 gnd.n4843 585
R9985 gnd.n4845 gnd.n4844 585
R9986 gnd.n4822 gnd.n3595 585
R9987 gnd.n4847 gnd.n3595 585
R9988 gnd.n4821 gnd.n4820 585
R9989 gnd.n4820 gnd.n4819 585
R9990 gnd.n3597 gnd.n3596 585
R9991 gnd.n4803 gnd.n3597 585
R9992 gnd.n4800 gnd.n4799 585
R9993 gnd.n4801 gnd.n4800 585
R9994 gnd.n4798 gnd.n3605 585
R9995 gnd.n4809 gnd.n3605 585
R9996 gnd.n4797 gnd.n4796 585
R9997 gnd.n4796 gnd.n4795 585
R9998 gnd.n3612 gnd.n3611 585
R9999 gnd.n4793 gnd.n3612 585
R10000 gnd.n4770 gnd.n4769 585
R10001 gnd.n4769 gnd.n3619 585
R10002 gnd.n4771 gnd.n3617 585
R10003 gnd.n4787 gnd.n3617 585
R10004 gnd.n4773 gnd.n4772 585
R10005 gnd.n4774 gnd.n4773 585
R10006 gnd.n4768 gnd.n3627 585
R10007 gnd.n3627 gnd.n3625 585
R10008 gnd.n4767 gnd.n4766 585
R10009 gnd.n4766 gnd.n4765 585
R10010 gnd.n3629 gnd.n3628 585
R10011 gnd.n3638 gnd.n3629 585
R10012 gnd.n4644 gnd.n3637 585
R10013 gnd.n4758 gnd.n3637 585
R10014 gnd.n4647 gnd.n4646 585
R10015 gnd.n4646 gnd.n4645 585
R10016 gnd.n4648 gnd.n3647 585
R10017 gnd.n4746 gnd.n3647 585
R10018 gnd.n4650 gnd.n4649 585
R10019 gnd.n4649 gnd.n3645 585
R10020 gnd.n4651 gnd.n3653 585
R10021 gnd.n4740 gnd.n3653 585
R10022 gnd.n4655 gnd.n4654 585
R10023 gnd.n4654 gnd.n4653 585
R10024 gnd.n4656 gnd.n3660 585
R10025 gnd.n4694 gnd.n3660 585
R10026 gnd.n4658 gnd.n4657 585
R10027 gnd.n4657 gnd.n3666 585
R10028 gnd.n4659 gnd.n3665 585
R10029 gnd.n4688 gnd.n3665 585
R10030 gnd.n4663 gnd.n4662 585
R10031 gnd.n4662 gnd.n4661 585
R10032 gnd.n4664 gnd.n3674 585
R10033 gnd.n4675 gnd.n3674 585
R10034 gnd.n4666 gnd.n4665 585
R10035 gnd.n4667 gnd.n4666 585
R10036 gnd.n4643 gnd.n3680 585
R10037 gnd.n4669 gnd.n3680 585
R10038 gnd.n4642 gnd.n4641 585
R10039 gnd.n4641 gnd.n4640 585
R10040 gnd.n3682 gnd.n3681 585
R10041 gnd.n4624 gnd.n3682 585
R10042 gnd.n4574 gnd.n4573 585
R10043 gnd.n4573 gnd.n4572 585
R10044 gnd.n4575 gnd.n3689 585
R10045 gnd.n4630 gnd.n3689 585
R10046 gnd.n4578 gnd.n4577 585
R10047 gnd.n4577 gnd.n4576 585
R10048 gnd.n4579 gnd.n3701 585
R10049 gnd.n4605 gnd.n3701 585
R10050 gnd.n4581 gnd.n4580 585
R10051 gnd.n4580 gnd.n3707 585
R10052 gnd.n4582 gnd.n3706 585
R10053 gnd.n4599 gnd.n3706 585
R10054 gnd.n4584 gnd.n4583 585
R10055 gnd.n4586 gnd.n4584 585
R10056 gnd.n4571 gnd.n3715 585
R10057 gnd.n3715 gnd.n3713 585
R10058 gnd.n4570 gnd.n4569 585
R10059 gnd.n4569 gnd.n4568 585
R10060 gnd.n3717 gnd.n3716 585
R10061 gnd.n4554 gnd.n3717 585
R10062 gnd.n4523 gnd.n3725 585
R10063 gnd.n4561 gnd.n3725 585
R10064 gnd.n4527 gnd.n4524 585
R10065 gnd.n4527 gnd.n4526 585
R10066 gnd.n4529 gnd.n4528 585
R10067 gnd.n4528 gnd.n2942 585
R10068 gnd.n4530 gnd.n3736 585
R10069 gnd.n3736 gnd.n2940 585
R10070 gnd.n4532 gnd.n4531 585
R10071 gnd.n4539 gnd.n4532 585
R10072 gnd.n4522 gnd.n3735 585
R10073 gnd.n3735 gnd.n3734 585
R10074 gnd.n4521 gnd.n2931 585
R10075 gnd.n6136 gnd.n2931 585
R10076 gnd.n4520 gnd.n4519 585
R10077 gnd.n4519 gnd.n4518 585
R10078 gnd.n3737 gnd.n2922 585
R10079 gnd.n6142 gnd.n2922 585
R10080 gnd.n4506 gnd.n4505 585
R10081 gnd.n4507 gnd.n4506 585
R10082 gnd.n4504 gnd.n3749 585
R10083 gnd.n3749 gnd.n3747 585
R10084 gnd.n4503 gnd.n4502 585
R10085 gnd.n4502 gnd.n4501 585
R10086 gnd.n3750 gnd.n2913 585
R10087 gnd.n6150 gnd.n2913 585
R10088 gnd.n3823 gnd.n3822 585
R10089 gnd.n3824 gnd.n3823 585
R10090 gnd.n6359 gnd.n6358 585
R10091 gnd.n6358 gnd.n6357 585
R10092 gnd.n6360 gnd.n2565 585
R10093 gnd.n6350 gnd.n2565 585
R10094 gnd.n6362 gnd.n6361 585
R10095 gnd.n6363 gnd.n6362 585
R10096 gnd.n2550 gnd.n2549 585
R10097 gnd.n4425 gnd.n2550 585
R10098 gnd.n6371 gnd.n6370 585
R10099 gnd.n6370 gnd.n6369 585
R10100 gnd.n6372 gnd.n2544 585
R10101 gnd.n4419 gnd.n2544 585
R10102 gnd.n6374 gnd.n6373 585
R10103 gnd.n6375 gnd.n6374 585
R10104 gnd.n2530 gnd.n2529 585
R10105 gnd.n4436 gnd.n2530 585
R10106 gnd.n6383 gnd.n6382 585
R10107 gnd.n6382 gnd.n6381 585
R10108 gnd.n6384 gnd.n2524 585
R10109 gnd.n4412 gnd.n2524 585
R10110 gnd.n6386 gnd.n6385 585
R10111 gnd.n6387 gnd.n6386 585
R10112 gnd.n2510 gnd.n2509 585
R10113 gnd.n4404 gnd.n2510 585
R10114 gnd.n6395 gnd.n6394 585
R10115 gnd.n6394 gnd.n6393 585
R10116 gnd.n6396 gnd.n2504 585
R10117 gnd.n4398 gnd.n2504 585
R10118 gnd.n6398 gnd.n6397 585
R10119 gnd.n6399 gnd.n6398 585
R10120 gnd.n2490 gnd.n2489 585
R10121 gnd.n4390 gnd.n2490 585
R10122 gnd.n6407 gnd.n6406 585
R10123 gnd.n6406 gnd.n6405 585
R10124 gnd.n6408 gnd.n2487 585
R10125 gnd.n4341 gnd.n2487 585
R10126 gnd.n6411 gnd.n6410 585
R10127 gnd.n6412 gnd.n6411 585
R10128 gnd.n2488 gnd.n2473 585
R10129 gnd.n4332 gnd.n2473 585
R10130 gnd.n6420 gnd.n6419 585
R10131 gnd.n6419 gnd.n6418 585
R10132 gnd.n6421 gnd.n2470 585
R10133 gnd.n4317 gnd.n2470 585
R10134 gnd.n6424 gnd.n6423 585
R10135 gnd.n6425 gnd.n6424 585
R10136 gnd.n2471 gnd.n2456 585
R10137 gnd.n4354 gnd.n2456 585
R10138 gnd.n6433 gnd.n6432 585
R10139 gnd.n6432 gnd.n6431 585
R10140 gnd.n6434 gnd.n2452 585
R10141 gnd.n4310 gnd.n2452 585
R10142 gnd.n6437 gnd.n6436 585
R10143 gnd.n6438 gnd.n6437 585
R10144 gnd.n2437 gnd.n2436 585
R10145 gnd.n4301 gnd.n2437 585
R10146 gnd.n6446 gnd.n6445 585
R10147 gnd.n6445 gnd.n6444 585
R10148 gnd.n6447 gnd.n2431 585
R10149 gnd.n4295 gnd.n2431 585
R10150 gnd.n6449 gnd.n6448 585
R10151 gnd.n6450 gnd.n6449 585
R10152 gnd.n2417 gnd.n2416 585
R10153 gnd.n4287 gnd.n2417 585
R10154 gnd.n6458 gnd.n6457 585
R10155 gnd.n6457 gnd.n6456 585
R10156 gnd.n6459 gnd.n2411 585
R10157 gnd.n4232 gnd.n2411 585
R10158 gnd.n6461 gnd.n6460 585
R10159 gnd.n6462 gnd.n6461 585
R10160 gnd.n2396 gnd.n2395 585
R10161 gnd.n4238 gnd.n2396 585
R10162 gnd.n6470 gnd.n6469 585
R10163 gnd.n6469 gnd.n6468 585
R10164 gnd.n6471 gnd.n2390 585
R10165 gnd.n4244 gnd.n2390 585
R10166 gnd.n6473 gnd.n6472 585
R10167 gnd.n6474 gnd.n6473 585
R10168 gnd.n2374 gnd.n2373 585
R10169 gnd.n4250 gnd.n2374 585
R10170 gnd.n6482 gnd.n6481 585
R10171 gnd.n6481 gnd.n6480 585
R10172 gnd.n6483 gnd.n2369 585
R10173 gnd.n4256 gnd.n2369 585
R10174 gnd.n6485 gnd.n6484 585
R10175 gnd.n6486 gnd.n6485 585
R10176 gnd.n4063 gnd.n2368 585
R10177 gnd.n4066 gnd.n4065 585
R10178 gnd.n4061 gnd.n4060 585
R10179 gnd.n4060 gnd.n2363 585
R10180 gnd.n4071 gnd.n4070 585
R10181 gnd.n4073 gnd.n4059 585
R10182 gnd.n4076 gnd.n4075 585
R10183 gnd.n4057 gnd.n4056 585
R10184 gnd.n4081 gnd.n4080 585
R10185 gnd.n4083 gnd.n4055 585
R10186 gnd.n4086 gnd.n4085 585
R10187 gnd.n4053 gnd.n4052 585
R10188 gnd.n4091 gnd.n4090 585
R10189 gnd.n4093 gnd.n4051 585
R10190 gnd.n4096 gnd.n4095 585
R10191 gnd.n4049 gnd.n4048 585
R10192 gnd.n4101 gnd.n4100 585
R10193 gnd.n4103 gnd.n4044 585
R10194 gnd.n4106 gnd.n4105 585
R10195 gnd.n4042 gnd.n4041 585
R10196 gnd.n4111 gnd.n4110 585
R10197 gnd.n4113 gnd.n4040 585
R10198 gnd.n4116 gnd.n4115 585
R10199 gnd.n4038 gnd.n4037 585
R10200 gnd.n4121 gnd.n4120 585
R10201 gnd.n4123 gnd.n4036 585
R10202 gnd.n4126 gnd.n4125 585
R10203 gnd.n4034 gnd.n4033 585
R10204 gnd.n4131 gnd.n4130 585
R10205 gnd.n4133 gnd.n4032 585
R10206 gnd.n4136 gnd.n4135 585
R10207 gnd.n4030 gnd.n4029 585
R10208 gnd.n4141 gnd.n4140 585
R10209 gnd.n4143 gnd.n4028 585
R10210 gnd.n4146 gnd.n4145 585
R10211 gnd.n4026 gnd.n4025 585
R10212 gnd.n4151 gnd.n4150 585
R10213 gnd.n4153 gnd.n4024 585
R10214 gnd.n4158 gnd.n4155 585
R10215 gnd.n4022 gnd.n4021 585
R10216 gnd.n4163 gnd.n4162 585
R10217 gnd.n4165 gnd.n4020 585
R10218 gnd.n4168 gnd.n4167 585
R10219 gnd.n4018 gnd.n4017 585
R10220 gnd.n4173 gnd.n4172 585
R10221 gnd.n4175 gnd.n4016 585
R10222 gnd.n4178 gnd.n4177 585
R10223 gnd.n4014 gnd.n4013 585
R10224 gnd.n4183 gnd.n4182 585
R10225 gnd.n4185 gnd.n4012 585
R10226 gnd.n4188 gnd.n4187 585
R10227 gnd.n4010 gnd.n4009 585
R10228 gnd.n4193 gnd.n4192 585
R10229 gnd.n4195 gnd.n4008 585
R10230 gnd.n4198 gnd.n4197 585
R10231 gnd.n4006 gnd.n4005 585
R10232 gnd.n4204 gnd.n4203 585
R10233 gnd.n4206 gnd.n4004 585
R10234 gnd.n4207 gnd.n4003 585
R10235 gnd.n4210 gnd.n4209 585
R10236 gnd.n2781 gnd.n2780 585
R10237 gnd.n2787 gnd.n2786 585
R10238 gnd.n2789 gnd.n2788 585
R10239 gnd.n2791 gnd.n2790 585
R10240 gnd.n2793 gnd.n2792 585
R10241 gnd.n2795 gnd.n2794 585
R10242 gnd.n2797 gnd.n2796 585
R10243 gnd.n2799 gnd.n2798 585
R10244 gnd.n2801 gnd.n2800 585
R10245 gnd.n2803 gnd.n2802 585
R10246 gnd.n2805 gnd.n2804 585
R10247 gnd.n2807 gnd.n2806 585
R10248 gnd.n2809 gnd.n2808 585
R10249 gnd.n2811 gnd.n2810 585
R10250 gnd.n2813 gnd.n2812 585
R10251 gnd.n2815 gnd.n2814 585
R10252 gnd.n2817 gnd.n2816 585
R10253 gnd.n2819 gnd.n2818 585
R10254 gnd.n2821 gnd.n2820 585
R10255 gnd.n2824 gnd.n2823 585
R10256 gnd.n2822 gnd.n2760 585
R10257 gnd.n2829 gnd.n2828 585
R10258 gnd.n2831 gnd.n2830 585
R10259 gnd.n2833 gnd.n2832 585
R10260 gnd.n2835 gnd.n2834 585
R10261 gnd.n2837 gnd.n2836 585
R10262 gnd.n2839 gnd.n2838 585
R10263 gnd.n2841 gnd.n2840 585
R10264 gnd.n2843 gnd.n2842 585
R10265 gnd.n2846 gnd.n2845 585
R10266 gnd.n2844 gnd.n2751 585
R10267 gnd.n6226 gnd.n6225 585
R10268 gnd.n6228 gnd.n6227 585
R10269 gnd.n6230 gnd.n6229 585
R10270 gnd.n6232 gnd.n6231 585
R10271 gnd.n6234 gnd.n6233 585
R10272 gnd.n6236 gnd.n6235 585
R10273 gnd.n6238 gnd.n6237 585
R10274 gnd.n6240 gnd.n6239 585
R10275 gnd.n6243 gnd.n6242 585
R10276 gnd.n6245 gnd.n6244 585
R10277 gnd.n6247 gnd.n6246 585
R10278 gnd.n6249 gnd.n6248 585
R10279 gnd.n6251 gnd.n6250 585
R10280 gnd.n6253 gnd.n6252 585
R10281 gnd.n6255 gnd.n6254 585
R10282 gnd.n6257 gnd.n6256 585
R10283 gnd.n6259 gnd.n6258 585
R10284 gnd.n6261 gnd.n6260 585
R10285 gnd.n6263 gnd.n6262 585
R10286 gnd.n6265 gnd.n6264 585
R10287 gnd.n6267 gnd.n6266 585
R10288 gnd.n6269 gnd.n6268 585
R10289 gnd.n6270 gnd.n2720 585
R10290 gnd.n6272 gnd.n6271 585
R10291 gnd.n2721 gnd.n2719 585
R10292 gnd.n2722 gnd.n2570 585
R10293 gnd.n6274 gnd.n2570 585
R10294 gnd.n6353 gnd.n2572 585
R10295 gnd.n6357 gnd.n2572 585
R10296 gnd.n6352 gnd.n6351 585
R10297 gnd.n6351 gnd.n6350 585
R10298 gnd.n2578 gnd.n2562 585
R10299 gnd.n6363 gnd.n2562 585
R10300 gnd.n4424 gnd.n4423 585
R10301 gnd.n4425 gnd.n4424 585
R10302 gnd.n4422 gnd.n2552 585
R10303 gnd.n6369 gnd.n2552 585
R10304 gnd.n4421 gnd.n4420 585
R10305 gnd.n4420 gnd.n4419 585
R10306 gnd.n4417 gnd.n2541 585
R10307 gnd.n6375 gnd.n2541 585
R10308 gnd.n4416 gnd.n3857 585
R10309 gnd.n4436 gnd.n3857 585
R10310 gnd.n4415 gnd.n2532 585
R10311 gnd.n6381 gnd.n2532 585
R10312 gnd.n4414 gnd.n4413 585
R10313 gnd.n4413 gnd.n4412 585
R10314 gnd.n3863 gnd.n2521 585
R10315 gnd.n6387 gnd.n2521 585
R10316 gnd.n4403 gnd.n4402 585
R10317 gnd.n4404 gnd.n4403 585
R10318 gnd.n4401 gnd.n2512 585
R10319 gnd.n6393 gnd.n2512 585
R10320 gnd.n4400 gnd.n4399 585
R10321 gnd.n4399 gnd.n4398 585
R10322 gnd.n3869 gnd.n2501 585
R10323 gnd.n6399 gnd.n2501 585
R10324 gnd.n4337 gnd.n3874 585
R10325 gnd.n4390 gnd.n3874 585
R10326 gnd.n4338 gnd.n2492 585
R10327 gnd.n6405 gnd.n2492 585
R10328 gnd.n4340 gnd.n4339 585
R10329 gnd.n4341 gnd.n4340 585
R10330 gnd.n4335 gnd.n2484 585
R10331 gnd.n6412 gnd.n2484 585
R10332 gnd.n4334 gnd.n4333 585
R10333 gnd.n4333 gnd.n4332 585
R10334 gnd.n4320 gnd.n2475 585
R10335 gnd.n6418 gnd.n2475 585
R10336 gnd.n4319 gnd.n4318 585
R10337 gnd.n4318 gnd.n4317 585
R10338 gnd.n4315 gnd.n2467 585
R10339 gnd.n6425 gnd.n2467 585
R10340 gnd.n4314 gnd.n3890 585
R10341 gnd.n4354 gnd.n3890 585
R10342 gnd.n4313 gnd.n2458 585
R10343 gnd.n6431 gnd.n2458 585
R10344 gnd.n4312 gnd.n4311 585
R10345 gnd.n4311 gnd.n4310 585
R10346 gnd.n3898 gnd.n2449 585
R10347 gnd.n6438 gnd.n2449 585
R10348 gnd.n4300 gnd.n4299 585
R10349 gnd.n4301 gnd.n4300 585
R10350 gnd.n4298 gnd.n2439 585
R10351 gnd.n6444 gnd.n2439 585
R10352 gnd.n4297 gnd.n4296 585
R10353 gnd.n4296 gnd.n4295 585
R10354 gnd.n3903 gnd.n2428 585
R10355 gnd.n6450 gnd.n2428 585
R10356 gnd.n4226 gnd.n3908 585
R10357 gnd.n4287 gnd.n3908 585
R10358 gnd.n4227 gnd.n2419 585
R10359 gnd.n6456 gnd.n2419 585
R10360 gnd.n4234 gnd.n4233 585
R10361 gnd.n4233 gnd.n4232 585
R10362 gnd.n4235 gnd.n2408 585
R10363 gnd.n6462 gnd.n2408 585
R10364 gnd.n4237 gnd.n4236 585
R10365 gnd.n4238 gnd.n4237 585
R10366 gnd.n4219 gnd.n2398 585
R10367 gnd.n6468 gnd.n2398 585
R10368 gnd.n4246 gnd.n4245 585
R10369 gnd.n4245 gnd.n4244 585
R10370 gnd.n4247 gnd.n2387 585
R10371 gnd.n6474 gnd.n2387 585
R10372 gnd.n4249 gnd.n4248 585
R10373 gnd.n4250 gnd.n4249 585
R10374 gnd.n4217 gnd.n2375 585
R10375 gnd.n6480 gnd.n2375 585
R10376 gnd.n4216 gnd.n3924 585
R10377 gnd.n4256 gnd.n3924 585
R10378 gnd.n3930 gnd.n2364 585
R10379 gnd.n6486 gnd.n2364 585
R10380 gnd.n7677 gnd.n7676 585
R10381 gnd.n7676 gnd.n7675 585
R10382 gnd.n7678 gnd.n162 585
R10383 gnd.n7668 gnd.n162 585
R10384 gnd.n7680 gnd.n7679 585
R10385 gnd.n7681 gnd.n7680 585
R10386 gnd.n148 gnd.n147 585
R10387 gnd.n5889 gnd.n148 585
R10388 gnd.n7689 gnd.n7688 585
R10389 gnd.n7688 gnd.n7687 585
R10390 gnd.n7690 gnd.n142 585
R10391 gnd.n5895 gnd.n142 585
R10392 gnd.n7692 gnd.n7691 585
R10393 gnd.n7693 gnd.n7692 585
R10394 gnd.n127 gnd.n126 585
R10395 gnd.n5901 gnd.n127 585
R10396 gnd.n7701 gnd.n7700 585
R10397 gnd.n7700 gnd.n7699 585
R10398 gnd.n7702 gnd.n121 585
R10399 gnd.n5907 gnd.n121 585
R10400 gnd.n7704 gnd.n7703 585
R10401 gnd.n7705 gnd.n7704 585
R10402 gnd.n107 gnd.n106 585
R10403 gnd.n5913 gnd.n107 585
R10404 gnd.n7713 gnd.n7712 585
R10405 gnd.n7712 gnd.n7711 585
R10406 gnd.n7714 gnd.n102 585
R10407 gnd.n5870 gnd.n102 585
R10408 gnd.n7716 gnd.n7715 585
R10409 gnd.n7717 gnd.n7716 585
R10410 gnd.n85 gnd.n83 585
R10411 gnd.n5861 gnd.n85 585
R10412 gnd.n7725 gnd.n7724 585
R10413 gnd.n7724 gnd.n7723 585
R10414 gnd.n84 gnd.n76 585
R10415 gnd.n5855 gnd.n84 585
R10416 gnd.n7728 gnd.n74 585
R10417 gnd.n5928 gnd.n74 585
R10418 gnd.n7730 gnd.n7729 585
R10419 gnd.n7731 gnd.n7730 585
R10420 gnd.n3162 gnd.n73 585
R10421 gnd.n5845 gnd.n73 585
R10422 gnd.n5936 gnd.n3163 585
R10423 gnd.n5936 gnd.n5935 585
R10424 gnd.n5939 gnd.n5938 585
R10425 gnd.n5940 gnd.n5939 585
R10426 gnd.n5937 gnd.n3161 585
R10427 gnd.n3161 gnd.n3156 585
R10428 gnd.n3145 gnd.n3144 585
R10429 gnd.n3149 gnd.n3144 585
R10430 gnd.n5950 gnd.n3146 585
R10431 gnd.n5950 gnd.n5949 585
R10432 gnd.n5952 gnd.n5951 585
R10433 gnd.n5953 gnd.n5952 585
R10434 gnd.n3130 gnd.n3129 585
R10435 gnd.n5828 gnd.n3130 585
R10436 gnd.n5961 gnd.n5960 585
R10437 gnd.n5960 gnd.n5959 585
R10438 gnd.n5962 gnd.n3124 585
R10439 gnd.n5810 gnd.n3124 585
R10440 gnd.n5964 gnd.n5963 585
R10441 gnd.n5965 gnd.n5964 585
R10442 gnd.n3110 gnd.n3109 585
R10443 gnd.n5803 gnd.n3110 585
R10444 gnd.n5973 gnd.n5972 585
R10445 gnd.n5972 gnd.n5971 585
R10446 gnd.n5974 gnd.n3104 585
R10447 gnd.n5747 gnd.n3104 585
R10448 gnd.n5976 gnd.n5975 585
R10449 gnd.n5977 gnd.n5976 585
R10450 gnd.n3090 gnd.n3089 585
R10451 gnd.n5758 gnd.n3090 585
R10452 gnd.n5985 gnd.n5984 585
R10453 gnd.n5984 gnd.n5983 585
R10454 gnd.n5986 gnd.n3084 585
R10455 gnd.n5738 gnd.n3084 585
R10456 gnd.n5988 gnd.n5987 585
R10457 gnd.n5989 gnd.n5988 585
R10458 gnd.n3067 gnd.n3066 585
R10459 gnd.n5730 gnd.n3067 585
R10460 gnd.n5997 gnd.n5996 585
R10461 gnd.n5996 gnd.n5995 585
R10462 gnd.n5998 gnd.n3062 585
R10463 gnd.n5195 gnd.n3062 585
R10464 gnd.n6000 gnd.n5999 585
R10465 gnd.n6001 gnd.n6000 585
R10466 gnd.n5571 gnd.n3061 585
R10467 gnd.n5576 gnd.n5574 585
R10468 gnd.n5577 gnd.n5570 585
R10469 gnd.n5577 gnd.n3048 585
R10470 gnd.n5580 gnd.n5579 585
R10471 gnd.n5568 gnd.n5567 585
R10472 gnd.n5585 gnd.n5584 585
R10473 gnd.n5587 gnd.n5566 585
R10474 gnd.n5590 gnd.n5589 585
R10475 gnd.n5564 gnd.n5563 585
R10476 gnd.n5595 gnd.n5594 585
R10477 gnd.n5597 gnd.n5562 585
R10478 gnd.n5600 gnd.n5599 585
R10479 gnd.n5560 gnd.n5559 585
R10480 gnd.n5605 gnd.n5604 585
R10481 gnd.n5607 gnd.n5558 585
R10482 gnd.n5610 gnd.n5609 585
R10483 gnd.n5556 gnd.n5555 585
R10484 gnd.n5618 gnd.n5617 585
R10485 gnd.n5620 gnd.n5554 585
R10486 gnd.n5623 gnd.n5622 585
R10487 gnd.n5552 gnd.n5551 585
R10488 gnd.n5628 gnd.n5627 585
R10489 gnd.n5630 gnd.n5550 585
R10490 gnd.n5633 gnd.n5632 585
R10491 gnd.n5548 gnd.n5547 585
R10492 gnd.n5639 gnd.n5638 585
R10493 gnd.n5643 gnd.n3298 585
R10494 gnd.n5646 gnd.n5645 585
R10495 gnd.n3296 gnd.n3295 585
R10496 gnd.n5651 gnd.n5650 585
R10497 gnd.n5653 gnd.n3294 585
R10498 gnd.n5656 gnd.n5655 585
R10499 gnd.n3292 gnd.n3291 585
R10500 gnd.n5661 gnd.n5660 585
R10501 gnd.n5663 gnd.n3290 585
R10502 gnd.n5668 gnd.n5665 585
R10503 gnd.n3288 gnd.n3287 585
R10504 gnd.n5673 gnd.n5672 585
R10505 gnd.n5675 gnd.n3286 585
R10506 gnd.n5678 gnd.n5677 585
R10507 gnd.n3284 gnd.n3283 585
R10508 gnd.n5683 gnd.n5682 585
R10509 gnd.n5685 gnd.n3282 585
R10510 gnd.n5688 gnd.n5687 585
R10511 gnd.n3280 gnd.n3279 585
R10512 gnd.n5693 gnd.n5692 585
R10513 gnd.n5695 gnd.n3278 585
R10514 gnd.n5698 gnd.n5697 585
R10515 gnd.n3276 gnd.n3275 585
R10516 gnd.n5703 gnd.n5702 585
R10517 gnd.n5705 gnd.n3274 585
R10518 gnd.n5708 gnd.n5707 585
R10519 gnd.n3272 gnd.n3271 585
R10520 gnd.n5714 gnd.n5713 585
R10521 gnd.n5716 gnd.n3270 585
R10522 gnd.n5717 gnd.n3269 585
R10523 gnd.n5720 gnd.n5719 585
R10524 gnd.n7537 gnd.n7536 585
R10525 gnd.n7543 gnd.n7542 585
R10526 gnd.n7545 gnd.n7544 585
R10527 gnd.n7547 gnd.n7546 585
R10528 gnd.n7549 gnd.n7548 585
R10529 gnd.n7551 gnd.n7550 585
R10530 gnd.n7553 gnd.n7552 585
R10531 gnd.n7555 gnd.n7554 585
R10532 gnd.n7557 gnd.n7556 585
R10533 gnd.n7559 gnd.n7558 585
R10534 gnd.n7561 gnd.n7560 585
R10535 gnd.n7563 gnd.n7562 585
R10536 gnd.n7565 gnd.n7564 585
R10537 gnd.n7567 gnd.n7566 585
R10538 gnd.n7569 gnd.n7568 585
R10539 gnd.n7571 gnd.n7570 585
R10540 gnd.n7573 gnd.n7572 585
R10541 gnd.n7575 gnd.n7574 585
R10542 gnd.n7577 gnd.n7576 585
R10543 gnd.n7580 gnd.n7579 585
R10544 gnd.n7578 gnd.n7516 585
R10545 gnd.n7585 gnd.n7584 585
R10546 gnd.n7587 gnd.n7586 585
R10547 gnd.n7589 gnd.n7588 585
R10548 gnd.n7591 gnd.n7590 585
R10549 gnd.n7593 gnd.n7592 585
R10550 gnd.n7595 gnd.n7594 585
R10551 gnd.n7597 gnd.n7596 585
R10552 gnd.n7599 gnd.n7598 585
R10553 gnd.n7601 gnd.n7600 585
R10554 gnd.n7603 gnd.n7602 585
R10555 gnd.n7605 gnd.n7604 585
R10556 gnd.n7607 gnd.n7606 585
R10557 gnd.n7609 gnd.n7608 585
R10558 gnd.n7611 gnd.n7610 585
R10559 gnd.n7613 gnd.n7612 585
R10560 gnd.n7615 gnd.n7614 585
R10561 gnd.n7617 gnd.n7616 585
R10562 gnd.n7619 gnd.n7618 585
R10563 gnd.n7621 gnd.n7620 585
R10564 gnd.n7623 gnd.n7622 585
R10565 gnd.n7628 gnd.n7627 585
R10566 gnd.n7630 gnd.n7629 585
R10567 gnd.n7632 gnd.n7631 585
R10568 gnd.n7634 gnd.n7633 585
R10569 gnd.n7636 gnd.n7635 585
R10570 gnd.n7638 gnd.n7637 585
R10571 gnd.n7640 gnd.n7639 585
R10572 gnd.n7642 gnd.n7641 585
R10573 gnd.n7644 gnd.n7643 585
R10574 gnd.n7646 gnd.n7645 585
R10575 gnd.n7648 gnd.n7647 585
R10576 gnd.n7650 gnd.n7649 585
R10577 gnd.n7652 gnd.n7651 585
R10578 gnd.n7654 gnd.n7653 585
R10579 gnd.n7655 gnd.n7476 585
R10580 gnd.n7657 gnd.n7656 585
R10581 gnd.n7477 gnd.n7475 585
R10582 gnd.n7478 gnd.n167 585
R10583 gnd.n7659 gnd.n167 585
R10584 gnd.n7671 gnd.n169 585
R10585 gnd.n7675 gnd.n169 585
R10586 gnd.n7670 gnd.n7669 585
R10587 gnd.n7669 gnd.n7668 585
R10588 gnd.n175 gnd.n160 585
R10589 gnd.n7681 gnd.n160 585
R10590 gnd.n5891 gnd.n5890 585
R10591 gnd.n5890 gnd.n5889 585
R10592 gnd.n5892 gnd.n150 585
R10593 gnd.n7687 gnd.n150 585
R10594 gnd.n5894 gnd.n5893 585
R10595 gnd.n5895 gnd.n5894 585
R10596 gnd.n5877 gnd.n139 585
R10597 gnd.n7693 gnd.n139 585
R10598 gnd.n5903 gnd.n5902 585
R10599 gnd.n5902 gnd.n5901 585
R10600 gnd.n5904 gnd.n129 585
R10601 gnd.n7699 gnd.n129 585
R10602 gnd.n5906 gnd.n5905 585
R10603 gnd.n5907 gnd.n5906 585
R10604 gnd.n5875 gnd.n118 585
R10605 gnd.n7705 gnd.n118 585
R10606 gnd.n5874 gnd.n3227 585
R10607 gnd.n5913 gnd.n3227 585
R10608 gnd.n5873 gnd.n109 585
R10609 gnd.n7711 gnd.n109 585
R10610 gnd.n5872 gnd.n5871 585
R10611 gnd.n5871 gnd.n5870 585
R10612 gnd.n3233 gnd.n99 585
R10613 gnd.n7717 gnd.n99 585
R10614 gnd.n5860 gnd.n5859 585
R10615 gnd.n5861 gnd.n5860 585
R10616 gnd.n5858 gnd.n87 585
R10617 gnd.n7723 gnd.n87 585
R10618 gnd.n5857 gnd.n5856 585
R10619 gnd.n5856 gnd.n5855 585
R10620 gnd.n5849 gnd.n3173 585
R10621 gnd.n5928 gnd.n3173 585
R10622 gnd.n5848 gnd.n70 585
R10623 gnd.n7731 gnd.n70 585
R10624 gnd.n5847 gnd.n5846 585
R10625 gnd.n5846 gnd.n5845 585
R10626 gnd.n5844 gnd.n3164 585
R10627 gnd.n5935 gnd.n3164 585
R10628 gnd.n5843 gnd.n3157 585
R10629 gnd.n5940 gnd.n3157 585
R10630 gnd.n5833 gnd.n3238 585
R10631 gnd.n5833 gnd.n3156 585
R10632 gnd.n5835 gnd.n5834 585
R10633 gnd.n5834 gnd.n3149 585
R10634 gnd.n5832 gnd.n3147 585
R10635 gnd.n5949 gnd.n3147 585
R10636 gnd.n5831 gnd.n3141 585
R10637 gnd.n5953 gnd.n3141 585
R10638 gnd.n5830 gnd.n5829 585
R10639 gnd.n5829 gnd.n5828 585
R10640 gnd.n3240 gnd.n3132 585
R10641 gnd.n5959 gnd.n3132 585
R10642 gnd.n5809 gnd.n5808 585
R10643 gnd.n5810 gnd.n5809 585
R10644 gnd.n5806 gnd.n3121 585
R10645 gnd.n5965 gnd.n3121 585
R10646 gnd.n5805 gnd.n5804 585
R10647 gnd.n5804 gnd.n5803 585
R10648 gnd.n3246 gnd.n3112 585
R10649 gnd.n5971 gnd.n3112 585
R10650 gnd.n5746 gnd.n5745 585
R10651 gnd.n5747 gnd.n5746 585
R10652 gnd.n5743 gnd.n3101 585
R10653 gnd.n5977 gnd.n3101 585
R10654 gnd.n5742 gnd.n3253 585
R10655 gnd.n5758 gnd.n3253 585
R10656 gnd.n5741 gnd.n3092 585
R10657 gnd.n5983 gnd.n3092 585
R10658 gnd.n5740 gnd.n5739 585
R10659 gnd.n5739 gnd.n5738 585
R10660 gnd.n3258 gnd.n3081 585
R10661 gnd.n5989 gnd.n3081 585
R10662 gnd.n5729 gnd.n5728 585
R10663 gnd.n5730 gnd.n5729 585
R10664 gnd.n5727 gnd.n3069 585
R10665 gnd.n5995 gnd.n3069 585
R10666 gnd.n5726 gnd.n3264 585
R10667 gnd.n5195 gnd.n3264 585
R10668 gnd.n3263 gnd.n3057 585
R10669 gnd.n6001 gnd.n3057 585
R10670 gnd.n6517 gnd.n871 585
R10671 gnd.n2339 gnd.n871 585
R10672 gnd.n7421 gnd.n7420 585
R10673 gnd.n7422 gnd.n7421 585
R10674 gnd.n267 gnd.n266 585
R10675 gnd.n7423 gnd.n267 585
R10676 gnd.n7426 gnd.n7425 585
R10677 gnd.n7425 gnd.n7424 585
R10678 gnd.n7427 gnd.n261 585
R10679 gnd.n261 gnd.n260 585
R10680 gnd.n7429 gnd.n7428 585
R10681 gnd.n7430 gnd.n7429 585
R10682 gnd.n259 gnd.n258 585
R10683 gnd.n7431 gnd.n259 585
R10684 gnd.n7434 gnd.n7433 585
R10685 gnd.n7433 gnd.n7432 585
R10686 gnd.n7435 gnd.n253 585
R10687 gnd.n253 gnd.n252 585
R10688 gnd.n7437 gnd.n7436 585
R10689 gnd.n7438 gnd.n7437 585
R10690 gnd.n251 gnd.n250 585
R10691 gnd.n7439 gnd.n251 585
R10692 gnd.n7442 gnd.n7441 585
R10693 gnd.n7441 gnd.n7440 585
R10694 gnd.n7443 gnd.n245 585
R10695 gnd.n245 gnd.n243 585
R10696 gnd.n7445 gnd.n7444 585
R10697 gnd.n7446 gnd.n7445 585
R10698 gnd.n246 gnd.n244 585
R10699 gnd.n244 gnd.n184 585
R10700 gnd.n3210 gnd.n3209 585
R10701 gnd.n3209 gnd.n171 585
R10702 gnd.n3211 gnd.n3203 585
R10703 gnd.n3203 gnd.n168 585
R10704 gnd.n3213 gnd.n3212 585
R10705 gnd.n3213 gnd.n176 585
R10706 gnd.n3214 gnd.n3202 585
R10707 gnd.n3214 gnd.n159 585
R10708 gnd.n3216 gnd.n3215 585
R10709 gnd.n3215 gnd.n152 585
R10710 gnd.n3217 gnd.n3197 585
R10711 gnd.n3197 gnd.n149 585
R10712 gnd.n3219 gnd.n3218 585
R10713 gnd.n3219 gnd.n141 585
R10714 gnd.n3220 gnd.n3196 585
R10715 gnd.n3220 gnd.n138 585
R10716 gnd.n3222 gnd.n3221 585
R10717 gnd.n3221 gnd.n131 585
R10718 gnd.n3223 gnd.n3191 585
R10719 gnd.n3191 gnd.n128 585
R10720 gnd.n3225 gnd.n3224 585
R10721 gnd.n3225 gnd.n120 585
R10722 gnd.n3226 gnd.n3190 585
R10723 gnd.n3226 gnd.n117 585
R10724 gnd.n5916 gnd.n5915 585
R10725 gnd.n5915 gnd.n5914 585
R10726 gnd.n5917 gnd.n3185 585
R10727 gnd.n3185 gnd.n108 585
R10728 gnd.n5919 gnd.n5918 585
R10729 gnd.n5919 gnd.n101 585
R10730 gnd.n5920 gnd.n3184 585
R10731 gnd.n5920 gnd.n98 585
R10732 gnd.n5922 gnd.n5921 585
R10733 gnd.n5921 gnd.n89 585
R10734 gnd.n5923 gnd.n3175 585
R10735 gnd.n3175 gnd.n86 585
R10736 gnd.n5926 gnd.n5925 585
R10737 gnd.n5927 gnd.n5926 585
R10738 gnd.n3182 gnd.n3174 585
R10739 gnd.n3174 gnd.n71 585
R10740 gnd.n3180 gnd.n3179 585
R10741 gnd.n3179 gnd.n69 585
R10742 gnd.n3178 gnd.n3177 585
R10743 gnd.n3178 gnd.n3166 585
R10744 gnd.n3154 gnd.n3153 585
R10745 gnd.n3159 gnd.n3154 585
R10746 gnd.n5943 gnd.n5942 585
R10747 gnd.n5942 gnd.n5941 585
R10748 gnd.n5945 gnd.n3151 585
R10749 gnd.n3155 gnd.n3151 585
R10750 gnd.n5947 gnd.n5946 585
R10751 gnd.n5948 gnd.n5947 585
R10752 gnd.n5793 gnd.n3150 585
R10753 gnd.n3150 gnd.n3143 585
R10754 gnd.n5795 gnd.n5794 585
R10755 gnd.n5795 gnd.n3140 585
R10756 gnd.n5796 gnd.n5790 585
R10757 gnd.n5796 gnd.n3241 585
R10758 gnd.n5798 gnd.n5797 585
R10759 gnd.n5797 gnd.n3131 585
R10760 gnd.n5799 gnd.n3249 585
R10761 gnd.n3249 gnd.n3123 585
R10762 gnd.n5801 gnd.n5800 585
R10763 gnd.n5802 gnd.n5801 585
R10764 gnd.n3250 gnd.n3248 585
R10765 gnd.n3248 gnd.n3114 585
R10766 gnd.n5784 gnd.n5783 585
R10767 gnd.n5783 gnd.n3111 585
R10768 gnd.n5782 gnd.n3252 585
R10769 gnd.n5782 gnd.n3103 585
R10770 gnd.n5781 gnd.n5780 585
R10771 gnd.n5781 gnd.n3100 585
R10772 gnd.n5761 gnd.n5760 585
R10773 gnd.n5760 gnd.n5759 585
R10774 gnd.n5776 gnd.n5775 585
R10775 gnd.n5775 gnd.n3091 585
R10776 gnd.n5774 gnd.n5763 585
R10777 gnd.n5774 gnd.n3083 585
R10778 gnd.n5773 gnd.n5772 585
R10779 gnd.n5773 gnd.n3080 585
R10780 gnd.n5765 gnd.n5764 585
R10781 gnd.n5764 gnd.n3071 585
R10782 gnd.n5768 gnd.n5767 585
R10783 gnd.n5767 gnd.n3068 585
R10784 gnd.n3055 gnd.n3054 585
R10785 gnd.n3059 gnd.n3055 585
R10786 gnd.n6004 gnd.n6003 585
R10787 gnd.n6003 gnd.n6002 585
R10788 gnd.n6005 gnd.n3049 585
R10789 gnd.n3056 gnd.n3049 585
R10790 gnd.n6007 gnd.n6006 585
R10791 gnd.n6008 gnd.n6007 585
R10792 gnd.n3046 gnd.n3045 585
R10793 gnd.n6009 gnd.n3046 585
R10794 gnd.n6012 gnd.n6011 585
R10795 gnd.n6011 gnd.n6010 585
R10796 gnd.n6013 gnd.n3040 585
R10797 gnd.n3040 gnd.n3038 585
R10798 gnd.n6015 gnd.n6014 585
R10799 gnd.n6016 gnd.n6015 585
R10800 gnd.n3041 gnd.n3039 585
R10801 gnd.n3039 gnd.n3036 585
R10802 gnd.n5378 gnd.n3356 585
R10803 gnd.n5378 gnd.n5377 585
R10804 gnd.n5380 gnd.n5379 585
R10805 gnd.n5379 gnd.n3303 585
R10806 gnd.n5381 gnd.n3349 585
R10807 gnd.n3349 gnd.n3340 585
R10808 gnd.n5383 gnd.n5382 585
R10809 gnd.n5384 gnd.n5383 585
R10810 gnd.n3350 gnd.n3348 585
R10811 gnd.n3433 gnd.n3348 585
R10812 gnd.n5166 gnd.n3378 585
R10813 gnd.n3432 gnd.n3378 585
R10814 gnd.n5168 gnd.n5167 585
R10815 gnd.n5169 gnd.n5168 585
R10816 gnd.n3379 gnd.n3377 585
R10817 gnd.n3377 gnd.n3374 585
R10818 gnd.n5160 gnd.n5159 585
R10819 gnd.n5159 gnd.n5158 585
R10820 gnd.n3382 gnd.n3381 585
R10821 gnd.n5147 gnd.n3382 585
R10822 gnd.n5137 gnd.n5136 585
R10823 gnd.n5138 gnd.n5137 585
R10824 gnd.n3401 gnd.n3400 585
R10825 gnd.n3450 gnd.n3400 585
R10826 gnd.n5132 gnd.n5131 585
R10827 gnd.n5131 gnd.n5130 585
R10828 gnd.n3404 gnd.n3403 585
R10829 gnd.n3411 gnd.n3404 585
R10830 gnd.n5094 gnd.n5093 585
R10831 gnd.n5095 gnd.n5094 585
R10832 gnd.n3459 gnd.n3458 585
R10833 gnd.n3458 gnd.n3420 585
R10834 gnd.n5089 gnd.n5088 585
R10835 gnd.n5088 gnd.n3425 585
R10836 gnd.n5087 gnd.n3461 585
R10837 gnd.n5087 gnd.n5086 585
R10838 gnd.n5066 gnd.n3462 585
R10839 gnd.n3468 gnd.n3462 585
R10840 gnd.n5068 gnd.n5067 585
R10841 gnd.n5069 gnd.n5068 585
R10842 gnd.n3476 gnd.n3475 585
R10843 gnd.n3483 gnd.n3475 585
R10844 gnd.n5061 gnd.n5060 585
R10845 gnd.n5060 gnd.n5059 585
R10846 gnd.n3479 gnd.n3478 585
R10847 gnd.n3487 gnd.n3479 585
R10848 gnd.n5014 gnd.n3503 585
R10849 gnd.n3503 gnd.n3497 585
R10850 gnd.n5016 gnd.n5015 585
R10851 gnd.n5017 gnd.n5016 585
R10852 gnd.n3504 gnd.n3502 585
R10853 gnd.n4991 gnd.n3502 585
R10854 gnd.n5009 gnd.n5008 585
R10855 gnd.n5008 gnd.n5007 585
R10856 gnd.n3507 gnd.n3506 585
R10857 gnd.n4999 gnd.n3507 585
R10858 gnd.n4945 gnd.n4944 585
R10859 gnd.n4944 gnd.n4943 585
R10860 gnd.n4946 gnd.n3534 585
R10861 gnd.n3534 gnd.n3525 585
R10862 gnd.n4948 gnd.n4947 585
R10863 gnd.n4949 gnd.n4948 585
R10864 gnd.n3535 gnd.n3533 585
R10865 gnd.n3533 gnd.n3530 585
R10866 gnd.n4934 gnd.n4933 585
R10867 gnd.n4933 gnd.n4932 585
R10868 gnd.n3538 gnd.n3537 585
R10869 gnd.n3544 gnd.n3538 585
R10870 gnd.n4911 gnd.n4910 585
R10871 gnd.n4912 gnd.n4911 585
R10872 gnd.n3554 gnd.n3553 585
R10873 gnd.n3561 gnd.n3553 585
R10874 gnd.n4906 gnd.n4905 585
R10875 gnd.n4905 gnd.n4904 585
R10876 gnd.n3557 gnd.n3556 585
R10877 gnd.n3565 gnd.n3557 585
R10878 gnd.n4861 gnd.n3582 585
R10879 gnd.n3582 gnd.n3575 585
R10880 gnd.n4863 gnd.n4862 585
R10881 gnd.n4864 gnd.n4863 585
R10882 gnd.n3583 gnd.n3581 585
R10883 gnd.n3581 gnd.n3579 585
R10884 gnd.n4856 gnd.n4855 585
R10885 gnd.n4855 gnd.n4854 585
R10886 gnd.n3586 gnd.n3585 585
R10887 gnd.n4846 gnd.n3586 585
R10888 gnd.n4817 gnd.n4816 585
R10889 gnd.n4818 gnd.n4817 585
R10890 gnd.n3600 gnd.n3599 585
R10891 gnd.n4802 gnd.n3599 585
R10892 gnd.n4812 gnd.n4811 585
R10893 gnd.n4811 gnd.n4810 585
R10894 gnd.n3603 gnd.n3602 585
R10895 gnd.n4794 gnd.n3603 585
R10896 gnd.n4784 gnd.n4783 585
R10897 gnd.n4785 gnd.n4784 585
R10898 gnd.n3621 gnd.n3620 585
R10899 gnd.n3620 gnd.n3616 585
R10900 gnd.n4779 gnd.n4778 585
R10901 gnd.n4778 gnd.n4777 585
R10902 gnd.n3624 gnd.n3623 585
R10903 gnd.n3630 gnd.n3624 585
R10904 gnd.n4756 gnd.n4755 585
R10905 gnd.n4757 gnd.n4756 585
R10906 gnd.n3641 gnd.n3640 585
R10907 gnd.n3648 gnd.n3640 585
R10908 gnd.n4751 gnd.n4750 585
R10909 gnd.n4750 gnd.n4749 585
R10910 gnd.n3644 gnd.n3643 585
R10911 gnd.n3652 gnd.n3644 585
R10912 gnd.n4683 gnd.n3668 585
R10913 gnd.n3668 gnd.n3661 585
R10914 gnd.n4685 gnd.n4684 585
R10915 gnd.n4686 gnd.n4685 585
R10916 gnd.n3669 gnd.n3667 585
R10917 gnd.n4660 gnd.n3667 585
R10918 gnd.n4678 gnd.n4677 585
R10919 gnd.n4677 gnd.n4676 585
R10920 gnd.n3672 gnd.n3671 585
R10921 gnd.n4668 gnd.n3672 585
R10922 gnd.n4638 gnd.n4637 585
R10923 gnd.n4639 gnd.n4638 585
R10924 gnd.n3684 gnd.n3683 585
R10925 gnd.n3693 gnd.n3683 585
R10926 gnd.n4633 gnd.n4632 585
R10927 gnd.n4632 gnd.n4631 585
R10928 gnd.n3687 gnd.n3686 585
R10929 gnd.n3702 gnd.n3687 585
R10930 gnd.n4595 gnd.n4594 585
R10931 gnd.n4596 gnd.n4595 585
R10932 gnd.n3709 gnd.n3708 585
R10933 gnd.n4585 gnd.n3708 585
R10934 gnd.n4590 gnd.n4589 585
R10935 gnd.n4589 gnd.n4588 585
R10936 gnd.n3712 gnd.n3711 585
R10937 gnd.n3718 gnd.n3712 585
R10938 gnd.n4559 gnd.n4558 585
R10939 gnd.n4560 gnd.n4559 585
R10940 gnd.n2939 gnd.n2938 585
R10941 gnd.n4525 gnd.n2939 585
R10942 gnd.n6131 gnd.n6130 585
R10943 gnd.n6130 gnd.n6129 585
R10944 gnd.n6132 gnd.n2933 585
R10945 gnd.n3733 gnd.n2933 585
R10946 gnd.n6134 gnd.n6133 585
R10947 gnd.n6135 gnd.n6134 585
R10948 gnd.n2921 gnd.n2920 585
R10949 gnd.n2924 gnd.n2921 585
R10950 gnd.n6145 gnd.n6144 585
R10951 gnd.n6144 gnd.n6143 585
R10952 gnd.n6146 gnd.n2915 585
R10953 gnd.n4499 gnd.n2915 585
R10954 gnd.n6148 gnd.n6147 585
R10955 gnd.n6149 gnd.n6148 585
R10956 gnd.n2916 gnd.n2914 585
R10957 gnd.n3825 gnd.n2914 585
R10958 gnd.n4472 gnd.n3839 585
R10959 gnd.n3839 gnd.n2886 585
R10960 gnd.n4474 gnd.n4473 585
R10961 gnd.n4475 gnd.n4474 585
R10962 gnd.n3840 gnd.n3838 585
R10963 gnd.n3838 gnd.n3832 585
R10964 gnd.n4466 gnd.n4465 585
R10965 gnd.n4465 gnd.n4464 585
R10966 gnd.n4462 gnd.n3842 585
R10967 gnd.n4462 gnd.n2601 585
R10968 gnd.n4461 gnd.n4460 585
R10969 gnd.n4461 gnd.n2587 585
R10970 gnd.n3845 gnd.n3844 585
R10971 gnd.n3844 gnd.n3843 585
R10972 gnd.n4456 gnd.n4455 585
R10973 gnd.n4455 gnd.n2690 585
R10974 gnd.n4454 gnd.n3847 585
R10975 gnd.n4454 gnd.n2676 585
R10976 gnd.n4453 gnd.n4452 585
R10977 gnd.n4453 gnd.n2574 585
R10978 gnd.n3849 gnd.n3848 585
R10979 gnd.n3848 gnd.n2571 585
R10980 gnd.n4448 gnd.n4447 585
R10981 gnd.n4447 gnd.n2564 585
R10982 gnd.n4446 gnd.n3851 585
R10983 gnd.n4446 gnd.n2561 585
R10984 gnd.n4445 gnd.n4444 585
R10985 gnd.n4445 gnd.n2554 585
R10986 gnd.n3853 gnd.n3852 585
R10987 gnd.n3852 gnd.n2551 585
R10988 gnd.n4440 gnd.n4439 585
R10989 gnd.n4439 gnd.n2543 585
R10990 gnd.n4438 gnd.n3855 585
R10991 gnd.n4438 gnd.n4437 585
R10992 gnd.n4377 gnd.n3856 585
R10993 gnd.n3856 gnd.n2534 585
R10994 gnd.n4379 gnd.n4378 585
R10995 gnd.n4378 gnd.n2531 585
R10996 gnd.n4380 gnd.n4371 585
R10997 gnd.n4371 gnd.n2523 585
R10998 gnd.n4382 gnd.n4381 585
R10999 gnd.n4382 gnd.n2520 585
R11000 gnd.n4383 gnd.n4370 585
R11001 gnd.n4383 gnd.n3868 585
R11002 gnd.n4385 gnd.n4384 585
R11003 gnd.n4384 gnd.n2511 585
R11004 gnd.n4386 gnd.n3876 585
R11005 gnd.n3876 gnd.n2503 585
R11006 gnd.n4388 gnd.n4387 585
R11007 gnd.n4389 gnd.n4388 585
R11008 gnd.n3877 gnd.n3875 585
R11009 gnd.n3875 gnd.n2494 585
R11010 gnd.n4323 gnd.n4322 585
R11011 gnd.n4323 gnd.n2491 585
R11012 gnd.n4325 gnd.n4324 585
R11013 gnd.n4324 gnd.n2486 585
R11014 gnd.n4327 gnd.n4326 585
R11015 gnd.n4327 gnd.n2483 585
R11016 gnd.n4330 gnd.n4329 585
R11017 gnd.n4331 gnd.n4330 585
R11018 gnd.n4328 gnd.n4321 585
R11019 gnd.n4321 gnd.n2474 585
R11020 gnd.n3888 gnd.n3887 585
R11021 gnd.n3887 gnd.n2469 585
R11022 gnd.n4356 gnd.n3889 585
R11023 gnd.n4356 gnd.n4355 585
R11024 gnd.n4358 gnd.n4357 585
R11025 gnd.n4357 gnd.n2460 585
R11026 gnd.n4360 gnd.n4359 585
R11027 gnd.n4360 gnd.n2457 585
R11028 gnd.n4361 gnd.n3885 585
R11029 gnd.n4361 gnd.n2451 585
R11030 gnd.n4363 gnd.n4362 585
R11031 gnd.n4362 gnd.n2448 585
R11032 gnd.n3886 gnd.n3884 585
R11033 gnd.n3886 gnd.n2441 585
R11034 gnd.n4282 gnd.n4281 585
R11035 gnd.n4281 gnd.n2438 585
R11036 gnd.n4283 gnd.n3910 585
R11037 gnd.n3910 gnd.n2430 585
R11038 gnd.n4285 gnd.n4284 585
R11039 gnd.n4286 gnd.n4285 585
R11040 gnd.n3911 gnd.n3909 585
R11041 gnd.n3909 gnd.n2421 585
R11042 gnd.n4275 gnd.n4274 585
R11043 gnd.n4274 gnd.n2418 585
R11044 gnd.n4273 gnd.n3913 585
R11045 gnd.n4273 gnd.n2410 585
R11046 gnd.n4272 gnd.n4271 585
R11047 gnd.n4272 gnd.n2407 585
R11048 gnd.n3915 gnd.n3914 585
R11049 gnd.n3914 gnd.n2400 585
R11050 gnd.n4267 gnd.n4266 585
R11051 gnd.n4266 gnd.n2397 585
R11052 gnd.n4265 gnd.n3917 585
R11053 gnd.n4265 gnd.n2389 585
R11054 gnd.n4264 gnd.n4263 585
R11055 gnd.n4264 gnd.n2386 585
R11056 gnd.n3919 gnd.n3918 585
R11057 gnd.n3918 gnd.n2377 585
R11058 gnd.n4259 gnd.n4258 585
R11059 gnd.n4258 gnd.n4257 585
R11060 gnd.n3923 gnd.n3922 585
R11061 gnd.n3923 gnd.n2366 585
R11062 gnd.n2362 gnd.n2361 585
R11063 gnd.n6487 gnd.n2362 585
R11064 gnd.n6490 gnd.n6489 585
R11065 gnd.n6489 gnd.n6488 585
R11066 gnd.n6491 gnd.n2356 585
R11067 gnd.n2356 gnd.n2355 585
R11068 gnd.n6493 gnd.n6492 585
R11069 gnd.n6494 gnd.n6493 585
R11070 gnd.n2354 gnd.n2353 585
R11071 gnd.n6495 gnd.n2354 585
R11072 gnd.n6498 gnd.n6497 585
R11073 gnd.n6497 gnd.n6496 585
R11074 gnd.n6499 gnd.n2348 585
R11075 gnd.n2348 gnd.n2347 585
R11076 gnd.n6501 gnd.n6500 585
R11077 gnd.n6502 gnd.n6501 585
R11078 gnd.n2346 gnd.n2345 585
R11079 gnd.n6503 gnd.n2346 585
R11080 gnd.n6506 gnd.n6505 585
R11081 gnd.n6505 gnd.n6504 585
R11082 gnd.n6507 gnd.n2341 585
R11083 gnd.n2341 gnd.n2340 585
R11084 gnd.n6509 gnd.n6508 585
R11085 gnd.n6510 gnd.n6509 585
R11086 gnd.n876 gnd.n875 585
R11087 gnd.n6511 gnd.n876 585
R11088 gnd.n6514 gnd.n6513 585
R11089 gnd.n6513 gnd.n6512 585
R11090 gnd.n6019 gnd.n6018 585
R11091 gnd.n6018 gnd.n6017 585
R11092 gnd.n6020 gnd.n3034 585
R11093 gnd.n5376 gnd.n3034 585
R11094 gnd.n3357 gnd.n3032 585
R11095 gnd.n3358 gnd.n3357 585
R11096 gnd.n6024 gnd.n3031 585
R11097 gnd.n5189 gnd.n3031 585
R11098 gnd.n6025 gnd.n3030 585
R11099 gnd.n5187 gnd.n3030 585
R11100 gnd.n6026 gnd.n3029 585
R11101 gnd.n3345 gnd.n3029 585
R11102 gnd.n3435 gnd.n3027 585
R11103 gnd.n3436 gnd.n3435 585
R11104 gnd.n6030 gnd.n3026 585
R11105 gnd.n5179 gnd.n3026 585
R11106 gnd.n6031 gnd.n3025 585
R11107 gnd.n5171 gnd.n3025 585
R11108 gnd.n6032 gnd.n3024 585
R11109 gnd.n5156 gnd.n3024 585
R11110 gnd.n3392 gnd.n3022 585
R11111 gnd.n3393 gnd.n3392 585
R11112 gnd.n6036 gnd.n3021 585
R11113 gnd.n5148 gnd.n3021 585
R11114 gnd.n6037 gnd.n3020 585
R11115 gnd.n3398 gnd.n3020 585
R11116 gnd.n6038 gnd.n3019 585
R11117 gnd.n3407 gnd.n3019 585
R11118 gnd.n5121 gnd.n3017 585
R11119 gnd.n5122 gnd.n5121 585
R11120 gnd.n6042 gnd.n3016 585
R11121 gnd.n5096 gnd.n3016 585
R11122 gnd.n6043 gnd.n3015 585
R11123 gnd.n5112 gnd.n3015 585
R11124 gnd.n6044 gnd.n3014 585
R11125 gnd.n5104 gnd.n3014 585
R11126 gnd.n5084 gnd.n3012 585
R11127 gnd.n5085 gnd.n5084 585
R11128 gnd.n6048 gnd.n3011 585
R11129 gnd.t9 gnd.n3011 585
R11130 gnd.n6049 gnd.n3010 585
R11131 gnd.n5035 gnd.n3010 585
R11132 gnd.n6050 gnd.n3009 585
R11133 gnd.n3473 gnd.n3009 585
R11134 gnd.n5057 gnd.n3007 585
R11135 gnd.n5058 gnd.n5057 585
R11136 gnd.n6054 gnd.n3006 585
R11137 gnd.n5049 gnd.n3006 585
R11138 gnd.n6055 gnd.n3005 585
R11139 gnd.n4984 gnd.n3005 585
R11140 gnd.n6056 gnd.n3004 585
R11141 gnd.n5027 gnd.n3004 585
R11142 gnd.n5018 gnd.n3002 585
R11143 gnd.n5019 gnd.n5018 585
R11144 gnd.n6060 gnd.n3001 585
R11145 gnd.n3510 gnd.n3001 585
R11146 gnd.n6061 gnd.n3000 585
R11147 gnd.n3508 gnd.n3000 585
R11148 gnd.n6062 gnd.n2999 585
R11149 gnd.n4971 gnd.n2999 585
R11150 gnd.n4941 gnd.n2997 585
R11151 gnd.n4942 gnd.n4941 585
R11152 gnd.n6066 gnd.n2996 585
R11153 gnd.n4959 gnd.n2996 585
R11154 gnd.n6067 gnd.n2995 585
R11155 gnd.n4950 gnd.n2995 585
R11156 gnd.n6068 gnd.n2994 585
R11157 gnd.n4931 gnd.n2994 585
R11158 gnd.n4880 gnd.n2992 585
R11159 gnd.n4881 gnd.n4880 585
R11160 gnd.n6072 gnd.n2991 585
R11161 gnd.n3552 gnd.n2991 585
R11162 gnd.n6073 gnd.n2990 585
R11163 gnd.n3549 gnd.n2990 585
R11164 gnd.n6074 gnd.n2989 585
R11165 gnd.n4903 gnd.n2989 585
R11166 gnd.n4894 gnd.n2987 585
R11167 gnd.n4895 gnd.n4894 585
R11168 gnd.n6078 gnd.n2986 585
R11169 gnd.n4831 gnd.n2986 585
R11170 gnd.n6079 gnd.n2985 585
R11171 gnd.n4872 gnd.n2985 585
R11172 gnd.n6080 gnd.n2984 585
R11173 gnd.n4865 gnd.n2984 585
R11174 gnd.n3589 gnd.n2982 585
R11175 gnd.n3590 gnd.n3589 585
R11176 gnd.n6084 gnd.n2981 585
R11177 gnd.n3587 gnd.n2981 585
R11178 gnd.n6085 gnd.n2980 585
R11179 gnd.n3594 gnd.n2980 585
R11180 gnd.n6086 gnd.n2979 585
R11181 gnd.n3598 gnd.n2979 585
R11182 gnd.n3606 gnd.n2977 585
R11183 gnd.n3607 gnd.n3606 585
R11184 gnd.n6090 gnd.n2976 585
R11185 gnd.n3604 gnd.n2976 585
R11186 gnd.n6091 gnd.n2975 585
R11187 gnd.n4706 gnd.n2975 585
R11188 gnd.n6092 gnd.n2974 585
R11189 gnd.n4786 gnd.n2974 585
R11190 gnd.n4775 gnd.n2972 585
R11191 gnd.n4776 gnd.n4775 585
R11192 gnd.n6096 gnd.n2971 585
R11193 gnd.n3631 gnd.n2971 585
R11194 gnd.n6097 gnd.n2970 585
R11195 gnd.n3639 gnd.n2970 585
R11196 gnd.n6098 gnd.n2969 585
R11197 gnd.n3636 gnd.n2969 585
R11198 gnd.n4747 gnd.n2967 585
R11199 gnd.n4748 gnd.n4747 585
R11200 gnd.n6102 gnd.n2966 585
R11201 gnd.n4739 gnd.n2966 585
R11202 gnd.n6103 gnd.n2965 585
R11203 gnd.n4652 gnd.n2965 585
R11204 gnd.n6104 gnd.n2964 585
R11205 gnd.n4695 gnd.n2964 585
R11206 gnd.n4687 gnd.n2962 585
R11207 gnd.n4688 gnd.n4687 585
R11208 gnd.n6108 gnd.n2961 585
R11209 gnd.n3675 gnd.n2961 585
R11210 gnd.n6109 gnd.n2960 585
R11211 gnd.n3673 gnd.n2960 585
R11212 gnd.n6110 gnd.n2959 585
R11213 gnd.n3679 gnd.n2959 585
R11214 gnd.n4622 gnd.n2957 585
R11215 gnd.n4623 gnd.n4622 585
R11216 gnd.n6114 gnd.n2956 585
R11217 gnd.t189 gnd.n2956 585
R11218 gnd.n6115 gnd.n2955 585
R11219 gnd.n3688 gnd.n2955 585
R11220 gnd.n6116 gnd.n2954 585
R11221 gnd.n4606 gnd.n2954 585
R11222 gnd.n4597 gnd.n2952 585
R11223 gnd.n4598 gnd.n4597 585
R11224 gnd.n6120 gnd.n2951 585
R11225 gnd.n4587 gnd.n2951 585
R11226 gnd.n6121 gnd.n2950 585
R11227 gnd.n3719 gnd.n2950 585
R11228 gnd.n6122 gnd.n2949 585
R11229 gnd.n4555 gnd.n2949 585
R11230 gnd.n2946 gnd.n2944 585
R11231 gnd.n3724 gnd.n2944 585
R11232 gnd.n6127 gnd.n6126 585
R11233 gnd.n6128 gnd.n6127 585
R11234 gnd.n2945 gnd.n2943 585
R11235 gnd.n4540 gnd.n2943 585
R11236 gnd.n3741 gnd.n3739 585
R11237 gnd.n3739 gnd.n2932 585
R11238 gnd.n4516 gnd.n4515 585
R11239 gnd.n4517 gnd.n4516 585
R11240 gnd.n3740 gnd.n2925 585
R11241 gnd.n6142 gnd.n2925 585
R11242 gnd.n4510 gnd.n4509 585
R11243 gnd.n4509 gnd.n4508 585
R11244 gnd.n3744 gnd.n3743 585
R11245 gnd.n4500 gnd.n3744 585
R11246 gnd.n3829 gnd.n3827 585
R11247 gnd.n3827 gnd.n2912 585
R11248 gnd.n4484 gnd.n4483 585
R11249 gnd.n4485 gnd.n4484 585
R11250 gnd.n3828 gnd.n3826 585
R11251 gnd.n3826 gnd.n2854 585
R11252 gnd.n4478 gnd.n4477 585
R11253 gnd.n4477 gnd.n4476 585
R11254 gnd.n3831 gnd.n2604 585
R11255 gnd.n4463 gnd.n2604 585
R11256 gnd.n6337 gnd.n6336 585
R11257 gnd.n6335 gnd.n2603 585
R11258 gnd.n2606 gnd.n2602 585
R11259 gnd.n6339 gnd.n2602 585
R11260 gnd.n6331 gnd.n2608 585
R11261 gnd.n6330 gnd.n2609 585
R11262 gnd.n6329 gnd.n2610 585
R11263 gnd.n2613 gnd.n2611 585
R11264 gnd.n6324 gnd.n2614 585
R11265 gnd.n6323 gnd.n2615 585
R11266 gnd.n6322 gnd.n2616 585
R11267 gnd.n2625 gnd.n2617 585
R11268 gnd.n6315 gnd.n2626 585
R11269 gnd.n6314 gnd.n2627 585
R11270 gnd.n2629 gnd.n2628 585
R11271 gnd.n6307 gnd.n2635 585
R11272 gnd.n6306 gnd.n2636 585
R11273 gnd.n2643 gnd.n2637 585
R11274 gnd.n6299 gnd.n2644 585
R11275 gnd.n6298 gnd.n2645 585
R11276 gnd.n2647 gnd.n2646 585
R11277 gnd.n6291 gnd.n2653 585
R11278 gnd.n6290 gnd.n2654 585
R11279 gnd.n2661 gnd.n2655 585
R11280 gnd.n6283 gnd.n2662 585
R11281 gnd.n6282 gnd.n2663 585
R11282 gnd.n2668 gnd.n2667 585
R11283 gnd.n2599 gnd.n2584 585
R11284 gnd.n6343 gnd.n2585 585
R11285 gnd.n6342 gnd.n6341 585
R11286 gnd.n3361 gnd.n3037 585
R11287 gnd.n6017 gnd.n3037 585
R11288 gnd.n5375 gnd.n5374 585
R11289 gnd.n5376 gnd.n5375 585
R11290 gnd.n3360 gnd.n3359 585
R11291 gnd.n3359 gnd.n3358 585
R11292 gnd.n5191 gnd.n5190 585
R11293 gnd.n5190 gnd.n5189 585
R11294 gnd.n5188 gnd.n3363 585
R11295 gnd.n5188 gnd.n5187 585
R11296 gnd.n5186 gnd.n5185 585
R11297 gnd.n5186 gnd.n3345 585
R11298 gnd.n3365 gnd.n3364 585
R11299 gnd.n3436 gnd.n3364 585
R11300 gnd.n5181 gnd.n5180 585
R11301 gnd.n5180 gnd.n5179 585
R11302 gnd.n3368 gnd.n3367 585
R11303 gnd.n5171 gnd.n3368 585
R11304 gnd.n5155 gnd.n5154 585
R11305 gnd.n5156 gnd.n5155 585
R11306 gnd.n3386 gnd.n3385 585
R11307 gnd.n3393 gnd.n3385 585
R11308 gnd.n5150 gnd.n5149 585
R11309 gnd.n5149 gnd.n5148 585
R11310 gnd.n3389 gnd.n3388 585
R11311 gnd.n3398 gnd.n3389 585
R11312 gnd.n3416 gnd.n3414 585
R11313 gnd.n3414 gnd.n3407 585
R11314 gnd.n5120 gnd.n5119 585
R11315 gnd.n5122 gnd.n5120 585
R11316 gnd.n3415 gnd.n3413 585
R11317 gnd.n5096 gnd.n3413 585
R11318 gnd.n5114 gnd.n5113 585
R11319 gnd.n5113 gnd.n5112 585
R11320 gnd.n3419 gnd.n3418 585
R11321 gnd.n5104 gnd.n3419 585
R11322 gnd.n5038 gnd.n3464 585
R11323 gnd.n5085 gnd.n3464 585
R11324 gnd.n5041 gnd.n5037 585
R11325 gnd.n5037 gnd.t9 585
R11326 gnd.n5042 gnd.n5036 585
R11327 gnd.n5036 gnd.n5035 585
R11328 gnd.n5043 gnd.n5033 585
R11329 gnd.n5033 gnd.n3473 585
R11330 gnd.n3491 gnd.n3481 585
R11331 gnd.n5058 gnd.n3481 585
R11332 gnd.n5048 gnd.n5047 585
R11333 gnd.n5049 gnd.n5048 585
R11334 gnd.n3490 gnd.n3489 585
R11335 gnd.n4984 gnd.n3489 585
R11336 gnd.n5029 gnd.n5028 585
R11337 gnd.n5028 gnd.n5027 585
R11338 gnd.n3494 gnd.n3493 585
R11339 gnd.n5019 gnd.n3494 585
R11340 gnd.n4965 gnd.n4964 585
R11341 gnd.n4964 gnd.n3510 585
R11342 gnd.n3520 gnd.n3518 585
R11343 gnd.n3518 gnd.n3508 585
R11344 gnd.n4970 gnd.n4969 585
R11345 gnd.n4971 gnd.n4970 585
R11346 gnd.n3519 gnd.n3517 585
R11347 gnd.n4942 gnd.n3517 585
R11348 gnd.n4961 gnd.n4960 585
R11349 gnd.n4960 gnd.n4959 585
R11350 gnd.n3523 gnd.n3522 585
R11351 gnd.n4950 gnd.n3523 585
R11352 gnd.n4883 gnd.n3540 585
R11353 gnd.n4931 gnd.n3540 585
R11354 gnd.n4886 gnd.n4882 585
R11355 gnd.n4882 gnd.n4881 585
R11356 gnd.n4887 gnd.n4879 585
R11357 gnd.n4879 gnd.n3552 585
R11358 gnd.n4888 gnd.n4878 585
R11359 gnd.n4878 gnd.n3549 585
R11360 gnd.n3569 gnd.n3559 585
R11361 gnd.n4903 gnd.n3559 585
R11362 gnd.n4893 gnd.n4892 585
R11363 gnd.n4895 gnd.n4893 585
R11364 gnd.n3568 gnd.n3567 585
R11365 gnd.n4831 gnd.n3567 585
R11366 gnd.n4874 gnd.n4873 585
R11367 gnd.n4873 gnd.n4872 585
R11368 gnd.n3572 gnd.n3571 585
R11369 gnd.n4865 gnd.n3572 585
R11370 gnd.n4716 gnd.n4715 585
R11371 gnd.n4715 gnd.n3590 585
R11372 gnd.n4719 gnd.n4714 585
R11373 gnd.n4714 gnd.n3587 585
R11374 gnd.n4720 gnd.n4713 585
R11375 gnd.n4713 gnd.n3594 585
R11376 gnd.n4721 gnd.n4712 585
R11377 gnd.n4712 gnd.n3598 585
R11378 gnd.n4711 gnd.n4709 585
R11379 gnd.n4711 gnd.n3607 585
R11380 gnd.n4725 gnd.n4708 585
R11381 gnd.n4708 gnd.n3604 585
R11382 gnd.n4726 gnd.n4707 585
R11383 gnd.n4707 gnd.n4706 585
R11384 gnd.n4727 gnd.n3618 585
R11385 gnd.n4786 gnd.n3618 585
R11386 gnd.n4704 gnd.n3626 585
R11387 gnd.n4776 gnd.n3626 585
R11388 gnd.n4731 gnd.n4703 585
R11389 gnd.n4703 gnd.n3631 585
R11390 gnd.n4732 gnd.n4702 585
R11391 gnd.n4702 gnd.n3639 585
R11392 gnd.n4733 gnd.n4701 585
R11393 gnd.n4701 gnd.n3636 585
R11394 gnd.n3656 gnd.n3646 585
R11395 gnd.n4748 gnd.n3646 585
R11396 gnd.n4738 gnd.n4737 585
R11397 gnd.n4739 gnd.n4738 585
R11398 gnd.n3655 gnd.n3654 585
R11399 gnd.n4652 gnd.n3654 585
R11400 gnd.n4697 gnd.n4696 585
R11401 gnd.n4696 gnd.n4695 585
R11402 gnd.n3659 gnd.n3658 585
R11403 gnd.n4688 gnd.n3659 585
R11404 gnd.n4615 gnd.n4614 585
R11405 gnd.n4614 gnd.n3675 585
R11406 gnd.n4616 gnd.n4613 585
R11407 gnd.n4613 gnd.n3673 585
R11408 gnd.n3697 gnd.n3695 585
R11409 gnd.n3695 gnd.n3679 585
R11410 gnd.n4621 gnd.n4620 585
R11411 gnd.n4623 gnd.n4621 585
R11412 gnd.n3696 gnd.n3694 585
R11413 gnd.n3694 gnd.t189 585
R11414 gnd.n4609 gnd.n4608 585
R11415 gnd.n4608 gnd.n3688 585
R11416 gnd.n4607 gnd.n3699 585
R11417 gnd.n4607 gnd.n4606 585
R11418 gnd.n4547 gnd.n3700 585
R11419 gnd.n4598 gnd.n3700 585
R11420 gnd.n4548 gnd.n3714 585
R11421 gnd.n4587 gnd.n3714 585
R11422 gnd.n3729 gnd.n3727 585
R11423 gnd.n3727 gnd.n3719 585
R11424 gnd.n4553 gnd.n4552 585
R11425 gnd.n4555 gnd.n4553 585
R11426 gnd.n3728 gnd.n3726 585
R11427 gnd.n3726 gnd.n3724 585
R11428 gnd.n4543 gnd.n2941 585
R11429 gnd.n6128 gnd.n2941 585
R11430 gnd.n4542 gnd.n4541 585
R11431 gnd.n4541 gnd.n4540 585
R11432 gnd.n3732 gnd.n3731 585
R11433 gnd.n3732 gnd.n2932 585
R11434 gnd.n4492 gnd.n3738 585
R11435 gnd.n4517 gnd.n3738 585
R11436 gnd.n4493 gnd.n2923 585
R11437 gnd.n6142 gnd.n2923 585
R11438 gnd.n3753 gnd.n3748 585
R11439 gnd.n4508 gnd.n3748 585
R11440 gnd.n4498 gnd.n4497 585
R11441 gnd.n4500 gnd.n4498 585
R11442 gnd.n3752 gnd.n3751 585
R11443 gnd.n3751 gnd.n2912 585
R11444 gnd.n4487 gnd.n4486 585
R11445 gnd.n4486 gnd.n4485 585
R11446 gnd.n3756 gnd.n3755 585
R11447 gnd.n3756 gnd.n2854 585
R11448 gnd.n3837 gnd.n3836 585
R11449 gnd.n4476 gnd.n3837 585
R11450 gnd.n3833 gnd.n2586 585
R11451 gnd.n4463 gnd.n2586 585
R11452 gnd.n5349 gnd.n5203 585
R11453 gnd.n5203 gnd.n3047 585
R11454 gnd.n5350 gnd.n5347 585
R11455 gnd.n5345 gnd.n5221 585
R11456 gnd.n5344 gnd.n5343 585
R11457 gnd.n5328 gnd.n5223 585
R11458 gnd.n5330 gnd.n5329 585
R11459 gnd.n5326 gnd.n5230 585
R11460 gnd.n5325 gnd.n5324 585
R11461 gnd.n5309 gnd.n5232 585
R11462 gnd.n5311 gnd.n5310 585
R11463 gnd.n5307 gnd.n5239 585
R11464 gnd.n5306 gnd.n5305 585
R11465 gnd.n5290 gnd.n5241 585
R11466 gnd.n5292 gnd.n5291 585
R11467 gnd.n5288 gnd.n5248 585
R11468 gnd.n5287 gnd.n5286 585
R11469 gnd.n5275 gnd.n5250 585
R11470 gnd.n5277 gnd.n5276 585
R11471 gnd.n5273 gnd.n5251 585
R11472 gnd.n5272 gnd.n5271 585
R11473 gnd.n5264 gnd.n5253 585
R11474 gnd.n5266 gnd.n5265 585
R11475 gnd.n5262 gnd.n5255 585
R11476 gnd.n5261 gnd.n5260 585
R11477 gnd.n5257 gnd.n3035 585
R11478 gnd.n5370 gnd.n5369 585
R11479 gnd.n5367 gnd.n5201 585
R11480 gnd.n5366 gnd.n5202 585
R11481 gnd.n5364 gnd.n5363 585
R11482 gnd.n6690 gnd.n705 540.215
R11483 gnd.n5474 gnd.n3342 506.916
R11484 gnd.n5477 gnd.n5476 506.916
R11485 gnd.n3823 gnd.n3757 506.916
R11486 gnd.n6218 gnd.n2889 506.916
R11487 gnd.n3758 gnd.t148 389.64
R11488 gnd.n3336 gnd.t75 389.64
R11489 gnd.n6155 gnd.t82 389.64
R11490 gnd.n5408 gnd.t129 389.64
R11491 gnd.n2664 gnd.t112 371.625
R11492 gnd.n5214 gnd.t135 371.625
R11493 gnd.n2671 gnd.t151 371.625
R11494 gnd.n5614 gnd.t132 371.625
R11495 gnd.n5666 gnd.t120 371.625
R11496 gnd.n3267 gnd.t62 371.625
R11497 gnd.n7538 gnd.t69 371.625
R11498 gnd.n7517 gnd.t58 371.625
R11499 gnd.n7624 gnd.t126 371.625
R11500 gnd.n180 gnd.t145 371.625
R11501 gnd.n4045 gnd.t97 371.625
R11502 gnd.n4156 gnd.t79 371.625
R11503 gnd.n4001 gnd.t103 371.625
R11504 gnd.n3961 gnd.t54 371.625
R11505 gnd.n2741 gnd.t138 371.625
R11506 gnd.n2782 gnd.t86 371.625
R11507 gnd.n2761 gnd.t106 371.625
R11508 gnd.n5204 gnd.t93 371.625
R11509 gnd.n7422 gnd.n268 368.44
R11510 gnd.n1356 gnd.t116 323.425
R11511 gnd.n916 gnd.t141 323.425
R11512 gnd.n7212 gnd.n7211 301.784
R11513 gnd.n7213 gnd.n7212 301.784
R11514 gnd.n7213 gnd.n388 301.784
R11515 gnd.n7221 gnd.n388 301.784
R11516 gnd.n7222 gnd.n7221 301.784
R11517 gnd.n7223 gnd.n7222 301.784
R11518 gnd.n7223 gnd.n382 301.784
R11519 gnd.n7231 gnd.n382 301.784
R11520 gnd.n7232 gnd.n7231 301.784
R11521 gnd.n7233 gnd.n7232 301.784
R11522 gnd.n7233 gnd.n376 301.784
R11523 gnd.n7241 gnd.n376 301.784
R11524 gnd.n7242 gnd.n7241 301.784
R11525 gnd.n7243 gnd.n7242 301.784
R11526 gnd.n7243 gnd.n370 301.784
R11527 gnd.n7251 gnd.n370 301.784
R11528 gnd.n7252 gnd.n7251 301.784
R11529 gnd.n7253 gnd.n7252 301.784
R11530 gnd.n7253 gnd.n364 301.784
R11531 gnd.n7261 gnd.n364 301.784
R11532 gnd.n7262 gnd.n7261 301.784
R11533 gnd.n7263 gnd.n7262 301.784
R11534 gnd.n7263 gnd.n358 301.784
R11535 gnd.n7271 gnd.n358 301.784
R11536 gnd.n7272 gnd.n7271 301.784
R11537 gnd.n7273 gnd.n7272 301.784
R11538 gnd.n7273 gnd.n352 301.784
R11539 gnd.n7281 gnd.n352 301.784
R11540 gnd.n7282 gnd.n7281 301.784
R11541 gnd.n7283 gnd.n7282 301.784
R11542 gnd.n7283 gnd.n346 301.784
R11543 gnd.n7291 gnd.n346 301.784
R11544 gnd.n7292 gnd.n7291 301.784
R11545 gnd.n7293 gnd.n7292 301.784
R11546 gnd.n7293 gnd.n340 301.784
R11547 gnd.n7301 gnd.n340 301.784
R11548 gnd.n7302 gnd.n7301 301.784
R11549 gnd.n7303 gnd.n7302 301.784
R11550 gnd.n7303 gnd.n334 301.784
R11551 gnd.n7311 gnd.n334 301.784
R11552 gnd.n7312 gnd.n7311 301.784
R11553 gnd.n7313 gnd.n7312 301.784
R11554 gnd.n7313 gnd.n328 301.784
R11555 gnd.n7321 gnd.n328 301.784
R11556 gnd.n7322 gnd.n7321 301.784
R11557 gnd.n7323 gnd.n7322 301.784
R11558 gnd.n7323 gnd.n322 301.784
R11559 gnd.n7331 gnd.n322 301.784
R11560 gnd.n7332 gnd.n7331 301.784
R11561 gnd.n7333 gnd.n7332 301.784
R11562 gnd.n7333 gnd.n316 301.784
R11563 gnd.n7341 gnd.n316 301.784
R11564 gnd.n7342 gnd.n7341 301.784
R11565 gnd.n7343 gnd.n7342 301.784
R11566 gnd.n7343 gnd.n310 301.784
R11567 gnd.n7351 gnd.n310 301.784
R11568 gnd.n7352 gnd.n7351 301.784
R11569 gnd.n7353 gnd.n7352 301.784
R11570 gnd.n7353 gnd.n304 301.784
R11571 gnd.n7361 gnd.n304 301.784
R11572 gnd.n7362 gnd.n7361 301.784
R11573 gnd.n7363 gnd.n7362 301.784
R11574 gnd.n7363 gnd.n298 301.784
R11575 gnd.n7371 gnd.n298 301.784
R11576 gnd.n7372 gnd.n7371 301.784
R11577 gnd.n7373 gnd.n7372 301.784
R11578 gnd.n7373 gnd.n292 301.784
R11579 gnd.n7381 gnd.n292 301.784
R11580 gnd.n7382 gnd.n7381 301.784
R11581 gnd.n7383 gnd.n7382 301.784
R11582 gnd.n7383 gnd.n286 301.784
R11583 gnd.n7391 gnd.n286 301.784
R11584 gnd.n7392 gnd.n7391 301.784
R11585 gnd.n7393 gnd.n7392 301.784
R11586 gnd.n7393 gnd.n280 301.784
R11587 gnd.n7401 gnd.n280 301.784
R11588 gnd.n7402 gnd.n7401 301.784
R11589 gnd.n7403 gnd.n7402 301.784
R11590 gnd.n7403 gnd.n274 301.784
R11591 gnd.n7411 gnd.n274 301.784
R11592 gnd.n7412 gnd.n7411 301.784
R11593 gnd.n7413 gnd.n7412 301.784
R11594 gnd.n7413 gnd.n268 301.784
R11595 gnd.n2206 gnd.n2180 289.615
R11596 gnd.n2174 gnd.n2148 289.615
R11597 gnd.n2142 gnd.n2116 289.615
R11598 gnd.n2111 gnd.n2085 289.615
R11599 gnd.n2079 gnd.n2053 289.615
R11600 gnd.n2047 gnd.n2021 289.615
R11601 gnd.n2015 gnd.n1989 289.615
R11602 gnd.n1984 gnd.n1958 289.615
R11603 gnd.n1430 gnd.t47 279.217
R11604 gnd.n942 gnd.t37 279.217
R11605 gnd.n2896 gnd.t111 260.649
R11606 gnd.n5400 gnd.t125 260.649
R11607 gnd.n6220 gnd.n6219 256.663
R11608 gnd.n6220 gnd.n2855 256.663
R11609 gnd.n6220 gnd.n2856 256.663
R11610 gnd.n6220 gnd.n2857 256.663
R11611 gnd.n6220 gnd.n2858 256.663
R11612 gnd.n6220 gnd.n2859 256.663
R11613 gnd.n6220 gnd.n2860 256.663
R11614 gnd.n6220 gnd.n2861 256.663
R11615 gnd.n6220 gnd.n2862 256.663
R11616 gnd.n6220 gnd.n2863 256.663
R11617 gnd.n6220 gnd.n2864 256.663
R11618 gnd.n6220 gnd.n2865 256.663
R11619 gnd.n6220 gnd.n2866 256.663
R11620 gnd.n6220 gnd.n2867 256.663
R11621 gnd.n6220 gnd.n2868 256.663
R11622 gnd.n6220 gnd.n2869 256.663
R11623 gnd.n6223 gnd.n2852 256.663
R11624 gnd.n6221 gnd.n6220 256.663
R11625 gnd.n6220 gnd.n2870 256.663
R11626 gnd.n6220 gnd.n2871 256.663
R11627 gnd.n6220 gnd.n2872 256.663
R11628 gnd.n6220 gnd.n2873 256.663
R11629 gnd.n6220 gnd.n2874 256.663
R11630 gnd.n6220 gnd.n2875 256.663
R11631 gnd.n6220 gnd.n2876 256.663
R11632 gnd.n6220 gnd.n2877 256.663
R11633 gnd.n6220 gnd.n2878 256.663
R11634 gnd.n6220 gnd.n2879 256.663
R11635 gnd.n6220 gnd.n2880 256.663
R11636 gnd.n6220 gnd.n2881 256.663
R11637 gnd.n6220 gnd.n2882 256.663
R11638 gnd.n6220 gnd.n2883 256.663
R11639 gnd.n6220 gnd.n2884 256.663
R11640 gnd.n6220 gnd.n2885 256.663
R11641 gnd.n5542 gnd.n3320 256.663
R11642 gnd.n5542 gnd.n3321 256.663
R11643 gnd.n5542 gnd.n3322 256.663
R11644 gnd.n5542 gnd.n3323 256.663
R11645 gnd.n5542 gnd.n3324 256.663
R11646 gnd.n5542 gnd.n3325 256.663
R11647 gnd.n5542 gnd.n3326 256.663
R11648 gnd.n5542 gnd.n3327 256.663
R11649 gnd.n5542 gnd.n3328 256.663
R11650 gnd.n5542 gnd.n3329 256.663
R11651 gnd.n5542 gnd.n3330 256.663
R11652 gnd.n5542 gnd.n3331 256.663
R11653 gnd.n5542 gnd.n3332 256.663
R11654 gnd.n5542 gnd.n3333 256.663
R11655 gnd.n5542 gnd.n3334 256.663
R11656 gnd.n5542 gnd.n5539 256.663
R11657 gnd.n5545 gnd.n3301 256.663
R11658 gnd.n5543 gnd.n5542 256.663
R11659 gnd.n5542 gnd.n3319 256.663
R11660 gnd.n5542 gnd.n3318 256.663
R11661 gnd.n5542 gnd.n3317 256.663
R11662 gnd.n5542 gnd.n3316 256.663
R11663 gnd.n5542 gnd.n3315 256.663
R11664 gnd.n5542 gnd.n3314 256.663
R11665 gnd.n5542 gnd.n3313 256.663
R11666 gnd.n5542 gnd.n3312 256.663
R11667 gnd.n5542 gnd.n3311 256.663
R11668 gnd.n5542 gnd.n3310 256.663
R11669 gnd.n5542 gnd.n3309 256.663
R11670 gnd.n5542 gnd.n3308 256.663
R11671 gnd.n5542 gnd.n3307 256.663
R11672 gnd.n5542 gnd.n3306 256.663
R11673 gnd.n5542 gnd.n3305 256.663
R11674 gnd.n5542 gnd.n3304 256.663
R11675 gnd.n3996 gnd.n2363 242.672
R11676 gnd.n3933 gnd.n2363 242.672
R11677 gnd.n3989 gnd.n2363 242.672
R11678 gnd.n3983 gnd.n2363 242.672
R11679 gnd.n3981 gnd.n2363 242.672
R11680 gnd.n3975 gnd.n2363 242.672
R11681 gnd.n3973 gnd.n2363 242.672
R11682 gnd.n3967 gnd.n2363 242.672
R11683 gnd.n3965 gnd.n2363 242.672
R11684 gnd.n6275 gnd.n6274 242.672
R11685 gnd.n6274 gnd.n2689 242.672
R11686 gnd.n6274 gnd.n2687 242.672
R11687 gnd.n6274 gnd.n2686 242.672
R11688 gnd.n6274 gnd.n2684 242.672
R11689 gnd.n6274 gnd.n2682 242.672
R11690 gnd.n6274 gnd.n2681 242.672
R11691 gnd.n6274 gnd.n2679 242.672
R11692 gnd.n6274 gnd.n2677 242.672
R11693 gnd.n1484 gnd.n1483 242.672
R11694 gnd.n1484 gnd.n1394 242.672
R11695 gnd.n1484 gnd.n1395 242.672
R11696 gnd.n1484 gnd.n1396 242.672
R11697 gnd.n1484 gnd.n1397 242.672
R11698 gnd.n1484 gnd.n1398 242.672
R11699 gnd.n1484 gnd.n1399 242.672
R11700 gnd.n1484 gnd.n1400 242.672
R11701 gnd.n1484 gnd.n1401 242.672
R11702 gnd.n1484 gnd.n1402 242.672
R11703 gnd.n1484 gnd.n1403 242.672
R11704 gnd.n1484 gnd.n1404 242.672
R11705 gnd.n1485 gnd.n1484 242.672
R11706 gnd.n2338 gnd.n891 242.672
R11707 gnd.n2338 gnd.n890 242.672
R11708 gnd.n2338 gnd.n889 242.672
R11709 gnd.n2338 gnd.n888 242.672
R11710 gnd.n2338 gnd.n887 242.672
R11711 gnd.n2338 gnd.n886 242.672
R11712 gnd.n2338 gnd.n885 242.672
R11713 gnd.n2338 gnd.n884 242.672
R11714 gnd.n2338 gnd.n883 242.672
R11715 gnd.n2338 gnd.n882 242.672
R11716 gnd.n2338 gnd.n881 242.672
R11717 gnd.n2338 gnd.n880 242.672
R11718 gnd.n2338 gnd.n879 242.672
R11719 gnd.n5280 gnd.n3048 242.672
R11720 gnd.n5297 gnd.n3048 242.672
R11721 gnd.n5299 gnd.n3048 242.672
R11722 gnd.n5316 gnd.n3048 242.672
R11723 gnd.n5318 gnd.n3048 242.672
R11724 gnd.n5335 gnd.n3048 242.672
R11725 gnd.n5337 gnd.n3048 242.672
R11726 gnd.n5355 gnd.n3048 242.672
R11727 gnd.n5357 gnd.n3048 242.672
R11728 gnd.n7660 gnd.n7659 242.672
R11729 gnd.n7659 gnd.n242 242.672
R11730 gnd.n7659 gnd.n191 242.672
R11731 gnd.n7659 gnd.n190 242.672
R11732 gnd.n7659 gnd.n189 242.672
R11733 gnd.n7659 gnd.n188 242.672
R11734 gnd.n7659 gnd.n187 242.672
R11735 gnd.n7659 gnd.n186 242.672
R11736 gnd.n7659 gnd.n185 242.672
R11737 gnd.n1568 gnd.n1567 242.672
R11738 gnd.n1567 gnd.n1306 242.672
R11739 gnd.n1567 gnd.n1307 242.672
R11740 gnd.n1567 gnd.n1308 242.672
R11741 gnd.n1567 gnd.n1309 242.672
R11742 gnd.n1567 gnd.n1310 242.672
R11743 gnd.n1567 gnd.n1311 242.672
R11744 gnd.n1567 gnd.n1312 242.672
R11745 gnd.n2338 gnd.n892 242.672
R11746 gnd.n2338 gnd.n893 242.672
R11747 gnd.n2338 gnd.n894 242.672
R11748 gnd.n2338 gnd.n895 242.672
R11749 gnd.n2338 gnd.n896 242.672
R11750 gnd.n2338 gnd.n897 242.672
R11751 gnd.n2338 gnd.n898 242.672
R11752 gnd.n2338 gnd.n899 242.672
R11753 gnd.n4064 gnd.n2363 242.672
R11754 gnd.n4072 gnd.n2363 242.672
R11755 gnd.n4074 gnd.n2363 242.672
R11756 gnd.n4082 gnd.n2363 242.672
R11757 gnd.n4084 gnd.n2363 242.672
R11758 gnd.n4092 gnd.n2363 242.672
R11759 gnd.n4094 gnd.n2363 242.672
R11760 gnd.n4102 gnd.n2363 242.672
R11761 gnd.n4104 gnd.n2363 242.672
R11762 gnd.n4112 gnd.n2363 242.672
R11763 gnd.n4114 gnd.n2363 242.672
R11764 gnd.n4122 gnd.n2363 242.672
R11765 gnd.n4124 gnd.n2363 242.672
R11766 gnd.n4132 gnd.n2363 242.672
R11767 gnd.n4134 gnd.n2363 242.672
R11768 gnd.n4142 gnd.n2363 242.672
R11769 gnd.n4144 gnd.n2363 242.672
R11770 gnd.n4152 gnd.n2363 242.672
R11771 gnd.n4154 gnd.n2363 242.672
R11772 gnd.n4164 gnd.n2363 242.672
R11773 gnd.n4166 gnd.n2363 242.672
R11774 gnd.n4174 gnd.n2363 242.672
R11775 gnd.n4176 gnd.n2363 242.672
R11776 gnd.n4184 gnd.n2363 242.672
R11777 gnd.n4186 gnd.n2363 242.672
R11778 gnd.n4194 gnd.n2363 242.672
R11779 gnd.n4196 gnd.n2363 242.672
R11780 gnd.n4205 gnd.n2363 242.672
R11781 gnd.n4208 gnd.n2363 242.672
R11782 gnd.n6274 gnd.n2691 242.672
R11783 gnd.n6274 gnd.n2692 242.672
R11784 gnd.n6274 gnd.n2693 242.672
R11785 gnd.n6274 gnd.n2694 242.672
R11786 gnd.n6274 gnd.n2695 242.672
R11787 gnd.n6274 gnd.n2696 242.672
R11788 gnd.n6274 gnd.n2697 242.672
R11789 gnd.n6274 gnd.n2698 242.672
R11790 gnd.n6274 gnd.n2699 242.672
R11791 gnd.n6274 gnd.n2700 242.672
R11792 gnd.n6274 gnd.n2701 242.672
R11793 gnd.n6274 gnd.n2702 242.672
R11794 gnd.n6274 gnd.n2703 242.672
R11795 gnd.n6274 gnd.n2704 242.672
R11796 gnd.n6274 gnd.n2705 242.672
R11797 gnd.n6274 gnd.n2706 242.672
R11798 gnd.n6224 gnd.n2752 242.672
R11799 gnd.n6274 gnd.n2707 242.672
R11800 gnd.n6274 gnd.n2708 242.672
R11801 gnd.n6274 gnd.n2709 242.672
R11802 gnd.n6274 gnd.n2710 242.672
R11803 gnd.n6274 gnd.n2711 242.672
R11804 gnd.n6274 gnd.n2712 242.672
R11805 gnd.n6274 gnd.n2713 242.672
R11806 gnd.n6274 gnd.n2714 242.672
R11807 gnd.n6274 gnd.n2715 242.672
R11808 gnd.n6274 gnd.n2716 242.672
R11809 gnd.n6274 gnd.n2717 242.672
R11810 gnd.n6274 gnd.n2718 242.672
R11811 gnd.n6274 gnd.n6273 242.672
R11812 gnd.n5575 gnd.n3048 242.672
R11813 gnd.n5578 gnd.n3048 242.672
R11814 gnd.n5586 gnd.n3048 242.672
R11815 gnd.n5588 gnd.n3048 242.672
R11816 gnd.n5596 gnd.n3048 242.672
R11817 gnd.n5598 gnd.n3048 242.672
R11818 gnd.n5606 gnd.n3048 242.672
R11819 gnd.n5608 gnd.n3048 242.672
R11820 gnd.n5619 gnd.n3048 242.672
R11821 gnd.n5621 gnd.n3048 242.672
R11822 gnd.n5629 gnd.n3048 242.672
R11823 gnd.n5631 gnd.n3048 242.672
R11824 gnd.n5640 gnd.n3048 242.672
R11825 gnd.n5641 gnd.n5546 242.672
R11826 gnd.n5642 gnd.n3048 242.672
R11827 gnd.n5644 gnd.n3048 242.672
R11828 gnd.n5652 gnd.n3048 242.672
R11829 gnd.n5654 gnd.n3048 242.672
R11830 gnd.n5662 gnd.n3048 242.672
R11831 gnd.n5664 gnd.n3048 242.672
R11832 gnd.n5674 gnd.n3048 242.672
R11833 gnd.n5676 gnd.n3048 242.672
R11834 gnd.n5684 gnd.n3048 242.672
R11835 gnd.n5686 gnd.n3048 242.672
R11836 gnd.n5694 gnd.n3048 242.672
R11837 gnd.n5696 gnd.n3048 242.672
R11838 gnd.n5704 gnd.n3048 242.672
R11839 gnd.n5706 gnd.n3048 242.672
R11840 gnd.n5715 gnd.n3048 242.672
R11841 gnd.n5718 gnd.n3048 242.672
R11842 gnd.n7659 gnd.n7447 242.672
R11843 gnd.n7659 gnd.n7448 242.672
R11844 gnd.n7659 gnd.n7449 242.672
R11845 gnd.n7659 gnd.n7450 242.672
R11846 gnd.n7659 gnd.n7451 242.672
R11847 gnd.n7659 gnd.n7452 242.672
R11848 gnd.n7659 gnd.n7453 242.672
R11849 gnd.n7659 gnd.n7454 242.672
R11850 gnd.n7659 gnd.n7455 242.672
R11851 gnd.n7659 gnd.n7456 242.672
R11852 gnd.n7659 gnd.n7457 242.672
R11853 gnd.n7659 gnd.n7458 242.672
R11854 gnd.n7659 gnd.n7459 242.672
R11855 gnd.n7659 gnd.n7460 242.672
R11856 gnd.n7659 gnd.n7461 242.672
R11857 gnd.n7659 gnd.n7462 242.672
R11858 gnd.n7659 gnd.n7463 242.672
R11859 gnd.n7659 gnd.n7464 242.672
R11860 gnd.n7659 gnd.n7465 242.672
R11861 gnd.n7659 gnd.n7466 242.672
R11862 gnd.n7659 gnd.n7467 242.672
R11863 gnd.n7659 gnd.n7468 242.672
R11864 gnd.n7659 gnd.n7469 242.672
R11865 gnd.n7659 gnd.n7470 242.672
R11866 gnd.n7659 gnd.n7471 242.672
R11867 gnd.n7659 gnd.n7472 242.672
R11868 gnd.n7659 gnd.n7473 242.672
R11869 gnd.n7659 gnd.n7474 242.672
R11870 gnd.n7659 gnd.n7658 242.672
R11871 gnd.n6339 gnd.n6338 242.672
R11872 gnd.n6339 gnd.n2588 242.672
R11873 gnd.n6339 gnd.n2589 242.672
R11874 gnd.n6339 gnd.n2590 242.672
R11875 gnd.n6339 gnd.n2591 242.672
R11876 gnd.n6339 gnd.n2592 242.672
R11877 gnd.n6339 gnd.n2593 242.672
R11878 gnd.n6339 gnd.n2594 242.672
R11879 gnd.n6339 gnd.n2595 242.672
R11880 gnd.n6339 gnd.n2596 242.672
R11881 gnd.n6339 gnd.n2597 242.672
R11882 gnd.n6339 gnd.n2598 242.672
R11883 gnd.n6339 gnd.n2600 242.672
R11884 gnd.n6340 gnd.n6339 242.672
R11885 gnd.n5346 gnd.n3047 242.672
R11886 gnd.n5222 gnd.n3047 242.672
R11887 gnd.n5327 gnd.n3047 242.672
R11888 gnd.n5231 gnd.n3047 242.672
R11889 gnd.n5308 gnd.n3047 242.672
R11890 gnd.n5240 gnd.n3047 242.672
R11891 gnd.n5289 gnd.n3047 242.672
R11892 gnd.n5249 gnd.n3047 242.672
R11893 gnd.n5274 gnd.n3047 242.672
R11894 gnd.n5252 gnd.n3047 242.672
R11895 gnd.n5263 gnd.n3047 242.672
R11896 gnd.n5256 gnd.n3047 242.672
R11897 gnd.n5368 gnd.n3047 242.672
R11898 gnd.n5365 gnd.n3047 242.672
R11899 gnd.n7475 gnd.n167 240.244
R11900 gnd.n7657 gnd.n7476 240.244
R11901 gnd.n7653 gnd.n7652 240.244
R11902 gnd.n7649 gnd.n7648 240.244
R11903 gnd.n7645 gnd.n7644 240.244
R11904 gnd.n7641 gnd.n7640 240.244
R11905 gnd.n7637 gnd.n7636 240.244
R11906 gnd.n7633 gnd.n7632 240.244
R11907 gnd.n7629 gnd.n7628 240.244
R11908 gnd.n7622 gnd.n7621 240.244
R11909 gnd.n7618 gnd.n7617 240.244
R11910 gnd.n7614 gnd.n7613 240.244
R11911 gnd.n7610 gnd.n7609 240.244
R11912 gnd.n7606 gnd.n7605 240.244
R11913 gnd.n7602 gnd.n7601 240.244
R11914 gnd.n7598 gnd.n7597 240.244
R11915 gnd.n7594 gnd.n7593 240.244
R11916 gnd.n7590 gnd.n7589 240.244
R11917 gnd.n7586 gnd.n7585 240.244
R11918 gnd.n7579 gnd.n7578 240.244
R11919 gnd.n7576 gnd.n7575 240.244
R11920 gnd.n7572 gnd.n7571 240.244
R11921 gnd.n7568 gnd.n7567 240.244
R11922 gnd.n7564 gnd.n7563 240.244
R11923 gnd.n7560 gnd.n7559 240.244
R11924 gnd.n7556 gnd.n7555 240.244
R11925 gnd.n7552 gnd.n7551 240.244
R11926 gnd.n7548 gnd.n7547 240.244
R11927 gnd.n7544 gnd.n7543 240.244
R11928 gnd.n3264 gnd.n3057 240.244
R11929 gnd.n3264 gnd.n3069 240.244
R11930 gnd.n5729 gnd.n3069 240.244
R11931 gnd.n5729 gnd.n3081 240.244
R11932 gnd.n5739 gnd.n3081 240.244
R11933 gnd.n5739 gnd.n3092 240.244
R11934 gnd.n3253 gnd.n3092 240.244
R11935 gnd.n3253 gnd.n3101 240.244
R11936 gnd.n5746 gnd.n3101 240.244
R11937 gnd.n5746 gnd.n3112 240.244
R11938 gnd.n5804 gnd.n3112 240.244
R11939 gnd.n5804 gnd.n3121 240.244
R11940 gnd.n5809 gnd.n3121 240.244
R11941 gnd.n5809 gnd.n3132 240.244
R11942 gnd.n5829 gnd.n3132 240.244
R11943 gnd.n5829 gnd.n3141 240.244
R11944 gnd.n3147 gnd.n3141 240.244
R11945 gnd.n5834 gnd.n3147 240.244
R11946 gnd.n5834 gnd.n5833 240.244
R11947 gnd.n5833 gnd.n3157 240.244
R11948 gnd.n3164 gnd.n3157 240.244
R11949 gnd.n5846 gnd.n3164 240.244
R11950 gnd.n5846 gnd.n70 240.244
R11951 gnd.n3173 gnd.n70 240.244
R11952 gnd.n5856 gnd.n3173 240.244
R11953 gnd.n5856 gnd.n87 240.244
R11954 gnd.n5860 gnd.n87 240.244
R11955 gnd.n5860 gnd.n99 240.244
R11956 gnd.n5871 gnd.n99 240.244
R11957 gnd.n5871 gnd.n109 240.244
R11958 gnd.n3227 gnd.n109 240.244
R11959 gnd.n3227 gnd.n118 240.244
R11960 gnd.n5906 gnd.n118 240.244
R11961 gnd.n5906 gnd.n129 240.244
R11962 gnd.n5902 gnd.n129 240.244
R11963 gnd.n5902 gnd.n139 240.244
R11964 gnd.n5894 gnd.n139 240.244
R11965 gnd.n5894 gnd.n150 240.244
R11966 gnd.n5890 gnd.n150 240.244
R11967 gnd.n5890 gnd.n160 240.244
R11968 gnd.n7669 gnd.n160 240.244
R11969 gnd.n7669 gnd.n169 240.244
R11970 gnd.n5577 gnd.n5576 240.244
R11971 gnd.n5579 gnd.n5577 240.244
R11972 gnd.n5585 gnd.n5567 240.244
R11973 gnd.n5589 gnd.n5587 240.244
R11974 gnd.n5595 gnd.n5563 240.244
R11975 gnd.n5599 gnd.n5597 240.244
R11976 gnd.n5605 gnd.n5559 240.244
R11977 gnd.n5609 gnd.n5607 240.244
R11978 gnd.n5618 gnd.n5555 240.244
R11979 gnd.n5622 gnd.n5620 240.244
R11980 gnd.n5628 gnd.n5551 240.244
R11981 gnd.n5632 gnd.n5630 240.244
R11982 gnd.n5639 gnd.n5547 240.244
R11983 gnd.n5645 gnd.n5643 240.244
R11984 gnd.n5651 gnd.n3295 240.244
R11985 gnd.n5655 gnd.n5653 240.244
R11986 gnd.n5661 gnd.n3291 240.244
R11987 gnd.n5665 gnd.n5663 240.244
R11988 gnd.n5673 gnd.n3287 240.244
R11989 gnd.n5677 gnd.n5675 240.244
R11990 gnd.n5683 gnd.n3283 240.244
R11991 gnd.n5687 gnd.n5685 240.244
R11992 gnd.n5693 gnd.n3279 240.244
R11993 gnd.n5697 gnd.n5695 240.244
R11994 gnd.n5703 gnd.n3275 240.244
R11995 gnd.n5707 gnd.n5705 240.244
R11996 gnd.n5714 gnd.n3271 240.244
R11997 gnd.n5717 gnd.n5716 240.244
R11998 gnd.n6000 gnd.n3062 240.244
R11999 gnd.n5996 gnd.n3062 240.244
R12000 gnd.n5996 gnd.n3067 240.244
R12001 gnd.n5988 gnd.n3067 240.244
R12002 gnd.n5988 gnd.n3084 240.244
R12003 gnd.n5984 gnd.n3084 240.244
R12004 gnd.n5984 gnd.n3090 240.244
R12005 gnd.n5976 gnd.n3090 240.244
R12006 gnd.n5976 gnd.n3104 240.244
R12007 gnd.n5972 gnd.n3104 240.244
R12008 gnd.n5972 gnd.n3110 240.244
R12009 gnd.n5964 gnd.n3110 240.244
R12010 gnd.n5964 gnd.n3124 240.244
R12011 gnd.n5960 gnd.n3124 240.244
R12012 gnd.n5960 gnd.n3130 240.244
R12013 gnd.n5952 gnd.n3130 240.244
R12014 gnd.n5952 gnd.n5950 240.244
R12015 gnd.n5950 gnd.n3144 240.244
R12016 gnd.n3161 gnd.n3144 240.244
R12017 gnd.n5939 gnd.n3161 240.244
R12018 gnd.n5939 gnd.n5936 240.244
R12019 gnd.n5936 gnd.n73 240.244
R12020 gnd.n7730 gnd.n73 240.244
R12021 gnd.n7730 gnd.n74 240.244
R12022 gnd.n84 gnd.n74 240.244
R12023 gnd.n7724 gnd.n84 240.244
R12024 gnd.n7724 gnd.n85 240.244
R12025 gnd.n7716 gnd.n85 240.244
R12026 gnd.n7716 gnd.n102 240.244
R12027 gnd.n7712 gnd.n102 240.244
R12028 gnd.n7712 gnd.n107 240.244
R12029 gnd.n7704 gnd.n107 240.244
R12030 gnd.n7704 gnd.n121 240.244
R12031 gnd.n7700 gnd.n121 240.244
R12032 gnd.n7700 gnd.n127 240.244
R12033 gnd.n7692 gnd.n127 240.244
R12034 gnd.n7692 gnd.n142 240.244
R12035 gnd.n7688 gnd.n142 240.244
R12036 gnd.n7688 gnd.n148 240.244
R12037 gnd.n7680 gnd.n148 240.244
R12038 gnd.n7680 gnd.n162 240.244
R12039 gnd.n7676 gnd.n162 240.244
R12040 gnd.n2719 gnd.n2570 240.244
R12041 gnd.n6272 gnd.n2720 240.244
R12042 gnd.n6268 gnd.n6267 240.244
R12043 gnd.n6264 gnd.n6263 240.244
R12044 gnd.n6260 gnd.n6259 240.244
R12045 gnd.n6256 gnd.n6255 240.244
R12046 gnd.n6252 gnd.n6251 240.244
R12047 gnd.n6248 gnd.n6247 240.244
R12048 gnd.n6244 gnd.n6243 240.244
R12049 gnd.n6239 gnd.n6238 240.244
R12050 gnd.n6235 gnd.n6234 240.244
R12051 gnd.n6231 gnd.n6230 240.244
R12052 gnd.n6227 gnd.n6226 240.244
R12053 gnd.n2845 gnd.n2844 240.244
R12054 gnd.n2842 gnd.n2841 240.244
R12055 gnd.n2838 gnd.n2837 240.244
R12056 gnd.n2834 gnd.n2833 240.244
R12057 gnd.n2830 gnd.n2829 240.244
R12058 gnd.n2823 gnd.n2822 240.244
R12059 gnd.n2820 gnd.n2819 240.244
R12060 gnd.n2816 gnd.n2815 240.244
R12061 gnd.n2812 gnd.n2811 240.244
R12062 gnd.n2808 gnd.n2807 240.244
R12063 gnd.n2804 gnd.n2803 240.244
R12064 gnd.n2800 gnd.n2799 240.244
R12065 gnd.n2796 gnd.n2795 240.244
R12066 gnd.n2792 gnd.n2791 240.244
R12067 gnd.n2788 gnd.n2787 240.244
R12068 gnd.n3924 gnd.n2364 240.244
R12069 gnd.n3924 gnd.n2375 240.244
R12070 gnd.n4249 gnd.n2375 240.244
R12071 gnd.n4249 gnd.n2387 240.244
R12072 gnd.n4245 gnd.n2387 240.244
R12073 gnd.n4245 gnd.n2398 240.244
R12074 gnd.n4237 gnd.n2398 240.244
R12075 gnd.n4237 gnd.n2408 240.244
R12076 gnd.n4233 gnd.n2408 240.244
R12077 gnd.n4233 gnd.n2419 240.244
R12078 gnd.n3908 gnd.n2419 240.244
R12079 gnd.n3908 gnd.n2428 240.244
R12080 gnd.n4296 gnd.n2428 240.244
R12081 gnd.n4296 gnd.n2439 240.244
R12082 gnd.n4300 gnd.n2439 240.244
R12083 gnd.n4300 gnd.n2449 240.244
R12084 gnd.n4311 gnd.n2449 240.244
R12085 gnd.n4311 gnd.n2458 240.244
R12086 gnd.n3890 gnd.n2458 240.244
R12087 gnd.n3890 gnd.n2467 240.244
R12088 gnd.n4318 gnd.n2467 240.244
R12089 gnd.n4318 gnd.n2475 240.244
R12090 gnd.n4333 gnd.n2475 240.244
R12091 gnd.n4333 gnd.n2484 240.244
R12092 gnd.n4340 gnd.n2484 240.244
R12093 gnd.n4340 gnd.n2492 240.244
R12094 gnd.n3874 gnd.n2492 240.244
R12095 gnd.n3874 gnd.n2501 240.244
R12096 gnd.n4399 gnd.n2501 240.244
R12097 gnd.n4399 gnd.n2512 240.244
R12098 gnd.n4403 gnd.n2512 240.244
R12099 gnd.n4403 gnd.n2521 240.244
R12100 gnd.n4413 gnd.n2521 240.244
R12101 gnd.n4413 gnd.n2532 240.244
R12102 gnd.n3857 gnd.n2532 240.244
R12103 gnd.n3857 gnd.n2541 240.244
R12104 gnd.n4420 gnd.n2541 240.244
R12105 gnd.n4420 gnd.n2552 240.244
R12106 gnd.n4424 gnd.n2552 240.244
R12107 gnd.n4424 gnd.n2562 240.244
R12108 gnd.n6351 gnd.n2562 240.244
R12109 gnd.n6351 gnd.n2572 240.244
R12110 gnd.n4065 gnd.n4060 240.244
R12111 gnd.n4071 gnd.n4060 240.244
R12112 gnd.n4075 gnd.n4073 240.244
R12113 gnd.n4081 gnd.n4056 240.244
R12114 gnd.n4085 gnd.n4083 240.244
R12115 gnd.n4091 gnd.n4052 240.244
R12116 gnd.n4095 gnd.n4093 240.244
R12117 gnd.n4101 gnd.n4048 240.244
R12118 gnd.n4105 gnd.n4103 240.244
R12119 gnd.n4111 gnd.n4041 240.244
R12120 gnd.n4115 gnd.n4113 240.244
R12121 gnd.n4121 gnd.n4037 240.244
R12122 gnd.n4125 gnd.n4123 240.244
R12123 gnd.n4131 gnd.n4033 240.244
R12124 gnd.n4135 gnd.n4133 240.244
R12125 gnd.n4141 gnd.n4029 240.244
R12126 gnd.n4145 gnd.n4143 240.244
R12127 gnd.n4151 gnd.n4025 240.244
R12128 gnd.n4155 gnd.n4153 240.244
R12129 gnd.n4163 gnd.n4021 240.244
R12130 gnd.n4167 gnd.n4165 240.244
R12131 gnd.n4173 gnd.n4017 240.244
R12132 gnd.n4177 gnd.n4175 240.244
R12133 gnd.n4183 gnd.n4013 240.244
R12134 gnd.n4187 gnd.n4185 240.244
R12135 gnd.n4193 gnd.n4009 240.244
R12136 gnd.n4197 gnd.n4195 240.244
R12137 gnd.n4204 gnd.n4005 240.244
R12138 gnd.n4207 gnd.n4206 240.244
R12139 gnd.n6485 gnd.n2369 240.244
R12140 gnd.n6481 gnd.n2369 240.244
R12141 gnd.n6481 gnd.n2374 240.244
R12142 gnd.n6473 gnd.n2374 240.244
R12143 gnd.n6473 gnd.n2390 240.244
R12144 gnd.n6469 gnd.n2390 240.244
R12145 gnd.n6469 gnd.n2396 240.244
R12146 gnd.n6461 gnd.n2396 240.244
R12147 gnd.n6461 gnd.n2411 240.244
R12148 gnd.n6457 gnd.n2411 240.244
R12149 gnd.n6457 gnd.n2417 240.244
R12150 gnd.n6449 gnd.n2417 240.244
R12151 gnd.n6449 gnd.n2431 240.244
R12152 gnd.n6445 gnd.n2431 240.244
R12153 gnd.n6445 gnd.n2437 240.244
R12154 gnd.n6437 gnd.n2437 240.244
R12155 gnd.n6437 gnd.n2452 240.244
R12156 gnd.n6432 gnd.n2452 240.244
R12157 gnd.n6432 gnd.n2456 240.244
R12158 gnd.n6424 gnd.n2456 240.244
R12159 gnd.n6424 gnd.n2470 240.244
R12160 gnd.n6419 gnd.n2470 240.244
R12161 gnd.n6419 gnd.n2473 240.244
R12162 gnd.n6411 gnd.n2473 240.244
R12163 gnd.n6411 gnd.n2487 240.244
R12164 gnd.n6406 gnd.n2487 240.244
R12165 gnd.n6406 gnd.n2490 240.244
R12166 gnd.n6398 gnd.n2490 240.244
R12167 gnd.n6398 gnd.n2504 240.244
R12168 gnd.n6394 gnd.n2504 240.244
R12169 gnd.n6394 gnd.n2510 240.244
R12170 gnd.n6386 gnd.n2510 240.244
R12171 gnd.n6386 gnd.n2524 240.244
R12172 gnd.n6382 gnd.n2524 240.244
R12173 gnd.n6382 gnd.n2530 240.244
R12174 gnd.n6374 gnd.n2530 240.244
R12175 gnd.n6374 gnd.n2544 240.244
R12176 gnd.n6370 gnd.n2544 240.244
R12177 gnd.n6370 gnd.n2550 240.244
R12178 gnd.n6362 gnd.n2550 240.244
R12179 gnd.n6362 gnd.n2565 240.244
R12180 gnd.n6358 gnd.n2565 240.244
R12181 gnd.n2337 gnd.n901 240.244
R12182 gnd.n2330 gnd.n2329 240.244
R12183 gnd.n2327 gnd.n2326 240.244
R12184 gnd.n2323 gnd.n2322 240.244
R12185 gnd.n2319 gnd.n2318 240.244
R12186 gnd.n2315 gnd.n2314 240.244
R12187 gnd.n2311 gnd.n2310 240.244
R12188 gnd.n2307 gnd.n2306 240.244
R12189 gnd.n1579 gnd.n1291 240.244
R12190 gnd.n1589 gnd.n1291 240.244
R12191 gnd.n1589 gnd.n1282 240.244
R12192 gnd.n1282 gnd.n1271 240.244
R12193 gnd.n1610 gnd.n1271 240.244
R12194 gnd.n1610 gnd.n1265 240.244
R12195 gnd.n1620 gnd.n1265 240.244
R12196 gnd.n1620 gnd.n1254 240.244
R12197 gnd.n1254 gnd.n1246 240.244
R12198 gnd.n1638 gnd.n1246 240.244
R12199 gnd.n1639 gnd.n1638 240.244
R12200 gnd.n1639 gnd.n1231 240.244
R12201 gnd.n1641 gnd.n1231 240.244
R12202 gnd.n1641 gnd.n1217 240.244
R12203 gnd.n1683 gnd.n1217 240.244
R12204 gnd.n1684 gnd.n1683 240.244
R12205 gnd.n1687 gnd.n1684 240.244
R12206 gnd.n1687 gnd.n1172 240.244
R12207 gnd.n1212 gnd.n1172 240.244
R12208 gnd.n1212 gnd.n1182 240.244
R12209 gnd.n1697 gnd.n1182 240.244
R12210 gnd.n1697 gnd.n1203 240.244
R12211 gnd.n1707 gnd.n1203 240.244
R12212 gnd.n1707 gnd.n1101 240.244
R12213 gnd.n1752 gnd.n1101 240.244
R12214 gnd.n1752 gnd.n1087 240.244
R12215 gnd.n1774 gnd.n1087 240.244
R12216 gnd.n1775 gnd.n1774 240.244
R12217 gnd.n1775 gnd.n1074 240.244
R12218 gnd.n1074 gnd.n1063 240.244
R12219 gnd.n1806 gnd.n1063 240.244
R12220 gnd.n1807 gnd.n1806 240.244
R12221 gnd.n1808 gnd.n1807 240.244
R12222 gnd.n1808 gnd.n1048 240.244
R12223 gnd.n1839 gnd.n1048 240.244
R12224 gnd.n1839 gnd.n1034 240.244
R12225 gnd.n1861 gnd.n1034 240.244
R12226 gnd.n1862 gnd.n1861 240.244
R12227 gnd.n1862 gnd.n1021 240.244
R12228 gnd.n1021 gnd.n1010 240.244
R12229 gnd.n1893 gnd.n1010 240.244
R12230 gnd.n1894 gnd.n1893 240.244
R12231 gnd.n1895 gnd.n1894 240.244
R12232 gnd.n1895 gnd.n994 240.244
R12233 gnd.n994 gnd.n993 240.244
R12234 gnd.n993 gnd.n980 240.244
R12235 gnd.n1950 gnd.n980 240.244
R12236 gnd.n1951 gnd.n1950 240.244
R12237 gnd.n1951 gnd.n967 240.244
R12238 gnd.n967 gnd.n957 240.244
R12239 gnd.n2238 gnd.n957 240.244
R12240 gnd.n2241 gnd.n2238 240.244
R12241 gnd.n2241 gnd.n2240 240.244
R12242 gnd.n1569 gnd.n1304 240.244
R12243 gnd.n1325 gnd.n1304 240.244
R12244 gnd.n1328 gnd.n1327 240.244
R12245 gnd.n1335 gnd.n1334 240.244
R12246 gnd.n1338 gnd.n1337 240.244
R12247 gnd.n1345 gnd.n1344 240.244
R12248 gnd.n1348 gnd.n1347 240.244
R12249 gnd.n1355 gnd.n1354 240.244
R12250 gnd.n1577 gnd.n1301 240.244
R12251 gnd.n1301 gnd.n1280 240.244
R12252 gnd.n1600 gnd.n1280 240.244
R12253 gnd.n1600 gnd.n1274 240.244
R12254 gnd.n1608 gnd.n1274 240.244
R12255 gnd.n1608 gnd.n1276 240.244
R12256 gnd.n1276 gnd.n1252 240.244
R12257 gnd.n1630 gnd.n1252 240.244
R12258 gnd.n1630 gnd.n1248 240.244
R12259 gnd.n1636 gnd.n1248 240.244
R12260 gnd.n1636 gnd.n1230 240.244
R12261 gnd.n1661 gnd.n1230 240.244
R12262 gnd.n1661 gnd.n1225 240.244
R12263 gnd.n1673 gnd.n1225 240.244
R12264 gnd.n1673 gnd.n1226 240.244
R12265 gnd.n1669 gnd.n1226 240.244
R12266 gnd.n1669 gnd.n1174 240.244
R12267 gnd.n1721 gnd.n1174 240.244
R12268 gnd.n1721 gnd.n1175 240.244
R12269 gnd.n1717 gnd.n1175 240.244
R12270 gnd.n1717 gnd.n1181 240.244
R12271 gnd.n1201 gnd.n1181 240.244
R12272 gnd.n1201 gnd.n1099 240.244
R12273 gnd.n1756 gnd.n1099 240.244
R12274 gnd.n1756 gnd.n1094 240.244
R12275 gnd.n1764 gnd.n1094 240.244
R12276 gnd.n1764 gnd.n1095 240.244
R12277 gnd.n1095 gnd.n1072 240.244
R12278 gnd.n1796 gnd.n1072 240.244
R12279 gnd.n1796 gnd.n1067 240.244
R12280 gnd.n1804 gnd.n1067 240.244
R12281 gnd.n1804 gnd.n1068 240.244
R12282 gnd.n1068 gnd.n1046 240.244
R12283 gnd.n1843 gnd.n1046 240.244
R12284 gnd.n1843 gnd.n1041 240.244
R12285 gnd.n1851 gnd.n1041 240.244
R12286 gnd.n1851 gnd.n1042 240.244
R12287 gnd.n1042 gnd.n1019 240.244
R12288 gnd.n1883 gnd.n1019 240.244
R12289 gnd.n1883 gnd.n1014 240.244
R12290 gnd.n1891 gnd.n1014 240.244
R12291 gnd.n1891 gnd.n1015 240.244
R12292 gnd.n1015 gnd.n992 240.244
R12293 gnd.n1932 gnd.n992 240.244
R12294 gnd.n1932 gnd.n987 240.244
R12295 gnd.n1940 gnd.n987 240.244
R12296 gnd.n1940 gnd.n988 240.244
R12297 gnd.n988 gnd.n965 240.244
R12298 gnd.n2226 gnd.n965 240.244
R12299 gnd.n2226 gnd.n960 240.244
R12300 gnd.n2236 gnd.n960 240.244
R12301 gnd.n2236 gnd.n961 240.244
R12302 gnd.n961 gnd.n900 240.244
R12303 gnd.n203 gnd.n172 240.244
R12304 gnd.n206 gnd.n205 240.244
R12305 gnd.n213 gnd.n212 240.244
R12306 gnd.n216 gnd.n215 240.244
R12307 gnd.n223 gnd.n222 240.244
R12308 gnd.n226 gnd.n225 240.244
R12309 gnd.n233 gnd.n232 240.244
R12310 gnd.n235 gnd.n192 240.244
R12311 gnd.n241 gnd.n183 240.244
R12312 gnd.n5196 gnd.n3058 240.244
R12313 gnd.n5196 gnd.n3070 240.244
R12314 gnd.n5731 gnd.n3070 240.244
R12315 gnd.n5731 gnd.n3082 240.244
R12316 gnd.n5737 gnd.n3082 240.244
R12317 gnd.n5737 gnd.n3093 240.244
R12318 gnd.n5757 gnd.n3093 240.244
R12319 gnd.n5757 gnd.n3102 240.244
R12320 gnd.n5748 gnd.n3102 240.244
R12321 gnd.n5748 gnd.n3113 240.244
R12322 gnd.n3247 gnd.n3113 240.244
R12323 gnd.n3247 gnd.n3122 240.244
R12324 gnd.n5811 gnd.n3122 240.244
R12325 gnd.n5811 gnd.n3133 240.244
R12326 gnd.n5827 gnd.n3133 240.244
R12327 gnd.n5827 gnd.n3142 240.244
R12328 gnd.n3148 gnd.n3142 240.244
R12329 gnd.n5816 gnd.n3148 240.244
R12330 gnd.n5817 gnd.n5816 240.244
R12331 gnd.n5817 gnd.n3158 240.244
R12332 gnd.n3165 gnd.n3158 240.244
R12333 gnd.n3165 gnd.n66 240.244
R12334 gnd.n7732 gnd.n66 240.244
R12335 gnd.n7732 gnd.n68 240.244
R12336 gnd.n5854 gnd.n68 240.244
R12337 gnd.n5854 gnd.n88 240.244
R12338 gnd.n5862 gnd.n88 240.244
R12339 gnd.n5862 gnd.n100 240.244
R12340 gnd.n5869 gnd.n100 240.244
R12341 gnd.n5869 gnd.n110 240.244
R12342 gnd.n5912 gnd.n110 240.244
R12343 gnd.n5912 gnd.n119 240.244
R12344 gnd.n5908 gnd.n119 240.244
R12345 gnd.n5908 gnd.n130 240.244
R12346 gnd.n5900 gnd.n130 240.244
R12347 gnd.n5900 gnd.n140 240.244
R12348 gnd.n5896 gnd.n140 240.244
R12349 gnd.n5896 gnd.n151 240.244
R12350 gnd.n5888 gnd.n151 240.244
R12351 gnd.n5888 gnd.n161 240.244
R12352 gnd.n7667 gnd.n161 240.244
R12353 gnd.n7667 gnd.n170 240.244
R12354 gnd.n5296 gnd.n5244 240.244
R12355 gnd.n5300 gnd.n5298 240.244
R12356 gnd.n5315 gnd.n5235 240.244
R12357 gnd.n5319 gnd.n5317 240.244
R12358 gnd.n5334 gnd.n5226 240.244
R12359 gnd.n5338 gnd.n5336 240.244
R12360 gnd.n5354 gnd.n5217 240.244
R12361 gnd.n5358 gnd.n5356 240.244
R12362 gnd.n5213 gnd.n5212 240.244
R12363 gnd.n3072 gnd.n3060 240.244
R12364 gnd.n5994 gnd.n3072 240.244
R12365 gnd.n5994 gnd.n3073 240.244
R12366 gnd.n5990 gnd.n3073 240.244
R12367 gnd.n5990 gnd.n3079 240.244
R12368 gnd.n5982 gnd.n3079 240.244
R12369 gnd.n5982 gnd.n3094 240.244
R12370 gnd.n5978 gnd.n3094 240.244
R12371 gnd.n5978 gnd.n3099 240.244
R12372 gnd.n5970 gnd.n3099 240.244
R12373 gnd.n5970 gnd.n3115 240.244
R12374 gnd.n5966 gnd.n3115 240.244
R12375 gnd.n5966 gnd.n3120 240.244
R12376 gnd.n5958 gnd.n3120 240.244
R12377 gnd.n5958 gnd.n3134 240.244
R12378 gnd.n5954 gnd.n3134 240.244
R12379 gnd.n5954 gnd.n3139 240.244
R12380 gnd.n5838 gnd.n3139 240.244
R12381 gnd.n5839 gnd.n5838 240.244
R12382 gnd.n5839 gnd.n3160 240.244
R12383 gnd.n5934 gnd.n3160 240.244
R12384 gnd.n5934 gnd.n3167 240.244
R12385 gnd.n3167 gnd.n72 240.244
R12386 gnd.n5929 gnd.n72 240.244
R12387 gnd.n5929 gnd.n90 240.244
R12388 gnd.n7722 gnd.n90 240.244
R12389 gnd.n7722 gnd.n91 240.244
R12390 gnd.n7718 gnd.n91 240.244
R12391 gnd.n7718 gnd.n97 240.244
R12392 gnd.n7710 gnd.n97 240.244
R12393 gnd.n7710 gnd.n111 240.244
R12394 gnd.n7706 gnd.n111 240.244
R12395 gnd.n7706 gnd.n116 240.244
R12396 gnd.n7698 gnd.n116 240.244
R12397 gnd.n7698 gnd.n132 240.244
R12398 gnd.n7694 gnd.n132 240.244
R12399 gnd.n7694 gnd.n137 240.244
R12400 gnd.n7686 gnd.n137 240.244
R12401 gnd.n7686 gnd.n153 240.244
R12402 gnd.n7682 gnd.n153 240.244
R12403 gnd.n7682 gnd.n158 240.244
R12404 gnd.n7674 gnd.n158 240.244
R12405 gnd.n920 gnd.n878 240.244
R12406 gnd.n2297 gnd.n2296 240.244
R12407 gnd.n2293 gnd.n2292 240.244
R12408 gnd.n2289 gnd.n2288 240.244
R12409 gnd.n2285 gnd.n2284 240.244
R12410 gnd.n2281 gnd.n2280 240.244
R12411 gnd.n2277 gnd.n2276 240.244
R12412 gnd.n2273 gnd.n2272 240.244
R12413 gnd.n2269 gnd.n2268 240.244
R12414 gnd.n2265 gnd.n2264 240.244
R12415 gnd.n2261 gnd.n2260 240.244
R12416 gnd.n2257 gnd.n2256 240.244
R12417 gnd.n2253 gnd.n2252 240.244
R12418 gnd.n1492 gnd.n1389 240.244
R12419 gnd.n1492 gnd.n1382 240.244
R12420 gnd.n1503 gnd.n1382 240.244
R12421 gnd.n1503 gnd.n1378 240.244
R12422 gnd.n1509 gnd.n1378 240.244
R12423 gnd.n1509 gnd.n1370 240.244
R12424 gnd.n1519 gnd.n1370 240.244
R12425 gnd.n1519 gnd.n1365 240.244
R12426 gnd.n1555 gnd.n1365 240.244
R12427 gnd.n1555 gnd.n1366 240.244
R12428 gnd.n1366 gnd.n1313 240.244
R12429 gnd.n1550 gnd.n1313 240.244
R12430 gnd.n1550 gnd.n1549 240.244
R12431 gnd.n1549 gnd.n1292 240.244
R12432 gnd.n1545 gnd.n1292 240.244
R12433 gnd.n1545 gnd.n1283 240.244
R12434 gnd.n1542 gnd.n1283 240.244
R12435 gnd.n1542 gnd.n1541 240.244
R12436 gnd.n1541 gnd.n1266 240.244
R12437 gnd.n1537 gnd.n1266 240.244
R12438 gnd.n1537 gnd.n1255 240.244
R12439 gnd.n1255 gnd.n1236 240.244
R12440 gnd.n1650 gnd.n1236 240.244
R12441 gnd.n1650 gnd.n1232 240.244
R12442 gnd.n1658 gnd.n1232 240.244
R12443 gnd.n1658 gnd.n1223 240.244
R12444 gnd.n1223 gnd.n1159 240.244
R12445 gnd.n1730 gnd.n1159 240.244
R12446 gnd.n1730 gnd.n1160 240.244
R12447 gnd.n1171 gnd.n1160 240.244
R12448 gnd.n1206 gnd.n1171 240.244
R12449 gnd.n1209 gnd.n1206 240.244
R12450 gnd.n1209 gnd.n1183 240.244
R12451 gnd.n1196 gnd.n1183 240.244
R12452 gnd.n1196 gnd.n1193 240.244
R12453 gnd.n1193 gnd.n1102 240.244
R12454 gnd.n1751 gnd.n1102 240.244
R12455 gnd.n1751 gnd.n1092 240.244
R12456 gnd.n1747 gnd.n1092 240.244
R12457 gnd.n1747 gnd.n1086 240.244
R12458 gnd.n1744 gnd.n1086 240.244
R12459 gnd.n1744 gnd.n1075 240.244
R12460 gnd.n1741 gnd.n1075 240.244
R12461 gnd.n1741 gnd.n1053 240.244
R12462 gnd.n1817 gnd.n1053 240.244
R12463 gnd.n1817 gnd.n1049 240.244
R12464 gnd.n1838 gnd.n1049 240.244
R12465 gnd.n1838 gnd.n1039 240.244
R12466 gnd.n1834 gnd.n1039 240.244
R12467 gnd.n1834 gnd.n1033 240.244
R12468 gnd.n1831 gnd.n1033 240.244
R12469 gnd.n1831 gnd.n1022 240.244
R12470 gnd.n1828 gnd.n1022 240.244
R12471 gnd.n1828 gnd.n999 240.244
R12472 gnd.n1904 gnd.n999 240.244
R12473 gnd.n1904 gnd.n995 240.244
R12474 gnd.n1929 gnd.n995 240.244
R12475 gnd.n1929 gnd.n986 240.244
R12476 gnd.n1925 gnd.n986 240.244
R12477 gnd.n1925 gnd.n979 240.244
R12478 gnd.n1921 gnd.n979 240.244
R12479 gnd.n1921 gnd.n968 240.244
R12480 gnd.n1918 gnd.n968 240.244
R12481 gnd.n1918 gnd.n949 240.244
R12482 gnd.n2248 gnd.n949 240.244
R12483 gnd.n1406 gnd.n1405 240.244
R12484 gnd.n1477 gnd.n1405 240.244
R12485 gnd.n1475 gnd.n1474 240.244
R12486 gnd.n1471 gnd.n1470 240.244
R12487 gnd.n1467 gnd.n1466 240.244
R12488 gnd.n1463 gnd.n1462 240.244
R12489 gnd.n1459 gnd.n1458 240.244
R12490 gnd.n1455 gnd.n1454 240.244
R12491 gnd.n1451 gnd.n1450 240.244
R12492 gnd.n1447 gnd.n1446 240.244
R12493 gnd.n1443 gnd.n1442 240.244
R12494 gnd.n1439 gnd.n1438 240.244
R12495 gnd.n1435 gnd.n1393 240.244
R12496 gnd.n1495 gnd.n1387 240.244
R12497 gnd.n1495 gnd.n1383 240.244
R12498 gnd.n1501 gnd.n1383 240.244
R12499 gnd.n1501 gnd.n1376 240.244
R12500 gnd.n1511 gnd.n1376 240.244
R12501 gnd.n1511 gnd.n1372 240.244
R12502 gnd.n1517 gnd.n1372 240.244
R12503 gnd.n1517 gnd.n1363 240.244
R12504 gnd.n1557 gnd.n1363 240.244
R12505 gnd.n1557 gnd.n1314 240.244
R12506 gnd.n1565 gnd.n1314 240.244
R12507 gnd.n1565 gnd.n1315 240.244
R12508 gnd.n1315 gnd.n1293 240.244
R12509 gnd.n1586 gnd.n1293 240.244
R12510 gnd.n1586 gnd.n1285 240.244
R12511 gnd.n1597 gnd.n1285 240.244
R12512 gnd.n1597 gnd.n1286 240.244
R12513 gnd.n1286 gnd.n1267 240.244
R12514 gnd.n1617 gnd.n1267 240.244
R12515 gnd.n1617 gnd.n1257 240.244
R12516 gnd.n1627 gnd.n1257 240.244
R12517 gnd.n1627 gnd.n1238 240.244
R12518 gnd.n1648 gnd.n1238 240.244
R12519 gnd.n1648 gnd.n1240 240.244
R12520 gnd.n1240 gnd.n1221 240.244
R12521 gnd.n1676 gnd.n1221 240.244
R12522 gnd.n1676 gnd.n1163 240.244
R12523 gnd.n1728 gnd.n1163 240.244
R12524 gnd.n1728 gnd.n1164 240.244
R12525 gnd.n1724 gnd.n1164 240.244
R12526 gnd.n1724 gnd.n1170 240.244
R12527 gnd.n1185 gnd.n1170 240.244
R12528 gnd.n1714 gnd.n1185 240.244
R12529 gnd.n1714 gnd.n1186 240.244
R12530 gnd.n1710 gnd.n1186 240.244
R12531 gnd.n1710 gnd.n1192 240.244
R12532 gnd.n1192 gnd.n1091 240.244
R12533 gnd.n1767 gnd.n1091 240.244
R12534 gnd.n1767 gnd.n1084 240.244
R12535 gnd.n1778 gnd.n1084 240.244
R12536 gnd.n1778 gnd.n1077 240.244
R12537 gnd.n1793 gnd.n1077 240.244
R12538 gnd.n1793 gnd.n1078 240.244
R12539 gnd.n1078 gnd.n1056 240.244
R12540 gnd.n1815 gnd.n1056 240.244
R12541 gnd.n1815 gnd.n1057 240.244
R12542 gnd.n1057 gnd.n1038 240.244
R12543 gnd.n1854 gnd.n1038 240.244
R12544 gnd.n1854 gnd.n1031 240.244
R12545 gnd.n1865 gnd.n1031 240.244
R12546 gnd.n1865 gnd.n1024 240.244
R12547 gnd.n1880 gnd.n1024 240.244
R12548 gnd.n1880 gnd.n1025 240.244
R12549 gnd.n1025 gnd.n1002 240.244
R12550 gnd.n1902 gnd.n1002 240.244
R12551 gnd.n1902 gnd.n1004 240.244
R12552 gnd.n1004 gnd.n984 240.244
R12553 gnd.n1943 gnd.n984 240.244
R12554 gnd.n1943 gnd.n977 240.244
R12555 gnd.n1954 gnd.n977 240.244
R12556 gnd.n1954 gnd.n970 240.244
R12557 gnd.n2223 gnd.n970 240.244
R12558 gnd.n2223 gnd.n971 240.244
R12559 gnd.n971 gnd.n952 240.244
R12560 gnd.n2246 gnd.n952 240.244
R12561 gnd.n2621 gnd.n2575 240.244
R12562 gnd.n2678 gnd.n2622 240.244
R12563 gnd.n2632 gnd.n2631 240.244
R12564 gnd.n2680 gnd.n2639 240.244
R12565 gnd.n2683 gnd.n2640 240.244
R12566 gnd.n2650 gnd.n2649 240.244
R12567 gnd.n2685 gnd.n2657 240.244
R12568 gnd.n2688 gnd.n2658 240.244
R12569 gnd.n2675 gnd.n2670 240.244
R12570 gnd.n4255 gnd.n2365 240.244
R12571 gnd.n4255 gnd.n2376 240.244
R12572 gnd.n4251 gnd.n2376 240.244
R12573 gnd.n4251 gnd.n2388 240.244
R12574 gnd.n4243 gnd.n2388 240.244
R12575 gnd.n4243 gnd.n2399 240.244
R12576 gnd.n4239 gnd.n2399 240.244
R12577 gnd.n4239 gnd.n2409 240.244
R12578 gnd.n4231 gnd.n2409 240.244
R12579 gnd.n4231 gnd.n2420 240.244
R12580 gnd.n4288 gnd.n2420 240.244
R12581 gnd.n4288 gnd.n2429 240.244
R12582 gnd.n4294 gnd.n2429 240.244
R12583 gnd.n4294 gnd.n2440 240.244
R12584 gnd.n4302 gnd.n2440 240.244
R12585 gnd.n4302 gnd.n2450 240.244
R12586 gnd.n4309 gnd.n2450 240.244
R12587 gnd.n4309 gnd.n2459 240.244
R12588 gnd.n4353 gnd.n2459 240.244
R12589 gnd.n4353 gnd.n2468 240.244
R12590 gnd.n3894 gnd.n2468 240.244
R12591 gnd.n3894 gnd.n2476 240.244
R12592 gnd.n3897 gnd.n2476 240.244
R12593 gnd.n3897 gnd.n2485 240.244
R12594 gnd.n4342 gnd.n2485 240.244
R12595 gnd.n4342 gnd.n2493 240.244
R12596 gnd.n4391 gnd.n2493 240.244
R12597 gnd.n4391 gnd.n2502 240.244
R12598 gnd.n4397 gnd.n2502 240.244
R12599 gnd.n4397 gnd.n2513 240.244
R12600 gnd.n4405 gnd.n2513 240.244
R12601 gnd.n4405 gnd.n2522 240.244
R12602 gnd.n4411 gnd.n2522 240.244
R12603 gnd.n4411 gnd.n2533 240.244
R12604 gnd.n4435 gnd.n2533 240.244
R12605 gnd.n4435 gnd.n2542 240.244
R12606 gnd.n3862 gnd.n2542 240.244
R12607 gnd.n3862 gnd.n2553 240.244
R12608 gnd.n4426 gnd.n2553 240.244
R12609 gnd.n4426 gnd.n2563 240.244
R12610 gnd.n6349 gnd.n2563 240.244
R12611 gnd.n6349 gnd.n2573 240.244
R12612 gnd.n3995 gnd.n3994 240.244
R12613 gnd.n3991 gnd.n3990 240.244
R12614 gnd.n3988 gnd.n3937 240.244
R12615 gnd.n3984 gnd.n3982 240.244
R12616 gnd.n3980 gnd.n3943 240.244
R12617 gnd.n3976 gnd.n3974 240.244
R12618 gnd.n3972 gnd.n3949 240.244
R12619 gnd.n3968 gnd.n3966 240.244
R12620 gnd.n3964 gnd.n3955 240.244
R12621 gnd.n2378 gnd.n2367 240.244
R12622 gnd.n6479 gnd.n2378 240.244
R12623 gnd.n6479 gnd.n2379 240.244
R12624 gnd.n6475 gnd.n2379 240.244
R12625 gnd.n6475 gnd.n2385 240.244
R12626 gnd.n6467 gnd.n2385 240.244
R12627 gnd.n6467 gnd.n2401 240.244
R12628 gnd.n6463 gnd.n2401 240.244
R12629 gnd.n6463 gnd.n2406 240.244
R12630 gnd.n6455 gnd.n2406 240.244
R12631 gnd.n6455 gnd.n2422 240.244
R12632 gnd.n6451 gnd.n2422 240.244
R12633 gnd.n6451 gnd.n2427 240.244
R12634 gnd.n6443 gnd.n2427 240.244
R12635 gnd.n6443 gnd.n2442 240.244
R12636 gnd.n6439 gnd.n2442 240.244
R12637 gnd.n6439 gnd.n2447 240.244
R12638 gnd.n6430 gnd.n2447 240.244
R12639 gnd.n6430 gnd.n2461 240.244
R12640 gnd.n6426 gnd.n2461 240.244
R12641 gnd.n6426 gnd.n2466 240.244
R12642 gnd.n6417 gnd.n2466 240.244
R12643 gnd.n6417 gnd.n2477 240.244
R12644 gnd.n6413 gnd.n2477 240.244
R12645 gnd.n6413 gnd.n2482 240.244
R12646 gnd.n6404 gnd.n2482 240.244
R12647 gnd.n6404 gnd.n2495 240.244
R12648 gnd.n6400 gnd.n2495 240.244
R12649 gnd.n6400 gnd.n2500 240.244
R12650 gnd.n6392 gnd.n2500 240.244
R12651 gnd.n6392 gnd.n2514 240.244
R12652 gnd.n6388 gnd.n2514 240.244
R12653 gnd.n6388 gnd.n2519 240.244
R12654 gnd.n6380 gnd.n2519 240.244
R12655 gnd.n6380 gnd.n2535 240.244
R12656 gnd.n6376 gnd.n2535 240.244
R12657 gnd.n6376 gnd.n2540 240.244
R12658 gnd.n6368 gnd.n2540 240.244
R12659 gnd.n6368 gnd.n2555 240.244
R12660 gnd.n6364 gnd.n2555 240.244
R12661 gnd.n6364 gnd.n2560 240.244
R12662 gnd.n6356 gnd.n2560 240.244
R12663 gnd.n6689 gnd.n704 240.244
R12664 gnd.n6693 gnd.n704 240.244
R12665 gnd.n6693 gnd.n700 240.244
R12666 gnd.n6699 gnd.n700 240.244
R12667 gnd.n6699 gnd.n698 240.244
R12668 gnd.n6703 gnd.n698 240.244
R12669 gnd.n6703 gnd.n694 240.244
R12670 gnd.n6709 gnd.n694 240.244
R12671 gnd.n6709 gnd.n692 240.244
R12672 gnd.n6713 gnd.n692 240.244
R12673 gnd.n6713 gnd.n688 240.244
R12674 gnd.n6719 gnd.n688 240.244
R12675 gnd.n6719 gnd.n686 240.244
R12676 gnd.n6723 gnd.n686 240.244
R12677 gnd.n6723 gnd.n682 240.244
R12678 gnd.n6729 gnd.n682 240.244
R12679 gnd.n6729 gnd.n680 240.244
R12680 gnd.n6733 gnd.n680 240.244
R12681 gnd.n6733 gnd.n676 240.244
R12682 gnd.n6739 gnd.n676 240.244
R12683 gnd.n6739 gnd.n674 240.244
R12684 gnd.n6743 gnd.n674 240.244
R12685 gnd.n6743 gnd.n670 240.244
R12686 gnd.n6749 gnd.n670 240.244
R12687 gnd.n6749 gnd.n668 240.244
R12688 gnd.n6753 gnd.n668 240.244
R12689 gnd.n6753 gnd.n664 240.244
R12690 gnd.n6759 gnd.n664 240.244
R12691 gnd.n6759 gnd.n662 240.244
R12692 gnd.n6763 gnd.n662 240.244
R12693 gnd.n6763 gnd.n658 240.244
R12694 gnd.n6769 gnd.n658 240.244
R12695 gnd.n6769 gnd.n656 240.244
R12696 gnd.n6773 gnd.n656 240.244
R12697 gnd.n6773 gnd.n652 240.244
R12698 gnd.n6779 gnd.n652 240.244
R12699 gnd.n6779 gnd.n650 240.244
R12700 gnd.n6783 gnd.n650 240.244
R12701 gnd.n6783 gnd.n646 240.244
R12702 gnd.n6789 gnd.n646 240.244
R12703 gnd.n6789 gnd.n644 240.244
R12704 gnd.n6793 gnd.n644 240.244
R12705 gnd.n6793 gnd.n640 240.244
R12706 gnd.n6799 gnd.n640 240.244
R12707 gnd.n6799 gnd.n638 240.244
R12708 gnd.n6803 gnd.n638 240.244
R12709 gnd.n6803 gnd.n634 240.244
R12710 gnd.n6809 gnd.n634 240.244
R12711 gnd.n6809 gnd.n632 240.244
R12712 gnd.n6813 gnd.n632 240.244
R12713 gnd.n6813 gnd.n628 240.244
R12714 gnd.n6819 gnd.n628 240.244
R12715 gnd.n6819 gnd.n626 240.244
R12716 gnd.n6823 gnd.n626 240.244
R12717 gnd.n6823 gnd.n622 240.244
R12718 gnd.n6829 gnd.n622 240.244
R12719 gnd.n6829 gnd.n620 240.244
R12720 gnd.n6833 gnd.n620 240.244
R12721 gnd.n6833 gnd.n616 240.244
R12722 gnd.n6839 gnd.n616 240.244
R12723 gnd.n6839 gnd.n614 240.244
R12724 gnd.n6843 gnd.n614 240.244
R12725 gnd.n6843 gnd.n610 240.244
R12726 gnd.n6849 gnd.n610 240.244
R12727 gnd.n6849 gnd.n608 240.244
R12728 gnd.n6853 gnd.n608 240.244
R12729 gnd.n6853 gnd.n604 240.244
R12730 gnd.n6859 gnd.n604 240.244
R12731 gnd.n6859 gnd.n602 240.244
R12732 gnd.n6863 gnd.n602 240.244
R12733 gnd.n6863 gnd.n598 240.244
R12734 gnd.n6869 gnd.n598 240.244
R12735 gnd.n6869 gnd.n596 240.244
R12736 gnd.n6873 gnd.n596 240.244
R12737 gnd.n6873 gnd.n592 240.244
R12738 gnd.n6879 gnd.n592 240.244
R12739 gnd.n6879 gnd.n590 240.244
R12740 gnd.n6883 gnd.n590 240.244
R12741 gnd.n6883 gnd.n586 240.244
R12742 gnd.n6889 gnd.n586 240.244
R12743 gnd.n6889 gnd.n584 240.244
R12744 gnd.n6893 gnd.n584 240.244
R12745 gnd.n6893 gnd.n580 240.244
R12746 gnd.n6899 gnd.n580 240.244
R12747 gnd.n6899 gnd.n578 240.244
R12748 gnd.n6903 gnd.n578 240.244
R12749 gnd.n6903 gnd.n574 240.244
R12750 gnd.n6909 gnd.n574 240.244
R12751 gnd.n6909 gnd.n572 240.244
R12752 gnd.n6913 gnd.n572 240.244
R12753 gnd.n6913 gnd.n568 240.244
R12754 gnd.n6919 gnd.n568 240.244
R12755 gnd.n6919 gnd.n566 240.244
R12756 gnd.n6923 gnd.n566 240.244
R12757 gnd.n6923 gnd.n562 240.244
R12758 gnd.n6929 gnd.n562 240.244
R12759 gnd.n6929 gnd.n560 240.244
R12760 gnd.n6933 gnd.n560 240.244
R12761 gnd.n6933 gnd.n556 240.244
R12762 gnd.n6939 gnd.n556 240.244
R12763 gnd.n6939 gnd.n554 240.244
R12764 gnd.n6943 gnd.n554 240.244
R12765 gnd.n6943 gnd.n550 240.244
R12766 gnd.n6949 gnd.n550 240.244
R12767 gnd.n6949 gnd.n548 240.244
R12768 gnd.n6953 gnd.n548 240.244
R12769 gnd.n6953 gnd.n544 240.244
R12770 gnd.n6959 gnd.n544 240.244
R12771 gnd.n6959 gnd.n542 240.244
R12772 gnd.n6963 gnd.n542 240.244
R12773 gnd.n6963 gnd.n538 240.244
R12774 gnd.n6969 gnd.n538 240.244
R12775 gnd.n6969 gnd.n536 240.244
R12776 gnd.n6973 gnd.n536 240.244
R12777 gnd.n6973 gnd.n532 240.244
R12778 gnd.n6979 gnd.n532 240.244
R12779 gnd.n6979 gnd.n530 240.244
R12780 gnd.n6983 gnd.n530 240.244
R12781 gnd.n6983 gnd.n526 240.244
R12782 gnd.n6989 gnd.n526 240.244
R12783 gnd.n6989 gnd.n524 240.244
R12784 gnd.n6993 gnd.n524 240.244
R12785 gnd.n6993 gnd.n520 240.244
R12786 gnd.n6999 gnd.n520 240.244
R12787 gnd.n6999 gnd.n518 240.244
R12788 gnd.n7003 gnd.n518 240.244
R12789 gnd.n7003 gnd.n514 240.244
R12790 gnd.n7009 gnd.n514 240.244
R12791 gnd.n7009 gnd.n512 240.244
R12792 gnd.n7013 gnd.n512 240.244
R12793 gnd.n7013 gnd.n508 240.244
R12794 gnd.n7019 gnd.n508 240.244
R12795 gnd.n7019 gnd.n506 240.244
R12796 gnd.n7023 gnd.n506 240.244
R12797 gnd.n7023 gnd.n502 240.244
R12798 gnd.n7029 gnd.n502 240.244
R12799 gnd.n7029 gnd.n500 240.244
R12800 gnd.n7033 gnd.n500 240.244
R12801 gnd.n7033 gnd.n496 240.244
R12802 gnd.n7039 gnd.n496 240.244
R12803 gnd.n7039 gnd.n494 240.244
R12804 gnd.n7043 gnd.n494 240.244
R12805 gnd.n7043 gnd.n490 240.244
R12806 gnd.n7049 gnd.n490 240.244
R12807 gnd.n7049 gnd.n488 240.244
R12808 gnd.n7053 gnd.n488 240.244
R12809 gnd.n7053 gnd.n484 240.244
R12810 gnd.n7059 gnd.n484 240.244
R12811 gnd.n7059 gnd.n482 240.244
R12812 gnd.n7063 gnd.n482 240.244
R12813 gnd.n7063 gnd.n478 240.244
R12814 gnd.n7069 gnd.n478 240.244
R12815 gnd.n7069 gnd.n476 240.244
R12816 gnd.n7073 gnd.n476 240.244
R12817 gnd.n7073 gnd.n472 240.244
R12818 gnd.n7079 gnd.n472 240.244
R12819 gnd.n7079 gnd.n470 240.244
R12820 gnd.n7083 gnd.n470 240.244
R12821 gnd.n7083 gnd.n466 240.244
R12822 gnd.n7089 gnd.n466 240.244
R12823 gnd.n7089 gnd.n464 240.244
R12824 gnd.n7093 gnd.n464 240.244
R12825 gnd.n7093 gnd.n460 240.244
R12826 gnd.n7099 gnd.n460 240.244
R12827 gnd.n7099 gnd.n458 240.244
R12828 gnd.n7103 gnd.n458 240.244
R12829 gnd.n7103 gnd.n454 240.244
R12830 gnd.n7109 gnd.n454 240.244
R12831 gnd.n7109 gnd.n452 240.244
R12832 gnd.n7113 gnd.n452 240.244
R12833 gnd.n7113 gnd.n448 240.244
R12834 gnd.n7119 gnd.n448 240.244
R12835 gnd.n7119 gnd.n446 240.244
R12836 gnd.n7123 gnd.n446 240.244
R12837 gnd.n7123 gnd.n442 240.244
R12838 gnd.n7129 gnd.n442 240.244
R12839 gnd.n7129 gnd.n440 240.244
R12840 gnd.n7133 gnd.n440 240.244
R12841 gnd.n7133 gnd.n436 240.244
R12842 gnd.n7139 gnd.n436 240.244
R12843 gnd.n7139 gnd.n434 240.244
R12844 gnd.n7143 gnd.n434 240.244
R12845 gnd.n7143 gnd.n430 240.244
R12846 gnd.n7149 gnd.n430 240.244
R12847 gnd.n7149 gnd.n428 240.244
R12848 gnd.n7153 gnd.n428 240.244
R12849 gnd.n7153 gnd.n424 240.244
R12850 gnd.n7159 gnd.n424 240.244
R12851 gnd.n7159 gnd.n422 240.244
R12852 gnd.n7163 gnd.n422 240.244
R12853 gnd.n7163 gnd.n418 240.244
R12854 gnd.n7169 gnd.n418 240.244
R12855 gnd.n7169 gnd.n416 240.244
R12856 gnd.n7173 gnd.n416 240.244
R12857 gnd.n7173 gnd.n412 240.244
R12858 gnd.n7179 gnd.n412 240.244
R12859 gnd.n7179 gnd.n410 240.244
R12860 gnd.n7183 gnd.n410 240.244
R12861 gnd.n7183 gnd.n406 240.244
R12862 gnd.n7189 gnd.n406 240.244
R12863 gnd.n7189 gnd.n404 240.244
R12864 gnd.n7193 gnd.n404 240.244
R12865 gnd.n7193 gnd.n400 240.244
R12866 gnd.n7200 gnd.n400 240.244
R12867 gnd.n7200 gnd.n398 240.244
R12868 gnd.n7204 gnd.n398 240.244
R12869 gnd.n7204 gnd.n395 240.244
R12870 gnd.n7210 gnd.n393 240.244
R12871 gnd.n7214 gnd.n393 240.244
R12872 gnd.n7214 gnd.n389 240.244
R12873 gnd.n7220 gnd.n389 240.244
R12874 gnd.n7220 gnd.n387 240.244
R12875 gnd.n7224 gnd.n387 240.244
R12876 gnd.n7224 gnd.n383 240.244
R12877 gnd.n7230 gnd.n383 240.244
R12878 gnd.n7230 gnd.n381 240.244
R12879 gnd.n7234 gnd.n381 240.244
R12880 gnd.n7234 gnd.n377 240.244
R12881 gnd.n7240 gnd.n377 240.244
R12882 gnd.n7240 gnd.n375 240.244
R12883 gnd.n7244 gnd.n375 240.244
R12884 gnd.n7244 gnd.n371 240.244
R12885 gnd.n7250 gnd.n371 240.244
R12886 gnd.n7250 gnd.n369 240.244
R12887 gnd.n7254 gnd.n369 240.244
R12888 gnd.n7254 gnd.n365 240.244
R12889 gnd.n7260 gnd.n365 240.244
R12890 gnd.n7260 gnd.n363 240.244
R12891 gnd.n7264 gnd.n363 240.244
R12892 gnd.n7264 gnd.n359 240.244
R12893 gnd.n7270 gnd.n359 240.244
R12894 gnd.n7270 gnd.n357 240.244
R12895 gnd.n7274 gnd.n357 240.244
R12896 gnd.n7274 gnd.n353 240.244
R12897 gnd.n7280 gnd.n353 240.244
R12898 gnd.n7280 gnd.n351 240.244
R12899 gnd.n7284 gnd.n351 240.244
R12900 gnd.n7284 gnd.n347 240.244
R12901 gnd.n7290 gnd.n347 240.244
R12902 gnd.n7290 gnd.n345 240.244
R12903 gnd.n7294 gnd.n345 240.244
R12904 gnd.n7294 gnd.n341 240.244
R12905 gnd.n7300 gnd.n341 240.244
R12906 gnd.n7300 gnd.n339 240.244
R12907 gnd.n7304 gnd.n339 240.244
R12908 gnd.n7304 gnd.n335 240.244
R12909 gnd.n7310 gnd.n335 240.244
R12910 gnd.n7310 gnd.n333 240.244
R12911 gnd.n7314 gnd.n333 240.244
R12912 gnd.n7314 gnd.n329 240.244
R12913 gnd.n7320 gnd.n329 240.244
R12914 gnd.n7320 gnd.n327 240.244
R12915 gnd.n7324 gnd.n327 240.244
R12916 gnd.n7324 gnd.n323 240.244
R12917 gnd.n7330 gnd.n323 240.244
R12918 gnd.n7330 gnd.n321 240.244
R12919 gnd.n7334 gnd.n321 240.244
R12920 gnd.n7334 gnd.n317 240.244
R12921 gnd.n7340 gnd.n317 240.244
R12922 gnd.n7340 gnd.n315 240.244
R12923 gnd.n7344 gnd.n315 240.244
R12924 gnd.n7344 gnd.n311 240.244
R12925 gnd.n7350 gnd.n311 240.244
R12926 gnd.n7350 gnd.n309 240.244
R12927 gnd.n7354 gnd.n309 240.244
R12928 gnd.n7354 gnd.n305 240.244
R12929 gnd.n7360 gnd.n305 240.244
R12930 gnd.n7360 gnd.n303 240.244
R12931 gnd.n7364 gnd.n303 240.244
R12932 gnd.n7364 gnd.n299 240.244
R12933 gnd.n7370 gnd.n299 240.244
R12934 gnd.n7370 gnd.n297 240.244
R12935 gnd.n7374 gnd.n297 240.244
R12936 gnd.n7374 gnd.n293 240.244
R12937 gnd.n7380 gnd.n293 240.244
R12938 gnd.n7380 gnd.n291 240.244
R12939 gnd.n7384 gnd.n291 240.244
R12940 gnd.n7384 gnd.n287 240.244
R12941 gnd.n7390 gnd.n287 240.244
R12942 gnd.n7390 gnd.n285 240.244
R12943 gnd.n7394 gnd.n285 240.244
R12944 gnd.n7394 gnd.n281 240.244
R12945 gnd.n7400 gnd.n281 240.244
R12946 gnd.n7400 gnd.n279 240.244
R12947 gnd.n7404 gnd.n279 240.244
R12948 gnd.n7404 gnd.n275 240.244
R12949 gnd.n7410 gnd.n275 240.244
R12950 gnd.n7410 gnd.n273 240.244
R12951 gnd.n7414 gnd.n273 240.244
R12952 gnd.n7414 gnd.n269 240.244
R12953 gnd.n7421 gnd.n269 240.244
R12954 gnd.n6513 gnd.n876 240.244
R12955 gnd.n6509 gnd.n876 240.244
R12956 gnd.n6509 gnd.n2341 240.244
R12957 gnd.n6505 gnd.n2341 240.244
R12958 gnd.n6505 gnd.n2346 240.244
R12959 gnd.n6501 gnd.n2346 240.244
R12960 gnd.n6501 gnd.n2348 240.244
R12961 gnd.n6497 gnd.n2348 240.244
R12962 gnd.n6497 gnd.n2354 240.244
R12963 gnd.n6493 gnd.n2354 240.244
R12964 gnd.n6493 gnd.n2356 240.244
R12965 gnd.n6489 gnd.n2356 240.244
R12966 gnd.n6489 gnd.n2362 240.244
R12967 gnd.n3923 gnd.n2362 240.244
R12968 gnd.n4258 gnd.n3923 240.244
R12969 gnd.n4258 gnd.n3918 240.244
R12970 gnd.n4264 gnd.n3918 240.244
R12971 gnd.n4265 gnd.n4264 240.244
R12972 gnd.n4266 gnd.n4265 240.244
R12973 gnd.n4266 gnd.n3914 240.244
R12974 gnd.n4272 gnd.n3914 240.244
R12975 gnd.n4273 gnd.n4272 240.244
R12976 gnd.n4274 gnd.n4273 240.244
R12977 gnd.n4274 gnd.n3909 240.244
R12978 gnd.n4285 gnd.n3909 240.244
R12979 gnd.n4285 gnd.n3910 240.244
R12980 gnd.n4281 gnd.n3910 240.244
R12981 gnd.n4281 gnd.n3886 240.244
R12982 gnd.n4362 gnd.n3886 240.244
R12983 gnd.n4362 gnd.n4361 240.244
R12984 gnd.n4361 gnd.n4360 240.244
R12985 gnd.n4360 gnd.n4357 240.244
R12986 gnd.n4357 gnd.n4356 240.244
R12987 gnd.n4356 gnd.n3887 240.244
R12988 gnd.n4321 gnd.n3887 240.244
R12989 gnd.n4330 gnd.n4321 240.244
R12990 gnd.n4330 gnd.n4327 240.244
R12991 gnd.n4327 gnd.n4324 240.244
R12992 gnd.n4324 gnd.n4323 240.244
R12993 gnd.n4323 gnd.n3875 240.244
R12994 gnd.n4388 gnd.n3875 240.244
R12995 gnd.n4388 gnd.n3876 240.244
R12996 gnd.n4384 gnd.n3876 240.244
R12997 gnd.n4384 gnd.n4383 240.244
R12998 gnd.n4383 gnd.n4382 240.244
R12999 gnd.n4382 gnd.n4371 240.244
R13000 gnd.n4378 gnd.n4371 240.244
R13001 gnd.n4378 gnd.n3856 240.244
R13002 gnd.n4438 gnd.n3856 240.244
R13003 gnd.n4439 gnd.n4438 240.244
R13004 gnd.n4439 gnd.n3852 240.244
R13005 gnd.n4445 gnd.n3852 240.244
R13006 gnd.n4446 gnd.n4445 240.244
R13007 gnd.n4447 gnd.n4446 240.244
R13008 gnd.n4447 gnd.n3848 240.244
R13009 gnd.n4453 gnd.n3848 240.244
R13010 gnd.n4454 gnd.n4453 240.244
R13011 gnd.n4455 gnd.n4454 240.244
R13012 gnd.n4455 gnd.n3844 240.244
R13013 gnd.n4461 gnd.n3844 240.244
R13014 gnd.n4462 gnd.n4461 240.244
R13015 gnd.n4465 gnd.n4462 240.244
R13016 gnd.n4465 gnd.n3838 240.244
R13017 gnd.n4474 gnd.n3838 240.244
R13018 gnd.n4474 gnd.n3839 240.244
R13019 gnd.n3839 gnd.n2914 240.244
R13020 gnd.n6148 gnd.n2914 240.244
R13021 gnd.n6148 gnd.n2915 240.244
R13022 gnd.n6144 gnd.n2915 240.244
R13023 gnd.n6144 gnd.n2921 240.244
R13024 gnd.n6134 gnd.n2921 240.244
R13025 gnd.n6134 gnd.n2933 240.244
R13026 gnd.n6130 gnd.n2933 240.244
R13027 gnd.n6130 gnd.n2939 240.244
R13028 gnd.n4559 gnd.n2939 240.244
R13029 gnd.n4559 gnd.n3712 240.244
R13030 gnd.n4589 gnd.n3712 240.244
R13031 gnd.n4589 gnd.n3708 240.244
R13032 gnd.n4595 gnd.n3708 240.244
R13033 gnd.n4595 gnd.n3687 240.244
R13034 gnd.n4632 gnd.n3687 240.244
R13035 gnd.n4632 gnd.n3683 240.244
R13036 gnd.n4638 gnd.n3683 240.244
R13037 gnd.n4638 gnd.n3672 240.244
R13038 gnd.n4677 gnd.n3672 240.244
R13039 gnd.n4677 gnd.n3667 240.244
R13040 gnd.n4685 gnd.n3667 240.244
R13041 gnd.n4685 gnd.n3668 240.244
R13042 gnd.n3668 gnd.n3644 240.244
R13043 gnd.n4750 gnd.n3644 240.244
R13044 gnd.n4750 gnd.n3640 240.244
R13045 gnd.n4756 gnd.n3640 240.244
R13046 gnd.n4756 gnd.n3624 240.244
R13047 gnd.n4778 gnd.n3624 240.244
R13048 gnd.n4778 gnd.n3620 240.244
R13049 gnd.n4784 gnd.n3620 240.244
R13050 gnd.n4784 gnd.n3603 240.244
R13051 gnd.n4811 gnd.n3603 240.244
R13052 gnd.n4811 gnd.n3599 240.244
R13053 gnd.n4817 gnd.n3599 240.244
R13054 gnd.n4817 gnd.n3586 240.244
R13055 gnd.n4855 gnd.n3586 240.244
R13056 gnd.n4855 gnd.n3581 240.244
R13057 gnd.n4863 gnd.n3581 240.244
R13058 gnd.n4863 gnd.n3582 240.244
R13059 gnd.n3582 gnd.n3557 240.244
R13060 gnd.n4905 gnd.n3557 240.244
R13061 gnd.n4905 gnd.n3553 240.244
R13062 gnd.n4911 gnd.n3553 240.244
R13063 gnd.n4911 gnd.n3538 240.244
R13064 gnd.n4933 gnd.n3538 240.244
R13065 gnd.n4933 gnd.n3533 240.244
R13066 gnd.n4948 gnd.n3533 240.244
R13067 gnd.n4948 gnd.n3534 240.244
R13068 gnd.n4944 gnd.n3534 240.244
R13069 gnd.n4944 gnd.n3507 240.244
R13070 gnd.n5008 gnd.n3507 240.244
R13071 gnd.n5008 gnd.n3502 240.244
R13072 gnd.n5016 gnd.n3502 240.244
R13073 gnd.n5016 gnd.n3503 240.244
R13074 gnd.n3503 gnd.n3479 240.244
R13075 gnd.n5060 gnd.n3479 240.244
R13076 gnd.n5060 gnd.n3475 240.244
R13077 gnd.n5068 gnd.n3475 240.244
R13078 gnd.n5068 gnd.n3462 240.244
R13079 gnd.n5087 gnd.n3462 240.244
R13080 gnd.n5088 gnd.n5087 240.244
R13081 gnd.n5088 gnd.n3458 240.244
R13082 gnd.n5094 gnd.n3458 240.244
R13083 gnd.n5094 gnd.n3404 240.244
R13084 gnd.n5131 gnd.n3404 240.244
R13085 gnd.n5131 gnd.n3400 240.244
R13086 gnd.n5137 gnd.n3400 240.244
R13087 gnd.n5137 gnd.n3382 240.244
R13088 gnd.n5159 gnd.n3382 240.244
R13089 gnd.n5159 gnd.n3377 240.244
R13090 gnd.n5168 gnd.n3377 240.244
R13091 gnd.n5168 gnd.n3378 240.244
R13092 gnd.n3378 gnd.n3348 240.244
R13093 gnd.n5383 gnd.n3348 240.244
R13094 gnd.n5383 gnd.n3349 240.244
R13095 gnd.n5379 gnd.n3349 240.244
R13096 gnd.n5379 gnd.n5378 240.244
R13097 gnd.n5378 gnd.n3039 240.244
R13098 gnd.n6015 gnd.n3039 240.244
R13099 gnd.n6015 gnd.n3040 240.244
R13100 gnd.n6011 gnd.n3040 240.244
R13101 gnd.n6011 gnd.n3046 240.244
R13102 gnd.n6007 gnd.n3046 240.244
R13103 gnd.n6007 gnd.n3049 240.244
R13104 gnd.n6003 gnd.n3049 240.244
R13105 gnd.n6003 gnd.n3055 240.244
R13106 gnd.n5767 gnd.n3055 240.244
R13107 gnd.n5767 gnd.n5764 240.244
R13108 gnd.n5773 gnd.n5764 240.244
R13109 gnd.n5774 gnd.n5773 240.244
R13110 gnd.n5775 gnd.n5774 240.244
R13111 gnd.n5775 gnd.n5760 240.244
R13112 gnd.n5781 gnd.n5760 240.244
R13113 gnd.n5782 gnd.n5781 240.244
R13114 gnd.n5783 gnd.n5782 240.244
R13115 gnd.n5783 gnd.n3248 240.244
R13116 gnd.n5801 gnd.n3248 240.244
R13117 gnd.n5801 gnd.n3249 240.244
R13118 gnd.n5797 gnd.n3249 240.244
R13119 gnd.n5797 gnd.n5796 240.244
R13120 gnd.n5796 gnd.n5795 240.244
R13121 gnd.n5795 gnd.n3150 240.244
R13122 gnd.n5947 gnd.n3150 240.244
R13123 gnd.n5947 gnd.n3151 240.244
R13124 gnd.n5942 gnd.n3151 240.244
R13125 gnd.n5942 gnd.n3154 240.244
R13126 gnd.n3178 gnd.n3154 240.244
R13127 gnd.n3179 gnd.n3178 240.244
R13128 gnd.n3179 gnd.n3174 240.244
R13129 gnd.n5926 gnd.n3174 240.244
R13130 gnd.n5926 gnd.n3175 240.244
R13131 gnd.n5921 gnd.n3175 240.244
R13132 gnd.n5921 gnd.n5920 240.244
R13133 gnd.n5920 gnd.n5919 240.244
R13134 gnd.n5919 gnd.n3185 240.244
R13135 gnd.n5915 gnd.n3185 240.244
R13136 gnd.n5915 gnd.n3226 240.244
R13137 gnd.n3226 gnd.n3225 240.244
R13138 gnd.n3225 gnd.n3191 240.244
R13139 gnd.n3221 gnd.n3191 240.244
R13140 gnd.n3221 gnd.n3220 240.244
R13141 gnd.n3220 gnd.n3219 240.244
R13142 gnd.n3219 gnd.n3197 240.244
R13143 gnd.n3215 gnd.n3197 240.244
R13144 gnd.n3215 gnd.n3214 240.244
R13145 gnd.n3214 gnd.n3213 240.244
R13146 gnd.n3213 gnd.n3203 240.244
R13147 gnd.n3209 gnd.n3203 240.244
R13148 gnd.n3209 gnd.n244 240.244
R13149 gnd.n7445 gnd.n244 240.244
R13150 gnd.n7445 gnd.n245 240.244
R13151 gnd.n7441 gnd.n245 240.244
R13152 gnd.n7441 gnd.n251 240.244
R13153 gnd.n7437 gnd.n251 240.244
R13154 gnd.n7437 gnd.n253 240.244
R13155 gnd.n7433 gnd.n253 240.244
R13156 gnd.n7433 gnd.n259 240.244
R13157 gnd.n7429 gnd.n259 240.244
R13158 gnd.n7429 gnd.n261 240.244
R13159 gnd.n7425 gnd.n261 240.244
R13160 gnd.n7425 gnd.n267 240.244
R13161 gnd.n6683 gnd.n706 240.244
R13162 gnd.n6683 gnd.n709 240.244
R13163 gnd.n6679 gnd.n709 240.244
R13164 gnd.n6679 gnd.n711 240.244
R13165 gnd.n6675 gnd.n711 240.244
R13166 gnd.n6675 gnd.n717 240.244
R13167 gnd.n6671 gnd.n717 240.244
R13168 gnd.n6671 gnd.n719 240.244
R13169 gnd.n6667 gnd.n719 240.244
R13170 gnd.n6667 gnd.n725 240.244
R13171 gnd.n6663 gnd.n725 240.244
R13172 gnd.n6663 gnd.n727 240.244
R13173 gnd.n6659 gnd.n727 240.244
R13174 gnd.n6659 gnd.n733 240.244
R13175 gnd.n6655 gnd.n733 240.244
R13176 gnd.n6655 gnd.n735 240.244
R13177 gnd.n6651 gnd.n735 240.244
R13178 gnd.n6651 gnd.n741 240.244
R13179 gnd.n6647 gnd.n741 240.244
R13180 gnd.n6647 gnd.n743 240.244
R13181 gnd.n6643 gnd.n743 240.244
R13182 gnd.n6643 gnd.n749 240.244
R13183 gnd.n6639 gnd.n749 240.244
R13184 gnd.n6639 gnd.n751 240.244
R13185 gnd.n6635 gnd.n751 240.244
R13186 gnd.n6635 gnd.n757 240.244
R13187 gnd.n6631 gnd.n757 240.244
R13188 gnd.n6631 gnd.n759 240.244
R13189 gnd.n6627 gnd.n759 240.244
R13190 gnd.n6627 gnd.n765 240.244
R13191 gnd.n6623 gnd.n765 240.244
R13192 gnd.n6623 gnd.n767 240.244
R13193 gnd.n6619 gnd.n767 240.244
R13194 gnd.n6619 gnd.n773 240.244
R13195 gnd.n6615 gnd.n773 240.244
R13196 gnd.n6615 gnd.n775 240.244
R13197 gnd.n6611 gnd.n775 240.244
R13198 gnd.n6611 gnd.n781 240.244
R13199 gnd.n6607 gnd.n781 240.244
R13200 gnd.n6607 gnd.n783 240.244
R13201 gnd.n6603 gnd.n783 240.244
R13202 gnd.n6603 gnd.n789 240.244
R13203 gnd.n6599 gnd.n789 240.244
R13204 gnd.n6599 gnd.n791 240.244
R13205 gnd.n6595 gnd.n791 240.244
R13206 gnd.n6595 gnd.n797 240.244
R13207 gnd.n6591 gnd.n797 240.244
R13208 gnd.n6591 gnd.n799 240.244
R13209 gnd.n6587 gnd.n799 240.244
R13210 gnd.n6587 gnd.n805 240.244
R13211 gnd.n6583 gnd.n805 240.244
R13212 gnd.n6583 gnd.n807 240.244
R13213 gnd.n6579 gnd.n807 240.244
R13214 gnd.n6579 gnd.n813 240.244
R13215 gnd.n6575 gnd.n813 240.244
R13216 gnd.n6575 gnd.n815 240.244
R13217 gnd.n6571 gnd.n815 240.244
R13218 gnd.n6571 gnd.n821 240.244
R13219 gnd.n6567 gnd.n821 240.244
R13220 gnd.n6567 gnd.n823 240.244
R13221 gnd.n6563 gnd.n823 240.244
R13222 gnd.n6563 gnd.n829 240.244
R13223 gnd.n6559 gnd.n829 240.244
R13224 gnd.n6559 gnd.n831 240.244
R13225 gnd.n6555 gnd.n831 240.244
R13226 gnd.n6555 gnd.n837 240.244
R13227 gnd.n6551 gnd.n837 240.244
R13228 gnd.n6551 gnd.n839 240.244
R13229 gnd.n6547 gnd.n839 240.244
R13230 gnd.n6547 gnd.n845 240.244
R13231 gnd.n6543 gnd.n845 240.244
R13232 gnd.n6543 gnd.n847 240.244
R13233 gnd.n6539 gnd.n847 240.244
R13234 gnd.n6539 gnd.n853 240.244
R13235 gnd.n6535 gnd.n853 240.244
R13236 gnd.n6535 gnd.n855 240.244
R13237 gnd.n6531 gnd.n855 240.244
R13238 gnd.n6531 gnd.n861 240.244
R13239 gnd.n6527 gnd.n861 240.244
R13240 gnd.n6527 gnd.n863 240.244
R13241 gnd.n6523 gnd.n863 240.244
R13242 gnd.n6523 gnd.n869 240.244
R13243 gnd.n6519 gnd.n869 240.244
R13244 gnd.n6519 gnd.n871 240.244
R13245 gnd.n4477 gnd.n2604 240.244
R13246 gnd.n4477 gnd.n3826 240.244
R13247 gnd.n4484 gnd.n3826 240.244
R13248 gnd.n4484 gnd.n3827 240.244
R13249 gnd.n3827 gnd.n3744 240.244
R13250 gnd.n4509 gnd.n3744 240.244
R13251 gnd.n4509 gnd.n2925 240.244
R13252 gnd.n4516 gnd.n2925 240.244
R13253 gnd.n4516 gnd.n3739 240.244
R13254 gnd.n3739 gnd.n2943 240.244
R13255 gnd.n6127 gnd.n2943 240.244
R13256 gnd.n6127 gnd.n2944 240.244
R13257 gnd.n2949 gnd.n2944 240.244
R13258 gnd.n2950 gnd.n2949 240.244
R13259 gnd.n2951 gnd.n2950 240.244
R13260 gnd.n4597 gnd.n2951 240.244
R13261 gnd.n4597 gnd.n2954 240.244
R13262 gnd.n2955 gnd.n2954 240.244
R13263 gnd.n2956 gnd.n2955 240.244
R13264 gnd.n4622 gnd.n2956 240.244
R13265 gnd.n4622 gnd.n2959 240.244
R13266 gnd.n2960 gnd.n2959 240.244
R13267 gnd.n2961 gnd.n2960 240.244
R13268 gnd.n4687 gnd.n2961 240.244
R13269 gnd.n4687 gnd.n2964 240.244
R13270 gnd.n2965 gnd.n2964 240.244
R13271 gnd.n2966 gnd.n2965 240.244
R13272 gnd.n4747 gnd.n2966 240.244
R13273 gnd.n4747 gnd.n2969 240.244
R13274 gnd.n2970 gnd.n2969 240.244
R13275 gnd.n2971 gnd.n2970 240.244
R13276 gnd.n4775 gnd.n2971 240.244
R13277 gnd.n4775 gnd.n2974 240.244
R13278 gnd.n2975 gnd.n2974 240.244
R13279 gnd.n2976 gnd.n2975 240.244
R13280 gnd.n3606 gnd.n2976 240.244
R13281 gnd.n3606 gnd.n2979 240.244
R13282 gnd.n2980 gnd.n2979 240.244
R13283 gnd.n2981 gnd.n2980 240.244
R13284 gnd.n3589 gnd.n2981 240.244
R13285 gnd.n3589 gnd.n2984 240.244
R13286 gnd.n2985 gnd.n2984 240.244
R13287 gnd.n2986 gnd.n2985 240.244
R13288 gnd.n4894 gnd.n2986 240.244
R13289 gnd.n4894 gnd.n2989 240.244
R13290 gnd.n2990 gnd.n2989 240.244
R13291 gnd.n2991 gnd.n2990 240.244
R13292 gnd.n4880 gnd.n2991 240.244
R13293 gnd.n4880 gnd.n2994 240.244
R13294 gnd.n2995 gnd.n2994 240.244
R13295 gnd.n2996 gnd.n2995 240.244
R13296 gnd.n4941 gnd.n2996 240.244
R13297 gnd.n4941 gnd.n2999 240.244
R13298 gnd.n3000 gnd.n2999 240.244
R13299 gnd.n3001 gnd.n3000 240.244
R13300 gnd.n5018 gnd.n3001 240.244
R13301 gnd.n5018 gnd.n3004 240.244
R13302 gnd.n3005 gnd.n3004 240.244
R13303 gnd.n3006 gnd.n3005 240.244
R13304 gnd.n5057 gnd.n3006 240.244
R13305 gnd.n5057 gnd.n3009 240.244
R13306 gnd.n3010 gnd.n3009 240.244
R13307 gnd.n3011 gnd.n3010 240.244
R13308 gnd.n5084 gnd.n3011 240.244
R13309 gnd.n5084 gnd.n3014 240.244
R13310 gnd.n3015 gnd.n3014 240.244
R13311 gnd.n3016 gnd.n3015 240.244
R13312 gnd.n5121 gnd.n3016 240.244
R13313 gnd.n5121 gnd.n3019 240.244
R13314 gnd.n3020 gnd.n3019 240.244
R13315 gnd.n3021 gnd.n3020 240.244
R13316 gnd.n3392 gnd.n3021 240.244
R13317 gnd.n3392 gnd.n3024 240.244
R13318 gnd.n3025 gnd.n3024 240.244
R13319 gnd.n3026 gnd.n3025 240.244
R13320 gnd.n3435 gnd.n3026 240.244
R13321 gnd.n3435 gnd.n3029 240.244
R13322 gnd.n3030 gnd.n3029 240.244
R13323 gnd.n3031 gnd.n3030 240.244
R13324 gnd.n3357 gnd.n3031 240.244
R13325 gnd.n3357 gnd.n3034 240.244
R13326 gnd.n6018 gnd.n3034 240.244
R13327 gnd.n2603 gnd.n2602 240.244
R13328 gnd.n2608 gnd.n2602 240.244
R13329 gnd.n2610 gnd.n2609 240.244
R13330 gnd.n2614 gnd.n2613 240.244
R13331 gnd.n2616 gnd.n2615 240.244
R13332 gnd.n2626 gnd.n2625 240.244
R13333 gnd.n2628 gnd.n2627 240.244
R13334 gnd.n2636 gnd.n2635 240.244
R13335 gnd.n2644 gnd.n2643 240.244
R13336 gnd.n2646 gnd.n2645 240.244
R13337 gnd.n2654 gnd.n2653 240.244
R13338 gnd.n2662 gnd.n2661 240.244
R13339 gnd.n2667 gnd.n2663 240.244
R13340 gnd.n2599 gnd.n2585 240.244
R13341 gnd.n3837 gnd.n2586 240.244
R13342 gnd.n3837 gnd.n3756 240.244
R13343 gnd.n4486 gnd.n3756 240.244
R13344 gnd.n4486 gnd.n3751 240.244
R13345 gnd.n4498 gnd.n3751 240.244
R13346 gnd.n4498 gnd.n3748 240.244
R13347 gnd.n3748 gnd.n2923 240.244
R13348 gnd.n3738 gnd.n2923 240.244
R13349 gnd.n3738 gnd.n3732 240.244
R13350 gnd.n4541 gnd.n3732 240.244
R13351 gnd.n4541 gnd.n2941 240.244
R13352 gnd.n3726 gnd.n2941 240.244
R13353 gnd.n4553 gnd.n3726 240.244
R13354 gnd.n4553 gnd.n3727 240.244
R13355 gnd.n3727 gnd.n3714 240.244
R13356 gnd.n3714 gnd.n3700 240.244
R13357 gnd.n4607 gnd.n3700 240.244
R13358 gnd.n4608 gnd.n4607 240.244
R13359 gnd.n4608 gnd.n3694 240.244
R13360 gnd.n4621 gnd.n3694 240.244
R13361 gnd.n4621 gnd.n3695 240.244
R13362 gnd.n4613 gnd.n3695 240.244
R13363 gnd.n4614 gnd.n4613 240.244
R13364 gnd.n4614 gnd.n3659 240.244
R13365 gnd.n4696 gnd.n3659 240.244
R13366 gnd.n4696 gnd.n3654 240.244
R13367 gnd.n4738 gnd.n3654 240.244
R13368 gnd.n4738 gnd.n3646 240.244
R13369 gnd.n4701 gnd.n3646 240.244
R13370 gnd.n4702 gnd.n4701 240.244
R13371 gnd.n4703 gnd.n4702 240.244
R13372 gnd.n4703 gnd.n3626 240.244
R13373 gnd.n3626 gnd.n3618 240.244
R13374 gnd.n4707 gnd.n3618 240.244
R13375 gnd.n4708 gnd.n4707 240.244
R13376 gnd.n4711 gnd.n4708 240.244
R13377 gnd.n4712 gnd.n4711 240.244
R13378 gnd.n4713 gnd.n4712 240.244
R13379 gnd.n4714 gnd.n4713 240.244
R13380 gnd.n4715 gnd.n4714 240.244
R13381 gnd.n4715 gnd.n3572 240.244
R13382 gnd.n4873 gnd.n3572 240.244
R13383 gnd.n4873 gnd.n3567 240.244
R13384 gnd.n4893 gnd.n3567 240.244
R13385 gnd.n4893 gnd.n3559 240.244
R13386 gnd.n4878 gnd.n3559 240.244
R13387 gnd.n4879 gnd.n4878 240.244
R13388 gnd.n4882 gnd.n4879 240.244
R13389 gnd.n4882 gnd.n3540 240.244
R13390 gnd.n3540 gnd.n3523 240.244
R13391 gnd.n4960 gnd.n3523 240.244
R13392 gnd.n4960 gnd.n3517 240.244
R13393 gnd.n4970 gnd.n3517 240.244
R13394 gnd.n4970 gnd.n3518 240.244
R13395 gnd.n4964 gnd.n3518 240.244
R13396 gnd.n4964 gnd.n3494 240.244
R13397 gnd.n5028 gnd.n3494 240.244
R13398 gnd.n5028 gnd.n3489 240.244
R13399 gnd.n5048 gnd.n3489 240.244
R13400 gnd.n5048 gnd.n3481 240.244
R13401 gnd.n5033 gnd.n3481 240.244
R13402 gnd.n5036 gnd.n5033 240.244
R13403 gnd.n5037 gnd.n5036 240.244
R13404 gnd.n5037 gnd.n3464 240.244
R13405 gnd.n3464 gnd.n3419 240.244
R13406 gnd.n5113 gnd.n3419 240.244
R13407 gnd.n5113 gnd.n3413 240.244
R13408 gnd.n5120 gnd.n3413 240.244
R13409 gnd.n5120 gnd.n3414 240.244
R13410 gnd.n3414 gnd.n3389 240.244
R13411 gnd.n5149 gnd.n3389 240.244
R13412 gnd.n5149 gnd.n3385 240.244
R13413 gnd.n5155 gnd.n3385 240.244
R13414 gnd.n5155 gnd.n3368 240.244
R13415 gnd.n5180 gnd.n3368 240.244
R13416 gnd.n5180 gnd.n3364 240.244
R13417 gnd.n5186 gnd.n3364 240.244
R13418 gnd.n5188 gnd.n5186 240.244
R13419 gnd.n5190 gnd.n5188 240.244
R13420 gnd.n5190 gnd.n3359 240.244
R13421 gnd.n5375 gnd.n3359 240.244
R13422 gnd.n5375 gnd.n3037 240.244
R13423 gnd.n5262 gnd.n5261 240.244
R13424 gnd.n5265 gnd.n5264 240.244
R13425 gnd.n5273 gnd.n5272 240.244
R13426 gnd.n5276 gnd.n5275 240.244
R13427 gnd.n5288 gnd.n5287 240.244
R13428 gnd.n5291 gnd.n5290 240.244
R13429 gnd.n5307 gnd.n5306 240.244
R13430 gnd.n5310 gnd.n5309 240.244
R13431 gnd.n5326 gnd.n5325 240.244
R13432 gnd.n5329 gnd.n5328 240.244
R13433 gnd.n5345 gnd.n5344 240.244
R13434 gnd.n5347 gnd.n5203 240.244
R13435 gnd.n5364 gnd.n5203 240.244
R13436 gnd.n5367 gnd.n5366 240.244
R13437 gnd.n2896 gnd.n2895 240.132
R13438 gnd.n5400 gnd.n5399 240.132
R13439 gnd.n6691 gnd.n6690 225.874
R13440 gnd.n6692 gnd.n6691 225.874
R13441 gnd.n6692 gnd.n699 225.874
R13442 gnd.n6700 gnd.n699 225.874
R13443 gnd.n6701 gnd.n6700 225.874
R13444 gnd.n6702 gnd.n6701 225.874
R13445 gnd.n6702 gnd.n693 225.874
R13446 gnd.n6710 gnd.n693 225.874
R13447 gnd.n6711 gnd.n6710 225.874
R13448 gnd.n6712 gnd.n6711 225.874
R13449 gnd.n6712 gnd.n687 225.874
R13450 gnd.n6720 gnd.n687 225.874
R13451 gnd.n6721 gnd.n6720 225.874
R13452 gnd.n6722 gnd.n6721 225.874
R13453 gnd.n6722 gnd.n681 225.874
R13454 gnd.n6730 gnd.n681 225.874
R13455 gnd.n6731 gnd.n6730 225.874
R13456 gnd.n6732 gnd.n6731 225.874
R13457 gnd.n6732 gnd.n675 225.874
R13458 gnd.n6740 gnd.n675 225.874
R13459 gnd.n6741 gnd.n6740 225.874
R13460 gnd.n6742 gnd.n6741 225.874
R13461 gnd.n6742 gnd.n669 225.874
R13462 gnd.n6750 gnd.n669 225.874
R13463 gnd.n6751 gnd.n6750 225.874
R13464 gnd.n6752 gnd.n6751 225.874
R13465 gnd.n6752 gnd.n663 225.874
R13466 gnd.n6760 gnd.n663 225.874
R13467 gnd.n6761 gnd.n6760 225.874
R13468 gnd.n6762 gnd.n6761 225.874
R13469 gnd.n6762 gnd.n657 225.874
R13470 gnd.n6770 gnd.n657 225.874
R13471 gnd.n6771 gnd.n6770 225.874
R13472 gnd.n6772 gnd.n6771 225.874
R13473 gnd.n6772 gnd.n651 225.874
R13474 gnd.n6780 gnd.n651 225.874
R13475 gnd.n6781 gnd.n6780 225.874
R13476 gnd.n6782 gnd.n6781 225.874
R13477 gnd.n6782 gnd.n645 225.874
R13478 gnd.n6790 gnd.n645 225.874
R13479 gnd.n6791 gnd.n6790 225.874
R13480 gnd.n6792 gnd.n6791 225.874
R13481 gnd.n6792 gnd.n639 225.874
R13482 gnd.n6800 gnd.n639 225.874
R13483 gnd.n6801 gnd.n6800 225.874
R13484 gnd.n6802 gnd.n6801 225.874
R13485 gnd.n6802 gnd.n633 225.874
R13486 gnd.n6810 gnd.n633 225.874
R13487 gnd.n6811 gnd.n6810 225.874
R13488 gnd.n6812 gnd.n6811 225.874
R13489 gnd.n6812 gnd.n627 225.874
R13490 gnd.n6820 gnd.n627 225.874
R13491 gnd.n6821 gnd.n6820 225.874
R13492 gnd.n6822 gnd.n6821 225.874
R13493 gnd.n6822 gnd.n621 225.874
R13494 gnd.n6830 gnd.n621 225.874
R13495 gnd.n6831 gnd.n6830 225.874
R13496 gnd.n6832 gnd.n6831 225.874
R13497 gnd.n6832 gnd.n615 225.874
R13498 gnd.n6840 gnd.n615 225.874
R13499 gnd.n6841 gnd.n6840 225.874
R13500 gnd.n6842 gnd.n6841 225.874
R13501 gnd.n6842 gnd.n609 225.874
R13502 gnd.n6850 gnd.n609 225.874
R13503 gnd.n6851 gnd.n6850 225.874
R13504 gnd.n6852 gnd.n6851 225.874
R13505 gnd.n6852 gnd.n603 225.874
R13506 gnd.n6860 gnd.n603 225.874
R13507 gnd.n6861 gnd.n6860 225.874
R13508 gnd.n6862 gnd.n6861 225.874
R13509 gnd.n6862 gnd.n597 225.874
R13510 gnd.n6870 gnd.n597 225.874
R13511 gnd.n6871 gnd.n6870 225.874
R13512 gnd.n6872 gnd.n6871 225.874
R13513 gnd.n6872 gnd.n591 225.874
R13514 gnd.n6880 gnd.n591 225.874
R13515 gnd.n6881 gnd.n6880 225.874
R13516 gnd.n6882 gnd.n6881 225.874
R13517 gnd.n6882 gnd.n585 225.874
R13518 gnd.n6890 gnd.n585 225.874
R13519 gnd.n6891 gnd.n6890 225.874
R13520 gnd.n6892 gnd.n6891 225.874
R13521 gnd.n6892 gnd.n579 225.874
R13522 gnd.n6900 gnd.n579 225.874
R13523 gnd.n6901 gnd.n6900 225.874
R13524 gnd.n6902 gnd.n6901 225.874
R13525 gnd.n6902 gnd.n573 225.874
R13526 gnd.n6910 gnd.n573 225.874
R13527 gnd.n6911 gnd.n6910 225.874
R13528 gnd.n6912 gnd.n6911 225.874
R13529 gnd.n6912 gnd.n567 225.874
R13530 gnd.n6920 gnd.n567 225.874
R13531 gnd.n6921 gnd.n6920 225.874
R13532 gnd.n6922 gnd.n6921 225.874
R13533 gnd.n6922 gnd.n561 225.874
R13534 gnd.n6930 gnd.n561 225.874
R13535 gnd.n6931 gnd.n6930 225.874
R13536 gnd.n6932 gnd.n6931 225.874
R13537 gnd.n6932 gnd.n555 225.874
R13538 gnd.n6940 gnd.n555 225.874
R13539 gnd.n6941 gnd.n6940 225.874
R13540 gnd.n6942 gnd.n6941 225.874
R13541 gnd.n6942 gnd.n549 225.874
R13542 gnd.n6950 gnd.n549 225.874
R13543 gnd.n6951 gnd.n6950 225.874
R13544 gnd.n6952 gnd.n6951 225.874
R13545 gnd.n6952 gnd.n543 225.874
R13546 gnd.n6960 gnd.n543 225.874
R13547 gnd.n6961 gnd.n6960 225.874
R13548 gnd.n6962 gnd.n6961 225.874
R13549 gnd.n6962 gnd.n537 225.874
R13550 gnd.n6970 gnd.n537 225.874
R13551 gnd.n6971 gnd.n6970 225.874
R13552 gnd.n6972 gnd.n6971 225.874
R13553 gnd.n6972 gnd.n531 225.874
R13554 gnd.n6980 gnd.n531 225.874
R13555 gnd.n6981 gnd.n6980 225.874
R13556 gnd.n6982 gnd.n6981 225.874
R13557 gnd.n6982 gnd.n525 225.874
R13558 gnd.n6990 gnd.n525 225.874
R13559 gnd.n6991 gnd.n6990 225.874
R13560 gnd.n6992 gnd.n6991 225.874
R13561 gnd.n6992 gnd.n519 225.874
R13562 gnd.n7000 gnd.n519 225.874
R13563 gnd.n7001 gnd.n7000 225.874
R13564 gnd.n7002 gnd.n7001 225.874
R13565 gnd.n7002 gnd.n513 225.874
R13566 gnd.n7010 gnd.n513 225.874
R13567 gnd.n7011 gnd.n7010 225.874
R13568 gnd.n7012 gnd.n7011 225.874
R13569 gnd.n7012 gnd.n507 225.874
R13570 gnd.n7020 gnd.n507 225.874
R13571 gnd.n7021 gnd.n7020 225.874
R13572 gnd.n7022 gnd.n7021 225.874
R13573 gnd.n7022 gnd.n501 225.874
R13574 gnd.n7030 gnd.n501 225.874
R13575 gnd.n7031 gnd.n7030 225.874
R13576 gnd.n7032 gnd.n7031 225.874
R13577 gnd.n7032 gnd.n495 225.874
R13578 gnd.n7040 gnd.n495 225.874
R13579 gnd.n7041 gnd.n7040 225.874
R13580 gnd.n7042 gnd.n7041 225.874
R13581 gnd.n7042 gnd.n489 225.874
R13582 gnd.n7050 gnd.n489 225.874
R13583 gnd.n7051 gnd.n7050 225.874
R13584 gnd.n7052 gnd.n7051 225.874
R13585 gnd.n7052 gnd.n483 225.874
R13586 gnd.n7060 gnd.n483 225.874
R13587 gnd.n7061 gnd.n7060 225.874
R13588 gnd.n7062 gnd.n7061 225.874
R13589 gnd.n7062 gnd.n477 225.874
R13590 gnd.n7070 gnd.n477 225.874
R13591 gnd.n7071 gnd.n7070 225.874
R13592 gnd.n7072 gnd.n7071 225.874
R13593 gnd.n7072 gnd.n471 225.874
R13594 gnd.n7080 gnd.n471 225.874
R13595 gnd.n7081 gnd.n7080 225.874
R13596 gnd.n7082 gnd.n7081 225.874
R13597 gnd.n7082 gnd.n465 225.874
R13598 gnd.n7090 gnd.n465 225.874
R13599 gnd.n7091 gnd.n7090 225.874
R13600 gnd.n7092 gnd.n7091 225.874
R13601 gnd.n7092 gnd.n459 225.874
R13602 gnd.n7100 gnd.n459 225.874
R13603 gnd.n7101 gnd.n7100 225.874
R13604 gnd.n7102 gnd.n7101 225.874
R13605 gnd.n7102 gnd.n453 225.874
R13606 gnd.n7110 gnd.n453 225.874
R13607 gnd.n7111 gnd.n7110 225.874
R13608 gnd.n7112 gnd.n7111 225.874
R13609 gnd.n7112 gnd.n447 225.874
R13610 gnd.n7120 gnd.n447 225.874
R13611 gnd.n7121 gnd.n7120 225.874
R13612 gnd.n7122 gnd.n7121 225.874
R13613 gnd.n7122 gnd.n441 225.874
R13614 gnd.n7130 gnd.n441 225.874
R13615 gnd.n7131 gnd.n7130 225.874
R13616 gnd.n7132 gnd.n7131 225.874
R13617 gnd.n7132 gnd.n435 225.874
R13618 gnd.n7140 gnd.n435 225.874
R13619 gnd.n7141 gnd.n7140 225.874
R13620 gnd.n7142 gnd.n7141 225.874
R13621 gnd.n7142 gnd.n429 225.874
R13622 gnd.n7150 gnd.n429 225.874
R13623 gnd.n7151 gnd.n7150 225.874
R13624 gnd.n7152 gnd.n7151 225.874
R13625 gnd.n7152 gnd.n423 225.874
R13626 gnd.n7160 gnd.n423 225.874
R13627 gnd.n7161 gnd.n7160 225.874
R13628 gnd.n7162 gnd.n7161 225.874
R13629 gnd.n7162 gnd.n417 225.874
R13630 gnd.n7170 gnd.n417 225.874
R13631 gnd.n7171 gnd.n7170 225.874
R13632 gnd.n7172 gnd.n7171 225.874
R13633 gnd.n7172 gnd.n411 225.874
R13634 gnd.n7180 gnd.n411 225.874
R13635 gnd.n7181 gnd.n7180 225.874
R13636 gnd.n7182 gnd.n7181 225.874
R13637 gnd.n7182 gnd.n405 225.874
R13638 gnd.n7190 gnd.n405 225.874
R13639 gnd.n7191 gnd.n7190 225.874
R13640 gnd.n7192 gnd.n7191 225.874
R13641 gnd.n7192 gnd.n399 225.874
R13642 gnd.n7201 gnd.n399 225.874
R13643 gnd.n7202 gnd.n7201 225.874
R13644 gnd.n7203 gnd.n7202 225.874
R13645 gnd.n7203 gnd.n394 225.874
R13646 gnd.n1430 gnd.t50 224.174
R13647 gnd.n942 gnd.t39 224.174
R13648 gnd.n5641 gnd.n5640 199.319
R13649 gnd.n5642 gnd.n5641 199.319
R13650 gnd.n2752 gnd.n2707 199.319
R13651 gnd.n2752 gnd.n2706 199.319
R13652 gnd.n2897 gnd.n2894 186.49
R13653 gnd.n5401 gnd.n5398 186.49
R13654 gnd.n2207 gnd.n2206 185
R13655 gnd.n2205 gnd.n2204 185
R13656 gnd.n2184 gnd.n2183 185
R13657 gnd.n2199 gnd.n2198 185
R13658 gnd.n2197 gnd.n2196 185
R13659 gnd.n2188 gnd.n2187 185
R13660 gnd.n2191 gnd.n2190 185
R13661 gnd.n2175 gnd.n2174 185
R13662 gnd.n2173 gnd.n2172 185
R13663 gnd.n2152 gnd.n2151 185
R13664 gnd.n2167 gnd.n2166 185
R13665 gnd.n2165 gnd.n2164 185
R13666 gnd.n2156 gnd.n2155 185
R13667 gnd.n2159 gnd.n2158 185
R13668 gnd.n2143 gnd.n2142 185
R13669 gnd.n2141 gnd.n2140 185
R13670 gnd.n2120 gnd.n2119 185
R13671 gnd.n2135 gnd.n2134 185
R13672 gnd.n2133 gnd.n2132 185
R13673 gnd.n2124 gnd.n2123 185
R13674 gnd.n2127 gnd.n2126 185
R13675 gnd.n2112 gnd.n2111 185
R13676 gnd.n2110 gnd.n2109 185
R13677 gnd.n2089 gnd.n2088 185
R13678 gnd.n2104 gnd.n2103 185
R13679 gnd.n2102 gnd.n2101 185
R13680 gnd.n2093 gnd.n2092 185
R13681 gnd.n2096 gnd.n2095 185
R13682 gnd.n2080 gnd.n2079 185
R13683 gnd.n2078 gnd.n2077 185
R13684 gnd.n2057 gnd.n2056 185
R13685 gnd.n2072 gnd.n2071 185
R13686 gnd.n2070 gnd.n2069 185
R13687 gnd.n2061 gnd.n2060 185
R13688 gnd.n2064 gnd.n2063 185
R13689 gnd.n2048 gnd.n2047 185
R13690 gnd.n2046 gnd.n2045 185
R13691 gnd.n2025 gnd.n2024 185
R13692 gnd.n2040 gnd.n2039 185
R13693 gnd.n2038 gnd.n2037 185
R13694 gnd.n2029 gnd.n2028 185
R13695 gnd.n2032 gnd.n2031 185
R13696 gnd.n2016 gnd.n2015 185
R13697 gnd.n2014 gnd.n2013 185
R13698 gnd.n1993 gnd.n1992 185
R13699 gnd.n2008 gnd.n2007 185
R13700 gnd.n2006 gnd.n2005 185
R13701 gnd.n1997 gnd.n1996 185
R13702 gnd.n2000 gnd.n1999 185
R13703 gnd.n1985 gnd.n1984 185
R13704 gnd.n1983 gnd.n1982 185
R13705 gnd.n1962 gnd.n1961 185
R13706 gnd.n1977 gnd.n1976 185
R13707 gnd.n1975 gnd.n1974 185
R13708 gnd.n1966 gnd.n1965 185
R13709 gnd.n1969 gnd.n1968 185
R13710 gnd.n1431 gnd.t49 178.987
R13711 gnd.n943 gnd.t40 178.987
R13712 gnd.n1 gnd.t8 170.774
R13713 gnd.n7 gnd.t186 170.103
R13714 gnd.n6 gnd.t313 170.103
R13715 gnd.n5 gnd.t183 170.103
R13716 gnd.n4 gnd.t323 170.103
R13717 gnd.n3 gnd.t315 170.103
R13718 gnd.n2 gnd.t19 170.103
R13719 gnd.n1 gnd.t176 170.103
R13720 gnd.n5469 gnd.n5468 163.367
R13721 gnd.n5465 gnd.n5464 163.367
R13722 gnd.n5461 gnd.n5460 163.367
R13723 gnd.n5457 gnd.n5456 163.367
R13724 gnd.n5453 gnd.n5452 163.367
R13725 gnd.n5449 gnd.n5448 163.367
R13726 gnd.n5445 gnd.n5444 163.367
R13727 gnd.n5441 gnd.n5440 163.367
R13728 gnd.n5437 gnd.n5436 163.367
R13729 gnd.n5433 gnd.n5432 163.367
R13730 gnd.n5429 gnd.n5428 163.367
R13731 gnd.n5425 gnd.n5424 163.367
R13732 gnd.n5421 gnd.n5420 163.367
R13733 gnd.n5417 gnd.n5416 163.367
R13734 gnd.n5412 gnd.n5411 163.367
R13735 gnd.n5544 gnd.n3302 163.367
R13736 gnd.n5541 gnd.n5540 163.367
R13737 gnd.n5538 gnd.n3335 163.367
R13738 gnd.n5533 gnd.n5532 163.367
R13739 gnd.n5529 gnd.n5528 163.367
R13740 gnd.n5525 gnd.n5524 163.367
R13741 gnd.n5521 gnd.n5520 163.367
R13742 gnd.n5517 gnd.n5516 163.367
R13743 gnd.n5513 gnd.n5512 163.367
R13744 gnd.n5509 gnd.n5508 163.367
R13745 gnd.n5505 gnd.n5504 163.367
R13746 gnd.n5501 gnd.n5500 163.367
R13747 gnd.n5497 gnd.n5496 163.367
R13748 gnd.n5493 gnd.n5492 163.367
R13749 gnd.n5489 gnd.n5488 163.367
R13750 gnd.n5485 gnd.n5484 163.367
R13751 gnd.n5481 gnd.n5480 163.367
R13752 gnd.n3823 gnd.n2913 163.367
R13753 gnd.n4502 gnd.n2913 163.367
R13754 gnd.n4502 gnd.n3749 163.367
R13755 gnd.n4506 gnd.n3749 163.367
R13756 gnd.n4506 gnd.n2922 163.367
R13757 gnd.n4519 gnd.n2922 163.367
R13758 gnd.n4519 gnd.n2931 163.367
R13759 gnd.n3735 gnd.n2931 163.367
R13760 gnd.n4532 gnd.n3735 163.367
R13761 gnd.n4532 gnd.n3736 163.367
R13762 gnd.n4528 gnd.n3736 163.367
R13763 gnd.n4528 gnd.n4527 163.367
R13764 gnd.n4527 gnd.n3725 163.367
R13765 gnd.n3725 gnd.n3717 163.367
R13766 gnd.n4569 gnd.n3717 163.367
R13767 gnd.n4569 gnd.n3715 163.367
R13768 gnd.n4584 gnd.n3715 163.367
R13769 gnd.n4584 gnd.n3706 163.367
R13770 gnd.n4580 gnd.n3706 163.367
R13771 gnd.n4580 gnd.n3701 163.367
R13772 gnd.n4577 gnd.n3701 163.367
R13773 gnd.n4577 gnd.n3689 163.367
R13774 gnd.n4573 gnd.n3689 163.367
R13775 gnd.n4573 gnd.n3682 163.367
R13776 gnd.n4641 gnd.n3682 163.367
R13777 gnd.n4641 gnd.n3680 163.367
R13778 gnd.n4666 gnd.n3680 163.367
R13779 gnd.n4666 gnd.n3674 163.367
R13780 gnd.n4662 gnd.n3674 163.367
R13781 gnd.n4662 gnd.n3665 163.367
R13782 gnd.n4657 gnd.n3665 163.367
R13783 gnd.n4657 gnd.n3660 163.367
R13784 gnd.n4654 gnd.n3660 163.367
R13785 gnd.n4654 gnd.n3653 163.367
R13786 gnd.n4649 gnd.n3653 163.367
R13787 gnd.n4649 gnd.n3647 163.367
R13788 gnd.n4646 gnd.n3647 163.367
R13789 gnd.n4646 gnd.n3637 163.367
R13790 gnd.n3637 gnd.n3629 163.367
R13791 gnd.n4766 gnd.n3629 163.367
R13792 gnd.n4766 gnd.n3627 163.367
R13793 gnd.n4773 gnd.n3627 163.367
R13794 gnd.n4773 gnd.n3617 163.367
R13795 gnd.n4769 gnd.n3617 163.367
R13796 gnd.n4769 gnd.n3612 163.367
R13797 gnd.n4796 gnd.n3612 163.367
R13798 gnd.n4796 gnd.n3605 163.367
R13799 gnd.n4800 gnd.n3605 163.367
R13800 gnd.n4800 gnd.n3597 163.367
R13801 gnd.n4820 gnd.n3597 163.367
R13802 gnd.n4820 gnd.n3595 163.367
R13803 gnd.n4844 gnd.n3595 163.367
R13804 gnd.n4844 gnd.n3588 163.367
R13805 gnd.n4840 gnd.n3588 163.367
R13806 gnd.n4840 gnd.n3580 163.367
R13807 gnd.n4836 gnd.n3580 163.367
R13808 gnd.n4836 gnd.n3574 163.367
R13809 gnd.n4833 gnd.n3574 163.367
R13810 gnd.n4833 gnd.n3566 163.367
R13811 gnd.n4828 gnd.n3566 163.367
R13812 gnd.n4828 gnd.n3560 163.367
R13813 gnd.n4825 gnd.n3560 163.367
R13814 gnd.n4825 gnd.n3550 163.367
R13815 gnd.n3550 gnd.n3543 163.367
R13816 gnd.n4921 gnd.n3543 163.367
R13817 gnd.n4921 gnd.n3541 163.367
R13818 gnd.n4929 gnd.n3541 163.367
R13819 gnd.n4929 gnd.n3531 163.367
R13820 gnd.n4925 gnd.n3531 163.367
R13821 gnd.n4925 gnd.n3524 163.367
R13822 gnd.n3524 gnd.n3516 163.367
R13823 gnd.n4973 gnd.n3516 163.367
R13824 gnd.n4973 gnd.n3514 163.367
R13825 gnd.n4997 gnd.n3514 163.367
R13826 gnd.n4997 gnd.n3509 163.367
R13827 gnd.n4993 gnd.n3509 163.367
R13828 gnd.n4993 gnd.n3501 163.367
R13829 gnd.n4988 gnd.n3501 163.367
R13830 gnd.n4988 gnd.n3496 163.367
R13831 gnd.n4985 gnd.n3496 163.367
R13832 gnd.n4985 gnd.n3488 163.367
R13833 gnd.n4981 gnd.n3488 163.367
R13834 gnd.n4981 gnd.n3482 163.367
R13835 gnd.n4978 gnd.n3482 163.367
R13836 gnd.n4978 gnd.n3474 163.367
R13837 gnd.n3474 gnd.n3467 163.367
R13838 gnd.n5078 gnd.n3467 163.367
R13839 gnd.n5078 gnd.n3465 163.367
R13840 gnd.n5082 gnd.n3465 163.367
R13841 gnd.n5082 gnd.n3426 163.367
R13842 gnd.n5102 gnd.n3426 163.367
R13843 gnd.n5102 gnd.n3421 163.367
R13844 gnd.n5098 gnd.n3421 163.367
R13845 gnd.n5098 gnd.n3412 163.367
R13846 gnd.n3455 gnd.n3412 163.367
R13847 gnd.n3455 gnd.n3406 163.367
R13848 gnd.n3452 gnd.n3406 163.367
R13849 gnd.n3452 gnd.n3399 163.367
R13850 gnd.n3447 gnd.n3399 163.367
R13851 gnd.n3447 gnd.n3391 163.367
R13852 gnd.n3444 gnd.n3391 163.367
R13853 gnd.n3444 gnd.n3384 163.367
R13854 gnd.n3384 gnd.n3375 163.367
R13855 gnd.n3376 gnd.n3375 163.367
R13856 gnd.n3376 gnd.n3369 163.367
R13857 gnd.n3438 gnd.n3369 163.367
R13858 gnd.n3438 gnd.n3431 163.367
R13859 gnd.n3431 gnd.n3346 163.367
R13860 gnd.n3346 gnd.n3339 163.367
R13861 gnd.n5476 gnd.n3339 163.367
R13862 gnd.n2888 gnd.n2887 163.367
R13863 gnd.n6213 gnd.n2887 163.367
R13864 gnd.n6211 gnd.n6210 163.367
R13865 gnd.n6207 gnd.n6206 163.367
R13866 gnd.n6203 gnd.n6202 163.367
R13867 gnd.n6199 gnd.n6198 163.367
R13868 gnd.n6195 gnd.n6194 163.367
R13869 gnd.n6191 gnd.n6190 163.367
R13870 gnd.n6187 gnd.n6186 163.367
R13871 gnd.n6183 gnd.n6182 163.367
R13872 gnd.n6179 gnd.n6178 163.367
R13873 gnd.n6175 gnd.n6174 163.367
R13874 gnd.n6171 gnd.n6170 163.367
R13875 gnd.n6167 gnd.n6166 163.367
R13876 gnd.n6163 gnd.n6162 163.367
R13877 gnd.n6159 gnd.n6158 163.367
R13878 gnd.n6222 gnd.n2853 163.367
R13879 gnd.n3762 gnd.n3761 163.367
R13880 gnd.n3767 gnd.n3766 163.367
R13881 gnd.n3771 gnd.n3770 163.367
R13882 gnd.n3775 gnd.n3774 163.367
R13883 gnd.n3779 gnd.n3778 163.367
R13884 gnd.n3783 gnd.n3782 163.367
R13885 gnd.n3787 gnd.n3786 163.367
R13886 gnd.n3791 gnd.n3790 163.367
R13887 gnd.n3795 gnd.n3794 163.367
R13888 gnd.n3799 gnd.n3798 163.367
R13889 gnd.n3803 gnd.n3802 163.367
R13890 gnd.n3807 gnd.n3806 163.367
R13891 gnd.n3811 gnd.n3810 163.367
R13892 gnd.n3815 gnd.n3814 163.367
R13893 gnd.n3819 gnd.n3818 163.367
R13894 gnd.n6151 gnd.n2889 163.367
R13895 gnd.n6151 gnd.n2911 163.367
R13896 gnd.n3746 gnd.n2911 163.367
R13897 gnd.n3746 gnd.n2926 163.367
R13898 gnd.n6141 gnd.n2926 163.367
R13899 gnd.n6141 gnd.n2927 163.367
R13900 gnd.n6137 gnd.n2927 163.367
R13901 gnd.n6137 gnd.n2930 163.367
R13902 gnd.n4538 gnd.n2930 163.367
R13903 gnd.n4538 gnd.n4533 163.367
R13904 gnd.n4534 gnd.n4533 163.367
R13905 gnd.n4534 gnd.n3723 163.367
R13906 gnd.n4562 gnd.n3723 163.367
R13907 gnd.n4562 gnd.n3720 163.367
R13908 gnd.n4567 gnd.n3720 163.367
R13909 gnd.n4567 gnd.n3721 163.367
R13910 gnd.n3721 gnd.n3705 163.367
R13911 gnd.n4600 gnd.n3705 163.367
R13912 gnd.n4600 gnd.n3703 163.367
R13913 gnd.n4604 gnd.n3703 163.367
R13914 gnd.n4604 gnd.n3690 163.367
R13915 gnd.n4629 gnd.n3690 163.367
R13916 gnd.n4629 gnd.n3691 163.367
R13917 gnd.n4625 gnd.n3691 163.367
R13918 gnd.n4625 gnd.n3678 163.367
R13919 gnd.n4670 gnd.n3678 163.367
R13920 gnd.n4670 gnd.n3676 163.367
R13921 gnd.n4674 gnd.n3676 163.367
R13922 gnd.n4674 gnd.n3664 163.367
R13923 gnd.n4689 gnd.n3664 163.367
R13924 gnd.n4689 gnd.n3662 163.367
R13925 gnd.n4693 gnd.n3662 163.367
R13926 gnd.n4693 gnd.n3651 163.367
R13927 gnd.n4741 gnd.n3651 163.367
R13928 gnd.n4741 gnd.n3649 163.367
R13929 gnd.n4745 gnd.n3649 163.367
R13930 gnd.n4745 gnd.n3635 163.367
R13931 gnd.n4759 gnd.n3635 163.367
R13932 gnd.n4759 gnd.n3632 163.367
R13933 gnd.n4764 gnd.n3632 163.367
R13934 gnd.n4764 gnd.n3633 163.367
R13935 gnd.n3633 gnd.n3615 163.367
R13936 gnd.n4788 gnd.n3615 163.367
R13937 gnd.n4788 gnd.n3613 163.367
R13938 gnd.n4792 gnd.n3613 163.367
R13939 gnd.n4792 gnd.n3608 163.367
R13940 gnd.n4808 gnd.n3608 163.367
R13941 gnd.n4808 gnd.n3609 163.367
R13942 gnd.n4804 gnd.n3609 163.367
R13943 gnd.n4804 gnd.n3593 163.367
R13944 gnd.n4848 gnd.n3593 163.367
R13945 gnd.n4848 gnd.n3591 163.367
R13946 gnd.n4852 gnd.n3591 163.367
R13947 gnd.n4852 gnd.n3578 163.367
R13948 gnd.n4866 gnd.n3578 163.367
R13949 gnd.n4866 gnd.n3576 163.367
R13950 gnd.n4870 gnd.n3576 163.367
R13951 gnd.n4870 gnd.n3564 163.367
R13952 gnd.n4897 gnd.n3564 163.367
R13953 gnd.n4897 gnd.n3562 163.367
R13954 gnd.n4901 gnd.n3562 163.367
R13955 gnd.n4901 gnd.n3548 163.367
R13956 gnd.n4914 gnd.n3548 163.367
R13957 gnd.n4914 gnd.n3545 163.367
R13958 gnd.n4919 gnd.n3545 163.367
R13959 gnd.n4919 gnd.n3546 163.367
R13960 gnd.n3546 gnd.n3529 163.367
R13961 gnd.n4952 gnd.n3529 163.367
R13962 gnd.n4952 gnd.n3526 163.367
R13963 gnd.n4957 gnd.n3526 163.367
R13964 gnd.n4957 gnd.n3527 163.367
R13965 gnd.n3527 gnd.n3513 163.367
R13966 gnd.n5001 gnd.n3513 163.367
R13967 gnd.n5001 gnd.n3511 163.367
R13968 gnd.n5005 gnd.n3511 163.367
R13969 gnd.n5005 gnd.n3500 163.367
R13970 gnd.n5021 gnd.n3500 163.367
R13971 gnd.n5021 gnd.n3498 163.367
R13972 gnd.n5025 gnd.n3498 163.367
R13973 gnd.n5025 gnd.n3486 163.367
R13974 gnd.n5051 gnd.n3486 163.367
R13975 gnd.n5051 gnd.n3484 163.367
R13976 gnd.n5055 gnd.n3484 163.367
R13977 gnd.n5055 gnd.n3472 163.367
R13978 gnd.n5071 gnd.n3472 163.367
R13979 gnd.n5071 gnd.n3469 163.367
R13980 gnd.n5076 gnd.n3469 163.367
R13981 gnd.n5076 gnd.n3470 163.367
R13982 gnd.n3470 gnd.n3424 163.367
R13983 gnd.n5106 gnd.n3424 163.367
R13984 gnd.n5106 gnd.n3422 163.367
R13985 gnd.n5110 gnd.n3422 163.367
R13986 gnd.n5110 gnd.n3410 163.367
R13987 gnd.n5124 gnd.n3410 163.367
R13988 gnd.n5124 gnd.n3408 163.367
R13989 gnd.n5128 gnd.n3408 163.367
R13990 gnd.n5128 gnd.n3397 163.367
R13991 gnd.n5140 gnd.n3397 163.367
R13992 gnd.n5140 gnd.n3394 163.367
R13993 gnd.n5145 gnd.n3394 163.367
R13994 gnd.n5145 gnd.n3395 163.367
R13995 gnd.n3395 gnd.n3373 163.367
R13996 gnd.n5173 gnd.n3373 163.367
R13997 gnd.n5173 gnd.n3370 163.367
R13998 gnd.n5178 gnd.n3370 163.367
R13999 gnd.n5178 gnd.n3371 163.367
R14000 gnd.n3371 gnd.n3344 163.367
R14001 gnd.n5386 gnd.n3344 163.367
R14002 gnd.n5386 gnd.n3341 163.367
R14003 gnd.n5474 gnd.n3341 163.367
R14004 gnd.n5407 gnd.n5406 156.462
R14005 gnd.n2147 gnd.n2115 153.042
R14006 gnd.n2211 gnd.n2210 152.079
R14007 gnd.n2179 gnd.n2178 152.079
R14008 gnd.n2147 gnd.n2146 152.079
R14009 gnd.n2902 gnd.n2901 152
R14010 gnd.n2903 gnd.n2892 152
R14011 gnd.n2905 gnd.n2904 152
R14012 gnd.n2907 gnd.n2890 152
R14013 gnd.n2909 gnd.n2908 152
R14014 gnd.n5405 gnd.n5389 152
R14015 gnd.n5397 gnd.n5390 152
R14016 gnd.n5396 gnd.n5395 152
R14017 gnd.n5394 gnd.n5391 152
R14018 gnd.n5392 gnd.t123 150.546
R14019 gnd.t21 gnd.n2189 147.661
R14020 gnd.t317 gnd.n2157 147.661
R14021 gnd.t162 gnd.n2125 147.661
R14022 gnd.t188 gnd.n2094 147.661
R14023 gnd.t169 gnd.n2062 147.661
R14024 gnd.t327 gnd.n2030 147.661
R14025 gnd.t179 gnd.n1998 147.661
R14026 gnd.t15 gnd.n1967 147.661
R14027 gnd.n5543 gnd.n3301 143.351
R14028 gnd.n2869 gnd.n2852 143.351
R14029 gnd.n6221 gnd.n2852 143.351
R14030 gnd.n2899 gnd.t51 130.484
R14031 gnd.n2908 gnd.t109 126.766
R14032 gnd.n2906 gnd.t44 126.766
R14033 gnd.n2892 gnd.t72 126.766
R14034 gnd.n2900 gnd.t154 126.766
R14035 gnd.n5393 gnd.t100 126.766
R14036 gnd.n5395 gnd.t41 126.766
R14037 gnd.n5404 gnd.t90 126.766
R14038 gnd.n5406 gnd.t66 126.766
R14039 gnd.n2206 gnd.n2205 104.615
R14040 gnd.n2205 gnd.n2183 104.615
R14041 gnd.n2198 gnd.n2183 104.615
R14042 gnd.n2198 gnd.n2197 104.615
R14043 gnd.n2197 gnd.n2187 104.615
R14044 gnd.n2190 gnd.n2187 104.615
R14045 gnd.n2174 gnd.n2173 104.615
R14046 gnd.n2173 gnd.n2151 104.615
R14047 gnd.n2166 gnd.n2151 104.615
R14048 gnd.n2166 gnd.n2165 104.615
R14049 gnd.n2165 gnd.n2155 104.615
R14050 gnd.n2158 gnd.n2155 104.615
R14051 gnd.n2142 gnd.n2141 104.615
R14052 gnd.n2141 gnd.n2119 104.615
R14053 gnd.n2134 gnd.n2119 104.615
R14054 gnd.n2134 gnd.n2133 104.615
R14055 gnd.n2133 gnd.n2123 104.615
R14056 gnd.n2126 gnd.n2123 104.615
R14057 gnd.n2111 gnd.n2110 104.615
R14058 gnd.n2110 gnd.n2088 104.615
R14059 gnd.n2103 gnd.n2088 104.615
R14060 gnd.n2103 gnd.n2102 104.615
R14061 gnd.n2102 gnd.n2092 104.615
R14062 gnd.n2095 gnd.n2092 104.615
R14063 gnd.n2079 gnd.n2078 104.615
R14064 gnd.n2078 gnd.n2056 104.615
R14065 gnd.n2071 gnd.n2056 104.615
R14066 gnd.n2071 gnd.n2070 104.615
R14067 gnd.n2070 gnd.n2060 104.615
R14068 gnd.n2063 gnd.n2060 104.615
R14069 gnd.n2047 gnd.n2046 104.615
R14070 gnd.n2046 gnd.n2024 104.615
R14071 gnd.n2039 gnd.n2024 104.615
R14072 gnd.n2039 gnd.n2038 104.615
R14073 gnd.n2038 gnd.n2028 104.615
R14074 gnd.n2031 gnd.n2028 104.615
R14075 gnd.n2015 gnd.n2014 104.615
R14076 gnd.n2014 gnd.n1992 104.615
R14077 gnd.n2007 gnd.n1992 104.615
R14078 gnd.n2007 gnd.n2006 104.615
R14079 gnd.n2006 gnd.n1996 104.615
R14080 gnd.n1999 gnd.n1996 104.615
R14081 gnd.n1984 gnd.n1983 104.615
R14082 gnd.n1983 gnd.n1961 104.615
R14083 gnd.n1976 gnd.n1961 104.615
R14084 gnd.n1976 gnd.n1975 104.615
R14085 gnd.n1975 gnd.n1965 104.615
R14086 gnd.n1968 gnd.n1965 104.615
R14087 gnd.n1356 gnd.t119 100.632
R14088 gnd.n916 gnd.t143 100.632
R14089 gnd.n7658 gnd.n7657 99.6594
R14090 gnd.n7653 gnd.n7474 99.6594
R14091 gnd.n7649 gnd.n7473 99.6594
R14092 gnd.n7645 gnd.n7472 99.6594
R14093 gnd.n7641 gnd.n7471 99.6594
R14094 gnd.n7637 gnd.n7470 99.6594
R14095 gnd.n7633 gnd.n7469 99.6594
R14096 gnd.n7629 gnd.n7468 99.6594
R14097 gnd.n7622 gnd.n7467 99.6594
R14098 gnd.n7618 gnd.n7466 99.6594
R14099 gnd.n7614 gnd.n7465 99.6594
R14100 gnd.n7610 gnd.n7464 99.6594
R14101 gnd.n7606 gnd.n7463 99.6594
R14102 gnd.n7602 gnd.n7462 99.6594
R14103 gnd.n7598 gnd.n7461 99.6594
R14104 gnd.n7594 gnd.n7460 99.6594
R14105 gnd.n7590 gnd.n7459 99.6594
R14106 gnd.n7586 gnd.n7458 99.6594
R14107 gnd.n7578 gnd.n7457 99.6594
R14108 gnd.n7576 gnd.n7456 99.6594
R14109 gnd.n7572 gnd.n7455 99.6594
R14110 gnd.n7568 gnd.n7454 99.6594
R14111 gnd.n7564 gnd.n7453 99.6594
R14112 gnd.n7560 gnd.n7452 99.6594
R14113 gnd.n7556 gnd.n7451 99.6594
R14114 gnd.n7552 gnd.n7450 99.6594
R14115 gnd.n7548 gnd.n7449 99.6594
R14116 gnd.n7544 gnd.n7448 99.6594
R14117 gnd.n7536 gnd.n7447 99.6594
R14118 gnd.n5575 gnd.n3061 99.6594
R14119 gnd.n5579 gnd.n5578 99.6594
R14120 gnd.n5586 gnd.n5585 99.6594
R14121 gnd.n5589 gnd.n5588 99.6594
R14122 gnd.n5596 gnd.n5595 99.6594
R14123 gnd.n5599 gnd.n5598 99.6594
R14124 gnd.n5606 gnd.n5605 99.6594
R14125 gnd.n5609 gnd.n5608 99.6594
R14126 gnd.n5619 gnd.n5618 99.6594
R14127 gnd.n5622 gnd.n5621 99.6594
R14128 gnd.n5629 gnd.n5628 99.6594
R14129 gnd.n5632 gnd.n5631 99.6594
R14130 gnd.n5640 gnd.n5639 99.6594
R14131 gnd.n5645 gnd.n5644 99.6594
R14132 gnd.n5652 gnd.n5651 99.6594
R14133 gnd.n5655 gnd.n5654 99.6594
R14134 gnd.n5662 gnd.n5661 99.6594
R14135 gnd.n5665 gnd.n5664 99.6594
R14136 gnd.n5674 gnd.n5673 99.6594
R14137 gnd.n5677 gnd.n5676 99.6594
R14138 gnd.n5684 gnd.n5683 99.6594
R14139 gnd.n5687 gnd.n5686 99.6594
R14140 gnd.n5694 gnd.n5693 99.6594
R14141 gnd.n5697 gnd.n5696 99.6594
R14142 gnd.n5704 gnd.n5703 99.6594
R14143 gnd.n5707 gnd.n5706 99.6594
R14144 gnd.n5715 gnd.n5714 99.6594
R14145 gnd.n5718 gnd.n5717 99.6594
R14146 gnd.n6273 gnd.n6272 99.6594
R14147 gnd.n6268 gnd.n2718 99.6594
R14148 gnd.n6264 gnd.n2717 99.6594
R14149 gnd.n6260 gnd.n2716 99.6594
R14150 gnd.n6256 gnd.n2715 99.6594
R14151 gnd.n6252 gnd.n2714 99.6594
R14152 gnd.n6248 gnd.n2713 99.6594
R14153 gnd.n6244 gnd.n2712 99.6594
R14154 gnd.n6239 gnd.n2711 99.6594
R14155 gnd.n6235 gnd.n2710 99.6594
R14156 gnd.n6231 gnd.n2709 99.6594
R14157 gnd.n6227 gnd.n2708 99.6594
R14158 gnd.n2844 gnd.n2706 99.6594
R14159 gnd.n2842 gnd.n2705 99.6594
R14160 gnd.n2838 gnd.n2704 99.6594
R14161 gnd.n2834 gnd.n2703 99.6594
R14162 gnd.n2830 gnd.n2702 99.6594
R14163 gnd.n2822 gnd.n2701 99.6594
R14164 gnd.n2820 gnd.n2700 99.6594
R14165 gnd.n2816 gnd.n2699 99.6594
R14166 gnd.n2812 gnd.n2698 99.6594
R14167 gnd.n2808 gnd.n2697 99.6594
R14168 gnd.n2804 gnd.n2696 99.6594
R14169 gnd.n2800 gnd.n2695 99.6594
R14170 gnd.n2796 gnd.n2694 99.6594
R14171 gnd.n2792 gnd.n2693 99.6594
R14172 gnd.n2788 gnd.n2692 99.6594
R14173 gnd.n2780 gnd.n2691 99.6594
R14174 gnd.n4064 gnd.n2368 99.6594
R14175 gnd.n4072 gnd.n4071 99.6594
R14176 gnd.n4075 gnd.n4074 99.6594
R14177 gnd.n4082 gnd.n4081 99.6594
R14178 gnd.n4085 gnd.n4084 99.6594
R14179 gnd.n4092 gnd.n4091 99.6594
R14180 gnd.n4095 gnd.n4094 99.6594
R14181 gnd.n4102 gnd.n4101 99.6594
R14182 gnd.n4105 gnd.n4104 99.6594
R14183 gnd.n4112 gnd.n4111 99.6594
R14184 gnd.n4115 gnd.n4114 99.6594
R14185 gnd.n4122 gnd.n4121 99.6594
R14186 gnd.n4125 gnd.n4124 99.6594
R14187 gnd.n4132 gnd.n4131 99.6594
R14188 gnd.n4135 gnd.n4134 99.6594
R14189 gnd.n4142 gnd.n4141 99.6594
R14190 gnd.n4145 gnd.n4144 99.6594
R14191 gnd.n4152 gnd.n4151 99.6594
R14192 gnd.n4155 gnd.n4154 99.6594
R14193 gnd.n4164 gnd.n4163 99.6594
R14194 gnd.n4167 gnd.n4166 99.6594
R14195 gnd.n4174 gnd.n4173 99.6594
R14196 gnd.n4177 gnd.n4176 99.6594
R14197 gnd.n4184 gnd.n4183 99.6594
R14198 gnd.n4187 gnd.n4186 99.6594
R14199 gnd.n4194 gnd.n4193 99.6594
R14200 gnd.n4197 gnd.n4196 99.6594
R14201 gnd.n4205 gnd.n4204 99.6594
R14202 gnd.n4208 gnd.n4207 99.6594
R14203 gnd.n2329 gnd.n899 99.6594
R14204 gnd.n2327 gnd.n898 99.6594
R14205 gnd.n2323 gnd.n897 99.6594
R14206 gnd.n2319 gnd.n896 99.6594
R14207 gnd.n2315 gnd.n895 99.6594
R14208 gnd.n2311 gnd.n894 99.6594
R14209 gnd.n2307 gnd.n893 99.6594
R14210 gnd.n2239 gnd.n892 99.6594
R14211 gnd.n1568 gnd.n1299 99.6594
R14212 gnd.n1325 gnd.n1306 99.6594
R14213 gnd.n1327 gnd.n1307 99.6594
R14214 gnd.n1335 gnd.n1308 99.6594
R14215 gnd.n1337 gnd.n1309 99.6594
R14216 gnd.n1345 gnd.n1310 99.6594
R14217 gnd.n1347 gnd.n1311 99.6594
R14218 gnd.n1355 gnd.n1312 99.6594
R14219 gnd.n206 gnd.n185 99.6594
R14220 gnd.n212 gnd.n186 99.6594
R14221 gnd.n216 gnd.n187 99.6594
R14222 gnd.n222 gnd.n188 99.6594
R14223 gnd.n226 gnd.n189 99.6594
R14224 gnd.n232 gnd.n190 99.6594
R14225 gnd.n235 gnd.n191 99.6594
R14226 gnd.n242 gnd.n241 99.6594
R14227 gnd.n7661 gnd.n7660 99.6594
R14228 gnd.n5281 gnd.n5280 99.6594
R14229 gnd.n5297 gnd.n5296 99.6594
R14230 gnd.n5300 gnd.n5299 99.6594
R14231 gnd.n5316 gnd.n5315 99.6594
R14232 gnd.n5319 gnd.n5318 99.6594
R14233 gnd.n5335 gnd.n5334 99.6594
R14234 gnd.n5338 gnd.n5337 99.6594
R14235 gnd.n5355 gnd.n5354 99.6594
R14236 gnd.n5358 gnd.n5357 99.6594
R14237 gnd.n2297 gnd.n879 99.6594
R14238 gnd.n2293 gnd.n880 99.6594
R14239 gnd.n2289 gnd.n881 99.6594
R14240 gnd.n2285 gnd.n882 99.6594
R14241 gnd.n2281 gnd.n883 99.6594
R14242 gnd.n2277 gnd.n884 99.6594
R14243 gnd.n2273 gnd.n885 99.6594
R14244 gnd.n2269 gnd.n886 99.6594
R14245 gnd.n2265 gnd.n887 99.6594
R14246 gnd.n2261 gnd.n888 99.6594
R14247 gnd.n2257 gnd.n889 99.6594
R14248 gnd.n2253 gnd.n890 99.6594
R14249 gnd.n2249 gnd.n891 99.6594
R14250 gnd.n1483 gnd.n1482 99.6594
R14251 gnd.n1477 gnd.n1394 99.6594
R14252 gnd.n1474 gnd.n1395 99.6594
R14253 gnd.n1470 gnd.n1396 99.6594
R14254 gnd.n1466 gnd.n1397 99.6594
R14255 gnd.n1462 gnd.n1398 99.6594
R14256 gnd.n1458 gnd.n1399 99.6594
R14257 gnd.n1454 gnd.n1400 99.6594
R14258 gnd.n1450 gnd.n1401 99.6594
R14259 gnd.n1446 gnd.n1402 99.6594
R14260 gnd.n1442 gnd.n1403 99.6594
R14261 gnd.n1438 gnd.n1404 99.6594
R14262 gnd.n1485 gnd.n1393 99.6594
R14263 gnd.n2677 gnd.n2622 99.6594
R14264 gnd.n2679 gnd.n2631 99.6594
R14265 gnd.n2681 gnd.n2680 99.6594
R14266 gnd.n2682 gnd.n2640 99.6594
R14267 gnd.n2684 gnd.n2649 99.6594
R14268 gnd.n2686 gnd.n2685 99.6594
R14269 gnd.n2687 gnd.n2658 99.6594
R14270 gnd.n2689 gnd.n2670 99.6594
R14271 gnd.n6276 gnd.n6275 99.6594
R14272 gnd.n3997 gnd.n3996 99.6594
R14273 gnd.n3994 gnd.n3933 99.6594
R14274 gnd.n3990 gnd.n3989 99.6594
R14275 gnd.n3983 gnd.n3937 99.6594
R14276 gnd.n3982 gnd.n3981 99.6594
R14277 gnd.n3975 gnd.n3943 99.6594
R14278 gnd.n3974 gnd.n3973 99.6594
R14279 gnd.n3967 gnd.n3949 99.6594
R14280 gnd.n3966 gnd.n3965 99.6594
R14281 gnd.n3996 gnd.n3995 99.6594
R14282 gnd.n3991 gnd.n3933 99.6594
R14283 gnd.n3989 gnd.n3988 99.6594
R14284 gnd.n3984 gnd.n3983 99.6594
R14285 gnd.n3981 gnd.n3980 99.6594
R14286 gnd.n3976 gnd.n3975 99.6594
R14287 gnd.n3973 gnd.n3972 99.6594
R14288 gnd.n3968 gnd.n3967 99.6594
R14289 gnd.n3965 gnd.n3964 99.6594
R14290 gnd.n6275 gnd.n2675 99.6594
R14291 gnd.n2689 gnd.n2688 99.6594
R14292 gnd.n2687 gnd.n2657 99.6594
R14293 gnd.n2686 gnd.n2650 99.6594
R14294 gnd.n2684 gnd.n2683 99.6594
R14295 gnd.n2682 gnd.n2639 99.6594
R14296 gnd.n2681 gnd.n2632 99.6594
R14297 gnd.n2679 gnd.n2678 99.6594
R14298 gnd.n2677 gnd.n2621 99.6594
R14299 gnd.n1483 gnd.n1406 99.6594
R14300 gnd.n1475 gnd.n1394 99.6594
R14301 gnd.n1471 gnd.n1395 99.6594
R14302 gnd.n1467 gnd.n1396 99.6594
R14303 gnd.n1463 gnd.n1397 99.6594
R14304 gnd.n1459 gnd.n1398 99.6594
R14305 gnd.n1455 gnd.n1399 99.6594
R14306 gnd.n1451 gnd.n1400 99.6594
R14307 gnd.n1447 gnd.n1401 99.6594
R14308 gnd.n1443 gnd.n1402 99.6594
R14309 gnd.n1439 gnd.n1403 99.6594
R14310 gnd.n1435 gnd.n1404 99.6594
R14311 gnd.n1486 gnd.n1485 99.6594
R14312 gnd.n2252 gnd.n891 99.6594
R14313 gnd.n2256 gnd.n890 99.6594
R14314 gnd.n2260 gnd.n889 99.6594
R14315 gnd.n2264 gnd.n888 99.6594
R14316 gnd.n2268 gnd.n887 99.6594
R14317 gnd.n2272 gnd.n886 99.6594
R14318 gnd.n2276 gnd.n885 99.6594
R14319 gnd.n2280 gnd.n884 99.6594
R14320 gnd.n2284 gnd.n883 99.6594
R14321 gnd.n2288 gnd.n882 99.6594
R14322 gnd.n2292 gnd.n881 99.6594
R14323 gnd.n2296 gnd.n880 99.6594
R14324 gnd.n920 gnd.n879 99.6594
R14325 gnd.n5280 gnd.n5244 99.6594
R14326 gnd.n5298 gnd.n5297 99.6594
R14327 gnd.n5299 gnd.n5235 99.6594
R14328 gnd.n5317 gnd.n5316 99.6594
R14329 gnd.n5318 gnd.n5226 99.6594
R14330 gnd.n5336 gnd.n5335 99.6594
R14331 gnd.n5337 gnd.n5217 99.6594
R14332 gnd.n5356 gnd.n5355 99.6594
R14333 gnd.n5357 gnd.n5213 99.6594
R14334 gnd.n7660 gnd.n183 99.6594
R14335 gnd.n242 gnd.n192 99.6594
R14336 gnd.n233 gnd.n191 99.6594
R14337 gnd.n225 gnd.n190 99.6594
R14338 gnd.n223 gnd.n189 99.6594
R14339 gnd.n215 gnd.n188 99.6594
R14340 gnd.n213 gnd.n187 99.6594
R14341 gnd.n205 gnd.n186 99.6594
R14342 gnd.n203 gnd.n185 99.6594
R14343 gnd.n1569 gnd.n1568 99.6594
R14344 gnd.n1328 gnd.n1306 99.6594
R14345 gnd.n1334 gnd.n1307 99.6594
R14346 gnd.n1338 gnd.n1308 99.6594
R14347 gnd.n1344 gnd.n1309 99.6594
R14348 gnd.n1348 gnd.n1310 99.6594
R14349 gnd.n1354 gnd.n1311 99.6594
R14350 gnd.n1312 gnd.n1296 99.6594
R14351 gnd.n2306 gnd.n892 99.6594
R14352 gnd.n2310 gnd.n893 99.6594
R14353 gnd.n2314 gnd.n894 99.6594
R14354 gnd.n2318 gnd.n895 99.6594
R14355 gnd.n2322 gnd.n896 99.6594
R14356 gnd.n2326 gnd.n897 99.6594
R14357 gnd.n2330 gnd.n898 99.6594
R14358 gnd.n901 gnd.n899 99.6594
R14359 gnd.n4065 gnd.n4064 99.6594
R14360 gnd.n4073 gnd.n4072 99.6594
R14361 gnd.n4074 gnd.n4056 99.6594
R14362 gnd.n4083 gnd.n4082 99.6594
R14363 gnd.n4084 gnd.n4052 99.6594
R14364 gnd.n4093 gnd.n4092 99.6594
R14365 gnd.n4094 gnd.n4048 99.6594
R14366 gnd.n4103 gnd.n4102 99.6594
R14367 gnd.n4104 gnd.n4041 99.6594
R14368 gnd.n4113 gnd.n4112 99.6594
R14369 gnd.n4114 gnd.n4037 99.6594
R14370 gnd.n4123 gnd.n4122 99.6594
R14371 gnd.n4124 gnd.n4033 99.6594
R14372 gnd.n4133 gnd.n4132 99.6594
R14373 gnd.n4134 gnd.n4029 99.6594
R14374 gnd.n4143 gnd.n4142 99.6594
R14375 gnd.n4144 gnd.n4025 99.6594
R14376 gnd.n4153 gnd.n4152 99.6594
R14377 gnd.n4154 gnd.n4021 99.6594
R14378 gnd.n4165 gnd.n4164 99.6594
R14379 gnd.n4166 gnd.n4017 99.6594
R14380 gnd.n4175 gnd.n4174 99.6594
R14381 gnd.n4176 gnd.n4013 99.6594
R14382 gnd.n4185 gnd.n4184 99.6594
R14383 gnd.n4186 gnd.n4009 99.6594
R14384 gnd.n4195 gnd.n4194 99.6594
R14385 gnd.n4196 gnd.n4005 99.6594
R14386 gnd.n4206 gnd.n4205 99.6594
R14387 gnd.n4209 gnd.n4208 99.6594
R14388 gnd.n2787 gnd.n2691 99.6594
R14389 gnd.n2791 gnd.n2692 99.6594
R14390 gnd.n2795 gnd.n2693 99.6594
R14391 gnd.n2799 gnd.n2694 99.6594
R14392 gnd.n2803 gnd.n2695 99.6594
R14393 gnd.n2807 gnd.n2696 99.6594
R14394 gnd.n2811 gnd.n2697 99.6594
R14395 gnd.n2815 gnd.n2698 99.6594
R14396 gnd.n2819 gnd.n2699 99.6594
R14397 gnd.n2823 gnd.n2700 99.6594
R14398 gnd.n2829 gnd.n2701 99.6594
R14399 gnd.n2833 gnd.n2702 99.6594
R14400 gnd.n2837 gnd.n2703 99.6594
R14401 gnd.n2841 gnd.n2704 99.6594
R14402 gnd.n2845 gnd.n2705 99.6594
R14403 gnd.n6226 gnd.n2707 99.6594
R14404 gnd.n6230 gnd.n2708 99.6594
R14405 gnd.n6234 gnd.n2709 99.6594
R14406 gnd.n6238 gnd.n2710 99.6594
R14407 gnd.n6243 gnd.n2711 99.6594
R14408 gnd.n6247 gnd.n2712 99.6594
R14409 gnd.n6251 gnd.n2713 99.6594
R14410 gnd.n6255 gnd.n2714 99.6594
R14411 gnd.n6259 gnd.n2715 99.6594
R14412 gnd.n6263 gnd.n2716 99.6594
R14413 gnd.n6267 gnd.n2717 99.6594
R14414 gnd.n2720 gnd.n2718 99.6594
R14415 gnd.n6273 gnd.n2719 99.6594
R14416 gnd.n5576 gnd.n5575 99.6594
R14417 gnd.n5578 gnd.n5567 99.6594
R14418 gnd.n5587 gnd.n5586 99.6594
R14419 gnd.n5588 gnd.n5563 99.6594
R14420 gnd.n5597 gnd.n5596 99.6594
R14421 gnd.n5598 gnd.n5559 99.6594
R14422 gnd.n5607 gnd.n5606 99.6594
R14423 gnd.n5608 gnd.n5555 99.6594
R14424 gnd.n5620 gnd.n5619 99.6594
R14425 gnd.n5621 gnd.n5551 99.6594
R14426 gnd.n5630 gnd.n5629 99.6594
R14427 gnd.n5631 gnd.n5547 99.6594
R14428 gnd.n5643 gnd.n5642 99.6594
R14429 gnd.n5644 gnd.n3295 99.6594
R14430 gnd.n5653 gnd.n5652 99.6594
R14431 gnd.n5654 gnd.n3291 99.6594
R14432 gnd.n5663 gnd.n5662 99.6594
R14433 gnd.n5664 gnd.n3287 99.6594
R14434 gnd.n5675 gnd.n5674 99.6594
R14435 gnd.n5676 gnd.n3283 99.6594
R14436 gnd.n5685 gnd.n5684 99.6594
R14437 gnd.n5686 gnd.n3279 99.6594
R14438 gnd.n5695 gnd.n5694 99.6594
R14439 gnd.n5696 gnd.n3275 99.6594
R14440 gnd.n5705 gnd.n5704 99.6594
R14441 gnd.n5706 gnd.n3271 99.6594
R14442 gnd.n5716 gnd.n5715 99.6594
R14443 gnd.n5719 gnd.n5718 99.6594
R14444 gnd.n7543 gnd.n7447 99.6594
R14445 gnd.n7547 gnd.n7448 99.6594
R14446 gnd.n7551 gnd.n7449 99.6594
R14447 gnd.n7555 gnd.n7450 99.6594
R14448 gnd.n7559 gnd.n7451 99.6594
R14449 gnd.n7563 gnd.n7452 99.6594
R14450 gnd.n7567 gnd.n7453 99.6594
R14451 gnd.n7571 gnd.n7454 99.6594
R14452 gnd.n7575 gnd.n7455 99.6594
R14453 gnd.n7579 gnd.n7456 99.6594
R14454 gnd.n7585 gnd.n7457 99.6594
R14455 gnd.n7589 gnd.n7458 99.6594
R14456 gnd.n7593 gnd.n7459 99.6594
R14457 gnd.n7597 gnd.n7460 99.6594
R14458 gnd.n7601 gnd.n7461 99.6594
R14459 gnd.n7605 gnd.n7462 99.6594
R14460 gnd.n7609 gnd.n7463 99.6594
R14461 gnd.n7613 gnd.n7464 99.6594
R14462 gnd.n7617 gnd.n7465 99.6594
R14463 gnd.n7621 gnd.n7466 99.6594
R14464 gnd.n7628 gnd.n7467 99.6594
R14465 gnd.n7632 gnd.n7468 99.6594
R14466 gnd.n7636 gnd.n7469 99.6594
R14467 gnd.n7640 gnd.n7470 99.6594
R14468 gnd.n7644 gnd.n7471 99.6594
R14469 gnd.n7648 gnd.n7472 99.6594
R14470 gnd.n7652 gnd.n7473 99.6594
R14471 gnd.n7476 gnd.n7474 99.6594
R14472 gnd.n7658 gnd.n7475 99.6594
R14473 gnd.n6338 gnd.n6337 99.6594
R14474 gnd.n2608 gnd.n2588 99.6594
R14475 gnd.n2610 gnd.n2589 99.6594
R14476 gnd.n2614 gnd.n2590 99.6594
R14477 gnd.n2616 gnd.n2591 99.6594
R14478 gnd.n2626 gnd.n2592 99.6594
R14479 gnd.n2628 gnd.n2593 99.6594
R14480 gnd.n2636 gnd.n2594 99.6594
R14481 gnd.n2644 gnd.n2595 99.6594
R14482 gnd.n2646 gnd.n2596 99.6594
R14483 gnd.n2654 gnd.n2597 99.6594
R14484 gnd.n2662 gnd.n2598 99.6594
R14485 gnd.n2667 gnd.n2600 99.6594
R14486 gnd.n6340 gnd.n2585 99.6594
R14487 gnd.n6338 gnd.n2603 99.6594
R14488 gnd.n2609 gnd.n2588 99.6594
R14489 gnd.n2613 gnd.n2589 99.6594
R14490 gnd.n2615 gnd.n2590 99.6594
R14491 gnd.n2625 gnd.n2591 99.6594
R14492 gnd.n2627 gnd.n2592 99.6594
R14493 gnd.n2635 gnd.n2593 99.6594
R14494 gnd.n2643 gnd.n2594 99.6594
R14495 gnd.n2645 gnd.n2595 99.6594
R14496 gnd.n2653 gnd.n2596 99.6594
R14497 gnd.n2661 gnd.n2597 99.6594
R14498 gnd.n2663 gnd.n2598 99.6594
R14499 gnd.n2600 gnd.n2599 99.6594
R14500 gnd.n6341 gnd.n6340 99.6594
R14501 gnd.n5261 gnd.n5256 99.6594
R14502 gnd.n5265 gnd.n5263 99.6594
R14503 gnd.n5272 gnd.n5252 99.6594
R14504 gnd.n5276 gnd.n5274 99.6594
R14505 gnd.n5287 gnd.n5249 99.6594
R14506 gnd.n5291 gnd.n5289 99.6594
R14507 gnd.n5306 gnd.n5240 99.6594
R14508 gnd.n5310 gnd.n5308 99.6594
R14509 gnd.n5325 gnd.n5231 99.6594
R14510 gnd.n5329 gnd.n5327 99.6594
R14511 gnd.n5344 gnd.n5222 99.6594
R14512 gnd.n5347 gnd.n5346 99.6594
R14513 gnd.n5365 gnd.n5364 99.6594
R14514 gnd.n5368 gnd.n5367 99.6594
R14515 gnd.n5346 gnd.n5345 99.6594
R14516 gnd.n5328 gnd.n5222 99.6594
R14517 gnd.n5327 gnd.n5326 99.6594
R14518 gnd.n5309 gnd.n5231 99.6594
R14519 gnd.n5308 gnd.n5307 99.6594
R14520 gnd.n5290 gnd.n5240 99.6594
R14521 gnd.n5289 gnd.n5288 99.6594
R14522 gnd.n5275 gnd.n5249 99.6594
R14523 gnd.n5274 gnd.n5273 99.6594
R14524 gnd.n5264 gnd.n5252 99.6594
R14525 gnd.n5263 gnd.n5262 99.6594
R14526 gnd.n5256 gnd.n3035 99.6594
R14527 gnd.n5369 gnd.n5368 99.6594
R14528 gnd.n5366 gnd.n5365 99.6594
R14529 gnd.n2664 gnd.t115 98.63
R14530 gnd.n5214 gnd.t137 98.63
R14531 gnd.n2671 gnd.t152 98.63
R14532 gnd.n5614 gnd.t134 98.63
R14533 gnd.n5666 gnd.t122 98.63
R14534 gnd.n3267 gnd.t65 98.63
R14535 gnd.n7538 gnd.t70 98.63
R14536 gnd.n7517 gnd.t60 98.63
R14537 gnd.n7624 gnd.t127 98.63
R14538 gnd.n180 gnd.t146 98.63
R14539 gnd.n4045 gnd.t99 98.63
R14540 gnd.n4156 gnd.t81 98.63
R14541 gnd.n4001 gnd.t105 98.63
R14542 gnd.n3961 gnd.t57 98.63
R14543 gnd.n2741 gnd.t139 98.63
R14544 gnd.n2782 gnd.t88 98.63
R14545 gnd.n2761 gnd.t107 98.63
R14546 gnd.n5204 gnd.t95 98.63
R14547 gnd.n3758 gnd.t150 96.6984
R14548 gnd.n3336 gnd.t77 96.6984
R14549 gnd.n6155 gnd.t85 96.6906
R14550 gnd.n5408 gnd.t130 96.6906
R14551 gnd.n2899 gnd.n2898 81.8399
R14552 gnd.n1357 gnd.t118 74.8376
R14553 gnd.n917 gnd.t144 74.8376
R14554 gnd.n3759 gnd.t149 72.8438
R14555 gnd.n3337 gnd.t78 72.8438
R14556 gnd.n2900 gnd.n2893 72.8411
R14557 gnd.n2906 gnd.n2891 72.8411
R14558 gnd.n5404 gnd.n5403 72.8411
R14559 gnd.n2665 gnd.t114 72.836
R14560 gnd.n6156 gnd.t84 72.836
R14561 gnd.n5409 gnd.t131 72.836
R14562 gnd.n5215 gnd.t136 72.836
R14563 gnd.n2672 gnd.t153 72.836
R14564 gnd.n5615 gnd.t133 72.836
R14565 gnd.n5667 gnd.t121 72.836
R14566 gnd.n3268 gnd.t64 72.836
R14567 gnd.n7539 gnd.t71 72.836
R14568 gnd.n7518 gnd.t61 72.836
R14569 gnd.n7625 gnd.t128 72.836
R14570 gnd.n181 gnd.t147 72.836
R14571 gnd.n4046 gnd.t98 72.836
R14572 gnd.n4157 gnd.t80 72.836
R14573 gnd.n4002 gnd.t104 72.836
R14574 gnd.n3962 gnd.t56 72.836
R14575 gnd.n2742 gnd.t140 72.836
R14576 gnd.n2783 gnd.t89 72.836
R14577 gnd.n2762 gnd.t108 72.836
R14578 gnd.n5205 gnd.t96 72.836
R14579 gnd.n5469 gnd.n3304 71.676
R14580 gnd.n5465 gnd.n3305 71.676
R14581 gnd.n5461 gnd.n3306 71.676
R14582 gnd.n5457 gnd.n3307 71.676
R14583 gnd.n5453 gnd.n3308 71.676
R14584 gnd.n5449 gnd.n3309 71.676
R14585 gnd.n5445 gnd.n3310 71.676
R14586 gnd.n5441 gnd.n3311 71.676
R14587 gnd.n5437 gnd.n3312 71.676
R14588 gnd.n5433 gnd.n3313 71.676
R14589 gnd.n5429 gnd.n3314 71.676
R14590 gnd.n5425 gnd.n3315 71.676
R14591 gnd.n5421 gnd.n3316 71.676
R14592 gnd.n5417 gnd.n3317 71.676
R14593 gnd.n5412 gnd.n3318 71.676
R14594 gnd.n3319 gnd.n3302 71.676
R14595 gnd.n5541 gnd.n3301 71.676
R14596 gnd.n5539 gnd.n5538 71.676
R14597 gnd.n5533 gnd.n3334 71.676
R14598 gnd.n5529 gnd.n3333 71.676
R14599 gnd.n5525 gnd.n3332 71.676
R14600 gnd.n5521 gnd.n3331 71.676
R14601 gnd.n5517 gnd.n3330 71.676
R14602 gnd.n5513 gnd.n3329 71.676
R14603 gnd.n5509 gnd.n3328 71.676
R14604 gnd.n5505 gnd.n3327 71.676
R14605 gnd.n5501 gnd.n3326 71.676
R14606 gnd.n5497 gnd.n3325 71.676
R14607 gnd.n5493 gnd.n3324 71.676
R14608 gnd.n5489 gnd.n3323 71.676
R14609 gnd.n5485 gnd.n3322 71.676
R14610 gnd.n5481 gnd.n3321 71.676
R14611 gnd.n5477 gnd.n3320 71.676
R14612 gnd.n6219 gnd.n6218 71.676
R14613 gnd.n6213 gnd.n2855 71.676
R14614 gnd.n6210 gnd.n2856 71.676
R14615 gnd.n6206 gnd.n2857 71.676
R14616 gnd.n6202 gnd.n2858 71.676
R14617 gnd.n6198 gnd.n2859 71.676
R14618 gnd.n6194 gnd.n2860 71.676
R14619 gnd.n6190 gnd.n2861 71.676
R14620 gnd.n6186 gnd.n2862 71.676
R14621 gnd.n6182 gnd.n2863 71.676
R14622 gnd.n6178 gnd.n2864 71.676
R14623 gnd.n6174 gnd.n2865 71.676
R14624 gnd.n6170 gnd.n2866 71.676
R14625 gnd.n6166 gnd.n2867 71.676
R14626 gnd.n6162 gnd.n2868 71.676
R14627 gnd.n6158 gnd.n2869 71.676
R14628 gnd.n2870 gnd.n2853 71.676
R14629 gnd.n3762 gnd.n2871 71.676
R14630 gnd.n3767 gnd.n2872 71.676
R14631 gnd.n3771 gnd.n2873 71.676
R14632 gnd.n3775 gnd.n2874 71.676
R14633 gnd.n3779 gnd.n2875 71.676
R14634 gnd.n3783 gnd.n2876 71.676
R14635 gnd.n3787 gnd.n2877 71.676
R14636 gnd.n3791 gnd.n2878 71.676
R14637 gnd.n3795 gnd.n2879 71.676
R14638 gnd.n3799 gnd.n2880 71.676
R14639 gnd.n3803 gnd.n2881 71.676
R14640 gnd.n3807 gnd.n2882 71.676
R14641 gnd.n3811 gnd.n2883 71.676
R14642 gnd.n3815 gnd.n2884 71.676
R14643 gnd.n3819 gnd.n2885 71.676
R14644 gnd.n6219 gnd.n2888 71.676
R14645 gnd.n6211 gnd.n2855 71.676
R14646 gnd.n6207 gnd.n2856 71.676
R14647 gnd.n6203 gnd.n2857 71.676
R14648 gnd.n6199 gnd.n2858 71.676
R14649 gnd.n6195 gnd.n2859 71.676
R14650 gnd.n6191 gnd.n2860 71.676
R14651 gnd.n6187 gnd.n2861 71.676
R14652 gnd.n6183 gnd.n2862 71.676
R14653 gnd.n6179 gnd.n2863 71.676
R14654 gnd.n6175 gnd.n2864 71.676
R14655 gnd.n6171 gnd.n2865 71.676
R14656 gnd.n6167 gnd.n2866 71.676
R14657 gnd.n6163 gnd.n2867 71.676
R14658 gnd.n6159 gnd.n2868 71.676
R14659 gnd.n6222 gnd.n6221 71.676
R14660 gnd.n3761 gnd.n2870 71.676
R14661 gnd.n3766 gnd.n2871 71.676
R14662 gnd.n3770 gnd.n2872 71.676
R14663 gnd.n3774 gnd.n2873 71.676
R14664 gnd.n3778 gnd.n2874 71.676
R14665 gnd.n3782 gnd.n2875 71.676
R14666 gnd.n3786 gnd.n2876 71.676
R14667 gnd.n3790 gnd.n2877 71.676
R14668 gnd.n3794 gnd.n2878 71.676
R14669 gnd.n3798 gnd.n2879 71.676
R14670 gnd.n3802 gnd.n2880 71.676
R14671 gnd.n3806 gnd.n2881 71.676
R14672 gnd.n3810 gnd.n2882 71.676
R14673 gnd.n3814 gnd.n2883 71.676
R14674 gnd.n3818 gnd.n2884 71.676
R14675 gnd.n3757 gnd.n2885 71.676
R14676 gnd.n5480 gnd.n3320 71.676
R14677 gnd.n5484 gnd.n3321 71.676
R14678 gnd.n5488 gnd.n3322 71.676
R14679 gnd.n5492 gnd.n3323 71.676
R14680 gnd.n5496 gnd.n3324 71.676
R14681 gnd.n5500 gnd.n3325 71.676
R14682 gnd.n5504 gnd.n3326 71.676
R14683 gnd.n5508 gnd.n3327 71.676
R14684 gnd.n5512 gnd.n3328 71.676
R14685 gnd.n5516 gnd.n3329 71.676
R14686 gnd.n5520 gnd.n3330 71.676
R14687 gnd.n5524 gnd.n3331 71.676
R14688 gnd.n5528 gnd.n3332 71.676
R14689 gnd.n5532 gnd.n3333 71.676
R14690 gnd.n3335 gnd.n3334 71.676
R14691 gnd.n5540 gnd.n5539 71.676
R14692 gnd.n5544 gnd.n5543 71.676
R14693 gnd.n5411 gnd.n3319 71.676
R14694 gnd.n5416 gnd.n3318 71.676
R14695 gnd.n5420 gnd.n3317 71.676
R14696 gnd.n5424 gnd.n3316 71.676
R14697 gnd.n5428 gnd.n3315 71.676
R14698 gnd.n5432 gnd.n3314 71.676
R14699 gnd.n5436 gnd.n3313 71.676
R14700 gnd.n5440 gnd.n3312 71.676
R14701 gnd.n5444 gnd.n3311 71.676
R14702 gnd.n5448 gnd.n3310 71.676
R14703 gnd.n5452 gnd.n3309 71.676
R14704 gnd.n5456 gnd.n3308 71.676
R14705 gnd.n5460 gnd.n3307 71.676
R14706 gnd.n5464 gnd.n3306 71.676
R14707 gnd.n5468 gnd.n3305 71.676
R14708 gnd.n3342 gnd.n3304 71.676
R14709 gnd.n8 gnd.t2 69.1507
R14710 gnd.n14 gnd.t26 68.4792
R14711 gnd.n13 gnd.t321 68.4792
R14712 gnd.n12 gnd.t325 68.4792
R14713 gnd.n11 gnd.t36 68.4792
R14714 gnd.n10 gnd.t31 68.4792
R14715 gnd.n9 gnd.t319 68.4792
R14716 gnd.n8 gnd.t24 68.4792
R14717 gnd.n1484 gnd.n1388 64.369
R14718 gnd.n6512 gnd.n2339 59.5891
R14719 gnd.n7423 gnd.n7422 59.5891
R14720 gnd.n3764 gnd.n3759 59.5399
R14721 gnd.n5535 gnd.n3337 59.5399
R14722 gnd.n6157 gnd.n6156 59.5399
R14723 gnd.n5414 gnd.n5409 59.5399
R14724 gnd.n6154 gnd.n2909 59.1804
R14725 gnd.n2338 gnd.n877 57.3586
R14726 gnd.n1143 gnd.t249 56.407
R14727 gnd.n1108 gnd.t296 56.407
R14728 gnd.n1119 gnd.t208 56.407
R14729 gnd.n1131 gnd.t288 56.407
R14730 gnd.n52 gnd.t224 56.407
R14731 gnd.n17 gnd.t215 56.407
R14732 gnd.n28 gnd.t305 56.407
R14733 gnd.n40 gnd.t263 56.407
R14734 gnd.n1152 gnd.t275 55.8337
R14735 gnd.n1117 gnd.t204 55.8337
R14736 gnd.n1128 gnd.t307 55.8337
R14737 gnd.n1140 gnd.t210 55.8337
R14738 gnd.n61 gnd.t247 55.8337
R14739 gnd.n26 gnd.t239 55.8337
R14740 gnd.n37 gnd.t287 55.8337
R14741 gnd.n49 gnd.t285 55.8337
R14742 gnd.n2897 gnd.n2896 54.358
R14743 gnd.n5401 gnd.n5400 54.358
R14744 gnd.n1143 gnd.n1142 53.0052
R14745 gnd.n1145 gnd.n1144 53.0052
R14746 gnd.n1147 gnd.n1146 53.0052
R14747 gnd.n1149 gnd.n1148 53.0052
R14748 gnd.n1151 gnd.n1150 53.0052
R14749 gnd.n1108 gnd.n1107 53.0052
R14750 gnd.n1110 gnd.n1109 53.0052
R14751 gnd.n1112 gnd.n1111 53.0052
R14752 gnd.n1114 gnd.n1113 53.0052
R14753 gnd.n1116 gnd.n1115 53.0052
R14754 gnd.n1119 gnd.n1118 53.0052
R14755 gnd.n1121 gnd.n1120 53.0052
R14756 gnd.n1123 gnd.n1122 53.0052
R14757 gnd.n1125 gnd.n1124 53.0052
R14758 gnd.n1127 gnd.n1126 53.0052
R14759 gnd.n1131 gnd.n1130 53.0052
R14760 gnd.n1133 gnd.n1132 53.0052
R14761 gnd.n1135 gnd.n1134 53.0052
R14762 gnd.n1137 gnd.n1136 53.0052
R14763 gnd.n1139 gnd.n1138 53.0052
R14764 gnd.n60 gnd.n59 53.0052
R14765 gnd.n58 gnd.n57 53.0052
R14766 gnd.n56 gnd.n55 53.0052
R14767 gnd.n54 gnd.n53 53.0052
R14768 gnd.n52 gnd.n51 53.0052
R14769 gnd.n25 gnd.n24 53.0052
R14770 gnd.n23 gnd.n22 53.0052
R14771 gnd.n21 gnd.n20 53.0052
R14772 gnd.n19 gnd.n18 53.0052
R14773 gnd.n17 gnd.n16 53.0052
R14774 gnd.n36 gnd.n35 53.0052
R14775 gnd.n34 gnd.n33 53.0052
R14776 gnd.n32 gnd.n31 53.0052
R14777 gnd.n30 gnd.n29 53.0052
R14778 gnd.n28 gnd.n27 53.0052
R14779 gnd.n48 gnd.n47 53.0052
R14780 gnd.n46 gnd.n45 53.0052
R14781 gnd.n44 gnd.n43 53.0052
R14782 gnd.n42 gnd.n41 53.0052
R14783 gnd.n40 gnd.n39 53.0052
R14784 gnd.n5392 gnd.n5391 52.4801
R14785 gnd.n2190 gnd.t21 52.3082
R14786 gnd.n2158 gnd.t317 52.3082
R14787 gnd.n2126 gnd.t162 52.3082
R14788 gnd.n2095 gnd.t188 52.3082
R14789 gnd.n2063 gnd.t169 52.3082
R14790 gnd.n2031 gnd.t327 52.3082
R14791 gnd.n1999 gnd.t179 52.3082
R14792 gnd.n1968 gnd.t15 52.3082
R14793 gnd.n2020 gnd.n1988 51.4173
R14794 gnd.n2084 gnd.n2083 50.455
R14795 gnd.n2052 gnd.n2051 50.455
R14796 gnd.n2020 gnd.n2019 50.455
R14797 gnd.n5546 gnd.n5545 45.6325
R14798 gnd.n6224 gnd.n6223 45.6325
R14799 gnd.n1431 gnd.n1430 45.1884
R14800 gnd.n943 gnd.n942 45.1884
R14801 gnd.n5472 gnd.n5407 44.3322
R14802 gnd.n2900 gnd.n2899 44.3189
R14803 gnd.n6682 gnd.n705 43.8952
R14804 gnd.n6682 gnd.n6681 43.8952
R14805 gnd.n6681 gnd.n6680 43.8952
R14806 gnd.n6680 gnd.n710 43.8952
R14807 gnd.n6674 gnd.n710 43.8952
R14808 gnd.n6674 gnd.n6673 43.8952
R14809 gnd.n6673 gnd.n6672 43.8952
R14810 gnd.n6672 gnd.n718 43.8952
R14811 gnd.n6666 gnd.n718 43.8952
R14812 gnd.n6666 gnd.n6665 43.8952
R14813 gnd.n6665 gnd.n6664 43.8952
R14814 gnd.n6664 gnd.n726 43.8952
R14815 gnd.n6658 gnd.n726 43.8952
R14816 gnd.n6658 gnd.n6657 43.8952
R14817 gnd.n6657 gnd.n6656 43.8952
R14818 gnd.n6656 gnd.n734 43.8952
R14819 gnd.n6650 gnd.n734 43.8952
R14820 gnd.n6650 gnd.n6649 43.8952
R14821 gnd.n6649 gnd.n6648 43.8952
R14822 gnd.n6648 gnd.n742 43.8952
R14823 gnd.n6642 gnd.n742 43.8952
R14824 gnd.n6642 gnd.n6641 43.8952
R14825 gnd.n6641 gnd.n6640 43.8952
R14826 gnd.n6640 gnd.n750 43.8952
R14827 gnd.n6634 gnd.n750 43.8952
R14828 gnd.n6634 gnd.n6633 43.8952
R14829 gnd.n6633 gnd.n6632 43.8952
R14830 gnd.n6632 gnd.n758 43.8952
R14831 gnd.n6626 gnd.n758 43.8952
R14832 gnd.n6626 gnd.n6625 43.8952
R14833 gnd.n6625 gnd.n6624 43.8952
R14834 gnd.n6624 gnd.n766 43.8952
R14835 gnd.n6618 gnd.n766 43.8952
R14836 gnd.n6618 gnd.n6617 43.8952
R14837 gnd.n6617 gnd.n6616 43.8952
R14838 gnd.n6616 gnd.n774 43.8952
R14839 gnd.n6610 gnd.n774 43.8952
R14840 gnd.n6610 gnd.n6609 43.8952
R14841 gnd.n6609 gnd.n6608 43.8952
R14842 gnd.n6608 gnd.n782 43.8952
R14843 gnd.n6602 gnd.n782 43.8952
R14844 gnd.n6602 gnd.n6601 43.8952
R14845 gnd.n6601 gnd.n6600 43.8952
R14846 gnd.n6600 gnd.n790 43.8952
R14847 gnd.n6594 gnd.n790 43.8952
R14848 gnd.n6594 gnd.n6593 43.8952
R14849 gnd.n6593 gnd.n6592 43.8952
R14850 gnd.n6592 gnd.n798 43.8952
R14851 gnd.n6586 gnd.n798 43.8952
R14852 gnd.n6586 gnd.n6585 43.8952
R14853 gnd.n6585 gnd.n6584 43.8952
R14854 gnd.n6584 gnd.n806 43.8952
R14855 gnd.n6578 gnd.n806 43.8952
R14856 gnd.n6578 gnd.n6577 43.8952
R14857 gnd.n6577 gnd.n6576 43.8952
R14858 gnd.n6576 gnd.n814 43.8952
R14859 gnd.n6570 gnd.n814 43.8952
R14860 gnd.n6570 gnd.n6569 43.8952
R14861 gnd.n6569 gnd.n6568 43.8952
R14862 gnd.n6568 gnd.n822 43.8952
R14863 gnd.n6562 gnd.n822 43.8952
R14864 gnd.n6562 gnd.n6561 43.8952
R14865 gnd.n6561 gnd.n6560 43.8952
R14866 gnd.n6560 gnd.n830 43.8952
R14867 gnd.n6554 gnd.n830 43.8952
R14868 gnd.n6554 gnd.n6553 43.8952
R14869 gnd.n6553 gnd.n6552 43.8952
R14870 gnd.n6552 gnd.n838 43.8952
R14871 gnd.n6546 gnd.n838 43.8952
R14872 gnd.n6546 gnd.n6545 43.8952
R14873 gnd.n6545 gnd.n6544 43.8952
R14874 gnd.n6544 gnd.n846 43.8952
R14875 gnd.n6538 gnd.n846 43.8952
R14876 gnd.n6538 gnd.n6537 43.8952
R14877 gnd.n6537 gnd.n6536 43.8952
R14878 gnd.n6536 gnd.n854 43.8952
R14879 gnd.n6530 gnd.n854 43.8952
R14880 gnd.n6530 gnd.n6529 43.8952
R14881 gnd.n6529 gnd.n6528 43.8952
R14882 gnd.n6528 gnd.n862 43.8952
R14883 gnd.n6522 gnd.n862 43.8952
R14884 gnd.n6522 gnd.n6521 43.8952
R14885 gnd.n6521 gnd.n6520 43.8952
R14886 gnd.n2666 gnd.n2665 42.2793
R14887 gnd.n5360 gnd.n5215 42.2793
R14888 gnd.n1432 gnd.n1431 42.2793
R14889 gnd.n944 gnd.n943 42.2793
R14890 gnd.n1358 gnd.n1357 42.2793
R14891 gnd.n2305 gnd.n917 42.2793
R14892 gnd.n6278 gnd.n2672 42.2793
R14893 gnd.n5616 gnd.n5615 42.2793
R14894 gnd.n5668 gnd.n5667 42.2793
R14895 gnd.n3269 gnd.n3268 42.2793
R14896 gnd.n7542 gnd.n7539 42.2793
R14897 gnd.n7584 gnd.n7518 42.2793
R14898 gnd.n7626 gnd.n7625 42.2793
R14899 gnd.n182 gnd.n181 42.2793
R14900 gnd.n4047 gnd.n4046 42.2793
R14901 gnd.n4158 gnd.n4157 42.2793
R14902 gnd.n4003 gnd.n4002 42.2793
R14903 gnd.n3963 gnd.n3962 42.2793
R14904 gnd.n6241 gnd.n2742 42.2793
R14905 gnd.n2786 gnd.n2783 42.2793
R14906 gnd.n2828 gnd.n2762 42.2793
R14907 gnd.n5206 gnd.n5205 42.2793
R14908 gnd.n2898 gnd.n2897 41.6274
R14909 gnd.n5402 gnd.n5401 41.6274
R14910 gnd.n2907 gnd.n2906 40.8975
R14911 gnd.n5405 gnd.n5404 40.8975
R14912 gnd.n2906 gnd.n2905 35.055
R14913 gnd.n2901 gnd.n2900 35.055
R14914 gnd.n5394 gnd.n5393 35.055
R14915 gnd.n5404 gnd.n5390 35.055
R14916 gnd.n5478 gnd.n3338 32.9371
R14917 gnd.n3822 gnd.n3821 32.9371
R14918 gnd.n1494 gnd.n1388 31.8661
R14919 gnd.n1494 gnd.n1493 31.8661
R14920 gnd.n1502 gnd.n1377 31.8661
R14921 gnd.n1510 gnd.n1377 31.8661
R14922 gnd.n1510 gnd.n1371 31.8661
R14923 gnd.n1518 gnd.n1371 31.8661
R14924 gnd.n1518 gnd.n1364 31.8661
R14925 gnd.n1556 gnd.n1364 31.8661
R14926 gnd.n1566 gnd.n1297 31.8661
R14927 gnd.n6512 gnd.n6511 31.8661
R14928 gnd.n6511 gnd.n6510 31.8661
R14929 gnd.n6510 gnd.n2340 31.8661
R14930 gnd.n6504 gnd.n2340 31.8661
R14931 gnd.n6504 gnd.n6503 31.8661
R14932 gnd.n6503 gnd.n6502 31.8661
R14933 gnd.n6502 gnd.n2347 31.8661
R14934 gnd.n6496 gnd.n2347 31.8661
R14935 gnd.n6496 gnd.n6495 31.8661
R14936 gnd.n6495 gnd.n6494 31.8661
R14937 gnd.n6494 gnd.n2355 31.8661
R14938 gnd.n6488 gnd.n6487 31.8661
R14939 gnd.n2676 gnd.n2574 31.8661
R14940 gnd.n3843 gnd.n2690 31.8661
R14941 gnd.n3843 gnd.n2587 31.8661
R14942 gnd.n4464 gnd.n2601 31.8661
R14943 gnd.n6016 gnd.n3038 31.8661
R14944 gnd.n6010 gnd.n6009 31.8661
R14945 gnd.n6009 gnd.n6008 31.8661
R14946 gnd.n6002 gnd.n3056 31.8661
R14947 gnd.n184 gnd.n171 31.8661
R14948 gnd.n7446 gnd.n243 31.8661
R14949 gnd.n7440 gnd.n243 31.8661
R14950 gnd.n7440 gnd.n7439 31.8661
R14951 gnd.n7439 gnd.n7438 31.8661
R14952 gnd.n7438 gnd.n252 31.8661
R14953 gnd.n7432 gnd.n252 31.8661
R14954 gnd.n7432 gnd.n7431 31.8661
R14955 gnd.n7431 gnd.n7430 31.8661
R14956 gnd.n7430 gnd.n260 31.8661
R14957 gnd.n7424 gnd.n260 31.8661
R14958 gnd.n7424 gnd.n7423 31.8661
R14959 gnd.n6520 gnd.n870 26.3373
R14960 gnd.n2665 gnd.n2664 25.7944
R14961 gnd.n5215 gnd.n5214 25.7944
R14962 gnd.n1357 gnd.n1356 25.7944
R14963 gnd.n917 gnd.n916 25.7944
R14964 gnd.n2672 gnd.n2671 25.7944
R14965 gnd.n5615 gnd.n5614 25.7944
R14966 gnd.n5667 gnd.n5666 25.7944
R14967 gnd.n3268 gnd.n3267 25.7944
R14968 gnd.n7539 gnd.n7538 25.7944
R14969 gnd.n7518 gnd.n7517 25.7944
R14970 gnd.n7625 gnd.n7624 25.7944
R14971 gnd.n181 gnd.n180 25.7944
R14972 gnd.n4046 gnd.n4045 25.7944
R14973 gnd.n4157 gnd.n4156 25.7944
R14974 gnd.n4002 gnd.n4001 25.7944
R14975 gnd.n3962 gnd.n3961 25.7944
R14976 gnd.n2742 gnd.n2741 25.7944
R14977 gnd.n2783 gnd.n2782 25.7944
R14978 gnd.n2762 gnd.n2761 25.7944
R14979 gnd.n5205 gnd.n5204 25.7944
R14980 gnd.n1578 gnd.n1298 24.8557
R14981 gnd.n1588 gnd.n1281 24.8557
R14982 gnd.n1284 gnd.n1272 24.8557
R14983 gnd.n1609 gnd.n1273 24.8557
R14984 gnd.n1619 gnd.n1253 24.8557
R14985 gnd.n1629 gnd.n1628 24.8557
R14986 gnd.n1239 gnd.n1237 24.8557
R14987 gnd.n1660 gnd.n1659 24.8557
R14988 gnd.n1675 gnd.n1222 24.8557
R14989 gnd.n1729 gnd.n1161 24.8557
R14990 gnd.n1685 gnd.n1162 24.8557
R14991 gnd.n1722 gnd.n1173 24.8557
R14992 gnd.n1211 gnd.n1210 24.8557
R14993 gnd.n1716 gnd.n1715 24.8557
R14994 gnd.n1197 gnd.n1184 24.8557
R14995 gnd.n1755 gnd.n1754 24.8557
R14996 gnd.n1765 gnd.n1093 24.8557
R14997 gnd.n1777 gnd.n1085 24.8557
R14998 gnd.n1776 gnd.n1073 24.8557
R14999 gnd.n1795 gnd.n1794 24.8557
R15000 gnd.n1805 gnd.n1066 24.8557
R15001 gnd.n1816 gnd.n1054 24.8557
R15002 gnd.n1842 gnd.n1841 24.8557
R15003 gnd.n1852 gnd.n1040 24.8557
R15004 gnd.n1864 gnd.n1032 24.8557
R15005 gnd.n1882 gnd.n1881 24.8557
R15006 gnd.n1023 gnd.n1012 24.8557
R15007 gnd.n1903 gnd.n1000 24.8557
R15008 gnd.n1931 gnd.n1930 24.8557
R15009 gnd.n1942 gnd.n985 24.8557
R15010 gnd.n1953 gnd.n978 24.8557
R15011 gnd.n1952 gnd.n966 24.8557
R15012 gnd.n2225 gnd.n2224 24.8557
R15013 gnd.n2247 gnd.n951 24.8557
R15014 gnd.n3759 gnd.n3758 23.855
R15015 gnd.n3337 gnd.n3336 23.855
R15016 gnd.n6156 gnd.n6155 23.855
R15017 gnd.n5409 gnd.n5408 23.855
R15018 gnd.n1599 gnd.t14 23.2624
R15019 gnd.n1300 gnd.t117 22.6251
R15020 gnd.n2363 gnd.n2355 21.6691
R15021 gnd.n7659 gnd.n7446 21.6691
R15022 gnd.t187 gnd.n1305 21.3504
R15023 gnd.n6487 gnd.n6486 21.0318
R15024 gnd.n4256 gnd.n2366 21.0318
R15025 gnd.n4250 gnd.n2377 21.0318
R15026 gnd.n6474 gnd.n2386 21.0318
R15027 gnd.n4244 gnd.n2389 21.0318
R15028 gnd.n6468 gnd.n2397 21.0318
R15029 gnd.n6462 gnd.n2407 21.0318
R15030 gnd.n4232 gnd.n2410 21.0318
R15031 gnd.n6456 gnd.n2418 21.0318
R15032 gnd.n4287 gnd.n2421 21.0318
R15033 gnd.n4295 gnd.n2430 21.0318
R15034 gnd.n6444 gnd.n2438 21.0318
R15035 gnd.n6438 gnd.n2448 21.0318
R15036 gnd.n4310 gnd.n2451 21.0318
R15037 gnd.n6431 gnd.n2457 21.0318
R15038 gnd.n4354 gnd.n2460 21.0318
R15039 gnd.n4317 gnd.n2469 21.0318
R15040 gnd.n6418 gnd.n2474 21.0318
R15041 gnd.n4332 gnd.n4331 21.0318
R15042 gnd.n6412 gnd.n2483 21.0318
R15043 gnd.n6405 gnd.n2491 21.0318
R15044 gnd.n4390 gnd.n2494 21.0318
R15045 gnd.n4398 gnd.n2503 21.0318
R15046 gnd.n6393 gnd.n2511 21.0318
R15047 gnd.n4404 gnd.n3868 21.0318
R15048 gnd.n6387 gnd.n2520 21.0318
R15049 gnd.n6381 gnd.n2531 21.0318
R15050 gnd.n4436 gnd.n2534 21.0318
R15051 gnd.n4419 gnd.n2543 21.0318
R15052 gnd.n6369 gnd.n2551 21.0318
R15053 gnd.n4425 gnd.n2554 21.0318
R15054 gnd.n6363 gnd.n2561 21.0318
R15055 gnd.n6357 gnd.n2571 21.0318
R15056 gnd.n6001 gnd.n3059 21.0318
R15057 gnd.n5995 gnd.n3071 21.0318
R15058 gnd.n5730 gnd.n3080 21.0318
R15059 gnd.n5989 gnd.n3083 21.0318
R15060 gnd.n5738 gnd.n3091 21.0318
R15061 gnd.n5758 gnd.n3100 21.0318
R15062 gnd.n5977 gnd.n3103 21.0318
R15063 gnd.n5971 gnd.n3114 21.0318
R15064 gnd.n5803 gnd.n5802 21.0318
R15065 gnd.n5965 gnd.n3123 21.0318
R15066 gnd.n5810 gnd.n3131 21.0318
R15067 gnd.n5828 gnd.n3140 21.0318
R15068 gnd.n5953 gnd.n3143 21.0318
R15069 gnd.n3155 gnd.n3149 21.0318
R15070 gnd.n5941 gnd.n3156 21.0318
R15071 gnd.n5940 gnd.n3159 21.0318
R15072 gnd.n5935 gnd.n3166 21.0318
R15073 gnd.n7731 gnd.n71 21.0318
R15074 gnd.n5928 gnd.n5927 21.0318
R15075 gnd.n5855 gnd.n86 21.0318
R15076 gnd.n7723 gnd.n89 21.0318
R15077 gnd.n7717 gnd.n101 21.0318
R15078 gnd.n5870 gnd.n108 21.0318
R15079 gnd.n5913 gnd.n117 21.0318
R15080 gnd.n7705 gnd.n120 21.0318
R15081 gnd.n5907 gnd.n128 21.0318
R15082 gnd.n7699 gnd.n131 21.0318
R15083 gnd.n7693 gnd.n141 21.0318
R15084 gnd.n5895 gnd.n149 21.0318
R15085 gnd.n7687 gnd.n152 21.0318
R15086 gnd.n5889 gnd.n159 21.0318
R15087 gnd.n7668 gnd.n168 21.0318
R15088 gnd.n7675 gnd.n171 21.0318
R15089 gnd.n6154 gnd.n6153 20.7615
R15090 gnd.n5473 gnd.n5472 20.7615
R15091 gnd.t166 gnd.n1013 20.7131
R15092 gnd.n4301 gnd.t251 20.7131
R15093 gnd.t212 gnd.n2486 20.7131
R15094 gnd.t196 gnd.n5948 20.7131
R15095 gnd.n5861 gnd.t225 20.7131
R15096 gnd.n6274 gnd.n2676 20.3945
R15097 gnd.n3056 gnd.n3048 20.3945
R15098 gnd.t174 gnd.n1047 20.0758
R15099 gnd.n4238 gnd.t203 20.0758
R15100 gnd.t217 gnd.n2523 20.0758
R15101 gnd.t192 gnd.n3111 20.0758
R15102 gnd.n5901 gnd.t238 20.0758
R15103 gnd.n2895 gnd.t46 19.8005
R15104 gnd.n2895 gnd.t74 19.8005
R15105 gnd.n2894 gnd.t156 19.8005
R15106 gnd.n2894 gnd.t53 19.8005
R15107 gnd.n5399 gnd.t102 19.8005
R15108 gnd.n5399 gnd.t43 19.8005
R15109 gnd.n5398 gnd.t92 19.8005
R15110 gnd.n5398 gnd.t68 19.8005
R15111 gnd.n2891 gnd.n2890 19.5087
R15112 gnd.n2904 gnd.n2891 19.5087
R15113 gnd.n2902 gnd.n2893 19.5087
R15114 gnd.n5403 gnd.n5397 19.5087
R15115 gnd.n1766 gnd.t4 19.4385
R15116 gnd.n3836 gnd.n3833 19.3944
R15117 gnd.n3836 gnd.n3755 19.3944
R15118 gnd.n4487 gnd.n3755 19.3944
R15119 gnd.n4487 gnd.n3752 19.3944
R15120 gnd.n4497 gnd.n3752 19.3944
R15121 gnd.n4497 gnd.n3753 19.3944
R15122 gnd.n4493 gnd.n3753 19.3944
R15123 gnd.n4493 gnd.n4492 19.3944
R15124 gnd.n4492 gnd.n3731 19.3944
R15125 gnd.n4542 gnd.n3731 19.3944
R15126 gnd.n4543 gnd.n4542 19.3944
R15127 gnd.n4543 gnd.n3728 19.3944
R15128 gnd.n4552 gnd.n3728 19.3944
R15129 gnd.n4552 gnd.n3729 19.3944
R15130 gnd.n4548 gnd.n3729 19.3944
R15131 gnd.n4548 gnd.n4547 19.3944
R15132 gnd.n4547 gnd.n3699 19.3944
R15133 gnd.n4609 gnd.n3699 19.3944
R15134 gnd.n4609 gnd.n3696 19.3944
R15135 gnd.n4620 gnd.n3696 19.3944
R15136 gnd.n4620 gnd.n3697 19.3944
R15137 gnd.n4616 gnd.n3697 19.3944
R15138 gnd.n4616 gnd.n4615 19.3944
R15139 gnd.n4615 gnd.n3658 19.3944
R15140 gnd.n4697 gnd.n3658 19.3944
R15141 gnd.n4697 gnd.n3655 19.3944
R15142 gnd.n4737 gnd.n3655 19.3944
R15143 gnd.n4737 gnd.n3656 19.3944
R15144 gnd.n4733 gnd.n3656 19.3944
R15145 gnd.n4733 gnd.n4732 19.3944
R15146 gnd.n4732 gnd.n4731 19.3944
R15147 gnd.n4731 gnd.n4704 19.3944
R15148 gnd.n4727 gnd.n4704 19.3944
R15149 gnd.n4727 gnd.n4726 19.3944
R15150 gnd.n4726 gnd.n4725 19.3944
R15151 gnd.n4725 gnd.n4709 19.3944
R15152 gnd.n4721 gnd.n4709 19.3944
R15153 gnd.n4721 gnd.n4720 19.3944
R15154 gnd.n4720 gnd.n4719 19.3944
R15155 gnd.n4719 gnd.n4716 19.3944
R15156 gnd.n4716 gnd.n3571 19.3944
R15157 gnd.n4874 gnd.n3571 19.3944
R15158 gnd.n4874 gnd.n3568 19.3944
R15159 gnd.n4892 gnd.n3568 19.3944
R15160 gnd.n4892 gnd.n3569 19.3944
R15161 gnd.n4888 gnd.n3569 19.3944
R15162 gnd.n4888 gnd.n4887 19.3944
R15163 gnd.n4887 gnd.n4886 19.3944
R15164 gnd.n4886 gnd.n4883 19.3944
R15165 gnd.n4883 gnd.n3522 19.3944
R15166 gnd.n4961 gnd.n3522 19.3944
R15167 gnd.n4961 gnd.n3519 19.3944
R15168 gnd.n4969 gnd.n3519 19.3944
R15169 gnd.n4969 gnd.n3520 19.3944
R15170 gnd.n4965 gnd.n3520 19.3944
R15171 gnd.n4965 gnd.n3493 19.3944
R15172 gnd.n5029 gnd.n3493 19.3944
R15173 gnd.n5029 gnd.n3490 19.3944
R15174 gnd.n5047 gnd.n3490 19.3944
R15175 gnd.n5047 gnd.n3491 19.3944
R15176 gnd.n5043 gnd.n3491 19.3944
R15177 gnd.n5043 gnd.n5042 19.3944
R15178 gnd.n5042 gnd.n5041 19.3944
R15179 gnd.n5041 gnd.n5038 19.3944
R15180 gnd.n5038 gnd.n3418 19.3944
R15181 gnd.n5114 gnd.n3418 19.3944
R15182 gnd.n5114 gnd.n3415 19.3944
R15183 gnd.n5119 gnd.n3415 19.3944
R15184 gnd.n5119 gnd.n3416 19.3944
R15185 gnd.n3416 gnd.n3388 19.3944
R15186 gnd.n5150 gnd.n3388 19.3944
R15187 gnd.n5150 gnd.n3386 19.3944
R15188 gnd.n5154 gnd.n3386 19.3944
R15189 gnd.n5154 gnd.n3367 19.3944
R15190 gnd.n5181 gnd.n3367 19.3944
R15191 gnd.n5181 gnd.n3365 19.3944
R15192 gnd.n5185 gnd.n3365 19.3944
R15193 gnd.n5185 gnd.n3363 19.3944
R15194 gnd.n5191 gnd.n3363 19.3944
R15195 gnd.n5191 gnd.n3360 19.3944
R15196 gnd.n5374 gnd.n3360 19.3944
R15197 gnd.n5374 gnd.n3361 19.3944
R15198 gnd.n2668 gnd.n2584 19.3944
R15199 gnd.n6343 gnd.n2584 19.3944
R15200 gnd.n6343 gnd.n6342 19.3944
R15201 gnd.n6336 gnd.n6335 19.3944
R15202 gnd.n6335 gnd.n2606 19.3944
R15203 gnd.n6331 gnd.n2606 19.3944
R15204 gnd.n6331 gnd.n6330 19.3944
R15205 gnd.n6330 gnd.n6329 19.3944
R15206 gnd.n6329 gnd.n2611 19.3944
R15207 gnd.n6324 gnd.n2611 19.3944
R15208 gnd.n6324 gnd.n6323 19.3944
R15209 gnd.n6323 gnd.n6322 19.3944
R15210 gnd.n6322 gnd.n2617 19.3944
R15211 gnd.n6315 gnd.n2617 19.3944
R15212 gnd.n6315 gnd.n6314 19.3944
R15213 gnd.n6314 gnd.n2629 19.3944
R15214 gnd.n6307 gnd.n2629 19.3944
R15215 gnd.n6307 gnd.n6306 19.3944
R15216 gnd.n6306 gnd.n2637 19.3944
R15217 gnd.n6299 gnd.n2637 19.3944
R15218 gnd.n6299 gnd.n6298 19.3944
R15219 gnd.n6298 gnd.n2647 19.3944
R15220 gnd.n6291 gnd.n2647 19.3944
R15221 gnd.n6291 gnd.n6290 19.3944
R15222 gnd.n6290 gnd.n2655 19.3944
R15223 gnd.n6283 gnd.n2655 19.3944
R15224 gnd.n6283 gnd.n6282 19.3944
R15225 gnd.n5282 gnd.n5245 19.3944
R15226 gnd.n5295 gnd.n5245 19.3944
R15227 gnd.n5295 gnd.n5243 19.3944
R15228 gnd.n5301 gnd.n5243 19.3944
R15229 gnd.n5301 gnd.n5236 19.3944
R15230 gnd.n5314 gnd.n5236 19.3944
R15231 gnd.n5314 gnd.n5234 19.3944
R15232 gnd.n5320 gnd.n5234 19.3944
R15233 gnd.n5320 gnd.n5227 19.3944
R15234 gnd.n5333 gnd.n5227 19.3944
R15235 gnd.n5333 gnd.n5225 19.3944
R15236 gnd.n5339 gnd.n5225 19.3944
R15237 gnd.n5339 gnd.n5218 19.3944
R15238 gnd.n5353 gnd.n5218 19.3944
R15239 gnd.n5353 gnd.n5216 19.3944
R15240 gnd.n5359 gnd.n5216 19.3944
R15241 gnd.n1481 gnd.n1480 19.3944
R15242 gnd.n1480 gnd.n1479 19.3944
R15243 gnd.n1479 gnd.n1478 19.3944
R15244 gnd.n1478 gnd.n1476 19.3944
R15245 gnd.n1476 gnd.n1473 19.3944
R15246 gnd.n1473 gnd.n1472 19.3944
R15247 gnd.n1472 gnd.n1469 19.3944
R15248 gnd.n1469 gnd.n1468 19.3944
R15249 gnd.n1468 gnd.n1465 19.3944
R15250 gnd.n1465 gnd.n1464 19.3944
R15251 gnd.n1464 gnd.n1461 19.3944
R15252 gnd.n1461 gnd.n1460 19.3944
R15253 gnd.n1460 gnd.n1457 19.3944
R15254 gnd.n1457 gnd.n1456 19.3944
R15255 gnd.n1456 gnd.n1453 19.3944
R15256 gnd.n1453 gnd.n1452 19.3944
R15257 gnd.n1452 gnd.n1449 19.3944
R15258 gnd.n1449 gnd.n1448 19.3944
R15259 gnd.n1448 gnd.n1445 19.3944
R15260 gnd.n1445 gnd.n1444 19.3944
R15261 gnd.n1444 gnd.n1441 19.3944
R15262 gnd.n1441 gnd.n1440 19.3944
R15263 gnd.n1437 gnd.n1436 19.3944
R15264 gnd.n1436 gnd.n1392 19.3944
R15265 gnd.n1487 gnd.n1392 19.3944
R15266 gnd.n2255 gnd.n2254 19.3944
R15267 gnd.n2254 gnd.n2251 19.3944
R15268 gnd.n2251 gnd.n2250 19.3944
R15269 gnd.n2300 gnd.n2299 19.3944
R15270 gnd.n2299 gnd.n2298 19.3944
R15271 gnd.n2298 gnd.n2295 19.3944
R15272 gnd.n2295 gnd.n2294 19.3944
R15273 gnd.n2294 gnd.n2291 19.3944
R15274 gnd.n2291 gnd.n2290 19.3944
R15275 gnd.n2290 gnd.n2287 19.3944
R15276 gnd.n2287 gnd.n2286 19.3944
R15277 gnd.n2286 gnd.n2283 19.3944
R15278 gnd.n2283 gnd.n2282 19.3944
R15279 gnd.n2282 gnd.n2279 19.3944
R15280 gnd.n2279 gnd.n2278 19.3944
R15281 gnd.n2278 gnd.n2275 19.3944
R15282 gnd.n2275 gnd.n2274 19.3944
R15283 gnd.n2274 gnd.n2271 19.3944
R15284 gnd.n2271 gnd.n2270 19.3944
R15285 gnd.n2270 gnd.n2267 19.3944
R15286 gnd.n2267 gnd.n2266 19.3944
R15287 gnd.n2266 gnd.n2263 19.3944
R15288 gnd.n2263 gnd.n2262 19.3944
R15289 gnd.n2262 gnd.n2259 19.3944
R15290 gnd.n2259 gnd.n2258 19.3944
R15291 gnd.n1580 gnd.n1289 19.3944
R15292 gnd.n1590 gnd.n1289 19.3944
R15293 gnd.n1591 gnd.n1590 19.3944
R15294 gnd.n1591 gnd.n1270 19.3944
R15295 gnd.n1611 gnd.n1270 19.3944
R15296 gnd.n1611 gnd.n1262 19.3944
R15297 gnd.n1621 gnd.n1262 19.3944
R15298 gnd.n1622 gnd.n1621 19.3944
R15299 gnd.n1623 gnd.n1622 19.3944
R15300 gnd.n1623 gnd.n1245 19.3944
R15301 gnd.n1640 gnd.n1245 19.3944
R15302 gnd.n1643 gnd.n1640 19.3944
R15303 gnd.n1643 gnd.n1642 19.3944
R15304 gnd.n1642 gnd.n1218 19.3944
R15305 gnd.n1682 gnd.n1218 19.3944
R15306 gnd.n1682 gnd.n1215 19.3944
R15307 gnd.n1688 gnd.n1215 19.3944
R15308 gnd.n1689 gnd.n1688 19.3944
R15309 gnd.n1689 gnd.n1213 19.3944
R15310 gnd.n1695 gnd.n1213 19.3944
R15311 gnd.n1698 gnd.n1695 19.3944
R15312 gnd.n1700 gnd.n1698 19.3944
R15313 gnd.n1706 gnd.n1700 19.3944
R15314 gnd.n1706 gnd.n1705 19.3944
R15315 gnd.n1705 gnd.n1088 19.3944
R15316 gnd.n1772 gnd.n1088 19.3944
R15317 gnd.n1773 gnd.n1772 19.3944
R15318 gnd.n1773 gnd.n1081 19.3944
R15319 gnd.n1784 gnd.n1081 19.3944
R15320 gnd.n1785 gnd.n1784 19.3944
R15321 gnd.n1785 gnd.n1064 19.3944
R15322 gnd.n1064 gnd.n1062 19.3944
R15323 gnd.n1809 gnd.n1062 19.3944
R15324 gnd.n1810 gnd.n1809 19.3944
R15325 gnd.n1810 gnd.n1035 19.3944
R15326 gnd.n1859 gnd.n1035 19.3944
R15327 gnd.n1860 gnd.n1859 19.3944
R15328 gnd.n1860 gnd.n1028 19.3944
R15329 gnd.n1871 gnd.n1028 19.3944
R15330 gnd.n1872 gnd.n1871 19.3944
R15331 gnd.n1872 gnd.n1011 19.3944
R15332 gnd.n1011 gnd.n1009 19.3944
R15333 gnd.n1896 gnd.n1009 19.3944
R15334 gnd.n1897 gnd.n1896 19.3944
R15335 gnd.n1897 gnd.n981 19.3944
R15336 gnd.n1948 gnd.n981 19.3944
R15337 gnd.n1949 gnd.n1948 19.3944
R15338 gnd.n1949 gnd.n974 19.3944
R15339 gnd.n2216 gnd.n974 19.3944
R15340 gnd.n2217 gnd.n2216 19.3944
R15341 gnd.n2217 gnd.n955 19.3944
R15342 gnd.n2242 gnd.n955 19.3944
R15343 gnd.n2242 gnd.n956 19.3944
R15344 gnd.n1571 gnd.n1570 19.3944
R15345 gnd.n1570 gnd.n1303 19.3944
R15346 gnd.n1326 gnd.n1303 19.3944
R15347 gnd.n1329 gnd.n1326 19.3944
R15348 gnd.n1329 gnd.n1322 19.3944
R15349 gnd.n1333 gnd.n1322 19.3944
R15350 gnd.n1336 gnd.n1333 19.3944
R15351 gnd.n1339 gnd.n1336 19.3944
R15352 gnd.n1339 gnd.n1320 19.3944
R15353 gnd.n1343 gnd.n1320 19.3944
R15354 gnd.n1346 gnd.n1343 19.3944
R15355 gnd.n1349 gnd.n1346 19.3944
R15356 gnd.n1349 gnd.n1318 19.3944
R15357 gnd.n1353 gnd.n1318 19.3944
R15358 gnd.n1576 gnd.n1575 19.3944
R15359 gnd.n1575 gnd.n1279 19.3944
R15360 gnd.n1601 gnd.n1279 19.3944
R15361 gnd.n1601 gnd.n1277 19.3944
R15362 gnd.n1607 gnd.n1277 19.3944
R15363 gnd.n1607 gnd.n1606 19.3944
R15364 gnd.n1606 gnd.n1251 19.3944
R15365 gnd.n1631 gnd.n1251 19.3944
R15366 gnd.n1631 gnd.n1249 19.3944
R15367 gnd.n1635 gnd.n1249 19.3944
R15368 gnd.n1635 gnd.n1229 19.3944
R15369 gnd.n1662 gnd.n1229 19.3944
R15370 gnd.n1662 gnd.n1227 19.3944
R15371 gnd.n1672 gnd.n1227 19.3944
R15372 gnd.n1672 gnd.n1671 19.3944
R15373 gnd.n1671 gnd.n1670 19.3944
R15374 gnd.n1670 gnd.n1176 19.3944
R15375 gnd.n1720 gnd.n1176 19.3944
R15376 gnd.n1720 gnd.n1719 19.3944
R15377 gnd.n1719 gnd.n1718 19.3944
R15378 gnd.n1718 gnd.n1180 19.3944
R15379 gnd.n1200 gnd.n1180 19.3944
R15380 gnd.n1200 gnd.n1098 19.3944
R15381 gnd.n1757 gnd.n1098 19.3944
R15382 gnd.n1757 gnd.n1096 19.3944
R15383 gnd.n1763 gnd.n1096 19.3944
R15384 gnd.n1763 gnd.n1762 19.3944
R15385 gnd.n1762 gnd.n1071 19.3944
R15386 gnd.n1797 gnd.n1071 19.3944
R15387 gnd.n1797 gnd.n1069 19.3944
R15388 gnd.n1803 gnd.n1069 19.3944
R15389 gnd.n1803 gnd.n1802 19.3944
R15390 gnd.n1802 gnd.n1045 19.3944
R15391 gnd.n1844 gnd.n1045 19.3944
R15392 gnd.n1844 gnd.n1043 19.3944
R15393 gnd.n1850 gnd.n1043 19.3944
R15394 gnd.n1850 gnd.n1849 19.3944
R15395 gnd.n1849 gnd.n1018 19.3944
R15396 gnd.n1884 gnd.n1018 19.3944
R15397 gnd.n1884 gnd.n1016 19.3944
R15398 gnd.n1890 gnd.n1016 19.3944
R15399 gnd.n1890 gnd.n1889 19.3944
R15400 gnd.n1889 gnd.n991 19.3944
R15401 gnd.n1933 gnd.n991 19.3944
R15402 gnd.n1933 gnd.n989 19.3944
R15403 gnd.n1939 gnd.n989 19.3944
R15404 gnd.n1939 gnd.n1938 19.3944
R15405 gnd.n1938 gnd.n964 19.3944
R15406 gnd.n2227 gnd.n964 19.3944
R15407 gnd.n2227 gnd.n962 19.3944
R15408 gnd.n2235 gnd.n962 19.3944
R15409 gnd.n2235 gnd.n2234 19.3944
R15410 gnd.n2234 gnd.n2233 19.3944
R15411 gnd.n2336 gnd.n2335 19.3944
R15412 gnd.n2335 gnd.n903 19.3944
R15413 gnd.n2331 gnd.n903 19.3944
R15414 gnd.n2331 gnd.n2328 19.3944
R15415 gnd.n2328 gnd.n2325 19.3944
R15416 gnd.n2325 gnd.n2324 19.3944
R15417 gnd.n2324 gnd.n2321 19.3944
R15418 gnd.n2321 gnd.n2320 19.3944
R15419 gnd.n2320 gnd.n2317 19.3944
R15420 gnd.n2317 gnd.n2316 19.3944
R15421 gnd.n2316 gnd.n2313 19.3944
R15422 gnd.n2313 gnd.n2312 19.3944
R15423 gnd.n2312 gnd.n2309 19.3944
R15424 gnd.n2309 gnd.n2308 19.3944
R15425 gnd.n1491 gnd.n1390 19.3944
R15426 gnd.n1491 gnd.n1381 19.3944
R15427 gnd.n1504 gnd.n1381 19.3944
R15428 gnd.n1504 gnd.n1379 19.3944
R15429 gnd.n1508 gnd.n1379 19.3944
R15430 gnd.n1508 gnd.n1369 19.3944
R15431 gnd.n1520 gnd.n1369 19.3944
R15432 gnd.n1520 gnd.n1367 19.3944
R15433 gnd.n1554 gnd.n1367 19.3944
R15434 gnd.n1554 gnd.n1553 19.3944
R15435 gnd.n1553 gnd.n1552 19.3944
R15436 gnd.n1552 gnd.n1551 19.3944
R15437 gnd.n1551 gnd.n1548 19.3944
R15438 gnd.n1548 gnd.n1547 19.3944
R15439 gnd.n1547 gnd.n1546 19.3944
R15440 gnd.n1546 gnd.n1544 19.3944
R15441 gnd.n1544 gnd.n1543 19.3944
R15442 gnd.n1543 gnd.n1540 19.3944
R15443 gnd.n1540 gnd.n1539 19.3944
R15444 gnd.n1539 gnd.n1538 19.3944
R15445 gnd.n1538 gnd.n1536 19.3944
R15446 gnd.n1536 gnd.n1235 19.3944
R15447 gnd.n1651 gnd.n1235 19.3944
R15448 gnd.n1651 gnd.n1233 19.3944
R15449 gnd.n1657 gnd.n1233 19.3944
R15450 gnd.n1657 gnd.n1656 19.3944
R15451 gnd.n1656 gnd.n1157 19.3944
R15452 gnd.n1731 gnd.n1157 19.3944
R15453 gnd.n1731 gnd.n1158 19.3944
R15454 gnd.n1205 gnd.n1204 19.3944
R15455 gnd.n1208 gnd.n1207 19.3944
R15456 gnd.n1195 gnd.n1194 19.3944
R15457 gnd.n1750 gnd.n1103 19.3944
R15458 gnd.n1750 gnd.n1749 19.3944
R15459 gnd.n1749 gnd.n1748 19.3944
R15460 gnd.n1748 gnd.n1746 19.3944
R15461 gnd.n1746 gnd.n1745 19.3944
R15462 gnd.n1745 gnd.n1743 19.3944
R15463 gnd.n1743 gnd.n1742 19.3944
R15464 gnd.n1742 gnd.n1052 19.3944
R15465 gnd.n1818 gnd.n1052 19.3944
R15466 gnd.n1818 gnd.n1050 19.3944
R15467 gnd.n1837 gnd.n1050 19.3944
R15468 gnd.n1837 gnd.n1836 19.3944
R15469 gnd.n1836 gnd.n1835 19.3944
R15470 gnd.n1835 gnd.n1833 19.3944
R15471 gnd.n1833 gnd.n1832 19.3944
R15472 gnd.n1832 gnd.n1830 19.3944
R15473 gnd.n1830 gnd.n1829 19.3944
R15474 gnd.n1829 gnd.n998 19.3944
R15475 gnd.n1905 gnd.n998 19.3944
R15476 gnd.n1905 gnd.n996 19.3944
R15477 gnd.n1928 gnd.n996 19.3944
R15478 gnd.n1928 gnd.n1927 19.3944
R15479 gnd.n1927 gnd.n1926 19.3944
R15480 gnd.n1926 gnd.n1923 19.3944
R15481 gnd.n1923 gnd.n1922 19.3944
R15482 gnd.n1922 gnd.n1920 19.3944
R15483 gnd.n1920 gnd.n1919 19.3944
R15484 gnd.n1919 gnd.n1917 19.3944
R15485 gnd.n1917 gnd.n950 19.3944
R15486 gnd.n1496 gnd.n1386 19.3944
R15487 gnd.n1496 gnd.n1384 19.3944
R15488 gnd.n1500 gnd.n1384 19.3944
R15489 gnd.n1500 gnd.n1375 19.3944
R15490 gnd.n1512 gnd.n1375 19.3944
R15491 gnd.n1512 gnd.n1373 19.3944
R15492 gnd.n1516 gnd.n1373 19.3944
R15493 gnd.n1516 gnd.n1362 19.3944
R15494 gnd.n1558 gnd.n1362 19.3944
R15495 gnd.n1558 gnd.n1316 19.3944
R15496 gnd.n1564 gnd.n1316 19.3944
R15497 gnd.n1564 gnd.n1563 19.3944
R15498 gnd.n1563 gnd.n1294 19.3944
R15499 gnd.n1585 gnd.n1294 19.3944
R15500 gnd.n1585 gnd.n1287 19.3944
R15501 gnd.n1596 gnd.n1287 19.3944
R15502 gnd.n1596 gnd.n1595 19.3944
R15503 gnd.n1595 gnd.n1268 19.3944
R15504 gnd.n1616 gnd.n1268 19.3944
R15505 gnd.n1616 gnd.n1258 19.3944
R15506 gnd.n1626 gnd.n1258 19.3944
R15507 gnd.n1626 gnd.n1241 19.3944
R15508 gnd.n1647 gnd.n1241 19.3944
R15509 gnd.n1647 gnd.n1646 19.3944
R15510 gnd.n1646 gnd.n1220 19.3944
R15511 gnd.n1677 gnd.n1220 19.3944
R15512 gnd.n1677 gnd.n1165 19.3944
R15513 gnd.n1727 gnd.n1165 19.3944
R15514 gnd.n1727 gnd.n1726 19.3944
R15515 gnd.n1726 gnd.n1725 19.3944
R15516 gnd.n1725 gnd.n1169 19.3944
R15517 gnd.n1187 gnd.n1169 19.3944
R15518 gnd.n1713 gnd.n1187 19.3944
R15519 gnd.n1713 gnd.n1712 19.3944
R15520 gnd.n1712 gnd.n1711 19.3944
R15521 gnd.n1711 gnd.n1191 19.3944
R15522 gnd.n1191 gnd.n1090 19.3944
R15523 gnd.n1768 gnd.n1090 19.3944
R15524 gnd.n1768 gnd.n1083 19.3944
R15525 gnd.n1779 gnd.n1083 19.3944
R15526 gnd.n1779 gnd.n1079 19.3944
R15527 gnd.n1792 gnd.n1079 19.3944
R15528 gnd.n1792 gnd.n1791 19.3944
R15529 gnd.n1791 gnd.n1058 19.3944
R15530 gnd.n1814 gnd.n1058 19.3944
R15531 gnd.n1814 gnd.n1813 19.3944
R15532 gnd.n1813 gnd.n1037 19.3944
R15533 gnd.n1855 gnd.n1037 19.3944
R15534 gnd.n1855 gnd.n1030 19.3944
R15535 gnd.n1866 gnd.n1030 19.3944
R15536 gnd.n1866 gnd.n1026 19.3944
R15537 gnd.n1879 gnd.n1026 19.3944
R15538 gnd.n1879 gnd.n1878 19.3944
R15539 gnd.n1878 gnd.n1005 19.3944
R15540 gnd.n1901 gnd.n1005 19.3944
R15541 gnd.n1901 gnd.n1900 19.3944
R15542 gnd.n1900 gnd.n983 19.3944
R15543 gnd.n1944 gnd.n983 19.3944
R15544 gnd.n1944 gnd.n976 19.3944
R15545 gnd.n1955 gnd.n976 19.3944
R15546 gnd.n1955 gnd.n972 19.3944
R15547 gnd.n2222 gnd.n972 19.3944
R15548 gnd.n2222 gnd.n2221 19.3944
R15549 gnd.n2221 gnd.n953 19.3944
R15550 gnd.n2245 gnd.n953 19.3944
R15551 gnd.n6319 gnd.n2620 19.3944
R15552 gnd.n6319 gnd.n6318 19.3944
R15553 gnd.n6318 gnd.n2623 19.3944
R15554 gnd.n6311 gnd.n2623 19.3944
R15555 gnd.n6311 gnd.n6310 19.3944
R15556 gnd.n6310 gnd.n2633 19.3944
R15557 gnd.n6303 gnd.n2633 19.3944
R15558 gnd.n6303 gnd.n6302 19.3944
R15559 gnd.n6302 gnd.n2641 19.3944
R15560 gnd.n6295 gnd.n2641 19.3944
R15561 gnd.n6295 gnd.n6294 19.3944
R15562 gnd.n6294 gnd.n2651 19.3944
R15563 gnd.n6287 gnd.n2651 19.3944
R15564 gnd.n6287 gnd.n6286 19.3944
R15565 gnd.n6286 gnd.n2659 19.3944
R15566 gnd.n6279 gnd.n2659 19.3944
R15567 gnd.n7209 gnd.n392 19.3944
R15568 gnd.n7215 gnd.n392 19.3944
R15569 gnd.n7215 gnd.n390 19.3944
R15570 gnd.n7219 gnd.n390 19.3944
R15571 gnd.n7219 gnd.n386 19.3944
R15572 gnd.n7225 gnd.n386 19.3944
R15573 gnd.n7225 gnd.n384 19.3944
R15574 gnd.n7229 gnd.n384 19.3944
R15575 gnd.n7229 gnd.n380 19.3944
R15576 gnd.n7235 gnd.n380 19.3944
R15577 gnd.n7235 gnd.n378 19.3944
R15578 gnd.n7239 gnd.n378 19.3944
R15579 gnd.n7239 gnd.n374 19.3944
R15580 gnd.n7245 gnd.n374 19.3944
R15581 gnd.n7245 gnd.n372 19.3944
R15582 gnd.n7249 gnd.n372 19.3944
R15583 gnd.n7249 gnd.n368 19.3944
R15584 gnd.n7255 gnd.n368 19.3944
R15585 gnd.n7255 gnd.n366 19.3944
R15586 gnd.n7259 gnd.n366 19.3944
R15587 gnd.n7259 gnd.n362 19.3944
R15588 gnd.n7265 gnd.n362 19.3944
R15589 gnd.n7265 gnd.n360 19.3944
R15590 gnd.n7269 gnd.n360 19.3944
R15591 gnd.n7269 gnd.n356 19.3944
R15592 gnd.n7275 gnd.n356 19.3944
R15593 gnd.n7275 gnd.n354 19.3944
R15594 gnd.n7279 gnd.n354 19.3944
R15595 gnd.n7279 gnd.n350 19.3944
R15596 gnd.n7285 gnd.n350 19.3944
R15597 gnd.n7285 gnd.n348 19.3944
R15598 gnd.n7289 gnd.n348 19.3944
R15599 gnd.n7289 gnd.n344 19.3944
R15600 gnd.n7295 gnd.n344 19.3944
R15601 gnd.n7295 gnd.n342 19.3944
R15602 gnd.n7299 gnd.n342 19.3944
R15603 gnd.n7299 gnd.n338 19.3944
R15604 gnd.n7305 gnd.n338 19.3944
R15605 gnd.n7305 gnd.n336 19.3944
R15606 gnd.n7309 gnd.n336 19.3944
R15607 gnd.n7309 gnd.n332 19.3944
R15608 gnd.n7315 gnd.n332 19.3944
R15609 gnd.n7315 gnd.n330 19.3944
R15610 gnd.n7319 gnd.n330 19.3944
R15611 gnd.n7319 gnd.n326 19.3944
R15612 gnd.n7325 gnd.n326 19.3944
R15613 gnd.n7325 gnd.n324 19.3944
R15614 gnd.n7329 gnd.n324 19.3944
R15615 gnd.n7329 gnd.n320 19.3944
R15616 gnd.n7335 gnd.n320 19.3944
R15617 gnd.n7335 gnd.n318 19.3944
R15618 gnd.n7339 gnd.n318 19.3944
R15619 gnd.n7339 gnd.n314 19.3944
R15620 gnd.n7345 gnd.n314 19.3944
R15621 gnd.n7345 gnd.n312 19.3944
R15622 gnd.n7349 gnd.n312 19.3944
R15623 gnd.n7349 gnd.n308 19.3944
R15624 gnd.n7355 gnd.n308 19.3944
R15625 gnd.n7355 gnd.n306 19.3944
R15626 gnd.n7359 gnd.n306 19.3944
R15627 gnd.n7359 gnd.n302 19.3944
R15628 gnd.n7365 gnd.n302 19.3944
R15629 gnd.n7365 gnd.n300 19.3944
R15630 gnd.n7369 gnd.n300 19.3944
R15631 gnd.n7369 gnd.n296 19.3944
R15632 gnd.n7375 gnd.n296 19.3944
R15633 gnd.n7375 gnd.n294 19.3944
R15634 gnd.n7379 gnd.n294 19.3944
R15635 gnd.n7379 gnd.n290 19.3944
R15636 gnd.n7385 gnd.n290 19.3944
R15637 gnd.n7385 gnd.n288 19.3944
R15638 gnd.n7389 gnd.n288 19.3944
R15639 gnd.n7389 gnd.n284 19.3944
R15640 gnd.n7395 gnd.n284 19.3944
R15641 gnd.n7395 gnd.n282 19.3944
R15642 gnd.n7399 gnd.n282 19.3944
R15643 gnd.n7399 gnd.n278 19.3944
R15644 gnd.n7405 gnd.n278 19.3944
R15645 gnd.n7405 gnd.n276 19.3944
R15646 gnd.n7409 gnd.n276 19.3944
R15647 gnd.n7409 gnd.n272 19.3944
R15648 gnd.n7415 gnd.n272 19.3944
R15649 gnd.n7415 gnd.n270 19.3944
R15650 gnd.n7420 gnd.n270 19.3944
R15651 gnd.n6688 gnd.n703 19.3944
R15652 gnd.n6694 gnd.n703 19.3944
R15653 gnd.n6694 gnd.n701 19.3944
R15654 gnd.n6698 gnd.n701 19.3944
R15655 gnd.n6698 gnd.n697 19.3944
R15656 gnd.n6704 gnd.n697 19.3944
R15657 gnd.n6704 gnd.n695 19.3944
R15658 gnd.n6708 gnd.n695 19.3944
R15659 gnd.n6708 gnd.n691 19.3944
R15660 gnd.n6714 gnd.n691 19.3944
R15661 gnd.n6714 gnd.n689 19.3944
R15662 gnd.n6718 gnd.n689 19.3944
R15663 gnd.n6718 gnd.n685 19.3944
R15664 gnd.n6724 gnd.n685 19.3944
R15665 gnd.n6724 gnd.n683 19.3944
R15666 gnd.n6728 gnd.n683 19.3944
R15667 gnd.n6728 gnd.n679 19.3944
R15668 gnd.n6734 gnd.n679 19.3944
R15669 gnd.n6734 gnd.n677 19.3944
R15670 gnd.n6738 gnd.n677 19.3944
R15671 gnd.n6738 gnd.n673 19.3944
R15672 gnd.n6744 gnd.n673 19.3944
R15673 gnd.n6744 gnd.n671 19.3944
R15674 gnd.n6748 gnd.n671 19.3944
R15675 gnd.n6748 gnd.n667 19.3944
R15676 gnd.n6754 gnd.n667 19.3944
R15677 gnd.n6754 gnd.n665 19.3944
R15678 gnd.n6758 gnd.n665 19.3944
R15679 gnd.n6758 gnd.n661 19.3944
R15680 gnd.n6764 gnd.n661 19.3944
R15681 gnd.n6764 gnd.n659 19.3944
R15682 gnd.n6768 gnd.n659 19.3944
R15683 gnd.n6768 gnd.n655 19.3944
R15684 gnd.n6774 gnd.n655 19.3944
R15685 gnd.n6774 gnd.n653 19.3944
R15686 gnd.n6778 gnd.n653 19.3944
R15687 gnd.n6778 gnd.n649 19.3944
R15688 gnd.n6784 gnd.n649 19.3944
R15689 gnd.n6784 gnd.n647 19.3944
R15690 gnd.n6788 gnd.n647 19.3944
R15691 gnd.n6788 gnd.n643 19.3944
R15692 gnd.n6794 gnd.n643 19.3944
R15693 gnd.n6794 gnd.n641 19.3944
R15694 gnd.n6798 gnd.n641 19.3944
R15695 gnd.n6798 gnd.n637 19.3944
R15696 gnd.n6804 gnd.n637 19.3944
R15697 gnd.n6804 gnd.n635 19.3944
R15698 gnd.n6808 gnd.n635 19.3944
R15699 gnd.n6808 gnd.n631 19.3944
R15700 gnd.n6814 gnd.n631 19.3944
R15701 gnd.n6814 gnd.n629 19.3944
R15702 gnd.n6818 gnd.n629 19.3944
R15703 gnd.n6818 gnd.n625 19.3944
R15704 gnd.n6824 gnd.n625 19.3944
R15705 gnd.n6824 gnd.n623 19.3944
R15706 gnd.n6828 gnd.n623 19.3944
R15707 gnd.n6828 gnd.n619 19.3944
R15708 gnd.n6834 gnd.n619 19.3944
R15709 gnd.n6834 gnd.n617 19.3944
R15710 gnd.n6838 gnd.n617 19.3944
R15711 gnd.n6838 gnd.n613 19.3944
R15712 gnd.n6844 gnd.n613 19.3944
R15713 gnd.n6844 gnd.n611 19.3944
R15714 gnd.n6848 gnd.n611 19.3944
R15715 gnd.n6848 gnd.n607 19.3944
R15716 gnd.n6854 gnd.n607 19.3944
R15717 gnd.n6854 gnd.n605 19.3944
R15718 gnd.n6858 gnd.n605 19.3944
R15719 gnd.n6858 gnd.n601 19.3944
R15720 gnd.n6864 gnd.n601 19.3944
R15721 gnd.n6864 gnd.n599 19.3944
R15722 gnd.n6868 gnd.n599 19.3944
R15723 gnd.n6868 gnd.n595 19.3944
R15724 gnd.n6874 gnd.n595 19.3944
R15725 gnd.n6874 gnd.n593 19.3944
R15726 gnd.n6878 gnd.n593 19.3944
R15727 gnd.n6878 gnd.n589 19.3944
R15728 gnd.n6884 gnd.n589 19.3944
R15729 gnd.n6884 gnd.n587 19.3944
R15730 gnd.n6888 gnd.n587 19.3944
R15731 gnd.n6888 gnd.n583 19.3944
R15732 gnd.n6894 gnd.n583 19.3944
R15733 gnd.n6894 gnd.n581 19.3944
R15734 gnd.n6898 gnd.n581 19.3944
R15735 gnd.n6898 gnd.n577 19.3944
R15736 gnd.n6904 gnd.n577 19.3944
R15737 gnd.n6904 gnd.n575 19.3944
R15738 gnd.n6908 gnd.n575 19.3944
R15739 gnd.n6908 gnd.n571 19.3944
R15740 gnd.n6914 gnd.n571 19.3944
R15741 gnd.n6914 gnd.n569 19.3944
R15742 gnd.n6918 gnd.n569 19.3944
R15743 gnd.n6918 gnd.n565 19.3944
R15744 gnd.n6924 gnd.n565 19.3944
R15745 gnd.n6924 gnd.n563 19.3944
R15746 gnd.n6928 gnd.n563 19.3944
R15747 gnd.n6928 gnd.n559 19.3944
R15748 gnd.n6934 gnd.n559 19.3944
R15749 gnd.n6934 gnd.n557 19.3944
R15750 gnd.n6938 gnd.n557 19.3944
R15751 gnd.n6938 gnd.n553 19.3944
R15752 gnd.n6944 gnd.n553 19.3944
R15753 gnd.n6944 gnd.n551 19.3944
R15754 gnd.n6948 gnd.n551 19.3944
R15755 gnd.n6948 gnd.n547 19.3944
R15756 gnd.n6954 gnd.n547 19.3944
R15757 gnd.n6954 gnd.n545 19.3944
R15758 gnd.n6958 gnd.n545 19.3944
R15759 gnd.n6958 gnd.n541 19.3944
R15760 gnd.n6964 gnd.n541 19.3944
R15761 gnd.n6964 gnd.n539 19.3944
R15762 gnd.n6968 gnd.n539 19.3944
R15763 gnd.n6968 gnd.n535 19.3944
R15764 gnd.n6974 gnd.n535 19.3944
R15765 gnd.n6974 gnd.n533 19.3944
R15766 gnd.n6978 gnd.n533 19.3944
R15767 gnd.n6978 gnd.n529 19.3944
R15768 gnd.n6984 gnd.n529 19.3944
R15769 gnd.n6984 gnd.n527 19.3944
R15770 gnd.n6988 gnd.n527 19.3944
R15771 gnd.n6988 gnd.n523 19.3944
R15772 gnd.n6994 gnd.n523 19.3944
R15773 gnd.n6994 gnd.n521 19.3944
R15774 gnd.n6998 gnd.n521 19.3944
R15775 gnd.n6998 gnd.n517 19.3944
R15776 gnd.n7004 gnd.n517 19.3944
R15777 gnd.n7004 gnd.n515 19.3944
R15778 gnd.n7008 gnd.n515 19.3944
R15779 gnd.n7008 gnd.n511 19.3944
R15780 gnd.n7014 gnd.n511 19.3944
R15781 gnd.n7014 gnd.n509 19.3944
R15782 gnd.n7018 gnd.n509 19.3944
R15783 gnd.n7018 gnd.n505 19.3944
R15784 gnd.n7024 gnd.n505 19.3944
R15785 gnd.n7024 gnd.n503 19.3944
R15786 gnd.n7028 gnd.n503 19.3944
R15787 gnd.n7028 gnd.n499 19.3944
R15788 gnd.n7034 gnd.n499 19.3944
R15789 gnd.n7034 gnd.n497 19.3944
R15790 gnd.n7038 gnd.n497 19.3944
R15791 gnd.n7038 gnd.n493 19.3944
R15792 gnd.n7044 gnd.n493 19.3944
R15793 gnd.n7044 gnd.n491 19.3944
R15794 gnd.n7048 gnd.n491 19.3944
R15795 gnd.n7048 gnd.n487 19.3944
R15796 gnd.n7054 gnd.n487 19.3944
R15797 gnd.n7054 gnd.n485 19.3944
R15798 gnd.n7058 gnd.n485 19.3944
R15799 gnd.n7058 gnd.n481 19.3944
R15800 gnd.n7064 gnd.n481 19.3944
R15801 gnd.n7064 gnd.n479 19.3944
R15802 gnd.n7068 gnd.n479 19.3944
R15803 gnd.n7068 gnd.n475 19.3944
R15804 gnd.n7074 gnd.n475 19.3944
R15805 gnd.n7074 gnd.n473 19.3944
R15806 gnd.n7078 gnd.n473 19.3944
R15807 gnd.n7078 gnd.n469 19.3944
R15808 gnd.n7084 gnd.n469 19.3944
R15809 gnd.n7084 gnd.n467 19.3944
R15810 gnd.n7088 gnd.n467 19.3944
R15811 gnd.n7088 gnd.n463 19.3944
R15812 gnd.n7094 gnd.n463 19.3944
R15813 gnd.n7094 gnd.n461 19.3944
R15814 gnd.n7098 gnd.n461 19.3944
R15815 gnd.n7098 gnd.n457 19.3944
R15816 gnd.n7104 gnd.n457 19.3944
R15817 gnd.n7104 gnd.n455 19.3944
R15818 gnd.n7108 gnd.n455 19.3944
R15819 gnd.n7108 gnd.n451 19.3944
R15820 gnd.n7114 gnd.n451 19.3944
R15821 gnd.n7114 gnd.n449 19.3944
R15822 gnd.n7118 gnd.n449 19.3944
R15823 gnd.n7118 gnd.n445 19.3944
R15824 gnd.n7124 gnd.n445 19.3944
R15825 gnd.n7124 gnd.n443 19.3944
R15826 gnd.n7128 gnd.n443 19.3944
R15827 gnd.n7128 gnd.n439 19.3944
R15828 gnd.n7134 gnd.n439 19.3944
R15829 gnd.n7134 gnd.n437 19.3944
R15830 gnd.n7138 gnd.n437 19.3944
R15831 gnd.n7138 gnd.n433 19.3944
R15832 gnd.n7144 gnd.n433 19.3944
R15833 gnd.n7144 gnd.n431 19.3944
R15834 gnd.n7148 gnd.n431 19.3944
R15835 gnd.n7148 gnd.n427 19.3944
R15836 gnd.n7154 gnd.n427 19.3944
R15837 gnd.n7154 gnd.n425 19.3944
R15838 gnd.n7158 gnd.n425 19.3944
R15839 gnd.n7158 gnd.n421 19.3944
R15840 gnd.n7164 gnd.n421 19.3944
R15841 gnd.n7164 gnd.n419 19.3944
R15842 gnd.n7168 gnd.n419 19.3944
R15843 gnd.n7168 gnd.n415 19.3944
R15844 gnd.n7174 gnd.n415 19.3944
R15845 gnd.n7174 gnd.n413 19.3944
R15846 gnd.n7178 gnd.n413 19.3944
R15847 gnd.n7178 gnd.n409 19.3944
R15848 gnd.n7184 gnd.n409 19.3944
R15849 gnd.n7184 gnd.n407 19.3944
R15850 gnd.n7188 gnd.n407 19.3944
R15851 gnd.n7188 gnd.n403 19.3944
R15852 gnd.n7194 gnd.n403 19.3944
R15853 gnd.n7194 gnd.n401 19.3944
R15854 gnd.n7199 gnd.n401 19.3944
R15855 gnd.n7199 gnd.n397 19.3944
R15856 gnd.n7205 gnd.n397 19.3944
R15857 gnd.n7206 gnd.n7205 19.3944
R15858 gnd.n5574 gnd.n5571 19.3944
R15859 gnd.n5574 gnd.n5570 19.3944
R15860 gnd.n5580 gnd.n5570 19.3944
R15861 gnd.n5580 gnd.n5568 19.3944
R15862 gnd.n5584 gnd.n5568 19.3944
R15863 gnd.n5584 gnd.n5566 19.3944
R15864 gnd.n5590 gnd.n5566 19.3944
R15865 gnd.n5590 gnd.n5564 19.3944
R15866 gnd.n5594 gnd.n5564 19.3944
R15867 gnd.n5594 gnd.n5562 19.3944
R15868 gnd.n5600 gnd.n5562 19.3944
R15869 gnd.n5600 gnd.n5560 19.3944
R15870 gnd.n5604 gnd.n5560 19.3944
R15871 gnd.n5604 gnd.n5558 19.3944
R15872 gnd.n5610 gnd.n5558 19.3944
R15873 gnd.n5610 gnd.n5556 19.3944
R15874 gnd.n5617 gnd.n5556 19.3944
R15875 gnd.n5623 gnd.n5554 19.3944
R15876 gnd.n5623 gnd.n5552 19.3944
R15877 gnd.n5627 gnd.n5552 19.3944
R15878 gnd.n5627 gnd.n5550 19.3944
R15879 gnd.n5633 gnd.n5550 19.3944
R15880 gnd.n5633 gnd.n5548 19.3944
R15881 gnd.n5638 gnd.n5548 19.3944
R15882 gnd.n5646 gnd.n3298 19.3944
R15883 gnd.n5646 gnd.n3296 19.3944
R15884 gnd.n5650 gnd.n3296 19.3944
R15885 gnd.n5650 gnd.n3294 19.3944
R15886 gnd.n5656 gnd.n3294 19.3944
R15887 gnd.n5656 gnd.n3292 19.3944
R15888 gnd.n5660 gnd.n3292 19.3944
R15889 gnd.n5660 gnd.n3290 19.3944
R15890 gnd.n5672 gnd.n3288 19.3944
R15891 gnd.n5672 gnd.n3286 19.3944
R15892 gnd.n5678 gnd.n3286 19.3944
R15893 gnd.n5678 gnd.n3284 19.3944
R15894 gnd.n5682 gnd.n3284 19.3944
R15895 gnd.n5682 gnd.n3282 19.3944
R15896 gnd.n5688 gnd.n3282 19.3944
R15897 gnd.n5688 gnd.n3280 19.3944
R15898 gnd.n5692 gnd.n3280 19.3944
R15899 gnd.n5692 gnd.n3278 19.3944
R15900 gnd.n5698 gnd.n3278 19.3944
R15901 gnd.n5698 gnd.n3276 19.3944
R15902 gnd.n5702 gnd.n3276 19.3944
R15903 gnd.n5702 gnd.n3274 19.3944
R15904 gnd.n5708 gnd.n3274 19.3944
R15905 gnd.n5708 gnd.n3272 19.3944
R15906 gnd.n5713 gnd.n3272 19.3944
R15907 gnd.n5713 gnd.n3270 19.3944
R15908 gnd.n5726 gnd.n3263 19.3944
R15909 gnd.n5727 gnd.n5726 19.3944
R15910 gnd.n5728 gnd.n5727 19.3944
R15911 gnd.n5728 gnd.n3258 19.3944
R15912 gnd.n5740 gnd.n3258 19.3944
R15913 gnd.n5741 gnd.n5740 19.3944
R15914 gnd.n5742 gnd.n5741 19.3944
R15915 gnd.n5743 gnd.n5742 19.3944
R15916 gnd.n5745 gnd.n5743 19.3944
R15917 gnd.n5745 gnd.n3246 19.3944
R15918 gnd.n5805 gnd.n3246 19.3944
R15919 gnd.n5806 gnd.n5805 19.3944
R15920 gnd.n5808 gnd.n5806 19.3944
R15921 gnd.n5808 gnd.n3240 19.3944
R15922 gnd.n5830 gnd.n3240 19.3944
R15923 gnd.n5831 gnd.n5830 19.3944
R15924 gnd.n5832 gnd.n5831 19.3944
R15925 gnd.n5835 gnd.n5832 19.3944
R15926 gnd.n5835 gnd.n3238 19.3944
R15927 gnd.n5843 gnd.n3238 19.3944
R15928 gnd.n5844 gnd.n5843 19.3944
R15929 gnd.n5847 gnd.n5844 19.3944
R15930 gnd.n5848 gnd.n5847 19.3944
R15931 gnd.n5849 gnd.n5848 19.3944
R15932 gnd.n5857 gnd.n5849 19.3944
R15933 gnd.n5858 gnd.n5857 19.3944
R15934 gnd.n5859 gnd.n5858 19.3944
R15935 gnd.n5859 gnd.n3233 19.3944
R15936 gnd.n5872 gnd.n3233 19.3944
R15937 gnd.n5873 gnd.n5872 19.3944
R15938 gnd.n5874 gnd.n5873 19.3944
R15939 gnd.n5875 gnd.n5874 19.3944
R15940 gnd.n5905 gnd.n5875 19.3944
R15941 gnd.n5905 gnd.n5904 19.3944
R15942 gnd.n5904 gnd.n5903 19.3944
R15943 gnd.n5903 gnd.n5877 19.3944
R15944 gnd.n5893 gnd.n5877 19.3944
R15945 gnd.n5893 gnd.n5892 19.3944
R15946 gnd.n5892 gnd.n5891 19.3944
R15947 gnd.n5891 gnd.n175 19.3944
R15948 gnd.n7670 gnd.n175 19.3944
R15949 gnd.n7671 gnd.n7670 19.3944
R15950 gnd.n5723 gnd.n3074 19.3944
R15951 gnd.n5993 gnd.n3074 19.3944
R15952 gnd.n5993 gnd.n5992 19.3944
R15953 gnd.n5992 gnd.n5991 19.3944
R15954 gnd.n5991 gnd.n3078 19.3944
R15955 gnd.n5981 gnd.n3078 19.3944
R15956 gnd.n5981 gnd.n5980 19.3944
R15957 gnd.n5980 gnd.n5979 19.3944
R15958 gnd.n5979 gnd.n3098 19.3944
R15959 gnd.n5969 gnd.n3098 19.3944
R15960 gnd.n5969 gnd.n5968 19.3944
R15961 gnd.n5968 gnd.n5967 19.3944
R15962 gnd.n5967 gnd.n3119 19.3944
R15963 gnd.n5957 gnd.n3119 19.3944
R15964 gnd.n5957 gnd.n5956 19.3944
R15965 gnd.n5956 gnd.n5955 19.3944
R15966 gnd.n5955 gnd.n3138 19.3944
R15967 gnd.n5837 gnd.n3138 19.3944
R15968 gnd.n5840 gnd.n5837 19.3944
R15969 gnd.n5840 gnd.n3168 19.3944
R15970 gnd.n5933 gnd.n3168 19.3944
R15971 gnd.n5933 gnd.n5932 19.3944
R15972 gnd.n5932 gnd.n5931 19.3944
R15973 gnd.n5931 gnd.n5930 19.3944
R15974 gnd.n5930 gnd.n92 19.3944
R15975 gnd.n7721 gnd.n92 19.3944
R15976 gnd.n7721 gnd.n7720 19.3944
R15977 gnd.n7720 gnd.n7719 19.3944
R15978 gnd.n7719 gnd.n96 19.3944
R15979 gnd.n7709 gnd.n96 19.3944
R15980 gnd.n7709 gnd.n7708 19.3944
R15981 gnd.n7708 gnd.n7707 19.3944
R15982 gnd.n7707 gnd.n115 19.3944
R15983 gnd.n7697 gnd.n115 19.3944
R15984 gnd.n7697 gnd.n7696 19.3944
R15985 gnd.n7696 gnd.n7695 19.3944
R15986 gnd.n7695 gnd.n136 19.3944
R15987 gnd.n7685 gnd.n136 19.3944
R15988 gnd.n7685 gnd.n7684 19.3944
R15989 gnd.n7684 gnd.n7683 19.3944
R15990 gnd.n7683 gnd.n157 19.3944
R15991 gnd.n7673 gnd.n157 19.3944
R15992 gnd.n7580 gnd.n7516 19.3944
R15993 gnd.n7580 gnd.n7577 19.3944
R15994 gnd.n7577 gnd.n7574 19.3944
R15995 gnd.n7574 gnd.n7573 19.3944
R15996 gnd.n7573 gnd.n7570 19.3944
R15997 gnd.n7570 gnd.n7569 19.3944
R15998 gnd.n7569 gnd.n7566 19.3944
R15999 gnd.n7566 gnd.n7565 19.3944
R16000 gnd.n7565 gnd.n7562 19.3944
R16001 gnd.n7562 gnd.n7561 19.3944
R16002 gnd.n7561 gnd.n7558 19.3944
R16003 gnd.n7558 gnd.n7557 19.3944
R16004 gnd.n7557 gnd.n7554 19.3944
R16005 gnd.n7554 gnd.n7553 19.3944
R16006 gnd.n7553 gnd.n7550 19.3944
R16007 gnd.n7550 gnd.n7549 19.3944
R16008 gnd.n7549 gnd.n7546 19.3944
R16009 gnd.n7546 gnd.n7545 19.3944
R16010 gnd.n7623 gnd.n7620 19.3944
R16011 gnd.n7620 gnd.n7619 19.3944
R16012 gnd.n7619 gnd.n7616 19.3944
R16013 gnd.n7616 gnd.n7615 19.3944
R16014 gnd.n7615 gnd.n7612 19.3944
R16015 gnd.n7612 gnd.n7611 19.3944
R16016 gnd.n7611 gnd.n7608 19.3944
R16017 gnd.n7608 gnd.n7607 19.3944
R16018 gnd.n7607 gnd.n7604 19.3944
R16019 gnd.n7604 gnd.n7603 19.3944
R16020 gnd.n7603 gnd.n7600 19.3944
R16021 gnd.n7600 gnd.n7599 19.3944
R16022 gnd.n7599 gnd.n7596 19.3944
R16023 gnd.n7596 gnd.n7595 19.3944
R16024 gnd.n7595 gnd.n7592 19.3944
R16025 gnd.n7592 gnd.n7591 19.3944
R16026 gnd.n7591 gnd.n7588 19.3944
R16027 gnd.n7588 gnd.n7587 19.3944
R16028 gnd.n7478 gnd.n7477 19.3944
R16029 gnd.n7656 gnd.n7477 19.3944
R16030 gnd.n7656 gnd.n7655 19.3944
R16031 gnd.n7655 gnd.n7654 19.3944
R16032 gnd.n7654 gnd.n7651 19.3944
R16033 gnd.n7651 gnd.n7650 19.3944
R16034 gnd.n7650 gnd.n7647 19.3944
R16035 gnd.n7647 gnd.n7646 19.3944
R16036 gnd.n7646 gnd.n7643 19.3944
R16037 gnd.n7643 gnd.n7642 19.3944
R16038 gnd.n7642 gnd.n7639 19.3944
R16039 gnd.n7639 gnd.n7638 19.3944
R16040 gnd.n7638 gnd.n7635 19.3944
R16041 gnd.n7635 gnd.n7634 19.3944
R16042 gnd.n7634 gnd.n7631 19.3944
R16043 gnd.n7631 gnd.n7630 19.3944
R16044 gnd.n7630 gnd.n7627 19.3944
R16045 gnd.n204 gnd.n202 19.3944
R16046 gnd.n207 gnd.n204 19.3944
R16047 gnd.n207 gnd.n199 19.3944
R16048 gnd.n211 gnd.n199 19.3944
R16049 gnd.n214 gnd.n211 19.3944
R16050 gnd.n217 gnd.n214 19.3944
R16051 gnd.n217 gnd.n197 19.3944
R16052 gnd.n221 gnd.n197 19.3944
R16053 gnd.n224 gnd.n221 19.3944
R16054 gnd.n227 gnd.n224 19.3944
R16055 gnd.n227 gnd.n195 19.3944
R16056 gnd.n231 gnd.n195 19.3944
R16057 gnd.n234 gnd.n231 19.3944
R16058 gnd.n236 gnd.n234 19.3944
R16059 gnd.n236 gnd.n193 19.3944
R16060 gnd.n240 gnd.n193 19.3944
R16061 gnd.n5198 gnd.n5197 19.3944
R16062 gnd.n5197 gnd.n3262 19.3944
R16063 gnd.n5732 gnd.n3262 19.3944
R16064 gnd.n5732 gnd.n3260 19.3944
R16065 gnd.n5736 gnd.n3260 19.3944
R16066 gnd.n5736 gnd.n3254 19.3944
R16067 gnd.n5756 gnd.n3254 19.3944
R16068 gnd.n5756 gnd.n3255 19.3944
R16069 gnd.n5752 gnd.n3255 19.3944
R16070 gnd.n5752 gnd.n5751 19.3944
R16071 gnd.n5751 gnd.n5750 19.3944
R16072 gnd.n5750 gnd.n3245 19.3944
R16073 gnd.n5812 gnd.n3245 19.3944
R16074 gnd.n5812 gnd.n3242 19.3944
R16075 gnd.n5826 gnd.n3242 19.3944
R16076 gnd.n5826 gnd.n3243 19.3944
R16077 gnd.n5822 gnd.n3243 19.3944
R16078 gnd.n5822 gnd.n5821 19.3944
R16079 gnd.n5821 gnd.n5820 19.3944
R16080 gnd.n5820 gnd.n5818 19.3944
R16081 gnd.n5818 gnd.n64 19.3944
R16082 gnd.n7734 gnd.n64 19.3944
R16083 gnd.n7734 gnd.n7733 19.3944
R16084 gnd.n7733 gnd.n67 19.3944
R16085 gnd.n5853 gnd.n67 19.3944
R16086 gnd.n5853 gnd.n3237 19.3944
R16087 gnd.n5863 gnd.n3237 19.3944
R16088 gnd.n5863 gnd.n3235 19.3944
R16089 gnd.n5868 gnd.n3235 19.3944
R16090 gnd.n5868 gnd.n3228 19.3944
R16091 gnd.n5911 gnd.n3228 19.3944
R16092 gnd.n5911 gnd.n5910 19.3944
R16093 gnd.n5910 gnd.n5909 19.3944
R16094 gnd.n5909 gnd.n3232 19.3944
R16095 gnd.n5899 gnd.n3232 19.3944
R16096 gnd.n5899 gnd.n5898 19.3944
R16097 gnd.n5898 gnd.n5897 19.3944
R16098 gnd.n5897 gnd.n5882 19.3944
R16099 gnd.n5887 gnd.n5882 19.3944
R16100 gnd.n5887 gnd.n177 19.3944
R16101 gnd.n7666 gnd.n177 19.3944
R16102 gnd.n7666 gnd.n7665 19.3944
R16103 gnd.n5999 gnd.n5998 19.3944
R16104 gnd.n5998 gnd.n5997 19.3944
R16105 gnd.n5997 gnd.n3066 19.3944
R16106 gnd.n5987 gnd.n3066 19.3944
R16107 gnd.n5987 gnd.n5986 19.3944
R16108 gnd.n5986 gnd.n5985 19.3944
R16109 gnd.n5985 gnd.n3089 19.3944
R16110 gnd.n5975 gnd.n3089 19.3944
R16111 gnd.n5975 gnd.n5974 19.3944
R16112 gnd.n5974 gnd.n5973 19.3944
R16113 gnd.n5973 gnd.n3109 19.3944
R16114 gnd.n5963 gnd.n3109 19.3944
R16115 gnd.n5963 gnd.n5962 19.3944
R16116 gnd.n5962 gnd.n5961 19.3944
R16117 gnd.n5961 gnd.n3129 19.3944
R16118 gnd.n5951 gnd.n3129 19.3944
R16119 gnd.n3146 gnd.n3145 19.3944
R16120 gnd.n5938 gnd.n5937 19.3944
R16121 gnd.n3163 gnd.n3162 19.3944
R16122 gnd.n7729 gnd.n7728 19.3944
R16123 gnd.n7725 gnd.n76 19.3944
R16124 gnd.n7725 gnd.n83 19.3944
R16125 gnd.n7715 gnd.n83 19.3944
R16126 gnd.n7715 gnd.n7714 19.3944
R16127 gnd.n7714 gnd.n7713 19.3944
R16128 gnd.n7713 gnd.n106 19.3944
R16129 gnd.n7703 gnd.n106 19.3944
R16130 gnd.n7703 gnd.n7702 19.3944
R16131 gnd.n7702 gnd.n7701 19.3944
R16132 gnd.n7701 gnd.n126 19.3944
R16133 gnd.n7691 gnd.n126 19.3944
R16134 gnd.n7691 gnd.n7690 19.3944
R16135 gnd.n7690 gnd.n7689 19.3944
R16136 gnd.n7689 gnd.n147 19.3944
R16137 gnd.n7679 gnd.n147 19.3944
R16138 gnd.n7679 gnd.n7678 19.3944
R16139 gnd.n7678 gnd.n7677 19.3944
R16140 gnd.n6514 gnd.n875 19.3944
R16141 gnd.n6508 gnd.n875 19.3944
R16142 gnd.n6508 gnd.n6507 19.3944
R16143 gnd.n6507 gnd.n6506 19.3944
R16144 gnd.n6506 gnd.n2345 19.3944
R16145 gnd.n6500 gnd.n2345 19.3944
R16146 gnd.n6500 gnd.n6499 19.3944
R16147 gnd.n6499 gnd.n6498 19.3944
R16148 gnd.n6498 gnd.n2353 19.3944
R16149 gnd.n6492 gnd.n2353 19.3944
R16150 gnd.n6492 gnd.n6491 19.3944
R16151 gnd.n6491 gnd.n6490 19.3944
R16152 gnd.n6490 gnd.n2361 19.3944
R16153 gnd.n3922 gnd.n2361 19.3944
R16154 gnd.n4259 gnd.n3922 19.3944
R16155 gnd.n4259 gnd.n3919 19.3944
R16156 gnd.n4263 gnd.n3919 19.3944
R16157 gnd.n4263 gnd.n3917 19.3944
R16158 gnd.n4267 gnd.n3917 19.3944
R16159 gnd.n4267 gnd.n3915 19.3944
R16160 gnd.n4271 gnd.n3915 19.3944
R16161 gnd.n4271 gnd.n3913 19.3944
R16162 gnd.n4275 gnd.n3913 19.3944
R16163 gnd.n4275 gnd.n3911 19.3944
R16164 gnd.n4284 gnd.n3911 19.3944
R16165 gnd.n4284 gnd.n4283 19.3944
R16166 gnd.n4283 gnd.n4282 19.3944
R16167 gnd.n4282 gnd.n3884 19.3944
R16168 gnd.n4363 gnd.n3884 19.3944
R16169 gnd.n4363 gnd.n3885 19.3944
R16170 gnd.n4359 gnd.n4358 19.3944
R16171 gnd.n3889 gnd.n3888 19.3944
R16172 gnd.n4329 gnd.n4328 19.3944
R16173 gnd.n4326 gnd.n4325 19.3944
R16174 gnd.n4322 gnd.n3877 19.3944
R16175 gnd.n4387 gnd.n3877 19.3944
R16176 gnd.n4387 gnd.n4386 19.3944
R16177 gnd.n4386 gnd.n4385 19.3944
R16178 gnd.n4385 gnd.n4370 19.3944
R16179 gnd.n4381 gnd.n4370 19.3944
R16180 gnd.n4381 gnd.n4380 19.3944
R16181 gnd.n4380 gnd.n4379 19.3944
R16182 gnd.n4379 gnd.n4377 19.3944
R16183 gnd.n4377 gnd.n3855 19.3944
R16184 gnd.n4440 gnd.n3855 19.3944
R16185 gnd.n4440 gnd.n3853 19.3944
R16186 gnd.n4444 gnd.n3853 19.3944
R16187 gnd.n4444 gnd.n3851 19.3944
R16188 gnd.n4448 gnd.n3851 19.3944
R16189 gnd.n4448 gnd.n3849 19.3944
R16190 gnd.n4452 gnd.n3849 19.3944
R16191 gnd.n4452 gnd.n3847 19.3944
R16192 gnd.n4456 gnd.n3847 19.3944
R16193 gnd.n4456 gnd.n3845 19.3944
R16194 gnd.n4460 gnd.n3845 19.3944
R16195 gnd.n4460 gnd.n3842 19.3944
R16196 gnd.n4466 gnd.n3842 19.3944
R16197 gnd.n4466 gnd.n3840 19.3944
R16198 gnd.n4473 gnd.n3840 19.3944
R16199 gnd.n4473 gnd.n4472 19.3944
R16200 gnd.n4472 gnd.n2916 19.3944
R16201 gnd.n6147 gnd.n2916 19.3944
R16202 gnd.n6147 gnd.n6146 19.3944
R16203 gnd.n6146 gnd.n6145 19.3944
R16204 gnd.n6145 gnd.n2920 19.3944
R16205 gnd.n6133 gnd.n2920 19.3944
R16206 gnd.n6133 gnd.n6132 19.3944
R16207 gnd.n6132 gnd.n6131 19.3944
R16208 gnd.n6131 gnd.n2938 19.3944
R16209 gnd.n4558 gnd.n2938 19.3944
R16210 gnd.n4558 gnd.n3711 19.3944
R16211 gnd.n4590 gnd.n3711 19.3944
R16212 gnd.n4590 gnd.n3709 19.3944
R16213 gnd.n4594 gnd.n3709 19.3944
R16214 gnd.n4594 gnd.n3686 19.3944
R16215 gnd.n4633 gnd.n3686 19.3944
R16216 gnd.n4633 gnd.n3684 19.3944
R16217 gnd.n4637 gnd.n3684 19.3944
R16218 gnd.n4637 gnd.n3671 19.3944
R16219 gnd.n4678 gnd.n3671 19.3944
R16220 gnd.n4678 gnd.n3669 19.3944
R16221 gnd.n4684 gnd.n3669 19.3944
R16222 gnd.n4684 gnd.n4683 19.3944
R16223 gnd.n4683 gnd.n3643 19.3944
R16224 gnd.n4751 gnd.n3643 19.3944
R16225 gnd.n4751 gnd.n3641 19.3944
R16226 gnd.n4755 gnd.n3641 19.3944
R16227 gnd.n4755 gnd.n3623 19.3944
R16228 gnd.n4779 gnd.n3623 19.3944
R16229 gnd.n4779 gnd.n3621 19.3944
R16230 gnd.n4783 gnd.n3621 19.3944
R16231 gnd.n4783 gnd.n3602 19.3944
R16232 gnd.n4812 gnd.n3602 19.3944
R16233 gnd.n4812 gnd.n3600 19.3944
R16234 gnd.n4816 gnd.n3600 19.3944
R16235 gnd.n4816 gnd.n3585 19.3944
R16236 gnd.n4856 gnd.n3585 19.3944
R16237 gnd.n4856 gnd.n3583 19.3944
R16238 gnd.n4862 gnd.n3583 19.3944
R16239 gnd.n4862 gnd.n4861 19.3944
R16240 gnd.n4861 gnd.n3556 19.3944
R16241 gnd.n4906 gnd.n3556 19.3944
R16242 gnd.n4906 gnd.n3554 19.3944
R16243 gnd.n4910 gnd.n3554 19.3944
R16244 gnd.n4910 gnd.n3537 19.3944
R16245 gnd.n4934 gnd.n3537 19.3944
R16246 gnd.n4934 gnd.n3535 19.3944
R16247 gnd.n4947 gnd.n3535 19.3944
R16248 gnd.n4947 gnd.n4946 19.3944
R16249 gnd.n4946 gnd.n4945 19.3944
R16250 gnd.n4945 gnd.n3506 19.3944
R16251 gnd.n5009 gnd.n3506 19.3944
R16252 gnd.n5009 gnd.n3504 19.3944
R16253 gnd.n5015 gnd.n3504 19.3944
R16254 gnd.n5015 gnd.n5014 19.3944
R16255 gnd.n5014 gnd.n3478 19.3944
R16256 gnd.n5061 gnd.n3478 19.3944
R16257 gnd.n5061 gnd.n3476 19.3944
R16258 gnd.n5067 gnd.n3476 19.3944
R16259 gnd.n5067 gnd.n5066 19.3944
R16260 gnd.n5066 gnd.n3461 19.3944
R16261 gnd.n5089 gnd.n3461 19.3944
R16262 gnd.n5089 gnd.n3459 19.3944
R16263 gnd.n5093 gnd.n3459 19.3944
R16264 gnd.n5093 gnd.n3403 19.3944
R16265 gnd.n5132 gnd.n3403 19.3944
R16266 gnd.n5132 gnd.n3401 19.3944
R16267 gnd.n5136 gnd.n3401 19.3944
R16268 gnd.n5136 gnd.n3381 19.3944
R16269 gnd.n5160 gnd.n3381 19.3944
R16270 gnd.n5160 gnd.n3379 19.3944
R16271 gnd.n5167 gnd.n3379 19.3944
R16272 gnd.n5167 gnd.n5166 19.3944
R16273 gnd.n5166 gnd.n3350 19.3944
R16274 gnd.n5382 gnd.n3350 19.3944
R16275 gnd.n5382 gnd.n5381 19.3944
R16276 gnd.n5381 gnd.n5380 19.3944
R16277 gnd.n5380 gnd.n3356 19.3944
R16278 gnd.n3356 gnd.n3041 19.3944
R16279 gnd.n6014 gnd.n3041 19.3944
R16280 gnd.n6014 gnd.n6013 19.3944
R16281 gnd.n6013 gnd.n6012 19.3944
R16282 gnd.n6012 gnd.n3045 19.3944
R16283 gnd.n6006 gnd.n3045 19.3944
R16284 gnd.n6006 gnd.n6005 19.3944
R16285 gnd.n6005 gnd.n6004 19.3944
R16286 gnd.n6004 gnd.n3054 19.3944
R16287 gnd.n5768 gnd.n3054 19.3944
R16288 gnd.n5768 gnd.n5765 19.3944
R16289 gnd.n5772 gnd.n5765 19.3944
R16290 gnd.n5772 gnd.n5763 19.3944
R16291 gnd.n5776 gnd.n5763 19.3944
R16292 gnd.n5776 gnd.n5761 19.3944
R16293 gnd.n5780 gnd.n5761 19.3944
R16294 gnd.n5780 gnd.n3252 19.3944
R16295 gnd.n5784 gnd.n3252 19.3944
R16296 gnd.n5784 gnd.n3250 19.3944
R16297 gnd.n5800 gnd.n3250 19.3944
R16298 gnd.n5800 gnd.n5799 19.3944
R16299 gnd.n5799 gnd.n5798 19.3944
R16300 gnd.n5798 gnd.n5790 19.3944
R16301 gnd.n5794 gnd.n5790 19.3944
R16302 gnd.n5794 gnd.n5793 19.3944
R16303 gnd.n5946 gnd.n5945 19.3944
R16304 gnd.n5943 gnd.n3153 19.3944
R16305 gnd.n3180 gnd.n3177 19.3944
R16306 gnd.n5925 gnd.n3182 19.3944
R16307 gnd.n5923 gnd.n5922 19.3944
R16308 gnd.n5922 gnd.n3184 19.3944
R16309 gnd.n5918 gnd.n3184 19.3944
R16310 gnd.n5918 gnd.n5917 19.3944
R16311 gnd.n5917 gnd.n5916 19.3944
R16312 gnd.n5916 gnd.n3190 19.3944
R16313 gnd.n3224 gnd.n3190 19.3944
R16314 gnd.n3224 gnd.n3223 19.3944
R16315 gnd.n3223 gnd.n3222 19.3944
R16316 gnd.n3222 gnd.n3196 19.3944
R16317 gnd.n3218 gnd.n3196 19.3944
R16318 gnd.n3218 gnd.n3217 19.3944
R16319 gnd.n3217 gnd.n3216 19.3944
R16320 gnd.n3216 gnd.n3202 19.3944
R16321 gnd.n3212 gnd.n3202 19.3944
R16322 gnd.n3212 gnd.n3211 19.3944
R16323 gnd.n3211 gnd.n3210 19.3944
R16324 gnd.n3210 gnd.n246 19.3944
R16325 gnd.n7444 gnd.n246 19.3944
R16326 gnd.n7444 gnd.n7443 19.3944
R16327 gnd.n7443 gnd.n7442 19.3944
R16328 gnd.n7442 gnd.n250 19.3944
R16329 gnd.n7436 gnd.n250 19.3944
R16330 gnd.n7436 gnd.n7435 19.3944
R16331 gnd.n7435 gnd.n7434 19.3944
R16332 gnd.n7434 gnd.n258 19.3944
R16333 gnd.n7428 gnd.n258 19.3944
R16334 gnd.n7428 gnd.n7427 19.3944
R16335 gnd.n7427 gnd.n7426 19.3944
R16336 gnd.n7426 gnd.n266 19.3944
R16337 gnd.n4066 gnd.n4063 19.3944
R16338 gnd.n4066 gnd.n4061 19.3944
R16339 gnd.n4070 gnd.n4061 19.3944
R16340 gnd.n4070 gnd.n4059 19.3944
R16341 gnd.n4076 gnd.n4059 19.3944
R16342 gnd.n4076 gnd.n4057 19.3944
R16343 gnd.n4080 gnd.n4057 19.3944
R16344 gnd.n4080 gnd.n4055 19.3944
R16345 gnd.n4086 gnd.n4055 19.3944
R16346 gnd.n4086 gnd.n4053 19.3944
R16347 gnd.n4090 gnd.n4053 19.3944
R16348 gnd.n4090 gnd.n4051 19.3944
R16349 gnd.n4096 gnd.n4051 19.3944
R16350 gnd.n4096 gnd.n4049 19.3944
R16351 gnd.n4100 gnd.n4049 19.3944
R16352 gnd.n4100 gnd.n4044 19.3944
R16353 gnd.n4106 gnd.n4044 19.3944
R16354 gnd.n4110 gnd.n4042 19.3944
R16355 gnd.n4110 gnd.n4040 19.3944
R16356 gnd.n4116 gnd.n4040 19.3944
R16357 gnd.n4116 gnd.n4038 19.3944
R16358 gnd.n4120 gnd.n4038 19.3944
R16359 gnd.n4120 gnd.n4036 19.3944
R16360 gnd.n4126 gnd.n4036 19.3944
R16361 gnd.n4126 gnd.n4034 19.3944
R16362 gnd.n4130 gnd.n4034 19.3944
R16363 gnd.n4130 gnd.n4032 19.3944
R16364 gnd.n4136 gnd.n4032 19.3944
R16365 gnd.n4136 gnd.n4030 19.3944
R16366 gnd.n4140 gnd.n4030 19.3944
R16367 gnd.n4140 gnd.n4028 19.3944
R16368 gnd.n4146 gnd.n4028 19.3944
R16369 gnd.n4146 gnd.n4026 19.3944
R16370 gnd.n4150 gnd.n4026 19.3944
R16371 gnd.n4150 gnd.n4024 19.3944
R16372 gnd.n4162 gnd.n4022 19.3944
R16373 gnd.n4162 gnd.n4020 19.3944
R16374 gnd.n4168 gnd.n4020 19.3944
R16375 gnd.n4168 gnd.n4018 19.3944
R16376 gnd.n4172 gnd.n4018 19.3944
R16377 gnd.n4172 gnd.n4016 19.3944
R16378 gnd.n4178 gnd.n4016 19.3944
R16379 gnd.n4178 gnd.n4014 19.3944
R16380 gnd.n4182 gnd.n4014 19.3944
R16381 gnd.n4182 gnd.n4012 19.3944
R16382 gnd.n4188 gnd.n4012 19.3944
R16383 gnd.n4188 gnd.n4010 19.3944
R16384 gnd.n4192 gnd.n4010 19.3944
R16385 gnd.n4192 gnd.n4008 19.3944
R16386 gnd.n4198 gnd.n4008 19.3944
R16387 gnd.n4198 gnd.n4006 19.3944
R16388 gnd.n4203 gnd.n4006 19.3944
R16389 gnd.n4203 gnd.n4004 19.3944
R16390 gnd.n3998 gnd.n3932 19.3944
R16391 gnd.n3993 gnd.n3932 19.3944
R16392 gnd.n3993 gnd.n3992 19.3944
R16393 gnd.n3992 gnd.n3936 19.3944
R16394 gnd.n3987 gnd.n3936 19.3944
R16395 gnd.n3987 gnd.n3986 19.3944
R16396 gnd.n3986 gnd.n3985 19.3944
R16397 gnd.n3985 gnd.n3942 19.3944
R16398 gnd.n3979 gnd.n3942 19.3944
R16399 gnd.n3979 gnd.n3978 19.3944
R16400 gnd.n3978 gnd.n3977 19.3944
R16401 gnd.n3977 gnd.n3948 19.3944
R16402 gnd.n3971 gnd.n3948 19.3944
R16403 gnd.n3971 gnd.n3970 19.3944
R16404 gnd.n3970 gnd.n3969 19.3944
R16405 gnd.n3969 gnd.n3954 19.3944
R16406 gnd.n4254 gnd.n3925 19.3944
R16407 gnd.n4254 gnd.n4253 19.3944
R16408 gnd.n4253 gnd.n4252 19.3944
R16409 gnd.n4252 gnd.n3929 19.3944
R16410 gnd.n4242 gnd.n3929 19.3944
R16411 gnd.n4242 gnd.n4241 19.3944
R16412 gnd.n4241 gnd.n4240 19.3944
R16413 gnd.n4240 gnd.n4224 19.3944
R16414 gnd.n4230 gnd.n4224 19.3944
R16415 gnd.n4230 gnd.n3907 19.3944
R16416 gnd.n4289 gnd.n3907 19.3944
R16417 gnd.n4289 gnd.n3905 19.3944
R16418 gnd.n4293 gnd.n3905 19.3944
R16419 gnd.n4293 gnd.n3902 19.3944
R16420 gnd.n4303 gnd.n3902 19.3944
R16421 gnd.n4303 gnd.n3900 19.3944
R16422 gnd.n4308 gnd.n3900 19.3944
R16423 gnd.n4308 gnd.n3891 19.3944
R16424 gnd.n4352 gnd.n3891 19.3944
R16425 gnd.n4352 gnd.n4351 19.3944
R16426 gnd.n4351 gnd.n4350 19.3944
R16427 gnd.n4350 gnd.n3895 19.3944
R16428 gnd.n4346 gnd.n3895 19.3944
R16429 gnd.n4346 gnd.n4345 19.3944
R16430 gnd.n4345 gnd.n4344 19.3944
R16431 gnd.n4344 gnd.n3873 19.3944
R16432 gnd.n4392 gnd.n3873 19.3944
R16433 gnd.n4392 gnd.n3871 19.3944
R16434 gnd.n4396 gnd.n3871 19.3944
R16435 gnd.n4396 gnd.n3867 19.3944
R16436 gnd.n4406 gnd.n3867 19.3944
R16437 gnd.n4406 gnd.n3865 19.3944
R16438 gnd.n4410 gnd.n3865 19.3944
R16439 gnd.n4410 gnd.n3858 19.3944
R16440 gnd.n4434 gnd.n3858 19.3944
R16441 gnd.n4434 gnd.n3859 19.3944
R16442 gnd.n4430 gnd.n3859 19.3944
R16443 gnd.n4430 gnd.n4429 19.3944
R16444 gnd.n4429 gnd.n4428 19.3944
R16445 gnd.n4428 gnd.n2579 19.3944
R16446 gnd.n6348 gnd.n2579 19.3944
R16447 gnd.n6348 gnd.n2580 19.3944
R16448 gnd.n4216 gnd.n3930 19.3944
R16449 gnd.n4217 gnd.n4216 19.3944
R16450 gnd.n4248 gnd.n4217 19.3944
R16451 gnd.n4248 gnd.n4247 19.3944
R16452 gnd.n4247 gnd.n4246 19.3944
R16453 gnd.n4246 gnd.n4219 19.3944
R16454 gnd.n4236 gnd.n4219 19.3944
R16455 gnd.n4236 gnd.n4235 19.3944
R16456 gnd.n4235 gnd.n4234 19.3944
R16457 gnd.n4234 gnd.n4227 19.3944
R16458 gnd.n4227 gnd.n4226 19.3944
R16459 gnd.n4226 gnd.n3903 19.3944
R16460 gnd.n4297 gnd.n3903 19.3944
R16461 gnd.n4298 gnd.n4297 19.3944
R16462 gnd.n4299 gnd.n4298 19.3944
R16463 gnd.n4299 gnd.n3898 19.3944
R16464 gnd.n4312 gnd.n3898 19.3944
R16465 gnd.n4313 gnd.n4312 19.3944
R16466 gnd.n4314 gnd.n4313 19.3944
R16467 gnd.n4315 gnd.n4314 19.3944
R16468 gnd.n4319 gnd.n4315 19.3944
R16469 gnd.n4320 gnd.n4319 19.3944
R16470 gnd.n4334 gnd.n4320 19.3944
R16471 gnd.n4335 gnd.n4334 19.3944
R16472 gnd.n4339 gnd.n4335 19.3944
R16473 gnd.n4339 gnd.n4338 19.3944
R16474 gnd.n4338 gnd.n4337 19.3944
R16475 gnd.n4337 gnd.n3869 19.3944
R16476 gnd.n4400 gnd.n3869 19.3944
R16477 gnd.n4401 gnd.n4400 19.3944
R16478 gnd.n4402 gnd.n4401 19.3944
R16479 gnd.n4402 gnd.n3863 19.3944
R16480 gnd.n4414 gnd.n3863 19.3944
R16481 gnd.n4415 gnd.n4414 19.3944
R16482 gnd.n4416 gnd.n4415 19.3944
R16483 gnd.n4417 gnd.n4416 19.3944
R16484 gnd.n4421 gnd.n4417 19.3944
R16485 gnd.n4422 gnd.n4421 19.3944
R16486 gnd.n4423 gnd.n4422 19.3944
R16487 gnd.n4423 gnd.n2578 19.3944
R16488 gnd.n6352 gnd.n2578 19.3944
R16489 gnd.n6353 gnd.n6352 19.3944
R16490 gnd.n4213 gnd.n2380 19.3944
R16491 gnd.n6478 gnd.n2380 19.3944
R16492 gnd.n6478 gnd.n6477 19.3944
R16493 gnd.n6477 gnd.n6476 19.3944
R16494 gnd.n6476 gnd.n2384 19.3944
R16495 gnd.n6466 gnd.n2384 19.3944
R16496 gnd.n6466 gnd.n6465 19.3944
R16497 gnd.n6465 gnd.n6464 19.3944
R16498 gnd.n6464 gnd.n2405 19.3944
R16499 gnd.n6454 gnd.n2405 19.3944
R16500 gnd.n6454 gnd.n6453 19.3944
R16501 gnd.n6453 gnd.n6452 19.3944
R16502 gnd.n6452 gnd.n2426 19.3944
R16503 gnd.n6442 gnd.n2426 19.3944
R16504 gnd.n6442 gnd.n6441 19.3944
R16505 gnd.n6441 gnd.n6440 19.3944
R16506 gnd.n6440 gnd.n2446 19.3944
R16507 gnd.n6429 gnd.n2446 19.3944
R16508 gnd.n6429 gnd.n6428 19.3944
R16509 gnd.n6428 gnd.n6427 19.3944
R16510 gnd.n6427 gnd.n2465 19.3944
R16511 gnd.n6416 gnd.n2465 19.3944
R16512 gnd.n6416 gnd.n6415 19.3944
R16513 gnd.n6415 gnd.n6414 19.3944
R16514 gnd.n6414 gnd.n2481 19.3944
R16515 gnd.n6403 gnd.n2481 19.3944
R16516 gnd.n6403 gnd.n6402 19.3944
R16517 gnd.n6402 gnd.n6401 19.3944
R16518 gnd.n6401 gnd.n2499 19.3944
R16519 gnd.n6391 gnd.n2499 19.3944
R16520 gnd.n6391 gnd.n6390 19.3944
R16521 gnd.n6390 gnd.n6389 19.3944
R16522 gnd.n6389 gnd.n2518 19.3944
R16523 gnd.n6379 gnd.n2518 19.3944
R16524 gnd.n6379 gnd.n6378 19.3944
R16525 gnd.n6378 gnd.n6377 19.3944
R16526 gnd.n6377 gnd.n2539 19.3944
R16527 gnd.n6367 gnd.n2539 19.3944
R16528 gnd.n6367 gnd.n6366 19.3944
R16529 gnd.n6366 gnd.n6365 19.3944
R16530 gnd.n6365 gnd.n2559 19.3944
R16531 gnd.n6355 gnd.n2559 19.3944
R16532 gnd.n2722 gnd.n2721 19.3944
R16533 gnd.n6271 gnd.n2721 19.3944
R16534 gnd.n6271 gnd.n6270 19.3944
R16535 gnd.n6270 gnd.n6269 19.3944
R16536 gnd.n6269 gnd.n6266 19.3944
R16537 gnd.n6266 gnd.n6265 19.3944
R16538 gnd.n6265 gnd.n6262 19.3944
R16539 gnd.n6262 gnd.n6261 19.3944
R16540 gnd.n6261 gnd.n6258 19.3944
R16541 gnd.n6258 gnd.n6257 19.3944
R16542 gnd.n6257 gnd.n6254 19.3944
R16543 gnd.n6254 gnd.n6253 19.3944
R16544 gnd.n6253 gnd.n6250 19.3944
R16545 gnd.n6250 gnd.n6249 19.3944
R16546 gnd.n6249 gnd.n6246 19.3944
R16547 gnd.n6246 gnd.n6245 19.3944
R16548 gnd.n6245 gnd.n6242 19.3944
R16549 gnd.n2824 gnd.n2760 19.3944
R16550 gnd.n2824 gnd.n2821 19.3944
R16551 gnd.n2821 gnd.n2818 19.3944
R16552 gnd.n2818 gnd.n2817 19.3944
R16553 gnd.n2817 gnd.n2814 19.3944
R16554 gnd.n2814 gnd.n2813 19.3944
R16555 gnd.n2813 gnd.n2810 19.3944
R16556 gnd.n2810 gnd.n2809 19.3944
R16557 gnd.n2809 gnd.n2806 19.3944
R16558 gnd.n2806 gnd.n2805 19.3944
R16559 gnd.n2805 gnd.n2802 19.3944
R16560 gnd.n2802 gnd.n2801 19.3944
R16561 gnd.n2801 gnd.n2798 19.3944
R16562 gnd.n2798 gnd.n2797 19.3944
R16563 gnd.n2797 gnd.n2794 19.3944
R16564 gnd.n2794 gnd.n2793 19.3944
R16565 gnd.n2793 gnd.n2790 19.3944
R16566 gnd.n2790 gnd.n2789 19.3944
R16567 gnd.n2846 gnd.n2751 19.3944
R16568 gnd.n2846 gnd.n2843 19.3944
R16569 gnd.n2843 gnd.n2840 19.3944
R16570 gnd.n2840 gnd.n2839 19.3944
R16571 gnd.n2839 gnd.n2836 19.3944
R16572 gnd.n2836 gnd.n2835 19.3944
R16573 gnd.n2835 gnd.n2832 19.3944
R16574 gnd.n2832 gnd.n2831 19.3944
R16575 gnd.n6240 gnd.n6237 19.3944
R16576 gnd.n6237 gnd.n6236 19.3944
R16577 gnd.n6236 gnd.n6233 19.3944
R16578 gnd.n6233 gnd.n6232 19.3944
R16579 gnd.n6232 gnd.n6229 19.3944
R16580 gnd.n6229 gnd.n6228 19.3944
R16581 gnd.n6228 gnd.n6225 19.3944
R16582 gnd.n6484 gnd.n6483 19.3944
R16583 gnd.n6483 gnd.n6482 19.3944
R16584 gnd.n6482 gnd.n2373 19.3944
R16585 gnd.n6472 gnd.n2373 19.3944
R16586 gnd.n6472 gnd.n6471 19.3944
R16587 gnd.n6471 gnd.n6470 19.3944
R16588 gnd.n6470 gnd.n2395 19.3944
R16589 gnd.n6460 gnd.n2395 19.3944
R16590 gnd.n6460 gnd.n6459 19.3944
R16591 gnd.n6459 gnd.n6458 19.3944
R16592 gnd.n6458 gnd.n2416 19.3944
R16593 gnd.n6448 gnd.n2416 19.3944
R16594 gnd.n6448 gnd.n6447 19.3944
R16595 gnd.n6447 gnd.n6446 19.3944
R16596 gnd.n6446 gnd.n2436 19.3944
R16597 gnd.n6436 gnd.n2436 19.3944
R16598 gnd.n6434 gnd.n6433 19.3944
R16599 gnd.n6423 gnd.n2471 19.3944
R16600 gnd.n6421 gnd.n6420 19.3944
R16601 gnd.n6410 gnd.n2488 19.3944
R16602 gnd.n6408 gnd.n6407 19.3944
R16603 gnd.n6407 gnd.n2489 19.3944
R16604 gnd.n6397 gnd.n2489 19.3944
R16605 gnd.n6397 gnd.n6396 19.3944
R16606 gnd.n6396 gnd.n6395 19.3944
R16607 gnd.n6395 gnd.n2509 19.3944
R16608 gnd.n6385 gnd.n2509 19.3944
R16609 gnd.n6385 gnd.n6384 19.3944
R16610 gnd.n6384 gnd.n6383 19.3944
R16611 gnd.n6383 gnd.n2529 19.3944
R16612 gnd.n6373 gnd.n2529 19.3944
R16613 gnd.n6373 gnd.n6372 19.3944
R16614 gnd.n6372 gnd.n6371 19.3944
R16615 gnd.n6371 gnd.n2549 19.3944
R16616 gnd.n6361 gnd.n2549 19.3944
R16617 gnd.n6361 gnd.n6360 19.3944
R16618 gnd.n6360 gnd.n6359 19.3944
R16619 gnd.n6685 gnd.n6684 19.3944
R16620 gnd.n6684 gnd.n708 19.3944
R16621 gnd.n6678 gnd.n708 19.3944
R16622 gnd.n6678 gnd.n6677 19.3944
R16623 gnd.n6677 gnd.n6676 19.3944
R16624 gnd.n6676 gnd.n716 19.3944
R16625 gnd.n6670 gnd.n716 19.3944
R16626 gnd.n6670 gnd.n6669 19.3944
R16627 gnd.n6669 gnd.n6668 19.3944
R16628 gnd.n6668 gnd.n724 19.3944
R16629 gnd.n6662 gnd.n724 19.3944
R16630 gnd.n6662 gnd.n6661 19.3944
R16631 gnd.n6661 gnd.n6660 19.3944
R16632 gnd.n6660 gnd.n732 19.3944
R16633 gnd.n6654 gnd.n732 19.3944
R16634 gnd.n6654 gnd.n6653 19.3944
R16635 gnd.n6653 gnd.n6652 19.3944
R16636 gnd.n6652 gnd.n740 19.3944
R16637 gnd.n6646 gnd.n740 19.3944
R16638 gnd.n6646 gnd.n6645 19.3944
R16639 gnd.n6645 gnd.n6644 19.3944
R16640 gnd.n6644 gnd.n748 19.3944
R16641 gnd.n6638 gnd.n748 19.3944
R16642 gnd.n6638 gnd.n6637 19.3944
R16643 gnd.n6637 gnd.n6636 19.3944
R16644 gnd.n6636 gnd.n756 19.3944
R16645 gnd.n6630 gnd.n756 19.3944
R16646 gnd.n6630 gnd.n6629 19.3944
R16647 gnd.n6629 gnd.n6628 19.3944
R16648 gnd.n6628 gnd.n764 19.3944
R16649 gnd.n6622 gnd.n764 19.3944
R16650 gnd.n6622 gnd.n6621 19.3944
R16651 gnd.n6621 gnd.n6620 19.3944
R16652 gnd.n6620 gnd.n772 19.3944
R16653 gnd.n6614 gnd.n772 19.3944
R16654 gnd.n6614 gnd.n6613 19.3944
R16655 gnd.n6613 gnd.n6612 19.3944
R16656 gnd.n6612 gnd.n780 19.3944
R16657 gnd.n6606 gnd.n780 19.3944
R16658 gnd.n6606 gnd.n6605 19.3944
R16659 gnd.n6605 gnd.n6604 19.3944
R16660 gnd.n6604 gnd.n788 19.3944
R16661 gnd.n6598 gnd.n788 19.3944
R16662 gnd.n6598 gnd.n6597 19.3944
R16663 gnd.n6597 gnd.n6596 19.3944
R16664 gnd.n6596 gnd.n796 19.3944
R16665 gnd.n6590 gnd.n796 19.3944
R16666 gnd.n6590 gnd.n6589 19.3944
R16667 gnd.n6589 gnd.n6588 19.3944
R16668 gnd.n6588 gnd.n804 19.3944
R16669 gnd.n6582 gnd.n804 19.3944
R16670 gnd.n6582 gnd.n6581 19.3944
R16671 gnd.n6581 gnd.n6580 19.3944
R16672 gnd.n6580 gnd.n812 19.3944
R16673 gnd.n6574 gnd.n812 19.3944
R16674 gnd.n6574 gnd.n6573 19.3944
R16675 gnd.n6573 gnd.n6572 19.3944
R16676 gnd.n6572 gnd.n820 19.3944
R16677 gnd.n6566 gnd.n820 19.3944
R16678 gnd.n6566 gnd.n6565 19.3944
R16679 gnd.n6565 gnd.n6564 19.3944
R16680 gnd.n6564 gnd.n828 19.3944
R16681 gnd.n6558 gnd.n828 19.3944
R16682 gnd.n6558 gnd.n6557 19.3944
R16683 gnd.n6557 gnd.n6556 19.3944
R16684 gnd.n6556 gnd.n836 19.3944
R16685 gnd.n6550 gnd.n836 19.3944
R16686 gnd.n6550 gnd.n6549 19.3944
R16687 gnd.n6549 gnd.n6548 19.3944
R16688 gnd.n6548 gnd.n844 19.3944
R16689 gnd.n6542 gnd.n844 19.3944
R16690 gnd.n6542 gnd.n6541 19.3944
R16691 gnd.n6541 gnd.n6540 19.3944
R16692 gnd.n6540 gnd.n852 19.3944
R16693 gnd.n6534 gnd.n852 19.3944
R16694 gnd.n6534 gnd.n6533 19.3944
R16695 gnd.n6533 gnd.n6532 19.3944
R16696 gnd.n6532 gnd.n860 19.3944
R16697 gnd.n6526 gnd.n860 19.3944
R16698 gnd.n6526 gnd.n6525 19.3944
R16699 gnd.n6525 gnd.n6524 19.3944
R16700 gnd.n6524 gnd.n868 19.3944
R16701 gnd.n6518 gnd.n868 19.3944
R16702 gnd.n6518 gnd.n6517 19.3944
R16703 gnd.n4478 gnd.n3831 19.3944
R16704 gnd.n4478 gnd.n3828 19.3944
R16705 gnd.n4483 gnd.n3828 19.3944
R16706 gnd.n4483 gnd.n3829 19.3944
R16707 gnd.n3829 gnd.n3743 19.3944
R16708 gnd.n4510 gnd.n3743 19.3944
R16709 gnd.n4510 gnd.n3740 19.3944
R16710 gnd.n4515 gnd.n3740 19.3944
R16711 gnd.n4515 gnd.n3741 19.3944
R16712 gnd.n3741 gnd.n2945 19.3944
R16713 gnd.n6126 gnd.n2945 19.3944
R16714 gnd.n6126 gnd.n2946 19.3944
R16715 gnd.n6122 gnd.n2946 19.3944
R16716 gnd.n6122 gnd.n6121 19.3944
R16717 gnd.n6121 gnd.n6120 19.3944
R16718 gnd.n6120 gnd.n2952 19.3944
R16719 gnd.n6116 gnd.n2952 19.3944
R16720 gnd.n6116 gnd.n6115 19.3944
R16721 gnd.n6115 gnd.n6114 19.3944
R16722 gnd.n6114 gnd.n2957 19.3944
R16723 gnd.n6110 gnd.n2957 19.3944
R16724 gnd.n6110 gnd.n6109 19.3944
R16725 gnd.n6109 gnd.n6108 19.3944
R16726 gnd.n6108 gnd.n2962 19.3944
R16727 gnd.n6104 gnd.n2962 19.3944
R16728 gnd.n6104 gnd.n6103 19.3944
R16729 gnd.n6103 gnd.n6102 19.3944
R16730 gnd.n6102 gnd.n2967 19.3944
R16731 gnd.n6098 gnd.n2967 19.3944
R16732 gnd.n6098 gnd.n6097 19.3944
R16733 gnd.n6097 gnd.n6096 19.3944
R16734 gnd.n6096 gnd.n2972 19.3944
R16735 gnd.n6092 gnd.n2972 19.3944
R16736 gnd.n6092 gnd.n6091 19.3944
R16737 gnd.n6091 gnd.n6090 19.3944
R16738 gnd.n6090 gnd.n2977 19.3944
R16739 gnd.n6086 gnd.n2977 19.3944
R16740 gnd.n6086 gnd.n6085 19.3944
R16741 gnd.n6085 gnd.n6084 19.3944
R16742 gnd.n6084 gnd.n2982 19.3944
R16743 gnd.n6080 gnd.n2982 19.3944
R16744 gnd.n6080 gnd.n6079 19.3944
R16745 gnd.n6079 gnd.n6078 19.3944
R16746 gnd.n6078 gnd.n2987 19.3944
R16747 gnd.n6074 gnd.n2987 19.3944
R16748 gnd.n6074 gnd.n6073 19.3944
R16749 gnd.n6073 gnd.n6072 19.3944
R16750 gnd.n6072 gnd.n2992 19.3944
R16751 gnd.n6068 gnd.n2992 19.3944
R16752 gnd.n6068 gnd.n6067 19.3944
R16753 gnd.n6067 gnd.n6066 19.3944
R16754 gnd.n6066 gnd.n2997 19.3944
R16755 gnd.n6062 gnd.n2997 19.3944
R16756 gnd.n6062 gnd.n6061 19.3944
R16757 gnd.n6061 gnd.n6060 19.3944
R16758 gnd.n6060 gnd.n3002 19.3944
R16759 gnd.n6056 gnd.n3002 19.3944
R16760 gnd.n6056 gnd.n6055 19.3944
R16761 gnd.n6055 gnd.n6054 19.3944
R16762 gnd.n6054 gnd.n3007 19.3944
R16763 gnd.n6050 gnd.n3007 19.3944
R16764 gnd.n6050 gnd.n6049 19.3944
R16765 gnd.n6049 gnd.n6048 19.3944
R16766 gnd.n6048 gnd.n3012 19.3944
R16767 gnd.n6044 gnd.n3012 19.3944
R16768 gnd.n6044 gnd.n6043 19.3944
R16769 gnd.n6043 gnd.n6042 19.3944
R16770 gnd.n6042 gnd.n3017 19.3944
R16771 gnd.n6038 gnd.n3017 19.3944
R16772 gnd.n6038 gnd.n6037 19.3944
R16773 gnd.n6037 gnd.n6036 19.3944
R16774 gnd.n6036 gnd.n3022 19.3944
R16775 gnd.n6032 gnd.n3022 19.3944
R16776 gnd.n6032 gnd.n6031 19.3944
R16777 gnd.n6031 gnd.n6030 19.3944
R16778 gnd.n6030 gnd.n3027 19.3944
R16779 gnd.n6026 gnd.n3027 19.3944
R16780 gnd.n6026 gnd.n6025 19.3944
R16781 gnd.n6025 gnd.n6024 19.3944
R16782 gnd.n6024 gnd.n3032 19.3944
R16783 gnd.n6020 gnd.n3032 19.3944
R16784 gnd.n6020 gnd.n6019 19.3944
R16785 gnd.n5260 gnd.n5257 19.3944
R16786 gnd.n5260 gnd.n5255 19.3944
R16787 gnd.n5266 gnd.n5255 19.3944
R16788 gnd.n5266 gnd.n5253 19.3944
R16789 gnd.n5271 gnd.n5253 19.3944
R16790 gnd.n5271 gnd.n5251 19.3944
R16791 gnd.n5277 gnd.n5251 19.3944
R16792 gnd.n5277 gnd.n5250 19.3944
R16793 gnd.n5286 gnd.n5250 19.3944
R16794 gnd.n5286 gnd.n5248 19.3944
R16795 gnd.n5292 gnd.n5248 19.3944
R16796 gnd.n5292 gnd.n5241 19.3944
R16797 gnd.n5305 gnd.n5241 19.3944
R16798 gnd.n5305 gnd.n5239 19.3944
R16799 gnd.n5311 gnd.n5239 19.3944
R16800 gnd.n5311 gnd.n5232 19.3944
R16801 gnd.n5324 gnd.n5232 19.3944
R16802 gnd.n5324 gnd.n5230 19.3944
R16803 gnd.n5330 gnd.n5230 19.3944
R16804 gnd.n5330 gnd.n5223 19.3944
R16805 gnd.n5343 gnd.n5223 19.3944
R16806 gnd.n5343 gnd.n5221 19.3944
R16807 gnd.n5350 gnd.n5221 19.3944
R16808 gnd.n5350 gnd.n5349 19.3944
R16809 gnd.n5363 gnd.n5202 19.3944
R16810 gnd.n5202 gnd.n5201 19.3944
R16811 gnd.n5370 gnd.n5201 19.3944
R16812 gnd.n1723 gnd.t159 18.8012
R16813 gnd.n1708 gnd.t316 18.8012
R16814 gnd.n1567 gnd.n1566 18.4825
R16815 gnd.n5638 gnd.n5546 18.4247
R16816 gnd.n6225 gnd.n6224 18.4247
R16817 gnd.n5360 gnd.n5359 18.2308
R16818 gnd.n6279 gnd.n6278 18.2308
R16819 gnd.n240 gnd.n182 18.2308
R16820 gnd.n3963 gnd.n3954 18.2308
R16821 gnd.t167 gnd.n1247 18.1639
R16822 gnd.n1853 gnd.n870 18.1639
R16823 gnd.n1275 gnd.t3 17.5266
R16824 gnd.n1674 gnd.t173 16.8893
R16825 gnd.n6350 gnd.t87 16.8893
R16826 gnd.n5195 gnd.t63 16.8893
R16827 gnd.n5668 gnd.n3290 16.6793
R16828 gnd.n7587 gnd.n7584 16.6793
R16829 gnd.n4158 gnd.n4024 16.6793
R16830 gnd.n2831 gnd.n2828 16.6793
R16831 gnd.n1502 gnd.t48 16.2519
R16832 gnd.n1202 gnd.t165 16.2519
R16833 gnd.n6339 gnd.n2587 15.9333
R16834 gnd.n6339 gnd.n2601 15.9333
R16835 gnd.n4464 gnd.n4463 15.9333
R16836 gnd.n4463 gnd.n3832 15.9333
R16837 gnd.n4476 gnd.n3832 15.9333
R16838 gnd.n4476 gnd.n4475 15.9333
R16839 gnd.n4485 gnd.n2886 15.9333
R16840 gnd.n4500 gnd.n4499 15.9333
R16841 gnd.n6142 gnd.n2924 15.9333
R16842 gnd.n6135 gnd.n2932 15.9333
R16843 gnd.n4560 gnd.n4555 15.9333
R16844 gnd.n4588 gnd.n4587 15.9333
R16845 gnd.n4598 gnd.n4596 15.9333
R16846 gnd.n4631 gnd.n3688 15.9333
R16847 gnd.n4676 gnd.n3673 15.9333
R16848 gnd.n4688 gnd.n4686 15.9333
R16849 gnd.n4652 gnd.n3661 15.9333
R16850 gnd.n4749 gnd.n4748 15.9333
R16851 gnd.n4757 gnd.n3639 15.9333
R16852 gnd.n4777 gnd.n4776 15.9333
R16853 gnd.n4786 gnd.n4785 15.9333
R16854 gnd.n4810 gnd.n3604 15.9333
R16855 gnd.n4818 gnd.n3598 15.9333
R16856 gnd.n4854 gnd.n3587 15.9333
R16857 gnd.n4865 gnd.n3579 15.9333
R16858 gnd.n4865 gnd.n4864 15.9333
R16859 gnd.n4831 gnd.n3575 15.9333
R16860 gnd.n4904 gnd.n4903 15.9333
R16861 gnd.n4912 gnd.n3552 15.9333
R16862 gnd.n4932 gnd.n4931 15.9333
R16863 gnd.n4950 gnd.n4949 15.9333
R16864 gnd.n4943 gnd.n4942 15.9333
R16865 gnd.n5007 gnd.n3508 15.9333
R16866 gnd.n5019 gnd.n5017 15.9333
R16867 gnd.n4984 gnd.n3497 15.9333
R16868 gnd.n5059 gnd.n5058 15.9333
R16869 gnd.n5086 gnd.n5085 15.9333
R16870 gnd.n5112 gnd.n3420 15.9333
R16871 gnd.n5096 gnd.n3411 15.9333
R16872 gnd.n3450 gnd.n3407 15.9333
R16873 gnd.n5189 gnd.n3340 15.9333
R16874 gnd.n5189 gnd.n3303 15.9333
R16875 gnd.n5377 gnd.n5376 15.9333
R16876 gnd.n5376 gnd.n3036 15.9333
R16877 gnd.n6017 gnd.n3036 15.9333
R16878 gnd.n6017 gnd.n6016 15.9333
R16879 gnd.n3047 gnd.n3038 15.9333
R16880 gnd.n6010 gnd.n3047 15.9333
R16881 gnd.n2191 gnd.n2189 15.6674
R16882 gnd.n2159 gnd.n2157 15.6674
R16883 gnd.n2127 gnd.n2125 15.6674
R16884 gnd.n2096 gnd.n2094 15.6674
R16885 gnd.n2064 gnd.n2062 15.6674
R16886 gnd.n2032 gnd.n2030 15.6674
R16887 gnd.n2000 gnd.n1998 15.6674
R16888 gnd.n1969 gnd.n1967 15.6674
R16889 gnd.n1493 gnd.t48 15.6146
R16890 gnd.t38 gnd.n958 15.6146
R16891 gnd.t142 gnd.n959 15.6146
R16892 gnd.t113 gnd.n2854 15.6146
R16893 gnd.n3358 gnd.t94 15.6146
R16894 gnd.n5720 gnd.n3269 15.3217
R16895 gnd.n7542 gnd.n7537 15.3217
R16896 gnd.n4210 gnd.n4003 15.3217
R16897 gnd.n2786 gnd.n2781 15.3217
R16898 gnd.n3432 gnd.t76 15.296
R16899 gnd.n5393 gnd.n5392 15.0827
R16900 gnd.n2898 gnd.n2893 15.0481
R16901 gnd.n5403 gnd.n5402 15.0481
R16902 gnd.n1863 gnd.t171 14.9773
R16903 gnd.n6480 gnd.t55 14.9773
R16904 gnd.n6129 gnd.t1 14.9773
R16905 gnd.t185 gnd.n5147 14.9773
R16906 gnd.n7681 gnd.t59 14.9773
R16907 gnd.n3734 gnd.n3733 14.6587
R16908 gnd.n4606 gnd.t0 14.6587
R16909 gnd.n4668 gnd.n4667 14.6587
R16910 gnd.n5056 gnd.n3483 14.6587
R16911 gnd.n5104 gnd.t191 14.6587
R16912 gnd.n5158 gnd.n5157 14.6587
R16913 gnd.n5385 gnd.n5384 14.6587
R16914 gnd.t168 gnd.n1001 14.34
R16915 gnd.n1941 gnd.t172 14.34
R16916 gnd.n4561 gnd.n3724 14.0214
R16917 gnd.n4630 gnd.t189 14.0214
R16918 gnd.n4758 gnd.n3636 14.0214
R16919 gnd.n4809 gnd.n3607 14.0214
R16920 gnd.n4913 gnd.n3549 14.0214
R16921 gnd.n4972 gnd.n4971 14.0214
R16922 gnd.t9 gnd.n3463 14.0214
R16923 gnd.n3451 gnd.n3398 14.0214
R16924 gnd.t42 gnd.n3345 14.0214
R16925 gnd.n1649 gnd.t161 13.7027
R16926 gnd.n1359 gnd.n1358 13.5763
R16927 gnd.n2305 gnd.n915 13.5763
R16928 gnd.n1567 gnd.n1305 13.384
R16929 gnd.n6149 gnd.t45 13.384
R16930 gnd.n4525 gnd.n2942 13.384
R16931 gnd.n4624 gnd.n3693 13.384
R16932 gnd.n4660 gnd.t27 13.384
R16933 gnd.n4746 gnd.n3648 13.384
R16934 gnd.n4803 gnd.n4802 13.384
R16935 gnd.n4902 gnd.n3561 13.384
R16936 gnd.n4999 gnd.n4998 13.384
R16937 gnd.t164 gnd.n3487 13.384
R16938 gnd.n5034 gnd.n3468 13.384
R16939 gnd.n5138 gnd.n3390 13.384
R16940 gnd.n2909 gnd.n2890 13.1884
R16941 gnd.n2904 gnd.n2903 13.1884
R16942 gnd.n2903 gnd.n2902 13.1884
R16943 gnd.n5396 gnd.n5391 13.1884
R16944 gnd.n5397 gnd.n5396 13.1884
R16945 gnd.n2905 gnd.n2892 13.146
R16946 gnd.n2901 gnd.n2892 13.146
R16947 gnd.n5395 gnd.n5394 13.146
R16948 gnd.n5395 gnd.n5390 13.146
R16949 gnd.n2192 gnd.n2188 12.8005
R16950 gnd.n2160 gnd.n2156 12.8005
R16951 gnd.n2128 gnd.n2124 12.8005
R16952 gnd.n2097 gnd.n2093 12.8005
R16953 gnd.n2065 gnd.n2061 12.8005
R16954 gnd.n2033 gnd.n2029 12.8005
R16955 gnd.n2001 gnd.n1997 12.8005
R16956 gnd.n1970 gnd.n1966 12.8005
R16957 gnd.n3824 gnd.n2912 12.7467
R16958 gnd.t73 gnd.t83 12.7467
R16959 gnd.n4540 gnd.n2940 12.7467
R16960 gnd.t6 gnd.n3713 12.7467
R16961 gnd.n4640 gnd.n3679 12.7467
R16962 gnd.n4739 gnd.n3645 12.7467
R16963 gnd.n4819 gnd.n3594 12.7467
R16964 gnd.n4895 gnd.n3558 12.7467
R16965 gnd.n5006 gnd.n3510 12.7467
R16966 gnd.n5070 gnd.n3473 12.7467
R16967 gnd.n5123 gnd.t160 12.7467
R16968 gnd.n5146 gnd.n3393 12.7467
R16969 gnd.n5169 gnd.t101 12.7467
R16970 gnd.n1358 gnd.n1353 12.4126
R16971 gnd.n2308 gnd.n2305 12.4126
R16972 gnd.n6217 gnd.n6154 12.1761
R16973 gnd.n5472 gnd.n5471 12.1761
R16974 gnd.n4554 gnd.n3718 12.1094
R16975 gnd.n4576 gnd.n3702 12.1094
R16976 gnd.n3638 gnd.n3630 12.1094
R16977 gnd.n4795 gnd.n4794 12.1094
R16978 gnd.n3551 gnd.n3544 12.1094
R16979 gnd.n4940 gnd.n3525 12.1094
R16980 gnd.n5083 gnd.n3425 12.1094
R16981 gnd.n5130 gnd.n5129 12.1094
R16982 gnd.n2196 gnd.n2195 12.0247
R16983 gnd.n2164 gnd.n2163 12.0247
R16984 gnd.n2132 gnd.n2131 12.0247
R16985 gnd.n2101 gnd.n2100 12.0247
R16986 gnd.n2069 gnd.n2068 12.0247
R16987 gnd.n2037 gnd.n2036 12.0247
R16988 gnd.n2005 gnd.n2004 12.0247
R16989 gnd.n1974 gnd.n1973 12.0247
R16990 gnd.n6375 gnd.t207 11.7908
R16991 gnd.n5983 gnd.t214 11.7908
R16992 gnd.n6274 gnd.n2690 11.4721
R16993 gnd.n4508 gnd.n3747 11.4721
R16994 gnd.n4675 gnd.n3675 11.4721
R16995 gnd.n4695 gnd.n4694 11.4721
R16996 gnd.n4853 gnd.n3590 11.4721
R16997 gnd.n4872 gnd.n4871 11.4721
R16998 gnd.n5027 gnd.n3495 11.4721
R16999 gnd.n5049 gnd.n3480 11.4721
R17000 gnd.n5172 gnd.n5171 11.4721
R17001 gnd.n3436 gnd.n3434 11.4721
R17002 gnd.n6008 gnd.n3048 11.4721
R17003 gnd.n2199 gnd.n2186 11.249
R17004 gnd.n2167 gnd.n2154 11.249
R17005 gnd.n2135 gnd.n2122 11.249
R17006 gnd.n2104 gnd.n2091 11.249
R17007 gnd.n2072 gnd.n2059 11.249
R17008 gnd.n2040 gnd.n2027 11.249
R17009 gnd.n2008 gnd.n1995 11.249
R17010 gnd.n1977 gnd.n1964 11.249
R17011 gnd.n1637 gnd.t161 11.1535
R17012 gnd.n4286 gnd.t227 11.1535
R17013 gnd.n6399 gnd.t201 11.1535
R17014 gnd.n5959 gnd.t222 11.1535
R17015 gnd.n5914 gnd.t260 11.1535
R17016 gnd.n6486 gnd.n2366 10.8348
R17017 gnd.n4257 gnd.n4256 10.8348
R17018 gnd.n6480 gnd.n2377 10.8348
R17019 gnd.n4250 gnd.n2386 10.8348
R17020 gnd.n6474 gnd.n2389 10.8348
R17021 gnd.n4244 gnd.n2397 10.8348
R17022 gnd.n6468 gnd.n2400 10.8348
R17023 gnd.n4238 gnd.n2407 10.8348
R17024 gnd.n6462 gnd.n2410 10.8348
R17025 gnd.n6456 gnd.n2421 10.8348
R17026 gnd.n4287 gnd.n4286 10.8348
R17027 gnd.n6450 gnd.n2430 10.8348
R17028 gnd.n4295 gnd.n2438 10.8348
R17029 gnd.n6444 gnd.n2441 10.8348
R17030 gnd.n4301 gnd.n2448 10.8348
R17031 gnd.n6438 gnd.n2451 10.8348
R17032 gnd.n6431 gnd.n2460 10.8348
R17033 gnd.n4355 gnd.n4354 10.8348
R17034 gnd.n6425 gnd.n2469 10.8348
R17035 gnd.n4317 gnd.n2474 10.8348
R17036 gnd.n4332 gnd.n2483 10.8348
R17037 gnd.n6412 gnd.n2486 10.8348
R17038 gnd.n4341 gnd.n2491 10.8348
R17039 gnd.n6405 gnd.n2494 10.8348
R17040 gnd.n4390 gnd.n4389 10.8348
R17041 gnd.n6399 gnd.n2503 10.8348
R17042 gnd.n4398 gnd.n2511 10.8348
R17043 gnd.n4404 gnd.n2520 10.8348
R17044 gnd.n6387 gnd.n2523 10.8348
R17045 gnd.n4412 gnd.n2531 10.8348
R17046 gnd.n6381 gnd.n2534 10.8348
R17047 gnd.n4437 gnd.n4436 10.8348
R17048 gnd.n6375 gnd.n2543 10.8348
R17049 gnd.n4419 gnd.n2551 10.8348
R17050 gnd.n6369 gnd.n2554 10.8348
R17051 gnd.n4425 gnd.n2561 10.8348
R17052 gnd.n6363 gnd.n2564 10.8348
R17053 gnd.n6350 gnd.n2571 10.8348
R17054 gnd.n6357 gnd.n2574 10.8348
R17055 gnd.n4586 gnd.n4585 10.8348
R17056 gnd.n4653 gnd.t22 10.8348
R17057 gnd.n4774 gnd.n3616 10.8348
R17058 gnd.n4787 gnd.n3616 10.8348
R17059 gnd.n4930 gnd.n3530 10.8348
R17060 gnd.n4951 gnd.n3530 10.8348
R17061 gnd.n5020 gnd.t29 10.8348
R17062 gnd.n5097 gnd.n5095 10.8348
R17063 gnd.n6002 gnd.n6001 10.8348
R17064 gnd.n5195 gnd.n3059 10.8348
R17065 gnd.n5995 gnd.n3068 10.8348
R17066 gnd.n5730 gnd.n3071 10.8348
R17067 gnd.n5989 gnd.n3080 10.8348
R17068 gnd.n5738 gnd.n3083 10.8348
R17069 gnd.n5983 gnd.n3091 10.8348
R17070 gnd.n5759 gnd.n5758 10.8348
R17071 gnd.n5977 gnd.n3100 10.8348
R17072 gnd.n5747 gnd.n3103 10.8348
R17073 gnd.n5971 gnd.n3111 10.8348
R17074 gnd.n5803 gnd.n3114 10.8348
R17075 gnd.n5810 gnd.n3123 10.8348
R17076 gnd.n5959 gnd.n3131 10.8348
R17077 gnd.n5828 gnd.n3241 10.8348
R17078 gnd.n5953 gnd.n3140 10.8348
R17079 gnd.n5949 gnd.n3143 10.8348
R17080 gnd.n5948 gnd.n3149 10.8348
R17081 gnd.n3156 gnd.n3155 10.8348
R17082 gnd.n5935 gnd.n3159 10.8348
R17083 gnd.n5845 gnd.n3166 10.8348
R17084 gnd.n7731 gnd.n69 10.8348
R17085 gnd.n5928 gnd.n71 10.8348
R17086 gnd.n7723 gnd.n86 10.8348
R17087 gnd.n5861 gnd.n89 10.8348
R17088 gnd.n7717 gnd.n98 10.8348
R17089 gnd.n5870 gnd.n101 10.8348
R17090 gnd.n7711 gnd.n108 10.8348
R17091 gnd.n5914 gnd.n5913 10.8348
R17092 gnd.n7705 gnd.n117 10.8348
R17093 gnd.n7699 gnd.n128 10.8348
R17094 gnd.n5901 gnd.n131 10.8348
R17095 gnd.n7693 gnd.n138 10.8348
R17096 gnd.n5895 gnd.n141 10.8348
R17097 gnd.n7687 gnd.n149 10.8348
R17098 gnd.n5889 gnd.n152 10.8348
R17099 gnd.n7681 gnd.n159 10.8348
R17100 gnd.n7668 gnd.n176 10.8348
R17101 gnd.n7675 gnd.n168 10.8348
R17102 gnd.n3270 gnd.n3269 10.6672
R17103 gnd.n7545 gnd.n7542 10.6672
R17104 gnd.n4004 gnd.n4003 10.6672
R17105 gnd.n2789 gnd.n2786 10.6672
R17106 gnd.n5537 gnd.n3299 10.6151
R17107 gnd.n5537 gnd.n5536 10.6151
R17108 gnd.n5534 gnd.n5531 10.6151
R17109 gnd.n5531 gnd.n5530 10.6151
R17110 gnd.n5530 gnd.n5527 10.6151
R17111 gnd.n5527 gnd.n5526 10.6151
R17112 gnd.n5526 gnd.n5523 10.6151
R17113 gnd.n5523 gnd.n5522 10.6151
R17114 gnd.n5522 gnd.n5519 10.6151
R17115 gnd.n5519 gnd.n5518 10.6151
R17116 gnd.n5518 gnd.n5515 10.6151
R17117 gnd.n5515 gnd.n5514 10.6151
R17118 gnd.n5514 gnd.n5511 10.6151
R17119 gnd.n5511 gnd.n5510 10.6151
R17120 gnd.n5510 gnd.n5507 10.6151
R17121 gnd.n5507 gnd.n5506 10.6151
R17122 gnd.n5506 gnd.n5503 10.6151
R17123 gnd.n5503 gnd.n5502 10.6151
R17124 gnd.n5502 gnd.n5499 10.6151
R17125 gnd.n5499 gnd.n5498 10.6151
R17126 gnd.n5498 gnd.n5495 10.6151
R17127 gnd.n5495 gnd.n5494 10.6151
R17128 gnd.n5494 gnd.n5491 10.6151
R17129 gnd.n5491 gnd.n5490 10.6151
R17130 gnd.n5490 gnd.n5487 10.6151
R17131 gnd.n5487 gnd.n5486 10.6151
R17132 gnd.n5486 gnd.n5483 10.6151
R17133 gnd.n5483 gnd.n5482 10.6151
R17134 gnd.n5482 gnd.n5479 10.6151
R17135 gnd.n5479 gnd.n5478 10.6151
R17136 gnd.n3822 gnd.n3750 10.6151
R17137 gnd.n4503 gnd.n3750 10.6151
R17138 gnd.n4504 gnd.n4503 10.6151
R17139 gnd.n4505 gnd.n4504 10.6151
R17140 gnd.n4505 gnd.n3737 10.6151
R17141 gnd.n4520 gnd.n3737 10.6151
R17142 gnd.n4521 gnd.n4520 10.6151
R17143 gnd.n4522 gnd.n4521 10.6151
R17144 gnd.n4531 gnd.n4522 10.6151
R17145 gnd.n4531 gnd.n4530 10.6151
R17146 gnd.n4530 gnd.n4529 10.6151
R17147 gnd.n4529 gnd.n4524 10.6151
R17148 gnd.n4524 gnd.n4523 10.6151
R17149 gnd.n4523 gnd.n3716 10.6151
R17150 gnd.n4570 gnd.n3716 10.6151
R17151 gnd.n4571 gnd.n4570 10.6151
R17152 gnd.n4583 gnd.n4571 10.6151
R17153 gnd.n4583 gnd.n4582 10.6151
R17154 gnd.n4582 gnd.n4581 10.6151
R17155 gnd.n4581 gnd.n4579 10.6151
R17156 gnd.n4579 gnd.n4578 10.6151
R17157 gnd.n4578 gnd.n4575 10.6151
R17158 gnd.n4575 gnd.n4574 10.6151
R17159 gnd.n4574 gnd.n3681 10.6151
R17160 gnd.n4642 gnd.n3681 10.6151
R17161 gnd.n4643 gnd.n4642 10.6151
R17162 gnd.n4665 gnd.n4643 10.6151
R17163 gnd.n4665 gnd.n4664 10.6151
R17164 gnd.n4664 gnd.n4663 10.6151
R17165 gnd.n4663 gnd.n4659 10.6151
R17166 gnd.n4659 gnd.n4658 10.6151
R17167 gnd.n4658 gnd.n4656 10.6151
R17168 gnd.n4656 gnd.n4655 10.6151
R17169 gnd.n4655 gnd.n4651 10.6151
R17170 gnd.n4651 gnd.n4650 10.6151
R17171 gnd.n4650 gnd.n4648 10.6151
R17172 gnd.n4648 gnd.n4647 10.6151
R17173 gnd.n4647 gnd.n4644 10.6151
R17174 gnd.n4644 gnd.n3628 10.6151
R17175 gnd.n4767 gnd.n3628 10.6151
R17176 gnd.n4768 gnd.n4767 10.6151
R17177 gnd.n4772 gnd.n4768 10.6151
R17178 gnd.n4772 gnd.n4771 10.6151
R17179 gnd.n4771 gnd.n4770 10.6151
R17180 gnd.n4770 gnd.n3611 10.6151
R17181 gnd.n4797 gnd.n3611 10.6151
R17182 gnd.n4798 gnd.n4797 10.6151
R17183 gnd.n4799 gnd.n4798 10.6151
R17184 gnd.n4799 gnd.n3596 10.6151
R17185 gnd.n4821 gnd.n3596 10.6151
R17186 gnd.n4822 gnd.n4821 10.6151
R17187 gnd.n4843 gnd.n4822 10.6151
R17188 gnd.n4843 gnd.n4842 10.6151
R17189 gnd.n4842 gnd.n4841 10.6151
R17190 gnd.n4841 gnd.n4838 10.6151
R17191 gnd.n4838 gnd.n4837 10.6151
R17192 gnd.n4837 gnd.n4835 10.6151
R17193 gnd.n4835 gnd.n4834 10.6151
R17194 gnd.n4834 gnd.n4830 10.6151
R17195 gnd.n4830 gnd.n4829 10.6151
R17196 gnd.n4829 gnd.n4827 10.6151
R17197 gnd.n4827 gnd.n4826 10.6151
R17198 gnd.n4826 gnd.n4823 10.6151
R17199 gnd.n4823 gnd.n3542 10.6151
R17200 gnd.n4922 gnd.n3542 10.6151
R17201 gnd.n4923 gnd.n4922 10.6151
R17202 gnd.n4928 gnd.n4923 10.6151
R17203 gnd.n4928 gnd.n4927 10.6151
R17204 gnd.n4927 gnd.n4926 10.6151
R17205 gnd.n4926 gnd.n4924 10.6151
R17206 gnd.n4924 gnd.n3515 10.6151
R17207 gnd.n4974 gnd.n3515 10.6151
R17208 gnd.n4975 gnd.n4974 10.6151
R17209 gnd.n4996 gnd.n4975 10.6151
R17210 gnd.n4996 gnd.n4995 10.6151
R17211 gnd.n4995 gnd.n4994 10.6151
R17212 gnd.n4994 gnd.n4990 10.6151
R17213 gnd.n4990 gnd.n4989 10.6151
R17214 gnd.n4989 gnd.n4987 10.6151
R17215 gnd.n4987 gnd.n4986 10.6151
R17216 gnd.n4986 gnd.n4983 10.6151
R17217 gnd.n4983 gnd.n4982 10.6151
R17218 gnd.n4982 gnd.n4980 10.6151
R17219 gnd.n4980 gnd.n4979 10.6151
R17220 gnd.n4979 gnd.n4976 10.6151
R17221 gnd.n4976 gnd.n3466 10.6151
R17222 gnd.n5079 gnd.n3466 10.6151
R17223 gnd.n5080 gnd.n5079 10.6151
R17224 gnd.n5081 gnd.n5080 10.6151
R17225 gnd.n5081 gnd.n3427 10.6151
R17226 gnd.n5101 gnd.n3427 10.6151
R17227 gnd.n5101 gnd.n5100 10.6151
R17228 gnd.n5100 gnd.n5099 10.6151
R17229 gnd.n5099 gnd.n3457 10.6151
R17230 gnd.n3457 gnd.n3456 10.6151
R17231 gnd.n3456 gnd.n3454 10.6151
R17232 gnd.n3454 gnd.n3453 10.6151
R17233 gnd.n3453 gnd.n3449 10.6151
R17234 gnd.n3449 gnd.n3448 10.6151
R17235 gnd.n3448 gnd.n3446 10.6151
R17236 gnd.n3446 gnd.n3445 10.6151
R17237 gnd.n3445 gnd.n3443 10.6151
R17238 gnd.n3443 gnd.n3442 10.6151
R17239 gnd.n3442 gnd.n3441 10.6151
R17240 gnd.n3441 gnd.n3440 10.6151
R17241 gnd.n3440 gnd.n3439 10.6151
R17242 gnd.n3439 gnd.n3430 10.6151
R17243 gnd.n3430 gnd.n3429 10.6151
R17244 gnd.n3429 gnd.n3428 10.6151
R17245 gnd.n3428 gnd.n3338 10.6151
R17246 gnd.n3760 gnd.n2850 10.6151
R17247 gnd.n3763 gnd.n3760 10.6151
R17248 gnd.n3768 gnd.n3765 10.6151
R17249 gnd.n3769 gnd.n3768 10.6151
R17250 gnd.n3772 gnd.n3769 10.6151
R17251 gnd.n3773 gnd.n3772 10.6151
R17252 gnd.n3776 gnd.n3773 10.6151
R17253 gnd.n3777 gnd.n3776 10.6151
R17254 gnd.n3780 gnd.n3777 10.6151
R17255 gnd.n3781 gnd.n3780 10.6151
R17256 gnd.n3784 gnd.n3781 10.6151
R17257 gnd.n3785 gnd.n3784 10.6151
R17258 gnd.n3788 gnd.n3785 10.6151
R17259 gnd.n3789 gnd.n3788 10.6151
R17260 gnd.n3792 gnd.n3789 10.6151
R17261 gnd.n3793 gnd.n3792 10.6151
R17262 gnd.n3796 gnd.n3793 10.6151
R17263 gnd.n3797 gnd.n3796 10.6151
R17264 gnd.n3800 gnd.n3797 10.6151
R17265 gnd.n3801 gnd.n3800 10.6151
R17266 gnd.n3804 gnd.n3801 10.6151
R17267 gnd.n3805 gnd.n3804 10.6151
R17268 gnd.n3808 gnd.n3805 10.6151
R17269 gnd.n3809 gnd.n3808 10.6151
R17270 gnd.n3812 gnd.n3809 10.6151
R17271 gnd.n3813 gnd.n3812 10.6151
R17272 gnd.n3816 gnd.n3813 10.6151
R17273 gnd.n3817 gnd.n3816 10.6151
R17274 gnd.n3820 gnd.n3817 10.6151
R17275 gnd.n3821 gnd.n3820 10.6151
R17276 gnd.n6217 gnd.n6216 10.6151
R17277 gnd.n6216 gnd.n6215 10.6151
R17278 gnd.n6215 gnd.n6214 10.6151
R17279 gnd.n6214 gnd.n6212 10.6151
R17280 gnd.n6212 gnd.n6209 10.6151
R17281 gnd.n6209 gnd.n6208 10.6151
R17282 gnd.n6208 gnd.n6205 10.6151
R17283 gnd.n6205 gnd.n6204 10.6151
R17284 gnd.n6204 gnd.n6201 10.6151
R17285 gnd.n6201 gnd.n6200 10.6151
R17286 gnd.n6200 gnd.n6197 10.6151
R17287 gnd.n6197 gnd.n6196 10.6151
R17288 gnd.n6196 gnd.n6193 10.6151
R17289 gnd.n6193 gnd.n6192 10.6151
R17290 gnd.n6192 gnd.n6189 10.6151
R17291 gnd.n6189 gnd.n6188 10.6151
R17292 gnd.n6188 gnd.n6185 10.6151
R17293 gnd.n6185 gnd.n6184 10.6151
R17294 gnd.n6184 gnd.n6181 10.6151
R17295 gnd.n6181 gnd.n6180 10.6151
R17296 gnd.n6180 gnd.n6177 10.6151
R17297 gnd.n6177 gnd.n6176 10.6151
R17298 gnd.n6176 gnd.n6173 10.6151
R17299 gnd.n6173 gnd.n6172 10.6151
R17300 gnd.n6172 gnd.n6169 10.6151
R17301 gnd.n6169 gnd.n6168 10.6151
R17302 gnd.n6168 gnd.n6165 10.6151
R17303 gnd.n6165 gnd.n6164 10.6151
R17304 gnd.n6161 gnd.n6160 10.6151
R17305 gnd.n6160 gnd.n2851 10.6151
R17306 gnd.n5471 gnd.n5470 10.6151
R17307 gnd.n5470 gnd.n5467 10.6151
R17308 gnd.n5467 gnd.n5466 10.6151
R17309 gnd.n5466 gnd.n5463 10.6151
R17310 gnd.n5463 gnd.n5462 10.6151
R17311 gnd.n5462 gnd.n5459 10.6151
R17312 gnd.n5459 gnd.n5458 10.6151
R17313 gnd.n5458 gnd.n5455 10.6151
R17314 gnd.n5455 gnd.n5454 10.6151
R17315 gnd.n5454 gnd.n5451 10.6151
R17316 gnd.n5451 gnd.n5450 10.6151
R17317 gnd.n5450 gnd.n5447 10.6151
R17318 gnd.n5447 gnd.n5446 10.6151
R17319 gnd.n5446 gnd.n5443 10.6151
R17320 gnd.n5443 gnd.n5442 10.6151
R17321 gnd.n5442 gnd.n5439 10.6151
R17322 gnd.n5439 gnd.n5438 10.6151
R17323 gnd.n5438 gnd.n5435 10.6151
R17324 gnd.n5435 gnd.n5434 10.6151
R17325 gnd.n5434 gnd.n5431 10.6151
R17326 gnd.n5431 gnd.n5430 10.6151
R17327 gnd.n5430 gnd.n5427 10.6151
R17328 gnd.n5427 gnd.n5426 10.6151
R17329 gnd.n5426 gnd.n5423 10.6151
R17330 gnd.n5423 gnd.n5422 10.6151
R17331 gnd.n5422 gnd.n5419 10.6151
R17332 gnd.n5419 gnd.n5418 10.6151
R17333 gnd.n5418 gnd.n5415 10.6151
R17334 gnd.n5413 gnd.n5410 10.6151
R17335 gnd.n5410 gnd.n3300 10.6151
R17336 gnd.n6153 gnd.n6152 10.6151
R17337 gnd.n6152 gnd.n2910 10.6151
R17338 gnd.n3745 gnd.n2910 10.6151
R17339 gnd.n3745 gnd.n2928 10.6151
R17340 gnd.n6140 gnd.n2928 10.6151
R17341 gnd.n6140 gnd.n6139 10.6151
R17342 gnd.n6139 gnd.n6138 10.6151
R17343 gnd.n6138 gnd.n2929 10.6151
R17344 gnd.n4537 gnd.n2929 10.6151
R17345 gnd.n4537 gnd.n4536 10.6151
R17346 gnd.n4536 gnd.n4535 10.6151
R17347 gnd.n4535 gnd.n3722 10.6151
R17348 gnd.n4563 gnd.n3722 10.6151
R17349 gnd.n4564 gnd.n4563 10.6151
R17350 gnd.n4566 gnd.n4564 10.6151
R17351 gnd.n4566 gnd.n4565 10.6151
R17352 gnd.n4565 gnd.n3704 10.6151
R17353 gnd.n4601 gnd.n3704 10.6151
R17354 gnd.n4602 gnd.n4601 10.6151
R17355 gnd.n4603 gnd.n4602 10.6151
R17356 gnd.n4603 gnd.n3692 10.6151
R17357 gnd.n4628 gnd.n3692 10.6151
R17358 gnd.n4628 gnd.n4627 10.6151
R17359 gnd.n4627 gnd.n4626 10.6151
R17360 gnd.n4626 gnd.n3677 10.6151
R17361 gnd.n4671 gnd.n3677 10.6151
R17362 gnd.n4672 gnd.n4671 10.6151
R17363 gnd.n4673 gnd.n4672 10.6151
R17364 gnd.n4673 gnd.n3663 10.6151
R17365 gnd.n4690 gnd.n3663 10.6151
R17366 gnd.n4691 gnd.n4690 10.6151
R17367 gnd.n4692 gnd.n4691 10.6151
R17368 gnd.n4692 gnd.n3650 10.6151
R17369 gnd.n4742 gnd.n3650 10.6151
R17370 gnd.n4743 gnd.n4742 10.6151
R17371 gnd.n4744 gnd.n4743 10.6151
R17372 gnd.n4744 gnd.n3634 10.6151
R17373 gnd.n4760 gnd.n3634 10.6151
R17374 gnd.n4761 gnd.n4760 10.6151
R17375 gnd.n4763 gnd.n4761 10.6151
R17376 gnd.n4763 gnd.n4762 10.6151
R17377 gnd.n4762 gnd.n3614 10.6151
R17378 gnd.n4789 gnd.n3614 10.6151
R17379 gnd.n4790 gnd.n4789 10.6151
R17380 gnd.n4791 gnd.n4790 10.6151
R17381 gnd.n4791 gnd.n3610 10.6151
R17382 gnd.n4807 gnd.n3610 10.6151
R17383 gnd.n4807 gnd.n4806 10.6151
R17384 gnd.n4806 gnd.n4805 10.6151
R17385 gnd.n4805 gnd.n3592 10.6151
R17386 gnd.n4849 gnd.n3592 10.6151
R17387 gnd.n4850 gnd.n4849 10.6151
R17388 gnd.n4851 gnd.n4850 10.6151
R17389 gnd.n4851 gnd.n3577 10.6151
R17390 gnd.n4867 gnd.n3577 10.6151
R17391 gnd.n4868 gnd.n4867 10.6151
R17392 gnd.n4869 gnd.n4868 10.6151
R17393 gnd.n4869 gnd.n3563 10.6151
R17394 gnd.n4898 gnd.n3563 10.6151
R17395 gnd.n4899 gnd.n4898 10.6151
R17396 gnd.n4900 gnd.n4899 10.6151
R17397 gnd.n4900 gnd.n3547 10.6151
R17398 gnd.n4915 gnd.n3547 10.6151
R17399 gnd.n4916 gnd.n4915 10.6151
R17400 gnd.n4918 gnd.n4916 10.6151
R17401 gnd.n4918 gnd.n4917 10.6151
R17402 gnd.n4917 gnd.n3528 10.6151
R17403 gnd.n4953 gnd.n3528 10.6151
R17404 gnd.n4954 gnd.n4953 10.6151
R17405 gnd.n4956 gnd.n4954 10.6151
R17406 gnd.n4956 gnd.n4955 10.6151
R17407 gnd.n4955 gnd.n3512 10.6151
R17408 gnd.n5002 gnd.n3512 10.6151
R17409 gnd.n5003 gnd.n5002 10.6151
R17410 gnd.n5004 gnd.n5003 10.6151
R17411 gnd.n5004 gnd.n3499 10.6151
R17412 gnd.n5022 gnd.n3499 10.6151
R17413 gnd.n5023 gnd.n5022 10.6151
R17414 gnd.n5024 gnd.n5023 10.6151
R17415 gnd.n5024 gnd.n3485 10.6151
R17416 gnd.n5052 gnd.n3485 10.6151
R17417 gnd.n5053 gnd.n5052 10.6151
R17418 gnd.n5054 gnd.n5053 10.6151
R17419 gnd.n5054 gnd.n3471 10.6151
R17420 gnd.n5072 gnd.n3471 10.6151
R17421 gnd.n5073 gnd.n5072 10.6151
R17422 gnd.n5075 gnd.n5073 10.6151
R17423 gnd.n5075 gnd.n5074 10.6151
R17424 gnd.n5074 gnd.n3423 10.6151
R17425 gnd.n5107 gnd.n3423 10.6151
R17426 gnd.n5108 gnd.n5107 10.6151
R17427 gnd.n5109 gnd.n5108 10.6151
R17428 gnd.n5109 gnd.n3409 10.6151
R17429 gnd.n5125 gnd.n3409 10.6151
R17430 gnd.n5126 gnd.n5125 10.6151
R17431 gnd.n5127 gnd.n5126 10.6151
R17432 gnd.n5127 gnd.n3396 10.6151
R17433 gnd.n5141 gnd.n3396 10.6151
R17434 gnd.n5142 gnd.n5141 10.6151
R17435 gnd.n5144 gnd.n5142 10.6151
R17436 gnd.n5144 gnd.n5143 10.6151
R17437 gnd.n5143 gnd.n3372 10.6151
R17438 gnd.n5174 gnd.n3372 10.6151
R17439 gnd.n5175 gnd.n5174 10.6151
R17440 gnd.n5177 gnd.n5175 10.6151
R17441 gnd.n5177 gnd.n5176 10.6151
R17442 gnd.n5176 gnd.n3343 10.6151
R17443 gnd.n5387 gnd.n3343 10.6151
R17444 gnd.n5388 gnd.n5387 10.6151
R17445 gnd.n5473 gnd.n5388 10.6151
R17446 gnd.n1556 gnd.t187 10.5161
R17447 gnd.n1003 gnd.t168 10.5161
R17448 gnd.n1924 gnd.t172 10.5161
R17449 gnd.t220 gnd.n2457 10.5161
R17450 gnd.n4355 gnd.t264 10.5161
R17451 gnd.n6425 gnd.t264 10.5161
R17452 gnd.n6418 gnd.t253 10.5161
R17453 gnd.t229 gnd.n5940 10.5161
R17454 gnd.n5845 gnd.t244 10.5161
R17455 gnd.t244 gnd.n69 10.5161
R17456 gnd.n5927 gnd.t194 10.5161
R17457 gnd.n2200 gnd.n2184 10.4732
R17458 gnd.n2168 gnd.n2152 10.4732
R17459 gnd.n2136 gnd.n2120 10.4732
R17460 gnd.n2105 gnd.n2089 10.4732
R17461 gnd.n2073 gnd.n2057 10.4732
R17462 gnd.n2041 gnd.n2025 10.4732
R17463 gnd.n2009 gnd.n1993 10.4732
R17464 gnd.n1978 gnd.n1962 10.4732
R17465 gnd.n6488 gnd.n2363 10.1975
R17466 gnd.n4508 gnd.n4507 10.1975
R17467 gnd.n4518 gnd.n4517 10.1975
R17468 gnd.n4661 gnd.n3675 10.1975
R17469 gnd.n4839 gnd.n3590 10.1975
R17470 gnd.n4872 gnd.n3573 10.1975
R17471 gnd.n5050 gnd.n5049 10.1975
R17472 gnd.n5171 gnd.n5170 10.1975
R17473 gnd.n3437 gnd.n3436 10.1975
R17474 gnd.n7659 gnd.n184 10.1975
R17475 gnd.t171 gnd.n1020 9.87883
R17476 gnd.t240 gnd.n2418 9.87883
R17477 gnd.n6450 gnd.t227 9.87883
R17478 gnd.n4389 gnd.t201 9.87883
R17479 gnd.n6393 gnd.t233 9.87883
R17480 gnd.n5965 gnd.t205 9.87883
R17481 gnd.n3241 gnd.t222 9.87883
R17482 gnd.n7711 gnd.t260 9.87883
R17483 gnd.t198 gnd.n120 9.87883
R17484 gnd.n2204 gnd.n2203 9.69747
R17485 gnd.n2172 gnd.n2171 9.69747
R17486 gnd.n2140 gnd.n2139 9.69747
R17487 gnd.n2109 gnd.n2108 9.69747
R17488 gnd.n2077 gnd.n2076 9.69747
R17489 gnd.n2045 gnd.n2044 9.69747
R17490 gnd.n2013 gnd.n2012 9.69747
R17491 gnd.n1982 gnd.n1981 9.69747
R17492 gnd.n4568 gnd.n3718 9.56018
R17493 gnd.n4605 gnd.n3702 9.56018
R17494 gnd.n4765 gnd.n3630 9.56018
R17495 gnd.n3631 gnd.t184 9.56018
R17496 gnd.n4794 gnd.n4793 9.56018
R17497 gnd.n4920 gnd.n3544 9.56018
R17498 gnd.n4959 gnd.t190 9.56018
R17499 gnd.n4958 gnd.n3525 9.56018
R17500 gnd.n5105 gnd.n3425 9.56018
R17501 gnd.n5130 gnd.n3405 9.56018
R17502 gnd.n2210 gnd.n2209 9.45567
R17503 gnd.n2178 gnd.n2177 9.45567
R17504 gnd.n2146 gnd.n2145 9.45567
R17505 gnd.n2115 gnd.n2114 9.45567
R17506 gnd.n2083 gnd.n2082 9.45567
R17507 gnd.n2051 gnd.n2050 9.45567
R17508 gnd.n2019 gnd.n2018 9.45567
R17509 gnd.n1988 gnd.n1987 9.45567
R17510 gnd.n5668 gnd.n3288 9.30959
R17511 gnd.n7584 gnd.n7516 9.30959
R17512 gnd.n4158 gnd.n4022 9.30959
R17513 gnd.n2828 gnd.n2760 9.30959
R17514 gnd.n2209 gnd.n2208 9.3005
R17515 gnd.n2182 gnd.n2181 9.3005
R17516 gnd.n2203 gnd.n2202 9.3005
R17517 gnd.n2201 gnd.n2200 9.3005
R17518 gnd.n2186 gnd.n2185 9.3005
R17519 gnd.n2195 gnd.n2194 9.3005
R17520 gnd.n2193 gnd.n2192 9.3005
R17521 gnd.n2177 gnd.n2176 9.3005
R17522 gnd.n2150 gnd.n2149 9.3005
R17523 gnd.n2171 gnd.n2170 9.3005
R17524 gnd.n2169 gnd.n2168 9.3005
R17525 gnd.n2154 gnd.n2153 9.3005
R17526 gnd.n2163 gnd.n2162 9.3005
R17527 gnd.n2161 gnd.n2160 9.3005
R17528 gnd.n2145 gnd.n2144 9.3005
R17529 gnd.n2118 gnd.n2117 9.3005
R17530 gnd.n2139 gnd.n2138 9.3005
R17531 gnd.n2137 gnd.n2136 9.3005
R17532 gnd.n2122 gnd.n2121 9.3005
R17533 gnd.n2131 gnd.n2130 9.3005
R17534 gnd.n2129 gnd.n2128 9.3005
R17535 gnd.n2114 gnd.n2113 9.3005
R17536 gnd.n2087 gnd.n2086 9.3005
R17537 gnd.n2108 gnd.n2107 9.3005
R17538 gnd.n2106 gnd.n2105 9.3005
R17539 gnd.n2091 gnd.n2090 9.3005
R17540 gnd.n2100 gnd.n2099 9.3005
R17541 gnd.n2098 gnd.n2097 9.3005
R17542 gnd.n2082 gnd.n2081 9.3005
R17543 gnd.n2055 gnd.n2054 9.3005
R17544 gnd.n2076 gnd.n2075 9.3005
R17545 gnd.n2074 gnd.n2073 9.3005
R17546 gnd.n2059 gnd.n2058 9.3005
R17547 gnd.n2068 gnd.n2067 9.3005
R17548 gnd.n2066 gnd.n2065 9.3005
R17549 gnd.n2050 gnd.n2049 9.3005
R17550 gnd.n2023 gnd.n2022 9.3005
R17551 gnd.n2044 gnd.n2043 9.3005
R17552 gnd.n2042 gnd.n2041 9.3005
R17553 gnd.n2027 gnd.n2026 9.3005
R17554 gnd.n2036 gnd.n2035 9.3005
R17555 gnd.n2034 gnd.n2033 9.3005
R17556 gnd.n2018 gnd.n2017 9.3005
R17557 gnd.n1991 gnd.n1990 9.3005
R17558 gnd.n2012 gnd.n2011 9.3005
R17559 gnd.n2010 gnd.n2009 9.3005
R17560 gnd.n1995 gnd.n1994 9.3005
R17561 gnd.n2004 gnd.n2003 9.3005
R17562 gnd.n2002 gnd.n2001 9.3005
R17563 gnd.n1987 gnd.n1986 9.3005
R17564 gnd.n1960 gnd.n1959 9.3005
R17565 gnd.n1981 gnd.n1980 9.3005
R17566 gnd.n1979 gnd.n1978 9.3005
R17567 gnd.n1964 gnd.n1963 9.3005
R17568 gnd.n1973 gnd.n1972 9.3005
R17569 gnd.n1971 gnd.n1970 9.3005
R17570 gnd.n2335 gnd.n2334 9.3005
R17571 gnd.n2333 gnd.n903 9.3005
R17572 gnd.n2332 gnd.n2331 9.3005
R17573 gnd.n2328 gnd.n904 9.3005
R17574 gnd.n2325 gnd.n905 9.3005
R17575 gnd.n2324 gnd.n906 9.3005
R17576 gnd.n2321 gnd.n907 9.3005
R17577 gnd.n2320 gnd.n908 9.3005
R17578 gnd.n2317 gnd.n909 9.3005
R17579 gnd.n2316 gnd.n910 9.3005
R17580 gnd.n2313 gnd.n911 9.3005
R17581 gnd.n2312 gnd.n912 9.3005
R17582 gnd.n2309 gnd.n913 9.3005
R17583 gnd.n2308 gnd.n914 9.3005
R17584 gnd.n2305 gnd.n2304 9.3005
R17585 gnd.n2303 gnd.n915 9.3005
R17586 gnd.n2336 gnd.n902 9.3005
R17587 gnd.n1575 gnd.n1574 9.3005
R17588 gnd.n1279 gnd.n1278 9.3005
R17589 gnd.n1602 gnd.n1601 9.3005
R17590 gnd.n1603 gnd.n1277 9.3005
R17591 gnd.n1607 gnd.n1604 9.3005
R17592 gnd.n1606 gnd.n1605 9.3005
R17593 gnd.n1251 gnd.n1250 9.3005
R17594 gnd.n1632 gnd.n1631 9.3005
R17595 gnd.n1633 gnd.n1249 9.3005
R17596 gnd.n1635 gnd.n1634 9.3005
R17597 gnd.n1229 gnd.n1228 9.3005
R17598 gnd.n1663 gnd.n1662 9.3005
R17599 gnd.n1664 gnd.n1227 9.3005
R17600 gnd.n1672 gnd.n1665 9.3005
R17601 gnd.n1671 gnd.n1666 9.3005
R17602 gnd.n1670 gnd.n1668 9.3005
R17603 gnd.n1667 gnd.n1176 9.3005
R17604 gnd.n1720 gnd.n1177 9.3005
R17605 gnd.n1719 gnd.n1178 9.3005
R17606 gnd.n1718 gnd.n1179 9.3005
R17607 gnd.n1198 gnd.n1180 9.3005
R17608 gnd.n1200 gnd.n1199 9.3005
R17609 gnd.n1098 gnd.n1097 9.3005
R17610 gnd.n1758 gnd.n1757 9.3005
R17611 gnd.n1759 gnd.n1096 9.3005
R17612 gnd.n1763 gnd.n1760 9.3005
R17613 gnd.n1762 gnd.n1761 9.3005
R17614 gnd.n1071 gnd.n1070 9.3005
R17615 gnd.n1798 gnd.n1797 9.3005
R17616 gnd.n1799 gnd.n1069 9.3005
R17617 gnd.n1803 gnd.n1800 9.3005
R17618 gnd.n1802 gnd.n1801 9.3005
R17619 gnd.n1045 gnd.n1044 9.3005
R17620 gnd.n1845 gnd.n1844 9.3005
R17621 gnd.n1846 gnd.n1043 9.3005
R17622 gnd.n1850 gnd.n1847 9.3005
R17623 gnd.n1849 gnd.n1848 9.3005
R17624 gnd.n1018 gnd.n1017 9.3005
R17625 gnd.n1885 gnd.n1884 9.3005
R17626 gnd.n1886 gnd.n1016 9.3005
R17627 gnd.n1890 gnd.n1887 9.3005
R17628 gnd.n1889 gnd.n1888 9.3005
R17629 gnd.n991 gnd.n990 9.3005
R17630 gnd.n1934 gnd.n1933 9.3005
R17631 gnd.n1935 gnd.n989 9.3005
R17632 gnd.n1939 gnd.n1936 9.3005
R17633 gnd.n1938 gnd.n1937 9.3005
R17634 gnd.n964 gnd.n963 9.3005
R17635 gnd.n2228 gnd.n2227 9.3005
R17636 gnd.n2229 gnd.n962 9.3005
R17637 gnd.n2235 gnd.n2230 9.3005
R17638 gnd.n2234 gnd.n2231 9.3005
R17639 gnd.n2233 gnd.n2232 9.3005
R17640 gnd.n1576 gnd.n1573 9.3005
R17641 gnd.n1358 gnd.n1317 9.3005
R17642 gnd.n1353 gnd.n1352 9.3005
R17643 gnd.n1351 gnd.n1318 9.3005
R17644 gnd.n1350 gnd.n1349 9.3005
R17645 gnd.n1346 gnd.n1319 9.3005
R17646 gnd.n1343 gnd.n1342 9.3005
R17647 gnd.n1341 gnd.n1320 9.3005
R17648 gnd.n1340 gnd.n1339 9.3005
R17649 gnd.n1336 gnd.n1321 9.3005
R17650 gnd.n1333 gnd.n1332 9.3005
R17651 gnd.n1331 gnd.n1322 9.3005
R17652 gnd.n1330 gnd.n1329 9.3005
R17653 gnd.n1326 gnd.n1324 9.3005
R17654 gnd.n1323 gnd.n1303 9.3005
R17655 gnd.n1570 gnd.n1302 9.3005
R17656 gnd.n1572 gnd.n1571 9.3005
R17657 gnd.n1360 gnd.n1359 9.3005
R17658 gnd.n1583 gnd.n1289 9.3005
R17659 gnd.n1590 gnd.n1290 9.3005
R17660 gnd.n1592 gnd.n1591 9.3005
R17661 gnd.n1593 gnd.n1270 9.3005
R17662 gnd.n1612 gnd.n1611 9.3005
R17663 gnd.n1614 gnd.n1262 9.3005
R17664 gnd.n1621 gnd.n1264 9.3005
R17665 gnd.n1622 gnd.n1259 9.3005
R17666 gnd.n1624 gnd.n1623 9.3005
R17667 gnd.n1260 gnd.n1245 9.3005
R17668 gnd.n1640 gnd.n1243 9.3005
R17669 gnd.n1644 gnd.n1643 9.3005
R17670 gnd.n1642 gnd.n1219 9.3005
R17671 gnd.n1679 gnd.n1218 9.3005
R17672 gnd.n1682 gnd.n1681 9.3005
R17673 gnd.n1215 gnd.n1214 9.3005
R17674 gnd.n1688 gnd.n1216 9.3005
R17675 gnd.n1690 gnd.n1689 9.3005
R17676 gnd.n1692 gnd.n1213 9.3005
R17677 gnd.n1695 gnd.n1694 9.3005
R17678 gnd.n1698 gnd.n1696 9.3005
R17679 gnd.n1700 gnd.n1699 9.3005
R17680 gnd.n1706 gnd.n1701 9.3005
R17681 gnd.n1705 gnd.n1704 9.3005
R17682 gnd.n1089 gnd.n1088 9.3005
R17683 gnd.n1772 gnd.n1771 9.3005
R17684 gnd.n1773 gnd.n1082 9.3005
R17685 gnd.n1781 gnd.n1081 9.3005
R17686 gnd.n1784 gnd.n1783 9.3005
R17687 gnd.n1786 gnd.n1785 9.3005
R17688 gnd.n1789 gnd.n1064 9.3005
R17689 gnd.n1787 gnd.n1062 9.3005
R17690 gnd.n1809 gnd.n1060 9.3005
R17691 gnd.n1811 gnd.n1810 9.3005
R17692 gnd.n1036 gnd.n1035 9.3005
R17693 gnd.n1859 gnd.n1858 9.3005
R17694 gnd.n1860 gnd.n1029 9.3005
R17695 gnd.n1868 gnd.n1028 9.3005
R17696 gnd.n1871 gnd.n1870 9.3005
R17697 gnd.n1873 gnd.n1872 9.3005
R17698 gnd.n1876 gnd.n1011 9.3005
R17699 gnd.n1874 gnd.n1009 9.3005
R17700 gnd.n1896 gnd.n1007 9.3005
R17701 gnd.n1898 gnd.n1897 9.3005
R17702 gnd.n982 gnd.n981 9.3005
R17703 gnd.n1948 gnd.n1947 9.3005
R17704 gnd.n1949 gnd.n975 9.3005
R17705 gnd.n1957 gnd.n974 9.3005
R17706 gnd.n2216 gnd.n2215 9.3005
R17707 gnd.n2218 gnd.n2217 9.3005
R17708 gnd.n2219 gnd.n955 9.3005
R17709 gnd.n2243 gnd.n2242 9.3005
R17710 gnd.n956 gnd.n918 9.3005
R17711 gnd.n1581 gnd.n1580 9.3005
R17712 gnd.n2299 gnd.n919 9.3005
R17713 gnd.n2298 gnd.n921 9.3005
R17714 gnd.n2295 gnd.n922 9.3005
R17715 gnd.n2294 gnd.n923 9.3005
R17716 gnd.n2291 gnd.n924 9.3005
R17717 gnd.n2290 gnd.n925 9.3005
R17718 gnd.n2287 gnd.n926 9.3005
R17719 gnd.n2286 gnd.n927 9.3005
R17720 gnd.n2283 gnd.n928 9.3005
R17721 gnd.n2282 gnd.n929 9.3005
R17722 gnd.n2279 gnd.n930 9.3005
R17723 gnd.n2278 gnd.n931 9.3005
R17724 gnd.n2275 gnd.n932 9.3005
R17725 gnd.n2274 gnd.n933 9.3005
R17726 gnd.n2271 gnd.n934 9.3005
R17727 gnd.n2270 gnd.n935 9.3005
R17728 gnd.n2267 gnd.n936 9.3005
R17729 gnd.n2266 gnd.n937 9.3005
R17730 gnd.n2263 gnd.n938 9.3005
R17731 gnd.n2262 gnd.n939 9.3005
R17732 gnd.n2259 gnd.n940 9.3005
R17733 gnd.n2258 gnd.n941 9.3005
R17734 gnd.n2255 gnd.n945 9.3005
R17735 gnd.n2254 gnd.n946 9.3005
R17736 gnd.n2251 gnd.n947 9.3005
R17737 gnd.n2250 gnd.n948 9.3005
R17738 gnd.n2301 gnd.n2300 9.3005
R17739 gnd.n1750 gnd.n1734 9.3005
R17740 gnd.n1749 gnd.n1735 9.3005
R17741 gnd.n1748 gnd.n1736 9.3005
R17742 gnd.n1746 gnd.n1737 9.3005
R17743 gnd.n1745 gnd.n1738 9.3005
R17744 gnd.n1743 gnd.n1739 9.3005
R17745 gnd.n1742 gnd.n1740 9.3005
R17746 gnd.n1052 gnd.n1051 9.3005
R17747 gnd.n1819 gnd.n1818 9.3005
R17748 gnd.n1820 gnd.n1050 9.3005
R17749 gnd.n1837 gnd.n1821 9.3005
R17750 gnd.n1836 gnd.n1822 9.3005
R17751 gnd.n1835 gnd.n1823 9.3005
R17752 gnd.n1833 gnd.n1824 9.3005
R17753 gnd.n1832 gnd.n1825 9.3005
R17754 gnd.n1830 gnd.n1826 9.3005
R17755 gnd.n1829 gnd.n1827 9.3005
R17756 gnd.n998 gnd.n997 9.3005
R17757 gnd.n1906 gnd.n1905 9.3005
R17758 gnd.n1907 gnd.n996 9.3005
R17759 gnd.n1928 gnd.n1908 9.3005
R17760 gnd.n1927 gnd.n1909 9.3005
R17761 gnd.n1926 gnd.n1910 9.3005
R17762 gnd.n1923 gnd.n1911 9.3005
R17763 gnd.n1922 gnd.n1912 9.3005
R17764 gnd.n1920 gnd.n1913 9.3005
R17765 gnd.n1919 gnd.n1914 9.3005
R17766 gnd.n1917 gnd.n1916 9.3005
R17767 gnd.n1915 gnd.n950 9.3005
R17768 gnd.n1491 gnd.n1490 9.3005
R17769 gnd.n1381 gnd.n1380 9.3005
R17770 gnd.n1505 gnd.n1504 9.3005
R17771 gnd.n1506 gnd.n1379 9.3005
R17772 gnd.n1508 gnd.n1507 9.3005
R17773 gnd.n1369 gnd.n1368 9.3005
R17774 gnd.n1521 gnd.n1520 9.3005
R17775 gnd.n1522 gnd.n1367 9.3005
R17776 gnd.n1554 gnd.n1523 9.3005
R17777 gnd.n1553 gnd.n1524 9.3005
R17778 gnd.n1552 gnd.n1525 9.3005
R17779 gnd.n1551 gnd.n1526 9.3005
R17780 gnd.n1548 gnd.n1527 9.3005
R17781 gnd.n1547 gnd.n1528 9.3005
R17782 gnd.n1546 gnd.n1529 9.3005
R17783 gnd.n1544 gnd.n1530 9.3005
R17784 gnd.n1543 gnd.n1531 9.3005
R17785 gnd.n1540 gnd.n1532 9.3005
R17786 gnd.n1539 gnd.n1533 9.3005
R17787 gnd.n1538 gnd.n1534 9.3005
R17788 gnd.n1536 gnd.n1535 9.3005
R17789 gnd.n1235 gnd.n1234 9.3005
R17790 gnd.n1652 gnd.n1651 9.3005
R17791 gnd.n1653 gnd.n1233 9.3005
R17792 gnd.n1657 gnd.n1654 9.3005
R17793 gnd.n1656 gnd.n1655 9.3005
R17794 gnd.n1157 gnd.n1156 9.3005
R17795 gnd.n1732 gnd.n1731 9.3005
R17796 gnd.n1489 gnd.n1390 9.3005
R17797 gnd.n1392 gnd.n1391 9.3005
R17798 gnd.n1436 gnd.n1434 9.3005
R17799 gnd.n1437 gnd.n1433 9.3005
R17800 gnd.n1440 gnd.n1429 9.3005
R17801 gnd.n1441 gnd.n1428 9.3005
R17802 gnd.n1444 gnd.n1427 9.3005
R17803 gnd.n1445 gnd.n1426 9.3005
R17804 gnd.n1448 gnd.n1425 9.3005
R17805 gnd.n1449 gnd.n1424 9.3005
R17806 gnd.n1452 gnd.n1423 9.3005
R17807 gnd.n1453 gnd.n1422 9.3005
R17808 gnd.n1456 gnd.n1421 9.3005
R17809 gnd.n1457 gnd.n1420 9.3005
R17810 gnd.n1460 gnd.n1419 9.3005
R17811 gnd.n1461 gnd.n1418 9.3005
R17812 gnd.n1464 gnd.n1417 9.3005
R17813 gnd.n1465 gnd.n1416 9.3005
R17814 gnd.n1468 gnd.n1415 9.3005
R17815 gnd.n1469 gnd.n1414 9.3005
R17816 gnd.n1472 gnd.n1413 9.3005
R17817 gnd.n1473 gnd.n1412 9.3005
R17818 gnd.n1476 gnd.n1411 9.3005
R17819 gnd.n1478 gnd.n1410 9.3005
R17820 gnd.n1479 gnd.n1409 9.3005
R17821 gnd.n1480 gnd.n1408 9.3005
R17822 gnd.n1481 gnd.n1407 9.3005
R17823 gnd.n1488 gnd.n1487 9.3005
R17824 gnd.n1497 gnd.n1496 9.3005
R17825 gnd.n1498 gnd.n1384 9.3005
R17826 gnd.n1500 gnd.n1499 9.3005
R17827 gnd.n1375 gnd.n1374 9.3005
R17828 gnd.n1513 gnd.n1512 9.3005
R17829 gnd.n1514 gnd.n1373 9.3005
R17830 gnd.n1516 gnd.n1515 9.3005
R17831 gnd.n1362 gnd.n1361 9.3005
R17832 gnd.n1559 gnd.n1558 9.3005
R17833 gnd.n1560 gnd.n1316 9.3005
R17834 gnd.n1564 gnd.n1562 9.3005
R17835 gnd.n1563 gnd.n1295 9.3005
R17836 gnd.n1582 gnd.n1294 9.3005
R17837 gnd.n1585 gnd.n1584 9.3005
R17838 gnd.n1288 gnd.n1287 9.3005
R17839 gnd.n1596 gnd.n1594 9.3005
R17840 gnd.n1595 gnd.n1269 9.3005
R17841 gnd.n1613 gnd.n1268 9.3005
R17842 gnd.n1616 gnd.n1615 9.3005
R17843 gnd.n1263 gnd.n1258 9.3005
R17844 gnd.n1626 gnd.n1625 9.3005
R17845 gnd.n1261 gnd.n1241 9.3005
R17846 gnd.n1647 gnd.n1242 9.3005
R17847 gnd.n1646 gnd.n1645 9.3005
R17848 gnd.n1244 gnd.n1220 9.3005
R17849 gnd.n1678 gnd.n1677 9.3005
R17850 gnd.n1680 gnd.n1165 9.3005
R17851 gnd.n1727 gnd.n1166 9.3005
R17852 gnd.n1726 gnd.n1167 9.3005
R17853 gnd.n1725 gnd.n1168 9.3005
R17854 gnd.n1691 gnd.n1169 9.3005
R17855 gnd.n1693 gnd.n1187 9.3005
R17856 gnd.n1713 gnd.n1188 9.3005
R17857 gnd.n1712 gnd.n1189 9.3005
R17858 gnd.n1711 gnd.n1190 9.3005
R17859 gnd.n1702 gnd.n1191 9.3005
R17860 gnd.n1703 gnd.n1090 9.3005
R17861 gnd.n1769 gnd.n1768 9.3005
R17862 gnd.n1770 gnd.n1083 9.3005
R17863 gnd.n1780 gnd.n1779 9.3005
R17864 gnd.n1782 gnd.n1079 9.3005
R17865 gnd.n1792 gnd.n1080 9.3005
R17866 gnd.n1791 gnd.n1790 9.3005
R17867 gnd.n1788 gnd.n1058 9.3005
R17868 gnd.n1814 gnd.n1059 9.3005
R17869 gnd.n1813 gnd.n1812 9.3005
R17870 gnd.n1061 gnd.n1037 9.3005
R17871 gnd.n1856 gnd.n1855 9.3005
R17872 gnd.n1857 gnd.n1030 9.3005
R17873 gnd.n1867 gnd.n1866 9.3005
R17874 gnd.n1869 gnd.n1026 9.3005
R17875 gnd.n1879 gnd.n1027 9.3005
R17876 gnd.n1878 gnd.n1877 9.3005
R17877 gnd.n1875 gnd.n1005 9.3005
R17878 gnd.n1901 gnd.n1006 9.3005
R17879 gnd.n1900 gnd.n1899 9.3005
R17880 gnd.n1008 gnd.n983 9.3005
R17881 gnd.n1945 gnd.n1944 9.3005
R17882 gnd.n1946 gnd.n976 9.3005
R17883 gnd.n1956 gnd.n1955 9.3005
R17884 gnd.n2214 gnd.n972 9.3005
R17885 gnd.n2222 gnd.n973 9.3005
R17886 gnd.n2221 gnd.n2220 9.3005
R17887 gnd.n954 gnd.n953 9.3005
R17888 gnd.n2245 gnd.n2244 9.3005
R17889 gnd.n1386 gnd.n1385 9.3005
R17890 gnd.n6688 gnd.n6687 9.3005
R17891 gnd.n703 gnd.n702 9.3005
R17892 gnd.n6695 gnd.n6694 9.3005
R17893 gnd.n6696 gnd.n701 9.3005
R17894 gnd.n6698 gnd.n6697 9.3005
R17895 gnd.n697 gnd.n696 9.3005
R17896 gnd.n6705 gnd.n6704 9.3005
R17897 gnd.n6706 gnd.n695 9.3005
R17898 gnd.n6708 gnd.n6707 9.3005
R17899 gnd.n691 gnd.n690 9.3005
R17900 gnd.n6715 gnd.n6714 9.3005
R17901 gnd.n6716 gnd.n689 9.3005
R17902 gnd.n6718 gnd.n6717 9.3005
R17903 gnd.n685 gnd.n684 9.3005
R17904 gnd.n6725 gnd.n6724 9.3005
R17905 gnd.n6726 gnd.n683 9.3005
R17906 gnd.n6728 gnd.n6727 9.3005
R17907 gnd.n679 gnd.n678 9.3005
R17908 gnd.n6735 gnd.n6734 9.3005
R17909 gnd.n6736 gnd.n677 9.3005
R17910 gnd.n6738 gnd.n6737 9.3005
R17911 gnd.n673 gnd.n672 9.3005
R17912 gnd.n6745 gnd.n6744 9.3005
R17913 gnd.n6746 gnd.n671 9.3005
R17914 gnd.n6748 gnd.n6747 9.3005
R17915 gnd.n667 gnd.n666 9.3005
R17916 gnd.n6755 gnd.n6754 9.3005
R17917 gnd.n6756 gnd.n665 9.3005
R17918 gnd.n6758 gnd.n6757 9.3005
R17919 gnd.n661 gnd.n660 9.3005
R17920 gnd.n6765 gnd.n6764 9.3005
R17921 gnd.n6766 gnd.n659 9.3005
R17922 gnd.n6768 gnd.n6767 9.3005
R17923 gnd.n655 gnd.n654 9.3005
R17924 gnd.n6775 gnd.n6774 9.3005
R17925 gnd.n6776 gnd.n653 9.3005
R17926 gnd.n6778 gnd.n6777 9.3005
R17927 gnd.n649 gnd.n648 9.3005
R17928 gnd.n6785 gnd.n6784 9.3005
R17929 gnd.n6786 gnd.n647 9.3005
R17930 gnd.n6788 gnd.n6787 9.3005
R17931 gnd.n643 gnd.n642 9.3005
R17932 gnd.n6795 gnd.n6794 9.3005
R17933 gnd.n6796 gnd.n641 9.3005
R17934 gnd.n6798 gnd.n6797 9.3005
R17935 gnd.n637 gnd.n636 9.3005
R17936 gnd.n6805 gnd.n6804 9.3005
R17937 gnd.n6806 gnd.n635 9.3005
R17938 gnd.n6808 gnd.n6807 9.3005
R17939 gnd.n631 gnd.n630 9.3005
R17940 gnd.n6815 gnd.n6814 9.3005
R17941 gnd.n6816 gnd.n629 9.3005
R17942 gnd.n6818 gnd.n6817 9.3005
R17943 gnd.n625 gnd.n624 9.3005
R17944 gnd.n6825 gnd.n6824 9.3005
R17945 gnd.n6826 gnd.n623 9.3005
R17946 gnd.n6828 gnd.n6827 9.3005
R17947 gnd.n619 gnd.n618 9.3005
R17948 gnd.n6835 gnd.n6834 9.3005
R17949 gnd.n6836 gnd.n617 9.3005
R17950 gnd.n6838 gnd.n6837 9.3005
R17951 gnd.n613 gnd.n612 9.3005
R17952 gnd.n6845 gnd.n6844 9.3005
R17953 gnd.n6846 gnd.n611 9.3005
R17954 gnd.n6848 gnd.n6847 9.3005
R17955 gnd.n607 gnd.n606 9.3005
R17956 gnd.n6855 gnd.n6854 9.3005
R17957 gnd.n6856 gnd.n605 9.3005
R17958 gnd.n6858 gnd.n6857 9.3005
R17959 gnd.n601 gnd.n600 9.3005
R17960 gnd.n6865 gnd.n6864 9.3005
R17961 gnd.n6866 gnd.n599 9.3005
R17962 gnd.n6868 gnd.n6867 9.3005
R17963 gnd.n595 gnd.n594 9.3005
R17964 gnd.n6875 gnd.n6874 9.3005
R17965 gnd.n6876 gnd.n593 9.3005
R17966 gnd.n6878 gnd.n6877 9.3005
R17967 gnd.n589 gnd.n588 9.3005
R17968 gnd.n6885 gnd.n6884 9.3005
R17969 gnd.n6886 gnd.n587 9.3005
R17970 gnd.n6888 gnd.n6887 9.3005
R17971 gnd.n583 gnd.n582 9.3005
R17972 gnd.n6895 gnd.n6894 9.3005
R17973 gnd.n6896 gnd.n581 9.3005
R17974 gnd.n6898 gnd.n6897 9.3005
R17975 gnd.n577 gnd.n576 9.3005
R17976 gnd.n6905 gnd.n6904 9.3005
R17977 gnd.n6906 gnd.n575 9.3005
R17978 gnd.n6908 gnd.n6907 9.3005
R17979 gnd.n571 gnd.n570 9.3005
R17980 gnd.n6915 gnd.n6914 9.3005
R17981 gnd.n6916 gnd.n569 9.3005
R17982 gnd.n6918 gnd.n6917 9.3005
R17983 gnd.n565 gnd.n564 9.3005
R17984 gnd.n6925 gnd.n6924 9.3005
R17985 gnd.n6926 gnd.n563 9.3005
R17986 gnd.n6928 gnd.n6927 9.3005
R17987 gnd.n559 gnd.n558 9.3005
R17988 gnd.n6935 gnd.n6934 9.3005
R17989 gnd.n6936 gnd.n557 9.3005
R17990 gnd.n6938 gnd.n6937 9.3005
R17991 gnd.n553 gnd.n552 9.3005
R17992 gnd.n6945 gnd.n6944 9.3005
R17993 gnd.n6946 gnd.n551 9.3005
R17994 gnd.n6948 gnd.n6947 9.3005
R17995 gnd.n547 gnd.n546 9.3005
R17996 gnd.n6955 gnd.n6954 9.3005
R17997 gnd.n6956 gnd.n545 9.3005
R17998 gnd.n6958 gnd.n6957 9.3005
R17999 gnd.n541 gnd.n540 9.3005
R18000 gnd.n6965 gnd.n6964 9.3005
R18001 gnd.n6966 gnd.n539 9.3005
R18002 gnd.n6968 gnd.n6967 9.3005
R18003 gnd.n535 gnd.n534 9.3005
R18004 gnd.n6975 gnd.n6974 9.3005
R18005 gnd.n6976 gnd.n533 9.3005
R18006 gnd.n6978 gnd.n6977 9.3005
R18007 gnd.n529 gnd.n528 9.3005
R18008 gnd.n6985 gnd.n6984 9.3005
R18009 gnd.n6986 gnd.n527 9.3005
R18010 gnd.n6988 gnd.n6987 9.3005
R18011 gnd.n523 gnd.n522 9.3005
R18012 gnd.n6995 gnd.n6994 9.3005
R18013 gnd.n6996 gnd.n521 9.3005
R18014 gnd.n6998 gnd.n6997 9.3005
R18015 gnd.n517 gnd.n516 9.3005
R18016 gnd.n7005 gnd.n7004 9.3005
R18017 gnd.n7006 gnd.n515 9.3005
R18018 gnd.n7008 gnd.n7007 9.3005
R18019 gnd.n511 gnd.n510 9.3005
R18020 gnd.n7015 gnd.n7014 9.3005
R18021 gnd.n7016 gnd.n509 9.3005
R18022 gnd.n7018 gnd.n7017 9.3005
R18023 gnd.n505 gnd.n504 9.3005
R18024 gnd.n7025 gnd.n7024 9.3005
R18025 gnd.n7026 gnd.n503 9.3005
R18026 gnd.n7028 gnd.n7027 9.3005
R18027 gnd.n499 gnd.n498 9.3005
R18028 gnd.n7035 gnd.n7034 9.3005
R18029 gnd.n7036 gnd.n497 9.3005
R18030 gnd.n7038 gnd.n7037 9.3005
R18031 gnd.n493 gnd.n492 9.3005
R18032 gnd.n7045 gnd.n7044 9.3005
R18033 gnd.n7046 gnd.n491 9.3005
R18034 gnd.n7048 gnd.n7047 9.3005
R18035 gnd.n487 gnd.n486 9.3005
R18036 gnd.n7055 gnd.n7054 9.3005
R18037 gnd.n7056 gnd.n485 9.3005
R18038 gnd.n7058 gnd.n7057 9.3005
R18039 gnd.n481 gnd.n480 9.3005
R18040 gnd.n7065 gnd.n7064 9.3005
R18041 gnd.n7066 gnd.n479 9.3005
R18042 gnd.n7068 gnd.n7067 9.3005
R18043 gnd.n475 gnd.n474 9.3005
R18044 gnd.n7075 gnd.n7074 9.3005
R18045 gnd.n7076 gnd.n473 9.3005
R18046 gnd.n7078 gnd.n7077 9.3005
R18047 gnd.n469 gnd.n468 9.3005
R18048 gnd.n7085 gnd.n7084 9.3005
R18049 gnd.n7086 gnd.n467 9.3005
R18050 gnd.n7088 gnd.n7087 9.3005
R18051 gnd.n463 gnd.n462 9.3005
R18052 gnd.n7095 gnd.n7094 9.3005
R18053 gnd.n7096 gnd.n461 9.3005
R18054 gnd.n7098 gnd.n7097 9.3005
R18055 gnd.n457 gnd.n456 9.3005
R18056 gnd.n7105 gnd.n7104 9.3005
R18057 gnd.n7106 gnd.n455 9.3005
R18058 gnd.n7108 gnd.n7107 9.3005
R18059 gnd.n451 gnd.n450 9.3005
R18060 gnd.n7115 gnd.n7114 9.3005
R18061 gnd.n7116 gnd.n449 9.3005
R18062 gnd.n7118 gnd.n7117 9.3005
R18063 gnd.n445 gnd.n444 9.3005
R18064 gnd.n7125 gnd.n7124 9.3005
R18065 gnd.n7126 gnd.n443 9.3005
R18066 gnd.n7128 gnd.n7127 9.3005
R18067 gnd.n439 gnd.n438 9.3005
R18068 gnd.n7135 gnd.n7134 9.3005
R18069 gnd.n7136 gnd.n437 9.3005
R18070 gnd.n7138 gnd.n7137 9.3005
R18071 gnd.n433 gnd.n432 9.3005
R18072 gnd.n7145 gnd.n7144 9.3005
R18073 gnd.n7146 gnd.n431 9.3005
R18074 gnd.n7148 gnd.n7147 9.3005
R18075 gnd.n427 gnd.n426 9.3005
R18076 gnd.n7155 gnd.n7154 9.3005
R18077 gnd.n7156 gnd.n425 9.3005
R18078 gnd.n7158 gnd.n7157 9.3005
R18079 gnd.n421 gnd.n420 9.3005
R18080 gnd.n7165 gnd.n7164 9.3005
R18081 gnd.n7166 gnd.n419 9.3005
R18082 gnd.n7168 gnd.n7167 9.3005
R18083 gnd.n415 gnd.n414 9.3005
R18084 gnd.n7175 gnd.n7174 9.3005
R18085 gnd.n7176 gnd.n413 9.3005
R18086 gnd.n7178 gnd.n7177 9.3005
R18087 gnd.n409 gnd.n408 9.3005
R18088 gnd.n7185 gnd.n7184 9.3005
R18089 gnd.n7186 gnd.n407 9.3005
R18090 gnd.n7188 gnd.n7187 9.3005
R18091 gnd.n403 gnd.n402 9.3005
R18092 gnd.n7195 gnd.n7194 9.3005
R18093 gnd.n7196 gnd.n401 9.3005
R18094 gnd.n7199 gnd.n7198 9.3005
R18095 gnd.n7197 gnd.n397 9.3005
R18096 gnd.n7205 gnd.n396 9.3005
R18097 gnd.n7207 gnd.n7206 9.3005
R18098 gnd.n392 gnd.n391 9.3005
R18099 gnd.n7216 gnd.n7215 9.3005
R18100 gnd.n7217 gnd.n390 9.3005
R18101 gnd.n7219 gnd.n7218 9.3005
R18102 gnd.n386 gnd.n385 9.3005
R18103 gnd.n7226 gnd.n7225 9.3005
R18104 gnd.n7227 gnd.n384 9.3005
R18105 gnd.n7229 gnd.n7228 9.3005
R18106 gnd.n380 gnd.n379 9.3005
R18107 gnd.n7236 gnd.n7235 9.3005
R18108 gnd.n7237 gnd.n378 9.3005
R18109 gnd.n7239 gnd.n7238 9.3005
R18110 gnd.n374 gnd.n373 9.3005
R18111 gnd.n7246 gnd.n7245 9.3005
R18112 gnd.n7247 gnd.n372 9.3005
R18113 gnd.n7249 gnd.n7248 9.3005
R18114 gnd.n368 gnd.n367 9.3005
R18115 gnd.n7256 gnd.n7255 9.3005
R18116 gnd.n7257 gnd.n366 9.3005
R18117 gnd.n7259 gnd.n7258 9.3005
R18118 gnd.n362 gnd.n361 9.3005
R18119 gnd.n7266 gnd.n7265 9.3005
R18120 gnd.n7267 gnd.n360 9.3005
R18121 gnd.n7269 gnd.n7268 9.3005
R18122 gnd.n356 gnd.n355 9.3005
R18123 gnd.n7276 gnd.n7275 9.3005
R18124 gnd.n7277 gnd.n354 9.3005
R18125 gnd.n7279 gnd.n7278 9.3005
R18126 gnd.n350 gnd.n349 9.3005
R18127 gnd.n7286 gnd.n7285 9.3005
R18128 gnd.n7287 gnd.n348 9.3005
R18129 gnd.n7289 gnd.n7288 9.3005
R18130 gnd.n344 gnd.n343 9.3005
R18131 gnd.n7296 gnd.n7295 9.3005
R18132 gnd.n7297 gnd.n342 9.3005
R18133 gnd.n7299 gnd.n7298 9.3005
R18134 gnd.n338 gnd.n337 9.3005
R18135 gnd.n7306 gnd.n7305 9.3005
R18136 gnd.n7307 gnd.n336 9.3005
R18137 gnd.n7309 gnd.n7308 9.3005
R18138 gnd.n332 gnd.n331 9.3005
R18139 gnd.n7316 gnd.n7315 9.3005
R18140 gnd.n7317 gnd.n330 9.3005
R18141 gnd.n7319 gnd.n7318 9.3005
R18142 gnd.n326 gnd.n325 9.3005
R18143 gnd.n7326 gnd.n7325 9.3005
R18144 gnd.n7327 gnd.n324 9.3005
R18145 gnd.n7329 gnd.n7328 9.3005
R18146 gnd.n320 gnd.n319 9.3005
R18147 gnd.n7336 gnd.n7335 9.3005
R18148 gnd.n7337 gnd.n318 9.3005
R18149 gnd.n7339 gnd.n7338 9.3005
R18150 gnd.n314 gnd.n313 9.3005
R18151 gnd.n7346 gnd.n7345 9.3005
R18152 gnd.n7347 gnd.n312 9.3005
R18153 gnd.n7349 gnd.n7348 9.3005
R18154 gnd.n308 gnd.n307 9.3005
R18155 gnd.n7356 gnd.n7355 9.3005
R18156 gnd.n7357 gnd.n306 9.3005
R18157 gnd.n7359 gnd.n7358 9.3005
R18158 gnd.n302 gnd.n301 9.3005
R18159 gnd.n7366 gnd.n7365 9.3005
R18160 gnd.n7367 gnd.n300 9.3005
R18161 gnd.n7369 gnd.n7368 9.3005
R18162 gnd.n296 gnd.n295 9.3005
R18163 gnd.n7376 gnd.n7375 9.3005
R18164 gnd.n7377 gnd.n294 9.3005
R18165 gnd.n7379 gnd.n7378 9.3005
R18166 gnd.n290 gnd.n289 9.3005
R18167 gnd.n7386 gnd.n7385 9.3005
R18168 gnd.n7387 gnd.n288 9.3005
R18169 gnd.n7389 gnd.n7388 9.3005
R18170 gnd.n284 gnd.n283 9.3005
R18171 gnd.n7396 gnd.n7395 9.3005
R18172 gnd.n7397 gnd.n282 9.3005
R18173 gnd.n7399 gnd.n7398 9.3005
R18174 gnd.n278 gnd.n277 9.3005
R18175 gnd.n7406 gnd.n7405 9.3005
R18176 gnd.n7407 gnd.n276 9.3005
R18177 gnd.n7409 gnd.n7408 9.3005
R18178 gnd.n272 gnd.n271 9.3005
R18179 gnd.n7416 gnd.n7415 9.3005
R18180 gnd.n7417 gnd.n270 9.3005
R18181 gnd.n7420 gnd.n7419 9.3005
R18182 gnd.n7209 gnd.n7208 9.3005
R18183 gnd.n7735 gnd.n7734 9.3005
R18184 gnd.n7733 gnd.n65 9.3005
R18185 gnd.n5851 gnd.n67 9.3005
R18186 gnd.n5853 gnd.n5852 9.3005
R18187 gnd.n3237 gnd.n3236 9.3005
R18188 gnd.n5864 gnd.n5863 9.3005
R18189 gnd.n5865 gnd.n3235 9.3005
R18190 gnd.n5868 gnd.n5867 9.3005
R18191 gnd.n5866 gnd.n3228 9.3005
R18192 gnd.n5911 gnd.n3229 9.3005
R18193 gnd.n5910 gnd.n3230 9.3005
R18194 gnd.n5909 gnd.n3231 9.3005
R18195 gnd.n5878 gnd.n3232 9.3005
R18196 gnd.n5899 gnd.n5879 9.3005
R18197 gnd.n5898 gnd.n5880 9.3005
R18198 gnd.n5897 gnd.n5881 9.3005
R18199 gnd.n5884 gnd.n5882 9.3005
R18200 gnd.n5887 gnd.n5886 9.3005
R18201 gnd.n5885 gnd.n177 9.3005
R18202 gnd.n7666 gnd.n178 9.3005
R18203 gnd.n7665 gnd.n7664 9.3005
R18204 gnd.n204 gnd.n200 9.3005
R18205 gnd.n208 gnd.n207 9.3005
R18206 gnd.n209 gnd.n199 9.3005
R18207 gnd.n211 gnd.n210 9.3005
R18208 gnd.n214 gnd.n198 9.3005
R18209 gnd.n218 gnd.n217 9.3005
R18210 gnd.n219 gnd.n197 9.3005
R18211 gnd.n221 gnd.n220 9.3005
R18212 gnd.n224 gnd.n196 9.3005
R18213 gnd.n228 gnd.n227 9.3005
R18214 gnd.n229 gnd.n195 9.3005
R18215 gnd.n231 gnd.n230 9.3005
R18216 gnd.n234 gnd.n194 9.3005
R18217 gnd.n237 gnd.n236 9.3005
R18218 gnd.n238 gnd.n193 9.3005
R18219 gnd.n240 gnd.n239 9.3005
R18220 gnd.n182 gnd.n179 9.3005
R18221 gnd.n7663 gnd.n7662 9.3005
R18222 gnd.n202 gnd.n201 9.3005
R18223 gnd.n7480 gnd.n7477 9.3005
R18224 gnd.n7656 gnd.n7481 9.3005
R18225 gnd.n7655 gnd.n7482 9.3005
R18226 gnd.n7654 gnd.n7483 9.3005
R18227 gnd.n7651 gnd.n7484 9.3005
R18228 gnd.n7650 gnd.n7485 9.3005
R18229 gnd.n7647 gnd.n7486 9.3005
R18230 gnd.n7646 gnd.n7487 9.3005
R18231 gnd.n7643 gnd.n7488 9.3005
R18232 gnd.n7642 gnd.n7489 9.3005
R18233 gnd.n7639 gnd.n7490 9.3005
R18234 gnd.n7638 gnd.n7491 9.3005
R18235 gnd.n7635 gnd.n7492 9.3005
R18236 gnd.n7634 gnd.n7493 9.3005
R18237 gnd.n7631 gnd.n7494 9.3005
R18238 gnd.n7630 gnd.n7495 9.3005
R18239 gnd.n7627 gnd.n7496 9.3005
R18240 gnd.n7623 gnd.n7497 9.3005
R18241 gnd.n7620 gnd.n7498 9.3005
R18242 gnd.n7619 gnd.n7499 9.3005
R18243 gnd.n7616 gnd.n7500 9.3005
R18244 gnd.n7615 gnd.n7501 9.3005
R18245 gnd.n7612 gnd.n7502 9.3005
R18246 gnd.n7611 gnd.n7503 9.3005
R18247 gnd.n7608 gnd.n7504 9.3005
R18248 gnd.n7607 gnd.n7505 9.3005
R18249 gnd.n7604 gnd.n7506 9.3005
R18250 gnd.n7603 gnd.n7507 9.3005
R18251 gnd.n7600 gnd.n7508 9.3005
R18252 gnd.n7599 gnd.n7509 9.3005
R18253 gnd.n7596 gnd.n7510 9.3005
R18254 gnd.n7595 gnd.n7511 9.3005
R18255 gnd.n7592 gnd.n7512 9.3005
R18256 gnd.n7591 gnd.n7513 9.3005
R18257 gnd.n7588 gnd.n7514 9.3005
R18258 gnd.n7587 gnd.n7515 9.3005
R18259 gnd.n7584 gnd.n7583 9.3005
R18260 gnd.n7582 gnd.n7516 9.3005
R18261 gnd.n7581 gnd.n7580 9.3005
R18262 gnd.n7577 gnd.n7519 9.3005
R18263 gnd.n7574 gnd.n7520 9.3005
R18264 gnd.n7573 gnd.n7521 9.3005
R18265 gnd.n7570 gnd.n7522 9.3005
R18266 gnd.n7569 gnd.n7523 9.3005
R18267 gnd.n7566 gnd.n7524 9.3005
R18268 gnd.n7565 gnd.n7525 9.3005
R18269 gnd.n7562 gnd.n7526 9.3005
R18270 gnd.n7561 gnd.n7527 9.3005
R18271 gnd.n7558 gnd.n7528 9.3005
R18272 gnd.n7557 gnd.n7529 9.3005
R18273 gnd.n7554 gnd.n7530 9.3005
R18274 gnd.n7553 gnd.n7531 9.3005
R18275 gnd.n7550 gnd.n7532 9.3005
R18276 gnd.n7549 gnd.n7533 9.3005
R18277 gnd.n7546 gnd.n7534 9.3005
R18278 gnd.n7545 gnd.n7535 9.3005
R18279 gnd.n7542 gnd.n7541 9.3005
R18280 gnd.n7540 gnd.n7537 9.3005
R18281 gnd.n7479 gnd.n7478 9.3005
R18282 gnd.n5725 gnd.n3074 9.3005
R18283 gnd.n5993 gnd.n3075 9.3005
R18284 gnd.n5992 gnd.n3076 9.3005
R18285 gnd.n5991 gnd.n3077 9.3005
R18286 gnd.n3259 gnd.n3078 9.3005
R18287 gnd.n5981 gnd.n3095 9.3005
R18288 gnd.n5980 gnd.n3096 9.3005
R18289 gnd.n5979 gnd.n3097 9.3005
R18290 gnd.n5744 gnd.n3098 9.3005
R18291 gnd.n5969 gnd.n3116 9.3005
R18292 gnd.n5968 gnd.n3117 9.3005
R18293 gnd.n5967 gnd.n3118 9.3005
R18294 gnd.n5807 gnd.n3119 9.3005
R18295 gnd.n5957 gnd.n3135 9.3005
R18296 gnd.n5956 gnd.n3136 9.3005
R18297 gnd.n5955 gnd.n3137 9.3005
R18298 gnd.n3239 gnd.n3138 9.3005
R18299 gnd.n5837 gnd.n5836 9.3005
R18300 gnd.n5841 gnd.n5840 9.3005
R18301 gnd.n5842 gnd.n3168 9.3005
R18302 gnd.n5933 gnd.n3169 9.3005
R18303 gnd.n5932 gnd.n3170 9.3005
R18304 gnd.n5931 gnd.n3171 9.3005
R18305 gnd.n5930 gnd.n3172 9.3005
R18306 gnd.n5850 gnd.n92 9.3005
R18307 gnd.n7721 gnd.n93 9.3005
R18308 gnd.n7720 gnd.n94 9.3005
R18309 gnd.n7719 gnd.n95 9.3005
R18310 gnd.n3234 gnd.n96 9.3005
R18311 gnd.n7709 gnd.n112 9.3005
R18312 gnd.n7708 gnd.n113 9.3005
R18313 gnd.n7707 gnd.n114 9.3005
R18314 gnd.n5876 gnd.n115 9.3005
R18315 gnd.n7697 gnd.n133 9.3005
R18316 gnd.n7696 gnd.n134 9.3005
R18317 gnd.n7695 gnd.n135 9.3005
R18318 gnd.n5883 gnd.n136 9.3005
R18319 gnd.n7685 gnd.n154 9.3005
R18320 gnd.n7684 gnd.n155 9.3005
R18321 gnd.n7683 gnd.n156 9.3005
R18322 gnd.n173 gnd.n157 9.3005
R18323 gnd.n7673 gnd.n7672 9.3005
R18324 gnd.n5724 gnd.n5723 9.3005
R18325 gnd.n5726 gnd.n5725 9.3005
R18326 gnd.n5727 gnd.n3075 9.3005
R18327 gnd.n5728 gnd.n3076 9.3005
R18328 gnd.n3258 gnd.n3077 9.3005
R18329 gnd.n5740 gnd.n3259 9.3005
R18330 gnd.n5741 gnd.n3095 9.3005
R18331 gnd.n5742 gnd.n3096 9.3005
R18332 gnd.n5743 gnd.n3097 9.3005
R18333 gnd.n5745 gnd.n5744 9.3005
R18334 gnd.n3246 gnd.n3116 9.3005
R18335 gnd.n5805 gnd.n3117 9.3005
R18336 gnd.n5806 gnd.n3118 9.3005
R18337 gnd.n5808 gnd.n5807 9.3005
R18338 gnd.n3240 gnd.n3135 9.3005
R18339 gnd.n5830 gnd.n3136 9.3005
R18340 gnd.n5831 gnd.n3137 9.3005
R18341 gnd.n5832 gnd.n3239 9.3005
R18342 gnd.n5836 gnd.n5835 9.3005
R18343 gnd.n5841 gnd.n3238 9.3005
R18344 gnd.n5843 gnd.n5842 9.3005
R18345 gnd.n5844 gnd.n3169 9.3005
R18346 gnd.n5847 gnd.n3170 9.3005
R18347 gnd.n5848 gnd.n3171 9.3005
R18348 gnd.n5849 gnd.n3172 9.3005
R18349 gnd.n5857 gnd.n5850 9.3005
R18350 gnd.n5858 gnd.n93 9.3005
R18351 gnd.n5859 gnd.n94 9.3005
R18352 gnd.n3233 gnd.n95 9.3005
R18353 gnd.n5872 gnd.n3234 9.3005
R18354 gnd.n5873 gnd.n112 9.3005
R18355 gnd.n5874 gnd.n113 9.3005
R18356 gnd.n5875 gnd.n114 9.3005
R18357 gnd.n5905 gnd.n5876 9.3005
R18358 gnd.n5904 gnd.n133 9.3005
R18359 gnd.n5903 gnd.n134 9.3005
R18360 gnd.n5877 gnd.n135 9.3005
R18361 gnd.n5893 gnd.n5883 9.3005
R18362 gnd.n5892 gnd.n154 9.3005
R18363 gnd.n5891 gnd.n155 9.3005
R18364 gnd.n175 gnd.n156 9.3005
R18365 gnd.n7670 gnd.n173 9.3005
R18366 gnd.n7672 gnd.n7671 9.3005
R18367 gnd.n5724 gnd.n3263 9.3005
R18368 gnd.n3269 gnd.n3266 9.3005
R18369 gnd.n5711 gnd.n3270 9.3005
R18370 gnd.n5713 gnd.n5712 9.3005
R18371 gnd.n5710 gnd.n3272 9.3005
R18372 gnd.n5709 gnd.n5708 9.3005
R18373 gnd.n3274 gnd.n3273 9.3005
R18374 gnd.n5702 gnd.n5701 9.3005
R18375 gnd.n5700 gnd.n3276 9.3005
R18376 gnd.n5699 gnd.n5698 9.3005
R18377 gnd.n3278 gnd.n3277 9.3005
R18378 gnd.n5692 gnd.n5691 9.3005
R18379 gnd.n5690 gnd.n3280 9.3005
R18380 gnd.n5689 gnd.n5688 9.3005
R18381 gnd.n3282 gnd.n3281 9.3005
R18382 gnd.n5682 gnd.n5681 9.3005
R18383 gnd.n5680 gnd.n3284 9.3005
R18384 gnd.n5679 gnd.n5678 9.3005
R18385 gnd.n3286 gnd.n3285 9.3005
R18386 gnd.n5672 gnd.n5671 9.3005
R18387 gnd.n5670 gnd.n3288 9.3005
R18388 gnd.n3290 gnd.n3289 9.3005
R18389 gnd.n5660 gnd.n5659 9.3005
R18390 gnd.n5658 gnd.n3292 9.3005
R18391 gnd.n5657 gnd.n5656 9.3005
R18392 gnd.n3294 gnd.n3293 9.3005
R18393 gnd.n5650 gnd.n5649 9.3005
R18394 gnd.n5648 gnd.n3296 9.3005
R18395 gnd.n5647 gnd.n5646 9.3005
R18396 gnd.n3298 gnd.n3297 9.3005
R18397 gnd.n5638 gnd.n5637 9.3005
R18398 gnd.n5635 gnd.n5548 9.3005
R18399 gnd.n5634 gnd.n5633 9.3005
R18400 gnd.n5550 gnd.n5549 9.3005
R18401 gnd.n5627 gnd.n5626 9.3005
R18402 gnd.n5625 gnd.n5552 9.3005
R18403 gnd.n5624 gnd.n5623 9.3005
R18404 gnd.n5554 gnd.n5553 9.3005
R18405 gnd.n5617 gnd.n5613 9.3005
R18406 gnd.n5612 gnd.n5556 9.3005
R18407 gnd.n5611 gnd.n5610 9.3005
R18408 gnd.n5558 gnd.n5557 9.3005
R18409 gnd.n5604 gnd.n5603 9.3005
R18410 gnd.n5602 gnd.n5560 9.3005
R18411 gnd.n5601 gnd.n5600 9.3005
R18412 gnd.n5562 gnd.n5561 9.3005
R18413 gnd.n5594 gnd.n5593 9.3005
R18414 gnd.n5592 gnd.n5564 9.3005
R18415 gnd.n5591 gnd.n5590 9.3005
R18416 gnd.n5566 gnd.n5565 9.3005
R18417 gnd.n5584 gnd.n5583 9.3005
R18418 gnd.n5582 gnd.n5568 9.3005
R18419 gnd.n5581 gnd.n5580 9.3005
R18420 gnd.n5570 gnd.n5569 9.3005
R18421 gnd.n5574 gnd.n5573 9.3005
R18422 gnd.n5572 gnd.n5571 9.3005
R18423 gnd.n5669 gnd.n5668 9.3005
R18424 gnd.n5721 gnd.n5720 9.3005
R18425 gnd.n5998 gnd.n3064 9.3005
R18426 gnd.n5997 gnd.n3065 9.3005
R18427 gnd.n3085 gnd.n3066 9.3005
R18428 gnd.n5987 gnd.n3086 9.3005
R18429 gnd.n5986 gnd.n3087 9.3005
R18430 gnd.n5985 gnd.n3088 9.3005
R18431 gnd.n3105 gnd.n3089 9.3005
R18432 gnd.n5975 gnd.n3106 9.3005
R18433 gnd.n5974 gnd.n3107 9.3005
R18434 gnd.n5973 gnd.n3108 9.3005
R18435 gnd.n3125 gnd.n3109 9.3005
R18436 gnd.n5963 gnd.n3126 9.3005
R18437 gnd.n5962 gnd.n3127 9.3005
R18438 gnd.n5961 gnd.n3128 9.3005
R18439 gnd.n3129 gnd.n78 9.3005
R18440 gnd.n83 gnd.n77 9.3005
R18441 gnd.n7715 gnd.n103 9.3005
R18442 gnd.n7714 gnd.n104 9.3005
R18443 gnd.n7713 gnd.n105 9.3005
R18444 gnd.n122 gnd.n106 9.3005
R18445 gnd.n7703 gnd.n123 9.3005
R18446 gnd.n7702 gnd.n124 9.3005
R18447 gnd.n7701 gnd.n125 9.3005
R18448 gnd.n143 gnd.n126 9.3005
R18449 gnd.n7691 gnd.n144 9.3005
R18450 gnd.n7690 gnd.n145 9.3005
R18451 gnd.n7689 gnd.n146 9.3005
R18452 gnd.n163 gnd.n147 9.3005
R18453 gnd.n7679 gnd.n164 9.3005
R18454 gnd.n7678 gnd.n165 9.3005
R18455 gnd.n7677 gnd.n166 9.3005
R18456 gnd.n5999 gnd.n3063 9.3005
R18457 gnd.n7726 gnd.n7725 9.3005
R18458 gnd.n4366 gnd.n3877 9.3005
R18459 gnd.n4387 gnd.n4367 9.3005
R18460 gnd.n4386 gnd.n4368 9.3005
R18461 gnd.n4385 gnd.n4369 9.3005
R18462 gnd.n4372 gnd.n4370 9.3005
R18463 gnd.n4381 gnd.n4373 9.3005
R18464 gnd.n4380 gnd.n4374 9.3005
R18465 gnd.n4379 gnd.n4375 9.3005
R18466 gnd.n4377 gnd.n4376 9.3005
R18467 gnd.n3855 gnd.n3854 9.3005
R18468 gnd.n4441 gnd.n4440 9.3005
R18469 gnd.n4442 gnd.n3853 9.3005
R18470 gnd.n4444 gnd.n4443 9.3005
R18471 gnd.n3851 gnd.n3850 9.3005
R18472 gnd.n4449 gnd.n4448 9.3005
R18473 gnd.n4450 gnd.n3849 9.3005
R18474 gnd.n4452 gnd.n4451 9.3005
R18475 gnd.n3847 gnd.n3846 9.3005
R18476 gnd.n4457 gnd.n4456 9.3005
R18477 gnd.n4458 gnd.n3845 9.3005
R18478 gnd.n4460 gnd.n4459 9.3005
R18479 gnd.n3842 gnd.n3841 9.3005
R18480 gnd.n4467 gnd.n4466 9.3005
R18481 gnd.n4468 gnd.n3840 9.3005
R18482 gnd.n4473 gnd.n4469 9.3005
R18483 gnd.n4472 gnd.n4471 9.3005
R18484 gnd.n4470 gnd.n2916 9.3005
R18485 gnd.n6147 gnd.n2917 9.3005
R18486 gnd.n6146 gnd.n2918 9.3005
R18487 gnd.n6145 gnd.n2919 9.3005
R18488 gnd.n2934 gnd.n2920 9.3005
R18489 gnd.n6133 gnd.n2935 9.3005
R18490 gnd.n6132 gnd.n2936 9.3005
R18491 gnd.n6131 gnd.n2937 9.3005
R18492 gnd.n4556 gnd.n2938 9.3005
R18493 gnd.n4558 gnd.n4557 9.3005
R18494 gnd.n3711 gnd.n3710 9.3005
R18495 gnd.n4591 gnd.n4590 9.3005
R18496 gnd.n4592 gnd.n3709 9.3005
R18497 gnd.n4594 gnd.n4593 9.3005
R18498 gnd.n3686 gnd.n3685 9.3005
R18499 gnd.n4634 gnd.n4633 9.3005
R18500 gnd.n4635 gnd.n3684 9.3005
R18501 gnd.n4637 gnd.n4636 9.3005
R18502 gnd.n3671 gnd.n3670 9.3005
R18503 gnd.n4679 gnd.n4678 9.3005
R18504 gnd.n4680 gnd.n3669 9.3005
R18505 gnd.n4684 gnd.n4681 9.3005
R18506 gnd.n4683 gnd.n4682 9.3005
R18507 gnd.n3643 gnd.n3642 9.3005
R18508 gnd.n4752 gnd.n4751 9.3005
R18509 gnd.n4753 gnd.n3641 9.3005
R18510 gnd.n4755 gnd.n4754 9.3005
R18511 gnd.n3623 gnd.n3622 9.3005
R18512 gnd.n4780 gnd.n4779 9.3005
R18513 gnd.n4781 gnd.n3621 9.3005
R18514 gnd.n4783 gnd.n4782 9.3005
R18515 gnd.n3602 gnd.n3601 9.3005
R18516 gnd.n4813 gnd.n4812 9.3005
R18517 gnd.n4814 gnd.n3600 9.3005
R18518 gnd.n4816 gnd.n4815 9.3005
R18519 gnd.n3585 gnd.n3584 9.3005
R18520 gnd.n4857 gnd.n4856 9.3005
R18521 gnd.n4858 gnd.n3583 9.3005
R18522 gnd.n4862 gnd.n4859 9.3005
R18523 gnd.n4861 gnd.n4860 9.3005
R18524 gnd.n3556 gnd.n3555 9.3005
R18525 gnd.n4907 gnd.n4906 9.3005
R18526 gnd.n4908 gnd.n3554 9.3005
R18527 gnd.n4910 gnd.n4909 9.3005
R18528 gnd.n3537 gnd.n3536 9.3005
R18529 gnd.n4935 gnd.n4934 9.3005
R18530 gnd.n4936 gnd.n3535 9.3005
R18531 gnd.n4947 gnd.n4937 9.3005
R18532 gnd.n4946 gnd.n4938 9.3005
R18533 gnd.n4945 gnd.n4939 9.3005
R18534 gnd.n3506 gnd.n3505 9.3005
R18535 gnd.n5010 gnd.n5009 9.3005
R18536 gnd.n5011 gnd.n3504 9.3005
R18537 gnd.n5015 gnd.n5012 9.3005
R18538 gnd.n5014 gnd.n5013 9.3005
R18539 gnd.n3478 gnd.n3477 9.3005
R18540 gnd.n5062 gnd.n5061 9.3005
R18541 gnd.n5063 gnd.n3476 9.3005
R18542 gnd.n5067 gnd.n5064 9.3005
R18543 gnd.n5066 gnd.n5065 9.3005
R18544 gnd.n3461 gnd.n3460 9.3005
R18545 gnd.n5090 gnd.n5089 9.3005
R18546 gnd.n5091 gnd.n3459 9.3005
R18547 gnd.n5093 gnd.n5092 9.3005
R18548 gnd.n3403 gnd.n3402 9.3005
R18549 gnd.n5133 gnd.n5132 9.3005
R18550 gnd.n5134 gnd.n3401 9.3005
R18551 gnd.n5136 gnd.n5135 9.3005
R18552 gnd.n3381 gnd.n3380 9.3005
R18553 gnd.n5161 gnd.n5160 9.3005
R18554 gnd.n5162 gnd.n3379 9.3005
R18555 gnd.n5167 gnd.n5163 9.3005
R18556 gnd.n5166 gnd.n5165 9.3005
R18557 gnd.n5164 gnd.n3350 9.3005
R18558 gnd.n5382 gnd.n3351 9.3005
R18559 gnd.n5381 gnd.n3352 9.3005
R18560 gnd.n5380 gnd.n3353 9.3005
R18561 gnd.n3356 gnd.n3355 9.3005
R18562 gnd.n3354 gnd.n3041 9.3005
R18563 gnd.n6014 gnd.n3042 9.3005
R18564 gnd.n6013 gnd.n3043 9.3005
R18565 gnd.n6012 gnd.n3044 9.3005
R18566 gnd.n3050 gnd.n3045 9.3005
R18567 gnd.n6006 gnd.n3051 9.3005
R18568 gnd.n6005 gnd.n3052 9.3005
R18569 gnd.n6004 gnd.n3053 9.3005
R18570 gnd.n5766 gnd.n3054 9.3005
R18571 gnd.n5769 gnd.n5768 9.3005
R18572 gnd.n5770 gnd.n5765 9.3005
R18573 gnd.n5772 gnd.n5771 9.3005
R18574 gnd.n5763 gnd.n5762 9.3005
R18575 gnd.n5777 gnd.n5776 9.3005
R18576 gnd.n5778 gnd.n5761 9.3005
R18577 gnd.n5780 gnd.n5779 9.3005
R18578 gnd.n3252 gnd.n3251 9.3005
R18579 gnd.n5785 gnd.n5784 9.3005
R18580 gnd.n5786 gnd.n3250 9.3005
R18581 gnd.n5800 gnd.n5787 9.3005
R18582 gnd.n5799 gnd.n5788 9.3005
R18583 gnd.n5798 gnd.n5789 9.3005
R18584 gnd.n5791 gnd.n5790 9.3005
R18585 gnd.n5794 gnd.n5792 9.3005
R18586 gnd.n5922 gnd.n3183 9.3005
R18587 gnd.n3186 gnd.n3184 9.3005
R18588 gnd.n5918 gnd.n3187 9.3005
R18589 gnd.n5917 gnd.n3188 9.3005
R18590 gnd.n5916 gnd.n3189 9.3005
R18591 gnd.n3192 gnd.n3190 9.3005
R18592 gnd.n3224 gnd.n3193 9.3005
R18593 gnd.n3223 gnd.n3194 9.3005
R18594 gnd.n3222 gnd.n3195 9.3005
R18595 gnd.n3198 gnd.n3196 9.3005
R18596 gnd.n3218 gnd.n3199 9.3005
R18597 gnd.n3217 gnd.n3200 9.3005
R18598 gnd.n3216 gnd.n3201 9.3005
R18599 gnd.n3204 gnd.n3202 9.3005
R18600 gnd.n3212 gnd.n3205 9.3005
R18601 gnd.n3211 gnd.n3206 9.3005
R18602 gnd.n3210 gnd.n3208 9.3005
R18603 gnd.n3207 gnd.n246 9.3005
R18604 gnd.n7444 gnd.n247 9.3005
R18605 gnd.n7443 gnd.n248 9.3005
R18606 gnd.n7442 gnd.n249 9.3005
R18607 gnd.n254 gnd.n250 9.3005
R18608 gnd.n7436 gnd.n255 9.3005
R18609 gnd.n7435 gnd.n256 9.3005
R18610 gnd.n7434 gnd.n257 9.3005
R18611 gnd.n262 gnd.n258 9.3005
R18612 gnd.n7428 gnd.n263 9.3005
R18613 gnd.n7427 gnd.n264 9.3005
R18614 gnd.n7426 gnd.n265 9.3005
R18615 gnd.n7418 gnd.n266 9.3005
R18616 gnd.n4350 gnd.n4349 9.3005
R18617 gnd.n4254 gnd.n3926 9.3005
R18618 gnd.n4253 gnd.n3927 9.3005
R18619 gnd.n4252 gnd.n3928 9.3005
R18620 gnd.n4220 gnd.n3929 9.3005
R18621 gnd.n4242 gnd.n4221 9.3005
R18622 gnd.n4241 gnd.n4222 9.3005
R18623 gnd.n4240 gnd.n4223 9.3005
R18624 gnd.n4228 gnd.n4224 9.3005
R18625 gnd.n4230 gnd.n4229 9.3005
R18626 gnd.n3907 gnd.n3906 9.3005
R18627 gnd.n4290 gnd.n4289 9.3005
R18628 gnd.n4291 gnd.n3905 9.3005
R18629 gnd.n4293 gnd.n4292 9.3005
R18630 gnd.n3902 gnd.n3901 9.3005
R18631 gnd.n4304 gnd.n4303 9.3005
R18632 gnd.n4305 gnd.n3900 9.3005
R18633 gnd.n4308 gnd.n4307 9.3005
R18634 gnd.n4306 gnd.n3891 9.3005
R18635 gnd.n4352 gnd.n3892 9.3005
R18636 gnd.n4351 gnd.n3893 9.3005
R18637 gnd.n3958 gnd.n3925 9.3005
R18638 gnd.n3957 gnd.n3954 9.3005
R18639 gnd.n3969 gnd.n3953 9.3005
R18640 gnd.n3970 gnd.n3952 9.3005
R18641 gnd.n3971 gnd.n3951 9.3005
R18642 gnd.n3950 gnd.n3948 9.3005
R18643 gnd.n3977 gnd.n3947 9.3005
R18644 gnd.n3978 gnd.n3946 9.3005
R18645 gnd.n3979 gnd.n3945 9.3005
R18646 gnd.n3944 gnd.n3942 9.3005
R18647 gnd.n3985 gnd.n3941 9.3005
R18648 gnd.n3986 gnd.n3940 9.3005
R18649 gnd.n3987 gnd.n3939 9.3005
R18650 gnd.n3938 gnd.n3936 9.3005
R18651 gnd.n3992 gnd.n3935 9.3005
R18652 gnd.n3993 gnd.n3934 9.3005
R18653 gnd.n3932 gnd.n3931 9.3005
R18654 gnd.n3999 gnd.n3998 9.3005
R18655 gnd.n3963 gnd.n3960 9.3005
R18656 gnd.n3959 gnd.n3956 9.3005
R18657 gnd.n6225 gnd.n2750 9.3005
R18658 gnd.n6228 gnd.n2749 9.3005
R18659 gnd.n6229 gnd.n2748 9.3005
R18660 gnd.n6232 gnd.n2747 9.3005
R18661 gnd.n6233 gnd.n2746 9.3005
R18662 gnd.n6236 gnd.n2745 9.3005
R18663 gnd.n6237 gnd.n2744 9.3005
R18664 gnd.n6240 gnd.n2743 9.3005
R18665 gnd.n6242 gnd.n2740 9.3005
R18666 gnd.n6245 gnd.n2739 9.3005
R18667 gnd.n6246 gnd.n2738 9.3005
R18668 gnd.n6249 gnd.n2737 9.3005
R18669 gnd.n6250 gnd.n2736 9.3005
R18670 gnd.n6253 gnd.n2735 9.3005
R18671 gnd.n6254 gnd.n2734 9.3005
R18672 gnd.n6257 gnd.n2733 9.3005
R18673 gnd.n6258 gnd.n2732 9.3005
R18674 gnd.n6261 gnd.n2731 9.3005
R18675 gnd.n6262 gnd.n2730 9.3005
R18676 gnd.n6265 gnd.n2729 9.3005
R18677 gnd.n6266 gnd.n2728 9.3005
R18678 gnd.n6269 gnd.n2727 9.3005
R18679 gnd.n6270 gnd.n2726 9.3005
R18680 gnd.n6271 gnd.n2725 9.3005
R18681 gnd.n2724 gnd.n2721 9.3005
R18682 gnd.n2723 gnd.n2722 9.3005
R18683 gnd.n2847 gnd.n2846 9.3005
R18684 gnd.n2843 gnd.n2753 9.3005
R18685 gnd.n2840 gnd.n2754 9.3005
R18686 gnd.n2839 gnd.n2755 9.3005
R18687 gnd.n2836 gnd.n2756 9.3005
R18688 gnd.n2835 gnd.n2757 9.3005
R18689 gnd.n2832 gnd.n2758 9.3005
R18690 gnd.n2831 gnd.n2759 9.3005
R18691 gnd.n2828 gnd.n2827 9.3005
R18692 gnd.n2826 gnd.n2760 9.3005
R18693 gnd.n2825 gnd.n2824 9.3005
R18694 gnd.n2821 gnd.n2763 9.3005
R18695 gnd.n2818 gnd.n2764 9.3005
R18696 gnd.n2817 gnd.n2765 9.3005
R18697 gnd.n2814 gnd.n2766 9.3005
R18698 gnd.n2813 gnd.n2767 9.3005
R18699 gnd.n2810 gnd.n2768 9.3005
R18700 gnd.n2809 gnd.n2769 9.3005
R18701 gnd.n2806 gnd.n2770 9.3005
R18702 gnd.n2805 gnd.n2771 9.3005
R18703 gnd.n2802 gnd.n2772 9.3005
R18704 gnd.n2801 gnd.n2773 9.3005
R18705 gnd.n2798 gnd.n2774 9.3005
R18706 gnd.n2797 gnd.n2775 9.3005
R18707 gnd.n2794 gnd.n2776 9.3005
R18708 gnd.n2793 gnd.n2777 9.3005
R18709 gnd.n2790 gnd.n2778 9.3005
R18710 gnd.n2789 gnd.n2779 9.3005
R18711 gnd.n2786 gnd.n2785 9.3005
R18712 gnd.n2784 gnd.n2781 9.3005
R18713 gnd.n2848 gnd.n2751 9.3005
R18714 gnd.n4215 gnd.n2380 9.3005
R18715 gnd.n6478 gnd.n2381 9.3005
R18716 gnd.n6477 gnd.n2382 9.3005
R18717 gnd.n6476 gnd.n2383 9.3005
R18718 gnd.n4218 gnd.n2384 9.3005
R18719 gnd.n6466 gnd.n2402 9.3005
R18720 gnd.n6465 gnd.n2403 9.3005
R18721 gnd.n6464 gnd.n2404 9.3005
R18722 gnd.n4225 gnd.n2405 9.3005
R18723 gnd.n6454 gnd.n2423 9.3005
R18724 gnd.n6453 gnd.n2424 9.3005
R18725 gnd.n6452 gnd.n2425 9.3005
R18726 gnd.n3904 gnd.n2426 9.3005
R18727 gnd.n6442 gnd.n2443 9.3005
R18728 gnd.n6441 gnd.n2444 9.3005
R18729 gnd.n6440 gnd.n2445 9.3005
R18730 gnd.n3899 gnd.n2446 9.3005
R18731 gnd.n6429 gnd.n2462 9.3005
R18732 gnd.n6428 gnd.n2463 9.3005
R18733 gnd.n6427 gnd.n2464 9.3005
R18734 gnd.n4316 gnd.n2465 9.3005
R18735 gnd.n6416 gnd.n2478 9.3005
R18736 gnd.n6415 gnd.n2479 9.3005
R18737 gnd.n6414 gnd.n2480 9.3005
R18738 gnd.n4336 gnd.n2481 9.3005
R18739 gnd.n6403 gnd.n2496 9.3005
R18740 gnd.n6402 gnd.n2497 9.3005
R18741 gnd.n6401 gnd.n2498 9.3005
R18742 gnd.n3870 gnd.n2499 9.3005
R18743 gnd.n6391 gnd.n2515 9.3005
R18744 gnd.n6390 gnd.n2516 9.3005
R18745 gnd.n6389 gnd.n2517 9.3005
R18746 gnd.n3864 gnd.n2518 9.3005
R18747 gnd.n6379 gnd.n2536 9.3005
R18748 gnd.n6378 gnd.n2537 9.3005
R18749 gnd.n6377 gnd.n2538 9.3005
R18750 gnd.n4418 gnd.n2539 9.3005
R18751 gnd.n6367 gnd.n2556 9.3005
R18752 gnd.n6366 gnd.n2557 9.3005
R18753 gnd.n6365 gnd.n2558 9.3005
R18754 gnd.n2576 gnd.n2559 9.3005
R18755 gnd.n6355 gnd.n6354 9.3005
R18756 gnd.n4214 gnd.n4213 9.3005
R18757 gnd.n4216 gnd.n4215 9.3005
R18758 gnd.n4217 gnd.n2381 9.3005
R18759 gnd.n4248 gnd.n2382 9.3005
R18760 gnd.n4247 gnd.n2383 9.3005
R18761 gnd.n4246 gnd.n4218 9.3005
R18762 gnd.n4219 gnd.n2402 9.3005
R18763 gnd.n4236 gnd.n2403 9.3005
R18764 gnd.n4235 gnd.n2404 9.3005
R18765 gnd.n4234 gnd.n4225 9.3005
R18766 gnd.n4227 gnd.n2423 9.3005
R18767 gnd.n4226 gnd.n2424 9.3005
R18768 gnd.n3903 gnd.n2425 9.3005
R18769 gnd.n4297 gnd.n3904 9.3005
R18770 gnd.n4298 gnd.n2443 9.3005
R18771 gnd.n4299 gnd.n2444 9.3005
R18772 gnd.n3898 gnd.n2445 9.3005
R18773 gnd.n4312 gnd.n3899 9.3005
R18774 gnd.n4313 gnd.n2462 9.3005
R18775 gnd.n4314 gnd.n2463 9.3005
R18776 gnd.n4315 gnd.n2464 9.3005
R18777 gnd.n4319 gnd.n4316 9.3005
R18778 gnd.n4320 gnd.n2478 9.3005
R18779 gnd.n4334 gnd.n2479 9.3005
R18780 gnd.n4335 gnd.n2480 9.3005
R18781 gnd.n4339 gnd.n4336 9.3005
R18782 gnd.n4338 gnd.n2496 9.3005
R18783 gnd.n4337 gnd.n2497 9.3005
R18784 gnd.n3869 gnd.n2498 9.3005
R18785 gnd.n4400 gnd.n3870 9.3005
R18786 gnd.n4401 gnd.n2515 9.3005
R18787 gnd.n4402 gnd.n2516 9.3005
R18788 gnd.n3863 gnd.n2517 9.3005
R18789 gnd.n4414 gnd.n3864 9.3005
R18790 gnd.n4415 gnd.n2536 9.3005
R18791 gnd.n4416 gnd.n2537 9.3005
R18792 gnd.n4417 gnd.n2538 9.3005
R18793 gnd.n4421 gnd.n4418 9.3005
R18794 gnd.n4422 gnd.n2556 9.3005
R18795 gnd.n4423 gnd.n2557 9.3005
R18796 gnd.n2578 gnd.n2558 9.3005
R18797 gnd.n6352 gnd.n2576 9.3005
R18798 gnd.n6354 gnd.n6353 9.3005
R18799 gnd.n4214 gnd.n3930 9.3005
R18800 gnd.n4003 gnd.n4000 9.3005
R18801 gnd.n4201 gnd.n4004 9.3005
R18802 gnd.n4203 gnd.n4202 9.3005
R18803 gnd.n4200 gnd.n4006 9.3005
R18804 gnd.n4199 gnd.n4198 9.3005
R18805 gnd.n4008 gnd.n4007 9.3005
R18806 gnd.n4192 gnd.n4191 9.3005
R18807 gnd.n4190 gnd.n4010 9.3005
R18808 gnd.n4189 gnd.n4188 9.3005
R18809 gnd.n4012 gnd.n4011 9.3005
R18810 gnd.n4182 gnd.n4181 9.3005
R18811 gnd.n4180 gnd.n4014 9.3005
R18812 gnd.n4179 gnd.n4178 9.3005
R18813 gnd.n4016 gnd.n4015 9.3005
R18814 gnd.n4172 gnd.n4171 9.3005
R18815 gnd.n4170 gnd.n4018 9.3005
R18816 gnd.n4169 gnd.n4168 9.3005
R18817 gnd.n4020 gnd.n4019 9.3005
R18818 gnd.n4162 gnd.n4161 9.3005
R18819 gnd.n4160 gnd.n4022 9.3005
R18820 gnd.n4024 gnd.n4023 9.3005
R18821 gnd.n4150 gnd.n4149 9.3005
R18822 gnd.n4148 gnd.n4026 9.3005
R18823 gnd.n4147 gnd.n4146 9.3005
R18824 gnd.n4028 gnd.n4027 9.3005
R18825 gnd.n4140 gnd.n4139 9.3005
R18826 gnd.n4138 gnd.n4030 9.3005
R18827 gnd.n4137 gnd.n4136 9.3005
R18828 gnd.n4032 gnd.n4031 9.3005
R18829 gnd.n4130 gnd.n4129 9.3005
R18830 gnd.n4128 gnd.n4034 9.3005
R18831 gnd.n4127 gnd.n4126 9.3005
R18832 gnd.n4036 gnd.n4035 9.3005
R18833 gnd.n4120 gnd.n4119 9.3005
R18834 gnd.n4118 gnd.n4038 9.3005
R18835 gnd.n4117 gnd.n4116 9.3005
R18836 gnd.n4040 gnd.n4039 9.3005
R18837 gnd.n4110 gnd.n4109 9.3005
R18838 gnd.n4108 gnd.n4042 9.3005
R18839 gnd.n4107 gnd.n4106 9.3005
R18840 gnd.n4044 gnd.n4043 9.3005
R18841 gnd.n4100 gnd.n4099 9.3005
R18842 gnd.n4098 gnd.n4049 9.3005
R18843 gnd.n4097 gnd.n4096 9.3005
R18844 gnd.n4051 gnd.n4050 9.3005
R18845 gnd.n4090 gnd.n4089 9.3005
R18846 gnd.n4088 gnd.n4053 9.3005
R18847 gnd.n4087 gnd.n4086 9.3005
R18848 gnd.n4055 gnd.n4054 9.3005
R18849 gnd.n4080 gnd.n4079 9.3005
R18850 gnd.n4078 gnd.n4057 9.3005
R18851 gnd.n4077 gnd.n4076 9.3005
R18852 gnd.n4059 gnd.n4058 9.3005
R18853 gnd.n4070 gnd.n4069 9.3005
R18854 gnd.n4068 gnd.n4061 9.3005
R18855 gnd.n4067 gnd.n4066 9.3005
R18856 gnd.n4063 gnd.n4062 9.3005
R18857 gnd.n4159 gnd.n4158 9.3005
R18858 gnd.n4211 gnd.n4210 9.3005
R18859 gnd.n6483 gnd.n2371 9.3005
R18860 gnd.n6482 gnd.n2372 9.3005
R18861 gnd.n2391 gnd.n2373 9.3005
R18862 gnd.n6472 gnd.n2392 9.3005
R18863 gnd.n6471 gnd.n2393 9.3005
R18864 gnd.n6470 gnd.n2394 9.3005
R18865 gnd.n2412 gnd.n2395 9.3005
R18866 gnd.n6460 gnd.n2413 9.3005
R18867 gnd.n6459 gnd.n2414 9.3005
R18868 gnd.n6458 gnd.n2415 9.3005
R18869 gnd.n2432 gnd.n2416 9.3005
R18870 gnd.n6448 gnd.n2433 9.3005
R18871 gnd.n6447 gnd.n2434 9.3005
R18872 gnd.n6446 gnd.n2435 9.3005
R18873 gnd.n2453 gnd.n2436 9.3005
R18874 gnd.n2505 gnd.n2489 9.3005
R18875 gnd.n6397 gnd.n2506 9.3005
R18876 gnd.n6396 gnd.n2507 9.3005
R18877 gnd.n6395 gnd.n2508 9.3005
R18878 gnd.n2525 gnd.n2509 9.3005
R18879 gnd.n6385 gnd.n2526 9.3005
R18880 gnd.n6384 gnd.n2527 9.3005
R18881 gnd.n6383 gnd.n2528 9.3005
R18882 gnd.n2545 gnd.n2529 9.3005
R18883 gnd.n6373 gnd.n2546 9.3005
R18884 gnd.n6372 gnd.n2547 9.3005
R18885 gnd.n6371 gnd.n2548 9.3005
R18886 gnd.n2566 gnd.n2549 9.3005
R18887 gnd.n6361 gnd.n2567 9.3005
R18888 gnd.n6360 gnd.n2568 9.3005
R18889 gnd.n6359 gnd.n2569 9.3005
R18890 gnd.n6484 gnd.n2370 9.3005
R18891 gnd.n6407 gnd.n2454 9.3005
R18892 gnd.n875 gnd.n874 9.3005
R18893 gnd.n6508 gnd.n2342 9.3005
R18894 gnd.n6507 gnd.n2343 9.3005
R18895 gnd.n6506 gnd.n2344 9.3005
R18896 gnd.n2349 gnd.n2345 9.3005
R18897 gnd.n6500 gnd.n2350 9.3005
R18898 gnd.n6499 gnd.n2351 9.3005
R18899 gnd.n6498 gnd.n2352 9.3005
R18900 gnd.n2357 gnd.n2353 9.3005
R18901 gnd.n6492 gnd.n2358 9.3005
R18902 gnd.n6491 gnd.n2359 9.3005
R18903 gnd.n6490 gnd.n2360 9.3005
R18904 gnd.n3920 gnd.n2361 9.3005
R18905 gnd.n3922 gnd.n3921 9.3005
R18906 gnd.n4260 gnd.n4259 9.3005
R18907 gnd.n4261 gnd.n3919 9.3005
R18908 gnd.n4263 gnd.n4262 9.3005
R18909 gnd.n3917 gnd.n3916 9.3005
R18910 gnd.n4268 gnd.n4267 9.3005
R18911 gnd.n4269 gnd.n3915 9.3005
R18912 gnd.n4271 gnd.n4270 9.3005
R18913 gnd.n3913 gnd.n3912 9.3005
R18914 gnd.n4276 gnd.n4275 9.3005
R18915 gnd.n4277 gnd.n3911 9.3005
R18916 gnd.n4284 gnd.n4278 9.3005
R18917 gnd.n4283 gnd.n4279 9.3005
R18918 gnd.n4282 gnd.n4280 9.3005
R18919 gnd.n3884 gnd.n3883 9.3005
R18920 gnd.n4364 gnd.n4363 9.3005
R18921 gnd.n6515 gnd.n6514 9.3005
R18922 gnd.n6518 gnd.n873 9.3005
R18923 gnd.n872 gnd.n868 9.3005
R18924 gnd.n6524 gnd.n867 9.3005
R18925 gnd.n6525 gnd.n866 9.3005
R18926 gnd.n6526 gnd.n865 9.3005
R18927 gnd.n864 gnd.n860 9.3005
R18928 gnd.n6532 gnd.n859 9.3005
R18929 gnd.n6533 gnd.n858 9.3005
R18930 gnd.n6534 gnd.n857 9.3005
R18931 gnd.n856 gnd.n852 9.3005
R18932 gnd.n6540 gnd.n851 9.3005
R18933 gnd.n6541 gnd.n850 9.3005
R18934 gnd.n6542 gnd.n849 9.3005
R18935 gnd.n848 gnd.n844 9.3005
R18936 gnd.n6548 gnd.n843 9.3005
R18937 gnd.n6549 gnd.n842 9.3005
R18938 gnd.n6550 gnd.n841 9.3005
R18939 gnd.n840 gnd.n836 9.3005
R18940 gnd.n6556 gnd.n835 9.3005
R18941 gnd.n6557 gnd.n834 9.3005
R18942 gnd.n6558 gnd.n833 9.3005
R18943 gnd.n832 gnd.n828 9.3005
R18944 gnd.n6564 gnd.n827 9.3005
R18945 gnd.n6565 gnd.n826 9.3005
R18946 gnd.n6566 gnd.n825 9.3005
R18947 gnd.n824 gnd.n820 9.3005
R18948 gnd.n6572 gnd.n819 9.3005
R18949 gnd.n6573 gnd.n818 9.3005
R18950 gnd.n6574 gnd.n817 9.3005
R18951 gnd.n816 gnd.n812 9.3005
R18952 gnd.n6580 gnd.n811 9.3005
R18953 gnd.n6581 gnd.n810 9.3005
R18954 gnd.n6582 gnd.n809 9.3005
R18955 gnd.n808 gnd.n804 9.3005
R18956 gnd.n6588 gnd.n803 9.3005
R18957 gnd.n6589 gnd.n802 9.3005
R18958 gnd.n6590 gnd.n801 9.3005
R18959 gnd.n800 gnd.n796 9.3005
R18960 gnd.n6596 gnd.n795 9.3005
R18961 gnd.n6597 gnd.n794 9.3005
R18962 gnd.n6598 gnd.n793 9.3005
R18963 gnd.n792 gnd.n788 9.3005
R18964 gnd.n6604 gnd.n787 9.3005
R18965 gnd.n6605 gnd.n786 9.3005
R18966 gnd.n6606 gnd.n785 9.3005
R18967 gnd.n784 gnd.n780 9.3005
R18968 gnd.n6612 gnd.n779 9.3005
R18969 gnd.n6613 gnd.n778 9.3005
R18970 gnd.n6614 gnd.n777 9.3005
R18971 gnd.n776 gnd.n772 9.3005
R18972 gnd.n6620 gnd.n771 9.3005
R18973 gnd.n6621 gnd.n770 9.3005
R18974 gnd.n6622 gnd.n769 9.3005
R18975 gnd.n768 gnd.n764 9.3005
R18976 gnd.n6628 gnd.n763 9.3005
R18977 gnd.n6629 gnd.n762 9.3005
R18978 gnd.n6630 gnd.n761 9.3005
R18979 gnd.n760 gnd.n756 9.3005
R18980 gnd.n6636 gnd.n755 9.3005
R18981 gnd.n6637 gnd.n754 9.3005
R18982 gnd.n6638 gnd.n753 9.3005
R18983 gnd.n752 gnd.n748 9.3005
R18984 gnd.n6644 gnd.n747 9.3005
R18985 gnd.n6645 gnd.n746 9.3005
R18986 gnd.n6646 gnd.n745 9.3005
R18987 gnd.n744 gnd.n740 9.3005
R18988 gnd.n6652 gnd.n739 9.3005
R18989 gnd.n6653 gnd.n738 9.3005
R18990 gnd.n6654 gnd.n737 9.3005
R18991 gnd.n736 gnd.n732 9.3005
R18992 gnd.n6660 gnd.n731 9.3005
R18993 gnd.n6661 gnd.n730 9.3005
R18994 gnd.n6662 gnd.n729 9.3005
R18995 gnd.n728 gnd.n724 9.3005
R18996 gnd.n6668 gnd.n723 9.3005
R18997 gnd.n6669 gnd.n722 9.3005
R18998 gnd.n6670 gnd.n721 9.3005
R18999 gnd.n720 gnd.n716 9.3005
R19000 gnd.n6676 gnd.n715 9.3005
R19001 gnd.n6677 gnd.n714 9.3005
R19002 gnd.n6678 gnd.n713 9.3005
R19003 gnd.n712 gnd.n708 9.3005
R19004 gnd.n6684 gnd.n707 9.3005
R19005 gnd.n6686 gnd.n6685 9.3005
R19006 gnd.n6517 gnd.n6516 9.3005
R19007 gnd.n5371 gnd.n5370 9.3005
R19008 gnd.n3836 gnd.n3835 9.3005
R19009 gnd.n3755 gnd.n3754 9.3005
R19010 gnd.n4488 gnd.n4487 9.3005
R19011 gnd.n4489 gnd.n3752 9.3005
R19012 gnd.n4497 gnd.n4496 9.3005
R19013 gnd.n4495 gnd.n3753 9.3005
R19014 gnd.n4494 gnd.n4493 9.3005
R19015 gnd.n4492 gnd.n4491 9.3005
R19016 gnd.n4490 gnd.n3731 9.3005
R19017 gnd.n4542 gnd.n3730 9.3005
R19018 gnd.n4544 gnd.n4543 9.3005
R19019 gnd.n4545 gnd.n3728 9.3005
R19020 gnd.n4552 gnd.n4551 9.3005
R19021 gnd.n4550 gnd.n3729 9.3005
R19022 gnd.n4549 gnd.n4548 9.3005
R19023 gnd.n4547 gnd.n4546 9.3005
R19024 gnd.n3699 gnd.n3698 9.3005
R19025 gnd.n4610 gnd.n4609 9.3005
R19026 gnd.n4611 gnd.n3696 9.3005
R19027 gnd.n4620 gnd.n4619 9.3005
R19028 gnd.n4618 gnd.n3697 9.3005
R19029 gnd.n4617 gnd.n4616 9.3005
R19030 gnd.n4615 gnd.n4612 9.3005
R19031 gnd.n3658 gnd.n3657 9.3005
R19032 gnd.n4698 gnd.n4697 9.3005
R19033 gnd.n4699 gnd.n3655 9.3005
R19034 gnd.n4737 gnd.n4736 9.3005
R19035 gnd.n4735 gnd.n3656 9.3005
R19036 gnd.n4734 gnd.n4733 9.3005
R19037 gnd.n4732 gnd.n4700 9.3005
R19038 gnd.n4731 gnd.n4730 9.3005
R19039 gnd.n4729 gnd.n4704 9.3005
R19040 gnd.n4728 gnd.n4727 9.3005
R19041 gnd.n4726 gnd.n4705 9.3005
R19042 gnd.n4725 gnd.n4724 9.3005
R19043 gnd.n4723 gnd.n4709 9.3005
R19044 gnd.n4722 gnd.n4721 9.3005
R19045 gnd.n4720 gnd.n4710 9.3005
R19046 gnd.n4719 gnd.n4718 9.3005
R19047 gnd.n4717 gnd.n4716 9.3005
R19048 gnd.n3571 gnd.n3570 9.3005
R19049 gnd.n4875 gnd.n4874 9.3005
R19050 gnd.n4876 gnd.n3568 9.3005
R19051 gnd.n4892 gnd.n4891 9.3005
R19052 gnd.n4890 gnd.n3569 9.3005
R19053 gnd.n4889 gnd.n4888 9.3005
R19054 gnd.n4887 gnd.n4877 9.3005
R19055 gnd.n4886 gnd.n4885 9.3005
R19056 gnd.n4884 gnd.n4883 9.3005
R19057 gnd.n3522 gnd.n3521 9.3005
R19058 gnd.n4962 gnd.n4961 9.3005
R19059 gnd.n4963 gnd.n3519 9.3005
R19060 gnd.n4969 gnd.n4968 9.3005
R19061 gnd.n4967 gnd.n3520 9.3005
R19062 gnd.n4966 gnd.n4965 9.3005
R19063 gnd.n3493 gnd.n3492 9.3005
R19064 gnd.n5030 gnd.n5029 9.3005
R19065 gnd.n5031 gnd.n3490 9.3005
R19066 gnd.n5047 gnd.n5046 9.3005
R19067 gnd.n5045 gnd.n3491 9.3005
R19068 gnd.n5044 gnd.n5043 9.3005
R19069 gnd.n5042 gnd.n5032 9.3005
R19070 gnd.n5041 gnd.n5040 9.3005
R19071 gnd.n5039 gnd.n5038 9.3005
R19072 gnd.n3418 gnd.n3417 9.3005
R19073 gnd.n5115 gnd.n5114 9.3005
R19074 gnd.n5116 gnd.n3415 9.3005
R19075 gnd.n5119 gnd.n5118 9.3005
R19076 gnd.n5117 gnd.n3416 9.3005
R19077 gnd.n3388 gnd.n3387 9.3005
R19078 gnd.n5151 gnd.n5150 9.3005
R19079 gnd.n5152 gnd.n3386 9.3005
R19080 gnd.n5154 gnd.n5153 9.3005
R19081 gnd.n3367 gnd.n3366 9.3005
R19082 gnd.n5182 gnd.n5181 9.3005
R19083 gnd.n5183 gnd.n3365 9.3005
R19084 gnd.n5185 gnd.n5184 9.3005
R19085 gnd.n3363 gnd.n3362 9.3005
R19086 gnd.n5192 gnd.n5191 9.3005
R19087 gnd.n5193 gnd.n3360 9.3005
R19088 gnd.n5374 gnd.n5373 9.3005
R19089 gnd.n5372 gnd.n3361 9.3005
R19090 gnd.n3834 gnd.n3833 9.3005
R19091 gnd.n6342 gnd.n2582 9.3005
R19092 gnd.n4348 gnd.n3895 9.3005
R19093 gnd.n4347 gnd.n4346 9.3005
R19094 gnd.n4345 gnd.n3896 9.3005
R19095 gnd.n4344 gnd.n4343 9.3005
R19096 gnd.n3873 gnd.n3872 9.3005
R19097 gnd.n4393 gnd.n4392 9.3005
R19098 gnd.n4394 gnd.n3871 9.3005
R19099 gnd.n4396 gnd.n4395 9.3005
R19100 gnd.n3867 gnd.n3866 9.3005
R19101 gnd.n4407 gnd.n4406 9.3005
R19102 gnd.n4408 gnd.n3865 9.3005
R19103 gnd.n4410 gnd.n4409 9.3005
R19104 gnd.n3860 gnd.n3858 9.3005
R19105 gnd.n4434 gnd.n4433 9.3005
R19106 gnd.n4432 gnd.n3859 9.3005
R19107 gnd.n4431 gnd.n4430 9.3005
R19108 gnd.n4429 gnd.n3861 9.3005
R19109 gnd.n4428 gnd.n4427 9.3005
R19110 gnd.n2581 gnd.n2579 9.3005
R19111 gnd.n6348 gnd.n6347 9.3005
R19112 gnd.n6346 gnd.n2580 9.3005
R19113 gnd.n6320 gnd.n6319 9.3005
R19114 gnd.n6318 gnd.n6317 9.3005
R19115 gnd.n2624 gnd.n2623 9.3005
R19116 gnd.n6312 gnd.n6311 9.3005
R19117 gnd.n6310 gnd.n6309 9.3005
R19118 gnd.n2634 gnd.n2633 9.3005
R19119 gnd.n6304 gnd.n6303 9.3005
R19120 gnd.n6302 gnd.n6301 9.3005
R19121 gnd.n2642 gnd.n2641 9.3005
R19122 gnd.n6296 gnd.n6295 9.3005
R19123 gnd.n6294 gnd.n6293 9.3005
R19124 gnd.n2652 gnd.n2651 9.3005
R19125 gnd.n6288 gnd.n6287 9.3005
R19126 gnd.n6286 gnd.n6285 9.3005
R19127 gnd.n2660 gnd.n2659 9.3005
R19128 gnd.n6280 gnd.n6279 9.3005
R19129 gnd.n6278 gnd.n2674 9.3005
R19130 gnd.n6277 gnd.n2583 9.3005
R19131 gnd.n2620 gnd.n2618 9.3005
R19132 gnd.n6344 gnd.n6343 9.3005
R19133 gnd.n2673 gnd.n2584 9.3005
R19134 gnd.n2669 gnd.n2668 9.3005
R19135 gnd.n6282 gnd.n6281 9.3005
R19136 gnd.n6284 gnd.n6283 9.3005
R19137 gnd.n2656 gnd.n2655 9.3005
R19138 gnd.n6290 gnd.n6289 9.3005
R19139 gnd.n6292 gnd.n6291 9.3005
R19140 gnd.n2648 gnd.n2647 9.3005
R19141 gnd.n6298 gnd.n6297 9.3005
R19142 gnd.n6300 gnd.n6299 9.3005
R19143 gnd.n2638 gnd.n2637 9.3005
R19144 gnd.n6306 gnd.n6305 9.3005
R19145 gnd.n6308 gnd.n6307 9.3005
R19146 gnd.n2630 gnd.n2629 9.3005
R19147 gnd.n6314 gnd.n6313 9.3005
R19148 gnd.n6316 gnd.n6315 9.3005
R19149 gnd.n2619 gnd.n2617 9.3005
R19150 gnd.n6322 gnd.n6321 9.3005
R19151 gnd.n6323 gnd.n2612 9.3005
R19152 gnd.n6325 gnd.n6324 9.3005
R19153 gnd.n6327 gnd.n2611 9.3005
R19154 gnd.n6329 gnd.n6328 9.3005
R19155 gnd.n6330 gnd.n2607 9.3005
R19156 gnd.n6332 gnd.n6331 9.3005
R19157 gnd.n6333 gnd.n2606 9.3005
R19158 gnd.n6335 gnd.n6334 9.3005
R19159 gnd.n6336 gnd.n2605 9.3005
R19160 gnd.n4479 gnd.n4478 9.3005
R19161 gnd.n4480 gnd.n3828 9.3005
R19162 gnd.n4483 gnd.n4482 9.3005
R19163 gnd.n4481 gnd.n3829 9.3005
R19164 gnd.n3743 gnd.n3742 9.3005
R19165 gnd.n4511 gnd.n4510 9.3005
R19166 gnd.n4512 gnd.n3740 9.3005
R19167 gnd.n4515 gnd.n4514 9.3005
R19168 gnd.n4513 gnd.n3741 9.3005
R19169 gnd.n2947 gnd.n2945 9.3005
R19170 gnd.n6126 gnd.n6125 9.3005
R19171 gnd.n6124 gnd.n2946 9.3005
R19172 gnd.n6123 gnd.n6122 9.3005
R19173 gnd.n6121 gnd.n2948 9.3005
R19174 gnd.n6120 gnd.n6119 9.3005
R19175 gnd.n6118 gnd.n2952 9.3005
R19176 gnd.n6117 gnd.n6116 9.3005
R19177 gnd.n6115 gnd.n2953 9.3005
R19178 gnd.n6114 gnd.n6113 9.3005
R19179 gnd.n6112 gnd.n2957 9.3005
R19180 gnd.n6111 gnd.n6110 9.3005
R19181 gnd.n6109 gnd.n2958 9.3005
R19182 gnd.n6108 gnd.n6107 9.3005
R19183 gnd.n6106 gnd.n2962 9.3005
R19184 gnd.n6105 gnd.n6104 9.3005
R19185 gnd.n6103 gnd.n2963 9.3005
R19186 gnd.n6102 gnd.n6101 9.3005
R19187 gnd.n6100 gnd.n2967 9.3005
R19188 gnd.n6099 gnd.n6098 9.3005
R19189 gnd.n6097 gnd.n2968 9.3005
R19190 gnd.n6096 gnd.n6095 9.3005
R19191 gnd.n6094 gnd.n2972 9.3005
R19192 gnd.n6093 gnd.n6092 9.3005
R19193 gnd.n6091 gnd.n2973 9.3005
R19194 gnd.n6090 gnd.n6089 9.3005
R19195 gnd.n6088 gnd.n2977 9.3005
R19196 gnd.n6087 gnd.n6086 9.3005
R19197 gnd.n6085 gnd.n2978 9.3005
R19198 gnd.n6084 gnd.n6083 9.3005
R19199 gnd.n6082 gnd.n2982 9.3005
R19200 gnd.n6081 gnd.n6080 9.3005
R19201 gnd.n6079 gnd.n2983 9.3005
R19202 gnd.n6078 gnd.n6077 9.3005
R19203 gnd.n6076 gnd.n2987 9.3005
R19204 gnd.n6075 gnd.n6074 9.3005
R19205 gnd.n6073 gnd.n2988 9.3005
R19206 gnd.n6072 gnd.n6071 9.3005
R19207 gnd.n6070 gnd.n2992 9.3005
R19208 gnd.n6069 gnd.n6068 9.3005
R19209 gnd.n6067 gnd.n2993 9.3005
R19210 gnd.n6066 gnd.n6065 9.3005
R19211 gnd.n6064 gnd.n2997 9.3005
R19212 gnd.n6063 gnd.n6062 9.3005
R19213 gnd.n6061 gnd.n2998 9.3005
R19214 gnd.n6060 gnd.n6059 9.3005
R19215 gnd.n6058 gnd.n3002 9.3005
R19216 gnd.n6057 gnd.n6056 9.3005
R19217 gnd.n6055 gnd.n3003 9.3005
R19218 gnd.n6054 gnd.n6053 9.3005
R19219 gnd.n6052 gnd.n3007 9.3005
R19220 gnd.n6051 gnd.n6050 9.3005
R19221 gnd.n6049 gnd.n3008 9.3005
R19222 gnd.n6048 gnd.n6047 9.3005
R19223 gnd.n6046 gnd.n3012 9.3005
R19224 gnd.n6045 gnd.n6044 9.3005
R19225 gnd.n6043 gnd.n3013 9.3005
R19226 gnd.n6042 gnd.n6041 9.3005
R19227 gnd.n6040 gnd.n3017 9.3005
R19228 gnd.n6039 gnd.n6038 9.3005
R19229 gnd.n6037 gnd.n3018 9.3005
R19230 gnd.n6036 gnd.n6035 9.3005
R19231 gnd.n6034 gnd.n3022 9.3005
R19232 gnd.n6033 gnd.n6032 9.3005
R19233 gnd.n6031 gnd.n3023 9.3005
R19234 gnd.n6030 gnd.n6029 9.3005
R19235 gnd.n6028 gnd.n3027 9.3005
R19236 gnd.n6027 gnd.n6026 9.3005
R19237 gnd.n6025 gnd.n3028 9.3005
R19238 gnd.n6024 gnd.n6023 9.3005
R19239 gnd.n6022 gnd.n3032 9.3005
R19240 gnd.n6021 gnd.n6020 9.3005
R19241 gnd.n6019 gnd.n3033 9.3005
R19242 gnd.n3831 gnd.n3830 9.3005
R19243 gnd.n5260 gnd.n5259 9.3005
R19244 gnd.n5255 gnd.n5254 9.3005
R19245 gnd.n5267 gnd.n5266 9.3005
R19246 gnd.n5268 gnd.n5253 9.3005
R19247 gnd.n5271 gnd.n5270 9.3005
R19248 gnd.n5269 gnd.n5251 9.3005
R19249 gnd.n5258 gnd.n5257 9.3005
R19250 gnd.n5359 gnd.n5207 9.3005
R19251 gnd.n5220 gnd.n5216 9.3005
R19252 gnd.n5353 gnd.n5352 9.3005
R19253 gnd.n5341 gnd.n5218 9.3005
R19254 gnd.n5340 gnd.n5339 9.3005
R19255 gnd.n5229 gnd.n5225 9.3005
R19256 gnd.n5333 gnd.n5332 9.3005
R19257 gnd.n5322 gnd.n5227 9.3005
R19258 gnd.n5321 gnd.n5320 9.3005
R19259 gnd.n5238 gnd.n5234 9.3005
R19260 gnd.n5314 gnd.n5313 9.3005
R19261 gnd.n5303 gnd.n5236 9.3005
R19262 gnd.n5302 gnd.n5301 9.3005
R19263 gnd.n5247 gnd.n5243 9.3005
R19264 gnd.n5295 gnd.n5294 9.3005
R19265 gnd.n5284 gnd.n5245 9.3005
R19266 gnd.n5283 gnd.n5282 9.3005
R19267 gnd.n5361 gnd.n5360 9.3005
R19268 gnd.n5211 gnd.n5210 9.3005
R19269 gnd.n5278 gnd.n5277 9.3005
R19270 gnd.n5279 gnd.n5250 9.3005
R19271 gnd.n5286 gnd.n5285 9.3005
R19272 gnd.n5248 gnd.n5246 9.3005
R19273 gnd.n5293 gnd.n5292 9.3005
R19274 gnd.n5242 gnd.n5241 9.3005
R19275 gnd.n5305 gnd.n5304 9.3005
R19276 gnd.n5239 gnd.n5237 9.3005
R19277 gnd.n5312 gnd.n5311 9.3005
R19278 gnd.n5233 gnd.n5232 9.3005
R19279 gnd.n5324 gnd.n5323 9.3005
R19280 gnd.n5230 gnd.n5228 9.3005
R19281 gnd.n5331 gnd.n5330 9.3005
R19282 gnd.n5224 gnd.n5223 9.3005
R19283 gnd.n5343 gnd.n5342 9.3005
R19284 gnd.n5221 gnd.n5219 9.3005
R19285 gnd.n5351 gnd.n5350 9.3005
R19286 gnd.n5349 gnd.n5348 9.3005
R19287 gnd.n5363 gnd.n5362 9.3005
R19288 gnd.n5208 gnd.n5202 9.3005
R19289 gnd.n5209 gnd.n5201 9.3005
R19290 gnd.n5197 gnd.n5194 9.3005
R19291 gnd.n3262 gnd.n3261 9.3005
R19292 gnd.n5733 gnd.n5732 9.3005
R19293 gnd.n5734 gnd.n3260 9.3005
R19294 gnd.n5736 gnd.n5735 9.3005
R19295 gnd.n3256 gnd.n3254 9.3005
R19296 gnd.n5756 gnd.n5755 9.3005
R19297 gnd.n5754 gnd.n3255 9.3005
R19298 gnd.n5753 gnd.n5752 9.3005
R19299 gnd.n5751 gnd.n3257 9.3005
R19300 gnd.n5750 gnd.n5749 9.3005
R19301 gnd.n3245 gnd.n3244 9.3005
R19302 gnd.n5813 gnd.n5812 9.3005
R19303 gnd.n5814 gnd.n3242 9.3005
R19304 gnd.n5826 gnd.n5825 9.3005
R19305 gnd.n5824 gnd.n3243 9.3005
R19306 gnd.n5823 gnd.n5822 9.3005
R19307 gnd.n5821 gnd.n5815 9.3005
R19308 gnd.n5820 gnd.n5819 9.3005
R19309 gnd.n5818 gnd.n63 9.3005
R19310 gnd.n5199 gnd.n5198 9.3005
R19311 gnd.n7736 gnd.n64 9.3005
R19312 gnd.t170 gnd.n1065 9.24152
R19313 gnd.n969 gnd.t38 9.24152
R19314 gnd.n2237 gnd.t142 9.24152
R19315 gnd.n4437 gnd.t207 9.24152
R19316 gnd.n4639 gnd.t23 9.24152
R19317 gnd.n5069 gnd.t312 9.24152
R19318 gnd.n5759 gnd.t214 9.24152
R19319 gnd.t326 gnd.t170 8.92286
R19320 gnd.n6150 gnd.n2912 8.92286
R19321 gnd.n4669 gnd.n3679 8.92286
R19322 gnd.n4740 gnd.n4739 8.92286
R19323 gnd.n4847 gnd.n3594 8.92286
R19324 gnd.n4896 gnd.n4895 8.92286
R19325 gnd.n4992 gnd.n3510 8.92286
R19326 gnd.n4977 gnd.n3473 8.92286
R19327 gnd.n3393 gnd.n3383 8.92286
R19328 gnd.n5187 gnd.n3347 8.92286
R19329 gnd.n2207 gnd.n2182 8.92171
R19330 gnd.n2175 gnd.n2150 8.92171
R19331 gnd.n2143 gnd.n2118 8.92171
R19332 gnd.n2112 gnd.n2087 8.92171
R19333 gnd.n2080 gnd.n2055 8.92171
R19334 gnd.n2048 gnd.n2023 8.92171
R19335 gnd.n2016 gnd.n1991 8.92171
R19336 gnd.n1985 gnd.n1960 8.92171
R19337 gnd.n5407 gnd.n5389 8.72777
R19338 gnd.n1709 gnd.t165 8.60421
R19339 gnd.n6220 gnd.n2854 8.60421
R19340 gnd.t30 gnd.n4845 8.60421
R19341 gnd.n4832 gnd.t322 8.60421
R19342 gnd.n1129 gnd.n1117 8.43656
R19343 gnd.n38 gnd.n26 8.43656
R19344 gnd.n4485 gnd.t110 8.28555
R19345 gnd.n4572 gnd.n3693 8.28555
R19346 gnd.n4645 gnd.n3648 8.28555
R19347 gnd.n4802 gnd.n4801 8.28555
R19348 gnd.n4824 gnd.n3561 8.28555
R19349 gnd.n5000 gnd.n4999 8.28555
R19350 gnd.n5077 gnd.n3468 8.28555
R19351 gnd.t124 gnd.n3374 8.28555
R19352 gnd.n2208 gnd.n2180 8.14595
R19353 gnd.n2176 gnd.n2148 8.14595
R19354 gnd.n2144 gnd.n2116 8.14595
R19355 gnd.n2113 gnd.n2085 8.14595
R19356 gnd.n2081 gnd.n2053 8.14595
R19357 gnd.n2049 gnd.n2021 8.14595
R19358 gnd.n2017 gnd.n1989 8.14595
R19359 gnd.n1986 gnd.n1958 8.14595
R19360 gnd.n4349 gnd.n0 8.10675
R19361 gnd.n7737 gnd.n7736 8.10675
R19362 gnd.n2213 gnd.n2212 7.97301
R19363 gnd.t173 gnd.n1224 7.9669
R19364 gnd.n4599 gnd.t175 7.9669
R19365 gnd.n5111 gnd.t320 7.9669
R19366 gnd.n7737 gnd.n62 7.78567
R19367 gnd.n5360 gnd.n5211 7.75808
R19368 gnd.n6278 gnd.n6277 7.75808
R19369 gnd.n7662 gnd.n182 7.75808
R19370 gnd.n3963 gnd.n3956 7.75808
R19371 gnd.t110 gnd.n3825 7.64824
R19372 gnd.n4517 gnd.t155 7.64824
R19373 gnd.n4526 gnd.n3724 7.64824
R19374 gnd.n4572 gnd.t189 7.64824
R19375 gnd.t163 gnd.n3619 7.64824
R19376 gnd.n4706 gnd.t163 7.64824
R19377 gnd.n4881 gnd.t13 7.64824
R19378 gnd.t13 gnd.n3539 7.64824
R19379 gnd.n5077 gnd.t9 7.64824
R19380 gnd.n5139 gnd.n3398 7.64824
R19381 gnd.n5156 gnd.t124 7.64824
R19382 gnd.n1154 gnd.n1153 7.53171
R19383 gnd.n1618 gnd.t3 7.32958
R19384 gnd.n6220 gnd.n2886 7.32958
R19385 gnd.n5542 gnd.n3303 7.32958
R19386 gnd.n2908 gnd.n2907 7.30353
R19387 gnd.n5406 gnd.n5405 7.30353
R19388 gnd.n1578 gnd.n1297 7.01093
R19389 gnd.n1300 gnd.n1298 7.01093
R19390 gnd.n1588 gnd.n1587 7.01093
R19391 gnd.n1599 gnd.n1281 7.01093
R19392 gnd.n1598 gnd.n1284 7.01093
R19393 gnd.n1609 gnd.n1272 7.01093
R19394 gnd.n1275 gnd.n1273 7.01093
R19395 gnd.n1619 gnd.n1618 7.01093
R19396 gnd.n1629 gnd.n1253 7.01093
R19397 gnd.n1628 gnd.n1256 7.01093
R19398 gnd.n1637 gnd.n1247 7.01093
R19399 gnd.n1649 gnd.n1237 7.01093
R19400 gnd.n1659 gnd.n1222 7.01093
R19401 gnd.n1675 gnd.n1674 7.01093
R19402 gnd.n1224 gnd.n1161 7.01093
R19403 gnd.n1729 gnd.n1162 7.01093
R19404 gnd.n1723 gnd.n1722 7.01093
R19405 gnd.n1211 gnd.n1173 7.01093
R19406 gnd.n1715 gnd.n1184 7.01093
R19407 gnd.n1202 gnd.n1197 7.01093
R19408 gnd.n1709 gnd.n1708 7.01093
R19409 gnd.n1755 gnd.n1100 7.01093
R19410 gnd.n1754 gnd.n1753 7.01093
R19411 gnd.n1766 gnd.n1765 7.01093
R19412 gnd.n1093 gnd.n1085 7.01093
R19413 gnd.n1795 gnd.n1073 7.01093
R19414 gnd.n1794 gnd.n1076 7.01093
R19415 gnd.n1805 gnd.n1065 7.01093
R19416 gnd.n1066 gnd.n1054 7.01093
R19417 gnd.n1816 gnd.n1055 7.01093
R19418 gnd.n1842 gnd.n1047 7.01093
R19419 gnd.n1841 gnd.n1840 7.01093
R19420 gnd.n1864 gnd.n1863 7.01093
R19421 gnd.n1882 gnd.n1020 7.01093
R19422 gnd.n1881 gnd.n1023 7.01093
R19423 gnd.n1892 gnd.n1012 7.01093
R19424 gnd.n1013 gnd.n1000 7.01093
R19425 gnd.n1903 gnd.n1001 7.01093
R19426 gnd.n1930 gnd.n985 7.01093
R19427 gnd.n1942 gnd.n1941 7.01093
R19428 gnd.n1924 gnd.n978 7.01093
R19429 gnd.n1953 gnd.n1952 7.01093
R19430 gnd.n2225 gnd.n966 7.01093
R19431 gnd.n2224 gnd.n969 7.01093
R19432 gnd.n2237 gnd.n958 7.01093
R19433 gnd.n959 gnd.n951 7.01093
R19434 gnd.n2247 gnd.n877 7.01093
R19435 gnd.n6150 gnd.n6149 7.01093
R19436 gnd.n4539 gnd.n3733 7.01093
R19437 gnd.n4740 gnd.n3652 7.01093
R19438 gnd.t16 gnd.n3607 7.01093
R19439 gnd.n4847 gnd.n4846 7.01093
R19440 gnd.n4896 gnd.n3565 7.01093
R19441 gnd.t17 gnd.n3549 7.01093
R19442 gnd.n4992 gnd.n4991 7.01093
R19443 gnd.n5158 gnd.n3383 7.01093
R19444 gnd.n5384 gnd.n3347 7.01093
R19445 gnd.n5187 gnd.t91 7.01093
R19446 gnd.n1256 gnd.t167 6.69227
R19447 gnd.n1076 gnd.t326 6.69227
R19448 gnd.n1840 gnd.n870 6.69227
R19449 gnd.n1931 gnd.t10 6.69227
R19450 gnd.n4623 gnd.t23 6.69227
R19451 gnd.n5035 gnd.t312 6.69227
R19452 gnd.n5536 gnd.n5535 6.5566
R19453 gnd.n3764 gnd.n3763 6.5566
R19454 gnd.n6161 gnd.n6157 6.5566
R19455 gnd.n5414 gnd.n5413 6.5566
R19456 gnd.n4568 gnd.n3719 6.37362
R19457 gnd.n4606 gnd.n4605 6.37362
R19458 gnd.n4765 gnd.n3631 6.37362
R19459 gnd.n4959 gnd.n4958 6.37362
R19460 gnd.n5105 gnd.n5104 6.37362
R19461 gnd.n5122 gnd.n3405 6.37362
R19462 gnd.n2668 gnd.n2666 6.20656
R19463 gnd.n5363 gnd.n5206 6.20656
R19464 gnd.t178 gnd.n1685 6.05496
R19465 gnd.n1686 gnd.t159 6.05496
R19466 gnd.t316 gnd.n1100 6.05496
R19467 gnd.t158 gnd.n1852 6.05496
R19468 gnd.n4257 gnd.t55 6.05496
R19469 gnd.n176 gnd.t59 6.05496
R19470 gnd.n2210 gnd.n2180 5.81868
R19471 gnd.n2178 gnd.n2148 5.81868
R19472 gnd.n2146 gnd.n2116 5.81868
R19473 gnd.n2115 gnd.n2085 5.81868
R19474 gnd.n2083 gnd.n2053 5.81868
R19475 gnd.n2051 gnd.n2021 5.81868
R19476 gnd.n2019 gnd.n1989 5.81868
R19477 gnd.n1988 gnd.n1958 5.81868
R19478 gnd.n4518 gnd.n2924 5.73631
R19479 gnd.t52 gnd.n4539 5.73631
R19480 gnd.n4669 gnd.t33 5.73631
R19481 gnd.n4661 gnd.n4660 5.73631
R19482 gnd.n4686 gnd.n3666 5.73631
R19483 gnd.t184 gnd.n3625 5.73631
R19484 gnd.n4846 gnd.t177 5.73631
R19485 gnd.n4839 gnd.n3579 5.73631
R19486 gnd.n4864 gnd.n3573 5.73631
R19487 gnd.t28 gnd.n3565 5.73631
R19488 gnd.n3532 gnd.t190 5.73631
R19489 gnd.n5026 gnd.n3497 5.73631
R19490 gnd.n5050 gnd.n3487 5.73631
R19491 gnd.n4977 gnd.t5 5.73631
R19492 gnd.n5170 gnd.n5169 5.73631
R19493 gnd.n5475 gnd.t91 5.73631
R19494 gnd.n5545 gnd.n3299 5.62001
R19495 gnd.n6223 gnd.n2850 5.62001
R19496 gnd.n6223 gnd.n2851 5.62001
R19497 gnd.n5545 gnd.n3300 5.62001
R19498 gnd.n1437 gnd.n1432 5.4308
R19499 gnd.n2255 gnd.n944 5.4308
R19500 gnd.n1753 gnd.t4 5.41765
R19501 gnd.t157 gnd.n1776 5.41765
R19502 gnd.t20 gnd.n1032 5.41765
R19503 gnd.n4695 gnd.t18 5.41765
R19504 gnd.n5027 gnd.t324 5.41765
R19505 gnd.n4587 gnd.n4586 5.09899
R19506 gnd.n4599 gnd.n4598 5.09899
R19507 gnd.t32 gnd.n3636 5.09899
R19508 gnd.n4776 gnd.n4774 5.09899
R19509 gnd.n4787 gnd.n4786 5.09899
R19510 gnd.n4931 gnd.n4930 5.09899
R19511 gnd.n4951 gnd.n4950 5.09899
R19512 gnd.n4971 gnd.t34 5.09899
R19513 gnd.n5112 gnd.n5111 5.09899
R19514 gnd.n5097 gnd.n5096 5.09899
R19515 gnd.n2208 gnd.n2207 5.04292
R19516 gnd.n2176 gnd.n2175 5.04292
R19517 gnd.n2144 gnd.n2143 5.04292
R19518 gnd.n2113 gnd.n2112 5.04292
R19519 gnd.n2081 gnd.n2080 5.04292
R19520 gnd.n2049 gnd.n2048 5.04292
R19521 gnd.n2017 gnd.n2016 5.04292
R19522 gnd.n1986 gnd.n1985 5.04292
R19523 gnd.n1716 gnd.t12 4.78034
R19524 gnd.n1055 gnd.t174 4.78034
R19525 gnd.n6143 gnd.t7 4.78034
R19526 gnd.n3666 gnd.t18 4.78034
R19527 gnd.t324 gnd.n5026 4.78034
R19528 gnd.t25 gnd.n3432 4.78034
R19529 gnd.n5542 gnd.t67 4.78034
R19530 gnd.n1158 gnd.n1155 4.74817
R19531 gnd.n1208 gnd.n1106 4.74817
R19532 gnd.n1195 gnd.n1105 4.74817
R19533 gnd.n1104 gnd.n1103 4.74817
R19534 gnd.n1204 gnd.n1155 4.74817
R19535 gnd.n1205 gnd.n1106 4.74817
R19536 gnd.n1207 gnd.n1105 4.74817
R19537 gnd.n1194 gnd.n1104 4.74817
R19538 gnd.n3146 gnd.n82 4.74817
R19539 gnd.n5937 gnd.n81 4.74817
R19540 gnd.n3163 gnd.n80 4.74817
R19541 gnd.n7729 gnd.n75 4.74817
R19542 gnd.n7727 gnd.n76 4.74817
R19543 gnd.n5951 gnd.n82 4.74817
R19544 gnd.n3145 gnd.n81 4.74817
R19545 gnd.n5938 gnd.n80 4.74817
R19546 gnd.n3162 gnd.n75 4.74817
R19547 gnd.n7728 gnd.n7727 4.74817
R19548 gnd.n3885 gnd.n3882 4.74817
R19549 gnd.n3889 gnd.n3881 4.74817
R19550 gnd.n4328 gnd.n3880 4.74817
R19551 gnd.n4326 gnd.n3879 4.74817
R19552 gnd.n4322 gnd.n3878 4.74817
R19553 gnd.n5946 gnd.n3152 4.74817
R19554 gnd.n5944 gnd.n5943 4.74817
R19555 gnd.n3177 gnd.n3176 4.74817
R19556 gnd.n3182 gnd.n3181 4.74817
R19557 gnd.n5924 gnd.n5923 4.74817
R19558 gnd.n5793 gnd.n3152 4.74817
R19559 gnd.n5945 gnd.n5944 4.74817
R19560 gnd.n3176 gnd.n3153 4.74817
R19561 gnd.n3181 gnd.n3180 4.74817
R19562 gnd.n5925 gnd.n5924 4.74817
R19563 gnd.n6435 gnd.n6434 4.74817
R19564 gnd.n2471 gnd.n2455 4.74817
R19565 gnd.n6422 gnd.n6421 4.74817
R19566 gnd.n2488 gnd.n2472 4.74817
R19567 gnd.n6409 gnd.n6408 4.74817
R19568 gnd.n6436 gnd.n6435 4.74817
R19569 gnd.n6433 gnd.n2455 4.74817
R19570 gnd.n6423 gnd.n6422 4.74817
R19571 gnd.n6420 gnd.n2472 4.74817
R19572 gnd.n6410 gnd.n6409 4.74817
R19573 gnd.n4359 gnd.n3882 4.74817
R19574 gnd.n4358 gnd.n3881 4.74817
R19575 gnd.n3888 gnd.n3880 4.74817
R19576 gnd.n4329 gnd.n3879 4.74817
R19577 gnd.n4325 gnd.n3878 4.74817
R19578 gnd.n1153 gnd.n1152 4.74296
R19579 gnd.n62 gnd.n61 4.74296
R19580 gnd.n1129 gnd.n1128 4.7074
R19581 gnd.n1141 gnd.n1140 4.7074
R19582 gnd.n38 gnd.n37 4.7074
R19583 gnd.n50 gnd.n49 4.7074
R19584 gnd.n1153 gnd.n1141 4.65959
R19585 gnd.n62 gnd.n50 4.65959
R19586 gnd.n5636 gnd.n5546 4.6132
R19587 gnd.n6224 gnd.n2849 4.6132
R19588 gnd.n4499 gnd.n3747 4.46168
R19589 gnd.n6136 gnd.n6135 4.46168
R19590 gnd.n4526 gnd.t181 4.46168
R19591 gnd.n4676 gnd.n4675 4.46168
R19592 gnd.n4694 gnd.n3661 4.46168
R19593 gnd.n4854 gnd.n4853 4.46168
R19594 gnd.n4871 gnd.n3575 4.46168
R19595 gnd.n5017 gnd.n3495 4.46168
R19596 gnd.n5059 gnd.n3480 4.46168
R19597 gnd.n5139 gnd.t180 4.46168
R19598 gnd.n5172 gnd.n3374 4.46168
R19599 gnd.n3434 gnd.n3433 4.46168
R19600 gnd.n5402 gnd.n5389 4.46111
R19601 gnd.n2193 gnd.n2189 4.38594
R19602 gnd.n2161 gnd.n2157 4.38594
R19603 gnd.n2129 gnd.n2125 4.38594
R19604 gnd.n2098 gnd.n2094 4.38594
R19605 gnd.n2066 gnd.n2062 4.38594
R19606 gnd.n2034 gnd.n2030 4.38594
R19607 gnd.n2002 gnd.n1998 4.38594
R19608 gnd.n1971 gnd.n1967 4.38594
R19609 gnd.n2204 gnd.n2182 4.26717
R19610 gnd.n2172 gnd.n2150 4.26717
R19611 gnd.n2140 gnd.n2118 4.26717
R19612 gnd.n2109 gnd.n2087 4.26717
R19613 gnd.n2077 gnd.n2055 4.26717
R19614 gnd.n2045 gnd.n2023 4.26717
R19615 gnd.n2013 gnd.n1991 4.26717
R19616 gnd.n1982 gnd.n1960 4.26717
R19617 gnd.n1660 gnd.t11 4.14303
R19618 gnd.n1892 gnd.t166 4.14303
R19619 gnd.t87 gnd.n2564 4.14303
R19620 gnd.n4793 gnd.t314 4.14303
R19621 gnd.n4920 gnd.t35 4.14303
R19622 gnd.t63 gnd.n3068 4.14303
R19623 gnd.n2212 gnd.n2211 4.08274
R19624 gnd.n5535 gnd.n5534 4.05904
R19625 gnd.n3765 gnd.n3764 4.05904
R19626 gnd.n6164 gnd.n6157 4.05904
R19627 gnd.n5415 gnd.n5414 4.05904
R19628 gnd.n15 gnd.n7 3.99943
R19629 gnd.n1733 gnd.n1154 3.9165
R19630 gnd.n6136 gnd.t155 3.82437
R19631 gnd.t181 gnd.n4525 3.82437
R19632 gnd.n4555 gnd.n4554 3.82437
R19633 gnd.n4576 gnd.n3688 3.82437
R19634 gnd.t22 gnd.n3652 3.82437
R19635 gnd.n3639 gnd.n3638 3.82437
R19636 gnd.n4795 gnd.n3604 3.82437
R19637 gnd.n3552 gnd.n3551 3.82437
R19638 gnd.n4942 gnd.n4940 3.82437
R19639 gnd.n4991 gnd.t29 3.82437
R19640 gnd.n5085 gnd.n5083 3.82437
R19641 gnd.n5129 gnd.n3407 3.82437
R19642 gnd.t180 gnd.n5138 3.82437
R19643 gnd.n3358 gnd.t67 3.82437
R19644 gnd.n1141 gnd.n1129 3.72967
R19645 gnd.n50 gnd.n38 3.72967
R19646 gnd.n2212 gnd.n2084 3.70378
R19647 gnd.n15 gnd.n14 3.60163
R19648 gnd.n2203 gnd.n2184 3.49141
R19649 gnd.n2171 gnd.n2152 3.49141
R19650 gnd.n2139 gnd.n2120 3.49141
R19651 gnd.n2108 gnd.n2089 3.49141
R19652 gnd.n2076 gnd.n2057 3.49141
R19653 gnd.n2044 gnd.n2025 3.49141
R19654 gnd.n2012 gnd.n1993 3.49141
R19655 gnd.n1981 gnd.n1962 3.49141
R19656 gnd.n5617 gnd.n5616 3.29747
R19657 gnd.n5616 gnd.n5554 3.29747
R19658 gnd.n7626 gnd.n7623 3.29747
R19659 gnd.n7627 gnd.n7626 3.29747
R19660 gnd.n4106 gnd.n4047 3.29747
R19661 gnd.n4047 gnd.n4042 3.29747
R19662 gnd.n6242 gnd.n6241 3.29747
R19663 gnd.n6241 gnd.n6240 3.29747
R19664 gnd.n3825 gnd.n3824 3.18706
R19665 gnd.n4540 gnd.t52 3.18706
R19666 gnd.n6129 gnd.n2940 3.18706
R19667 gnd.n4640 gnd.n4639 3.18706
R19668 gnd.n4749 gnd.n3645 3.18706
R19669 gnd.n4819 gnd.n4818 3.18706
R19670 gnd.n4904 gnd.n3558 3.18706
R19671 gnd.n5007 gnd.n5006 3.18706
R19672 gnd.n5070 gnd.n5069 3.18706
R19673 gnd.n5147 gnd.n5146 3.18706
R19674 gnd.n5179 gnd.t101 3.18706
R19675 gnd.n5475 gnd.n3340 3.18706
R19676 gnd.n1239 gnd.t11 2.8684
R19677 gnd.n4585 gnd.t175 2.8684
R19678 gnd.n5095 gnd.t320 2.8684
R19679 gnd.n1142 gnd.t234 2.82907
R19680 gnd.n1142 gnd.t295 2.82907
R19681 gnd.n1144 gnd.t213 2.82907
R19682 gnd.n1144 gnd.t248 2.82907
R19683 gnd.n1146 gnd.t265 2.82907
R19684 gnd.n1146 gnd.t254 2.82907
R19685 gnd.n1148 gnd.t252 2.82907
R19686 gnd.n1148 gnd.t243 2.82907
R19687 gnd.n1150 gnd.t257 2.82907
R19688 gnd.n1150 gnd.t284 2.82907
R19689 gnd.n1107 gnd.t259 2.82907
R19690 gnd.n1107 gnd.t274 2.82907
R19691 gnd.n1109 gnd.t280 2.82907
R19692 gnd.n1109 gnd.t236 2.82907
R19693 gnd.n1111 gnd.t273 2.82907
R19694 gnd.n1111 gnd.t269 2.82907
R19695 gnd.n1113 gnd.t306 2.82907
R19696 gnd.n1113 gnd.t297 2.82907
R19697 gnd.n1115 gnd.t241 2.82907
R19698 gnd.n1115 gnd.t278 2.82907
R19699 gnd.n1118 gnd.t309 2.82907
R19700 gnd.n1118 gnd.t218 2.82907
R19701 gnd.n1120 gnd.t219 2.82907
R19702 gnd.n1120 gnd.t202 2.82907
R19703 gnd.n1122 gnd.t283 2.82907
R19704 gnd.n1122 gnd.t310 2.82907
R19705 gnd.n1124 gnd.t304 2.82907
R19706 gnd.n1124 gnd.t221 2.82907
R19707 gnd.n1126 gnd.t298 2.82907
R19708 gnd.n1126 gnd.t282 2.82907
R19709 gnd.n1130 gnd.t271 2.82907
R19710 gnd.n1130 gnd.t237 2.82907
R19711 gnd.n1132 gnd.t258 2.82907
R19712 gnd.n1132 gnd.t281 2.82907
R19713 gnd.n1134 gnd.t303 2.82907
R19714 gnd.n1134 gnd.t292 2.82907
R19715 gnd.n1136 gnd.t290 2.82907
R19716 gnd.n1136 gnd.t277 2.82907
R19717 gnd.n1138 gnd.t294 2.82907
R19718 gnd.n1138 gnd.t228 2.82907
R19719 gnd.n59 gnd.t261 2.82907
R19720 gnd.n59 gnd.t242 2.82907
R19721 gnd.n57 gnd.t209 2.82907
R19722 gnd.n57 gnd.t226 2.82907
R19723 gnd.n55 gnd.t230 2.82907
R19724 gnd.n55 gnd.t245 2.82907
R19725 gnd.n53 gnd.t223 2.82907
R19726 gnd.n53 gnd.t291 2.82907
R19727 gnd.n51 gnd.t270 2.82907
R19728 gnd.n51 gnd.t206 2.82907
R19729 gnd.n24 gnd.t311 2.82907
R19730 gnd.n24 gnd.t232 2.82907
R19731 gnd.n22 gnd.t216 2.82907
R19732 gnd.n22 gnd.t231 2.82907
R19733 gnd.n20 gnd.t289 2.82907
R19734 gnd.n20 gnd.t266 2.82907
R19735 gnd.n18 gnd.t256 2.82907
R19736 gnd.n18 gnd.t200 2.82907
R19737 gnd.n16 gnd.t302 2.82907
R19738 gnd.n16 gnd.t246 2.82907
R19739 gnd.n35 gnd.t272 2.82907
R19740 gnd.n35 gnd.t199 2.82907
R19741 gnd.n33 gnd.t195 2.82907
R19742 gnd.n33 gnd.t286 2.82907
R19743 gnd.n31 gnd.t293 2.82907
R19744 gnd.n31 gnd.t300 2.82907
R19745 gnd.n29 gnd.t299 2.82907
R19746 gnd.n29 gnd.t197 2.82907
R19747 gnd.n27 gnd.t193 2.82907
R19748 gnd.n27 gnd.t211 2.82907
R19749 gnd.n47 gnd.t301 2.82907
R19750 gnd.n47 gnd.t276 2.82907
R19751 gnd.n45 gnd.t255 2.82907
R19752 gnd.n45 gnd.t267 2.82907
R19753 gnd.n43 gnd.t268 2.82907
R19754 gnd.n43 gnd.t279 2.82907
R19755 gnd.n41 gnd.t262 2.82907
R19756 gnd.n41 gnd.t235 2.82907
R19757 gnd.n39 gnd.t308 2.82907
R19758 gnd.n39 gnd.t250 2.82907
R19759 gnd.n2200 gnd.n2199 2.71565
R19760 gnd.n2168 gnd.n2167 2.71565
R19761 gnd.n2136 gnd.n2135 2.71565
R19762 gnd.n2105 gnd.n2104 2.71565
R19763 gnd.n2073 gnd.n2072 2.71565
R19764 gnd.n2041 gnd.n2040 2.71565
R19765 gnd.n2009 gnd.n2008 2.71565
R19766 gnd.n1978 gnd.n1977 2.71565
R19767 gnd.n6143 gnd.t73 2.54975
R19768 gnd.n6128 gnd.n2942 2.54975
R19769 gnd.n3719 gnd.t6 2.54975
R19770 gnd.n4624 gnd.n4623 2.54975
R19771 gnd.n4688 gnd.t27 2.54975
R19772 gnd.n4748 gnd.n4746 2.54975
R19773 gnd.n4645 gnd.t32 2.54975
R19774 gnd.n4803 gnd.n3598 2.54975
R19775 gnd.n4903 gnd.n4902 2.54975
R19776 gnd.n5000 gnd.t34 2.54975
R19777 gnd.n4998 gnd.n3508 2.54975
R19778 gnd.n4984 gnd.t164 2.54975
R19779 gnd.n5035 gnd.n5034 2.54975
R19780 gnd.t160 gnd.n5122 2.54975
R19781 gnd.n5148 gnd.n3390 2.54975
R19782 gnd.n1733 gnd.n1155 2.27742
R19783 gnd.n1733 gnd.n1106 2.27742
R19784 gnd.n1733 gnd.n1105 2.27742
R19785 gnd.n1733 gnd.n1104 2.27742
R19786 gnd.n7726 gnd.n82 2.27742
R19787 gnd.n7726 gnd.n81 2.27742
R19788 gnd.n7726 gnd.n80 2.27742
R19789 gnd.n7726 gnd.n75 2.27742
R19790 gnd.n7727 gnd.n7726 2.27742
R19791 gnd.n3152 gnd.n79 2.27742
R19792 gnd.n5944 gnd.n79 2.27742
R19793 gnd.n3176 gnd.n79 2.27742
R19794 gnd.n3181 gnd.n79 2.27742
R19795 gnd.n5924 gnd.n79 2.27742
R19796 gnd.n6435 gnd.n2454 2.27742
R19797 gnd.n2455 gnd.n2454 2.27742
R19798 gnd.n6422 gnd.n2454 2.27742
R19799 gnd.n2472 gnd.n2454 2.27742
R19800 gnd.n6409 gnd.n2454 2.27742
R19801 gnd.n4365 gnd.n3882 2.27742
R19802 gnd.n4365 gnd.n3881 2.27742
R19803 gnd.n4365 gnd.n3880 2.27742
R19804 gnd.n4365 gnd.n3879 2.27742
R19805 gnd.n4365 gnd.n3878 2.27742
R19806 gnd.n1587 gnd.t117 2.23109
R19807 gnd.n1210 gnd.t12 2.23109
R19808 gnd.n4706 gnd.t314 2.23109
R19809 gnd.n4881 gnd.t35 2.23109
R19810 gnd.n2196 gnd.n2186 1.93989
R19811 gnd.n2164 gnd.n2154 1.93989
R19812 gnd.n2132 gnd.n2122 1.93989
R19813 gnd.n2101 gnd.n2091 1.93989
R19814 gnd.n2069 gnd.n2059 1.93989
R19815 gnd.n2037 gnd.n2027 1.93989
R19816 gnd.n2005 gnd.n1995 1.93989
R19817 gnd.n1974 gnd.n1964 1.93989
R19818 gnd.n4561 gnd.n4560 1.91244
R19819 gnd.n4631 gnd.n4630 1.91244
R19820 gnd.n4810 gnd.n4809 1.91244
R19821 gnd.n4913 gnd.n4912 1.91244
R19822 gnd.n5086 gnd.n3463 1.91244
R19823 gnd.n3451 gnd.n3450 1.91244
R19824 gnd.n3433 gnd.t42 1.91244
R19825 gnd.t14 gnd.n1598 1.59378
R19826 gnd.n1777 gnd.t157 1.59378
R19827 gnd.n1040 gnd.t20 1.59378
R19828 gnd.t318 gnd.n4757 1.59378
R19829 gnd.n4943 gnd.t182 1.59378
R19830 gnd.n4501 gnd.t45 1.27512
R19831 gnd.n4501 gnd.n4500 1.27512
R19832 gnd.n3734 gnd.n2932 1.27512
R19833 gnd.t33 gnd.n4668 1.27512
R19834 gnd.n4667 gnd.n3673 1.27512
R19835 gnd.n4653 gnd.n4652 1.27512
R19836 gnd.n4845 gnd.n3587 1.27512
R19837 gnd.n4832 gnd.n4831 1.27512
R19838 gnd.n5020 gnd.n5019 1.27512
R19839 gnd.n5058 gnd.n5056 1.27512
R19840 gnd.t5 gnd.n3483 1.27512
R19841 gnd.n5157 gnd.n5156 1.27512
R19842 gnd.n5385 gnd.n3345 1.27512
R19843 gnd.n1440 gnd.n1432 1.16414
R19844 gnd.n2258 gnd.n944 1.16414
R19845 gnd.n2195 gnd.n2188 1.16414
R19846 gnd.n2163 gnd.n2156 1.16414
R19847 gnd.n2131 gnd.n2124 1.16414
R19848 gnd.n2100 gnd.n2093 1.16414
R19849 gnd.n2068 gnd.n2061 1.16414
R19850 gnd.n2036 gnd.n2029 1.16414
R19851 gnd.n2004 gnd.n1997 1.16414
R19852 gnd.n1973 gnd.n1966 1.16414
R19853 gnd.n5546 gnd.n3298 0.970197
R19854 gnd.n6224 gnd.n2751 0.970197
R19855 gnd.n2179 gnd.n2147 0.962709
R19856 gnd.n2211 gnd.n2179 0.962709
R19857 gnd.n2052 gnd.n2020 0.962709
R19858 gnd.n2084 gnd.n2052 0.962709
R19859 gnd.n1686 gnd.t178 0.956468
R19860 gnd.n1853 gnd.t158 0.956468
R19861 gnd.t203 gnd.n2400 0.956468
R19862 gnd.n4232 gnd.t240 0.956468
R19863 gnd.n3868 gnd.t233 0.956468
R19864 gnd.n4412 gnd.t217 0.956468
R19865 gnd.n4507 gnd.t7 0.956468
R19866 gnd.t1 gnd.n6128 0.956468
R19867 gnd.n5148 gnd.t185 0.956468
R19868 gnd.n3437 gnd.t25 0.956468
R19869 gnd.n5747 gnd.t192 0.956468
R19870 gnd.n5802 gnd.t205 0.956468
R19871 gnd.n5907 gnd.t198 0.956468
R19872 gnd.t238 gnd.n138 0.956468
R19873 gnd.n2 gnd.n1 0.672012
R19874 gnd.n3 gnd.n2 0.672012
R19875 gnd.n4 gnd.n3 0.672012
R19876 gnd.n5 gnd.n4 0.672012
R19877 gnd.n6 gnd.n5 0.672012
R19878 gnd.n7 gnd.n6 0.672012
R19879 gnd.n9 gnd.n8 0.672012
R19880 gnd.n10 gnd.n9 0.672012
R19881 gnd.n11 gnd.n10 0.672012
R19882 gnd.n12 gnd.n11 0.672012
R19883 gnd.n13 gnd.n12 0.672012
R19884 gnd.n14 gnd.n13 0.672012
R19885 gnd.t83 gnd.n6142 0.637812
R19886 gnd.n4588 gnd.n3713 0.637812
R19887 gnd.n4596 gnd.n3707 0.637812
R19888 gnd.n3707 gnd.t0 0.637812
R19889 gnd.n4777 gnd.n3625 0.637812
R19890 gnd.n4785 gnd.n3619 0.637812
R19891 gnd.n4801 gnd.t16 0.637812
R19892 gnd.n4824 gnd.t17 0.637812
R19893 gnd.n4932 gnd.n3539 0.637812
R19894 gnd.n4949 gnd.n3532 0.637812
R19895 gnd.t191 gnd.n5103 0.637812
R19896 gnd.n5103 gnd.n3420 0.637812
R19897 gnd.n5123 gnd.n3411 0.637812
R19898 gnd.n5179 gnd.t76 0.637812
R19899 gnd.n1152 gnd.n1151 0.573776
R19900 gnd.n1151 gnd.n1149 0.573776
R19901 gnd.n1149 gnd.n1147 0.573776
R19902 gnd.n1147 gnd.n1145 0.573776
R19903 gnd.n1145 gnd.n1143 0.573776
R19904 gnd.n1117 gnd.n1116 0.573776
R19905 gnd.n1116 gnd.n1114 0.573776
R19906 gnd.n1114 gnd.n1112 0.573776
R19907 gnd.n1112 gnd.n1110 0.573776
R19908 gnd.n1110 gnd.n1108 0.573776
R19909 gnd.n1128 gnd.n1127 0.573776
R19910 gnd.n1127 gnd.n1125 0.573776
R19911 gnd.n1125 gnd.n1123 0.573776
R19912 gnd.n1123 gnd.n1121 0.573776
R19913 gnd.n1121 gnd.n1119 0.573776
R19914 gnd.n1140 gnd.n1139 0.573776
R19915 gnd.n1139 gnd.n1137 0.573776
R19916 gnd.n1137 gnd.n1135 0.573776
R19917 gnd.n1135 gnd.n1133 0.573776
R19918 gnd.n1133 gnd.n1131 0.573776
R19919 gnd.n54 gnd.n52 0.573776
R19920 gnd.n56 gnd.n54 0.573776
R19921 gnd.n58 gnd.n56 0.573776
R19922 gnd.n60 gnd.n58 0.573776
R19923 gnd.n61 gnd.n60 0.573776
R19924 gnd.n19 gnd.n17 0.573776
R19925 gnd.n21 gnd.n19 0.573776
R19926 gnd.n23 gnd.n21 0.573776
R19927 gnd.n25 gnd.n23 0.573776
R19928 gnd.n26 gnd.n25 0.573776
R19929 gnd.n30 gnd.n28 0.573776
R19930 gnd.n32 gnd.n30 0.573776
R19931 gnd.n34 gnd.n32 0.573776
R19932 gnd.n36 gnd.n34 0.573776
R19933 gnd.n37 gnd.n36 0.573776
R19934 gnd.n42 gnd.n40 0.573776
R19935 gnd.n44 gnd.n42 0.573776
R19936 gnd.n46 gnd.n44 0.573776
R19937 gnd.n48 gnd.n46 0.573776
R19938 gnd.n49 gnd.n48 0.573776
R19939 gnd gnd.n0 0.551497
R19940 gnd.n7664 gnd.n7663 0.532512
R19941 gnd.n3959 gnd.n3958 0.532512
R19942 gnd.n7479 gnd.n166 0.497451
R19943 gnd.n2723 gnd.n2569 0.497451
R19944 gnd.n5572 gnd.n3063 0.497451
R19945 gnd.n4062 gnd.n2370 0.497451
R19946 gnd.n5372 gnd.n5371 0.489829
R19947 gnd.n3834 gnd.n2582 0.489829
R19948 gnd.n3830 gnd.n2605 0.489829
R19949 gnd.n5258 gnd.n3033 0.489829
R19950 gnd.n1915 gnd.n948 0.486781
R19951 gnd.n1489 gnd.n1488 0.48678
R19952 gnd.n2232 gnd.n902 0.480683
R19953 gnd.n1573 gnd.n1572 0.480683
R19954 gnd.n7738 gnd.n7737 0.470187
R19955 gnd.n6687 gnd.n6686 0.468488
R19956 gnd.n7208 gnd.n7207 0.468488
R19957 gnd.n7419 gnd.n7418 0.468488
R19958 gnd.n6516 gnd.n6515 0.468488
R19959 gnd.n7726 gnd.n79 0.4255
R19960 gnd.n4365 gnd.n2454 0.4255
R19961 gnd.n6282 gnd.n2666 0.388379
R19962 gnd.n2192 gnd.n2191 0.388379
R19963 gnd.n2160 gnd.n2159 0.388379
R19964 gnd.n2128 gnd.n2127 0.388379
R19965 gnd.n2097 gnd.n2096 0.388379
R19966 gnd.n2065 gnd.n2064 0.388379
R19967 gnd.n2033 gnd.n2032 0.388379
R19968 gnd.n2001 gnd.n2000 0.388379
R19969 gnd.n1970 gnd.n1969 0.388379
R19970 gnd.n5349 gnd.n5206 0.388379
R19971 gnd.n7738 gnd.n15 0.374463
R19972 gnd.n1003 gnd.t10 0.319156
R19973 gnd.t251 gnd.n2441 0.319156
R19974 gnd.n4310 gnd.t220 0.319156
R19975 gnd.n4331 gnd.t253 0.319156
R19976 gnd.n4341 gnd.t212 0.319156
R19977 gnd.n4475 gnd.t113 0.319156
R19978 gnd.n4758 gnd.t318 0.319156
R19979 gnd.t177 gnd.t30 0.319156
R19980 gnd.t322 gnd.t28 0.319156
R19981 gnd.n4972 gnd.t182 0.319156
R19982 gnd.n5377 gnd.t94 0.319156
R19983 gnd.n5949 gnd.t196 0.319156
R19984 gnd.n5941 gnd.t229 0.319156
R19985 gnd.n5855 gnd.t194 0.319156
R19986 gnd.t225 gnd.n98 0.319156
R19987 gnd.n1407 gnd.n1385 0.311721
R19988 gnd.n6346 gnd.n6345 0.302329
R19989 gnd.n5200 gnd.n5199 0.302329
R19990 gnd gnd.n7738 0.295112
R19991 gnd.n201 gnd.n174 0.293183
R19992 gnd.n4212 gnd.n3999 0.293183
R19993 gnd.n2303 gnd.n2302 0.268793
R19994 gnd.n7540 gnd.n174 0.258122
R19995 gnd.n5722 gnd.n5721 0.258122
R19996 gnd.n2784 gnd.n2577 0.258122
R19997 gnd.n4212 gnd.n4211 0.258122
R19998 gnd.n2302 gnd.n2301 0.241354
R19999 gnd.n5637 gnd.n5636 0.229039
R20000 gnd.n5636 gnd.n3297 0.229039
R20001 gnd.n2849 gnd.n2750 0.229039
R20002 gnd.n2849 gnd.n2848 0.229039
R20003 gnd.n1561 gnd.n1360 0.206293
R20004 gnd.n2209 gnd.n2181 0.155672
R20005 gnd.n2202 gnd.n2181 0.155672
R20006 gnd.n2202 gnd.n2201 0.155672
R20007 gnd.n2201 gnd.n2185 0.155672
R20008 gnd.n2194 gnd.n2185 0.155672
R20009 gnd.n2194 gnd.n2193 0.155672
R20010 gnd.n2177 gnd.n2149 0.155672
R20011 gnd.n2170 gnd.n2149 0.155672
R20012 gnd.n2170 gnd.n2169 0.155672
R20013 gnd.n2169 gnd.n2153 0.155672
R20014 gnd.n2162 gnd.n2153 0.155672
R20015 gnd.n2162 gnd.n2161 0.155672
R20016 gnd.n2145 gnd.n2117 0.155672
R20017 gnd.n2138 gnd.n2117 0.155672
R20018 gnd.n2138 gnd.n2137 0.155672
R20019 gnd.n2137 gnd.n2121 0.155672
R20020 gnd.n2130 gnd.n2121 0.155672
R20021 gnd.n2130 gnd.n2129 0.155672
R20022 gnd.n2114 gnd.n2086 0.155672
R20023 gnd.n2107 gnd.n2086 0.155672
R20024 gnd.n2107 gnd.n2106 0.155672
R20025 gnd.n2106 gnd.n2090 0.155672
R20026 gnd.n2099 gnd.n2090 0.155672
R20027 gnd.n2099 gnd.n2098 0.155672
R20028 gnd.n2082 gnd.n2054 0.155672
R20029 gnd.n2075 gnd.n2054 0.155672
R20030 gnd.n2075 gnd.n2074 0.155672
R20031 gnd.n2074 gnd.n2058 0.155672
R20032 gnd.n2067 gnd.n2058 0.155672
R20033 gnd.n2067 gnd.n2066 0.155672
R20034 gnd.n2050 gnd.n2022 0.155672
R20035 gnd.n2043 gnd.n2022 0.155672
R20036 gnd.n2043 gnd.n2042 0.155672
R20037 gnd.n2042 gnd.n2026 0.155672
R20038 gnd.n2035 gnd.n2026 0.155672
R20039 gnd.n2035 gnd.n2034 0.155672
R20040 gnd.n2018 gnd.n1990 0.155672
R20041 gnd.n2011 gnd.n1990 0.155672
R20042 gnd.n2011 gnd.n2010 0.155672
R20043 gnd.n2010 gnd.n1994 0.155672
R20044 gnd.n2003 gnd.n1994 0.155672
R20045 gnd.n2003 gnd.n2002 0.155672
R20046 gnd.n1987 gnd.n1959 0.155672
R20047 gnd.n1980 gnd.n1959 0.155672
R20048 gnd.n1980 gnd.n1979 0.155672
R20049 gnd.n1979 gnd.n1963 0.155672
R20050 gnd.n1972 gnd.n1963 0.155672
R20051 gnd.n1972 gnd.n1971 0.155672
R20052 gnd.n2334 gnd.n902 0.152939
R20053 gnd.n2334 gnd.n2333 0.152939
R20054 gnd.n2333 gnd.n2332 0.152939
R20055 gnd.n2332 gnd.n904 0.152939
R20056 gnd.n905 gnd.n904 0.152939
R20057 gnd.n906 gnd.n905 0.152939
R20058 gnd.n907 gnd.n906 0.152939
R20059 gnd.n908 gnd.n907 0.152939
R20060 gnd.n909 gnd.n908 0.152939
R20061 gnd.n910 gnd.n909 0.152939
R20062 gnd.n911 gnd.n910 0.152939
R20063 gnd.n912 gnd.n911 0.152939
R20064 gnd.n913 gnd.n912 0.152939
R20065 gnd.n914 gnd.n913 0.152939
R20066 gnd.n2304 gnd.n914 0.152939
R20067 gnd.n2304 gnd.n2303 0.152939
R20068 gnd.n1574 gnd.n1573 0.152939
R20069 gnd.n1574 gnd.n1278 0.152939
R20070 gnd.n1602 gnd.n1278 0.152939
R20071 gnd.n1603 gnd.n1602 0.152939
R20072 gnd.n1604 gnd.n1603 0.152939
R20073 gnd.n1605 gnd.n1604 0.152939
R20074 gnd.n1605 gnd.n1250 0.152939
R20075 gnd.n1632 gnd.n1250 0.152939
R20076 gnd.n1633 gnd.n1632 0.152939
R20077 gnd.n1634 gnd.n1633 0.152939
R20078 gnd.n1634 gnd.n1228 0.152939
R20079 gnd.n1663 gnd.n1228 0.152939
R20080 gnd.n1664 gnd.n1663 0.152939
R20081 gnd.n1665 gnd.n1664 0.152939
R20082 gnd.n1666 gnd.n1665 0.152939
R20083 gnd.n1668 gnd.n1666 0.152939
R20084 gnd.n1668 gnd.n1667 0.152939
R20085 gnd.n1667 gnd.n1177 0.152939
R20086 gnd.n1178 gnd.n1177 0.152939
R20087 gnd.n1179 gnd.n1178 0.152939
R20088 gnd.n1198 gnd.n1179 0.152939
R20089 gnd.n1199 gnd.n1198 0.152939
R20090 gnd.n1199 gnd.n1097 0.152939
R20091 gnd.n1758 gnd.n1097 0.152939
R20092 gnd.n1759 gnd.n1758 0.152939
R20093 gnd.n1760 gnd.n1759 0.152939
R20094 gnd.n1761 gnd.n1760 0.152939
R20095 gnd.n1761 gnd.n1070 0.152939
R20096 gnd.n1798 gnd.n1070 0.152939
R20097 gnd.n1799 gnd.n1798 0.152939
R20098 gnd.n1800 gnd.n1799 0.152939
R20099 gnd.n1801 gnd.n1800 0.152939
R20100 gnd.n1801 gnd.n1044 0.152939
R20101 gnd.n1845 gnd.n1044 0.152939
R20102 gnd.n1846 gnd.n1845 0.152939
R20103 gnd.n1847 gnd.n1846 0.152939
R20104 gnd.n1848 gnd.n1847 0.152939
R20105 gnd.n1848 gnd.n1017 0.152939
R20106 gnd.n1885 gnd.n1017 0.152939
R20107 gnd.n1886 gnd.n1885 0.152939
R20108 gnd.n1887 gnd.n1886 0.152939
R20109 gnd.n1888 gnd.n1887 0.152939
R20110 gnd.n1888 gnd.n990 0.152939
R20111 gnd.n1934 gnd.n990 0.152939
R20112 gnd.n1935 gnd.n1934 0.152939
R20113 gnd.n1936 gnd.n1935 0.152939
R20114 gnd.n1937 gnd.n1936 0.152939
R20115 gnd.n1937 gnd.n963 0.152939
R20116 gnd.n2228 gnd.n963 0.152939
R20117 gnd.n2229 gnd.n2228 0.152939
R20118 gnd.n2230 gnd.n2229 0.152939
R20119 gnd.n2231 gnd.n2230 0.152939
R20120 gnd.n2232 gnd.n2231 0.152939
R20121 gnd.n1572 gnd.n1302 0.152939
R20122 gnd.n1323 gnd.n1302 0.152939
R20123 gnd.n1324 gnd.n1323 0.152939
R20124 gnd.n1330 gnd.n1324 0.152939
R20125 gnd.n1331 gnd.n1330 0.152939
R20126 gnd.n1332 gnd.n1331 0.152939
R20127 gnd.n1332 gnd.n1321 0.152939
R20128 gnd.n1340 gnd.n1321 0.152939
R20129 gnd.n1341 gnd.n1340 0.152939
R20130 gnd.n1342 gnd.n1341 0.152939
R20131 gnd.n1342 gnd.n1319 0.152939
R20132 gnd.n1350 gnd.n1319 0.152939
R20133 gnd.n1351 gnd.n1350 0.152939
R20134 gnd.n1352 gnd.n1351 0.152939
R20135 gnd.n1352 gnd.n1317 0.152939
R20136 gnd.n1360 gnd.n1317 0.152939
R20137 gnd.n2301 gnd.n919 0.152939
R20138 gnd.n921 gnd.n919 0.152939
R20139 gnd.n922 gnd.n921 0.152939
R20140 gnd.n923 gnd.n922 0.152939
R20141 gnd.n924 gnd.n923 0.152939
R20142 gnd.n925 gnd.n924 0.152939
R20143 gnd.n926 gnd.n925 0.152939
R20144 gnd.n927 gnd.n926 0.152939
R20145 gnd.n928 gnd.n927 0.152939
R20146 gnd.n929 gnd.n928 0.152939
R20147 gnd.n930 gnd.n929 0.152939
R20148 gnd.n931 gnd.n930 0.152939
R20149 gnd.n932 gnd.n931 0.152939
R20150 gnd.n933 gnd.n932 0.152939
R20151 gnd.n934 gnd.n933 0.152939
R20152 gnd.n935 gnd.n934 0.152939
R20153 gnd.n936 gnd.n935 0.152939
R20154 gnd.n937 gnd.n936 0.152939
R20155 gnd.n938 gnd.n937 0.152939
R20156 gnd.n939 gnd.n938 0.152939
R20157 gnd.n940 gnd.n939 0.152939
R20158 gnd.n941 gnd.n940 0.152939
R20159 gnd.n945 gnd.n941 0.152939
R20160 gnd.n946 gnd.n945 0.152939
R20161 gnd.n947 gnd.n946 0.152939
R20162 gnd.n948 gnd.n947 0.152939
R20163 gnd.n1735 gnd.n1734 0.152939
R20164 gnd.n1736 gnd.n1735 0.152939
R20165 gnd.n1737 gnd.n1736 0.152939
R20166 gnd.n1738 gnd.n1737 0.152939
R20167 gnd.n1739 gnd.n1738 0.152939
R20168 gnd.n1740 gnd.n1739 0.152939
R20169 gnd.n1740 gnd.n1051 0.152939
R20170 gnd.n1819 gnd.n1051 0.152939
R20171 gnd.n1820 gnd.n1819 0.152939
R20172 gnd.n1821 gnd.n1820 0.152939
R20173 gnd.n1822 gnd.n1821 0.152939
R20174 gnd.n1823 gnd.n1822 0.152939
R20175 gnd.n1824 gnd.n1823 0.152939
R20176 gnd.n1825 gnd.n1824 0.152939
R20177 gnd.n1826 gnd.n1825 0.152939
R20178 gnd.n1827 gnd.n1826 0.152939
R20179 gnd.n1827 gnd.n997 0.152939
R20180 gnd.n1906 gnd.n997 0.152939
R20181 gnd.n1907 gnd.n1906 0.152939
R20182 gnd.n1908 gnd.n1907 0.152939
R20183 gnd.n1909 gnd.n1908 0.152939
R20184 gnd.n1910 gnd.n1909 0.152939
R20185 gnd.n1911 gnd.n1910 0.152939
R20186 gnd.n1912 gnd.n1911 0.152939
R20187 gnd.n1913 gnd.n1912 0.152939
R20188 gnd.n1914 gnd.n1913 0.152939
R20189 gnd.n1916 gnd.n1914 0.152939
R20190 gnd.n1916 gnd.n1915 0.152939
R20191 gnd.n1490 gnd.n1489 0.152939
R20192 gnd.n1490 gnd.n1380 0.152939
R20193 gnd.n1505 gnd.n1380 0.152939
R20194 gnd.n1506 gnd.n1505 0.152939
R20195 gnd.n1507 gnd.n1506 0.152939
R20196 gnd.n1507 gnd.n1368 0.152939
R20197 gnd.n1521 gnd.n1368 0.152939
R20198 gnd.n1522 gnd.n1521 0.152939
R20199 gnd.n1523 gnd.n1522 0.152939
R20200 gnd.n1524 gnd.n1523 0.152939
R20201 gnd.n1525 gnd.n1524 0.152939
R20202 gnd.n1526 gnd.n1525 0.152939
R20203 gnd.n1527 gnd.n1526 0.152939
R20204 gnd.n1528 gnd.n1527 0.152939
R20205 gnd.n1529 gnd.n1528 0.152939
R20206 gnd.n1530 gnd.n1529 0.152939
R20207 gnd.n1531 gnd.n1530 0.152939
R20208 gnd.n1532 gnd.n1531 0.152939
R20209 gnd.n1533 gnd.n1532 0.152939
R20210 gnd.n1534 gnd.n1533 0.152939
R20211 gnd.n1535 gnd.n1534 0.152939
R20212 gnd.n1535 gnd.n1234 0.152939
R20213 gnd.n1652 gnd.n1234 0.152939
R20214 gnd.n1653 gnd.n1652 0.152939
R20215 gnd.n1654 gnd.n1653 0.152939
R20216 gnd.n1655 gnd.n1654 0.152939
R20217 gnd.n1655 gnd.n1156 0.152939
R20218 gnd.n1732 gnd.n1156 0.152939
R20219 gnd.n1408 gnd.n1407 0.152939
R20220 gnd.n1409 gnd.n1408 0.152939
R20221 gnd.n1410 gnd.n1409 0.152939
R20222 gnd.n1411 gnd.n1410 0.152939
R20223 gnd.n1412 gnd.n1411 0.152939
R20224 gnd.n1413 gnd.n1412 0.152939
R20225 gnd.n1414 gnd.n1413 0.152939
R20226 gnd.n1415 gnd.n1414 0.152939
R20227 gnd.n1416 gnd.n1415 0.152939
R20228 gnd.n1417 gnd.n1416 0.152939
R20229 gnd.n1418 gnd.n1417 0.152939
R20230 gnd.n1419 gnd.n1418 0.152939
R20231 gnd.n1420 gnd.n1419 0.152939
R20232 gnd.n1421 gnd.n1420 0.152939
R20233 gnd.n1422 gnd.n1421 0.152939
R20234 gnd.n1423 gnd.n1422 0.152939
R20235 gnd.n1424 gnd.n1423 0.152939
R20236 gnd.n1425 gnd.n1424 0.152939
R20237 gnd.n1426 gnd.n1425 0.152939
R20238 gnd.n1427 gnd.n1426 0.152939
R20239 gnd.n1428 gnd.n1427 0.152939
R20240 gnd.n1429 gnd.n1428 0.152939
R20241 gnd.n1433 gnd.n1429 0.152939
R20242 gnd.n1434 gnd.n1433 0.152939
R20243 gnd.n1434 gnd.n1391 0.152939
R20244 gnd.n1488 gnd.n1391 0.152939
R20245 gnd.n6687 gnd.n702 0.152939
R20246 gnd.n6695 gnd.n702 0.152939
R20247 gnd.n6696 gnd.n6695 0.152939
R20248 gnd.n6697 gnd.n6696 0.152939
R20249 gnd.n6697 gnd.n696 0.152939
R20250 gnd.n6705 gnd.n696 0.152939
R20251 gnd.n6706 gnd.n6705 0.152939
R20252 gnd.n6707 gnd.n6706 0.152939
R20253 gnd.n6707 gnd.n690 0.152939
R20254 gnd.n6715 gnd.n690 0.152939
R20255 gnd.n6716 gnd.n6715 0.152939
R20256 gnd.n6717 gnd.n6716 0.152939
R20257 gnd.n6717 gnd.n684 0.152939
R20258 gnd.n6725 gnd.n684 0.152939
R20259 gnd.n6726 gnd.n6725 0.152939
R20260 gnd.n6727 gnd.n6726 0.152939
R20261 gnd.n6727 gnd.n678 0.152939
R20262 gnd.n6735 gnd.n678 0.152939
R20263 gnd.n6736 gnd.n6735 0.152939
R20264 gnd.n6737 gnd.n6736 0.152939
R20265 gnd.n6737 gnd.n672 0.152939
R20266 gnd.n6745 gnd.n672 0.152939
R20267 gnd.n6746 gnd.n6745 0.152939
R20268 gnd.n6747 gnd.n6746 0.152939
R20269 gnd.n6747 gnd.n666 0.152939
R20270 gnd.n6755 gnd.n666 0.152939
R20271 gnd.n6756 gnd.n6755 0.152939
R20272 gnd.n6757 gnd.n6756 0.152939
R20273 gnd.n6757 gnd.n660 0.152939
R20274 gnd.n6765 gnd.n660 0.152939
R20275 gnd.n6766 gnd.n6765 0.152939
R20276 gnd.n6767 gnd.n6766 0.152939
R20277 gnd.n6767 gnd.n654 0.152939
R20278 gnd.n6775 gnd.n654 0.152939
R20279 gnd.n6776 gnd.n6775 0.152939
R20280 gnd.n6777 gnd.n6776 0.152939
R20281 gnd.n6777 gnd.n648 0.152939
R20282 gnd.n6785 gnd.n648 0.152939
R20283 gnd.n6786 gnd.n6785 0.152939
R20284 gnd.n6787 gnd.n6786 0.152939
R20285 gnd.n6787 gnd.n642 0.152939
R20286 gnd.n6795 gnd.n642 0.152939
R20287 gnd.n6796 gnd.n6795 0.152939
R20288 gnd.n6797 gnd.n6796 0.152939
R20289 gnd.n6797 gnd.n636 0.152939
R20290 gnd.n6805 gnd.n636 0.152939
R20291 gnd.n6806 gnd.n6805 0.152939
R20292 gnd.n6807 gnd.n6806 0.152939
R20293 gnd.n6807 gnd.n630 0.152939
R20294 gnd.n6815 gnd.n630 0.152939
R20295 gnd.n6816 gnd.n6815 0.152939
R20296 gnd.n6817 gnd.n6816 0.152939
R20297 gnd.n6817 gnd.n624 0.152939
R20298 gnd.n6825 gnd.n624 0.152939
R20299 gnd.n6826 gnd.n6825 0.152939
R20300 gnd.n6827 gnd.n6826 0.152939
R20301 gnd.n6827 gnd.n618 0.152939
R20302 gnd.n6835 gnd.n618 0.152939
R20303 gnd.n6836 gnd.n6835 0.152939
R20304 gnd.n6837 gnd.n6836 0.152939
R20305 gnd.n6837 gnd.n612 0.152939
R20306 gnd.n6845 gnd.n612 0.152939
R20307 gnd.n6846 gnd.n6845 0.152939
R20308 gnd.n6847 gnd.n6846 0.152939
R20309 gnd.n6847 gnd.n606 0.152939
R20310 gnd.n6855 gnd.n606 0.152939
R20311 gnd.n6856 gnd.n6855 0.152939
R20312 gnd.n6857 gnd.n6856 0.152939
R20313 gnd.n6857 gnd.n600 0.152939
R20314 gnd.n6865 gnd.n600 0.152939
R20315 gnd.n6866 gnd.n6865 0.152939
R20316 gnd.n6867 gnd.n6866 0.152939
R20317 gnd.n6867 gnd.n594 0.152939
R20318 gnd.n6875 gnd.n594 0.152939
R20319 gnd.n6876 gnd.n6875 0.152939
R20320 gnd.n6877 gnd.n6876 0.152939
R20321 gnd.n6877 gnd.n588 0.152939
R20322 gnd.n6885 gnd.n588 0.152939
R20323 gnd.n6886 gnd.n6885 0.152939
R20324 gnd.n6887 gnd.n6886 0.152939
R20325 gnd.n6887 gnd.n582 0.152939
R20326 gnd.n6895 gnd.n582 0.152939
R20327 gnd.n6896 gnd.n6895 0.152939
R20328 gnd.n6897 gnd.n6896 0.152939
R20329 gnd.n6897 gnd.n576 0.152939
R20330 gnd.n6905 gnd.n576 0.152939
R20331 gnd.n6906 gnd.n6905 0.152939
R20332 gnd.n6907 gnd.n6906 0.152939
R20333 gnd.n6907 gnd.n570 0.152939
R20334 gnd.n6915 gnd.n570 0.152939
R20335 gnd.n6916 gnd.n6915 0.152939
R20336 gnd.n6917 gnd.n6916 0.152939
R20337 gnd.n6917 gnd.n564 0.152939
R20338 gnd.n6925 gnd.n564 0.152939
R20339 gnd.n6926 gnd.n6925 0.152939
R20340 gnd.n6927 gnd.n6926 0.152939
R20341 gnd.n6927 gnd.n558 0.152939
R20342 gnd.n6935 gnd.n558 0.152939
R20343 gnd.n6936 gnd.n6935 0.152939
R20344 gnd.n6937 gnd.n6936 0.152939
R20345 gnd.n6937 gnd.n552 0.152939
R20346 gnd.n6945 gnd.n552 0.152939
R20347 gnd.n6946 gnd.n6945 0.152939
R20348 gnd.n6947 gnd.n6946 0.152939
R20349 gnd.n6947 gnd.n546 0.152939
R20350 gnd.n6955 gnd.n546 0.152939
R20351 gnd.n6956 gnd.n6955 0.152939
R20352 gnd.n6957 gnd.n6956 0.152939
R20353 gnd.n6957 gnd.n540 0.152939
R20354 gnd.n6965 gnd.n540 0.152939
R20355 gnd.n6966 gnd.n6965 0.152939
R20356 gnd.n6967 gnd.n6966 0.152939
R20357 gnd.n6967 gnd.n534 0.152939
R20358 gnd.n6975 gnd.n534 0.152939
R20359 gnd.n6976 gnd.n6975 0.152939
R20360 gnd.n6977 gnd.n6976 0.152939
R20361 gnd.n6977 gnd.n528 0.152939
R20362 gnd.n6985 gnd.n528 0.152939
R20363 gnd.n6986 gnd.n6985 0.152939
R20364 gnd.n6987 gnd.n6986 0.152939
R20365 gnd.n6987 gnd.n522 0.152939
R20366 gnd.n6995 gnd.n522 0.152939
R20367 gnd.n6996 gnd.n6995 0.152939
R20368 gnd.n6997 gnd.n6996 0.152939
R20369 gnd.n6997 gnd.n516 0.152939
R20370 gnd.n7005 gnd.n516 0.152939
R20371 gnd.n7006 gnd.n7005 0.152939
R20372 gnd.n7007 gnd.n7006 0.152939
R20373 gnd.n7007 gnd.n510 0.152939
R20374 gnd.n7015 gnd.n510 0.152939
R20375 gnd.n7016 gnd.n7015 0.152939
R20376 gnd.n7017 gnd.n7016 0.152939
R20377 gnd.n7017 gnd.n504 0.152939
R20378 gnd.n7025 gnd.n504 0.152939
R20379 gnd.n7026 gnd.n7025 0.152939
R20380 gnd.n7027 gnd.n7026 0.152939
R20381 gnd.n7027 gnd.n498 0.152939
R20382 gnd.n7035 gnd.n498 0.152939
R20383 gnd.n7036 gnd.n7035 0.152939
R20384 gnd.n7037 gnd.n7036 0.152939
R20385 gnd.n7037 gnd.n492 0.152939
R20386 gnd.n7045 gnd.n492 0.152939
R20387 gnd.n7046 gnd.n7045 0.152939
R20388 gnd.n7047 gnd.n7046 0.152939
R20389 gnd.n7047 gnd.n486 0.152939
R20390 gnd.n7055 gnd.n486 0.152939
R20391 gnd.n7056 gnd.n7055 0.152939
R20392 gnd.n7057 gnd.n7056 0.152939
R20393 gnd.n7057 gnd.n480 0.152939
R20394 gnd.n7065 gnd.n480 0.152939
R20395 gnd.n7066 gnd.n7065 0.152939
R20396 gnd.n7067 gnd.n7066 0.152939
R20397 gnd.n7067 gnd.n474 0.152939
R20398 gnd.n7075 gnd.n474 0.152939
R20399 gnd.n7076 gnd.n7075 0.152939
R20400 gnd.n7077 gnd.n7076 0.152939
R20401 gnd.n7077 gnd.n468 0.152939
R20402 gnd.n7085 gnd.n468 0.152939
R20403 gnd.n7086 gnd.n7085 0.152939
R20404 gnd.n7087 gnd.n7086 0.152939
R20405 gnd.n7087 gnd.n462 0.152939
R20406 gnd.n7095 gnd.n462 0.152939
R20407 gnd.n7096 gnd.n7095 0.152939
R20408 gnd.n7097 gnd.n7096 0.152939
R20409 gnd.n7097 gnd.n456 0.152939
R20410 gnd.n7105 gnd.n456 0.152939
R20411 gnd.n7106 gnd.n7105 0.152939
R20412 gnd.n7107 gnd.n7106 0.152939
R20413 gnd.n7107 gnd.n450 0.152939
R20414 gnd.n7115 gnd.n450 0.152939
R20415 gnd.n7116 gnd.n7115 0.152939
R20416 gnd.n7117 gnd.n7116 0.152939
R20417 gnd.n7117 gnd.n444 0.152939
R20418 gnd.n7125 gnd.n444 0.152939
R20419 gnd.n7126 gnd.n7125 0.152939
R20420 gnd.n7127 gnd.n7126 0.152939
R20421 gnd.n7127 gnd.n438 0.152939
R20422 gnd.n7135 gnd.n438 0.152939
R20423 gnd.n7136 gnd.n7135 0.152939
R20424 gnd.n7137 gnd.n7136 0.152939
R20425 gnd.n7137 gnd.n432 0.152939
R20426 gnd.n7145 gnd.n432 0.152939
R20427 gnd.n7146 gnd.n7145 0.152939
R20428 gnd.n7147 gnd.n7146 0.152939
R20429 gnd.n7147 gnd.n426 0.152939
R20430 gnd.n7155 gnd.n426 0.152939
R20431 gnd.n7156 gnd.n7155 0.152939
R20432 gnd.n7157 gnd.n7156 0.152939
R20433 gnd.n7157 gnd.n420 0.152939
R20434 gnd.n7165 gnd.n420 0.152939
R20435 gnd.n7166 gnd.n7165 0.152939
R20436 gnd.n7167 gnd.n7166 0.152939
R20437 gnd.n7167 gnd.n414 0.152939
R20438 gnd.n7175 gnd.n414 0.152939
R20439 gnd.n7176 gnd.n7175 0.152939
R20440 gnd.n7177 gnd.n7176 0.152939
R20441 gnd.n7177 gnd.n408 0.152939
R20442 gnd.n7185 gnd.n408 0.152939
R20443 gnd.n7186 gnd.n7185 0.152939
R20444 gnd.n7187 gnd.n7186 0.152939
R20445 gnd.n7187 gnd.n402 0.152939
R20446 gnd.n7195 gnd.n402 0.152939
R20447 gnd.n7196 gnd.n7195 0.152939
R20448 gnd.n7198 gnd.n7196 0.152939
R20449 gnd.n7198 gnd.n7197 0.152939
R20450 gnd.n7197 gnd.n396 0.152939
R20451 gnd.n7207 gnd.n396 0.152939
R20452 gnd.n7208 gnd.n391 0.152939
R20453 gnd.n7216 gnd.n391 0.152939
R20454 gnd.n7217 gnd.n7216 0.152939
R20455 gnd.n7218 gnd.n7217 0.152939
R20456 gnd.n7218 gnd.n385 0.152939
R20457 gnd.n7226 gnd.n385 0.152939
R20458 gnd.n7227 gnd.n7226 0.152939
R20459 gnd.n7228 gnd.n7227 0.152939
R20460 gnd.n7228 gnd.n379 0.152939
R20461 gnd.n7236 gnd.n379 0.152939
R20462 gnd.n7237 gnd.n7236 0.152939
R20463 gnd.n7238 gnd.n7237 0.152939
R20464 gnd.n7238 gnd.n373 0.152939
R20465 gnd.n7246 gnd.n373 0.152939
R20466 gnd.n7247 gnd.n7246 0.152939
R20467 gnd.n7248 gnd.n7247 0.152939
R20468 gnd.n7248 gnd.n367 0.152939
R20469 gnd.n7256 gnd.n367 0.152939
R20470 gnd.n7257 gnd.n7256 0.152939
R20471 gnd.n7258 gnd.n7257 0.152939
R20472 gnd.n7258 gnd.n361 0.152939
R20473 gnd.n7266 gnd.n361 0.152939
R20474 gnd.n7267 gnd.n7266 0.152939
R20475 gnd.n7268 gnd.n7267 0.152939
R20476 gnd.n7268 gnd.n355 0.152939
R20477 gnd.n7276 gnd.n355 0.152939
R20478 gnd.n7277 gnd.n7276 0.152939
R20479 gnd.n7278 gnd.n7277 0.152939
R20480 gnd.n7278 gnd.n349 0.152939
R20481 gnd.n7286 gnd.n349 0.152939
R20482 gnd.n7287 gnd.n7286 0.152939
R20483 gnd.n7288 gnd.n7287 0.152939
R20484 gnd.n7288 gnd.n343 0.152939
R20485 gnd.n7296 gnd.n343 0.152939
R20486 gnd.n7297 gnd.n7296 0.152939
R20487 gnd.n7298 gnd.n7297 0.152939
R20488 gnd.n7298 gnd.n337 0.152939
R20489 gnd.n7306 gnd.n337 0.152939
R20490 gnd.n7307 gnd.n7306 0.152939
R20491 gnd.n7308 gnd.n7307 0.152939
R20492 gnd.n7308 gnd.n331 0.152939
R20493 gnd.n7316 gnd.n331 0.152939
R20494 gnd.n7317 gnd.n7316 0.152939
R20495 gnd.n7318 gnd.n7317 0.152939
R20496 gnd.n7318 gnd.n325 0.152939
R20497 gnd.n7326 gnd.n325 0.152939
R20498 gnd.n7327 gnd.n7326 0.152939
R20499 gnd.n7328 gnd.n7327 0.152939
R20500 gnd.n7328 gnd.n319 0.152939
R20501 gnd.n7336 gnd.n319 0.152939
R20502 gnd.n7337 gnd.n7336 0.152939
R20503 gnd.n7338 gnd.n7337 0.152939
R20504 gnd.n7338 gnd.n313 0.152939
R20505 gnd.n7346 gnd.n313 0.152939
R20506 gnd.n7347 gnd.n7346 0.152939
R20507 gnd.n7348 gnd.n7347 0.152939
R20508 gnd.n7348 gnd.n307 0.152939
R20509 gnd.n7356 gnd.n307 0.152939
R20510 gnd.n7357 gnd.n7356 0.152939
R20511 gnd.n7358 gnd.n7357 0.152939
R20512 gnd.n7358 gnd.n301 0.152939
R20513 gnd.n7366 gnd.n301 0.152939
R20514 gnd.n7367 gnd.n7366 0.152939
R20515 gnd.n7368 gnd.n7367 0.152939
R20516 gnd.n7368 gnd.n295 0.152939
R20517 gnd.n7376 gnd.n295 0.152939
R20518 gnd.n7377 gnd.n7376 0.152939
R20519 gnd.n7378 gnd.n7377 0.152939
R20520 gnd.n7378 gnd.n289 0.152939
R20521 gnd.n7386 gnd.n289 0.152939
R20522 gnd.n7387 gnd.n7386 0.152939
R20523 gnd.n7388 gnd.n7387 0.152939
R20524 gnd.n7388 gnd.n283 0.152939
R20525 gnd.n7396 gnd.n283 0.152939
R20526 gnd.n7397 gnd.n7396 0.152939
R20527 gnd.n7398 gnd.n7397 0.152939
R20528 gnd.n7398 gnd.n277 0.152939
R20529 gnd.n7406 gnd.n277 0.152939
R20530 gnd.n7407 gnd.n7406 0.152939
R20531 gnd.n7408 gnd.n7407 0.152939
R20532 gnd.n7408 gnd.n271 0.152939
R20533 gnd.n7416 gnd.n271 0.152939
R20534 gnd.n7417 gnd.n7416 0.152939
R20535 gnd.n7419 gnd.n7417 0.152939
R20536 gnd.n3186 gnd.n3183 0.152939
R20537 gnd.n3187 gnd.n3186 0.152939
R20538 gnd.n3188 gnd.n3187 0.152939
R20539 gnd.n3189 gnd.n3188 0.152939
R20540 gnd.n3192 gnd.n3189 0.152939
R20541 gnd.n3193 gnd.n3192 0.152939
R20542 gnd.n3194 gnd.n3193 0.152939
R20543 gnd.n3195 gnd.n3194 0.152939
R20544 gnd.n3198 gnd.n3195 0.152939
R20545 gnd.n3199 gnd.n3198 0.152939
R20546 gnd.n3200 gnd.n3199 0.152939
R20547 gnd.n3201 gnd.n3200 0.152939
R20548 gnd.n3204 gnd.n3201 0.152939
R20549 gnd.n3205 gnd.n3204 0.152939
R20550 gnd.n3206 gnd.n3205 0.152939
R20551 gnd.n3208 gnd.n3206 0.152939
R20552 gnd.n3208 gnd.n3207 0.152939
R20553 gnd.n3207 gnd.n247 0.152939
R20554 gnd.n248 gnd.n247 0.152939
R20555 gnd.n249 gnd.n248 0.152939
R20556 gnd.n254 gnd.n249 0.152939
R20557 gnd.n255 gnd.n254 0.152939
R20558 gnd.n256 gnd.n255 0.152939
R20559 gnd.n257 gnd.n256 0.152939
R20560 gnd.n262 gnd.n257 0.152939
R20561 gnd.n263 gnd.n262 0.152939
R20562 gnd.n264 gnd.n263 0.152939
R20563 gnd.n265 gnd.n264 0.152939
R20564 gnd.n7418 gnd.n265 0.152939
R20565 gnd.n7726 gnd.n77 0.152939
R20566 gnd.n103 gnd.n77 0.152939
R20567 gnd.n104 gnd.n103 0.152939
R20568 gnd.n105 gnd.n104 0.152939
R20569 gnd.n122 gnd.n105 0.152939
R20570 gnd.n123 gnd.n122 0.152939
R20571 gnd.n124 gnd.n123 0.152939
R20572 gnd.n125 gnd.n124 0.152939
R20573 gnd.n143 gnd.n125 0.152939
R20574 gnd.n144 gnd.n143 0.152939
R20575 gnd.n145 gnd.n144 0.152939
R20576 gnd.n146 gnd.n145 0.152939
R20577 gnd.n163 gnd.n146 0.152939
R20578 gnd.n164 gnd.n163 0.152939
R20579 gnd.n165 gnd.n164 0.152939
R20580 gnd.n166 gnd.n165 0.152939
R20581 gnd.n7735 gnd.n65 0.152939
R20582 gnd.n5851 gnd.n65 0.152939
R20583 gnd.n5852 gnd.n5851 0.152939
R20584 gnd.n5852 gnd.n3236 0.152939
R20585 gnd.n5864 gnd.n3236 0.152939
R20586 gnd.n5865 gnd.n5864 0.152939
R20587 gnd.n5867 gnd.n5865 0.152939
R20588 gnd.n5867 gnd.n5866 0.152939
R20589 gnd.n5866 gnd.n3229 0.152939
R20590 gnd.n3230 gnd.n3229 0.152939
R20591 gnd.n3231 gnd.n3230 0.152939
R20592 gnd.n5878 gnd.n3231 0.152939
R20593 gnd.n5879 gnd.n5878 0.152939
R20594 gnd.n5880 gnd.n5879 0.152939
R20595 gnd.n5881 gnd.n5880 0.152939
R20596 gnd.n5884 gnd.n5881 0.152939
R20597 gnd.n5886 gnd.n5884 0.152939
R20598 gnd.n5886 gnd.n5885 0.152939
R20599 gnd.n5885 gnd.n178 0.152939
R20600 gnd.n7664 gnd.n178 0.152939
R20601 gnd.n201 gnd.n200 0.152939
R20602 gnd.n208 gnd.n200 0.152939
R20603 gnd.n209 gnd.n208 0.152939
R20604 gnd.n210 gnd.n209 0.152939
R20605 gnd.n210 gnd.n198 0.152939
R20606 gnd.n218 gnd.n198 0.152939
R20607 gnd.n219 gnd.n218 0.152939
R20608 gnd.n220 gnd.n219 0.152939
R20609 gnd.n220 gnd.n196 0.152939
R20610 gnd.n228 gnd.n196 0.152939
R20611 gnd.n229 gnd.n228 0.152939
R20612 gnd.n230 gnd.n229 0.152939
R20613 gnd.n230 gnd.n194 0.152939
R20614 gnd.n237 gnd.n194 0.152939
R20615 gnd.n238 gnd.n237 0.152939
R20616 gnd.n239 gnd.n238 0.152939
R20617 gnd.n239 gnd.n179 0.152939
R20618 gnd.n7663 gnd.n179 0.152939
R20619 gnd.n7480 gnd.n7479 0.152939
R20620 gnd.n7481 gnd.n7480 0.152939
R20621 gnd.n7482 gnd.n7481 0.152939
R20622 gnd.n7483 gnd.n7482 0.152939
R20623 gnd.n7484 gnd.n7483 0.152939
R20624 gnd.n7485 gnd.n7484 0.152939
R20625 gnd.n7486 gnd.n7485 0.152939
R20626 gnd.n7487 gnd.n7486 0.152939
R20627 gnd.n7488 gnd.n7487 0.152939
R20628 gnd.n7489 gnd.n7488 0.152939
R20629 gnd.n7490 gnd.n7489 0.152939
R20630 gnd.n7491 gnd.n7490 0.152939
R20631 gnd.n7492 gnd.n7491 0.152939
R20632 gnd.n7493 gnd.n7492 0.152939
R20633 gnd.n7494 gnd.n7493 0.152939
R20634 gnd.n7495 gnd.n7494 0.152939
R20635 gnd.n7496 gnd.n7495 0.152939
R20636 gnd.n7497 gnd.n7496 0.152939
R20637 gnd.n7498 gnd.n7497 0.152939
R20638 gnd.n7499 gnd.n7498 0.152939
R20639 gnd.n7500 gnd.n7499 0.152939
R20640 gnd.n7501 gnd.n7500 0.152939
R20641 gnd.n7502 gnd.n7501 0.152939
R20642 gnd.n7503 gnd.n7502 0.152939
R20643 gnd.n7504 gnd.n7503 0.152939
R20644 gnd.n7505 gnd.n7504 0.152939
R20645 gnd.n7506 gnd.n7505 0.152939
R20646 gnd.n7507 gnd.n7506 0.152939
R20647 gnd.n7508 gnd.n7507 0.152939
R20648 gnd.n7509 gnd.n7508 0.152939
R20649 gnd.n7510 gnd.n7509 0.152939
R20650 gnd.n7511 gnd.n7510 0.152939
R20651 gnd.n7512 gnd.n7511 0.152939
R20652 gnd.n7513 gnd.n7512 0.152939
R20653 gnd.n7514 gnd.n7513 0.152939
R20654 gnd.n7515 gnd.n7514 0.152939
R20655 gnd.n7583 gnd.n7515 0.152939
R20656 gnd.n7583 gnd.n7582 0.152939
R20657 gnd.n7582 gnd.n7581 0.152939
R20658 gnd.n7581 gnd.n7519 0.152939
R20659 gnd.n7520 gnd.n7519 0.152939
R20660 gnd.n7521 gnd.n7520 0.152939
R20661 gnd.n7522 gnd.n7521 0.152939
R20662 gnd.n7523 gnd.n7522 0.152939
R20663 gnd.n7524 gnd.n7523 0.152939
R20664 gnd.n7525 gnd.n7524 0.152939
R20665 gnd.n7526 gnd.n7525 0.152939
R20666 gnd.n7527 gnd.n7526 0.152939
R20667 gnd.n7528 gnd.n7527 0.152939
R20668 gnd.n7529 gnd.n7528 0.152939
R20669 gnd.n7530 gnd.n7529 0.152939
R20670 gnd.n7531 gnd.n7530 0.152939
R20671 gnd.n7532 gnd.n7531 0.152939
R20672 gnd.n7533 gnd.n7532 0.152939
R20673 gnd.n7534 gnd.n7533 0.152939
R20674 gnd.n7535 gnd.n7534 0.152939
R20675 gnd.n7541 gnd.n7535 0.152939
R20676 gnd.n7541 gnd.n7540 0.152939
R20677 gnd.n5573 gnd.n5572 0.152939
R20678 gnd.n5573 gnd.n5569 0.152939
R20679 gnd.n5581 gnd.n5569 0.152939
R20680 gnd.n5582 gnd.n5581 0.152939
R20681 gnd.n5583 gnd.n5582 0.152939
R20682 gnd.n5583 gnd.n5565 0.152939
R20683 gnd.n5591 gnd.n5565 0.152939
R20684 gnd.n5592 gnd.n5591 0.152939
R20685 gnd.n5593 gnd.n5592 0.152939
R20686 gnd.n5593 gnd.n5561 0.152939
R20687 gnd.n5601 gnd.n5561 0.152939
R20688 gnd.n5602 gnd.n5601 0.152939
R20689 gnd.n5603 gnd.n5602 0.152939
R20690 gnd.n5603 gnd.n5557 0.152939
R20691 gnd.n5611 gnd.n5557 0.152939
R20692 gnd.n5612 gnd.n5611 0.152939
R20693 gnd.n5613 gnd.n5612 0.152939
R20694 gnd.n5613 gnd.n5553 0.152939
R20695 gnd.n5624 gnd.n5553 0.152939
R20696 gnd.n5625 gnd.n5624 0.152939
R20697 gnd.n5626 gnd.n5625 0.152939
R20698 gnd.n5626 gnd.n5549 0.152939
R20699 gnd.n5634 gnd.n5549 0.152939
R20700 gnd.n5635 gnd.n5634 0.152939
R20701 gnd.n5637 gnd.n5635 0.152939
R20702 gnd.n5647 gnd.n3297 0.152939
R20703 gnd.n5648 gnd.n5647 0.152939
R20704 gnd.n5649 gnd.n5648 0.152939
R20705 gnd.n5649 gnd.n3293 0.152939
R20706 gnd.n5657 gnd.n3293 0.152939
R20707 gnd.n5658 gnd.n5657 0.152939
R20708 gnd.n5659 gnd.n5658 0.152939
R20709 gnd.n5659 gnd.n3289 0.152939
R20710 gnd.n5669 gnd.n3289 0.152939
R20711 gnd.n5670 gnd.n5669 0.152939
R20712 gnd.n5671 gnd.n5670 0.152939
R20713 gnd.n5671 gnd.n3285 0.152939
R20714 gnd.n5679 gnd.n3285 0.152939
R20715 gnd.n5680 gnd.n5679 0.152939
R20716 gnd.n5681 gnd.n5680 0.152939
R20717 gnd.n5681 gnd.n3281 0.152939
R20718 gnd.n5689 gnd.n3281 0.152939
R20719 gnd.n5690 gnd.n5689 0.152939
R20720 gnd.n5691 gnd.n5690 0.152939
R20721 gnd.n5691 gnd.n3277 0.152939
R20722 gnd.n5699 gnd.n3277 0.152939
R20723 gnd.n5700 gnd.n5699 0.152939
R20724 gnd.n5701 gnd.n5700 0.152939
R20725 gnd.n5701 gnd.n3273 0.152939
R20726 gnd.n5709 gnd.n3273 0.152939
R20727 gnd.n5710 gnd.n5709 0.152939
R20728 gnd.n5712 gnd.n5710 0.152939
R20729 gnd.n5712 gnd.n5711 0.152939
R20730 gnd.n5711 gnd.n3266 0.152939
R20731 gnd.n5721 gnd.n3266 0.152939
R20732 gnd.n3064 gnd.n3063 0.152939
R20733 gnd.n3065 gnd.n3064 0.152939
R20734 gnd.n3085 gnd.n3065 0.152939
R20735 gnd.n3086 gnd.n3085 0.152939
R20736 gnd.n3087 gnd.n3086 0.152939
R20737 gnd.n3088 gnd.n3087 0.152939
R20738 gnd.n3105 gnd.n3088 0.152939
R20739 gnd.n3106 gnd.n3105 0.152939
R20740 gnd.n3107 gnd.n3106 0.152939
R20741 gnd.n3108 gnd.n3107 0.152939
R20742 gnd.n3125 gnd.n3108 0.152939
R20743 gnd.n3126 gnd.n3125 0.152939
R20744 gnd.n3127 gnd.n3126 0.152939
R20745 gnd.n3128 gnd.n3127 0.152939
R20746 gnd.n3128 gnd.n78 0.152939
R20747 gnd.n7726 gnd.n78 0.152939
R20748 gnd.n4367 gnd.n4366 0.152939
R20749 gnd.n4368 gnd.n4367 0.152939
R20750 gnd.n4369 gnd.n4368 0.152939
R20751 gnd.n4372 gnd.n4369 0.152939
R20752 gnd.n4373 gnd.n4372 0.152939
R20753 gnd.n4374 gnd.n4373 0.152939
R20754 gnd.n4375 gnd.n4374 0.152939
R20755 gnd.n4376 gnd.n4375 0.152939
R20756 gnd.n4376 gnd.n3854 0.152939
R20757 gnd.n4441 gnd.n3854 0.152939
R20758 gnd.n4442 gnd.n4441 0.152939
R20759 gnd.n4443 gnd.n4442 0.152939
R20760 gnd.n4443 gnd.n3850 0.152939
R20761 gnd.n4449 gnd.n3850 0.152939
R20762 gnd.n4450 gnd.n4449 0.152939
R20763 gnd.n4451 gnd.n4450 0.152939
R20764 gnd.n4451 gnd.n3846 0.152939
R20765 gnd.n4457 gnd.n3846 0.152939
R20766 gnd.n4458 gnd.n4457 0.152939
R20767 gnd.n4459 gnd.n4458 0.152939
R20768 gnd.n4459 gnd.n3841 0.152939
R20769 gnd.n4467 gnd.n3841 0.152939
R20770 gnd.n4468 gnd.n4467 0.152939
R20771 gnd.n4469 gnd.n4468 0.152939
R20772 gnd.n4471 gnd.n4469 0.152939
R20773 gnd.n4471 gnd.n4470 0.152939
R20774 gnd.n4470 gnd.n2917 0.152939
R20775 gnd.n2918 gnd.n2917 0.152939
R20776 gnd.n2919 gnd.n2918 0.152939
R20777 gnd.n2934 gnd.n2919 0.152939
R20778 gnd.n2935 gnd.n2934 0.152939
R20779 gnd.n2936 gnd.n2935 0.152939
R20780 gnd.n2937 gnd.n2936 0.152939
R20781 gnd.n4556 gnd.n2937 0.152939
R20782 gnd.n4557 gnd.n4556 0.152939
R20783 gnd.n4557 gnd.n3710 0.152939
R20784 gnd.n4591 gnd.n3710 0.152939
R20785 gnd.n4592 gnd.n4591 0.152939
R20786 gnd.n4593 gnd.n4592 0.152939
R20787 gnd.n4593 gnd.n3685 0.152939
R20788 gnd.n4634 gnd.n3685 0.152939
R20789 gnd.n4635 gnd.n4634 0.152939
R20790 gnd.n4636 gnd.n4635 0.152939
R20791 gnd.n4636 gnd.n3670 0.152939
R20792 gnd.n4679 gnd.n3670 0.152939
R20793 gnd.n4680 gnd.n4679 0.152939
R20794 gnd.n4681 gnd.n4680 0.152939
R20795 gnd.n4682 gnd.n4681 0.152939
R20796 gnd.n4682 gnd.n3642 0.152939
R20797 gnd.n4752 gnd.n3642 0.152939
R20798 gnd.n4753 gnd.n4752 0.152939
R20799 gnd.n4754 gnd.n4753 0.152939
R20800 gnd.n4754 gnd.n3622 0.152939
R20801 gnd.n4780 gnd.n3622 0.152939
R20802 gnd.n4781 gnd.n4780 0.152939
R20803 gnd.n4782 gnd.n4781 0.152939
R20804 gnd.n4782 gnd.n3601 0.152939
R20805 gnd.n4813 gnd.n3601 0.152939
R20806 gnd.n4814 gnd.n4813 0.152939
R20807 gnd.n4815 gnd.n4814 0.152939
R20808 gnd.n4815 gnd.n3584 0.152939
R20809 gnd.n4857 gnd.n3584 0.152939
R20810 gnd.n4858 gnd.n4857 0.152939
R20811 gnd.n4859 gnd.n4858 0.152939
R20812 gnd.n4860 gnd.n4859 0.152939
R20813 gnd.n4860 gnd.n3555 0.152939
R20814 gnd.n4907 gnd.n3555 0.152939
R20815 gnd.n4908 gnd.n4907 0.152939
R20816 gnd.n4909 gnd.n4908 0.152939
R20817 gnd.n4909 gnd.n3536 0.152939
R20818 gnd.n4935 gnd.n3536 0.152939
R20819 gnd.n4936 gnd.n4935 0.152939
R20820 gnd.n4937 gnd.n4936 0.152939
R20821 gnd.n4938 gnd.n4937 0.152939
R20822 gnd.n4939 gnd.n4938 0.152939
R20823 gnd.n4939 gnd.n3505 0.152939
R20824 gnd.n5010 gnd.n3505 0.152939
R20825 gnd.n5011 gnd.n5010 0.152939
R20826 gnd.n5012 gnd.n5011 0.152939
R20827 gnd.n5013 gnd.n5012 0.152939
R20828 gnd.n5013 gnd.n3477 0.152939
R20829 gnd.n5062 gnd.n3477 0.152939
R20830 gnd.n5063 gnd.n5062 0.152939
R20831 gnd.n5064 gnd.n5063 0.152939
R20832 gnd.n5065 gnd.n5064 0.152939
R20833 gnd.n5065 gnd.n3460 0.152939
R20834 gnd.n5090 gnd.n3460 0.152939
R20835 gnd.n5091 gnd.n5090 0.152939
R20836 gnd.n5092 gnd.n5091 0.152939
R20837 gnd.n5092 gnd.n3402 0.152939
R20838 gnd.n5133 gnd.n3402 0.152939
R20839 gnd.n5134 gnd.n5133 0.152939
R20840 gnd.n5135 gnd.n5134 0.152939
R20841 gnd.n5135 gnd.n3380 0.152939
R20842 gnd.n5161 gnd.n3380 0.152939
R20843 gnd.n5162 gnd.n5161 0.152939
R20844 gnd.n5163 gnd.n5162 0.152939
R20845 gnd.n5165 gnd.n5163 0.152939
R20846 gnd.n5165 gnd.n5164 0.152939
R20847 gnd.n5164 gnd.n3351 0.152939
R20848 gnd.n3352 gnd.n3351 0.152939
R20849 gnd.n3353 gnd.n3352 0.152939
R20850 gnd.n3355 gnd.n3353 0.152939
R20851 gnd.n3355 gnd.n3354 0.152939
R20852 gnd.n3354 gnd.n3042 0.152939
R20853 gnd.n3043 gnd.n3042 0.152939
R20854 gnd.n3044 gnd.n3043 0.152939
R20855 gnd.n3050 gnd.n3044 0.152939
R20856 gnd.n3051 gnd.n3050 0.152939
R20857 gnd.n3052 gnd.n3051 0.152939
R20858 gnd.n3053 gnd.n3052 0.152939
R20859 gnd.n5766 gnd.n3053 0.152939
R20860 gnd.n5769 gnd.n5766 0.152939
R20861 gnd.n5770 gnd.n5769 0.152939
R20862 gnd.n5771 gnd.n5770 0.152939
R20863 gnd.n5771 gnd.n5762 0.152939
R20864 gnd.n5777 gnd.n5762 0.152939
R20865 gnd.n5778 gnd.n5777 0.152939
R20866 gnd.n5779 gnd.n5778 0.152939
R20867 gnd.n5779 gnd.n3251 0.152939
R20868 gnd.n5785 gnd.n3251 0.152939
R20869 gnd.n5786 gnd.n5785 0.152939
R20870 gnd.n5787 gnd.n5786 0.152939
R20871 gnd.n5788 gnd.n5787 0.152939
R20872 gnd.n5789 gnd.n5788 0.152939
R20873 gnd.n5791 gnd.n5789 0.152939
R20874 gnd.n5792 gnd.n5791 0.152939
R20875 gnd.n3958 gnd.n3926 0.152939
R20876 gnd.n3927 gnd.n3926 0.152939
R20877 gnd.n3928 gnd.n3927 0.152939
R20878 gnd.n4220 gnd.n3928 0.152939
R20879 gnd.n4221 gnd.n4220 0.152939
R20880 gnd.n4222 gnd.n4221 0.152939
R20881 gnd.n4223 gnd.n4222 0.152939
R20882 gnd.n4228 gnd.n4223 0.152939
R20883 gnd.n4229 gnd.n4228 0.152939
R20884 gnd.n4229 gnd.n3906 0.152939
R20885 gnd.n4290 gnd.n3906 0.152939
R20886 gnd.n4291 gnd.n4290 0.152939
R20887 gnd.n4292 gnd.n4291 0.152939
R20888 gnd.n4292 gnd.n3901 0.152939
R20889 gnd.n4304 gnd.n3901 0.152939
R20890 gnd.n4305 gnd.n4304 0.152939
R20891 gnd.n4307 gnd.n4305 0.152939
R20892 gnd.n4307 gnd.n4306 0.152939
R20893 gnd.n4306 gnd.n3892 0.152939
R20894 gnd.n3893 gnd.n3892 0.152939
R20895 gnd.n3999 gnd.n3931 0.152939
R20896 gnd.n3934 gnd.n3931 0.152939
R20897 gnd.n3935 gnd.n3934 0.152939
R20898 gnd.n3938 gnd.n3935 0.152939
R20899 gnd.n3939 gnd.n3938 0.152939
R20900 gnd.n3940 gnd.n3939 0.152939
R20901 gnd.n3941 gnd.n3940 0.152939
R20902 gnd.n3944 gnd.n3941 0.152939
R20903 gnd.n3945 gnd.n3944 0.152939
R20904 gnd.n3946 gnd.n3945 0.152939
R20905 gnd.n3947 gnd.n3946 0.152939
R20906 gnd.n3950 gnd.n3947 0.152939
R20907 gnd.n3951 gnd.n3950 0.152939
R20908 gnd.n3952 gnd.n3951 0.152939
R20909 gnd.n3953 gnd.n3952 0.152939
R20910 gnd.n3957 gnd.n3953 0.152939
R20911 gnd.n3960 gnd.n3957 0.152939
R20912 gnd.n3960 gnd.n3959 0.152939
R20913 gnd.n2505 gnd.n2454 0.152939
R20914 gnd.n2506 gnd.n2505 0.152939
R20915 gnd.n2507 gnd.n2506 0.152939
R20916 gnd.n2508 gnd.n2507 0.152939
R20917 gnd.n2525 gnd.n2508 0.152939
R20918 gnd.n2526 gnd.n2525 0.152939
R20919 gnd.n2527 gnd.n2526 0.152939
R20920 gnd.n2528 gnd.n2527 0.152939
R20921 gnd.n2545 gnd.n2528 0.152939
R20922 gnd.n2546 gnd.n2545 0.152939
R20923 gnd.n2547 gnd.n2546 0.152939
R20924 gnd.n2548 gnd.n2547 0.152939
R20925 gnd.n2566 gnd.n2548 0.152939
R20926 gnd.n2567 gnd.n2566 0.152939
R20927 gnd.n2568 gnd.n2567 0.152939
R20928 gnd.n2569 gnd.n2568 0.152939
R20929 gnd.n2724 gnd.n2723 0.152939
R20930 gnd.n2725 gnd.n2724 0.152939
R20931 gnd.n2726 gnd.n2725 0.152939
R20932 gnd.n2727 gnd.n2726 0.152939
R20933 gnd.n2728 gnd.n2727 0.152939
R20934 gnd.n2729 gnd.n2728 0.152939
R20935 gnd.n2730 gnd.n2729 0.152939
R20936 gnd.n2731 gnd.n2730 0.152939
R20937 gnd.n2732 gnd.n2731 0.152939
R20938 gnd.n2733 gnd.n2732 0.152939
R20939 gnd.n2734 gnd.n2733 0.152939
R20940 gnd.n2735 gnd.n2734 0.152939
R20941 gnd.n2736 gnd.n2735 0.152939
R20942 gnd.n2737 gnd.n2736 0.152939
R20943 gnd.n2738 gnd.n2737 0.152939
R20944 gnd.n2739 gnd.n2738 0.152939
R20945 gnd.n2740 gnd.n2739 0.152939
R20946 gnd.n2743 gnd.n2740 0.152939
R20947 gnd.n2744 gnd.n2743 0.152939
R20948 gnd.n2745 gnd.n2744 0.152939
R20949 gnd.n2746 gnd.n2745 0.152939
R20950 gnd.n2747 gnd.n2746 0.152939
R20951 gnd.n2748 gnd.n2747 0.152939
R20952 gnd.n2749 gnd.n2748 0.152939
R20953 gnd.n2750 gnd.n2749 0.152939
R20954 gnd.n2848 gnd.n2847 0.152939
R20955 gnd.n2847 gnd.n2753 0.152939
R20956 gnd.n2754 gnd.n2753 0.152939
R20957 gnd.n2755 gnd.n2754 0.152939
R20958 gnd.n2756 gnd.n2755 0.152939
R20959 gnd.n2757 gnd.n2756 0.152939
R20960 gnd.n2758 gnd.n2757 0.152939
R20961 gnd.n2759 gnd.n2758 0.152939
R20962 gnd.n2827 gnd.n2759 0.152939
R20963 gnd.n2827 gnd.n2826 0.152939
R20964 gnd.n2826 gnd.n2825 0.152939
R20965 gnd.n2825 gnd.n2763 0.152939
R20966 gnd.n2764 gnd.n2763 0.152939
R20967 gnd.n2765 gnd.n2764 0.152939
R20968 gnd.n2766 gnd.n2765 0.152939
R20969 gnd.n2767 gnd.n2766 0.152939
R20970 gnd.n2768 gnd.n2767 0.152939
R20971 gnd.n2769 gnd.n2768 0.152939
R20972 gnd.n2770 gnd.n2769 0.152939
R20973 gnd.n2771 gnd.n2770 0.152939
R20974 gnd.n2772 gnd.n2771 0.152939
R20975 gnd.n2773 gnd.n2772 0.152939
R20976 gnd.n2774 gnd.n2773 0.152939
R20977 gnd.n2775 gnd.n2774 0.152939
R20978 gnd.n2776 gnd.n2775 0.152939
R20979 gnd.n2777 gnd.n2776 0.152939
R20980 gnd.n2778 gnd.n2777 0.152939
R20981 gnd.n2779 gnd.n2778 0.152939
R20982 gnd.n2785 gnd.n2779 0.152939
R20983 gnd.n2785 gnd.n2784 0.152939
R20984 gnd.n4067 gnd.n4062 0.152939
R20985 gnd.n4068 gnd.n4067 0.152939
R20986 gnd.n4069 gnd.n4068 0.152939
R20987 gnd.n4069 gnd.n4058 0.152939
R20988 gnd.n4077 gnd.n4058 0.152939
R20989 gnd.n4078 gnd.n4077 0.152939
R20990 gnd.n4079 gnd.n4078 0.152939
R20991 gnd.n4079 gnd.n4054 0.152939
R20992 gnd.n4087 gnd.n4054 0.152939
R20993 gnd.n4088 gnd.n4087 0.152939
R20994 gnd.n4089 gnd.n4088 0.152939
R20995 gnd.n4089 gnd.n4050 0.152939
R20996 gnd.n4097 gnd.n4050 0.152939
R20997 gnd.n4098 gnd.n4097 0.152939
R20998 gnd.n4099 gnd.n4098 0.152939
R20999 gnd.n4099 gnd.n4043 0.152939
R21000 gnd.n4107 gnd.n4043 0.152939
R21001 gnd.n4108 gnd.n4107 0.152939
R21002 gnd.n4109 gnd.n4108 0.152939
R21003 gnd.n4109 gnd.n4039 0.152939
R21004 gnd.n4117 gnd.n4039 0.152939
R21005 gnd.n4118 gnd.n4117 0.152939
R21006 gnd.n4119 gnd.n4118 0.152939
R21007 gnd.n4119 gnd.n4035 0.152939
R21008 gnd.n4127 gnd.n4035 0.152939
R21009 gnd.n4128 gnd.n4127 0.152939
R21010 gnd.n4129 gnd.n4128 0.152939
R21011 gnd.n4129 gnd.n4031 0.152939
R21012 gnd.n4137 gnd.n4031 0.152939
R21013 gnd.n4138 gnd.n4137 0.152939
R21014 gnd.n4139 gnd.n4138 0.152939
R21015 gnd.n4139 gnd.n4027 0.152939
R21016 gnd.n4147 gnd.n4027 0.152939
R21017 gnd.n4148 gnd.n4147 0.152939
R21018 gnd.n4149 gnd.n4148 0.152939
R21019 gnd.n4149 gnd.n4023 0.152939
R21020 gnd.n4159 gnd.n4023 0.152939
R21021 gnd.n4160 gnd.n4159 0.152939
R21022 gnd.n4161 gnd.n4160 0.152939
R21023 gnd.n4161 gnd.n4019 0.152939
R21024 gnd.n4169 gnd.n4019 0.152939
R21025 gnd.n4170 gnd.n4169 0.152939
R21026 gnd.n4171 gnd.n4170 0.152939
R21027 gnd.n4171 gnd.n4015 0.152939
R21028 gnd.n4179 gnd.n4015 0.152939
R21029 gnd.n4180 gnd.n4179 0.152939
R21030 gnd.n4181 gnd.n4180 0.152939
R21031 gnd.n4181 gnd.n4011 0.152939
R21032 gnd.n4189 gnd.n4011 0.152939
R21033 gnd.n4190 gnd.n4189 0.152939
R21034 gnd.n4191 gnd.n4190 0.152939
R21035 gnd.n4191 gnd.n4007 0.152939
R21036 gnd.n4199 gnd.n4007 0.152939
R21037 gnd.n4200 gnd.n4199 0.152939
R21038 gnd.n4202 gnd.n4200 0.152939
R21039 gnd.n4202 gnd.n4201 0.152939
R21040 gnd.n4201 gnd.n4000 0.152939
R21041 gnd.n4211 gnd.n4000 0.152939
R21042 gnd.n2371 gnd.n2370 0.152939
R21043 gnd.n2372 gnd.n2371 0.152939
R21044 gnd.n2391 gnd.n2372 0.152939
R21045 gnd.n2392 gnd.n2391 0.152939
R21046 gnd.n2393 gnd.n2392 0.152939
R21047 gnd.n2394 gnd.n2393 0.152939
R21048 gnd.n2412 gnd.n2394 0.152939
R21049 gnd.n2413 gnd.n2412 0.152939
R21050 gnd.n2414 gnd.n2413 0.152939
R21051 gnd.n2415 gnd.n2414 0.152939
R21052 gnd.n2432 gnd.n2415 0.152939
R21053 gnd.n2433 gnd.n2432 0.152939
R21054 gnd.n2434 gnd.n2433 0.152939
R21055 gnd.n2435 gnd.n2434 0.152939
R21056 gnd.n2453 gnd.n2435 0.152939
R21057 gnd.n2454 gnd.n2453 0.152939
R21058 gnd.n6515 gnd.n874 0.152939
R21059 gnd.n2342 gnd.n874 0.152939
R21060 gnd.n2343 gnd.n2342 0.152939
R21061 gnd.n2344 gnd.n2343 0.152939
R21062 gnd.n2349 gnd.n2344 0.152939
R21063 gnd.n2350 gnd.n2349 0.152939
R21064 gnd.n2351 gnd.n2350 0.152939
R21065 gnd.n2352 gnd.n2351 0.152939
R21066 gnd.n2357 gnd.n2352 0.152939
R21067 gnd.n2358 gnd.n2357 0.152939
R21068 gnd.n2359 gnd.n2358 0.152939
R21069 gnd.n2360 gnd.n2359 0.152939
R21070 gnd.n3920 gnd.n2360 0.152939
R21071 gnd.n3921 gnd.n3920 0.152939
R21072 gnd.n4260 gnd.n3921 0.152939
R21073 gnd.n4261 gnd.n4260 0.152939
R21074 gnd.n4262 gnd.n4261 0.152939
R21075 gnd.n4262 gnd.n3916 0.152939
R21076 gnd.n4268 gnd.n3916 0.152939
R21077 gnd.n4269 gnd.n4268 0.152939
R21078 gnd.n4270 gnd.n4269 0.152939
R21079 gnd.n4270 gnd.n3912 0.152939
R21080 gnd.n4276 gnd.n3912 0.152939
R21081 gnd.n4277 gnd.n4276 0.152939
R21082 gnd.n4278 gnd.n4277 0.152939
R21083 gnd.n4279 gnd.n4278 0.152939
R21084 gnd.n4280 gnd.n4279 0.152939
R21085 gnd.n4280 gnd.n3883 0.152939
R21086 gnd.n4364 gnd.n3883 0.152939
R21087 gnd.n6686 gnd.n707 0.152939
R21088 gnd.n712 gnd.n707 0.152939
R21089 gnd.n713 gnd.n712 0.152939
R21090 gnd.n714 gnd.n713 0.152939
R21091 gnd.n715 gnd.n714 0.152939
R21092 gnd.n720 gnd.n715 0.152939
R21093 gnd.n721 gnd.n720 0.152939
R21094 gnd.n722 gnd.n721 0.152939
R21095 gnd.n723 gnd.n722 0.152939
R21096 gnd.n728 gnd.n723 0.152939
R21097 gnd.n729 gnd.n728 0.152939
R21098 gnd.n730 gnd.n729 0.152939
R21099 gnd.n731 gnd.n730 0.152939
R21100 gnd.n736 gnd.n731 0.152939
R21101 gnd.n737 gnd.n736 0.152939
R21102 gnd.n738 gnd.n737 0.152939
R21103 gnd.n739 gnd.n738 0.152939
R21104 gnd.n744 gnd.n739 0.152939
R21105 gnd.n745 gnd.n744 0.152939
R21106 gnd.n746 gnd.n745 0.152939
R21107 gnd.n747 gnd.n746 0.152939
R21108 gnd.n752 gnd.n747 0.152939
R21109 gnd.n753 gnd.n752 0.152939
R21110 gnd.n754 gnd.n753 0.152939
R21111 gnd.n755 gnd.n754 0.152939
R21112 gnd.n760 gnd.n755 0.152939
R21113 gnd.n761 gnd.n760 0.152939
R21114 gnd.n762 gnd.n761 0.152939
R21115 gnd.n763 gnd.n762 0.152939
R21116 gnd.n768 gnd.n763 0.152939
R21117 gnd.n769 gnd.n768 0.152939
R21118 gnd.n770 gnd.n769 0.152939
R21119 gnd.n771 gnd.n770 0.152939
R21120 gnd.n776 gnd.n771 0.152939
R21121 gnd.n777 gnd.n776 0.152939
R21122 gnd.n778 gnd.n777 0.152939
R21123 gnd.n779 gnd.n778 0.152939
R21124 gnd.n784 gnd.n779 0.152939
R21125 gnd.n785 gnd.n784 0.152939
R21126 gnd.n786 gnd.n785 0.152939
R21127 gnd.n787 gnd.n786 0.152939
R21128 gnd.n792 gnd.n787 0.152939
R21129 gnd.n793 gnd.n792 0.152939
R21130 gnd.n794 gnd.n793 0.152939
R21131 gnd.n795 gnd.n794 0.152939
R21132 gnd.n800 gnd.n795 0.152939
R21133 gnd.n801 gnd.n800 0.152939
R21134 gnd.n802 gnd.n801 0.152939
R21135 gnd.n803 gnd.n802 0.152939
R21136 gnd.n808 gnd.n803 0.152939
R21137 gnd.n809 gnd.n808 0.152939
R21138 gnd.n810 gnd.n809 0.152939
R21139 gnd.n811 gnd.n810 0.152939
R21140 gnd.n816 gnd.n811 0.152939
R21141 gnd.n817 gnd.n816 0.152939
R21142 gnd.n818 gnd.n817 0.152939
R21143 gnd.n819 gnd.n818 0.152939
R21144 gnd.n824 gnd.n819 0.152939
R21145 gnd.n825 gnd.n824 0.152939
R21146 gnd.n826 gnd.n825 0.152939
R21147 gnd.n827 gnd.n826 0.152939
R21148 gnd.n832 gnd.n827 0.152939
R21149 gnd.n833 gnd.n832 0.152939
R21150 gnd.n834 gnd.n833 0.152939
R21151 gnd.n835 gnd.n834 0.152939
R21152 gnd.n840 gnd.n835 0.152939
R21153 gnd.n841 gnd.n840 0.152939
R21154 gnd.n842 gnd.n841 0.152939
R21155 gnd.n843 gnd.n842 0.152939
R21156 gnd.n848 gnd.n843 0.152939
R21157 gnd.n849 gnd.n848 0.152939
R21158 gnd.n850 gnd.n849 0.152939
R21159 gnd.n851 gnd.n850 0.152939
R21160 gnd.n856 gnd.n851 0.152939
R21161 gnd.n857 gnd.n856 0.152939
R21162 gnd.n858 gnd.n857 0.152939
R21163 gnd.n859 gnd.n858 0.152939
R21164 gnd.n864 gnd.n859 0.152939
R21165 gnd.n865 gnd.n864 0.152939
R21166 gnd.n866 gnd.n865 0.152939
R21167 gnd.n867 gnd.n866 0.152939
R21168 gnd.n872 gnd.n867 0.152939
R21169 gnd.n873 gnd.n872 0.152939
R21170 gnd.n6516 gnd.n873 0.152939
R21171 gnd.n3835 gnd.n3834 0.152939
R21172 gnd.n3835 gnd.n3754 0.152939
R21173 gnd.n4488 gnd.n3754 0.152939
R21174 gnd.n4489 gnd.n4488 0.152939
R21175 gnd.n4496 gnd.n4489 0.152939
R21176 gnd.n4496 gnd.n4495 0.152939
R21177 gnd.n4495 gnd.n4494 0.152939
R21178 gnd.n4494 gnd.n4491 0.152939
R21179 gnd.n4491 gnd.n4490 0.152939
R21180 gnd.n4490 gnd.n3730 0.152939
R21181 gnd.n4544 gnd.n3730 0.152939
R21182 gnd.n4545 gnd.n4544 0.152939
R21183 gnd.n4551 gnd.n4545 0.152939
R21184 gnd.n4551 gnd.n4550 0.152939
R21185 gnd.n4550 gnd.n4549 0.152939
R21186 gnd.n4549 gnd.n4546 0.152939
R21187 gnd.n4546 gnd.n3698 0.152939
R21188 gnd.n4610 gnd.n3698 0.152939
R21189 gnd.n4611 gnd.n4610 0.152939
R21190 gnd.n4619 gnd.n4611 0.152939
R21191 gnd.n4619 gnd.n4618 0.152939
R21192 gnd.n4618 gnd.n4617 0.152939
R21193 gnd.n4617 gnd.n4612 0.152939
R21194 gnd.n4612 gnd.n3657 0.152939
R21195 gnd.n4698 gnd.n3657 0.152939
R21196 gnd.n4699 gnd.n4698 0.152939
R21197 gnd.n4736 gnd.n4699 0.152939
R21198 gnd.n4736 gnd.n4735 0.152939
R21199 gnd.n4735 gnd.n4734 0.152939
R21200 gnd.n4734 gnd.n4700 0.152939
R21201 gnd.n4730 gnd.n4700 0.152939
R21202 gnd.n4730 gnd.n4729 0.152939
R21203 gnd.n4729 gnd.n4728 0.152939
R21204 gnd.n4728 gnd.n4705 0.152939
R21205 gnd.n4724 gnd.n4705 0.152939
R21206 gnd.n4724 gnd.n4723 0.152939
R21207 gnd.n4723 gnd.n4722 0.152939
R21208 gnd.n4722 gnd.n4710 0.152939
R21209 gnd.n4718 gnd.n4710 0.152939
R21210 gnd.n4718 gnd.n4717 0.152939
R21211 gnd.n4717 gnd.n3570 0.152939
R21212 gnd.n4875 gnd.n3570 0.152939
R21213 gnd.n4876 gnd.n4875 0.152939
R21214 gnd.n4891 gnd.n4876 0.152939
R21215 gnd.n4891 gnd.n4890 0.152939
R21216 gnd.n4890 gnd.n4889 0.152939
R21217 gnd.n4889 gnd.n4877 0.152939
R21218 gnd.n4885 gnd.n4877 0.152939
R21219 gnd.n4885 gnd.n4884 0.152939
R21220 gnd.n4884 gnd.n3521 0.152939
R21221 gnd.n4962 gnd.n3521 0.152939
R21222 gnd.n4963 gnd.n4962 0.152939
R21223 gnd.n4968 gnd.n4963 0.152939
R21224 gnd.n4968 gnd.n4967 0.152939
R21225 gnd.n4967 gnd.n4966 0.152939
R21226 gnd.n4966 gnd.n3492 0.152939
R21227 gnd.n5030 gnd.n3492 0.152939
R21228 gnd.n5031 gnd.n5030 0.152939
R21229 gnd.n5046 gnd.n5031 0.152939
R21230 gnd.n5046 gnd.n5045 0.152939
R21231 gnd.n5045 gnd.n5044 0.152939
R21232 gnd.n5044 gnd.n5032 0.152939
R21233 gnd.n5040 gnd.n5032 0.152939
R21234 gnd.n5040 gnd.n5039 0.152939
R21235 gnd.n5039 gnd.n3417 0.152939
R21236 gnd.n5115 gnd.n3417 0.152939
R21237 gnd.n5116 gnd.n5115 0.152939
R21238 gnd.n5118 gnd.n5116 0.152939
R21239 gnd.n5118 gnd.n5117 0.152939
R21240 gnd.n5117 gnd.n3387 0.152939
R21241 gnd.n5151 gnd.n3387 0.152939
R21242 gnd.n5152 gnd.n5151 0.152939
R21243 gnd.n5153 gnd.n5152 0.152939
R21244 gnd.n5153 gnd.n3366 0.152939
R21245 gnd.n5182 gnd.n3366 0.152939
R21246 gnd.n5183 gnd.n5182 0.152939
R21247 gnd.n5184 gnd.n5183 0.152939
R21248 gnd.n5184 gnd.n3362 0.152939
R21249 gnd.n5192 gnd.n3362 0.152939
R21250 gnd.n5193 gnd.n5192 0.152939
R21251 gnd.n5373 gnd.n5193 0.152939
R21252 gnd.n5373 gnd.n5372 0.152939
R21253 gnd.n4348 gnd.n4347 0.152939
R21254 gnd.n4347 gnd.n3896 0.152939
R21255 gnd.n4343 gnd.n3896 0.152939
R21256 gnd.n4343 gnd.n3872 0.152939
R21257 gnd.n4393 gnd.n3872 0.152939
R21258 gnd.n4394 gnd.n4393 0.152939
R21259 gnd.n4395 gnd.n4394 0.152939
R21260 gnd.n4395 gnd.n3866 0.152939
R21261 gnd.n4407 gnd.n3866 0.152939
R21262 gnd.n4408 gnd.n4407 0.152939
R21263 gnd.n4409 gnd.n4408 0.152939
R21264 gnd.n4409 gnd.n3860 0.152939
R21265 gnd.n4433 gnd.n3860 0.152939
R21266 gnd.n4433 gnd.n4432 0.152939
R21267 gnd.n4432 gnd.n4431 0.152939
R21268 gnd.n4431 gnd.n3861 0.152939
R21269 gnd.n4427 gnd.n3861 0.152939
R21270 gnd.n4427 gnd.n2581 0.152939
R21271 gnd.n6347 gnd.n2581 0.152939
R21272 gnd.n6347 gnd.n6346 0.152939
R21273 gnd.n6334 gnd.n2605 0.152939
R21274 gnd.n6334 gnd.n6333 0.152939
R21275 gnd.n6333 gnd.n6332 0.152939
R21276 gnd.n6332 gnd.n2607 0.152939
R21277 gnd.n6328 gnd.n2607 0.152939
R21278 gnd.n6328 gnd.n6327 0.152939
R21279 gnd.n4479 gnd.n3830 0.152939
R21280 gnd.n4480 gnd.n4479 0.152939
R21281 gnd.n4482 gnd.n4480 0.152939
R21282 gnd.n4482 gnd.n4481 0.152939
R21283 gnd.n4481 gnd.n3742 0.152939
R21284 gnd.n4511 gnd.n3742 0.152939
R21285 gnd.n4512 gnd.n4511 0.152939
R21286 gnd.n4514 gnd.n4512 0.152939
R21287 gnd.n4514 gnd.n4513 0.152939
R21288 gnd.n4513 gnd.n2947 0.152939
R21289 gnd.n6125 gnd.n2947 0.152939
R21290 gnd.n6125 gnd.n6124 0.152939
R21291 gnd.n6124 gnd.n6123 0.152939
R21292 gnd.n6123 gnd.n2948 0.152939
R21293 gnd.n6119 gnd.n2948 0.152939
R21294 gnd.n6119 gnd.n6118 0.152939
R21295 gnd.n6118 gnd.n6117 0.152939
R21296 gnd.n6117 gnd.n2953 0.152939
R21297 gnd.n6113 gnd.n2953 0.152939
R21298 gnd.n6113 gnd.n6112 0.152939
R21299 gnd.n6112 gnd.n6111 0.152939
R21300 gnd.n6111 gnd.n2958 0.152939
R21301 gnd.n6107 gnd.n2958 0.152939
R21302 gnd.n6107 gnd.n6106 0.152939
R21303 gnd.n6106 gnd.n6105 0.152939
R21304 gnd.n6105 gnd.n2963 0.152939
R21305 gnd.n6101 gnd.n2963 0.152939
R21306 gnd.n6101 gnd.n6100 0.152939
R21307 gnd.n6100 gnd.n6099 0.152939
R21308 gnd.n6099 gnd.n2968 0.152939
R21309 gnd.n6095 gnd.n2968 0.152939
R21310 gnd.n6095 gnd.n6094 0.152939
R21311 gnd.n6094 gnd.n6093 0.152939
R21312 gnd.n6093 gnd.n2973 0.152939
R21313 gnd.n6089 gnd.n2973 0.152939
R21314 gnd.n6089 gnd.n6088 0.152939
R21315 gnd.n6088 gnd.n6087 0.152939
R21316 gnd.n6087 gnd.n2978 0.152939
R21317 gnd.n6083 gnd.n2978 0.152939
R21318 gnd.n6083 gnd.n6082 0.152939
R21319 gnd.n6082 gnd.n6081 0.152939
R21320 gnd.n6081 gnd.n2983 0.152939
R21321 gnd.n6077 gnd.n2983 0.152939
R21322 gnd.n6077 gnd.n6076 0.152939
R21323 gnd.n6076 gnd.n6075 0.152939
R21324 gnd.n6075 gnd.n2988 0.152939
R21325 gnd.n6071 gnd.n2988 0.152939
R21326 gnd.n6071 gnd.n6070 0.152939
R21327 gnd.n6070 gnd.n6069 0.152939
R21328 gnd.n6069 gnd.n2993 0.152939
R21329 gnd.n6065 gnd.n2993 0.152939
R21330 gnd.n6065 gnd.n6064 0.152939
R21331 gnd.n6064 gnd.n6063 0.152939
R21332 gnd.n6063 gnd.n2998 0.152939
R21333 gnd.n6059 gnd.n2998 0.152939
R21334 gnd.n6059 gnd.n6058 0.152939
R21335 gnd.n6058 gnd.n6057 0.152939
R21336 gnd.n6057 gnd.n3003 0.152939
R21337 gnd.n6053 gnd.n3003 0.152939
R21338 gnd.n6053 gnd.n6052 0.152939
R21339 gnd.n6052 gnd.n6051 0.152939
R21340 gnd.n6051 gnd.n3008 0.152939
R21341 gnd.n6047 gnd.n3008 0.152939
R21342 gnd.n6047 gnd.n6046 0.152939
R21343 gnd.n6046 gnd.n6045 0.152939
R21344 gnd.n6045 gnd.n3013 0.152939
R21345 gnd.n6041 gnd.n3013 0.152939
R21346 gnd.n6041 gnd.n6040 0.152939
R21347 gnd.n6040 gnd.n6039 0.152939
R21348 gnd.n6039 gnd.n3018 0.152939
R21349 gnd.n6035 gnd.n3018 0.152939
R21350 gnd.n6035 gnd.n6034 0.152939
R21351 gnd.n6034 gnd.n6033 0.152939
R21352 gnd.n6033 gnd.n3023 0.152939
R21353 gnd.n6029 gnd.n3023 0.152939
R21354 gnd.n6029 gnd.n6028 0.152939
R21355 gnd.n6028 gnd.n6027 0.152939
R21356 gnd.n6027 gnd.n3028 0.152939
R21357 gnd.n6023 gnd.n3028 0.152939
R21358 gnd.n6023 gnd.n6022 0.152939
R21359 gnd.n6022 gnd.n6021 0.152939
R21360 gnd.n6021 gnd.n3033 0.152939
R21361 gnd.n5259 gnd.n5258 0.152939
R21362 gnd.n5259 gnd.n5254 0.152939
R21363 gnd.n5267 gnd.n5254 0.152939
R21364 gnd.n5268 gnd.n5267 0.152939
R21365 gnd.n5270 gnd.n5268 0.152939
R21366 gnd.n5270 gnd.n5269 0.152939
R21367 gnd.n5199 gnd.n5194 0.152939
R21368 gnd.n5194 gnd.n3261 0.152939
R21369 gnd.n5733 gnd.n3261 0.152939
R21370 gnd.n5734 gnd.n5733 0.152939
R21371 gnd.n5735 gnd.n5734 0.152939
R21372 gnd.n5735 gnd.n3256 0.152939
R21373 gnd.n5755 gnd.n3256 0.152939
R21374 gnd.n5755 gnd.n5754 0.152939
R21375 gnd.n5754 gnd.n5753 0.152939
R21376 gnd.n5753 gnd.n3257 0.152939
R21377 gnd.n5749 gnd.n3257 0.152939
R21378 gnd.n5749 gnd.n3244 0.152939
R21379 gnd.n5813 gnd.n3244 0.152939
R21380 gnd.n5814 gnd.n5813 0.152939
R21381 gnd.n5825 gnd.n5814 0.152939
R21382 gnd.n5825 gnd.n5824 0.152939
R21383 gnd.n5824 gnd.n5823 0.152939
R21384 gnd.n5823 gnd.n5815 0.152939
R21385 gnd.n5819 gnd.n5815 0.152939
R21386 gnd.n5819 gnd.n63 0.152939
R21387 gnd.n7736 gnd.n7735 0.145814
R21388 gnd.n4349 gnd.n3893 0.145814
R21389 gnd.n4349 gnd.n4348 0.145814
R21390 gnd.n7736 gnd.n63 0.145814
R21391 gnd.n6327 gnd.n6326 0.128549
R21392 gnd.n5269 gnd.n3265 0.128549
R21393 gnd.n1154 gnd.n0 0.127478
R21394 gnd.n3183 gnd.n79 0.10111
R21395 gnd.n4365 gnd.n4364 0.10111
R21396 gnd.n1734 gnd.n1733 0.0767195
R21397 gnd.n1733 gnd.n1732 0.0767195
R21398 gnd.n6326 gnd.n2577 0.063
R21399 gnd.n5722 gnd.n3265 0.063
R21400 gnd.n5724 gnd.n5722 0.0538288
R21401 gnd.n7672 gnd.n174 0.0538288
R21402 gnd.n4214 gnd.n4212 0.0538288
R21403 gnd.n6354 gnd.n2577 0.0538288
R21404 gnd.n4366 gnd.n4365 0.0523293
R21405 gnd.n5792 gnd.n79 0.0523293
R21406 gnd.n2302 gnd.n918 0.0477147
R21407 gnd.n1497 gnd.n1385 0.0442063
R21408 gnd.n1498 gnd.n1497 0.0442063
R21409 gnd.n1499 gnd.n1498 0.0442063
R21410 gnd.n1499 gnd.n1374 0.0442063
R21411 gnd.n1513 gnd.n1374 0.0442063
R21412 gnd.n1514 gnd.n1513 0.0442063
R21413 gnd.n1515 gnd.n1514 0.0442063
R21414 gnd.n1515 gnd.n1361 0.0442063
R21415 gnd.n1559 gnd.n1361 0.0442063
R21416 gnd.n1560 gnd.n1559 0.0442063
R21417 gnd.n1562 gnd.n1295 0.0344674
R21418 gnd.n5725 gnd.n5724 0.0344674
R21419 gnd.n5725 gnd.n3075 0.0344674
R21420 gnd.n3076 gnd.n3075 0.0344674
R21421 gnd.n3077 gnd.n3076 0.0344674
R21422 gnd.n3259 gnd.n3077 0.0344674
R21423 gnd.n3259 gnd.n3095 0.0344674
R21424 gnd.n3096 gnd.n3095 0.0344674
R21425 gnd.n3097 gnd.n3096 0.0344674
R21426 gnd.n5744 gnd.n3097 0.0344674
R21427 gnd.n5744 gnd.n3116 0.0344674
R21428 gnd.n3117 gnd.n3116 0.0344674
R21429 gnd.n3118 gnd.n3117 0.0344674
R21430 gnd.n5807 gnd.n3118 0.0344674
R21431 gnd.n5807 gnd.n3135 0.0344674
R21432 gnd.n3136 gnd.n3135 0.0344674
R21433 gnd.n3137 gnd.n3136 0.0344674
R21434 gnd.n3239 gnd.n3137 0.0344674
R21435 gnd.n5836 gnd.n3239 0.0344674
R21436 gnd.n5841 gnd.n5836 0.0344674
R21437 gnd.n5842 gnd.n5841 0.0344674
R21438 gnd.n5842 gnd.n3169 0.0344674
R21439 gnd.n3170 gnd.n3169 0.0344674
R21440 gnd.n3171 gnd.n3170 0.0344674
R21441 gnd.n3172 gnd.n3171 0.0344674
R21442 gnd.n5850 gnd.n3172 0.0344674
R21443 gnd.n5850 gnd.n93 0.0344674
R21444 gnd.n94 gnd.n93 0.0344674
R21445 gnd.n95 gnd.n94 0.0344674
R21446 gnd.n3234 gnd.n95 0.0344674
R21447 gnd.n3234 gnd.n112 0.0344674
R21448 gnd.n113 gnd.n112 0.0344674
R21449 gnd.n114 gnd.n113 0.0344674
R21450 gnd.n5876 gnd.n114 0.0344674
R21451 gnd.n5876 gnd.n133 0.0344674
R21452 gnd.n134 gnd.n133 0.0344674
R21453 gnd.n135 gnd.n134 0.0344674
R21454 gnd.n5883 gnd.n135 0.0344674
R21455 gnd.n5883 gnd.n154 0.0344674
R21456 gnd.n155 gnd.n154 0.0344674
R21457 gnd.n156 gnd.n155 0.0344674
R21458 gnd.n173 gnd.n156 0.0344674
R21459 gnd.n7672 gnd.n173 0.0344674
R21460 gnd.n4215 gnd.n4214 0.0344674
R21461 gnd.n4215 gnd.n2381 0.0344674
R21462 gnd.n2382 gnd.n2381 0.0344674
R21463 gnd.n2383 gnd.n2382 0.0344674
R21464 gnd.n4218 gnd.n2383 0.0344674
R21465 gnd.n4218 gnd.n2402 0.0344674
R21466 gnd.n2403 gnd.n2402 0.0344674
R21467 gnd.n2404 gnd.n2403 0.0344674
R21468 gnd.n4225 gnd.n2404 0.0344674
R21469 gnd.n4225 gnd.n2423 0.0344674
R21470 gnd.n2424 gnd.n2423 0.0344674
R21471 gnd.n2425 gnd.n2424 0.0344674
R21472 gnd.n3904 gnd.n2425 0.0344674
R21473 gnd.n3904 gnd.n2443 0.0344674
R21474 gnd.n2444 gnd.n2443 0.0344674
R21475 gnd.n2445 gnd.n2444 0.0344674
R21476 gnd.n3899 gnd.n2445 0.0344674
R21477 gnd.n3899 gnd.n2462 0.0344674
R21478 gnd.n2463 gnd.n2462 0.0344674
R21479 gnd.n2464 gnd.n2463 0.0344674
R21480 gnd.n4316 gnd.n2464 0.0344674
R21481 gnd.n4316 gnd.n2478 0.0344674
R21482 gnd.n2479 gnd.n2478 0.0344674
R21483 gnd.n2480 gnd.n2479 0.0344674
R21484 gnd.n4336 gnd.n2480 0.0344674
R21485 gnd.n4336 gnd.n2496 0.0344674
R21486 gnd.n2497 gnd.n2496 0.0344674
R21487 gnd.n2498 gnd.n2497 0.0344674
R21488 gnd.n3870 gnd.n2498 0.0344674
R21489 gnd.n3870 gnd.n2515 0.0344674
R21490 gnd.n2516 gnd.n2515 0.0344674
R21491 gnd.n2517 gnd.n2516 0.0344674
R21492 gnd.n3864 gnd.n2517 0.0344674
R21493 gnd.n3864 gnd.n2536 0.0344674
R21494 gnd.n2537 gnd.n2536 0.0344674
R21495 gnd.n2538 gnd.n2537 0.0344674
R21496 gnd.n4418 gnd.n2538 0.0344674
R21497 gnd.n4418 gnd.n2556 0.0344674
R21498 gnd.n2557 gnd.n2556 0.0344674
R21499 gnd.n2558 gnd.n2557 0.0344674
R21500 gnd.n2576 gnd.n2558 0.0344674
R21501 gnd.n6354 gnd.n2576 0.0344674
R21502 gnd.n6325 gnd.n2612 0.0344674
R21503 gnd.n5279 gnd.n5278 0.0344674
R21504 gnd.n6345 gnd.n6344 0.029712
R21505 gnd.n5209 gnd.n5200 0.029712
R21506 gnd.n1582 gnd.n1581 0.0269946
R21507 gnd.n1584 gnd.n1583 0.0269946
R21508 gnd.n1290 gnd.n1288 0.0269946
R21509 gnd.n1594 gnd.n1592 0.0269946
R21510 gnd.n1593 gnd.n1269 0.0269946
R21511 gnd.n1613 gnd.n1612 0.0269946
R21512 gnd.n1615 gnd.n1614 0.0269946
R21513 gnd.n1264 gnd.n1263 0.0269946
R21514 gnd.n1625 gnd.n1259 0.0269946
R21515 gnd.n1624 gnd.n1261 0.0269946
R21516 gnd.n1260 gnd.n1242 0.0269946
R21517 gnd.n1645 gnd.n1243 0.0269946
R21518 gnd.n1644 gnd.n1244 0.0269946
R21519 gnd.n1678 gnd.n1219 0.0269946
R21520 gnd.n1680 gnd.n1679 0.0269946
R21521 gnd.n1681 gnd.n1166 0.0269946
R21522 gnd.n1214 gnd.n1167 0.0269946
R21523 gnd.n1216 gnd.n1168 0.0269946
R21524 gnd.n1691 gnd.n1690 0.0269946
R21525 gnd.n1693 gnd.n1692 0.0269946
R21526 gnd.n1694 gnd.n1188 0.0269946
R21527 gnd.n1696 gnd.n1189 0.0269946
R21528 gnd.n1699 gnd.n1190 0.0269946
R21529 gnd.n1702 gnd.n1701 0.0269946
R21530 gnd.n1704 gnd.n1703 0.0269946
R21531 gnd.n1769 gnd.n1089 0.0269946
R21532 gnd.n1771 gnd.n1770 0.0269946
R21533 gnd.n1780 gnd.n1082 0.0269946
R21534 gnd.n1782 gnd.n1781 0.0269946
R21535 gnd.n1783 gnd.n1080 0.0269946
R21536 gnd.n1790 gnd.n1786 0.0269946
R21537 gnd.n1789 gnd.n1788 0.0269946
R21538 gnd.n1787 gnd.n1059 0.0269946
R21539 gnd.n1812 gnd.n1060 0.0269946
R21540 gnd.n1811 gnd.n1061 0.0269946
R21541 gnd.n1856 gnd.n1036 0.0269946
R21542 gnd.n1858 gnd.n1857 0.0269946
R21543 gnd.n1867 gnd.n1029 0.0269946
R21544 gnd.n1869 gnd.n1868 0.0269946
R21545 gnd.n1870 gnd.n1027 0.0269946
R21546 gnd.n1877 gnd.n1873 0.0269946
R21547 gnd.n1876 gnd.n1875 0.0269946
R21548 gnd.n1874 gnd.n1006 0.0269946
R21549 gnd.n1899 gnd.n1007 0.0269946
R21550 gnd.n1898 gnd.n1008 0.0269946
R21551 gnd.n1945 gnd.n982 0.0269946
R21552 gnd.n1947 gnd.n1946 0.0269946
R21553 gnd.n1956 gnd.n975 0.0269946
R21554 gnd.n2215 gnd.n973 0.0269946
R21555 gnd.n2220 gnd.n2218 0.0269946
R21556 gnd.n2219 gnd.n954 0.0269946
R21557 gnd.n2244 gnd.n2243 0.0269946
R21558 gnd.n6321 gnd.n2618 0.0225788
R21559 gnd.n6320 gnd.n2619 0.0225788
R21560 gnd.n6317 gnd.n6316 0.0225788
R21561 gnd.n6313 gnd.n2624 0.0225788
R21562 gnd.n6312 gnd.n2630 0.0225788
R21563 gnd.n6309 gnd.n6308 0.0225788
R21564 gnd.n6305 gnd.n2634 0.0225788
R21565 gnd.n6304 gnd.n2638 0.0225788
R21566 gnd.n6301 gnd.n6300 0.0225788
R21567 gnd.n6297 gnd.n2642 0.0225788
R21568 gnd.n6296 gnd.n2648 0.0225788
R21569 gnd.n6293 gnd.n6292 0.0225788
R21570 gnd.n6289 gnd.n2652 0.0225788
R21571 gnd.n6288 gnd.n2656 0.0225788
R21572 gnd.n6285 gnd.n6284 0.0225788
R21573 gnd.n6281 gnd.n2660 0.0225788
R21574 gnd.n6280 gnd.n2669 0.0225788
R21575 gnd.n2674 gnd.n2673 0.0225788
R21576 gnd.n6344 gnd.n2583 0.0225788
R21577 gnd.n5285 gnd.n5283 0.0225788
R21578 gnd.n5284 gnd.n5246 0.0225788
R21579 gnd.n5294 gnd.n5293 0.0225788
R21580 gnd.n5247 gnd.n5242 0.0225788
R21581 gnd.n5304 gnd.n5302 0.0225788
R21582 gnd.n5303 gnd.n5237 0.0225788
R21583 gnd.n5313 gnd.n5312 0.0225788
R21584 gnd.n5238 gnd.n5233 0.0225788
R21585 gnd.n5323 gnd.n5321 0.0225788
R21586 gnd.n5322 gnd.n5228 0.0225788
R21587 gnd.n5332 gnd.n5331 0.0225788
R21588 gnd.n5229 gnd.n5224 0.0225788
R21589 gnd.n5342 gnd.n5340 0.0225788
R21590 gnd.n5341 gnd.n5219 0.0225788
R21591 gnd.n5352 gnd.n5351 0.0225788
R21592 gnd.n5348 gnd.n5220 0.0225788
R21593 gnd.n5362 gnd.n5207 0.0225788
R21594 gnd.n5361 gnd.n5208 0.0225788
R21595 gnd.n5210 gnd.n5209 0.0225788
R21596 gnd.n5371 gnd.n5200 0.0218415
R21597 gnd.n6345 gnd.n2582 0.0218415
R21598 gnd.n1562 gnd.n1561 0.0202011
R21599 gnd.n1561 gnd.n1560 0.0148637
R21600 gnd.n2213 gnd.n1957 0.0144266
R21601 gnd.n2214 gnd.n2213 0.0130679
R21602 gnd.n2618 gnd.n2612 0.0123886
R21603 gnd.n6321 gnd.n6320 0.0123886
R21604 gnd.n6317 gnd.n2619 0.0123886
R21605 gnd.n6316 gnd.n2624 0.0123886
R21606 gnd.n6313 gnd.n6312 0.0123886
R21607 gnd.n6309 gnd.n2630 0.0123886
R21608 gnd.n6308 gnd.n2634 0.0123886
R21609 gnd.n6305 gnd.n6304 0.0123886
R21610 gnd.n6301 gnd.n2638 0.0123886
R21611 gnd.n6300 gnd.n2642 0.0123886
R21612 gnd.n6297 gnd.n6296 0.0123886
R21613 gnd.n6293 gnd.n2648 0.0123886
R21614 gnd.n6292 gnd.n2652 0.0123886
R21615 gnd.n6289 gnd.n6288 0.0123886
R21616 gnd.n6285 gnd.n2656 0.0123886
R21617 gnd.n6284 gnd.n2660 0.0123886
R21618 gnd.n6281 gnd.n6280 0.0123886
R21619 gnd.n2674 gnd.n2669 0.0123886
R21620 gnd.n2673 gnd.n2583 0.0123886
R21621 gnd.n5283 gnd.n5279 0.0123886
R21622 gnd.n5285 gnd.n5284 0.0123886
R21623 gnd.n5294 gnd.n5246 0.0123886
R21624 gnd.n5293 gnd.n5247 0.0123886
R21625 gnd.n5302 gnd.n5242 0.0123886
R21626 gnd.n5304 gnd.n5303 0.0123886
R21627 gnd.n5313 gnd.n5237 0.0123886
R21628 gnd.n5312 gnd.n5238 0.0123886
R21629 gnd.n5321 gnd.n5233 0.0123886
R21630 gnd.n5323 gnd.n5322 0.0123886
R21631 gnd.n5332 gnd.n5228 0.0123886
R21632 gnd.n5331 gnd.n5229 0.0123886
R21633 gnd.n5340 gnd.n5224 0.0123886
R21634 gnd.n5342 gnd.n5341 0.0123886
R21635 gnd.n5352 gnd.n5219 0.0123886
R21636 gnd.n5351 gnd.n5220 0.0123886
R21637 gnd.n5348 gnd.n5207 0.0123886
R21638 gnd.n5362 gnd.n5361 0.0123886
R21639 gnd.n5210 gnd.n5208 0.0123886
R21640 gnd.n1581 gnd.n1295 0.00797283
R21641 gnd.n1583 gnd.n1582 0.00797283
R21642 gnd.n1584 gnd.n1290 0.00797283
R21643 gnd.n1592 gnd.n1288 0.00797283
R21644 gnd.n1594 gnd.n1593 0.00797283
R21645 gnd.n1612 gnd.n1269 0.00797283
R21646 gnd.n1614 gnd.n1613 0.00797283
R21647 gnd.n1615 gnd.n1264 0.00797283
R21648 gnd.n1263 gnd.n1259 0.00797283
R21649 gnd.n1625 gnd.n1624 0.00797283
R21650 gnd.n1261 gnd.n1260 0.00797283
R21651 gnd.n1243 gnd.n1242 0.00797283
R21652 gnd.n1645 gnd.n1644 0.00797283
R21653 gnd.n1244 gnd.n1219 0.00797283
R21654 gnd.n1679 gnd.n1678 0.00797283
R21655 gnd.n1681 gnd.n1680 0.00797283
R21656 gnd.n1214 gnd.n1166 0.00797283
R21657 gnd.n1216 gnd.n1167 0.00797283
R21658 gnd.n1690 gnd.n1168 0.00797283
R21659 gnd.n1692 gnd.n1691 0.00797283
R21660 gnd.n1694 gnd.n1693 0.00797283
R21661 gnd.n1696 gnd.n1188 0.00797283
R21662 gnd.n1699 gnd.n1189 0.00797283
R21663 gnd.n1701 gnd.n1190 0.00797283
R21664 gnd.n1704 gnd.n1702 0.00797283
R21665 gnd.n1703 gnd.n1089 0.00797283
R21666 gnd.n1771 gnd.n1769 0.00797283
R21667 gnd.n1770 gnd.n1082 0.00797283
R21668 gnd.n1781 gnd.n1780 0.00797283
R21669 gnd.n1783 gnd.n1782 0.00797283
R21670 gnd.n1786 gnd.n1080 0.00797283
R21671 gnd.n1790 gnd.n1789 0.00797283
R21672 gnd.n1788 gnd.n1787 0.00797283
R21673 gnd.n1060 gnd.n1059 0.00797283
R21674 gnd.n1812 gnd.n1811 0.00797283
R21675 gnd.n1061 gnd.n1036 0.00797283
R21676 gnd.n1858 gnd.n1856 0.00797283
R21677 gnd.n1857 gnd.n1029 0.00797283
R21678 gnd.n1868 gnd.n1867 0.00797283
R21679 gnd.n1870 gnd.n1869 0.00797283
R21680 gnd.n1873 gnd.n1027 0.00797283
R21681 gnd.n1877 gnd.n1876 0.00797283
R21682 gnd.n1875 gnd.n1874 0.00797283
R21683 gnd.n1007 gnd.n1006 0.00797283
R21684 gnd.n1899 gnd.n1898 0.00797283
R21685 gnd.n1008 gnd.n982 0.00797283
R21686 gnd.n1947 gnd.n1945 0.00797283
R21687 gnd.n1946 gnd.n975 0.00797283
R21688 gnd.n1957 gnd.n1956 0.00797283
R21689 gnd.n2215 gnd.n2214 0.00797283
R21690 gnd.n2218 gnd.n973 0.00797283
R21691 gnd.n2220 gnd.n2219 0.00797283
R21692 gnd.n2243 gnd.n954 0.00797283
R21693 gnd.n2244 gnd.n918 0.00797283
R21694 gnd.n6326 gnd.n6325 0.00593478
R21695 gnd.n5278 gnd.n3265 0.00593478
R21696 CSoutput.n19 CSoutput.t192 184.661
R21697 CSoutput.n78 CSoutput.n77 165.8
R21698 CSoutput.n76 CSoutput.n0 165.8
R21699 CSoutput.n75 CSoutput.n74 165.8
R21700 CSoutput.n73 CSoutput.n72 165.8
R21701 CSoutput.n71 CSoutput.n2 165.8
R21702 CSoutput.n69 CSoutput.n68 165.8
R21703 CSoutput.n67 CSoutput.n3 165.8
R21704 CSoutput.n66 CSoutput.n65 165.8
R21705 CSoutput.n63 CSoutput.n4 165.8
R21706 CSoutput.n61 CSoutput.n60 165.8
R21707 CSoutput.n59 CSoutput.n5 165.8
R21708 CSoutput.n58 CSoutput.n57 165.8
R21709 CSoutput.n55 CSoutput.n6 165.8
R21710 CSoutput.n54 CSoutput.n53 165.8
R21711 CSoutput.n52 CSoutput.n51 165.8
R21712 CSoutput.n50 CSoutput.n8 165.8
R21713 CSoutput.n48 CSoutput.n47 165.8
R21714 CSoutput.n46 CSoutput.n9 165.8
R21715 CSoutput.n45 CSoutput.n44 165.8
R21716 CSoutput.n42 CSoutput.n10 165.8
R21717 CSoutput.n41 CSoutput.n40 165.8
R21718 CSoutput.n39 CSoutput.n38 165.8
R21719 CSoutput.n37 CSoutput.n12 165.8
R21720 CSoutput.n35 CSoutput.n34 165.8
R21721 CSoutput.n33 CSoutput.n13 165.8
R21722 CSoutput.n32 CSoutput.n31 165.8
R21723 CSoutput.n29 CSoutput.n14 165.8
R21724 CSoutput.n28 CSoutput.n27 165.8
R21725 CSoutput.n26 CSoutput.n25 165.8
R21726 CSoutput.n24 CSoutput.n16 165.8
R21727 CSoutput.n22 CSoutput.n21 165.8
R21728 CSoutput.n20 CSoutput.n17 165.8
R21729 CSoutput.n77 CSoutput.t194 162.194
R21730 CSoutput.n18 CSoutput.t201 120.501
R21731 CSoutput.n23 CSoutput.t203 120.501
R21732 CSoutput.n15 CSoutput.t196 120.501
R21733 CSoutput.n30 CSoutput.t213 120.501
R21734 CSoutput.n36 CSoutput.t204 120.501
R21735 CSoutput.n11 CSoutput.t199 120.501
R21736 CSoutput.n43 CSoutput.t193 120.501
R21737 CSoutput.n49 CSoutput.t210 120.501
R21738 CSoutput.n7 CSoutput.t207 120.501
R21739 CSoutput.n56 CSoutput.t197 120.501
R21740 CSoutput.n62 CSoutput.t212 120.501
R21741 CSoutput.n64 CSoutput.t208 120.501
R21742 CSoutput.n70 CSoutput.t200 120.501
R21743 CSoutput.n1 CSoutput.t202 120.501
R21744 CSoutput.n330 CSoutput.n328 103.469
R21745 CSoutput.n310 CSoutput.n308 103.469
R21746 CSoutput.n291 CSoutput.n289 103.469
R21747 CSoutput.n120 CSoutput.n118 103.469
R21748 CSoutput.n100 CSoutput.n98 103.469
R21749 CSoutput.n81 CSoutput.n79 103.469
R21750 CSoutput.n344 CSoutput.n343 103.111
R21751 CSoutput.n342 CSoutput.n341 103.111
R21752 CSoutput.n340 CSoutput.n339 103.111
R21753 CSoutput.n338 CSoutput.n337 103.111
R21754 CSoutput.n336 CSoutput.n335 103.111
R21755 CSoutput.n334 CSoutput.n333 103.111
R21756 CSoutput.n332 CSoutput.n331 103.111
R21757 CSoutput.n330 CSoutput.n329 103.111
R21758 CSoutput.n326 CSoutput.n325 103.111
R21759 CSoutput.n324 CSoutput.n323 103.111
R21760 CSoutput.n322 CSoutput.n321 103.111
R21761 CSoutput.n320 CSoutput.n319 103.111
R21762 CSoutput.n318 CSoutput.n317 103.111
R21763 CSoutput.n316 CSoutput.n315 103.111
R21764 CSoutput.n314 CSoutput.n313 103.111
R21765 CSoutput.n312 CSoutput.n311 103.111
R21766 CSoutput.n310 CSoutput.n309 103.111
R21767 CSoutput.n307 CSoutput.n306 103.111
R21768 CSoutput.n305 CSoutput.n304 103.111
R21769 CSoutput.n303 CSoutput.n302 103.111
R21770 CSoutput.n301 CSoutput.n300 103.111
R21771 CSoutput.n299 CSoutput.n298 103.111
R21772 CSoutput.n297 CSoutput.n296 103.111
R21773 CSoutput.n295 CSoutput.n294 103.111
R21774 CSoutput.n293 CSoutput.n292 103.111
R21775 CSoutput.n291 CSoutput.n290 103.111
R21776 CSoutput.n120 CSoutput.n119 103.111
R21777 CSoutput.n122 CSoutput.n121 103.111
R21778 CSoutput.n124 CSoutput.n123 103.111
R21779 CSoutput.n126 CSoutput.n125 103.111
R21780 CSoutput.n128 CSoutput.n127 103.111
R21781 CSoutput.n130 CSoutput.n129 103.111
R21782 CSoutput.n132 CSoutput.n131 103.111
R21783 CSoutput.n134 CSoutput.n133 103.111
R21784 CSoutput.n136 CSoutput.n135 103.111
R21785 CSoutput.n100 CSoutput.n99 103.111
R21786 CSoutput.n102 CSoutput.n101 103.111
R21787 CSoutput.n104 CSoutput.n103 103.111
R21788 CSoutput.n106 CSoutput.n105 103.111
R21789 CSoutput.n108 CSoutput.n107 103.111
R21790 CSoutput.n110 CSoutput.n109 103.111
R21791 CSoutput.n112 CSoutput.n111 103.111
R21792 CSoutput.n114 CSoutput.n113 103.111
R21793 CSoutput.n116 CSoutput.n115 103.111
R21794 CSoutput.n81 CSoutput.n80 103.111
R21795 CSoutput.n83 CSoutput.n82 103.111
R21796 CSoutput.n85 CSoutput.n84 103.111
R21797 CSoutput.n87 CSoutput.n86 103.111
R21798 CSoutput.n89 CSoutput.n88 103.111
R21799 CSoutput.n91 CSoutput.n90 103.111
R21800 CSoutput.n93 CSoutput.n92 103.111
R21801 CSoutput.n95 CSoutput.n94 103.111
R21802 CSoutput.n97 CSoutput.n96 103.111
R21803 CSoutput.n346 CSoutput.n345 103.111
R21804 CSoutput.n374 CSoutput.n372 81.5057
R21805 CSoutput.n362 CSoutput.n360 81.5057
R21806 CSoutput.n351 CSoutput.n349 81.5057
R21807 CSoutput.n410 CSoutput.n408 81.5057
R21808 CSoutput.n398 CSoutput.n396 81.5057
R21809 CSoutput.n387 CSoutput.n385 81.5057
R21810 CSoutput.n382 CSoutput.n381 80.9324
R21811 CSoutput.n380 CSoutput.n379 80.9324
R21812 CSoutput.n378 CSoutput.n377 80.9324
R21813 CSoutput.n376 CSoutput.n375 80.9324
R21814 CSoutput.n374 CSoutput.n373 80.9324
R21815 CSoutput.n370 CSoutput.n369 80.9324
R21816 CSoutput.n368 CSoutput.n367 80.9324
R21817 CSoutput.n366 CSoutput.n365 80.9324
R21818 CSoutput.n364 CSoutput.n363 80.9324
R21819 CSoutput.n362 CSoutput.n361 80.9324
R21820 CSoutput.n359 CSoutput.n358 80.9324
R21821 CSoutput.n357 CSoutput.n356 80.9324
R21822 CSoutput.n355 CSoutput.n354 80.9324
R21823 CSoutput.n353 CSoutput.n352 80.9324
R21824 CSoutput.n351 CSoutput.n350 80.9324
R21825 CSoutput.n410 CSoutput.n409 80.9324
R21826 CSoutput.n412 CSoutput.n411 80.9324
R21827 CSoutput.n414 CSoutput.n413 80.9324
R21828 CSoutput.n416 CSoutput.n415 80.9324
R21829 CSoutput.n418 CSoutput.n417 80.9324
R21830 CSoutput.n398 CSoutput.n397 80.9324
R21831 CSoutput.n400 CSoutput.n399 80.9324
R21832 CSoutput.n402 CSoutput.n401 80.9324
R21833 CSoutput.n404 CSoutput.n403 80.9324
R21834 CSoutput.n406 CSoutput.n405 80.9324
R21835 CSoutput.n387 CSoutput.n386 80.9324
R21836 CSoutput.n389 CSoutput.n388 80.9324
R21837 CSoutput.n391 CSoutput.n390 80.9324
R21838 CSoutput.n393 CSoutput.n392 80.9324
R21839 CSoutput.n395 CSoutput.n394 80.9324
R21840 CSoutput.n25 CSoutput.n24 48.1486
R21841 CSoutput.n69 CSoutput.n3 48.1486
R21842 CSoutput.n38 CSoutput.n37 48.1486
R21843 CSoutput.n42 CSoutput.n41 48.1486
R21844 CSoutput.n51 CSoutput.n50 48.1486
R21845 CSoutput.n55 CSoutput.n54 48.1486
R21846 CSoutput.n22 CSoutput.n17 46.462
R21847 CSoutput.n72 CSoutput.n71 46.462
R21848 CSoutput.n20 CSoutput.n19 44.9055
R21849 CSoutput.n29 CSoutput.n28 43.7635
R21850 CSoutput.n65 CSoutput.n63 43.7635
R21851 CSoutput.n35 CSoutput.n13 41.7396
R21852 CSoutput.n57 CSoutput.n5 41.7396
R21853 CSoutput.n44 CSoutput.n9 37.0171
R21854 CSoutput.n48 CSoutput.n9 37.0171
R21855 CSoutput.n76 CSoutput.n75 34.9932
R21856 CSoutput.n31 CSoutput.n13 32.2947
R21857 CSoutput.n61 CSoutput.n5 32.2947
R21858 CSoutput.n30 CSoutput.n29 29.6014
R21859 CSoutput.n63 CSoutput.n62 29.6014
R21860 CSoutput.n19 CSoutput.n18 28.4085
R21861 CSoutput.n18 CSoutput.n17 25.1176
R21862 CSoutput.n72 CSoutput.n1 25.1176
R21863 CSoutput.n43 CSoutput.n42 22.0922
R21864 CSoutput.n50 CSoutput.n49 22.0922
R21865 CSoutput.n77 CSoutput.n76 21.8586
R21866 CSoutput.n37 CSoutput.n36 18.9681
R21867 CSoutput.n56 CSoutput.n55 18.9681
R21868 CSoutput.n25 CSoutput.n15 17.6292
R21869 CSoutput.n64 CSoutput.n3 17.6292
R21870 CSoutput.n24 CSoutput.n23 15.844
R21871 CSoutput.n70 CSoutput.n69 15.844
R21872 CSoutput.n38 CSoutput.n11 14.5051
R21873 CSoutput.n54 CSoutput.n7 14.5051
R21874 CSoutput.n421 CSoutput.n78 11.4967
R21875 CSoutput.n41 CSoutput.n11 11.3811
R21876 CSoutput.n51 CSoutput.n7 11.3811
R21877 CSoutput.n23 CSoutput.n22 10.0422
R21878 CSoutput.n71 CSoutput.n70 10.0422
R21879 CSoutput.n327 CSoutput.n307 9.25285
R21880 CSoutput.n117 CSoutput.n97 9.25285
R21881 CSoutput.n371 CSoutput.n359 8.98182
R21882 CSoutput.n407 CSoutput.n395 8.98182
R21883 CSoutput.n384 CSoutput.n348 8.71742
R21884 CSoutput.n28 CSoutput.n15 8.25698
R21885 CSoutput.n65 CSoutput.n64 8.25698
R21886 CSoutput.n348 CSoutput.n347 7.12641
R21887 CSoutput.n138 CSoutput.n137 7.12641
R21888 CSoutput.n36 CSoutput.n35 6.91809
R21889 CSoutput.n57 CSoutput.n56 6.91809
R21890 CSoutput.n384 CSoutput.n383 6.02792
R21891 CSoutput.n420 CSoutput.n419 6.02792
R21892 CSoutput.n383 CSoutput.n382 5.25266
R21893 CSoutput.n371 CSoutput.n370 5.25266
R21894 CSoutput.n419 CSoutput.n418 5.25266
R21895 CSoutput.n407 CSoutput.n406 5.25266
R21896 CSoutput.n347 CSoutput.n346 5.1449
R21897 CSoutput.n327 CSoutput.n326 5.1449
R21898 CSoutput.n137 CSoutput.n136 5.1449
R21899 CSoutput.n117 CSoutput.n116 5.1449
R21900 CSoutput.n421 CSoutput.n138 4.91834
R21901 CSoutput.n229 CSoutput.n182 4.5005
R21902 CSoutput.n198 CSoutput.n182 4.5005
R21903 CSoutput.n193 CSoutput.n177 4.5005
R21904 CSoutput.n193 CSoutput.n179 4.5005
R21905 CSoutput.n193 CSoutput.n176 4.5005
R21906 CSoutput.n193 CSoutput.n180 4.5005
R21907 CSoutput.n193 CSoutput.n175 4.5005
R21908 CSoutput.n193 CSoutput.t198 4.5005
R21909 CSoutput.n193 CSoutput.n174 4.5005
R21910 CSoutput.n193 CSoutput.n181 4.5005
R21911 CSoutput.n193 CSoutput.n182 4.5005
R21912 CSoutput.n191 CSoutput.n177 4.5005
R21913 CSoutput.n191 CSoutput.n179 4.5005
R21914 CSoutput.n191 CSoutput.n176 4.5005
R21915 CSoutput.n191 CSoutput.n180 4.5005
R21916 CSoutput.n191 CSoutput.n175 4.5005
R21917 CSoutput.n191 CSoutput.t198 4.5005
R21918 CSoutput.n191 CSoutput.n174 4.5005
R21919 CSoutput.n191 CSoutput.n181 4.5005
R21920 CSoutput.n191 CSoutput.n182 4.5005
R21921 CSoutput.n190 CSoutput.n177 4.5005
R21922 CSoutput.n190 CSoutput.n179 4.5005
R21923 CSoutput.n190 CSoutput.n176 4.5005
R21924 CSoutput.n190 CSoutput.n180 4.5005
R21925 CSoutput.n190 CSoutput.n175 4.5005
R21926 CSoutput.n190 CSoutput.t198 4.5005
R21927 CSoutput.n190 CSoutput.n174 4.5005
R21928 CSoutput.n190 CSoutput.n181 4.5005
R21929 CSoutput.n190 CSoutput.n182 4.5005
R21930 CSoutput.n275 CSoutput.n177 4.5005
R21931 CSoutput.n275 CSoutput.n179 4.5005
R21932 CSoutput.n275 CSoutput.n176 4.5005
R21933 CSoutput.n275 CSoutput.n180 4.5005
R21934 CSoutput.n275 CSoutput.n175 4.5005
R21935 CSoutput.n275 CSoutput.t198 4.5005
R21936 CSoutput.n275 CSoutput.n174 4.5005
R21937 CSoutput.n275 CSoutput.n181 4.5005
R21938 CSoutput.n275 CSoutput.n182 4.5005
R21939 CSoutput.n273 CSoutput.n177 4.5005
R21940 CSoutput.n273 CSoutput.n179 4.5005
R21941 CSoutput.n273 CSoutput.n176 4.5005
R21942 CSoutput.n273 CSoutput.n180 4.5005
R21943 CSoutput.n273 CSoutput.n175 4.5005
R21944 CSoutput.n273 CSoutput.t198 4.5005
R21945 CSoutput.n273 CSoutput.n174 4.5005
R21946 CSoutput.n273 CSoutput.n181 4.5005
R21947 CSoutput.n271 CSoutput.n177 4.5005
R21948 CSoutput.n271 CSoutput.n179 4.5005
R21949 CSoutput.n271 CSoutput.n176 4.5005
R21950 CSoutput.n271 CSoutput.n180 4.5005
R21951 CSoutput.n271 CSoutput.n175 4.5005
R21952 CSoutput.n271 CSoutput.t198 4.5005
R21953 CSoutput.n271 CSoutput.n174 4.5005
R21954 CSoutput.n271 CSoutput.n181 4.5005
R21955 CSoutput.n201 CSoutput.n177 4.5005
R21956 CSoutput.n201 CSoutput.n179 4.5005
R21957 CSoutput.n201 CSoutput.n176 4.5005
R21958 CSoutput.n201 CSoutput.n180 4.5005
R21959 CSoutput.n201 CSoutput.n175 4.5005
R21960 CSoutput.n201 CSoutput.t198 4.5005
R21961 CSoutput.n201 CSoutput.n174 4.5005
R21962 CSoutput.n201 CSoutput.n181 4.5005
R21963 CSoutput.n201 CSoutput.n182 4.5005
R21964 CSoutput.n200 CSoutput.n177 4.5005
R21965 CSoutput.n200 CSoutput.n179 4.5005
R21966 CSoutput.n200 CSoutput.n176 4.5005
R21967 CSoutput.n200 CSoutput.n180 4.5005
R21968 CSoutput.n200 CSoutput.n175 4.5005
R21969 CSoutput.n200 CSoutput.t198 4.5005
R21970 CSoutput.n200 CSoutput.n174 4.5005
R21971 CSoutput.n200 CSoutput.n181 4.5005
R21972 CSoutput.n200 CSoutput.n182 4.5005
R21973 CSoutput.n204 CSoutput.n177 4.5005
R21974 CSoutput.n204 CSoutput.n179 4.5005
R21975 CSoutput.n204 CSoutput.n176 4.5005
R21976 CSoutput.n204 CSoutput.n180 4.5005
R21977 CSoutput.n204 CSoutput.n175 4.5005
R21978 CSoutput.n204 CSoutput.t198 4.5005
R21979 CSoutput.n204 CSoutput.n174 4.5005
R21980 CSoutput.n204 CSoutput.n181 4.5005
R21981 CSoutput.n204 CSoutput.n182 4.5005
R21982 CSoutput.n203 CSoutput.n177 4.5005
R21983 CSoutput.n203 CSoutput.n179 4.5005
R21984 CSoutput.n203 CSoutput.n176 4.5005
R21985 CSoutput.n203 CSoutput.n180 4.5005
R21986 CSoutput.n203 CSoutput.n175 4.5005
R21987 CSoutput.n203 CSoutput.t198 4.5005
R21988 CSoutput.n203 CSoutput.n174 4.5005
R21989 CSoutput.n203 CSoutput.n181 4.5005
R21990 CSoutput.n203 CSoutput.n182 4.5005
R21991 CSoutput.n186 CSoutput.n177 4.5005
R21992 CSoutput.n186 CSoutput.n179 4.5005
R21993 CSoutput.n186 CSoutput.n176 4.5005
R21994 CSoutput.n186 CSoutput.n180 4.5005
R21995 CSoutput.n186 CSoutput.n175 4.5005
R21996 CSoutput.n186 CSoutput.t198 4.5005
R21997 CSoutput.n186 CSoutput.n174 4.5005
R21998 CSoutput.n186 CSoutput.n181 4.5005
R21999 CSoutput.n186 CSoutput.n182 4.5005
R22000 CSoutput.n278 CSoutput.n177 4.5005
R22001 CSoutput.n278 CSoutput.n179 4.5005
R22002 CSoutput.n278 CSoutput.n176 4.5005
R22003 CSoutput.n278 CSoutput.n180 4.5005
R22004 CSoutput.n278 CSoutput.n175 4.5005
R22005 CSoutput.n278 CSoutput.t198 4.5005
R22006 CSoutput.n278 CSoutput.n174 4.5005
R22007 CSoutput.n278 CSoutput.n181 4.5005
R22008 CSoutput.n278 CSoutput.n182 4.5005
R22009 CSoutput.n265 CSoutput.n236 4.5005
R22010 CSoutput.n265 CSoutput.n242 4.5005
R22011 CSoutput.n223 CSoutput.n212 4.5005
R22012 CSoutput.n223 CSoutput.n214 4.5005
R22013 CSoutput.n223 CSoutput.n211 4.5005
R22014 CSoutput.n223 CSoutput.n215 4.5005
R22015 CSoutput.n223 CSoutput.n210 4.5005
R22016 CSoutput.n223 CSoutput.t206 4.5005
R22017 CSoutput.n223 CSoutput.n209 4.5005
R22018 CSoutput.n223 CSoutput.n216 4.5005
R22019 CSoutput.n265 CSoutput.n223 4.5005
R22020 CSoutput.n244 CSoutput.n212 4.5005
R22021 CSoutput.n244 CSoutput.n214 4.5005
R22022 CSoutput.n244 CSoutput.n211 4.5005
R22023 CSoutput.n244 CSoutput.n215 4.5005
R22024 CSoutput.n244 CSoutput.n210 4.5005
R22025 CSoutput.n244 CSoutput.t206 4.5005
R22026 CSoutput.n244 CSoutput.n209 4.5005
R22027 CSoutput.n244 CSoutput.n216 4.5005
R22028 CSoutput.n265 CSoutput.n244 4.5005
R22029 CSoutput.n222 CSoutput.n212 4.5005
R22030 CSoutput.n222 CSoutput.n214 4.5005
R22031 CSoutput.n222 CSoutput.n211 4.5005
R22032 CSoutput.n222 CSoutput.n215 4.5005
R22033 CSoutput.n222 CSoutput.n210 4.5005
R22034 CSoutput.n222 CSoutput.t206 4.5005
R22035 CSoutput.n222 CSoutput.n209 4.5005
R22036 CSoutput.n222 CSoutput.n216 4.5005
R22037 CSoutput.n265 CSoutput.n222 4.5005
R22038 CSoutput.n246 CSoutput.n212 4.5005
R22039 CSoutput.n246 CSoutput.n214 4.5005
R22040 CSoutput.n246 CSoutput.n211 4.5005
R22041 CSoutput.n246 CSoutput.n215 4.5005
R22042 CSoutput.n246 CSoutput.n210 4.5005
R22043 CSoutput.n246 CSoutput.t206 4.5005
R22044 CSoutput.n246 CSoutput.n209 4.5005
R22045 CSoutput.n246 CSoutput.n216 4.5005
R22046 CSoutput.n265 CSoutput.n246 4.5005
R22047 CSoutput.n212 CSoutput.n207 4.5005
R22048 CSoutput.n214 CSoutput.n207 4.5005
R22049 CSoutput.n211 CSoutput.n207 4.5005
R22050 CSoutput.n215 CSoutput.n207 4.5005
R22051 CSoutput.n210 CSoutput.n207 4.5005
R22052 CSoutput.t206 CSoutput.n207 4.5005
R22053 CSoutput.n209 CSoutput.n207 4.5005
R22054 CSoutput.n216 CSoutput.n207 4.5005
R22055 CSoutput.n268 CSoutput.n212 4.5005
R22056 CSoutput.n268 CSoutput.n214 4.5005
R22057 CSoutput.n268 CSoutput.n211 4.5005
R22058 CSoutput.n268 CSoutput.n215 4.5005
R22059 CSoutput.n268 CSoutput.n210 4.5005
R22060 CSoutput.n268 CSoutput.t206 4.5005
R22061 CSoutput.n268 CSoutput.n209 4.5005
R22062 CSoutput.n268 CSoutput.n216 4.5005
R22063 CSoutput.n266 CSoutput.n212 4.5005
R22064 CSoutput.n266 CSoutput.n214 4.5005
R22065 CSoutput.n266 CSoutput.n211 4.5005
R22066 CSoutput.n266 CSoutput.n215 4.5005
R22067 CSoutput.n266 CSoutput.n210 4.5005
R22068 CSoutput.n266 CSoutput.t206 4.5005
R22069 CSoutput.n266 CSoutput.n209 4.5005
R22070 CSoutput.n266 CSoutput.n216 4.5005
R22071 CSoutput.n266 CSoutput.n265 4.5005
R22072 CSoutput.n248 CSoutput.n212 4.5005
R22073 CSoutput.n248 CSoutput.n214 4.5005
R22074 CSoutput.n248 CSoutput.n211 4.5005
R22075 CSoutput.n248 CSoutput.n215 4.5005
R22076 CSoutput.n248 CSoutput.n210 4.5005
R22077 CSoutput.n248 CSoutput.t206 4.5005
R22078 CSoutput.n248 CSoutput.n209 4.5005
R22079 CSoutput.n248 CSoutput.n216 4.5005
R22080 CSoutput.n265 CSoutput.n248 4.5005
R22081 CSoutput.n220 CSoutput.n212 4.5005
R22082 CSoutput.n220 CSoutput.n214 4.5005
R22083 CSoutput.n220 CSoutput.n211 4.5005
R22084 CSoutput.n220 CSoutput.n215 4.5005
R22085 CSoutput.n220 CSoutput.n210 4.5005
R22086 CSoutput.n220 CSoutput.t206 4.5005
R22087 CSoutput.n220 CSoutput.n209 4.5005
R22088 CSoutput.n220 CSoutput.n216 4.5005
R22089 CSoutput.n265 CSoutput.n220 4.5005
R22090 CSoutput.n250 CSoutput.n212 4.5005
R22091 CSoutput.n250 CSoutput.n214 4.5005
R22092 CSoutput.n250 CSoutput.n211 4.5005
R22093 CSoutput.n250 CSoutput.n215 4.5005
R22094 CSoutput.n250 CSoutput.n210 4.5005
R22095 CSoutput.n250 CSoutput.t206 4.5005
R22096 CSoutput.n250 CSoutput.n209 4.5005
R22097 CSoutput.n250 CSoutput.n216 4.5005
R22098 CSoutput.n265 CSoutput.n250 4.5005
R22099 CSoutput.n219 CSoutput.n212 4.5005
R22100 CSoutput.n219 CSoutput.n214 4.5005
R22101 CSoutput.n219 CSoutput.n211 4.5005
R22102 CSoutput.n219 CSoutput.n215 4.5005
R22103 CSoutput.n219 CSoutput.n210 4.5005
R22104 CSoutput.n219 CSoutput.t206 4.5005
R22105 CSoutput.n219 CSoutput.n209 4.5005
R22106 CSoutput.n219 CSoutput.n216 4.5005
R22107 CSoutput.n265 CSoutput.n219 4.5005
R22108 CSoutput.n264 CSoutput.n212 4.5005
R22109 CSoutput.n264 CSoutput.n214 4.5005
R22110 CSoutput.n264 CSoutput.n211 4.5005
R22111 CSoutput.n264 CSoutput.n215 4.5005
R22112 CSoutput.n264 CSoutput.n210 4.5005
R22113 CSoutput.n264 CSoutput.t206 4.5005
R22114 CSoutput.n264 CSoutput.n209 4.5005
R22115 CSoutput.n264 CSoutput.n216 4.5005
R22116 CSoutput.n265 CSoutput.n264 4.5005
R22117 CSoutput.n263 CSoutput.n148 4.5005
R22118 CSoutput.n164 CSoutput.n148 4.5005
R22119 CSoutput.n159 CSoutput.n143 4.5005
R22120 CSoutput.n159 CSoutput.n145 4.5005
R22121 CSoutput.n159 CSoutput.n142 4.5005
R22122 CSoutput.n159 CSoutput.n146 4.5005
R22123 CSoutput.n159 CSoutput.n141 4.5005
R22124 CSoutput.n159 CSoutput.t209 4.5005
R22125 CSoutput.n159 CSoutput.n140 4.5005
R22126 CSoutput.n159 CSoutput.n147 4.5005
R22127 CSoutput.n159 CSoutput.n148 4.5005
R22128 CSoutput.n157 CSoutput.n143 4.5005
R22129 CSoutput.n157 CSoutput.n145 4.5005
R22130 CSoutput.n157 CSoutput.n142 4.5005
R22131 CSoutput.n157 CSoutput.n146 4.5005
R22132 CSoutput.n157 CSoutput.n141 4.5005
R22133 CSoutput.n157 CSoutput.t209 4.5005
R22134 CSoutput.n157 CSoutput.n140 4.5005
R22135 CSoutput.n157 CSoutput.n147 4.5005
R22136 CSoutput.n157 CSoutput.n148 4.5005
R22137 CSoutput.n156 CSoutput.n143 4.5005
R22138 CSoutput.n156 CSoutput.n145 4.5005
R22139 CSoutput.n156 CSoutput.n142 4.5005
R22140 CSoutput.n156 CSoutput.n146 4.5005
R22141 CSoutput.n156 CSoutput.n141 4.5005
R22142 CSoutput.n156 CSoutput.t209 4.5005
R22143 CSoutput.n156 CSoutput.n140 4.5005
R22144 CSoutput.n156 CSoutput.n147 4.5005
R22145 CSoutput.n156 CSoutput.n148 4.5005
R22146 CSoutput.n285 CSoutput.n143 4.5005
R22147 CSoutput.n285 CSoutput.n145 4.5005
R22148 CSoutput.n285 CSoutput.n142 4.5005
R22149 CSoutput.n285 CSoutput.n146 4.5005
R22150 CSoutput.n285 CSoutput.n141 4.5005
R22151 CSoutput.n285 CSoutput.t209 4.5005
R22152 CSoutput.n285 CSoutput.n140 4.5005
R22153 CSoutput.n285 CSoutput.n147 4.5005
R22154 CSoutput.n285 CSoutput.n148 4.5005
R22155 CSoutput.n283 CSoutput.n143 4.5005
R22156 CSoutput.n283 CSoutput.n145 4.5005
R22157 CSoutput.n283 CSoutput.n142 4.5005
R22158 CSoutput.n283 CSoutput.n146 4.5005
R22159 CSoutput.n283 CSoutput.n141 4.5005
R22160 CSoutput.n283 CSoutput.t209 4.5005
R22161 CSoutput.n283 CSoutput.n140 4.5005
R22162 CSoutput.n283 CSoutput.n147 4.5005
R22163 CSoutput.n281 CSoutput.n143 4.5005
R22164 CSoutput.n281 CSoutput.n145 4.5005
R22165 CSoutput.n281 CSoutput.n142 4.5005
R22166 CSoutput.n281 CSoutput.n146 4.5005
R22167 CSoutput.n281 CSoutput.n141 4.5005
R22168 CSoutput.n281 CSoutput.t209 4.5005
R22169 CSoutput.n281 CSoutput.n140 4.5005
R22170 CSoutput.n281 CSoutput.n147 4.5005
R22171 CSoutput.n167 CSoutput.n143 4.5005
R22172 CSoutput.n167 CSoutput.n145 4.5005
R22173 CSoutput.n167 CSoutput.n142 4.5005
R22174 CSoutput.n167 CSoutput.n146 4.5005
R22175 CSoutput.n167 CSoutput.n141 4.5005
R22176 CSoutput.n167 CSoutput.t209 4.5005
R22177 CSoutput.n167 CSoutput.n140 4.5005
R22178 CSoutput.n167 CSoutput.n147 4.5005
R22179 CSoutput.n167 CSoutput.n148 4.5005
R22180 CSoutput.n166 CSoutput.n143 4.5005
R22181 CSoutput.n166 CSoutput.n145 4.5005
R22182 CSoutput.n166 CSoutput.n142 4.5005
R22183 CSoutput.n166 CSoutput.n146 4.5005
R22184 CSoutput.n166 CSoutput.n141 4.5005
R22185 CSoutput.n166 CSoutput.t209 4.5005
R22186 CSoutput.n166 CSoutput.n140 4.5005
R22187 CSoutput.n166 CSoutput.n147 4.5005
R22188 CSoutput.n166 CSoutput.n148 4.5005
R22189 CSoutput.n170 CSoutput.n143 4.5005
R22190 CSoutput.n170 CSoutput.n145 4.5005
R22191 CSoutput.n170 CSoutput.n142 4.5005
R22192 CSoutput.n170 CSoutput.n146 4.5005
R22193 CSoutput.n170 CSoutput.n141 4.5005
R22194 CSoutput.n170 CSoutput.t209 4.5005
R22195 CSoutput.n170 CSoutput.n140 4.5005
R22196 CSoutput.n170 CSoutput.n147 4.5005
R22197 CSoutput.n170 CSoutput.n148 4.5005
R22198 CSoutput.n169 CSoutput.n143 4.5005
R22199 CSoutput.n169 CSoutput.n145 4.5005
R22200 CSoutput.n169 CSoutput.n142 4.5005
R22201 CSoutput.n169 CSoutput.n146 4.5005
R22202 CSoutput.n169 CSoutput.n141 4.5005
R22203 CSoutput.n169 CSoutput.t209 4.5005
R22204 CSoutput.n169 CSoutput.n140 4.5005
R22205 CSoutput.n169 CSoutput.n147 4.5005
R22206 CSoutput.n169 CSoutput.n148 4.5005
R22207 CSoutput.n152 CSoutput.n143 4.5005
R22208 CSoutput.n152 CSoutput.n145 4.5005
R22209 CSoutput.n152 CSoutput.n142 4.5005
R22210 CSoutput.n152 CSoutput.n146 4.5005
R22211 CSoutput.n152 CSoutput.n141 4.5005
R22212 CSoutput.n152 CSoutput.t209 4.5005
R22213 CSoutput.n152 CSoutput.n140 4.5005
R22214 CSoutput.n152 CSoutput.n147 4.5005
R22215 CSoutput.n152 CSoutput.n148 4.5005
R22216 CSoutput.n288 CSoutput.n143 4.5005
R22217 CSoutput.n288 CSoutput.n145 4.5005
R22218 CSoutput.n288 CSoutput.n142 4.5005
R22219 CSoutput.n288 CSoutput.n146 4.5005
R22220 CSoutput.n288 CSoutput.n141 4.5005
R22221 CSoutput.n288 CSoutput.t209 4.5005
R22222 CSoutput.n288 CSoutput.n140 4.5005
R22223 CSoutput.n288 CSoutput.n147 4.5005
R22224 CSoutput.n288 CSoutput.n148 4.5005
R22225 CSoutput.n347 CSoutput.n327 4.10845
R22226 CSoutput.n137 CSoutput.n117 4.10845
R22227 CSoutput.n345 CSoutput.t183 4.06363
R22228 CSoutput.n345 CSoutput.t39 4.06363
R22229 CSoutput.n343 CSoutput.t85 4.06363
R22230 CSoutput.n343 CSoutput.t9 4.06363
R22231 CSoutput.n341 CSoutput.t52 4.06363
R22232 CSoutput.n341 CSoutput.t26 4.06363
R22233 CSoutput.n339 CSoutput.t79 4.06363
R22234 CSoutput.n339 CSoutput.t21 4.06363
R22235 CSoutput.n337 CSoutput.t23 4.06363
R22236 CSoutput.n337 CSoutput.t54 4.06363
R22237 CSoutput.n335 CSoutput.t80 4.06363
R22238 CSoutput.n335 CSoutput.t87 4.06363
R22239 CSoutput.n333 CSoutput.t29 4.06363
R22240 CSoutput.n333 CSoutput.t164 4.06363
R22241 CSoutput.n331 CSoutput.t8 4.06363
R22242 CSoutput.n331 CSoutput.t172 4.06363
R22243 CSoutput.n329 CSoutput.t35 4.06363
R22244 CSoutput.n329 CSoutput.t1 4.06363
R22245 CSoutput.n328 CSoutput.t53 4.06363
R22246 CSoutput.n328 CSoutput.t47 4.06363
R22247 CSoutput.n325 CSoutput.t83 4.06363
R22248 CSoutput.n325 CSoutput.t82 4.06363
R22249 CSoutput.n323 CSoutput.t34 4.06363
R22250 CSoutput.n323 CSoutput.t0 4.06363
R22251 CSoutput.n321 CSoutput.t91 4.06363
R22252 CSoutput.n321 CSoutput.t15 4.06363
R22253 CSoutput.n319 CSoutput.t11 4.06363
R22254 CSoutput.n319 CSoutput.t43 4.06363
R22255 CSoutput.n317 CSoutput.t60 4.06363
R22256 CSoutput.n317 CSoutput.t181 4.06363
R22257 CSoutput.n315 CSoutput.t167 4.06363
R22258 CSoutput.n315 CSoutput.t40 4.06363
R22259 CSoutput.n313 CSoutput.t19 4.06363
R22260 CSoutput.n313 CSoutput.t191 4.06363
R22261 CSoutput.n311 CSoutput.t69 4.06363
R22262 CSoutput.n311 CSoutput.t55 4.06363
R22263 CSoutput.n309 CSoutput.t14 4.06363
R22264 CSoutput.n309 CSoutput.t178 4.06363
R22265 CSoutput.n308 CSoutput.t90 4.06363
R22266 CSoutput.n308 CSoutput.t63 4.06363
R22267 CSoutput.n306 CSoutput.t66 4.06363
R22268 CSoutput.n306 CSoutput.t89 4.06363
R22269 CSoutput.n304 CSoutput.t72 4.06363
R22270 CSoutput.n304 CSoutput.t77 4.06363
R22271 CSoutput.n302 CSoutput.t46 4.06363
R22272 CSoutput.n302 CSoutput.t42 4.06363
R22273 CSoutput.n300 CSoutput.t6 4.06363
R22274 CSoutput.n300 CSoutput.t86 4.06363
R22275 CSoutput.n298 CSoutput.t190 4.06363
R22276 CSoutput.n298 CSoutput.t16 4.06363
R22277 CSoutput.n296 CSoutput.t67 4.06363
R22278 CSoutput.n296 CSoutput.t51 4.06363
R22279 CSoutput.n294 CSoutput.t22 4.06363
R22280 CSoutput.n294 CSoutput.t174 4.06363
R22281 CSoutput.n292 CSoutput.t45 4.06363
R22282 CSoutput.n292 CSoutput.t173 4.06363
R22283 CSoutput.n290 CSoutput.t68 4.06363
R22284 CSoutput.n290 CSoutput.t2 4.06363
R22285 CSoutput.n289 CSoutput.t18 4.06363
R22286 CSoutput.n289 CSoutput.t10 4.06363
R22287 CSoutput.n118 CSoutput.t36 4.06363
R22288 CSoutput.n118 CSoutput.t188 4.06363
R22289 CSoutput.n119 CSoutput.t48 4.06363
R22290 CSoutput.n119 CSoutput.t12 4.06363
R22291 CSoutput.n121 CSoutput.t32 4.06363
R22292 CSoutput.n121 CSoutput.t56 4.06363
R22293 CSoutput.n123 CSoutput.t49 4.06363
R22294 CSoutput.n123 CSoutput.t168 4.06363
R22295 CSoutput.n125 CSoutput.t64 4.06363
R22296 CSoutput.n125 CSoutput.t58 4.06363
R22297 CSoutput.n127 CSoutput.t78 4.06363
R22298 CSoutput.n127 CSoutput.t3 4.06363
R22299 CSoutput.n129 CSoutput.t186 4.06363
R22300 CSoutput.n129 CSoutput.t88 4.06363
R22301 CSoutput.n131 CSoutput.t13 4.06363
R22302 CSoutput.n131 CSoutput.t175 4.06363
R22303 CSoutput.n133 CSoutput.t57 4.06363
R22304 CSoutput.n133 CSoutput.t166 4.06363
R22305 CSoutput.n135 CSoutput.t37 4.06363
R22306 CSoutput.n135 CSoutput.t33 4.06363
R22307 CSoutput.n98 CSoutput.t185 4.06363
R22308 CSoutput.n98 CSoutput.t31 4.06363
R22309 CSoutput.n99 CSoutput.t74 4.06363
R22310 CSoutput.n99 CSoutput.t177 4.06363
R22311 CSoutput.n101 CSoutput.t171 4.06363
R22312 CSoutput.n101 CSoutput.t38 4.06363
R22313 CSoutput.n103 CSoutput.t75 4.06363
R22314 CSoutput.n103 CSoutput.t81 4.06363
R22315 CSoutput.n105 CSoutput.t61 4.06363
R22316 CSoutput.n105 CSoutput.t189 4.06363
R22317 CSoutput.n107 CSoutput.t41 4.06363
R22318 CSoutput.n107 CSoutput.t73 4.06363
R22319 CSoutput.n109 CSoutput.t62 4.06363
R22320 CSoutput.n109 CSoutput.t20 4.06363
R22321 CSoutput.n111 CSoutput.t184 4.06363
R22322 CSoutput.n111 CSoutput.t30 4.06363
R22323 CSoutput.n113 CSoutput.t182 4.06363
R22324 CSoutput.n113 CSoutput.t70 4.06363
R22325 CSoutput.n115 CSoutput.t170 4.06363
R22326 CSoutput.n115 CSoutput.t4 4.06363
R22327 CSoutput.n79 CSoutput.t180 4.06363
R22328 CSoutput.n79 CSoutput.t5 4.06363
R22329 CSoutput.n80 CSoutput.t169 4.06363
R22330 CSoutput.n80 CSoutput.t7 4.06363
R22331 CSoutput.n82 CSoutput.t27 4.06363
R22332 CSoutput.n82 CSoutput.t44 4.06363
R22333 CSoutput.n84 CSoutput.t76 4.06363
R22334 CSoutput.n84 CSoutput.t176 4.06363
R22335 CSoutput.n86 CSoutput.t50 4.06363
R22336 CSoutput.n86 CSoutput.t25 4.06363
R22337 CSoutput.n88 CSoutput.t17 4.06363
R22338 CSoutput.n88 CSoutput.t179 4.06363
R22339 CSoutput.n90 CSoutput.t59 4.06363
R22340 CSoutput.n90 CSoutput.t71 4.06363
R22341 CSoutput.n92 CSoutput.t28 4.06363
R22342 CSoutput.n92 CSoutput.t187 4.06363
R22343 CSoutput.n94 CSoutput.t84 4.06363
R22344 CSoutput.n94 CSoutput.t165 4.06363
R22345 CSoutput.n96 CSoutput.t65 4.06363
R22346 CSoutput.n96 CSoutput.t24 4.06363
R22347 CSoutput.n44 CSoutput.n43 3.79402
R22348 CSoutput.n49 CSoutput.n48 3.79402
R22349 CSoutput.n421 CSoutput.n420 3.78008
R22350 CSoutput.n383 CSoutput.n371 3.72967
R22351 CSoutput.n419 CSoutput.n407 3.72967
R22352 CSoutput.n348 CSoutput.n138 3.19963
R22353 CSoutput.n381 CSoutput.t109 2.82907
R22354 CSoutput.n381 CSoutput.t113 2.82907
R22355 CSoutput.n379 CSoutput.t108 2.82907
R22356 CSoutput.n379 CSoutput.t163 2.82907
R22357 CSoutput.n377 CSoutput.t123 2.82907
R22358 CSoutput.n377 CSoutput.t103 2.82907
R22359 CSoutput.n375 CSoutput.t96 2.82907
R22360 CSoutput.n375 CSoutput.t143 2.82907
R22361 CSoutput.n373 CSoutput.t115 2.82907
R22362 CSoutput.n373 CSoutput.t118 2.82907
R22363 CSoutput.n372 CSoutput.t102 2.82907
R22364 CSoutput.n372 CSoutput.t154 2.82907
R22365 CSoutput.n369 CSoutput.t95 2.82907
R22366 CSoutput.n369 CSoutput.t141 2.82907
R22367 CSoutput.n367 CSoutput.t140 2.82907
R22368 CSoutput.n367 CSoutput.t128 2.82907
R22369 CSoutput.n365 CSoutput.t152 2.82907
R22370 CSoutput.n365 CSoutput.t93 2.82907
R22371 CSoutput.n363 CSoutput.t94 2.82907
R22372 CSoutput.n363 CSoutput.t146 2.82907
R22373 CSoutput.n361 CSoutput.t101 2.82907
R22374 CSoutput.n361 CSoutput.t151 2.82907
R22375 CSoutput.n360 CSoutput.t157 2.82907
R22376 CSoutput.n360 CSoutput.t92 2.82907
R22377 CSoutput.n358 CSoutput.t131 2.82907
R22378 CSoutput.n358 CSoutput.t138 2.82907
R22379 CSoutput.n356 CSoutput.t124 2.82907
R22380 CSoutput.n356 CSoutput.t153 2.82907
R22381 CSoutput.n354 CSoutput.t134 2.82907
R22382 CSoutput.n354 CSoutput.t117 2.82907
R22383 CSoutput.n352 CSoutput.t110 2.82907
R22384 CSoutput.n352 CSoutput.t125 2.82907
R22385 CSoutput.n350 CSoutput.t116 2.82907
R22386 CSoutput.n350 CSoutput.t121 2.82907
R22387 CSoutput.n349 CSoutput.t122 2.82907
R22388 CSoutput.n349 CSoutput.t160 2.82907
R22389 CSoutput.n408 CSoutput.t130 2.82907
R22390 CSoutput.n408 CSoutput.t148 2.82907
R22391 CSoutput.n409 CSoutput.t111 2.82907
R22392 CSoutput.n409 CSoutput.t120 2.82907
R22393 CSoutput.n411 CSoutput.t126 2.82907
R22394 CSoutput.n411 CSoutput.t135 2.82907
R22395 CSoutput.n413 CSoutput.t149 2.82907
R22396 CSoutput.n413 CSoutput.t129 2.82907
R22397 CSoutput.n415 CSoutput.t133 2.82907
R22398 CSoutput.n415 CSoutput.t158 2.82907
R22399 CSoutput.n417 CSoutput.t98 2.82907
R22400 CSoutput.n417 CSoutput.t114 2.82907
R22401 CSoutput.n396 CSoutput.t104 2.82907
R22402 CSoutput.n396 CSoutput.t99 2.82907
R22403 CSoutput.n397 CSoutput.t97 2.82907
R22404 CSoutput.n397 CSoutput.t161 2.82907
R22405 CSoutput.n399 CSoutput.t162 2.82907
R22406 CSoutput.n399 CSoutput.t105 2.82907
R22407 CSoutput.n401 CSoutput.t106 2.82907
R22408 CSoutput.n401 CSoutput.t137 2.82907
R22409 CSoutput.n403 CSoutput.t136 2.82907
R22410 CSoutput.n403 CSoutput.t156 2.82907
R22411 CSoutput.n405 CSoutput.t159 2.82907
R22412 CSoutput.n405 CSoutput.t150 2.82907
R22413 CSoutput.n385 CSoutput.t112 2.82907
R22414 CSoutput.n385 CSoutput.t142 2.82907
R22415 CSoutput.n386 CSoutput.t139 2.82907
R22416 CSoutput.n386 CSoutput.t127 2.82907
R22417 CSoutput.n388 CSoutput.t145 2.82907
R22418 CSoutput.n388 CSoutput.t119 2.82907
R22419 CSoutput.n390 CSoutput.t132 2.82907
R22420 CSoutput.n390 CSoutput.t155 2.82907
R22421 CSoutput.n392 CSoutput.t107 2.82907
R22422 CSoutput.n392 CSoutput.t144 2.82907
R22423 CSoutput.n394 CSoutput.t100 2.82907
R22424 CSoutput.n394 CSoutput.t147 2.82907
R22425 CSoutput.n420 CSoutput.n384 2.75627
R22426 CSoutput.n75 CSoutput.n1 2.45513
R22427 CSoutput.n229 CSoutput.n227 2.251
R22428 CSoutput.n229 CSoutput.n226 2.251
R22429 CSoutput.n229 CSoutput.n225 2.251
R22430 CSoutput.n229 CSoutput.n224 2.251
R22431 CSoutput.n198 CSoutput.n197 2.251
R22432 CSoutput.n198 CSoutput.n196 2.251
R22433 CSoutput.n198 CSoutput.n195 2.251
R22434 CSoutput.n198 CSoutput.n194 2.251
R22435 CSoutput.n271 CSoutput.n270 2.251
R22436 CSoutput.n236 CSoutput.n234 2.251
R22437 CSoutput.n236 CSoutput.n233 2.251
R22438 CSoutput.n236 CSoutput.n232 2.251
R22439 CSoutput.n254 CSoutput.n236 2.251
R22440 CSoutput.n242 CSoutput.n241 2.251
R22441 CSoutput.n242 CSoutput.n240 2.251
R22442 CSoutput.n242 CSoutput.n239 2.251
R22443 CSoutput.n242 CSoutput.n238 2.251
R22444 CSoutput.n268 CSoutput.n208 2.251
R22445 CSoutput.n263 CSoutput.n261 2.251
R22446 CSoutput.n263 CSoutput.n260 2.251
R22447 CSoutput.n263 CSoutput.n259 2.251
R22448 CSoutput.n263 CSoutput.n258 2.251
R22449 CSoutput.n164 CSoutput.n163 2.251
R22450 CSoutput.n164 CSoutput.n162 2.251
R22451 CSoutput.n164 CSoutput.n161 2.251
R22452 CSoutput.n164 CSoutput.n160 2.251
R22453 CSoutput.n281 CSoutput.n280 2.251
R22454 CSoutput.n198 CSoutput.n178 2.2505
R22455 CSoutput.n193 CSoutput.n178 2.2505
R22456 CSoutput.n191 CSoutput.n178 2.2505
R22457 CSoutput.n190 CSoutput.n178 2.2505
R22458 CSoutput.n275 CSoutput.n178 2.2505
R22459 CSoutput.n273 CSoutput.n178 2.2505
R22460 CSoutput.n271 CSoutput.n178 2.2505
R22461 CSoutput.n201 CSoutput.n178 2.2505
R22462 CSoutput.n200 CSoutput.n178 2.2505
R22463 CSoutput.n204 CSoutput.n178 2.2505
R22464 CSoutput.n203 CSoutput.n178 2.2505
R22465 CSoutput.n186 CSoutput.n178 2.2505
R22466 CSoutput.n278 CSoutput.n178 2.2505
R22467 CSoutput.n278 CSoutput.n277 2.2505
R22468 CSoutput.n242 CSoutput.n213 2.2505
R22469 CSoutput.n223 CSoutput.n213 2.2505
R22470 CSoutput.n244 CSoutput.n213 2.2505
R22471 CSoutput.n222 CSoutput.n213 2.2505
R22472 CSoutput.n246 CSoutput.n213 2.2505
R22473 CSoutput.n213 CSoutput.n207 2.2505
R22474 CSoutput.n268 CSoutput.n213 2.2505
R22475 CSoutput.n266 CSoutput.n213 2.2505
R22476 CSoutput.n248 CSoutput.n213 2.2505
R22477 CSoutput.n220 CSoutput.n213 2.2505
R22478 CSoutput.n250 CSoutput.n213 2.2505
R22479 CSoutput.n219 CSoutput.n213 2.2505
R22480 CSoutput.n264 CSoutput.n213 2.2505
R22481 CSoutput.n264 CSoutput.n217 2.2505
R22482 CSoutput.n164 CSoutput.n144 2.2505
R22483 CSoutput.n159 CSoutput.n144 2.2505
R22484 CSoutput.n157 CSoutput.n144 2.2505
R22485 CSoutput.n156 CSoutput.n144 2.2505
R22486 CSoutput.n285 CSoutput.n144 2.2505
R22487 CSoutput.n283 CSoutput.n144 2.2505
R22488 CSoutput.n281 CSoutput.n144 2.2505
R22489 CSoutput.n167 CSoutput.n144 2.2505
R22490 CSoutput.n166 CSoutput.n144 2.2505
R22491 CSoutput.n170 CSoutput.n144 2.2505
R22492 CSoutput.n169 CSoutput.n144 2.2505
R22493 CSoutput.n152 CSoutput.n144 2.2505
R22494 CSoutput.n288 CSoutput.n144 2.2505
R22495 CSoutput.n288 CSoutput.n287 2.2505
R22496 CSoutput.n206 CSoutput.n199 2.25024
R22497 CSoutput.n206 CSoutput.n192 2.25024
R22498 CSoutput.n274 CSoutput.n206 2.25024
R22499 CSoutput.n206 CSoutput.n202 2.25024
R22500 CSoutput.n206 CSoutput.n205 2.25024
R22501 CSoutput.n206 CSoutput.n173 2.25024
R22502 CSoutput.n256 CSoutput.n253 2.25024
R22503 CSoutput.n256 CSoutput.n252 2.25024
R22504 CSoutput.n256 CSoutput.n251 2.25024
R22505 CSoutput.n256 CSoutput.n218 2.25024
R22506 CSoutput.n256 CSoutput.n255 2.25024
R22507 CSoutput.n257 CSoutput.n256 2.25024
R22508 CSoutput.n172 CSoutput.n165 2.25024
R22509 CSoutput.n172 CSoutput.n158 2.25024
R22510 CSoutput.n284 CSoutput.n172 2.25024
R22511 CSoutput.n172 CSoutput.n168 2.25024
R22512 CSoutput.n172 CSoutput.n171 2.25024
R22513 CSoutput.n172 CSoutput.n139 2.25024
R22514 CSoutput.n273 CSoutput.n183 1.50111
R22515 CSoutput.n221 CSoutput.n207 1.50111
R22516 CSoutput.n283 CSoutput.n149 1.50111
R22517 CSoutput.n229 CSoutput.n228 1.501
R22518 CSoutput.n236 CSoutput.n235 1.501
R22519 CSoutput.n263 CSoutput.n262 1.501
R22520 CSoutput.n277 CSoutput.n188 1.12536
R22521 CSoutput.n277 CSoutput.n189 1.12536
R22522 CSoutput.n277 CSoutput.n276 1.12536
R22523 CSoutput.n237 CSoutput.n217 1.12536
R22524 CSoutput.n243 CSoutput.n217 1.12536
R22525 CSoutput.n245 CSoutput.n217 1.12536
R22526 CSoutput.n287 CSoutput.n154 1.12536
R22527 CSoutput.n287 CSoutput.n155 1.12536
R22528 CSoutput.n287 CSoutput.n286 1.12536
R22529 CSoutput.n277 CSoutput.n184 1.12536
R22530 CSoutput.n277 CSoutput.n185 1.12536
R22531 CSoutput.n277 CSoutput.n187 1.12536
R22532 CSoutput.n267 CSoutput.n217 1.12536
R22533 CSoutput.n247 CSoutput.n217 1.12536
R22534 CSoutput.n249 CSoutput.n217 1.12536
R22535 CSoutput.n287 CSoutput.n150 1.12536
R22536 CSoutput.n287 CSoutput.n151 1.12536
R22537 CSoutput.n287 CSoutput.n153 1.12536
R22538 CSoutput.n31 CSoutput.n30 0.669944
R22539 CSoutput.n62 CSoutput.n61 0.669944
R22540 CSoutput.n376 CSoutput.n374 0.573776
R22541 CSoutput.n378 CSoutput.n376 0.573776
R22542 CSoutput.n380 CSoutput.n378 0.573776
R22543 CSoutput.n382 CSoutput.n380 0.573776
R22544 CSoutput.n364 CSoutput.n362 0.573776
R22545 CSoutput.n366 CSoutput.n364 0.573776
R22546 CSoutput.n368 CSoutput.n366 0.573776
R22547 CSoutput.n370 CSoutput.n368 0.573776
R22548 CSoutput.n353 CSoutput.n351 0.573776
R22549 CSoutput.n355 CSoutput.n353 0.573776
R22550 CSoutput.n357 CSoutput.n355 0.573776
R22551 CSoutput.n359 CSoutput.n357 0.573776
R22552 CSoutput.n418 CSoutput.n416 0.573776
R22553 CSoutput.n416 CSoutput.n414 0.573776
R22554 CSoutput.n414 CSoutput.n412 0.573776
R22555 CSoutput.n412 CSoutput.n410 0.573776
R22556 CSoutput.n406 CSoutput.n404 0.573776
R22557 CSoutput.n404 CSoutput.n402 0.573776
R22558 CSoutput.n402 CSoutput.n400 0.573776
R22559 CSoutput.n400 CSoutput.n398 0.573776
R22560 CSoutput.n395 CSoutput.n393 0.573776
R22561 CSoutput.n393 CSoutput.n391 0.573776
R22562 CSoutput.n391 CSoutput.n389 0.573776
R22563 CSoutput.n389 CSoutput.n387 0.573776
R22564 CSoutput.n421 CSoutput.n288 0.534303
R22565 CSoutput.n332 CSoutput.n330 0.358259
R22566 CSoutput.n334 CSoutput.n332 0.358259
R22567 CSoutput.n336 CSoutput.n334 0.358259
R22568 CSoutput.n338 CSoutput.n336 0.358259
R22569 CSoutput.n340 CSoutput.n338 0.358259
R22570 CSoutput.n342 CSoutput.n340 0.358259
R22571 CSoutput.n344 CSoutput.n342 0.358259
R22572 CSoutput.n346 CSoutput.n344 0.358259
R22573 CSoutput.n312 CSoutput.n310 0.358259
R22574 CSoutput.n314 CSoutput.n312 0.358259
R22575 CSoutput.n316 CSoutput.n314 0.358259
R22576 CSoutput.n318 CSoutput.n316 0.358259
R22577 CSoutput.n320 CSoutput.n318 0.358259
R22578 CSoutput.n322 CSoutput.n320 0.358259
R22579 CSoutput.n324 CSoutput.n322 0.358259
R22580 CSoutput.n326 CSoutput.n324 0.358259
R22581 CSoutput.n293 CSoutput.n291 0.358259
R22582 CSoutput.n295 CSoutput.n293 0.358259
R22583 CSoutput.n297 CSoutput.n295 0.358259
R22584 CSoutput.n299 CSoutput.n297 0.358259
R22585 CSoutput.n301 CSoutput.n299 0.358259
R22586 CSoutput.n303 CSoutput.n301 0.358259
R22587 CSoutput.n305 CSoutput.n303 0.358259
R22588 CSoutput.n307 CSoutput.n305 0.358259
R22589 CSoutput.n136 CSoutput.n134 0.358259
R22590 CSoutput.n134 CSoutput.n132 0.358259
R22591 CSoutput.n132 CSoutput.n130 0.358259
R22592 CSoutput.n130 CSoutput.n128 0.358259
R22593 CSoutput.n128 CSoutput.n126 0.358259
R22594 CSoutput.n126 CSoutput.n124 0.358259
R22595 CSoutput.n124 CSoutput.n122 0.358259
R22596 CSoutput.n122 CSoutput.n120 0.358259
R22597 CSoutput.n116 CSoutput.n114 0.358259
R22598 CSoutput.n114 CSoutput.n112 0.358259
R22599 CSoutput.n112 CSoutput.n110 0.358259
R22600 CSoutput.n110 CSoutput.n108 0.358259
R22601 CSoutput.n108 CSoutput.n106 0.358259
R22602 CSoutput.n106 CSoutput.n104 0.358259
R22603 CSoutput.n104 CSoutput.n102 0.358259
R22604 CSoutput.n102 CSoutput.n100 0.358259
R22605 CSoutput.n97 CSoutput.n95 0.358259
R22606 CSoutput.n95 CSoutput.n93 0.358259
R22607 CSoutput.n93 CSoutput.n91 0.358259
R22608 CSoutput.n91 CSoutput.n89 0.358259
R22609 CSoutput.n89 CSoutput.n87 0.358259
R22610 CSoutput.n87 CSoutput.n85 0.358259
R22611 CSoutput.n85 CSoutput.n83 0.358259
R22612 CSoutput.n83 CSoutput.n81 0.358259
R22613 CSoutput.n21 CSoutput.n20 0.169105
R22614 CSoutput.n21 CSoutput.n16 0.169105
R22615 CSoutput.n26 CSoutput.n16 0.169105
R22616 CSoutput.n27 CSoutput.n26 0.169105
R22617 CSoutput.n27 CSoutput.n14 0.169105
R22618 CSoutput.n32 CSoutput.n14 0.169105
R22619 CSoutput.n33 CSoutput.n32 0.169105
R22620 CSoutput.n34 CSoutput.n33 0.169105
R22621 CSoutput.n34 CSoutput.n12 0.169105
R22622 CSoutput.n39 CSoutput.n12 0.169105
R22623 CSoutput.n40 CSoutput.n39 0.169105
R22624 CSoutput.n40 CSoutput.n10 0.169105
R22625 CSoutput.n45 CSoutput.n10 0.169105
R22626 CSoutput.n46 CSoutput.n45 0.169105
R22627 CSoutput.n47 CSoutput.n46 0.169105
R22628 CSoutput.n47 CSoutput.n8 0.169105
R22629 CSoutput.n52 CSoutput.n8 0.169105
R22630 CSoutput.n53 CSoutput.n52 0.169105
R22631 CSoutput.n53 CSoutput.n6 0.169105
R22632 CSoutput.n58 CSoutput.n6 0.169105
R22633 CSoutput.n59 CSoutput.n58 0.169105
R22634 CSoutput.n60 CSoutput.n59 0.169105
R22635 CSoutput.n60 CSoutput.n4 0.169105
R22636 CSoutput.n66 CSoutput.n4 0.169105
R22637 CSoutput.n67 CSoutput.n66 0.169105
R22638 CSoutput.n68 CSoutput.n67 0.169105
R22639 CSoutput.n68 CSoutput.n2 0.169105
R22640 CSoutput.n73 CSoutput.n2 0.169105
R22641 CSoutput.n74 CSoutput.n73 0.169105
R22642 CSoutput.n74 CSoutput.n0 0.169105
R22643 CSoutput.n78 CSoutput.n0 0.169105
R22644 CSoutput.n231 CSoutput.n230 0.0910737
R22645 CSoutput.n282 CSoutput.n279 0.0723685
R22646 CSoutput.n236 CSoutput.n231 0.0522944
R22647 CSoutput.n279 CSoutput.n278 0.0499135
R22648 CSoutput.n230 CSoutput.n229 0.0499135
R22649 CSoutput.n264 CSoutput.n263 0.0464294
R22650 CSoutput.n272 CSoutput.n269 0.0391444
R22651 CSoutput.n231 CSoutput.t211 0.023435
R22652 CSoutput.n279 CSoutput.t195 0.02262
R22653 CSoutput.n230 CSoutput.t205 0.02262
R22654 CSoutput CSoutput.n421 0.0052
R22655 CSoutput.n201 CSoutput.n184 0.00365111
R22656 CSoutput.n204 CSoutput.n185 0.00365111
R22657 CSoutput.n187 CSoutput.n186 0.00365111
R22658 CSoutput.n229 CSoutput.n188 0.00365111
R22659 CSoutput.n193 CSoutput.n189 0.00365111
R22660 CSoutput.n276 CSoutput.n190 0.00365111
R22661 CSoutput.n267 CSoutput.n266 0.00365111
R22662 CSoutput.n247 CSoutput.n220 0.00365111
R22663 CSoutput.n249 CSoutput.n219 0.00365111
R22664 CSoutput.n237 CSoutput.n236 0.00365111
R22665 CSoutput.n243 CSoutput.n223 0.00365111
R22666 CSoutput.n245 CSoutput.n222 0.00365111
R22667 CSoutput.n167 CSoutput.n150 0.00365111
R22668 CSoutput.n170 CSoutput.n151 0.00365111
R22669 CSoutput.n153 CSoutput.n152 0.00365111
R22670 CSoutput.n263 CSoutput.n154 0.00365111
R22671 CSoutput.n159 CSoutput.n155 0.00365111
R22672 CSoutput.n286 CSoutput.n156 0.00365111
R22673 CSoutput.n198 CSoutput.n188 0.00340054
R22674 CSoutput.n191 CSoutput.n189 0.00340054
R22675 CSoutput.n276 CSoutput.n275 0.00340054
R22676 CSoutput.n271 CSoutput.n184 0.00340054
R22677 CSoutput.n200 CSoutput.n185 0.00340054
R22678 CSoutput.n203 CSoutput.n187 0.00340054
R22679 CSoutput.n242 CSoutput.n237 0.00340054
R22680 CSoutput.n244 CSoutput.n243 0.00340054
R22681 CSoutput.n246 CSoutput.n245 0.00340054
R22682 CSoutput.n268 CSoutput.n267 0.00340054
R22683 CSoutput.n248 CSoutput.n247 0.00340054
R22684 CSoutput.n250 CSoutput.n249 0.00340054
R22685 CSoutput.n164 CSoutput.n154 0.00340054
R22686 CSoutput.n157 CSoutput.n155 0.00340054
R22687 CSoutput.n286 CSoutput.n285 0.00340054
R22688 CSoutput.n281 CSoutput.n150 0.00340054
R22689 CSoutput.n166 CSoutput.n151 0.00340054
R22690 CSoutput.n169 CSoutput.n153 0.00340054
R22691 CSoutput.n199 CSoutput.n193 0.00252698
R22692 CSoutput.n192 CSoutput.n190 0.00252698
R22693 CSoutput.n274 CSoutput.n273 0.00252698
R22694 CSoutput.n202 CSoutput.n200 0.00252698
R22695 CSoutput.n205 CSoutput.n203 0.00252698
R22696 CSoutput.n278 CSoutput.n173 0.00252698
R22697 CSoutput.n199 CSoutput.n198 0.00252698
R22698 CSoutput.n192 CSoutput.n191 0.00252698
R22699 CSoutput.n275 CSoutput.n274 0.00252698
R22700 CSoutput.n202 CSoutput.n201 0.00252698
R22701 CSoutput.n205 CSoutput.n204 0.00252698
R22702 CSoutput.n186 CSoutput.n173 0.00252698
R22703 CSoutput.n253 CSoutput.n223 0.00252698
R22704 CSoutput.n252 CSoutput.n222 0.00252698
R22705 CSoutput.n251 CSoutput.n207 0.00252698
R22706 CSoutput.n248 CSoutput.n218 0.00252698
R22707 CSoutput.n255 CSoutput.n250 0.00252698
R22708 CSoutput.n264 CSoutput.n257 0.00252698
R22709 CSoutput.n253 CSoutput.n242 0.00252698
R22710 CSoutput.n252 CSoutput.n244 0.00252698
R22711 CSoutput.n251 CSoutput.n246 0.00252698
R22712 CSoutput.n266 CSoutput.n218 0.00252698
R22713 CSoutput.n255 CSoutput.n220 0.00252698
R22714 CSoutput.n257 CSoutput.n219 0.00252698
R22715 CSoutput.n165 CSoutput.n159 0.00252698
R22716 CSoutput.n158 CSoutput.n156 0.00252698
R22717 CSoutput.n284 CSoutput.n283 0.00252698
R22718 CSoutput.n168 CSoutput.n166 0.00252698
R22719 CSoutput.n171 CSoutput.n169 0.00252698
R22720 CSoutput.n288 CSoutput.n139 0.00252698
R22721 CSoutput.n165 CSoutput.n164 0.00252698
R22722 CSoutput.n158 CSoutput.n157 0.00252698
R22723 CSoutput.n285 CSoutput.n284 0.00252698
R22724 CSoutput.n168 CSoutput.n167 0.00252698
R22725 CSoutput.n171 CSoutput.n170 0.00252698
R22726 CSoutput.n152 CSoutput.n139 0.00252698
R22727 CSoutput.n273 CSoutput.n272 0.0020275
R22728 CSoutput.n272 CSoutput.n271 0.0020275
R22729 CSoutput.n269 CSoutput.n207 0.0020275
R22730 CSoutput.n269 CSoutput.n268 0.0020275
R22731 CSoutput.n283 CSoutput.n282 0.0020275
R22732 CSoutput.n282 CSoutput.n281 0.0020275
R22733 CSoutput.n183 CSoutput.n182 0.00166668
R22734 CSoutput.n265 CSoutput.n221 0.00166668
R22735 CSoutput.n149 CSoutput.n148 0.00166668
R22736 CSoutput.n287 CSoutput.n149 0.00133328
R22737 CSoutput.n221 CSoutput.n217 0.00133328
R22738 CSoutput.n277 CSoutput.n183 0.00133328
R22739 CSoutput.n280 CSoutput.n172 0.001
R22740 CSoutput.n258 CSoutput.n172 0.001
R22741 CSoutput.n160 CSoutput.n140 0.001
R22742 CSoutput.n259 CSoutput.n140 0.001
R22743 CSoutput.n161 CSoutput.n141 0.001
R22744 CSoutput.n260 CSoutput.n141 0.001
R22745 CSoutput.n162 CSoutput.n142 0.001
R22746 CSoutput.n261 CSoutput.n142 0.001
R22747 CSoutput.n163 CSoutput.n143 0.001
R22748 CSoutput.n262 CSoutput.n143 0.001
R22749 CSoutput.n256 CSoutput.n208 0.001
R22750 CSoutput.n256 CSoutput.n254 0.001
R22751 CSoutput.n238 CSoutput.n209 0.001
R22752 CSoutput.n232 CSoutput.n209 0.001
R22753 CSoutput.n239 CSoutput.n210 0.001
R22754 CSoutput.n233 CSoutput.n210 0.001
R22755 CSoutput.n240 CSoutput.n211 0.001
R22756 CSoutput.n234 CSoutput.n211 0.001
R22757 CSoutput.n241 CSoutput.n212 0.001
R22758 CSoutput.n235 CSoutput.n212 0.001
R22759 CSoutput.n270 CSoutput.n206 0.001
R22760 CSoutput.n224 CSoutput.n206 0.001
R22761 CSoutput.n194 CSoutput.n174 0.001
R22762 CSoutput.n225 CSoutput.n174 0.001
R22763 CSoutput.n195 CSoutput.n175 0.001
R22764 CSoutput.n226 CSoutput.n175 0.001
R22765 CSoutput.n196 CSoutput.n176 0.001
R22766 CSoutput.n227 CSoutput.n176 0.001
R22767 CSoutput.n197 CSoutput.n177 0.001
R22768 CSoutput.n228 CSoutput.n177 0.001
R22769 CSoutput.n228 CSoutput.n178 0.001
R22770 CSoutput.n227 CSoutput.n179 0.001
R22771 CSoutput.n226 CSoutput.n180 0.001
R22772 CSoutput.n225 CSoutput.t198 0.001
R22773 CSoutput.n224 CSoutput.n181 0.001
R22774 CSoutput.n197 CSoutput.n179 0.001
R22775 CSoutput.n196 CSoutput.n180 0.001
R22776 CSoutput.n195 CSoutput.t198 0.001
R22777 CSoutput.n194 CSoutput.n181 0.001
R22778 CSoutput.n270 CSoutput.n182 0.001
R22779 CSoutput.n235 CSoutput.n213 0.001
R22780 CSoutput.n234 CSoutput.n214 0.001
R22781 CSoutput.n233 CSoutput.n215 0.001
R22782 CSoutput.n232 CSoutput.t206 0.001
R22783 CSoutput.n254 CSoutput.n216 0.001
R22784 CSoutput.n241 CSoutput.n214 0.001
R22785 CSoutput.n240 CSoutput.n215 0.001
R22786 CSoutput.n239 CSoutput.t206 0.001
R22787 CSoutput.n238 CSoutput.n216 0.001
R22788 CSoutput.n265 CSoutput.n208 0.001
R22789 CSoutput.n262 CSoutput.n144 0.001
R22790 CSoutput.n261 CSoutput.n145 0.001
R22791 CSoutput.n260 CSoutput.n146 0.001
R22792 CSoutput.n259 CSoutput.t209 0.001
R22793 CSoutput.n258 CSoutput.n147 0.001
R22794 CSoutput.n163 CSoutput.n145 0.001
R22795 CSoutput.n162 CSoutput.n146 0.001
R22796 CSoutput.n161 CSoutput.t209 0.001
R22797 CSoutput.n160 CSoutput.n147 0.001
R22798 CSoutput.n280 CSoutput.n148 0.001
R22799 a_n9628_8799.n231 a_n9628_8799.t145 485.149
R22800 a_n9628_8799.n250 a_n9628_8799.t160 485.149
R22801 a_n9628_8799.n270 a_n9628_8799.t83 485.149
R22802 a_n9628_8799.n170 a_n9628_8799.t97 485.149
R22803 a_n9628_8799.n189 a_n9628_8799.t110 485.149
R22804 a_n9628_8799.n209 a_n9628_8799.t81 485.149
R22805 a_n9628_8799.n58 a_n9628_8799.t55 485.135
R22806 a_n9628_8799.n243 a_n9628_8799.t53 464.166
R22807 a_n9628_8799.n225 a_n9628_8799.t139 464.166
R22808 a_n9628_8799.n242 a_n9628_8799.t75 464.166
R22809 a_n9628_8799.n241 a_n9628_8799.t58 464.166
R22810 a_n9628_8799.n226 a_n9628_8799.t146 464.166
R22811 a_n9628_8799.n240 a_n9628_8799.t101 464.166
R22812 a_n9628_8799.n239 a_n9628_8799.t76 464.166
R22813 a_n9628_8799.n227 a_n9628_8799.t164 464.166
R22814 a_n9628_8799.n238 a_n9628_8799.t119 464.166
R22815 a_n9628_8799.n237 a_n9628_8799.t79 464.166
R22816 a_n9628_8799.n228 a_n9628_8799.t158 464.166
R22817 a_n9628_8799.n236 a_n9628_8799.t121 464.166
R22818 a_n9628_8799.n235 a_n9628_8799.t93 464.166
R22819 a_n9628_8799.n229 a_n9628_8799.t54 464.166
R22820 a_n9628_8799.n234 a_n9628_8799.t142 464.166
R22821 a_n9628_8799.n233 a_n9628_8799.t123 464.166
R22822 a_n9628_8799.n230 a_n9628_8799.t59 464.166
R22823 a_n9628_8799.n232 a_n9628_8799.t149 464.166
R22824 a_n9628_8799.n73 a_n9628_8799.t66 485.135
R22825 a_n9628_8799.n262 a_n9628_8799.t65 464.166
R22826 a_n9628_8799.n244 a_n9628_8799.t156 464.166
R22827 a_n9628_8799.n261 a_n9628_8799.t84 464.166
R22828 a_n9628_8799.n260 a_n9628_8799.t73 464.166
R22829 a_n9628_8799.n245 a_n9628_8799.t159 464.166
R22830 a_n9628_8799.n259 a_n9628_8799.t115 464.166
R22831 a_n9628_8799.n258 a_n9628_8799.t87 464.166
R22832 a_n9628_8799.n246 a_n9628_8799.t57 464.166
R22833 a_n9628_8799.n257 a_n9628_8799.t132 464.166
R22834 a_n9628_8799.n256 a_n9628_8799.t88 464.166
R22835 a_n9628_8799.n247 a_n9628_8799.t49 464.166
R22836 a_n9628_8799.n255 a_n9628_8799.t137 464.166
R22837 a_n9628_8799.n254 a_n9628_8799.t103 464.166
R22838 a_n9628_8799.n248 a_n9628_8799.t67 464.166
R22839 a_n9628_8799.n253 a_n9628_8799.t157 464.166
R22840 a_n9628_8799.n252 a_n9628_8799.t138 464.166
R22841 a_n9628_8799.n249 a_n9628_8799.t74 464.166
R22842 a_n9628_8799.n251 a_n9628_8799.t161 464.166
R22843 a_n9628_8799.n88 a_n9628_8799.t114 485.135
R22844 a_n9628_8799.n282 a_n9628_8799.t136 464.166
R22845 a_n9628_8799.n264 a_n9628_8799.t72 464.166
R22846 a_n9628_8799.n281 a_n9628_8799.t154 464.166
R22847 a_n9628_8799.n280 a_n9628_8799.t91 464.166
R22848 a_n9628_8799.n265 a_n9628_8799.t147 464.166
R22849 a_n9628_8799.n279 a_n9628_8799.t78 464.166
R22850 a_n9628_8799.n278 a_n9628_8799.t126 464.166
R22851 a_n9628_8799.n266 a_n9628_8799.t63 464.166
R22852 a_n9628_8799.n277 a_n9628_8799.t109 464.166
R22853 a_n9628_8799.n276 a_n9628_8799.t86 464.166
R22854 a_n9628_8799.n267 a_n9628_8799.t134 464.166
R22855 a_n9628_8799.n275 a_n9628_8799.t70 464.166
R22856 a_n9628_8799.n274 a_n9628_8799.t118 464.166
R22857 a_n9628_8799.n268 a_n9628_8799.t52 464.166
R22858 a_n9628_8799.n273 a_n9628_8799.t102 464.166
R22859 a_n9628_8799.n272 a_n9628_8799.t166 464.166
R22860 a_n9628_8799.n269 a_n9628_8799.t125 464.166
R22861 a_n9628_8799.n271 a_n9628_8799.t62 464.166
R22862 a_n9628_8799.n171 a_n9628_8799.t99 464.166
R22863 a_n9628_8799.n172 a_n9628_8799.t131 464.166
R22864 a_n9628_8799.n173 a_n9628_8799.t56 464.166
R22865 a_n9628_8799.n174 a_n9628_8799.t95 464.166
R22866 a_n9628_8799.n169 a_n9628_8799.t127 464.166
R22867 a_n9628_8799.n175 a_n9628_8799.t50 464.166
R22868 a_n9628_8799.n176 a_n9628_8799.t82 464.166
R22869 a_n9628_8799.n177 a_n9628_8799.t120 464.166
R22870 a_n9628_8799.n178 a_n9628_8799.t155 464.166
R22871 a_n9628_8799.n168 a_n9628_8799.t80 464.166
R22872 a_n9628_8799.n179 a_n9628_8799.t116 464.166
R22873 a_n9628_8799.n167 a_n9628_8799.t151 464.166
R22874 a_n9628_8799.n180 a_n9628_8799.t152 464.166
R22875 a_n9628_8799.n181 a_n9628_8799.t98 464.166
R22876 a_n9628_8799.n182 a_n9628_8799.t130 464.166
R22877 a_n9628_8799.n183 a_n9628_8799.t150 464.166
R22878 a_n9628_8799.n166 a_n9628_8799.t94 464.166
R22879 a_n9628_8799.n184 a_n9628_8799.t96 464.166
R22880 a_n9628_8799.n190 a_n9628_8799.t112 464.166
R22881 a_n9628_8799.n191 a_n9628_8799.t148 464.166
R22882 a_n9628_8799.n192 a_n9628_8799.t68 464.166
R22883 a_n9628_8799.n193 a_n9628_8799.t106 464.166
R22884 a_n9628_8799.n188 a_n9628_8799.t140 464.166
R22885 a_n9628_8799.n194 a_n9628_8799.t64 464.166
R22886 a_n9628_8799.n195 a_n9628_8799.t92 464.166
R22887 a_n9628_8799.n196 a_n9628_8799.t133 464.166
R22888 a_n9628_8799.n197 a_n9628_8799.t167 464.166
R22889 a_n9628_8799.n187 a_n9628_8799.t89 464.166
R22890 a_n9628_8799.n198 a_n9628_8799.t129 464.166
R22891 a_n9628_8799.n186 a_n9628_8799.t163 464.166
R22892 a_n9628_8799.n199 a_n9628_8799.t165 464.166
R22893 a_n9628_8799.n200 a_n9628_8799.t111 464.166
R22894 a_n9628_8799.n201 a_n9628_8799.t144 464.166
R22895 a_n9628_8799.n202 a_n9628_8799.t162 464.166
R22896 a_n9628_8799.n185 a_n9628_8799.t105 464.166
R22897 a_n9628_8799.n203 a_n9628_8799.t107 464.166
R22898 a_n9628_8799.n210 a_n9628_8799.t60 464.166
R22899 a_n9628_8799.n211 a_n9628_8799.t122 464.166
R22900 a_n9628_8799.n212 a_n9628_8799.t77 464.166
R22901 a_n9628_8799.n213 a_n9628_8799.t100 464.166
R22902 a_n9628_8799.n208 a_n9628_8799.t51 464.166
R22903 a_n9628_8799.n214 a_n9628_8799.t117 464.166
R22904 a_n9628_8799.n215 a_n9628_8799.t69 464.166
R22905 a_n9628_8799.n216 a_n9628_8799.t135 464.166
R22906 a_n9628_8799.n217 a_n9628_8799.t85 464.166
R22907 a_n9628_8799.n207 a_n9628_8799.t108 464.166
R22908 a_n9628_8799.n218 a_n9628_8799.t61 464.166
R22909 a_n9628_8799.n206 a_n9628_8799.t124 464.166
R22910 a_n9628_8799.n219 a_n9628_8799.t104 464.166
R22911 a_n9628_8799.n220 a_n9628_8799.t143 464.166
R22912 a_n9628_8799.n221 a_n9628_8799.t90 464.166
R22913 a_n9628_8799.n222 a_n9628_8799.t153 464.166
R22914 a_n9628_8799.n205 a_n9628_8799.t71 464.166
R22915 a_n9628_8799.n223 a_n9628_8799.t48 464.166
R22916 a_n9628_8799.n45 a_n9628_8799.n72 71.7212
R22917 a_n9628_8799.n72 a_n9628_8799.n230 17.8606
R22918 a_n9628_8799.n71 a_n9628_8799.n45 76.9909
R22919 a_n9628_8799.n233 a_n9628_8799.n71 7.32118
R22920 a_n9628_8799.n70 a_n9628_8799.n44 78.3454
R22921 a_n9628_8799.n44 a_n9628_8799.n69 72.8951
R22922 a_n9628_8799.n68 a_n9628_8799.n46 70.1674
R22923 a_n9628_8799.n236 a_n9628_8799.n68 20.9683
R22924 a_n9628_8799.n46 a_n9628_8799.n67 72.3034
R22925 a_n9628_8799.n67 a_n9628_8799.n228 16.6962
R22926 a_n9628_8799.n66 a_n9628_8799.n47 77.6622
R22927 a_n9628_8799.n237 a_n9628_8799.n66 5.97853
R22928 a_n9628_8799.n65 a_n9628_8799.n47 77.6622
R22929 a_n9628_8799.n48 a_n9628_8799.n64 72.3034
R22930 a_n9628_8799.n63 a_n9628_8799.n48 70.1674
R22931 a_n9628_8799.n240 a_n9628_8799.n63 20.9683
R22932 a_n9628_8799.n50 a_n9628_8799.n62 72.8951
R22933 a_n9628_8799.n62 a_n9628_8799.n226 15.5127
R22934 a_n9628_8799.n61 a_n9628_8799.n50 78.3454
R22935 a_n9628_8799.n241 a_n9628_8799.n61 4.61226
R22936 a_n9628_8799.n60 a_n9628_8799.n49 76.9909
R22937 a_n9628_8799.n49 a_n9628_8799.n59 71.7212
R22938 a_n9628_8799.n243 a_n9628_8799.n58 20.9683
R22939 a_n9628_8799.n51 a_n9628_8799.n58 70.1674
R22940 a_n9628_8799.n37 a_n9628_8799.n87 71.7212
R22941 a_n9628_8799.n87 a_n9628_8799.n249 17.8606
R22942 a_n9628_8799.n86 a_n9628_8799.n37 76.9909
R22943 a_n9628_8799.n252 a_n9628_8799.n86 7.32118
R22944 a_n9628_8799.n85 a_n9628_8799.n36 78.3454
R22945 a_n9628_8799.n36 a_n9628_8799.n84 72.8951
R22946 a_n9628_8799.n83 a_n9628_8799.n38 70.1674
R22947 a_n9628_8799.n255 a_n9628_8799.n83 20.9683
R22948 a_n9628_8799.n38 a_n9628_8799.n82 72.3034
R22949 a_n9628_8799.n82 a_n9628_8799.n247 16.6962
R22950 a_n9628_8799.n81 a_n9628_8799.n39 77.6622
R22951 a_n9628_8799.n256 a_n9628_8799.n81 5.97853
R22952 a_n9628_8799.n80 a_n9628_8799.n39 77.6622
R22953 a_n9628_8799.n40 a_n9628_8799.n79 72.3034
R22954 a_n9628_8799.n78 a_n9628_8799.n40 70.1674
R22955 a_n9628_8799.n259 a_n9628_8799.n78 20.9683
R22956 a_n9628_8799.n42 a_n9628_8799.n77 72.8951
R22957 a_n9628_8799.n77 a_n9628_8799.n245 15.5127
R22958 a_n9628_8799.n76 a_n9628_8799.n42 78.3454
R22959 a_n9628_8799.n260 a_n9628_8799.n76 4.61226
R22960 a_n9628_8799.n75 a_n9628_8799.n41 76.9909
R22961 a_n9628_8799.n41 a_n9628_8799.n74 71.7212
R22962 a_n9628_8799.n262 a_n9628_8799.n73 20.9683
R22963 a_n9628_8799.n43 a_n9628_8799.n73 70.1674
R22964 a_n9628_8799.n29 a_n9628_8799.n102 71.7212
R22965 a_n9628_8799.n102 a_n9628_8799.n269 17.8606
R22966 a_n9628_8799.n101 a_n9628_8799.n29 76.9909
R22967 a_n9628_8799.n272 a_n9628_8799.n101 7.32118
R22968 a_n9628_8799.n100 a_n9628_8799.n28 78.3454
R22969 a_n9628_8799.n28 a_n9628_8799.n99 72.8951
R22970 a_n9628_8799.n98 a_n9628_8799.n30 70.1674
R22971 a_n9628_8799.n275 a_n9628_8799.n98 20.9683
R22972 a_n9628_8799.n30 a_n9628_8799.n97 72.3034
R22973 a_n9628_8799.n97 a_n9628_8799.n267 16.6962
R22974 a_n9628_8799.n96 a_n9628_8799.n31 77.6622
R22975 a_n9628_8799.n276 a_n9628_8799.n96 5.97853
R22976 a_n9628_8799.n95 a_n9628_8799.n31 77.6622
R22977 a_n9628_8799.n32 a_n9628_8799.n94 72.3034
R22978 a_n9628_8799.n93 a_n9628_8799.n32 70.1674
R22979 a_n9628_8799.n279 a_n9628_8799.n93 20.9683
R22980 a_n9628_8799.n34 a_n9628_8799.n92 72.8951
R22981 a_n9628_8799.n92 a_n9628_8799.n265 15.5127
R22982 a_n9628_8799.n91 a_n9628_8799.n34 78.3454
R22983 a_n9628_8799.n280 a_n9628_8799.n91 4.61226
R22984 a_n9628_8799.n90 a_n9628_8799.n33 76.9909
R22985 a_n9628_8799.n33 a_n9628_8799.n89 71.7212
R22986 a_n9628_8799.n282 a_n9628_8799.n88 20.9683
R22987 a_n9628_8799.n35 a_n9628_8799.n88 70.1674
R22988 a_n9628_8799.n21 a_n9628_8799.n117 70.1674
R22989 a_n9628_8799.n184 a_n9628_8799.n117 20.9683
R22990 a_n9628_8799.n116 a_n9628_8799.n21 71.7212
R22991 a_n9628_8799.n116 a_n9628_8799.n166 17.8606
R22992 a_n9628_8799.n20 a_n9628_8799.n115 76.9909
R22993 a_n9628_8799.n183 a_n9628_8799.n115 7.32118
R22994 a_n9628_8799.n114 a_n9628_8799.n20 78.3454
R22995 a_n9628_8799.n22 a_n9628_8799.n113 72.8951
R22996 a_n9628_8799.n112 a_n9628_8799.n22 70.1674
R22997 a_n9628_8799.n112 a_n9628_8799.n167 20.9683
R22998 a_n9628_8799.n23 a_n9628_8799.n111 72.3034
R22999 a_n9628_8799.n179 a_n9628_8799.n111 16.6962
R23000 a_n9628_8799.n110 a_n9628_8799.n23 77.6622
R23001 a_n9628_8799.n110 a_n9628_8799.n168 5.97853
R23002 a_n9628_8799.n24 a_n9628_8799.n109 77.6622
R23003 a_n9628_8799.n108 a_n9628_8799.n24 72.3034
R23004 a_n9628_8799.n25 a_n9628_8799.n107 70.1674
R23005 a_n9628_8799.n175 a_n9628_8799.n107 20.9683
R23006 a_n9628_8799.n106 a_n9628_8799.n25 72.8951
R23007 a_n9628_8799.n106 a_n9628_8799.n169 15.5127
R23008 a_n9628_8799.n26 a_n9628_8799.n105 78.3454
R23009 a_n9628_8799.n174 a_n9628_8799.n105 4.61226
R23010 a_n9628_8799.n104 a_n9628_8799.n26 76.9909
R23011 a_n9628_8799.n103 a_n9628_8799.n172 17.8606
R23012 a_n9628_8799.n103 a_n9628_8799.n27 71.7212
R23013 a_n9628_8799.n13 a_n9628_8799.n132 70.1674
R23014 a_n9628_8799.n203 a_n9628_8799.n132 20.9683
R23015 a_n9628_8799.n131 a_n9628_8799.n13 71.7212
R23016 a_n9628_8799.n131 a_n9628_8799.n185 17.8606
R23017 a_n9628_8799.n12 a_n9628_8799.n130 76.9909
R23018 a_n9628_8799.n202 a_n9628_8799.n130 7.32118
R23019 a_n9628_8799.n129 a_n9628_8799.n12 78.3454
R23020 a_n9628_8799.n14 a_n9628_8799.n128 72.8951
R23021 a_n9628_8799.n127 a_n9628_8799.n14 70.1674
R23022 a_n9628_8799.n127 a_n9628_8799.n186 20.9683
R23023 a_n9628_8799.n15 a_n9628_8799.n126 72.3034
R23024 a_n9628_8799.n198 a_n9628_8799.n126 16.6962
R23025 a_n9628_8799.n125 a_n9628_8799.n15 77.6622
R23026 a_n9628_8799.n125 a_n9628_8799.n187 5.97853
R23027 a_n9628_8799.n16 a_n9628_8799.n124 77.6622
R23028 a_n9628_8799.n123 a_n9628_8799.n16 72.3034
R23029 a_n9628_8799.n17 a_n9628_8799.n122 70.1674
R23030 a_n9628_8799.n194 a_n9628_8799.n122 20.9683
R23031 a_n9628_8799.n121 a_n9628_8799.n17 72.8951
R23032 a_n9628_8799.n121 a_n9628_8799.n188 15.5127
R23033 a_n9628_8799.n18 a_n9628_8799.n120 78.3454
R23034 a_n9628_8799.n193 a_n9628_8799.n120 4.61226
R23035 a_n9628_8799.n119 a_n9628_8799.n18 76.9909
R23036 a_n9628_8799.n118 a_n9628_8799.n191 17.8606
R23037 a_n9628_8799.n118 a_n9628_8799.n19 71.7212
R23038 a_n9628_8799.n5 a_n9628_8799.n147 70.1674
R23039 a_n9628_8799.n223 a_n9628_8799.n147 20.9683
R23040 a_n9628_8799.n146 a_n9628_8799.n5 71.7212
R23041 a_n9628_8799.n146 a_n9628_8799.n205 17.8606
R23042 a_n9628_8799.n4 a_n9628_8799.n145 76.9909
R23043 a_n9628_8799.n222 a_n9628_8799.n145 7.32118
R23044 a_n9628_8799.n144 a_n9628_8799.n4 78.3454
R23045 a_n9628_8799.n6 a_n9628_8799.n143 72.8951
R23046 a_n9628_8799.n142 a_n9628_8799.n6 70.1674
R23047 a_n9628_8799.n142 a_n9628_8799.n206 20.9683
R23048 a_n9628_8799.n7 a_n9628_8799.n141 72.3034
R23049 a_n9628_8799.n218 a_n9628_8799.n141 16.6962
R23050 a_n9628_8799.n140 a_n9628_8799.n7 77.6622
R23051 a_n9628_8799.n140 a_n9628_8799.n207 5.97853
R23052 a_n9628_8799.n8 a_n9628_8799.n139 77.6622
R23053 a_n9628_8799.n138 a_n9628_8799.n8 72.3034
R23054 a_n9628_8799.n9 a_n9628_8799.n137 70.1674
R23055 a_n9628_8799.n214 a_n9628_8799.n137 20.9683
R23056 a_n9628_8799.n136 a_n9628_8799.n9 72.8951
R23057 a_n9628_8799.n136 a_n9628_8799.n208 15.5127
R23058 a_n9628_8799.n10 a_n9628_8799.n135 78.3454
R23059 a_n9628_8799.n213 a_n9628_8799.n135 4.61226
R23060 a_n9628_8799.n134 a_n9628_8799.n10 76.9909
R23061 a_n9628_8799.n133 a_n9628_8799.n211 17.8606
R23062 a_n9628_8799.n133 a_n9628_8799.n11 71.7212
R23063 a_n9628_8799.n52 a_n9628_8799.n148 98.9633
R23064 a_n9628_8799.n55 a_n9628_8799.n288 98.9631
R23065 a_n9628_8799.n55 a_n9628_8799.n289 98.6055
R23066 a_n9628_8799.n55 a_n9628_8799.n290 98.6055
R23067 a_n9628_8799.n57 a_n9628_8799.n291 98.6055
R23068 a_n9628_8799.n56 a_n9628_8799.n287 98.6055
R23069 a_n9628_8799.n54 a_n9628_8799.n153 98.6055
R23070 a_n9628_8799.n54 a_n9628_8799.n152 98.6055
R23071 a_n9628_8799.n53 a_n9628_8799.n151 98.6055
R23072 a_n9628_8799.n53 a_n9628_8799.n150 98.6055
R23073 a_n9628_8799.n52 a_n9628_8799.n149 98.6055
R23074 a_n9628_8799.n292 a_n9628_8799.n57 98.6054
R23075 a_n9628_8799.n1 a_n9628_8799.n154 81.4626
R23076 a_n9628_8799.n3 a_n9628_8799.n160 81.4626
R23077 a_n9628_8799.n0 a_n9628_8799.n157 81.4626
R23078 a_n9628_8799.n2 a_n9628_8799.n163 80.9324
R23079 a_n9628_8799.n2 a_n9628_8799.n164 80.9324
R23080 a_n9628_8799.n1 a_n9628_8799.n165 80.9324
R23081 a_n9628_8799.n1 a_n9628_8799.n156 80.9324
R23082 a_n9628_8799.n1 a_n9628_8799.n155 80.9324
R23083 a_n9628_8799.n3 a_n9628_8799.n161 80.9324
R23084 a_n9628_8799.n0 a_n9628_8799.n162 80.9324
R23085 a_n9628_8799.n0 a_n9628_8799.n159 80.9324
R23086 a_n9628_8799.n0 a_n9628_8799.n158 80.9324
R23087 a_n9628_8799.n45 a_n9628_8799.n231 70.4033
R23088 a_n9628_8799.n37 a_n9628_8799.n250 70.4033
R23089 a_n9628_8799.n29 a_n9628_8799.n270 70.4033
R23090 a_n9628_8799.n170 a_n9628_8799.n27 70.4033
R23091 a_n9628_8799.n189 a_n9628_8799.n19 70.4033
R23092 a_n9628_8799.n209 a_n9628_8799.n11 70.4033
R23093 a_n9628_8799.n242 a_n9628_8799.n241 48.2005
R23094 a_n9628_8799.n63 a_n9628_8799.n239 20.9683
R23095 a_n9628_8799.n238 a_n9628_8799.n237 48.2005
R23096 a_n9628_8799.n68 a_n9628_8799.n235 20.9683
R23097 a_n9628_8799.n234 a_n9628_8799.n233 48.2005
R23098 a_n9628_8799.n261 a_n9628_8799.n260 48.2005
R23099 a_n9628_8799.n78 a_n9628_8799.n258 20.9683
R23100 a_n9628_8799.n257 a_n9628_8799.n256 48.2005
R23101 a_n9628_8799.n83 a_n9628_8799.n254 20.9683
R23102 a_n9628_8799.n253 a_n9628_8799.n252 48.2005
R23103 a_n9628_8799.n281 a_n9628_8799.n280 48.2005
R23104 a_n9628_8799.n93 a_n9628_8799.n278 20.9683
R23105 a_n9628_8799.n277 a_n9628_8799.n276 48.2005
R23106 a_n9628_8799.n98 a_n9628_8799.n274 20.9683
R23107 a_n9628_8799.n273 a_n9628_8799.n272 48.2005
R23108 a_n9628_8799.n174 a_n9628_8799.n173 48.2005
R23109 a_n9628_8799.n176 a_n9628_8799.n107 20.9683
R23110 a_n9628_8799.n178 a_n9628_8799.n168 48.2005
R23111 a_n9628_8799.n180 a_n9628_8799.n112 20.9683
R23112 a_n9628_8799.n183 a_n9628_8799.n182 48.2005
R23113 a_n9628_8799.t128 a_n9628_8799.n117 485.135
R23114 a_n9628_8799.n193 a_n9628_8799.n192 48.2005
R23115 a_n9628_8799.n195 a_n9628_8799.n122 20.9683
R23116 a_n9628_8799.n197 a_n9628_8799.n187 48.2005
R23117 a_n9628_8799.n199 a_n9628_8799.n127 20.9683
R23118 a_n9628_8799.n202 a_n9628_8799.n201 48.2005
R23119 a_n9628_8799.t141 a_n9628_8799.n132 485.135
R23120 a_n9628_8799.n213 a_n9628_8799.n212 48.2005
R23121 a_n9628_8799.n215 a_n9628_8799.n137 20.9683
R23122 a_n9628_8799.n217 a_n9628_8799.n207 48.2005
R23123 a_n9628_8799.n219 a_n9628_8799.n142 20.9683
R23124 a_n9628_8799.n222 a_n9628_8799.n221 48.2005
R23125 a_n9628_8799.t113 a_n9628_8799.n147 485.135
R23126 a_n9628_8799.n59 a_n9628_8799.n225 17.8606
R23127 a_n9628_8799.n232 a_n9628_8799.n72 25.894
R23128 a_n9628_8799.n74 a_n9628_8799.n244 17.8606
R23129 a_n9628_8799.n251 a_n9628_8799.n87 25.894
R23130 a_n9628_8799.n89 a_n9628_8799.n264 17.8606
R23131 a_n9628_8799.n271 a_n9628_8799.n102 25.894
R23132 a_n9628_8799.n184 a_n9628_8799.n116 25.894
R23133 a_n9628_8799.n203 a_n9628_8799.n131 25.894
R23134 a_n9628_8799.n223 a_n9628_8799.n146 25.894
R23135 a_n9628_8799.n70 a_n9628_8799.n229 43.3183
R23136 a_n9628_8799.n85 a_n9628_8799.n248 43.3183
R23137 a_n9628_8799.n100 a_n9628_8799.n268 43.3183
R23138 a_n9628_8799.n181 a_n9628_8799.n114 43.3183
R23139 a_n9628_8799.n200 a_n9628_8799.n129 43.3183
R23140 a_n9628_8799.n220 a_n9628_8799.n144 43.3183
R23141 a_n9628_8799.n64 a_n9628_8799.n227 16.6962
R23142 a_n9628_8799.n236 a_n9628_8799.n67 27.6507
R23143 a_n9628_8799.n79 a_n9628_8799.n246 16.6962
R23144 a_n9628_8799.n255 a_n9628_8799.n82 27.6507
R23145 a_n9628_8799.n94 a_n9628_8799.n266 16.6962
R23146 a_n9628_8799.n275 a_n9628_8799.n97 27.6507
R23147 a_n9628_8799.n177 a_n9628_8799.n108 16.6962
R23148 a_n9628_8799.n167 a_n9628_8799.n111 27.6507
R23149 a_n9628_8799.n196 a_n9628_8799.n123 16.6962
R23150 a_n9628_8799.n186 a_n9628_8799.n126 27.6507
R23151 a_n9628_8799.n216 a_n9628_8799.n138 16.6962
R23152 a_n9628_8799.n206 a_n9628_8799.n141 27.6507
R23153 a_n9628_8799.n65 a_n9628_8799.n227 41.7634
R23154 a_n9628_8799.n80 a_n9628_8799.n246 41.7634
R23155 a_n9628_8799.n95 a_n9628_8799.n266 41.7634
R23156 a_n9628_8799.n109 a_n9628_8799.n177 41.7634
R23157 a_n9628_8799.n124 a_n9628_8799.n196 41.7634
R23158 a_n9628_8799.n139 a_n9628_8799.n216 41.7634
R23159 a_n9628_8799.n56 a_n9628_8799.n286 34.414
R23160 a_n9628_8799.n240 a_n9628_8799.n62 29.3885
R23161 a_n9628_8799.n69 a_n9628_8799.n229 15.5127
R23162 a_n9628_8799.n259 a_n9628_8799.n77 29.3885
R23163 a_n9628_8799.n84 a_n9628_8799.n248 15.5127
R23164 a_n9628_8799.n279 a_n9628_8799.n92 29.3885
R23165 a_n9628_8799.n99 a_n9628_8799.n268 15.5127
R23166 a_n9628_8799.n175 a_n9628_8799.n106 29.3885
R23167 a_n9628_8799.n181 a_n9628_8799.n113 15.5127
R23168 a_n9628_8799.n194 a_n9628_8799.n121 29.3885
R23169 a_n9628_8799.n200 a_n9628_8799.n128 15.5127
R23170 a_n9628_8799.n214 a_n9628_8799.n136 29.3885
R23171 a_n9628_8799.n220 a_n9628_8799.n143 15.5127
R23172 a_n9628_8799.n2 a_n9628_8799.n0 34.3237
R23173 a_n9628_8799.n60 a_n9628_8799.n225 40.1848
R23174 a_n9628_8799.n75 a_n9628_8799.n244 40.1848
R23175 a_n9628_8799.n90 a_n9628_8799.n264 40.1848
R23176 a_n9628_8799.n172 a_n9628_8799.n104 40.1848
R23177 a_n9628_8799.n191 a_n9628_8799.n119 40.1848
R23178 a_n9628_8799.n211 a_n9628_8799.n134 40.1848
R23179 a_n9628_8799.n232 a_n9628_8799.n231 20.9576
R23180 a_n9628_8799.n251 a_n9628_8799.n250 20.9576
R23181 a_n9628_8799.n271 a_n9628_8799.n270 20.9576
R23182 a_n9628_8799.n171 a_n9628_8799.n170 20.9576
R23183 a_n9628_8799.n190 a_n9628_8799.n189 20.9576
R23184 a_n9628_8799.n210 a_n9628_8799.n209 20.9576
R23185 a_n9628_8799.n286 a_n9628_8799.n54 20.4753
R23186 a_n9628_8799.n60 a_n9628_8799.n242 7.32118
R23187 a_n9628_8799.n71 a_n9628_8799.n230 40.1848
R23188 a_n9628_8799.n75 a_n9628_8799.n261 7.32118
R23189 a_n9628_8799.n86 a_n9628_8799.n249 40.1848
R23190 a_n9628_8799.n90 a_n9628_8799.n281 7.32118
R23191 a_n9628_8799.n101 a_n9628_8799.n269 40.1848
R23192 a_n9628_8799.n173 a_n9628_8799.n104 7.32118
R23193 a_n9628_8799.n166 a_n9628_8799.n115 40.1848
R23194 a_n9628_8799.n192 a_n9628_8799.n119 7.32118
R23195 a_n9628_8799.n185 a_n9628_8799.n130 40.1848
R23196 a_n9628_8799.n212 a_n9628_8799.n134 7.32118
R23197 a_n9628_8799.n205 a_n9628_8799.n145 40.1848
R23198 a_n9628_8799.n235 a_n9628_8799.n69 29.3885
R23199 a_n9628_8799.n254 a_n9628_8799.n84 29.3885
R23200 a_n9628_8799.n274 a_n9628_8799.n99 29.3885
R23201 a_n9628_8799.n113 a_n9628_8799.n180 29.3885
R23202 a_n9628_8799.n128 a_n9628_8799.n199 29.3885
R23203 a_n9628_8799.n143 a_n9628_8799.n219 29.3885
R23204 a_n9628_8799.n65 a_n9628_8799.n238 5.97853
R23205 a_n9628_8799.n66 a_n9628_8799.n228 41.7634
R23206 a_n9628_8799.n80 a_n9628_8799.n257 5.97853
R23207 a_n9628_8799.n81 a_n9628_8799.n247 41.7634
R23208 a_n9628_8799.n95 a_n9628_8799.n277 5.97853
R23209 a_n9628_8799.n96 a_n9628_8799.n267 41.7634
R23210 a_n9628_8799.n178 a_n9628_8799.n109 5.97853
R23211 a_n9628_8799.n179 a_n9628_8799.n110 41.7634
R23212 a_n9628_8799.n197 a_n9628_8799.n124 5.97853
R23213 a_n9628_8799.n198 a_n9628_8799.n125 41.7634
R23214 a_n9628_8799.n217 a_n9628_8799.n139 5.97853
R23215 a_n9628_8799.n218 a_n9628_8799.n140 41.7634
R23216 a_n9628_8799.n285 a_n9628_8799.n1 12.3339
R23217 a_n9628_8799.n286 a_n9628_8799.n285 11.4887
R23218 a_n9628_8799.n239 a_n9628_8799.n64 27.6507
R23219 a_n9628_8799.n258 a_n9628_8799.n79 27.6507
R23220 a_n9628_8799.n278 a_n9628_8799.n94 27.6507
R23221 a_n9628_8799.n176 a_n9628_8799.n108 27.6507
R23222 a_n9628_8799.n195 a_n9628_8799.n123 27.6507
R23223 a_n9628_8799.n215 a_n9628_8799.n138 27.6507
R23224 a_n9628_8799.n61 a_n9628_8799.n226 43.3183
R23225 a_n9628_8799.n70 a_n9628_8799.n234 4.61226
R23226 a_n9628_8799.n76 a_n9628_8799.n245 43.3183
R23227 a_n9628_8799.n85 a_n9628_8799.n253 4.61226
R23228 a_n9628_8799.n91 a_n9628_8799.n265 43.3183
R23229 a_n9628_8799.n100 a_n9628_8799.n273 4.61226
R23230 a_n9628_8799.n169 a_n9628_8799.n105 43.3183
R23231 a_n9628_8799.n182 a_n9628_8799.n114 4.61226
R23232 a_n9628_8799.n188 a_n9628_8799.n120 43.3183
R23233 a_n9628_8799.n201 a_n9628_8799.n129 4.61226
R23234 a_n9628_8799.n208 a_n9628_8799.n135 43.3183
R23235 a_n9628_8799.n221 a_n9628_8799.n144 4.61226
R23236 a_n9628_8799.n263 a_n9628_8799.n51 9.04406
R23237 a_n9628_8799.n204 a_n9628_8799.n21 9.04406
R23238 a_n9628_8799.n243 a_n9628_8799.n59 25.894
R23239 a_n9628_8799.n262 a_n9628_8799.n74 25.894
R23240 a_n9628_8799.n282 a_n9628_8799.n89 25.894
R23241 a_n9628_8799.n103 a_n9628_8799.n171 25.894
R23242 a_n9628_8799.n118 a_n9628_8799.n190 25.894
R23243 a_n9628_8799.n133 a_n9628_8799.n210 25.894
R23244 a_n9628_8799.n284 a_n9628_8799.n224 7.2518
R23245 a_n9628_8799.n284 a_n9628_8799.n283 6.75517
R23246 a_n9628_8799.n263 a_n9628_8799.n43 4.93611
R23247 a_n9628_8799.n283 a_n9628_8799.n35 4.93611
R23248 a_n9628_8799.n204 a_n9628_8799.n13 4.93611
R23249 a_n9628_8799.n224 a_n9628_8799.n5 4.93611
R23250 a_n9628_8799.n283 a_n9628_8799.n263 4.10845
R23251 a_n9628_8799.n224 a_n9628_8799.n204 4.10845
R23252 a_n9628_8799.n288 a_n9628_8799.t27 3.61217
R23253 a_n9628_8799.n288 a_n9628_8799.t41 3.61217
R23254 a_n9628_8799.n289 a_n9628_8799.t43 3.61217
R23255 a_n9628_8799.n289 a_n9628_8799.t23 3.61217
R23256 a_n9628_8799.n290 a_n9628_8799.t33 3.61217
R23257 a_n9628_8799.n290 a_n9628_8799.t32 3.61217
R23258 a_n9628_8799.n291 a_n9628_8799.t31 3.61217
R23259 a_n9628_8799.n291 a_n9628_8799.t36 3.61217
R23260 a_n9628_8799.n287 a_n9628_8799.t28 3.61217
R23261 a_n9628_8799.n287 a_n9628_8799.t38 3.61217
R23262 a_n9628_8799.n153 a_n9628_8799.t39 3.61217
R23263 a_n9628_8799.n153 a_n9628_8799.t21 3.61217
R23264 a_n9628_8799.n152 a_n9628_8799.t25 3.61217
R23265 a_n9628_8799.n152 a_n9628_8799.t35 3.61217
R23266 a_n9628_8799.n151 a_n9628_8799.t29 3.61217
R23267 a_n9628_8799.n151 a_n9628_8799.t42 3.61217
R23268 a_n9628_8799.n150 a_n9628_8799.t26 3.61217
R23269 a_n9628_8799.n150 a_n9628_8799.t30 3.61217
R23270 a_n9628_8799.n149 a_n9628_8799.t24 3.61217
R23271 a_n9628_8799.n149 a_n9628_8799.t40 3.61217
R23272 a_n9628_8799.n148 a_n9628_8799.t34 3.61217
R23273 a_n9628_8799.n148 a_n9628_8799.t22 3.61217
R23274 a_n9628_8799.n292 a_n9628_8799.t37 3.61217
R23275 a_n9628_8799.t20 a_n9628_8799.n292 3.61217
R23276 a_n9628_8799.n285 a_n9628_8799.n284 3.4105
R23277 a_n9628_8799.n163 a_n9628_8799.t9 2.82907
R23278 a_n9628_8799.n163 a_n9628_8799.t11 2.82907
R23279 a_n9628_8799.n164 a_n9628_8799.t13 2.82907
R23280 a_n9628_8799.n164 a_n9628_8799.t45 2.82907
R23281 a_n9628_8799.n165 a_n9628_8799.t14 2.82907
R23282 a_n9628_8799.n165 a_n9628_8799.t1 2.82907
R23283 a_n9628_8799.n156 a_n9628_8799.t16 2.82907
R23284 a_n9628_8799.n156 a_n9628_8799.t7 2.82907
R23285 a_n9628_8799.n155 a_n9628_8799.t3 2.82907
R23286 a_n9628_8799.n155 a_n9628_8799.t18 2.82907
R23287 a_n9628_8799.n154 a_n9628_8799.t19 2.82907
R23288 a_n9628_8799.n154 a_n9628_8799.t5 2.82907
R23289 a_n9628_8799.n160 a_n9628_8799.t4 2.82907
R23290 a_n9628_8799.n160 a_n9628_8799.t10 2.82907
R23291 a_n9628_8799.n161 a_n9628_8799.t47 2.82907
R23292 a_n9628_8799.n161 a_n9628_8799.t46 2.82907
R23293 a_n9628_8799.n162 a_n9628_8799.t6 2.82907
R23294 a_n9628_8799.n162 a_n9628_8799.t44 2.82907
R23295 a_n9628_8799.n159 a_n9628_8799.t8 2.82907
R23296 a_n9628_8799.n159 a_n9628_8799.t15 2.82907
R23297 a_n9628_8799.n158 a_n9628_8799.t0 2.82907
R23298 a_n9628_8799.n158 a_n9628_8799.t17 2.82907
R23299 a_n9628_8799.n157 a_n9628_8799.t12 2.82907
R23300 a_n9628_8799.n157 a_n9628_8799.t2 2.82907
R23301 a_n9628_8799.n1 a_n9628_8799.n2 2.12119
R23302 a_n9628_8799.n0 a_n9628_8799.n3 1.59102
R23303 a_n9628_8799.n45 a_n9628_8799.n44 1.13686
R23304 a_n9628_8799.n37 a_n9628_8799.n36 1.13686
R23305 a_n9628_8799.n29 a_n9628_8799.n28 1.13686
R23306 a_n9628_8799.n21 a_n9628_8799.n20 1.13686
R23307 a_n9628_8799.n13 a_n9628_8799.n12 1.13686
R23308 a_n9628_8799.n5 a_n9628_8799.n4 1.13686
R23309 a_n9628_8799.n50 a_n9628_8799.n49 0.758076
R23310 a_n9628_8799.n50 a_n9628_8799.n48 0.758076
R23311 a_n9628_8799.n48 a_n9628_8799.n47 0.758076
R23312 a_n9628_8799.n47 a_n9628_8799.n46 0.758076
R23313 a_n9628_8799.n44 a_n9628_8799.n46 0.758076
R23314 a_n9628_8799.n42 a_n9628_8799.n41 0.758076
R23315 a_n9628_8799.n42 a_n9628_8799.n40 0.758076
R23316 a_n9628_8799.n40 a_n9628_8799.n39 0.758076
R23317 a_n9628_8799.n39 a_n9628_8799.n38 0.758076
R23318 a_n9628_8799.n36 a_n9628_8799.n38 0.758076
R23319 a_n9628_8799.n34 a_n9628_8799.n33 0.758076
R23320 a_n9628_8799.n34 a_n9628_8799.n32 0.758076
R23321 a_n9628_8799.n32 a_n9628_8799.n31 0.758076
R23322 a_n9628_8799.n31 a_n9628_8799.n30 0.758076
R23323 a_n9628_8799.n28 a_n9628_8799.n30 0.758076
R23324 a_n9628_8799.n25 a_n9628_8799.n26 0.758076
R23325 a_n9628_8799.n24 a_n9628_8799.n25 0.758076
R23326 a_n9628_8799.n23 a_n9628_8799.n24 0.758076
R23327 a_n9628_8799.n22 a_n9628_8799.n23 0.758076
R23328 a_n9628_8799.n20 a_n9628_8799.n22 0.758076
R23329 a_n9628_8799.n17 a_n9628_8799.n18 0.758076
R23330 a_n9628_8799.n16 a_n9628_8799.n17 0.758076
R23331 a_n9628_8799.n15 a_n9628_8799.n16 0.758076
R23332 a_n9628_8799.n14 a_n9628_8799.n15 0.758076
R23333 a_n9628_8799.n12 a_n9628_8799.n14 0.758076
R23334 a_n9628_8799.n9 a_n9628_8799.n10 0.758076
R23335 a_n9628_8799.n8 a_n9628_8799.n9 0.758076
R23336 a_n9628_8799.n7 a_n9628_8799.n8 0.758076
R23337 a_n9628_8799.n6 a_n9628_8799.n7 0.758076
R23338 a_n9628_8799.n4 a_n9628_8799.n6 0.758076
R23339 a_n9628_8799.n57 a_n9628_8799.n55 0.716017
R23340 a_n9628_8799.n57 a_n9628_8799.n56 0.716017
R23341 a_n9628_8799.n54 a_n9628_8799.n53 0.716017
R23342 a_n9628_8799.n53 a_n9628_8799.n52 0.716017
R23343 a_n9628_8799.n10 a_n9628_8799.n11 0.568682
R23344 a_n9628_8799.n18 a_n9628_8799.n19 0.568682
R23345 a_n9628_8799.n26 a_n9628_8799.n27 0.568682
R23346 a_n9628_8799.n33 a_n9628_8799.n35 0.568682
R23347 a_n9628_8799.n41 a_n9628_8799.n43 0.568682
R23348 a_n9628_8799.n49 a_n9628_8799.n51 0.568682
R23349 plus.n76 plus.t11 250.337
R23350 plus.n15 plus.t14 250.337
R23351 plus.n124 plus.t1 243.97
R23352 plus.n120 plus.t24 231.093
R23353 plus.n59 plus.t20 231.093
R23354 plus.n124 plus.n123 223.454
R23355 plus.n126 plus.n125 223.454
R23356 plus.n77 plus.t5 187.445
R23357 plus.n74 plus.t22 187.445
R23358 plus.n72 plus.t21 187.445
R23359 plus.n89 plus.t16 187.445
R23360 plus.n95 plus.t17 187.445
R23361 plus.n68 plus.t13 187.445
R23362 plus.n66 plus.t15 187.445
R23363 plus.n107 plus.t10 187.445
R23364 plus.n113 plus.t26 187.445
R23365 plus.n62 plus.t28 187.445
R23366 plus.n1 plus.t23 187.445
R23367 plus.n52 plus.t6 187.445
R23368 plus.n46 plus.t12 187.445
R23369 plus.n5 plus.t8 187.445
R23370 plus.n7 plus.t7 187.445
R23371 plus.n34 plus.t19 187.445
R23372 plus.n28 plus.t18 187.445
R23373 plus.n11 plus.t27 187.445
R23374 plus.n13 plus.t25 187.445
R23375 plus.n16 plus.t9 187.445
R23376 plus.n121 plus.n120 161.3
R23377 plus.n119 plus.n61 161.3
R23378 plus.n118 plus.n117 161.3
R23379 plus.n116 plus.n115 161.3
R23380 plus.n114 plus.n63 161.3
R23381 plus.n112 plus.n111 161.3
R23382 plus.n110 plus.n64 161.3
R23383 plus.n109 plus.n108 161.3
R23384 plus.n106 plus.n65 161.3
R23385 plus.n105 plus.n104 161.3
R23386 plus.n103 plus.n102 161.3
R23387 plus.n101 plus.n67 161.3
R23388 plus.n100 plus.n99 161.3
R23389 plus.n98 plus.n97 161.3
R23390 plus.n96 plus.n69 161.3
R23391 plus.n94 plus.n93 161.3
R23392 plus.n92 plus.n70 161.3
R23393 plus.n91 plus.n90 161.3
R23394 plus.n88 plus.n71 161.3
R23395 plus.n87 plus.n86 161.3
R23396 plus.n85 plus.n84 161.3
R23397 plus.n83 plus.n73 161.3
R23398 plus.n82 plus.n81 161.3
R23399 plus.n80 plus.n79 161.3
R23400 plus.n78 plus.n75 161.3
R23401 plus.n17 plus.n14 161.3
R23402 plus.n19 plus.n18 161.3
R23403 plus.n21 plus.n20 161.3
R23404 plus.n22 plus.n12 161.3
R23405 plus.n24 plus.n23 161.3
R23406 plus.n26 plus.n25 161.3
R23407 plus.n27 plus.n10 161.3
R23408 plus.n30 plus.n29 161.3
R23409 plus.n31 plus.n9 161.3
R23410 plus.n33 plus.n32 161.3
R23411 plus.n35 plus.n8 161.3
R23412 plus.n37 plus.n36 161.3
R23413 plus.n39 plus.n38 161.3
R23414 plus.n40 plus.n6 161.3
R23415 plus.n42 plus.n41 161.3
R23416 plus.n44 plus.n43 161.3
R23417 plus.n45 plus.n4 161.3
R23418 plus.n48 plus.n47 161.3
R23419 plus.n49 plus.n3 161.3
R23420 plus.n51 plus.n50 161.3
R23421 plus.n53 plus.n2 161.3
R23422 plus.n55 plus.n54 161.3
R23423 plus.n57 plus.n56 161.3
R23424 plus.n58 plus.n0 161.3
R23425 plus.n60 plus.n59 161.3
R23426 plus.n88 plus.n87 56.5617
R23427 plus.n97 plus.n96 56.5617
R23428 plus.n106 plus.n105 56.5617
R23429 plus.n45 plus.n44 56.5617
R23430 plus.n36 plus.n35 56.5617
R23431 plus.n27 plus.n26 56.5617
R23432 plus.n79 plus.n78 56.5617
R23433 plus.n115 plus.n114 56.5617
R23434 plus.n54 plus.n53 56.5617
R23435 plus.n18 plus.n17 56.5617
R23436 plus.n119 plus.n118 50.2647
R23437 plus.n58 plus.n57 50.2647
R23438 plus.n84 plus.n83 46.3896
R23439 plus.n108 plus.n64 46.3896
R23440 plus.n47 plus.n3 46.3896
R23441 plus.n23 plus.n22 46.3896
R23442 plus.n76 plus.n75 43.1929
R23443 plus.n15 plus.n14 43.1929
R23444 plus.n94 plus.n70 42.5146
R23445 plus.n101 plus.n100 42.5146
R23446 plus.n40 plus.n39 42.5146
R23447 plus.n33 plus.n9 42.5146
R23448 plus.n77 plus.n76 40.6041
R23449 plus.n16 plus.n15 40.6041
R23450 plus.n90 plus.n70 38.6395
R23451 plus.n102 plus.n101 38.6395
R23452 plus.n41 plus.n40 38.6395
R23453 plus.n29 plus.n9 38.6395
R23454 plus.n122 plus.n121 35.2031
R23455 plus.n83 plus.n82 34.7644
R23456 plus.n112 plus.n64 34.7644
R23457 plus.n51 plus.n3 34.7644
R23458 plus.n22 plus.n21 34.7644
R23459 plus.n79 plus.n74 21.8872
R23460 plus.n114 plus.n113 21.8872
R23461 plus.n53 plus.n52 21.8872
R23462 plus.n18 plus.n13 21.8872
R23463 plus.n89 plus.n88 19.9199
R23464 plus.n105 plus.n66 19.9199
R23465 plus.n44 plus.n5 19.9199
R23466 plus.n28 plus.n27 19.9199
R23467 plus.n123 plus.t2 19.8005
R23468 plus.n123 plus.t4 19.8005
R23469 plus.n125 plus.t3 19.8005
R23470 plus.n125 plus.t0 19.8005
R23471 plus.n96 plus.n95 17.9525
R23472 plus.n97 plus.n68 17.9525
R23473 plus.n36 plus.n7 17.9525
R23474 plus.n35 plus.n34 17.9525
R23475 plus.n87 plus.n72 15.9852
R23476 plus.n107 plus.n106 15.9852
R23477 plus.n46 plus.n45 15.9852
R23478 plus.n26 plus.n11 15.9852
R23479 plus plus.n127 14.8156
R23480 plus.n78 plus.n77 14.0178
R23481 plus.n115 plus.n62 14.0178
R23482 plus.n54 plus.n1 14.0178
R23483 plus.n17 plus.n16 14.0178
R23484 plus.n122 plus.n60 11.9342
R23485 plus.n118 plus.n62 10.575
R23486 plus.n57 plus.n1 10.575
R23487 plus.n120 plus.n119 9.49444
R23488 plus.n59 plus.n58 9.49444
R23489 plus.n84 plus.n72 8.60764
R23490 plus.n108 plus.n107 8.60764
R23491 plus.n47 plus.n46 8.60764
R23492 plus.n23 plus.n11 8.60764
R23493 plus.n95 plus.n94 6.6403
R23494 plus.n100 plus.n68 6.6403
R23495 plus.n39 plus.n7 6.6403
R23496 plus.n34 plus.n33 6.6403
R23497 plus.n127 plus.n126 5.40567
R23498 plus.n90 plus.n89 4.67295
R23499 plus.n102 plus.n66 4.67295
R23500 plus.n41 plus.n5 4.67295
R23501 plus.n29 plus.n28 4.67295
R23502 plus.n82 plus.n74 2.7056
R23503 plus.n113 plus.n112 2.7056
R23504 plus.n52 plus.n51 2.7056
R23505 plus.n21 plus.n13 2.7056
R23506 plus.n127 plus.n122 1.188
R23507 plus.n126 plus.n124 0.716017
R23508 plus.n80 plus.n75 0.189894
R23509 plus.n81 plus.n80 0.189894
R23510 plus.n81 plus.n73 0.189894
R23511 plus.n85 plus.n73 0.189894
R23512 plus.n86 plus.n85 0.189894
R23513 plus.n86 plus.n71 0.189894
R23514 plus.n91 plus.n71 0.189894
R23515 plus.n92 plus.n91 0.189894
R23516 plus.n93 plus.n92 0.189894
R23517 plus.n93 plus.n69 0.189894
R23518 plus.n98 plus.n69 0.189894
R23519 plus.n99 plus.n98 0.189894
R23520 plus.n99 plus.n67 0.189894
R23521 plus.n103 plus.n67 0.189894
R23522 plus.n104 plus.n103 0.189894
R23523 plus.n104 plus.n65 0.189894
R23524 plus.n109 plus.n65 0.189894
R23525 plus.n110 plus.n109 0.189894
R23526 plus.n111 plus.n110 0.189894
R23527 plus.n111 plus.n63 0.189894
R23528 plus.n116 plus.n63 0.189894
R23529 plus.n117 plus.n116 0.189894
R23530 plus.n117 plus.n61 0.189894
R23531 plus.n121 plus.n61 0.189894
R23532 plus.n60 plus.n0 0.189894
R23533 plus.n56 plus.n0 0.189894
R23534 plus.n56 plus.n55 0.189894
R23535 plus.n55 plus.n2 0.189894
R23536 plus.n50 plus.n2 0.189894
R23537 plus.n50 plus.n49 0.189894
R23538 plus.n49 plus.n48 0.189894
R23539 plus.n48 plus.n4 0.189894
R23540 plus.n43 plus.n4 0.189894
R23541 plus.n43 plus.n42 0.189894
R23542 plus.n42 plus.n6 0.189894
R23543 plus.n38 plus.n6 0.189894
R23544 plus.n38 plus.n37 0.189894
R23545 plus.n37 plus.n8 0.189894
R23546 plus.n32 plus.n8 0.189894
R23547 plus.n32 plus.n31 0.189894
R23548 plus.n31 plus.n30 0.189894
R23549 plus.n30 plus.n10 0.189894
R23550 plus.n25 plus.n10 0.189894
R23551 plus.n25 plus.n24 0.189894
R23552 plus.n24 plus.n12 0.189894
R23553 plus.n20 plus.n12 0.189894
R23554 plus.n20 plus.n19 0.189894
R23555 plus.n19 plus.n14 0.189894
R23556 a_n3106_n452.n33 a_n3106_n452.t24 214.321
R23557 a_n3106_n452.n32 a_n3106_n452.t26 214.321
R23558 a_n3106_n452.n31 a_n3106_n452.t17 214.321
R23559 a_n3106_n452.n30 a_n3106_n452.t30 214.321
R23560 a_n3106_n452.n29 a_n3106_n452.t27 214.321
R23561 a_n3106_n452.n28 a_n3106_n452.t2 214.321
R23562 a_n3106_n452.n27 a_n3106_n452.t15 214.321
R23563 a_n3106_n452.n26 a_n3106_n452.t0 214.321
R23564 a_n3106_n452.n12 a_n3106_n452.t49 55.8337
R23565 a_n3106_n452.n13 a_n3106_n452.t21 55.8337
R23566 a_n3106_n452.n24 a_n3106_n452.t29 55.8337
R23567 a_n3106_n452.n1 a_n3106_n452.t36 55.8335
R23568 a_n3106_n452.n35 a_n3106_n452.t22 55.8335
R23569 a_n3106_n452.n46 a_n3106_n452.t5 55.8335
R23570 a_n3106_n452.n47 a_n3106_n452.t46 55.8335
R23571 a_n3106_n452.n0 a_n3106_n452.t40 55.8335
R23572 a_n3106_n452.n57 a_n3106_n452.n56 53.0054
R23573 a_n3106_n452.n3 a_n3106_n452.n2 53.0052
R23574 a_n3106_n452.n5 a_n3106_n452.n4 53.0052
R23575 a_n3106_n452.n7 a_n3106_n452.n6 53.0052
R23576 a_n3106_n452.n9 a_n3106_n452.n8 53.0052
R23577 a_n3106_n452.n11 a_n3106_n452.n10 53.0052
R23578 a_n3106_n452.n15 a_n3106_n452.n14 53.0052
R23579 a_n3106_n452.n17 a_n3106_n452.n16 53.0052
R23580 a_n3106_n452.n19 a_n3106_n452.n18 53.0052
R23581 a_n3106_n452.n21 a_n3106_n452.n20 53.0052
R23582 a_n3106_n452.n23 a_n3106_n452.n22 53.0052
R23583 a_n3106_n452.n37 a_n3106_n452.n36 53.0051
R23584 a_n3106_n452.n39 a_n3106_n452.n38 53.0051
R23585 a_n3106_n452.n41 a_n3106_n452.n40 53.0051
R23586 a_n3106_n452.n43 a_n3106_n452.n42 53.0051
R23587 a_n3106_n452.n45 a_n3106_n452.n44 53.0051
R23588 a_n3106_n452.n49 a_n3106_n452.n48 53.0051
R23589 a_n3106_n452.n51 a_n3106_n452.n50 53.0051
R23590 a_n3106_n452.n53 a_n3106_n452.n52 53.0051
R23591 a_n3106_n452.n55 a_n3106_n452.n54 53.0051
R23592 a_n3106_n452.n25 a_n3106_n452.n24 12.2417
R23593 a_n3106_n452.n34 a_n3106_n452.n1 12.2417
R23594 a_n3106_n452.n25 a_n3106_n452.n0 5.16214
R23595 a_n3106_n452.n35 a_n3106_n452.n34 5.16214
R23596 a_n3106_n452.n36 a_n3106_n452.t25 2.82907
R23597 a_n3106_n452.n36 a_n3106_n452.t10 2.82907
R23598 a_n3106_n452.n38 a_n3106_n452.t6 2.82907
R23599 a_n3106_n452.n38 a_n3106_n452.t1 2.82907
R23600 a_n3106_n452.n40 a_n3106_n452.t14 2.82907
R23601 a_n3106_n452.n40 a_n3106_n452.t13 2.82907
R23602 a_n3106_n452.n42 a_n3106_n452.t31 2.82907
R23603 a_n3106_n452.n42 a_n3106_n452.t8 2.82907
R23604 a_n3106_n452.n44 a_n3106_n452.t9 2.82907
R23605 a_n3106_n452.n44 a_n3106_n452.t19 2.82907
R23606 a_n3106_n452.n48 a_n3106_n452.t35 2.82907
R23607 a_n3106_n452.n48 a_n3106_n452.t51 2.82907
R23608 a_n3106_n452.n50 a_n3106_n452.t42 2.82907
R23609 a_n3106_n452.n50 a_n3106_n452.t33 2.82907
R23610 a_n3106_n452.n52 a_n3106_n452.t53 2.82907
R23611 a_n3106_n452.n52 a_n3106_n452.t41 2.82907
R23612 a_n3106_n452.n54 a_n3106_n452.t48 2.82907
R23613 a_n3106_n452.n54 a_n3106_n452.t52 2.82907
R23614 a_n3106_n452.n2 a_n3106_n452.t34 2.82907
R23615 a_n3106_n452.n2 a_n3106_n452.t32 2.82907
R23616 a_n3106_n452.n4 a_n3106_n452.t45 2.82907
R23617 a_n3106_n452.n4 a_n3106_n452.t50 2.82907
R23618 a_n3106_n452.n6 a_n3106_n452.t43 2.82907
R23619 a_n3106_n452.n6 a_n3106_n452.t47 2.82907
R23620 a_n3106_n452.n8 a_n3106_n452.t39 2.82907
R23621 a_n3106_n452.n8 a_n3106_n452.t44 2.82907
R23622 a_n3106_n452.n10 a_n3106_n452.t55 2.82907
R23623 a_n3106_n452.n10 a_n3106_n452.t38 2.82907
R23624 a_n3106_n452.n14 a_n3106_n452.t12 2.82907
R23625 a_n3106_n452.n14 a_n3106_n452.t16 2.82907
R23626 a_n3106_n452.n16 a_n3106_n452.t7 2.82907
R23627 a_n3106_n452.n16 a_n3106_n452.t18 2.82907
R23628 a_n3106_n452.n18 a_n3106_n452.t4 2.82907
R23629 a_n3106_n452.n18 a_n3106_n452.t23 2.82907
R23630 a_n3106_n452.n20 a_n3106_n452.t28 2.82907
R23631 a_n3106_n452.n20 a_n3106_n452.t11 2.82907
R23632 a_n3106_n452.n22 a_n3106_n452.t3 2.82907
R23633 a_n3106_n452.n22 a_n3106_n452.t20 2.82907
R23634 a_n3106_n452.n57 a_n3106_n452.t37 2.82907
R23635 a_n3106_n452.t54 a_n3106_n452.n57 2.82907
R23636 a_n3106_n452.n34 a_n3106_n452.n33 2.54197
R23637 a_n3106_n452.n26 a_n3106_n452.n25 2.0129
R23638 a_n3106_n452.n27 a_n3106_n452.n26 0.672012
R23639 a_n3106_n452.n28 a_n3106_n452.n27 0.672012
R23640 a_n3106_n452.n29 a_n3106_n452.n28 0.672012
R23641 a_n3106_n452.n30 a_n3106_n452.n29 0.672012
R23642 a_n3106_n452.n31 a_n3106_n452.n30 0.672012
R23643 a_n3106_n452.n32 a_n3106_n452.n31 0.672012
R23644 a_n3106_n452.n33 a_n3106_n452.n32 0.672012
R23645 a_n3106_n452.n24 a_n3106_n452.n23 0.530672
R23646 a_n3106_n452.n23 a_n3106_n452.n21 0.530672
R23647 a_n3106_n452.n21 a_n3106_n452.n19 0.530672
R23648 a_n3106_n452.n19 a_n3106_n452.n17 0.530672
R23649 a_n3106_n452.n17 a_n3106_n452.n15 0.530672
R23650 a_n3106_n452.n15 a_n3106_n452.n13 0.530672
R23651 a_n3106_n452.n12 a_n3106_n452.n11 0.530672
R23652 a_n3106_n452.n11 a_n3106_n452.n9 0.530672
R23653 a_n3106_n452.n9 a_n3106_n452.n7 0.530672
R23654 a_n3106_n452.n7 a_n3106_n452.n5 0.530672
R23655 a_n3106_n452.n5 a_n3106_n452.n3 0.530672
R23656 a_n3106_n452.n3 a_n3106_n452.n1 0.530672
R23657 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R23658 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R23659 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R23660 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R23661 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R23662 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R23663 a_n3106_n452.n46 a_n3106_n452.n45 0.530672
R23664 a_n3106_n452.n45 a_n3106_n452.n43 0.530672
R23665 a_n3106_n452.n43 a_n3106_n452.n41 0.530672
R23666 a_n3106_n452.n41 a_n3106_n452.n39 0.530672
R23667 a_n3106_n452.n39 a_n3106_n452.n37 0.530672
R23668 a_n3106_n452.n37 a_n3106_n452.n35 0.530672
R23669 a_n3106_n452.n13 a_n3106_n452.n12 0.235414
R23670 a_n3106_n452.n47 a_n3106_n452.n46 0.235414
R23671 a_n2982_8322.n28 a_n2982_8322.t20 74.6477
R23672 a_n2982_8322.n13 a_n2982_8322.t9 74.6477
R23673 a_n2982_8322.n1 a_n2982_8322.t35 74.6474
R23674 a_n2982_8322.n20 a_n2982_8322.t14 74.2899
R23675 a_n2982_8322.n10 a_n2982_8322.t15 74.2899
R23676 a_n2982_8322.n14 a_n2982_8322.t7 74.2899
R23677 a_n2982_8322.n15 a_n2982_8322.t10 74.2899
R23678 a_n2982_8322.n18 a_n2982_8322.t11 74.2899
R23679 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R23680 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R23681 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R23682 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R23683 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R23684 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R23685 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R23686 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R23687 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R23688 a_n2982_8322.n13 a_n2982_8322.n12 70.6783
R23689 a_n2982_8322.n17 a_n2982_8322.n16 70.6783
R23690 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R23691 a_n2982_8322.n20 a_n2982_8322.n19 24.9022
R23692 a_n2982_8322.n11 a_n2982_8322.t0 9.69161
R23693 a_n2982_8322.n19 a_n2982_8322.n18 8.38735
R23694 a_n2982_8322.n11 a_n2982_8322.n10 6.90998
R23695 a_n2982_8322.n19 a_n2982_8322.n11 5.3452
R23696 a_n2982_8322.n27 a_n2982_8322.t33 3.61217
R23697 a_n2982_8322.n27 a_n2982_8322.t29 3.61217
R23698 a_n2982_8322.n25 a_n2982_8322.t17 3.61217
R23699 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R23700 a_n2982_8322.n23 a_n2982_8322.t30 3.61217
R23701 a_n2982_8322.n23 a_n2982_8322.t23 3.61217
R23702 a_n2982_8322.n21 a_n2982_8322.t27 3.61217
R23703 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R23704 a_n2982_8322.n0 a_n2982_8322.t28 3.61217
R23705 a_n2982_8322.n0 a_n2982_8322.t24 3.61217
R23706 a_n2982_8322.n2 a_n2982_8322.t21 3.61217
R23707 a_n2982_8322.n2 a_n2982_8322.t37 3.61217
R23708 a_n2982_8322.n4 a_n2982_8322.t34 3.61217
R23709 a_n2982_8322.n4 a_n2982_8322.t22 3.61217
R23710 a_n2982_8322.n6 a_n2982_8322.t19 3.61217
R23711 a_n2982_8322.n6 a_n2982_8322.t18 3.61217
R23712 a_n2982_8322.n8 a_n2982_8322.t32 3.61217
R23713 a_n2982_8322.n8 a_n2982_8322.t31 3.61217
R23714 a_n2982_8322.n12 a_n2982_8322.t13 3.61217
R23715 a_n2982_8322.n12 a_n2982_8322.t12 3.61217
R23716 a_n2982_8322.n16 a_n2982_8322.t8 3.61217
R23717 a_n2982_8322.n16 a_n2982_8322.t6 3.61217
R23718 a_n2982_8322.t36 a_n2982_8322.n30 3.61217
R23719 a_n2982_8322.n30 a_n2982_8322.t26 3.61217
R23720 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R23721 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R23722 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R23723 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R23724 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R23725 a_n2982_8322.n18 a_n2982_8322.n17 0.358259
R23726 a_n2982_8322.n17 a_n2982_8322.n15 0.358259
R23727 a_n2982_8322.n14 a_n2982_8322.n13 0.358259
R23728 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R23729 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R23730 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R23731 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R23732 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R23733 a_n2982_8322.n15 a_n2982_8322.n14 0.101793
R23734 a_n2982_8322.t5 a_n2982_8322.t1 0.0788333
R23735 a_n2982_8322.t4 a_n2982_8322.t2 0.0788333
R23736 a_n2982_8322.t0 a_n2982_8322.t3 0.0788333
R23737 a_n2982_8322.t4 a_n2982_8322.t5 0.0318333
R23738 a_n2982_8322.t0 a_n2982_8322.t2 0.0318333
R23739 a_n2982_8322.t1 a_n2982_8322.t2 0.0318333
R23740 a_n2982_8322.t3 a_n2982_8322.t4 0.0318333
R23741 output.n41 output.n15 289.615
R23742 output.n72 output.n46 289.615
R23743 output.n104 output.n78 289.615
R23744 output.n136 output.n110 289.615
R23745 output.n77 output.n45 197.26
R23746 output.n77 output.n76 196.298
R23747 output.n109 output.n108 196.298
R23748 output.n141 output.n140 196.298
R23749 output.n42 output.n41 185
R23750 output.n40 output.n39 185
R23751 output.n19 output.n18 185
R23752 output.n34 output.n33 185
R23753 output.n32 output.n31 185
R23754 output.n23 output.n22 185
R23755 output.n26 output.n25 185
R23756 output.n73 output.n72 185
R23757 output.n71 output.n70 185
R23758 output.n50 output.n49 185
R23759 output.n65 output.n64 185
R23760 output.n63 output.n62 185
R23761 output.n54 output.n53 185
R23762 output.n57 output.n56 185
R23763 output.n105 output.n104 185
R23764 output.n103 output.n102 185
R23765 output.n82 output.n81 185
R23766 output.n97 output.n96 185
R23767 output.n95 output.n94 185
R23768 output.n86 output.n85 185
R23769 output.n89 output.n88 185
R23770 output.n137 output.n136 185
R23771 output.n135 output.n134 185
R23772 output.n114 output.n113 185
R23773 output.n129 output.n128 185
R23774 output.n127 output.n126 185
R23775 output.n118 output.n117 185
R23776 output.n121 output.n120 185
R23777 output.t0 output.n24 147.661
R23778 output.t19 output.n55 147.661
R23779 output.t17 output.n87 147.661
R23780 output.t18 output.n119 147.661
R23781 output.n41 output.n40 104.615
R23782 output.n40 output.n18 104.615
R23783 output.n33 output.n18 104.615
R23784 output.n33 output.n32 104.615
R23785 output.n32 output.n22 104.615
R23786 output.n25 output.n22 104.615
R23787 output.n72 output.n71 104.615
R23788 output.n71 output.n49 104.615
R23789 output.n64 output.n49 104.615
R23790 output.n64 output.n63 104.615
R23791 output.n63 output.n53 104.615
R23792 output.n56 output.n53 104.615
R23793 output.n104 output.n103 104.615
R23794 output.n103 output.n81 104.615
R23795 output.n96 output.n81 104.615
R23796 output.n96 output.n95 104.615
R23797 output.n95 output.n85 104.615
R23798 output.n88 output.n85 104.615
R23799 output.n136 output.n135 104.615
R23800 output.n135 output.n113 104.615
R23801 output.n128 output.n113 104.615
R23802 output.n128 output.n127 104.615
R23803 output.n127 output.n117 104.615
R23804 output.n120 output.n117 104.615
R23805 output.n1 output.t14 77.056
R23806 output.n14 output.t16 76.6694
R23807 output.n1 output.n0 72.7095
R23808 output.n3 output.n2 72.7095
R23809 output.n5 output.n4 72.7095
R23810 output.n7 output.n6 72.7095
R23811 output.n9 output.n8 72.7095
R23812 output.n11 output.n10 72.7095
R23813 output.n13 output.n12 72.7095
R23814 output.n25 output.t0 52.3082
R23815 output.n56 output.t19 52.3082
R23816 output.n88 output.t17 52.3082
R23817 output.n120 output.t18 52.3082
R23818 output.n26 output.n24 15.6674
R23819 output.n57 output.n55 15.6674
R23820 output.n89 output.n87 15.6674
R23821 output.n121 output.n119 15.6674
R23822 output.n27 output.n23 12.8005
R23823 output.n58 output.n54 12.8005
R23824 output.n90 output.n86 12.8005
R23825 output.n122 output.n118 12.8005
R23826 output.n31 output.n30 12.0247
R23827 output.n62 output.n61 12.0247
R23828 output.n94 output.n93 12.0247
R23829 output.n126 output.n125 12.0247
R23830 output.n34 output.n21 11.249
R23831 output.n65 output.n52 11.249
R23832 output.n97 output.n84 11.249
R23833 output.n129 output.n116 11.249
R23834 output.n35 output.n19 10.4732
R23835 output.n66 output.n50 10.4732
R23836 output.n98 output.n82 10.4732
R23837 output.n130 output.n114 10.4732
R23838 output.n39 output.n38 9.69747
R23839 output.n70 output.n69 9.69747
R23840 output.n102 output.n101 9.69747
R23841 output.n134 output.n133 9.69747
R23842 output.n45 output.n44 9.45567
R23843 output.n76 output.n75 9.45567
R23844 output.n108 output.n107 9.45567
R23845 output.n140 output.n139 9.45567
R23846 output.n44 output.n43 9.3005
R23847 output.n17 output.n16 9.3005
R23848 output.n38 output.n37 9.3005
R23849 output.n36 output.n35 9.3005
R23850 output.n21 output.n20 9.3005
R23851 output.n30 output.n29 9.3005
R23852 output.n28 output.n27 9.3005
R23853 output.n75 output.n74 9.3005
R23854 output.n48 output.n47 9.3005
R23855 output.n69 output.n68 9.3005
R23856 output.n67 output.n66 9.3005
R23857 output.n52 output.n51 9.3005
R23858 output.n61 output.n60 9.3005
R23859 output.n59 output.n58 9.3005
R23860 output.n107 output.n106 9.3005
R23861 output.n80 output.n79 9.3005
R23862 output.n101 output.n100 9.3005
R23863 output.n99 output.n98 9.3005
R23864 output.n84 output.n83 9.3005
R23865 output.n93 output.n92 9.3005
R23866 output.n91 output.n90 9.3005
R23867 output.n139 output.n138 9.3005
R23868 output.n112 output.n111 9.3005
R23869 output.n133 output.n132 9.3005
R23870 output.n131 output.n130 9.3005
R23871 output.n116 output.n115 9.3005
R23872 output.n125 output.n124 9.3005
R23873 output.n123 output.n122 9.3005
R23874 output.n42 output.n17 8.92171
R23875 output.n73 output.n48 8.92171
R23876 output.n105 output.n80 8.92171
R23877 output.n137 output.n112 8.92171
R23878 output output.n141 8.15037
R23879 output.n43 output.n15 8.14595
R23880 output.n74 output.n46 8.14595
R23881 output.n106 output.n78 8.14595
R23882 output.n138 output.n110 8.14595
R23883 output.n45 output.n15 5.81868
R23884 output.n76 output.n46 5.81868
R23885 output.n108 output.n78 5.81868
R23886 output.n140 output.n110 5.81868
R23887 output.n43 output.n42 5.04292
R23888 output.n74 output.n73 5.04292
R23889 output.n106 output.n105 5.04292
R23890 output.n138 output.n137 5.04292
R23891 output.n28 output.n24 4.38594
R23892 output.n59 output.n55 4.38594
R23893 output.n91 output.n87 4.38594
R23894 output.n123 output.n119 4.38594
R23895 output.n39 output.n17 4.26717
R23896 output.n70 output.n48 4.26717
R23897 output.n102 output.n80 4.26717
R23898 output.n134 output.n112 4.26717
R23899 output.n0 output.t10 3.9605
R23900 output.n0 output.t8 3.9605
R23901 output.n2 output.t2 3.9605
R23902 output.n2 output.t4 3.9605
R23903 output.n4 output.t5 3.9605
R23904 output.n4 output.t12 3.9605
R23905 output.n6 output.t15 3.9605
R23906 output.n6 output.t3 3.9605
R23907 output.n8 output.t6 3.9605
R23908 output.n8 output.t11 3.9605
R23909 output.n10 output.t13 3.9605
R23910 output.n10 output.t1 3.9605
R23911 output.n12 output.t9 3.9605
R23912 output.n12 output.t7 3.9605
R23913 output.n38 output.n19 3.49141
R23914 output.n69 output.n50 3.49141
R23915 output.n101 output.n82 3.49141
R23916 output.n133 output.n114 3.49141
R23917 output.n35 output.n34 2.71565
R23918 output.n66 output.n65 2.71565
R23919 output.n98 output.n97 2.71565
R23920 output.n130 output.n129 2.71565
R23921 output.n31 output.n21 1.93989
R23922 output.n62 output.n52 1.93989
R23923 output.n94 output.n84 1.93989
R23924 output.n126 output.n116 1.93989
R23925 output.n30 output.n23 1.16414
R23926 output.n61 output.n54 1.16414
R23927 output.n93 output.n86 1.16414
R23928 output.n125 output.n118 1.16414
R23929 output.n141 output.n109 0.962709
R23930 output.n109 output.n77 0.962709
R23931 output.n27 output.n26 0.388379
R23932 output.n58 output.n57 0.388379
R23933 output.n90 output.n89 0.388379
R23934 output.n122 output.n121 0.388379
R23935 output.n14 output.n13 0.387128
R23936 output.n13 output.n11 0.387128
R23937 output.n11 output.n9 0.387128
R23938 output.n9 output.n7 0.387128
R23939 output.n7 output.n5 0.387128
R23940 output.n5 output.n3 0.387128
R23941 output.n3 output.n1 0.387128
R23942 output.n44 output.n16 0.155672
R23943 output.n37 output.n16 0.155672
R23944 output.n37 output.n36 0.155672
R23945 output.n36 output.n20 0.155672
R23946 output.n29 output.n20 0.155672
R23947 output.n29 output.n28 0.155672
R23948 output.n75 output.n47 0.155672
R23949 output.n68 output.n47 0.155672
R23950 output.n68 output.n67 0.155672
R23951 output.n67 output.n51 0.155672
R23952 output.n60 output.n51 0.155672
R23953 output.n60 output.n59 0.155672
R23954 output.n107 output.n79 0.155672
R23955 output.n100 output.n79 0.155672
R23956 output.n100 output.n99 0.155672
R23957 output.n99 output.n83 0.155672
R23958 output.n92 output.n83 0.155672
R23959 output.n92 output.n91 0.155672
R23960 output.n139 output.n111 0.155672
R23961 output.n132 output.n111 0.155672
R23962 output.n132 output.n131 0.155672
R23963 output.n131 output.n115 0.155672
R23964 output.n124 output.n115 0.155672
R23965 output.n124 output.n123 0.155672
R23966 output output.n14 0.126227
R23967 minus.n76 minus.t28 250.337
R23968 minus.n15 minus.t20 250.337
R23969 minus.n126 minus.t1 243.255
R23970 minus.n120 minus.t8 231.093
R23971 minus.n59 minus.t10 231.093
R23972 minus.n125 minus.n123 224.169
R23973 minus.n125 minus.n124 223.454
R23974 minus.n62 minus.t12 187.445
R23975 minus.n113 minus.t18 187.445
R23976 minus.n107 minus.t25 187.445
R23977 minus.n66 minus.t22 187.445
R23978 minus.n68 minus.t19 187.445
R23979 minus.n95 minus.t7 187.445
R23980 minus.n89 minus.t6 187.445
R23981 minus.n72 minus.t16 187.445
R23982 minus.n74 minus.t15 187.445
R23983 minus.n77 minus.t23 187.445
R23984 minus.n16 minus.t14 187.445
R23985 minus.n13 minus.t9 187.445
R23986 minus.n11 minus.t5 187.445
R23987 minus.n28 minus.t26 187.445
R23988 minus.n34 minus.t27 187.445
R23989 minus.n7 minus.t21 187.445
R23990 minus.n5 minus.t24 187.445
R23991 minus.n46 minus.t17 187.445
R23992 minus.n52 minus.t11 187.445
R23993 minus.n1 minus.t13 187.445
R23994 minus.n78 minus.n75 161.3
R23995 minus.n80 minus.n79 161.3
R23996 minus.n82 minus.n81 161.3
R23997 minus.n83 minus.n73 161.3
R23998 minus.n85 minus.n84 161.3
R23999 minus.n87 minus.n86 161.3
R24000 minus.n88 minus.n71 161.3
R24001 minus.n91 minus.n90 161.3
R24002 minus.n92 minus.n70 161.3
R24003 minus.n94 minus.n93 161.3
R24004 minus.n96 minus.n69 161.3
R24005 minus.n98 minus.n97 161.3
R24006 minus.n100 minus.n99 161.3
R24007 minus.n101 minus.n67 161.3
R24008 minus.n103 minus.n102 161.3
R24009 minus.n105 minus.n104 161.3
R24010 minus.n106 minus.n65 161.3
R24011 minus.n109 minus.n108 161.3
R24012 minus.n110 minus.n64 161.3
R24013 minus.n112 minus.n111 161.3
R24014 minus.n114 minus.n63 161.3
R24015 minus.n116 minus.n115 161.3
R24016 minus.n118 minus.n117 161.3
R24017 minus.n119 minus.n61 161.3
R24018 minus.n121 minus.n120 161.3
R24019 minus.n60 minus.n59 161.3
R24020 minus.n58 minus.n0 161.3
R24021 minus.n57 minus.n56 161.3
R24022 minus.n55 minus.n54 161.3
R24023 minus.n53 minus.n2 161.3
R24024 minus.n51 minus.n50 161.3
R24025 minus.n49 minus.n3 161.3
R24026 minus.n48 minus.n47 161.3
R24027 minus.n45 minus.n4 161.3
R24028 minus.n44 minus.n43 161.3
R24029 minus.n42 minus.n41 161.3
R24030 minus.n40 minus.n6 161.3
R24031 minus.n39 minus.n38 161.3
R24032 minus.n37 minus.n36 161.3
R24033 minus.n35 minus.n8 161.3
R24034 minus.n33 minus.n32 161.3
R24035 minus.n31 minus.n9 161.3
R24036 minus.n30 minus.n29 161.3
R24037 minus.n27 minus.n10 161.3
R24038 minus.n26 minus.n25 161.3
R24039 minus.n24 minus.n23 161.3
R24040 minus.n22 minus.n12 161.3
R24041 minus.n21 minus.n20 161.3
R24042 minus.n19 minus.n18 161.3
R24043 minus.n17 minus.n14 161.3
R24044 minus.n106 minus.n105 56.5617
R24045 minus.n97 minus.n96 56.5617
R24046 minus.n88 minus.n87 56.5617
R24047 minus.n27 minus.n26 56.5617
R24048 minus.n36 minus.n35 56.5617
R24049 minus.n45 minus.n44 56.5617
R24050 minus.n115 minus.n114 56.5617
R24051 minus.n79 minus.n78 56.5617
R24052 minus.n18 minus.n17 56.5617
R24053 minus.n54 minus.n53 56.5617
R24054 minus.n119 minus.n118 50.2647
R24055 minus.n58 minus.n57 50.2647
R24056 minus.n108 minus.n64 46.3896
R24057 minus.n84 minus.n83 46.3896
R24058 minus.n23 minus.n22 46.3896
R24059 minus.n47 minus.n3 46.3896
R24060 minus.n76 minus.n75 43.1929
R24061 minus.n15 minus.n14 43.1929
R24062 minus.n101 minus.n100 42.5146
R24063 minus.n94 minus.n70 42.5146
R24064 minus.n33 minus.n9 42.5146
R24065 minus.n40 minus.n39 42.5146
R24066 minus.n77 minus.n76 40.6041
R24067 minus.n16 minus.n15 40.6041
R24068 minus.n102 minus.n101 38.6395
R24069 minus.n90 minus.n70 38.6395
R24070 minus.n29 minus.n9 38.6395
R24071 minus.n41 minus.n40 38.6395
R24072 minus.n122 minus.n121 35.4191
R24073 minus.n112 minus.n64 34.7644
R24074 minus.n83 minus.n82 34.7644
R24075 minus.n22 minus.n21 34.7644
R24076 minus.n51 minus.n3 34.7644
R24077 minus.n114 minus.n113 21.8872
R24078 minus.n79 minus.n74 21.8872
R24079 minus.n18 minus.n13 21.8872
R24080 minus.n53 minus.n52 21.8872
R24081 minus.n105 minus.n66 19.9199
R24082 minus.n89 minus.n88 19.9199
R24083 minus.n28 minus.n27 19.9199
R24084 minus.n44 minus.n5 19.9199
R24085 minus.n124 minus.t0 19.8005
R24086 minus.n124 minus.t2 19.8005
R24087 minus.n123 minus.t4 19.8005
R24088 minus.n123 minus.t3 19.8005
R24089 minus.n97 minus.n68 17.9525
R24090 minus.n96 minus.n95 17.9525
R24091 minus.n35 minus.n34 17.9525
R24092 minus.n36 minus.n7 17.9525
R24093 minus.n107 minus.n106 15.9852
R24094 minus.n87 minus.n72 15.9852
R24095 minus.n26 minus.n11 15.9852
R24096 minus.n46 minus.n45 15.9852
R24097 minus.n115 minus.n62 14.0178
R24098 minus.n78 minus.n77 14.0178
R24099 minus.n17 minus.n16 14.0178
R24100 minus.n54 minus.n1 14.0178
R24101 minus.n122 minus.n60 12.1501
R24102 minus minus.n127 11.3284
R24103 minus.n118 minus.n62 10.575
R24104 minus.n57 minus.n1 10.575
R24105 minus.n120 minus.n119 9.49444
R24106 minus.n59 minus.n58 9.49444
R24107 minus.n108 minus.n107 8.60764
R24108 minus.n84 minus.n72 8.60764
R24109 minus.n23 minus.n11 8.60764
R24110 minus.n47 minus.n46 8.60764
R24111 minus.n100 minus.n68 6.6403
R24112 minus.n95 minus.n94 6.6403
R24113 minus.n34 minus.n33 6.6403
R24114 minus.n39 minus.n7 6.6403
R24115 minus.n127 minus.n126 4.80222
R24116 minus.n102 minus.n66 4.67295
R24117 minus.n90 minus.n89 4.67295
R24118 minus.n29 minus.n28 4.67295
R24119 minus.n41 minus.n5 4.67295
R24120 minus.n113 minus.n112 2.7056
R24121 minus.n82 minus.n74 2.7056
R24122 minus.n21 minus.n13 2.7056
R24123 minus.n52 minus.n51 2.7056
R24124 minus.n127 minus.n122 0.972091
R24125 minus.n126 minus.n125 0.716017
R24126 minus.n121 minus.n61 0.189894
R24127 minus.n117 minus.n61 0.189894
R24128 minus.n117 minus.n116 0.189894
R24129 minus.n116 minus.n63 0.189894
R24130 minus.n111 minus.n63 0.189894
R24131 minus.n111 minus.n110 0.189894
R24132 minus.n110 minus.n109 0.189894
R24133 minus.n109 minus.n65 0.189894
R24134 minus.n104 minus.n65 0.189894
R24135 minus.n104 minus.n103 0.189894
R24136 minus.n103 minus.n67 0.189894
R24137 minus.n99 minus.n67 0.189894
R24138 minus.n99 minus.n98 0.189894
R24139 minus.n98 minus.n69 0.189894
R24140 minus.n93 minus.n69 0.189894
R24141 minus.n93 minus.n92 0.189894
R24142 minus.n92 minus.n91 0.189894
R24143 minus.n91 minus.n71 0.189894
R24144 minus.n86 minus.n71 0.189894
R24145 minus.n86 minus.n85 0.189894
R24146 minus.n85 minus.n73 0.189894
R24147 minus.n81 minus.n73 0.189894
R24148 minus.n81 minus.n80 0.189894
R24149 minus.n80 minus.n75 0.189894
R24150 minus.n19 minus.n14 0.189894
R24151 minus.n20 minus.n19 0.189894
R24152 minus.n20 minus.n12 0.189894
R24153 minus.n24 minus.n12 0.189894
R24154 minus.n25 minus.n24 0.189894
R24155 minus.n25 minus.n10 0.189894
R24156 minus.n30 minus.n10 0.189894
R24157 minus.n31 minus.n30 0.189894
R24158 minus.n32 minus.n31 0.189894
R24159 minus.n32 minus.n8 0.189894
R24160 minus.n37 minus.n8 0.189894
R24161 minus.n38 minus.n37 0.189894
R24162 minus.n38 minus.n6 0.189894
R24163 minus.n42 minus.n6 0.189894
R24164 minus.n43 minus.n42 0.189894
R24165 minus.n43 minus.n4 0.189894
R24166 minus.n48 minus.n4 0.189894
R24167 minus.n49 minus.n48 0.189894
R24168 minus.n50 minus.n49 0.189894
R24169 minus.n50 minus.n2 0.189894
R24170 minus.n55 minus.n2 0.189894
R24171 minus.n56 minus.n55 0.189894
R24172 minus.n56 minus.n0 0.189894
R24173 minus.n60 minus.n0 0.189894
R24174 diffpairibias.n0 diffpairibias.t18 436.822
R24175 diffpairibias.n21 diffpairibias.t19 435.479
R24176 diffpairibias.n20 diffpairibias.t16 435.479
R24177 diffpairibias.n19 diffpairibias.t17 435.479
R24178 diffpairibias.n18 diffpairibias.t21 435.479
R24179 diffpairibias.n0 diffpairibias.t22 435.479
R24180 diffpairibias.n1 diffpairibias.t20 435.479
R24181 diffpairibias.n2 diffpairibias.t23 435.479
R24182 diffpairibias.n10 diffpairibias.t0 377.536
R24183 diffpairibias.n10 diffpairibias.t8 376.193
R24184 diffpairibias.n11 diffpairibias.t10 376.193
R24185 diffpairibias.n12 diffpairibias.t6 376.193
R24186 diffpairibias.n13 diffpairibias.t2 376.193
R24187 diffpairibias.n14 diffpairibias.t12 376.193
R24188 diffpairibias.n15 diffpairibias.t4 376.193
R24189 diffpairibias.n16 diffpairibias.t14 376.193
R24190 diffpairibias.n3 diffpairibias.t1 113.368
R24191 diffpairibias.n3 diffpairibias.t9 112.698
R24192 diffpairibias.n4 diffpairibias.t11 112.698
R24193 diffpairibias.n5 diffpairibias.t7 112.698
R24194 diffpairibias.n6 diffpairibias.t3 112.698
R24195 diffpairibias.n7 diffpairibias.t13 112.698
R24196 diffpairibias.n8 diffpairibias.t5 112.698
R24197 diffpairibias.n9 diffpairibias.t15 112.698
R24198 diffpairibias.n17 diffpairibias.n16 4.77242
R24199 diffpairibias.n17 diffpairibias.n9 4.30807
R24200 diffpairibias.n18 diffpairibias.n17 4.13945
R24201 diffpairibias.n16 diffpairibias.n15 1.34352
R24202 diffpairibias.n15 diffpairibias.n14 1.34352
R24203 diffpairibias.n14 diffpairibias.n13 1.34352
R24204 diffpairibias.n13 diffpairibias.n12 1.34352
R24205 diffpairibias.n12 diffpairibias.n11 1.34352
R24206 diffpairibias.n11 diffpairibias.n10 1.34352
R24207 diffpairibias.n2 diffpairibias.n1 1.34352
R24208 diffpairibias.n1 diffpairibias.n0 1.34352
R24209 diffpairibias.n19 diffpairibias.n18 1.34352
R24210 diffpairibias.n20 diffpairibias.n19 1.34352
R24211 diffpairibias.n21 diffpairibias.n20 1.34352
R24212 diffpairibias.n22 diffpairibias.n21 0.862419
R24213 diffpairibias diffpairibias.n22 0.684875
R24214 diffpairibias.n9 diffpairibias.n8 0.672012
R24215 diffpairibias.n8 diffpairibias.n7 0.672012
R24216 diffpairibias.n7 diffpairibias.n6 0.672012
R24217 diffpairibias.n6 diffpairibias.n5 0.672012
R24218 diffpairibias.n5 diffpairibias.n4 0.672012
R24219 diffpairibias.n4 diffpairibias.n3 0.672012
R24220 diffpairibias.n22 diffpairibias.n2 0.190907
R24221 outputibias.n27 outputibias.n1 289.615
R24222 outputibias.n58 outputibias.n32 289.615
R24223 outputibias.n90 outputibias.n64 289.615
R24224 outputibias.n122 outputibias.n96 289.615
R24225 outputibias.n28 outputibias.n27 185
R24226 outputibias.n26 outputibias.n25 185
R24227 outputibias.n5 outputibias.n4 185
R24228 outputibias.n20 outputibias.n19 185
R24229 outputibias.n18 outputibias.n17 185
R24230 outputibias.n9 outputibias.n8 185
R24231 outputibias.n12 outputibias.n11 185
R24232 outputibias.n59 outputibias.n58 185
R24233 outputibias.n57 outputibias.n56 185
R24234 outputibias.n36 outputibias.n35 185
R24235 outputibias.n51 outputibias.n50 185
R24236 outputibias.n49 outputibias.n48 185
R24237 outputibias.n40 outputibias.n39 185
R24238 outputibias.n43 outputibias.n42 185
R24239 outputibias.n91 outputibias.n90 185
R24240 outputibias.n89 outputibias.n88 185
R24241 outputibias.n68 outputibias.n67 185
R24242 outputibias.n83 outputibias.n82 185
R24243 outputibias.n81 outputibias.n80 185
R24244 outputibias.n72 outputibias.n71 185
R24245 outputibias.n75 outputibias.n74 185
R24246 outputibias.n123 outputibias.n122 185
R24247 outputibias.n121 outputibias.n120 185
R24248 outputibias.n100 outputibias.n99 185
R24249 outputibias.n115 outputibias.n114 185
R24250 outputibias.n113 outputibias.n112 185
R24251 outputibias.n104 outputibias.n103 185
R24252 outputibias.n107 outputibias.n106 185
R24253 outputibias.n0 outputibias.t10 178.945
R24254 outputibias.n133 outputibias.t8 177.018
R24255 outputibias.n132 outputibias.t11 177.018
R24256 outputibias.n0 outputibias.t9 177.018
R24257 outputibias.t7 outputibias.n10 147.661
R24258 outputibias.t3 outputibias.n41 147.661
R24259 outputibias.t1 outputibias.n73 147.661
R24260 outputibias.t5 outputibias.n105 147.661
R24261 outputibias.n128 outputibias.t6 132.363
R24262 outputibias.n128 outputibias.t2 130.436
R24263 outputibias.n129 outputibias.t0 130.436
R24264 outputibias.n130 outputibias.t4 130.436
R24265 outputibias.n27 outputibias.n26 104.615
R24266 outputibias.n26 outputibias.n4 104.615
R24267 outputibias.n19 outputibias.n4 104.615
R24268 outputibias.n19 outputibias.n18 104.615
R24269 outputibias.n18 outputibias.n8 104.615
R24270 outputibias.n11 outputibias.n8 104.615
R24271 outputibias.n58 outputibias.n57 104.615
R24272 outputibias.n57 outputibias.n35 104.615
R24273 outputibias.n50 outputibias.n35 104.615
R24274 outputibias.n50 outputibias.n49 104.615
R24275 outputibias.n49 outputibias.n39 104.615
R24276 outputibias.n42 outputibias.n39 104.615
R24277 outputibias.n90 outputibias.n89 104.615
R24278 outputibias.n89 outputibias.n67 104.615
R24279 outputibias.n82 outputibias.n67 104.615
R24280 outputibias.n82 outputibias.n81 104.615
R24281 outputibias.n81 outputibias.n71 104.615
R24282 outputibias.n74 outputibias.n71 104.615
R24283 outputibias.n122 outputibias.n121 104.615
R24284 outputibias.n121 outputibias.n99 104.615
R24285 outputibias.n114 outputibias.n99 104.615
R24286 outputibias.n114 outputibias.n113 104.615
R24287 outputibias.n113 outputibias.n103 104.615
R24288 outputibias.n106 outputibias.n103 104.615
R24289 outputibias.n63 outputibias.n31 95.6354
R24290 outputibias.n63 outputibias.n62 94.6732
R24291 outputibias.n95 outputibias.n94 94.6732
R24292 outputibias.n127 outputibias.n126 94.6732
R24293 outputibias.n11 outputibias.t7 52.3082
R24294 outputibias.n42 outputibias.t3 52.3082
R24295 outputibias.n74 outputibias.t1 52.3082
R24296 outputibias.n106 outputibias.t5 52.3082
R24297 outputibias.n12 outputibias.n10 15.6674
R24298 outputibias.n43 outputibias.n41 15.6674
R24299 outputibias.n75 outputibias.n73 15.6674
R24300 outputibias.n107 outputibias.n105 15.6674
R24301 outputibias.n13 outputibias.n9 12.8005
R24302 outputibias.n44 outputibias.n40 12.8005
R24303 outputibias.n76 outputibias.n72 12.8005
R24304 outputibias.n108 outputibias.n104 12.8005
R24305 outputibias.n17 outputibias.n16 12.0247
R24306 outputibias.n48 outputibias.n47 12.0247
R24307 outputibias.n80 outputibias.n79 12.0247
R24308 outputibias.n112 outputibias.n111 12.0247
R24309 outputibias.n20 outputibias.n7 11.249
R24310 outputibias.n51 outputibias.n38 11.249
R24311 outputibias.n83 outputibias.n70 11.249
R24312 outputibias.n115 outputibias.n102 11.249
R24313 outputibias.n21 outputibias.n5 10.4732
R24314 outputibias.n52 outputibias.n36 10.4732
R24315 outputibias.n84 outputibias.n68 10.4732
R24316 outputibias.n116 outputibias.n100 10.4732
R24317 outputibias.n25 outputibias.n24 9.69747
R24318 outputibias.n56 outputibias.n55 9.69747
R24319 outputibias.n88 outputibias.n87 9.69747
R24320 outputibias.n120 outputibias.n119 9.69747
R24321 outputibias.n31 outputibias.n30 9.45567
R24322 outputibias.n62 outputibias.n61 9.45567
R24323 outputibias.n94 outputibias.n93 9.45567
R24324 outputibias.n126 outputibias.n125 9.45567
R24325 outputibias.n30 outputibias.n29 9.3005
R24326 outputibias.n3 outputibias.n2 9.3005
R24327 outputibias.n24 outputibias.n23 9.3005
R24328 outputibias.n22 outputibias.n21 9.3005
R24329 outputibias.n7 outputibias.n6 9.3005
R24330 outputibias.n16 outputibias.n15 9.3005
R24331 outputibias.n14 outputibias.n13 9.3005
R24332 outputibias.n61 outputibias.n60 9.3005
R24333 outputibias.n34 outputibias.n33 9.3005
R24334 outputibias.n55 outputibias.n54 9.3005
R24335 outputibias.n53 outputibias.n52 9.3005
R24336 outputibias.n38 outputibias.n37 9.3005
R24337 outputibias.n47 outputibias.n46 9.3005
R24338 outputibias.n45 outputibias.n44 9.3005
R24339 outputibias.n93 outputibias.n92 9.3005
R24340 outputibias.n66 outputibias.n65 9.3005
R24341 outputibias.n87 outputibias.n86 9.3005
R24342 outputibias.n85 outputibias.n84 9.3005
R24343 outputibias.n70 outputibias.n69 9.3005
R24344 outputibias.n79 outputibias.n78 9.3005
R24345 outputibias.n77 outputibias.n76 9.3005
R24346 outputibias.n125 outputibias.n124 9.3005
R24347 outputibias.n98 outputibias.n97 9.3005
R24348 outputibias.n119 outputibias.n118 9.3005
R24349 outputibias.n117 outputibias.n116 9.3005
R24350 outputibias.n102 outputibias.n101 9.3005
R24351 outputibias.n111 outputibias.n110 9.3005
R24352 outputibias.n109 outputibias.n108 9.3005
R24353 outputibias.n28 outputibias.n3 8.92171
R24354 outputibias.n59 outputibias.n34 8.92171
R24355 outputibias.n91 outputibias.n66 8.92171
R24356 outputibias.n123 outputibias.n98 8.92171
R24357 outputibias.n29 outputibias.n1 8.14595
R24358 outputibias.n60 outputibias.n32 8.14595
R24359 outputibias.n92 outputibias.n64 8.14595
R24360 outputibias.n124 outputibias.n96 8.14595
R24361 outputibias.n31 outputibias.n1 5.81868
R24362 outputibias.n62 outputibias.n32 5.81868
R24363 outputibias.n94 outputibias.n64 5.81868
R24364 outputibias.n126 outputibias.n96 5.81868
R24365 outputibias.n131 outputibias.n130 5.20947
R24366 outputibias.n29 outputibias.n28 5.04292
R24367 outputibias.n60 outputibias.n59 5.04292
R24368 outputibias.n92 outputibias.n91 5.04292
R24369 outputibias.n124 outputibias.n123 5.04292
R24370 outputibias.n131 outputibias.n127 4.42209
R24371 outputibias.n14 outputibias.n10 4.38594
R24372 outputibias.n45 outputibias.n41 4.38594
R24373 outputibias.n77 outputibias.n73 4.38594
R24374 outputibias.n109 outputibias.n105 4.38594
R24375 outputibias.n132 outputibias.n131 4.28454
R24376 outputibias.n25 outputibias.n3 4.26717
R24377 outputibias.n56 outputibias.n34 4.26717
R24378 outputibias.n88 outputibias.n66 4.26717
R24379 outputibias.n120 outputibias.n98 4.26717
R24380 outputibias.n24 outputibias.n5 3.49141
R24381 outputibias.n55 outputibias.n36 3.49141
R24382 outputibias.n87 outputibias.n68 3.49141
R24383 outputibias.n119 outputibias.n100 3.49141
R24384 outputibias.n21 outputibias.n20 2.71565
R24385 outputibias.n52 outputibias.n51 2.71565
R24386 outputibias.n84 outputibias.n83 2.71565
R24387 outputibias.n116 outputibias.n115 2.71565
R24388 outputibias.n17 outputibias.n7 1.93989
R24389 outputibias.n48 outputibias.n38 1.93989
R24390 outputibias.n80 outputibias.n70 1.93989
R24391 outputibias.n112 outputibias.n102 1.93989
R24392 outputibias.n130 outputibias.n129 1.9266
R24393 outputibias.n129 outputibias.n128 1.9266
R24394 outputibias.n133 outputibias.n132 1.92658
R24395 outputibias.n134 outputibias.n133 1.29913
R24396 outputibias.n16 outputibias.n9 1.16414
R24397 outputibias.n47 outputibias.n40 1.16414
R24398 outputibias.n79 outputibias.n72 1.16414
R24399 outputibias.n111 outputibias.n104 1.16414
R24400 outputibias.n127 outputibias.n95 0.962709
R24401 outputibias.n95 outputibias.n63 0.962709
R24402 outputibias.n13 outputibias.n12 0.388379
R24403 outputibias.n44 outputibias.n43 0.388379
R24404 outputibias.n76 outputibias.n75 0.388379
R24405 outputibias.n108 outputibias.n107 0.388379
R24406 outputibias.n134 outputibias.n0 0.337251
R24407 outputibias outputibias.n134 0.302375
R24408 outputibias.n30 outputibias.n2 0.155672
R24409 outputibias.n23 outputibias.n2 0.155672
R24410 outputibias.n23 outputibias.n22 0.155672
R24411 outputibias.n22 outputibias.n6 0.155672
R24412 outputibias.n15 outputibias.n6 0.155672
R24413 outputibias.n15 outputibias.n14 0.155672
R24414 outputibias.n61 outputibias.n33 0.155672
R24415 outputibias.n54 outputibias.n33 0.155672
R24416 outputibias.n54 outputibias.n53 0.155672
R24417 outputibias.n53 outputibias.n37 0.155672
R24418 outputibias.n46 outputibias.n37 0.155672
R24419 outputibias.n46 outputibias.n45 0.155672
R24420 outputibias.n93 outputibias.n65 0.155672
R24421 outputibias.n86 outputibias.n65 0.155672
R24422 outputibias.n86 outputibias.n85 0.155672
R24423 outputibias.n85 outputibias.n69 0.155672
R24424 outputibias.n78 outputibias.n69 0.155672
R24425 outputibias.n78 outputibias.n77 0.155672
R24426 outputibias.n125 outputibias.n97 0.155672
R24427 outputibias.n118 outputibias.n97 0.155672
R24428 outputibias.n118 outputibias.n117 0.155672
R24429 outputibias.n117 outputibias.n101 0.155672
R24430 outputibias.n110 outputibias.n101 0.155672
R24431 outputibias.n110 outputibias.n109 0.155672
C0 vdd output 7.23429f
C1 CSoutput output 6.13881f
C2 CSoutput outputibias 0.032386f
C3 vdd CSoutput 0.14236p
C4 minus diffpairibias 5.39e-19
C5 commonsourceibias output 0.006829f
C6 CSoutput minus 2.59304f
C7 vdd plus 0.106505f
C8 commonsourceibias outputibias 0.003902f
C9 plus diffpairibias 4.4e-19
C10 vdd commonsourceibias 0.004262f
C11 CSoutput plus 0.899588f
C12 commonsourceibias diffpairibias 0.06482f
C13 CSoutput commonsourceibias 42.168602f
C14 minus plus 10.1452f
C15 minus commonsourceibias 0.515277f
C16 plus commonsourceibias 0.49873f
C17 output outputibias 2.34152f
C18 diffpairibias gnd 48.964737f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144169p
C22 plus gnd 38.6522f
C23 minus gnd 30.23477f
C24 CSoutput gnd 0.107452p
C25 vdd gnd 0.542244p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t3 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t2 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.031048f
C221 minus.t13 gnd 0.52206f
C222 minus.n1 gnd 0.211144f
C223 minus.n2 gnd 0.031048f
C224 minus.t11 gnd 0.52206f
C225 minus.n3 gnd 0.026531f
C226 minus.n4 gnd 0.031048f
C227 minus.t17 gnd 0.52206f
C228 minus.t24 gnd 0.52206f
C229 minus.n5 gnd 0.211144f
C230 minus.n6 gnd 0.031048f
C231 minus.t21 gnd 0.52206f
C232 minus.n7 gnd 0.211144f
C233 minus.n8 gnd 0.031048f
C234 minus.t27 gnd 0.52206f
C235 minus.n9 gnd 0.025235f
C236 minus.n10 gnd 0.031048f
C237 minus.t26 gnd 0.52206f
C238 minus.t5 gnd 0.52206f
C239 minus.n11 gnd 0.211144f
C240 minus.n12 gnd 0.031048f
C241 minus.t9 gnd 0.52206f
C242 minus.n13 gnd 0.211144f
C243 minus.n14 gnd 0.131763f
C244 minus.t14 gnd 0.52206f
C245 minus.t20 gnd 0.584019f
C246 minus.n15 gnd 0.246849f
C247 minus.n16 gnd 0.2418f
C248 minus.n17 gnd 0.039783f
C249 minus.n18 gnd 0.035134f
C250 minus.n19 gnd 0.031048f
C251 minus.n20 gnd 0.031048f
C252 minus.n21 gnd 0.037102f
C253 minus.n22 gnd 0.026531f
C254 minus.n23 gnd 0.040435f
C255 minus.n24 gnd 0.031048f
C256 minus.n25 gnd 0.031048f
C257 minus.n26 gnd 0.03862f
C258 minus.n27 gnd 0.036296f
C259 minus.n28 gnd 0.211144f
C260 minus.n29 gnd 0.038892f
C261 minus.n30 gnd 0.031048f
C262 minus.n31 gnd 0.031048f
C263 minus.n32 gnd 0.031048f
C264 minus.n33 gnd 0.039941f
C265 minus.n34 gnd 0.211144f
C266 minus.n35 gnd 0.037458f
C267 minus.n36 gnd 0.037458f
C268 minus.n37 gnd 0.031048f
C269 minus.n38 gnd 0.031048f
C270 minus.n39 gnd 0.039941f
C271 minus.n40 gnd 0.025235f
C272 minus.n41 gnd 0.038892f
C273 minus.n42 gnd 0.031048f
C274 minus.n43 gnd 0.031048f
C275 minus.n44 gnd 0.036296f
C276 minus.n45 gnd 0.03862f
C277 minus.n46 gnd 0.211144f
C278 minus.n47 gnd 0.040435f
C279 minus.n48 gnd 0.031048f
C280 minus.n49 gnd 0.031048f
C281 minus.n50 gnd 0.031048f
C282 minus.n51 gnd 0.037102f
C283 minus.n52 gnd 0.211144f
C284 minus.n53 gnd 0.035134f
C285 minus.n54 gnd 0.039783f
C286 minus.n55 gnd 0.031048f
C287 minus.n56 gnd 0.031048f
C288 minus.n57 gnd 0.040503f
C289 minus.n58 gnd 0.011284f
C290 minus.t10 gnd 0.564608f
C291 minus.n59 gnd 0.24447f
C292 minus.n60 gnd 0.36371f
C293 minus.n61 gnd 0.031048f
C294 minus.t8 gnd 0.564608f
C295 minus.t12 gnd 0.52206f
C296 minus.n62 gnd 0.211144f
C297 minus.n63 gnd 0.031048f
C298 minus.t18 gnd 0.52206f
C299 minus.n64 gnd 0.026531f
C300 minus.n65 gnd 0.031048f
C301 minus.t25 gnd 0.52206f
C302 minus.t22 gnd 0.52206f
C303 minus.n66 gnd 0.211144f
C304 minus.n67 gnd 0.031048f
C305 minus.t19 gnd 0.52206f
C306 minus.n68 gnd 0.211144f
C307 minus.n69 gnd 0.031048f
C308 minus.t7 gnd 0.52206f
C309 minus.n70 gnd 0.025235f
C310 minus.n71 gnd 0.031048f
C311 minus.t6 gnd 0.52206f
C312 minus.t16 gnd 0.52206f
C313 minus.n72 gnd 0.211144f
C314 minus.n73 gnd 0.031048f
C315 minus.t15 gnd 0.52206f
C316 minus.n74 gnd 0.211144f
C317 minus.n75 gnd 0.131763f
C318 minus.t23 gnd 0.52206f
C319 minus.t28 gnd 0.584019f
C320 minus.n76 gnd 0.246849f
C321 minus.n77 gnd 0.2418f
C322 minus.n78 gnd 0.039783f
C323 minus.n79 gnd 0.035134f
C324 minus.n80 gnd 0.031048f
C325 minus.n81 gnd 0.031048f
C326 minus.n82 gnd 0.037102f
C327 minus.n83 gnd 0.026531f
C328 minus.n84 gnd 0.040435f
C329 minus.n85 gnd 0.031048f
C330 minus.n86 gnd 0.031048f
C331 minus.n87 gnd 0.03862f
C332 minus.n88 gnd 0.036296f
C333 minus.n89 gnd 0.211144f
C334 minus.n90 gnd 0.038892f
C335 minus.n91 gnd 0.031048f
C336 minus.n92 gnd 0.031048f
C337 minus.n93 gnd 0.031048f
C338 minus.n94 gnd 0.039941f
C339 minus.n95 gnd 0.211144f
C340 minus.n96 gnd 0.037458f
C341 minus.n97 gnd 0.037458f
C342 minus.n98 gnd 0.031048f
C343 minus.n99 gnd 0.031048f
C344 minus.n100 gnd 0.039941f
C345 minus.n101 gnd 0.025235f
C346 minus.n102 gnd 0.038892f
C347 minus.n103 gnd 0.031048f
C348 minus.n104 gnd 0.031048f
C349 minus.n105 gnd 0.036296f
C350 minus.n106 gnd 0.03862f
C351 minus.n107 gnd 0.211144f
C352 minus.n108 gnd 0.040435f
C353 minus.n109 gnd 0.031048f
C354 minus.n110 gnd 0.031048f
C355 minus.n111 gnd 0.031048f
C356 minus.n112 gnd 0.037102f
C357 minus.n113 gnd 0.211144f
C358 minus.n114 gnd 0.035134f
C359 minus.n115 gnd 0.039783f
C360 minus.n116 gnd 0.031048f
C361 minus.n117 gnd 0.031048f
C362 minus.n118 gnd 0.040503f
C363 minus.n119 gnd 0.011284f
C364 minus.n120 gnd 0.24447f
C365 minus.n121 gnd 1.1326f
C366 minus.n122 gnd 1.66371f
C367 minus.t4 gnd 0.009571f
C368 minus.t3 gnd 0.009571f
C369 minus.n123 gnd 0.031472f
C370 minus.t0 gnd 0.009571f
C371 minus.t2 gnd 0.009571f
C372 minus.n124 gnd 0.031041f
C373 minus.n125 gnd 0.264918f
C374 minus.t1 gnd 0.053271f
C375 minus.n126 gnd 0.144563f
C376 minus.n127 gnd 1.81446f
C377 output.t14 gnd 0.464308f
C378 output.t10 gnd 0.044422f
C379 output.t8 gnd 0.044422f
C380 output.n0 gnd 0.364624f
C381 output.n1 gnd 0.614102f
C382 output.t2 gnd 0.044422f
C383 output.t4 gnd 0.044422f
C384 output.n2 gnd 0.364624f
C385 output.n3 gnd 0.350265f
C386 output.t5 gnd 0.044422f
C387 output.t12 gnd 0.044422f
C388 output.n4 gnd 0.364624f
C389 output.n5 gnd 0.350265f
C390 output.t15 gnd 0.044422f
C391 output.t3 gnd 0.044422f
C392 output.n6 gnd 0.364624f
C393 output.n7 gnd 0.350265f
C394 output.t6 gnd 0.044422f
C395 output.t11 gnd 0.044422f
C396 output.n8 gnd 0.364624f
C397 output.n9 gnd 0.350265f
C398 output.t13 gnd 0.044422f
C399 output.t1 gnd 0.044422f
C400 output.n10 gnd 0.364624f
C401 output.n11 gnd 0.350265f
C402 output.t9 gnd 0.044422f
C403 output.t7 gnd 0.044422f
C404 output.n12 gnd 0.364624f
C405 output.n13 gnd 0.350265f
C406 output.t16 gnd 0.462979f
C407 output.n14 gnd 0.28994f
C408 output.n15 gnd 0.015803f
C409 output.n16 gnd 0.011243f
C410 output.n17 gnd 0.006041f
C411 output.n18 gnd 0.01428f
C412 output.n19 gnd 0.006397f
C413 output.n20 gnd 0.011243f
C414 output.n21 gnd 0.006041f
C415 output.n22 gnd 0.01428f
C416 output.n23 gnd 0.006397f
C417 output.n24 gnd 0.048111f
C418 output.t0 gnd 0.023274f
C419 output.n25 gnd 0.01071f
C420 output.n26 gnd 0.008435f
C421 output.n27 gnd 0.006041f
C422 output.n28 gnd 0.267512f
C423 output.n29 gnd 0.011243f
C424 output.n30 gnd 0.006041f
C425 output.n31 gnd 0.006397f
C426 output.n32 gnd 0.01428f
C427 output.n33 gnd 0.01428f
C428 output.n34 gnd 0.006397f
C429 output.n35 gnd 0.006041f
C430 output.n36 gnd 0.011243f
C431 output.n37 gnd 0.011243f
C432 output.n38 gnd 0.006041f
C433 output.n39 gnd 0.006397f
C434 output.n40 gnd 0.01428f
C435 output.n41 gnd 0.030913f
C436 output.n42 gnd 0.006397f
C437 output.n43 gnd 0.006041f
C438 output.n44 gnd 0.025987f
C439 output.n45 gnd 0.097665f
C440 output.n46 gnd 0.015803f
C441 output.n47 gnd 0.011243f
C442 output.n48 gnd 0.006041f
C443 output.n49 gnd 0.01428f
C444 output.n50 gnd 0.006397f
C445 output.n51 gnd 0.011243f
C446 output.n52 gnd 0.006041f
C447 output.n53 gnd 0.01428f
C448 output.n54 gnd 0.006397f
C449 output.n55 gnd 0.048111f
C450 output.t19 gnd 0.023274f
C451 output.n56 gnd 0.01071f
C452 output.n57 gnd 0.008435f
C453 output.n58 gnd 0.006041f
C454 output.n59 gnd 0.267512f
C455 output.n60 gnd 0.011243f
C456 output.n61 gnd 0.006041f
C457 output.n62 gnd 0.006397f
C458 output.n63 gnd 0.01428f
C459 output.n64 gnd 0.01428f
C460 output.n65 gnd 0.006397f
C461 output.n66 gnd 0.006041f
C462 output.n67 gnd 0.011243f
C463 output.n68 gnd 0.011243f
C464 output.n69 gnd 0.006041f
C465 output.n70 gnd 0.006397f
C466 output.n71 gnd 0.01428f
C467 output.n72 gnd 0.030913f
C468 output.n73 gnd 0.006397f
C469 output.n74 gnd 0.006041f
C470 output.n75 gnd 0.025987f
C471 output.n76 gnd 0.09306f
C472 output.n77 gnd 1.65264f
C473 output.n78 gnd 0.015803f
C474 output.n79 gnd 0.011243f
C475 output.n80 gnd 0.006041f
C476 output.n81 gnd 0.01428f
C477 output.n82 gnd 0.006397f
C478 output.n83 gnd 0.011243f
C479 output.n84 gnd 0.006041f
C480 output.n85 gnd 0.01428f
C481 output.n86 gnd 0.006397f
C482 output.n87 gnd 0.048111f
C483 output.t17 gnd 0.023274f
C484 output.n88 gnd 0.01071f
C485 output.n89 gnd 0.008435f
C486 output.n90 gnd 0.006041f
C487 output.n91 gnd 0.267512f
C488 output.n92 gnd 0.011243f
C489 output.n93 gnd 0.006041f
C490 output.n94 gnd 0.006397f
C491 output.n95 gnd 0.01428f
C492 output.n96 gnd 0.01428f
C493 output.n97 gnd 0.006397f
C494 output.n98 gnd 0.006041f
C495 output.n99 gnd 0.011243f
C496 output.n100 gnd 0.011243f
C497 output.n101 gnd 0.006041f
C498 output.n102 gnd 0.006397f
C499 output.n103 gnd 0.01428f
C500 output.n104 gnd 0.030913f
C501 output.n105 gnd 0.006397f
C502 output.n106 gnd 0.006041f
C503 output.n107 gnd 0.025987f
C504 output.n108 gnd 0.09306f
C505 output.n109 gnd 0.713089f
C506 output.n110 gnd 0.015803f
C507 output.n111 gnd 0.011243f
C508 output.n112 gnd 0.006041f
C509 output.n113 gnd 0.01428f
C510 output.n114 gnd 0.006397f
C511 output.n115 gnd 0.011243f
C512 output.n116 gnd 0.006041f
C513 output.n117 gnd 0.01428f
C514 output.n118 gnd 0.006397f
C515 output.n119 gnd 0.048111f
C516 output.t18 gnd 0.023274f
C517 output.n120 gnd 0.01071f
C518 output.n121 gnd 0.008435f
C519 output.n122 gnd 0.006041f
C520 output.n123 gnd 0.267512f
C521 output.n124 gnd 0.011243f
C522 output.n125 gnd 0.006041f
C523 output.n126 gnd 0.006397f
C524 output.n127 gnd 0.01428f
C525 output.n128 gnd 0.01428f
C526 output.n129 gnd 0.006397f
C527 output.n130 gnd 0.006041f
C528 output.n131 gnd 0.011243f
C529 output.n132 gnd 0.011243f
C530 output.n133 gnd 0.006041f
C531 output.n134 gnd 0.006397f
C532 output.n135 gnd 0.01428f
C533 output.n136 gnd 0.030913f
C534 output.n137 gnd 0.006397f
C535 output.n138 gnd 0.006041f
C536 output.n139 gnd 0.025987f
C537 output.n140 gnd 0.09306f
C538 output.n141 gnd 1.67353f
C539 a_n2982_8322.t26 gnd 0.100161f
C540 a_n2982_8322.t2 gnd 20.7793f
C541 a_n2982_8322.t1 gnd 20.633598f
C542 a_n2982_8322.t5 gnd 20.633598f
C543 a_n2982_8322.t4 gnd 20.7793f
C544 a_n2982_8322.t3 gnd 20.633598f
C545 a_n2982_8322.t0 gnd 28.9697f
C546 a_n2982_8322.t35 gnd 0.937854f
C547 a_n2982_8322.t28 gnd 0.100161f
C548 a_n2982_8322.t24 gnd 0.100161f
C549 a_n2982_8322.n0 gnd 0.705534f
C550 a_n2982_8322.n1 gnd 0.788332f
C551 a_n2982_8322.t21 gnd 0.100161f
C552 a_n2982_8322.t37 gnd 0.100161f
C553 a_n2982_8322.n2 gnd 0.705534f
C554 a_n2982_8322.n3 gnd 0.40054f
C555 a_n2982_8322.t34 gnd 0.100161f
C556 a_n2982_8322.t22 gnd 0.100161f
C557 a_n2982_8322.n4 gnd 0.705534f
C558 a_n2982_8322.n5 gnd 0.40054f
C559 a_n2982_8322.t19 gnd 0.100161f
C560 a_n2982_8322.t18 gnd 0.100161f
C561 a_n2982_8322.n6 gnd 0.705534f
C562 a_n2982_8322.n7 gnd 0.40054f
C563 a_n2982_8322.t32 gnd 0.100161f
C564 a_n2982_8322.t31 gnd 0.100161f
C565 a_n2982_8322.n8 gnd 0.705534f
C566 a_n2982_8322.n9 gnd 0.40054f
C567 a_n2982_8322.t15 gnd 0.935989f
C568 a_n2982_8322.n10 gnd 1.11148f
C569 a_n2982_8322.n11 gnd 3.33814f
C570 a_n2982_8322.t9 gnd 0.937857f
C571 a_n2982_8322.t13 gnd 0.100161f
C572 a_n2982_8322.t12 gnd 0.100161f
C573 a_n2982_8322.n12 gnd 0.705534f
C574 a_n2982_8322.n13 gnd 0.78833f
C575 a_n2982_8322.t7 gnd 0.935989f
C576 a_n2982_8322.n14 gnd 0.396699f
C577 a_n2982_8322.t10 gnd 0.935989f
C578 a_n2982_8322.n15 gnd 0.396699f
C579 a_n2982_8322.t8 gnd 0.100161f
C580 a_n2982_8322.t6 gnd 0.100161f
C581 a_n2982_8322.n16 gnd 0.705534f
C582 a_n2982_8322.n17 gnd 0.40054f
C583 a_n2982_8322.t11 gnd 0.935989f
C584 a_n2982_8322.n18 gnd 1.47142f
C585 a_n2982_8322.n19 gnd 2.35138f
C586 a_n2982_8322.t14 gnd 0.935989f
C587 a_n2982_8322.n20 gnd 1.87142f
C588 a_n2982_8322.t27 gnd 0.100161f
C589 a_n2982_8322.t25 gnd 0.100161f
C590 a_n2982_8322.n21 gnd 0.705534f
C591 a_n2982_8322.n22 gnd 0.40054f
C592 a_n2982_8322.t30 gnd 0.100161f
C593 a_n2982_8322.t23 gnd 0.100161f
C594 a_n2982_8322.n23 gnd 0.705534f
C595 a_n2982_8322.n24 gnd 0.40054f
C596 a_n2982_8322.t17 gnd 0.100161f
C597 a_n2982_8322.t16 gnd 0.100161f
C598 a_n2982_8322.n25 gnd 0.705534f
C599 a_n2982_8322.n26 gnd 0.40054f
C600 a_n2982_8322.t20 gnd 0.937857f
C601 a_n2982_8322.t33 gnd 0.100161f
C602 a_n2982_8322.t29 gnd 0.100161f
C603 a_n2982_8322.n27 gnd 0.705534f
C604 a_n2982_8322.n28 gnd 0.78833f
C605 a_n2982_8322.n29 gnd 0.400539f
C606 a_n2982_8322.n30 gnd 0.705536f
C607 a_n2982_8322.t36 gnd 0.100161f
C608 a_n3106_n452.t37 gnd 0.10001f
C609 a_n3106_n452.t40 gnd 1.03941f
C610 a_n3106_n452.n0 gnd 0.645631f
C611 a_n3106_n452.t36 gnd 1.03941f
C612 a_n3106_n452.n1 gnd 0.972978f
C613 a_n3106_n452.t34 gnd 0.10001f
C614 a_n3106_n452.t32 gnd 0.10001f
C615 a_n3106_n452.n2 gnd 0.816794f
C616 a_n3106_n452.n3 gnd 0.411618f
C617 a_n3106_n452.t45 gnd 0.10001f
C618 a_n3106_n452.t50 gnd 0.10001f
C619 a_n3106_n452.n4 gnd 0.816794f
C620 a_n3106_n452.n5 gnd 0.411618f
C621 a_n3106_n452.t43 gnd 0.10001f
C622 a_n3106_n452.t47 gnd 0.10001f
C623 a_n3106_n452.n6 gnd 0.816794f
C624 a_n3106_n452.n7 gnd 0.411618f
C625 a_n3106_n452.t39 gnd 0.10001f
C626 a_n3106_n452.t44 gnd 0.10001f
C627 a_n3106_n452.n8 gnd 0.816794f
C628 a_n3106_n452.n9 gnd 0.411618f
C629 a_n3106_n452.t55 gnd 0.10001f
C630 a_n3106_n452.t38 gnd 0.10001f
C631 a_n3106_n452.n10 gnd 0.816794f
C632 a_n3106_n452.n11 gnd 0.411618f
C633 a_n3106_n452.t49 gnd 1.03942f
C634 a_n3106_n452.n12 gnd 0.392946f
C635 a_n3106_n452.t21 gnd 1.03942f
C636 a_n3106_n452.n13 gnd 0.392946f
C637 a_n3106_n452.t12 gnd 0.10001f
C638 a_n3106_n452.t16 gnd 0.10001f
C639 a_n3106_n452.n14 gnd 0.816794f
C640 a_n3106_n452.n15 gnd 0.411618f
C641 a_n3106_n452.t7 gnd 0.10001f
C642 a_n3106_n452.t18 gnd 0.10001f
C643 a_n3106_n452.n16 gnd 0.816794f
C644 a_n3106_n452.n17 gnd 0.411618f
C645 a_n3106_n452.t4 gnd 0.10001f
C646 a_n3106_n452.t23 gnd 0.10001f
C647 a_n3106_n452.n18 gnd 0.816794f
C648 a_n3106_n452.n19 gnd 0.411618f
C649 a_n3106_n452.t28 gnd 0.10001f
C650 a_n3106_n452.t11 gnd 0.10001f
C651 a_n3106_n452.n20 gnd 0.816794f
C652 a_n3106_n452.n21 gnd 0.411618f
C653 a_n3106_n452.t3 gnd 0.10001f
C654 a_n3106_n452.t20 gnd 0.10001f
C655 a_n3106_n452.n22 gnd 0.816794f
C656 a_n3106_n452.n23 gnd 0.411618f
C657 a_n3106_n452.t29 gnd 1.03942f
C658 a_n3106_n452.n24 gnd 0.972974f
C659 a_n3106_n452.n25 gnd 0.948418f
C660 a_n3106_n452.t0 gnd 1.29145f
C661 a_n3106_n452.n26 gnd 0.789472f
C662 a_n3106_n452.t15 gnd 1.29145f
C663 a_n3106_n452.n27 gnd 0.909591f
C664 a_n3106_n452.t2 gnd 1.29145f
C665 a_n3106_n452.n28 gnd 0.909591f
C666 a_n3106_n452.t27 gnd 1.29145f
C667 a_n3106_n452.n29 gnd 0.909591f
C668 a_n3106_n452.t30 gnd 1.29145f
C669 a_n3106_n452.n30 gnd 0.909591f
C670 a_n3106_n452.t17 gnd 1.29145f
C671 a_n3106_n452.n31 gnd 0.909591f
C672 a_n3106_n452.t26 gnd 1.29145f
C673 a_n3106_n452.n32 gnd 0.909591f
C674 a_n3106_n452.t24 gnd 1.29145f
C675 a_n3106_n452.n33 gnd 1.22854f
C676 a_n3106_n452.n34 gnd 1.05146f
C677 a_n3106_n452.t22 gnd 1.03941f
C678 a_n3106_n452.n35 gnd 0.645631f
C679 a_n3106_n452.t25 gnd 0.10001f
C680 a_n3106_n452.t10 gnd 0.10001f
C681 a_n3106_n452.n36 gnd 0.816793f
C682 a_n3106_n452.n37 gnd 0.411619f
C683 a_n3106_n452.t6 gnd 0.10001f
C684 a_n3106_n452.t1 gnd 0.10001f
C685 a_n3106_n452.n38 gnd 0.816793f
C686 a_n3106_n452.n39 gnd 0.411619f
C687 a_n3106_n452.t14 gnd 0.10001f
C688 a_n3106_n452.t13 gnd 0.10001f
C689 a_n3106_n452.n40 gnd 0.816793f
C690 a_n3106_n452.n41 gnd 0.411619f
C691 a_n3106_n452.t31 gnd 0.10001f
C692 a_n3106_n452.t8 gnd 0.10001f
C693 a_n3106_n452.n42 gnd 0.816793f
C694 a_n3106_n452.n43 gnd 0.411619f
C695 a_n3106_n452.t9 gnd 0.10001f
C696 a_n3106_n452.t19 gnd 0.10001f
C697 a_n3106_n452.n44 gnd 0.816793f
C698 a_n3106_n452.n45 gnd 0.411619f
C699 a_n3106_n452.t5 gnd 1.03941f
C700 a_n3106_n452.n46 gnd 0.39295f
C701 a_n3106_n452.t46 gnd 1.03941f
C702 a_n3106_n452.n47 gnd 0.39295f
C703 a_n3106_n452.t35 gnd 0.10001f
C704 a_n3106_n452.t51 gnd 0.10001f
C705 a_n3106_n452.n48 gnd 0.816793f
C706 a_n3106_n452.n49 gnd 0.411619f
C707 a_n3106_n452.t42 gnd 0.10001f
C708 a_n3106_n452.t33 gnd 0.10001f
C709 a_n3106_n452.n50 gnd 0.816793f
C710 a_n3106_n452.n51 gnd 0.411619f
C711 a_n3106_n452.t53 gnd 0.10001f
C712 a_n3106_n452.t41 gnd 0.10001f
C713 a_n3106_n452.n52 gnd 0.816793f
C714 a_n3106_n452.n53 gnd 0.411619f
C715 a_n3106_n452.t48 gnd 0.10001f
C716 a_n3106_n452.t52 gnd 0.10001f
C717 a_n3106_n452.n54 gnd 0.816793f
C718 a_n3106_n452.n55 gnd 0.411619f
C719 a_n3106_n452.n56 gnd 0.411623f
C720 a_n3106_n452.n57 gnd 0.81679f
C721 a_n3106_n452.t54 gnd 0.10001f
C722 plus.n0 gnd 0.023113f
C723 plus.t20 gnd 0.420313f
C724 plus.t23 gnd 0.388639f
C725 plus.n1 gnd 0.157183f
C726 plus.n2 gnd 0.023113f
C727 plus.t6 gnd 0.388639f
C728 plus.n3 gnd 0.01975f
C729 plus.n4 gnd 0.023113f
C730 plus.t12 gnd 0.388639f
C731 plus.t8 gnd 0.388639f
C732 plus.n5 gnd 0.157183f
C733 plus.n6 gnd 0.023113f
C734 plus.t7 gnd 0.388639f
C735 plus.n7 gnd 0.157183f
C736 plus.n8 gnd 0.023113f
C737 plus.t19 gnd 0.388639f
C738 plus.n9 gnd 0.018786f
C739 plus.n10 gnd 0.023113f
C740 plus.t18 gnd 0.388639f
C741 plus.t27 gnd 0.388639f
C742 plus.n11 gnd 0.157183f
C743 plus.n12 gnd 0.023113f
C744 plus.t25 gnd 0.388639f
C745 plus.n13 gnd 0.157183f
C746 plus.n14 gnd 0.098089f
C747 plus.t9 gnd 0.388639f
C748 plus.t14 gnd 0.434763f
C749 plus.n15 gnd 0.183763f
C750 plus.n16 gnd 0.180004f
C751 plus.n17 gnd 0.029616f
C752 plus.n18 gnd 0.026155f
C753 plus.n19 gnd 0.023113f
C754 plus.n20 gnd 0.023113f
C755 plus.n21 gnd 0.02762f
C756 plus.n22 gnd 0.01975f
C757 plus.n23 gnd 0.030102f
C758 plus.n24 gnd 0.023113f
C759 plus.n25 gnd 0.023113f
C760 plus.n26 gnd 0.02875f
C761 plus.n27 gnd 0.02702f
C762 plus.n28 gnd 0.157183f
C763 plus.n29 gnd 0.028953f
C764 plus.n30 gnd 0.023113f
C765 plus.n31 gnd 0.023113f
C766 plus.n32 gnd 0.023113f
C767 plus.n33 gnd 0.029734f
C768 plus.n34 gnd 0.157183f
C769 plus.n35 gnd 0.027885f
C770 plus.n36 gnd 0.027885f
C771 plus.n37 gnd 0.023113f
C772 plus.n38 gnd 0.023113f
C773 plus.n39 gnd 0.029734f
C774 plus.n40 gnd 0.018786f
C775 plus.n41 gnd 0.028953f
C776 plus.n42 gnd 0.023113f
C777 plus.n43 gnd 0.023113f
C778 plus.n44 gnd 0.02702f
C779 plus.n45 gnd 0.02875f
C780 plus.n46 gnd 0.157183f
C781 plus.n47 gnd 0.030102f
C782 plus.n48 gnd 0.023113f
C783 plus.n49 gnd 0.023113f
C784 plus.n50 gnd 0.023113f
C785 plus.n51 gnd 0.02762f
C786 plus.n52 gnd 0.157183f
C787 plus.n53 gnd 0.026155f
C788 plus.n54 gnd 0.029616f
C789 plus.n55 gnd 0.023113f
C790 plus.n56 gnd 0.023113f
C791 plus.n57 gnd 0.030152f
C792 plus.n58 gnd 0.0084f
C793 plus.n59 gnd 0.181991f
C794 plus.n60 gnd 0.264812f
C795 plus.n61 gnd 0.023113f
C796 plus.t28 gnd 0.388639f
C797 plus.n62 gnd 0.157183f
C798 plus.n63 gnd 0.023113f
C799 plus.t26 gnd 0.388639f
C800 plus.n64 gnd 0.01975f
C801 plus.n65 gnd 0.023113f
C802 plus.t10 gnd 0.388639f
C803 plus.t15 gnd 0.388639f
C804 plus.n66 gnd 0.157183f
C805 plus.n67 gnd 0.023113f
C806 plus.t13 gnd 0.388639f
C807 plus.n68 gnd 0.157183f
C808 plus.n69 gnd 0.023113f
C809 plus.t17 gnd 0.388639f
C810 plus.n70 gnd 0.018786f
C811 plus.n71 gnd 0.023113f
C812 plus.t16 gnd 0.388639f
C813 plus.t21 gnd 0.388639f
C814 plus.n72 gnd 0.157183f
C815 plus.n73 gnd 0.023113f
C816 plus.t22 gnd 0.388639f
C817 plus.n74 gnd 0.157183f
C818 plus.n75 gnd 0.098089f
C819 plus.t5 gnd 0.388639f
C820 plus.t11 gnd 0.434763f
C821 plus.n76 gnd 0.183763f
C822 plus.n77 gnd 0.180004f
C823 plus.n78 gnd 0.029616f
C824 plus.n79 gnd 0.026155f
C825 plus.n80 gnd 0.023113f
C826 plus.n81 gnd 0.023113f
C827 plus.n82 gnd 0.02762f
C828 plus.n83 gnd 0.01975f
C829 plus.n84 gnd 0.030102f
C830 plus.n85 gnd 0.023113f
C831 plus.n86 gnd 0.023113f
C832 plus.n87 gnd 0.02875f
C833 plus.n88 gnd 0.02702f
C834 plus.n89 gnd 0.157183f
C835 plus.n90 gnd 0.028953f
C836 plus.n91 gnd 0.023113f
C837 plus.n92 gnd 0.023113f
C838 plus.n93 gnd 0.023113f
C839 plus.n94 gnd 0.029734f
C840 plus.n95 gnd 0.157183f
C841 plus.n96 gnd 0.027885f
C842 plus.n97 gnd 0.027885f
C843 plus.n98 gnd 0.023113f
C844 plus.n99 gnd 0.023113f
C845 plus.n100 gnd 0.029734f
C846 plus.n101 gnd 0.018786f
C847 plus.n102 gnd 0.028953f
C848 plus.n103 gnd 0.023113f
C849 plus.n104 gnd 0.023113f
C850 plus.n105 gnd 0.02702f
C851 plus.n106 gnd 0.02875f
C852 plus.n107 gnd 0.157183f
C853 plus.n108 gnd 0.030102f
C854 plus.n109 gnd 0.023113f
C855 plus.n110 gnd 0.023113f
C856 plus.n111 gnd 0.023113f
C857 plus.n112 gnd 0.02762f
C858 plus.n113 gnd 0.157183f
C859 plus.n114 gnd 0.026155f
C860 plus.n115 gnd 0.029616f
C861 plus.n116 gnd 0.023113f
C862 plus.n117 gnd 0.023113f
C863 plus.n118 gnd 0.030152f
C864 plus.n119 gnd 0.0084f
C865 plus.t24 gnd 0.420313f
C866 plus.n120 gnd 0.181991f
C867 plus.n121 gnd 0.833903f
C868 plus.n122 gnd 1.22934f
C869 plus.t1 gnd 0.0399f
C870 plus.t2 gnd 0.007125f
C871 plus.t4 gnd 0.007125f
C872 plus.n123 gnd 0.023108f
C873 plus.n124 gnd 0.179387f
C874 plus.t3 gnd 0.007125f
C875 plus.t0 gnd 0.007125f
C876 plus.n125 gnd 0.023108f
C877 plus.n126 gnd 0.134652f
C878 plus.n127 gnd 2.87855f
C879 a_n9628_8799.n0 gnd 4.33507f
C880 a_n9628_8799.n1 gnd 2.12179f
C881 a_n9628_8799.n2 gnd 3.56287f
C882 a_n9628_8799.n3 gnd 0.888441f
C883 a_n9628_8799.n4 gnd 0.210176f
C884 a_n9628_8799.n5 gnd 0.288599f
C885 a_n9628_8799.n6 gnd 0.210176f
C886 a_n9628_8799.n7 gnd 0.210176f
C887 a_n9628_8799.n8 gnd 0.210176f
C888 a_n9628_8799.n9 gnd 0.210176f
C889 a_n9628_8799.n10 gnd 0.210176f
C890 a_n9628_8799.n11 gnd 0.218545f
C891 a_n9628_8799.n12 gnd 0.210176f
C892 a_n9628_8799.n13 gnd 0.288599f
C893 a_n9628_8799.n14 gnd 0.210176f
C894 a_n9628_8799.n15 gnd 0.210176f
C895 a_n9628_8799.n16 gnd 0.210176f
C896 a_n9628_8799.n17 gnd 0.210176f
C897 a_n9628_8799.n18 gnd 0.210176f
C898 a_n9628_8799.n19 gnd 0.218545f
C899 a_n9628_8799.n20 gnd 0.210176f
C900 a_n9628_8799.n21 gnd 0.455543f
C901 a_n9628_8799.n22 gnd 0.210176f
C902 a_n9628_8799.n23 gnd 0.210176f
C903 a_n9628_8799.n24 gnd 0.210176f
C904 a_n9628_8799.n25 gnd 0.210176f
C905 a_n9628_8799.n26 gnd 0.210176f
C906 a_n9628_8799.n27 gnd 0.218545f
C907 a_n9628_8799.n28 gnd 0.210176f
C908 a_n9628_8799.n29 gnd 0.323633f
C909 a_n9628_8799.n30 gnd 0.210176f
C910 a_n9628_8799.n31 gnd 0.210176f
C911 a_n9628_8799.n32 gnd 0.210176f
C912 a_n9628_8799.n33 gnd 0.210176f
C913 a_n9628_8799.n34 gnd 0.210176f
C914 a_n9628_8799.n35 gnd 0.183511f
C915 a_n9628_8799.n36 gnd 0.210176f
C916 a_n9628_8799.n37 gnd 0.323633f
C917 a_n9628_8799.n38 gnd 0.210176f
C918 a_n9628_8799.n39 gnd 0.210176f
C919 a_n9628_8799.n40 gnd 0.210176f
C920 a_n9628_8799.n41 gnd 0.210176f
C921 a_n9628_8799.n42 gnd 0.210176f
C922 a_n9628_8799.n43 gnd 0.183511f
C923 a_n9628_8799.n44 gnd 0.210176f
C924 a_n9628_8799.n45 gnd 0.323633f
C925 a_n9628_8799.n46 gnd 0.210176f
C926 a_n9628_8799.n47 gnd 0.210176f
C927 a_n9628_8799.n48 gnd 0.210176f
C928 a_n9628_8799.n49 gnd 0.210176f
C929 a_n9628_8799.n50 gnd 0.210176f
C930 a_n9628_8799.n51 gnd 0.350455f
C931 a_n9628_8799.n52 gnd 1.03182f
C932 a_n9628_8799.n53 gnd 1.0172f
C933 a_n9628_8799.n54 gnd 2.9877f
C934 a_n9628_8799.n55 gnd 1.54042f
C935 a_n9628_8799.n56 gnd 3.79021f
C936 a_n9628_8799.n57 gnd 1.0172f
C937 a_n9628_8799.n58 gnd 0.253032f
C938 a_n9628_8799.n59 gnd 0.003699f
C939 a_n9628_8799.n60 gnd 0.009751f
C940 a_n9628_8799.n61 gnd 0.010654f
C941 a_n9628_8799.n62 gnd 0.00563f
C942 a_n9628_8799.n64 gnd 0.004724f
C943 a_n9628_8799.n65 gnd 0.010217f
C944 a_n9628_8799.n66 gnd 0.010217f
C945 a_n9628_8799.n67 gnd 0.004724f
C946 a_n9628_8799.n69 gnd 0.00563f
C947 a_n9628_8799.n70 gnd 0.010654f
C948 a_n9628_8799.n71 gnd 0.009751f
C949 a_n9628_8799.n72 gnd 0.003699f
C950 a_n9628_8799.n73 gnd 0.253032f
C951 a_n9628_8799.n74 gnd 0.003699f
C952 a_n9628_8799.n75 gnd 0.009751f
C953 a_n9628_8799.n76 gnd 0.010654f
C954 a_n9628_8799.n77 gnd 0.00563f
C955 a_n9628_8799.n79 gnd 0.004724f
C956 a_n9628_8799.n80 gnd 0.010217f
C957 a_n9628_8799.n81 gnd 0.010217f
C958 a_n9628_8799.n82 gnd 0.004724f
C959 a_n9628_8799.n84 gnd 0.00563f
C960 a_n9628_8799.n85 gnd 0.010654f
C961 a_n9628_8799.n86 gnd 0.009751f
C962 a_n9628_8799.n87 gnd 0.003699f
C963 a_n9628_8799.n88 gnd 0.253032f
C964 a_n9628_8799.n89 gnd 0.003699f
C965 a_n9628_8799.n90 gnd 0.009751f
C966 a_n9628_8799.n91 gnd 0.010654f
C967 a_n9628_8799.n92 gnd 0.00563f
C968 a_n9628_8799.n94 gnd 0.004724f
C969 a_n9628_8799.n95 gnd 0.010217f
C970 a_n9628_8799.n96 gnd 0.010217f
C971 a_n9628_8799.n97 gnd 0.004724f
C972 a_n9628_8799.n99 gnd 0.00563f
C973 a_n9628_8799.n100 gnd 0.010654f
C974 a_n9628_8799.n101 gnd 0.009751f
C975 a_n9628_8799.n102 gnd 0.003699f
C976 a_n9628_8799.n103 gnd 0.003699f
C977 a_n9628_8799.n104 gnd 0.009751f
C978 a_n9628_8799.n105 gnd 0.010654f
C979 a_n9628_8799.n106 gnd 0.00563f
C980 a_n9628_8799.n108 gnd 0.004724f
C981 a_n9628_8799.n109 gnd 0.010217f
C982 a_n9628_8799.n110 gnd 0.010217f
C983 a_n9628_8799.n111 gnd 0.004724f
C984 a_n9628_8799.n113 gnd 0.00563f
C985 a_n9628_8799.n114 gnd 0.010654f
C986 a_n9628_8799.n115 gnd 0.009751f
C987 a_n9628_8799.n116 gnd 0.003699f
C988 a_n9628_8799.n117 gnd 0.253032f
C989 a_n9628_8799.n118 gnd 0.003699f
C990 a_n9628_8799.n119 gnd 0.009751f
C991 a_n9628_8799.n120 gnd 0.010654f
C992 a_n9628_8799.n121 gnd 0.00563f
C993 a_n9628_8799.n123 gnd 0.004724f
C994 a_n9628_8799.n124 gnd 0.010217f
C995 a_n9628_8799.n125 gnd 0.010217f
C996 a_n9628_8799.n126 gnd 0.004724f
C997 a_n9628_8799.n128 gnd 0.00563f
C998 a_n9628_8799.n129 gnd 0.010654f
C999 a_n9628_8799.n130 gnd 0.009751f
C1000 a_n9628_8799.n131 gnd 0.003699f
C1001 a_n9628_8799.n132 gnd 0.253032f
C1002 a_n9628_8799.n133 gnd 0.003699f
C1003 a_n9628_8799.n134 gnd 0.009751f
C1004 a_n9628_8799.n135 gnd 0.010654f
C1005 a_n9628_8799.n136 gnd 0.00563f
C1006 a_n9628_8799.n138 gnd 0.004724f
C1007 a_n9628_8799.n139 gnd 0.010217f
C1008 a_n9628_8799.n140 gnd 0.010217f
C1009 a_n9628_8799.n141 gnd 0.004724f
C1010 a_n9628_8799.n143 gnd 0.00563f
C1011 a_n9628_8799.n144 gnd 0.010654f
C1012 a_n9628_8799.n145 gnd 0.009751f
C1013 a_n9628_8799.n146 gnd 0.003699f
C1014 a_n9628_8799.n147 gnd 0.253032f
C1015 a_n9628_8799.t37 gnd 0.14578f
C1016 a_n9628_8799.t34 gnd 0.14578f
C1017 a_n9628_8799.t22 gnd 0.14578f
C1018 a_n9628_8799.n148 gnd 1.14979f
C1019 a_n9628_8799.t24 gnd 0.14578f
C1020 a_n9628_8799.t40 gnd 0.14578f
C1021 a_n9628_8799.n149 gnd 1.14789f
C1022 a_n9628_8799.t26 gnd 0.14578f
C1023 a_n9628_8799.t30 gnd 0.14578f
C1024 a_n9628_8799.n150 gnd 1.14789f
C1025 a_n9628_8799.t29 gnd 0.14578f
C1026 a_n9628_8799.t42 gnd 0.14578f
C1027 a_n9628_8799.n151 gnd 1.14789f
C1028 a_n9628_8799.t25 gnd 0.14578f
C1029 a_n9628_8799.t35 gnd 0.14578f
C1030 a_n9628_8799.n152 gnd 1.14789f
C1031 a_n9628_8799.t39 gnd 0.14578f
C1032 a_n9628_8799.t21 gnd 0.14578f
C1033 a_n9628_8799.n153 gnd 1.14789f
C1034 a_n9628_8799.t19 gnd 0.113385f
C1035 a_n9628_8799.t5 gnd 0.113385f
C1036 a_n9628_8799.n154 gnd 1.00486f
C1037 a_n9628_8799.t3 gnd 0.113385f
C1038 a_n9628_8799.t18 gnd 0.113385f
C1039 a_n9628_8799.n155 gnd 1.00191f
C1040 a_n9628_8799.t16 gnd 0.113385f
C1041 a_n9628_8799.t7 gnd 0.113385f
C1042 a_n9628_8799.n156 gnd 1.00191f
C1043 a_n9628_8799.t12 gnd 0.113385f
C1044 a_n9628_8799.t2 gnd 0.113385f
C1045 a_n9628_8799.n157 gnd 1.00486f
C1046 a_n9628_8799.t0 gnd 0.113385f
C1047 a_n9628_8799.t17 gnd 0.113385f
C1048 a_n9628_8799.n158 gnd 1.00191f
C1049 a_n9628_8799.t8 gnd 0.113385f
C1050 a_n9628_8799.t15 gnd 0.113385f
C1051 a_n9628_8799.n159 gnd 1.00191f
C1052 a_n9628_8799.t4 gnd 0.113385f
C1053 a_n9628_8799.t10 gnd 0.113385f
C1054 a_n9628_8799.n160 gnd 1.00486f
C1055 a_n9628_8799.t47 gnd 0.113385f
C1056 a_n9628_8799.t46 gnd 0.113385f
C1057 a_n9628_8799.n161 gnd 1.00191f
C1058 a_n9628_8799.t6 gnd 0.113385f
C1059 a_n9628_8799.t44 gnd 0.113385f
C1060 a_n9628_8799.n162 gnd 1.00191f
C1061 a_n9628_8799.t9 gnd 0.113385f
C1062 a_n9628_8799.t11 gnd 0.113385f
C1063 a_n9628_8799.n163 gnd 1.00191f
C1064 a_n9628_8799.t13 gnd 0.113385f
C1065 a_n9628_8799.t45 gnd 0.113385f
C1066 a_n9628_8799.n164 gnd 1.00191f
C1067 a_n9628_8799.t14 gnd 0.113385f
C1068 a_n9628_8799.t1 gnd 0.113385f
C1069 a_n9628_8799.n165 gnd 1.00191f
C1070 a_n9628_8799.t94 gnd 0.604473f
C1071 a_n9628_8799.n166 gnd 0.272141f
C1072 a_n9628_8799.t130 gnd 0.604473f
C1073 a_n9628_8799.t151 gnd 0.604473f
C1074 a_n9628_8799.n167 gnd 0.274091f
C1075 a_n9628_8799.t152 gnd 0.604473f
C1076 a_n9628_8799.t80 gnd 0.604473f
C1077 a_n9628_8799.n168 gnd 0.267216f
C1078 a_n9628_8799.t120 gnd 0.604473f
C1079 a_n9628_8799.t127 gnd 0.604473f
C1080 a_n9628_8799.n169 gnd 0.271239f
C1081 a_n9628_8799.t56 gnd 0.604473f
C1082 a_n9628_8799.t99 gnd 0.604473f
C1083 a_n9628_8799.t97 gnd 0.615913f
C1084 a_n9628_8799.n170 gnd 0.253399f
C1085 a_n9628_8799.n171 gnd 0.274468f
C1086 a_n9628_8799.t131 gnd 0.604473f
C1087 a_n9628_8799.n172 gnd 0.272141f
C1088 a_n9628_8799.n173 gnd 0.267863f
C1089 a_n9628_8799.t95 gnd 0.604473f
C1090 a_n9628_8799.n174 gnd 0.266568f
C1091 a_n9628_8799.t50 gnd 0.604473f
C1092 a_n9628_8799.n175 gnd 0.273833f
C1093 a_n9628_8799.t82 gnd 0.604473f
C1094 a_n9628_8799.n176 gnd 0.274091f
C1095 a_n9628_8799.n177 gnd 0.271676f
C1096 a_n9628_8799.t155 gnd 0.604473f
C1097 a_n9628_8799.n178 gnd 0.267216f
C1098 a_n9628_8799.t116 gnd 0.604473f
C1099 a_n9628_8799.n179 gnd 0.271676f
C1100 a_n9628_8799.n180 gnd 0.273833f
C1101 a_n9628_8799.t98 gnd 0.604473f
C1102 a_n9628_8799.n181 gnd 0.271239f
C1103 a_n9628_8799.n182 gnd 0.266568f
C1104 a_n9628_8799.t150 gnd 0.604473f
C1105 a_n9628_8799.n183 gnd 0.267863f
C1106 a_n9628_8799.t96 gnd 0.604473f
C1107 a_n9628_8799.n184 gnd 0.274468f
C1108 a_n9628_8799.t128 gnd 0.615903f
C1109 a_n9628_8799.t105 gnd 0.604473f
C1110 a_n9628_8799.n185 gnd 0.272141f
C1111 a_n9628_8799.t144 gnd 0.604473f
C1112 a_n9628_8799.t163 gnd 0.604473f
C1113 a_n9628_8799.n186 gnd 0.274091f
C1114 a_n9628_8799.t165 gnd 0.604473f
C1115 a_n9628_8799.t89 gnd 0.604473f
C1116 a_n9628_8799.n187 gnd 0.267216f
C1117 a_n9628_8799.t133 gnd 0.604473f
C1118 a_n9628_8799.t140 gnd 0.604473f
C1119 a_n9628_8799.n188 gnd 0.271239f
C1120 a_n9628_8799.t68 gnd 0.604473f
C1121 a_n9628_8799.t112 gnd 0.604473f
C1122 a_n9628_8799.t110 gnd 0.615913f
C1123 a_n9628_8799.n189 gnd 0.253399f
C1124 a_n9628_8799.n190 gnd 0.274468f
C1125 a_n9628_8799.t148 gnd 0.604473f
C1126 a_n9628_8799.n191 gnd 0.272141f
C1127 a_n9628_8799.n192 gnd 0.267863f
C1128 a_n9628_8799.t106 gnd 0.604473f
C1129 a_n9628_8799.n193 gnd 0.266568f
C1130 a_n9628_8799.t64 gnd 0.604473f
C1131 a_n9628_8799.n194 gnd 0.273833f
C1132 a_n9628_8799.t92 gnd 0.604473f
C1133 a_n9628_8799.n195 gnd 0.274091f
C1134 a_n9628_8799.n196 gnd 0.271676f
C1135 a_n9628_8799.t167 gnd 0.604473f
C1136 a_n9628_8799.n197 gnd 0.267216f
C1137 a_n9628_8799.t129 gnd 0.604473f
C1138 a_n9628_8799.n198 gnd 0.271676f
C1139 a_n9628_8799.n199 gnd 0.273833f
C1140 a_n9628_8799.t111 gnd 0.604473f
C1141 a_n9628_8799.n200 gnd 0.271239f
C1142 a_n9628_8799.n201 gnd 0.266568f
C1143 a_n9628_8799.t162 gnd 0.604473f
C1144 a_n9628_8799.n202 gnd 0.267863f
C1145 a_n9628_8799.t107 gnd 0.604473f
C1146 a_n9628_8799.n203 gnd 0.274468f
C1147 a_n9628_8799.t141 gnd 0.615903f
C1148 a_n9628_8799.n204 gnd 0.908741f
C1149 a_n9628_8799.t71 gnd 0.604473f
C1150 a_n9628_8799.n205 gnd 0.272141f
C1151 a_n9628_8799.t90 gnd 0.604473f
C1152 a_n9628_8799.t124 gnd 0.604473f
C1153 a_n9628_8799.n206 gnd 0.274091f
C1154 a_n9628_8799.t104 gnd 0.604473f
C1155 a_n9628_8799.t108 gnd 0.604473f
C1156 a_n9628_8799.n207 gnd 0.267216f
C1157 a_n9628_8799.t135 gnd 0.604473f
C1158 a_n9628_8799.t51 gnd 0.604473f
C1159 a_n9628_8799.n208 gnd 0.271239f
C1160 a_n9628_8799.t77 gnd 0.604473f
C1161 a_n9628_8799.t60 gnd 0.604473f
C1162 a_n9628_8799.t81 gnd 0.615913f
C1163 a_n9628_8799.n209 gnd 0.253399f
C1164 a_n9628_8799.n210 gnd 0.274468f
C1165 a_n9628_8799.t122 gnd 0.604473f
C1166 a_n9628_8799.n211 gnd 0.272141f
C1167 a_n9628_8799.n212 gnd 0.267863f
C1168 a_n9628_8799.t100 gnd 0.604473f
C1169 a_n9628_8799.n213 gnd 0.266568f
C1170 a_n9628_8799.t117 gnd 0.604473f
C1171 a_n9628_8799.n214 gnd 0.273833f
C1172 a_n9628_8799.t69 gnd 0.604473f
C1173 a_n9628_8799.n215 gnd 0.274091f
C1174 a_n9628_8799.n216 gnd 0.271676f
C1175 a_n9628_8799.t85 gnd 0.604473f
C1176 a_n9628_8799.n217 gnd 0.267216f
C1177 a_n9628_8799.t61 gnd 0.604473f
C1178 a_n9628_8799.n218 gnd 0.271676f
C1179 a_n9628_8799.n219 gnd 0.273833f
C1180 a_n9628_8799.t143 gnd 0.604473f
C1181 a_n9628_8799.n220 gnd 0.271239f
C1182 a_n9628_8799.n221 gnd 0.266568f
C1183 a_n9628_8799.t153 gnd 0.604473f
C1184 a_n9628_8799.n222 gnd 0.267863f
C1185 a_n9628_8799.t48 gnd 0.604473f
C1186 a_n9628_8799.n223 gnd 0.274468f
C1187 a_n9628_8799.t113 gnd 0.615903f
C1188 a_n9628_8799.n224 gnd 1.97579f
C1189 a_n9628_8799.t55 gnd 0.615903f
C1190 a_n9628_8799.t53 gnd 0.604473f
C1191 a_n9628_8799.t139 gnd 0.604473f
C1192 a_n9628_8799.n225 gnd 0.272141f
C1193 a_n9628_8799.t75 gnd 0.604473f
C1194 a_n9628_8799.t58 gnd 0.604473f
C1195 a_n9628_8799.t146 gnd 0.604473f
C1196 a_n9628_8799.n226 gnd 0.271239f
C1197 a_n9628_8799.t101 gnd 0.604473f
C1198 a_n9628_8799.t76 gnd 0.604473f
C1199 a_n9628_8799.t164 gnd 0.604473f
C1200 a_n9628_8799.n227 gnd 0.271676f
C1201 a_n9628_8799.t119 gnd 0.604473f
C1202 a_n9628_8799.t79 gnd 0.604473f
C1203 a_n9628_8799.t158 gnd 0.604473f
C1204 a_n9628_8799.n228 gnd 0.271676f
C1205 a_n9628_8799.t121 gnd 0.604473f
C1206 a_n9628_8799.t93 gnd 0.604473f
C1207 a_n9628_8799.t54 gnd 0.604473f
C1208 a_n9628_8799.n229 gnd 0.271239f
C1209 a_n9628_8799.t142 gnd 0.604473f
C1210 a_n9628_8799.t123 gnd 0.604473f
C1211 a_n9628_8799.t59 gnd 0.604473f
C1212 a_n9628_8799.n230 gnd 0.272141f
C1213 a_n9628_8799.t145 gnd 0.615913f
C1214 a_n9628_8799.n231 gnd 0.253399f
C1215 a_n9628_8799.t149 gnd 0.604473f
C1216 a_n9628_8799.n232 gnd 0.274468f
C1217 a_n9628_8799.n233 gnd 0.267863f
C1218 a_n9628_8799.n234 gnd 0.266568f
C1219 a_n9628_8799.n235 gnd 0.273833f
C1220 a_n9628_8799.n236 gnd 0.274091f
C1221 a_n9628_8799.n237 gnd 0.267216f
C1222 a_n9628_8799.n238 gnd 0.267216f
C1223 a_n9628_8799.n239 gnd 0.274091f
C1224 a_n9628_8799.n240 gnd 0.273833f
C1225 a_n9628_8799.n241 gnd 0.266568f
C1226 a_n9628_8799.n242 gnd 0.267863f
C1227 a_n9628_8799.n243 gnd 0.274468f
C1228 a_n9628_8799.t66 gnd 0.615903f
C1229 a_n9628_8799.t65 gnd 0.604473f
C1230 a_n9628_8799.t156 gnd 0.604473f
C1231 a_n9628_8799.n244 gnd 0.272141f
C1232 a_n9628_8799.t84 gnd 0.604473f
C1233 a_n9628_8799.t73 gnd 0.604473f
C1234 a_n9628_8799.t159 gnd 0.604473f
C1235 a_n9628_8799.n245 gnd 0.271239f
C1236 a_n9628_8799.t115 gnd 0.604473f
C1237 a_n9628_8799.t87 gnd 0.604473f
C1238 a_n9628_8799.t57 gnd 0.604473f
C1239 a_n9628_8799.n246 gnd 0.271676f
C1240 a_n9628_8799.t132 gnd 0.604473f
C1241 a_n9628_8799.t88 gnd 0.604473f
C1242 a_n9628_8799.t49 gnd 0.604473f
C1243 a_n9628_8799.n247 gnd 0.271676f
C1244 a_n9628_8799.t137 gnd 0.604473f
C1245 a_n9628_8799.t103 gnd 0.604473f
C1246 a_n9628_8799.t67 gnd 0.604473f
C1247 a_n9628_8799.n248 gnd 0.271239f
C1248 a_n9628_8799.t157 gnd 0.604473f
C1249 a_n9628_8799.t138 gnd 0.604473f
C1250 a_n9628_8799.t74 gnd 0.604473f
C1251 a_n9628_8799.n249 gnd 0.272141f
C1252 a_n9628_8799.t160 gnd 0.615913f
C1253 a_n9628_8799.n250 gnd 0.253399f
C1254 a_n9628_8799.t161 gnd 0.604473f
C1255 a_n9628_8799.n251 gnd 0.274468f
C1256 a_n9628_8799.n252 gnd 0.267863f
C1257 a_n9628_8799.n253 gnd 0.266568f
C1258 a_n9628_8799.n254 gnd 0.273833f
C1259 a_n9628_8799.n255 gnd 0.274091f
C1260 a_n9628_8799.n256 gnd 0.267216f
C1261 a_n9628_8799.n257 gnd 0.267216f
C1262 a_n9628_8799.n258 gnd 0.274091f
C1263 a_n9628_8799.n259 gnd 0.273833f
C1264 a_n9628_8799.n260 gnd 0.266568f
C1265 a_n9628_8799.n261 gnd 0.267863f
C1266 a_n9628_8799.n262 gnd 0.274468f
C1267 a_n9628_8799.n263 gnd 0.908741f
C1268 a_n9628_8799.t114 gnd 0.615903f
C1269 a_n9628_8799.t136 gnd 0.604473f
C1270 a_n9628_8799.t72 gnd 0.604473f
C1271 a_n9628_8799.n264 gnd 0.272141f
C1272 a_n9628_8799.t154 gnd 0.604473f
C1273 a_n9628_8799.t91 gnd 0.604473f
C1274 a_n9628_8799.t147 gnd 0.604473f
C1275 a_n9628_8799.n265 gnd 0.271239f
C1276 a_n9628_8799.t78 gnd 0.604473f
C1277 a_n9628_8799.t126 gnd 0.604473f
C1278 a_n9628_8799.t63 gnd 0.604473f
C1279 a_n9628_8799.n266 gnd 0.271676f
C1280 a_n9628_8799.t109 gnd 0.604473f
C1281 a_n9628_8799.t86 gnd 0.604473f
C1282 a_n9628_8799.t134 gnd 0.604473f
C1283 a_n9628_8799.n267 gnd 0.271676f
C1284 a_n9628_8799.t70 gnd 0.604473f
C1285 a_n9628_8799.t118 gnd 0.604473f
C1286 a_n9628_8799.t52 gnd 0.604473f
C1287 a_n9628_8799.n268 gnd 0.271239f
C1288 a_n9628_8799.t102 gnd 0.604473f
C1289 a_n9628_8799.t166 gnd 0.604473f
C1290 a_n9628_8799.t125 gnd 0.604473f
C1291 a_n9628_8799.n269 gnd 0.272141f
C1292 a_n9628_8799.t83 gnd 0.615913f
C1293 a_n9628_8799.n270 gnd 0.253399f
C1294 a_n9628_8799.t62 gnd 0.604473f
C1295 a_n9628_8799.n271 gnd 0.274468f
C1296 a_n9628_8799.n272 gnd 0.267863f
C1297 a_n9628_8799.n273 gnd 0.266568f
C1298 a_n9628_8799.n274 gnd 0.273833f
C1299 a_n9628_8799.n275 gnd 0.274091f
C1300 a_n9628_8799.n276 gnd 0.267216f
C1301 a_n9628_8799.n277 gnd 0.267216f
C1302 a_n9628_8799.n278 gnd 0.274091f
C1303 a_n9628_8799.n279 gnd 0.273833f
C1304 a_n9628_8799.n280 gnd 0.266568f
C1305 a_n9628_8799.n281 gnd 0.267863f
C1306 a_n9628_8799.n282 gnd 0.274468f
C1307 a_n9628_8799.n283 gnd 1.35394f
C1308 a_n9628_8799.n284 gnd 17.5375f
C1309 a_n9628_8799.n285 gnd 4.42387f
C1310 a_n9628_8799.n286 gnd 7.70781f
C1311 a_n9628_8799.t28 gnd 0.14578f
C1312 a_n9628_8799.t38 gnd 0.14578f
C1313 a_n9628_8799.n287 gnd 1.14789f
C1314 a_n9628_8799.t27 gnd 0.14578f
C1315 a_n9628_8799.t41 gnd 0.14578f
C1316 a_n9628_8799.n288 gnd 1.14979f
C1317 a_n9628_8799.t43 gnd 0.14578f
C1318 a_n9628_8799.t23 gnd 0.14578f
C1319 a_n9628_8799.n289 gnd 1.14789f
C1320 a_n9628_8799.t33 gnd 0.14578f
C1321 a_n9628_8799.t32 gnd 0.14578f
C1322 a_n9628_8799.n290 gnd 1.14789f
C1323 a_n9628_8799.t31 gnd 0.14578f
C1324 a_n9628_8799.t36 gnd 0.14578f
C1325 a_n9628_8799.n291 gnd 1.14789f
C1326 a_n9628_8799.n292 gnd 1.1479f
C1327 a_n9628_8799.t20 gnd 0.14578f
C1328 CSoutput.n0 gnd 0.04891f
C1329 CSoutput.t202 gnd 0.323528f
C1330 CSoutput.n1 gnd 0.146089f
C1331 CSoutput.n2 gnd 0.04891f
C1332 CSoutput.t200 gnd 0.323528f
C1333 CSoutput.n3 gnd 0.038765f
C1334 CSoutput.n4 gnd 0.04891f
C1335 CSoutput.t212 gnd 0.323528f
C1336 CSoutput.n5 gnd 0.033427f
C1337 CSoutput.n6 gnd 0.04891f
C1338 CSoutput.t197 gnd 0.323528f
C1339 CSoutput.t207 gnd 0.323528f
C1340 CSoutput.n7 gnd 0.144497f
C1341 CSoutput.n8 gnd 0.04891f
C1342 CSoutput.t210 gnd 0.323528f
C1343 CSoutput.n9 gnd 0.031871f
C1344 CSoutput.n10 gnd 0.04891f
C1345 CSoutput.t193 gnd 0.323528f
C1346 CSoutput.t199 gnd 0.323528f
C1347 CSoutput.n11 gnd 0.144497f
C1348 CSoutput.n12 gnd 0.04891f
C1349 CSoutput.t204 gnd 0.323528f
C1350 CSoutput.n13 gnd 0.033427f
C1351 CSoutput.n14 gnd 0.04891f
C1352 CSoutput.t213 gnd 0.323528f
C1353 CSoutput.t196 gnd 0.323528f
C1354 CSoutput.n15 gnd 0.144497f
C1355 CSoutput.n16 gnd 0.04891f
C1356 CSoutput.t203 gnd 0.323528f
C1357 CSoutput.n17 gnd 0.035702f
C1358 CSoutput.t192 gnd 0.386624f
C1359 CSoutput.t201 gnd 0.323528f
C1360 CSoutput.n18 gnd 0.184466f
C1361 CSoutput.n19 gnd 0.178996f
C1362 CSoutput.n20 gnd 0.207657f
C1363 CSoutput.n21 gnd 0.04891f
C1364 CSoutput.n22 gnd 0.040821f
C1365 CSoutput.n23 gnd 0.144497f
C1366 CSoutput.n24 gnd 0.03935f
C1367 CSoutput.n25 gnd 0.038765f
C1368 CSoutput.n26 gnd 0.04891f
C1369 CSoutput.n27 gnd 0.04891f
C1370 CSoutput.n28 gnd 0.040507f
C1371 CSoutput.n29 gnd 0.034391f
C1372 CSoutput.n30 gnd 0.147713f
C1373 CSoutput.n31 gnd 0.034865f
C1374 CSoutput.n32 gnd 0.04891f
C1375 CSoutput.n33 gnd 0.04891f
C1376 CSoutput.n34 gnd 0.04891f
C1377 CSoutput.n35 gnd 0.040075f
C1378 CSoutput.n36 gnd 0.144497f
C1379 CSoutput.n37 gnd 0.038326f
C1380 CSoutput.n38 gnd 0.039789f
C1381 CSoutput.n39 gnd 0.04891f
C1382 CSoutput.n40 gnd 0.04891f
C1383 CSoutput.n41 gnd 0.040812f
C1384 CSoutput.n42 gnd 0.037303f
C1385 CSoutput.n43 gnd 0.144497f
C1386 CSoutput.n44 gnd 0.038248f
C1387 CSoutput.n45 gnd 0.04891f
C1388 CSoutput.n46 gnd 0.04891f
C1389 CSoutput.n47 gnd 0.04891f
C1390 CSoutput.n48 gnd 0.038248f
C1391 CSoutput.n49 gnd 0.144497f
C1392 CSoutput.n50 gnd 0.037303f
C1393 CSoutput.n51 gnd 0.040812f
C1394 CSoutput.n52 gnd 0.04891f
C1395 CSoutput.n53 gnd 0.04891f
C1396 CSoutput.n54 gnd 0.039789f
C1397 CSoutput.n55 gnd 0.038326f
C1398 CSoutput.n56 gnd 0.144497f
C1399 CSoutput.n57 gnd 0.040075f
C1400 CSoutput.n58 gnd 0.04891f
C1401 CSoutput.n59 gnd 0.04891f
C1402 CSoutput.n60 gnd 0.04891f
C1403 CSoutput.n61 gnd 0.034865f
C1404 CSoutput.n62 gnd 0.147713f
C1405 CSoutput.n63 gnd 0.034391f
C1406 CSoutput.t208 gnd 0.323528f
C1407 CSoutput.n64 gnd 0.144497f
C1408 CSoutput.n65 gnd 0.040507f
C1409 CSoutput.n66 gnd 0.04891f
C1410 CSoutput.n67 gnd 0.04891f
C1411 CSoutput.n68 gnd 0.04891f
C1412 CSoutput.n69 gnd 0.03935f
C1413 CSoutput.n70 gnd 0.144497f
C1414 CSoutput.n71 gnd 0.040821f
C1415 CSoutput.n72 gnd 0.035702f
C1416 CSoutput.n73 gnd 0.04891f
C1417 CSoutput.n74 gnd 0.04891f
C1418 CSoutput.n75 gnd 0.037026f
C1419 CSoutput.n76 gnd 0.02199f
C1420 CSoutput.t194 gnd 0.363506f
C1421 CSoutput.n77 gnd 0.180575f
C1422 CSoutput.n78 gnd 0.738615f
C1423 CSoutput.t180 gnd 0.061008f
C1424 CSoutput.t5 gnd 0.061008f
C1425 CSoutput.n79 gnd 0.472345f
C1426 CSoutput.t169 gnd 0.061008f
C1427 CSoutput.t7 gnd 0.061008f
C1428 CSoutput.n80 gnd 0.471503f
C1429 CSoutput.n81 gnd 0.478574f
C1430 CSoutput.t27 gnd 0.061008f
C1431 CSoutput.t44 gnd 0.061008f
C1432 CSoutput.n82 gnd 0.471503f
C1433 CSoutput.n83 gnd 0.235821f
C1434 CSoutput.t76 gnd 0.061008f
C1435 CSoutput.t176 gnd 0.061008f
C1436 CSoutput.n84 gnd 0.471503f
C1437 CSoutput.n85 gnd 0.235821f
C1438 CSoutput.t50 gnd 0.061008f
C1439 CSoutput.t25 gnd 0.061008f
C1440 CSoutput.n86 gnd 0.471503f
C1441 CSoutput.n87 gnd 0.235821f
C1442 CSoutput.t17 gnd 0.061008f
C1443 CSoutput.t179 gnd 0.061008f
C1444 CSoutput.n88 gnd 0.471503f
C1445 CSoutput.n89 gnd 0.235821f
C1446 CSoutput.t59 gnd 0.061008f
C1447 CSoutput.t71 gnd 0.061008f
C1448 CSoutput.n90 gnd 0.471503f
C1449 CSoutput.n91 gnd 0.235821f
C1450 CSoutput.t28 gnd 0.061008f
C1451 CSoutput.t187 gnd 0.061008f
C1452 CSoutput.n92 gnd 0.471503f
C1453 CSoutput.n93 gnd 0.235821f
C1454 CSoutput.t84 gnd 0.061008f
C1455 CSoutput.t165 gnd 0.061008f
C1456 CSoutput.n94 gnd 0.471503f
C1457 CSoutput.n95 gnd 0.235821f
C1458 CSoutput.t65 gnd 0.061008f
C1459 CSoutput.t24 gnd 0.061008f
C1460 CSoutput.n96 gnd 0.471503f
C1461 CSoutput.n97 gnd 0.432442f
C1462 CSoutput.t185 gnd 0.061008f
C1463 CSoutput.t31 gnd 0.061008f
C1464 CSoutput.n98 gnd 0.472345f
C1465 CSoutput.t74 gnd 0.061008f
C1466 CSoutput.t177 gnd 0.061008f
C1467 CSoutput.n99 gnd 0.471503f
C1468 CSoutput.n100 gnd 0.478574f
C1469 CSoutput.t171 gnd 0.061008f
C1470 CSoutput.t38 gnd 0.061008f
C1471 CSoutput.n101 gnd 0.471503f
C1472 CSoutput.n102 gnd 0.235821f
C1473 CSoutput.t75 gnd 0.061008f
C1474 CSoutput.t81 gnd 0.061008f
C1475 CSoutput.n103 gnd 0.471503f
C1476 CSoutput.n104 gnd 0.235821f
C1477 CSoutput.t61 gnd 0.061008f
C1478 CSoutput.t189 gnd 0.061008f
C1479 CSoutput.n105 gnd 0.471503f
C1480 CSoutput.n106 gnd 0.235821f
C1481 CSoutput.t41 gnd 0.061008f
C1482 CSoutput.t73 gnd 0.061008f
C1483 CSoutput.n107 gnd 0.471503f
C1484 CSoutput.n108 gnd 0.235821f
C1485 CSoutput.t62 gnd 0.061008f
C1486 CSoutput.t20 gnd 0.061008f
C1487 CSoutput.n109 gnd 0.471503f
C1488 CSoutput.n110 gnd 0.235821f
C1489 CSoutput.t184 gnd 0.061008f
C1490 CSoutput.t30 gnd 0.061008f
C1491 CSoutput.n111 gnd 0.471503f
C1492 CSoutput.n112 gnd 0.235821f
C1493 CSoutput.t182 gnd 0.061008f
C1494 CSoutput.t70 gnd 0.061008f
C1495 CSoutput.n113 gnd 0.471503f
C1496 CSoutput.n114 gnd 0.235821f
C1497 CSoutput.t170 gnd 0.061008f
C1498 CSoutput.t4 gnd 0.061008f
C1499 CSoutput.n115 gnd 0.471503f
C1500 CSoutput.n116 gnd 0.351669f
C1501 CSoutput.n117 gnd 0.443452f
C1502 CSoutput.t36 gnd 0.061008f
C1503 CSoutput.t188 gnd 0.061008f
C1504 CSoutput.n118 gnd 0.472345f
C1505 CSoutput.t48 gnd 0.061008f
C1506 CSoutput.t12 gnd 0.061008f
C1507 CSoutput.n119 gnd 0.471503f
C1508 CSoutput.n120 gnd 0.478574f
C1509 CSoutput.t32 gnd 0.061008f
C1510 CSoutput.t56 gnd 0.061008f
C1511 CSoutput.n121 gnd 0.471503f
C1512 CSoutput.n122 gnd 0.235821f
C1513 CSoutput.t49 gnd 0.061008f
C1514 CSoutput.t168 gnd 0.061008f
C1515 CSoutput.n123 gnd 0.471503f
C1516 CSoutput.n124 gnd 0.235821f
C1517 CSoutput.t64 gnd 0.061008f
C1518 CSoutput.t58 gnd 0.061008f
C1519 CSoutput.n125 gnd 0.471503f
C1520 CSoutput.n126 gnd 0.235821f
C1521 CSoutput.t78 gnd 0.061008f
C1522 CSoutput.t3 gnd 0.061008f
C1523 CSoutput.n127 gnd 0.471503f
C1524 CSoutput.n128 gnd 0.235821f
C1525 CSoutput.t186 gnd 0.061008f
C1526 CSoutput.t88 gnd 0.061008f
C1527 CSoutput.n129 gnd 0.471503f
C1528 CSoutput.n130 gnd 0.235821f
C1529 CSoutput.t13 gnd 0.061008f
C1530 CSoutput.t175 gnd 0.061008f
C1531 CSoutput.n131 gnd 0.471503f
C1532 CSoutput.n132 gnd 0.235821f
C1533 CSoutput.t57 gnd 0.061008f
C1534 CSoutput.t166 gnd 0.061008f
C1535 CSoutput.n133 gnd 0.471503f
C1536 CSoutput.n134 gnd 0.235821f
C1537 CSoutput.t37 gnd 0.061008f
C1538 CSoutput.t33 gnd 0.061008f
C1539 CSoutput.n135 gnd 0.471503f
C1540 CSoutput.n136 gnd 0.351669f
C1541 CSoutput.n137 gnd 0.495666f
C1542 CSoutput.n138 gnd 9.49517f
C1543 CSoutput.n140 gnd 0.865206f
C1544 CSoutput.n141 gnd 0.648904f
C1545 CSoutput.n142 gnd 0.865206f
C1546 CSoutput.n143 gnd 0.865206f
C1547 CSoutput.n144 gnd 2.3294f
C1548 CSoutput.n145 gnd 0.865206f
C1549 CSoutput.n146 gnd 0.865206f
C1550 CSoutput.t209 gnd 1.08151f
C1551 CSoutput.n147 gnd 0.865206f
C1552 CSoutput.n148 gnd 0.865206f
C1553 CSoutput.n152 gnd 0.865206f
C1554 CSoutput.n156 gnd 0.865206f
C1555 CSoutput.n157 gnd 0.865206f
C1556 CSoutput.n159 gnd 0.865206f
C1557 CSoutput.n164 gnd 0.865206f
C1558 CSoutput.n166 gnd 0.865206f
C1559 CSoutput.n167 gnd 0.865206f
C1560 CSoutput.n169 gnd 0.865206f
C1561 CSoutput.n170 gnd 0.865206f
C1562 CSoutput.n172 gnd 0.865206f
C1563 CSoutput.t195 gnd 14.4575f
C1564 CSoutput.n174 gnd 0.865206f
C1565 CSoutput.n175 gnd 0.648904f
C1566 CSoutput.n176 gnd 0.865206f
C1567 CSoutput.n177 gnd 0.865206f
C1568 CSoutput.n178 gnd 2.3294f
C1569 CSoutput.n179 gnd 0.865206f
C1570 CSoutput.n180 gnd 0.865206f
C1571 CSoutput.t198 gnd 1.08151f
C1572 CSoutput.n181 gnd 0.865206f
C1573 CSoutput.n182 gnd 0.865206f
C1574 CSoutput.n186 gnd 0.865206f
C1575 CSoutput.n190 gnd 0.865206f
C1576 CSoutput.n191 gnd 0.865206f
C1577 CSoutput.n193 gnd 0.865206f
C1578 CSoutput.n198 gnd 0.865206f
C1579 CSoutput.n200 gnd 0.865206f
C1580 CSoutput.n201 gnd 0.865206f
C1581 CSoutput.n203 gnd 0.865206f
C1582 CSoutput.n204 gnd 0.865206f
C1583 CSoutput.n206 gnd 0.865206f
C1584 CSoutput.n207 gnd 0.648904f
C1585 CSoutput.n209 gnd 0.865206f
C1586 CSoutput.n210 gnd 0.648904f
C1587 CSoutput.n211 gnd 0.865206f
C1588 CSoutput.n212 gnd 0.865206f
C1589 CSoutput.n213 gnd 2.3294f
C1590 CSoutput.n214 gnd 0.865206f
C1591 CSoutput.n215 gnd 0.865206f
C1592 CSoutput.t206 gnd 1.08151f
C1593 CSoutput.n216 gnd 0.865206f
C1594 CSoutput.n217 gnd 2.3294f
C1595 CSoutput.n219 gnd 0.865206f
C1596 CSoutput.n220 gnd 0.865206f
C1597 CSoutput.n222 gnd 0.865206f
C1598 CSoutput.n223 gnd 0.865206f
C1599 CSoutput.t211 gnd 14.2219f
C1600 CSoutput.t205 gnd 14.4575f
C1601 CSoutput.n229 gnd 2.71428f
C1602 CSoutput.n230 gnd 11.057f
C1603 CSoutput.n231 gnd 11.5196f
C1604 CSoutput.n236 gnd 2.94029f
C1605 CSoutput.n242 gnd 0.865206f
C1606 CSoutput.n244 gnd 0.865206f
C1607 CSoutput.n246 gnd 0.865206f
C1608 CSoutput.n248 gnd 0.865206f
C1609 CSoutput.n250 gnd 0.865206f
C1610 CSoutput.n256 gnd 0.865206f
C1611 CSoutput.n263 gnd 1.58732f
C1612 CSoutput.n264 gnd 1.58732f
C1613 CSoutput.n265 gnd 0.865206f
C1614 CSoutput.n266 gnd 0.865206f
C1615 CSoutput.n268 gnd 0.648904f
C1616 CSoutput.n269 gnd 0.555728f
C1617 CSoutput.n271 gnd 0.648904f
C1618 CSoutput.n272 gnd 0.555728f
C1619 CSoutput.n273 gnd 0.648904f
C1620 CSoutput.n275 gnd 0.865206f
C1621 CSoutput.n277 gnd 2.3294f
C1622 CSoutput.n278 gnd 2.71428f
C1623 CSoutput.n279 gnd 10.1696f
C1624 CSoutput.n281 gnd 0.648904f
C1625 CSoutput.n282 gnd 1.66967f
C1626 CSoutput.n283 gnd 0.648904f
C1627 CSoutput.n285 gnd 0.865206f
C1628 CSoutput.n287 gnd 2.3294f
C1629 CSoutput.n288 gnd 5.07327f
C1630 CSoutput.t18 gnd 0.061008f
C1631 CSoutput.t10 gnd 0.061008f
C1632 CSoutput.n289 gnd 0.472345f
C1633 CSoutput.t68 gnd 0.061008f
C1634 CSoutput.t2 gnd 0.061008f
C1635 CSoutput.n290 gnd 0.471503f
C1636 CSoutput.n291 gnd 0.478574f
C1637 CSoutput.t45 gnd 0.061008f
C1638 CSoutput.t173 gnd 0.061008f
C1639 CSoutput.n292 gnd 0.471503f
C1640 CSoutput.n293 gnd 0.235821f
C1641 CSoutput.t22 gnd 0.061008f
C1642 CSoutput.t174 gnd 0.061008f
C1643 CSoutput.n294 gnd 0.471503f
C1644 CSoutput.n295 gnd 0.235821f
C1645 CSoutput.t67 gnd 0.061008f
C1646 CSoutput.t51 gnd 0.061008f
C1647 CSoutput.n296 gnd 0.471503f
C1648 CSoutput.n297 gnd 0.235821f
C1649 CSoutput.t190 gnd 0.061008f
C1650 CSoutput.t16 gnd 0.061008f
C1651 CSoutput.n298 gnd 0.471503f
C1652 CSoutput.n299 gnd 0.235821f
C1653 CSoutput.t6 gnd 0.061008f
C1654 CSoutput.t86 gnd 0.061008f
C1655 CSoutput.n300 gnd 0.471503f
C1656 CSoutput.n301 gnd 0.235821f
C1657 CSoutput.t46 gnd 0.061008f
C1658 CSoutput.t42 gnd 0.061008f
C1659 CSoutput.n302 gnd 0.471503f
C1660 CSoutput.n303 gnd 0.235821f
C1661 CSoutput.t72 gnd 0.061008f
C1662 CSoutput.t77 gnd 0.061008f
C1663 CSoutput.n304 gnd 0.471503f
C1664 CSoutput.n305 gnd 0.235821f
C1665 CSoutput.t66 gnd 0.061008f
C1666 CSoutput.t89 gnd 0.061008f
C1667 CSoutput.n306 gnd 0.471503f
C1668 CSoutput.n307 gnd 0.432442f
C1669 CSoutput.t90 gnd 0.061008f
C1670 CSoutput.t63 gnd 0.061008f
C1671 CSoutput.n308 gnd 0.472345f
C1672 CSoutput.t14 gnd 0.061008f
C1673 CSoutput.t178 gnd 0.061008f
C1674 CSoutput.n309 gnd 0.471503f
C1675 CSoutput.n310 gnd 0.478574f
C1676 CSoutput.t69 gnd 0.061008f
C1677 CSoutput.t55 gnd 0.061008f
C1678 CSoutput.n311 gnd 0.471503f
C1679 CSoutput.n312 gnd 0.235821f
C1680 CSoutput.t19 gnd 0.061008f
C1681 CSoutput.t191 gnd 0.061008f
C1682 CSoutput.n313 gnd 0.471503f
C1683 CSoutput.n314 gnd 0.235821f
C1684 CSoutput.t167 gnd 0.061008f
C1685 CSoutput.t40 gnd 0.061008f
C1686 CSoutput.n315 gnd 0.471503f
C1687 CSoutput.n316 gnd 0.235821f
C1688 CSoutput.t60 gnd 0.061008f
C1689 CSoutput.t181 gnd 0.061008f
C1690 CSoutput.n317 gnd 0.471503f
C1691 CSoutput.n318 gnd 0.235821f
C1692 CSoutput.t11 gnd 0.061008f
C1693 CSoutput.t43 gnd 0.061008f
C1694 CSoutput.n319 gnd 0.471503f
C1695 CSoutput.n320 gnd 0.235821f
C1696 CSoutput.t91 gnd 0.061008f
C1697 CSoutput.t15 gnd 0.061008f
C1698 CSoutput.n321 gnd 0.471503f
C1699 CSoutput.n322 gnd 0.235821f
C1700 CSoutput.t34 gnd 0.061008f
C1701 CSoutput.t0 gnd 0.061008f
C1702 CSoutput.n323 gnd 0.471503f
C1703 CSoutput.n324 gnd 0.235821f
C1704 CSoutput.t83 gnd 0.061008f
C1705 CSoutput.t82 gnd 0.061008f
C1706 CSoutput.n325 gnd 0.471503f
C1707 CSoutput.n326 gnd 0.351669f
C1708 CSoutput.n327 gnd 0.443452f
C1709 CSoutput.t53 gnd 0.061008f
C1710 CSoutput.t47 gnd 0.061008f
C1711 CSoutput.n328 gnd 0.472345f
C1712 CSoutput.t35 gnd 0.061008f
C1713 CSoutput.t1 gnd 0.061008f
C1714 CSoutput.n329 gnd 0.471503f
C1715 CSoutput.n330 gnd 0.478574f
C1716 CSoutput.t8 gnd 0.061008f
C1717 CSoutput.t172 gnd 0.061008f
C1718 CSoutput.n331 gnd 0.471503f
C1719 CSoutput.n332 gnd 0.235821f
C1720 CSoutput.t29 gnd 0.061008f
C1721 CSoutput.t164 gnd 0.061008f
C1722 CSoutput.n333 gnd 0.471503f
C1723 CSoutput.n334 gnd 0.235821f
C1724 CSoutput.t80 gnd 0.061008f
C1725 CSoutput.t87 gnd 0.061008f
C1726 CSoutput.n335 gnd 0.471503f
C1727 CSoutput.n336 gnd 0.235821f
C1728 CSoutput.t23 gnd 0.061008f
C1729 CSoutput.t54 gnd 0.061008f
C1730 CSoutput.n337 gnd 0.471503f
C1731 CSoutput.n338 gnd 0.235821f
C1732 CSoutput.t79 gnd 0.061008f
C1733 CSoutput.t21 gnd 0.061008f
C1734 CSoutput.n339 gnd 0.471503f
C1735 CSoutput.n340 gnd 0.235821f
C1736 CSoutput.t52 gnd 0.061008f
C1737 CSoutput.t26 gnd 0.061008f
C1738 CSoutput.n341 gnd 0.471503f
C1739 CSoutput.n342 gnd 0.235821f
C1740 CSoutput.t85 gnd 0.061008f
C1741 CSoutput.t9 gnd 0.061008f
C1742 CSoutput.n343 gnd 0.471503f
C1743 CSoutput.n344 gnd 0.235821f
C1744 CSoutput.t183 gnd 0.061008f
C1745 CSoutput.t39 gnd 0.061008f
C1746 CSoutput.n345 gnd 0.471501f
C1747 CSoutput.n346 gnd 0.351671f
C1748 CSoutput.n347 gnd 0.495666f
C1749 CSoutput.n348 gnd 13.6482f
C1750 CSoutput.t122 gnd 0.053382f
C1751 CSoutput.t160 gnd 0.053382f
C1752 CSoutput.n349 gnd 0.473281f
C1753 CSoutput.t116 gnd 0.053382f
C1754 CSoutput.t121 gnd 0.053382f
C1755 CSoutput.n350 gnd 0.471703f
C1756 CSoutput.n351 gnd 0.439539f
C1757 CSoutput.t110 gnd 0.053382f
C1758 CSoutput.t125 gnd 0.053382f
C1759 CSoutput.n352 gnd 0.471703f
C1760 CSoutput.n353 gnd 0.216672f
C1761 CSoutput.t134 gnd 0.053382f
C1762 CSoutput.t117 gnd 0.053382f
C1763 CSoutput.n354 gnd 0.471703f
C1764 CSoutput.n355 gnd 0.216672f
C1765 CSoutput.t124 gnd 0.053382f
C1766 CSoutput.t153 gnd 0.053382f
C1767 CSoutput.n356 gnd 0.471703f
C1768 CSoutput.n357 gnd 0.216672f
C1769 CSoutput.t131 gnd 0.053382f
C1770 CSoutput.t138 gnd 0.053382f
C1771 CSoutput.n358 gnd 0.471703f
C1772 CSoutput.n359 gnd 0.399639f
C1773 CSoutput.t157 gnd 0.053382f
C1774 CSoutput.t92 gnd 0.053382f
C1775 CSoutput.n360 gnd 0.473281f
C1776 CSoutput.t101 gnd 0.053382f
C1777 CSoutput.t151 gnd 0.053382f
C1778 CSoutput.n361 gnd 0.471703f
C1779 CSoutput.n362 gnd 0.439539f
C1780 CSoutput.t94 gnd 0.053382f
C1781 CSoutput.t146 gnd 0.053382f
C1782 CSoutput.n363 gnd 0.471703f
C1783 CSoutput.n364 gnd 0.216672f
C1784 CSoutput.t152 gnd 0.053382f
C1785 CSoutput.t93 gnd 0.053382f
C1786 CSoutput.n365 gnd 0.471703f
C1787 CSoutput.n366 gnd 0.216672f
C1788 CSoutput.t140 gnd 0.053382f
C1789 CSoutput.t128 gnd 0.053382f
C1790 CSoutput.n367 gnd 0.471703f
C1791 CSoutput.n368 gnd 0.216672f
C1792 CSoutput.t95 gnd 0.053382f
C1793 CSoutput.t141 gnd 0.053382f
C1794 CSoutput.n369 gnd 0.471703f
C1795 CSoutput.n370 gnd 0.328954f
C1796 CSoutput.n371 gnd 0.414914f
C1797 CSoutput.t102 gnd 0.053382f
C1798 CSoutput.t154 gnd 0.053382f
C1799 CSoutput.n372 gnd 0.473281f
C1800 CSoutput.t115 gnd 0.053382f
C1801 CSoutput.t118 gnd 0.053382f
C1802 CSoutput.n373 gnd 0.471703f
C1803 CSoutput.n374 gnd 0.439539f
C1804 CSoutput.t96 gnd 0.053382f
C1805 CSoutput.t143 gnd 0.053382f
C1806 CSoutput.n375 gnd 0.471703f
C1807 CSoutput.n376 gnd 0.216672f
C1808 CSoutput.t123 gnd 0.053382f
C1809 CSoutput.t103 gnd 0.053382f
C1810 CSoutput.n377 gnd 0.471703f
C1811 CSoutput.n378 gnd 0.216672f
C1812 CSoutput.t108 gnd 0.053382f
C1813 CSoutput.t163 gnd 0.053382f
C1814 CSoutput.n379 gnd 0.471703f
C1815 CSoutput.n380 gnd 0.216672f
C1816 CSoutput.t109 gnd 0.053382f
C1817 CSoutput.t113 gnd 0.053382f
C1818 CSoutput.n381 gnd 0.471703f
C1819 CSoutput.n382 gnd 0.328954f
C1820 CSoutput.n383 gnd 0.445552f
C1821 CSoutput.n384 gnd 13.257f
C1822 CSoutput.t112 gnd 0.053382f
C1823 CSoutput.t142 gnd 0.053382f
C1824 CSoutput.n385 gnd 0.473281f
C1825 CSoutput.t139 gnd 0.053382f
C1826 CSoutput.t127 gnd 0.053382f
C1827 CSoutput.n386 gnd 0.471703f
C1828 CSoutput.n387 gnd 0.439539f
C1829 CSoutput.t145 gnd 0.053382f
C1830 CSoutput.t119 gnd 0.053382f
C1831 CSoutput.n388 gnd 0.471703f
C1832 CSoutput.n389 gnd 0.216672f
C1833 CSoutput.t132 gnd 0.053382f
C1834 CSoutput.t155 gnd 0.053382f
C1835 CSoutput.n390 gnd 0.471703f
C1836 CSoutput.n391 gnd 0.216672f
C1837 CSoutput.t107 gnd 0.053382f
C1838 CSoutput.t144 gnd 0.053382f
C1839 CSoutput.n392 gnd 0.471703f
C1840 CSoutput.n393 gnd 0.216672f
C1841 CSoutput.t100 gnd 0.053382f
C1842 CSoutput.t147 gnd 0.053382f
C1843 CSoutput.n394 gnd 0.471703f
C1844 CSoutput.n395 gnd 0.399639f
C1845 CSoutput.t104 gnd 0.053382f
C1846 CSoutput.t99 gnd 0.053382f
C1847 CSoutput.n396 gnd 0.473281f
C1848 CSoutput.t97 gnd 0.053382f
C1849 CSoutput.t161 gnd 0.053382f
C1850 CSoutput.n397 gnd 0.471703f
C1851 CSoutput.n398 gnd 0.439539f
C1852 CSoutput.t162 gnd 0.053382f
C1853 CSoutput.t105 gnd 0.053382f
C1854 CSoutput.n399 gnd 0.471703f
C1855 CSoutput.n400 gnd 0.216672f
C1856 CSoutput.t106 gnd 0.053382f
C1857 CSoutput.t137 gnd 0.053382f
C1858 CSoutput.n401 gnd 0.471703f
C1859 CSoutput.n402 gnd 0.216672f
C1860 CSoutput.t136 gnd 0.053382f
C1861 CSoutput.t156 gnd 0.053382f
C1862 CSoutput.n403 gnd 0.471703f
C1863 CSoutput.n404 gnd 0.216672f
C1864 CSoutput.t159 gnd 0.053382f
C1865 CSoutput.t150 gnd 0.053382f
C1866 CSoutput.n405 gnd 0.471703f
C1867 CSoutput.n406 gnd 0.328954f
C1868 CSoutput.n407 gnd 0.414914f
C1869 CSoutput.t130 gnd 0.053382f
C1870 CSoutput.t148 gnd 0.053382f
C1871 CSoutput.n408 gnd 0.473281f
C1872 CSoutput.t111 gnd 0.053382f
C1873 CSoutput.t120 gnd 0.053382f
C1874 CSoutput.n409 gnd 0.471703f
C1875 CSoutput.n410 gnd 0.439539f
C1876 CSoutput.t126 gnd 0.053382f
C1877 CSoutput.t135 gnd 0.053382f
C1878 CSoutput.n411 gnd 0.471703f
C1879 CSoutput.n412 gnd 0.216672f
C1880 CSoutput.t149 gnd 0.053382f
C1881 CSoutput.t129 gnd 0.053382f
C1882 CSoutput.n413 gnd 0.471703f
C1883 CSoutput.n414 gnd 0.216672f
C1884 CSoutput.t133 gnd 0.053382f
C1885 CSoutput.t158 gnd 0.053382f
C1886 CSoutput.n415 gnd 0.471703f
C1887 CSoutput.n416 gnd 0.216672f
C1888 CSoutput.t98 gnd 0.053382f
C1889 CSoutput.t114 gnd 0.053382f
C1890 CSoutput.n417 gnd 0.471703f
C1891 CSoutput.n418 gnd 0.328954f
C1892 CSoutput.n419 gnd 0.445552f
C1893 CSoutput.n420 gnd 7.88002f
C1894 CSoutput.n421 gnd 14.761401f
C1895 commonsourceibias.n0 gnd 0.01231f
C1896 commonsourceibias.t89 gnd 0.186396f
C1897 commonsourceibias.t51 gnd 0.17235f
C1898 commonsourceibias.n1 gnd 0.068768f
C1899 commonsourceibias.n2 gnd 0.009225f
C1900 commonsourceibias.t95 gnd 0.17235f
C1901 commonsourceibias.n3 gnd 0.007462f
C1902 commonsourceibias.n4 gnd 0.009225f
C1903 commonsourceibias.t90 gnd 0.17235f
C1904 commonsourceibias.n5 gnd 0.008906f
C1905 commonsourceibias.n6 gnd 0.009225f
C1906 commonsourceibias.t101 gnd 0.17235f
C1907 commonsourceibias.n7 gnd 0.068768f
C1908 commonsourceibias.t86 gnd 0.17235f
C1909 commonsourceibias.n8 gnd 0.007451f
C1910 commonsourceibias.n9 gnd 0.01231f
C1911 commonsourceibias.t20 gnd 0.186396f
C1912 commonsourceibias.t28 gnd 0.17235f
C1913 commonsourceibias.n10 gnd 0.068768f
C1914 commonsourceibias.n11 gnd 0.009225f
C1915 commonsourceibias.t2 gnd 0.17235f
C1916 commonsourceibias.n12 gnd 0.007462f
C1917 commonsourceibias.n13 gnd 0.009225f
C1918 commonsourceibias.t18 gnd 0.17235f
C1919 commonsourceibias.n14 gnd 0.008906f
C1920 commonsourceibias.n15 gnd 0.009225f
C1921 commonsourceibias.t32 gnd 0.17235f
C1922 commonsourceibias.n16 gnd 0.068768f
C1923 commonsourceibias.t14 gnd 0.17235f
C1924 commonsourceibias.n17 gnd 0.007451f
C1925 commonsourceibias.n18 gnd 0.009225f
C1926 commonsourceibias.t12 gnd 0.17235f
C1927 commonsourceibias.t44 gnd 0.17235f
C1928 commonsourceibias.n19 gnd 0.068768f
C1929 commonsourceibias.n20 gnd 0.009225f
C1930 commonsourceibias.t22 gnd 0.17235f
C1931 commonsourceibias.n21 gnd 0.068768f
C1932 commonsourceibias.n22 gnd 0.009225f
C1933 commonsourceibias.t6 gnd 0.17235f
C1934 commonsourceibias.n23 gnd 0.068768f
C1935 commonsourceibias.n24 gnd 0.046441f
C1936 commonsourceibias.t8 gnd 0.17235f
C1937 commonsourceibias.t34 gnd 0.194477f
C1938 commonsourceibias.n25 gnd 0.079804f
C1939 commonsourceibias.n26 gnd 0.082619f
C1940 commonsourceibias.n27 gnd 0.01137f
C1941 commonsourceibias.n28 gnd 0.012578f
C1942 commonsourceibias.n29 gnd 0.009225f
C1943 commonsourceibias.n30 gnd 0.009225f
C1944 commonsourceibias.n31 gnd 0.012496f
C1945 commonsourceibias.n32 gnd 0.007462f
C1946 commonsourceibias.n33 gnd 0.012651f
C1947 commonsourceibias.n34 gnd 0.009225f
C1948 commonsourceibias.n35 gnd 0.009225f
C1949 commonsourceibias.n36 gnd 0.012728f
C1950 commonsourceibias.n37 gnd 0.010975f
C1951 commonsourceibias.n38 gnd 0.008906f
C1952 commonsourceibias.n39 gnd 0.009225f
C1953 commonsourceibias.n40 gnd 0.009225f
C1954 commonsourceibias.n41 gnd 0.011283f
C1955 commonsourceibias.n42 gnd 0.012665f
C1956 commonsourceibias.n43 gnd 0.068768f
C1957 commonsourceibias.n44 gnd 0.01258f
C1958 commonsourceibias.n45 gnd 0.009225f
C1959 commonsourceibias.n46 gnd 0.009225f
C1960 commonsourceibias.n47 gnd 0.009225f
C1961 commonsourceibias.n48 gnd 0.01258f
C1962 commonsourceibias.n49 gnd 0.068768f
C1963 commonsourceibias.n50 gnd 0.012665f
C1964 commonsourceibias.n51 gnd 0.011283f
C1965 commonsourceibias.n52 gnd 0.009225f
C1966 commonsourceibias.n53 gnd 0.009225f
C1967 commonsourceibias.n54 gnd 0.009225f
C1968 commonsourceibias.n55 gnd 0.010975f
C1969 commonsourceibias.n56 gnd 0.012728f
C1970 commonsourceibias.n57 gnd 0.068768f
C1971 commonsourceibias.n58 gnd 0.012651f
C1972 commonsourceibias.n59 gnd 0.009225f
C1973 commonsourceibias.n60 gnd 0.009225f
C1974 commonsourceibias.n61 gnd 0.009225f
C1975 commonsourceibias.n62 gnd 0.012496f
C1976 commonsourceibias.n63 gnd 0.068768f
C1977 commonsourceibias.n64 gnd 0.012578f
C1978 commonsourceibias.n65 gnd 0.01137f
C1979 commonsourceibias.n66 gnd 0.009225f
C1980 commonsourceibias.n67 gnd 0.009225f
C1981 commonsourceibias.n68 gnd 0.009358f
C1982 commonsourceibias.n69 gnd 0.009674f
C1983 commonsourceibias.n70 gnd 0.082281f
C1984 commonsourceibias.n71 gnd 0.091278f
C1985 commonsourceibias.t21 gnd 0.019906f
C1986 commonsourceibias.t29 gnd 0.019906f
C1987 commonsourceibias.n72 gnd 0.1759f
C1988 commonsourceibias.n73 gnd 0.151991f
C1989 commonsourceibias.t3 gnd 0.019906f
C1990 commonsourceibias.t19 gnd 0.019906f
C1991 commonsourceibias.n74 gnd 0.1759f
C1992 commonsourceibias.n75 gnd 0.080798f
C1993 commonsourceibias.t33 gnd 0.019906f
C1994 commonsourceibias.t15 gnd 0.019906f
C1995 commonsourceibias.n76 gnd 0.1759f
C1996 commonsourceibias.n77 gnd 0.067503f
C1997 commonsourceibias.t9 gnd 0.019906f
C1998 commonsourceibias.t35 gnd 0.019906f
C1999 commonsourceibias.n78 gnd 0.176489f
C2000 commonsourceibias.t23 gnd 0.019906f
C2001 commonsourceibias.t7 gnd 0.019906f
C2002 commonsourceibias.n79 gnd 0.1759f
C2003 commonsourceibias.n80 gnd 0.163906f
C2004 commonsourceibias.t13 gnd 0.019906f
C2005 commonsourceibias.t45 gnd 0.019906f
C2006 commonsourceibias.n81 gnd 0.1759f
C2007 commonsourceibias.n82 gnd 0.067503f
C2008 commonsourceibias.n83 gnd 0.081739f
C2009 commonsourceibias.n84 gnd 0.009225f
C2010 commonsourceibias.t77 gnd 0.17235f
C2011 commonsourceibias.t94 gnd 0.17235f
C2012 commonsourceibias.n85 gnd 0.068768f
C2013 commonsourceibias.n86 gnd 0.009225f
C2014 commonsourceibias.t87 gnd 0.17235f
C2015 commonsourceibias.n87 gnd 0.068768f
C2016 commonsourceibias.n88 gnd 0.009225f
C2017 commonsourceibias.t58 gnd 0.17235f
C2018 commonsourceibias.n89 gnd 0.068768f
C2019 commonsourceibias.n90 gnd 0.046441f
C2020 commonsourceibias.t80 gnd 0.17235f
C2021 commonsourceibias.t73 gnd 0.194477f
C2022 commonsourceibias.n91 gnd 0.079804f
C2023 commonsourceibias.n92 gnd 0.082619f
C2024 commonsourceibias.n93 gnd 0.01137f
C2025 commonsourceibias.n94 gnd 0.012578f
C2026 commonsourceibias.n95 gnd 0.009225f
C2027 commonsourceibias.n96 gnd 0.009225f
C2028 commonsourceibias.n97 gnd 0.012496f
C2029 commonsourceibias.n98 gnd 0.007462f
C2030 commonsourceibias.n99 gnd 0.012651f
C2031 commonsourceibias.n100 gnd 0.009225f
C2032 commonsourceibias.n101 gnd 0.009225f
C2033 commonsourceibias.n102 gnd 0.012728f
C2034 commonsourceibias.n103 gnd 0.010975f
C2035 commonsourceibias.n104 gnd 0.008906f
C2036 commonsourceibias.n105 gnd 0.009225f
C2037 commonsourceibias.n106 gnd 0.009225f
C2038 commonsourceibias.n107 gnd 0.011283f
C2039 commonsourceibias.n108 gnd 0.012665f
C2040 commonsourceibias.n109 gnd 0.068768f
C2041 commonsourceibias.n110 gnd 0.01258f
C2042 commonsourceibias.n111 gnd 0.009181f
C2043 commonsourceibias.n112 gnd 0.066685f
C2044 commonsourceibias.n113 gnd 0.009181f
C2045 commonsourceibias.n114 gnd 0.01258f
C2046 commonsourceibias.n115 gnd 0.068768f
C2047 commonsourceibias.n116 gnd 0.012665f
C2048 commonsourceibias.n117 gnd 0.011283f
C2049 commonsourceibias.n118 gnd 0.009225f
C2050 commonsourceibias.n119 gnd 0.009225f
C2051 commonsourceibias.n120 gnd 0.009225f
C2052 commonsourceibias.n121 gnd 0.010975f
C2053 commonsourceibias.n122 gnd 0.012728f
C2054 commonsourceibias.n123 gnd 0.068768f
C2055 commonsourceibias.n124 gnd 0.012651f
C2056 commonsourceibias.n125 gnd 0.009225f
C2057 commonsourceibias.n126 gnd 0.009225f
C2058 commonsourceibias.n127 gnd 0.009225f
C2059 commonsourceibias.n128 gnd 0.012496f
C2060 commonsourceibias.n129 gnd 0.068768f
C2061 commonsourceibias.n130 gnd 0.012578f
C2062 commonsourceibias.n131 gnd 0.01137f
C2063 commonsourceibias.n132 gnd 0.009225f
C2064 commonsourceibias.n133 gnd 0.009225f
C2065 commonsourceibias.n134 gnd 0.009358f
C2066 commonsourceibias.n135 gnd 0.009674f
C2067 commonsourceibias.n136 gnd 0.082281f
C2068 commonsourceibias.n137 gnd 0.053268f
C2069 commonsourceibias.n138 gnd 0.01231f
C2070 commonsourceibias.t54 gnd 0.186396f
C2071 commonsourceibias.t119 gnd 0.17235f
C2072 commonsourceibias.n139 gnd 0.068768f
C2073 commonsourceibias.n140 gnd 0.009225f
C2074 commonsourceibias.t110 gnd 0.17235f
C2075 commonsourceibias.n141 gnd 0.007462f
C2076 commonsourceibias.n142 gnd 0.009225f
C2077 commonsourceibias.t60 gnd 0.17235f
C2078 commonsourceibias.n143 gnd 0.008906f
C2079 commonsourceibias.n144 gnd 0.009225f
C2080 commonsourceibias.t117 gnd 0.17235f
C2081 commonsourceibias.n145 gnd 0.068768f
C2082 commonsourceibias.t65 gnd 0.17235f
C2083 commonsourceibias.n146 gnd 0.007451f
C2084 commonsourceibias.n147 gnd 0.009225f
C2085 commonsourceibias.t59 gnd 0.17235f
C2086 commonsourceibias.t118 gnd 0.17235f
C2087 commonsourceibias.n148 gnd 0.068768f
C2088 commonsourceibias.n149 gnd 0.009225f
C2089 commonsourceibias.t71 gnd 0.17235f
C2090 commonsourceibias.n150 gnd 0.068768f
C2091 commonsourceibias.n151 gnd 0.009225f
C2092 commonsourceibias.t83 gnd 0.17235f
C2093 commonsourceibias.n152 gnd 0.068768f
C2094 commonsourceibias.n153 gnd 0.046441f
C2095 commonsourceibias.t116 gnd 0.17235f
C2096 commonsourceibias.t70 gnd 0.194477f
C2097 commonsourceibias.n154 gnd 0.079804f
C2098 commonsourceibias.n155 gnd 0.082619f
C2099 commonsourceibias.n156 gnd 0.01137f
C2100 commonsourceibias.n157 gnd 0.012578f
C2101 commonsourceibias.n158 gnd 0.009225f
C2102 commonsourceibias.n159 gnd 0.009225f
C2103 commonsourceibias.n160 gnd 0.012496f
C2104 commonsourceibias.n161 gnd 0.007462f
C2105 commonsourceibias.n162 gnd 0.012651f
C2106 commonsourceibias.n163 gnd 0.009225f
C2107 commonsourceibias.n164 gnd 0.009225f
C2108 commonsourceibias.n165 gnd 0.012728f
C2109 commonsourceibias.n166 gnd 0.010975f
C2110 commonsourceibias.n167 gnd 0.008906f
C2111 commonsourceibias.n168 gnd 0.009225f
C2112 commonsourceibias.n169 gnd 0.009225f
C2113 commonsourceibias.n170 gnd 0.011283f
C2114 commonsourceibias.n171 gnd 0.012665f
C2115 commonsourceibias.n172 gnd 0.068768f
C2116 commonsourceibias.n173 gnd 0.01258f
C2117 commonsourceibias.n174 gnd 0.009225f
C2118 commonsourceibias.n175 gnd 0.009225f
C2119 commonsourceibias.n176 gnd 0.009225f
C2120 commonsourceibias.n177 gnd 0.01258f
C2121 commonsourceibias.n178 gnd 0.068768f
C2122 commonsourceibias.n179 gnd 0.012665f
C2123 commonsourceibias.n180 gnd 0.011283f
C2124 commonsourceibias.n181 gnd 0.009225f
C2125 commonsourceibias.n182 gnd 0.009225f
C2126 commonsourceibias.n183 gnd 0.009225f
C2127 commonsourceibias.n184 gnd 0.010975f
C2128 commonsourceibias.n185 gnd 0.012728f
C2129 commonsourceibias.n186 gnd 0.068768f
C2130 commonsourceibias.n187 gnd 0.012651f
C2131 commonsourceibias.n188 gnd 0.009225f
C2132 commonsourceibias.n189 gnd 0.009225f
C2133 commonsourceibias.n190 gnd 0.009225f
C2134 commonsourceibias.n191 gnd 0.012496f
C2135 commonsourceibias.n192 gnd 0.068768f
C2136 commonsourceibias.n193 gnd 0.012578f
C2137 commonsourceibias.n194 gnd 0.01137f
C2138 commonsourceibias.n195 gnd 0.009225f
C2139 commonsourceibias.n196 gnd 0.009225f
C2140 commonsourceibias.n197 gnd 0.009358f
C2141 commonsourceibias.n198 gnd 0.009674f
C2142 commonsourceibias.n199 gnd 0.082281f
C2143 commonsourceibias.n200 gnd 0.028001f
C2144 commonsourceibias.n201 gnd 0.147196f
C2145 commonsourceibias.n202 gnd 0.01231f
C2146 commonsourceibias.t57 gnd 0.17235f
C2147 commonsourceibias.n203 gnd 0.068768f
C2148 commonsourceibias.n204 gnd 0.009225f
C2149 commonsourceibias.t96 gnd 0.17235f
C2150 commonsourceibias.n205 gnd 0.007462f
C2151 commonsourceibias.n206 gnd 0.009225f
C2152 commonsourceibias.t93 gnd 0.17235f
C2153 commonsourceibias.n207 gnd 0.008906f
C2154 commonsourceibias.n208 gnd 0.009225f
C2155 commonsourceibias.t115 gnd 0.17235f
C2156 commonsourceibias.n209 gnd 0.068768f
C2157 commonsourceibias.t68 gnd 0.17235f
C2158 commonsourceibias.n210 gnd 0.007451f
C2159 commonsourceibias.n211 gnd 0.009225f
C2160 commonsourceibias.t88 gnd 0.17235f
C2161 commonsourceibias.t108 gnd 0.17235f
C2162 commonsourceibias.n212 gnd 0.068768f
C2163 commonsourceibias.n213 gnd 0.009225f
C2164 commonsourceibias.t103 gnd 0.17235f
C2165 commonsourceibias.n214 gnd 0.068768f
C2166 commonsourceibias.n215 gnd 0.009225f
C2167 commonsourceibias.t48 gnd 0.17235f
C2168 commonsourceibias.n216 gnd 0.068768f
C2169 commonsourceibias.n217 gnd 0.046441f
C2170 commonsourceibias.t102 gnd 0.17235f
C2171 commonsourceibias.t98 gnd 0.194477f
C2172 commonsourceibias.n218 gnd 0.079804f
C2173 commonsourceibias.n219 gnd 0.082619f
C2174 commonsourceibias.n220 gnd 0.01137f
C2175 commonsourceibias.n221 gnd 0.012578f
C2176 commonsourceibias.n222 gnd 0.009225f
C2177 commonsourceibias.n223 gnd 0.009225f
C2178 commonsourceibias.n224 gnd 0.012496f
C2179 commonsourceibias.n225 gnd 0.007462f
C2180 commonsourceibias.n226 gnd 0.012651f
C2181 commonsourceibias.n227 gnd 0.009225f
C2182 commonsourceibias.n228 gnd 0.009225f
C2183 commonsourceibias.n229 gnd 0.012728f
C2184 commonsourceibias.n230 gnd 0.010975f
C2185 commonsourceibias.n231 gnd 0.008906f
C2186 commonsourceibias.n232 gnd 0.009225f
C2187 commonsourceibias.n233 gnd 0.009225f
C2188 commonsourceibias.n234 gnd 0.011283f
C2189 commonsourceibias.n235 gnd 0.012665f
C2190 commonsourceibias.n236 gnd 0.068768f
C2191 commonsourceibias.n237 gnd 0.01258f
C2192 commonsourceibias.n238 gnd 0.009225f
C2193 commonsourceibias.n239 gnd 0.009225f
C2194 commonsourceibias.n240 gnd 0.009225f
C2195 commonsourceibias.n241 gnd 0.01258f
C2196 commonsourceibias.n242 gnd 0.068768f
C2197 commonsourceibias.n243 gnd 0.012665f
C2198 commonsourceibias.n244 gnd 0.011283f
C2199 commonsourceibias.n245 gnd 0.009225f
C2200 commonsourceibias.n246 gnd 0.009225f
C2201 commonsourceibias.n247 gnd 0.009225f
C2202 commonsourceibias.n248 gnd 0.010975f
C2203 commonsourceibias.n249 gnd 0.012728f
C2204 commonsourceibias.n250 gnd 0.068768f
C2205 commonsourceibias.n251 gnd 0.012651f
C2206 commonsourceibias.n252 gnd 0.009225f
C2207 commonsourceibias.n253 gnd 0.009225f
C2208 commonsourceibias.n254 gnd 0.009225f
C2209 commonsourceibias.n255 gnd 0.012496f
C2210 commonsourceibias.n256 gnd 0.068768f
C2211 commonsourceibias.n257 gnd 0.012578f
C2212 commonsourceibias.n258 gnd 0.01137f
C2213 commonsourceibias.n259 gnd 0.009225f
C2214 commonsourceibias.n260 gnd 0.009225f
C2215 commonsourceibias.n261 gnd 0.009358f
C2216 commonsourceibias.n262 gnd 0.009674f
C2217 commonsourceibias.t109 gnd 0.186396f
C2218 commonsourceibias.n263 gnd 0.082281f
C2219 commonsourceibias.n264 gnd 0.028001f
C2220 commonsourceibias.n265 gnd 0.438243f
C2221 commonsourceibias.n266 gnd 0.01231f
C2222 commonsourceibias.t69 gnd 0.186396f
C2223 commonsourceibias.t99 gnd 0.17235f
C2224 commonsourceibias.n267 gnd 0.068768f
C2225 commonsourceibias.n268 gnd 0.009225f
C2226 commonsourceibias.t84 gnd 0.17235f
C2227 commonsourceibias.n269 gnd 0.007462f
C2228 commonsourceibias.n270 gnd 0.009225f
C2229 commonsourceibias.t72 gnd 0.17235f
C2230 commonsourceibias.n271 gnd 0.008906f
C2231 commonsourceibias.n272 gnd 0.009225f
C2232 commonsourceibias.t66 gnd 0.17235f
C2233 commonsourceibias.n273 gnd 0.007451f
C2234 commonsourceibias.n274 gnd 0.009225f
C2235 commonsourceibias.t56 gnd 0.17235f
C2236 commonsourceibias.t79 gnd 0.17235f
C2237 commonsourceibias.n275 gnd 0.068768f
C2238 commonsourceibias.n276 gnd 0.009225f
C2239 commonsourceibias.t67 gnd 0.17235f
C2240 commonsourceibias.n277 gnd 0.068768f
C2241 commonsourceibias.n278 gnd 0.009225f
C2242 commonsourceibias.t104 gnd 0.17235f
C2243 commonsourceibias.n279 gnd 0.068768f
C2244 commonsourceibias.n280 gnd 0.046441f
C2245 commonsourceibias.t64 gnd 0.17235f
C2246 commonsourceibias.t111 gnd 0.194477f
C2247 commonsourceibias.n281 gnd 0.079804f
C2248 commonsourceibias.n282 gnd 0.082619f
C2249 commonsourceibias.n283 gnd 0.01137f
C2250 commonsourceibias.n284 gnd 0.012578f
C2251 commonsourceibias.n285 gnd 0.009225f
C2252 commonsourceibias.n286 gnd 0.009225f
C2253 commonsourceibias.n287 gnd 0.012496f
C2254 commonsourceibias.n288 gnd 0.007462f
C2255 commonsourceibias.n289 gnd 0.012651f
C2256 commonsourceibias.n290 gnd 0.009225f
C2257 commonsourceibias.n291 gnd 0.009225f
C2258 commonsourceibias.n292 gnd 0.012728f
C2259 commonsourceibias.n293 gnd 0.010975f
C2260 commonsourceibias.n294 gnd 0.008906f
C2261 commonsourceibias.n295 gnd 0.009225f
C2262 commonsourceibias.n296 gnd 0.009225f
C2263 commonsourceibias.n297 gnd 0.011283f
C2264 commonsourceibias.n298 gnd 0.012665f
C2265 commonsourceibias.n299 gnd 0.068768f
C2266 commonsourceibias.n300 gnd 0.01258f
C2267 commonsourceibias.n301 gnd 0.009181f
C2268 commonsourceibias.t25 gnd 0.019906f
C2269 commonsourceibias.t5 gnd 0.019906f
C2270 commonsourceibias.n302 gnd 0.176489f
C2271 commonsourceibias.t31 gnd 0.019906f
C2272 commonsourceibias.t41 gnd 0.019906f
C2273 commonsourceibias.n303 gnd 0.1759f
C2274 commonsourceibias.n304 gnd 0.163906f
C2275 commonsourceibias.t11 gnd 0.019906f
C2276 commonsourceibias.t27 gnd 0.019906f
C2277 commonsourceibias.n305 gnd 0.1759f
C2278 commonsourceibias.n306 gnd 0.067503f
C2279 commonsourceibias.n307 gnd 0.01231f
C2280 commonsourceibias.t0 gnd 0.17235f
C2281 commonsourceibias.n308 gnd 0.068768f
C2282 commonsourceibias.n309 gnd 0.009225f
C2283 commonsourceibias.t16 gnd 0.17235f
C2284 commonsourceibias.n310 gnd 0.007462f
C2285 commonsourceibias.n311 gnd 0.009225f
C2286 commonsourceibias.t36 gnd 0.17235f
C2287 commonsourceibias.n312 gnd 0.008906f
C2288 commonsourceibias.n313 gnd 0.009225f
C2289 commonsourceibias.t42 gnd 0.17235f
C2290 commonsourceibias.n314 gnd 0.007451f
C2291 commonsourceibias.n315 gnd 0.009225f
C2292 commonsourceibias.t26 gnd 0.17235f
C2293 commonsourceibias.t10 gnd 0.17235f
C2294 commonsourceibias.n316 gnd 0.068768f
C2295 commonsourceibias.n317 gnd 0.009225f
C2296 commonsourceibias.t40 gnd 0.17235f
C2297 commonsourceibias.n318 gnd 0.068768f
C2298 commonsourceibias.n319 gnd 0.009225f
C2299 commonsourceibias.t30 gnd 0.17235f
C2300 commonsourceibias.n320 gnd 0.068768f
C2301 commonsourceibias.n321 gnd 0.046441f
C2302 commonsourceibias.t4 gnd 0.17235f
C2303 commonsourceibias.t24 gnd 0.194477f
C2304 commonsourceibias.n322 gnd 0.079804f
C2305 commonsourceibias.n323 gnd 0.082619f
C2306 commonsourceibias.n324 gnd 0.01137f
C2307 commonsourceibias.n325 gnd 0.012578f
C2308 commonsourceibias.n326 gnd 0.009225f
C2309 commonsourceibias.n327 gnd 0.009225f
C2310 commonsourceibias.n328 gnd 0.012496f
C2311 commonsourceibias.n329 gnd 0.007462f
C2312 commonsourceibias.n330 gnd 0.012651f
C2313 commonsourceibias.n331 gnd 0.009225f
C2314 commonsourceibias.n332 gnd 0.009225f
C2315 commonsourceibias.n333 gnd 0.012728f
C2316 commonsourceibias.n334 gnd 0.010975f
C2317 commonsourceibias.n335 gnd 0.008906f
C2318 commonsourceibias.n336 gnd 0.009225f
C2319 commonsourceibias.n337 gnd 0.009225f
C2320 commonsourceibias.n338 gnd 0.011283f
C2321 commonsourceibias.n339 gnd 0.012665f
C2322 commonsourceibias.n340 gnd 0.068768f
C2323 commonsourceibias.n341 gnd 0.01258f
C2324 commonsourceibias.n342 gnd 0.009225f
C2325 commonsourceibias.n343 gnd 0.009225f
C2326 commonsourceibias.n344 gnd 0.009225f
C2327 commonsourceibias.n345 gnd 0.01258f
C2328 commonsourceibias.n346 gnd 0.068768f
C2329 commonsourceibias.n347 gnd 0.012665f
C2330 commonsourceibias.t46 gnd 0.17235f
C2331 commonsourceibias.n348 gnd 0.068768f
C2332 commonsourceibias.n349 gnd 0.011283f
C2333 commonsourceibias.n350 gnd 0.009225f
C2334 commonsourceibias.n351 gnd 0.009225f
C2335 commonsourceibias.n352 gnd 0.009225f
C2336 commonsourceibias.n353 gnd 0.010975f
C2337 commonsourceibias.n354 gnd 0.012728f
C2338 commonsourceibias.n355 gnd 0.068768f
C2339 commonsourceibias.n356 gnd 0.012651f
C2340 commonsourceibias.n357 gnd 0.009225f
C2341 commonsourceibias.n358 gnd 0.009225f
C2342 commonsourceibias.n359 gnd 0.009225f
C2343 commonsourceibias.n360 gnd 0.012496f
C2344 commonsourceibias.n361 gnd 0.068768f
C2345 commonsourceibias.n362 gnd 0.012578f
C2346 commonsourceibias.n363 gnd 0.01137f
C2347 commonsourceibias.n364 gnd 0.009225f
C2348 commonsourceibias.n365 gnd 0.009225f
C2349 commonsourceibias.n366 gnd 0.009358f
C2350 commonsourceibias.n367 gnd 0.009674f
C2351 commonsourceibias.t38 gnd 0.186396f
C2352 commonsourceibias.n368 gnd 0.082281f
C2353 commonsourceibias.n369 gnd 0.091278f
C2354 commonsourceibias.t1 gnd 0.019906f
C2355 commonsourceibias.t39 gnd 0.019906f
C2356 commonsourceibias.n370 gnd 0.1759f
C2357 commonsourceibias.n371 gnd 0.151991f
C2358 commonsourceibias.t37 gnd 0.019906f
C2359 commonsourceibias.t17 gnd 0.019906f
C2360 commonsourceibias.n372 gnd 0.1759f
C2361 commonsourceibias.n373 gnd 0.080798f
C2362 commonsourceibias.t43 gnd 0.019906f
C2363 commonsourceibias.t47 gnd 0.019906f
C2364 commonsourceibias.n374 gnd 0.1759f
C2365 commonsourceibias.n375 gnd 0.067503f
C2366 commonsourceibias.n376 gnd 0.081739f
C2367 commonsourceibias.n377 gnd 0.066685f
C2368 commonsourceibias.n378 gnd 0.009181f
C2369 commonsourceibias.n379 gnd 0.01258f
C2370 commonsourceibias.n380 gnd 0.068768f
C2371 commonsourceibias.n381 gnd 0.012665f
C2372 commonsourceibias.t92 gnd 0.17235f
C2373 commonsourceibias.n382 gnd 0.068768f
C2374 commonsourceibias.n383 gnd 0.011283f
C2375 commonsourceibias.n384 gnd 0.009225f
C2376 commonsourceibias.n385 gnd 0.009225f
C2377 commonsourceibias.n386 gnd 0.009225f
C2378 commonsourceibias.n387 gnd 0.010975f
C2379 commonsourceibias.n388 gnd 0.012728f
C2380 commonsourceibias.n389 gnd 0.068768f
C2381 commonsourceibias.n390 gnd 0.012651f
C2382 commonsourceibias.n391 gnd 0.009225f
C2383 commonsourceibias.n392 gnd 0.009225f
C2384 commonsourceibias.n393 gnd 0.009225f
C2385 commonsourceibias.n394 gnd 0.012496f
C2386 commonsourceibias.n395 gnd 0.068768f
C2387 commonsourceibias.n396 gnd 0.012578f
C2388 commonsourceibias.n397 gnd 0.01137f
C2389 commonsourceibias.n398 gnd 0.009225f
C2390 commonsourceibias.n399 gnd 0.009225f
C2391 commonsourceibias.n400 gnd 0.009358f
C2392 commonsourceibias.n401 gnd 0.009674f
C2393 commonsourceibias.n402 gnd 0.082281f
C2394 commonsourceibias.n403 gnd 0.053268f
C2395 commonsourceibias.n404 gnd 0.01231f
C2396 commonsourceibias.t107 gnd 0.17235f
C2397 commonsourceibias.n405 gnd 0.068768f
C2398 commonsourceibias.n406 gnd 0.009225f
C2399 commonsourceibias.t50 gnd 0.17235f
C2400 commonsourceibias.n407 gnd 0.007462f
C2401 commonsourceibias.n408 gnd 0.009225f
C2402 commonsourceibias.t114 gnd 0.17235f
C2403 commonsourceibias.n409 gnd 0.008906f
C2404 commonsourceibias.n410 gnd 0.009225f
C2405 commonsourceibias.t49 gnd 0.17235f
C2406 commonsourceibias.n411 gnd 0.007451f
C2407 commonsourceibias.n412 gnd 0.009225f
C2408 commonsourceibias.t74 gnd 0.17235f
C2409 commonsourceibias.t105 gnd 0.17235f
C2410 commonsourceibias.n413 gnd 0.068768f
C2411 commonsourceibias.n414 gnd 0.009225f
C2412 commonsourceibias.t55 gnd 0.17235f
C2413 commonsourceibias.n415 gnd 0.068768f
C2414 commonsourceibias.n416 gnd 0.009225f
C2415 commonsourceibias.t75 gnd 0.17235f
C2416 commonsourceibias.n417 gnd 0.068768f
C2417 commonsourceibias.n418 gnd 0.046441f
C2418 commonsourceibias.t61 gnd 0.17235f
C2419 commonsourceibias.t52 gnd 0.194477f
C2420 commonsourceibias.n419 gnd 0.079804f
C2421 commonsourceibias.n420 gnd 0.082619f
C2422 commonsourceibias.n421 gnd 0.01137f
C2423 commonsourceibias.n422 gnd 0.012578f
C2424 commonsourceibias.n423 gnd 0.009225f
C2425 commonsourceibias.n424 gnd 0.009225f
C2426 commonsourceibias.n425 gnd 0.012496f
C2427 commonsourceibias.n426 gnd 0.007462f
C2428 commonsourceibias.n427 gnd 0.012651f
C2429 commonsourceibias.n428 gnd 0.009225f
C2430 commonsourceibias.n429 gnd 0.009225f
C2431 commonsourceibias.n430 gnd 0.012728f
C2432 commonsourceibias.n431 gnd 0.010975f
C2433 commonsourceibias.n432 gnd 0.008906f
C2434 commonsourceibias.n433 gnd 0.009225f
C2435 commonsourceibias.n434 gnd 0.009225f
C2436 commonsourceibias.n435 gnd 0.011283f
C2437 commonsourceibias.n436 gnd 0.012665f
C2438 commonsourceibias.n437 gnd 0.068768f
C2439 commonsourceibias.n438 gnd 0.01258f
C2440 commonsourceibias.n439 gnd 0.009225f
C2441 commonsourceibias.n440 gnd 0.009225f
C2442 commonsourceibias.n441 gnd 0.009225f
C2443 commonsourceibias.n442 gnd 0.01258f
C2444 commonsourceibias.n443 gnd 0.068768f
C2445 commonsourceibias.n444 gnd 0.012665f
C2446 commonsourceibias.t106 gnd 0.17235f
C2447 commonsourceibias.n445 gnd 0.068768f
C2448 commonsourceibias.n446 gnd 0.011283f
C2449 commonsourceibias.n447 gnd 0.009225f
C2450 commonsourceibias.n448 gnd 0.009225f
C2451 commonsourceibias.n449 gnd 0.009225f
C2452 commonsourceibias.n450 gnd 0.010975f
C2453 commonsourceibias.n451 gnd 0.012728f
C2454 commonsourceibias.n452 gnd 0.068768f
C2455 commonsourceibias.n453 gnd 0.012651f
C2456 commonsourceibias.n454 gnd 0.009225f
C2457 commonsourceibias.n455 gnd 0.009225f
C2458 commonsourceibias.n456 gnd 0.009225f
C2459 commonsourceibias.n457 gnd 0.012496f
C2460 commonsourceibias.n458 gnd 0.068768f
C2461 commonsourceibias.n459 gnd 0.012578f
C2462 commonsourceibias.n460 gnd 0.01137f
C2463 commonsourceibias.n461 gnd 0.009225f
C2464 commonsourceibias.n462 gnd 0.009225f
C2465 commonsourceibias.n463 gnd 0.009358f
C2466 commonsourceibias.n464 gnd 0.009674f
C2467 commonsourceibias.t112 gnd 0.186396f
C2468 commonsourceibias.n465 gnd 0.082281f
C2469 commonsourceibias.n466 gnd 0.028001f
C2470 commonsourceibias.n467 gnd 0.147196f
C2471 commonsourceibias.n468 gnd 0.01231f
C2472 commonsourceibias.t81 gnd 0.17235f
C2473 commonsourceibias.n469 gnd 0.068768f
C2474 commonsourceibias.n470 gnd 0.009225f
C2475 commonsourceibias.t91 gnd 0.17235f
C2476 commonsourceibias.n471 gnd 0.007462f
C2477 commonsourceibias.n472 gnd 0.009225f
C2478 commonsourceibias.t100 gnd 0.17235f
C2479 commonsourceibias.n473 gnd 0.008906f
C2480 commonsourceibias.n474 gnd 0.009225f
C2481 commonsourceibias.t85 gnd 0.17235f
C2482 commonsourceibias.n475 gnd 0.007451f
C2483 commonsourceibias.n476 gnd 0.009225f
C2484 commonsourceibias.t82 gnd 0.17235f
C2485 commonsourceibias.t62 gnd 0.17235f
C2486 commonsourceibias.n477 gnd 0.068768f
C2487 commonsourceibias.n478 gnd 0.009225f
C2488 commonsourceibias.t53 gnd 0.17235f
C2489 commonsourceibias.n479 gnd 0.068768f
C2490 commonsourceibias.n480 gnd 0.009225f
C2491 commonsourceibias.t78 gnd 0.17235f
C2492 commonsourceibias.n481 gnd 0.068768f
C2493 commonsourceibias.n482 gnd 0.046441f
C2494 commonsourceibias.t97 gnd 0.17235f
C2495 commonsourceibias.t113 gnd 0.194477f
C2496 commonsourceibias.n483 gnd 0.079804f
C2497 commonsourceibias.n484 gnd 0.082619f
C2498 commonsourceibias.n485 gnd 0.01137f
C2499 commonsourceibias.n486 gnd 0.012578f
C2500 commonsourceibias.n487 gnd 0.009225f
C2501 commonsourceibias.n488 gnd 0.009225f
C2502 commonsourceibias.n489 gnd 0.012496f
C2503 commonsourceibias.n490 gnd 0.007462f
C2504 commonsourceibias.n491 gnd 0.012651f
C2505 commonsourceibias.n492 gnd 0.009225f
C2506 commonsourceibias.n493 gnd 0.009225f
C2507 commonsourceibias.n494 gnd 0.012728f
C2508 commonsourceibias.n495 gnd 0.010975f
C2509 commonsourceibias.n496 gnd 0.008906f
C2510 commonsourceibias.n497 gnd 0.009225f
C2511 commonsourceibias.n498 gnd 0.009225f
C2512 commonsourceibias.n499 gnd 0.011283f
C2513 commonsourceibias.n500 gnd 0.012665f
C2514 commonsourceibias.n501 gnd 0.068768f
C2515 commonsourceibias.n502 gnd 0.01258f
C2516 commonsourceibias.n503 gnd 0.009225f
C2517 commonsourceibias.n504 gnd 0.009225f
C2518 commonsourceibias.n505 gnd 0.009225f
C2519 commonsourceibias.n506 gnd 0.01258f
C2520 commonsourceibias.n507 gnd 0.068768f
C2521 commonsourceibias.n508 gnd 0.012665f
C2522 commonsourceibias.t76 gnd 0.17235f
C2523 commonsourceibias.n509 gnd 0.068768f
C2524 commonsourceibias.n510 gnd 0.011283f
C2525 commonsourceibias.n511 gnd 0.009225f
C2526 commonsourceibias.n512 gnd 0.009225f
C2527 commonsourceibias.n513 gnd 0.009225f
C2528 commonsourceibias.n514 gnd 0.010975f
C2529 commonsourceibias.n515 gnd 0.012728f
C2530 commonsourceibias.n516 gnd 0.068768f
C2531 commonsourceibias.n517 gnd 0.012651f
C2532 commonsourceibias.n518 gnd 0.009225f
C2533 commonsourceibias.n519 gnd 0.009225f
C2534 commonsourceibias.n520 gnd 0.009225f
C2535 commonsourceibias.n521 gnd 0.012496f
C2536 commonsourceibias.n522 gnd 0.068768f
C2537 commonsourceibias.n523 gnd 0.012578f
C2538 commonsourceibias.n524 gnd 0.01137f
C2539 commonsourceibias.n525 gnd 0.009225f
C2540 commonsourceibias.n526 gnd 0.009225f
C2541 commonsourceibias.n527 gnd 0.009358f
C2542 commonsourceibias.n528 gnd 0.009674f
C2543 commonsourceibias.t63 gnd 0.186396f
C2544 commonsourceibias.n529 gnd 0.082281f
C2545 commonsourceibias.n530 gnd 0.028001f
C2546 commonsourceibias.n531 gnd 0.194447f
C2547 commonsourceibias.n532 gnd 4.93338f
C2548 vdd.t267 gnd 0.037058f
C2549 vdd.t247 gnd 0.037058f
C2550 vdd.n0 gnd 0.29228f
C2551 vdd.t226 gnd 0.037058f
C2552 vdd.t263 gnd 0.037058f
C2553 vdd.n1 gnd 0.291797f
C2554 vdd.n2 gnd 0.269092f
C2555 vdd.t244 gnd 0.037058f
C2556 vdd.t274 gnd 0.037058f
C2557 vdd.n3 gnd 0.291797f
C2558 vdd.n4 gnd 0.13609f
C2559 vdd.t272 gnd 0.037058f
C2560 vdd.t252 gnd 0.037058f
C2561 vdd.n5 gnd 0.291797f
C2562 vdd.n6 gnd 0.127695f
C2563 vdd.t278 gnd 0.037058f
C2564 vdd.t242 gnd 0.037058f
C2565 vdd.n7 gnd 0.29228f
C2566 vdd.t250 gnd 0.037058f
C2567 vdd.t270 gnd 0.037058f
C2568 vdd.n8 gnd 0.291797f
C2569 vdd.n9 gnd 0.269093f
C2570 vdd.t259 gnd 0.037058f
C2571 vdd.t230 gnd 0.037058f
C2572 vdd.n10 gnd 0.291797f
C2573 vdd.n11 gnd 0.13609f
C2574 vdd.t239 gnd 0.037058f
C2575 vdd.t257 gnd 0.037058f
C2576 vdd.n12 gnd 0.291797f
C2577 vdd.n13 gnd 0.127695f
C2578 vdd.n14 gnd 0.090278f
C2579 vdd.t26 gnd 0.020588f
C2580 vdd.t99 gnd 0.020588f
C2581 vdd.n15 gnd 0.1895f
C2582 vdd.t98 gnd 0.020588f
C2583 vdd.t95 gnd 0.020588f
C2584 vdd.n16 gnd 0.188945f
C2585 vdd.n17 gnd 0.328824f
C2586 vdd.t101 gnd 0.020588f
C2587 vdd.t83 gnd 0.020588f
C2588 vdd.n18 gnd 0.188945f
C2589 vdd.n19 gnd 0.136039f
C2590 vdd.t4 gnd 0.020588f
C2591 vdd.t96 gnd 0.020588f
C2592 vdd.n20 gnd 0.1895f
C2593 vdd.t27 gnd 0.020588f
C2594 vdd.t100 gnd 0.020588f
C2595 vdd.n21 gnd 0.188945f
C2596 vdd.n22 gnd 0.328824f
C2597 vdd.t84 gnd 0.020588f
C2598 vdd.t28 gnd 0.020588f
C2599 vdd.n23 gnd 0.188945f
C2600 vdd.n24 gnd 0.136039f
C2601 vdd.t94 gnd 0.020588f
C2602 vdd.t5 gnd 0.020588f
C2603 vdd.n25 gnd 0.188945f
C2604 vdd.t82 gnd 0.020588f
C2605 vdd.t97 gnd 0.020588f
C2606 vdd.n26 gnd 0.188945f
C2607 vdd.n27 gnd 20.7697f
C2608 vdd.n28 gnd 8.3397f
C2609 vdd.n29 gnd 0.005615f
C2610 vdd.n30 gnd 0.005211f
C2611 vdd.n31 gnd 0.002882f
C2612 vdd.n32 gnd 0.006618f
C2613 vdd.n33 gnd 0.0028f
C2614 vdd.n34 gnd 0.002965f
C2615 vdd.n35 gnd 0.005211f
C2616 vdd.n36 gnd 0.0028f
C2617 vdd.n37 gnd 0.006618f
C2618 vdd.n38 gnd 0.002965f
C2619 vdd.n39 gnd 0.005211f
C2620 vdd.n40 gnd 0.0028f
C2621 vdd.n41 gnd 0.004963f
C2622 vdd.n42 gnd 0.004978f
C2623 vdd.t38 gnd 0.014218f
C2624 vdd.n43 gnd 0.031635f
C2625 vdd.n44 gnd 0.164637f
C2626 vdd.n45 gnd 0.0028f
C2627 vdd.n46 gnd 0.002965f
C2628 vdd.n47 gnd 0.006618f
C2629 vdd.n48 gnd 0.006618f
C2630 vdd.n49 gnd 0.002965f
C2631 vdd.n50 gnd 0.0028f
C2632 vdd.n51 gnd 0.005211f
C2633 vdd.n52 gnd 0.005211f
C2634 vdd.n53 gnd 0.0028f
C2635 vdd.n54 gnd 0.002965f
C2636 vdd.n55 gnd 0.006618f
C2637 vdd.n56 gnd 0.006618f
C2638 vdd.n57 gnd 0.002965f
C2639 vdd.n58 gnd 0.0028f
C2640 vdd.n59 gnd 0.005211f
C2641 vdd.n60 gnd 0.005211f
C2642 vdd.n61 gnd 0.0028f
C2643 vdd.n62 gnd 0.002965f
C2644 vdd.n63 gnd 0.006618f
C2645 vdd.n64 gnd 0.006618f
C2646 vdd.n65 gnd 0.015646f
C2647 vdd.n66 gnd 0.002882f
C2648 vdd.n67 gnd 0.0028f
C2649 vdd.n68 gnd 0.013467f
C2650 vdd.n69 gnd 0.009402f
C2651 vdd.t21 gnd 0.03294f
C2652 vdd.t121 gnd 0.03294f
C2653 vdd.n70 gnd 0.226387f
C2654 vdd.n71 gnd 0.178019f
C2655 vdd.t6 gnd 0.03294f
C2656 vdd.t78 gnd 0.03294f
C2657 vdd.n72 gnd 0.226387f
C2658 vdd.n73 gnd 0.14366f
C2659 vdd.t289 gnd 0.03294f
C2660 vdd.t45 gnd 0.03294f
C2661 vdd.n74 gnd 0.226387f
C2662 vdd.n75 gnd 0.14366f
C2663 vdd.t290 gnd 0.03294f
C2664 vdd.t120 gnd 0.03294f
C2665 vdd.n76 gnd 0.226387f
C2666 vdd.n77 gnd 0.14366f
C2667 vdd.t91 gnd 0.03294f
C2668 vdd.t306 gnd 0.03294f
C2669 vdd.n78 gnd 0.226387f
C2670 vdd.n79 gnd 0.14366f
C2671 vdd.t34 gnd 0.03294f
C2672 vdd.t14 gnd 0.03294f
C2673 vdd.n80 gnd 0.226387f
C2674 vdd.n81 gnd 0.14366f
C2675 vdd.t141 gnd 0.03294f
C2676 vdd.t80 gnd 0.03294f
C2677 vdd.n82 gnd 0.226387f
C2678 vdd.n83 gnd 0.14366f
C2679 vdd.t75 gnd 0.03294f
C2680 vdd.t126 gnd 0.03294f
C2681 vdd.n84 gnd 0.226387f
C2682 vdd.n85 gnd 0.14366f
C2683 vdd.t131 gnd 0.03294f
C2684 vdd.t118 gnd 0.03294f
C2685 vdd.n86 gnd 0.226387f
C2686 vdd.n87 gnd 0.14366f
C2687 vdd.n88 gnd 0.005615f
C2688 vdd.n89 gnd 0.005211f
C2689 vdd.n90 gnd 0.002882f
C2690 vdd.n91 gnd 0.006618f
C2691 vdd.n92 gnd 0.0028f
C2692 vdd.n93 gnd 0.002965f
C2693 vdd.n94 gnd 0.005211f
C2694 vdd.n95 gnd 0.0028f
C2695 vdd.n96 gnd 0.006618f
C2696 vdd.n97 gnd 0.002965f
C2697 vdd.n98 gnd 0.005211f
C2698 vdd.n99 gnd 0.0028f
C2699 vdd.n100 gnd 0.004963f
C2700 vdd.n101 gnd 0.004978f
C2701 vdd.t144 gnd 0.014218f
C2702 vdd.n102 gnd 0.031635f
C2703 vdd.n103 gnd 0.164637f
C2704 vdd.n104 gnd 0.0028f
C2705 vdd.n105 gnd 0.002965f
C2706 vdd.n106 gnd 0.006618f
C2707 vdd.n107 gnd 0.006618f
C2708 vdd.n108 gnd 0.002965f
C2709 vdd.n109 gnd 0.0028f
C2710 vdd.n110 gnd 0.005211f
C2711 vdd.n111 gnd 0.005211f
C2712 vdd.n112 gnd 0.0028f
C2713 vdd.n113 gnd 0.002965f
C2714 vdd.n114 gnd 0.006618f
C2715 vdd.n115 gnd 0.006618f
C2716 vdd.n116 gnd 0.002965f
C2717 vdd.n117 gnd 0.0028f
C2718 vdd.n118 gnd 0.005211f
C2719 vdd.n119 gnd 0.005211f
C2720 vdd.n120 gnd 0.0028f
C2721 vdd.n121 gnd 0.002965f
C2722 vdd.n122 gnd 0.006618f
C2723 vdd.n123 gnd 0.006618f
C2724 vdd.n124 gnd 0.015646f
C2725 vdd.n125 gnd 0.002882f
C2726 vdd.n126 gnd 0.0028f
C2727 vdd.n127 gnd 0.013467f
C2728 vdd.n128 gnd 0.009107f
C2729 vdd.n129 gnd 0.106884f
C2730 vdd.n130 gnd 0.005615f
C2731 vdd.n131 gnd 0.005211f
C2732 vdd.n132 gnd 0.002882f
C2733 vdd.n133 gnd 0.006618f
C2734 vdd.n134 gnd 0.0028f
C2735 vdd.n135 gnd 0.002965f
C2736 vdd.n136 gnd 0.005211f
C2737 vdd.n137 gnd 0.0028f
C2738 vdd.n138 gnd 0.006618f
C2739 vdd.n139 gnd 0.002965f
C2740 vdd.n140 gnd 0.005211f
C2741 vdd.n141 gnd 0.0028f
C2742 vdd.n142 gnd 0.004963f
C2743 vdd.n143 gnd 0.004978f
C2744 vdd.t145 gnd 0.014218f
C2745 vdd.n144 gnd 0.031635f
C2746 vdd.n145 gnd 0.164637f
C2747 vdd.n146 gnd 0.0028f
C2748 vdd.n147 gnd 0.002965f
C2749 vdd.n148 gnd 0.006618f
C2750 vdd.n149 gnd 0.006618f
C2751 vdd.n150 gnd 0.002965f
C2752 vdd.n151 gnd 0.0028f
C2753 vdd.n152 gnd 0.005211f
C2754 vdd.n153 gnd 0.005211f
C2755 vdd.n154 gnd 0.0028f
C2756 vdd.n155 gnd 0.002965f
C2757 vdd.n156 gnd 0.006618f
C2758 vdd.n157 gnd 0.006618f
C2759 vdd.n158 gnd 0.002965f
C2760 vdd.n159 gnd 0.0028f
C2761 vdd.n160 gnd 0.005211f
C2762 vdd.n161 gnd 0.005211f
C2763 vdd.n162 gnd 0.0028f
C2764 vdd.n163 gnd 0.002965f
C2765 vdd.n164 gnd 0.006618f
C2766 vdd.n165 gnd 0.006618f
C2767 vdd.n166 gnd 0.015646f
C2768 vdd.n167 gnd 0.002882f
C2769 vdd.n168 gnd 0.0028f
C2770 vdd.n169 gnd 0.013467f
C2771 vdd.n170 gnd 0.009402f
C2772 vdd.t114 gnd 0.03294f
C2773 vdd.t30 gnd 0.03294f
C2774 vdd.n171 gnd 0.226387f
C2775 vdd.n172 gnd 0.178019f
C2776 vdd.t294 gnd 0.03294f
C2777 vdd.t122 gnd 0.03294f
C2778 vdd.n173 gnd 0.226387f
C2779 vdd.n174 gnd 0.14366f
C2780 vdd.t104 gnd 0.03294f
C2781 vdd.t40 gnd 0.03294f
C2782 vdd.n175 gnd 0.226387f
C2783 vdd.n176 gnd 0.14366f
C2784 vdd.t307 gnd 0.03294f
C2785 vdd.t283 gnd 0.03294f
C2786 vdd.n177 gnd 0.226387f
C2787 vdd.n178 gnd 0.14366f
C2788 vdd.t73 gnd 0.03294f
C2789 vdd.t111 gnd 0.03294f
C2790 vdd.n179 gnd 0.226387f
C2791 vdd.n180 gnd 0.14366f
C2792 vdd.t297 gnd 0.03294f
C2793 vdd.t22 gnd 0.03294f
C2794 vdd.n181 gnd 0.226387f
C2795 vdd.n182 gnd 0.14366f
C2796 vdd.t76 gnd 0.03294f
C2797 vdd.t146 gnd 0.03294f
C2798 vdd.n183 gnd 0.226387f
C2799 vdd.n184 gnd 0.14366f
C2800 vdd.t32 gnd 0.03294f
C2801 vdd.t62 gnd 0.03294f
C2802 vdd.n185 gnd 0.226387f
C2803 vdd.n186 gnd 0.14366f
C2804 vdd.t1 gnd 0.03294f
C2805 vdd.t138 gnd 0.03294f
C2806 vdd.n187 gnd 0.226387f
C2807 vdd.n188 gnd 0.14366f
C2808 vdd.n189 gnd 0.005615f
C2809 vdd.n190 gnd 0.005211f
C2810 vdd.n191 gnd 0.002882f
C2811 vdd.n192 gnd 0.006618f
C2812 vdd.n193 gnd 0.0028f
C2813 vdd.n194 gnd 0.002965f
C2814 vdd.n195 gnd 0.005211f
C2815 vdd.n196 gnd 0.0028f
C2816 vdd.n197 gnd 0.006618f
C2817 vdd.n198 gnd 0.002965f
C2818 vdd.n199 gnd 0.005211f
C2819 vdd.n200 gnd 0.0028f
C2820 vdd.n201 gnd 0.004963f
C2821 vdd.n202 gnd 0.004978f
C2822 vdd.t137 gnd 0.014218f
C2823 vdd.n203 gnd 0.031635f
C2824 vdd.n204 gnd 0.164637f
C2825 vdd.n205 gnd 0.0028f
C2826 vdd.n206 gnd 0.002965f
C2827 vdd.n207 gnd 0.006618f
C2828 vdd.n208 gnd 0.006618f
C2829 vdd.n209 gnd 0.002965f
C2830 vdd.n210 gnd 0.0028f
C2831 vdd.n211 gnd 0.005211f
C2832 vdd.n212 gnd 0.005211f
C2833 vdd.n213 gnd 0.0028f
C2834 vdd.n214 gnd 0.002965f
C2835 vdd.n215 gnd 0.006618f
C2836 vdd.n216 gnd 0.006618f
C2837 vdd.n217 gnd 0.002965f
C2838 vdd.n218 gnd 0.0028f
C2839 vdd.n219 gnd 0.005211f
C2840 vdd.n220 gnd 0.005211f
C2841 vdd.n221 gnd 0.0028f
C2842 vdd.n222 gnd 0.002965f
C2843 vdd.n223 gnd 0.006618f
C2844 vdd.n224 gnd 0.006618f
C2845 vdd.n225 gnd 0.015646f
C2846 vdd.n226 gnd 0.002882f
C2847 vdd.n227 gnd 0.0028f
C2848 vdd.n228 gnd 0.013467f
C2849 vdd.n229 gnd 0.009107f
C2850 vdd.n230 gnd 0.063585f
C2851 vdd.n231 gnd 0.229114f
C2852 vdd.n232 gnd 0.005615f
C2853 vdd.n233 gnd 0.005211f
C2854 vdd.n234 gnd 0.002882f
C2855 vdd.n235 gnd 0.006618f
C2856 vdd.n236 gnd 0.0028f
C2857 vdd.n237 gnd 0.002965f
C2858 vdd.n238 gnd 0.005211f
C2859 vdd.n239 gnd 0.0028f
C2860 vdd.n240 gnd 0.006618f
C2861 vdd.n241 gnd 0.002965f
C2862 vdd.n242 gnd 0.005211f
C2863 vdd.n243 gnd 0.0028f
C2864 vdd.n244 gnd 0.004963f
C2865 vdd.n245 gnd 0.004978f
C2866 vdd.t93 gnd 0.014218f
C2867 vdd.n246 gnd 0.031635f
C2868 vdd.n247 gnd 0.164637f
C2869 vdd.n248 gnd 0.0028f
C2870 vdd.n249 gnd 0.002965f
C2871 vdd.n250 gnd 0.006618f
C2872 vdd.n251 gnd 0.006618f
C2873 vdd.n252 gnd 0.002965f
C2874 vdd.n253 gnd 0.0028f
C2875 vdd.n254 gnd 0.005211f
C2876 vdd.n255 gnd 0.005211f
C2877 vdd.n256 gnd 0.0028f
C2878 vdd.n257 gnd 0.002965f
C2879 vdd.n258 gnd 0.006618f
C2880 vdd.n259 gnd 0.006618f
C2881 vdd.n260 gnd 0.002965f
C2882 vdd.n261 gnd 0.0028f
C2883 vdd.n262 gnd 0.005211f
C2884 vdd.n263 gnd 0.005211f
C2885 vdd.n264 gnd 0.0028f
C2886 vdd.n265 gnd 0.002965f
C2887 vdd.n266 gnd 0.006618f
C2888 vdd.n267 gnd 0.006618f
C2889 vdd.n268 gnd 0.015646f
C2890 vdd.n269 gnd 0.002882f
C2891 vdd.n270 gnd 0.0028f
C2892 vdd.n271 gnd 0.013467f
C2893 vdd.n272 gnd 0.009402f
C2894 vdd.t81 gnd 0.03294f
C2895 vdd.t63 gnd 0.03294f
C2896 vdd.n273 gnd 0.226387f
C2897 vdd.n274 gnd 0.178019f
C2898 vdd.t3 gnd 0.03294f
C2899 vdd.t18 gnd 0.03294f
C2900 vdd.n275 gnd 0.226387f
C2901 vdd.n276 gnd 0.14366f
C2902 vdd.t288 gnd 0.03294f
C2903 vdd.t55 gnd 0.03294f
C2904 vdd.n277 gnd 0.226387f
C2905 vdd.n278 gnd 0.14366f
C2906 vdd.t280 gnd 0.03294f
C2907 vdd.t134 gnd 0.03294f
C2908 vdd.n279 gnd 0.226387f
C2909 vdd.n280 gnd 0.14366f
C2910 vdd.t142 gnd 0.03294f
C2911 vdd.t47 gnd 0.03294f
C2912 vdd.n281 gnd 0.226387f
C2913 vdd.n282 gnd 0.14366f
C2914 vdd.t102 gnd 0.03294f
C2915 vdd.t133 gnd 0.03294f
C2916 vdd.n283 gnd 0.226387f
C2917 vdd.n284 gnd 0.14366f
C2918 vdd.t44 gnd 0.03294f
C2919 vdd.t92 gnd 0.03294f
C2920 vdd.n285 gnd 0.226387f
C2921 vdd.n286 gnd 0.14366f
C2922 vdd.t51 gnd 0.03294f
C2923 vdd.t140 gnd 0.03294f
C2924 vdd.n287 gnd 0.226387f
C2925 vdd.n288 gnd 0.14366f
C2926 vdd.t19 gnd 0.03294f
C2927 vdd.t299 gnd 0.03294f
C2928 vdd.n289 gnd 0.226387f
C2929 vdd.n290 gnd 0.14366f
C2930 vdd.n291 gnd 0.005615f
C2931 vdd.n292 gnd 0.005211f
C2932 vdd.n293 gnd 0.002882f
C2933 vdd.n294 gnd 0.006618f
C2934 vdd.n295 gnd 0.0028f
C2935 vdd.n296 gnd 0.002965f
C2936 vdd.n297 gnd 0.005211f
C2937 vdd.n298 gnd 0.0028f
C2938 vdd.n299 gnd 0.006618f
C2939 vdd.n300 gnd 0.002965f
C2940 vdd.n301 gnd 0.005211f
C2941 vdd.n302 gnd 0.0028f
C2942 vdd.n303 gnd 0.004963f
C2943 vdd.n304 gnd 0.004978f
C2944 vdd.t71 gnd 0.014218f
C2945 vdd.n305 gnd 0.031635f
C2946 vdd.n306 gnd 0.164637f
C2947 vdd.n307 gnd 0.0028f
C2948 vdd.n308 gnd 0.002965f
C2949 vdd.n309 gnd 0.006618f
C2950 vdd.n310 gnd 0.006618f
C2951 vdd.n311 gnd 0.002965f
C2952 vdd.n312 gnd 0.0028f
C2953 vdd.n313 gnd 0.005211f
C2954 vdd.n314 gnd 0.005211f
C2955 vdd.n315 gnd 0.0028f
C2956 vdd.n316 gnd 0.002965f
C2957 vdd.n317 gnd 0.006618f
C2958 vdd.n318 gnd 0.006618f
C2959 vdd.n319 gnd 0.002965f
C2960 vdd.n320 gnd 0.0028f
C2961 vdd.n321 gnd 0.005211f
C2962 vdd.n322 gnd 0.005211f
C2963 vdd.n323 gnd 0.0028f
C2964 vdd.n324 gnd 0.002965f
C2965 vdd.n325 gnd 0.006618f
C2966 vdd.n326 gnd 0.006618f
C2967 vdd.n327 gnd 0.015646f
C2968 vdd.n328 gnd 0.002882f
C2969 vdd.n329 gnd 0.0028f
C2970 vdd.n330 gnd 0.013467f
C2971 vdd.n331 gnd 0.009107f
C2972 vdd.n332 gnd 0.063585f
C2973 vdd.n333 gnd 0.262286f
C2974 vdd.n334 gnd 0.007863f
C2975 vdd.n335 gnd 0.010231f
C2976 vdd.n336 gnd 0.008235f
C2977 vdd.n337 gnd 0.008235f
C2978 vdd.n338 gnd 0.010231f
C2979 vdd.n339 gnd 0.010231f
C2980 vdd.n340 gnd 0.747604f
C2981 vdd.n341 gnd 0.010231f
C2982 vdd.n342 gnd 0.010231f
C2983 vdd.n343 gnd 0.010231f
C2984 vdd.n344 gnd 0.810339f
C2985 vdd.n345 gnd 0.010231f
C2986 vdd.n346 gnd 0.010231f
C2987 vdd.n347 gnd 0.010231f
C2988 vdd.n348 gnd 0.010231f
C2989 vdd.n349 gnd 0.008235f
C2990 vdd.n350 gnd 0.010231f
C2991 vdd.t13 gnd 0.5228f
C2992 vdd.n351 gnd 0.010231f
C2993 vdd.n352 gnd 0.010231f
C2994 vdd.n353 gnd 0.010231f
C2995 vdd.t79 gnd 0.5228f
C2996 vdd.n354 gnd 0.010231f
C2997 vdd.n355 gnd 0.010231f
C2998 vdd.n356 gnd 0.010231f
C2999 vdd.n357 gnd 0.010231f
C3000 vdd.n358 gnd 0.010231f
C3001 vdd.n359 gnd 0.008235f
C3002 vdd.n360 gnd 0.010231f
C3003 vdd.n361 gnd 0.590764f
C3004 vdd.n362 gnd 0.010231f
C3005 vdd.n363 gnd 0.010231f
C3006 vdd.n364 gnd 0.010231f
C3007 vdd.t61 gnd 0.5228f
C3008 vdd.n365 gnd 0.010231f
C3009 vdd.n366 gnd 0.010231f
C3010 vdd.n367 gnd 0.010231f
C3011 vdd.n368 gnd 0.010231f
C3012 vdd.n369 gnd 0.010231f
C3013 vdd.n370 gnd 0.008235f
C3014 vdd.n371 gnd 0.010231f
C3015 vdd.t0 gnd 0.5228f
C3016 vdd.n372 gnd 0.010231f
C3017 vdd.n373 gnd 0.010231f
C3018 vdd.n374 gnd 0.010231f
C3019 vdd.n375 gnd 0.611676f
C3020 vdd.n376 gnd 0.010231f
C3021 vdd.n377 gnd 0.010231f
C3022 vdd.n378 gnd 0.010231f
C3023 vdd.n379 gnd 0.010231f
C3024 vdd.n380 gnd 0.010231f
C3025 vdd.n381 gnd 0.008235f
C3026 vdd.n382 gnd 0.010231f
C3027 vdd.t70 gnd 0.5228f
C3028 vdd.n383 gnd 0.010231f
C3029 vdd.n384 gnd 0.010231f
C3030 vdd.n385 gnd 0.010231f
C3031 vdd.n386 gnd 0.528028f
C3032 vdd.n387 gnd 0.010231f
C3033 vdd.n388 gnd 0.010231f
C3034 vdd.n389 gnd 0.010231f
C3035 vdd.n390 gnd 0.010231f
C3036 vdd.n391 gnd 0.024751f
C3037 vdd.n392 gnd 0.025281f
C3038 vdd.t160 gnd 0.5228f
C3039 vdd.n393 gnd 0.024751f
C3040 vdd.n425 gnd 0.010231f
C3041 vdd.t188 gnd 0.125873f
C3042 vdd.t187 gnd 0.134524f
C3043 vdd.t186 gnd 0.164388f
C3044 vdd.n426 gnd 0.210723f
C3045 vdd.n427 gnd 0.177869f
C3046 vdd.n428 gnd 0.013505f
C3047 vdd.n429 gnd 0.010231f
C3048 vdd.n430 gnd 0.008235f
C3049 vdd.n431 gnd 0.010231f
C3050 vdd.n432 gnd 0.008235f
C3051 vdd.n433 gnd 0.010231f
C3052 vdd.n434 gnd 0.008235f
C3053 vdd.n435 gnd 0.010231f
C3054 vdd.n436 gnd 0.008235f
C3055 vdd.n437 gnd 0.010231f
C3056 vdd.n438 gnd 0.008235f
C3057 vdd.n439 gnd 0.010231f
C3058 vdd.t162 gnd 0.125873f
C3059 vdd.t161 gnd 0.134524f
C3060 vdd.t159 gnd 0.164388f
C3061 vdd.n440 gnd 0.210723f
C3062 vdd.n441 gnd 0.177869f
C3063 vdd.n442 gnd 0.008235f
C3064 vdd.n443 gnd 0.010231f
C3065 vdd.n444 gnd 0.008235f
C3066 vdd.n445 gnd 0.010231f
C3067 vdd.n446 gnd 0.008235f
C3068 vdd.n447 gnd 0.010231f
C3069 vdd.n448 gnd 0.008235f
C3070 vdd.n449 gnd 0.010231f
C3071 vdd.n450 gnd 0.008235f
C3072 vdd.n451 gnd 0.010231f
C3073 vdd.t168 gnd 0.125873f
C3074 vdd.t167 gnd 0.134524f
C3075 vdd.t166 gnd 0.164388f
C3076 vdd.n452 gnd 0.210723f
C3077 vdd.n453 gnd 0.177869f
C3078 vdd.n454 gnd 0.017623f
C3079 vdd.n455 gnd 0.010231f
C3080 vdd.n456 gnd 0.008235f
C3081 vdd.n457 gnd 0.010231f
C3082 vdd.n458 gnd 0.008235f
C3083 vdd.n459 gnd 0.010231f
C3084 vdd.n460 gnd 0.008235f
C3085 vdd.n461 gnd 0.010231f
C3086 vdd.n462 gnd 0.008235f
C3087 vdd.n463 gnd 0.010231f
C3088 vdd.n464 gnd 0.025281f
C3089 vdd.n465 gnd 0.006835f
C3090 vdd.n466 gnd 0.008235f
C3091 vdd.n467 gnd 0.010231f
C3092 vdd.n468 gnd 0.010231f
C3093 vdd.n469 gnd 0.008235f
C3094 vdd.n470 gnd 0.010231f
C3095 vdd.n471 gnd 0.010231f
C3096 vdd.n472 gnd 0.010231f
C3097 vdd.n473 gnd 0.010231f
C3098 vdd.n474 gnd 0.010231f
C3099 vdd.n475 gnd 0.008235f
C3100 vdd.n476 gnd 0.008235f
C3101 vdd.n477 gnd 0.010231f
C3102 vdd.n478 gnd 0.010231f
C3103 vdd.n479 gnd 0.008235f
C3104 vdd.n480 gnd 0.010231f
C3105 vdd.n481 gnd 0.010231f
C3106 vdd.n482 gnd 0.010231f
C3107 vdd.n483 gnd 0.010231f
C3108 vdd.n484 gnd 0.010231f
C3109 vdd.n485 gnd 0.008235f
C3110 vdd.n486 gnd 0.008235f
C3111 vdd.n487 gnd 0.010231f
C3112 vdd.n488 gnd 0.010231f
C3113 vdd.n489 gnd 0.008235f
C3114 vdd.n490 gnd 0.010231f
C3115 vdd.n491 gnd 0.010231f
C3116 vdd.n492 gnd 0.010231f
C3117 vdd.n493 gnd 0.010231f
C3118 vdd.n494 gnd 0.010231f
C3119 vdd.n495 gnd 0.008235f
C3120 vdd.n496 gnd 0.008235f
C3121 vdd.n497 gnd 0.010231f
C3122 vdd.n498 gnd 0.010231f
C3123 vdd.n499 gnd 0.008235f
C3124 vdd.n500 gnd 0.010231f
C3125 vdd.n501 gnd 0.010231f
C3126 vdd.n502 gnd 0.010231f
C3127 vdd.n503 gnd 0.010231f
C3128 vdd.n504 gnd 0.010231f
C3129 vdd.n505 gnd 0.008235f
C3130 vdd.n506 gnd 0.008235f
C3131 vdd.n507 gnd 0.010231f
C3132 vdd.n508 gnd 0.010231f
C3133 vdd.n509 gnd 0.006876f
C3134 vdd.n510 gnd 0.010231f
C3135 vdd.n511 gnd 0.010231f
C3136 vdd.n512 gnd 0.010231f
C3137 vdd.n513 gnd 0.010231f
C3138 vdd.n514 gnd 0.010231f
C3139 vdd.n515 gnd 0.006876f
C3140 vdd.n516 gnd 0.008235f
C3141 vdd.n517 gnd 0.010231f
C3142 vdd.n518 gnd 0.010231f
C3143 vdd.n519 gnd 0.008235f
C3144 vdd.n520 gnd 0.010231f
C3145 vdd.n521 gnd 0.010231f
C3146 vdd.n522 gnd 0.010231f
C3147 vdd.n523 gnd 0.010231f
C3148 vdd.n524 gnd 0.010231f
C3149 vdd.n525 gnd 0.008235f
C3150 vdd.n526 gnd 0.008235f
C3151 vdd.n527 gnd 0.010231f
C3152 vdd.n528 gnd 0.010231f
C3153 vdd.n529 gnd 0.008235f
C3154 vdd.n530 gnd 0.010231f
C3155 vdd.n531 gnd 0.010231f
C3156 vdd.n532 gnd 0.010231f
C3157 vdd.n533 gnd 0.010231f
C3158 vdd.n534 gnd 0.010231f
C3159 vdd.n535 gnd 0.008235f
C3160 vdd.n536 gnd 0.008235f
C3161 vdd.n537 gnd 0.010231f
C3162 vdd.n538 gnd 0.010231f
C3163 vdd.n539 gnd 0.008235f
C3164 vdd.n540 gnd 0.010231f
C3165 vdd.n541 gnd 0.010231f
C3166 vdd.n542 gnd 0.010231f
C3167 vdd.n543 gnd 0.010231f
C3168 vdd.n544 gnd 0.010231f
C3169 vdd.n545 gnd 0.008235f
C3170 vdd.n546 gnd 0.008235f
C3171 vdd.n547 gnd 0.010231f
C3172 vdd.n548 gnd 0.010231f
C3173 vdd.n549 gnd 0.008235f
C3174 vdd.n550 gnd 0.010231f
C3175 vdd.n551 gnd 0.010231f
C3176 vdd.n552 gnd 0.010231f
C3177 vdd.n553 gnd 0.010231f
C3178 vdd.n554 gnd 0.010231f
C3179 vdd.n555 gnd 0.008235f
C3180 vdd.n556 gnd 0.008235f
C3181 vdd.n557 gnd 0.010231f
C3182 vdd.n558 gnd 0.010231f
C3183 vdd.n559 gnd 0.008235f
C3184 vdd.n560 gnd 0.010231f
C3185 vdd.n561 gnd 0.010231f
C3186 vdd.n562 gnd 0.010231f
C3187 vdd.n563 gnd 0.010231f
C3188 vdd.n564 gnd 0.010231f
C3189 vdd.n565 gnd 0.0056f
C3190 vdd.n566 gnd 0.017623f
C3191 vdd.n567 gnd 0.010231f
C3192 vdd.n568 gnd 0.010231f
C3193 vdd.n569 gnd 0.008153f
C3194 vdd.n570 gnd 0.010231f
C3195 vdd.n571 gnd 0.010231f
C3196 vdd.n572 gnd 0.010231f
C3197 vdd.n573 gnd 0.010231f
C3198 vdd.n574 gnd 0.010231f
C3199 vdd.n575 gnd 0.008235f
C3200 vdd.n576 gnd 0.008235f
C3201 vdd.n577 gnd 0.010231f
C3202 vdd.n578 gnd 0.010231f
C3203 vdd.n579 gnd 0.008235f
C3204 vdd.n580 gnd 0.010231f
C3205 vdd.n581 gnd 0.010231f
C3206 vdd.n582 gnd 0.010231f
C3207 vdd.n583 gnd 0.010231f
C3208 vdd.n584 gnd 0.010231f
C3209 vdd.n585 gnd 0.008235f
C3210 vdd.n586 gnd 0.008235f
C3211 vdd.n587 gnd 0.010231f
C3212 vdd.n588 gnd 0.010231f
C3213 vdd.n589 gnd 0.008235f
C3214 vdd.n590 gnd 0.010231f
C3215 vdd.n591 gnd 0.010231f
C3216 vdd.n592 gnd 0.010231f
C3217 vdd.n593 gnd 0.010231f
C3218 vdd.n594 gnd 0.010231f
C3219 vdd.n595 gnd 0.008235f
C3220 vdd.n596 gnd 0.008235f
C3221 vdd.n597 gnd 0.010231f
C3222 vdd.n598 gnd 0.010231f
C3223 vdd.n599 gnd 0.008235f
C3224 vdd.n600 gnd 0.010231f
C3225 vdd.n601 gnd 0.010231f
C3226 vdd.n602 gnd 0.010231f
C3227 vdd.n603 gnd 0.010231f
C3228 vdd.n604 gnd 0.010231f
C3229 vdd.n605 gnd 0.008235f
C3230 vdd.n606 gnd 0.008235f
C3231 vdd.n607 gnd 0.010231f
C3232 vdd.n608 gnd 0.010231f
C3233 vdd.n609 gnd 0.008235f
C3234 vdd.n610 gnd 0.010231f
C3235 vdd.n611 gnd 0.010231f
C3236 vdd.n612 gnd 0.010231f
C3237 vdd.n613 gnd 0.010231f
C3238 vdd.n614 gnd 0.010231f
C3239 vdd.n615 gnd 0.008235f
C3240 vdd.n616 gnd 0.010231f
C3241 vdd.n617 gnd 0.008235f
C3242 vdd.n618 gnd 0.004323f
C3243 vdd.n619 gnd 0.010231f
C3244 vdd.n620 gnd 0.010231f
C3245 vdd.n621 gnd 0.008235f
C3246 vdd.n622 gnd 0.010231f
C3247 vdd.n623 gnd 0.008235f
C3248 vdd.n624 gnd 0.010231f
C3249 vdd.n625 gnd 0.008235f
C3250 vdd.n626 gnd 0.010231f
C3251 vdd.n627 gnd 0.008235f
C3252 vdd.n628 gnd 0.010231f
C3253 vdd.n629 gnd 0.008235f
C3254 vdd.n630 gnd 0.010231f
C3255 vdd.n631 gnd 0.008235f
C3256 vdd.n632 gnd 0.010231f
C3257 vdd.n633 gnd 0.569852f
C3258 vdd.t72 gnd 0.5228f
C3259 vdd.n634 gnd 0.010231f
C3260 vdd.n635 gnd 0.008235f
C3261 vdd.n636 gnd 0.010231f
C3262 vdd.n637 gnd 0.008235f
C3263 vdd.n638 gnd 0.010231f
C3264 vdd.t279 gnd 0.5228f
C3265 vdd.n639 gnd 0.010231f
C3266 vdd.n640 gnd 0.008235f
C3267 vdd.n641 gnd 0.010231f
C3268 vdd.n642 gnd 0.008235f
C3269 vdd.n643 gnd 0.010231f
C3270 vdd.t39 gnd 0.5228f
C3271 vdd.n644 gnd 0.6535f
C3272 vdd.n645 gnd 0.010231f
C3273 vdd.n646 gnd 0.008235f
C3274 vdd.n647 gnd 0.010231f
C3275 vdd.n648 gnd 0.008235f
C3276 vdd.n649 gnd 0.010231f
C3277 vdd.t103 gnd 0.5228f
C3278 vdd.n650 gnd 0.010231f
C3279 vdd.n651 gnd 0.008235f
C3280 vdd.n652 gnd 0.010231f
C3281 vdd.n653 gnd 0.008235f
C3282 vdd.n654 gnd 0.010231f
C3283 vdd.n655 gnd 0.726692f
C3284 vdd.n656 gnd 0.867847f
C3285 vdd.t17 gnd 0.5228f
C3286 vdd.n657 gnd 0.010231f
C3287 vdd.n658 gnd 0.008235f
C3288 vdd.n659 gnd 0.010231f
C3289 vdd.n660 gnd 0.008235f
C3290 vdd.n661 gnd 0.010231f
C3291 vdd.n662 gnd 0.54894f
C3292 vdd.n663 gnd 0.010231f
C3293 vdd.n664 gnd 0.008235f
C3294 vdd.n665 gnd 0.010231f
C3295 vdd.n666 gnd 0.008235f
C3296 vdd.n667 gnd 0.010231f
C3297 vdd.t20 gnd 0.5228f
C3298 vdd.t29 gnd 0.5228f
C3299 vdd.n668 gnd 0.010231f
C3300 vdd.n669 gnd 0.008235f
C3301 vdd.n670 gnd 0.010231f
C3302 vdd.n671 gnd 0.008235f
C3303 vdd.n672 gnd 0.010231f
C3304 vdd.t37 gnd 0.5228f
C3305 vdd.n673 gnd 0.010231f
C3306 vdd.n674 gnd 0.008235f
C3307 vdd.n675 gnd 0.010231f
C3308 vdd.n676 gnd 0.008235f
C3309 vdd.n677 gnd 0.010231f
C3310 vdd.n678 gnd 1.0456f
C3311 vdd.n679 gnd 0.852163f
C3312 vdd.n680 gnd 0.010231f
C3313 vdd.n681 gnd 0.008235f
C3314 vdd.n682 gnd 0.024751f
C3315 vdd.n683 gnd 0.006835f
C3316 vdd.n684 gnd 0.024751f
C3317 vdd.t173 gnd 0.5228f
C3318 vdd.n685 gnd 0.024751f
C3319 vdd.n686 gnd 0.006835f
C3320 vdd.n687 gnd 0.008799f
C3321 vdd.t174 gnd 0.125873f
C3322 vdd.t175 gnd 0.134524f
C3323 vdd.t172 gnd 0.164388f
C3324 vdd.n688 gnd 0.210723f
C3325 vdd.n689 gnd 0.177045f
C3326 vdd.n690 gnd 0.012682f
C3327 vdd.n691 gnd 0.010231f
C3328 vdd.n692 gnd 12.3485f
C3329 vdd.n723 gnd 1.4377f
C3330 vdd.n724 gnd 0.010231f
C3331 vdd.n725 gnd 0.010231f
C3332 vdd.n726 gnd 0.025281f
C3333 vdd.n727 gnd 0.008799f
C3334 vdd.n728 gnd 0.010231f
C3335 vdd.n729 gnd 0.008235f
C3336 vdd.n730 gnd 0.006548f
C3337 vdd.n731 gnd 0.042961f
C3338 vdd.n732 gnd 0.008235f
C3339 vdd.n733 gnd 0.010231f
C3340 vdd.n734 gnd 0.010231f
C3341 vdd.n735 gnd 0.010231f
C3342 vdd.n736 gnd 0.010231f
C3343 vdd.n737 gnd 0.010231f
C3344 vdd.n738 gnd 0.010231f
C3345 vdd.n739 gnd 0.010231f
C3346 vdd.n740 gnd 0.010231f
C3347 vdd.n741 gnd 0.010231f
C3348 vdd.n742 gnd 0.010231f
C3349 vdd.n743 gnd 0.010231f
C3350 vdd.n744 gnd 0.010231f
C3351 vdd.n745 gnd 0.010231f
C3352 vdd.n746 gnd 0.010231f
C3353 vdd.n747 gnd 0.006876f
C3354 vdd.n748 gnd 0.010231f
C3355 vdd.n749 gnd 0.010231f
C3356 vdd.n750 gnd 0.010231f
C3357 vdd.n751 gnd 0.010231f
C3358 vdd.n752 gnd 0.010231f
C3359 vdd.n753 gnd 0.010231f
C3360 vdd.n754 gnd 0.010231f
C3361 vdd.n755 gnd 0.010231f
C3362 vdd.n756 gnd 0.010231f
C3363 vdd.n757 gnd 0.010231f
C3364 vdd.n758 gnd 0.010231f
C3365 vdd.n759 gnd 0.010231f
C3366 vdd.n760 gnd 0.010231f
C3367 vdd.n761 gnd 0.010231f
C3368 vdd.n762 gnd 0.010231f
C3369 vdd.n763 gnd 0.010231f
C3370 vdd.n764 gnd 0.010231f
C3371 vdd.n765 gnd 0.010231f
C3372 vdd.n766 gnd 0.010231f
C3373 vdd.n767 gnd 0.008153f
C3374 vdd.t184 gnd 0.125873f
C3375 vdd.t185 gnd 0.134524f
C3376 vdd.t183 gnd 0.164388f
C3377 vdd.n768 gnd 0.210723f
C3378 vdd.n769 gnd 0.177045f
C3379 vdd.n770 gnd 0.010231f
C3380 vdd.n771 gnd 0.010231f
C3381 vdd.n772 gnd 0.010231f
C3382 vdd.n773 gnd 0.010231f
C3383 vdd.n774 gnd 0.010231f
C3384 vdd.n775 gnd 0.010231f
C3385 vdd.n776 gnd 0.010231f
C3386 vdd.n777 gnd 0.010231f
C3387 vdd.n778 gnd 0.010231f
C3388 vdd.n779 gnd 0.010231f
C3389 vdd.n780 gnd 0.010231f
C3390 vdd.n781 gnd 0.010231f
C3391 vdd.n782 gnd 0.010231f
C3392 vdd.n783 gnd 0.006548f
C3393 vdd.n785 gnd 0.006957f
C3394 vdd.n786 gnd 0.006957f
C3395 vdd.n787 gnd 0.006957f
C3396 vdd.n788 gnd 0.006957f
C3397 vdd.n789 gnd 0.006957f
C3398 vdd.n790 gnd 0.006957f
C3399 vdd.n792 gnd 0.006957f
C3400 vdd.n793 gnd 0.006957f
C3401 vdd.n795 gnd 0.006957f
C3402 vdd.n796 gnd 0.005065f
C3403 vdd.n798 gnd 0.006957f
C3404 vdd.t150 gnd 0.281145f
C3405 vdd.t149 gnd 0.287787f
C3406 vdd.t147 gnd 0.183542f
C3407 vdd.n799 gnd 0.099195f
C3408 vdd.n800 gnd 0.056266f
C3409 vdd.n801 gnd 0.009943f
C3410 vdd.n802 gnd 0.015797f
C3411 vdd.n804 gnd 0.006957f
C3412 vdd.n805 gnd 0.711008f
C3413 vdd.n806 gnd 0.014897f
C3414 vdd.n807 gnd 0.014897f
C3415 vdd.n808 gnd 0.006957f
C3416 vdd.n809 gnd 0.015797f
C3417 vdd.n810 gnd 0.006957f
C3418 vdd.n811 gnd 0.006957f
C3419 vdd.n812 gnd 0.006957f
C3420 vdd.n813 gnd 0.006957f
C3421 vdd.n814 gnd 0.006957f
C3422 vdd.n816 gnd 0.006957f
C3423 vdd.n817 gnd 0.006957f
C3424 vdd.n819 gnd 0.006957f
C3425 vdd.n820 gnd 0.006957f
C3426 vdd.n822 gnd 0.006957f
C3427 vdd.n823 gnd 0.006957f
C3428 vdd.n825 gnd 0.006957f
C3429 vdd.n826 gnd 0.006957f
C3430 vdd.n828 gnd 0.006957f
C3431 vdd.n829 gnd 0.006957f
C3432 vdd.n831 gnd 0.006957f
C3433 vdd.t171 gnd 0.281145f
C3434 vdd.t170 gnd 0.287787f
C3435 vdd.t169 gnd 0.183542f
C3436 vdd.n832 gnd 0.099195f
C3437 vdd.n833 gnd 0.056266f
C3438 vdd.n834 gnd 0.006957f
C3439 vdd.n836 gnd 0.006957f
C3440 vdd.n837 gnd 0.006957f
C3441 vdd.t148 gnd 0.355504f
C3442 vdd.n838 gnd 0.006957f
C3443 vdd.n839 gnd 0.006957f
C3444 vdd.n840 gnd 0.006957f
C3445 vdd.n841 gnd 0.006957f
C3446 vdd.n842 gnd 0.006957f
C3447 vdd.n843 gnd 0.711008f
C3448 vdd.n844 gnd 0.006957f
C3449 vdd.n845 gnd 0.006957f
C3450 vdd.n846 gnd 0.559396f
C3451 vdd.n847 gnd 0.006957f
C3452 vdd.n848 gnd 0.006957f
C3453 vdd.n849 gnd 0.006957f
C3454 vdd.n850 gnd 0.006957f
C3455 vdd.n851 gnd 0.711008f
C3456 vdd.n852 gnd 0.006957f
C3457 vdd.n853 gnd 0.006957f
C3458 vdd.n854 gnd 0.006957f
C3459 vdd.n855 gnd 0.006957f
C3460 vdd.n856 gnd 0.006957f
C3461 vdd.t237 gnd 0.355504f
C3462 vdd.n857 gnd 0.006957f
C3463 vdd.n858 gnd 0.006957f
C3464 vdd.n859 gnd 0.006957f
C3465 vdd.n860 gnd 0.006957f
C3466 vdd.n861 gnd 0.006957f
C3467 vdd.t254 gnd 0.355504f
C3468 vdd.n862 gnd 0.006957f
C3469 vdd.n863 gnd 0.006957f
C3470 vdd.n864 gnd 0.684868f
C3471 vdd.n865 gnd 0.006957f
C3472 vdd.n866 gnd 0.006957f
C3473 vdd.n867 gnd 0.006957f
C3474 vdd.t253 gnd 0.355504f
C3475 vdd.n868 gnd 0.006957f
C3476 vdd.n869 gnd 0.006957f
C3477 vdd.n870 gnd 0.528028f
C3478 vdd.n871 gnd 0.006957f
C3479 vdd.n872 gnd 0.006957f
C3480 vdd.n873 gnd 0.006957f
C3481 vdd.n874 gnd 0.49666f
C3482 vdd.n875 gnd 0.006957f
C3483 vdd.n876 gnd 0.006957f
C3484 vdd.n877 gnd 0.371188f
C3485 vdd.n878 gnd 0.006957f
C3486 vdd.n879 gnd 0.006957f
C3487 vdd.n880 gnd 0.006957f
C3488 vdd.n881 gnd 0.6535f
C3489 vdd.n882 gnd 0.006957f
C3490 vdd.n883 gnd 0.006957f
C3491 vdd.t260 gnd 0.355504f
C3492 vdd.n884 gnd 0.006957f
C3493 vdd.n885 gnd 0.006957f
C3494 vdd.n886 gnd 0.006957f
C3495 vdd.n887 gnd 0.711008f
C3496 vdd.n888 gnd 0.006957f
C3497 vdd.n889 gnd 0.006957f
C3498 vdd.t261 gnd 0.355504f
C3499 vdd.n890 gnd 0.006957f
C3500 vdd.n891 gnd 0.006957f
C3501 vdd.n892 gnd 0.006957f
C3502 vdd.t231 gnd 0.355504f
C3503 vdd.n893 gnd 0.006957f
C3504 vdd.n894 gnd 0.006957f
C3505 vdd.n895 gnd 0.006957f
C3506 vdd.t178 gnd 0.287787f
C3507 vdd.t176 gnd 0.183542f
C3508 vdd.t179 gnd 0.287787f
C3509 vdd.n896 gnd 0.161748f
C3510 vdd.n897 gnd 0.020155f
C3511 vdd.n898 gnd 0.006957f
C3512 vdd.t177 gnd 0.256172f
C3513 vdd.n899 gnd 0.006957f
C3514 vdd.n900 gnd 0.006957f
C3515 vdd.n901 gnd 0.611676f
C3516 vdd.n902 gnd 0.006957f
C3517 vdd.n903 gnd 0.006957f
C3518 vdd.n904 gnd 0.006957f
C3519 vdd.n905 gnd 0.413012f
C3520 vdd.n906 gnd 0.006957f
C3521 vdd.n907 gnd 0.006957f
C3522 vdd.t232 gnd 0.146384f
C3523 vdd.n908 gnd 0.454836f
C3524 vdd.n909 gnd 0.006957f
C3525 vdd.n910 gnd 0.006957f
C3526 vdd.n911 gnd 0.006957f
C3527 vdd.n912 gnd 0.569852f
C3528 vdd.n913 gnd 0.006957f
C3529 vdd.n914 gnd 0.006957f
C3530 vdd.t245 gnd 0.355504f
C3531 vdd.n915 gnd 0.006957f
C3532 vdd.n916 gnd 0.006957f
C3533 vdd.n917 gnd 0.006957f
C3534 vdd.t241 gnd 0.355504f
C3535 vdd.n918 gnd 0.006957f
C3536 vdd.n919 gnd 0.006957f
C3537 vdd.t264 gnd 0.355504f
C3538 vdd.n920 gnd 0.006957f
C3539 vdd.n921 gnd 0.006957f
C3540 vdd.n922 gnd 0.006957f
C3541 vdd.t223 gnd 0.240488f
C3542 vdd.n923 gnd 0.006957f
C3543 vdd.n924 gnd 0.006957f
C3544 vdd.n925 gnd 0.62736f
C3545 vdd.n926 gnd 0.006957f
C3546 vdd.n927 gnd 0.006957f
C3547 vdd.n928 gnd 0.006957f
C3548 vdd.t265 gnd 0.355504f
C3549 vdd.n929 gnd 0.006957f
C3550 vdd.n930 gnd 0.006957f
C3551 vdd.t277 gnd 0.33982f
C3552 vdd.n931 gnd 0.47052f
C3553 vdd.n932 gnd 0.006957f
C3554 vdd.n933 gnd 0.006957f
C3555 vdd.n934 gnd 0.006957f
C3556 vdd.t227 gnd 0.355504f
C3557 vdd.n935 gnd 0.006957f
C3558 vdd.n936 gnd 0.006957f
C3559 vdd.t269 gnd 0.355504f
C3560 vdd.n937 gnd 0.006957f
C3561 vdd.n938 gnd 0.006957f
C3562 vdd.n939 gnd 0.006957f
C3563 vdd.n940 gnd 0.711008f
C3564 vdd.n941 gnd 0.006957f
C3565 vdd.n942 gnd 0.006957f
C3566 vdd.t249 gnd 0.355504f
C3567 vdd.n943 gnd 0.006957f
C3568 vdd.n944 gnd 0.006957f
C3569 vdd.n945 gnd 0.006957f
C3570 vdd.n946 gnd 0.491432f
C3571 vdd.n947 gnd 0.006957f
C3572 vdd.n948 gnd 0.006957f
C3573 vdd.n949 gnd 0.006957f
C3574 vdd.n950 gnd 0.006957f
C3575 vdd.n951 gnd 0.006957f
C3576 vdd.t200 gnd 0.355504f
C3577 vdd.n952 gnd 0.006957f
C3578 vdd.n953 gnd 0.006957f
C3579 vdd.t229 gnd 0.355504f
C3580 vdd.n954 gnd 0.006957f
C3581 vdd.n955 gnd 0.014897f
C3582 vdd.n956 gnd 0.014897f
C3583 vdd.n957 gnd 0.805111f
C3584 vdd.n958 gnd 0.006957f
C3585 vdd.n959 gnd 0.006957f
C3586 vdd.t258 gnd 0.355504f
C3587 vdd.n960 gnd 0.014897f
C3588 vdd.n961 gnd 0.006957f
C3589 vdd.n962 gnd 0.006957f
C3590 vdd.t271 gnd 0.606448f
C3591 vdd.n980 gnd 0.015797f
C3592 vdd.n998 gnd 0.014897f
C3593 vdd.n999 gnd 0.006957f
C3594 vdd.n1000 gnd 0.014897f
C3595 vdd.t216 gnd 0.281145f
C3596 vdd.t215 gnd 0.287787f
C3597 vdd.t214 gnd 0.183542f
C3598 vdd.n1001 gnd 0.099195f
C3599 vdd.n1002 gnd 0.056266f
C3600 vdd.n1003 gnd 0.015797f
C3601 vdd.n1004 gnd 0.006957f
C3602 vdd.n1005 gnd 0.41824f
C3603 vdd.n1006 gnd 0.014897f
C3604 vdd.n1007 gnd 0.006957f
C3605 vdd.n1008 gnd 0.015797f
C3606 vdd.n1009 gnd 0.006957f
C3607 vdd.t195 gnd 0.281145f
C3608 vdd.t194 gnd 0.287787f
C3609 vdd.t192 gnd 0.183542f
C3610 vdd.n1010 gnd 0.099195f
C3611 vdd.n1011 gnd 0.056266f
C3612 vdd.n1012 gnd 0.009943f
C3613 vdd.n1013 gnd 0.006957f
C3614 vdd.n1014 gnd 0.006957f
C3615 vdd.t193 gnd 0.355504f
C3616 vdd.n1015 gnd 0.006957f
C3617 vdd.t273 gnd 0.355504f
C3618 vdd.n1016 gnd 0.006957f
C3619 vdd.n1017 gnd 0.006957f
C3620 vdd.n1018 gnd 0.006957f
C3621 vdd.n1019 gnd 0.006957f
C3622 vdd.n1020 gnd 0.006957f
C3623 vdd.n1021 gnd 0.711008f
C3624 vdd.n1022 gnd 0.006957f
C3625 vdd.n1023 gnd 0.006957f
C3626 vdd.t243 gnd 0.355504f
C3627 vdd.n1024 gnd 0.006957f
C3628 vdd.n1025 gnd 0.006957f
C3629 vdd.n1026 gnd 0.006957f
C3630 vdd.n1027 gnd 0.006957f
C3631 vdd.n1028 gnd 0.512344f
C3632 vdd.n1029 gnd 0.006957f
C3633 vdd.n1030 gnd 0.006957f
C3634 vdd.n1031 gnd 0.006957f
C3635 vdd.n1032 gnd 0.006957f
C3636 vdd.n1033 gnd 0.006957f
C3637 vdd.t224 gnd 0.355504f
C3638 vdd.n1034 gnd 0.006957f
C3639 vdd.n1035 gnd 0.006957f
C3640 vdd.t262 gnd 0.355504f
C3641 vdd.n1036 gnd 0.006957f
C3642 vdd.n1037 gnd 0.006957f
C3643 vdd.n1038 gnd 0.006957f
C3644 vdd.t248 gnd 0.355504f
C3645 vdd.n1039 gnd 0.006957f
C3646 vdd.n1040 gnd 0.006957f
C3647 vdd.t225 gnd 0.355504f
C3648 vdd.n1041 gnd 0.006957f
C3649 vdd.n1042 gnd 0.006957f
C3650 vdd.n1043 gnd 0.006957f
C3651 vdd.t246 gnd 0.33982f
C3652 vdd.n1044 gnd 0.006957f
C3653 vdd.n1045 gnd 0.006957f
C3654 vdd.n1046 gnd 0.528028f
C3655 vdd.n1047 gnd 0.006957f
C3656 vdd.n1048 gnd 0.006957f
C3657 vdd.n1049 gnd 0.006957f
C3658 vdd.t266 gnd 0.355504f
C3659 vdd.n1050 gnd 0.006957f
C3660 vdd.n1051 gnd 0.006957f
C3661 vdd.t234 gnd 0.240488f
C3662 vdd.n1052 gnd 0.371188f
C3663 vdd.n1053 gnd 0.006957f
C3664 vdd.n1054 gnd 0.006957f
C3665 vdd.n1055 gnd 0.006957f
C3666 vdd.n1056 gnd 0.6535f
C3667 vdd.n1057 gnd 0.006957f
C3668 vdd.n1058 gnd 0.006957f
C3669 vdd.t275 gnd 0.355504f
C3670 vdd.n1059 gnd 0.006957f
C3671 vdd.n1060 gnd 0.006957f
C3672 vdd.n1061 gnd 0.006957f
C3673 vdd.n1062 gnd 0.711008f
C3674 vdd.n1063 gnd 0.006957f
C3675 vdd.n1064 gnd 0.006957f
C3676 vdd.t240 gnd 0.355504f
C3677 vdd.n1065 gnd 0.006957f
C3678 vdd.n1066 gnd 0.006957f
C3679 vdd.n1067 gnd 0.006957f
C3680 vdd.t233 gnd 0.146384f
C3681 vdd.n1068 gnd 0.006957f
C3682 vdd.n1069 gnd 0.006957f
C3683 vdd.n1070 gnd 0.006957f
C3684 vdd.t205 gnd 0.287787f
C3685 vdd.t203 gnd 0.183542f
C3686 vdd.t206 gnd 0.287787f
C3687 vdd.n1071 gnd 0.161748f
C3688 vdd.n1072 gnd 0.006957f
C3689 vdd.n1073 gnd 0.006957f
C3690 vdd.t255 gnd 0.355504f
C3691 vdd.n1074 gnd 0.006957f
C3692 vdd.n1075 gnd 0.006957f
C3693 vdd.t204 gnd 0.256172f
C3694 vdd.n1076 gnd 0.564624f
C3695 vdd.n1077 gnd 0.006957f
C3696 vdd.n1078 gnd 0.006957f
C3697 vdd.n1079 gnd 0.006957f
C3698 vdd.n1080 gnd 0.413012f
C3699 vdd.n1081 gnd 0.006957f
C3700 vdd.n1082 gnd 0.006957f
C3701 vdd.n1083 gnd 0.454836f
C3702 vdd.n1084 gnd 0.006957f
C3703 vdd.n1085 gnd 0.006957f
C3704 vdd.n1086 gnd 0.006957f
C3705 vdd.n1087 gnd 0.569852f
C3706 vdd.n1088 gnd 0.006957f
C3707 vdd.n1089 gnd 0.006957f
C3708 vdd.t235 gnd 0.355504f
C3709 vdd.n1090 gnd 0.006957f
C3710 vdd.n1091 gnd 0.006957f
C3711 vdd.n1092 gnd 0.006957f
C3712 vdd.n1093 gnd 0.711008f
C3713 vdd.n1094 gnd 0.006957f
C3714 vdd.n1095 gnd 0.006957f
C3715 vdd.t236 gnd 0.355504f
C3716 vdd.n1096 gnd 0.006957f
C3717 vdd.n1097 gnd 0.006957f
C3718 vdd.n1098 gnd 0.006957f
C3719 vdd.t276 gnd 0.355504f
C3720 vdd.n1099 gnd 0.006957f
C3721 vdd.n1100 gnd 0.006957f
C3722 vdd.n1101 gnd 0.006957f
C3723 vdd.n1102 gnd 0.006957f
C3724 vdd.n1103 gnd 0.006957f
C3725 vdd.t268 gnd 0.355504f
C3726 vdd.n1104 gnd 0.006957f
C3727 vdd.n1105 gnd 0.006957f
C3728 vdd.n1106 gnd 0.695324f
C3729 vdd.n1107 gnd 0.006957f
C3730 vdd.n1108 gnd 0.006957f
C3731 vdd.n1109 gnd 0.006957f
C3732 vdd.t228 gnd 0.355504f
C3733 vdd.n1110 gnd 0.006957f
C3734 vdd.n1111 gnd 0.006957f
C3735 vdd.n1112 gnd 0.538484f
C3736 vdd.n1113 gnd 0.006957f
C3737 vdd.n1114 gnd 0.006957f
C3738 vdd.n1115 gnd 0.006957f
C3739 vdd.n1116 gnd 0.711008f
C3740 vdd.n1117 gnd 0.006957f
C3741 vdd.n1118 gnd 0.006957f
C3742 vdd.n1119 gnd 0.381644f
C3743 vdd.n1120 gnd 0.006957f
C3744 vdd.n1121 gnd 0.006957f
C3745 vdd.n1122 gnd 0.006957f
C3746 vdd.n1123 gnd 0.711008f
C3747 vdd.n1124 gnd 0.006957f
C3748 vdd.n1125 gnd 0.006957f
C3749 vdd.n1126 gnd 0.006957f
C3750 vdd.n1127 gnd 0.006957f
C3751 vdd.n1128 gnd 0.006957f
C3752 vdd.t152 gnd 0.355504f
C3753 vdd.n1129 gnd 0.006957f
C3754 vdd.n1130 gnd 0.006957f
C3755 vdd.n1131 gnd 0.006957f
C3756 vdd.n1132 gnd 0.014897f
C3757 vdd.n1133 gnd 0.014897f
C3758 vdd.n1134 gnd 0.961951f
C3759 vdd.n1135 gnd 0.006957f
C3760 vdd.n1136 gnd 0.006957f
C3761 vdd.n1137 gnd 0.507116f
C3762 vdd.n1138 gnd 0.014897f
C3763 vdd.n1139 gnd 0.006957f
C3764 vdd.n1140 gnd 0.006957f
C3765 vdd.n1141 gnd 12.7668f
C3766 vdd.n1175 gnd 0.015797f
C3767 vdd.n1176 gnd 0.006957f
C3768 vdd.n1177 gnd 0.006957f
C3769 vdd.n1178 gnd 0.006548f
C3770 vdd.n1181 gnd 0.025281f
C3771 vdd.n1182 gnd 0.006835f
C3772 vdd.n1183 gnd 0.008235f
C3773 vdd.n1185 gnd 0.010231f
C3774 vdd.n1186 gnd 0.010231f
C3775 vdd.n1187 gnd 0.008235f
C3776 vdd.n1189 gnd 0.010231f
C3777 vdd.n1190 gnd 0.010231f
C3778 vdd.n1191 gnd 0.010231f
C3779 vdd.n1192 gnd 0.010231f
C3780 vdd.n1193 gnd 0.010231f
C3781 vdd.n1194 gnd 0.008235f
C3782 vdd.n1196 gnd 0.010231f
C3783 vdd.n1197 gnd 0.010231f
C3784 vdd.n1198 gnd 0.010231f
C3785 vdd.n1199 gnd 0.010231f
C3786 vdd.n1200 gnd 0.010231f
C3787 vdd.n1201 gnd 0.008235f
C3788 vdd.n1203 gnd 0.010231f
C3789 vdd.n1204 gnd 0.010231f
C3790 vdd.n1205 gnd 0.010231f
C3791 vdd.n1206 gnd 0.010231f
C3792 vdd.n1207 gnd 0.006876f
C3793 vdd.t165 gnd 0.125873f
C3794 vdd.t164 gnd 0.134524f
C3795 vdd.t163 gnd 0.164388f
C3796 vdd.n1208 gnd 0.210723f
C3797 vdd.n1209 gnd 0.177045f
C3798 vdd.n1211 gnd 0.010231f
C3799 vdd.n1212 gnd 0.010231f
C3800 vdd.n1213 gnd 0.008235f
C3801 vdd.n1214 gnd 0.010231f
C3802 vdd.n1216 gnd 0.010231f
C3803 vdd.n1217 gnd 0.010231f
C3804 vdd.n1218 gnd 0.010231f
C3805 vdd.n1219 gnd 0.010231f
C3806 vdd.n1220 gnd 0.008235f
C3807 vdd.n1222 gnd 0.010231f
C3808 vdd.n1223 gnd 0.010231f
C3809 vdd.n1224 gnd 0.010231f
C3810 vdd.n1225 gnd 0.010231f
C3811 vdd.n1226 gnd 0.010231f
C3812 vdd.n1227 gnd 0.008235f
C3813 vdd.n1229 gnd 0.010231f
C3814 vdd.n1230 gnd 0.010231f
C3815 vdd.n1231 gnd 0.010231f
C3816 vdd.n1232 gnd 0.010231f
C3817 vdd.n1233 gnd 0.010231f
C3818 vdd.n1234 gnd 0.008235f
C3819 vdd.n1236 gnd 0.010231f
C3820 vdd.n1237 gnd 0.010231f
C3821 vdd.n1238 gnd 0.010231f
C3822 vdd.n1239 gnd 0.010231f
C3823 vdd.n1240 gnd 0.010231f
C3824 vdd.n1241 gnd 0.008235f
C3825 vdd.n1243 gnd 0.010231f
C3826 vdd.n1244 gnd 0.010231f
C3827 vdd.n1245 gnd 0.010231f
C3828 vdd.n1246 gnd 0.010231f
C3829 vdd.n1247 gnd 0.008153f
C3830 vdd.t158 gnd 0.125873f
C3831 vdd.t157 gnd 0.134524f
C3832 vdd.t155 gnd 0.164388f
C3833 vdd.n1248 gnd 0.210723f
C3834 vdd.n1249 gnd 0.177045f
C3835 vdd.n1251 gnd 0.010231f
C3836 vdd.n1252 gnd 0.010231f
C3837 vdd.n1253 gnd 0.008235f
C3838 vdd.n1254 gnd 0.010231f
C3839 vdd.n1256 gnd 0.010231f
C3840 vdd.n1257 gnd 0.010231f
C3841 vdd.n1258 gnd 0.010231f
C3842 vdd.n1259 gnd 0.010231f
C3843 vdd.n1260 gnd 0.008235f
C3844 vdd.n1262 gnd 0.010231f
C3845 vdd.n1263 gnd 0.010231f
C3846 vdd.n1264 gnd 0.010231f
C3847 vdd.n1265 gnd 0.010231f
C3848 vdd.n1266 gnd 0.010231f
C3849 vdd.n1267 gnd 0.008235f
C3850 vdd.n1269 gnd 0.010231f
C3851 vdd.n1270 gnd 0.010231f
C3852 vdd.n1271 gnd 0.010231f
C3853 vdd.n1272 gnd 0.010231f
C3854 vdd.n1273 gnd 0.010231f
C3855 vdd.n1274 gnd 0.008235f
C3856 vdd.n1276 gnd 0.010231f
C3857 vdd.n1277 gnd 0.010231f
C3858 vdd.n1278 gnd 0.006548f
C3859 vdd.n1279 gnd 0.008235f
C3860 vdd.n1280 gnd 0.015797f
C3861 vdd.n1281 gnd 0.015797f
C3862 vdd.n1282 gnd 0.006957f
C3863 vdd.n1283 gnd 0.006957f
C3864 vdd.n1284 gnd 0.006957f
C3865 vdd.n1285 gnd 0.006957f
C3866 vdd.n1286 gnd 0.006957f
C3867 vdd.n1287 gnd 0.006957f
C3868 vdd.n1288 gnd 0.006957f
C3869 vdd.n1289 gnd 0.006957f
C3870 vdd.n1290 gnd 0.006957f
C3871 vdd.n1291 gnd 0.006957f
C3872 vdd.n1292 gnd 0.006957f
C3873 vdd.n1293 gnd 0.006957f
C3874 vdd.n1294 gnd 0.006957f
C3875 vdd.n1295 gnd 0.006957f
C3876 vdd.n1296 gnd 0.006957f
C3877 vdd.n1297 gnd 0.006957f
C3878 vdd.n1298 gnd 0.006957f
C3879 vdd.n1299 gnd 0.006957f
C3880 vdd.n1300 gnd 0.006957f
C3881 vdd.n1301 gnd 0.006957f
C3882 vdd.n1302 gnd 0.006957f
C3883 vdd.n1303 gnd 0.006957f
C3884 vdd.n1304 gnd 0.006957f
C3885 vdd.n1305 gnd 0.006957f
C3886 vdd.n1306 gnd 0.006957f
C3887 vdd.n1307 gnd 0.006957f
C3888 vdd.n1308 gnd 0.006957f
C3889 vdd.n1309 gnd 0.006957f
C3890 vdd.n1310 gnd 0.006957f
C3891 vdd.n1311 gnd 0.006957f
C3892 vdd.n1312 gnd 0.006957f
C3893 vdd.n1313 gnd 0.006957f
C3894 vdd.n1314 gnd 0.006957f
C3895 vdd.t153 gnd 0.281145f
C3896 vdd.t154 gnd 0.287787f
C3897 vdd.t151 gnd 0.183542f
C3898 vdd.n1315 gnd 0.099195f
C3899 vdd.n1316 gnd 0.056266f
C3900 vdd.n1317 gnd 0.009943f
C3901 vdd.n1318 gnd 0.006957f
C3902 vdd.t190 gnd 0.281145f
C3903 vdd.t191 gnd 0.287787f
C3904 vdd.t189 gnd 0.183542f
C3905 vdd.n1319 gnd 0.099195f
C3906 vdd.n1320 gnd 0.056266f
C3907 vdd.n1321 gnd 0.006957f
C3908 vdd.n1322 gnd 0.006957f
C3909 vdd.n1323 gnd 0.006957f
C3910 vdd.n1324 gnd 0.006957f
C3911 vdd.n1325 gnd 0.006957f
C3912 vdd.n1326 gnd 0.006957f
C3913 vdd.n1327 gnd 0.006957f
C3914 vdd.n1328 gnd 0.006957f
C3915 vdd.n1329 gnd 0.006957f
C3916 vdd.n1330 gnd 0.006957f
C3917 vdd.n1331 gnd 0.006957f
C3918 vdd.n1332 gnd 0.006957f
C3919 vdd.n1333 gnd 0.006957f
C3920 vdd.n1334 gnd 0.006957f
C3921 vdd.n1335 gnd 0.006957f
C3922 vdd.n1336 gnd 0.006957f
C3923 vdd.n1337 gnd 0.006957f
C3924 vdd.n1338 gnd 0.006957f
C3925 vdd.n1339 gnd 0.006957f
C3926 vdd.n1340 gnd 0.006957f
C3927 vdd.n1341 gnd 0.006957f
C3928 vdd.n1342 gnd 0.006957f
C3929 vdd.n1343 gnd 0.006957f
C3930 vdd.n1344 gnd 0.006957f
C3931 vdd.n1345 gnd 0.006957f
C3932 vdd.n1346 gnd 0.006957f
C3933 vdd.n1347 gnd 0.005065f
C3934 vdd.n1348 gnd 0.009943f
C3935 vdd.n1349 gnd 0.005371f
C3936 vdd.n1350 gnd 0.006957f
C3937 vdd.n1351 gnd 0.006957f
C3938 vdd.n1352 gnd 0.006957f
C3939 vdd.n1353 gnd 0.015797f
C3940 vdd.n1354 gnd 0.015797f
C3941 vdd.n1355 gnd 0.014897f
C3942 vdd.n1356 gnd 0.014897f
C3943 vdd.n1357 gnd 0.006957f
C3944 vdd.n1358 gnd 0.006957f
C3945 vdd.n1359 gnd 0.006957f
C3946 vdd.n1360 gnd 0.006957f
C3947 vdd.n1361 gnd 0.006957f
C3948 vdd.n1362 gnd 0.006957f
C3949 vdd.n1363 gnd 0.006957f
C3950 vdd.n1364 gnd 0.006957f
C3951 vdd.n1365 gnd 0.006957f
C3952 vdd.n1366 gnd 0.006957f
C3953 vdd.n1367 gnd 0.006957f
C3954 vdd.n1368 gnd 0.006957f
C3955 vdd.n1369 gnd 0.006957f
C3956 vdd.n1370 gnd 0.006957f
C3957 vdd.n1371 gnd 0.006957f
C3958 vdd.n1372 gnd 0.006957f
C3959 vdd.n1373 gnd 0.006957f
C3960 vdd.n1374 gnd 0.006957f
C3961 vdd.n1375 gnd 0.006957f
C3962 vdd.n1376 gnd 0.006957f
C3963 vdd.n1377 gnd 0.006957f
C3964 vdd.n1378 gnd 0.006957f
C3965 vdd.n1379 gnd 0.006957f
C3966 vdd.n1380 gnd 0.006957f
C3967 vdd.n1381 gnd 0.006957f
C3968 vdd.n1382 gnd 0.006957f
C3969 vdd.n1383 gnd 0.006957f
C3970 vdd.n1384 gnd 0.006957f
C3971 vdd.n1385 gnd 0.006957f
C3972 vdd.n1386 gnd 0.006957f
C3973 vdd.n1387 gnd 0.006957f
C3974 vdd.n1388 gnd 0.006957f
C3975 vdd.n1389 gnd 0.006957f
C3976 vdd.n1390 gnd 0.006957f
C3977 vdd.n1391 gnd 0.006957f
C3978 vdd.n1392 gnd 0.006957f
C3979 vdd.n1393 gnd 0.006957f
C3980 vdd.n1394 gnd 0.006957f
C3981 vdd.n1395 gnd 0.006957f
C3982 vdd.n1396 gnd 0.006957f
C3983 vdd.n1397 gnd 0.006957f
C3984 vdd.n1398 gnd 0.006957f
C3985 vdd.n1399 gnd 0.423468f
C3986 vdd.n1400 gnd 0.006957f
C3987 vdd.n1401 gnd 0.006957f
C3988 vdd.n1402 gnd 0.006957f
C3989 vdd.n1403 gnd 0.006957f
C3990 vdd.n1404 gnd 0.006957f
C3991 vdd.n1405 gnd 0.006957f
C3992 vdd.n1406 gnd 0.006957f
C3993 vdd.n1407 gnd 0.006957f
C3994 vdd.n1408 gnd 0.006957f
C3995 vdd.n1409 gnd 0.006957f
C3996 vdd.n1410 gnd 0.006957f
C3997 vdd.n1411 gnd 0.006957f
C3998 vdd.n1412 gnd 0.006957f
C3999 vdd.n1413 gnd 0.006957f
C4000 vdd.n1414 gnd 0.006957f
C4001 vdd.n1415 gnd 0.006957f
C4002 vdd.n1416 gnd 0.006957f
C4003 vdd.n1417 gnd 0.006957f
C4004 vdd.n1418 gnd 0.006957f
C4005 vdd.n1419 gnd 0.006957f
C4006 vdd.n1420 gnd 0.006957f
C4007 vdd.n1421 gnd 0.006957f
C4008 vdd.n1422 gnd 0.006957f
C4009 vdd.n1423 gnd 0.006957f
C4010 vdd.n1424 gnd 0.006957f
C4011 vdd.n1425 gnd 0.643044f
C4012 vdd.n1426 gnd 0.006957f
C4013 vdd.n1427 gnd 0.006957f
C4014 vdd.n1428 gnd 0.006957f
C4015 vdd.n1429 gnd 0.006957f
C4016 vdd.n1430 gnd 0.006957f
C4017 vdd.n1431 gnd 0.006957f
C4018 vdd.n1432 gnd 0.006957f
C4019 vdd.n1433 gnd 0.006957f
C4020 vdd.n1434 gnd 0.006957f
C4021 vdd.n1435 gnd 0.006957f
C4022 vdd.n1436 gnd 0.006957f
C4023 vdd.n1437 gnd 0.224804f
C4024 vdd.n1438 gnd 0.006957f
C4025 vdd.n1439 gnd 0.006957f
C4026 vdd.n1440 gnd 0.006957f
C4027 vdd.n1441 gnd 0.006957f
C4028 vdd.n1442 gnd 0.006957f
C4029 vdd.n1443 gnd 0.006957f
C4030 vdd.n1444 gnd 0.006957f
C4031 vdd.n1445 gnd 0.006957f
C4032 vdd.n1446 gnd 0.006957f
C4033 vdd.n1447 gnd 0.006957f
C4034 vdd.n1448 gnd 0.006957f
C4035 vdd.n1449 gnd 0.006957f
C4036 vdd.n1450 gnd 0.006957f
C4037 vdd.n1451 gnd 0.006957f
C4038 vdd.n1452 gnd 0.006957f
C4039 vdd.n1453 gnd 0.006957f
C4040 vdd.n1454 gnd 0.006957f
C4041 vdd.n1455 gnd 0.006957f
C4042 vdd.n1456 gnd 0.006957f
C4043 vdd.n1457 gnd 0.006957f
C4044 vdd.n1458 gnd 0.006957f
C4045 vdd.n1459 gnd 0.006957f
C4046 vdd.n1460 gnd 0.006957f
C4047 vdd.n1461 gnd 0.006957f
C4048 vdd.n1462 gnd 0.006957f
C4049 vdd.n1463 gnd 0.006957f
C4050 vdd.n1464 gnd 0.006957f
C4051 vdd.n1465 gnd 0.006957f
C4052 vdd.n1466 gnd 0.006957f
C4053 vdd.n1467 gnd 0.006957f
C4054 vdd.n1468 gnd 0.006957f
C4055 vdd.n1469 gnd 0.006957f
C4056 vdd.n1470 gnd 0.006957f
C4057 vdd.n1471 gnd 0.006957f
C4058 vdd.n1472 gnd 0.006957f
C4059 vdd.n1473 gnd 0.006957f
C4060 vdd.n1474 gnd 0.006957f
C4061 vdd.n1475 gnd 0.006957f
C4062 vdd.n1476 gnd 0.006957f
C4063 vdd.n1477 gnd 0.006957f
C4064 vdd.n1478 gnd 0.006957f
C4065 vdd.n1479 gnd 0.006957f
C4066 vdd.n1480 gnd 0.014897f
C4067 vdd.n1481 gnd 0.014897f
C4068 vdd.n1482 gnd 0.015797f
C4069 vdd.n1483 gnd 0.006957f
C4070 vdd.n1484 gnd 0.006957f
C4071 vdd.n1485 gnd 0.005371f
C4072 vdd.n1486 gnd 0.006957f
C4073 vdd.n1487 gnd 0.006957f
C4074 vdd.n1488 gnd 0.005065f
C4075 vdd.n1489 gnd 0.006957f
C4076 vdd.n1490 gnd 0.006957f
C4077 vdd.n1491 gnd 0.006957f
C4078 vdd.n1492 gnd 0.006957f
C4079 vdd.n1493 gnd 0.006957f
C4080 vdd.n1494 gnd 0.006957f
C4081 vdd.n1495 gnd 0.006957f
C4082 vdd.n1496 gnd 0.006957f
C4083 vdd.n1497 gnd 0.006957f
C4084 vdd.n1498 gnd 0.006957f
C4085 vdd.n1499 gnd 0.006957f
C4086 vdd.n1500 gnd 0.006957f
C4087 vdd.n1501 gnd 0.006957f
C4088 vdd.n1502 gnd 0.006957f
C4089 vdd.n1503 gnd 0.006957f
C4090 vdd.n1504 gnd 0.006957f
C4091 vdd.n1505 gnd 0.006957f
C4092 vdd.n1506 gnd 0.006957f
C4093 vdd.n1507 gnd 0.006957f
C4094 vdd.n1508 gnd 0.006957f
C4095 vdd.n1509 gnd 0.006957f
C4096 vdd.n1510 gnd 0.006957f
C4097 vdd.n1511 gnd 0.006957f
C4098 vdd.n1512 gnd 0.006957f
C4099 vdd.n1513 gnd 0.006957f
C4100 vdd.n1514 gnd 0.006957f
C4101 vdd.n1515 gnd 0.046868f
C4102 vdd.n1517 gnd 0.025281f
C4103 vdd.n1518 gnd 0.008235f
C4104 vdd.n1520 gnd 0.010231f
C4105 vdd.n1521 gnd 0.008235f
C4106 vdd.n1522 gnd 0.010231f
C4107 vdd.n1524 gnd 0.010231f
C4108 vdd.n1525 gnd 0.010231f
C4109 vdd.n1527 gnd 0.010231f
C4110 vdd.n1528 gnd 0.006835f
C4111 vdd.t156 gnd 0.5228f
C4112 vdd.n1529 gnd 0.010231f
C4113 vdd.n1530 gnd 0.025281f
C4114 vdd.n1531 gnd 0.008235f
C4115 vdd.n1532 gnd 0.010231f
C4116 vdd.n1533 gnd 0.008235f
C4117 vdd.n1534 gnd 0.010231f
C4118 vdd.n1535 gnd 1.0456f
C4119 vdd.n1536 gnd 0.010231f
C4120 vdd.n1537 gnd 0.008235f
C4121 vdd.n1538 gnd 0.008235f
C4122 vdd.n1539 gnd 0.010231f
C4123 vdd.n1540 gnd 0.008235f
C4124 vdd.n1541 gnd 0.010231f
C4125 vdd.t11 gnd 0.5228f
C4126 vdd.n1542 gnd 0.010231f
C4127 vdd.n1543 gnd 0.008235f
C4128 vdd.n1544 gnd 0.010231f
C4129 vdd.n1545 gnd 0.008235f
C4130 vdd.n1546 gnd 0.010231f
C4131 vdd.t64 gnd 0.5228f
C4132 vdd.n1547 gnd 0.010231f
C4133 vdd.n1548 gnd 0.008235f
C4134 vdd.n1549 gnd 0.010231f
C4135 vdd.n1550 gnd 0.008235f
C4136 vdd.n1551 gnd 0.010231f
C4137 vdd.n1552 gnd 0.841707f
C4138 vdd.n1553 gnd 0.867847f
C4139 vdd.t15 gnd 0.5228f
C4140 vdd.n1554 gnd 0.010231f
C4141 vdd.n1555 gnd 0.008235f
C4142 vdd.n1556 gnd 0.010231f
C4143 vdd.n1557 gnd 0.008235f
C4144 vdd.n1558 gnd 0.010231f
C4145 vdd.n1559 gnd 0.663956f
C4146 vdd.n1560 gnd 0.010231f
C4147 vdd.n1561 gnd 0.008235f
C4148 vdd.n1562 gnd 0.010231f
C4149 vdd.n1563 gnd 0.008235f
C4150 vdd.n1564 gnd 0.010231f
C4151 vdd.t52 gnd 0.5228f
C4152 vdd.t68 gnd 0.5228f
C4153 vdd.n1565 gnd 0.010231f
C4154 vdd.n1566 gnd 0.008235f
C4155 vdd.n1567 gnd 0.010231f
C4156 vdd.n1568 gnd 0.008235f
C4157 vdd.n1569 gnd 0.010231f
C4158 vdd.t135 gnd 0.5228f
C4159 vdd.n1570 gnd 0.010231f
C4160 vdd.n1571 gnd 0.008235f
C4161 vdd.n1572 gnd 0.010231f
C4162 vdd.n1573 gnd 0.008235f
C4163 vdd.n1574 gnd 0.010231f
C4164 vdd.t87 gnd 0.5228f
C4165 vdd.n1575 gnd 0.737148f
C4166 vdd.n1576 gnd 0.010231f
C4167 vdd.n1577 gnd 0.008235f
C4168 vdd.n1578 gnd 0.010231f
C4169 vdd.n1579 gnd 0.008235f
C4170 vdd.n1580 gnd 0.010231f
C4171 vdd.n1581 gnd 0.820795f
C4172 vdd.n1582 gnd 0.010231f
C4173 vdd.n1583 gnd 0.008235f
C4174 vdd.n1584 gnd 0.010231f
C4175 vdd.n1585 gnd 0.008235f
C4176 vdd.n1586 gnd 0.010231f
C4177 vdd.n1587 gnd 0.643044f
C4178 vdd.t89 gnd 0.5228f
C4179 vdd.n1588 gnd 0.010231f
C4180 vdd.n1589 gnd 0.008235f
C4181 vdd.n1590 gnd 0.010231f
C4182 vdd.n1591 gnd 0.008235f
C4183 vdd.n1592 gnd 0.010231f
C4184 vdd.t35 gnd 0.5228f
C4185 vdd.n1593 gnd 0.010231f
C4186 vdd.n1594 gnd 0.008235f
C4187 vdd.n1595 gnd 0.010231f
C4188 vdd.n1596 gnd 0.008235f
C4189 vdd.n1597 gnd 0.010231f
C4190 vdd.t41 gnd 0.5228f
C4191 vdd.n1598 gnd 0.580308f
C4192 vdd.n1599 gnd 0.010231f
C4193 vdd.n1600 gnd 0.008235f
C4194 vdd.n1601 gnd 0.010231f
C4195 vdd.n1602 gnd 0.008235f
C4196 vdd.n1603 gnd 0.010231f
C4197 vdd.t109 gnd 0.5228f
C4198 vdd.n1604 gnd 0.010231f
C4199 vdd.n1605 gnd 0.008235f
C4200 vdd.n1606 gnd 0.010231f
C4201 vdd.n1607 gnd 0.008235f
C4202 vdd.n1608 gnd 0.010231f
C4203 vdd.n1609 gnd 0.799883f
C4204 vdd.n1610 gnd 0.867847f
C4205 vdd.t56 gnd 0.5228f
C4206 vdd.n1611 gnd 0.010231f
C4207 vdd.n1612 gnd 0.008235f
C4208 vdd.n1613 gnd 0.010231f
C4209 vdd.n1614 gnd 0.008235f
C4210 vdd.n1615 gnd 0.010231f
C4211 vdd.n1616 gnd 0.622132f
C4212 vdd.n1617 gnd 0.010231f
C4213 vdd.n1618 gnd 0.008235f
C4214 vdd.n1619 gnd 0.010231f
C4215 vdd.n1620 gnd 0.008235f
C4216 vdd.n1621 gnd 0.010231f
C4217 vdd.t106 gnd 0.5228f
C4218 vdd.t123 gnd 0.5228f
C4219 vdd.n1622 gnd 0.010231f
C4220 vdd.n1623 gnd 0.008235f
C4221 vdd.n1624 gnd 0.010231f
C4222 vdd.n1625 gnd 0.008235f
C4223 vdd.n1626 gnd 0.010231f
C4224 vdd.t9 gnd 0.5228f
C4225 vdd.n1627 gnd 0.010231f
C4226 vdd.n1628 gnd 0.008235f
C4227 vdd.n1629 gnd 0.010231f
C4228 vdd.n1630 gnd 0.008235f
C4229 vdd.n1631 gnd 0.010231f
C4230 vdd.t66 gnd 0.5228f
C4231 vdd.n1632 gnd 0.778971f
C4232 vdd.n1633 gnd 0.010231f
C4233 vdd.n1634 gnd 0.008235f
C4234 vdd.n1635 gnd 0.010231f
C4235 vdd.n1636 gnd 0.008235f
C4236 vdd.n1637 gnd 0.010231f
C4237 vdd.n1638 gnd 1.0456f
C4238 vdd.n1639 gnd 0.010231f
C4239 vdd.n1640 gnd 0.008235f
C4240 vdd.n1641 gnd 0.024751f
C4241 vdd.n1642 gnd 0.006835f
C4242 vdd.n1643 gnd 0.024751f
C4243 vdd.t211 gnd 0.5228f
C4244 vdd.n1644 gnd 0.024751f
C4245 vdd.n1645 gnd 0.006835f
C4246 vdd.n1646 gnd 0.010231f
C4247 vdd.n1647 gnd 0.008235f
C4248 vdd.n1648 gnd 0.010231f
C4249 vdd.n1679 gnd 0.025281f
C4250 vdd.n1680 gnd 1.54226f
C4251 vdd.n1681 gnd 0.010231f
C4252 vdd.n1682 gnd 0.008235f
C4253 vdd.n1683 gnd 0.010231f
C4254 vdd.n1684 gnd 0.010231f
C4255 vdd.n1685 gnd 0.010231f
C4256 vdd.n1686 gnd 0.010231f
C4257 vdd.n1687 gnd 0.010231f
C4258 vdd.n1688 gnd 0.008235f
C4259 vdd.n1689 gnd 0.010231f
C4260 vdd.n1690 gnd 0.010231f
C4261 vdd.n1691 gnd 0.010231f
C4262 vdd.n1692 gnd 0.010231f
C4263 vdd.n1693 gnd 0.010231f
C4264 vdd.n1694 gnd 0.008235f
C4265 vdd.n1695 gnd 0.010231f
C4266 vdd.n1696 gnd 0.010231f
C4267 vdd.n1697 gnd 0.010231f
C4268 vdd.n1698 gnd 0.010231f
C4269 vdd.n1699 gnd 0.010231f
C4270 vdd.n1700 gnd 0.008235f
C4271 vdd.n1701 gnd 0.010231f
C4272 vdd.n1702 gnd 0.010231f
C4273 vdd.n1703 gnd 0.010231f
C4274 vdd.n1704 gnd 0.010231f
C4275 vdd.n1705 gnd 0.010231f
C4276 vdd.t221 gnd 0.125873f
C4277 vdd.t222 gnd 0.134524f
C4278 vdd.t220 gnd 0.164388f
C4279 vdd.n1706 gnd 0.210723f
C4280 vdd.n1707 gnd 0.177869f
C4281 vdd.n1708 gnd 0.017623f
C4282 vdd.n1709 gnd 0.010231f
C4283 vdd.n1710 gnd 0.010231f
C4284 vdd.n1711 gnd 0.010231f
C4285 vdd.n1712 gnd 0.010231f
C4286 vdd.n1713 gnd 0.010231f
C4287 vdd.n1714 gnd 0.008235f
C4288 vdd.n1715 gnd 0.010231f
C4289 vdd.n1716 gnd 0.010231f
C4290 vdd.n1717 gnd 0.010231f
C4291 vdd.n1718 gnd 0.010231f
C4292 vdd.n1719 gnd 0.010231f
C4293 vdd.n1720 gnd 0.008235f
C4294 vdd.n1721 gnd 0.010231f
C4295 vdd.n1722 gnd 0.010231f
C4296 vdd.n1723 gnd 0.010231f
C4297 vdd.n1724 gnd 0.010231f
C4298 vdd.n1725 gnd 0.010231f
C4299 vdd.n1726 gnd 0.008235f
C4300 vdd.n1727 gnd 0.010231f
C4301 vdd.n1728 gnd 0.010231f
C4302 vdd.n1729 gnd 0.010231f
C4303 vdd.n1730 gnd 0.010231f
C4304 vdd.n1731 gnd 0.010231f
C4305 vdd.n1732 gnd 0.008235f
C4306 vdd.n1733 gnd 0.010231f
C4307 vdd.n1734 gnd 0.010231f
C4308 vdd.n1735 gnd 0.010231f
C4309 vdd.n1736 gnd 0.010231f
C4310 vdd.n1737 gnd 0.010231f
C4311 vdd.n1738 gnd 0.008235f
C4312 vdd.n1739 gnd 0.010231f
C4313 vdd.n1740 gnd 0.010231f
C4314 vdd.n1741 gnd 0.010231f
C4315 vdd.n1742 gnd 0.010231f
C4316 vdd.n1743 gnd 0.008235f
C4317 vdd.n1744 gnd 0.010231f
C4318 vdd.n1745 gnd 0.010231f
C4319 vdd.n1746 gnd 0.010231f
C4320 vdd.n1747 gnd 0.010231f
C4321 vdd.n1748 gnd 0.010231f
C4322 vdd.n1749 gnd 0.008235f
C4323 vdd.n1750 gnd 0.010231f
C4324 vdd.n1751 gnd 0.010231f
C4325 vdd.n1752 gnd 0.010231f
C4326 vdd.n1753 gnd 0.010231f
C4327 vdd.n1754 gnd 0.010231f
C4328 vdd.n1755 gnd 0.008235f
C4329 vdd.n1756 gnd 0.010231f
C4330 vdd.n1757 gnd 0.010231f
C4331 vdd.n1758 gnd 0.010231f
C4332 vdd.n1759 gnd 0.010231f
C4333 vdd.n1760 gnd 0.010231f
C4334 vdd.n1761 gnd 0.008235f
C4335 vdd.n1762 gnd 0.010231f
C4336 vdd.n1763 gnd 0.010231f
C4337 vdd.n1764 gnd 0.010231f
C4338 vdd.n1765 gnd 0.010231f
C4339 vdd.n1766 gnd 0.010231f
C4340 vdd.n1767 gnd 0.008235f
C4341 vdd.n1768 gnd 0.010231f
C4342 vdd.n1769 gnd 0.010231f
C4343 vdd.n1770 gnd 0.010231f
C4344 vdd.n1771 gnd 0.010231f
C4345 vdd.t218 gnd 0.125873f
C4346 vdd.t219 gnd 0.134524f
C4347 vdd.t217 gnd 0.164388f
C4348 vdd.n1772 gnd 0.210723f
C4349 vdd.n1773 gnd 0.177869f
C4350 vdd.n1774 gnd 0.013505f
C4351 vdd.n1775 gnd 0.003912f
C4352 vdd.n1776 gnd 0.025281f
C4353 vdd.n1777 gnd 0.010231f
C4354 vdd.n1778 gnd 0.004323f
C4355 vdd.n1779 gnd 0.008235f
C4356 vdd.n1780 gnd 0.008235f
C4357 vdd.n1781 gnd 0.010231f
C4358 vdd.n1782 gnd 0.010231f
C4359 vdd.n1783 gnd 0.010231f
C4360 vdd.n1784 gnd 0.008235f
C4361 vdd.n1785 gnd 0.008235f
C4362 vdd.n1786 gnd 0.008235f
C4363 vdd.n1787 gnd 0.010231f
C4364 vdd.n1788 gnd 0.010231f
C4365 vdd.n1789 gnd 0.010231f
C4366 vdd.n1790 gnd 0.008235f
C4367 vdd.n1791 gnd 0.008235f
C4368 vdd.n1792 gnd 0.008235f
C4369 vdd.n1793 gnd 0.010231f
C4370 vdd.n1794 gnd 0.010231f
C4371 vdd.n1795 gnd 0.010231f
C4372 vdd.n1796 gnd 0.008235f
C4373 vdd.n1797 gnd 0.008235f
C4374 vdd.n1798 gnd 0.008235f
C4375 vdd.n1799 gnd 0.010231f
C4376 vdd.n1800 gnd 0.010231f
C4377 vdd.n1801 gnd 0.010231f
C4378 vdd.n1802 gnd 0.008235f
C4379 vdd.n1803 gnd 0.008235f
C4380 vdd.n1804 gnd 0.008235f
C4381 vdd.n1805 gnd 0.010231f
C4382 vdd.n1806 gnd 0.010231f
C4383 vdd.n1807 gnd 0.010231f
C4384 vdd.n1808 gnd 0.008153f
C4385 vdd.n1809 gnd 0.010231f
C4386 vdd.t212 gnd 0.125873f
C4387 vdd.t213 gnd 0.134524f
C4388 vdd.t210 gnd 0.164388f
C4389 vdd.n1810 gnd 0.210723f
C4390 vdd.n1811 gnd 0.177869f
C4391 vdd.n1812 gnd 0.017623f
C4392 vdd.n1813 gnd 0.0056f
C4393 vdd.n1814 gnd 0.010231f
C4394 vdd.n1815 gnd 0.010231f
C4395 vdd.n1816 gnd 0.010231f
C4396 vdd.n1817 gnd 0.008235f
C4397 vdd.n1818 gnd 0.008235f
C4398 vdd.n1819 gnd 0.008235f
C4399 vdd.n1820 gnd 0.010231f
C4400 vdd.n1821 gnd 0.010231f
C4401 vdd.n1822 gnd 0.010231f
C4402 vdd.n1823 gnd 0.008235f
C4403 vdd.n1824 gnd 0.008235f
C4404 vdd.n1825 gnd 0.008235f
C4405 vdd.n1826 gnd 0.010231f
C4406 vdd.n1827 gnd 0.010231f
C4407 vdd.n1828 gnd 0.010231f
C4408 vdd.n1829 gnd 0.008235f
C4409 vdd.n1830 gnd 0.008235f
C4410 vdd.n1831 gnd 0.008235f
C4411 vdd.n1832 gnd 0.010231f
C4412 vdd.n1833 gnd 0.010231f
C4413 vdd.n1834 gnd 0.010231f
C4414 vdd.n1835 gnd 0.008235f
C4415 vdd.n1836 gnd 0.008235f
C4416 vdd.n1837 gnd 0.008235f
C4417 vdd.n1838 gnd 0.010231f
C4418 vdd.n1839 gnd 0.010231f
C4419 vdd.n1840 gnd 0.010231f
C4420 vdd.n1841 gnd 0.008235f
C4421 vdd.n1842 gnd 0.008235f
C4422 vdd.n1843 gnd 0.006876f
C4423 vdd.n1844 gnd 0.010231f
C4424 vdd.n1845 gnd 0.010231f
C4425 vdd.n1846 gnd 0.010231f
C4426 vdd.n1847 gnd 0.006876f
C4427 vdd.n1848 gnd 0.008235f
C4428 vdd.n1849 gnd 0.008235f
C4429 vdd.n1850 gnd 0.010231f
C4430 vdd.n1851 gnd 0.010231f
C4431 vdd.n1852 gnd 0.010231f
C4432 vdd.n1853 gnd 0.008235f
C4433 vdd.n1854 gnd 0.008235f
C4434 vdd.n1855 gnd 0.008235f
C4435 vdd.n1856 gnd 0.010231f
C4436 vdd.n1857 gnd 0.010231f
C4437 vdd.n1858 gnd 0.010231f
C4438 vdd.n1859 gnd 0.008235f
C4439 vdd.n1860 gnd 0.008235f
C4440 vdd.n1861 gnd 0.008235f
C4441 vdd.n1862 gnd 0.010231f
C4442 vdd.n1863 gnd 0.010231f
C4443 vdd.n1864 gnd 0.010231f
C4444 vdd.n1865 gnd 0.008235f
C4445 vdd.n1866 gnd 0.008235f
C4446 vdd.n1867 gnd 0.008235f
C4447 vdd.n1868 gnd 0.010231f
C4448 vdd.n1869 gnd 0.010231f
C4449 vdd.n1870 gnd 0.010231f
C4450 vdd.n1871 gnd 0.008235f
C4451 vdd.n1872 gnd 0.010231f
C4452 vdd.n1873 gnd 2.47807f
C4453 vdd.n1875 gnd 0.025281f
C4454 vdd.n1876 gnd 0.006835f
C4455 vdd.n1877 gnd 0.025281f
C4456 vdd.n1878 gnd 0.024751f
C4457 vdd.n1879 gnd 0.010231f
C4458 vdd.n1880 gnd 0.008235f
C4459 vdd.n1881 gnd 0.010231f
C4460 vdd.n1882 gnd 0.528028f
C4461 vdd.n1883 gnd 0.010231f
C4462 vdd.n1884 gnd 0.008235f
C4463 vdd.n1885 gnd 0.010231f
C4464 vdd.n1886 gnd 0.010231f
C4465 vdd.n1887 gnd 0.010231f
C4466 vdd.n1888 gnd 0.008235f
C4467 vdd.n1889 gnd 0.010231f
C4468 vdd.n1890 gnd 0.956723f
C4469 vdd.n1891 gnd 1.0456f
C4470 vdd.n1892 gnd 0.010231f
C4471 vdd.n1893 gnd 0.008235f
C4472 vdd.n1894 gnd 0.010231f
C4473 vdd.n1895 gnd 0.010231f
C4474 vdd.n1896 gnd 0.010231f
C4475 vdd.n1897 gnd 0.008235f
C4476 vdd.n1898 gnd 0.010231f
C4477 vdd.n1899 gnd 0.611676f
C4478 vdd.n1900 gnd 0.010231f
C4479 vdd.n1901 gnd 0.008235f
C4480 vdd.n1902 gnd 0.010231f
C4481 vdd.n1903 gnd 0.010231f
C4482 vdd.n1904 gnd 0.010231f
C4483 vdd.n1905 gnd 0.008235f
C4484 vdd.n1906 gnd 0.010231f
C4485 vdd.n1907 gnd 0.60122f
C4486 vdd.n1908 gnd 0.789427f
C4487 vdd.n1909 gnd 0.010231f
C4488 vdd.n1910 gnd 0.008235f
C4489 vdd.n1911 gnd 0.010231f
C4490 vdd.n1912 gnd 0.010231f
C4491 vdd.n1913 gnd 0.010231f
C4492 vdd.n1914 gnd 0.008235f
C4493 vdd.n1915 gnd 0.010231f
C4494 vdd.n1916 gnd 0.867847f
C4495 vdd.n1917 gnd 0.010231f
C4496 vdd.n1918 gnd 0.008235f
C4497 vdd.n1919 gnd 0.010231f
C4498 vdd.n1920 gnd 0.010231f
C4499 vdd.n1921 gnd 0.010231f
C4500 vdd.n1922 gnd 0.008235f
C4501 vdd.n1923 gnd 0.010231f
C4502 vdd.t24 gnd 0.5228f
C4503 vdd.n1924 gnd 0.768516f
C4504 vdd.n1925 gnd 0.010231f
C4505 vdd.n1926 gnd 0.008235f
C4506 vdd.n1927 gnd 0.010231f
C4507 vdd.n1928 gnd 0.010231f
C4508 vdd.n1929 gnd 0.010231f
C4509 vdd.n1930 gnd 0.008235f
C4510 vdd.n1931 gnd 0.010231f
C4511 vdd.n1932 gnd 0.590764f
C4512 vdd.n1933 gnd 0.010231f
C4513 vdd.n1934 gnd 0.008235f
C4514 vdd.n1935 gnd 0.010231f
C4515 vdd.n1936 gnd 0.010231f
C4516 vdd.n1937 gnd 0.010231f
C4517 vdd.n1938 gnd 0.008235f
C4518 vdd.n1939 gnd 0.010231f
C4519 vdd.n1940 gnd 0.75806f
C4520 vdd.n1941 gnd 0.632588f
C4521 vdd.n1942 gnd 0.010231f
C4522 vdd.n1943 gnd 0.008235f
C4523 vdd.n1944 gnd 0.010231f
C4524 vdd.n1945 gnd 0.010231f
C4525 vdd.n1946 gnd 0.010231f
C4526 vdd.n1947 gnd 0.008235f
C4527 vdd.n1948 gnd 0.010231f
C4528 vdd.n1949 gnd 0.810339f
C4529 vdd.n1950 gnd 0.010231f
C4530 vdd.n1951 gnd 0.008235f
C4531 vdd.n1952 gnd 0.010231f
C4532 vdd.n1953 gnd 0.010231f
C4533 vdd.n1954 gnd 0.010231f
C4534 vdd.n1955 gnd 0.008235f
C4535 vdd.n1956 gnd 0.010231f
C4536 vdd.t7 gnd 0.5228f
C4537 vdd.n1957 gnd 0.867847f
C4538 vdd.n1958 gnd 0.010231f
C4539 vdd.n1959 gnd 0.008235f
C4540 vdd.n1960 gnd 0.010231f
C4541 vdd.n1961 gnd 0.007863f
C4542 vdd.n1962 gnd 0.005615f
C4543 vdd.n1963 gnd 0.005211f
C4544 vdd.n1964 gnd 0.002882f
C4545 vdd.n1965 gnd 0.006618f
C4546 vdd.n1966 gnd 0.0028f
C4547 vdd.n1967 gnd 0.002965f
C4548 vdd.n1968 gnd 0.005211f
C4549 vdd.n1969 gnd 0.0028f
C4550 vdd.n1970 gnd 0.006618f
C4551 vdd.n1971 gnd 0.002965f
C4552 vdd.n1972 gnd 0.005211f
C4553 vdd.n1973 gnd 0.0028f
C4554 vdd.n1974 gnd 0.004963f
C4555 vdd.n1975 gnd 0.004978f
C4556 vdd.t12 gnd 0.014218f
C4557 vdd.n1976 gnd 0.031635f
C4558 vdd.n1977 gnd 0.164637f
C4559 vdd.n1978 gnd 0.0028f
C4560 vdd.n1979 gnd 0.002965f
C4561 vdd.n1980 gnd 0.006618f
C4562 vdd.n1981 gnd 0.006618f
C4563 vdd.n1982 gnd 0.002965f
C4564 vdd.n1983 gnd 0.0028f
C4565 vdd.n1984 gnd 0.005211f
C4566 vdd.n1985 gnd 0.005211f
C4567 vdd.n1986 gnd 0.0028f
C4568 vdd.n1987 gnd 0.002965f
C4569 vdd.n1988 gnd 0.006618f
C4570 vdd.n1989 gnd 0.006618f
C4571 vdd.n1990 gnd 0.002965f
C4572 vdd.n1991 gnd 0.0028f
C4573 vdd.n1992 gnd 0.005211f
C4574 vdd.n1993 gnd 0.005211f
C4575 vdd.n1994 gnd 0.0028f
C4576 vdd.n1995 gnd 0.002965f
C4577 vdd.n1996 gnd 0.006618f
C4578 vdd.n1997 gnd 0.006618f
C4579 vdd.n1998 gnd 0.015646f
C4580 vdd.n1999 gnd 0.002882f
C4581 vdd.n2000 gnd 0.0028f
C4582 vdd.n2001 gnd 0.013467f
C4583 vdd.n2002 gnd 0.009402f
C4584 vdd.t16 gnd 0.03294f
C4585 vdd.t296 gnd 0.03294f
C4586 vdd.n2003 gnd 0.226387f
C4587 vdd.n2004 gnd 0.178019f
C4588 vdd.t77 gnd 0.03294f
C4589 vdd.t285 gnd 0.03294f
C4590 vdd.n2005 gnd 0.226387f
C4591 vdd.n2006 gnd 0.14366f
C4592 vdd.t292 gnd 0.03294f
C4593 vdd.t53 gnd 0.03294f
C4594 vdd.n2007 gnd 0.226387f
C4595 vdd.n2008 gnd 0.14366f
C4596 vdd.t50 gnd 0.03294f
C4597 vdd.t130 gnd 0.03294f
C4598 vdd.n2009 gnd 0.226387f
C4599 vdd.n2010 gnd 0.14366f
C4600 vdd.t295 gnd 0.03294f
C4601 vdd.t90 gnd 0.03294f
C4602 vdd.n2011 gnd 0.226387f
C4603 vdd.n2012 gnd 0.14366f
C4604 vdd.t125 gnd 0.03294f
C4605 vdd.t36 gnd 0.03294f
C4606 vdd.n2013 gnd 0.226387f
C4607 vdd.n2014 gnd 0.14366f
C4608 vdd.t303 gnd 0.03294f
C4609 vdd.t110 gnd 0.03294f
C4610 vdd.n2015 gnd 0.226387f
C4611 vdd.n2016 gnd 0.14366f
C4612 vdd.t281 gnd 0.03294f
C4613 vdd.t54 gnd 0.03294f
C4614 vdd.n2017 gnd 0.226387f
C4615 vdd.n2018 gnd 0.14366f
C4616 vdd.t48 gnd 0.03294f
C4617 vdd.t139 gnd 0.03294f
C4618 vdd.n2019 gnd 0.226387f
C4619 vdd.n2020 gnd 0.14366f
C4620 vdd.n2021 gnd 0.005615f
C4621 vdd.n2022 gnd 0.005211f
C4622 vdd.n2023 gnd 0.002882f
C4623 vdd.n2024 gnd 0.006618f
C4624 vdd.n2025 gnd 0.0028f
C4625 vdd.n2026 gnd 0.002965f
C4626 vdd.n2027 gnd 0.005211f
C4627 vdd.n2028 gnd 0.0028f
C4628 vdd.n2029 gnd 0.006618f
C4629 vdd.n2030 gnd 0.002965f
C4630 vdd.n2031 gnd 0.005211f
C4631 vdd.n2032 gnd 0.0028f
C4632 vdd.n2033 gnd 0.004963f
C4633 vdd.n2034 gnd 0.004978f
C4634 vdd.t116 gnd 0.014218f
C4635 vdd.n2035 gnd 0.031635f
C4636 vdd.n2036 gnd 0.164637f
C4637 vdd.n2037 gnd 0.0028f
C4638 vdd.n2038 gnd 0.002965f
C4639 vdd.n2039 gnd 0.006618f
C4640 vdd.n2040 gnd 0.006618f
C4641 vdd.n2041 gnd 0.002965f
C4642 vdd.n2042 gnd 0.0028f
C4643 vdd.n2043 gnd 0.005211f
C4644 vdd.n2044 gnd 0.005211f
C4645 vdd.n2045 gnd 0.0028f
C4646 vdd.n2046 gnd 0.002965f
C4647 vdd.n2047 gnd 0.006618f
C4648 vdd.n2048 gnd 0.006618f
C4649 vdd.n2049 gnd 0.002965f
C4650 vdd.n2050 gnd 0.0028f
C4651 vdd.n2051 gnd 0.005211f
C4652 vdd.n2052 gnd 0.005211f
C4653 vdd.n2053 gnd 0.0028f
C4654 vdd.n2054 gnd 0.002965f
C4655 vdd.n2055 gnd 0.006618f
C4656 vdd.n2056 gnd 0.006618f
C4657 vdd.n2057 gnd 0.015646f
C4658 vdd.n2058 gnd 0.002882f
C4659 vdd.n2059 gnd 0.0028f
C4660 vdd.n2060 gnd 0.013467f
C4661 vdd.n2061 gnd 0.009107f
C4662 vdd.n2062 gnd 0.106884f
C4663 vdd.n2063 gnd 0.005615f
C4664 vdd.n2064 gnd 0.005211f
C4665 vdd.n2065 gnd 0.002882f
C4666 vdd.n2066 gnd 0.006618f
C4667 vdd.n2067 gnd 0.0028f
C4668 vdd.n2068 gnd 0.002965f
C4669 vdd.n2069 gnd 0.005211f
C4670 vdd.n2070 gnd 0.0028f
C4671 vdd.n2071 gnd 0.006618f
C4672 vdd.n2072 gnd 0.002965f
C4673 vdd.n2073 gnd 0.005211f
C4674 vdd.n2074 gnd 0.0028f
C4675 vdd.n2075 gnd 0.004963f
C4676 vdd.n2076 gnd 0.004978f
C4677 vdd.t58 gnd 0.014218f
C4678 vdd.n2077 gnd 0.031635f
C4679 vdd.n2078 gnd 0.164637f
C4680 vdd.n2079 gnd 0.0028f
C4681 vdd.n2080 gnd 0.002965f
C4682 vdd.n2081 gnd 0.006618f
C4683 vdd.n2082 gnd 0.006618f
C4684 vdd.n2083 gnd 0.002965f
C4685 vdd.n2084 gnd 0.0028f
C4686 vdd.n2085 gnd 0.005211f
C4687 vdd.n2086 gnd 0.005211f
C4688 vdd.n2087 gnd 0.0028f
C4689 vdd.n2088 gnd 0.002965f
C4690 vdd.n2089 gnd 0.006618f
C4691 vdd.n2090 gnd 0.006618f
C4692 vdd.n2091 gnd 0.002965f
C4693 vdd.n2092 gnd 0.0028f
C4694 vdd.n2093 gnd 0.005211f
C4695 vdd.n2094 gnd 0.005211f
C4696 vdd.n2095 gnd 0.0028f
C4697 vdd.n2096 gnd 0.002965f
C4698 vdd.n2097 gnd 0.006618f
C4699 vdd.n2098 gnd 0.006618f
C4700 vdd.n2099 gnd 0.015646f
C4701 vdd.n2100 gnd 0.002882f
C4702 vdd.n2101 gnd 0.0028f
C4703 vdd.n2102 gnd 0.013467f
C4704 vdd.n2103 gnd 0.009402f
C4705 vdd.t293 gnd 0.03294f
C4706 vdd.t301 gnd 0.03294f
C4707 vdd.n2104 gnd 0.226387f
C4708 vdd.n2105 gnd 0.178019f
C4709 vdd.t69 gnd 0.03294f
C4710 vdd.t128 gnd 0.03294f
C4711 vdd.n2106 gnd 0.226387f
C4712 vdd.n2107 gnd 0.14366f
C4713 vdd.t136 gnd 0.03294f
C4714 vdd.t287 gnd 0.03294f
C4715 vdd.n2108 gnd 0.226387f
C4716 vdd.n2109 gnd 0.14366f
C4717 vdd.t305 gnd 0.03294f
C4718 vdd.t129 gnd 0.03294f
C4719 vdd.n2110 gnd 0.226387f
C4720 vdd.n2111 gnd 0.14366f
C4721 vdd.t127 gnd 0.03294f
C4722 vdd.t112 gnd 0.03294f
C4723 vdd.n2112 gnd 0.226387f
C4724 vdd.n2113 gnd 0.14366f
C4725 vdd.t42 gnd 0.03294f
C4726 vdd.t74 gnd 0.03294f
C4727 vdd.n2114 gnd 0.226387f
C4728 vdd.n2115 gnd 0.14366f
C4729 vdd.t57 gnd 0.03294f
C4730 vdd.t113 gnd 0.03294f
C4731 vdd.n2116 gnd 0.226387f
C4732 vdd.n2117 gnd 0.14366f
C4733 vdd.t124 gnd 0.03294f
C4734 vdd.t300 gnd 0.03294f
C4735 vdd.n2118 gnd 0.226387f
C4736 vdd.n2119 gnd 0.14366f
C4737 vdd.t10 gnd 0.03294f
C4738 vdd.t298 gnd 0.03294f
C4739 vdd.n2120 gnd 0.226387f
C4740 vdd.n2121 gnd 0.14366f
C4741 vdd.n2122 gnd 0.005615f
C4742 vdd.n2123 gnd 0.005211f
C4743 vdd.n2124 gnd 0.002882f
C4744 vdd.n2125 gnd 0.006618f
C4745 vdd.n2126 gnd 0.0028f
C4746 vdd.n2127 gnd 0.002965f
C4747 vdd.n2128 gnd 0.005211f
C4748 vdd.n2129 gnd 0.0028f
C4749 vdd.n2130 gnd 0.006618f
C4750 vdd.n2131 gnd 0.002965f
C4751 vdd.n2132 gnd 0.005211f
C4752 vdd.n2133 gnd 0.0028f
C4753 vdd.n2134 gnd 0.004963f
C4754 vdd.n2135 gnd 0.004978f
C4755 vdd.t286 gnd 0.014218f
C4756 vdd.n2136 gnd 0.031635f
C4757 vdd.n2137 gnd 0.164637f
C4758 vdd.n2138 gnd 0.0028f
C4759 vdd.n2139 gnd 0.002965f
C4760 vdd.n2140 gnd 0.006618f
C4761 vdd.n2141 gnd 0.006618f
C4762 vdd.n2142 gnd 0.002965f
C4763 vdd.n2143 gnd 0.0028f
C4764 vdd.n2144 gnd 0.005211f
C4765 vdd.n2145 gnd 0.005211f
C4766 vdd.n2146 gnd 0.0028f
C4767 vdd.n2147 gnd 0.002965f
C4768 vdd.n2148 gnd 0.006618f
C4769 vdd.n2149 gnd 0.006618f
C4770 vdd.n2150 gnd 0.002965f
C4771 vdd.n2151 gnd 0.0028f
C4772 vdd.n2152 gnd 0.005211f
C4773 vdd.n2153 gnd 0.005211f
C4774 vdd.n2154 gnd 0.0028f
C4775 vdd.n2155 gnd 0.002965f
C4776 vdd.n2156 gnd 0.006618f
C4777 vdd.n2157 gnd 0.006618f
C4778 vdd.n2158 gnd 0.015646f
C4779 vdd.n2159 gnd 0.002882f
C4780 vdd.n2160 gnd 0.0028f
C4781 vdd.n2161 gnd 0.013467f
C4782 vdd.n2162 gnd 0.009107f
C4783 vdd.n2163 gnd 0.063585f
C4784 vdd.n2164 gnd 0.229114f
C4785 vdd.n2165 gnd 0.005615f
C4786 vdd.n2166 gnd 0.005211f
C4787 vdd.n2167 gnd 0.002882f
C4788 vdd.n2168 gnd 0.006618f
C4789 vdd.n2169 gnd 0.0028f
C4790 vdd.n2170 gnd 0.002965f
C4791 vdd.n2171 gnd 0.005211f
C4792 vdd.n2172 gnd 0.0028f
C4793 vdd.n2173 gnd 0.006618f
C4794 vdd.n2174 gnd 0.002965f
C4795 vdd.n2175 gnd 0.005211f
C4796 vdd.n2176 gnd 0.0028f
C4797 vdd.n2177 gnd 0.004963f
C4798 vdd.n2178 gnd 0.004978f
C4799 vdd.t304 gnd 0.014218f
C4800 vdd.n2179 gnd 0.031635f
C4801 vdd.n2180 gnd 0.164637f
C4802 vdd.n2181 gnd 0.0028f
C4803 vdd.n2182 gnd 0.002965f
C4804 vdd.n2183 gnd 0.006618f
C4805 vdd.n2184 gnd 0.006618f
C4806 vdd.n2185 gnd 0.002965f
C4807 vdd.n2186 gnd 0.0028f
C4808 vdd.n2187 gnd 0.005211f
C4809 vdd.n2188 gnd 0.005211f
C4810 vdd.n2189 gnd 0.0028f
C4811 vdd.n2190 gnd 0.002965f
C4812 vdd.n2191 gnd 0.006618f
C4813 vdd.n2192 gnd 0.006618f
C4814 vdd.n2193 gnd 0.002965f
C4815 vdd.n2194 gnd 0.0028f
C4816 vdd.n2195 gnd 0.005211f
C4817 vdd.n2196 gnd 0.005211f
C4818 vdd.n2197 gnd 0.0028f
C4819 vdd.n2198 gnd 0.002965f
C4820 vdd.n2199 gnd 0.006618f
C4821 vdd.n2200 gnd 0.006618f
C4822 vdd.n2201 gnd 0.015646f
C4823 vdd.n2202 gnd 0.002882f
C4824 vdd.n2203 gnd 0.0028f
C4825 vdd.n2204 gnd 0.013467f
C4826 vdd.n2205 gnd 0.009402f
C4827 vdd.t23 gnd 0.03294f
C4828 vdd.t65 gnd 0.03294f
C4829 vdd.n2206 gnd 0.226387f
C4830 vdd.n2207 gnd 0.178019f
C4831 vdd.t105 gnd 0.03294f
C4832 vdd.t86 gnd 0.03294f
C4833 vdd.n2208 gnd 0.226387f
C4834 vdd.n2209 gnd 0.14366f
C4835 vdd.t284 gnd 0.03294f
C4836 vdd.t59 gnd 0.03294f
C4837 vdd.n2210 gnd 0.226387f
C4838 vdd.n2211 gnd 0.14366f
C4839 vdd.t108 gnd 0.03294f
C4840 vdd.t88 gnd 0.03294f
C4841 vdd.n2212 gnd 0.226387f
C4842 vdd.n2213 gnd 0.14366f
C4843 vdd.t8 gnd 0.03294f
C4844 vdd.t115 gnd 0.03294f
C4845 vdd.n2214 gnd 0.226387f
C4846 vdd.n2215 gnd 0.14366f
C4847 vdd.t143 gnd 0.03294f
C4848 vdd.t132 gnd 0.03294f
C4849 vdd.n2216 gnd 0.226387f
C4850 vdd.n2217 gnd 0.14366f
C4851 vdd.t291 gnd 0.03294f
C4852 vdd.t302 gnd 0.03294f
C4853 vdd.n2218 gnd 0.226387f
C4854 vdd.n2219 gnd 0.14366f
C4855 vdd.t282 gnd 0.03294f
C4856 vdd.t25 gnd 0.03294f
C4857 vdd.n2220 gnd 0.226387f
C4858 vdd.n2221 gnd 0.14366f
C4859 vdd.t60 gnd 0.03294f
C4860 vdd.t107 gnd 0.03294f
C4861 vdd.n2222 gnd 0.226387f
C4862 vdd.n2223 gnd 0.14366f
C4863 vdd.n2224 gnd 0.005615f
C4864 vdd.n2225 gnd 0.005211f
C4865 vdd.n2226 gnd 0.002882f
C4866 vdd.n2227 gnd 0.006618f
C4867 vdd.n2228 gnd 0.0028f
C4868 vdd.n2229 gnd 0.002965f
C4869 vdd.n2230 gnd 0.005211f
C4870 vdd.n2231 gnd 0.0028f
C4871 vdd.n2232 gnd 0.006618f
C4872 vdd.n2233 gnd 0.002965f
C4873 vdd.n2234 gnd 0.005211f
C4874 vdd.n2235 gnd 0.0028f
C4875 vdd.n2236 gnd 0.004963f
C4876 vdd.n2237 gnd 0.004978f
C4877 vdd.t67 gnd 0.014218f
C4878 vdd.n2238 gnd 0.031635f
C4879 vdd.n2239 gnd 0.164637f
C4880 vdd.n2240 gnd 0.0028f
C4881 vdd.n2241 gnd 0.002965f
C4882 vdd.n2242 gnd 0.006618f
C4883 vdd.n2243 gnd 0.006618f
C4884 vdd.n2244 gnd 0.002965f
C4885 vdd.n2245 gnd 0.0028f
C4886 vdd.n2246 gnd 0.005211f
C4887 vdd.n2247 gnd 0.005211f
C4888 vdd.n2248 gnd 0.0028f
C4889 vdd.n2249 gnd 0.002965f
C4890 vdd.n2250 gnd 0.006618f
C4891 vdd.n2251 gnd 0.006618f
C4892 vdd.n2252 gnd 0.002965f
C4893 vdd.n2253 gnd 0.0028f
C4894 vdd.n2254 gnd 0.005211f
C4895 vdd.n2255 gnd 0.005211f
C4896 vdd.n2256 gnd 0.0028f
C4897 vdd.n2257 gnd 0.002965f
C4898 vdd.n2258 gnd 0.006618f
C4899 vdd.n2259 gnd 0.006618f
C4900 vdd.n2260 gnd 0.015646f
C4901 vdd.n2261 gnd 0.002882f
C4902 vdd.n2262 gnd 0.0028f
C4903 vdd.n2263 gnd 0.013467f
C4904 vdd.n2264 gnd 0.009107f
C4905 vdd.n2265 gnd 0.063585f
C4906 vdd.n2266 gnd 0.262286f
C4907 vdd.n2267 gnd 2.99909f
C4908 vdd.n2268 gnd 0.603486f
C4909 vdd.n2269 gnd 0.007863f
C4910 vdd.n2270 gnd 0.008235f
C4911 vdd.n2271 gnd 0.010231f
C4912 vdd.n2272 gnd 0.747604f
C4913 vdd.n2273 gnd 0.010231f
C4914 vdd.n2274 gnd 0.008235f
C4915 vdd.n2275 gnd 0.010231f
C4916 vdd.n2276 gnd 0.010231f
C4917 vdd.n2277 gnd 0.010231f
C4918 vdd.n2278 gnd 0.008235f
C4919 vdd.n2279 gnd 0.010231f
C4920 vdd.n2280 gnd 0.867847f
C4921 vdd.t49 gnd 0.5228f
C4922 vdd.n2281 gnd 0.569852f
C4923 vdd.n2282 gnd 0.010231f
C4924 vdd.n2283 gnd 0.008235f
C4925 vdd.n2284 gnd 0.010231f
C4926 vdd.n2285 gnd 0.010231f
C4927 vdd.n2286 gnd 0.010231f
C4928 vdd.n2287 gnd 0.008235f
C4929 vdd.n2288 gnd 0.010231f
C4930 vdd.n2289 gnd 0.6535f
C4931 vdd.n2290 gnd 0.010231f
C4932 vdd.n2291 gnd 0.008235f
C4933 vdd.n2292 gnd 0.010231f
C4934 vdd.n2293 gnd 0.010231f
C4935 vdd.n2294 gnd 0.010231f
C4936 vdd.n2295 gnd 0.008235f
C4937 vdd.n2296 gnd 0.010231f
C4938 vdd.n2297 gnd 0.559396f
C4939 vdd.n2298 gnd 0.831251f
C4940 vdd.n2299 gnd 0.010231f
C4941 vdd.n2300 gnd 0.008235f
C4942 vdd.n2301 gnd 0.010231f
C4943 vdd.n2302 gnd 0.010231f
C4944 vdd.n2303 gnd 0.010231f
C4945 vdd.n2304 gnd 0.008235f
C4946 vdd.n2305 gnd 0.010231f
C4947 vdd.n2306 gnd 0.867847f
C4948 vdd.n2307 gnd 0.010231f
C4949 vdd.n2308 gnd 0.008235f
C4950 vdd.n2309 gnd 0.010231f
C4951 vdd.n2310 gnd 0.010231f
C4952 vdd.n2311 gnd 0.010231f
C4953 vdd.n2312 gnd 0.008235f
C4954 vdd.n2313 gnd 0.010231f
C4955 vdd.t85 gnd 0.5228f
C4956 vdd.n2314 gnd 0.726692f
C4957 vdd.n2315 gnd 0.010231f
C4958 vdd.n2316 gnd 0.008235f
C4959 vdd.n2317 gnd 0.010231f
C4960 vdd.n2318 gnd 0.010231f
C4961 vdd.n2319 gnd 0.010231f
C4962 vdd.n2320 gnd 0.008235f
C4963 vdd.n2321 gnd 0.010231f
C4964 vdd.n2322 gnd 0.54894f
C4965 vdd.n2323 gnd 0.010231f
C4966 vdd.n2324 gnd 0.008235f
C4967 vdd.n2325 gnd 0.010231f
C4968 vdd.n2326 gnd 0.010231f
C4969 vdd.n2327 gnd 0.010231f
C4970 vdd.n2328 gnd 0.008235f
C4971 vdd.n2329 gnd 0.010231f
C4972 vdd.n2330 gnd 0.716236f
C4973 vdd.n2331 gnd 0.674412f
C4974 vdd.n2332 gnd 0.010231f
C4975 vdd.n2333 gnd 0.008235f
C4976 vdd.n2334 gnd 0.010231f
C4977 vdd.n2335 gnd 0.010231f
C4978 vdd.n2336 gnd 0.010231f
C4979 vdd.n2337 gnd 0.008235f
C4980 vdd.n2338 gnd 0.010231f
C4981 vdd.n2339 gnd 0.852163f
C4982 vdd.n2340 gnd 0.010231f
C4983 vdd.n2341 gnd 0.008235f
C4984 vdd.n2342 gnd 0.010231f
C4985 vdd.n2343 gnd 0.010231f
C4986 vdd.n2344 gnd 0.024751f
C4987 vdd.n2345 gnd 0.010231f
C4988 vdd.n2346 gnd 0.010231f
C4989 vdd.n2347 gnd 0.008235f
C4990 vdd.n2348 gnd 0.010231f
C4991 vdd.n2349 gnd 0.632588f
C4992 vdd.n2350 gnd 1.0456f
C4993 vdd.n2351 gnd 0.010231f
C4994 vdd.n2352 gnd 0.008235f
C4995 vdd.n2353 gnd 0.010231f
C4996 vdd.n2354 gnd 0.010231f
C4997 vdd.n2355 gnd 0.024751f
C4998 vdd.n2356 gnd 0.006835f
C4999 vdd.n2357 gnd 0.024751f
C5000 vdd.n2358 gnd 1.4377f
C5001 vdd.n2359 gnd 0.024751f
C5002 vdd.n2360 gnd 0.025281f
C5003 vdd.n2361 gnd 0.003912f
C5004 vdd.t182 gnd 0.125873f
C5005 vdd.t181 gnd 0.134524f
C5006 vdd.t180 gnd 0.164388f
C5007 vdd.n2362 gnd 0.210723f
C5008 vdd.n2363 gnd 0.177045f
C5009 vdd.n2364 gnd 0.012682f
C5010 vdd.n2365 gnd 0.004323f
C5011 vdd.n2366 gnd 0.008799f
C5012 vdd.n2367 gnd 1.08617f
C5013 vdd.n2369 gnd 0.008235f
C5014 vdd.n2370 gnd 0.008235f
C5015 vdd.n2371 gnd 0.010231f
C5016 vdd.n2373 gnd 0.010231f
C5017 vdd.n2374 gnd 0.010231f
C5018 vdd.n2375 gnd 0.008235f
C5019 vdd.n2376 gnd 0.008235f
C5020 vdd.n2377 gnd 0.008235f
C5021 vdd.n2378 gnd 0.010231f
C5022 vdd.n2380 gnd 0.010231f
C5023 vdd.n2381 gnd 0.010231f
C5024 vdd.n2382 gnd 0.008235f
C5025 vdd.n2383 gnd 0.008235f
C5026 vdd.n2384 gnd 0.008235f
C5027 vdd.n2385 gnd 0.010231f
C5028 vdd.n2387 gnd 0.010231f
C5029 vdd.n2388 gnd 0.010231f
C5030 vdd.n2389 gnd 0.008235f
C5031 vdd.n2390 gnd 0.008235f
C5032 vdd.n2391 gnd 0.008235f
C5033 vdd.n2392 gnd 0.010231f
C5034 vdd.n2394 gnd 0.010231f
C5035 vdd.n2395 gnd 0.010231f
C5036 vdd.n2396 gnd 0.008235f
C5037 vdd.n2397 gnd 0.010231f
C5038 vdd.n2398 gnd 0.010231f
C5039 vdd.n2399 gnd 0.010231f
C5040 vdd.n2400 gnd 0.016799f
C5041 vdd.n2401 gnd 0.0056f
C5042 vdd.n2402 gnd 0.008235f
C5043 vdd.n2403 gnd 0.010231f
C5044 vdd.n2405 gnd 0.010231f
C5045 vdd.n2406 gnd 0.010231f
C5046 vdd.n2407 gnd 0.008235f
C5047 vdd.n2408 gnd 0.008235f
C5048 vdd.n2409 gnd 0.008235f
C5049 vdd.n2410 gnd 0.010231f
C5050 vdd.n2412 gnd 0.010231f
C5051 vdd.n2413 gnd 0.010231f
C5052 vdd.n2414 gnd 0.008235f
C5053 vdd.n2415 gnd 0.008235f
C5054 vdd.n2416 gnd 0.008235f
C5055 vdd.n2417 gnd 0.010231f
C5056 vdd.n2419 gnd 0.010231f
C5057 vdd.n2420 gnd 0.010231f
C5058 vdd.n2421 gnd 0.008235f
C5059 vdd.n2422 gnd 0.008235f
C5060 vdd.n2423 gnd 0.008235f
C5061 vdd.n2424 gnd 0.010231f
C5062 vdd.n2426 gnd 0.010231f
C5063 vdd.n2427 gnd 0.010231f
C5064 vdd.n2428 gnd 0.008235f
C5065 vdd.n2429 gnd 0.008235f
C5066 vdd.n2430 gnd 0.008235f
C5067 vdd.n2431 gnd 0.010231f
C5068 vdd.n2433 gnd 0.010231f
C5069 vdd.n2434 gnd 0.010231f
C5070 vdd.n2435 gnd 0.008235f
C5071 vdd.n2436 gnd 0.010231f
C5072 vdd.n2437 gnd 0.010231f
C5073 vdd.n2438 gnd 0.010231f
C5074 vdd.n2439 gnd 0.016799f
C5075 vdd.n2440 gnd 0.006876f
C5076 vdd.n2441 gnd 0.008235f
C5077 vdd.n2442 gnd 0.010231f
C5078 vdd.n2444 gnd 0.010231f
C5079 vdd.n2445 gnd 0.010231f
C5080 vdd.n2446 gnd 0.008235f
C5081 vdd.n2447 gnd 0.008235f
C5082 vdd.n2448 gnd 0.008235f
C5083 vdd.n2449 gnd 0.010231f
C5084 vdd.n2451 gnd 0.010231f
C5085 vdd.n2452 gnd 0.010231f
C5086 vdd.n2453 gnd 0.008235f
C5087 vdd.n2454 gnd 0.008235f
C5088 vdd.n2455 gnd 0.008235f
C5089 vdd.n2456 gnd 0.010231f
C5090 vdd.n2458 gnd 0.010231f
C5091 vdd.n2459 gnd 0.010231f
C5092 vdd.n2460 gnd 0.008235f
C5093 vdd.n2461 gnd 0.008235f
C5094 vdd.n2462 gnd 0.008235f
C5095 vdd.n2463 gnd 0.010231f
C5096 vdd.n2465 gnd 0.010231f
C5097 vdd.n2466 gnd 0.008235f
C5098 vdd.n2467 gnd 0.008235f
C5099 vdd.n2468 gnd 0.010231f
C5100 vdd.n2470 gnd 0.010231f
C5101 vdd.n2471 gnd 0.010231f
C5102 vdd.n2472 gnd 0.008235f
C5103 vdd.n2473 gnd 0.008799f
C5104 vdd.n2474 gnd 1.08617f
C5105 vdd.n2475 gnd 0.046868f
C5106 vdd.n2476 gnd 0.006957f
C5107 vdd.n2477 gnd 0.006957f
C5108 vdd.n2478 gnd 0.006957f
C5109 vdd.n2479 gnd 0.006957f
C5110 vdd.n2480 gnd 0.006957f
C5111 vdd.n2481 gnd 0.006957f
C5112 vdd.n2482 gnd 0.006957f
C5113 vdd.n2483 gnd 0.006957f
C5114 vdd.n2484 gnd 0.006957f
C5115 vdd.n2485 gnd 0.006957f
C5116 vdd.n2486 gnd 0.006957f
C5117 vdd.n2487 gnd 0.006957f
C5118 vdd.n2488 gnd 0.006957f
C5119 vdd.n2489 gnd 0.006957f
C5120 vdd.n2490 gnd 0.006957f
C5121 vdd.n2491 gnd 0.006957f
C5122 vdd.n2492 gnd 0.006957f
C5123 vdd.n2493 gnd 0.006957f
C5124 vdd.n2494 gnd 0.006957f
C5125 vdd.n2495 gnd 0.006957f
C5126 vdd.n2496 gnd 0.006957f
C5127 vdd.n2497 gnd 0.006957f
C5128 vdd.n2498 gnd 0.006957f
C5129 vdd.n2499 gnd 0.006957f
C5130 vdd.n2500 gnd 0.006957f
C5131 vdd.n2501 gnd 0.006957f
C5132 vdd.n2502 gnd 0.006957f
C5133 vdd.n2503 gnd 0.006957f
C5134 vdd.n2504 gnd 0.006957f
C5135 vdd.n2505 gnd 0.006957f
C5136 vdd.n2506 gnd 12.3485f
C5137 vdd.n2508 gnd 0.015797f
C5138 vdd.n2509 gnd 0.015797f
C5139 vdd.n2510 gnd 0.014897f
C5140 vdd.n2511 gnd 0.006957f
C5141 vdd.n2512 gnd 0.006957f
C5142 vdd.n2513 gnd 0.711008f
C5143 vdd.n2514 gnd 0.006957f
C5144 vdd.n2515 gnd 0.006957f
C5145 vdd.n2516 gnd 0.006957f
C5146 vdd.n2517 gnd 0.006957f
C5147 vdd.n2518 gnd 0.006957f
C5148 vdd.n2519 gnd 0.559396f
C5149 vdd.n2520 gnd 0.006957f
C5150 vdd.n2521 gnd 0.006957f
C5151 vdd.n2522 gnd 0.006957f
C5152 vdd.n2523 gnd 0.006957f
C5153 vdd.n2524 gnd 0.006957f
C5154 vdd.n2525 gnd 0.711008f
C5155 vdd.n2526 gnd 0.006957f
C5156 vdd.n2527 gnd 0.006957f
C5157 vdd.n2528 gnd 0.006957f
C5158 vdd.n2529 gnd 0.006957f
C5159 vdd.n2530 gnd 0.006957f
C5160 vdd.n2531 gnd 0.711008f
C5161 vdd.n2532 gnd 0.006957f
C5162 vdd.n2533 gnd 0.006957f
C5163 vdd.n2534 gnd 0.006957f
C5164 vdd.n2535 gnd 0.006957f
C5165 vdd.n2536 gnd 0.006957f
C5166 vdd.n2537 gnd 0.684868f
C5167 vdd.n2538 gnd 0.006957f
C5168 vdd.n2539 gnd 0.006957f
C5169 vdd.n2540 gnd 0.006957f
C5170 vdd.n2541 gnd 0.006957f
C5171 vdd.n2542 gnd 0.006957f
C5172 vdd.n2543 gnd 0.528028f
C5173 vdd.n2544 gnd 0.006957f
C5174 vdd.n2545 gnd 0.006957f
C5175 vdd.n2546 gnd 0.006957f
C5176 vdd.n2547 gnd 0.006957f
C5177 vdd.n2548 gnd 0.006957f
C5178 vdd.n2549 gnd 0.371188f
C5179 vdd.n2550 gnd 0.006957f
C5180 vdd.n2551 gnd 0.006957f
C5181 vdd.n2552 gnd 0.006957f
C5182 vdd.n2553 gnd 0.006957f
C5183 vdd.n2554 gnd 0.006957f
C5184 vdd.n2555 gnd 0.49666f
C5185 vdd.n2556 gnd 0.006957f
C5186 vdd.n2557 gnd 0.006957f
C5187 vdd.n2558 gnd 0.006957f
C5188 vdd.n2559 gnd 0.006957f
C5189 vdd.n2560 gnd 0.006957f
C5190 vdd.n2561 gnd 0.6535f
C5191 vdd.n2562 gnd 0.006957f
C5192 vdd.n2563 gnd 0.006957f
C5193 vdd.n2564 gnd 0.006957f
C5194 vdd.n2565 gnd 0.006957f
C5195 vdd.n2566 gnd 0.006957f
C5196 vdd.n2567 gnd 0.711008f
C5197 vdd.n2568 gnd 0.006957f
C5198 vdd.n2569 gnd 0.006957f
C5199 vdd.n2570 gnd 0.006957f
C5200 vdd.n2571 gnd 0.006957f
C5201 vdd.n2572 gnd 0.006957f
C5202 vdd.n2573 gnd 0.611676f
C5203 vdd.n2574 gnd 0.006957f
C5204 vdd.n2575 gnd 0.006957f
C5205 vdd.n2576 gnd 0.005525f
C5206 vdd.n2577 gnd 0.020155f
C5207 vdd.n2578 gnd 0.004911f
C5208 vdd.n2579 gnd 0.006957f
C5209 vdd.n2580 gnd 0.454836f
C5210 vdd.n2581 gnd 0.006957f
C5211 vdd.n2582 gnd 0.006957f
C5212 vdd.n2583 gnd 0.006957f
C5213 vdd.n2584 gnd 0.006957f
C5214 vdd.n2585 gnd 0.006957f
C5215 vdd.n2586 gnd 0.413012f
C5216 vdd.n2587 gnd 0.006957f
C5217 vdd.n2588 gnd 0.006957f
C5218 vdd.n2589 gnd 0.006957f
C5219 vdd.n2590 gnd 0.006957f
C5220 vdd.n2591 gnd 0.006957f
C5221 vdd.n2592 gnd 0.569852f
C5222 vdd.n2593 gnd 0.006957f
C5223 vdd.n2594 gnd 0.006957f
C5224 vdd.n2595 gnd 0.006957f
C5225 vdd.n2596 gnd 0.006957f
C5226 vdd.n2597 gnd 0.006957f
C5227 vdd.n2598 gnd 0.62736f
C5228 vdd.n2599 gnd 0.006957f
C5229 vdd.n2600 gnd 0.006957f
C5230 vdd.n2601 gnd 0.006957f
C5231 vdd.n2602 gnd 0.006957f
C5232 vdd.n2603 gnd 0.006957f
C5233 vdd.n2604 gnd 0.47052f
C5234 vdd.n2605 gnd 0.006957f
C5235 vdd.n2606 gnd 0.006957f
C5236 vdd.n2607 gnd 0.006957f
C5237 vdd.n2608 gnd 0.006957f
C5238 vdd.n2609 gnd 0.006957f
C5239 vdd.n2610 gnd 0.224804f
C5240 vdd.n2611 gnd 0.006957f
C5241 vdd.n2612 gnd 0.006957f
C5242 vdd.n2613 gnd 0.006957f
C5243 vdd.n2614 gnd 0.006957f
C5244 vdd.n2615 gnd 0.006957f
C5245 vdd.n2616 gnd 0.224804f
C5246 vdd.n2617 gnd 0.006957f
C5247 vdd.n2618 gnd 0.006957f
C5248 vdd.n2619 gnd 0.006957f
C5249 vdd.n2620 gnd 0.006957f
C5250 vdd.n2621 gnd 0.006957f
C5251 vdd.n2622 gnd 0.711008f
C5252 vdd.n2623 gnd 0.006957f
C5253 vdd.n2624 gnd 0.006957f
C5254 vdd.n2625 gnd 0.006957f
C5255 vdd.n2626 gnd 0.006957f
C5256 vdd.n2627 gnd 0.006957f
C5257 vdd.n2628 gnd 0.006957f
C5258 vdd.n2629 gnd 0.006957f
C5259 vdd.n2630 gnd 0.491432f
C5260 vdd.n2631 gnd 0.006957f
C5261 vdd.n2632 gnd 0.006957f
C5262 vdd.n2633 gnd 0.006957f
C5263 vdd.n2634 gnd 0.006957f
C5264 vdd.n2635 gnd 0.006957f
C5265 vdd.n2636 gnd 0.006957f
C5266 vdd.n2637 gnd 0.44438f
C5267 vdd.n2638 gnd 0.006957f
C5268 vdd.n2639 gnd 0.006957f
C5269 vdd.n2640 gnd 0.006957f
C5270 vdd.n2641 gnd 0.015797f
C5271 vdd.n2642 gnd 0.014897f
C5272 vdd.n2643 gnd 0.006957f
C5273 vdd.n2644 gnd 0.006957f
C5274 vdd.n2645 gnd 0.005371f
C5275 vdd.n2646 gnd 0.006957f
C5276 vdd.n2647 gnd 0.006957f
C5277 vdd.n2648 gnd 0.005065f
C5278 vdd.n2649 gnd 0.006957f
C5279 vdd.n2650 gnd 0.006957f
C5280 vdd.n2651 gnd 0.006957f
C5281 vdd.n2652 gnd 0.006957f
C5282 vdd.n2653 gnd 0.006957f
C5283 vdd.n2654 gnd 0.006957f
C5284 vdd.n2655 gnd 0.006957f
C5285 vdd.n2656 gnd 0.006957f
C5286 vdd.n2657 gnd 0.006957f
C5287 vdd.n2658 gnd 0.006957f
C5288 vdd.n2659 gnd 0.006957f
C5289 vdd.n2660 gnd 0.006957f
C5290 vdd.n2661 gnd 0.006957f
C5291 vdd.n2662 gnd 0.006957f
C5292 vdd.n2663 gnd 0.006957f
C5293 vdd.n2664 gnd 0.006957f
C5294 vdd.n2665 gnd 0.006957f
C5295 vdd.n2666 gnd 0.006957f
C5296 vdd.n2667 gnd 0.006957f
C5297 vdd.n2668 gnd 0.006957f
C5298 vdd.n2669 gnd 0.006957f
C5299 vdd.n2670 gnd 0.006957f
C5300 vdd.n2671 gnd 0.006957f
C5301 vdd.n2672 gnd 0.006957f
C5302 vdd.n2673 gnd 0.006957f
C5303 vdd.n2674 gnd 0.006957f
C5304 vdd.n2675 gnd 0.006957f
C5305 vdd.n2676 gnd 0.006957f
C5306 vdd.n2677 gnd 0.006957f
C5307 vdd.n2678 gnd 0.006957f
C5308 vdd.n2679 gnd 0.006957f
C5309 vdd.n2680 gnd 0.006957f
C5310 vdd.n2681 gnd 0.006957f
C5311 vdd.n2682 gnd 0.006957f
C5312 vdd.n2683 gnd 0.006957f
C5313 vdd.n2684 gnd 0.006957f
C5314 vdd.n2685 gnd 0.006957f
C5315 vdd.n2686 gnd 0.006957f
C5316 vdd.n2687 gnd 0.006957f
C5317 vdd.n2688 gnd 0.006957f
C5318 vdd.n2689 gnd 0.006957f
C5319 vdd.n2690 gnd 0.006957f
C5320 vdd.n2691 gnd 0.006957f
C5321 vdd.n2692 gnd 0.006957f
C5322 vdd.n2693 gnd 0.006957f
C5323 vdd.n2694 gnd 0.006957f
C5324 vdd.n2695 gnd 0.006957f
C5325 vdd.n2696 gnd 0.006957f
C5326 vdd.n2697 gnd 0.006957f
C5327 vdd.n2698 gnd 0.006957f
C5328 vdd.n2699 gnd 0.006957f
C5329 vdd.n2700 gnd 0.006957f
C5330 vdd.n2701 gnd 0.006957f
C5331 vdd.n2702 gnd 0.006957f
C5332 vdd.n2703 gnd 0.006957f
C5333 vdd.n2704 gnd 0.006957f
C5334 vdd.n2705 gnd 0.006957f
C5335 vdd.n2706 gnd 0.006957f
C5336 vdd.n2707 gnd 0.006957f
C5337 vdd.n2708 gnd 0.006957f
C5338 vdd.n2709 gnd 0.015797f
C5339 vdd.n2710 gnd 0.014897f
C5340 vdd.n2711 gnd 0.014897f
C5341 vdd.n2712 gnd 0.805111f
C5342 vdd.n2713 gnd 0.014897f
C5343 vdd.n2714 gnd 0.015797f
C5344 vdd.n2715 gnd 0.014897f
C5345 vdd.n2716 gnd 0.006957f
C5346 vdd.n2717 gnd 0.006957f
C5347 vdd.n2718 gnd 0.006957f
C5348 vdd.n2719 gnd 0.005371f
C5349 vdd.n2720 gnd 0.009943f
C5350 vdd.n2721 gnd 0.005065f
C5351 vdd.n2722 gnd 0.006957f
C5352 vdd.n2723 gnd 0.006957f
C5353 vdd.n2724 gnd 0.006957f
C5354 vdd.n2725 gnd 0.006957f
C5355 vdd.n2726 gnd 0.006957f
C5356 vdd.n2727 gnd 0.006957f
C5357 vdd.n2728 gnd 0.006957f
C5358 vdd.n2729 gnd 0.006957f
C5359 vdd.n2730 gnd 0.006957f
C5360 vdd.n2731 gnd 0.006957f
C5361 vdd.n2732 gnd 0.006957f
C5362 vdd.n2733 gnd 0.006957f
C5363 vdd.n2734 gnd 0.006957f
C5364 vdd.n2735 gnd 0.006957f
C5365 vdd.n2736 gnd 0.006957f
C5366 vdd.n2737 gnd 0.006957f
C5367 vdd.n2738 gnd 0.006957f
C5368 vdd.n2739 gnd 0.006957f
C5369 vdd.n2740 gnd 0.006957f
C5370 vdd.n2741 gnd 0.006957f
C5371 vdd.n2742 gnd 0.006957f
C5372 vdd.n2743 gnd 0.006957f
C5373 vdd.n2744 gnd 0.006957f
C5374 vdd.n2745 gnd 0.006957f
C5375 vdd.n2746 gnd 0.006957f
C5376 vdd.n2747 gnd 0.006957f
C5377 vdd.n2748 gnd 0.006957f
C5378 vdd.n2749 gnd 0.006957f
C5379 vdd.n2750 gnd 0.006957f
C5380 vdd.n2751 gnd 0.006957f
C5381 vdd.n2752 gnd 0.006957f
C5382 vdd.n2753 gnd 0.006957f
C5383 vdd.n2754 gnd 0.006957f
C5384 vdd.n2755 gnd 0.006957f
C5385 vdd.n2756 gnd 0.006957f
C5386 vdd.n2757 gnd 0.006957f
C5387 vdd.n2758 gnd 0.006957f
C5388 vdd.n2759 gnd 0.006957f
C5389 vdd.n2760 gnd 0.006957f
C5390 vdd.n2761 gnd 0.006957f
C5391 vdd.n2762 gnd 0.006957f
C5392 vdd.n2763 gnd 0.006957f
C5393 vdd.n2764 gnd 0.006957f
C5394 vdd.n2765 gnd 0.006957f
C5395 vdd.n2766 gnd 0.006957f
C5396 vdd.n2767 gnd 0.006957f
C5397 vdd.n2768 gnd 0.006957f
C5398 vdd.n2769 gnd 0.006957f
C5399 vdd.n2770 gnd 0.006957f
C5400 vdd.n2771 gnd 0.006957f
C5401 vdd.n2772 gnd 0.006957f
C5402 vdd.n2773 gnd 0.006957f
C5403 vdd.n2774 gnd 0.006957f
C5404 vdd.n2775 gnd 0.006957f
C5405 vdd.n2776 gnd 0.006957f
C5406 vdd.n2777 gnd 0.006957f
C5407 vdd.n2778 gnd 0.006957f
C5408 vdd.n2779 gnd 0.006957f
C5409 vdd.n2780 gnd 0.006957f
C5410 vdd.n2781 gnd 0.006957f
C5411 vdd.n2782 gnd 0.015797f
C5412 vdd.n2783 gnd 0.015797f
C5413 vdd.n2784 gnd 0.867847f
C5414 vdd.t251 gnd 3.08452f
C5415 vdd.t238 gnd 3.08452f
C5416 vdd.n2818 gnd 0.015797f
C5417 vdd.t256 gnd 0.606448f
C5418 vdd.n2819 gnd 0.006957f
C5419 vdd.t201 gnd 0.281145f
C5420 vdd.t202 gnd 0.287787f
C5421 vdd.t199 gnd 0.183542f
C5422 vdd.n2820 gnd 0.099195f
C5423 vdd.n2821 gnd 0.056266f
C5424 vdd.n2822 gnd 0.006957f
C5425 vdd.t208 gnd 0.281145f
C5426 vdd.t209 gnd 0.287787f
C5427 vdd.t207 gnd 0.183542f
C5428 vdd.n2823 gnd 0.099195f
C5429 vdd.n2824 gnd 0.056266f
C5430 vdd.n2825 gnd 0.009943f
C5431 vdd.n2826 gnd 0.015797f
C5432 vdd.n2827 gnd 0.015797f
C5433 vdd.n2828 gnd 0.006957f
C5434 vdd.n2829 gnd 0.006957f
C5435 vdd.n2830 gnd 0.006957f
C5436 vdd.n2831 gnd 0.006957f
C5437 vdd.n2832 gnd 0.006957f
C5438 vdd.n2833 gnd 0.006957f
C5439 vdd.n2834 gnd 0.006957f
C5440 vdd.n2835 gnd 0.006957f
C5441 vdd.n2836 gnd 0.006957f
C5442 vdd.n2837 gnd 0.006957f
C5443 vdd.n2838 gnd 0.006957f
C5444 vdd.n2839 gnd 0.006957f
C5445 vdd.n2840 gnd 0.006957f
C5446 vdd.n2841 gnd 0.006957f
C5447 vdd.n2842 gnd 0.006957f
C5448 vdd.n2843 gnd 0.006957f
C5449 vdd.n2844 gnd 0.006957f
C5450 vdd.n2845 gnd 0.006957f
C5451 vdd.n2846 gnd 0.006957f
C5452 vdd.n2847 gnd 0.006957f
C5453 vdd.n2848 gnd 0.006957f
C5454 vdd.n2849 gnd 0.006957f
C5455 vdd.n2850 gnd 0.006957f
C5456 vdd.n2851 gnd 0.006957f
C5457 vdd.n2852 gnd 0.006957f
C5458 vdd.n2853 gnd 0.006957f
C5459 vdd.n2854 gnd 0.006957f
C5460 vdd.n2855 gnd 0.006957f
C5461 vdd.n2856 gnd 0.006957f
C5462 vdd.n2857 gnd 0.006957f
C5463 vdd.n2858 gnd 0.006957f
C5464 vdd.n2859 gnd 0.006957f
C5465 vdd.n2860 gnd 0.006957f
C5466 vdd.n2861 gnd 0.006957f
C5467 vdd.n2862 gnd 0.006957f
C5468 vdd.n2863 gnd 0.006957f
C5469 vdd.n2864 gnd 0.006957f
C5470 vdd.n2865 gnd 0.006957f
C5471 vdd.n2866 gnd 0.006957f
C5472 vdd.n2867 gnd 0.006957f
C5473 vdd.n2868 gnd 0.006957f
C5474 vdd.n2869 gnd 0.006957f
C5475 vdd.n2870 gnd 0.006957f
C5476 vdd.n2871 gnd 0.006957f
C5477 vdd.n2872 gnd 0.006957f
C5478 vdd.n2873 gnd 0.006957f
C5479 vdd.n2874 gnd 0.006957f
C5480 vdd.n2875 gnd 0.006957f
C5481 vdd.n2876 gnd 0.006957f
C5482 vdd.n2877 gnd 0.006957f
C5483 vdd.n2878 gnd 0.006957f
C5484 vdd.n2879 gnd 0.006957f
C5485 vdd.n2880 gnd 0.006957f
C5486 vdd.n2881 gnd 0.006957f
C5487 vdd.n2882 gnd 0.006957f
C5488 vdd.n2883 gnd 0.006957f
C5489 vdd.n2884 gnd 0.006957f
C5490 vdd.n2885 gnd 0.006957f
C5491 vdd.n2886 gnd 0.006957f
C5492 vdd.n2887 gnd 0.006957f
C5493 vdd.n2888 gnd 0.005065f
C5494 vdd.n2889 gnd 0.006957f
C5495 vdd.n2890 gnd 0.006957f
C5496 vdd.n2891 gnd 0.005371f
C5497 vdd.n2892 gnd 0.006957f
C5498 vdd.n2893 gnd 0.006957f
C5499 vdd.n2894 gnd 0.015797f
C5500 vdd.n2895 gnd 0.014897f
C5501 vdd.n2896 gnd 0.014897f
C5502 vdd.n2897 gnd 0.006957f
C5503 vdd.n2898 gnd 0.006957f
C5504 vdd.n2899 gnd 0.006957f
C5505 vdd.n2900 gnd 0.006957f
C5506 vdd.n2901 gnd 0.006957f
C5507 vdd.n2902 gnd 0.006957f
C5508 vdd.n2903 gnd 0.006957f
C5509 vdd.n2904 gnd 0.006957f
C5510 vdd.n2905 gnd 0.006957f
C5511 vdd.n2906 gnd 0.006957f
C5512 vdd.n2907 gnd 0.006957f
C5513 vdd.n2908 gnd 0.006957f
C5514 vdd.n2909 gnd 0.006957f
C5515 vdd.n2910 gnd 0.006957f
C5516 vdd.n2911 gnd 0.006957f
C5517 vdd.n2912 gnd 0.006957f
C5518 vdd.n2913 gnd 0.006957f
C5519 vdd.n2914 gnd 0.006957f
C5520 vdd.n2915 gnd 0.006957f
C5521 vdd.n2916 gnd 0.006957f
C5522 vdd.n2917 gnd 0.006957f
C5523 vdd.n2918 gnd 0.006957f
C5524 vdd.n2919 gnd 0.006957f
C5525 vdd.n2920 gnd 0.006957f
C5526 vdd.n2921 gnd 0.006957f
C5527 vdd.n2922 gnd 0.006957f
C5528 vdd.n2923 gnd 0.006957f
C5529 vdd.n2924 gnd 0.006957f
C5530 vdd.n2925 gnd 0.006957f
C5531 vdd.n2926 gnd 0.006957f
C5532 vdd.n2927 gnd 0.006957f
C5533 vdd.n2928 gnd 0.006957f
C5534 vdd.n2929 gnd 0.006957f
C5535 vdd.n2930 gnd 0.006957f
C5536 vdd.n2931 gnd 0.006957f
C5537 vdd.n2932 gnd 0.006957f
C5538 vdd.n2933 gnd 0.006957f
C5539 vdd.n2934 gnd 0.006957f
C5540 vdd.n2935 gnd 0.006957f
C5541 vdd.n2936 gnd 0.006957f
C5542 vdd.n2937 gnd 0.006957f
C5543 vdd.n2938 gnd 0.006957f
C5544 vdd.n2939 gnd 0.006957f
C5545 vdd.n2940 gnd 0.006957f
C5546 vdd.n2941 gnd 0.006957f
C5547 vdd.n2942 gnd 0.006957f
C5548 vdd.n2943 gnd 0.006957f
C5549 vdd.n2944 gnd 0.006957f
C5550 vdd.n2945 gnd 0.006957f
C5551 vdd.n2946 gnd 0.006957f
C5552 vdd.n2947 gnd 0.006957f
C5553 vdd.n2948 gnd 0.006957f
C5554 vdd.n2949 gnd 0.006957f
C5555 vdd.n2950 gnd 0.006957f
C5556 vdd.n2951 gnd 0.006957f
C5557 vdd.n2952 gnd 0.006957f
C5558 vdd.n2953 gnd 0.006957f
C5559 vdd.n2954 gnd 0.006957f
C5560 vdd.n2955 gnd 0.006957f
C5561 vdd.n2956 gnd 0.006957f
C5562 vdd.n2957 gnd 0.006957f
C5563 vdd.n2958 gnd 0.006957f
C5564 vdd.n2959 gnd 0.006957f
C5565 vdd.n2960 gnd 0.006957f
C5566 vdd.n2961 gnd 0.006957f
C5567 vdd.n2962 gnd 0.006957f
C5568 vdd.n2963 gnd 0.006957f
C5569 vdd.n2964 gnd 0.006957f
C5570 vdd.n2965 gnd 0.006957f
C5571 vdd.n2966 gnd 0.006957f
C5572 vdd.n2967 gnd 0.006957f
C5573 vdd.n2968 gnd 0.006957f
C5574 vdd.n2969 gnd 0.006957f
C5575 vdd.n2970 gnd 0.006957f
C5576 vdd.n2971 gnd 0.006957f
C5577 vdd.n2972 gnd 0.006957f
C5578 vdd.n2973 gnd 0.006957f
C5579 vdd.n2974 gnd 0.006957f
C5580 vdd.n2975 gnd 0.006957f
C5581 vdd.n2976 gnd 0.006957f
C5582 vdd.n2977 gnd 0.006957f
C5583 vdd.n2978 gnd 0.006957f
C5584 vdd.n2979 gnd 0.006957f
C5585 vdd.n2980 gnd 0.006957f
C5586 vdd.n2981 gnd 0.006957f
C5587 vdd.n2982 gnd 0.006957f
C5588 vdd.n2983 gnd 0.006957f
C5589 vdd.n2984 gnd 0.006957f
C5590 vdd.n2985 gnd 0.006957f
C5591 vdd.n2986 gnd 0.006957f
C5592 vdd.n2987 gnd 0.006957f
C5593 vdd.n2988 gnd 0.006957f
C5594 vdd.n2989 gnd 0.006957f
C5595 vdd.n2990 gnd 0.006957f
C5596 vdd.n2991 gnd 0.006957f
C5597 vdd.n2992 gnd 0.006957f
C5598 vdd.n2993 gnd 0.006957f
C5599 vdd.n2994 gnd 0.006957f
C5600 vdd.n2995 gnd 0.006957f
C5601 vdd.n2996 gnd 0.006957f
C5602 vdd.n2997 gnd 0.006957f
C5603 vdd.n2998 gnd 0.224804f
C5604 vdd.n2999 gnd 0.006957f
C5605 vdd.n3000 gnd 0.006957f
C5606 vdd.n3001 gnd 0.006957f
C5607 vdd.n3002 gnd 0.006957f
C5608 vdd.n3003 gnd 0.006957f
C5609 vdd.n3004 gnd 0.224804f
C5610 vdd.n3005 gnd 0.006957f
C5611 vdd.n3006 gnd 0.006957f
C5612 vdd.n3007 gnd 0.006957f
C5613 vdd.n3008 gnd 0.006957f
C5614 vdd.n3009 gnd 0.006957f
C5615 vdd.n3010 gnd 0.006957f
C5616 vdd.n3011 gnd 0.006957f
C5617 vdd.n3012 gnd 0.006957f
C5618 vdd.n3013 gnd 0.006957f
C5619 vdd.n3014 gnd 0.006957f
C5620 vdd.n3015 gnd 0.006957f
C5621 vdd.n3016 gnd 0.44438f
C5622 vdd.n3017 gnd 0.006957f
C5623 vdd.n3018 gnd 0.006957f
C5624 vdd.n3019 gnd 0.006957f
C5625 vdd.n3020 gnd 0.014897f
C5626 vdd.n3021 gnd 0.014897f
C5627 vdd.n3022 gnd 0.015797f
C5628 vdd.n3023 gnd 0.015797f
C5629 vdd.n3024 gnd 0.006957f
C5630 vdd.n3025 gnd 0.006957f
C5631 vdd.n3026 gnd 0.006957f
C5632 vdd.n3027 gnd 0.005371f
C5633 vdd.n3028 gnd 0.009943f
C5634 vdd.n3029 gnd 0.005065f
C5635 vdd.n3030 gnd 0.006957f
C5636 vdd.n3031 gnd 0.006957f
C5637 vdd.n3032 gnd 0.006957f
C5638 vdd.n3033 gnd 0.006957f
C5639 vdd.n3034 gnd 0.006957f
C5640 vdd.n3035 gnd 0.006957f
C5641 vdd.n3036 gnd 0.006957f
C5642 vdd.n3037 gnd 0.006957f
C5643 vdd.n3038 gnd 0.006957f
C5644 vdd.n3039 gnd 0.006957f
C5645 vdd.n3040 gnd 0.006957f
C5646 vdd.n3041 gnd 0.006957f
C5647 vdd.n3042 gnd 0.006957f
C5648 vdd.n3043 gnd 0.006957f
C5649 vdd.n3044 gnd 0.006957f
C5650 vdd.n3045 gnd 0.006957f
C5651 vdd.n3046 gnd 0.006957f
C5652 vdd.n3047 gnd 0.006957f
C5653 vdd.n3048 gnd 0.006957f
C5654 vdd.n3049 gnd 0.006957f
C5655 vdd.n3050 gnd 0.006957f
C5656 vdd.n3051 gnd 0.006957f
C5657 vdd.n3052 gnd 0.006957f
C5658 vdd.n3053 gnd 0.006957f
C5659 vdd.n3054 gnd 0.006957f
C5660 vdd.n3055 gnd 0.006957f
C5661 vdd.n3056 gnd 0.006957f
C5662 vdd.n3057 gnd 0.006957f
C5663 vdd.n3058 gnd 0.006957f
C5664 vdd.n3059 gnd 0.006957f
C5665 vdd.n3060 gnd 0.006957f
C5666 vdd.n3061 gnd 0.006957f
C5667 vdd.n3062 gnd 0.006957f
C5668 vdd.n3063 gnd 0.006957f
C5669 vdd.n3064 gnd 0.006957f
C5670 vdd.n3065 gnd 0.006957f
C5671 vdd.n3066 gnd 0.006957f
C5672 vdd.n3067 gnd 0.006957f
C5673 vdd.n3068 gnd 0.006957f
C5674 vdd.n3069 gnd 0.006957f
C5675 vdd.n3070 gnd 0.006957f
C5676 vdd.n3071 gnd 0.006957f
C5677 vdd.n3072 gnd 0.006957f
C5678 vdd.n3073 gnd 0.006957f
C5679 vdd.n3074 gnd 0.006957f
C5680 vdd.n3075 gnd 0.006957f
C5681 vdd.n3076 gnd 0.006957f
C5682 vdd.n3077 gnd 0.006957f
C5683 vdd.n3078 gnd 0.006957f
C5684 vdd.n3079 gnd 0.006957f
C5685 vdd.n3080 gnd 0.006957f
C5686 vdd.n3081 gnd 0.006957f
C5687 vdd.n3082 gnd 0.006957f
C5688 vdd.n3083 gnd 0.006957f
C5689 vdd.n3084 gnd 0.006957f
C5690 vdd.n3085 gnd 0.006957f
C5691 vdd.n3086 gnd 0.006957f
C5692 vdd.n3087 gnd 0.006957f
C5693 vdd.n3088 gnd 0.867847f
C5694 vdd.n3090 gnd 0.015797f
C5695 vdd.n3091 gnd 0.015797f
C5696 vdd.n3092 gnd 0.014897f
C5697 vdd.n3093 gnd 0.006957f
C5698 vdd.n3094 gnd 0.006957f
C5699 vdd.n3095 gnd 0.41824f
C5700 vdd.n3096 gnd 0.006957f
C5701 vdd.n3097 gnd 0.006957f
C5702 vdd.n3098 gnd 0.006957f
C5703 vdd.n3099 gnd 0.006957f
C5704 vdd.n3100 gnd 0.006957f
C5705 vdd.n3101 gnd 0.423468f
C5706 vdd.n3102 gnd 0.006957f
C5707 vdd.n3103 gnd 0.006957f
C5708 vdd.n3104 gnd 0.006957f
C5709 vdd.n3105 gnd 0.006957f
C5710 vdd.n3106 gnd 0.006957f
C5711 vdd.n3107 gnd 0.711008f
C5712 vdd.n3108 gnd 0.006957f
C5713 vdd.n3109 gnd 0.006957f
C5714 vdd.n3110 gnd 0.006957f
C5715 vdd.n3111 gnd 0.006957f
C5716 vdd.n3112 gnd 0.006957f
C5717 vdd.n3113 gnd 0.512344f
C5718 vdd.n3114 gnd 0.006957f
C5719 vdd.n3115 gnd 0.006957f
C5720 vdd.n3116 gnd 0.006957f
C5721 vdd.n3117 gnd 0.006957f
C5722 vdd.n3118 gnd 0.006957f
C5723 vdd.n3119 gnd 0.643044f
C5724 vdd.n3120 gnd 0.006957f
C5725 vdd.n3121 gnd 0.006957f
C5726 vdd.n3122 gnd 0.006957f
C5727 vdd.n3123 gnd 0.006957f
C5728 vdd.n3124 gnd 0.006957f
C5729 vdd.n3125 gnd 0.528028f
C5730 vdd.n3126 gnd 0.006957f
C5731 vdd.n3127 gnd 0.006957f
C5732 vdd.n3128 gnd 0.006957f
C5733 vdd.n3129 gnd 0.006957f
C5734 vdd.n3130 gnd 0.006957f
C5735 vdd.n3131 gnd 0.371188f
C5736 vdd.n3132 gnd 0.006957f
C5737 vdd.n3133 gnd 0.006957f
C5738 vdd.n3134 gnd 0.006957f
C5739 vdd.n3135 gnd 0.006957f
C5740 vdd.n3136 gnd 0.006957f
C5741 vdd.n3137 gnd 0.224804f
C5742 vdd.n3138 gnd 0.006957f
C5743 vdd.n3139 gnd 0.006957f
C5744 vdd.n3140 gnd 0.006957f
C5745 vdd.n3141 gnd 0.006957f
C5746 vdd.n3142 gnd 0.006957f
C5747 vdd.n3143 gnd 0.6535f
C5748 vdd.n3144 gnd 0.006957f
C5749 vdd.n3145 gnd 0.006957f
C5750 vdd.n3146 gnd 0.006957f
C5751 vdd.n3147 gnd 0.004911f
C5752 vdd.n3148 gnd 0.006957f
C5753 vdd.n3149 gnd 0.006957f
C5754 vdd.n3150 gnd 0.711008f
C5755 vdd.n3151 gnd 0.006957f
C5756 vdd.n3152 gnd 0.006957f
C5757 vdd.n3153 gnd 0.006957f
C5758 vdd.n3154 gnd 0.006957f
C5759 vdd.n3155 gnd 0.006957f
C5760 vdd.n3156 gnd 0.564624f
C5761 vdd.n3157 gnd 0.006957f
C5762 vdd.n3158 gnd 0.005525f
C5763 vdd.n3159 gnd 0.006957f
C5764 vdd.n3160 gnd 0.006957f
C5765 vdd.n3161 gnd 0.006957f
C5766 vdd.n3162 gnd 0.454836f
C5767 vdd.n3163 gnd 0.006957f
C5768 vdd.n3164 gnd 0.006957f
C5769 vdd.n3165 gnd 0.006957f
C5770 vdd.n3166 gnd 0.006957f
C5771 vdd.n3167 gnd 0.006957f
C5772 vdd.n3168 gnd 0.413012f
C5773 vdd.n3169 gnd 0.006957f
C5774 vdd.n3170 gnd 0.006957f
C5775 vdd.n3171 gnd 0.006957f
C5776 vdd.n3172 gnd 0.006957f
C5777 vdd.n3173 gnd 0.006957f
C5778 vdd.n3174 gnd 0.569852f
C5779 vdd.n3175 gnd 0.006957f
C5780 vdd.n3176 gnd 0.006957f
C5781 vdd.n3177 gnd 0.006957f
C5782 vdd.n3178 gnd 0.006957f
C5783 vdd.n3179 gnd 0.006957f
C5784 vdd.n3180 gnd 0.711008f
C5785 vdd.n3181 gnd 0.006957f
C5786 vdd.n3182 gnd 0.006957f
C5787 vdd.n3183 gnd 0.006957f
C5788 vdd.n3184 gnd 0.006957f
C5789 vdd.n3185 gnd 0.006957f
C5790 vdd.n3186 gnd 0.695324f
C5791 vdd.n3187 gnd 0.006957f
C5792 vdd.n3188 gnd 0.006957f
C5793 vdd.n3189 gnd 0.006957f
C5794 vdd.n3190 gnd 0.006957f
C5795 vdd.n3191 gnd 0.006957f
C5796 vdd.n3192 gnd 0.538484f
C5797 vdd.n3193 gnd 0.006957f
C5798 vdd.n3194 gnd 0.006957f
C5799 vdd.n3195 gnd 0.006957f
C5800 vdd.n3196 gnd 0.006957f
C5801 vdd.n3197 gnd 0.006957f
C5802 vdd.n3198 gnd 0.381644f
C5803 vdd.n3199 gnd 0.006957f
C5804 vdd.n3200 gnd 0.006957f
C5805 vdd.n3201 gnd 0.006957f
C5806 vdd.n3202 gnd 0.006957f
C5807 vdd.n3203 gnd 0.006957f
C5808 vdd.n3204 gnd 0.711008f
C5809 vdd.n3205 gnd 0.006957f
C5810 vdd.n3206 gnd 0.006957f
C5811 vdd.n3207 gnd 0.006957f
C5812 vdd.n3208 gnd 0.006957f
C5813 vdd.n3209 gnd 0.006957f
C5814 vdd.n3210 gnd 0.006957f
C5815 vdd.n3212 gnd 0.006957f
C5816 vdd.n3213 gnd 0.006957f
C5817 vdd.n3215 gnd 0.006957f
C5818 vdd.n3216 gnd 0.006957f
C5819 vdd.n3219 gnd 0.006957f
C5820 vdd.n3220 gnd 0.006957f
C5821 vdd.n3221 gnd 0.006957f
C5822 vdd.n3222 gnd 0.006957f
C5823 vdd.n3224 gnd 0.006957f
C5824 vdd.n3225 gnd 0.006957f
C5825 vdd.n3226 gnd 0.006957f
C5826 vdd.n3227 gnd 0.006957f
C5827 vdd.n3228 gnd 0.006957f
C5828 vdd.n3229 gnd 0.006957f
C5829 vdd.n3231 gnd 0.006957f
C5830 vdd.n3232 gnd 0.006957f
C5831 vdd.n3233 gnd 0.006957f
C5832 vdd.n3234 gnd 0.006957f
C5833 vdd.n3235 gnd 0.006957f
C5834 vdd.n3236 gnd 0.006957f
C5835 vdd.n3238 gnd 0.006957f
C5836 vdd.n3239 gnd 0.006957f
C5837 vdd.n3240 gnd 0.006957f
C5838 vdd.n3241 gnd 0.006957f
C5839 vdd.n3242 gnd 0.006957f
C5840 vdd.n3243 gnd 0.006957f
C5841 vdd.n3245 gnd 0.006957f
C5842 vdd.n3246 gnd 0.015797f
C5843 vdd.n3247 gnd 0.015797f
C5844 vdd.n3248 gnd 0.014897f
C5845 vdd.n3249 gnd 0.006957f
C5846 vdd.n3250 gnd 0.006957f
C5847 vdd.n3251 gnd 0.006957f
C5848 vdd.n3252 gnd 0.006957f
C5849 vdd.n3253 gnd 0.006957f
C5850 vdd.n3254 gnd 0.006957f
C5851 vdd.n3255 gnd 0.711008f
C5852 vdd.n3256 gnd 0.006957f
C5853 vdd.n3257 gnd 0.006957f
C5854 vdd.n3258 gnd 0.006957f
C5855 vdd.n3259 gnd 0.006957f
C5856 vdd.n3260 gnd 0.006957f
C5857 vdd.n3261 gnd 0.507116f
C5858 vdd.n3262 gnd 0.006957f
C5859 vdd.n3263 gnd 0.006957f
C5860 vdd.n3264 gnd 0.006957f
C5861 vdd.n3265 gnd 0.015797f
C5862 vdd.n3266 gnd 0.014897f
C5863 vdd.n3267 gnd 0.015797f
C5864 vdd.n3269 gnd 0.006957f
C5865 vdd.n3270 gnd 0.006957f
C5866 vdd.n3271 gnd 0.005371f
C5867 vdd.n3272 gnd 0.009943f
C5868 vdd.n3273 gnd 0.005065f
C5869 vdd.n3274 gnd 0.006957f
C5870 vdd.n3275 gnd 0.006957f
C5871 vdd.n3277 gnd 0.006957f
C5872 vdd.n3278 gnd 0.006957f
C5873 vdd.n3279 gnd 0.006957f
C5874 vdd.n3280 gnd 0.006957f
C5875 vdd.n3281 gnd 0.006957f
C5876 vdd.n3282 gnd 0.006957f
C5877 vdd.n3284 gnd 0.006957f
C5878 vdd.n3285 gnd 0.006957f
C5879 vdd.n3286 gnd 0.006957f
C5880 vdd.n3287 gnd 0.006957f
C5881 vdd.n3288 gnd 0.006957f
C5882 vdd.n3289 gnd 0.006957f
C5883 vdd.n3291 gnd 0.006957f
C5884 vdd.n3292 gnd 0.006957f
C5885 vdd.n3293 gnd 0.006957f
C5886 vdd.n3294 gnd 0.006957f
C5887 vdd.n3295 gnd 0.006957f
C5888 vdd.n3296 gnd 0.006957f
C5889 vdd.n3298 gnd 0.006957f
C5890 vdd.n3299 gnd 0.006957f
C5891 vdd.n3300 gnd 0.006957f
C5892 vdd.n3302 gnd 0.006957f
C5893 vdd.n3303 gnd 0.006957f
C5894 vdd.n3304 gnd 0.006957f
C5895 vdd.n3305 gnd 0.006957f
C5896 vdd.n3306 gnd 0.006957f
C5897 vdd.n3307 gnd 0.006957f
C5898 vdd.n3309 gnd 0.006957f
C5899 vdd.n3310 gnd 0.006957f
C5900 vdd.n3311 gnd 0.006957f
C5901 vdd.n3312 gnd 0.006957f
C5902 vdd.n3313 gnd 0.006957f
C5903 vdd.n3314 gnd 0.006957f
C5904 vdd.n3316 gnd 0.006957f
C5905 vdd.n3317 gnd 0.006957f
C5906 vdd.n3318 gnd 0.006957f
C5907 vdd.n3319 gnd 0.006957f
C5908 vdd.n3320 gnd 0.006957f
C5909 vdd.n3321 gnd 0.006957f
C5910 vdd.n3323 gnd 0.006957f
C5911 vdd.n3324 gnd 0.006957f
C5912 vdd.n3326 gnd 0.006957f
C5913 vdd.n3327 gnd 0.006957f
C5914 vdd.n3328 gnd 0.015797f
C5915 vdd.n3329 gnd 0.014897f
C5916 vdd.n3330 gnd 0.014897f
C5917 vdd.n3331 gnd 0.961951f
C5918 vdd.n3332 gnd 0.014897f
C5919 vdd.n3333 gnd 0.015797f
C5920 vdd.n3334 gnd 0.014897f
C5921 vdd.n3335 gnd 0.006957f
C5922 vdd.n3336 gnd 0.005371f
C5923 vdd.n3337 gnd 0.006957f
C5924 vdd.n3339 gnd 0.006957f
C5925 vdd.n3340 gnd 0.006957f
C5926 vdd.n3341 gnd 0.006957f
C5927 vdd.n3342 gnd 0.006957f
C5928 vdd.n3343 gnd 0.006957f
C5929 vdd.n3344 gnd 0.006957f
C5930 vdd.n3346 gnd 0.006957f
C5931 vdd.n3347 gnd 0.006957f
C5932 vdd.n3348 gnd 0.006957f
C5933 vdd.n3349 gnd 0.006957f
C5934 vdd.n3350 gnd 0.006957f
C5935 vdd.n3351 gnd 0.006957f
C5936 vdd.n3353 gnd 0.006957f
C5937 vdd.n3354 gnd 0.006957f
C5938 vdd.n3355 gnd 0.006957f
C5939 vdd.n3356 gnd 0.006957f
C5940 vdd.n3357 gnd 0.006957f
C5941 vdd.n3358 gnd 0.006957f
C5942 vdd.n3360 gnd 0.006957f
C5943 vdd.n3361 gnd 0.006957f
C5944 vdd.n3363 gnd 0.006957f
C5945 vdd.n3364 gnd 0.042961f
C5946 vdd.n3365 gnd 1.09007f
C5947 vdd.n3367 gnd 0.004323f
C5948 vdd.n3368 gnd 0.008235f
C5949 vdd.n3369 gnd 0.010231f
C5950 vdd.n3370 gnd 0.010231f
C5951 vdd.n3371 gnd 0.008235f
C5952 vdd.n3372 gnd 0.008235f
C5953 vdd.n3373 gnd 0.010231f
C5954 vdd.n3374 gnd 0.010231f
C5955 vdd.n3375 gnd 0.008235f
C5956 vdd.n3376 gnd 0.008235f
C5957 vdd.n3377 gnd 0.010231f
C5958 vdd.n3378 gnd 0.010231f
C5959 vdd.n3379 gnd 0.008235f
C5960 vdd.n3380 gnd 0.008235f
C5961 vdd.n3381 gnd 0.010231f
C5962 vdd.n3382 gnd 0.010231f
C5963 vdd.n3383 gnd 0.008235f
C5964 vdd.n3384 gnd 0.008235f
C5965 vdd.n3385 gnd 0.010231f
C5966 vdd.n3386 gnd 0.010231f
C5967 vdd.n3387 gnd 0.008235f
C5968 vdd.n3388 gnd 0.008235f
C5969 vdd.n3389 gnd 0.010231f
C5970 vdd.n3390 gnd 0.010231f
C5971 vdd.n3391 gnd 0.008235f
C5972 vdd.n3392 gnd 0.008235f
C5973 vdd.n3393 gnd 0.010231f
C5974 vdd.n3394 gnd 0.010231f
C5975 vdd.n3395 gnd 0.008235f
C5976 vdd.n3396 gnd 0.008235f
C5977 vdd.n3397 gnd 0.010231f
C5978 vdd.n3398 gnd 0.010231f
C5979 vdd.n3399 gnd 0.008235f
C5980 vdd.n3400 gnd 0.008235f
C5981 vdd.n3401 gnd 0.010231f
C5982 vdd.n3402 gnd 0.010231f
C5983 vdd.n3403 gnd 0.008235f
C5984 vdd.n3404 gnd 0.010231f
C5985 vdd.n3405 gnd 0.010231f
C5986 vdd.n3406 gnd 0.008235f
C5987 vdd.n3407 gnd 0.010231f
C5988 vdd.n3408 gnd 0.010231f
C5989 vdd.n3409 gnd 0.010231f
C5990 vdd.n3410 gnd 0.016799f
C5991 vdd.n3411 gnd 0.010231f
C5992 vdd.n3412 gnd 0.010231f
C5993 vdd.n3413 gnd 0.0056f
C5994 vdd.n3414 gnd 0.008235f
C5995 vdd.n3415 gnd 0.010231f
C5996 vdd.n3416 gnd 0.010231f
C5997 vdd.n3417 gnd 0.008235f
C5998 vdd.n3418 gnd 0.008235f
C5999 vdd.n3419 gnd 0.010231f
C6000 vdd.n3420 gnd 0.010231f
C6001 vdd.n3421 gnd 0.008235f
C6002 vdd.n3422 gnd 0.008235f
C6003 vdd.n3423 gnd 0.010231f
C6004 vdd.n3424 gnd 0.010231f
C6005 vdd.n3425 gnd 0.008235f
C6006 vdd.n3426 gnd 0.008235f
C6007 vdd.n3427 gnd 0.010231f
C6008 vdd.n3428 gnd 0.010231f
C6009 vdd.n3429 gnd 0.008235f
C6010 vdd.n3430 gnd 0.008235f
C6011 vdd.n3431 gnd 0.010231f
C6012 vdd.n3432 gnd 0.010231f
C6013 vdd.n3433 gnd 0.008235f
C6014 vdd.n3434 gnd 0.008235f
C6015 vdd.n3435 gnd 0.010231f
C6016 vdd.n3436 gnd 0.010231f
C6017 vdd.n3437 gnd 0.008235f
C6018 vdd.n3438 gnd 0.008235f
C6019 vdd.n3439 gnd 0.010231f
C6020 vdd.n3440 gnd 0.010231f
C6021 vdd.n3441 gnd 0.008235f
C6022 vdd.n3442 gnd 0.008235f
C6023 vdd.n3443 gnd 0.010231f
C6024 vdd.n3444 gnd 0.010231f
C6025 vdd.n3445 gnd 0.008235f
C6026 vdd.n3446 gnd 0.008235f
C6027 vdd.n3447 gnd 0.010231f
C6028 vdd.n3448 gnd 0.010231f
C6029 vdd.n3449 gnd 0.008235f
C6030 vdd.n3450 gnd 0.010231f
C6031 vdd.n3451 gnd 0.010231f
C6032 vdd.n3452 gnd 0.008235f
C6033 vdd.n3453 gnd 0.010231f
C6034 vdd.n3454 gnd 0.010231f
C6035 vdd.n3455 gnd 0.010231f
C6036 vdd.t197 gnd 0.125873f
C6037 vdd.t198 gnd 0.134524f
C6038 vdd.t196 gnd 0.164388f
C6039 vdd.n3456 gnd 0.210723f
C6040 vdd.n3457 gnd 0.177045f
C6041 vdd.n3458 gnd 0.016799f
C6042 vdd.n3459 gnd 0.010231f
C6043 vdd.n3460 gnd 0.010231f
C6044 vdd.n3461 gnd 0.006876f
C6045 vdd.n3462 gnd 0.008235f
C6046 vdd.n3463 gnd 0.010231f
C6047 vdd.n3464 gnd 0.010231f
C6048 vdd.n3465 gnd 0.008235f
C6049 vdd.n3466 gnd 0.008235f
C6050 vdd.n3467 gnd 0.010231f
C6051 vdd.n3468 gnd 0.010231f
C6052 vdd.n3469 gnd 0.008235f
C6053 vdd.n3470 gnd 0.008235f
C6054 vdd.n3471 gnd 0.010231f
C6055 vdd.n3472 gnd 0.010231f
C6056 vdd.n3473 gnd 0.008235f
C6057 vdd.n3474 gnd 0.008235f
C6058 vdd.n3475 gnd 0.010231f
C6059 vdd.n3476 gnd 0.010231f
C6060 vdd.n3477 gnd 0.008235f
C6061 vdd.n3478 gnd 0.008235f
C6062 vdd.n3479 gnd 0.010231f
C6063 vdd.n3480 gnd 0.010231f
C6064 vdd.n3481 gnd 0.008235f
C6065 vdd.n3482 gnd 0.008235f
C6066 vdd.n3483 gnd 0.010231f
C6067 vdd.n3484 gnd 0.010231f
C6068 vdd.n3485 gnd 0.008235f
C6069 vdd.n3486 gnd 0.008235f
C6070 vdd.n3488 gnd 1.09007f
C6071 vdd.n3490 gnd 0.008235f
C6072 vdd.n3491 gnd 0.008235f
C6073 vdd.n3492 gnd 0.006835f
C6074 vdd.n3493 gnd 0.025281f
C6075 vdd.n3495 gnd 12.7668f
C6076 vdd.n3496 gnd 0.025281f
C6077 vdd.n3497 gnd 0.003912f
C6078 vdd.n3498 gnd 0.025281f
C6079 vdd.n3499 gnd 0.024751f
C6080 vdd.n3500 gnd 0.010231f
C6081 vdd.n3501 gnd 0.008235f
C6082 vdd.n3502 gnd 0.010231f
C6083 vdd.n3503 gnd 0.632588f
C6084 vdd.n3504 gnd 0.010231f
C6085 vdd.n3505 gnd 0.008235f
C6086 vdd.n3506 gnd 0.010231f
C6087 vdd.n3507 gnd 0.010231f
C6088 vdd.n3508 gnd 0.010231f
C6089 vdd.n3509 gnd 0.008235f
C6090 vdd.n3510 gnd 0.010231f
C6091 vdd.n3511 gnd 1.0456f
C6092 vdd.n3512 gnd 0.010231f
C6093 vdd.n3513 gnd 0.008235f
C6094 vdd.n3514 gnd 0.010231f
C6095 vdd.n3515 gnd 0.010231f
C6096 vdd.n3516 gnd 0.010231f
C6097 vdd.n3517 gnd 0.008235f
C6098 vdd.n3518 gnd 0.010231f
C6099 vdd.n3519 gnd 0.674412f
C6100 vdd.n3520 gnd 0.716236f
C6101 vdd.n3521 gnd 0.010231f
C6102 vdd.n3522 gnd 0.008235f
C6103 vdd.n3523 gnd 0.010231f
C6104 vdd.n3524 gnd 0.010231f
C6105 vdd.n3525 gnd 0.010231f
C6106 vdd.n3526 gnd 0.008235f
C6107 vdd.n3527 gnd 0.010231f
C6108 vdd.n3528 gnd 0.867847f
C6109 vdd.n3529 gnd 0.010231f
C6110 vdd.n3530 gnd 0.008235f
C6111 vdd.n3531 gnd 0.010231f
C6112 vdd.n3532 gnd 0.010231f
C6113 vdd.n3533 gnd 0.010231f
C6114 vdd.n3534 gnd 0.008235f
C6115 vdd.n3535 gnd 0.010231f
C6116 vdd.t2 gnd 0.5228f
C6117 vdd.n3536 gnd 0.841707f
C6118 vdd.n3537 gnd 0.010231f
C6119 vdd.n3538 gnd 0.008235f
C6120 vdd.n3539 gnd 0.010231f
C6121 vdd.n3540 gnd 0.010231f
C6122 vdd.n3541 gnd 0.010231f
C6123 vdd.n3542 gnd 0.008235f
C6124 vdd.n3543 gnd 0.010231f
C6125 vdd.n3544 gnd 0.663956f
C6126 vdd.n3545 gnd 0.010231f
C6127 vdd.n3546 gnd 0.008235f
C6128 vdd.n3547 gnd 0.010231f
C6129 vdd.n3548 gnd 0.010231f
C6130 vdd.n3549 gnd 0.010231f
C6131 vdd.n3550 gnd 0.008235f
C6132 vdd.n3551 gnd 0.010231f
C6133 vdd.n3552 gnd 0.831251f
C6134 vdd.n3553 gnd 0.559396f
C6135 vdd.n3554 gnd 0.010231f
C6136 vdd.n3555 gnd 0.008235f
C6137 vdd.n3556 gnd 0.010231f
C6138 vdd.n3557 gnd 0.010231f
C6139 vdd.n3558 gnd 0.010231f
C6140 vdd.n3559 gnd 0.008235f
C6141 vdd.n3560 gnd 0.010231f
C6142 vdd.n3561 gnd 0.737148f
C6143 vdd.n3562 gnd 0.010231f
C6144 vdd.n3563 gnd 0.008235f
C6145 vdd.n3564 gnd 0.010231f
C6146 vdd.n3565 gnd 0.010231f
C6147 vdd.n3566 gnd 0.010231f
C6148 vdd.n3567 gnd 0.010231f
C6149 vdd.n3568 gnd 0.010231f
C6150 vdd.n3569 gnd 0.008235f
C6151 vdd.n3570 gnd 0.008235f
C6152 vdd.n3571 gnd 0.010231f
C6153 vdd.t119 gnd 0.5228f
C6154 vdd.n3572 gnd 0.867847f
C6155 vdd.n3573 gnd 0.010231f
C6156 vdd.n3574 gnd 0.008235f
C6157 vdd.n3575 gnd 0.010231f
C6158 vdd.n3576 gnd 0.010231f
C6159 vdd.n3577 gnd 0.010231f
C6160 vdd.n3578 gnd 0.008235f
C6161 vdd.n3579 gnd 0.010231f
C6162 vdd.n3580 gnd 0.820795f
C6163 vdd.n3581 gnd 0.010231f
C6164 vdd.n3582 gnd 0.010231f
C6165 vdd.n3583 gnd 0.008235f
C6166 vdd.n3584 gnd 0.008235f
C6167 vdd.n3585 gnd 0.010231f
C6168 vdd.n3586 gnd 0.010231f
C6169 vdd.n3587 gnd 0.010231f
C6170 vdd.n3588 gnd 0.008235f
C6171 vdd.n3589 gnd 0.010231f
C6172 vdd.n3590 gnd 0.008235f
C6173 vdd.n3591 gnd 0.008235f
C6174 vdd.n3592 gnd 0.010231f
C6175 vdd.n3593 gnd 0.010231f
C6176 vdd.n3594 gnd 0.010231f
C6177 vdd.n3595 gnd 0.008235f
C6178 vdd.n3596 gnd 0.010231f
C6179 vdd.n3597 gnd 0.008235f
C6180 vdd.n3598 gnd 0.008235f
C6181 vdd.n3599 gnd 0.010231f
C6182 vdd.n3600 gnd 0.010231f
C6183 vdd.n3601 gnd 0.010231f
C6184 vdd.n3602 gnd 0.008235f
C6185 vdd.n3603 gnd 0.867847f
C6186 vdd.n3604 gnd 0.010231f
C6187 vdd.n3605 gnd 0.008235f
C6188 vdd.n3606 gnd 0.008235f
C6189 vdd.n3607 gnd 0.010231f
C6190 vdd.n3608 gnd 0.010231f
C6191 vdd.n3609 gnd 0.010231f
C6192 vdd.n3610 gnd 0.008235f
C6193 vdd.n3611 gnd 0.010231f
C6194 vdd.n3612 gnd 0.008235f
C6195 vdd.n3613 gnd 0.008235f
C6196 vdd.n3614 gnd 0.010231f
C6197 vdd.n3615 gnd 0.010231f
C6198 vdd.n3616 gnd 0.010231f
C6199 vdd.n3617 gnd 0.008235f
C6200 vdd.n3618 gnd 0.010231f
C6201 vdd.n3619 gnd 0.008235f
C6202 vdd.n3620 gnd 0.006835f
C6203 vdd.n3621 gnd 0.024751f
C6204 vdd.n3622 gnd 0.025281f
C6205 vdd.n3623 gnd 0.003912f
C6206 vdd.n3624 gnd 0.025281f
C6207 vdd.n3626 gnd 2.47807f
C6208 vdd.n3627 gnd 1.54226f
C6209 vdd.n3628 gnd 0.024751f
C6210 vdd.n3629 gnd 0.006835f
C6211 vdd.n3630 gnd 0.008235f
C6212 vdd.n3631 gnd 0.008235f
C6213 vdd.n3632 gnd 0.010231f
C6214 vdd.n3633 gnd 1.0456f
C6215 vdd.n3634 gnd 1.0456f
C6216 vdd.n3635 gnd 0.956723f
C6217 vdd.n3636 gnd 0.010231f
C6218 vdd.n3637 gnd 0.008235f
C6219 vdd.n3638 gnd 0.008235f
C6220 vdd.n3639 gnd 0.008235f
C6221 vdd.n3640 gnd 0.010231f
C6222 vdd.n3641 gnd 0.778971f
C6223 vdd.t117 gnd 0.5228f
C6224 vdd.n3642 gnd 0.789427f
C6225 vdd.n3643 gnd 0.60122f
C6226 vdd.n3644 gnd 0.010231f
C6227 vdd.n3645 gnd 0.008235f
C6228 vdd.n3646 gnd 0.008235f
C6229 vdd.n3647 gnd 0.008235f
C6230 vdd.n3648 gnd 0.010231f
C6231 vdd.n3649 gnd 0.622132f
C6232 vdd.n3650 gnd 0.768516f
C6233 vdd.t31 gnd 0.5228f
C6234 vdd.n3651 gnd 0.799883f
C6235 vdd.n3652 gnd 0.010231f
C6236 vdd.n3653 gnd 0.008235f
C6237 vdd.n3654 gnd 0.008235f
C6238 vdd.n3655 gnd 0.008235f
C6239 vdd.n3656 gnd 0.010231f
C6240 vdd.n3657 gnd 0.867847f
C6241 vdd.t43 gnd 0.5228f
C6242 vdd.n3658 gnd 0.632588f
C6243 vdd.n3659 gnd 0.75806f
C6244 vdd.n3660 gnd 0.010231f
C6245 vdd.n3661 gnd 0.008235f
C6246 vdd.n3662 gnd 0.008235f
C6247 vdd.n3663 gnd 0.008235f
C6248 vdd.n3664 gnd 0.010231f
C6249 vdd.n3665 gnd 0.580308f
C6250 vdd.t33 gnd 0.5228f
C6251 vdd.n3666 gnd 0.867847f
C6252 vdd.t46 gnd 0.5228f
C6253 vdd.n3667 gnd 0.643044f
C6254 vdd.n3668 gnd 0.010231f
C6255 vdd.n3669 gnd 0.008235f
C6256 vdd.n3670 gnd 0.007863f
C6257 vdd.n3671 gnd 0.603486f
C6258 vdd.n3672 gnd 2.98812f
C6259 a_n2804_13878.t29 gnd 0.194556f
C6260 a_n2804_13878.t25 gnd 0.194556f
C6261 a_n2804_13878.t31 gnd 0.194556f
C6262 a_n2804_13878.n0 gnd 1.53449f
C6263 a_n2804_13878.t8 gnd 0.194556f
C6264 a_n2804_13878.t20 gnd 0.194556f
C6265 a_n2804_13878.n1 gnd 1.53196f
C6266 a_n2804_13878.n2 gnd 1.37704f
C6267 a_n2804_13878.t12 gnd 0.194556f
C6268 a_n2804_13878.t22 gnd 0.194556f
C6269 a_n2804_13878.n3 gnd 1.53358f
C6270 a_n2804_13878.t27 gnd 0.194556f
C6271 a_n2804_13878.t17 gnd 0.194556f
C6272 a_n2804_13878.n4 gnd 1.53196f
C6273 a_n2804_13878.n5 gnd 2.14061f
C6274 a_n2804_13878.t23 gnd 0.194556f
C6275 a_n2804_13878.t16 gnd 0.194556f
C6276 a_n2804_13878.n6 gnd 1.53196f
C6277 a_n2804_13878.n7 gnd 1.04414f
C6278 a_n2804_13878.t10 gnd 0.194556f
C6279 a_n2804_13878.t13 gnd 0.194556f
C6280 a_n2804_13878.n8 gnd 1.53196f
C6281 a_n2804_13878.n9 gnd 1.04414f
C6282 a_n2804_13878.t26 gnd 0.194556f
C6283 a_n2804_13878.t11 gnd 0.194556f
C6284 a_n2804_13878.n10 gnd 1.53196f
C6285 a_n2804_13878.n11 gnd 1.04414f
C6286 a_n2804_13878.t21 gnd 0.194556f
C6287 a_n2804_13878.t9 gnd 0.194556f
C6288 a_n2804_13878.n12 gnd 1.53196f
C6289 a_n2804_13878.n13 gnd 4.90178f
C6290 a_n2804_13878.t3 gnd 1.82172f
C6291 a_n2804_13878.t5 gnd 0.194556f
C6292 a_n2804_13878.t6 gnd 0.194556f
C6293 a_n2804_13878.n14 gnd 1.37045f
C6294 a_n2804_13878.n15 gnd 1.53128f
C6295 a_n2804_13878.t2 gnd 1.81809f
C6296 a_n2804_13878.n16 gnd 0.770559f
C6297 a_n2804_13878.t7 gnd 1.81809f
C6298 a_n2804_13878.n17 gnd 0.770559f
C6299 a_n2804_13878.t0 gnd 0.194556f
C6300 a_n2804_13878.t1 gnd 0.194556f
C6301 a_n2804_13878.n18 gnd 1.37045f
C6302 a_n2804_13878.n19 gnd 0.778022f
C6303 a_n2804_13878.t4 gnd 1.81809f
C6304 a_n2804_13878.n20 gnd 2.85814f
C6305 a_n2804_13878.n21 gnd 3.74876f
C6306 a_n2804_13878.t15 gnd 0.194556f
C6307 a_n2804_13878.t24 gnd 0.194556f
C6308 a_n2804_13878.n22 gnd 1.53195f
C6309 a_n2804_13878.n23 gnd 2.50239f
C6310 a_n2804_13878.t28 gnd 0.194556f
C6311 a_n2804_13878.t14 gnd 0.194556f
C6312 a_n2804_13878.n24 gnd 1.53196f
C6313 a_n2804_13878.n25 gnd 0.678771f
C6314 a_n2804_13878.t18 gnd 0.194556f
C6315 a_n2804_13878.t19 gnd 0.194556f
C6316 a_n2804_13878.n26 gnd 1.53196f
C6317 a_n2804_13878.n27 gnd 0.678771f
C6318 a_n2804_13878.n28 gnd 0.678768f
C6319 a_n2804_13878.n29 gnd 1.53196f
C6320 a_n2804_13878.t30 gnd 0.194556f
C6321 a_n2982_13878.n0 gnd 4.29658f
C6322 a_n2982_13878.n1 gnd 3.072f
C6323 a_n2982_13878.n2 gnd 3.92841f
C6324 a_n2982_13878.n3 gnd 0.890133f
C6325 a_n2982_13878.n4 gnd 0.890135f
C6326 a_n2982_13878.n5 gnd 2.81212f
C6327 a_n2982_13878.n6 gnd 0.210577f
C6328 a_n2982_13878.n7 gnd 0.848479f
C6329 a_n2982_13878.n8 gnd 0.210577f
C6330 a_n2982_13878.n9 gnd 0.276098f
C6331 a_n2982_13878.n10 gnd 0.977046f
C6332 a_n2982_13878.n11 gnd 0.210577f
C6333 a_n2982_13878.n12 gnd 0.210577f
C6334 a_n2982_13878.n13 gnd 0.479585f
C6335 a_n2982_13878.n14 gnd 0.210577f
C6336 a_n2982_13878.n15 gnd 0.276098f
C6337 a_n2982_13878.n16 gnd 0.532229f
C6338 a_n2982_13878.n17 gnd 0.908905f
C6339 a_n2982_13878.n18 gnd 0.199803f
C6340 a_n2982_13878.n19 gnd 0.147158f
C6341 a_n2982_13878.n20 gnd 0.231286f
C6342 a_n2982_13878.n21 gnd 0.178642f
C6343 a_n2982_13878.n22 gnd 0.199803f
C6344 a_n2982_13878.n23 gnd 1.33098f
C6345 a_n2982_13878.n24 gnd 0.147158f
C6346 a_n2982_13878.n25 gnd 0.96155f
C6347 a_n2982_13878.n26 gnd 0.210577f
C6348 a_n2982_13878.n27 gnd 0.741157f
C6349 a_n2982_13878.n28 gnd 0.210577f
C6350 a_n2982_13878.n29 gnd 0.210577f
C6351 a_n2982_13878.n30 gnd 0.479585f
C6352 a_n2982_13878.n31 gnd 0.276098f
C6353 a_n2982_13878.n32 gnd 0.210577f
C6354 a_n2982_13878.n33 gnd 0.532229f
C6355 a_n2982_13878.n34 gnd 0.210577f
C6356 a_n2982_13878.n35 gnd 0.210577f
C6357 a_n2982_13878.n36 gnd 0.936913f
C6358 a_n2982_13878.n37 gnd 0.276098f
C6359 a_n2982_13878.n38 gnd 1.73365f
C6360 a_n2982_13878.n39 gnd 1.16816f
C6361 a_n2982_13878.n40 gnd 2.33309f
C6362 a_n2982_13878.n41 gnd 1.16816f
C6363 a_n2982_13878.n42 gnd 2.13309f
C6364 a_n2982_13878.n43 gnd 1.73365f
C6365 a_n2982_13878.n44 gnd 0.008449f
C6366 a_n2982_13878.n45 gnd 4.07e-19
C6367 a_n2982_13878.n47 gnd 0.008153f
C6368 a_n2982_13878.n48 gnd 0.011855f
C6369 a_n2982_13878.n49 gnd 0.007843f
C6370 a_n2982_13878.n51 gnd 0.279311f
C6371 a_n2982_13878.n52 gnd 0.008449f
C6372 a_n2982_13878.n53 gnd 4.07e-19
C6373 a_n2982_13878.n55 gnd 0.008153f
C6374 a_n2982_13878.n56 gnd 0.011855f
C6375 a_n2982_13878.n57 gnd 0.007843f
C6376 a_n2982_13878.n59 gnd 0.279311f
C6377 a_n2982_13878.n60 gnd 0.008153f
C6378 a_n2982_13878.n61 gnd 0.278171f
C6379 a_n2982_13878.n62 gnd 0.008153f
C6380 a_n2982_13878.n63 gnd 0.278171f
C6381 a_n2982_13878.n64 gnd 0.008153f
C6382 a_n2982_13878.n65 gnd 0.278171f
C6383 a_n2982_13878.n66 gnd 0.008153f
C6384 a_n2982_13878.n67 gnd 0.278171f
C6385 a_n2982_13878.n69 gnd 0.279311f
C6386 a_n2982_13878.n70 gnd 0.008449f
C6387 a_n2982_13878.n71 gnd 4.07e-19
C6388 a_n2982_13878.n73 gnd 0.008153f
C6389 a_n2982_13878.n74 gnd 0.011855f
C6390 a_n2982_13878.n75 gnd 0.007843f
C6391 a_n2982_13878.n77 gnd 0.279311f
C6392 a_n2982_13878.n78 gnd 0.008449f
C6393 a_n2982_13878.n79 gnd 4.07e-19
C6394 a_n2982_13878.n81 gnd 0.008153f
C6395 a_n2982_13878.n82 gnd 3.16e-19
C6396 a_n2982_13878.t50 gnd 0.146058f
C6397 a_n2982_13878.t65 gnd 0.693536f
C6398 a_n2982_13878.t21 gnd 0.679392f
C6399 a_n2982_13878.t49 gnd 0.679392f
C6400 a_n2982_13878.t25 gnd 0.679392f
C6401 a_n2982_13878.n83 gnd 0.29857f
C6402 a_n2982_13878.t35 gnd 0.679392f
C6403 a_n2982_13878.t29 gnd 0.679392f
C6404 a_n2982_13878.t61 gnd 0.679392f
C6405 a_n2982_13878.n84 gnd 0.294911f
C6406 a_n2982_13878.t43 gnd 0.679392f
C6407 a_n2982_13878.t57 gnd 0.679392f
C6408 a_n2982_13878.t3 gnd 0.113601f
C6409 a_n2982_13878.t7 gnd 0.113601f
C6410 a_n2982_13878.n85 gnd 1.00678f
C6411 a_n2982_13878.t15 gnd 0.113601f
C6412 a_n2982_13878.t71 gnd 0.113601f
C6413 a_n2982_13878.n86 gnd 1.00382f
C6414 a_n2982_13878.t6 gnd 0.113601f
C6415 a_n2982_13878.t12 gnd 0.113601f
C6416 a_n2982_13878.n87 gnd 1.00382f
C6417 a_n2982_13878.t8 gnd 0.113601f
C6418 a_n2982_13878.t18 gnd 0.113601f
C6419 a_n2982_13878.n88 gnd 1.00678f
C6420 a_n2982_13878.t0 gnd 0.113601f
C6421 a_n2982_13878.t20 gnd 0.113601f
C6422 a_n2982_13878.n89 gnd 1.00382f
C6423 a_n2982_13878.t11 gnd 0.113601f
C6424 a_n2982_13878.t4 gnd 0.113601f
C6425 a_n2982_13878.n90 gnd 1.00382f
C6426 a_n2982_13878.t70 gnd 0.113601f
C6427 a_n2982_13878.t1 gnd 0.113601f
C6428 a_n2982_13878.n91 gnd 1.00382f
C6429 a_n2982_13878.t16 gnd 0.113601f
C6430 a_n2982_13878.t69 gnd 0.113601f
C6431 a_n2982_13878.n92 gnd 1.00382f
C6432 a_n2982_13878.t9 gnd 0.113601f
C6433 a_n2982_13878.t2 gnd 0.113601f
C6434 a_n2982_13878.n93 gnd 1.00382f
C6435 a_n2982_13878.t13 gnd 0.113601f
C6436 a_n2982_13878.t17 gnd 0.113601f
C6437 a_n2982_13878.n94 gnd 1.00678f
C6438 a_n2982_13878.t14 gnd 0.113601f
C6439 a_n2982_13878.t10 gnd 0.113601f
C6440 a_n2982_13878.n95 gnd 1.00382f
C6441 a_n2982_13878.t19 gnd 0.113601f
C6442 a_n2982_13878.t5 gnd 0.113601f
C6443 a_n2982_13878.n96 gnd 1.00382f
C6444 a_n2982_13878.t39 gnd 0.679392f
C6445 a_n2982_13878.n97 gnd 0.294586f
C6446 a_n2982_13878.t41 gnd 0.679392f
C6447 a_n2982_13878.t53 gnd 0.690322f
C6448 a_n2982_13878.t110 gnd 0.693536f
C6449 a_n2982_13878.t87 gnd 0.679392f
C6450 a_n2982_13878.t92 gnd 0.679392f
C6451 a_n2982_13878.t80 gnd 0.679392f
C6452 a_n2982_13878.n98 gnd 0.29857f
C6453 a_n2982_13878.t97 gnd 0.679392f
C6454 a_n2982_13878.t106 gnd 0.679392f
C6455 a_n2982_13878.t107 gnd 0.679392f
C6456 a_n2982_13878.n99 gnd 0.294911f
C6457 a_n2982_13878.t74 gnd 0.679392f
C6458 a_n2982_13878.t89 gnd 0.679392f
C6459 a_n2982_13878.t77 gnd 0.679392f
C6460 a_n2982_13878.n100 gnd 0.298689f
C6461 a_n2982_13878.t84 gnd 0.679392f
C6462 a_n2982_13878.t103 gnd 0.690322f
C6463 a_n2982_13878.t64 gnd 1.36762f
C6464 a_n2982_13878.t38 gnd 0.146058f
C6465 a_n2982_13878.t32 gnd 0.146058f
C6466 a_n2982_13878.n101 gnd 1.02883f
C6467 a_n2982_13878.t46 gnd 0.146058f
C6468 a_n2982_13878.t28 gnd 0.146058f
C6469 a_n2982_13878.n102 gnd 1.02883f
C6470 a_n2982_13878.t60 gnd 0.146058f
C6471 a_n2982_13878.t48 gnd 0.146058f
C6472 a_n2982_13878.n103 gnd 1.02883f
C6473 a_n2982_13878.t68 gnd 0.146058f
C6474 a_n2982_13878.t52 gnd 0.146058f
C6475 a_n2982_13878.n104 gnd 1.02883f
C6476 a_n2982_13878.t56 gnd 0.146058f
C6477 a_n2982_13878.t34 gnd 0.146058f
C6478 a_n2982_13878.n105 gnd 1.02883f
C6479 a_n2982_13878.t24 gnd 1.36489f
C6480 a_n2982_13878.t55 gnd 0.679392f
C6481 a_n2982_13878.n106 gnd 0.298689f
C6482 a_n2982_13878.t33 gnd 0.679392f
C6483 a_n2982_13878.t67 gnd 0.679392f
C6484 a_n2982_13878.n107 gnd 0.289717f
C6485 a_n2982_13878.t27 gnd 0.679392f
C6486 a_n2982_13878.n108 gnd 0.301256f
C6487 a_n2982_13878.t59 gnd 0.679392f
C6488 a_n2982_13878.t31 gnd 0.679392f
C6489 a_n2982_13878.n109 gnd 0.294586f
C6490 a_n2982_13878.t63 gnd 0.693536f
C6491 a_n2982_13878.t86 gnd 0.679392f
C6492 a_n2982_13878.n110 gnd 0.298689f
C6493 a_n2982_13878.t95 gnd 0.679392f
C6494 a_n2982_13878.t101 gnd 0.679392f
C6495 a_n2982_13878.n111 gnd 0.289717f
C6496 a_n2982_13878.t105 gnd 0.679392f
C6497 a_n2982_13878.n112 gnd 0.301256f
C6498 a_n2982_13878.t76 gnd 0.679392f
C6499 a_n2982_13878.t79 gnd 0.679392f
C6500 a_n2982_13878.n113 gnd 0.294586f
C6501 a_n2982_13878.t109 gnd 0.693536f
C6502 a_n2982_13878.t78 gnd 0.679392f
C6503 a_n2982_13878.n114 gnd 0.300815f
C6504 a_n2982_13878.t104 gnd 0.679392f
C6505 a_n2982_13878.n115 gnd 0.29857f
C6506 a_n2982_13878.n116 gnd 0.298704f
C6507 a_n2982_13878.t100 gnd 0.679392f
C6508 a_n2982_13878.n117 gnd 0.294911f
C6509 a_n2982_13878.t73 gnd 0.679392f
C6510 a_n2982_13878.n118 gnd 0.295164f
C6511 a_n2982_13878.n119 gnd 0.300816f
C6512 a_n2982_13878.t75 gnd 0.690322f
C6513 a_n2982_13878.t37 gnd 0.679392f
C6514 a_n2982_13878.n120 gnd 0.300815f
C6515 a_n2982_13878.t45 gnd 0.679392f
C6516 a_n2982_13878.n121 gnd 0.29857f
C6517 a_n2982_13878.n122 gnd 0.298704f
C6518 a_n2982_13878.t47 gnd 0.679392f
C6519 a_n2982_13878.n123 gnd 0.294911f
C6520 a_n2982_13878.t51 gnd 0.679392f
C6521 a_n2982_13878.n124 gnd 0.295164f
C6522 a_n2982_13878.n125 gnd 0.300816f
C6523 a_n2982_13878.t23 gnd 0.690322f
C6524 a_n2982_13878.n126 gnd 1.31538f
C6525 a_n2982_13878.t83 gnd 0.679392f
C6526 a_n2982_13878.n127 gnd 0.294911f
C6527 a_n2982_13878.t91 gnd 0.679392f
C6528 a_n2982_13878.n128 gnd 0.294911f
C6529 a_n2982_13878.t81 gnd 0.679392f
C6530 a_n2982_13878.n129 gnd 0.294911f
C6531 a_n2982_13878.t96 gnd 0.679392f
C6532 a_n2982_13878.n130 gnd 0.294911f
C6533 a_n2982_13878.t85 gnd 0.679392f
C6534 a_n2982_13878.n131 gnd 0.289555f
C6535 a_n2982_13878.t111 gnd 0.679392f
C6536 a_n2982_13878.n132 gnd 0.298704f
C6537 a_n2982_13878.t88 gnd 0.690776f
C6538 a_n2982_13878.t98 gnd 0.679392f
C6539 a_n2982_13878.n133 gnd 0.289555f
C6540 a_n2982_13878.t82 gnd 0.679392f
C6541 a_n2982_13878.n134 gnd 0.298704f
C6542 a_n2982_13878.t93 gnd 0.690776f
C6543 a_n2982_13878.t102 gnd 0.679392f
C6544 a_n2982_13878.n135 gnd 0.289555f
C6545 a_n2982_13878.t90 gnd 0.679392f
C6546 a_n2982_13878.n136 gnd 0.298704f
C6547 a_n2982_13878.t108 gnd 0.690776f
C6548 a_n2982_13878.t94 gnd 0.679392f
C6549 a_n2982_13878.n137 gnd 0.289555f
C6550 a_n2982_13878.t72 gnd 0.679392f
C6551 a_n2982_13878.n138 gnd 0.298704f
C6552 a_n2982_13878.t99 gnd 0.690776f
C6553 a_n2982_13878.n139 gnd 1.65459f
C6554 a_n2982_13878.n140 gnd 0.300816f
C6555 a_n2982_13878.n141 gnd 0.295164f
C6556 a_n2982_13878.n142 gnd 0.289717f
C6557 a_n2982_13878.n143 gnd 0.298704f
C6558 a_n2982_13878.n144 gnd 0.301256f
C6559 a_n2982_13878.n145 gnd 0.294586f
C6560 a_n2982_13878.n146 gnd 0.300815f
C6561 a_n2982_13878.n147 gnd 0.300816f
C6562 a_n2982_13878.n148 gnd 0.011946f
C6563 a_n2982_13878.n149 gnd 0.295164f
C6564 a_n2982_13878.n150 gnd 0.301256f
C6565 a_n2982_13878.n151 gnd 0.298704f
C6566 a_n2982_13878.n152 gnd 0.301256f
C6567 a_n2982_13878.n153 gnd 0.294586f
C6568 a_n2982_13878.n154 gnd 0.300815f
C6569 a_n2982_13878.n155 gnd 1.00016f
C6570 a_n2982_13878.t66 gnd 1.36489f
C6571 a_n2982_13878.t54 gnd 1.36762f
C6572 a_n2982_13878.t40 gnd 0.146058f
C6573 a_n2982_13878.t42 gnd 0.146058f
C6574 a_n2982_13878.n156 gnd 1.02883f
C6575 a_n2982_13878.t44 gnd 0.146058f
C6576 a_n2982_13878.t58 gnd 0.146058f
C6577 a_n2982_13878.n157 gnd 1.02883f
C6578 a_n2982_13878.t30 gnd 0.146058f
C6579 a_n2982_13878.t62 gnd 0.146058f
C6580 a_n2982_13878.n158 gnd 1.02883f
C6581 a_n2982_13878.t26 gnd 0.146058f
C6582 a_n2982_13878.t36 gnd 0.146058f
C6583 a_n2982_13878.n159 gnd 1.02883f
C6584 a_n2982_13878.n160 gnd 1.02884f
C6585 a_n2982_13878.t22 gnd 0.146058f
.ends

