* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t136 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X1 commonsourceibias.t15 commonsourceibias.t14 gnd.t284 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 gnd.t283 commonsourceibias.t64 CSoutput.t19 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 vdd.t151 vdd.t149 vdd.t150 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X4 vdd.t174 a_n6308_8799.t28 CSoutput.t84 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 a_n1986_8322.t3 a_n1986_13878.t40 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 a_n1808_13878.t11 a_n1986_13878.t0 a_n1986_13878.t1 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X7 gnd.t282 commonsourceibias.t65 CSoutput.t106 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n1986_13878.t7 a_n1986_13878.t6 a_n1808_13878.t10 vdd.t158 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 a_n1808_13878.t9 a_n1986_13878.t16 a_n1986_13878.t17 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 vdd.t148 vdd.t146 vdd.t147 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X11 CSoutput.t85 a_n6308_8799.t29 vdd.t175 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 a_n1808_13878.t19 a_n1986_13878.t41 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 vdd.t145 vdd.t143 vdd.t144 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X14 vdd.t142 vdd.t140 vdd.t141 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X15 gnd.t144 gnd.t142 gnd.t143 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X16 gnd.t281 commonsourceibias.t12 commonsourceibias.t13 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 vdd.t213 CSoutput.t137 output.t18 gnd.t304 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 CSoutput.t82 a_n6308_8799.t30 vdd.t172 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 gnd.t280 commonsourceibias.t66 CSoutput.t27 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 CSoutput.t83 a_n6308_8799.t31 vdd.t173 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 gnd.t279 commonsourceibias.t67 CSoutput.t65 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 a_n6308_8799.t5 plus.t5 a_n2903_n3924.t15 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X23 output.t17 CSoutput.t138 vdd.t210 gnd.t303 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X24 a_n1986_8322.t13 a_n1986_13878.t42 a_n6308_8799.t17 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 gnd.t278 commonsourceibias.t10 commonsourceibias.t11 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 CSoutput.t139 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X27 output.t0 outputibias.t8 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X28 a_n6308_8799.t20 plus.t6 a_n2903_n3924.t14 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X29 gnd.t141 gnd.t139 gnd.t140 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X30 CSoutput.t114 commonsourceibias.t68 gnd.t277 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 gnd.t276 commonsourceibias.t8 commonsourceibias.t9 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 CSoutput.t80 a_n6308_8799.t32 vdd.t170 vdd.t164 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 vdd.t171 a_n6308_8799.t33 CSoutput.t81 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 output.t2 outputibias.t9 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X35 a_n6308_8799.t18 a_n1986_13878.t43 a_n1986_8322.t14 vdd.t182 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X36 CSoutput.t125 a_n6308_8799.t34 vdd.t208 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X37 vdd.t209 a_n6308_8799.t35 CSoutput.t126 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 gnd.t138 gnd.t136 plus.t4 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X39 a_n2903_n3924.t26 minus.t5 a_n1986_13878.t27 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X40 CSoutput.t41 commonsourceibias.t69 gnd.t275 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n2903_n3924.t20 diffpairibias.t16 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 vdd.t139 vdd.t136 vdd.t138 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X43 a_n1986_13878.t26 minus.t6 a_n2903_n3924.t25 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X44 a_n2903_n3924.t13 plus.t7 a_n6308_8799.t26 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X45 vdd.t223 CSoutput.t140 output.t16 gnd.t302 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X46 output.t15 CSoutput.t141 vdd.t221 gnd.t301 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 output.t1 outputibias.t10 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X48 CSoutput.t92 commonsourceibias.t70 gnd.t274 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n2903_n3924.t38 minus.t7 a_n1986_13878.t39 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X50 CSoutput.t104 a_n6308_8799.t36 vdd.t195 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 CSoutput.t105 a_n6308_8799.t37 vdd.t196 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 vdd.t135 vdd.t133 vdd.t134 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 gnd.t273 commonsourceibias.t22 commonsourceibias.t23 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X54 CSoutput.t119 commonsourceibias.t71 gnd.t272 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t78 a_n6308_8799.t38 vdd.t167 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 a_n2903_n3924.t23 minus.t8 a_n1986_13878.t24 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X57 a_n1808_13878.t8 a_n1986_13878.t10 a_n1986_13878.t11 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X58 vdd.t169 a_n6308_8799.t39 CSoutput.t79 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 diffpairibias.t15 diffpairibias.t14 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X60 a_n1986_13878.t15 a_n1986_13878.t14 a_n1808_13878.t7 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 CSoutput.t86 a_n6308_8799.t40 vdd.t176 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 vdd.t132 vdd.t130 vdd.t131 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 gnd.t135 gnd.t133 plus.t3 gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X64 minus.t4 gnd.t130 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X65 gnd.t271 commonsourceibias.t72 CSoutput.t111 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 gnd.t270 commonsourceibias.t73 CSoutput.t66 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 diffpairibias.t13 diffpairibias.t12 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X68 gnd.t269 commonsourceibias.t74 CSoutput.t120 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 commonsourceibias.t21 commonsourceibias.t20 gnd.t268 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t177 a_n6308_8799.t41 CSoutput.t87 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t219 CSoutput.t142 output.t14 gnd.t300 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X72 vdd.t53 a_n6308_8799.t42 CSoutput.t52 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 CSoutput.t53 a_n6308_8799.t43 vdd.t54 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X74 gnd.t267 commonsourceibias.t75 CSoutput.t58 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 CSoutput.t143 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X76 commonsourceibias.t19 commonsourceibias.t18 gnd.t266 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 vdd.t193 a_n6308_8799.t44 CSoutput.t102 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 gnd.t265 commonsourceibias.t76 CSoutput.t31 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 a_n6308_8799.t8 plus.t8 a_n2903_n3924.t12 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X80 commonsourceibias.t17 commonsourceibias.t16 gnd.t264 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 CSoutput.t103 a_n6308_8799.t45 vdd.t194 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t109 a_n6308_8799.t46 vdd.t202 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t2 commonsourceibias.t77 gnd.t263 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X84 a_n2903_n3924.t39 diffpairibias.t17 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 gnd.t262 commonsourceibias.t30 commonsourceibias.t31 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 CSoutput.t110 a_n6308_8799.t47 vdd.t203 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n2903_n3924.t24 minus.t9 a_n1986_13878.t25 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X88 vdd.t25 a_n6308_8799.t48 CSoutput.t23 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 a_n2903_n3924.t11 plus.t9 a_n6308_8799.t13 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X90 a_n1986_13878.t28 minus.t10 a_n2903_n3924.t27 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X91 gnd.t261 commonsourceibias.t28 commonsourceibias.t29 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t129 gnd.t127 gnd.t128 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 commonsourceibias.t27 commonsourceibias.t26 gnd.t260 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n1986_13878.t13 a_n1986_13878.t12 a_n1808_13878.t6 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 a_n1986_13878.t23 a_n1986_13878.t22 a_n1808_13878.t5 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X96 vdd.t27 a_n6308_8799.t49 CSoutput.t24 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 vdd.t20 a_n6308_8799.t50 CSoutput.t21 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 a_n6308_8799.t25 a_n1986_13878.t44 a_n1986_8322.t20 vdd.t199 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 CSoutput.t128 commonsourceibias.t78 gnd.t259 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 vdd.t22 a_n6308_8799.t51 CSoutput.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 a_n2903_n3924.t34 minus.t11 a_n1986_13878.t35 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X102 CSoutput.t3 commonsourceibias.t79 gnd.t258 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t20 commonsourceibias.t80 gnd.t257 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 vdd.t200 a_n6308_8799.t52 CSoutput.t107 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X105 gnd.t256 commonsourceibias.t81 CSoutput.t57 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X106 commonsourceibias.t25 commonsourceibias.t24 gnd.t255 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 CSoutput.t108 a_n6308_8799.t53 vdd.t201 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 CSoutput.t124 commonsourceibias.t82 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 CSoutput.t144 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X110 vdd.t190 a_n6308_8799.t54 CSoutput.t100 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 vdd.t129 vdd.t127 vdd.t128 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X112 vdd.t126 vdd.t123 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 gnd.t252 commonsourceibias.t83 CSoutput.t112 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n1986_13878.t34 minus.t12 a_n2903_n3924.t33 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X115 output.t19 outputibias.t11 gnd.t314 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X116 a_n2903_n3924.t16 diffpairibias.t18 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 vdd.t122 vdd.t119 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 CSoutput.t145 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X119 commonsourceibias.t37 commonsourceibias.t36 gnd.t251 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 vdd.t160 a_n1986_13878.t45 a_n1986_8322.t11 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X121 vdd.t118 vdd.t116 vdd.t117 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 a_n2903_n3924.t10 plus.t10 a_n6308_8799.t24 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X123 CSoutput.t101 a_n6308_8799.t55 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 a_n1986_8322.t10 a_n1986_13878.t46 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 vdd.t74 a_n6308_8799.t56 CSoutput.t71 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 gnd.t250 commonsourceibias.t34 commonsourceibias.t35 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t248 commonsourceibias.t84 CSoutput.t4 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 vdd.t227 a_n1986_13878.t47 a_n1808_13878.t18 vdd.t226 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t247 commonsourceibias.t85 CSoutput.t122 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 a_n6308_8799.t6 plus.t11 a_n2903_n3924.t9 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X131 gnd.t245 commonsourceibias.t86 CSoutput.t18 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 commonsourceibias.t33 commonsourceibias.t32 gnd.t244 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t115 vdd.t112 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X134 vdd.t224 CSoutput.t146 output.t13 gnd.t299 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X135 diffpairibias.t11 diffpairibias.t10 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X136 vdd.t111 vdd.t108 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X137 vdd.t75 a_n6308_8799.t57 CSoutput.t72 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 gnd.t243 commonsourceibias.t87 CSoutput.t40 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t126 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X140 a_n6308_8799.t0 a_n1986_13878.t48 a_n1986_8322.t0 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 a_n1986_8322.t1 a_n1986_13878.t49 vdd.t2 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X142 vdd.t107 vdd.t104 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X143 plus.t2 gnd.t120 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X144 CSoutput.t127 commonsourceibias.t88 gnd.t242 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X145 gnd.t241 commonsourceibias.t89 CSoutput.t45 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 vdd.t188 a_n6308_8799.t58 CSoutput.t98 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X147 a_n1986_13878.t9 a_n1986_13878.t8 a_n1808_13878.t4 vdd.t71 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X148 commonsourceibias.t1 commonsourceibias.t0 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X149 CSoutput.t99 a_n6308_8799.t59 vdd.t189 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 a_n6308_8799.t7 a_n1986_13878.t50 a_n1986_8322.t6 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 gnd.t119 gnd.t117 minus.t3 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X152 CSoutput.t44 commonsourceibias.t90 gnd.t237 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n1986_13878.t33 minus.t13 a_n2903_n3924.t32 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X154 a_n1808_13878.t3 a_n1986_13878.t4 a_n1986_13878.t5 vdd.t199 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 vdd.t44 a_n1986_13878.t51 a_n1986_8322.t4 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X156 gnd.t116 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 a_n2903_n3924.t17 diffpairibias.t19 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 CSoutput.t129 commonsourceibias.t91 gnd.t236 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 CSoutput.t36 a_n6308_8799.t60 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput.t77 commonsourceibias.t92 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n1986_13878.t32 minus.t14 a_n2903_n3924.t31 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X162 CSoutput.t17 commonsourceibias.t93 gnd.t233 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n2903_n3924.t19 diffpairibias.t20 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X164 vdd.t42 a_n6308_8799.t61 CSoutput.t37 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X165 gnd.t232 commonsourceibias.t94 CSoutput.t46 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X166 gnd.t230 commonsourceibias.t95 CSoutput.t15 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput.t56 commonsourceibias.t96 gnd.t229 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 commonsourceibias.t41 commonsourceibias.t40 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 vdd.t222 CSoutput.t147 output.t12 gnd.t298 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X170 vdd.t49 a_n6308_8799.t62 CSoutput.t49 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 gnd.t226 commonsourceibias.t97 CSoutput.t117 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 gnd.t112 gnd.t109 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X173 a_n1986_13878.t31 minus.t15 a_n2903_n3924.t30 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X174 CSoutput.t123 commonsourceibias.t98 gnd.t225 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t108 gnd.t106 gnd.t107 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X176 diffpairibias.t9 diffpairibias.t8 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X177 CSoutput.t50 a_n6308_8799.t63 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 a_n2903_n3924.t8 plus.t12 a_n6308_8799.t14 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X179 CSoutput.t134 a_n6308_8799.t64 vdd.t230 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 CSoutput.t51 commonsourceibias.t99 gnd.t224 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X181 gnd.t223 commonsourceibias.t100 CSoutput.t131 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 vdd.t103 vdd.t101 vdd.t102 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X183 a_n1808_13878.t17 a_n1986_13878.t52 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X184 vdd.t24 a_n1986_13878.t53 a_n1808_13878.t16 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 gnd.t105 gnd.t103 minus.t2 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X186 plus.t1 gnd.t100 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X187 gnd.t99 gnd.t97 gnd.t98 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X188 gnd.t96 gnd.t94 gnd.t95 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X189 a_n2903_n3924.t7 plus.t13 a_n6308_8799.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X190 gnd.t222 commonsourceibias.t38 commonsourceibias.t39 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 gnd.t221 commonsourceibias.t101 CSoutput.t91 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t220 commonsourceibias.t102 CSoutput.t0 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 CSoutput.t90 commonsourceibias.t103 gnd.t219 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 diffpairibias.t7 diffpairibias.t6 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X195 CSoutput.t135 a_n6308_8799.t65 vdd.t231 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 gnd.t215 commonsourceibias.t44 commonsourceibias.t45 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 output.t11 CSoutput.t148 vdd.t216 gnd.t297 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X198 vdd.t72 a_n6308_8799.t66 CSoutput.t69 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X199 CSoutput.t14 commonsourceibias.t104 gnd.t218 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 gnd.t93 gnd.t91 gnd.t92 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 a_n1986_8322.t12 a_n1986_13878.t54 a_n6308_8799.t16 vdd.t158 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 CSoutput.t118 commonsourceibias.t105 gnd.t217 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 vdd.t73 a_n6308_8799.t67 CSoutput.t70 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 CSoutput.t29 a_n6308_8799.t68 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 vdd.t33 a_n6308_8799.t69 CSoutput.t30 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 vdd.t205 a_n1986_13878.t55 a_n1986_8322.t18 vdd.t204 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X207 gnd.t90 gnd.t88 minus.t1 gnd.t89 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X208 gnd.t216 commonsourceibias.t46 commonsourceibias.t47 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 a_n1808_13878.t15 a_n1986_13878.t56 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X210 gnd.t87 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X211 CSoutput.t25 commonsourceibias.t106 gnd.t213 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 gnd.t83 gnd.t80 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X213 a_n2903_n3924.t21 diffpairibias.t21 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X214 vdd.t161 a_n6308_8799.t70 CSoutput.t73 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 vdd.t100 vdd.t98 vdd.t99 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X216 CSoutput.t74 a_n6308_8799.t71 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 output.t10 CSoutput.t149 vdd.t215 gnd.t296 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X218 CSoutput.t16 commonsourceibias.t107 gnd.t212 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 CSoutput.t75 a_n6308_8799.t72 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 gnd.t211 commonsourceibias.t108 CSoutput.t39 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X221 vdd.t97 vdd.t95 vdd.t96 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X222 CSoutput.t38 commonsourceibias.t109 gnd.t209 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 gnd.t79 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X224 gnd.t208 commonsourceibias.t42 commonsourceibias.t43 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 a_n1986_8322.t9 a_n1986_13878.t57 a_n6308_8799.t12 vdd.t71 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X226 vdd.t58 a_n1986_13878.t58 a_n1986_8322.t5 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X227 vdd.t166 a_n6308_8799.t73 CSoutput.t76 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 CSoutput.t115 a_n6308_8799.t74 vdd.t206 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 gnd.t206 commonsourceibias.t110 CSoutput.t26 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 CSoutput.t116 a_n6308_8799.t75 vdd.t207 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X231 a_n2903_n3924.t6 plus.t14 a_n6308_8799.t4 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X232 vdd.t220 CSoutput.t150 output.t9 gnd.t295 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X233 gnd.t75 gnd.t73 gnd.t74 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X234 output.t8 CSoutput.t151 vdd.t218 gnd.t294 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X235 vdd.t64 a_n6308_8799.t76 CSoutput.t62 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 vdd.t65 a_n6308_8799.t77 CSoutput.t63 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n2903_n3924.t29 minus.t16 a_n1986_13878.t30 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X238 a_n6308_8799.t15 plus.t15 a_n2903_n3924.t5 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X239 outputibias.t7 outputibias.t6 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X240 gnd.t72 gnd.t70 gnd.t71 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X241 CSoutput.t6 commonsourceibias.t111 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 diffpairibias.t5 diffpairibias.t4 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X243 vdd.t94 vdd.t91 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X244 a_n6308_8799.t27 plus.t16 a_n2903_n3924.t4 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X245 a_n2903_n3924.t28 minus.t17 a_n1986_13878.t29 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X246 outputibias.t5 outputibias.t4 gnd.t306 gnd.t305 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X247 a_n1808_13878.t2 a_n1986_13878.t2 a_n1986_13878.t3 vdd.t68 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 gnd.t203 commonsourceibias.t112 CSoutput.t121 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t67 commonsourceibias.t113 gnd.t201 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X250 a_n1986_8322.t8 a_n1986_13878.t59 a_n6308_8799.t11 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X251 outputibias.t3 outputibias.t2 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X252 gnd.t200 commonsourceibias.t114 CSoutput.t28 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 outputibias.t1 outputibias.t0 gnd.t310 gnd.t309 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X254 gnd.t170 commonsourceibias.t60 commonsourceibias.t61 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t185 a_n6308_8799.t78 CSoutput.t96 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 CSoutput.t97 a_n6308_8799.t79 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 a_n2903_n3924.t3 plus.t17 a_n6308_8799.t9 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X258 output.t7 CSoutput.t152 vdd.t225 gnd.t293 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X259 CSoutput.t113 commonsourceibias.t115 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t228 a_n6308_8799.t80 CSoutput.t132 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 CSoutput.t133 a_n6308_8799.t81 vdd.t229 vdd.t164 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 a_n1986_8322.t16 a_n1986_13878.t60 vdd.t198 vdd.t197 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X263 vdd.t90 vdd.t87 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X264 gnd.t69 gnd.t66 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X265 CSoutput.t64 commonsourceibias.t116 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 CSoutput.t59 commonsourceibias.t117 gnd.t195 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 gnd.t194 commonsourceibias.t118 CSoutput.t93 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 gnd.t193 commonsourceibias.t50 commonsourceibias.t51 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 gnd.t65 gnd.t62 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X270 a_n2903_n3924.t35 minus.t18 a_n1986_13878.t36 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X271 output.t6 CSoutput.t153 vdd.t217 gnd.t292 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X272 vdd.t4 a_n1986_13878.t61 a_n1808_13878.t14 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X273 CSoutput.t10 a_n6308_8799.t82 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X274 vdd.t13 a_n6308_8799.t83 CSoutput.t11 vdd.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t179 a_n6308_8799.t84 CSoutput.t88 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X277 a_n1986_8322.t15 a_n1986_13878.t62 a_n6308_8799.t19 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X278 vdd.t82 vdd.t80 vdd.t81 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X279 a_n6308_8799.t10 a_n1986_13878.t63 a_n1986_8322.t7 vdd.t68 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 a_n1808_13878.t13 a_n1986_13878.t64 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X281 vdd.t180 a_n6308_8799.t85 CSoutput.t89 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 CSoutput.t47 a_n6308_8799.t86 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 CSoutput.t54 commonsourceibias.t119 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 a_n1986_13878.t38 minus.t19 a_n2903_n3924.t37 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X285 commonsourceibias.t49 commonsourceibias.t48 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t187 commonsourceibias.t120 CSoutput.t68 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 vdd.t211 CSoutput.t154 output.t5 gnd.t291 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X288 gnd.t186 commonsourceibias.t121 CSoutput.t130 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 a_n6308_8799.t21 plus.t18 a_n2903_n3924.t2 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X290 CSoutput.t48 a_n6308_8799.t87 vdd.t48 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 a_n1808_13878.t1 a_n1986_13878.t18 a_n1986_13878.t19 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X292 gnd.t61 gnd.t59 gnd.t60 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X293 gnd.t58 gnd.t55 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X294 a_n2903_n3924.t18 diffpairibias.t22 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X295 gnd.t184 commonsourceibias.t122 CSoutput.t55 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 commonsourceibias.t7 commonsourceibias.t6 gnd.t182 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 vdd.t212 CSoutput.t155 output.t4 gnd.t290 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X298 a_n2903_n3924.t1 plus.t19 a_n6308_8799.t23 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X299 CSoutput.t94 a_n6308_8799.t88 vdd.t183 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t184 a_n6308_8799.t89 CSoutput.t95 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t156 a_n1986_8322.t19 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X302 diffpairibias.t3 diffpairibias.t2 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X303 a_n6308_8799.t22 a_n1986_13878.t65 a_n1986_8322.t17 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X304 a_n1986_13878.t21 a_n1986_13878.t20 a_n1808_13878.t0 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X305 vdd.t61 a_n6308_8799.t90 CSoutput.t60 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 commonsourceibias.t5 commonsourceibias.t4 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 gnd.t179 commonsourceibias.t123 CSoutput.t42 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X309 vdd.t63 a_n6308_8799.t91 CSoutput.t61 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X310 a_n6308_8799.t2 plus.t20 a_n2903_n3924.t0 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X311 diffpairibias.t1 diffpairibias.t0 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X312 gnd.t54 gnd.t51 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X313 CSoutput.t34 a_n6308_8799.t92 vdd.t38 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X314 CSoutput.t43 commonsourceibias.t124 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 gnd.t175 commonsourceibias.t125 CSoutput.t5 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 CSoutput.t1 commonsourceibias.t126 gnd.t174 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 commonsourceibias.t59 commonsourceibias.t58 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 gnd.t172 commonsourceibias.t2 commonsourceibias.t3 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 vdd.t70 a_n1986_13878.t66 a_n1808_13878.t12 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X320 CSoutput.t35 a_n6308_8799.t93 vdd.t39 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 CSoutput.t7 commonsourceibias.t127 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 a_n1986_13878.t37 minus.t20 a_n2903_n3924.t36 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X323 output.t3 CSoutput.t157 vdd.t214 gnd.t289 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X324 CSoutput.t32 a_n6308_8799.t94 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 vdd.t37 a_n6308_8799.t95 CSoutput.t33 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 gnd.t164 commonsourceibias.t56 commonsourceibias.t57 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 gnd.t50 gnd.t47 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X328 gnd.t46 gnd.t44 gnd.t45 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X329 commonsourceibias.t55 commonsourceibias.t54 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t8 a_n6308_8799.t96 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 gnd.t43 gnd.t41 plus.t0 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X332 vdd.t9 a_n6308_8799.t97 CSoutput.t9 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 a_n1986_8322.t2 a_n1986_13878.t67 a_n6308_8799.t1 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X334 minus.t0 gnd.t38 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X335 commonsourceibias.t53 commonsourceibias.t52 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X336 vdd.t16 a_n6308_8799.t98 CSoutput.t12 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t13 a_n6308_8799.t99 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X338 gnd.t158 commonsourceibias.t62 commonsourceibias.t63 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 a_n2903_n3924.t22 diffpairibias.t23 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 CSoutput.n19 CSoutput.t138 184.661
R1 CSoutput.n78 CSoutput.n77 165.8
R2 CSoutput.n76 CSoutput.n0 165.8
R3 CSoutput.n75 CSoutput.n74 165.8
R4 CSoutput.n73 CSoutput.n72 165.8
R5 CSoutput.n71 CSoutput.n2 165.8
R6 CSoutput.n69 CSoutput.n68 165.8
R7 CSoutput.n67 CSoutput.n3 165.8
R8 CSoutput.n66 CSoutput.n65 165.8
R9 CSoutput.n63 CSoutput.n4 165.8
R10 CSoutput.n61 CSoutput.n60 165.8
R11 CSoutput.n59 CSoutput.n5 165.8
R12 CSoutput.n58 CSoutput.n57 165.8
R13 CSoutput.n55 CSoutput.n6 165.8
R14 CSoutput.n54 CSoutput.n53 165.8
R15 CSoutput.n52 CSoutput.n51 165.8
R16 CSoutput.n50 CSoutput.n8 165.8
R17 CSoutput.n48 CSoutput.n47 165.8
R18 CSoutput.n46 CSoutput.n9 165.8
R19 CSoutput.n45 CSoutput.n44 165.8
R20 CSoutput.n42 CSoutput.n10 165.8
R21 CSoutput.n41 CSoutput.n40 165.8
R22 CSoutput.n39 CSoutput.n38 165.8
R23 CSoutput.n37 CSoutput.n12 165.8
R24 CSoutput.n35 CSoutput.n34 165.8
R25 CSoutput.n33 CSoutput.n13 165.8
R26 CSoutput.n32 CSoutput.n31 165.8
R27 CSoutput.n29 CSoutput.n14 165.8
R28 CSoutput.n28 CSoutput.n27 165.8
R29 CSoutput.n26 CSoutput.n25 165.8
R30 CSoutput.n24 CSoutput.n16 165.8
R31 CSoutput.n22 CSoutput.n21 165.8
R32 CSoutput.n20 CSoutput.n17 165.8
R33 CSoutput.n77 CSoutput.t140 162.194
R34 CSoutput.n18 CSoutput.t155 120.501
R35 CSoutput.n23 CSoutput.t151 120.501
R36 CSoutput.n15 CSoutput.t147 120.501
R37 CSoutput.n30 CSoutput.t157 120.501
R38 CSoutput.n36 CSoutput.t137 120.501
R39 CSoutput.n11 CSoutput.t148 120.501
R40 CSoutput.n43 CSoutput.t146 120.501
R41 CSoutput.n49 CSoutput.t141 120.501
R42 CSoutput.n7 CSoutput.t150 120.501
R43 CSoutput.n56 CSoutput.t152 120.501
R44 CSoutput.n62 CSoutput.t142 120.501
R45 CSoutput.n64 CSoutput.t153 120.501
R46 CSoutput.n70 CSoutput.t154 120.501
R47 CSoutput.n1 CSoutput.t149 120.501
R48 CSoutput.n290 CSoutput.n288 103.469
R49 CSoutput.n278 CSoutput.n276 103.469
R50 CSoutput.n267 CSoutput.n265 103.469
R51 CSoutput.n104 CSoutput.n102 103.469
R52 CSoutput.n92 CSoutput.n90 103.469
R53 CSoutput.n81 CSoutput.n79 103.469
R54 CSoutput.n296 CSoutput.n295 103.111
R55 CSoutput.n294 CSoutput.n293 103.111
R56 CSoutput.n292 CSoutput.n291 103.111
R57 CSoutput.n290 CSoutput.n289 103.111
R58 CSoutput.n286 CSoutput.n285 103.111
R59 CSoutput.n284 CSoutput.n283 103.111
R60 CSoutput.n282 CSoutput.n281 103.111
R61 CSoutput.n280 CSoutput.n279 103.111
R62 CSoutput.n278 CSoutput.n277 103.111
R63 CSoutput.n275 CSoutput.n274 103.111
R64 CSoutput.n273 CSoutput.n272 103.111
R65 CSoutput.n271 CSoutput.n270 103.111
R66 CSoutput.n269 CSoutput.n268 103.111
R67 CSoutput.n267 CSoutput.n266 103.111
R68 CSoutput.n104 CSoutput.n103 103.111
R69 CSoutput.n106 CSoutput.n105 103.111
R70 CSoutput.n108 CSoutput.n107 103.111
R71 CSoutput.n110 CSoutput.n109 103.111
R72 CSoutput.n112 CSoutput.n111 103.111
R73 CSoutput.n92 CSoutput.n91 103.111
R74 CSoutput.n94 CSoutput.n93 103.111
R75 CSoutput.n96 CSoutput.n95 103.111
R76 CSoutput.n98 CSoutput.n97 103.111
R77 CSoutput.n100 CSoutput.n99 103.111
R78 CSoutput.n81 CSoutput.n80 103.111
R79 CSoutput.n83 CSoutput.n82 103.111
R80 CSoutput.n85 CSoutput.n84 103.111
R81 CSoutput.n87 CSoutput.n86 103.111
R82 CSoutput.n89 CSoutput.n88 103.111
R83 CSoutput.n298 CSoutput.n297 103.111
R84 CSoutput.n318 CSoutput.n316 81.5057
R85 CSoutput.n303 CSoutput.n301 81.5057
R86 CSoutput.n350 CSoutput.n348 81.5057
R87 CSoutput.n335 CSoutput.n333 81.5057
R88 CSoutput.n330 CSoutput.n329 80.9324
R89 CSoutput.n328 CSoutput.n327 80.9324
R90 CSoutput.n326 CSoutput.n325 80.9324
R91 CSoutput.n324 CSoutput.n323 80.9324
R92 CSoutput.n322 CSoutput.n321 80.9324
R93 CSoutput.n320 CSoutput.n319 80.9324
R94 CSoutput.n318 CSoutput.n317 80.9324
R95 CSoutput.n315 CSoutput.n314 80.9324
R96 CSoutput.n313 CSoutput.n312 80.9324
R97 CSoutput.n311 CSoutput.n310 80.9324
R98 CSoutput.n309 CSoutput.n308 80.9324
R99 CSoutput.n307 CSoutput.n306 80.9324
R100 CSoutput.n305 CSoutput.n304 80.9324
R101 CSoutput.n303 CSoutput.n302 80.9324
R102 CSoutput.n350 CSoutput.n349 80.9324
R103 CSoutput.n352 CSoutput.n351 80.9324
R104 CSoutput.n354 CSoutput.n353 80.9324
R105 CSoutput.n356 CSoutput.n355 80.9324
R106 CSoutput.n358 CSoutput.n357 80.9324
R107 CSoutput.n360 CSoutput.n359 80.9324
R108 CSoutput.n362 CSoutput.n361 80.9324
R109 CSoutput.n335 CSoutput.n334 80.9324
R110 CSoutput.n337 CSoutput.n336 80.9324
R111 CSoutput.n339 CSoutput.n338 80.9324
R112 CSoutput.n341 CSoutput.n340 80.9324
R113 CSoutput.n343 CSoutput.n342 80.9324
R114 CSoutput.n345 CSoutput.n344 80.9324
R115 CSoutput.n347 CSoutput.n346 80.9324
R116 CSoutput.n25 CSoutput.n24 48.1486
R117 CSoutput.n69 CSoutput.n3 48.1486
R118 CSoutput.n38 CSoutput.n37 48.1486
R119 CSoutput.n42 CSoutput.n41 48.1486
R120 CSoutput.n51 CSoutput.n50 48.1486
R121 CSoutput.n55 CSoutput.n54 48.1486
R122 CSoutput.n22 CSoutput.n17 46.462
R123 CSoutput.n72 CSoutput.n71 46.462
R124 CSoutput.n20 CSoutput.n19 44.9055
R125 CSoutput.n29 CSoutput.n28 43.7635
R126 CSoutput.n65 CSoutput.n63 43.7635
R127 CSoutput.n35 CSoutput.n13 41.7396
R128 CSoutput.n57 CSoutput.n5 41.7396
R129 CSoutput.n44 CSoutput.n9 37.0171
R130 CSoutput.n48 CSoutput.n9 37.0171
R131 CSoutput.n76 CSoutput.n75 34.9932
R132 CSoutput.n31 CSoutput.n13 32.2947
R133 CSoutput.n61 CSoutput.n5 32.2947
R134 CSoutput.n30 CSoutput.n29 29.6014
R135 CSoutput.n63 CSoutput.n62 29.6014
R136 CSoutput.n19 CSoutput.n18 28.4085
R137 CSoutput.n18 CSoutput.n17 25.1176
R138 CSoutput.n72 CSoutput.n1 25.1176
R139 CSoutput.n43 CSoutput.n42 22.0922
R140 CSoutput.n50 CSoutput.n49 22.0922
R141 CSoutput.n77 CSoutput.n76 21.8586
R142 CSoutput.n37 CSoutput.n36 18.9681
R143 CSoutput.n56 CSoutput.n55 18.9681
R144 CSoutput.n25 CSoutput.n15 17.6292
R145 CSoutput.n64 CSoutput.n3 17.6292
R146 CSoutput.n24 CSoutput.n23 15.844
R147 CSoutput.n70 CSoutput.n69 15.844
R148 CSoutput.n38 CSoutput.n11 14.5051
R149 CSoutput.n54 CSoutput.n7 14.5051
R150 CSoutput.n365 CSoutput.n78 11.6139
R151 CSoutput.n41 CSoutput.n11 11.3811
R152 CSoutput.n51 CSoutput.n7 11.3811
R153 CSoutput.n23 CSoutput.n22 10.0422
R154 CSoutput.n71 CSoutput.n70 10.0422
R155 CSoutput.n287 CSoutput.n275 9.25285
R156 CSoutput.n101 CSoutput.n89 9.25285
R157 CSoutput.n332 CSoutput.n300 8.99096
R158 CSoutput.n331 CSoutput.n315 8.97993
R159 CSoutput.n363 CSoutput.n347 8.97993
R160 CSoutput.n28 CSoutput.n15 8.25698
R161 CSoutput.n65 CSoutput.n64 8.25698
R162 CSoutput.n332 CSoutput.n331 7.89345
R163 CSoutput.n364 CSoutput.n363 7.89345
R164 CSoutput.n300 CSoutput.n299 7.12641
R165 CSoutput.n114 CSoutput.n113 7.12641
R166 CSoutput.n36 CSoutput.n35 6.91809
R167 CSoutput.n57 CSoutput.n56 6.91809
R168 CSoutput.n365 CSoutput.n114 5.39852
R169 CSoutput.n331 CSoutput.n330 5.25266
R170 CSoutput.n363 CSoutput.n362 5.25266
R171 CSoutput.n299 CSoutput.n298 5.1449
R172 CSoutput.n287 CSoutput.n286 5.1449
R173 CSoutput.n113 CSoutput.n112 5.1449
R174 CSoutput.n101 CSoutput.n100 5.1449
R175 CSoutput.n205 CSoutput.n158 4.5005
R176 CSoutput.n174 CSoutput.n158 4.5005
R177 CSoutput.n169 CSoutput.n153 4.5005
R178 CSoutput.n169 CSoutput.n155 4.5005
R179 CSoutput.n169 CSoutput.n152 4.5005
R180 CSoutput.n169 CSoutput.n156 4.5005
R181 CSoutput.n169 CSoutput.n151 4.5005
R182 CSoutput.n169 CSoutput.t156 4.5005
R183 CSoutput.n169 CSoutput.n150 4.5005
R184 CSoutput.n169 CSoutput.n157 4.5005
R185 CSoutput.n169 CSoutput.n158 4.5005
R186 CSoutput.n167 CSoutput.n153 4.5005
R187 CSoutput.n167 CSoutput.n155 4.5005
R188 CSoutput.n167 CSoutput.n152 4.5005
R189 CSoutput.n167 CSoutput.n156 4.5005
R190 CSoutput.n167 CSoutput.n151 4.5005
R191 CSoutput.n167 CSoutput.t156 4.5005
R192 CSoutput.n167 CSoutput.n150 4.5005
R193 CSoutput.n167 CSoutput.n157 4.5005
R194 CSoutput.n167 CSoutput.n158 4.5005
R195 CSoutput.n166 CSoutput.n153 4.5005
R196 CSoutput.n166 CSoutput.n155 4.5005
R197 CSoutput.n166 CSoutput.n152 4.5005
R198 CSoutput.n166 CSoutput.n156 4.5005
R199 CSoutput.n166 CSoutput.n151 4.5005
R200 CSoutput.n166 CSoutput.t156 4.5005
R201 CSoutput.n166 CSoutput.n150 4.5005
R202 CSoutput.n166 CSoutput.n157 4.5005
R203 CSoutput.n166 CSoutput.n158 4.5005
R204 CSoutput.n251 CSoutput.n153 4.5005
R205 CSoutput.n251 CSoutput.n155 4.5005
R206 CSoutput.n251 CSoutput.n152 4.5005
R207 CSoutput.n251 CSoutput.n156 4.5005
R208 CSoutput.n251 CSoutput.n151 4.5005
R209 CSoutput.n251 CSoutput.t156 4.5005
R210 CSoutput.n251 CSoutput.n150 4.5005
R211 CSoutput.n251 CSoutput.n157 4.5005
R212 CSoutput.n251 CSoutput.n158 4.5005
R213 CSoutput.n249 CSoutput.n153 4.5005
R214 CSoutput.n249 CSoutput.n155 4.5005
R215 CSoutput.n249 CSoutput.n152 4.5005
R216 CSoutput.n249 CSoutput.n156 4.5005
R217 CSoutput.n249 CSoutput.n151 4.5005
R218 CSoutput.n249 CSoutput.t156 4.5005
R219 CSoutput.n249 CSoutput.n150 4.5005
R220 CSoutput.n249 CSoutput.n157 4.5005
R221 CSoutput.n247 CSoutput.n153 4.5005
R222 CSoutput.n247 CSoutput.n155 4.5005
R223 CSoutput.n247 CSoutput.n152 4.5005
R224 CSoutput.n247 CSoutput.n156 4.5005
R225 CSoutput.n247 CSoutput.n151 4.5005
R226 CSoutput.n247 CSoutput.t156 4.5005
R227 CSoutput.n247 CSoutput.n150 4.5005
R228 CSoutput.n247 CSoutput.n157 4.5005
R229 CSoutput.n177 CSoutput.n153 4.5005
R230 CSoutput.n177 CSoutput.n155 4.5005
R231 CSoutput.n177 CSoutput.n152 4.5005
R232 CSoutput.n177 CSoutput.n156 4.5005
R233 CSoutput.n177 CSoutput.n151 4.5005
R234 CSoutput.n177 CSoutput.t156 4.5005
R235 CSoutput.n177 CSoutput.n150 4.5005
R236 CSoutput.n177 CSoutput.n157 4.5005
R237 CSoutput.n177 CSoutput.n158 4.5005
R238 CSoutput.n176 CSoutput.n153 4.5005
R239 CSoutput.n176 CSoutput.n155 4.5005
R240 CSoutput.n176 CSoutput.n152 4.5005
R241 CSoutput.n176 CSoutput.n156 4.5005
R242 CSoutput.n176 CSoutput.n151 4.5005
R243 CSoutput.n176 CSoutput.t156 4.5005
R244 CSoutput.n176 CSoutput.n150 4.5005
R245 CSoutput.n176 CSoutput.n157 4.5005
R246 CSoutput.n176 CSoutput.n158 4.5005
R247 CSoutput.n180 CSoutput.n153 4.5005
R248 CSoutput.n180 CSoutput.n155 4.5005
R249 CSoutput.n180 CSoutput.n152 4.5005
R250 CSoutput.n180 CSoutput.n156 4.5005
R251 CSoutput.n180 CSoutput.n151 4.5005
R252 CSoutput.n180 CSoutput.t156 4.5005
R253 CSoutput.n180 CSoutput.n150 4.5005
R254 CSoutput.n180 CSoutput.n157 4.5005
R255 CSoutput.n180 CSoutput.n158 4.5005
R256 CSoutput.n179 CSoutput.n153 4.5005
R257 CSoutput.n179 CSoutput.n155 4.5005
R258 CSoutput.n179 CSoutput.n152 4.5005
R259 CSoutput.n179 CSoutput.n156 4.5005
R260 CSoutput.n179 CSoutput.n151 4.5005
R261 CSoutput.n179 CSoutput.t156 4.5005
R262 CSoutput.n179 CSoutput.n150 4.5005
R263 CSoutput.n179 CSoutput.n157 4.5005
R264 CSoutput.n179 CSoutput.n158 4.5005
R265 CSoutput.n162 CSoutput.n153 4.5005
R266 CSoutput.n162 CSoutput.n155 4.5005
R267 CSoutput.n162 CSoutput.n152 4.5005
R268 CSoutput.n162 CSoutput.n156 4.5005
R269 CSoutput.n162 CSoutput.n151 4.5005
R270 CSoutput.n162 CSoutput.t156 4.5005
R271 CSoutput.n162 CSoutput.n150 4.5005
R272 CSoutput.n162 CSoutput.n157 4.5005
R273 CSoutput.n162 CSoutput.n158 4.5005
R274 CSoutput.n254 CSoutput.n153 4.5005
R275 CSoutput.n254 CSoutput.n155 4.5005
R276 CSoutput.n254 CSoutput.n152 4.5005
R277 CSoutput.n254 CSoutput.n156 4.5005
R278 CSoutput.n254 CSoutput.n151 4.5005
R279 CSoutput.n254 CSoutput.t156 4.5005
R280 CSoutput.n254 CSoutput.n150 4.5005
R281 CSoutput.n254 CSoutput.n157 4.5005
R282 CSoutput.n254 CSoutput.n158 4.5005
R283 CSoutput.n241 CSoutput.n212 4.5005
R284 CSoutput.n241 CSoutput.n218 4.5005
R285 CSoutput.n199 CSoutput.n188 4.5005
R286 CSoutput.n199 CSoutput.n190 4.5005
R287 CSoutput.n199 CSoutput.n187 4.5005
R288 CSoutput.n199 CSoutput.n191 4.5005
R289 CSoutput.n199 CSoutput.n186 4.5005
R290 CSoutput.n199 CSoutput.t136 4.5005
R291 CSoutput.n199 CSoutput.n185 4.5005
R292 CSoutput.n199 CSoutput.n192 4.5005
R293 CSoutput.n241 CSoutput.n199 4.5005
R294 CSoutput.n220 CSoutput.n188 4.5005
R295 CSoutput.n220 CSoutput.n190 4.5005
R296 CSoutput.n220 CSoutput.n187 4.5005
R297 CSoutput.n220 CSoutput.n191 4.5005
R298 CSoutput.n220 CSoutput.n186 4.5005
R299 CSoutput.n220 CSoutput.t136 4.5005
R300 CSoutput.n220 CSoutput.n185 4.5005
R301 CSoutput.n220 CSoutput.n192 4.5005
R302 CSoutput.n241 CSoutput.n220 4.5005
R303 CSoutput.n198 CSoutput.n188 4.5005
R304 CSoutput.n198 CSoutput.n190 4.5005
R305 CSoutput.n198 CSoutput.n187 4.5005
R306 CSoutput.n198 CSoutput.n191 4.5005
R307 CSoutput.n198 CSoutput.n186 4.5005
R308 CSoutput.n198 CSoutput.t136 4.5005
R309 CSoutput.n198 CSoutput.n185 4.5005
R310 CSoutput.n198 CSoutput.n192 4.5005
R311 CSoutput.n241 CSoutput.n198 4.5005
R312 CSoutput.n222 CSoutput.n188 4.5005
R313 CSoutput.n222 CSoutput.n190 4.5005
R314 CSoutput.n222 CSoutput.n187 4.5005
R315 CSoutput.n222 CSoutput.n191 4.5005
R316 CSoutput.n222 CSoutput.n186 4.5005
R317 CSoutput.n222 CSoutput.t136 4.5005
R318 CSoutput.n222 CSoutput.n185 4.5005
R319 CSoutput.n222 CSoutput.n192 4.5005
R320 CSoutput.n241 CSoutput.n222 4.5005
R321 CSoutput.n188 CSoutput.n183 4.5005
R322 CSoutput.n190 CSoutput.n183 4.5005
R323 CSoutput.n187 CSoutput.n183 4.5005
R324 CSoutput.n191 CSoutput.n183 4.5005
R325 CSoutput.n186 CSoutput.n183 4.5005
R326 CSoutput.t136 CSoutput.n183 4.5005
R327 CSoutput.n185 CSoutput.n183 4.5005
R328 CSoutput.n192 CSoutput.n183 4.5005
R329 CSoutput.n244 CSoutput.n188 4.5005
R330 CSoutput.n244 CSoutput.n190 4.5005
R331 CSoutput.n244 CSoutput.n187 4.5005
R332 CSoutput.n244 CSoutput.n191 4.5005
R333 CSoutput.n244 CSoutput.n186 4.5005
R334 CSoutput.n244 CSoutput.t136 4.5005
R335 CSoutput.n244 CSoutput.n185 4.5005
R336 CSoutput.n244 CSoutput.n192 4.5005
R337 CSoutput.n242 CSoutput.n188 4.5005
R338 CSoutput.n242 CSoutput.n190 4.5005
R339 CSoutput.n242 CSoutput.n187 4.5005
R340 CSoutput.n242 CSoutput.n191 4.5005
R341 CSoutput.n242 CSoutput.n186 4.5005
R342 CSoutput.n242 CSoutput.t136 4.5005
R343 CSoutput.n242 CSoutput.n185 4.5005
R344 CSoutput.n242 CSoutput.n192 4.5005
R345 CSoutput.n242 CSoutput.n241 4.5005
R346 CSoutput.n224 CSoutput.n188 4.5005
R347 CSoutput.n224 CSoutput.n190 4.5005
R348 CSoutput.n224 CSoutput.n187 4.5005
R349 CSoutput.n224 CSoutput.n191 4.5005
R350 CSoutput.n224 CSoutput.n186 4.5005
R351 CSoutput.n224 CSoutput.t136 4.5005
R352 CSoutput.n224 CSoutput.n185 4.5005
R353 CSoutput.n224 CSoutput.n192 4.5005
R354 CSoutput.n241 CSoutput.n224 4.5005
R355 CSoutput.n196 CSoutput.n188 4.5005
R356 CSoutput.n196 CSoutput.n190 4.5005
R357 CSoutput.n196 CSoutput.n187 4.5005
R358 CSoutput.n196 CSoutput.n191 4.5005
R359 CSoutput.n196 CSoutput.n186 4.5005
R360 CSoutput.n196 CSoutput.t136 4.5005
R361 CSoutput.n196 CSoutput.n185 4.5005
R362 CSoutput.n196 CSoutput.n192 4.5005
R363 CSoutput.n241 CSoutput.n196 4.5005
R364 CSoutput.n226 CSoutput.n188 4.5005
R365 CSoutput.n226 CSoutput.n190 4.5005
R366 CSoutput.n226 CSoutput.n187 4.5005
R367 CSoutput.n226 CSoutput.n191 4.5005
R368 CSoutput.n226 CSoutput.n186 4.5005
R369 CSoutput.n226 CSoutput.t136 4.5005
R370 CSoutput.n226 CSoutput.n185 4.5005
R371 CSoutput.n226 CSoutput.n192 4.5005
R372 CSoutput.n241 CSoutput.n226 4.5005
R373 CSoutput.n195 CSoutput.n188 4.5005
R374 CSoutput.n195 CSoutput.n190 4.5005
R375 CSoutput.n195 CSoutput.n187 4.5005
R376 CSoutput.n195 CSoutput.n191 4.5005
R377 CSoutput.n195 CSoutput.n186 4.5005
R378 CSoutput.n195 CSoutput.t136 4.5005
R379 CSoutput.n195 CSoutput.n185 4.5005
R380 CSoutput.n195 CSoutput.n192 4.5005
R381 CSoutput.n241 CSoutput.n195 4.5005
R382 CSoutput.n240 CSoutput.n188 4.5005
R383 CSoutput.n240 CSoutput.n190 4.5005
R384 CSoutput.n240 CSoutput.n187 4.5005
R385 CSoutput.n240 CSoutput.n191 4.5005
R386 CSoutput.n240 CSoutput.n186 4.5005
R387 CSoutput.n240 CSoutput.t136 4.5005
R388 CSoutput.n240 CSoutput.n185 4.5005
R389 CSoutput.n240 CSoutput.n192 4.5005
R390 CSoutput.n241 CSoutput.n240 4.5005
R391 CSoutput.n239 CSoutput.n124 4.5005
R392 CSoutput.n140 CSoutput.n124 4.5005
R393 CSoutput.n135 CSoutput.n119 4.5005
R394 CSoutput.n135 CSoutput.n121 4.5005
R395 CSoutput.n135 CSoutput.n118 4.5005
R396 CSoutput.n135 CSoutput.n122 4.5005
R397 CSoutput.n135 CSoutput.n117 4.5005
R398 CSoutput.n135 CSoutput.t144 4.5005
R399 CSoutput.n135 CSoutput.n116 4.5005
R400 CSoutput.n135 CSoutput.n123 4.5005
R401 CSoutput.n135 CSoutput.n124 4.5005
R402 CSoutput.n133 CSoutput.n119 4.5005
R403 CSoutput.n133 CSoutput.n121 4.5005
R404 CSoutput.n133 CSoutput.n118 4.5005
R405 CSoutput.n133 CSoutput.n122 4.5005
R406 CSoutput.n133 CSoutput.n117 4.5005
R407 CSoutput.n133 CSoutput.t144 4.5005
R408 CSoutput.n133 CSoutput.n116 4.5005
R409 CSoutput.n133 CSoutput.n123 4.5005
R410 CSoutput.n133 CSoutput.n124 4.5005
R411 CSoutput.n132 CSoutput.n119 4.5005
R412 CSoutput.n132 CSoutput.n121 4.5005
R413 CSoutput.n132 CSoutput.n118 4.5005
R414 CSoutput.n132 CSoutput.n122 4.5005
R415 CSoutput.n132 CSoutput.n117 4.5005
R416 CSoutput.n132 CSoutput.t144 4.5005
R417 CSoutput.n132 CSoutput.n116 4.5005
R418 CSoutput.n132 CSoutput.n123 4.5005
R419 CSoutput.n132 CSoutput.n124 4.5005
R420 CSoutput.n261 CSoutput.n119 4.5005
R421 CSoutput.n261 CSoutput.n121 4.5005
R422 CSoutput.n261 CSoutput.n118 4.5005
R423 CSoutput.n261 CSoutput.n122 4.5005
R424 CSoutput.n261 CSoutput.n117 4.5005
R425 CSoutput.n261 CSoutput.t144 4.5005
R426 CSoutput.n261 CSoutput.n116 4.5005
R427 CSoutput.n261 CSoutput.n123 4.5005
R428 CSoutput.n261 CSoutput.n124 4.5005
R429 CSoutput.n259 CSoutput.n119 4.5005
R430 CSoutput.n259 CSoutput.n121 4.5005
R431 CSoutput.n259 CSoutput.n118 4.5005
R432 CSoutput.n259 CSoutput.n122 4.5005
R433 CSoutput.n259 CSoutput.n117 4.5005
R434 CSoutput.n259 CSoutput.t144 4.5005
R435 CSoutput.n259 CSoutput.n116 4.5005
R436 CSoutput.n259 CSoutput.n123 4.5005
R437 CSoutput.n257 CSoutput.n119 4.5005
R438 CSoutput.n257 CSoutput.n121 4.5005
R439 CSoutput.n257 CSoutput.n118 4.5005
R440 CSoutput.n257 CSoutput.n122 4.5005
R441 CSoutput.n257 CSoutput.n117 4.5005
R442 CSoutput.n257 CSoutput.t144 4.5005
R443 CSoutput.n257 CSoutput.n116 4.5005
R444 CSoutput.n257 CSoutput.n123 4.5005
R445 CSoutput.n143 CSoutput.n119 4.5005
R446 CSoutput.n143 CSoutput.n121 4.5005
R447 CSoutput.n143 CSoutput.n118 4.5005
R448 CSoutput.n143 CSoutput.n122 4.5005
R449 CSoutput.n143 CSoutput.n117 4.5005
R450 CSoutput.n143 CSoutput.t144 4.5005
R451 CSoutput.n143 CSoutput.n116 4.5005
R452 CSoutput.n143 CSoutput.n123 4.5005
R453 CSoutput.n143 CSoutput.n124 4.5005
R454 CSoutput.n142 CSoutput.n119 4.5005
R455 CSoutput.n142 CSoutput.n121 4.5005
R456 CSoutput.n142 CSoutput.n118 4.5005
R457 CSoutput.n142 CSoutput.n122 4.5005
R458 CSoutput.n142 CSoutput.n117 4.5005
R459 CSoutput.n142 CSoutput.t144 4.5005
R460 CSoutput.n142 CSoutput.n116 4.5005
R461 CSoutput.n142 CSoutput.n123 4.5005
R462 CSoutput.n142 CSoutput.n124 4.5005
R463 CSoutput.n146 CSoutput.n119 4.5005
R464 CSoutput.n146 CSoutput.n121 4.5005
R465 CSoutput.n146 CSoutput.n118 4.5005
R466 CSoutput.n146 CSoutput.n122 4.5005
R467 CSoutput.n146 CSoutput.n117 4.5005
R468 CSoutput.n146 CSoutput.t144 4.5005
R469 CSoutput.n146 CSoutput.n116 4.5005
R470 CSoutput.n146 CSoutput.n123 4.5005
R471 CSoutput.n146 CSoutput.n124 4.5005
R472 CSoutput.n145 CSoutput.n119 4.5005
R473 CSoutput.n145 CSoutput.n121 4.5005
R474 CSoutput.n145 CSoutput.n118 4.5005
R475 CSoutput.n145 CSoutput.n122 4.5005
R476 CSoutput.n145 CSoutput.n117 4.5005
R477 CSoutput.n145 CSoutput.t144 4.5005
R478 CSoutput.n145 CSoutput.n116 4.5005
R479 CSoutput.n145 CSoutput.n123 4.5005
R480 CSoutput.n145 CSoutput.n124 4.5005
R481 CSoutput.n128 CSoutput.n119 4.5005
R482 CSoutput.n128 CSoutput.n121 4.5005
R483 CSoutput.n128 CSoutput.n118 4.5005
R484 CSoutput.n128 CSoutput.n122 4.5005
R485 CSoutput.n128 CSoutput.n117 4.5005
R486 CSoutput.n128 CSoutput.t144 4.5005
R487 CSoutput.n128 CSoutput.n116 4.5005
R488 CSoutput.n128 CSoutput.n123 4.5005
R489 CSoutput.n128 CSoutput.n124 4.5005
R490 CSoutput.n264 CSoutput.n119 4.5005
R491 CSoutput.n264 CSoutput.n121 4.5005
R492 CSoutput.n264 CSoutput.n118 4.5005
R493 CSoutput.n264 CSoutput.n122 4.5005
R494 CSoutput.n264 CSoutput.n117 4.5005
R495 CSoutput.n264 CSoutput.t144 4.5005
R496 CSoutput.n264 CSoutput.n116 4.5005
R497 CSoutput.n264 CSoutput.n123 4.5005
R498 CSoutput.n264 CSoutput.n124 4.5005
R499 CSoutput.n299 CSoutput.n287 4.10845
R500 CSoutput.n113 CSoutput.n101 4.10845
R501 CSoutput.n297 CSoutput.t62 4.06363
R502 CSoutput.n297 CSoutput.t116 4.06363
R503 CSoutput.n295 CSoutput.t73 4.06363
R504 CSoutput.n295 CSoutput.t83 4.06363
R505 CSoutput.n293 CSoutput.t60 4.06363
R506 CSoutput.n293 CSoutput.t75 4.06363
R507 CSoutput.n291 CSoutput.t49 4.06363
R508 CSoutput.n291 CSoutput.t110 4.06363
R509 CSoutput.n289 CSoutput.t52 4.06363
R510 CSoutput.n289 CSoutput.t94 4.06363
R511 CSoutput.n288 CSoutput.t37 4.06363
R512 CSoutput.n288 CSoutput.t36 4.06363
R513 CSoutput.n285 CSoutput.t11 4.06363
R514 CSoutput.n285 CSoutput.t10 4.06363
R515 CSoutput.n283 CSoutput.t132 4.06363
R516 CSoutput.n283 CSoutput.t78 4.06363
R517 CSoutput.n281 CSoutput.t84 4.06363
R518 CSoutput.n281 CSoutput.t133 4.06363
R519 CSoutput.n279 CSoutput.t30 4.06363
R520 CSoutput.n279 CSoutput.t101 4.06363
R521 CSoutput.n277 CSoutput.t100 4.06363
R522 CSoutput.n277 CSoutput.t8 4.06363
R523 CSoutput.n276 CSoutput.t69 4.06363
R524 CSoutput.n276 CSoutput.t135 4.06363
R525 CSoutput.n274 CSoutput.t96 4.06363
R526 CSoutput.n274 CSoutput.t34 4.06363
R527 CSoutput.n272 CSoutput.t21 4.06363
R528 CSoutput.n272 CSoutput.t32 4.06363
R529 CSoutput.n270 CSoutput.t76 4.06363
R530 CSoutput.n270 CSoutput.t80 4.06363
R531 CSoutput.n268 CSoutput.t89 4.06363
R532 CSoutput.n268 CSoutput.t109 4.06363
R533 CSoutput.n266 CSoutput.t70 4.06363
R534 CSoutput.n266 CSoutput.t82 4.06363
R535 CSoutput.n265 CSoutput.t12 4.06363
R536 CSoutput.n265 CSoutput.t86 4.06363
R537 CSoutput.n102 CSoutput.t126 4.06363
R538 CSoutput.n102 CSoutput.t125 4.06363
R539 CSoutput.n103 CSoutput.t23 4.06363
R540 CSoutput.n103 CSoutput.t48 4.06363
R541 CSoutput.n105 CSoutput.t95 4.06363
R542 CSoutput.n105 CSoutput.t104 4.06363
R543 CSoutput.n107 CSoutput.t24 4.06363
R544 CSoutput.n107 CSoutput.t134 4.06363
R545 CSoutput.n109 CSoutput.t63 4.06363
R546 CSoutput.n109 CSoutput.t85 4.06363
R547 CSoutput.n111 CSoutput.t107 4.06363
R548 CSoutput.n111 CSoutput.t108 4.06363
R549 CSoutput.n90 CSoutput.t87 4.06363
R550 CSoutput.n90 CSoutput.t53 4.06363
R551 CSoutput.n91 CSoutput.t71 4.06363
R552 CSoutput.n91 CSoutput.t35 4.06363
R553 CSoutput.n93 CSoutput.t9 4.06363
R554 CSoutput.n93 CSoutput.t103 4.06363
R555 CSoutput.n95 CSoutput.t72 4.06363
R556 CSoutput.n95 CSoutput.t74 4.06363
R557 CSoutput.n97 CSoutput.t88 4.06363
R558 CSoutput.n97 CSoutput.t105 4.06363
R559 CSoutput.n99 CSoutput.t98 4.06363
R560 CSoutput.n99 CSoutput.t99 4.06363
R561 CSoutput.n79 CSoutput.t79 4.06363
R562 CSoutput.n79 CSoutput.t13 4.06363
R563 CSoutput.n80 CSoutput.t22 4.06363
R564 CSoutput.n80 CSoutput.t29 4.06363
R565 CSoutput.n82 CSoutput.t102 4.06363
R566 CSoutput.n82 CSoutput.t47 4.06363
R567 CSoutput.n84 CSoutput.t81 4.06363
R568 CSoutput.n84 CSoutput.t115 4.06363
R569 CSoutput.n86 CSoutput.t33 4.06363
R570 CSoutput.n86 CSoutput.t50 4.06363
R571 CSoutput.n88 CSoutput.t61 4.06363
R572 CSoutput.n88 CSoutput.t97 4.06363
R573 CSoutput.n44 CSoutput.n43 3.79402
R574 CSoutput.n49 CSoutput.n48 3.79402
R575 CSoutput.n365 CSoutput.n364 3.57343
R576 CSoutput.n364 CSoutput.n332 3.08965
R577 CSoutput.n329 CSoutput.t65 2.82907
R578 CSoutput.n329 CSoutput.t2 2.82907
R579 CSoutput.n327 CSoutput.t112 2.82907
R580 CSoutput.n327 CSoutput.t123 2.82907
R581 CSoutput.n325 CSoutput.t120 2.82907
R582 CSoutput.n325 CSoutput.t119 2.82907
R583 CSoutput.n323 CSoutput.t31 2.82907
R584 CSoutput.n323 CSoutput.t44 2.82907
R585 CSoutput.n321 CSoutput.t55 2.82907
R586 CSoutput.n321 CSoutput.t20 2.82907
R587 CSoutput.n319 CSoutput.t40 2.82907
R588 CSoutput.n319 CSoutput.t14 2.82907
R589 CSoutput.n317 CSoutput.t106 2.82907
R590 CSoutput.n317 CSoutput.t7 2.82907
R591 CSoutput.n316 CSoutput.t57 2.82907
R592 CSoutput.n316 CSoutput.t56 2.82907
R593 CSoutput.n314 CSoutput.t58 2.82907
R594 CSoutput.n314 CSoutput.t127 2.82907
R595 CSoutput.n312 CSoutput.t117 2.82907
R596 CSoutput.n312 CSoutput.t6 2.82907
R597 CSoutput.n310 CSoutput.t122 2.82907
R598 CSoutput.n310 CSoutput.t124 2.82907
R599 CSoutput.n308 CSoutput.t45 2.82907
R600 CSoutput.n308 CSoutput.t118 2.82907
R601 CSoutput.n306 CSoutput.t27 2.82907
R602 CSoutput.n306 CSoutput.t77 2.82907
R603 CSoutput.n304 CSoutput.t0 2.82907
R604 CSoutput.n304 CSoutput.t64 2.82907
R605 CSoutput.n302 CSoutput.t111 2.82907
R606 CSoutput.n302 CSoutput.t92 2.82907
R607 CSoutput.n301 CSoutput.t46 2.82907
R608 CSoutput.n301 CSoutput.t38 2.82907
R609 CSoutput.n348 CSoutput.t28 2.82907
R610 CSoutput.n348 CSoutput.t51 2.82907
R611 CSoutput.n349 CSoutput.t66 2.82907
R612 CSoutput.n349 CSoutput.t43 2.82907
R613 CSoutput.n351 CSoutput.t68 2.82907
R614 CSoutput.n351 CSoutput.t25 2.82907
R615 CSoutput.n353 CSoutput.t131 2.82907
R616 CSoutput.n353 CSoutput.t59 2.82907
R617 CSoutput.n355 CSoutput.t26 2.82907
R618 CSoutput.n355 CSoutput.t17 2.82907
R619 CSoutput.n357 CSoutput.t18 2.82907
R620 CSoutput.n357 CSoutput.t41 2.82907
R621 CSoutput.n359 CSoutput.t93 2.82907
R622 CSoutput.n359 CSoutput.t90 2.82907
R623 CSoutput.n361 CSoutput.t15 2.82907
R624 CSoutput.n361 CSoutput.t3 2.82907
R625 CSoutput.n333 CSoutput.t42 2.82907
R626 CSoutput.n333 CSoutput.t67 2.82907
R627 CSoutput.n334 CSoutput.t4 2.82907
R628 CSoutput.n334 CSoutput.t114 2.82907
R629 CSoutput.n336 CSoutput.t19 2.82907
R630 CSoutput.n336 CSoutput.t54 2.82907
R631 CSoutput.n338 CSoutput.t121 2.82907
R632 CSoutput.n338 CSoutput.t1 2.82907
R633 CSoutput.n340 CSoutput.t130 2.82907
R634 CSoutput.n340 CSoutput.t16 2.82907
R635 CSoutput.n342 CSoutput.t91 2.82907
R636 CSoutput.n342 CSoutput.t128 2.82907
R637 CSoutput.n344 CSoutput.t5 2.82907
R638 CSoutput.n344 CSoutput.t113 2.82907
R639 CSoutput.n346 CSoutput.t39 2.82907
R640 CSoutput.n346 CSoutput.t129 2.82907
R641 CSoutput.n75 CSoutput.n1 2.45513
R642 CSoutput.n205 CSoutput.n203 2.251
R643 CSoutput.n205 CSoutput.n202 2.251
R644 CSoutput.n205 CSoutput.n201 2.251
R645 CSoutput.n205 CSoutput.n200 2.251
R646 CSoutput.n174 CSoutput.n173 2.251
R647 CSoutput.n174 CSoutput.n172 2.251
R648 CSoutput.n174 CSoutput.n171 2.251
R649 CSoutput.n174 CSoutput.n170 2.251
R650 CSoutput.n247 CSoutput.n246 2.251
R651 CSoutput.n212 CSoutput.n210 2.251
R652 CSoutput.n212 CSoutput.n209 2.251
R653 CSoutput.n212 CSoutput.n208 2.251
R654 CSoutput.n230 CSoutput.n212 2.251
R655 CSoutput.n218 CSoutput.n217 2.251
R656 CSoutput.n218 CSoutput.n216 2.251
R657 CSoutput.n218 CSoutput.n215 2.251
R658 CSoutput.n218 CSoutput.n214 2.251
R659 CSoutput.n244 CSoutput.n184 2.251
R660 CSoutput.n239 CSoutput.n237 2.251
R661 CSoutput.n239 CSoutput.n236 2.251
R662 CSoutput.n239 CSoutput.n235 2.251
R663 CSoutput.n239 CSoutput.n234 2.251
R664 CSoutput.n140 CSoutput.n139 2.251
R665 CSoutput.n140 CSoutput.n138 2.251
R666 CSoutput.n140 CSoutput.n137 2.251
R667 CSoutput.n140 CSoutput.n136 2.251
R668 CSoutput.n257 CSoutput.n256 2.251
R669 CSoutput.n174 CSoutput.n154 2.2505
R670 CSoutput.n169 CSoutput.n154 2.2505
R671 CSoutput.n167 CSoutput.n154 2.2505
R672 CSoutput.n166 CSoutput.n154 2.2505
R673 CSoutput.n251 CSoutput.n154 2.2505
R674 CSoutput.n249 CSoutput.n154 2.2505
R675 CSoutput.n247 CSoutput.n154 2.2505
R676 CSoutput.n177 CSoutput.n154 2.2505
R677 CSoutput.n176 CSoutput.n154 2.2505
R678 CSoutput.n180 CSoutput.n154 2.2505
R679 CSoutput.n179 CSoutput.n154 2.2505
R680 CSoutput.n162 CSoutput.n154 2.2505
R681 CSoutput.n254 CSoutput.n154 2.2505
R682 CSoutput.n254 CSoutput.n253 2.2505
R683 CSoutput.n218 CSoutput.n189 2.2505
R684 CSoutput.n199 CSoutput.n189 2.2505
R685 CSoutput.n220 CSoutput.n189 2.2505
R686 CSoutput.n198 CSoutput.n189 2.2505
R687 CSoutput.n222 CSoutput.n189 2.2505
R688 CSoutput.n189 CSoutput.n183 2.2505
R689 CSoutput.n244 CSoutput.n189 2.2505
R690 CSoutput.n242 CSoutput.n189 2.2505
R691 CSoutput.n224 CSoutput.n189 2.2505
R692 CSoutput.n196 CSoutput.n189 2.2505
R693 CSoutput.n226 CSoutput.n189 2.2505
R694 CSoutput.n195 CSoutput.n189 2.2505
R695 CSoutput.n240 CSoutput.n189 2.2505
R696 CSoutput.n240 CSoutput.n193 2.2505
R697 CSoutput.n140 CSoutput.n120 2.2505
R698 CSoutput.n135 CSoutput.n120 2.2505
R699 CSoutput.n133 CSoutput.n120 2.2505
R700 CSoutput.n132 CSoutput.n120 2.2505
R701 CSoutput.n261 CSoutput.n120 2.2505
R702 CSoutput.n259 CSoutput.n120 2.2505
R703 CSoutput.n257 CSoutput.n120 2.2505
R704 CSoutput.n143 CSoutput.n120 2.2505
R705 CSoutput.n142 CSoutput.n120 2.2505
R706 CSoutput.n146 CSoutput.n120 2.2505
R707 CSoutput.n145 CSoutput.n120 2.2505
R708 CSoutput.n128 CSoutput.n120 2.2505
R709 CSoutput.n264 CSoutput.n120 2.2505
R710 CSoutput.n264 CSoutput.n263 2.2505
R711 CSoutput.n182 CSoutput.n175 2.25024
R712 CSoutput.n182 CSoutput.n168 2.25024
R713 CSoutput.n250 CSoutput.n182 2.25024
R714 CSoutput.n182 CSoutput.n178 2.25024
R715 CSoutput.n182 CSoutput.n181 2.25024
R716 CSoutput.n182 CSoutput.n149 2.25024
R717 CSoutput.n232 CSoutput.n229 2.25024
R718 CSoutput.n232 CSoutput.n228 2.25024
R719 CSoutput.n232 CSoutput.n227 2.25024
R720 CSoutput.n232 CSoutput.n194 2.25024
R721 CSoutput.n232 CSoutput.n231 2.25024
R722 CSoutput.n233 CSoutput.n232 2.25024
R723 CSoutput.n148 CSoutput.n141 2.25024
R724 CSoutput.n148 CSoutput.n134 2.25024
R725 CSoutput.n260 CSoutput.n148 2.25024
R726 CSoutput.n148 CSoutput.n144 2.25024
R727 CSoutput.n148 CSoutput.n147 2.25024
R728 CSoutput.n148 CSoutput.n115 2.25024
R729 CSoutput.n300 CSoutput.n114 2.15937
R730 CSoutput.n249 CSoutput.n159 1.50111
R731 CSoutput.n197 CSoutput.n183 1.50111
R732 CSoutput.n259 CSoutput.n125 1.50111
R733 CSoutput.n205 CSoutput.n204 1.501
R734 CSoutput.n212 CSoutput.n211 1.501
R735 CSoutput.n239 CSoutput.n238 1.501
R736 CSoutput.n253 CSoutput.n164 1.12536
R737 CSoutput.n253 CSoutput.n165 1.12536
R738 CSoutput.n253 CSoutput.n252 1.12536
R739 CSoutput.n213 CSoutput.n193 1.12536
R740 CSoutput.n219 CSoutput.n193 1.12536
R741 CSoutput.n221 CSoutput.n193 1.12536
R742 CSoutput.n263 CSoutput.n130 1.12536
R743 CSoutput.n263 CSoutput.n131 1.12536
R744 CSoutput.n263 CSoutput.n262 1.12536
R745 CSoutput.n253 CSoutput.n160 1.12536
R746 CSoutput.n253 CSoutput.n161 1.12536
R747 CSoutput.n253 CSoutput.n163 1.12536
R748 CSoutput.n243 CSoutput.n193 1.12536
R749 CSoutput.n223 CSoutput.n193 1.12536
R750 CSoutput.n225 CSoutput.n193 1.12536
R751 CSoutput.n263 CSoutput.n126 1.12536
R752 CSoutput.n263 CSoutput.n127 1.12536
R753 CSoutput.n263 CSoutput.n129 1.12536
R754 CSoutput.n31 CSoutput.n30 0.669944
R755 CSoutput.n62 CSoutput.n61 0.669944
R756 CSoutput.n320 CSoutput.n318 0.573776
R757 CSoutput.n322 CSoutput.n320 0.573776
R758 CSoutput.n324 CSoutput.n322 0.573776
R759 CSoutput.n326 CSoutput.n324 0.573776
R760 CSoutput.n328 CSoutput.n326 0.573776
R761 CSoutput.n330 CSoutput.n328 0.573776
R762 CSoutput.n305 CSoutput.n303 0.573776
R763 CSoutput.n307 CSoutput.n305 0.573776
R764 CSoutput.n309 CSoutput.n307 0.573776
R765 CSoutput.n311 CSoutput.n309 0.573776
R766 CSoutput.n313 CSoutput.n311 0.573776
R767 CSoutput.n315 CSoutput.n313 0.573776
R768 CSoutput.n362 CSoutput.n360 0.573776
R769 CSoutput.n360 CSoutput.n358 0.573776
R770 CSoutput.n358 CSoutput.n356 0.573776
R771 CSoutput.n356 CSoutput.n354 0.573776
R772 CSoutput.n354 CSoutput.n352 0.573776
R773 CSoutput.n352 CSoutput.n350 0.573776
R774 CSoutput.n347 CSoutput.n345 0.573776
R775 CSoutput.n345 CSoutput.n343 0.573776
R776 CSoutput.n343 CSoutput.n341 0.573776
R777 CSoutput.n341 CSoutput.n339 0.573776
R778 CSoutput.n339 CSoutput.n337 0.573776
R779 CSoutput.n337 CSoutput.n335 0.573776
R780 CSoutput.n365 CSoutput.n264 0.53442
R781 CSoutput.n292 CSoutput.n290 0.358259
R782 CSoutput.n294 CSoutput.n292 0.358259
R783 CSoutput.n296 CSoutput.n294 0.358259
R784 CSoutput.n298 CSoutput.n296 0.358259
R785 CSoutput.n280 CSoutput.n278 0.358259
R786 CSoutput.n282 CSoutput.n280 0.358259
R787 CSoutput.n284 CSoutput.n282 0.358259
R788 CSoutput.n286 CSoutput.n284 0.358259
R789 CSoutput.n269 CSoutput.n267 0.358259
R790 CSoutput.n271 CSoutput.n269 0.358259
R791 CSoutput.n273 CSoutput.n271 0.358259
R792 CSoutput.n275 CSoutput.n273 0.358259
R793 CSoutput.n112 CSoutput.n110 0.358259
R794 CSoutput.n110 CSoutput.n108 0.358259
R795 CSoutput.n108 CSoutput.n106 0.358259
R796 CSoutput.n106 CSoutput.n104 0.358259
R797 CSoutput.n100 CSoutput.n98 0.358259
R798 CSoutput.n98 CSoutput.n96 0.358259
R799 CSoutput.n96 CSoutput.n94 0.358259
R800 CSoutput.n94 CSoutput.n92 0.358259
R801 CSoutput.n89 CSoutput.n87 0.358259
R802 CSoutput.n87 CSoutput.n85 0.358259
R803 CSoutput.n85 CSoutput.n83 0.358259
R804 CSoutput.n83 CSoutput.n81 0.358259
R805 CSoutput.n21 CSoutput.n20 0.169105
R806 CSoutput.n21 CSoutput.n16 0.169105
R807 CSoutput.n26 CSoutput.n16 0.169105
R808 CSoutput.n27 CSoutput.n26 0.169105
R809 CSoutput.n27 CSoutput.n14 0.169105
R810 CSoutput.n32 CSoutput.n14 0.169105
R811 CSoutput.n33 CSoutput.n32 0.169105
R812 CSoutput.n34 CSoutput.n33 0.169105
R813 CSoutput.n34 CSoutput.n12 0.169105
R814 CSoutput.n39 CSoutput.n12 0.169105
R815 CSoutput.n40 CSoutput.n39 0.169105
R816 CSoutput.n40 CSoutput.n10 0.169105
R817 CSoutput.n45 CSoutput.n10 0.169105
R818 CSoutput.n46 CSoutput.n45 0.169105
R819 CSoutput.n47 CSoutput.n46 0.169105
R820 CSoutput.n47 CSoutput.n8 0.169105
R821 CSoutput.n52 CSoutput.n8 0.169105
R822 CSoutput.n53 CSoutput.n52 0.169105
R823 CSoutput.n53 CSoutput.n6 0.169105
R824 CSoutput.n58 CSoutput.n6 0.169105
R825 CSoutput.n59 CSoutput.n58 0.169105
R826 CSoutput.n60 CSoutput.n59 0.169105
R827 CSoutput.n60 CSoutput.n4 0.169105
R828 CSoutput.n66 CSoutput.n4 0.169105
R829 CSoutput.n67 CSoutput.n66 0.169105
R830 CSoutput.n68 CSoutput.n67 0.169105
R831 CSoutput.n68 CSoutput.n2 0.169105
R832 CSoutput.n73 CSoutput.n2 0.169105
R833 CSoutput.n74 CSoutput.n73 0.169105
R834 CSoutput.n74 CSoutput.n0 0.169105
R835 CSoutput.n78 CSoutput.n0 0.169105
R836 CSoutput.n207 CSoutput.n206 0.0910737
R837 CSoutput.n258 CSoutput.n255 0.0723685
R838 CSoutput.n212 CSoutput.n207 0.0522944
R839 CSoutput.n255 CSoutput.n254 0.0499135
R840 CSoutput.n206 CSoutput.n205 0.0499135
R841 CSoutput.n240 CSoutput.n239 0.0464294
R842 CSoutput.n248 CSoutput.n245 0.0391444
R843 CSoutput.n207 CSoutput.t145 0.023435
R844 CSoutput.n255 CSoutput.t139 0.02262
R845 CSoutput.n206 CSoutput.t143 0.02262
R846 CSoutput CSoutput.n365 0.0052
R847 CSoutput.n177 CSoutput.n160 0.00365111
R848 CSoutput.n180 CSoutput.n161 0.00365111
R849 CSoutput.n163 CSoutput.n162 0.00365111
R850 CSoutput.n205 CSoutput.n164 0.00365111
R851 CSoutput.n169 CSoutput.n165 0.00365111
R852 CSoutput.n252 CSoutput.n166 0.00365111
R853 CSoutput.n243 CSoutput.n242 0.00365111
R854 CSoutput.n223 CSoutput.n196 0.00365111
R855 CSoutput.n225 CSoutput.n195 0.00365111
R856 CSoutput.n213 CSoutput.n212 0.00365111
R857 CSoutput.n219 CSoutput.n199 0.00365111
R858 CSoutput.n221 CSoutput.n198 0.00365111
R859 CSoutput.n143 CSoutput.n126 0.00365111
R860 CSoutput.n146 CSoutput.n127 0.00365111
R861 CSoutput.n129 CSoutput.n128 0.00365111
R862 CSoutput.n239 CSoutput.n130 0.00365111
R863 CSoutput.n135 CSoutput.n131 0.00365111
R864 CSoutput.n262 CSoutput.n132 0.00365111
R865 CSoutput.n174 CSoutput.n164 0.00340054
R866 CSoutput.n167 CSoutput.n165 0.00340054
R867 CSoutput.n252 CSoutput.n251 0.00340054
R868 CSoutput.n247 CSoutput.n160 0.00340054
R869 CSoutput.n176 CSoutput.n161 0.00340054
R870 CSoutput.n179 CSoutput.n163 0.00340054
R871 CSoutput.n218 CSoutput.n213 0.00340054
R872 CSoutput.n220 CSoutput.n219 0.00340054
R873 CSoutput.n222 CSoutput.n221 0.00340054
R874 CSoutput.n244 CSoutput.n243 0.00340054
R875 CSoutput.n224 CSoutput.n223 0.00340054
R876 CSoutput.n226 CSoutput.n225 0.00340054
R877 CSoutput.n140 CSoutput.n130 0.00340054
R878 CSoutput.n133 CSoutput.n131 0.00340054
R879 CSoutput.n262 CSoutput.n261 0.00340054
R880 CSoutput.n257 CSoutput.n126 0.00340054
R881 CSoutput.n142 CSoutput.n127 0.00340054
R882 CSoutput.n145 CSoutput.n129 0.00340054
R883 CSoutput.n175 CSoutput.n169 0.00252698
R884 CSoutput.n168 CSoutput.n166 0.00252698
R885 CSoutput.n250 CSoutput.n249 0.00252698
R886 CSoutput.n178 CSoutput.n176 0.00252698
R887 CSoutput.n181 CSoutput.n179 0.00252698
R888 CSoutput.n254 CSoutput.n149 0.00252698
R889 CSoutput.n175 CSoutput.n174 0.00252698
R890 CSoutput.n168 CSoutput.n167 0.00252698
R891 CSoutput.n251 CSoutput.n250 0.00252698
R892 CSoutput.n178 CSoutput.n177 0.00252698
R893 CSoutput.n181 CSoutput.n180 0.00252698
R894 CSoutput.n162 CSoutput.n149 0.00252698
R895 CSoutput.n229 CSoutput.n199 0.00252698
R896 CSoutput.n228 CSoutput.n198 0.00252698
R897 CSoutput.n227 CSoutput.n183 0.00252698
R898 CSoutput.n224 CSoutput.n194 0.00252698
R899 CSoutput.n231 CSoutput.n226 0.00252698
R900 CSoutput.n240 CSoutput.n233 0.00252698
R901 CSoutput.n229 CSoutput.n218 0.00252698
R902 CSoutput.n228 CSoutput.n220 0.00252698
R903 CSoutput.n227 CSoutput.n222 0.00252698
R904 CSoutput.n242 CSoutput.n194 0.00252698
R905 CSoutput.n231 CSoutput.n196 0.00252698
R906 CSoutput.n233 CSoutput.n195 0.00252698
R907 CSoutput.n141 CSoutput.n135 0.00252698
R908 CSoutput.n134 CSoutput.n132 0.00252698
R909 CSoutput.n260 CSoutput.n259 0.00252698
R910 CSoutput.n144 CSoutput.n142 0.00252698
R911 CSoutput.n147 CSoutput.n145 0.00252698
R912 CSoutput.n264 CSoutput.n115 0.00252698
R913 CSoutput.n141 CSoutput.n140 0.00252698
R914 CSoutput.n134 CSoutput.n133 0.00252698
R915 CSoutput.n261 CSoutput.n260 0.00252698
R916 CSoutput.n144 CSoutput.n143 0.00252698
R917 CSoutput.n147 CSoutput.n146 0.00252698
R918 CSoutput.n128 CSoutput.n115 0.00252698
R919 CSoutput.n249 CSoutput.n248 0.0020275
R920 CSoutput.n248 CSoutput.n247 0.0020275
R921 CSoutput.n245 CSoutput.n183 0.0020275
R922 CSoutput.n245 CSoutput.n244 0.0020275
R923 CSoutput.n259 CSoutput.n258 0.0020275
R924 CSoutput.n258 CSoutput.n257 0.0020275
R925 CSoutput.n159 CSoutput.n158 0.00166668
R926 CSoutput.n241 CSoutput.n197 0.00166668
R927 CSoutput.n125 CSoutput.n124 0.00166668
R928 CSoutput.n263 CSoutput.n125 0.00133328
R929 CSoutput.n197 CSoutput.n193 0.00133328
R930 CSoutput.n253 CSoutput.n159 0.00133328
R931 CSoutput.n256 CSoutput.n148 0.001
R932 CSoutput.n234 CSoutput.n148 0.001
R933 CSoutput.n136 CSoutput.n116 0.001
R934 CSoutput.n235 CSoutput.n116 0.001
R935 CSoutput.n137 CSoutput.n117 0.001
R936 CSoutput.n236 CSoutput.n117 0.001
R937 CSoutput.n138 CSoutput.n118 0.001
R938 CSoutput.n237 CSoutput.n118 0.001
R939 CSoutput.n139 CSoutput.n119 0.001
R940 CSoutput.n238 CSoutput.n119 0.001
R941 CSoutput.n232 CSoutput.n184 0.001
R942 CSoutput.n232 CSoutput.n230 0.001
R943 CSoutput.n214 CSoutput.n185 0.001
R944 CSoutput.n208 CSoutput.n185 0.001
R945 CSoutput.n215 CSoutput.n186 0.001
R946 CSoutput.n209 CSoutput.n186 0.001
R947 CSoutput.n216 CSoutput.n187 0.001
R948 CSoutput.n210 CSoutput.n187 0.001
R949 CSoutput.n217 CSoutput.n188 0.001
R950 CSoutput.n211 CSoutput.n188 0.001
R951 CSoutput.n246 CSoutput.n182 0.001
R952 CSoutput.n200 CSoutput.n182 0.001
R953 CSoutput.n170 CSoutput.n150 0.001
R954 CSoutput.n201 CSoutput.n150 0.001
R955 CSoutput.n171 CSoutput.n151 0.001
R956 CSoutput.n202 CSoutput.n151 0.001
R957 CSoutput.n172 CSoutput.n152 0.001
R958 CSoutput.n203 CSoutput.n152 0.001
R959 CSoutput.n173 CSoutput.n153 0.001
R960 CSoutput.n204 CSoutput.n153 0.001
R961 CSoutput.n204 CSoutput.n154 0.001
R962 CSoutput.n203 CSoutput.n155 0.001
R963 CSoutput.n202 CSoutput.n156 0.001
R964 CSoutput.n201 CSoutput.t156 0.001
R965 CSoutput.n200 CSoutput.n157 0.001
R966 CSoutput.n173 CSoutput.n155 0.001
R967 CSoutput.n172 CSoutput.n156 0.001
R968 CSoutput.n171 CSoutput.t156 0.001
R969 CSoutput.n170 CSoutput.n157 0.001
R970 CSoutput.n246 CSoutput.n158 0.001
R971 CSoutput.n211 CSoutput.n189 0.001
R972 CSoutput.n210 CSoutput.n190 0.001
R973 CSoutput.n209 CSoutput.n191 0.001
R974 CSoutput.n208 CSoutput.t136 0.001
R975 CSoutput.n230 CSoutput.n192 0.001
R976 CSoutput.n217 CSoutput.n190 0.001
R977 CSoutput.n216 CSoutput.n191 0.001
R978 CSoutput.n215 CSoutput.t136 0.001
R979 CSoutput.n214 CSoutput.n192 0.001
R980 CSoutput.n241 CSoutput.n184 0.001
R981 CSoutput.n238 CSoutput.n120 0.001
R982 CSoutput.n237 CSoutput.n121 0.001
R983 CSoutput.n236 CSoutput.n122 0.001
R984 CSoutput.n235 CSoutput.t144 0.001
R985 CSoutput.n234 CSoutput.n123 0.001
R986 CSoutput.n139 CSoutput.n121 0.001
R987 CSoutput.n138 CSoutput.n122 0.001
R988 CSoutput.n137 CSoutput.t144 0.001
R989 CSoutput.n136 CSoutput.n123 0.001
R990 CSoutput.n256 CSoutput.n124 0.001
R991 a_n1986_8322.n0 a_n1986_8322.t18 74.6477
R992 a_n1986_8322.n2 a_n1986_8322.t17 74.6477
R993 a_n1986_8322.n4 a_n1986_8322.t14 74.6474
R994 a_n1986_8322.n3 a_n1986_8322.t15 74.2899
R995 a_n1986_8322.n0 a_n1986_8322.t16 74.2899
R996 a_n1986_8322.n0 a_n1986_8322.t4 74.2899
R997 a_n1986_8322.n1 a_n1986_8322.t1 74.2899
R998 a_n1986_8322.n7 a_n1986_8322.t2 74.2899
R999 a_n1986_8322.n4 a_n1986_8322.n12 70.6783
R1000 a_n1986_8322.n0 a_n1986_8322.n8 70.6783
R1001 a_n1986_8322.n1 a_n1986_8322.n9 70.6783
R1002 a_n1986_8322.n2 a_n1986_8322.n5 70.6783
R1003 a_n1986_8322.n2 a_n1986_8322.n6 70.6783
R1004 a_n1986_8322.n13 a_n1986_8322.n4 70.6782
R1005 a_n1986_8322.n10 a_n1986_8322.n7 22.7556
R1006 a_n1986_8322.n11 a_n1986_8322.t19 9.96389
R1007 a_n1986_8322.n10 a_n1986_8322.n1 6.2408
R1008 a_n1986_8322.n3 a_n1986_8322.n11 5.83671
R1009 a_n1986_8322.n11 a_n1986_8322.n10 5.3452
R1010 a_n1986_8322.n12 a_n1986_8322.t7 3.61217
R1011 a_n1986_8322.n12 a_n1986_8322.t13 3.61217
R1012 a_n1986_8322.n8 a_n1986_8322.t11 3.61217
R1013 a_n1986_8322.n8 a_n1986_8322.t10 3.61217
R1014 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R1015 a_n1986_8322.n9 a_n1986_8322.t3 3.61217
R1016 a_n1986_8322.n5 a_n1986_8322.t20 3.61217
R1017 a_n1986_8322.n5 a_n1986_8322.t8 3.61217
R1018 a_n1986_8322.n6 a_n1986_8322.t6 3.61217
R1019 a_n1986_8322.n6 a_n1986_8322.t12 3.61217
R1020 a_n1986_8322.t0 a_n1986_8322.n13 3.61217
R1021 a_n1986_8322.n13 a_n1986_8322.t9 3.61217
R1022 a_n1986_8322.n1 a_n1986_8322.n0 1.17507
R1023 a_n1986_8322.n4 a_n1986_8322.n3 0.716017
R1024 a_n1986_8322.n7 a_n1986_8322.n2 0.716017
R1025 commonsourceibias.n35 commonsourceibias.t0 223.028
R1026 commonsourceibias.n128 commonsourceibias.t88 223.028
R1027 commonsourceibias.n217 commonsourceibias.t77 223.028
R1028 commonsourceibias.n364 commonsourceibias.t22 223.028
R1029 commonsourceibias.n305 commonsourceibias.t108 223.028
R1030 commonsourceibias.n499 commonsourceibias.t95 223.028
R1031 commonsourceibias.n99 commonsourceibias.t28 207.983
R1032 commonsourceibias.n192 commonsourceibias.t94 207.983
R1033 commonsourceibias.n281 commonsourceibias.t81 207.983
R1034 commonsourceibias.n430 commonsourceibias.t52 207.983
R1035 commonsourceibias.n476 commonsourceibias.t113 207.983
R1036 commonsourceibias.n565 commonsourceibias.t99 207.983
R1037 commonsourceibias.n97 commonsourceibias.t48 168.701
R1038 commonsourceibias.n91 commonsourceibias.t34 168.701
R1039 commonsourceibias.n17 commonsourceibias.t26 168.701
R1040 commonsourceibias.n83 commonsourceibias.t44 168.701
R1041 commonsourceibias.n77 commonsourceibias.t16 168.701
R1042 commonsourceibias.n22 commonsourceibias.t12 168.701
R1043 commonsourceibias.n69 commonsourceibias.t36 168.701
R1044 commonsourceibias.n63 commonsourceibias.t30 168.701
R1045 commonsourceibias.n25 commonsourceibias.t4 168.701
R1046 commonsourceibias.n27 commonsourceibias.t8 168.701
R1047 commonsourceibias.n29 commonsourceibias.t14 168.701
R1048 commonsourceibias.n46 commonsourceibias.t42 168.701
R1049 commonsourceibias.n40 commonsourceibias.t18 168.701
R1050 commonsourceibias.n34 commonsourceibias.t50 168.701
R1051 commonsourceibias.n190 commonsourceibias.t109 168.701
R1052 commonsourceibias.n184 commonsourceibias.t72 168.701
R1053 commonsourceibias.n5 commonsourceibias.t70 168.701
R1054 commonsourceibias.n176 commonsourceibias.t102 168.701
R1055 commonsourceibias.n170 commonsourceibias.t116 168.701
R1056 commonsourceibias.n10 commonsourceibias.t66 168.701
R1057 commonsourceibias.n162 commonsourceibias.t92 168.701
R1058 commonsourceibias.n156 commonsourceibias.t89 168.701
R1059 commonsourceibias.n118 commonsourceibias.t105 168.701
R1060 commonsourceibias.n120 commonsourceibias.t85 168.701
R1061 commonsourceibias.n122 commonsourceibias.t82 168.701
R1062 commonsourceibias.n139 commonsourceibias.t97 168.701
R1063 commonsourceibias.n133 commonsourceibias.t111 168.701
R1064 commonsourceibias.n127 commonsourceibias.t75 168.701
R1065 commonsourceibias.n216 commonsourceibias.t67 168.701
R1066 commonsourceibias.n222 commonsourceibias.t98 168.701
R1067 commonsourceibias.n228 commonsourceibias.t83 168.701
R1068 commonsourceibias.n211 commonsourceibias.t71 168.701
R1069 commonsourceibias.n209 commonsourceibias.t74 168.701
R1070 commonsourceibias.n207 commonsourceibias.t90 168.701
R1071 commonsourceibias.n245 commonsourceibias.t76 168.701
R1072 commonsourceibias.n251 commonsourceibias.t80 168.701
R1073 commonsourceibias.n204 commonsourceibias.t122 168.701
R1074 commonsourceibias.n259 commonsourceibias.t104 168.701
R1075 commonsourceibias.n265 commonsourceibias.t87 168.701
R1076 commonsourceibias.n199 commonsourceibias.t127 168.701
R1077 commonsourceibias.n273 commonsourceibias.t65 168.701
R1078 commonsourceibias.n279 commonsourceibias.t96 168.701
R1079 commonsourceibias.n363 commonsourceibias.t40 168.701
R1080 commonsourceibias.n369 commonsourceibias.t2 168.701
R1081 commonsourceibias.n375 commonsourceibias.t32 168.701
R1082 commonsourceibias.n358 commonsourceibias.t60 168.701
R1083 commonsourceibias.n356 commonsourceibias.t58 168.701
R1084 commonsourceibias.n354 commonsourceibias.t46 168.701
R1085 commonsourceibias.n392 commonsourceibias.t54 168.701
R1086 commonsourceibias.n398 commonsourceibias.t10 168.701
R1087 commonsourceibias.n400 commonsourceibias.t6 168.701
R1088 commonsourceibias.n407 commonsourceibias.t56 168.701
R1089 commonsourceibias.n413 commonsourceibias.t24 168.701
R1090 commonsourceibias.n415 commonsourceibias.t62 168.701
R1091 commonsourceibias.n422 commonsourceibias.t20 168.701
R1092 commonsourceibias.n428 commonsourceibias.t38 168.701
R1093 commonsourceibias.n474 commonsourceibias.t123 168.701
R1094 commonsourceibias.n468 commonsourceibias.t68 168.701
R1095 commonsourceibias.n461 commonsourceibias.t84 168.701
R1096 commonsourceibias.n459 commonsourceibias.t119 168.701
R1097 commonsourceibias.n453 commonsourceibias.t64 168.701
R1098 commonsourceibias.n446 commonsourceibias.t126 168.701
R1099 commonsourceibias.n444 commonsourceibias.t112 168.701
R1100 commonsourceibias.n304 commonsourceibias.t91 168.701
R1101 commonsourceibias.n310 commonsourceibias.t125 168.701
R1102 commonsourceibias.n316 commonsourceibias.t115 168.701
R1103 commonsourceibias.n299 commonsourceibias.t101 168.701
R1104 commonsourceibias.n297 commonsourceibias.t78 168.701
R1105 commonsourceibias.n295 commonsourceibias.t121 168.701
R1106 commonsourceibias.n333 commonsourceibias.t107 168.701
R1107 commonsourceibias.n498 commonsourceibias.t79 168.701
R1108 commonsourceibias.n504 commonsourceibias.t118 168.701
R1109 commonsourceibias.n510 commonsourceibias.t103 168.701
R1110 commonsourceibias.n493 commonsourceibias.t86 168.701
R1111 commonsourceibias.n491 commonsourceibias.t69 168.701
R1112 commonsourceibias.n489 commonsourceibias.t110 168.701
R1113 commonsourceibias.n527 commonsourceibias.t93 168.701
R1114 commonsourceibias.n533 commonsourceibias.t100 168.701
R1115 commonsourceibias.n535 commonsourceibias.t117 168.701
R1116 commonsourceibias.n542 commonsourceibias.t120 168.701
R1117 commonsourceibias.n548 commonsourceibias.t106 168.701
R1118 commonsourceibias.n550 commonsourceibias.t73 168.701
R1119 commonsourceibias.n557 commonsourceibias.t124 168.701
R1120 commonsourceibias.n563 commonsourceibias.t114 168.701
R1121 commonsourceibias.n36 commonsourceibias.n33 161.3
R1122 commonsourceibias.n38 commonsourceibias.n37 161.3
R1123 commonsourceibias.n39 commonsourceibias.n32 161.3
R1124 commonsourceibias.n42 commonsourceibias.n41 161.3
R1125 commonsourceibias.n43 commonsourceibias.n31 161.3
R1126 commonsourceibias.n45 commonsourceibias.n44 161.3
R1127 commonsourceibias.n47 commonsourceibias.n30 161.3
R1128 commonsourceibias.n49 commonsourceibias.n48 161.3
R1129 commonsourceibias.n51 commonsourceibias.n50 161.3
R1130 commonsourceibias.n52 commonsourceibias.n28 161.3
R1131 commonsourceibias.n54 commonsourceibias.n53 161.3
R1132 commonsourceibias.n56 commonsourceibias.n55 161.3
R1133 commonsourceibias.n57 commonsourceibias.n26 161.3
R1134 commonsourceibias.n59 commonsourceibias.n58 161.3
R1135 commonsourceibias.n61 commonsourceibias.n60 161.3
R1136 commonsourceibias.n62 commonsourceibias.n24 161.3
R1137 commonsourceibias.n65 commonsourceibias.n64 161.3
R1138 commonsourceibias.n66 commonsourceibias.n23 161.3
R1139 commonsourceibias.n68 commonsourceibias.n67 161.3
R1140 commonsourceibias.n70 commonsourceibias.n21 161.3
R1141 commonsourceibias.n72 commonsourceibias.n71 161.3
R1142 commonsourceibias.n73 commonsourceibias.n20 161.3
R1143 commonsourceibias.n75 commonsourceibias.n74 161.3
R1144 commonsourceibias.n76 commonsourceibias.n19 161.3
R1145 commonsourceibias.n79 commonsourceibias.n78 161.3
R1146 commonsourceibias.n80 commonsourceibias.n18 161.3
R1147 commonsourceibias.n82 commonsourceibias.n81 161.3
R1148 commonsourceibias.n84 commonsourceibias.n16 161.3
R1149 commonsourceibias.n86 commonsourceibias.n85 161.3
R1150 commonsourceibias.n87 commonsourceibias.n15 161.3
R1151 commonsourceibias.n89 commonsourceibias.n88 161.3
R1152 commonsourceibias.n90 commonsourceibias.n14 161.3
R1153 commonsourceibias.n93 commonsourceibias.n92 161.3
R1154 commonsourceibias.n94 commonsourceibias.n13 161.3
R1155 commonsourceibias.n96 commonsourceibias.n95 161.3
R1156 commonsourceibias.n98 commonsourceibias.n12 161.3
R1157 commonsourceibias.n129 commonsourceibias.n126 161.3
R1158 commonsourceibias.n131 commonsourceibias.n130 161.3
R1159 commonsourceibias.n132 commonsourceibias.n125 161.3
R1160 commonsourceibias.n135 commonsourceibias.n134 161.3
R1161 commonsourceibias.n136 commonsourceibias.n124 161.3
R1162 commonsourceibias.n138 commonsourceibias.n137 161.3
R1163 commonsourceibias.n140 commonsourceibias.n123 161.3
R1164 commonsourceibias.n142 commonsourceibias.n141 161.3
R1165 commonsourceibias.n144 commonsourceibias.n143 161.3
R1166 commonsourceibias.n145 commonsourceibias.n121 161.3
R1167 commonsourceibias.n147 commonsourceibias.n146 161.3
R1168 commonsourceibias.n149 commonsourceibias.n148 161.3
R1169 commonsourceibias.n150 commonsourceibias.n119 161.3
R1170 commonsourceibias.n152 commonsourceibias.n151 161.3
R1171 commonsourceibias.n154 commonsourceibias.n153 161.3
R1172 commonsourceibias.n155 commonsourceibias.n117 161.3
R1173 commonsourceibias.n158 commonsourceibias.n157 161.3
R1174 commonsourceibias.n159 commonsourceibias.n11 161.3
R1175 commonsourceibias.n161 commonsourceibias.n160 161.3
R1176 commonsourceibias.n163 commonsourceibias.n9 161.3
R1177 commonsourceibias.n165 commonsourceibias.n164 161.3
R1178 commonsourceibias.n166 commonsourceibias.n8 161.3
R1179 commonsourceibias.n168 commonsourceibias.n167 161.3
R1180 commonsourceibias.n169 commonsourceibias.n7 161.3
R1181 commonsourceibias.n172 commonsourceibias.n171 161.3
R1182 commonsourceibias.n173 commonsourceibias.n6 161.3
R1183 commonsourceibias.n175 commonsourceibias.n174 161.3
R1184 commonsourceibias.n177 commonsourceibias.n4 161.3
R1185 commonsourceibias.n179 commonsourceibias.n178 161.3
R1186 commonsourceibias.n180 commonsourceibias.n3 161.3
R1187 commonsourceibias.n182 commonsourceibias.n181 161.3
R1188 commonsourceibias.n183 commonsourceibias.n2 161.3
R1189 commonsourceibias.n186 commonsourceibias.n185 161.3
R1190 commonsourceibias.n187 commonsourceibias.n1 161.3
R1191 commonsourceibias.n189 commonsourceibias.n188 161.3
R1192 commonsourceibias.n191 commonsourceibias.n0 161.3
R1193 commonsourceibias.n280 commonsourceibias.n194 161.3
R1194 commonsourceibias.n278 commonsourceibias.n277 161.3
R1195 commonsourceibias.n276 commonsourceibias.n195 161.3
R1196 commonsourceibias.n275 commonsourceibias.n274 161.3
R1197 commonsourceibias.n272 commonsourceibias.n196 161.3
R1198 commonsourceibias.n271 commonsourceibias.n270 161.3
R1199 commonsourceibias.n269 commonsourceibias.n197 161.3
R1200 commonsourceibias.n268 commonsourceibias.n267 161.3
R1201 commonsourceibias.n266 commonsourceibias.n198 161.3
R1202 commonsourceibias.n264 commonsourceibias.n263 161.3
R1203 commonsourceibias.n262 commonsourceibias.n200 161.3
R1204 commonsourceibias.n261 commonsourceibias.n260 161.3
R1205 commonsourceibias.n258 commonsourceibias.n201 161.3
R1206 commonsourceibias.n257 commonsourceibias.n256 161.3
R1207 commonsourceibias.n255 commonsourceibias.n202 161.3
R1208 commonsourceibias.n254 commonsourceibias.n253 161.3
R1209 commonsourceibias.n252 commonsourceibias.n203 161.3
R1210 commonsourceibias.n250 commonsourceibias.n249 161.3
R1211 commonsourceibias.n248 commonsourceibias.n205 161.3
R1212 commonsourceibias.n247 commonsourceibias.n246 161.3
R1213 commonsourceibias.n244 commonsourceibias.n206 161.3
R1214 commonsourceibias.n243 commonsourceibias.n242 161.3
R1215 commonsourceibias.n241 commonsourceibias.n240 161.3
R1216 commonsourceibias.n239 commonsourceibias.n208 161.3
R1217 commonsourceibias.n238 commonsourceibias.n237 161.3
R1218 commonsourceibias.n236 commonsourceibias.n235 161.3
R1219 commonsourceibias.n234 commonsourceibias.n210 161.3
R1220 commonsourceibias.n233 commonsourceibias.n232 161.3
R1221 commonsourceibias.n231 commonsourceibias.n230 161.3
R1222 commonsourceibias.n229 commonsourceibias.n212 161.3
R1223 commonsourceibias.n227 commonsourceibias.n226 161.3
R1224 commonsourceibias.n225 commonsourceibias.n213 161.3
R1225 commonsourceibias.n224 commonsourceibias.n223 161.3
R1226 commonsourceibias.n221 commonsourceibias.n214 161.3
R1227 commonsourceibias.n220 commonsourceibias.n219 161.3
R1228 commonsourceibias.n218 commonsourceibias.n215 161.3
R1229 commonsourceibias.n429 commonsourceibias.n343 161.3
R1230 commonsourceibias.n427 commonsourceibias.n426 161.3
R1231 commonsourceibias.n425 commonsourceibias.n344 161.3
R1232 commonsourceibias.n424 commonsourceibias.n423 161.3
R1233 commonsourceibias.n421 commonsourceibias.n345 161.3
R1234 commonsourceibias.n420 commonsourceibias.n419 161.3
R1235 commonsourceibias.n418 commonsourceibias.n346 161.3
R1236 commonsourceibias.n417 commonsourceibias.n416 161.3
R1237 commonsourceibias.n414 commonsourceibias.n347 161.3
R1238 commonsourceibias.n412 commonsourceibias.n411 161.3
R1239 commonsourceibias.n410 commonsourceibias.n348 161.3
R1240 commonsourceibias.n409 commonsourceibias.n408 161.3
R1241 commonsourceibias.n406 commonsourceibias.n349 161.3
R1242 commonsourceibias.n405 commonsourceibias.n404 161.3
R1243 commonsourceibias.n403 commonsourceibias.n350 161.3
R1244 commonsourceibias.n402 commonsourceibias.n401 161.3
R1245 commonsourceibias.n399 commonsourceibias.n351 161.3
R1246 commonsourceibias.n397 commonsourceibias.n396 161.3
R1247 commonsourceibias.n395 commonsourceibias.n352 161.3
R1248 commonsourceibias.n394 commonsourceibias.n393 161.3
R1249 commonsourceibias.n391 commonsourceibias.n353 161.3
R1250 commonsourceibias.n390 commonsourceibias.n389 161.3
R1251 commonsourceibias.n388 commonsourceibias.n387 161.3
R1252 commonsourceibias.n386 commonsourceibias.n355 161.3
R1253 commonsourceibias.n385 commonsourceibias.n384 161.3
R1254 commonsourceibias.n383 commonsourceibias.n382 161.3
R1255 commonsourceibias.n381 commonsourceibias.n357 161.3
R1256 commonsourceibias.n380 commonsourceibias.n379 161.3
R1257 commonsourceibias.n378 commonsourceibias.n377 161.3
R1258 commonsourceibias.n376 commonsourceibias.n359 161.3
R1259 commonsourceibias.n374 commonsourceibias.n373 161.3
R1260 commonsourceibias.n372 commonsourceibias.n360 161.3
R1261 commonsourceibias.n371 commonsourceibias.n370 161.3
R1262 commonsourceibias.n368 commonsourceibias.n361 161.3
R1263 commonsourceibias.n367 commonsourceibias.n366 161.3
R1264 commonsourceibias.n365 commonsourceibias.n362 161.3
R1265 commonsourceibias.n335 commonsourceibias.n334 161.3
R1266 commonsourceibias.n332 commonsourceibias.n294 161.3
R1267 commonsourceibias.n331 commonsourceibias.n330 161.3
R1268 commonsourceibias.n329 commonsourceibias.n328 161.3
R1269 commonsourceibias.n327 commonsourceibias.n296 161.3
R1270 commonsourceibias.n326 commonsourceibias.n325 161.3
R1271 commonsourceibias.n324 commonsourceibias.n323 161.3
R1272 commonsourceibias.n322 commonsourceibias.n298 161.3
R1273 commonsourceibias.n321 commonsourceibias.n320 161.3
R1274 commonsourceibias.n319 commonsourceibias.n318 161.3
R1275 commonsourceibias.n317 commonsourceibias.n300 161.3
R1276 commonsourceibias.n315 commonsourceibias.n314 161.3
R1277 commonsourceibias.n313 commonsourceibias.n301 161.3
R1278 commonsourceibias.n312 commonsourceibias.n311 161.3
R1279 commonsourceibias.n309 commonsourceibias.n302 161.3
R1280 commonsourceibias.n308 commonsourceibias.n307 161.3
R1281 commonsourceibias.n306 commonsourceibias.n303 161.3
R1282 commonsourceibias.n441 commonsourceibias.n293 161.3
R1283 commonsourceibias.n475 commonsourceibias.n284 161.3
R1284 commonsourceibias.n473 commonsourceibias.n472 161.3
R1285 commonsourceibias.n471 commonsourceibias.n285 161.3
R1286 commonsourceibias.n470 commonsourceibias.n469 161.3
R1287 commonsourceibias.n467 commonsourceibias.n286 161.3
R1288 commonsourceibias.n466 commonsourceibias.n465 161.3
R1289 commonsourceibias.n464 commonsourceibias.n287 161.3
R1290 commonsourceibias.n463 commonsourceibias.n462 161.3
R1291 commonsourceibias.n460 commonsourceibias.n288 161.3
R1292 commonsourceibias.n458 commonsourceibias.n457 161.3
R1293 commonsourceibias.n456 commonsourceibias.n289 161.3
R1294 commonsourceibias.n455 commonsourceibias.n454 161.3
R1295 commonsourceibias.n452 commonsourceibias.n290 161.3
R1296 commonsourceibias.n451 commonsourceibias.n450 161.3
R1297 commonsourceibias.n449 commonsourceibias.n291 161.3
R1298 commonsourceibias.n448 commonsourceibias.n447 161.3
R1299 commonsourceibias.n445 commonsourceibias.n292 161.3
R1300 commonsourceibias.n443 commonsourceibias.n442 161.3
R1301 commonsourceibias.n564 commonsourceibias.n478 161.3
R1302 commonsourceibias.n562 commonsourceibias.n561 161.3
R1303 commonsourceibias.n560 commonsourceibias.n479 161.3
R1304 commonsourceibias.n559 commonsourceibias.n558 161.3
R1305 commonsourceibias.n556 commonsourceibias.n480 161.3
R1306 commonsourceibias.n555 commonsourceibias.n554 161.3
R1307 commonsourceibias.n553 commonsourceibias.n481 161.3
R1308 commonsourceibias.n552 commonsourceibias.n551 161.3
R1309 commonsourceibias.n549 commonsourceibias.n482 161.3
R1310 commonsourceibias.n547 commonsourceibias.n546 161.3
R1311 commonsourceibias.n545 commonsourceibias.n483 161.3
R1312 commonsourceibias.n544 commonsourceibias.n543 161.3
R1313 commonsourceibias.n541 commonsourceibias.n484 161.3
R1314 commonsourceibias.n540 commonsourceibias.n539 161.3
R1315 commonsourceibias.n538 commonsourceibias.n485 161.3
R1316 commonsourceibias.n537 commonsourceibias.n536 161.3
R1317 commonsourceibias.n534 commonsourceibias.n486 161.3
R1318 commonsourceibias.n532 commonsourceibias.n531 161.3
R1319 commonsourceibias.n530 commonsourceibias.n487 161.3
R1320 commonsourceibias.n529 commonsourceibias.n528 161.3
R1321 commonsourceibias.n526 commonsourceibias.n488 161.3
R1322 commonsourceibias.n525 commonsourceibias.n524 161.3
R1323 commonsourceibias.n523 commonsourceibias.n522 161.3
R1324 commonsourceibias.n521 commonsourceibias.n490 161.3
R1325 commonsourceibias.n520 commonsourceibias.n519 161.3
R1326 commonsourceibias.n518 commonsourceibias.n517 161.3
R1327 commonsourceibias.n516 commonsourceibias.n492 161.3
R1328 commonsourceibias.n515 commonsourceibias.n514 161.3
R1329 commonsourceibias.n513 commonsourceibias.n512 161.3
R1330 commonsourceibias.n511 commonsourceibias.n494 161.3
R1331 commonsourceibias.n509 commonsourceibias.n508 161.3
R1332 commonsourceibias.n507 commonsourceibias.n495 161.3
R1333 commonsourceibias.n506 commonsourceibias.n505 161.3
R1334 commonsourceibias.n503 commonsourceibias.n496 161.3
R1335 commonsourceibias.n502 commonsourceibias.n501 161.3
R1336 commonsourceibias.n500 commonsourceibias.n497 161.3
R1337 commonsourceibias.n111 commonsourceibias.n109 81.5057
R1338 commonsourceibias.n338 commonsourceibias.n336 81.5057
R1339 commonsourceibias.n111 commonsourceibias.n110 80.9324
R1340 commonsourceibias.n113 commonsourceibias.n112 80.9324
R1341 commonsourceibias.n115 commonsourceibias.n114 80.9324
R1342 commonsourceibias.n108 commonsourceibias.n107 80.9324
R1343 commonsourceibias.n106 commonsourceibias.n105 80.9324
R1344 commonsourceibias.n104 commonsourceibias.n103 80.9324
R1345 commonsourceibias.n102 commonsourceibias.n101 80.9324
R1346 commonsourceibias.n433 commonsourceibias.n432 80.9324
R1347 commonsourceibias.n435 commonsourceibias.n434 80.9324
R1348 commonsourceibias.n437 commonsourceibias.n436 80.9324
R1349 commonsourceibias.n439 commonsourceibias.n438 80.9324
R1350 commonsourceibias.n342 commonsourceibias.n341 80.9324
R1351 commonsourceibias.n340 commonsourceibias.n339 80.9324
R1352 commonsourceibias.n338 commonsourceibias.n337 80.9324
R1353 commonsourceibias.n100 commonsourceibias.n99 80.6037
R1354 commonsourceibias.n193 commonsourceibias.n192 80.6037
R1355 commonsourceibias.n282 commonsourceibias.n281 80.6037
R1356 commonsourceibias.n431 commonsourceibias.n430 80.6037
R1357 commonsourceibias.n477 commonsourceibias.n476 80.6037
R1358 commonsourceibias.n566 commonsourceibias.n565 80.6037
R1359 commonsourceibias.n85 commonsourceibias.n84 56.5617
R1360 commonsourceibias.n71 commonsourceibias.n70 56.5617
R1361 commonsourceibias.n62 commonsourceibias.n61 56.5617
R1362 commonsourceibias.n48 commonsourceibias.n47 56.5617
R1363 commonsourceibias.n178 commonsourceibias.n177 56.5617
R1364 commonsourceibias.n164 commonsourceibias.n163 56.5617
R1365 commonsourceibias.n155 commonsourceibias.n154 56.5617
R1366 commonsourceibias.n141 commonsourceibias.n140 56.5617
R1367 commonsourceibias.n230 commonsourceibias.n229 56.5617
R1368 commonsourceibias.n244 commonsourceibias.n243 56.5617
R1369 commonsourceibias.n253 commonsourceibias.n252 56.5617
R1370 commonsourceibias.n267 commonsourceibias.n266 56.5617
R1371 commonsourceibias.n377 commonsourceibias.n376 56.5617
R1372 commonsourceibias.n391 commonsourceibias.n390 56.5617
R1373 commonsourceibias.n401 commonsourceibias.n399 56.5617
R1374 commonsourceibias.n416 commonsourceibias.n414 56.5617
R1375 commonsourceibias.n462 commonsourceibias.n460 56.5617
R1376 commonsourceibias.n447 commonsourceibias.n445 56.5617
R1377 commonsourceibias.n318 commonsourceibias.n317 56.5617
R1378 commonsourceibias.n332 commonsourceibias.n331 56.5617
R1379 commonsourceibias.n512 commonsourceibias.n511 56.5617
R1380 commonsourceibias.n526 commonsourceibias.n525 56.5617
R1381 commonsourceibias.n536 commonsourceibias.n534 56.5617
R1382 commonsourceibias.n551 commonsourceibias.n549 56.5617
R1383 commonsourceibias.n76 commonsourceibias.n75 56.0773
R1384 commonsourceibias.n57 commonsourceibias.n56 56.0773
R1385 commonsourceibias.n169 commonsourceibias.n168 56.0773
R1386 commonsourceibias.n150 commonsourceibias.n149 56.0773
R1387 commonsourceibias.n239 commonsourceibias.n238 56.0773
R1388 commonsourceibias.n258 commonsourceibias.n257 56.0773
R1389 commonsourceibias.n386 commonsourceibias.n385 56.0773
R1390 commonsourceibias.n406 commonsourceibias.n405 56.0773
R1391 commonsourceibias.n452 commonsourceibias.n451 56.0773
R1392 commonsourceibias.n327 commonsourceibias.n326 56.0773
R1393 commonsourceibias.n521 commonsourceibias.n520 56.0773
R1394 commonsourceibias.n541 commonsourceibias.n540 56.0773
R1395 commonsourceibias.n99 commonsourceibias.n98 55.3321
R1396 commonsourceibias.n192 commonsourceibias.n191 55.3321
R1397 commonsourceibias.n281 commonsourceibias.n280 55.3321
R1398 commonsourceibias.n430 commonsourceibias.n429 55.3321
R1399 commonsourceibias.n476 commonsourceibias.n475 55.3321
R1400 commonsourceibias.n565 commonsourceibias.n564 55.3321
R1401 commonsourceibias.n90 commonsourceibias.n89 55.1086
R1402 commonsourceibias.n41 commonsourceibias.n31 55.1086
R1403 commonsourceibias.n183 commonsourceibias.n182 55.1086
R1404 commonsourceibias.n134 commonsourceibias.n124 55.1086
R1405 commonsourceibias.n223 commonsourceibias.n213 55.1086
R1406 commonsourceibias.n272 commonsourceibias.n271 55.1086
R1407 commonsourceibias.n370 commonsourceibias.n360 55.1086
R1408 commonsourceibias.n421 commonsourceibias.n420 55.1086
R1409 commonsourceibias.n467 commonsourceibias.n466 55.1086
R1410 commonsourceibias.n311 commonsourceibias.n301 55.1086
R1411 commonsourceibias.n505 commonsourceibias.n495 55.1086
R1412 commonsourceibias.n556 commonsourceibias.n555 55.1086
R1413 commonsourceibias.n35 commonsourceibias.n34 47.4592
R1414 commonsourceibias.n128 commonsourceibias.n127 47.4592
R1415 commonsourceibias.n217 commonsourceibias.n216 47.4592
R1416 commonsourceibias.n364 commonsourceibias.n363 47.4592
R1417 commonsourceibias.n305 commonsourceibias.n304 47.4592
R1418 commonsourceibias.n499 commonsourceibias.n498 47.4592
R1419 commonsourceibias.n218 commonsourceibias.n217 44.0436
R1420 commonsourceibias.n365 commonsourceibias.n364 44.0436
R1421 commonsourceibias.n306 commonsourceibias.n305 44.0436
R1422 commonsourceibias.n500 commonsourceibias.n499 44.0436
R1423 commonsourceibias.n36 commonsourceibias.n35 44.0436
R1424 commonsourceibias.n129 commonsourceibias.n128 44.0436
R1425 commonsourceibias.n92 commonsourceibias.n13 42.5146
R1426 commonsourceibias.n39 commonsourceibias.n38 42.5146
R1427 commonsourceibias.n185 commonsourceibias.n1 42.5146
R1428 commonsourceibias.n132 commonsourceibias.n131 42.5146
R1429 commonsourceibias.n221 commonsourceibias.n220 42.5146
R1430 commonsourceibias.n274 commonsourceibias.n195 42.5146
R1431 commonsourceibias.n368 commonsourceibias.n367 42.5146
R1432 commonsourceibias.n423 commonsourceibias.n344 42.5146
R1433 commonsourceibias.n469 commonsourceibias.n285 42.5146
R1434 commonsourceibias.n309 commonsourceibias.n308 42.5146
R1435 commonsourceibias.n503 commonsourceibias.n502 42.5146
R1436 commonsourceibias.n558 commonsourceibias.n479 42.5146
R1437 commonsourceibias.n78 commonsourceibias.n18 41.5458
R1438 commonsourceibias.n53 commonsourceibias.n52 41.5458
R1439 commonsourceibias.n171 commonsourceibias.n6 41.5458
R1440 commonsourceibias.n146 commonsourceibias.n145 41.5458
R1441 commonsourceibias.n235 commonsourceibias.n234 41.5458
R1442 commonsourceibias.n260 commonsourceibias.n200 41.5458
R1443 commonsourceibias.n382 commonsourceibias.n381 41.5458
R1444 commonsourceibias.n408 commonsourceibias.n348 41.5458
R1445 commonsourceibias.n454 commonsourceibias.n289 41.5458
R1446 commonsourceibias.n323 commonsourceibias.n322 41.5458
R1447 commonsourceibias.n517 commonsourceibias.n516 41.5458
R1448 commonsourceibias.n543 commonsourceibias.n483 41.5458
R1449 commonsourceibias.n68 commonsourceibias.n23 40.577
R1450 commonsourceibias.n64 commonsourceibias.n23 40.577
R1451 commonsourceibias.n161 commonsourceibias.n11 40.577
R1452 commonsourceibias.n157 commonsourceibias.n11 40.577
R1453 commonsourceibias.n246 commonsourceibias.n205 40.577
R1454 commonsourceibias.n250 commonsourceibias.n205 40.577
R1455 commonsourceibias.n393 commonsourceibias.n352 40.577
R1456 commonsourceibias.n397 commonsourceibias.n352 40.577
R1457 commonsourceibias.n443 commonsourceibias.n293 40.577
R1458 commonsourceibias.n334 commonsourceibias.n293 40.577
R1459 commonsourceibias.n528 commonsourceibias.n487 40.577
R1460 commonsourceibias.n532 commonsourceibias.n487 40.577
R1461 commonsourceibias.n82 commonsourceibias.n18 39.6083
R1462 commonsourceibias.n52 commonsourceibias.n51 39.6083
R1463 commonsourceibias.n175 commonsourceibias.n6 39.6083
R1464 commonsourceibias.n145 commonsourceibias.n144 39.6083
R1465 commonsourceibias.n234 commonsourceibias.n233 39.6083
R1466 commonsourceibias.n264 commonsourceibias.n200 39.6083
R1467 commonsourceibias.n381 commonsourceibias.n380 39.6083
R1468 commonsourceibias.n412 commonsourceibias.n348 39.6083
R1469 commonsourceibias.n458 commonsourceibias.n289 39.6083
R1470 commonsourceibias.n322 commonsourceibias.n321 39.6083
R1471 commonsourceibias.n516 commonsourceibias.n515 39.6083
R1472 commonsourceibias.n547 commonsourceibias.n483 39.6083
R1473 commonsourceibias.n96 commonsourceibias.n13 38.6395
R1474 commonsourceibias.n38 commonsourceibias.n33 38.6395
R1475 commonsourceibias.n189 commonsourceibias.n1 38.6395
R1476 commonsourceibias.n131 commonsourceibias.n126 38.6395
R1477 commonsourceibias.n220 commonsourceibias.n215 38.6395
R1478 commonsourceibias.n278 commonsourceibias.n195 38.6395
R1479 commonsourceibias.n367 commonsourceibias.n362 38.6395
R1480 commonsourceibias.n427 commonsourceibias.n344 38.6395
R1481 commonsourceibias.n473 commonsourceibias.n285 38.6395
R1482 commonsourceibias.n308 commonsourceibias.n303 38.6395
R1483 commonsourceibias.n502 commonsourceibias.n497 38.6395
R1484 commonsourceibias.n562 commonsourceibias.n479 38.6395
R1485 commonsourceibias.n89 commonsourceibias.n15 26.0455
R1486 commonsourceibias.n45 commonsourceibias.n31 26.0455
R1487 commonsourceibias.n182 commonsourceibias.n3 26.0455
R1488 commonsourceibias.n138 commonsourceibias.n124 26.0455
R1489 commonsourceibias.n227 commonsourceibias.n213 26.0455
R1490 commonsourceibias.n271 commonsourceibias.n197 26.0455
R1491 commonsourceibias.n374 commonsourceibias.n360 26.0455
R1492 commonsourceibias.n420 commonsourceibias.n346 26.0455
R1493 commonsourceibias.n466 commonsourceibias.n287 26.0455
R1494 commonsourceibias.n315 commonsourceibias.n301 26.0455
R1495 commonsourceibias.n509 commonsourceibias.n495 26.0455
R1496 commonsourceibias.n555 commonsourceibias.n481 26.0455
R1497 commonsourceibias.n75 commonsourceibias.n20 25.0767
R1498 commonsourceibias.n58 commonsourceibias.n57 25.0767
R1499 commonsourceibias.n168 commonsourceibias.n8 25.0767
R1500 commonsourceibias.n151 commonsourceibias.n150 25.0767
R1501 commonsourceibias.n240 commonsourceibias.n239 25.0767
R1502 commonsourceibias.n257 commonsourceibias.n202 25.0767
R1503 commonsourceibias.n387 commonsourceibias.n386 25.0767
R1504 commonsourceibias.n405 commonsourceibias.n350 25.0767
R1505 commonsourceibias.n451 commonsourceibias.n291 25.0767
R1506 commonsourceibias.n328 commonsourceibias.n327 25.0767
R1507 commonsourceibias.n522 commonsourceibias.n521 25.0767
R1508 commonsourceibias.n540 commonsourceibias.n485 25.0767
R1509 commonsourceibias.n71 commonsourceibias.n22 24.3464
R1510 commonsourceibias.n61 commonsourceibias.n25 24.3464
R1511 commonsourceibias.n164 commonsourceibias.n10 24.3464
R1512 commonsourceibias.n154 commonsourceibias.n118 24.3464
R1513 commonsourceibias.n243 commonsourceibias.n207 24.3464
R1514 commonsourceibias.n253 commonsourceibias.n204 24.3464
R1515 commonsourceibias.n390 commonsourceibias.n354 24.3464
R1516 commonsourceibias.n401 commonsourceibias.n400 24.3464
R1517 commonsourceibias.n447 commonsourceibias.n446 24.3464
R1518 commonsourceibias.n331 commonsourceibias.n295 24.3464
R1519 commonsourceibias.n525 commonsourceibias.n489 24.3464
R1520 commonsourceibias.n536 commonsourceibias.n535 24.3464
R1521 commonsourceibias.n85 commonsourceibias.n17 23.8546
R1522 commonsourceibias.n47 commonsourceibias.n46 23.8546
R1523 commonsourceibias.n178 commonsourceibias.n5 23.8546
R1524 commonsourceibias.n140 commonsourceibias.n139 23.8546
R1525 commonsourceibias.n229 commonsourceibias.n228 23.8546
R1526 commonsourceibias.n267 commonsourceibias.n199 23.8546
R1527 commonsourceibias.n376 commonsourceibias.n375 23.8546
R1528 commonsourceibias.n416 commonsourceibias.n415 23.8546
R1529 commonsourceibias.n462 commonsourceibias.n461 23.8546
R1530 commonsourceibias.n317 commonsourceibias.n316 23.8546
R1531 commonsourceibias.n511 commonsourceibias.n510 23.8546
R1532 commonsourceibias.n551 commonsourceibias.n550 23.8546
R1533 commonsourceibias.n98 commonsourceibias.n97 17.4607
R1534 commonsourceibias.n191 commonsourceibias.n190 17.4607
R1535 commonsourceibias.n280 commonsourceibias.n279 17.4607
R1536 commonsourceibias.n429 commonsourceibias.n428 17.4607
R1537 commonsourceibias.n475 commonsourceibias.n474 17.4607
R1538 commonsourceibias.n564 commonsourceibias.n563 17.4607
R1539 commonsourceibias.n84 commonsourceibias.n83 16.9689
R1540 commonsourceibias.n48 commonsourceibias.n29 16.9689
R1541 commonsourceibias.n177 commonsourceibias.n176 16.9689
R1542 commonsourceibias.n141 commonsourceibias.n122 16.9689
R1543 commonsourceibias.n230 commonsourceibias.n211 16.9689
R1544 commonsourceibias.n266 commonsourceibias.n265 16.9689
R1545 commonsourceibias.n377 commonsourceibias.n358 16.9689
R1546 commonsourceibias.n414 commonsourceibias.n413 16.9689
R1547 commonsourceibias.n460 commonsourceibias.n459 16.9689
R1548 commonsourceibias.n318 commonsourceibias.n299 16.9689
R1549 commonsourceibias.n512 commonsourceibias.n493 16.9689
R1550 commonsourceibias.n549 commonsourceibias.n548 16.9689
R1551 commonsourceibias.n70 commonsourceibias.n69 16.477
R1552 commonsourceibias.n63 commonsourceibias.n62 16.477
R1553 commonsourceibias.n163 commonsourceibias.n162 16.477
R1554 commonsourceibias.n156 commonsourceibias.n155 16.477
R1555 commonsourceibias.n245 commonsourceibias.n244 16.477
R1556 commonsourceibias.n252 commonsourceibias.n251 16.477
R1557 commonsourceibias.n392 commonsourceibias.n391 16.477
R1558 commonsourceibias.n399 commonsourceibias.n398 16.477
R1559 commonsourceibias.n445 commonsourceibias.n444 16.477
R1560 commonsourceibias.n333 commonsourceibias.n332 16.477
R1561 commonsourceibias.n527 commonsourceibias.n526 16.477
R1562 commonsourceibias.n534 commonsourceibias.n533 16.477
R1563 commonsourceibias.n77 commonsourceibias.n76 15.9852
R1564 commonsourceibias.n56 commonsourceibias.n27 15.9852
R1565 commonsourceibias.n170 commonsourceibias.n169 15.9852
R1566 commonsourceibias.n149 commonsourceibias.n120 15.9852
R1567 commonsourceibias.n238 commonsourceibias.n209 15.9852
R1568 commonsourceibias.n259 commonsourceibias.n258 15.9852
R1569 commonsourceibias.n385 commonsourceibias.n356 15.9852
R1570 commonsourceibias.n407 commonsourceibias.n406 15.9852
R1571 commonsourceibias.n453 commonsourceibias.n452 15.9852
R1572 commonsourceibias.n326 commonsourceibias.n297 15.9852
R1573 commonsourceibias.n520 commonsourceibias.n491 15.9852
R1574 commonsourceibias.n542 commonsourceibias.n541 15.9852
R1575 commonsourceibias.n91 commonsourceibias.n90 15.4934
R1576 commonsourceibias.n41 commonsourceibias.n40 15.4934
R1577 commonsourceibias.n184 commonsourceibias.n183 15.4934
R1578 commonsourceibias.n134 commonsourceibias.n133 15.4934
R1579 commonsourceibias.n223 commonsourceibias.n222 15.4934
R1580 commonsourceibias.n273 commonsourceibias.n272 15.4934
R1581 commonsourceibias.n370 commonsourceibias.n369 15.4934
R1582 commonsourceibias.n422 commonsourceibias.n421 15.4934
R1583 commonsourceibias.n468 commonsourceibias.n467 15.4934
R1584 commonsourceibias.n311 commonsourceibias.n310 15.4934
R1585 commonsourceibias.n505 commonsourceibias.n504 15.4934
R1586 commonsourceibias.n557 commonsourceibias.n556 15.4934
R1587 commonsourceibias.n102 commonsourceibias.n100 13.2663
R1588 commonsourceibias.n433 commonsourceibias.n431 13.2663
R1589 commonsourceibias.n568 commonsourceibias.n283 11.9876
R1590 commonsourceibias.n568 commonsourceibias.n567 10.3347
R1591 commonsourceibias.n159 commonsourceibias.n116 9.50363
R1592 commonsourceibias.n441 commonsourceibias.n440 9.50363
R1593 commonsourceibias.n92 commonsourceibias.n91 9.09948
R1594 commonsourceibias.n40 commonsourceibias.n39 9.09948
R1595 commonsourceibias.n185 commonsourceibias.n184 9.09948
R1596 commonsourceibias.n133 commonsourceibias.n132 9.09948
R1597 commonsourceibias.n222 commonsourceibias.n221 9.09948
R1598 commonsourceibias.n274 commonsourceibias.n273 9.09948
R1599 commonsourceibias.n369 commonsourceibias.n368 9.09948
R1600 commonsourceibias.n423 commonsourceibias.n422 9.09948
R1601 commonsourceibias.n469 commonsourceibias.n468 9.09948
R1602 commonsourceibias.n310 commonsourceibias.n309 9.09948
R1603 commonsourceibias.n504 commonsourceibias.n503 9.09948
R1604 commonsourceibias.n558 commonsourceibias.n557 9.09948
R1605 commonsourceibias.n283 commonsourceibias.n193 8.79261
R1606 commonsourceibias.n567 commonsourceibias.n477 8.79261
R1607 commonsourceibias.n78 commonsourceibias.n77 8.60764
R1608 commonsourceibias.n53 commonsourceibias.n27 8.60764
R1609 commonsourceibias.n171 commonsourceibias.n170 8.60764
R1610 commonsourceibias.n146 commonsourceibias.n120 8.60764
R1611 commonsourceibias.n235 commonsourceibias.n209 8.60764
R1612 commonsourceibias.n260 commonsourceibias.n259 8.60764
R1613 commonsourceibias.n382 commonsourceibias.n356 8.60764
R1614 commonsourceibias.n408 commonsourceibias.n407 8.60764
R1615 commonsourceibias.n454 commonsourceibias.n453 8.60764
R1616 commonsourceibias.n323 commonsourceibias.n297 8.60764
R1617 commonsourceibias.n517 commonsourceibias.n491 8.60764
R1618 commonsourceibias.n543 commonsourceibias.n542 8.60764
R1619 commonsourceibias.n69 commonsourceibias.n68 8.11581
R1620 commonsourceibias.n64 commonsourceibias.n63 8.11581
R1621 commonsourceibias.n162 commonsourceibias.n161 8.11581
R1622 commonsourceibias.n157 commonsourceibias.n156 8.11581
R1623 commonsourceibias.n246 commonsourceibias.n245 8.11581
R1624 commonsourceibias.n251 commonsourceibias.n250 8.11581
R1625 commonsourceibias.n393 commonsourceibias.n392 8.11581
R1626 commonsourceibias.n398 commonsourceibias.n397 8.11581
R1627 commonsourceibias.n444 commonsourceibias.n443 8.11581
R1628 commonsourceibias.n334 commonsourceibias.n333 8.11581
R1629 commonsourceibias.n528 commonsourceibias.n527 8.11581
R1630 commonsourceibias.n533 commonsourceibias.n532 8.11581
R1631 commonsourceibias.n83 commonsourceibias.n82 7.62397
R1632 commonsourceibias.n51 commonsourceibias.n29 7.62397
R1633 commonsourceibias.n176 commonsourceibias.n175 7.62397
R1634 commonsourceibias.n144 commonsourceibias.n122 7.62397
R1635 commonsourceibias.n233 commonsourceibias.n211 7.62397
R1636 commonsourceibias.n265 commonsourceibias.n264 7.62397
R1637 commonsourceibias.n380 commonsourceibias.n358 7.62397
R1638 commonsourceibias.n413 commonsourceibias.n412 7.62397
R1639 commonsourceibias.n459 commonsourceibias.n458 7.62397
R1640 commonsourceibias.n321 commonsourceibias.n299 7.62397
R1641 commonsourceibias.n515 commonsourceibias.n493 7.62397
R1642 commonsourceibias.n548 commonsourceibias.n547 7.62397
R1643 commonsourceibias.n97 commonsourceibias.n96 7.13213
R1644 commonsourceibias.n34 commonsourceibias.n33 7.13213
R1645 commonsourceibias.n190 commonsourceibias.n189 7.13213
R1646 commonsourceibias.n127 commonsourceibias.n126 7.13213
R1647 commonsourceibias.n216 commonsourceibias.n215 7.13213
R1648 commonsourceibias.n279 commonsourceibias.n278 7.13213
R1649 commonsourceibias.n363 commonsourceibias.n362 7.13213
R1650 commonsourceibias.n428 commonsourceibias.n427 7.13213
R1651 commonsourceibias.n474 commonsourceibias.n473 7.13213
R1652 commonsourceibias.n304 commonsourceibias.n303 7.13213
R1653 commonsourceibias.n498 commonsourceibias.n497 7.13213
R1654 commonsourceibias.n563 commonsourceibias.n562 7.13213
R1655 commonsourceibias.n283 commonsourceibias.n282 5.06534
R1656 commonsourceibias.n567 commonsourceibias.n566 5.06534
R1657 commonsourceibias commonsourceibias.n568 4.04308
R1658 commonsourceibias.n109 commonsourceibias.t51 2.82907
R1659 commonsourceibias.n109 commonsourceibias.t1 2.82907
R1660 commonsourceibias.n110 commonsourceibias.t43 2.82907
R1661 commonsourceibias.n110 commonsourceibias.t19 2.82907
R1662 commonsourceibias.n112 commonsourceibias.t9 2.82907
R1663 commonsourceibias.n112 commonsourceibias.t15 2.82907
R1664 commonsourceibias.n114 commonsourceibias.t31 2.82907
R1665 commonsourceibias.n114 commonsourceibias.t5 2.82907
R1666 commonsourceibias.n107 commonsourceibias.t13 2.82907
R1667 commonsourceibias.n107 commonsourceibias.t37 2.82907
R1668 commonsourceibias.n105 commonsourceibias.t45 2.82907
R1669 commonsourceibias.n105 commonsourceibias.t17 2.82907
R1670 commonsourceibias.n103 commonsourceibias.t35 2.82907
R1671 commonsourceibias.n103 commonsourceibias.t27 2.82907
R1672 commonsourceibias.n101 commonsourceibias.t29 2.82907
R1673 commonsourceibias.n101 commonsourceibias.t49 2.82907
R1674 commonsourceibias.n432 commonsourceibias.t39 2.82907
R1675 commonsourceibias.n432 commonsourceibias.t53 2.82907
R1676 commonsourceibias.n434 commonsourceibias.t63 2.82907
R1677 commonsourceibias.n434 commonsourceibias.t21 2.82907
R1678 commonsourceibias.n436 commonsourceibias.t57 2.82907
R1679 commonsourceibias.n436 commonsourceibias.t25 2.82907
R1680 commonsourceibias.n438 commonsourceibias.t11 2.82907
R1681 commonsourceibias.n438 commonsourceibias.t7 2.82907
R1682 commonsourceibias.n341 commonsourceibias.t47 2.82907
R1683 commonsourceibias.n341 commonsourceibias.t55 2.82907
R1684 commonsourceibias.n339 commonsourceibias.t61 2.82907
R1685 commonsourceibias.n339 commonsourceibias.t59 2.82907
R1686 commonsourceibias.n337 commonsourceibias.t3 2.82907
R1687 commonsourceibias.n337 commonsourceibias.t33 2.82907
R1688 commonsourceibias.n336 commonsourceibias.t23 2.82907
R1689 commonsourceibias.n336 commonsourceibias.t41 2.82907
R1690 commonsourceibias.n17 commonsourceibias.n15 0.738255
R1691 commonsourceibias.n46 commonsourceibias.n45 0.738255
R1692 commonsourceibias.n5 commonsourceibias.n3 0.738255
R1693 commonsourceibias.n139 commonsourceibias.n138 0.738255
R1694 commonsourceibias.n228 commonsourceibias.n227 0.738255
R1695 commonsourceibias.n199 commonsourceibias.n197 0.738255
R1696 commonsourceibias.n375 commonsourceibias.n374 0.738255
R1697 commonsourceibias.n415 commonsourceibias.n346 0.738255
R1698 commonsourceibias.n461 commonsourceibias.n287 0.738255
R1699 commonsourceibias.n316 commonsourceibias.n315 0.738255
R1700 commonsourceibias.n510 commonsourceibias.n509 0.738255
R1701 commonsourceibias.n550 commonsourceibias.n481 0.738255
R1702 commonsourceibias.n104 commonsourceibias.n102 0.573776
R1703 commonsourceibias.n106 commonsourceibias.n104 0.573776
R1704 commonsourceibias.n108 commonsourceibias.n106 0.573776
R1705 commonsourceibias.n115 commonsourceibias.n113 0.573776
R1706 commonsourceibias.n113 commonsourceibias.n111 0.573776
R1707 commonsourceibias.n340 commonsourceibias.n338 0.573776
R1708 commonsourceibias.n342 commonsourceibias.n340 0.573776
R1709 commonsourceibias.n439 commonsourceibias.n437 0.573776
R1710 commonsourceibias.n437 commonsourceibias.n435 0.573776
R1711 commonsourceibias.n435 commonsourceibias.n433 0.573776
R1712 commonsourceibias.n116 commonsourceibias.n108 0.287138
R1713 commonsourceibias.n116 commonsourceibias.n115 0.287138
R1714 commonsourceibias.n440 commonsourceibias.n342 0.287138
R1715 commonsourceibias.n440 commonsourceibias.n439 0.287138
R1716 commonsourceibias.n100 commonsourceibias.n12 0.285035
R1717 commonsourceibias.n193 commonsourceibias.n0 0.285035
R1718 commonsourceibias.n282 commonsourceibias.n194 0.285035
R1719 commonsourceibias.n431 commonsourceibias.n343 0.285035
R1720 commonsourceibias.n477 commonsourceibias.n284 0.285035
R1721 commonsourceibias.n566 commonsourceibias.n478 0.285035
R1722 commonsourceibias.n22 commonsourceibias.n20 0.246418
R1723 commonsourceibias.n58 commonsourceibias.n25 0.246418
R1724 commonsourceibias.n10 commonsourceibias.n8 0.246418
R1725 commonsourceibias.n151 commonsourceibias.n118 0.246418
R1726 commonsourceibias.n240 commonsourceibias.n207 0.246418
R1727 commonsourceibias.n204 commonsourceibias.n202 0.246418
R1728 commonsourceibias.n387 commonsourceibias.n354 0.246418
R1729 commonsourceibias.n400 commonsourceibias.n350 0.246418
R1730 commonsourceibias.n446 commonsourceibias.n291 0.246418
R1731 commonsourceibias.n328 commonsourceibias.n295 0.246418
R1732 commonsourceibias.n522 commonsourceibias.n489 0.246418
R1733 commonsourceibias.n535 commonsourceibias.n485 0.246418
R1734 commonsourceibias.n95 commonsourceibias.n12 0.189894
R1735 commonsourceibias.n95 commonsourceibias.n94 0.189894
R1736 commonsourceibias.n94 commonsourceibias.n93 0.189894
R1737 commonsourceibias.n93 commonsourceibias.n14 0.189894
R1738 commonsourceibias.n88 commonsourceibias.n14 0.189894
R1739 commonsourceibias.n88 commonsourceibias.n87 0.189894
R1740 commonsourceibias.n87 commonsourceibias.n86 0.189894
R1741 commonsourceibias.n86 commonsourceibias.n16 0.189894
R1742 commonsourceibias.n81 commonsourceibias.n16 0.189894
R1743 commonsourceibias.n81 commonsourceibias.n80 0.189894
R1744 commonsourceibias.n80 commonsourceibias.n79 0.189894
R1745 commonsourceibias.n79 commonsourceibias.n19 0.189894
R1746 commonsourceibias.n74 commonsourceibias.n19 0.189894
R1747 commonsourceibias.n74 commonsourceibias.n73 0.189894
R1748 commonsourceibias.n73 commonsourceibias.n72 0.189894
R1749 commonsourceibias.n72 commonsourceibias.n21 0.189894
R1750 commonsourceibias.n67 commonsourceibias.n21 0.189894
R1751 commonsourceibias.n67 commonsourceibias.n66 0.189894
R1752 commonsourceibias.n66 commonsourceibias.n65 0.189894
R1753 commonsourceibias.n65 commonsourceibias.n24 0.189894
R1754 commonsourceibias.n60 commonsourceibias.n24 0.189894
R1755 commonsourceibias.n60 commonsourceibias.n59 0.189894
R1756 commonsourceibias.n59 commonsourceibias.n26 0.189894
R1757 commonsourceibias.n55 commonsourceibias.n26 0.189894
R1758 commonsourceibias.n55 commonsourceibias.n54 0.189894
R1759 commonsourceibias.n54 commonsourceibias.n28 0.189894
R1760 commonsourceibias.n50 commonsourceibias.n28 0.189894
R1761 commonsourceibias.n50 commonsourceibias.n49 0.189894
R1762 commonsourceibias.n49 commonsourceibias.n30 0.189894
R1763 commonsourceibias.n44 commonsourceibias.n30 0.189894
R1764 commonsourceibias.n44 commonsourceibias.n43 0.189894
R1765 commonsourceibias.n43 commonsourceibias.n42 0.189894
R1766 commonsourceibias.n42 commonsourceibias.n32 0.189894
R1767 commonsourceibias.n37 commonsourceibias.n32 0.189894
R1768 commonsourceibias.n37 commonsourceibias.n36 0.189894
R1769 commonsourceibias.n158 commonsourceibias.n117 0.189894
R1770 commonsourceibias.n153 commonsourceibias.n117 0.189894
R1771 commonsourceibias.n153 commonsourceibias.n152 0.189894
R1772 commonsourceibias.n152 commonsourceibias.n119 0.189894
R1773 commonsourceibias.n148 commonsourceibias.n119 0.189894
R1774 commonsourceibias.n148 commonsourceibias.n147 0.189894
R1775 commonsourceibias.n147 commonsourceibias.n121 0.189894
R1776 commonsourceibias.n143 commonsourceibias.n121 0.189894
R1777 commonsourceibias.n143 commonsourceibias.n142 0.189894
R1778 commonsourceibias.n142 commonsourceibias.n123 0.189894
R1779 commonsourceibias.n137 commonsourceibias.n123 0.189894
R1780 commonsourceibias.n137 commonsourceibias.n136 0.189894
R1781 commonsourceibias.n136 commonsourceibias.n135 0.189894
R1782 commonsourceibias.n135 commonsourceibias.n125 0.189894
R1783 commonsourceibias.n130 commonsourceibias.n125 0.189894
R1784 commonsourceibias.n130 commonsourceibias.n129 0.189894
R1785 commonsourceibias.n188 commonsourceibias.n0 0.189894
R1786 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1787 commonsourceibias.n187 commonsourceibias.n186 0.189894
R1788 commonsourceibias.n186 commonsourceibias.n2 0.189894
R1789 commonsourceibias.n181 commonsourceibias.n2 0.189894
R1790 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1791 commonsourceibias.n180 commonsourceibias.n179 0.189894
R1792 commonsourceibias.n179 commonsourceibias.n4 0.189894
R1793 commonsourceibias.n174 commonsourceibias.n4 0.189894
R1794 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1795 commonsourceibias.n173 commonsourceibias.n172 0.189894
R1796 commonsourceibias.n172 commonsourceibias.n7 0.189894
R1797 commonsourceibias.n167 commonsourceibias.n7 0.189894
R1798 commonsourceibias.n167 commonsourceibias.n166 0.189894
R1799 commonsourceibias.n166 commonsourceibias.n165 0.189894
R1800 commonsourceibias.n165 commonsourceibias.n9 0.189894
R1801 commonsourceibias.n160 commonsourceibias.n9 0.189894
R1802 commonsourceibias.n277 commonsourceibias.n194 0.189894
R1803 commonsourceibias.n277 commonsourceibias.n276 0.189894
R1804 commonsourceibias.n276 commonsourceibias.n275 0.189894
R1805 commonsourceibias.n275 commonsourceibias.n196 0.189894
R1806 commonsourceibias.n270 commonsourceibias.n196 0.189894
R1807 commonsourceibias.n270 commonsourceibias.n269 0.189894
R1808 commonsourceibias.n269 commonsourceibias.n268 0.189894
R1809 commonsourceibias.n268 commonsourceibias.n198 0.189894
R1810 commonsourceibias.n263 commonsourceibias.n198 0.189894
R1811 commonsourceibias.n263 commonsourceibias.n262 0.189894
R1812 commonsourceibias.n262 commonsourceibias.n261 0.189894
R1813 commonsourceibias.n261 commonsourceibias.n201 0.189894
R1814 commonsourceibias.n256 commonsourceibias.n201 0.189894
R1815 commonsourceibias.n256 commonsourceibias.n255 0.189894
R1816 commonsourceibias.n255 commonsourceibias.n254 0.189894
R1817 commonsourceibias.n254 commonsourceibias.n203 0.189894
R1818 commonsourceibias.n249 commonsourceibias.n203 0.189894
R1819 commonsourceibias.n249 commonsourceibias.n248 0.189894
R1820 commonsourceibias.n248 commonsourceibias.n247 0.189894
R1821 commonsourceibias.n247 commonsourceibias.n206 0.189894
R1822 commonsourceibias.n242 commonsourceibias.n206 0.189894
R1823 commonsourceibias.n242 commonsourceibias.n241 0.189894
R1824 commonsourceibias.n241 commonsourceibias.n208 0.189894
R1825 commonsourceibias.n237 commonsourceibias.n208 0.189894
R1826 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1827 commonsourceibias.n236 commonsourceibias.n210 0.189894
R1828 commonsourceibias.n232 commonsourceibias.n210 0.189894
R1829 commonsourceibias.n232 commonsourceibias.n231 0.189894
R1830 commonsourceibias.n231 commonsourceibias.n212 0.189894
R1831 commonsourceibias.n226 commonsourceibias.n212 0.189894
R1832 commonsourceibias.n226 commonsourceibias.n225 0.189894
R1833 commonsourceibias.n225 commonsourceibias.n224 0.189894
R1834 commonsourceibias.n224 commonsourceibias.n214 0.189894
R1835 commonsourceibias.n219 commonsourceibias.n214 0.189894
R1836 commonsourceibias.n219 commonsourceibias.n218 0.189894
R1837 commonsourceibias.n366 commonsourceibias.n365 0.189894
R1838 commonsourceibias.n366 commonsourceibias.n361 0.189894
R1839 commonsourceibias.n371 commonsourceibias.n361 0.189894
R1840 commonsourceibias.n372 commonsourceibias.n371 0.189894
R1841 commonsourceibias.n373 commonsourceibias.n372 0.189894
R1842 commonsourceibias.n373 commonsourceibias.n359 0.189894
R1843 commonsourceibias.n378 commonsourceibias.n359 0.189894
R1844 commonsourceibias.n379 commonsourceibias.n378 0.189894
R1845 commonsourceibias.n379 commonsourceibias.n357 0.189894
R1846 commonsourceibias.n383 commonsourceibias.n357 0.189894
R1847 commonsourceibias.n384 commonsourceibias.n383 0.189894
R1848 commonsourceibias.n384 commonsourceibias.n355 0.189894
R1849 commonsourceibias.n388 commonsourceibias.n355 0.189894
R1850 commonsourceibias.n389 commonsourceibias.n388 0.189894
R1851 commonsourceibias.n389 commonsourceibias.n353 0.189894
R1852 commonsourceibias.n394 commonsourceibias.n353 0.189894
R1853 commonsourceibias.n395 commonsourceibias.n394 0.189894
R1854 commonsourceibias.n396 commonsourceibias.n395 0.189894
R1855 commonsourceibias.n396 commonsourceibias.n351 0.189894
R1856 commonsourceibias.n402 commonsourceibias.n351 0.189894
R1857 commonsourceibias.n403 commonsourceibias.n402 0.189894
R1858 commonsourceibias.n404 commonsourceibias.n403 0.189894
R1859 commonsourceibias.n404 commonsourceibias.n349 0.189894
R1860 commonsourceibias.n409 commonsourceibias.n349 0.189894
R1861 commonsourceibias.n410 commonsourceibias.n409 0.189894
R1862 commonsourceibias.n411 commonsourceibias.n410 0.189894
R1863 commonsourceibias.n411 commonsourceibias.n347 0.189894
R1864 commonsourceibias.n417 commonsourceibias.n347 0.189894
R1865 commonsourceibias.n418 commonsourceibias.n417 0.189894
R1866 commonsourceibias.n419 commonsourceibias.n418 0.189894
R1867 commonsourceibias.n419 commonsourceibias.n345 0.189894
R1868 commonsourceibias.n424 commonsourceibias.n345 0.189894
R1869 commonsourceibias.n425 commonsourceibias.n424 0.189894
R1870 commonsourceibias.n426 commonsourceibias.n425 0.189894
R1871 commonsourceibias.n426 commonsourceibias.n343 0.189894
R1872 commonsourceibias.n307 commonsourceibias.n306 0.189894
R1873 commonsourceibias.n307 commonsourceibias.n302 0.189894
R1874 commonsourceibias.n312 commonsourceibias.n302 0.189894
R1875 commonsourceibias.n313 commonsourceibias.n312 0.189894
R1876 commonsourceibias.n314 commonsourceibias.n313 0.189894
R1877 commonsourceibias.n314 commonsourceibias.n300 0.189894
R1878 commonsourceibias.n319 commonsourceibias.n300 0.189894
R1879 commonsourceibias.n320 commonsourceibias.n319 0.189894
R1880 commonsourceibias.n320 commonsourceibias.n298 0.189894
R1881 commonsourceibias.n324 commonsourceibias.n298 0.189894
R1882 commonsourceibias.n325 commonsourceibias.n324 0.189894
R1883 commonsourceibias.n325 commonsourceibias.n296 0.189894
R1884 commonsourceibias.n329 commonsourceibias.n296 0.189894
R1885 commonsourceibias.n330 commonsourceibias.n329 0.189894
R1886 commonsourceibias.n330 commonsourceibias.n294 0.189894
R1887 commonsourceibias.n335 commonsourceibias.n294 0.189894
R1888 commonsourceibias.n442 commonsourceibias.n292 0.189894
R1889 commonsourceibias.n448 commonsourceibias.n292 0.189894
R1890 commonsourceibias.n449 commonsourceibias.n448 0.189894
R1891 commonsourceibias.n450 commonsourceibias.n449 0.189894
R1892 commonsourceibias.n450 commonsourceibias.n290 0.189894
R1893 commonsourceibias.n455 commonsourceibias.n290 0.189894
R1894 commonsourceibias.n456 commonsourceibias.n455 0.189894
R1895 commonsourceibias.n457 commonsourceibias.n456 0.189894
R1896 commonsourceibias.n457 commonsourceibias.n288 0.189894
R1897 commonsourceibias.n463 commonsourceibias.n288 0.189894
R1898 commonsourceibias.n464 commonsourceibias.n463 0.189894
R1899 commonsourceibias.n465 commonsourceibias.n464 0.189894
R1900 commonsourceibias.n465 commonsourceibias.n286 0.189894
R1901 commonsourceibias.n470 commonsourceibias.n286 0.189894
R1902 commonsourceibias.n471 commonsourceibias.n470 0.189894
R1903 commonsourceibias.n472 commonsourceibias.n471 0.189894
R1904 commonsourceibias.n472 commonsourceibias.n284 0.189894
R1905 commonsourceibias.n501 commonsourceibias.n500 0.189894
R1906 commonsourceibias.n501 commonsourceibias.n496 0.189894
R1907 commonsourceibias.n506 commonsourceibias.n496 0.189894
R1908 commonsourceibias.n507 commonsourceibias.n506 0.189894
R1909 commonsourceibias.n508 commonsourceibias.n507 0.189894
R1910 commonsourceibias.n508 commonsourceibias.n494 0.189894
R1911 commonsourceibias.n513 commonsourceibias.n494 0.189894
R1912 commonsourceibias.n514 commonsourceibias.n513 0.189894
R1913 commonsourceibias.n514 commonsourceibias.n492 0.189894
R1914 commonsourceibias.n518 commonsourceibias.n492 0.189894
R1915 commonsourceibias.n519 commonsourceibias.n518 0.189894
R1916 commonsourceibias.n519 commonsourceibias.n490 0.189894
R1917 commonsourceibias.n523 commonsourceibias.n490 0.189894
R1918 commonsourceibias.n524 commonsourceibias.n523 0.189894
R1919 commonsourceibias.n524 commonsourceibias.n488 0.189894
R1920 commonsourceibias.n529 commonsourceibias.n488 0.189894
R1921 commonsourceibias.n530 commonsourceibias.n529 0.189894
R1922 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1923 commonsourceibias.n531 commonsourceibias.n486 0.189894
R1924 commonsourceibias.n537 commonsourceibias.n486 0.189894
R1925 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1926 commonsourceibias.n539 commonsourceibias.n538 0.189894
R1927 commonsourceibias.n539 commonsourceibias.n484 0.189894
R1928 commonsourceibias.n544 commonsourceibias.n484 0.189894
R1929 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1930 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1931 commonsourceibias.n546 commonsourceibias.n482 0.189894
R1932 commonsourceibias.n552 commonsourceibias.n482 0.189894
R1933 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1934 commonsourceibias.n554 commonsourceibias.n553 0.189894
R1935 commonsourceibias.n554 commonsourceibias.n480 0.189894
R1936 commonsourceibias.n559 commonsourceibias.n480 0.189894
R1937 commonsourceibias.n560 commonsourceibias.n559 0.189894
R1938 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1939 commonsourceibias.n561 commonsourceibias.n478 0.189894
R1940 commonsourceibias.n159 commonsourceibias.n158 0.170955
R1941 commonsourceibias.n160 commonsourceibias.n159 0.170955
R1942 commonsourceibias.n441 commonsourceibias.n335 0.170955
R1943 commonsourceibias.n442 commonsourceibias.n441 0.170955
R1944 gnd.n6423 gnd.n463 1025.7
R1945 gnd.n4445 gnd.n4444 939.716
R1946 gnd.n6851 gnd.n103 795.207
R1947 gnd.n7015 gnd.n99 795.207
R1948 gnd.n3531 gnd.n1326 795.207
R1949 gnd.n3450 gnd.n1328 795.207
R1950 gnd.n4205 gnd.n1195 795.207
R1951 gnd.n2789 gnd.n1193 795.207
R1952 gnd.n2273 gnd.n884 795.207
R1953 gnd.n2335 gnd.n2274 795.207
R1954 gnd.n7013 gnd.n105 775.989
R1955 gnd.n173 gnd.n101 775.989
R1956 gnd.n3891 gnd.n1325 775.989
R1957 gnd.n4058 gnd.n1329 775.989
R1958 gnd.n4207 gnd.n1190 775.989
R1959 gnd.n2111 gnd.n1192 775.989
R1960 gnd.n4366 gnd.n4365 775.989
R1961 gnd.n4442 gnd.n888 775.989
R1962 gnd.n2835 gnd.n1200 771.183
R1963 gnd.n4076 gnd.n1303 771.183
R1964 gnd.n2849 gnd.n1959 771.183
R1965 gnd.n3564 gnd.n1305 771.183
R1966 gnd.n5889 gnd.n853 766.379
R1967 gnd.n5805 gnd.n855 766.379
R1968 gnd.n5201 gnd.n5100 766.379
R1969 gnd.n5199 gnd.n5102 766.379
R1970 gnd.n5886 gnd.n4447 756.769
R1971 gnd.n5855 gnd.n856 756.769
R1972 gnd.n5446 gnd.n5062 756.769
R1973 gnd.n5432 gnd.n5052 756.769
R1974 gnd.n6065 gnd.n676 689.5
R1975 gnd.n6422 gnd.n464 689.5
R1976 gnd.n6635 gnd.n6633 689.5
R1977 gnd.n2164 gnd.n844 689.5
R1978 gnd.n679 gnd.n676 585
R1979 gnd.n6063 gnd.n676 585
R1980 gnd.n6061 gnd.n6060 585
R1981 gnd.n6062 gnd.n6061 585
R1982 gnd.n6059 gnd.n678 585
R1983 gnd.n678 gnd.n677 585
R1984 gnd.n6058 gnd.n6057 585
R1985 gnd.n6057 gnd.n6056 585
R1986 gnd.n684 gnd.n683 585
R1987 gnd.n6055 gnd.n684 585
R1988 gnd.n6053 gnd.n6052 585
R1989 gnd.n6054 gnd.n6053 585
R1990 gnd.n6051 gnd.n686 585
R1991 gnd.n686 gnd.n685 585
R1992 gnd.n6050 gnd.n6049 585
R1993 gnd.n6049 gnd.n6048 585
R1994 gnd.n692 gnd.n691 585
R1995 gnd.n6047 gnd.n692 585
R1996 gnd.n6045 gnd.n6044 585
R1997 gnd.n6046 gnd.n6045 585
R1998 gnd.n6043 gnd.n694 585
R1999 gnd.n694 gnd.n693 585
R2000 gnd.n6042 gnd.n6041 585
R2001 gnd.n6041 gnd.n6040 585
R2002 gnd.n700 gnd.n699 585
R2003 gnd.n6039 gnd.n700 585
R2004 gnd.n6037 gnd.n6036 585
R2005 gnd.n6038 gnd.n6037 585
R2006 gnd.n6035 gnd.n702 585
R2007 gnd.n702 gnd.n701 585
R2008 gnd.n6034 gnd.n6033 585
R2009 gnd.n6033 gnd.n6032 585
R2010 gnd.n708 gnd.n707 585
R2011 gnd.n6031 gnd.n708 585
R2012 gnd.n6029 gnd.n6028 585
R2013 gnd.n6030 gnd.n6029 585
R2014 gnd.n6027 gnd.n710 585
R2015 gnd.n710 gnd.n709 585
R2016 gnd.n6026 gnd.n6025 585
R2017 gnd.n6025 gnd.n6024 585
R2018 gnd.n716 gnd.n715 585
R2019 gnd.n6023 gnd.n716 585
R2020 gnd.n6021 gnd.n6020 585
R2021 gnd.n6022 gnd.n6021 585
R2022 gnd.n6019 gnd.n718 585
R2023 gnd.n718 gnd.n717 585
R2024 gnd.n6018 gnd.n6017 585
R2025 gnd.n6017 gnd.n6016 585
R2026 gnd.n724 gnd.n723 585
R2027 gnd.n6015 gnd.n724 585
R2028 gnd.n6013 gnd.n6012 585
R2029 gnd.n6014 gnd.n6013 585
R2030 gnd.n6011 gnd.n726 585
R2031 gnd.n726 gnd.n725 585
R2032 gnd.n6010 gnd.n6009 585
R2033 gnd.n6009 gnd.n6008 585
R2034 gnd.n732 gnd.n731 585
R2035 gnd.n6007 gnd.n732 585
R2036 gnd.n6005 gnd.n6004 585
R2037 gnd.n6006 gnd.n6005 585
R2038 gnd.n6003 gnd.n734 585
R2039 gnd.n734 gnd.n733 585
R2040 gnd.n6002 gnd.n6001 585
R2041 gnd.n6001 gnd.n6000 585
R2042 gnd.n740 gnd.n739 585
R2043 gnd.n5999 gnd.n740 585
R2044 gnd.n5997 gnd.n5996 585
R2045 gnd.n5998 gnd.n5997 585
R2046 gnd.n5995 gnd.n742 585
R2047 gnd.n742 gnd.n741 585
R2048 gnd.n5994 gnd.n5993 585
R2049 gnd.n5993 gnd.n5992 585
R2050 gnd.n748 gnd.n747 585
R2051 gnd.n5991 gnd.n748 585
R2052 gnd.n5989 gnd.n5988 585
R2053 gnd.n5990 gnd.n5989 585
R2054 gnd.n5987 gnd.n750 585
R2055 gnd.n750 gnd.n749 585
R2056 gnd.n5986 gnd.n5985 585
R2057 gnd.n5985 gnd.n5984 585
R2058 gnd.n756 gnd.n755 585
R2059 gnd.n5983 gnd.n756 585
R2060 gnd.n5981 gnd.n5980 585
R2061 gnd.n5982 gnd.n5981 585
R2062 gnd.n5979 gnd.n758 585
R2063 gnd.n758 gnd.n757 585
R2064 gnd.n5978 gnd.n5977 585
R2065 gnd.n5977 gnd.n5976 585
R2066 gnd.n764 gnd.n763 585
R2067 gnd.n5975 gnd.n764 585
R2068 gnd.n5973 gnd.n5972 585
R2069 gnd.n5974 gnd.n5973 585
R2070 gnd.n5971 gnd.n766 585
R2071 gnd.n766 gnd.n765 585
R2072 gnd.n5970 gnd.n5969 585
R2073 gnd.n5969 gnd.n5968 585
R2074 gnd.n772 gnd.n771 585
R2075 gnd.n5967 gnd.n772 585
R2076 gnd.n5965 gnd.n5964 585
R2077 gnd.n5966 gnd.n5965 585
R2078 gnd.n5963 gnd.n774 585
R2079 gnd.n774 gnd.n773 585
R2080 gnd.n5962 gnd.n5961 585
R2081 gnd.n5961 gnd.n5960 585
R2082 gnd.n780 gnd.n779 585
R2083 gnd.n5959 gnd.n780 585
R2084 gnd.n5957 gnd.n5956 585
R2085 gnd.n5958 gnd.n5957 585
R2086 gnd.n5955 gnd.n782 585
R2087 gnd.n782 gnd.n781 585
R2088 gnd.n5954 gnd.n5953 585
R2089 gnd.n5953 gnd.n5952 585
R2090 gnd.n788 gnd.n787 585
R2091 gnd.n5951 gnd.n788 585
R2092 gnd.n5949 gnd.n5948 585
R2093 gnd.n5950 gnd.n5949 585
R2094 gnd.n5947 gnd.n790 585
R2095 gnd.n790 gnd.n789 585
R2096 gnd.n5946 gnd.n5945 585
R2097 gnd.n5945 gnd.n5944 585
R2098 gnd.n796 gnd.n795 585
R2099 gnd.n5943 gnd.n796 585
R2100 gnd.n5941 gnd.n5940 585
R2101 gnd.n5942 gnd.n5941 585
R2102 gnd.n5939 gnd.n798 585
R2103 gnd.n798 gnd.n797 585
R2104 gnd.n5938 gnd.n5937 585
R2105 gnd.n5937 gnd.n5936 585
R2106 gnd.n804 gnd.n803 585
R2107 gnd.n5935 gnd.n804 585
R2108 gnd.n5933 gnd.n5932 585
R2109 gnd.n5934 gnd.n5933 585
R2110 gnd.n5931 gnd.n806 585
R2111 gnd.n806 gnd.n805 585
R2112 gnd.n5930 gnd.n5929 585
R2113 gnd.n5929 gnd.n5928 585
R2114 gnd.n812 gnd.n811 585
R2115 gnd.n5927 gnd.n812 585
R2116 gnd.n5925 gnd.n5924 585
R2117 gnd.n5926 gnd.n5925 585
R2118 gnd.n5923 gnd.n814 585
R2119 gnd.n814 gnd.n813 585
R2120 gnd.n5922 gnd.n5921 585
R2121 gnd.n5921 gnd.n5920 585
R2122 gnd.n820 gnd.n819 585
R2123 gnd.n5919 gnd.n820 585
R2124 gnd.n5917 gnd.n5916 585
R2125 gnd.n5918 gnd.n5917 585
R2126 gnd.n5915 gnd.n822 585
R2127 gnd.n822 gnd.n821 585
R2128 gnd.n5914 gnd.n5913 585
R2129 gnd.n5913 gnd.n5912 585
R2130 gnd.n828 gnd.n827 585
R2131 gnd.n5911 gnd.n828 585
R2132 gnd.n5909 gnd.n5908 585
R2133 gnd.n5910 gnd.n5909 585
R2134 gnd.n5907 gnd.n830 585
R2135 gnd.n830 gnd.n829 585
R2136 gnd.n5906 gnd.n5905 585
R2137 gnd.n5905 gnd.n5904 585
R2138 gnd.n836 gnd.n835 585
R2139 gnd.n5903 gnd.n836 585
R2140 gnd.n5901 gnd.n5900 585
R2141 gnd.n5902 gnd.n5901 585
R2142 gnd.n5899 gnd.n838 585
R2143 gnd.n838 gnd.n837 585
R2144 gnd.n5898 gnd.n5897 585
R2145 gnd.n5897 gnd.n5896 585
R2146 gnd.n6066 gnd.n6065 585
R2147 gnd.n6065 gnd.n6064 585
R2148 gnd.n674 gnd.n673 585
R2149 gnd.n673 gnd.n672 585
R2150 gnd.n6071 gnd.n6070 585
R2151 gnd.n6072 gnd.n6071 585
R2152 gnd.n671 gnd.n670 585
R2153 gnd.n6073 gnd.n671 585
R2154 gnd.n6076 gnd.n6075 585
R2155 gnd.n6075 gnd.n6074 585
R2156 gnd.n668 gnd.n667 585
R2157 gnd.n667 gnd.n666 585
R2158 gnd.n6081 gnd.n6080 585
R2159 gnd.n6082 gnd.n6081 585
R2160 gnd.n665 gnd.n664 585
R2161 gnd.n6083 gnd.n665 585
R2162 gnd.n6086 gnd.n6085 585
R2163 gnd.n6085 gnd.n6084 585
R2164 gnd.n662 gnd.n661 585
R2165 gnd.n661 gnd.n660 585
R2166 gnd.n6091 gnd.n6090 585
R2167 gnd.n6092 gnd.n6091 585
R2168 gnd.n659 gnd.n658 585
R2169 gnd.n6093 gnd.n659 585
R2170 gnd.n6096 gnd.n6095 585
R2171 gnd.n6095 gnd.n6094 585
R2172 gnd.n656 gnd.n655 585
R2173 gnd.n655 gnd.n654 585
R2174 gnd.n6101 gnd.n6100 585
R2175 gnd.n6102 gnd.n6101 585
R2176 gnd.n653 gnd.n652 585
R2177 gnd.n6103 gnd.n653 585
R2178 gnd.n6106 gnd.n6105 585
R2179 gnd.n6105 gnd.n6104 585
R2180 gnd.n650 gnd.n649 585
R2181 gnd.n649 gnd.n648 585
R2182 gnd.n6111 gnd.n6110 585
R2183 gnd.n6112 gnd.n6111 585
R2184 gnd.n647 gnd.n646 585
R2185 gnd.n6113 gnd.n647 585
R2186 gnd.n6116 gnd.n6115 585
R2187 gnd.n6115 gnd.n6114 585
R2188 gnd.n644 gnd.n643 585
R2189 gnd.n643 gnd.n642 585
R2190 gnd.n6121 gnd.n6120 585
R2191 gnd.n6122 gnd.n6121 585
R2192 gnd.n641 gnd.n640 585
R2193 gnd.n6123 gnd.n641 585
R2194 gnd.n6126 gnd.n6125 585
R2195 gnd.n6125 gnd.n6124 585
R2196 gnd.n638 gnd.n637 585
R2197 gnd.n637 gnd.n636 585
R2198 gnd.n6131 gnd.n6130 585
R2199 gnd.n6132 gnd.n6131 585
R2200 gnd.n635 gnd.n634 585
R2201 gnd.n6133 gnd.n635 585
R2202 gnd.n6136 gnd.n6135 585
R2203 gnd.n6135 gnd.n6134 585
R2204 gnd.n632 gnd.n631 585
R2205 gnd.n631 gnd.n630 585
R2206 gnd.n6141 gnd.n6140 585
R2207 gnd.n6142 gnd.n6141 585
R2208 gnd.n629 gnd.n628 585
R2209 gnd.n6143 gnd.n629 585
R2210 gnd.n6146 gnd.n6145 585
R2211 gnd.n6145 gnd.n6144 585
R2212 gnd.n626 gnd.n625 585
R2213 gnd.n625 gnd.n624 585
R2214 gnd.n6151 gnd.n6150 585
R2215 gnd.n6152 gnd.n6151 585
R2216 gnd.n623 gnd.n622 585
R2217 gnd.n6153 gnd.n623 585
R2218 gnd.n6156 gnd.n6155 585
R2219 gnd.n6155 gnd.n6154 585
R2220 gnd.n620 gnd.n619 585
R2221 gnd.n619 gnd.n618 585
R2222 gnd.n6161 gnd.n6160 585
R2223 gnd.n6162 gnd.n6161 585
R2224 gnd.n617 gnd.n616 585
R2225 gnd.n6163 gnd.n617 585
R2226 gnd.n6166 gnd.n6165 585
R2227 gnd.n6165 gnd.n6164 585
R2228 gnd.n614 gnd.n613 585
R2229 gnd.n613 gnd.n612 585
R2230 gnd.n6171 gnd.n6170 585
R2231 gnd.n6172 gnd.n6171 585
R2232 gnd.n611 gnd.n610 585
R2233 gnd.n6173 gnd.n611 585
R2234 gnd.n6176 gnd.n6175 585
R2235 gnd.n6175 gnd.n6174 585
R2236 gnd.n608 gnd.n607 585
R2237 gnd.n607 gnd.n606 585
R2238 gnd.n6181 gnd.n6180 585
R2239 gnd.n6182 gnd.n6181 585
R2240 gnd.n605 gnd.n604 585
R2241 gnd.n6183 gnd.n605 585
R2242 gnd.n6186 gnd.n6185 585
R2243 gnd.n6185 gnd.n6184 585
R2244 gnd.n602 gnd.n601 585
R2245 gnd.n601 gnd.n600 585
R2246 gnd.n6191 gnd.n6190 585
R2247 gnd.n6192 gnd.n6191 585
R2248 gnd.n599 gnd.n598 585
R2249 gnd.n6193 gnd.n599 585
R2250 gnd.n6196 gnd.n6195 585
R2251 gnd.n6195 gnd.n6194 585
R2252 gnd.n596 gnd.n595 585
R2253 gnd.n595 gnd.n594 585
R2254 gnd.n6201 gnd.n6200 585
R2255 gnd.n6202 gnd.n6201 585
R2256 gnd.n593 gnd.n592 585
R2257 gnd.n6203 gnd.n593 585
R2258 gnd.n6206 gnd.n6205 585
R2259 gnd.n6205 gnd.n6204 585
R2260 gnd.n590 gnd.n589 585
R2261 gnd.n589 gnd.n588 585
R2262 gnd.n6211 gnd.n6210 585
R2263 gnd.n6212 gnd.n6211 585
R2264 gnd.n587 gnd.n586 585
R2265 gnd.n6213 gnd.n587 585
R2266 gnd.n6216 gnd.n6215 585
R2267 gnd.n6215 gnd.n6214 585
R2268 gnd.n584 gnd.n583 585
R2269 gnd.n583 gnd.n582 585
R2270 gnd.n6221 gnd.n6220 585
R2271 gnd.n6222 gnd.n6221 585
R2272 gnd.n581 gnd.n580 585
R2273 gnd.n6223 gnd.n581 585
R2274 gnd.n6226 gnd.n6225 585
R2275 gnd.n6225 gnd.n6224 585
R2276 gnd.n578 gnd.n577 585
R2277 gnd.n577 gnd.n576 585
R2278 gnd.n6231 gnd.n6230 585
R2279 gnd.n6232 gnd.n6231 585
R2280 gnd.n575 gnd.n574 585
R2281 gnd.n6233 gnd.n575 585
R2282 gnd.n6236 gnd.n6235 585
R2283 gnd.n6235 gnd.n6234 585
R2284 gnd.n572 gnd.n571 585
R2285 gnd.n571 gnd.n570 585
R2286 gnd.n6241 gnd.n6240 585
R2287 gnd.n6242 gnd.n6241 585
R2288 gnd.n569 gnd.n568 585
R2289 gnd.n6243 gnd.n569 585
R2290 gnd.n6246 gnd.n6245 585
R2291 gnd.n6245 gnd.n6244 585
R2292 gnd.n566 gnd.n565 585
R2293 gnd.n565 gnd.n564 585
R2294 gnd.n6251 gnd.n6250 585
R2295 gnd.n6252 gnd.n6251 585
R2296 gnd.n563 gnd.n562 585
R2297 gnd.n6253 gnd.n563 585
R2298 gnd.n6256 gnd.n6255 585
R2299 gnd.n6255 gnd.n6254 585
R2300 gnd.n560 gnd.n559 585
R2301 gnd.n559 gnd.n558 585
R2302 gnd.n6261 gnd.n6260 585
R2303 gnd.n6262 gnd.n6261 585
R2304 gnd.n557 gnd.n556 585
R2305 gnd.n6263 gnd.n557 585
R2306 gnd.n6266 gnd.n6265 585
R2307 gnd.n6265 gnd.n6264 585
R2308 gnd.n554 gnd.n553 585
R2309 gnd.n553 gnd.n552 585
R2310 gnd.n6271 gnd.n6270 585
R2311 gnd.n6272 gnd.n6271 585
R2312 gnd.n551 gnd.n550 585
R2313 gnd.n6273 gnd.n551 585
R2314 gnd.n6276 gnd.n6275 585
R2315 gnd.n6275 gnd.n6274 585
R2316 gnd.n548 gnd.n547 585
R2317 gnd.n547 gnd.n546 585
R2318 gnd.n6281 gnd.n6280 585
R2319 gnd.n6282 gnd.n6281 585
R2320 gnd.n545 gnd.n544 585
R2321 gnd.n6283 gnd.n545 585
R2322 gnd.n6286 gnd.n6285 585
R2323 gnd.n6285 gnd.n6284 585
R2324 gnd.n542 gnd.n541 585
R2325 gnd.n541 gnd.n540 585
R2326 gnd.n6291 gnd.n6290 585
R2327 gnd.n6292 gnd.n6291 585
R2328 gnd.n539 gnd.n538 585
R2329 gnd.n6293 gnd.n539 585
R2330 gnd.n6296 gnd.n6295 585
R2331 gnd.n6295 gnd.n6294 585
R2332 gnd.n536 gnd.n535 585
R2333 gnd.n535 gnd.n534 585
R2334 gnd.n6301 gnd.n6300 585
R2335 gnd.n6302 gnd.n6301 585
R2336 gnd.n533 gnd.n532 585
R2337 gnd.n6303 gnd.n533 585
R2338 gnd.n6306 gnd.n6305 585
R2339 gnd.n6305 gnd.n6304 585
R2340 gnd.n530 gnd.n529 585
R2341 gnd.n529 gnd.n528 585
R2342 gnd.n6311 gnd.n6310 585
R2343 gnd.n6312 gnd.n6311 585
R2344 gnd.n527 gnd.n526 585
R2345 gnd.n6313 gnd.n527 585
R2346 gnd.n6316 gnd.n6315 585
R2347 gnd.n6315 gnd.n6314 585
R2348 gnd.n524 gnd.n523 585
R2349 gnd.n523 gnd.n522 585
R2350 gnd.n6321 gnd.n6320 585
R2351 gnd.n6322 gnd.n6321 585
R2352 gnd.n521 gnd.n520 585
R2353 gnd.n6323 gnd.n521 585
R2354 gnd.n6326 gnd.n6325 585
R2355 gnd.n6325 gnd.n6324 585
R2356 gnd.n518 gnd.n517 585
R2357 gnd.n517 gnd.n516 585
R2358 gnd.n6331 gnd.n6330 585
R2359 gnd.n6332 gnd.n6331 585
R2360 gnd.n515 gnd.n514 585
R2361 gnd.n6333 gnd.n515 585
R2362 gnd.n6336 gnd.n6335 585
R2363 gnd.n6335 gnd.n6334 585
R2364 gnd.n512 gnd.n511 585
R2365 gnd.n511 gnd.n510 585
R2366 gnd.n6341 gnd.n6340 585
R2367 gnd.n6342 gnd.n6341 585
R2368 gnd.n509 gnd.n508 585
R2369 gnd.n6343 gnd.n509 585
R2370 gnd.n6346 gnd.n6345 585
R2371 gnd.n6345 gnd.n6344 585
R2372 gnd.n506 gnd.n505 585
R2373 gnd.n505 gnd.n504 585
R2374 gnd.n6351 gnd.n6350 585
R2375 gnd.n6352 gnd.n6351 585
R2376 gnd.n503 gnd.n502 585
R2377 gnd.n6353 gnd.n503 585
R2378 gnd.n6356 gnd.n6355 585
R2379 gnd.n6355 gnd.n6354 585
R2380 gnd.n500 gnd.n499 585
R2381 gnd.n499 gnd.n498 585
R2382 gnd.n6361 gnd.n6360 585
R2383 gnd.n6362 gnd.n6361 585
R2384 gnd.n497 gnd.n496 585
R2385 gnd.n6363 gnd.n497 585
R2386 gnd.n6366 gnd.n6365 585
R2387 gnd.n6365 gnd.n6364 585
R2388 gnd.n494 gnd.n493 585
R2389 gnd.n493 gnd.n492 585
R2390 gnd.n6371 gnd.n6370 585
R2391 gnd.n6372 gnd.n6371 585
R2392 gnd.n491 gnd.n490 585
R2393 gnd.n6373 gnd.n491 585
R2394 gnd.n6376 gnd.n6375 585
R2395 gnd.n6375 gnd.n6374 585
R2396 gnd.n488 gnd.n487 585
R2397 gnd.n487 gnd.n486 585
R2398 gnd.n6381 gnd.n6380 585
R2399 gnd.n6382 gnd.n6381 585
R2400 gnd.n485 gnd.n484 585
R2401 gnd.n6383 gnd.n485 585
R2402 gnd.n6386 gnd.n6385 585
R2403 gnd.n6385 gnd.n6384 585
R2404 gnd.n482 gnd.n481 585
R2405 gnd.n481 gnd.n480 585
R2406 gnd.n6391 gnd.n6390 585
R2407 gnd.n6392 gnd.n6391 585
R2408 gnd.n479 gnd.n478 585
R2409 gnd.n6393 gnd.n479 585
R2410 gnd.n6396 gnd.n6395 585
R2411 gnd.n6395 gnd.n6394 585
R2412 gnd.n476 gnd.n475 585
R2413 gnd.n475 gnd.n474 585
R2414 gnd.n6401 gnd.n6400 585
R2415 gnd.n6402 gnd.n6401 585
R2416 gnd.n473 gnd.n472 585
R2417 gnd.n6403 gnd.n473 585
R2418 gnd.n6406 gnd.n6405 585
R2419 gnd.n6405 gnd.n6404 585
R2420 gnd.n470 gnd.n469 585
R2421 gnd.n469 gnd.n468 585
R2422 gnd.n6412 gnd.n6411 585
R2423 gnd.n6413 gnd.n6412 585
R2424 gnd.n467 gnd.n466 585
R2425 gnd.n6414 gnd.n467 585
R2426 gnd.n6417 gnd.n6416 585
R2427 gnd.n6416 gnd.n6415 585
R2428 gnd.n6418 gnd.n464 585
R2429 gnd.n464 gnd.n463 585
R2430 gnd.n339 gnd.n338 585
R2431 gnd.n6625 gnd.n338 585
R2432 gnd.n6628 gnd.n6627 585
R2433 gnd.n6627 gnd.n6626 585
R2434 gnd.n342 gnd.n341 585
R2435 gnd.n6624 gnd.n342 585
R2436 gnd.n6622 gnd.n6621 585
R2437 gnd.n6623 gnd.n6622 585
R2438 gnd.n345 gnd.n344 585
R2439 gnd.n344 gnd.n343 585
R2440 gnd.n6617 gnd.n6616 585
R2441 gnd.n6616 gnd.n6615 585
R2442 gnd.n348 gnd.n347 585
R2443 gnd.n6614 gnd.n348 585
R2444 gnd.n6612 gnd.n6611 585
R2445 gnd.n6613 gnd.n6612 585
R2446 gnd.n351 gnd.n350 585
R2447 gnd.n350 gnd.n349 585
R2448 gnd.n6607 gnd.n6606 585
R2449 gnd.n6606 gnd.n6605 585
R2450 gnd.n354 gnd.n353 585
R2451 gnd.n6604 gnd.n354 585
R2452 gnd.n6602 gnd.n6601 585
R2453 gnd.n6603 gnd.n6602 585
R2454 gnd.n357 gnd.n356 585
R2455 gnd.n356 gnd.n355 585
R2456 gnd.n6597 gnd.n6596 585
R2457 gnd.n6596 gnd.n6595 585
R2458 gnd.n360 gnd.n359 585
R2459 gnd.n6594 gnd.n360 585
R2460 gnd.n6592 gnd.n6591 585
R2461 gnd.n6593 gnd.n6592 585
R2462 gnd.n363 gnd.n362 585
R2463 gnd.n362 gnd.n361 585
R2464 gnd.n6587 gnd.n6586 585
R2465 gnd.n6586 gnd.n6585 585
R2466 gnd.n366 gnd.n365 585
R2467 gnd.n6584 gnd.n366 585
R2468 gnd.n6582 gnd.n6581 585
R2469 gnd.n6583 gnd.n6582 585
R2470 gnd.n369 gnd.n368 585
R2471 gnd.n368 gnd.n367 585
R2472 gnd.n6577 gnd.n6576 585
R2473 gnd.n6576 gnd.n6575 585
R2474 gnd.n372 gnd.n371 585
R2475 gnd.n6574 gnd.n372 585
R2476 gnd.n6572 gnd.n6571 585
R2477 gnd.n6573 gnd.n6572 585
R2478 gnd.n375 gnd.n374 585
R2479 gnd.n374 gnd.n373 585
R2480 gnd.n6567 gnd.n6566 585
R2481 gnd.n6566 gnd.n6565 585
R2482 gnd.n378 gnd.n377 585
R2483 gnd.n6564 gnd.n378 585
R2484 gnd.n6562 gnd.n6561 585
R2485 gnd.n6563 gnd.n6562 585
R2486 gnd.n381 gnd.n380 585
R2487 gnd.n380 gnd.n379 585
R2488 gnd.n6557 gnd.n6556 585
R2489 gnd.n6556 gnd.n6555 585
R2490 gnd.n384 gnd.n383 585
R2491 gnd.n6554 gnd.n384 585
R2492 gnd.n6552 gnd.n6551 585
R2493 gnd.n6553 gnd.n6552 585
R2494 gnd.n387 gnd.n386 585
R2495 gnd.n386 gnd.n385 585
R2496 gnd.n6547 gnd.n6546 585
R2497 gnd.n6546 gnd.n6545 585
R2498 gnd.n390 gnd.n389 585
R2499 gnd.n6544 gnd.n390 585
R2500 gnd.n6542 gnd.n6541 585
R2501 gnd.n6543 gnd.n6542 585
R2502 gnd.n393 gnd.n392 585
R2503 gnd.n392 gnd.n391 585
R2504 gnd.n6537 gnd.n6536 585
R2505 gnd.n6536 gnd.n6535 585
R2506 gnd.n396 gnd.n395 585
R2507 gnd.n6534 gnd.n396 585
R2508 gnd.n6532 gnd.n6531 585
R2509 gnd.n6533 gnd.n6532 585
R2510 gnd.n399 gnd.n398 585
R2511 gnd.n398 gnd.n397 585
R2512 gnd.n6527 gnd.n6526 585
R2513 gnd.n6526 gnd.n6525 585
R2514 gnd.n402 gnd.n401 585
R2515 gnd.n6524 gnd.n402 585
R2516 gnd.n6522 gnd.n6521 585
R2517 gnd.n6523 gnd.n6522 585
R2518 gnd.n405 gnd.n404 585
R2519 gnd.n404 gnd.n403 585
R2520 gnd.n6517 gnd.n6516 585
R2521 gnd.n6516 gnd.n6515 585
R2522 gnd.n408 gnd.n407 585
R2523 gnd.n6514 gnd.n408 585
R2524 gnd.n6512 gnd.n6511 585
R2525 gnd.n6513 gnd.n6512 585
R2526 gnd.n411 gnd.n410 585
R2527 gnd.n410 gnd.n409 585
R2528 gnd.n6507 gnd.n6506 585
R2529 gnd.n6506 gnd.n6505 585
R2530 gnd.n414 gnd.n413 585
R2531 gnd.n6504 gnd.n414 585
R2532 gnd.n6502 gnd.n6501 585
R2533 gnd.n6503 gnd.n6502 585
R2534 gnd.n417 gnd.n416 585
R2535 gnd.n416 gnd.n415 585
R2536 gnd.n6497 gnd.n6496 585
R2537 gnd.n6496 gnd.n6495 585
R2538 gnd.n420 gnd.n419 585
R2539 gnd.n6494 gnd.n420 585
R2540 gnd.n6492 gnd.n6491 585
R2541 gnd.n6493 gnd.n6492 585
R2542 gnd.n423 gnd.n422 585
R2543 gnd.n422 gnd.n421 585
R2544 gnd.n6487 gnd.n6486 585
R2545 gnd.n6486 gnd.n6485 585
R2546 gnd.n426 gnd.n425 585
R2547 gnd.n6484 gnd.n426 585
R2548 gnd.n6482 gnd.n6481 585
R2549 gnd.n6483 gnd.n6482 585
R2550 gnd.n429 gnd.n428 585
R2551 gnd.n428 gnd.n427 585
R2552 gnd.n6477 gnd.n6476 585
R2553 gnd.n6476 gnd.n6475 585
R2554 gnd.n432 gnd.n431 585
R2555 gnd.n6474 gnd.n432 585
R2556 gnd.n6472 gnd.n6471 585
R2557 gnd.n6473 gnd.n6472 585
R2558 gnd.n435 gnd.n434 585
R2559 gnd.n434 gnd.n433 585
R2560 gnd.n6467 gnd.n6466 585
R2561 gnd.n6466 gnd.n6465 585
R2562 gnd.n438 gnd.n437 585
R2563 gnd.n6464 gnd.n438 585
R2564 gnd.n6462 gnd.n6461 585
R2565 gnd.n6463 gnd.n6462 585
R2566 gnd.n441 gnd.n440 585
R2567 gnd.n440 gnd.n439 585
R2568 gnd.n6457 gnd.n6456 585
R2569 gnd.n6456 gnd.n6455 585
R2570 gnd.n444 gnd.n443 585
R2571 gnd.n6454 gnd.n444 585
R2572 gnd.n6452 gnd.n6451 585
R2573 gnd.n6453 gnd.n6452 585
R2574 gnd.n447 gnd.n446 585
R2575 gnd.n446 gnd.n445 585
R2576 gnd.n6447 gnd.n6446 585
R2577 gnd.n6446 gnd.n6445 585
R2578 gnd.n450 gnd.n449 585
R2579 gnd.n6444 gnd.n450 585
R2580 gnd.n6442 gnd.n6441 585
R2581 gnd.n6443 gnd.n6442 585
R2582 gnd.n453 gnd.n452 585
R2583 gnd.n452 gnd.n451 585
R2584 gnd.n6437 gnd.n6436 585
R2585 gnd.n6436 gnd.n6435 585
R2586 gnd.n456 gnd.n455 585
R2587 gnd.n6434 gnd.n456 585
R2588 gnd.n6432 gnd.n6431 585
R2589 gnd.n6433 gnd.n6432 585
R2590 gnd.n459 gnd.n458 585
R2591 gnd.n458 gnd.n457 585
R2592 gnd.n6427 gnd.n6426 585
R2593 gnd.n6426 gnd.n6425 585
R2594 gnd.n462 gnd.n461 585
R2595 gnd.n6424 gnd.n462 585
R2596 gnd.n6422 gnd.n6421 585
R2597 gnd.n6423 gnd.n6422 585
R2598 gnd.n4205 gnd.n4204 585
R2599 gnd.n4206 gnd.n4205 585
R2600 gnd.n1180 gnd.n1179 585
R2601 gnd.n2580 gnd.n1180 585
R2602 gnd.n4214 gnd.n4213 585
R2603 gnd.n4213 gnd.n4212 585
R2604 gnd.n4215 gnd.n1174 585
R2605 gnd.n2536 gnd.n1174 585
R2606 gnd.n4217 gnd.n4216 585
R2607 gnd.n4218 gnd.n4217 585
R2608 gnd.n1159 gnd.n1158 585
R2609 gnd.n2527 gnd.n1159 585
R2610 gnd.n4226 gnd.n4225 585
R2611 gnd.n4225 gnd.n4224 585
R2612 gnd.n4227 gnd.n1153 585
R2613 gnd.n2519 gnd.n1153 585
R2614 gnd.n4229 gnd.n4228 585
R2615 gnd.n4230 gnd.n4229 585
R2616 gnd.n1137 gnd.n1136 585
R2617 gnd.n2459 gnd.n1137 585
R2618 gnd.n4238 gnd.n4237 585
R2619 gnd.n4237 gnd.n4236 585
R2620 gnd.n4239 gnd.n1131 585
R2621 gnd.n2447 gnd.n1131 585
R2622 gnd.n4241 gnd.n4240 585
R2623 gnd.n4242 gnd.n4241 585
R2624 gnd.n1117 gnd.n1116 585
R2625 gnd.n2442 gnd.n1117 585
R2626 gnd.n4250 gnd.n4249 585
R2627 gnd.n4249 gnd.n4248 585
R2628 gnd.n4251 gnd.n1111 585
R2629 gnd.n2473 gnd.n1111 585
R2630 gnd.n4253 gnd.n4252 585
R2631 gnd.n4254 gnd.n4253 585
R2632 gnd.n1095 gnd.n1094 585
R2633 gnd.n2434 gnd.n1095 585
R2634 gnd.n4262 gnd.n4261 585
R2635 gnd.n4261 gnd.n4260 585
R2636 gnd.n4263 gnd.n1089 585
R2637 gnd.n2426 gnd.n1089 585
R2638 gnd.n4265 gnd.n4264 585
R2639 gnd.n4266 gnd.n4265 585
R2640 gnd.n1076 gnd.n1075 585
R2641 gnd.n2417 gnd.n1076 585
R2642 gnd.n4274 gnd.n4273 585
R2643 gnd.n4273 gnd.n4272 585
R2644 gnd.n4275 gnd.n1070 585
R2645 gnd.n1070 gnd.n1069 585
R2646 gnd.n4277 gnd.n4276 585
R2647 gnd.n4278 gnd.n4277 585
R2648 gnd.n1058 gnd.n1057 585
R2649 gnd.n2257 gnd.n1058 585
R2650 gnd.n4287 gnd.n4286 585
R2651 gnd.n4286 gnd.n4285 585
R2652 gnd.n4288 gnd.n1052 585
R2653 gnd.n1059 gnd.n1052 585
R2654 gnd.n4290 gnd.n4289 585
R2655 gnd.n4291 gnd.n4290 585
R2656 gnd.n1041 gnd.n1040 585
R2657 gnd.n1044 gnd.n1041 585
R2658 gnd.n4299 gnd.n4298 585
R2659 gnd.n4298 gnd.n4297 585
R2660 gnd.n4300 gnd.n1035 585
R2661 gnd.n1035 gnd.n1034 585
R2662 gnd.n4302 gnd.n4301 585
R2663 gnd.n4303 gnd.n4302 585
R2664 gnd.n1020 gnd.n1019 585
R2665 gnd.n1031 gnd.n1020 585
R2666 gnd.n4311 gnd.n4310 585
R2667 gnd.n4310 gnd.n4309 585
R2668 gnd.n4312 gnd.n1014 585
R2669 gnd.n1021 gnd.n1014 585
R2670 gnd.n4314 gnd.n4313 585
R2671 gnd.n4315 gnd.n4314 585
R2672 gnd.n1001 gnd.n1000 585
R2673 gnd.n1004 gnd.n1001 585
R2674 gnd.n4323 gnd.n4322 585
R2675 gnd.n4322 gnd.n4321 585
R2676 gnd.n4324 gnd.n995 585
R2677 gnd.n995 gnd.n994 585
R2678 gnd.n4326 gnd.n4325 585
R2679 gnd.n4327 gnd.n4326 585
R2680 gnd.n980 gnd.n979 585
R2681 gnd.n991 gnd.n980 585
R2682 gnd.n4335 gnd.n4334 585
R2683 gnd.n4334 gnd.n4333 585
R2684 gnd.n4336 gnd.n974 585
R2685 gnd.n981 gnd.n974 585
R2686 gnd.n4338 gnd.n4337 585
R2687 gnd.n4339 gnd.n4338 585
R2688 gnd.n961 gnd.n960 585
R2689 gnd.n964 gnd.n961 585
R2690 gnd.n4347 gnd.n4346 585
R2691 gnd.n4346 gnd.n4345 585
R2692 gnd.n4348 gnd.n955 585
R2693 gnd.n955 gnd.n953 585
R2694 gnd.n4350 gnd.n4349 585
R2695 gnd.n4351 gnd.n4350 585
R2696 gnd.n956 gnd.n954 585
R2697 gnd.n954 gnd.n941 585
R2698 gnd.n2340 gnd.n942 585
R2699 gnd.n4357 gnd.n942 585
R2700 gnd.n2277 gnd.n2275 585
R2701 gnd.n2275 gnd.n939 585
R2702 gnd.n2345 gnd.n2344 585
R2703 gnd.n2352 gnd.n2345 585
R2704 gnd.n2276 gnd.n2274 585
R2705 gnd.n2274 gnd.n885 585
R2706 gnd.n2336 gnd.n2335 585
R2707 gnd.n2334 gnd.n2333 585
R2708 gnd.n2332 gnd.n2331 585
R2709 gnd.n2330 gnd.n2329 585
R2710 gnd.n2328 gnd.n2327 585
R2711 gnd.n2326 gnd.n2325 585
R2712 gnd.n2324 gnd.n2323 585
R2713 gnd.n2322 gnd.n2321 585
R2714 gnd.n2320 gnd.n2319 585
R2715 gnd.n2318 gnd.n2317 585
R2716 gnd.n2316 gnd.n2315 585
R2717 gnd.n2314 gnd.n2313 585
R2718 gnd.n2312 gnd.n2311 585
R2719 gnd.n2310 gnd.n2309 585
R2720 gnd.n2308 gnd.n2307 585
R2721 gnd.n2306 gnd.n2305 585
R2722 gnd.n2304 gnd.n2303 585
R2723 gnd.n2296 gnd.n2293 585
R2724 gnd.n2299 gnd.n884 585
R2725 gnd.n4444 gnd.n884 585
R2726 gnd.n2790 gnd.n2789 585
R2727 gnd.n2034 gnd.n2026 585
R2728 gnd.n2797 gnd.n2023 585
R2729 gnd.n2798 gnd.n2022 585
R2730 gnd.n2048 gnd.n2016 585
R2731 gnd.n2805 gnd.n2015 585
R2732 gnd.n2806 gnd.n2014 585
R2733 gnd.n2046 gnd.n2006 585
R2734 gnd.n2813 gnd.n2005 585
R2735 gnd.n2814 gnd.n2004 585
R2736 gnd.n2043 gnd.n1998 585
R2737 gnd.n2821 gnd.n1997 585
R2738 gnd.n2822 gnd.n1996 585
R2739 gnd.n2041 gnd.n1989 585
R2740 gnd.n2829 gnd.n1988 585
R2741 gnd.n2830 gnd.n1987 585
R2742 gnd.n2038 gnd.n1986 585
R2743 gnd.n2037 gnd.n2036 585
R2744 gnd.n1197 gnd.n1195 585
R2745 gnd.n2787 gnd.n1195 585
R2746 gnd.n2118 gnd.n1193 585
R2747 gnd.n4206 gnd.n1193 585
R2748 gnd.n2579 gnd.n2578 585
R2749 gnd.n2580 gnd.n2579 585
R2750 gnd.n2117 gnd.n1183 585
R2751 gnd.n4212 gnd.n1183 585
R2752 gnd.n2538 gnd.n2537 585
R2753 gnd.n2537 gnd.n2536 585
R2754 gnd.n2120 gnd.n1172 585
R2755 gnd.n4218 gnd.n1172 585
R2756 gnd.n2526 gnd.n2525 585
R2757 gnd.n2527 gnd.n2526 585
R2758 gnd.n2124 gnd.n1161 585
R2759 gnd.n4224 gnd.n1161 585
R2760 gnd.n2521 gnd.n2520 585
R2761 gnd.n2520 gnd.n2519 585
R2762 gnd.n2126 gnd.n1151 585
R2763 gnd.n4230 gnd.n1151 585
R2764 gnd.n2461 gnd.n2460 585
R2765 gnd.n2460 gnd.n2459 585
R2766 gnd.n2146 gnd.n1140 585
R2767 gnd.n4236 gnd.n1140 585
R2768 gnd.n2465 gnd.n2145 585
R2769 gnd.n2447 gnd.n2145 585
R2770 gnd.n2466 gnd.n1130 585
R2771 gnd.n4242 gnd.n1130 585
R2772 gnd.n2467 gnd.n2144 585
R2773 gnd.n2442 gnd.n2144 585
R2774 gnd.n2141 gnd.n1119 585
R2775 gnd.n4248 gnd.n1119 585
R2776 gnd.n2472 gnd.n2471 585
R2777 gnd.n2473 gnd.n2472 585
R2778 gnd.n2140 gnd.n1109 585
R2779 gnd.n4254 gnd.n1109 585
R2780 gnd.n2433 gnd.n2432 585
R2781 gnd.n2434 gnd.n2433 585
R2782 gnd.n2153 gnd.n1098 585
R2783 gnd.n4260 gnd.n1098 585
R2784 gnd.n2428 gnd.n2427 585
R2785 gnd.n2427 gnd.n2426 585
R2786 gnd.n2155 gnd.n1088 585
R2787 gnd.n4266 gnd.n1088 585
R2788 gnd.n2416 gnd.n2415 585
R2789 gnd.n2417 gnd.n2416 585
R2790 gnd.n2187 gnd.n1078 585
R2791 gnd.n4272 gnd.n1078 585
R2792 gnd.n2411 gnd.n2410 585
R2793 gnd.n2410 gnd.n1069 585
R2794 gnd.n2409 gnd.n1068 585
R2795 gnd.n4278 gnd.n1068 585
R2796 gnd.n2408 gnd.n2258 585
R2797 gnd.n2258 gnd.n2257 585
R2798 gnd.n2189 gnd.n1061 585
R2799 gnd.n4285 gnd.n1061 585
R2800 gnd.n2403 gnd.n2402 585
R2801 gnd.n2402 gnd.n1059 585
R2802 gnd.n2401 gnd.n1051 585
R2803 gnd.n4291 gnd.n1051 585
R2804 gnd.n2400 gnd.n2399 585
R2805 gnd.n2399 gnd.n1044 585
R2806 gnd.n2260 gnd.n1043 585
R2807 gnd.n4297 gnd.n1043 585
R2808 gnd.n2395 gnd.n2394 585
R2809 gnd.n2394 gnd.n1034 585
R2810 gnd.n2393 gnd.n1033 585
R2811 gnd.n4303 gnd.n1033 585
R2812 gnd.n2392 gnd.n2391 585
R2813 gnd.n2391 gnd.n1031 585
R2814 gnd.n2262 gnd.n1023 585
R2815 gnd.n4309 gnd.n1023 585
R2816 gnd.n2387 gnd.n2386 585
R2817 gnd.n2386 gnd.n1021 585
R2818 gnd.n2385 gnd.n1013 585
R2819 gnd.n4315 gnd.n1013 585
R2820 gnd.n2384 gnd.n2383 585
R2821 gnd.n2383 gnd.n1004 585
R2822 gnd.n2264 gnd.n1003 585
R2823 gnd.n4321 gnd.n1003 585
R2824 gnd.n2379 gnd.n2378 585
R2825 gnd.n2378 gnd.n994 585
R2826 gnd.n2377 gnd.n993 585
R2827 gnd.n4327 gnd.n993 585
R2828 gnd.n2376 gnd.n2375 585
R2829 gnd.n2375 gnd.n991 585
R2830 gnd.n2266 gnd.n983 585
R2831 gnd.n4333 gnd.n983 585
R2832 gnd.n2371 gnd.n2370 585
R2833 gnd.n2370 gnd.n981 585
R2834 gnd.n2369 gnd.n973 585
R2835 gnd.n4339 gnd.n973 585
R2836 gnd.n2368 gnd.n2367 585
R2837 gnd.n2367 gnd.n964 585
R2838 gnd.n2268 gnd.n963 585
R2839 gnd.n4345 gnd.n963 585
R2840 gnd.n2363 gnd.n2362 585
R2841 gnd.n2362 gnd.n953 585
R2842 gnd.n2361 gnd.n952 585
R2843 gnd.n4351 gnd.n952 585
R2844 gnd.n2360 gnd.n2359 585
R2845 gnd.n2359 gnd.n941 585
R2846 gnd.n2270 gnd.n940 585
R2847 gnd.n4357 gnd.n940 585
R2848 gnd.n2355 gnd.n2354 585
R2849 gnd.n2354 gnd.n939 585
R2850 gnd.n2353 gnd.n2272 585
R2851 gnd.n2353 gnd.n2352 585
R2852 gnd.n2297 gnd.n2273 585
R2853 gnd.n2273 gnd.n885 585
R2854 gnd.n6918 gnd.n103 585
R2855 gnd.n7014 gnd.n103 585
R2856 gnd.n6919 gnd.n6849 585
R2857 gnd.n6849 gnd.n100 585
R2858 gnd.n6920 gnd.n182 585
R2859 gnd.n6934 gnd.n182 585
R2860 gnd.n193 gnd.n191 585
R2861 gnd.n191 gnd.n181 585
R2862 gnd.n6925 gnd.n6924 585
R2863 gnd.n6926 gnd.n6925 585
R2864 gnd.n192 gnd.n190 585
R2865 gnd.n190 gnd.n188 585
R2866 gnd.n6845 gnd.n6844 585
R2867 gnd.n6844 gnd.n6843 585
R2868 gnd.n196 gnd.n195 585
R2869 gnd.n6718 gnd.n196 585
R2870 gnd.n6834 gnd.n6833 585
R2871 gnd.n6835 gnd.n6834 585
R2872 gnd.n207 gnd.n206 585
R2873 gnd.n206 gnd.n203 585
R2874 gnd.n6829 gnd.n6828 585
R2875 gnd.n6828 gnd.n6827 585
R2876 gnd.n210 gnd.n209 585
R2877 gnd.n212 gnd.n210 585
R2878 gnd.n6818 gnd.n6817 585
R2879 gnd.n6819 gnd.n6818 585
R2880 gnd.n222 gnd.n221 585
R2881 gnd.n221 gnd.n219 585
R2882 gnd.n6813 gnd.n6812 585
R2883 gnd.n6812 gnd.n6811 585
R2884 gnd.n225 gnd.n224 585
R2885 gnd.n235 gnd.n225 585
R2886 gnd.n6802 gnd.n6801 585
R2887 gnd.n6803 gnd.n6802 585
R2888 gnd.n237 gnd.n236 585
R2889 gnd.n236 gnd.n232 585
R2890 gnd.n6797 gnd.n6796 585
R2891 gnd.n6796 gnd.n6795 585
R2892 gnd.n240 gnd.n239 585
R2893 gnd.n242 gnd.n240 585
R2894 gnd.n6786 gnd.n6785 585
R2895 gnd.n6787 gnd.n6786 585
R2896 gnd.n252 gnd.n251 585
R2897 gnd.n251 gnd.n249 585
R2898 gnd.n6781 gnd.n6780 585
R2899 gnd.n6780 gnd.n6779 585
R2900 gnd.n255 gnd.n254 585
R2901 gnd.n288 gnd.n255 585
R2902 gnd.n6758 gnd.n6757 585
R2903 gnd.n6757 gnd.n6756 585
R2904 gnd.n6759 gnd.n284 585
R2905 gnd.n285 gnd.n284 585
R2906 gnd.n6749 gnd.n281 585
R2907 gnd.n6750 gnd.n6749 585
R2908 gnd.n6764 gnd.n280 585
R2909 gnd.n292 gnd.n280 585
R2910 gnd.n6765 gnd.n279 585
R2911 gnd.n6677 gnd.n279 585
R2912 gnd.n6766 gnd.n278 585
R2913 gnd.n6680 gnd.n278 585
R2914 gnd.n275 gnd.n273 585
R2915 gnd.n300 gnd.n273 585
R2916 gnd.n6771 gnd.n6770 585
R2917 gnd.n6772 gnd.n6771 585
R2918 gnd.n274 gnd.n272 585
R2919 gnd.n333 gnd.n272 585
R2920 gnd.n6645 gnd.n6644 585
R2921 gnd.n6644 gnd.n6643 585
R2922 gnd.n6646 gnd.n316 585
R2923 gnd.n6662 gnd.n316 585
R2924 gnd.n329 gnd.n327 585
R2925 gnd.n4010 gnd.n327 585
R2926 gnd.n6651 gnd.n6650 585
R2927 gnd.n6652 gnd.n6651 585
R2928 gnd.n328 gnd.n326 585
R2929 gnd.n3993 gnd.n326 585
R2930 gnd.n4030 gnd.n4029 585
R2931 gnd.n4029 gnd.n4028 585
R2932 gnd.n4033 gnd.n1358 585
R2933 gnd.n1371 gnd.n1358 585
R2934 gnd.n4034 gnd.n1357 585
R2935 gnd.n4020 gnd.n1357 585
R2936 gnd.n4035 gnd.n1356 585
R2937 gnd.n3958 gnd.n1356 585
R2938 gnd.n1420 gnd.n1354 585
R2939 gnd.n1421 gnd.n1420 585
R2940 gnd.n4039 gnd.n1353 585
R2941 gnd.n3977 gnd.n1353 585
R2942 gnd.n4040 gnd.n1352 585
R2943 gnd.n1410 gnd.n1352 585
R2944 gnd.n4041 gnd.n1351 585
R2945 gnd.n3967 gnd.n1351 585
R2946 gnd.n3921 gnd.n1349 585
R2947 gnd.n3922 gnd.n3921 585
R2948 gnd.n4045 gnd.n1348 585
R2949 gnd.n3938 gnd.n1348 585
R2950 gnd.n4046 gnd.n1347 585
R2951 gnd.n1438 gnd.n1347 585
R2952 gnd.n4047 gnd.n1346 585
R2953 gnd.n3930 gnd.n1346 585
R2954 gnd.n1343 gnd.n1341 585
R2955 gnd.n3897 gnd.n1341 585
R2956 gnd.n4052 gnd.n4051 585
R2957 gnd.n4053 gnd.n4052 585
R2958 gnd.n1342 gnd.n1340 585
R2959 gnd.n3905 gnd.n1340 585
R2960 gnd.n3446 gnd.n1328 585
R2961 gnd.n4059 gnd.n1328 585
R2962 gnd.n3450 gnd.n3449 585
R2963 gnd.n3452 gnd.n3443 585
R2964 gnd.n3455 gnd.n3454 585
R2965 gnd.n3436 gnd.n3435 585
R2966 gnd.n3469 gnd.n3468 585
R2967 gnd.n3471 gnd.n3434 585
R2968 gnd.n3474 gnd.n3473 585
R2969 gnd.n3427 gnd.n3426 585
R2970 gnd.n3488 gnd.n3487 585
R2971 gnd.n3490 gnd.n3425 585
R2972 gnd.n3493 gnd.n3492 585
R2973 gnd.n3418 gnd.n3417 585
R2974 gnd.n3507 gnd.n3506 585
R2975 gnd.n3509 gnd.n3416 585
R2976 gnd.n3512 gnd.n3511 585
R2977 gnd.n3409 gnd.n3408 585
R2978 gnd.n3528 gnd.n3527 585
R2979 gnd.n3530 gnd.n3407 585
R2980 gnd.n3532 gnd.n3531 585
R2981 gnd.n3531 gnd.n1316 585
R2982 gnd.n6889 gnd.n99 585
R2983 gnd.n6890 gnd.n6887 585
R2984 gnd.n6891 gnd.n6883 585
R2985 gnd.n6881 gnd.n6879 585
R2986 gnd.n6895 gnd.n6878 585
R2987 gnd.n6896 gnd.n6876 585
R2988 gnd.n6897 gnd.n6875 585
R2989 gnd.n6873 gnd.n6871 585
R2990 gnd.n6901 gnd.n6870 585
R2991 gnd.n6902 gnd.n6868 585
R2992 gnd.n6903 gnd.n6867 585
R2993 gnd.n6865 gnd.n6863 585
R2994 gnd.n6907 gnd.n6862 585
R2995 gnd.n6908 gnd.n6860 585
R2996 gnd.n6909 gnd.n6859 585
R2997 gnd.n6857 gnd.n6855 585
R2998 gnd.n6913 gnd.n6854 585
R2999 gnd.n6914 gnd.n6852 585
R3000 gnd.n6915 gnd.n6851 585
R3001 gnd.n6851 gnd.n102 585
R3002 gnd.n7016 gnd.n7015 585
R3003 gnd.n7015 gnd.n7014 585
R3004 gnd.n7017 gnd.n97 585
R3005 gnd.n100 gnd.n97 585
R3006 gnd.n7018 gnd.n96 585
R3007 gnd.n6934 gnd.n96 585
R3008 gnd.n180 gnd.n94 585
R3009 gnd.n181 gnd.n180 585
R3010 gnd.n7022 gnd.n93 585
R3011 gnd.n6926 gnd.n93 585
R3012 gnd.n7023 gnd.n92 585
R3013 gnd.n188 gnd.n92 585
R3014 gnd.n7024 gnd.n91 585
R3015 gnd.n6843 gnd.n91 585
R3016 gnd.n6717 gnd.n89 585
R3017 gnd.n6718 gnd.n6717 585
R3018 gnd.n7028 gnd.n88 585
R3019 gnd.n6835 gnd.n88 585
R3020 gnd.n7029 gnd.n87 585
R3021 gnd.n203 gnd.n87 585
R3022 gnd.n7030 gnd.n86 585
R3023 gnd.n6827 gnd.n86 585
R3024 gnd.n211 gnd.n84 585
R3025 gnd.n212 gnd.n211 585
R3026 gnd.n7034 gnd.n83 585
R3027 gnd.n6819 gnd.n83 585
R3028 gnd.n7035 gnd.n82 585
R3029 gnd.n219 gnd.n82 585
R3030 gnd.n7036 gnd.n81 585
R3031 gnd.n6811 gnd.n81 585
R3032 gnd.n234 gnd.n79 585
R3033 gnd.n235 gnd.n234 585
R3034 gnd.n7040 gnd.n78 585
R3035 gnd.n6803 gnd.n78 585
R3036 gnd.n7041 gnd.n77 585
R3037 gnd.n232 gnd.n77 585
R3038 gnd.n7042 gnd.n76 585
R3039 gnd.n6795 gnd.n76 585
R3040 gnd.n241 gnd.n74 585
R3041 gnd.n242 gnd.n241 585
R3042 gnd.n7046 gnd.n73 585
R3043 gnd.n6787 gnd.n73 585
R3044 gnd.n7047 gnd.n72 585
R3045 gnd.n249 gnd.n72 585
R3046 gnd.n7048 gnd.n71 585
R3047 gnd.n6779 gnd.n71 585
R3048 gnd.n287 gnd.n69 585
R3049 gnd.n288 gnd.n287 585
R3050 gnd.n7052 gnd.n68 585
R3051 gnd.n6756 gnd.n68 585
R3052 gnd.n7053 gnd.n67 585
R3053 gnd.n285 gnd.n67 585
R3054 gnd.n7054 gnd.n66 585
R3055 gnd.n6750 gnd.n66 585
R3056 gnd.n304 gnd.n65 585
R3057 gnd.n304 gnd.n292 585
R3058 gnd.n6676 gnd.n6675 585
R3059 gnd.n6677 gnd.n6676 585
R3060 gnd.n305 gnd.n301 585
R3061 gnd.n6680 gnd.n301 585
R3062 gnd.n6671 gnd.n6670 585
R3063 gnd.n6670 gnd.n300 585
R3064 gnd.n6669 gnd.n271 585
R3065 gnd.n6772 gnd.n271 585
R3066 gnd.n6668 gnd.n308 585
R3067 gnd.n333 gnd.n308 585
R3068 gnd.n312 gnd.n307 585
R3069 gnd.n6643 gnd.n312 585
R3070 gnd.n6664 gnd.n6663 585
R3071 gnd.n6663 gnd.n6662 585
R3072 gnd.n311 gnd.n310 585
R3073 gnd.n4010 gnd.n311 585
R3074 gnd.n1390 gnd.n325 585
R3075 gnd.n6652 gnd.n325 585
R3076 gnd.n3992 gnd.n3991 585
R3077 gnd.n3993 gnd.n3992 585
R3078 gnd.n1389 gnd.n1361 585
R3079 gnd.n4028 gnd.n1361 585
R3080 gnd.n3986 gnd.n3985 585
R3081 gnd.n3985 gnd.n1371 585
R3082 gnd.n3984 gnd.n1370 585
R3083 gnd.n4020 gnd.n1370 585
R3084 gnd.n3983 gnd.n1393 585
R3085 gnd.n3958 gnd.n1393 585
R3086 gnd.n1397 gnd.n1392 585
R3087 gnd.n1421 gnd.n1397 585
R3088 gnd.n3979 gnd.n3978 585
R3089 gnd.n3978 gnd.n3977 585
R3090 gnd.n1396 gnd.n1395 585
R3091 gnd.n1410 gnd.n1396 585
R3092 gnd.n1455 gnd.n1409 585
R3093 gnd.n3967 gnd.n1409 585
R3094 gnd.n3920 gnd.n3919 585
R3095 gnd.n3922 gnd.n3920 585
R3096 gnd.n1454 gnd.n1431 585
R3097 gnd.n3938 gnd.n1431 585
R3098 gnd.n3914 gnd.n3913 585
R3099 gnd.n3913 gnd.n1438 585
R3100 gnd.n3912 gnd.n1437 585
R3101 gnd.n3930 gnd.n1437 585
R3102 gnd.n3911 gnd.n1458 585
R3103 gnd.n3897 gnd.n1458 585
R3104 gnd.n1457 gnd.n1338 585
R3105 gnd.n4053 gnd.n1338 585
R3106 gnd.n3907 gnd.n3906 585
R3107 gnd.n3906 gnd.n3905 585
R3108 gnd.n1460 gnd.n1326 585
R3109 gnd.n4059 gnd.n1326 585
R3110 gnd.n5890 gnd.n5889 585
R3111 gnd.n5889 gnd.n5888 585
R3112 gnd.n5891 gnd.n848 585
R3113 gnd.n5798 gnd.n848 585
R3114 gnd.n5893 gnd.n5892 585
R3115 gnd.n5894 gnd.n5893 585
R3116 gnd.n849 gnd.n847 585
R3117 gnd.n4805 gnd.n847 585
R3118 gnd.n5790 gnd.n5789 585
R3119 gnd.n5791 gnd.n5790 585
R3120 gnd.n4536 gnd.n4535 585
R3121 gnd.n5771 gnd.n4535 585
R3122 gnd.n5764 gnd.n5763 585
R3123 gnd.n5763 gnd.n4812 585
R3124 gnd.n5762 gnd.n4816 585
R3125 gnd.n5762 gnd.n5761 585
R3126 gnd.n5747 gnd.n4817 585
R3127 gnd.n4832 gnd.n4817 585
R3128 gnd.n5749 gnd.n5748 585
R3129 gnd.n5750 gnd.n5749 585
R3130 gnd.n4826 gnd.n4825 585
R3131 gnd.n5728 gnd.n4825 585
R3132 gnd.n5719 gnd.n5718 585
R3133 gnd.n5718 gnd.n4839 585
R3134 gnd.n5717 gnd.n4843 585
R3135 gnd.n5717 gnd.n5716 585
R3136 gnd.n5702 gnd.n4844 585
R3137 gnd.n4852 gnd.n4844 585
R3138 gnd.n5704 gnd.n5703 585
R3139 gnd.n5705 gnd.n5704 585
R3140 gnd.n4855 gnd.n4854 585
R3141 gnd.n4862 gnd.n4854 585
R3142 gnd.n5680 gnd.n5679 585
R3143 gnd.n5681 gnd.n5680 585
R3144 gnd.n4873 gnd.n4872 585
R3145 gnd.n5671 gnd.n4872 585
R3146 gnd.n5658 gnd.n4889 585
R3147 gnd.n4889 gnd.n4881 585
R3148 gnd.n5660 gnd.n5659 585
R3149 gnd.n5661 gnd.n5660 585
R3150 gnd.n4890 gnd.n4888 585
R3151 gnd.n4894 gnd.n4888 585
R3152 gnd.n5639 gnd.n5638 585
R3153 gnd.n5640 gnd.n5639 585
R3154 gnd.n4906 gnd.n4905 585
R3155 gnd.n4905 gnd.n4901 585
R3156 gnd.n5629 gnd.n5628 585
R3157 gnd.n5630 gnd.n5629 585
R3158 gnd.n4914 gnd.n4913 585
R3159 gnd.n4918 gnd.n4913 585
R3160 gnd.n5607 gnd.n4930 585
R3161 gnd.n5272 gnd.n4930 585
R3162 gnd.n5609 gnd.n5608 585
R3163 gnd.n5610 gnd.n5609 585
R3164 gnd.n4931 gnd.n4929 585
R3165 gnd.n4929 gnd.n4925 585
R3166 gnd.n5598 gnd.n5597 585
R3167 gnd.n5599 gnd.n5598 585
R3168 gnd.n4939 gnd.n4938 585
R3169 gnd.n5280 gnd.n4938 585
R3170 gnd.n5576 gnd.n4955 585
R3171 gnd.n4955 gnd.n4943 585
R3172 gnd.n5578 gnd.n5577 585
R3173 gnd.n5579 gnd.n5578 585
R3174 gnd.n4956 gnd.n4954 585
R3175 gnd.n4954 gnd.n4950 585
R3176 gnd.n5567 gnd.n5566 585
R3177 gnd.n5568 gnd.n5567 585
R3178 gnd.n4964 gnd.n4963 585
R3179 gnd.n4969 gnd.n4963 585
R3180 gnd.n5545 gnd.n4981 585
R3181 gnd.n4981 gnd.n4968 585
R3182 gnd.n5547 gnd.n5546 585
R3183 gnd.n5548 gnd.n5547 585
R3184 gnd.n4982 gnd.n4980 585
R3185 gnd.n4980 gnd.n4976 585
R3186 gnd.n5536 gnd.n5535 585
R3187 gnd.n5537 gnd.n5536 585
R3188 gnd.n4989 gnd.n4988 585
R3189 gnd.n4994 gnd.n4988 585
R3190 gnd.n5514 gnd.n5007 585
R3191 gnd.n5007 gnd.n4993 585
R3192 gnd.n5516 gnd.n5515 585
R3193 gnd.n5517 gnd.n5516 585
R3194 gnd.n5008 gnd.n5006 585
R3195 gnd.n5006 gnd.n5002 585
R3196 gnd.n5505 gnd.n5504 585
R3197 gnd.n5506 gnd.n5505 585
R3198 gnd.n5015 gnd.n5014 585
R3199 gnd.n5020 gnd.n5014 585
R3200 gnd.n5483 gnd.n5033 585
R3201 gnd.n5033 gnd.n5019 585
R3202 gnd.n5485 gnd.n5484 585
R3203 gnd.n5486 gnd.n5485 585
R3204 gnd.n5034 gnd.n5032 585
R3205 gnd.n5032 gnd.n5028 585
R3206 gnd.n5474 gnd.n5473 585
R3207 gnd.n5475 gnd.n5474 585
R3208 gnd.n5042 gnd.n5041 585
R3209 gnd.n5364 gnd.n5041 585
R3210 gnd.n5452 gnd.n5058 585
R3211 gnd.n5058 gnd.n5046 585
R3212 gnd.n5454 gnd.n5453 585
R3213 gnd.n5455 gnd.n5454 585
R3214 gnd.n5059 gnd.n5057 585
R3215 gnd.n5057 gnd.n5053 585
R3216 gnd.n5443 gnd.n5442 585
R3217 gnd.n5444 gnd.n5443 585
R3218 gnd.n5066 gnd.n5065 585
R3219 gnd.n5065 gnd.n5063 585
R3220 gnd.n5437 gnd.n5436 585
R3221 gnd.n5436 gnd.n5435 585
R3222 gnd.n5070 gnd.n5069 585
R3223 gnd.n5078 gnd.n5070 585
R3224 gnd.n5231 gnd.n5230 585
R3225 gnd.n5232 gnd.n5231 585
R3226 gnd.n5080 gnd.n5079 585
R3227 gnd.n5079 gnd.n5077 585
R3228 gnd.n5226 gnd.n5225 585
R3229 gnd.n5225 gnd.n5224 585
R3230 gnd.n5083 gnd.n5082 585
R3231 gnd.n5084 gnd.n5083 585
R3232 gnd.n5215 gnd.n5214 585
R3233 gnd.n5216 gnd.n5215 585
R3234 gnd.n5092 gnd.n5091 585
R3235 gnd.n5091 gnd.n5090 585
R3236 gnd.n5210 gnd.n5209 585
R3237 gnd.n5209 gnd.n5208 585
R3238 gnd.n5095 gnd.n5094 585
R3239 gnd.n5096 gnd.n5095 585
R3240 gnd.n5199 gnd.n5198 585
R3241 gnd.n5200 gnd.n5199 585
R3242 gnd.n5195 gnd.n5102 585
R3243 gnd.n5194 gnd.n5193 585
R3244 gnd.n5191 gnd.n5104 585
R3245 gnd.n5191 gnd.n5101 585
R3246 gnd.n5190 gnd.n5189 585
R3247 gnd.n5188 gnd.n5187 585
R3248 gnd.n5186 gnd.n5109 585
R3249 gnd.n5184 gnd.n5183 585
R3250 gnd.n5182 gnd.n5110 585
R3251 gnd.n5181 gnd.n5180 585
R3252 gnd.n5178 gnd.n5115 585
R3253 gnd.n5176 gnd.n5175 585
R3254 gnd.n5174 gnd.n5116 585
R3255 gnd.n5173 gnd.n5172 585
R3256 gnd.n5170 gnd.n5121 585
R3257 gnd.n5168 gnd.n5167 585
R3258 gnd.n5166 gnd.n5122 585
R3259 gnd.n5165 gnd.n5164 585
R3260 gnd.n5162 gnd.n5127 585
R3261 gnd.n5160 gnd.n5159 585
R3262 gnd.n5158 gnd.n5128 585
R3263 gnd.n5157 gnd.n5156 585
R3264 gnd.n5154 gnd.n5133 585
R3265 gnd.n5152 gnd.n5151 585
R3266 gnd.n5149 gnd.n5134 585
R3267 gnd.n5148 gnd.n5147 585
R3268 gnd.n5145 gnd.n5143 585
R3269 gnd.n5141 gnd.n5100 585
R3270 gnd.n5806 gnd.n5805 585
R3271 gnd.n5807 gnd.n4523 585
R3272 gnd.n5809 gnd.n5808 585
R3273 gnd.n5811 gnd.n4522 585
R3274 gnd.n5813 gnd.n5812 585
R3275 gnd.n5814 gnd.n4513 585
R3276 gnd.n5816 gnd.n5815 585
R3277 gnd.n5818 gnd.n4511 585
R3278 gnd.n5820 gnd.n5819 585
R3279 gnd.n5821 gnd.n4506 585
R3280 gnd.n5823 gnd.n5822 585
R3281 gnd.n5825 gnd.n4504 585
R3282 gnd.n5827 gnd.n5826 585
R3283 gnd.n5828 gnd.n4499 585
R3284 gnd.n5830 gnd.n5829 585
R3285 gnd.n5832 gnd.n4497 585
R3286 gnd.n5834 gnd.n5833 585
R3287 gnd.n5835 gnd.n4492 585
R3288 gnd.n5837 gnd.n5836 585
R3289 gnd.n5839 gnd.n4490 585
R3290 gnd.n5841 gnd.n5840 585
R3291 gnd.n5842 gnd.n4485 585
R3292 gnd.n5844 gnd.n5843 585
R3293 gnd.n5846 gnd.n4483 585
R3294 gnd.n5848 gnd.n5847 585
R3295 gnd.n5849 gnd.n4481 585
R3296 gnd.n5850 gnd.n853 585
R3297 gnd.n4445 gnd.n853 585
R3298 gnd.n5801 gnd.n855 585
R3299 gnd.n5888 gnd.n855 585
R3300 gnd.n5800 gnd.n5799 585
R3301 gnd.n5799 gnd.n5798 585
R3302 gnd.n5797 gnd.n845 585
R3303 gnd.n5894 gnd.n845 585
R3304 gnd.n4532 gnd.n4528 585
R3305 gnd.n4805 gnd.n4532 585
R3306 gnd.n5793 gnd.n5792 585
R3307 gnd.n5792 gnd.n5791 585
R3308 gnd.n4531 gnd.n4530 585
R3309 gnd.n5771 gnd.n4531 585
R3310 gnd.n5757 gnd.n4820 585
R3311 gnd.n4820 gnd.n4812 585
R3312 gnd.n5759 gnd.n5758 585
R3313 gnd.n5761 gnd.n5759 585
R3314 gnd.n4821 gnd.n4819 585
R3315 gnd.n4832 gnd.n4819 585
R3316 gnd.n5752 gnd.n5751 585
R3317 gnd.n5751 gnd.n5750 585
R3318 gnd.n4824 gnd.n4823 585
R3319 gnd.n5728 gnd.n4824 585
R3320 gnd.n5712 gnd.n4847 585
R3321 gnd.n4847 gnd.n4839 585
R3322 gnd.n5714 gnd.n5713 585
R3323 gnd.n5716 gnd.n5714 585
R3324 gnd.n4848 gnd.n4846 585
R3325 gnd.n4852 gnd.n4846 585
R3326 gnd.n5707 gnd.n5706 585
R3327 gnd.n5706 gnd.n5705 585
R3328 gnd.n4851 gnd.n4850 585
R3329 gnd.n4862 gnd.n4851 585
R3330 gnd.n5668 gnd.n4870 585
R3331 gnd.n5681 gnd.n4870 585
R3332 gnd.n5670 gnd.n5669 585
R3333 gnd.n5671 gnd.n5670 585
R3334 gnd.n4883 gnd.n4882 585
R3335 gnd.n4882 gnd.n4881 585
R3336 gnd.n5663 gnd.n5662 585
R3337 gnd.n5662 gnd.n5661 585
R3338 gnd.n4886 gnd.n4885 585
R3339 gnd.n4894 gnd.n4886 585
R3340 gnd.n5266 gnd.n4903 585
R3341 gnd.n5640 gnd.n4903 585
R3342 gnd.n5268 gnd.n5267 585
R3343 gnd.n5267 gnd.n4901 585
R3344 gnd.n5269 gnd.n4912 585
R3345 gnd.n5630 gnd.n4912 585
R3346 gnd.n5271 gnd.n5270 585
R3347 gnd.n5271 gnd.n4918 585
R3348 gnd.n5274 gnd.n5273 585
R3349 gnd.n5273 gnd.n5272 585
R3350 gnd.n5275 gnd.n4927 585
R3351 gnd.n5610 gnd.n4927 585
R3352 gnd.n5277 gnd.n5276 585
R3353 gnd.n5276 gnd.n4925 585
R3354 gnd.n5278 gnd.n4937 585
R3355 gnd.n5599 gnd.n4937 585
R3356 gnd.n5281 gnd.n5279 585
R3357 gnd.n5281 gnd.n5280 585
R3358 gnd.n5283 gnd.n5282 585
R3359 gnd.n5282 gnd.n4943 585
R3360 gnd.n5284 gnd.n4952 585
R3361 gnd.n5579 gnd.n4952 585
R3362 gnd.n5287 gnd.n5286 585
R3363 gnd.n5286 gnd.n4950 585
R3364 gnd.n5288 gnd.n4962 585
R3365 gnd.n5568 gnd.n4962 585
R3366 gnd.n5291 gnd.n5290 585
R3367 gnd.n5290 gnd.n4969 585
R3368 gnd.n5289 gnd.n5256 585
R3369 gnd.n5289 gnd.n4968 585
R3370 gnd.n5343 gnd.n4978 585
R3371 gnd.n5548 gnd.n4978 585
R3372 gnd.n5345 gnd.n5344 585
R3373 gnd.n5344 gnd.n4976 585
R3374 gnd.n5346 gnd.n4987 585
R3375 gnd.n5537 gnd.n4987 585
R3376 gnd.n5348 gnd.n5347 585
R3377 gnd.n5348 gnd.n4994 585
R3378 gnd.n5350 gnd.n5349 585
R3379 gnd.n5349 gnd.n4993 585
R3380 gnd.n5351 gnd.n5004 585
R3381 gnd.n5517 gnd.n5004 585
R3382 gnd.n5353 gnd.n5352 585
R3383 gnd.n5352 gnd.n5002 585
R3384 gnd.n5354 gnd.n5013 585
R3385 gnd.n5506 gnd.n5013 585
R3386 gnd.n5356 gnd.n5355 585
R3387 gnd.n5356 gnd.n5020 585
R3388 gnd.n5358 gnd.n5357 585
R3389 gnd.n5357 gnd.n5019 585
R3390 gnd.n5359 gnd.n5030 585
R3391 gnd.n5486 gnd.n5030 585
R3392 gnd.n5361 gnd.n5360 585
R3393 gnd.n5360 gnd.n5028 585
R3394 gnd.n5362 gnd.n5040 585
R3395 gnd.n5475 gnd.n5040 585
R3396 gnd.n5365 gnd.n5363 585
R3397 gnd.n5365 gnd.n5364 585
R3398 gnd.n5367 gnd.n5366 585
R3399 gnd.n5366 gnd.n5046 585
R3400 gnd.n5368 gnd.n5055 585
R3401 gnd.n5455 gnd.n5055 585
R3402 gnd.n5370 gnd.n5369 585
R3403 gnd.n5369 gnd.n5053 585
R3404 gnd.n5371 gnd.n5064 585
R3405 gnd.n5444 gnd.n5064 585
R3406 gnd.n5372 gnd.n5072 585
R3407 gnd.n5072 gnd.n5063 585
R3408 gnd.n5374 gnd.n5373 585
R3409 gnd.n5435 gnd.n5374 585
R3410 gnd.n5073 gnd.n5071 585
R3411 gnd.n5078 gnd.n5071 585
R3412 gnd.n5234 gnd.n5233 585
R3413 gnd.n5233 gnd.n5232 585
R3414 gnd.n5076 gnd.n5075 585
R3415 gnd.n5077 gnd.n5076 585
R3416 gnd.n5223 gnd.n5222 585
R3417 gnd.n5224 gnd.n5223 585
R3418 gnd.n5086 gnd.n5085 585
R3419 gnd.n5085 gnd.n5084 585
R3420 gnd.n5218 gnd.n5217 585
R3421 gnd.n5217 gnd.n5216 585
R3422 gnd.n5089 gnd.n5088 585
R3423 gnd.n5090 gnd.n5089 585
R3424 gnd.n5207 gnd.n5206 585
R3425 gnd.n5208 gnd.n5207 585
R3426 gnd.n5098 gnd.n5097 585
R3427 gnd.n5097 gnd.n5096 585
R3428 gnd.n5202 gnd.n5201 585
R3429 gnd.n5201 gnd.n5200 585
R3430 gnd.n5886 gnd.n5885 585
R3431 gnd.n5887 gnd.n5886 585
R3432 gnd.n4448 gnd.n4446 585
R3433 gnd.n4446 gnd.n854 585
R3434 gnd.n5780 gnd.n4807 585
R3435 gnd.n4807 gnd.n846 585
R3436 gnd.n5782 gnd.n5781 585
R3437 gnd.n5783 gnd.n5782 585
R3438 gnd.n4808 gnd.n4806 585
R3439 gnd.n4806 gnd.n4534 585
R3440 gnd.n5775 gnd.n5774 585
R3441 gnd.n5774 gnd.n4533 585
R3442 gnd.n5773 gnd.n4810 585
R3443 gnd.n5773 gnd.n5772 585
R3444 gnd.n5737 gnd.n4811 585
R3445 gnd.n5760 gnd.n4811 585
R3446 gnd.n5738 gnd.n4834 585
R3447 gnd.n4834 gnd.n4818 585
R3448 gnd.n5740 gnd.n5739 585
R3449 gnd.n5741 gnd.n5740 585
R3450 gnd.n4835 gnd.n4833 585
R3451 gnd.n5727 gnd.n4833 585
R3452 gnd.n5731 gnd.n5730 585
R3453 gnd.n5730 gnd.n5729 585
R3454 gnd.n4838 gnd.n4837 585
R3455 gnd.n5715 gnd.n4838 585
R3456 gnd.n5691 gnd.n5690 585
R3457 gnd.n5690 gnd.n4845 585
R3458 gnd.n5692 gnd.n4864 585
R3459 gnd.n4864 gnd.n4853 585
R3460 gnd.n5694 gnd.n5693 585
R3461 gnd.n5695 gnd.n5694 585
R3462 gnd.n4865 gnd.n4863 585
R3463 gnd.n4871 gnd.n4863 585
R3464 gnd.n5684 gnd.n5683 585
R3465 gnd.n5683 gnd.n5682 585
R3466 gnd.n4868 gnd.n4867 585
R3467 gnd.n5672 gnd.n4868 585
R3468 gnd.n5648 gnd.n4896 585
R3469 gnd.n4896 gnd.n4887 585
R3470 gnd.n5650 gnd.n5649 585
R3471 gnd.n5651 gnd.n5650 585
R3472 gnd.n4897 gnd.n4895 585
R3473 gnd.n4904 gnd.n4895 585
R3474 gnd.n5643 gnd.n5642 585
R3475 gnd.n5642 gnd.n5641 585
R3476 gnd.n4900 gnd.n4899 585
R3477 gnd.n5631 gnd.n4900 585
R3478 gnd.n5618 gnd.n4920 585
R3479 gnd.n4920 gnd.n4911 585
R3480 gnd.n5620 gnd.n5619 585
R3481 gnd.n5621 gnd.n5620 585
R3482 gnd.n4921 gnd.n4919 585
R3483 gnd.n4928 gnd.n4919 585
R3484 gnd.n5613 gnd.n5612 585
R3485 gnd.n5612 gnd.n5611 585
R3486 gnd.n4924 gnd.n4923 585
R3487 gnd.n5600 gnd.n4924 585
R3488 gnd.n5587 gnd.n4945 585
R3489 gnd.n4945 gnd.n4936 585
R3490 gnd.n5589 gnd.n5588 585
R3491 gnd.n5590 gnd.n5589 585
R3492 gnd.n4946 gnd.n4944 585
R3493 gnd.n4953 gnd.n4944 585
R3494 gnd.n5582 gnd.n5581 585
R3495 gnd.n5581 gnd.n5580 585
R3496 gnd.n4949 gnd.n4948 585
R3497 gnd.n5569 gnd.n4949 585
R3498 gnd.n5556 gnd.n4971 585
R3499 gnd.n4971 gnd.n4961 585
R3500 gnd.n5558 gnd.n5557 585
R3501 gnd.n5559 gnd.n5558 585
R3502 gnd.n4972 gnd.n4970 585
R3503 gnd.n4979 gnd.n4970 585
R3504 gnd.n5551 gnd.n5550 585
R3505 gnd.n5550 gnd.n5549 585
R3506 gnd.n4975 gnd.n4974 585
R3507 gnd.n5538 gnd.n4975 585
R3508 gnd.n5525 gnd.n4997 585
R3509 gnd.n4997 gnd.n4996 585
R3510 gnd.n5527 gnd.n5526 585
R3511 gnd.n5528 gnd.n5527 585
R3512 gnd.n4998 gnd.n4995 585
R3513 gnd.n5005 gnd.n4995 585
R3514 gnd.n5520 gnd.n5519 585
R3515 gnd.n5519 gnd.n5518 585
R3516 gnd.n5001 gnd.n5000 585
R3517 gnd.n5507 gnd.n5001 585
R3518 gnd.n5494 gnd.n5023 585
R3519 gnd.n5023 gnd.n5022 585
R3520 gnd.n5496 gnd.n5495 585
R3521 gnd.n5497 gnd.n5496 585
R3522 gnd.n5024 gnd.n5021 585
R3523 gnd.n5031 gnd.n5021 585
R3524 gnd.n5489 gnd.n5488 585
R3525 gnd.n5488 gnd.n5487 585
R3526 gnd.n5027 gnd.n5026 585
R3527 gnd.n5476 gnd.n5027 585
R3528 gnd.n5463 gnd.n5048 585
R3529 gnd.n5048 gnd.n5039 585
R3530 gnd.n5465 gnd.n5464 585
R3531 gnd.n5466 gnd.n5465 585
R3532 gnd.n5049 gnd.n5047 585
R3533 gnd.n5056 gnd.n5047 585
R3534 gnd.n5458 gnd.n5457 585
R3535 gnd.n5457 gnd.n5456 585
R3536 gnd.n5052 gnd.n5051 585
R3537 gnd.n5445 gnd.n5052 585
R3538 gnd.n5432 gnd.n5431 585
R3539 gnd.n5430 gnd.n5383 585
R3540 gnd.n5429 gnd.n5382 585
R3541 gnd.n5434 gnd.n5382 585
R3542 gnd.n5428 gnd.n5427 585
R3543 gnd.n5426 gnd.n5425 585
R3544 gnd.n5424 gnd.n5423 585
R3545 gnd.n5422 gnd.n5421 585
R3546 gnd.n5420 gnd.n5419 585
R3547 gnd.n5418 gnd.n5417 585
R3548 gnd.n5416 gnd.n5415 585
R3549 gnd.n5414 gnd.n5413 585
R3550 gnd.n5412 gnd.n5411 585
R3551 gnd.n5410 gnd.n5409 585
R3552 gnd.n5408 gnd.n5407 585
R3553 gnd.n5406 gnd.n5405 585
R3554 gnd.n5404 gnd.n5403 585
R3555 gnd.n5399 gnd.n5062 585
R3556 gnd.n5855 gnd.n5854 585
R3557 gnd.n5857 gnd.n4476 585
R3558 gnd.n5859 gnd.n5858 585
R3559 gnd.n5860 gnd.n4469 585
R3560 gnd.n5862 gnd.n5861 585
R3561 gnd.n5864 gnd.n4467 585
R3562 gnd.n5866 gnd.n5865 585
R3563 gnd.n5867 gnd.n4462 585
R3564 gnd.n5869 gnd.n5868 585
R3565 gnd.n5871 gnd.n4460 585
R3566 gnd.n5873 gnd.n5872 585
R3567 gnd.n5874 gnd.n4455 585
R3568 gnd.n5876 gnd.n5875 585
R3569 gnd.n5878 gnd.n4453 585
R3570 gnd.n5880 gnd.n5879 585
R3571 gnd.n5881 gnd.n4451 585
R3572 gnd.n5882 gnd.n4447 585
R3573 gnd.n4447 gnd.n4445 585
R3574 gnd.n4801 gnd.n856 585
R3575 gnd.n5887 gnd.n856 585
R3576 gnd.n4802 gnd.n4798 585
R3577 gnd.n4798 gnd.n854 585
R3578 gnd.n4804 gnd.n4803 585
R3579 gnd.n4804 gnd.n846 585
R3580 gnd.n5784 gnd.n4796 585
R3581 gnd.n5784 gnd.n5783 585
R3582 gnd.n5786 gnd.n5785 585
R3583 gnd.n5785 gnd.n4534 585
R3584 gnd.n4797 gnd.n4794 585
R3585 gnd.n4797 gnd.n4533 585
R3586 gnd.n5770 gnd.n5769 585
R3587 gnd.n5772 gnd.n5770 585
R3588 gnd.n4814 gnd.n4813 585
R3589 gnd.n5760 gnd.n4813 585
R3590 gnd.n5744 gnd.n5743 585
R3591 gnd.n5743 gnd.n4818 585
R3592 gnd.n5742 gnd.n4830 585
R3593 gnd.n5742 gnd.n5741 585
R3594 gnd.n5724 gnd.n4831 585
R3595 gnd.n5727 gnd.n4831 585
R3596 gnd.n5726 gnd.n5725 585
R3597 gnd.n5729 gnd.n5726 585
R3598 gnd.n4841 gnd.n4840 585
R3599 gnd.n5715 gnd.n4840 585
R3600 gnd.n5699 gnd.n5698 585
R3601 gnd.n5698 gnd.n4845 585
R3602 gnd.n5697 gnd.n4859 585
R3603 gnd.n5697 gnd.n4853 585
R3604 gnd.n5696 gnd.n4861 585
R3605 gnd.n5696 gnd.n5695 585
R3606 gnd.n5676 gnd.n4860 585
R3607 gnd.n4871 gnd.n4860 585
R3608 gnd.n5675 gnd.n4869 585
R3609 gnd.n5682 gnd.n4869 585
R3610 gnd.n5674 gnd.n5673 585
R3611 gnd.n5673 gnd.n5672 585
R3612 gnd.n4880 gnd.n4877 585
R3613 gnd.n4887 gnd.n4880 585
R3614 gnd.n5653 gnd.n5652 585
R3615 gnd.n5652 gnd.n5651 585
R3616 gnd.n4893 gnd.n4892 585
R3617 gnd.n4904 gnd.n4893 585
R3618 gnd.n5634 gnd.n4902 585
R3619 gnd.n5641 gnd.n4902 585
R3620 gnd.n5633 gnd.n5632 585
R3621 gnd.n5632 gnd.n5631 585
R3622 gnd.n4910 gnd.n4908 585
R3623 gnd.n4911 gnd.n4910 585
R3624 gnd.n5623 gnd.n5622 585
R3625 gnd.n5622 gnd.n5621 585
R3626 gnd.n4917 gnd.n4916 585
R3627 gnd.n4928 gnd.n4917 585
R3628 gnd.n5603 gnd.n4926 585
R3629 gnd.n5611 gnd.n4926 585
R3630 gnd.n5602 gnd.n5601 585
R3631 gnd.n5601 gnd.n5600 585
R3632 gnd.n4935 gnd.n4933 585
R3633 gnd.n4936 gnd.n4935 585
R3634 gnd.n5592 gnd.n5591 585
R3635 gnd.n5591 gnd.n5590 585
R3636 gnd.n4942 gnd.n4941 585
R3637 gnd.n4953 gnd.n4942 585
R3638 gnd.n5572 gnd.n4951 585
R3639 gnd.n5580 gnd.n4951 585
R3640 gnd.n5571 gnd.n5570 585
R3641 gnd.n5570 gnd.n5569 585
R3642 gnd.n4960 gnd.n4958 585
R3643 gnd.n4961 gnd.n4960 585
R3644 gnd.n5561 gnd.n5560 585
R3645 gnd.n5560 gnd.n5559 585
R3646 gnd.n4967 gnd.n4966 585
R3647 gnd.n4979 gnd.n4967 585
R3648 gnd.n5541 gnd.n4977 585
R3649 gnd.n5549 gnd.n4977 585
R3650 gnd.n5540 gnd.n5539 585
R3651 gnd.n5539 gnd.n5538 585
R3652 gnd.n4986 gnd.n4984 585
R3653 gnd.n4996 gnd.n4986 585
R3654 gnd.n5530 gnd.n5529 585
R3655 gnd.n5529 gnd.n5528 585
R3656 gnd.n4992 gnd.n4991 585
R3657 gnd.n5005 gnd.n4992 585
R3658 gnd.n5510 gnd.n5003 585
R3659 gnd.n5518 gnd.n5003 585
R3660 gnd.n5509 gnd.n5508 585
R3661 gnd.n5508 gnd.n5507 585
R3662 gnd.n5012 gnd.n5010 585
R3663 gnd.n5022 gnd.n5012 585
R3664 gnd.n5499 gnd.n5498 585
R3665 gnd.n5498 gnd.n5497 585
R3666 gnd.n5018 gnd.n5017 585
R3667 gnd.n5031 gnd.n5018 585
R3668 gnd.n5479 gnd.n5029 585
R3669 gnd.n5487 gnd.n5029 585
R3670 gnd.n5478 gnd.n5477 585
R3671 gnd.n5477 gnd.n5476 585
R3672 gnd.n5038 gnd.n5036 585
R3673 gnd.n5039 gnd.n5038 585
R3674 gnd.n5468 gnd.n5467 585
R3675 gnd.n5467 gnd.n5466 585
R3676 gnd.n5045 gnd.n5044 585
R3677 gnd.n5056 gnd.n5045 585
R3678 gnd.n5448 gnd.n5054 585
R3679 gnd.n5456 gnd.n5054 585
R3680 gnd.n5447 gnd.n5446 585
R3681 gnd.n5446 gnd.n5445 585
R3682 gnd.n4208 gnd.n4207 585
R3683 gnd.n4207 gnd.n4206 585
R3684 gnd.n4209 gnd.n1185 585
R3685 gnd.n2580 gnd.n1185 585
R3686 gnd.n4211 gnd.n4210 585
R3687 gnd.n4212 gnd.n4211 585
R3688 gnd.n1169 gnd.n1168 585
R3689 gnd.n2536 gnd.n1169 585
R3690 gnd.n4220 gnd.n4219 585
R3691 gnd.n4219 gnd.n4218 585
R3692 gnd.n4221 gnd.n1163 585
R3693 gnd.n2527 gnd.n1163 585
R3694 gnd.n4223 gnd.n4222 585
R3695 gnd.n4224 gnd.n4223 585
R3696 gnd.n1148 gnd.n1147 585
R3697 gnd.n2519 gnd.n1148 585
R3698 gnd.n4232 gnd.n4231 585
R3699 gnd.n4231 gnd.n4230 585
R3700 gnd.n4233 gnd.n1142 585
R3701 gnd.n2459 gnd.n1142 585
R3702 gnd.n4235 gnd.n4234 585
R3703 gnd.n4236 gnd.n4235 585
R3704 gnd.n1127 gnd.n1126 585
R3705 gnd.n2447 gnd.n1127 585
R3706 gnd.n4244 gnd.n4243 585
R3707 gnd.n4243 gnd.n4242 585
R3708 gnd.n4245 gnd.n1121 585
R3709 gnd.n2442 gnd.n1121 585
R3710 gnd.n4247 gnd.n4246 585
R3711 gnd.n4248 gnd.n4247 585
R3712 gnd.n1106 gnd.n1105 585
R3713 gnd.n2473 gnd.n1106 585
R3714 gnd.n4256 gnd.n4255 585
R3715 gnd.n4255 gnd.n4254 585
R3716 gnd.n4257 gnd.n1100 585
R3717 gnd.n2434 gnd.n1100 585
R3718 gnd.n4259 gnd.n4258 585
R3719 gnd.n4260 gnd.n4259 585
R3720 gnd.n1085 gnd.n1084 585
R3721 gnd.n2426 gnd.n1085 585
R3722 gnd.n4268 gnd.n4267 585
R3723 gnd.n4267 gnd.n4266 585
R3724 gnd.n4269 gnd.n1080 585
R3725 gnd.n2417 gnd.n1080 585
R3726 gnd.n4271 gnd.n4270 585
R3727 gnd.n4272 gnd.n4271 585
R3728 gnd.n1081 gnd.n1065 585
R3729 gnd.n1069 gnd.n1065 585
R3730 gnd.n4280 gnd.n4279 585
R3731 gnd.n4279 gnd.n4278 585
R3732 gnd.n4281 gnd.n1062 585
R3733 gnd.n2257 gnd.n1062 585
R3734 gnd.n4284 gnd.n4283 585
R3735 gnd.n4285 gnd.n4284 585
R3736 gnd.n1063 gnd.n1049 585
R3737 gnd.n1059 gnd.n1049 585
R3738 gnd.n4293 gnd.n4292 585
R3739 gnd.n4292 gnd.n4291 585
R3740 gnd.n4294 gnd.n1045 585
R3741 gnd.n1045 gnd.n1044 585
R3742 gnd.n4296 gnd.n4295 585
R3743 gnd.n4297 gnd.n4296 585
R3744 gnd.n1030 gnd.n1029 585
R3745 gnd.n1034 gnd.n1030 585
R3746 gnd.n4305 gnd.n4304 585
R3747 gnd.n4304 gnd.n4303 585
R3748 gnd.n4306 gnd.n1024 585
R3749 gnd.n1031 gnd.n1024 585
R3750 gnd.n4308 gnd.n4307 585
R3751 gnd.n4309 gnd.n4308 585
R3752 gnd.n1011 gnd.n1010 585
R3753 gnd.n1021 gnd.n1011 585
R3754 gnd.n4317 gnd.n4316 585
R3755 gnd.n4316 gnd.n4315 585
R3756 gnd.n4318 gnd.n1005 585
R3757 gnd.n1005 gnd.n1004 585
R3758 gnd.n4320 gnd.n4319 585
R3759 gnd.n4321 gnd.n4320 585
R3760 gnd.n990 gnd.n989 585
R3761 gnd.n994 gnd.n990 585
R3762 gnd.n4329 gnd.n4328 585
R3763 gnd.n4328 gnd.n4327 585
R3764 gnd.n4330 gnd.n984 585
R3765 gnd.n991 gnd.n984 585
R3766 gnd.n4332 gnd.n4331 585
R3767 gnd.n4333 gnd.n4332 585
R3768 gnd.n971 gnd.n970 585
R3769 gnd.n981 gnd.n971 585
R3770 gnd.n4341 gnd.n4340 585
R3771 gnd.n4340 gnd.n4339 585
R3772 gnd.n4342 gnd.n965 585
R3773 gnd.n965 gnd.n964 585
R3774 gnd.n4344 gnd.n4343 585
R3775 gnd.n4345 gnd.n4344 585
R3776 gnd.n950 gnd.n949 585
R3777 gnd.n953 gnd.n950 585
R3778 gnd.n4353 gnd.n4352 585
R3779 gnd.n4352 gnd.n4351 585
R3780 gnd.n4354 gnd.n944 585
R3781 gnd.n944 gnd.n941 585
R3782 gnd.n4356 gnd.n4355 585
R3783 gnd.n4357 gnd.n4356 585
R3784 gnd.n945 gnd.n943 585
R3785 gnd.n943 gnd.n939 585
R3786 gnd.n2351 gnd.n2350 585
R3787 gnd.n2352 gnd.n2351 585
R3788 gnd.n2346 gnd.n888 585
R3789 gnd.n888 gnd.n885 585
R3790 gnd.n4442 gnd.n4441 585
R3791 gnd.n4440 gnd.n887 585
R3792 gnd.n4439 gnd.n886 585
R3793 gnd.n4444 gnd.n886 585
R3794 gnd.n4438 gnd.n4437 585
R3795 gnd.n4436 gnd.n4435 585
R3796 gnd.n4434 gnd.n4433 585
R3797 gnd.n4432 gnd.n4431 585
R3798 gnd.n4430 gnd.n4429 585
R3799 gnd.n4428 gnd.n4427 585
R3800 gnd.n4426 gnd.n4425 585
R3801 gnd.n4424 gnd.n4423 585
R3802 gnd.n4422 gnd.n4421 585
R3803 gnd.n4420 gnd.n4419 585
R3804 gnd.n4418 gnd.n4417 585
R3805 gnd.n4416 gnd.n4415 585
R3806 gnd.n4414 gnd.n4413 585
R3807 gnd.n4412 gnd.n4411 585
R3808 gnd.n4410 gnd.n4409 585
R3809 gnd.n4407 gnd.n4406 585
R3810 gnd.n4405 gnd.n4404 585
R3811 gnd.n4403 gnd.n4402 585
R3812 gnd.n4401 gnd.n4400 585
R3813 gnd.n4399 gnd.n4398 585
R3814 gnd.n4397 gnd.n4396 585
R3815 gnd.n4395 gnd.n4394 585
R3816 gnd.n4393 gnd.n4392 585
R3817 gnd.n4391 gnd.n4390 585
R3818 gnd.n4389 gnd.n4388 585
R3819 gnd.n4387 gnd.n4386 585
R3820 gnd.n4385 gnd.n4384 585
R3821 gnd.n4383 gnd.n4382 585
R3822 gnd.n4381 gnd.n4380 585
R3823 gnd.n4379 gnd.n4378 585
R3824 gnd.n4377 gnd.n4376 585
R3825 gnd.n4375 gnd.n4374 585
R3826 gnd.n4373 gnd.n4372 585
R3827 gnd.n4371 gnd.n927 585
R3828 gnd.n931 gnd.n928 585
R3829 gnd.n4367 gnd.n4366 585
R3830 gnd.n2112 gnd.n2111 585
R3831 gnd.n2588 gnd.n2587 585
R3832 gnd.n2590 gnd.n2589 585
R3833 gnd.n2592 gnd.n2591 585
R3834 gnd.n2594 gnd.n2593 585
R3835 gnd.n2596 gnd.n2595 585
R3836 gnd.n2598 gnd.n2597 585
R3837 gnd.n2600 gnd.n2599 585
R3838 gnd.n2602 gnd.n2601 585
R3839 gnd.n2604 gnd.n2603 585
R3840 gnd.n2606 gnd.n2605 585
R3841 gnd.n2608 gnd.n2607 585
R3842 gnd.n2610 gnd.n2609 585
R3843 gnd.n2612 gnd.n2611 585
R3844 gnd.n2614 gnd.n2613 585
R3845 gnd.n2616 gnd.n2615 585
R3846 gnd.n2618 gnd.n2617 585
R3847 gnd.n2620 gnd.n2619 585
R3848 gnd.n2622 gnd.n2621 585
R3849 gnd.n2625 gnd.n2624 585
R3850 gnd.n2623 gnd.n2090 585
R3851 gnd.n2760 gnd.n2759 585
R3852 gnd.n2762 gnd.n2761 585
R3853 gnd.n2764 gnd.n2763 585
R3854 gnd.n2766 gnd.n2765 585
R3855 gnd.n2768 gnd.n2767 585
R3856 gnd.n2770 gnd.n2769 585
R3857 gnd.n2772 gnd.n2771 585
R3858 gnd.n2774 gnd.n2773 585
R3859 gnd.n2776 gnd.n2775 585
R3860 gnd.n2778 gnd.n2777 585
R3861 gnd.n2780 gnd.n2779 585
R3862 gnd.n2782 gnd.n2781 585
R3863 gnd.n2783 gnd.n2071 585
R3864 gnd.n2785 gnd.n2784 585
R3865 gnd.n2072 gnd.n2070 585
R3866 gnd.n2073 gnd.n1190 585
R3867 gnd.n2787 gnd.n1190 585
R3868 gnd.n2583 gnd.n1192 585
R3869 gnd.n4206 gnd.n1192 585
R3870 gnd.n2582 gnd.n2581 585
R3871 gnd.n2581 gnd.n2580 585
R3872 gnd.n2116 gnd.n1182 585
R3873 gnd.n4212 gnd.n1182 585
R3874 gnd.n2535 gnd.n2534 585
R3875 gnd.n2536 gnd.n2535 585
R3876 gnd.n2121 gnd.n1171 585
R3877 gnd.n4218 gnd.n1171 585
R3878 gnd.n2529 gnd.n2528 585
R3879 gnd.n2528 gnd.n2527 585
R3880 gnd.n2123 gnd.n1160 585
R3881 gnd.n4224 gnd.n1160 585
R3882 gnd.n2455 gnd.n2127 585
R3883 gnd.n2519 gnd.n2127 585
R3884 gnd.n2456 gnd.n1150 585
R3885 gnd.n4230 gnd.n1150 585
R3886 gnd.n2458 gnd.n2457 585
R3887 gnd.n2459 gnd.n2458 585
R3888 gnd.n2147 gnd.n1139 585
R3889 gnd.n4236 gnd.n1139 585
R3890 gnd.n2449 gnd.n2448 585
R3891 gnd.n2448 gnd.n2447 585
R3892 gnd.n2445 gnd.n1129 585
R3893 gnd.n4242 gnd.n1129 585
R3894 gnd.n2444 gnd.n2443 585
R3895 gnd.n2443 gnd.n2442 585
R3896 gnd.n2149 gnd.n1118 585
R3897 gnd.n4248 gnd.n1118 585
R3898 gnd.n2438 gnd.n2139 585
R3899 gnd.n2473 gnd.n2139 585
R3900 gnd.n2437 gnd.n1108 585
R3901 gnd.n4254 gnd.n1108 585
R3902 gnd.n2436 gnd.n2435 585
R3903 gnd.n2435 gnd.n2434 585
R3904 gnd.n2151 gnd.n1097 585
R3905 gnd.n4260 gnd.n1097 585
R3906 gnd.n2425 gnd.n2424 585
R3907 gnd.n2426 gnd.n2425 585
R3908 gnd.n2184 gnd.n1087 585
R3909 gnd.n4266 gnd.n1087 585
R3910 gnd.n2419 gnd.n2418 585
R3911 gnd.n2418 gnd.n2417 585
R3912 gnd.n2186 gnd.n1077 585
R3913 gnd.n4272 gnd.n1077 585
R3914 gnd.n2253 gnd.n2252 585
R3915 gnd.n2252 gnd.n1069 585
R3916 gnd.n2254 gnd.n1067 585
R3917 gnd.n4278 gnd.n1067 585
R3918 gnd.n2256 gnd.n2255 585
R3919 gnd.n2257 gnd.n2256 585
R3920 gnd.n2190 gnd.n1060 585
R3921 gnd.n4285 gnd.n1060 585
R3922 gnd.n2245 gnd.n2244 585
R3923 gnd.n2244 gnd.n1059 585
R3924 gnd.n2243 gnd.n1050 585
R3925 gnd.n4291 gnd.n1050 585
R3926 gnd.n2242 gnd.n2241 585
R3927 gnd.n2241 gnd.n1044 585
R3928 gnd.n2193 gnd.n1042 585
R3929 gnd.n4297 gnd.n1042 585
R3930 gnd.n2237 gnd.n2236 585
R3931 gnd.n2236 gnd.n1034 585
R3932 gnd.n2235 gnd.n1032 585
R3933 gnd.n4303 gnd.n1032 585
R3934 gnd.n2234 gnd.n2233 585
R3935 gnd.n2233 gnd.n1031 585
R3936 gnd.n2195 gnd.n1022 585
R3937 gnd.n4309 gnd.n1022 585
R3938 gnd.n2229 gnd.n2228 585
R3939 gnd.n2228 gnd.n1021 585
R3940 gnd.n2227 gnd.n1012 585
R3941 gnd.n4315 gnd.n1012 585
R3942 gnd.n2226 gnd.n2225 585
R3943 gnd.n2225 gnd.n1004 585
R3944 gnd.n2197 gnd.n1002 585
R3945 gnd.n4321 gnd.n1002 585
R3946 gnd.n2221 gnd.n2220 585
R3947 gnd.n2220 gnd.n994 585
R3948 gnd.n2219 gnd.n992 585
R3949 gnd.n4327 gnd.n992 585
R3950 gnd.n2218 gnd.n2217 585
R3951 gnd.n2217 gnd.n991 585
R3952 gnd.n2199 gnd.n982 585
R3953 gnd.n4333 gnd.n982 585
R3954 gnd.n2213 gnd.n2212 585
R3955 gnd.n2212 gnd.n981 585
R3956 gnd.n2211 gnd.n972 585
R3957 gnd.n4339 gnd.n972 585
R3958 gnd.n2210 gnd.n2209 585
R3959 gnd.n2209 gnd.n964 585
R3960 gnd.n2201 gnd.n962 585
R3961 gnd.n4345 gnd.n962 585
R3962 gnd.n2205 gnd.n2204 585
R3963 gnd.n2204 gnd.n953 585
R3964 gnd.n2203 gnd.n951 585
R3965 gnd.n4351 gnd.n951 585
R3966 gnd.n938 gnd.n936 585
R3967 gnd.n941 gnd.n938 585
R3968 gnd.n4359 gnd.n4358 585
R3969 gnd.n4358 gnd.n4357 585
R3970 gnd.n937 gnd.n934 585
R3971 gnd.n939 gnd.n937 585
R3972 gnd.n4363 gnd.n933 585
R3973 gnd.n2352 gnd.n933 585
R3974 gnd.n4365 gnd.n4364 585
R3975 gnd.n4365 gnd.n885 585
R3976 gnd.n7013 gnd.n7012 585
R3977 gnd.n7014 gnd.n7013 585
R3978 gnd.n106 gnd.n104 585
R3979 gnd.n104 gnd.n100 585
R3980 gnd.n6933 gnd.n6932 585
R3981 gnd.n6934 gnd.n6933 585
R3982 gnd.n184 gnd.n183 585
R3983 gnd.n183 gnd.n181 585
R3984 gnd.n6928 gnd.n6927 585
R3985 gnd.n6927 gnd.n6926 585
R3986 gnd.n187 gnd.n186 585
R3987 gnd.n188 gnd.n187 585
R3988 gnd.n6842 gnd.n6841 585
R3989 gnd.n6843 gnd.n6842 585
R3990 gnd.n199 gnd.n198 585
R3991 gnd.n6718 gnd.n198 585
R3992 gnd.n6837 gnd.n6836 585
R3993 gnd.n6836 gnd.n6835 585
R3994 gnd.n202 gnd.n201 585
R3995 gnd.n203 gnd.n202 585
R3996 gnd.n6826 gnd.n6825 585
R3997 gnd.n6827 gnd.n6826 585
R3998 gnd.n215 gnd.n214 585
R3999 gnd.n214 gnd.n212 585
R4000 gnd.n6821 gnd.n6820 585
R4001 gnd.n6820 gnd.n6819 585
R4002 gnd.n218 gnd.n217 585
R4003 gnd.n219 gnd.n218 585
R4004 gnd.n6810 gnd.n6809 585
R4005 gnd.n6811 gnd.n6810 585
R4006 gnd.n228 gnd.n227 585
R4007 gnd.n235 gnd.n227 585
R4008 gnd.n6805 gnd.n6804 585
R4009 gnd.n6804 gnd.n6803 585
R4010 gnd.n231 gnd.n230 585
R4011 gnd.n232 gnd.n231 585
R4012 gnd.n6794 gnd.n6793 585
R4013 gnd.n6795 gnd.n6794 585
R4014 gnd.n245 gnd.n244 585
R4015 gnd.n244 gnd.n242 585
R4016 gnd.n6789 gnd.n6788 585
R4017 gnd.n6788 gnd.n6787 585
R4018 gnd.n248 gnd.n247 585
R4019 gnd.n249 gnd.n248 585
R4020 gnd.n6778 gnd.n6777 585
R4021 gnd.n6779 gnd.n6778 585
R4022 gnd.n258 gnd.n257 585
R4023 gnd.n288 gnd.n257 585
R4024 gnd.n6755 gnd.n6754 585
R4025 gnd.n6756 gnd.n6755 585
R4026 gnd.n6753 gnd.n6752 585
R4027 gnd.n6752 gnd.n285 585
R4028 gnd.n6751 gnd.n291 585
R4029 gnd.n6751 gnd.n6750 585
R4030 gnd.n290 gnd.n289 585
R4031 gnd.n292 gnd.n289 585
R4032 gnd.n6678 gnd.n303 585
R4033 gnd.n6678 gnd.n6677 585
R4034 gnd.n6679 gnd.n264 585
R4035 gnd.n6680 gnd.n6679 585
R4036 gnd.n268 gnd.n265 585
R4037 gnd.n300 gnd.n268 585
R4038 gnd.n6774 gnd.n6773 585
R4039 gnd.n6773 gnd.n6772 585
R4040 gnd.n267 gnd.n266 585
R4041 gnd.n333 gnd.n267 585
R4042 gnd.n6659 gnd.n318 585
R4043 gnd.n6643 gnd.n318 585
R4044 gnd.n6661 gnd.n6660 585
R4045 gnd.n6662 gnd.n6661 585
R4046 gnd.n319 gnd.n317 585
R4047 gnd.n4010 gnd.n317 585
R4048 gnd.n6654 gnd.n6653 585
R4049 gnd.n6653 gnd.n6652 585
R4050 gnd.n322 gnd.n321 585
R4051 gnd.n3993 gnd.n322 585
R4052 gnd.n4027 gnd.n4026 585
R4053 gnd.n4028 gnd.n4027 585
R4054 gnd.n1364 gnd.n1363 585
R4055 gnd.n1371 gnd.n1363 585
R4056 gnd.n4022 gnd.n4021 585
R4057 gnd.n4021 gnd.n4020 585
R4058 gnd.n1367 gnd.n1366 585
R4059 gnd.n3958 gnd.n1367 585
R4060 gnd.n3974 gnd.n1402 585
R4061 gnd.n1421 gnd.n1402 585
R4062 gnd.n3976 gnd.n3975 585
R4063 gnd.n3977 gnd.n3976 585
R4064 gnd.n1403 gnd.n1401 585
R4065 gnd.n1410 gnd.n1401 585
R4066 gnd.n3969 gnd.n3968 585
R4067 gnd.n3968 gnd.n3967 585
R4068 gnd.n1406 gnd.n1405 585
R4069 gnd.n3922 gnd.n1406 585
R4070 gnd.n3937 gnd.n3936 585
R4071 gnd.n3938 gnd.n3937 585
R4072 gnd.n1433 gnd.n1432 585
R4073 gnd.n1438 gnd.n1432 585
R4074 gnd.n3932 gnd.n3931 585
R4075 gnd.n3931 gnd.n3930 585
R4076 gnd.n1335 gnd.n1334 585
R4077 gnd.n3897 gnd.n1335 585
R4078 gnd.n4055 gnd.n4054 585
R4079 gnd.n4054 gnd.n4053 585
R4080 gnd.n4056 gnd.n1330 585
R4081 gnd.n3905 gnd.n1330 585
R4082 gnd.n4058 gnd.n4057 585
R4083 gnd.n4059 gnd.n4058 585
R4084 gnd.n3797 gnd.n1329 585
R4085 gnd.n3802 gnd.n3800 585
R4086 gnd.n3803 gnd.n3796 585
R4087 gnd.n3803 gnd.n1316 585
R4088 gnd.n3806 gnd.n3805 585
R4089 gnd.n3794 gnd.n3793 585
R4090 gnd.n3811 gnd.n3810 585
R4091 gnd.n3813 gnd.n3792 585
R4092 gnd.n3816 gnd.n3815 585
R4093 gnd.n3790 gnd.n3789 585
R4094 gnd.n3821 gnd.n3820 585
R4095 gnd.n3823 gnd.n3788 585
R4096 gnd.n3826 gnd.n3825 585
R4097 gnd.n3786 gnd.n3785 585
R4098 gnd.n3832 gnd.n3831 585
R4099 gnd.n3834 gnd.n3784 585
R4100 gnd.n3835 gnd.n1487 585
R4101 gnd.n1485 gnd.n1484 585
R4102 gnd.n3845 gnd.n3844 585
R4103 gnd.n3847 gnd.n1483 585
R4104 gnd.n3850 gnd.n3849 585
R4105 gnd.n1481 gnd.n1480 585
R4106 gnd.n3855 gnd.n3854 585
R4107 gnd.n3857 gnd.n1479 585
R4108 gnd.n3860 gnd.n3859 585
R4109 gnd.n1477 gnd.n1476 585
R4110 gnd.n3865 gnd.n3864 585
R4111 gnd.n3867 gnd.n1475 585
R4112 gnd.n3870 gnd.n3869 585
R4113 gnd.n1473 gnd.n1472 585
R4114 gnd.n3875 gnd.n3874 585
R4115 gnd.n3877 gnd.n1471 585
R4116 gnd.n3880 gnd.n3879 585
R4117 gnd.n1469 gnd.n1468 585
R4118 gnd.n3886 gnd.n3885 585
R4119 gnd.n3888 gnd.n1467 585
R4120 gnd.n3889 gnd.n1466 585
R4121 gnd.n3892 gnd.n3891 585
R4122 gnd.n174 gnd.n173 585
R4123 gnd.n6942 gnd.n169 585
R4124 gnd.n6944 gnd.n6943 585
R4125 gnd.n6946 gnd.n167 585
R4126 gnd.n6948 gnd.n6947 585
R4127 gnd.n6949 gnd.n162 585
R4128 gnd.n6951 gnd.n6950 585
R4129 gnd.n6953 gnd.n160 585
R4130 gnd.n6955 gnd.n6954 585
R4131 gnd.n6956 gnd.n155 585
R4132 gnd.n6958 gnd.n6957 585
R4133 gnd.n6960 gnd.n153 585
R4134 gnd.n6962 gnd.n6961 585
R4135 gnd.n6963 gnd.n148 585
R4136 gnd.n6965 gnd.n6964 585
R4137 gnd.n6967 gnd.n146 585
R4138 gnd.n6969 gnd.n6968 585
R4139 gnd.n6970 gnd.n141 585
R4140 gnd.n6972 gnd.n6971 585
R4141 gnd.n6974 gnd.n139 585
R4142 gnd.n6976 gnd.n6975 585
R4143 gnd.n6980 gnd.n134 585
R4144 gnd.n6982 gnd.n6981 585
R4145 gnd.n6984 gnd.n132 585
R4146 gnd.n6986 gnd.n6985 585
R4147 gnd.n6987 gnd.n127 585
R4148 gnd.n6989 gnd.n6988 585
R4149 gnd.n6991 gnd.n125 585
R4150 gnd.n6993 gnd.n6992 585
R4151 gnd.n6994 gnd.n120 585
R4152 gnd.n6996 gnd.n6995 585
R4153 gnd.n6998 gnd.n118 585
R4154 gnd.n7000 gnd.n6999 585
R4155 gnd.n7001 gnd.n113 585
R4156 gnd.n7003 gnd.n7002 585
R4157 gnd.n7005 gnd.n111 585
R4158 gnd.n7007 gnd.n7006 585
R4159 gnd.n7008 gnd.n109 585
R4160 gnd.n7009 gnd.n105 585
R4161 gnd.n105 gnd.n102 585
R4162 gnd.n6938 gnd.n101 585
R4163 gnd.n7014 gnd.n101 585
R4164 gnd.n6937 gnd.n6936 585
R4165 gnd.n6936 gnd.n100 585
R4166 gnd.n6935 gnd.n178 585
R4167 gnd.n6935 gnd.n6934 585
R4168 gnd.n6712 gnd.n179 585
R4169 gnd.n181 gnd.n179 585
R4170 gnd.n6713 gnd.n189 585
R4171 gnd.n6926 gnd.n189 585
R4172 gnd.n6715 gnd.n6714 585
R4173 gnd.n6714 gnd.n188 585
R4174 gnd.n6716 gnd.n197 585
R4175 gnd.n6843 gnd.n197 585
R4176 gnd.n6720 gnd.n6719 585
R4177 gnd.n6719 gnd.n6718 585
R4178 gnd.n6721 gnd.n204 585
R4179 gnd.n6835 gnd.n204 585
R4180 gnd.n6723 gnd.n6722 585
R4181 gnd.n6722 gnd.n203 585
R4182 gnd.n6724 gnd.n213 585
R4183 gnd.n6827 gnd.n213 585
R4184 gnd.n6726 gnd.n6725 585
R4185 gnd.n6725 gnd.n212 585
R4186 gnd.n6727 gnd.n220 585
R4187 gnd.n6819 gnd.n220 585
R4188 gnd.n6729 gnd.n6728 585
R4189 gnd.n6728 gnd.n219 585
R4190 gnd.n6730 gnd.n226 585
R4191 gnd.n6811 gnd.n226 585
R4192 gnd.n6732 gnd.n6731 585
R4193 gnd.n6731 gnd.n235 585
R4194 gnd.n6733 gnd.n233 585
R4195 gnd.n6803 gnd.n233 585
R4196 gnd.n6735 gnd.n6734 585
R4197 gnd.n6734 gnd.n232 585
R4198 gnd.n6736 gnd.n243 585
R4199 gnd.n6795 gnd.n243 585
R4200 gnd.n6738 gnd.n6737 585
R4201 gnd.n6737 gnd.n242 585
R4202 gnd.n6739 gnd.n250 585
R4203 gnd.n6787 gnd.n250 585
R4204 gnd.n6741 gnd.n6740 585
R4205 gnd.n6740 gnd.n249 585
R4206 gnd.n6742 gnd.n256 585
R4207 gnd.n6779 gnd.n256 585
R4208 gnd.n6744 gnd.n6743 585
R4209 gnd.n6743 gnd.n288 585
R4210 gnd.n6745 gnd.n286 585
R4211 gnd.n6756 gnd.n286 585
R4212 gnd.n6746 gnd.n294 585
R4213 gnd.n294 gnd.n285 585
R4214 gnd.n6748 gnd.n6747 585
R4215 gnd.n6750 gnd.n6748 585
R4216 gnd.n6686 gnd.n293 585
R4217 gnd.n293 gnd.n292 585
R4218 gnd.n299 gnd.n295 585
R4219 gnd.n6677 gnd.n299 585
R4220 gnd.n6682 gnd.n6681 585
R4221 gnd.n6681 gnd.n6680 585
R4222 gnd.n298 gnd.n297 585
R4223 gnd.n300 gnd.n298 585
R4224 gnd.n4003 gnd.n270 585
R4225 gnd.n6772 gnd.n270 585
R4226 gnd.n4005 gnd.n4004 585
R4227 gnd.n4004 gnd.n333 585
R4228 gnd.n4006 gnd.n332 585
R4229 gnd.n6643 gnd.n332 585
R4230 gnd.n4007 gnd.n314 585
R4231 gnd.n6662 gnd.n314 585
R4232 gnd.n4009 gnd.n4008 585
R4233 gnd.n4010 gnd.n4009 585
R4234 gnd.n1386 gnd.n324 585
R4235 gnd.n6652 gnd.n324 585
R4236 gnd.n3995 gnd.n3994 585
R4237 gnd.n3994 gnd.n3993 585
R4238 gnd.n1388 gnd.n1360 585
R4239 gnd.n4028 gnd.n1360 585
R4240 gnd.n3954 gnd.n3953 585
R4241 gnd.n3953 gnd.n1371 585
R4242 gnd.n3955 gnd.n1369 585
R4243 gnd.n4020 gnd.n1369 585
R4244 gnd.n3957 gnd.n3956 585
R4245 gnd.n3958 gnd.n3957 585
R4246 gnd.n1423 gnd.n1422 585
R4247 gnd.n1422 gnd.n1421 585
R4248 gnd.n3947 gnd.n1399 585
R4249 gnd.n3977 gnd.n1399 585
R4250 gnd.n3946 gnd.n3945 585
R4251 gnd.n3945 gnd.n1410 585
R4252 gnd.n3944 gnd.n1408 585
R4253 gnd.n3967 gnd.n1408 585
R4254 gnd.n1429 gnd.n1425 585
R4255 gnd.n3922 gnd.n1429 585
R4256 gnd.n3940 gnd.n3939 585
R4257 gnd.n3939 gnd.n3938 585
R4258 gnd.n1428 gnd.n1427 585
R4259 gnd.n1438 gnd.n1428 585
R4260 gnd.n3896 gnd.n1436 585
R4261 gnd.n3930 gnd.n1436 585
R4262 gnd.n3899 gnd.n3898 585
R4263 gnd.n3898 gnd.n3897 585
R4264 gnd.n1462 gnd.n1337 585
R4265 gnd.n4053 gnd.n1337 585
R4266 gnd.n3904 gnd.n3903 585
R4267 gnd.n3905 gnd.n3904 585
R4268 gnd.n1461 gnd.n1325 585
R4269 gnd.n4059 gnd.n1325 585
R4270 gnd.n3711 gnd.n3710 585
R4271 gnd.n3712 gnd.n3711 585
R4272 gnd.n3625 gnd.n1530 585
R4273 gnd.n1536 gnd.n1530 585
R4274 gnd.n3624 gnd.n3623 585
R4275 gnd.n3623 gnd.n3622 585
R4276 gnd.n1533 gnd.n1532 585
R4277 gnd.n3340 gnd.n1533 585
R4278 gnd.n3328 gnd.n1623 585
R4279 gnd.n1623 gnd.n1618 585
R4280 gnd.n3330 gnd.n3329 585
R4281 gnd.n3331 gnd.n3330 585
R4282 gnd.n3327 gnd.n1622 585
R4283 gnd.n3322 gnd.n1622 585
R4284 gnd.n3326 gnd.n3325 585
R4285 gnd.n3325 gnd.n3324 585
R4286 gnd.n1625 gnd.n1624 585
R4287 gnd.n3309 gnd.n1625 585
R4288 gnd.n3294 gnd.n1649 585
R4289 gnd.n1649 gnd.n1636 585
R4290 gnd.n3296 gnd.n3295 585
R4291 gnd.n3297 gnd.n3296 585
R4292 gnd.n3293 gnd.n1648 585
R4293 gnd.n1648 gnd.n1644 585
R4294 gnd.n3292 gnd.n3291 585
R4295 gnd.n3291 gnd.n3290 585
R4296 gnd.n1651 gnd.n1650 585
R4297 gnd.n3265 gnd.n1651 585
R4298 gnd.n3279 gnd.n3278 585
R4299 gnd.n3280 gnd.n3279 585
R4300 gnd.n3277 gnd.n1661 585
R4301 gnd.n3271 gnd.n1661 585
R4302 gnd.n3276 gnd.n3275 585
R4303 gnd.n3275 gnd.n3274 585
R4304 gnd.n1663 gnd.n1662 585
R4305 gnd.n3252 gnd.n1663 585
R4306 gnd.n3235 gnd.n1678 585
R4307 gnd.n3223 gnd.n1678 585
R4308 gnd.n3237 gnd.n3236 585
R4309 gnd.n3238 gnd.n3237 585
R4310 gnd.n3234 gnd.n1677 585
R4311 gnd.n1684 gnd.n1677 585
R4312 gnd.n3233 gnd.n3232 585
R4313 gnd.n3232 gnd.n3231 585
R4314 gnd.n1680 gnd.n1679 585
R4315 gnd.n3069 gnd.n1680 585
R4316 gnd.n3212 gnd.n3211 585
R4317 gnd.n3213 gnd.n3212 585
R4318 gnd.n3210 gnd.n1694 585
R4319 gnd.n1694 gnd.n1691 585
R4320 gnd.n3209 gnd.n3208 585
R4321 gnd.n3208 gnd.n3207 585
R4322 gnd.n1696 gnd.n1695 585
R4323 gnd.n3077 gnd.n1696 585
R4324 gnd.n3193 gnd.n3192 585
R4325 gnd.n3194 gnd.n3193 585
R4326 gnd.n3191 gnd.n1707 585
R4327 gnd.n3186 gnd.n1707 585
R4328 gnd.n3190 gnd.n3189 585
R4329 gnd.n3189 gnd.n3188 585
R4330 gnd.n1709 gnd.n1708 585
R4331 gnd.n3174 gnd.n1709 585
R4332 gnd.n3160 gnd.n1730 585
R4333 gnd.n1730 gnd.n1719 585
R4334 gnd.n3162 gnd.n3161 585
R4335 gnd.n3163 gnd.n3162 585
R4336 gnd.n3159 gnd.n1729 585
R4337 gnd.n1729 gnd.n1726 585
R4338 gnd.n3158 gnd.n3157 585
R4339 gnd.n3157 gnd.n3156 585
R4340 gnd.n1732 gnd.n1731 585
R4341 gnd.n3091 gnd.n1732 585
R4342 gnd.n3145 gnd.n3144 585
R4343 gnd.n3146 gnd.n3145 585
R4344 gnd.n3143 gnd.n1743 585
R4345 gnd.n1743 gnd.n1740 585
R4346 gnd.n3142 gnd.n3141 585
R4347 gnd.n3141 gnd.n3140 585
R4348 gnd.n1745 gnd.n1744 585
R4349 gnd.n3100 gnd.n1745 585
R4350 gnd.n3128 gnd.n3127 585
R4351 gnd.n3129 gnd.n3128 585
R4352 gnd.n3126 gnd.n1758 585
R4353 gnd.n1758 gnd.n1755 585
R4354 gnd.n3125 gnd.n3124 585
R4355 gnd.n3124 gnd.n3123 585
R4356 gnd.n1760 gnd.n1759 585
R4357 gnd.n3109 gnd.n1760 585
R4358 gnd.n3057 gnd.n1777 585
R4359 gnd.n1777 gnd.n1769 585
R4360 gnd.n3059 gnd.n3058 585
R4361 gnd.n3060 gnd.n3059 585
R4362 gnd.n3056 gnd.n1776 585
R4363 gnd.n1782 gnd.n1776 585
R4364 gnd.n3055 gnd.n3054 585
R4365 gnd.n3054 gnd.n3053 585
R4366 gnd.n1779 gnd.n1778 585
R4367 gnd.n3027 gnd.n1779 585
R4368 gnd.n3041 gnd.n3040 585
R4369 gnd.n3042 gnd.n3041 585
R4370 gnd.n3039 gnd.n1792 585
R4371 gnd.n3033 gnd.n1792 585
R4372 gnd.n3038 gnd.n3037 585
R4373 gnd.n3037 gnd.n3036 585
R4374 gnd.n1794 gnd.n1793 585
R4375 gnd.n3010 gnd.n1794 585
R4376 gnd.n3001 gnd.n1814 585
R4377 gnd.n1814 gnd.n1813 585
R4378 gnd.n3003 gnd.n3002 585
R4379 gnd.n3004 gnd.n3003 585
R4380 gnd.n3000 gnd.n1811 585
R4381 gnd.n2940 gnd.n1811 585
R4382 gnd.n2999 gnd.n2998 585
R4383 gnd.n2998 gnd.n2997 585
R4384 gnd.n1816 gnd.n1815 585
R4385 gnd.n1831 gnd.n1816 585
R4386 gnd.n2971 gnd.n1827 585
R4387 gnd.t121 gnd.n1827 585
R4388 gnd.n2972 gnd.n1838 585
R4389 gnd.n1838 gnd.n1826 585
R4390 gnd.n2974 gnd.n2973 585
R4391 gnd.n2975 gnd.n2974 585
R4392 gnd.n2969 gnd.n1837 585
R4393 gnd.n2968 gnd.n2967 585
R4394 gnd.n1860 gnd.n1859 585
R4395 gnd.n2965 gnd.n1860 585
R4396 gnd.n2697 gnd.n2696 585
R4397 gnd.n2699 gnd.n2698 585
R4398 gnd.n2701 gnd.n2700 585
R4399 gnd.n2703 gnd.n2702 585
R4400 gnd.n2705 gnd.n2704 585
R4401 gnd.n2707 gnd.n2706 585
R4402 gnd.n2709 gnd.n2708 585
R4403 gnd.n2711 gnd.n2710 585
R4404 gnd.n2713 gnd.n2712 585
R4405 gnd.n2715 gnd.n2714 585
R4406 gnd.n2717 gnd.n2716 585
R4407 gnd.n2719 gnd.n2718 585
R4408 gnd.n2721 gnd.n2720 585
R4409 gnd.n2723 gnd.n2722 585
R4410 gnd.n2725 gnd.n2724 585
R4411 gnd.n2727 gnd.n2726 585
R4412 gnd.n2729 gnd.n2728 585
R4413 gnd.n2731 gnd.n2730 585
R4414 gnd.n2733 gnd.n2732 585
R4415 gnd.n2735 gnd.n2734 585
R4416 gnd.n2737 gnd.n2736 585
R4417 gnd.n2739 gnd.n2738 585
R4418 gnd.n2741 gnd.n2740 585
R4419 gnd.n2743 gnd.n2742 585
R4420 gnd.n2745 gnd.n2744 585
R4421 gnd.n2747 gnd.n2746 585
R4422 gnd.n2749 gnd.n2748 585
R4423 gnd.n2751 gnd.n2750 585
R4424 gnd.n2753 gnd.n2752 585
R4425 gnd.n2757 gnd.n2756 585
R4426 gnd.n2755 gnd.n2692 585
R4427 gnd.n2691 gnd.n2690 585
R4428 gnd.n2689 gnd.n2688 585
R4429 gnd.n2686 gnd.n2685 585
R4430 gnd.n2684 gnd.n2683 585
R4431 gnd.n2682 gnd.n2681 585
R4432 gnd.n2680 gnd.n2679 585
R4433 gnd.n2678 gnd.n2677 585
R4434 gnd.n2676 gnd.n2675 585
R4435 gnd.n2674 gnd.n2673 585
R4436 gnd.n2672 gnd.n2671 585
R4437 gnd.n2670 gnd.n2669 585
R4438 gnd.n2668 gnd.n2667 585
R4439 gnd.n2666 gnd.n2665 585
R4440 gnd.n2664 gnd.n2663 585
R4441 gnd.n2662 gnd.n2661 585
R4442 gnd.n2660 gnd.n2659 585
R4443 gnd.n2658 gnd.n2657 585
R4444 gnd.n2656 gnd.n2655 585
R4445 gnd.n2654 gnd.n2653 585
R4446 gnd.n2652 gnd.n2651 585
R4447 gnd.n2650 gnd.n2649 585
R4448 gnd.n2648 gnd.n2647 585
R4449 gnd.n2646 gnd.n2645 585
R4450 gnd.n2644 gnd.n2643 585
R4451 gnd.n2642 gnd.n2641 585
R4452 gnd.n2640 gnd.n2639 585
R4453 gnd.n2638 gnd.n2637 585
R4454 gnd.n2636 gnd.n2635 585
R4455 gnd.n2634 gnd.n2633 585
R4456 gnd.n2632 gnd.n2631 585
R4457 gnd.n1834 gnd.n1833 585
R4458 gnd.n3715 gnd.n3714 585
R4459 gnd.n3717 gnd.n3716 585
R4460 gnd.n3719 gnd.n3718 585
R4461 gnd.n3721 gnd.n3720 585
R4462 gnd.n3723 gnd.n3722 585
R4463 gnd.n3725 gnd.n3724 585
R4464 gnd.n3727 gnd.n3726 585
R4465 gnd.n3729 gnd.n3728 585
R4466 gnd.n3731 gnd.n3730 585
R4467 gnd.n3733 gnd.n3732 585
R4468 gnd.n3735 gnd.n3734 585
R4469 gnd.n3737 gnd.n3736 585
R4470 gnd.n3739 gnd.n3738 585
R4471 gnd.n3741 gnd.n3740 585
R4472 gnd.n3743 gnd.n3742 585
R4473 gnd.n3745 gnd.n3744 585
R4474 gnd.n3747 gnd.n3746 585
R4475 gnd.n3749 gnd.n3748 585
R4476 gnd.n3751 gnd.n3750 585
R4477 gnd.n3753 gnd.n3752 585
R4478 gnd.n3755 gnd.n3754 585
R4479 gnd.n3757 gnd.n3756 585
R4480 gnd.n3759 gnd.n3758 585
R4481 gnd.n3761 gnd.n3760 585
R4482 gnd.n3763 gnd.n3762 585
R4483 gnd.n3765 gnd.n3764 585
R4484 gnd.n3767 gnd.n3766 585
R4485 gnd.n3769 gnd.n3768 585
R4486 gnd.n3771 gnd.n3770 585
R4487 gnd.n3773 gnd.n1524 585
R4488 gnd.n3775 gnd.n3774 585
R4489 gnd.n3777 gnd.n1488 585
R4490 gnd.n3779 gnd.n3778 585
R4491 gnd.n3782 gnd.n3781 585
R4492 gnd.n1491 gnd.n1489 585
R4493 gnd.n3648 gnd.n3647 585
R4494 gnd.n3650 gnd.n3649 585
R4495 gnd.n3653 gnd.n3652 585
R4496 gnd.n3655 gnd.n3654 585
R4497 gnd.n3657 gnd.n3656 585
R4498 gnd.n3659 gnd.n3658 585
R4499 gnd.n3661 gnd.n3660 585
R4500 gnd.n3663 gnd.n3662 585
R4501 gnd.n3665 gnd.n3664 585
R4502 gnd.n3667 gnd.n3666 585
R4503 gnd.n3669 gnd.n3668 585
R4504 gnd.n3671 gnd.n3670 585
R4505 gnd.n3673 gnd.n3672 585
R4506 gnd.n3675 gnd.n3674 585
R4507 gnd.n3677 gnd.n3676 585
R4508 gnd.n3679 gnd.n3678 585
R4509 gnd.n3681 gnd.n3680 585
R4510 gnd.n3683 gnd.n3682 585
R4511 gnd.n3685 gnd.n3684 585
R4512 gnd.n3687 gnd.n3686 585
R4513 gnd.n3689 gnd.n3688 585
R4514 gnd.n3691 gnd.n3690 585
R4515 gnd.n3693 gnd.n3692 585
R4516 gnd.n3695 gnd.n3694 585
R4517 gnd.n3697 gnd.n3696 585
R4518 gnd.n3699 gnd.n3698 585
R4519 gnd.n3701 gnd.n3700 585
R4520 gnd.n3703 gnd.n3702 585
R4521 gnd.n3705 gnd.n3704 585
R4522 gnd.n3707 gnd.n3706 585
R4523 gnd.n3708 gnd.n1531 585
R4524 gnd.n3713 gnd.n1527 585
R4525 gnd.n3713 gnd.n3712 585
R4526 gnd.n3335 gnd.n1528 585
R4527 gnd.n1536 gnd.n1528 585
R4528 gnd.n3336 gnd.n1535 585
R4529 gnd.n3622 gnd.n1535 585
R4530 gnd.n3338 gnd.n3337 585
R4531 gnd.n3340 gnd.n3338 585
R4532 gnd.n3334 gnd.n1619 585
R4533 gnd.n1619 gnd.n1618 585
R4534 gnd.n3333 gnd.n3332 585
R4535 gnd.n3332 gnd.n3331 585
R4536 gnd.n1621 gnd.n1620 585
R4537 gnd.n3322 gnd.n1621 585
R4538 gnd.n3256 gnd.n1627 585
R4539 gnd.n3324 gnd.n1627 585
R4540 gnd.n3257 gnd.n1637 585
R4541 gnd.n3309 gnd.n1637 585
R4542 gnd.n3259 gnd.n3258 585
R4543 gnd.n3258 gnd.n1636 585
R4544 gnd.n3260 gnd.n1645 585
R4545 gnd.n3297 gnd.n1645 585
R4546 gnd.n3262 gnd.n3261 585
R4547 gnd.n3261 gnd.n1644 585
R4548 gnd.n3263 gnd.n1653 585
R4549 gnd.n3290 gnd.n1653 585
R4550 gnd.n3267 gnd.n3266 585
R4551 gnd.n3266 gnd.n3265 585
R4552 gnd.n3268 gnd.n1659 585
R4553 gnd.n3280 gnd.n1659 585
R4554 gnd.n3270 gnd.n3269 585
R4555 gnd.n3271 gnd.n3270 585
R4556 gnd.n3255 gnd.n1665 585
R4557 gnd.n3274 gnd.n1665 585
R4558 gnd.n3254 gnd.n3253 585
R4559 gnd.n3253 gnd.n3252 585
R4560 gnd.n1668 gnd.n1667 585
R4561 gnd.n3223 gnd.n1668 585
R4562 gnd.n3064 gnd.n1675 585
R4563 gnd.n3238 gnd.n1675 585
R4564 gnd.n3066 gnd.n3065 585
R4565 gnd.n3065 gnd.n1684 585
R4566 gnd.n3067 gnd.n1683 585
R4567 gnd.n3231 gnd.n1683 585
R4568 gnd.n3071 gnd.n3070 585
R4569 gnd.n3070 gnd.n3069 585
R4570 gnd.n3072 gnd.n1692 585
R4571 gnd.n3213 gnd.n1692 585
R4572 gnd.n3074 gnd.n3073 585
R4573 gnd.n3073 gnd.n1691 585
R4574 gnd.n3075 gnd.n1698 585
R4575 gnd.n3207 gnd.n1698 585
R4576 gnd.n3079 gnd.n3078 585
R4577 gnd.n3078 gnd.n3077 585
R4578 gnd.n3080 gnd.n1706 585
R4579 gnd.n3194 gnd.n1706 585
R4580 gnd.n3081 gnd.n1712 585
R4581 gnd.n3186 gnd.n1712 585
R4582 gnd.n3082 gnd.n1711 585
R4583 gnd.n3188 gnd.n1711 585
R4584 gnd.n3083 gnd.n1720 585
R4585 gnd.n3174 gnd.n1720 585
R4586 gnd.n3085 gnd.n3084 585
R4587 gnd.n3084 gnd.n1719 585
R4588 gnd.n3086 gnd.n1727 585
R4589 gnd.n3163 gnd.n1727 585
R4590 gnd.n3088 gnd.n3087 585
R4591 gnd.n3087 gnd.n1726 585
R4592 gnd.n3089 gnd.n1734 585
R4593 gnd.n3156 gnd.n1734 585
R4594 gnd.n3093 gnd.n3092 585
R4595 gnd.n3092 gnd.n3091 585
R4596 gnd.n3094 gnd.n1741 585
R4597 gnd.n3146 gnd.n1741 585
R4598 gnd.n3096 gnd.n3095 585
R4599 gnd.n3095 gnd.n1740 585
R4600 gnd.n3097 gnd.n1747 585
R4601 gnd.n3140 gnd.n1747 585
R4602 gnd.n3102 gnd.n3101 585
R4603 gnd.n3101 gnd.n3100 585
R4604 gnd.n3103 gnd.n1756 585
R4605 gnd.n3129 gnd.n1756 585
R4606 gnd.n3105 gnd.n3104 585
R4607 gnd.n3104 gnd.n1755 585
R4608 gnd.n3106 gnd.n1762 585
R4609 gnd.n3123 gnd.n1762 585
R4610 gnd.n3108 gnd.n3107 585
R4611 gnd.n3109 gnd.n3108 585
R4612 gnd.n3063 gnd.n1771 585
R4613 gnd.n1771 gnd.n1769 585
R4614 gnd.n3062 gnd.n3061 585
R4615 gnd.n3061 gnd.n3060 585
R4616 gnd.n1773 gnd.n1772 585
R4617 gnd.n1782 gnd.n1773 585
R4618 gnd.n1799 gnd.n1780 585
R4619 gnd.n3053 gnd.n1780 585
R4620 gnd.n3029 gnd.n3028 585
R4621 gnd.n3028 gnd.n3027 585
R4622 gnd.n3030 gnd.n1790 585
R4623 gnd.n3042 gnd.n1790 585
R4624 gnd.n3032 gnd.n3031 585
R4625 gnd.n3033 gnd.n3032 585
R4626 gnd.n1798 gnd.n1796 585
R4627 gnd.n3036 gnd.n1796 585
R4628 gnd.n3009 gnd.n3008 585
R4629 gnd.n3010 gnd.n3009 585
R4630 gnd.n3007 gnd.n1807 585
R4631 gnd.n1813 gnd.n1807 585
R4632 gnd.n3006 gnd.n3005 585
R4633 gnd.n3005 gnd.n3004 585
R4634 gnd.n1809 gnd.n1808 585
R4635 gnd.n2940 gnd.n1809 585
R4636 gnd.n2979 gnd.n1819 585
R4637 gnd.n2997 gnd.n1819 585
R4638 gnd.n2980 gnd.n1832 585
R4639 gnd.n1832 gnd.n1831 585
R4640 gnd.n2982 gnd.n2981 585
R4641 gnd.t121 gnd.n2982 585
R4642 gnd.n2978 gnd.n1829 585
R4643 gnd.n1829 gnd.n1826 585
R4644 gnd.n2977 gnd.n2976 585
R4645 gnd.n2976 gnd.n2975 585
R4646 gnd.n844 gnd.n843 585
R4647 gnd.n1066 gnd.n844 585
R4648 gnd.n6633 gnd.n6632 585
R4649 gnd.n6633 gnd.n302 585
R4650 gnd.n6636 gnd.n6635 585
R4651 gnd.n6635 gnd.n6634 585
R4652 gnd.n6639 gnd.n335 585
R4653 gnd.n335 gnd.n269 585
R4654 gnd.n6641 gnd.n6640 585
R4655 gnd.n6642 gnd.n6641 585
R4656 gnd.n336 gnd.n334 585
R4657 gnd.n334 gnd.n315 585
R4658 gnd.n1384 gnd.n1379 585
R4659 gnd.n1379 gnd.n313 585
R4660 gnd.n4012 gnd.n1385 585
R4661 gnd.n4012 gnd.n4011 585
R4662 gnd.n4013 gnd.n1378 585
R4663 gnd.n4013 gnd.n323 585
R4664 gnd.n4015 gnd.n4014 585
R4665 gnd.n4014 gnd.n1362 585
R4666 gnd.n4016 gnd.n1373 585
R4667 gnd.n1373 gnd.n1359 585
R4668 gnd.n4018 gnd.n4017 585
R4669 gnd.n4019 gnd.n4018 585
R4670 gnd.n1374 gnd.n1372 585
R4671 gnd.n1372 gnd.n1368 585
R4672 gnd.n3960 gnd.n1419 585
R4673 gnd.n3960 gnd.n3959 585
R4674 gnd.n3962 gnd.n3961 585
R4675 gnd.n3961 gnd.n1400 585
R4676 gnd.n3963 gnd.n1412 585
R4677 gnd.n1412 gnd.n1398 585
R4678 gnd.n3965 gnd.n3964 585
R4679 gnd.n3966 gnd.n3965 585
R4680 gnd.n1413 gnd.n1411 585
R4681 gnd.n1411 gnd.n1407 585
R4682 gnd.n3925 gnd.n3924 585
R4683 gnd.n3924 gnd.n3923 585
R4684 gnd.n3926 gnd.n1440 585
R4685 gnd.n1440 gnd.n1430 585
R4686 gnd.n3928 gnd.n3927 585
R4687 gnd.n3929 gnd.n3928 585
R4688 gnd.n1441 gnd.n1439 585
R4689 gnd.n1439 gnd.n1435 585
R4690 gnd.n1447 gnd.n1446 585
R4691 gnd.n1446 gnd.n1339 585
R4692 gnd.n1445 gnd.n1444 585
R4693 gnd.n1445 gnd.n1336 585
R4694 gnd.n1323 gnd.n1322 585
R4695 gnd.n1327 gnd.n1323 585
R4696 gnd.n4062 gnd.n4061 585
R4697 gnd.n4061 gnd.n4060 585
R4698 gnd.n4063 gnd.n1317 585
R4699 gnd.n1324 gnd.n1317 585
R4700 gnd.n4065 gnd.n4064 585
R4701 gnd.n4066 gnd.n4065 585
R4702 gnd.n1314 gnd.n1313 585
R4703 gnd.n4067 gnd.n1314 585
R4704 gnd.n4070 gnd.n4069 585
R4705 gnd.n4069 gnd.n4068 585
R4706 gnd.n4071 gnd.n1308 585
R4707 gnd.n1308 gnd.n1306 585
R4708 gnd.n4073 gnd.n4072 585
R4709 gnd.n4074 gnd.n4073 585
R4710 gnd.n1309 gnd.n1307 585
R4711 gnd.n1307 gnd.n1304 585
R4712 gnd.n1596 gnd.n1595 585
R4713 gnd.n3572 gnd.n1596 585
R4714 gnd.n3576 gnd.n3575 585
R4715 gnd.n3575 gnd.n3574 585
R4716 gnd.n3577 gnd.n1588 585
R4717 gnd.n1597 gnd.n1588 585
R4718 gnd.n3579 gnd.n3578 585
R4719 gnd.n3580 gnd.n3579 585
R4720 gnd.n1581 gnd.n1580 585
R4721 gnd.n3582 gnd.n1581 585
R4722 gnd.n3586 gnd.n3585 585
R4723 gnd.n3585 gnd.n3584 585
R4724 gnd.n3587 gnd.n1575 585
R4725 gnd.n1582 gnd.n1575 585
R4726 gnd.n3589 gnd.n3588 585
R4727 gnd.n3590 gnd.n3589 585
R4728 gnd.n1571 gnd.n1570 585
R4729 gnd.n3592 gnd.n1571 585
R4730 gnd.n3596 gnd.n3595 585
R4731 gnd.n3595 gnd.n3594 585
R4732 gnd.n3597 gnd.n1565 585
R4733 gnd.n3369 gnd.n1565 585
R4734 gnd.n3599 gnd.n3598 585
R4735 gnd.n3600 gnd.n3599 585
R4736 gnd.n1558 gnd.n1557 585
R4737 gnd.n3602 gnd.n1558 585
R4738 gnd.n3606 gnd.n3605 585
R4739 gnd.n3605 gnd.n3604 585
R4740 gnd.n3607 gnd.n1550 585
R4741 gnd.n1559 gnd.n1550 585
R4742 gnd.n3609 gnd.n3608 585
R4743 gnd.n3610 gnd.n3609 585
R4744 gnd.n1551 gnd.n1544 585
R4745 gnd.n3612 gnd.n1544 585
R4746 gnd.n3615 gnd.n1543 585
R4747 gnd.n3615 gnd.n3614 585
R4748 gnd.n3617 gnd.n3616 585
R4749 gnd.n3616 gnd.n1492 585
R4750 gnd.n3618 gnd.n1538 585
R4751 gnd.n1538 gnd.n1529 585
R4752 gnd.n3620 gnd.n3619 585
R4753 gnd.n3621 gnd.n3620 585
R4754 gnd.n1539 gnd.n1537 585
R4755 gnd.n3339 gnd.n1537 585
R4756 gnd.n3318 gnd.n1631 585
R4757 gnd.n1631 gnd.n1630 585
R4758 gnd.n3320 gnd.n3319 585
R4759 gnd.n3321 gnd.n3320 585
R4760 gnd.n1632 gnd.n1629 585
R4761 gnd.n1629 gnd.n1626 585
R4762 gnd.n3312 gnd.n3311 585
R4763 gnd.n3311 gnd.n3310 585
R4764 gnd.n1635 gnd.n1634 585
R4765 gnd.n3298 gnd.n1635 585
R4766 gnd.n3288 gnd.n3287 585
R4767 gnd.n3289 gnd.n3288 585
R4768 gnd.n1655 gnd.n1654 585
R4769 gnd.n3264 gnd.n1654 585
R4770 gnd.n3283 gnd.n3282 585
R4771 gnd.n3282 gnd.n3281 585
R4772 gnd.n1658 gnd.n1657 585
R4773 gnd.n1664 gnd.n1658 585
R4774 gnd.n3226 gnd.n3225 585
R4775 gnd.n3225 gnd.n3224 585
R4776 gnd.n3227 gnd.n1686 585
R4777 gnd.n1686 gnd.n1676 585
R4778 gnd.n3229 gnd.n3228 585
R4779 gnd.n3230 gnd.n3229 585
R4780 gnd.n1687 gnd.n1685 585
R4781 gnd.n3068 gnd.n1685 585
R4782 gnd.n3216 gnd.n3215 585
R4783 gnd.n3215 gnd.n3214 585
R4784 gnd.n1690 gnd.n1689 585
R4785 gnd.n3206 gnd.n1690 585
R4786 gnd.n3182 gnd.n1714 585
R4787 gnd.n3076 gnd.n1714 585
R4788 gnd.n3184 gnd.n3183 585
R4789 gnd.n3185 gnd.n3184 585
R4790 gnd.n1715 gnd.n1713 585
R4791 gnd.n1713 gnd.n1710 585
R4792 gnd.n3177 gnd.n3176 585
R4793 gnd.n3176 gnd.n3175 585
R4794 gnd.n1718 gnd.n1717 585
R4795 gnd.n3164 gnd.n1718 585
R4796 gnd.n3154 gnd.n3153 585
R4797 gnd.n3155 gnd.n3154 585
R4798 gnd.n1736 gnd.n1735 585
R4799 gnd.n3090 gnd.n1735 585
R4800 gnd.n3149 gnd.n3148 585
R4801 gnd.n3148 gnd.n3147 585
R4802 gnd.n1739 gnd.n1738 585
R4803 gnd.n1746 gnd.n1739 585
R4804 gnd.n3118 gnd.n1764 585
R4805 gnd.n1764 gnd.n1757 585
R4806 gnd.n3120 gnd.n3119 585
R4807 gnd.n3121 gnd.n3120 585
R4808 gnd.n1765 gnd.n1763 585
R4809 gnd.n1763 gnd.n1761 585
R4810 gnd.n3113 gnd.n3112 585
R4811 gnd.n3112 gnd.n3111 585
R4812 gnd.n1768 gnd.n1767 585
R4813 gnd.n1781 gnd.n1768 585
R4814 gnd.n3051 gnd.n3050 585
R4815 gnd.n3052 gnd.n3051 585
R4816 gnd.n1785 gnd.n1784 585
R4817 gnd.n1791 gnd.n1784 585
R4818 gnd.n3046 gnd.n3045 585
R4819 gnd.n3045 gnd.n3044 585
R4820 gnd.n1788 gnd.n1787 585
R4821 gnd.n1795 gnd.n1788 585
R4822 gnd.n2992 gnd.n2991 585
R4823 gnd.n2991 gnd.n1806 585
R4824 gnd.n2993 gnd.n1821 585
R4825 gnd.n1821 gnd.n1810 585
R4826 gnd.n2995 gnd.n2994 585
R4827 gnd.n2996 gnd.n2995 585
R4828 gnd.n1822 gnd.n1820 585
R4829 gnd.n1830 gnd.n1820 585
R4830 gnd.n2985 gnd.n2984 585
R4831 gnd.n2984 gnd.n2983 585
R4832 gnd.n1825 gnd.n1824 585
R4833 gnd.n1835 gnd.n1825 585
R4834 gnd.n2963 gnd.n2962 585
R4835 gnd.n2964 gnd.n2963 585
R4836 gnd.n1897 gnd.n1896 585
R4837 gnd.n2954 gnd.n1896 585
R4838 gnd.n2958 gnd.n2957 585
R4839 gnd.n2957 gnd.n2956 585
R4840 gnd.n1900 gnd.n1899 585
R4841 gnd.n2927 gnd.n1900 585
R4842 gnd.n2925 gnd.n2924 585
R4843 gnd.n2926 gnd.n2925 585
R4844 gnd.n1912 gnd.n1911 585
R4845 gnd.n2916 gnd.n1911 585
R4846 gnd.n2920 gnd.n2919 585
R4847 gnd.n2919 gnd.n2918 585
R4848 gnd.n1915 gnd.n1914 585
R4849 gnd.n2907 gnd.n1915 585
R4850 gnd.n2905 gnd.n2904 585
R4851 gnd.n2906 gnd.n2905 585
R4852 gnd.n1925 gnd.n1924 585
R4853 gnd.n2896 gnd.n1924 585
R4854 gnd.n2900 gnd.n2899 585
R4855 gnd.n2899 gnd.n2898 585
R4856 gnd.n1928 gnd.n1927 585
R4857 gnd.n2887 gnd.n1928 585
R4858 gnd.n2885 gnd.n2884 585
R4859 gnd.n2886 gnd.n2885 585
R4860 gnd.n1938 gnd.n1937 585
R4861 gnd.n2876 gnd.n1937 585
R4862 gnd.n2880 gnd.n2879 585
R4863 gnd.n2879 gnd.n2878 585
R4864 gnd.n1941 gnd.n1940 585
R4865 gnd.n2867 gnd.n1941 585
R4866 gnd.n2865 gnd.n2864 585
R4867 gnd.n2866 gnd.n2865 585
R4868 gnd.n1951 gnd.n1950 585
R4869 gnd.n2856 gnd.n1950 585
R4870 gnd.n2860 gnd.n2859 585
R4871 gnd.n2859 gnd.n2858 585
R4872 gnd.n1954 gnd.n1953 585
R4873 gnd.n2847 gnd.n1954 585
R4874 gnd.n2845 gnd.n2844 585
R4875 gnd.n2846 gnd.n2845 585
R4876 gnd.n1962 gnd.n1961 585
R4877 gnd.n1961 gnd.n1960 585
R4878 gnd.n2840 gnd.n2839 585
R4879 gnd.n2839 gnd.n2838 585
R4880 gnd.n1965 gnd.n1964 585
R4881 gnd.n1966 gnd.n1965 585
R4882 gnd.n2503 gnd.n2499 585
R4883 gnd.n2499 gnd.n2051 585
R4884 gnd.n2505 gnd.n2504 585
R4885 gnd.n2505 gnd.n2035 585
R4886 gnd.n2506 gnd.n2498 585
R4887 gnd.n2506 gnd.n1194 585
R4888 gnd.n2508 gnd.n2507 585
R4889 gnd.n2507 gnd.n1191 585
R4890 gnd.n2509 gnd.n2493 585
R4891 gnd.n2493 gnd.n1184 585
R4892 gnd.n2511 gnd.n2510 585
R4893 gnd.n2511 gnd.n1181 585
R4894 gnd.n2512 gnd.n2492 585
R4895 gnd.n2512 gnd.n1173 585
R4896 gnd.n2514 gnd.n2513 585
R4897 gnd.n2513 gnd.n1170 585
R4898 gnd.n2515 gnd.n2129 585
R4899 gnd.n2129 gnd.n1162 585
R4900 gnd.n2517 gnd.n2516 585
R4901 gnd.n2518 gnd.n2517 585
R4902 gnd.n2130 gnd.n2128 585
R4903 gnd.n2128 gnd.n1152 585
R4904 gnd.n2486 gnd.n2485 585
R4905 gnd.n2485 gnd.n1149 585
R4906 gnd.n2484 gnd.n2132 585
R4907 gnd.n2484 gnd.n1141 585
R4908 gnd.n2483 gnd.n2482 585
R4909 gnd.n2483 gnd.n1138 585
R4910 gnd.n2134 gnd.n2133 585
R4911 gnd.n2446 gnd.n2133 585
R4912 gnd.n2478 gnd.n2477 585
R4913 gnd.n2477 gnd.n1128 585
R4914 gnd.n2476 gnd.n2136 585
R4915 gnd.n2476 gnd.n1120 585
R4916 gnd.n2475 gnd.n2138 585
R4917 gnd.n2475 gnd.n2474 585
R4918 gnd.n2175 gnd.n2137 585
R4919 gnd.n2137 gnd.n1110 585
R4920 gnd.n2177 gnd.n2176 585
R4921 gnd.n2177 gnd.n1107 585
R4922 gnd.n2179 gnd.n2178 585
R4923 gnd.n2178 gnd.n1099 585
R4924 gnd.n2180 gnd.n2157 585
R4925 gnd.n2157 gnd.n1096 585
R4926 gnd.n2182 gnd.n2181 585
R4927 gnd.n2183 gnd.n2182 585
R4928 gnd.n2158 gnd.n2156 585
R4929 gnd.n2156 gnd.n1086 585
R4930 gnd.n2166 gnd.n2165 585
R4931 gnd.n2165 gnd.n1079 585
R4932 gnd.n2164 gnd.n2162 585
R4933 gnd.n2164 gnd.n2163 585
R4934 gnd.n4077 gnd.n4076 585
R4935 gnd.n4076 gnd.n4075 585
R4936 gnd.n4078 gnd.n1301 585
R4937 gnd.n3571 gnd.n1301 585
R4938 gnd.n4079 gnd.n1300 585
R4939 gnd.n3573 gnd.n1300 585
R4940 gnd.n1598 gnd.n1298 585
R4941 gnd.n1599 gnd.n1598 585
R4942 gnd.n4083 gnd.n1297 585
R4943 gnd.n1587 gnd.n1297 585
R4944 gnd.n4084 gnd.n1296 585
R4945 gnd.n3581 gnd.n1296 585
R4946 gnd.n4085 gnd.n1295 585
R4947 gnd.n3583 gnd.n1295 585
R4948 gnd.n1583 gnd.n1293 585
R4949 gnd.n1584 gnd.n1583 585
R4950 gnd.n4089 gnd.n1292 585
R4951 gnd.n1574 gnd.n1292 585
R4952 gnd.n4090 gnd.n1291 585
R4953 gnd.n3591 gnd.n1291 585
R4954 gnd.n4091 gnd.n1290 585
R4955 gnd.n3593 gnd.n1290 585
R4956 gnd.n3370 gnd.n1288 585
R4957 gnd.n3371 gnd.n3370 585
R4958 gnd.n4095 gnd.n1287 585
R4959 gnd.n1564 gnd.n1287 585
R4960 gnd.n4096 gnd.n1286 585
R4961 gnd.n3601 gnd.n1286 585
R4962 gnd.n4097 gnd.n1285 585
R4963 gnd.n3603 gnd.n1285 585
R4964 gnd.n1560 gnd.n1283 585
R4965 gnd.n1561 gnd.n1560 585
R4966 gnd.n4101 gnd.n1282 585
R4967 gnd.n1549 gnd.n1282 585
R4968 gnd.n4102 gnd.n1281 585
R4969 gnd.n3611 gnd.n1281 585
R4970 gnd.n4103 gnd.n1280 585
R4971 gnd.n3613 gnd.n1280 585
R4972 gnd.n1545 gnd.n1278 585
R4973 gnd.n1546 gnd.n1545 585
R4974 gnd.n4107 gnd.n1277 585
R4975 gnd.n3351 gnd.n1277 585
R4976 gnd.n4108 gnd.n1276 585
R4977 gnd.n3349 gnd.n1276 585
R4978 gnd.n4109 gnd.n1275 585
R4979 gnd.n1534 gnd.n1275 585
R4980 gnd.n3341 gnd.n1273 585
R4981 gnd.n3342 gnd.n3341 585
R4982 gnd.n4113 gnd.n1272 585
R4983 gnd.n3331 gnd.n1272 585
R4984 gnd.n4114 gnd.n1271 585
R4985 gnd.n3323 gnd.n1271 585
R4986 gnd.n4115 gnd.n1270 585
R4987 gnd.n3308 gnd.n1270 585
R4988 gnd.n1646 gnd.n1268 585
R4989 gnd.n1647 gnd.n1646 585
R4990 gnd.n4119 gnd.n1267 585
R4991 gnd.n3299 gnd.n1267 585
R4992 gnd.n4120 gnd.n1266 585
R4993 gnd.n1652 gnd.n1266 585
R4994 gnd.n4121 gnd.n1265 585
R4995 gnd.n1660 gnd.n1265 585
R4996 gnd.n3272 gnd.n1263 585
R4997 gnd.n3273 gnd.n3272 585
R4998 gnd.n4125 gnd.n1262 585
R4999 gnd.n3251 gnd.n1262 585
R5000 gnd.n4126 gnd.n1261 585
R5001 gnd.n3222 gnd.n1261 585
R5002 gnd.n4127 gnd.n1260 585
R5003 gnd.n3239 gnd.n1260 585
R5004 gnd.n1681 gnd.n1258 585
R5005 gnd.n1682 gnd.n1681 585
R5006 gnd.n4131 gnd.n1257 585
R5007 gnd.n1693 gnd.n1257 585
R5008 gnd.n4132 gnd.n1256 585
R5009 gnd.n3205 gnd.n1256 585
R5010 gnd.n4133 gnd.n1255 585
R5011 gnd.n1697 gnd.n1255 585
R5012 gnd.n3195 gnd.n1253 585
R5013 gnd.n3196 gnd.n3195 585
R5014 gnd.n4137 gnd.n1252 585
R5015 gnd.n3187 gnd.n1252 585
R5016 gnd.n4138 gnd.n1251 585
R5017 gnd.n3174 gnd.n1251 585
R5018 gnd.n4139 gnd.n1250 585
R5019 gnd.n1728 gnd.n1250 585
R5020 gnd.n3165 gnd.n1248 585
R5021 gnd.n3166 gnd.n3165 585
R5022 gnd.n4143 gnd.n1247 585
R5023 gnd.n1733 gnd.n1247 585
R5024 gnd.n4144 gnd.n1246 585
R5025 gnd.n1742 gnd.n1246 585
R5026 gnd.n4145 gnd.n1245 585
R5027 gnd.n3139 gnd.n1245 585
R5028 gnd.n3098 gnd.n1243 585
R5029 gnd.n3099 gnd.n3098 585
R5030 gnd.n4149 gnd.n1242 585
R5031 gnd.n3130 gnd.n1242 585
R5032 gnd.n4150 gnd.n1241 585
R5033 gnd.n3122 gnd.n1241 585
R5034 gnd.n4151 gnd.n1240 585
R5035 gnd.n3110 gnd.n1240 585
R5036 gnd.n1774 gnd.n1238 585
R5037 gnd.n1775 gnd.n1774 585
R5038 gnd.n4155 gnd.n1237 585
R5039 gnd.n1783 gnd.n1237 585
R5040 gnd.n4156 gnd.n1236 585
R5041 gnd.n3026 gnd.n1236 585
R5042 gnd.n4157 gnd.n1235 585
R5043 gnd.n3043 gnd.n1235 585
R5044 gnd.n3034 gnd.n1233 585
R5045 gnd.n3035 gnd.n3034 585
R5046 gnd.n4161 gnd.n1232 585
R5047 gnd.n3011 gnd.n1232 585
R5048 gnd.n4162 gnd.n1231 585
R5049 gnd.n1812 gnd.n1231 585
R5050 gnd.n4163 gnd.n1230 585
R5051 gnd.n2940 gnd.n1230 585
R5052 gnd.n1817 gnd.n1228 585
R5053 gnd.n1818 gnd.n1817 585
R5054 gnd.n4167 gnd.n1227 585
R5055 gnd.n1828 gnd.n1227 585
R5056 gnd.n4168 gnd.n1226 585
R5057 gnd.n1836 gnd.n1226 585
R5058 gnd.n4169 gnd.n1225 585
R5059 gnd.n1895 gnd.n1225 585
R5060 gnd.n1861 gnd.n1223 585
R5061 gnd.n1862 gnd.n1861 585
R5062 gnd.n4173 gnd.n1222 585
R5063 gnd.n2955 gnd.n1222 585
R5064 gnd.n4174 gnd.n1221 585
R5065 gnd.n1901 gnd.n1221 585
R5066 gnd.n4175 gnd.n1220 585
R5067 gnd.n2928 gnd.n1220 585
R5068 gnd.n1909 gnd.n1218 585
R5069 gnd.n1910 gnd.n1909 585
R5070 gnd.n4179 gnd.n1217 585
R5071 gnd.n2917 gnd.n1217 585
R5072 gnd.n4180 gnd.n1216 585
R5073 gnd.n1916 gnd.n1216 585
R5074 gnd.n4181 gnd.n1215 585
R5075 gnd.n2908 gnd.n1215 585
R5076 gnd.n1922 gnd.n1213 585
R5077 gnd.n1923 gnd.n1922 585
R5078 gnd.n4185 gnd.n1212 585
R5079 gnd.n2897 gnd.n1212 585
R5080 gnd.n4186 gnd.n1211 585
R5081 gnd.n1929 gnd.n1211 585
R5082 gnd.n4187 gnd.n1210 585
R5083 gnd.n2888 gnd.n1210 585
R5084 gnd.n1935 gnd.n1208 585
R5085 gnd.n1936 gnd.n1935 585
R5086 gnd.n4191 gnd.n1207 585
R5087 gnd.n2877 gnd.n1207 585
R5088 gnd.n4192 gnd.n1206 585
R5089 gnd.n1942 gnd.n1206 585
R5090 gnd.n4193 gnd.n1205 585
R5091 gnd.n2868 gnd.n1205 585
R5092 gnd.n1948 gnd.n1203 585
R5093 gnd.n1949 gnd.n1948 585
R5094 gnd.n4197 gnd.n1202 585
R5095 gnd.n2857 gnd.n1202 585
R5096 gnd.n4198 gnd.n1201 585
R5097 gnd.n1955 gnd.n1201 585
R5098 gnd.n4199 gnd.n1200 585
R5099 gnd.n2848 gnd.n1200 585
R5100 gnd.n2835 gnd.n2834 585
R5101 gnd.n2833 gnd.n1981 585
R5102 gnd.n1983 gnd.n1980 585
R5103 gnd.n2837 gnd.n1980 585
R5104 gnd.n2826 gnd.n1991 585
R5105 gnd.n2825 gnd.n1992 585
R5106 gnd.n1994 gnd.n1993 585
R5107 gnd.n2818 gnd.n2000 585
R5108 gnd.n2817 gnd.n2001 585
R5109 gnd.n2008 gnd.n2002 585
R5110 gnd.n2810 gnd.n2009 585
R5111 gnd.n2809 gnd.n2010 585
R5112 gnd.n2012 gnd.n2011 585
R5113 gnd.n2802 gnd.n2018 585
R5114 gnd.n2801 gnd.n2019 585
R5115 gnd.n2028 gnd.n2020 585
R5116 gnd.n2794 gnd.n2029 585
R5117 gnd.n2793 gnd.n2030 585
R5118 gnd.n2032 gnd.n2031 585
R5119 gnd.n2573 gnd.n2542 585
R5120 gnd.n2572 gnd.n2543 585
R5121 gnd.n2571 gnd.n2544 585
R5122 gnd.n2546 gnd.n2545 585
R5123 gnd.n2567 gnd.n2548 585
R5124 gnd.n2566 gnd.n2549 585
R5125 gnd.n2565 gnd.n2550 585
R5126 gnd.n2562 gnd.n2555 585
R5127 gnd.n2561 gnd.n2556 585
R5128 gnd.n2560 gnd.n2557 585
R5129 gnd.n2558 gnd.n1959 585
R5130 gnd.n1602 gnd.n1305 585
R5131 gnd.n4075 gnd.n1305 585
R5132 gnd.n3570 gnd.n3569 585
R5133 gnd.n3571 gnd.n3570 585
R5134 gnd.n1601 gnd.n1600 585
R5135 gnd.n3573 gnd.n1600 585
R5136 gnd.n3389 gnd.n3388 585
R5137 gnd.n3388 gnd.n1599 585
R5138 gnd.n3387 gnd.n3386 585
R5139 gnd.n3387 gnd.n1587 585
R5140 gnd.n3385 gnd.n1586 585
R5141 gnd.n3581 gnd.n1586 585
R5142 gnd.n1604 gnd.n1585 585
R5143 gnd.n3583 gnd.n1585 585
R5144 gnd.n3381 gnd.n3380 585
R5145 gnd.n3380 gnd.n1584 585
R5146 gnd.n3379 gnd.n3378 585
R5147 gnd.n3379 gnd.n1574 585
R5148 gnd.n3377 gnd.n1573 585
R5149 gnd.n3591 gnd.n1573 585
R5150 gnd.n1606 gnd.n1572 585
R5151 gnd.n3593 gnd.n1572 585
R5152 gnd.n3373 gnd.n3372 585
R5153 gnd.n3372 gnd.n3371 585
R5154 gnd.n3368 gnd.n3367 585
R5155 gnd.n3368 gnd.n1564 585
R5156 gnd.n3366 gnd.n1563 585
R5157 gnd.n3601 gnd.n1563 585
R5158 gnd.n1608 gnd.n1562 585
R5159 gnd.n3603 gnd.n1562 585
R5160 gnd.n3362 gnd.n3361 585
R5161 gnd.n3361 gnd.n1561 585
R5162 gnd.n3360 gnd.n3359 585
R5163 gnd.n3360 gnd.n1549 585
R5164 gnd.n3358 gnd.n1548 585
R5165 gnd.n3611 gnd.n1548 585
R5166 gnd.n1610 gnd.n1547 585
R5167 gnd.n3613 gnd.n1547 585
R5168 gnd.n3354 gnd.n3353 585
R5169 gnd.n3353 gnd.n1546 585
R5170 gnd.n3352 gnd.n1612 585
R5171 gnd.n3352 gnd.n3351 585
R5172 gnd.n3350 gnd.n3348 585
R5173 gnd.n3350 gnd.n3349 585
R5174 gnd.n1614 gnd.n1613 585
R5175 gnd.n1613 gnd.n1534 585
R5176 gnd.n3344 gnd.n3343 585
R5177 gnd.n3343 gnd.n3342 585
R5178 gnd.n1617 gnd.n1616 585
R5179 gnd.n3331 gnd.n1617 585
R5180 gnd.n1640 gnd.n1628 585
R5181 gnd.n3323 gnd.n1628 585
R5182 gnd.n3307 gnd.n3306 585
R5183 gnd.n3308 gnd.n3307 585
R5184 gnd.n1639 gnd.n1638 585
R5185 gnd.n1647 gnd.n1638 585
R5186 gnd.n3301 gnd.n3300 585
R5187 gnd.n3300 gnd.n3299 585
R5188 gnd.n1643 gnd.n1642 585
R5189 gnd.n1652 gnd.n1643 585
R5190 gnd.n3245 gnd.n3244 585
R5191 gnd.n3244 gnd.n1660 585
R5192 gnd.n1671 gnd.n1666 585
R5193 gnd.n3273 gnd.n1666 585
R5194 gnd.n3250 gnd.n3249 585
R5195 gnd.n3251 gnd.n3250 585
R5196 gnd.n1670 gnd.n1669 585
R5197 gnd.n3222 gnd.n1669 585
R5198 gnd.n3241 gnd.n3240 585
R5199 gnd.n3240 gnd.n3239 585
R5200 gnd.n1674 gnd.n1673 585
R5201 gnd.n1682 gnd.n1674 585
R5202 gnd.n1702 gnd.n1700 585
R5203 gnd.n1700 gnd.n1693 585
R5204 gnd.n3204 gnd.n3203 585
R5205 gnd.n3205 gnd.n3204 585
R5206 gnd.n1701 gnd.n1699 585
R5207 gnd.n1699 gnd.n1697 585
R5208 gnd.n3198 gnd.n3197 585
R5209 gnd.n3197 gnd.n3196 585
R5210 gnd.n1705 gnd.n1704 585
R5211 gnd.n3187 gnd.n1705 585
R5212 gnd.n3173 gnd.n3172 585
R5213 gnd.n3174 gnd.n3173 585
R5214 gnd.n1722 gnd.n1721 585
R5215 gnd.n1728 gnd.n1721 585
R5216 gnd.n3168 gnd.n3167 585
R5217 gnd.n3167 gnd.n3166 585
R5218 gnd.n1725 gnd.n1724 585
R5219 gnd.n1733 gnd.n1725 585
R5220 gnd.n1751 gnd.n1749 585
R5221 gnd.n1749 gnd.n1742 585
R5222 gnd.n3138 gnd.n3137 585
R5223 gnd.n3139 gnd.n3138 585
R5224 gnd.n1750 gnd.n1748 585
R5225 gnd.n3099 gnd.n1748 585
R5226 gnd.n3132 gnd.n3131 585
R5227 gnd.n3131 gnd.n3130 585
R5228 gnd.n1754 gnd.n1753 585
R5229 gnd.n3122 gnd.n1754 585
R5230 gnd.n3019 gnd.n1770 585
R5231 gnd.n3110 gnd.n1770 585
R5232 gnd.n3020 gnd.n3018 585
R5233 gnd.n3018 gnd.n1775 585
R5234 gnd.n1802 gnd.n1800 585
R5235 gnd.n1800 gnd.n1783 585
R5236 gnd.n3025 gnd.n3024 585
R5237 gnd.n3026 gnd.n3025 585
R5238 gnd.n1801 gnd.n1789 585
R5239 gnd.n3043 gnd.n1789 585
R5240 gnd.n3014 gnd.n1797 585
R5241 gnd.n3035 gnd.n1797 585
R5242 gnd.n3013 gnd.n3012 585
R5243 gnd.n3012 gnd.n3011 585
R5244 gnd.n1805 gnd.n1804 585
R5245 gnd.n1812 gnd.n1805 585
R5246 gnd.n2942 gnd.n2941 585
R5247 gnd.n2941 gnd.n2940 585
R5248 gnd.n2939 gnd.n2937 585
R5249 gnd.n2939 gnd.n1818 585
R5250 gnd.n2946 gnd.n2936 585
R5251 gnd.n2936 gnd.n1828 585
R5252 gnd.n2947 gnd.n2935 585
R5253 gnd.n2935 gnd.n1836 585
R5254 gnd.n2948 gnd.n2934 585
R5255 gnd.n2934 gnd.n1895 585
R5256 gnd.n1905 gnd.n1903 585
R5257 gnd.n1903 gnd.n1862 585
R5258 gnd.n2953 gnd.n2952 585
R5259 gnd.n2955 gnd.n2953 585
R5260 gnd.n1904 gnd.n1902 585
R5261 gnd.n1902 gnd.n1901 585
R5262 gnd.n2930 gnd.n2929 585
R5263 gnd.n2929 gnd.n2928 585
R5264 gnd.n1908 gnd.n1907 585
R5265 gnd.n1910 gnd.n1908 585
R5266 gnd.n2915 gnd.n2914 585
R5267 gnd.n2917 gnd.n2915 585
R5268 gnd.n1918 gnd.n1917 585
R5269 gnd.n1917 gnd.n1916 585
R5270 gnd.n2910 gnd.n2909 585
R5271 gnd.n2909 gnd.n2908 585
R5272 gnd.n1921 gnd.n1920 585
R5273 gnd.n1923 gnd.n1921 585
R5274 gnd.n2895 gnd.n2894 585
R5275 gnd.n2897 gnd.n2895 585
R5276 gnd.n1931 gnd.n1930 585
R5277 gnd.n1930 gnd.n1929 585
R5278 gnd.n2890 gnd.n2889 585
R5279 gnd.n2889 gnd.n2888 585
R5280 gnd.n1934 gnd.n1933 585
R5281 gnd.n1936 gnd.n1934 585
R5282 gnd.n2875 gnd.n2874 585
R5283 gnd.n2877 gnd.n2875 585
R5284 gnd.n1944 gnd.n1943 585
R5285 gnd.n1943 gnd.n1942 585
R5286 gnd.n2870 gnd.n2869 585
R5287 gnd.n2869 gnd.n2868 585
R5288 gnd.n1947 gnd.n1946 585
R5289 gnd.n1949 gnd.n1947 585
R5290 gnd.n2855 gnd.n2854 585
R5291 gnd.n2857 gnd.n2855 585
R5292 gnd.n1957 gnd.n1956 585
R5293 gnd.n1956 gnd.n1955 585
R5294 gnd.n2850 gnd.n2849 585
R5295 gnd.n2849 gnd.n2848 585
R5296 gnd.n3565 gnd.n3564 585
R5297 gnd.n3564 gnd.n1315 585
R5298 gnd.n3563 gnd.n3393 585
R5299 gnd.n3561 gnd.n3560 585
R5300 gnd.n3395 gnd.n3394 585
R5301 gnd.n3556 gnd.n3552 585
R5302 gnd.n3550 gnd.n3397 585
R5303 gnd.n3548 gnd.n3547 585
R5304 gnd.n3399 gnd.n3398 585
R5305 gnd.n3543 gnd.n3542 585
R5306 gnd.n3540 gnd.n3401 585
R5307 gnd.n3538 gnd.n3537 585
R5308 gnd.n3403 gnd.n3402 585
R5309 gnd.n3523 gnd.n3522 585
R5310 gnd.n3524 gnd.n3520 585
R5311 gnd.n3518 gnd.n3412 585
R5312 gnd.n3517 gnd.n3516 585
R5313 gnd.n3501 gnd.n3414 585
R5314 gnd.n3503 gnd.n3502 585
R5315 gnd.n3499 gnd.n3421 585
R5316 gnd.n3498 gnd.n3497 585
R5317 gnd.n3482 gnd.n3423 585
R5318 gnd.n3484 gnd.n3483 585
R5319 gnd.n3480 gnd.n3430 585
R5320 gnd.n3479 gnd.n3478 585
R5321 gnd.n3463 gnd.n3432 585
R5322 gnd.n3465 gnd.n3464 585
R5323 gnd.n3461 gnd.n3439 585
R5324 gnd.n3460 gnd.n3459 585
R5325 gnd.n3441 gnd.n1303 585
R5326 gnd.n2629 gnd.t44 543.808
R5327 gnd.n1525 gnd.t47 543.808
R5328 gnd.n2693 gnd.t94 543.808
R5329 gnd.n3645 gnd.t97 543.808
R5330 gnd.n3711 gnd.n1531 497.305
R5331 gnd.n3714 gnd.n3713 497.305
R5332 gnd.n2976 gnd.n1834 497.305
R5333 gnd.n2974 gnd.n1837 497.305
R5334 gnd.n6064 gnd.n6063 392.846
R5335 gnd.n2551 gnd.t113 371.625
R5336 gnd.n6884 gnd.t51 371.625
R5337 gnd.n3405 gnd.t73 371.625
R5338 gnd.n2024 gnd.t106 371.625
R5339 gnd.n3838 gnd.t70 371.625
R5340 gnd.n1464 gnd.t55 371.625
R5341 gnd.n175 gnd.t142 371.625
R5342 gnd.n6977 gnd.t59 371.625
R5343 gnd.n907 gnd.t139 371.625
R5344 gnd.n929 gnd.t127 371.625
R5345 gnd.n2113 gnd.t62 371.625
R5346 gnd.n2091 gnd.t91 371.625
R5347 gnd.n2294 gnd.t80 371.625
R5348 gnd.n3553 gnd.t84 371.625
R5349 gnd.n5400 gnd.t66 323.425
R5350 gnd.n4474 gnd.t109 323.425
R5351 gnd.n4785 gnd.n4759 289.615
R5352 gnd.n4753 gnd.n4727 289.615
R5353 gnd.n4721 gnd.n4695 289.615
R5354 gnd.n4690 gnd.n4664 289.615
R5355 gnd.n4658 gnd.n4632 289.615
R5356 gnd.n4626 gnd.n4600 289.615
R5357 gnd.n4594 gnd.n4568 289.615
R5358 gnd.n4563 gnd.n4537 289.615
R5359 gnd.n5137 gnd.t76 279.217
R5360 gnd.n4518 gnd.t123 279.217
R5361 gnd.n1845 gnd.t135 260.649
R5362 gnd.n3637 gnd.t105 260.649
R5363 gnd.n2966 gnd.n2965 256.663
R5364 gnd.n2965 gnd.n1863 256.663
R5365 gnd.n2965 gnd.n1864 256.663
R5366 gnd.n2965 gnd.n1865 256.663
R5367 gnd.n2965 gnd.n1866 256.663
R5368 gnd.n2965 gnd.n1867 256.663
R5369 gnd.n2965 gnd.n1868 256.663
R5370 gnd.n2965 gnd.n1869 256.663
R5371 gnd.n2965 gnd.n1870 256.663
R5372 gnd.n2965 gnd.n1871 256.663
R5373 gnd.n2965 gnd.n1872 256.663
R5374 gnd.n2965 gnd.n1873 256.663
R5375 gnd.n2965 gnd.n1874 256.663
R5376 gnd.n2965 gnd.n1875 256.663
R5377 gnd.n2965 gnd.n1876 256.663
R5378 gnd.n2965 gnd.n1877 256.663
R5379 gnd.n2757 gnd.n2754 256.663
R5380 gnd.n2965 gnd.n1878 256.663
R5381 gnd.n2965 gnd.n1879 256.663
R5382 gnd.n2965 gnd.n1880 256.663
R5383 gnd.n2965 gnd.n1881 256.663
R5384 gnd.n2965 gnd.n1882 256.663
R5385 gnd.n2965 gnd.n1883 256.663
R5386 gnd.n2965 gnd.n1884 256.663
R5387 gnd.n2965 gnd.n1885 256.663
R5388 gnd.n2965 gnd.n1886 256.663
R5389 gnd.n2965 gnd.n1887 256.663
R5390 gnd.n2965 gnd.n1888 256.663
R5391 gnd.n2965 gnd.n1889 256.663
R5392 gnd.n2965 gnd.n1890 256.663
R5393 gnd.n2965 gnd.n1891 256.663
R5394 gnd.n2965 gnd.n1892 256.663
R5395 gnd.n2965 gnd.n1893 256.663
R5396 gnd.n2965 gnd.n1894 256.663
R5397 gnd.n3779 gnd.n1509 256.663
R5398 gnd.n3779 gnd.n1510 256.663
R5399 gnd.n3779 gnd.n1511 256.663
R5400 gnd.n3779 gnd.n1512 256.663
R5401 gnd.n3779 gnd.n1513 256.663
R5402 gnd.n3779 gnd.n1514 256.663
R5403 gnd.n3779 gnd.n1515 256.663
R5404 gnd.n3779 gnd.n1516 256.663
R5405 gnd.n3779 gnd.n1517 256.663
R5406 gnd.n3779 gnd.n1518 256.663
R5407 gnd.n3779 gnd.n1519 256.663
R5408 gnd.n3779 gnd.n1520 256.663
R5409 gnd.n3779 gnd.n1521 256.663
R5410 gnd.n3779 gnd.n1522 256.663
R5411 gnd.n3779 gnd.n1523 256.663
R5412 gnd.n3779 gnd.n3776 256.663
R5413 gnd.n3782 gnd.n1490 256.663
R5414 gnd.n3780 gnd.n3779 256.663
R5415 gnd.n3779 gnd.n1508 256.663
R5416 gnd.n3779 gnd.n1507 256.663
R5417 gnd.n3779 gnd.n1506 256.663
R5418 gnd.n3779 gnd.n1505 256.663
R5419 gnd.n3779 gnd.n1504 256.663
R5420 gnd.n3779 gnd.n1503 256.663
R5421 gnd.n3779 gnd.n1502 256.663
R5422 gnd.n3779 gnd.n1501 256.663
R5423 gnd.n3779 gnd.n1500 256.663
R5424 gnd.n3779 gnd.n1499 256.663
R5425 gnd.n3779 gnd.n1498 256.663
R5426 gnd.n3779 gnd.n1497 256.663
R5427 gnd.n3779 gnd.n1496 256.663
R5428 gnd.n3779 gnd.n1495 256.663
R5429 gnd.n3779 gnd.n1494 256.663
R5430 gnd.n3779 gnd.n1493 256.663
R5431 gnd.n4444 gnd.n875 242.672
R5432 gnd.n4444 gnd.n876 242.672
R5433 gnd.n4444 gnd.n877 242.672
R5434 gnd.n4444 gnd.n878 242.672
R5435 gnd.n4444 gnd.n879 242.672
R5436 gnd.n4444 gnd.n880 242.672
R5437 gnd.n4444 gnd.n881 242.672
R5438 gnd.n4444 gnd.n882 242.672
R5439 gnd.n4444 gnd.n883 242.672
R5440 gnd.n2788 gnd.n2787 242.672
R5441 gnd.n2787 gnd.n2050 242.672
R5442 gnd.n2787 gnd.n2049 242.672
R5443 gnd.n2787 gnd.n2047 242.672
R5444 gnd.n2787 gnd.n2045 242.672
R5445 gnd.n2787 gnd.n2044 242.672
R5446 gnd.n2787 gnd.n2042 242.672
R5447 gnd.n2787 gnd.n2040 242.672
R5448 gnd.n2787 gnd.n2039 242.672
R5449 gnd.n3451 gnd.n1316 242.672
R5450 gnd.n3453 gnd.n1316 242.672
R5451 gnd.n3470 gnd.n1316 242.672
R5452 gnd.n3472 gnd.n1316 242.672
R5453 gnd.n3489 gnd.n1316 242.672
R5454 gnd.n3491 gnd.n1316 242.672
R5455 gnd.n3508 gnd.n1316 242.672
R5456 gnd.n3510 gnd.n1316 242.672
R5457 gnd.n3529 gnd.n1316 242.672
R5458 gnd.n6886 gnd.n102 242.672
R5459 gnd.n6882 gnd.n102 242.672
R5460 gnd.n6877 gnd.n102 242.672
R5461 gnd.n6874 gnd.n102 242.672
R5462 gnd.n6869 gnd.n102 242.672
R5463 gnd.n6866 gnd.n102 242.672
R5464 gnd.n6861 gnd.n102 242.672
R5465 gnd.n6858 gnd.n102 242.672
R5466 gnd.n6853 gnd.n102 242.672
R5467 gnd.n5192 gnd.n5101 242.672
R5468 gnd.n5105 gnd.n5101 242.672
R5469 gnd.n5185 gnd.n5101 242.672
R5470 gnd.n5179 gnd.n5101 242.672
R5471 gnd.n5177 gnd.n5101 242.672
R5472 gnd.n5171 gnd.n5101 242.672
R5473 gnd.n5169 gnd.n5101 242.672
R5474 gnd.n5163 gnd.n5101 242.672
R5475 gnd.n5161 gnd.n5101 242.672
R5476 gnd.n5155 gnd.n5101 242.672
R5477 gnd.n5153 gnd.n5101 242.672
R5478 gnd.n5146 gnd.n5101 242.672
R5479 gnd.n5144 gnd.n5101 242.672
R5480 gnd.n5804 gnd.n4445 242.672
R5481 gnd.n5810 gnd.n4445 242.672
R5482 gnd.n4521 gnd.n4445 242.672
R5483 gnd.n5817 gnd.n4445 242.672
R5484 gnd.n4512 gnd.n4445 242.672
R5485 gnd.n5824 gnd.n4445 242.672
R5486 gnd.n4505 gnd.n4445 242.672
R5487 gnd.n5831 gnd.n4445 242.672
R5488 gnd.n4498 gnd.n4445 242.672
R5489 gnd.n5838 gnd.n4445 242.672
R5490 gnd.n4491 gnd.n4445 242.672
R5491 gnd.n5845 gnd.n4445 242.672
R5492 gnd.n4484 gnd.n4445 242.672
R5493 gnd.n5434 gnd.n5433 242.672
R5494 gnd.n5434 gnd.n5375 242.672
R5495 gnd.n5434 gnd.n5376 242.672
R5496 gnd.n5434 gnd.n5377 242.672
R5497 gnd.n5434 gnd.n5378 242.672
R5498 gnd.n5434 gnd.n5379 242.672
R5499 gnd.n5434 gnd.n5380 242.672
R5500 gnd.n5434 gnd.n5381 242.672
R5501 gnd.n5856 gnd.n4445 242.672
R5502 gnd.n4477 gnd.n4445 242.672
R5503 gnd.n5863 gnd.n4445 242.672
R5504 gnd.n4468 gnd.n4445 242.672
R5505 gnd.n5870 gnd.n4445 242.672
R5506 gnd.n4461 gnd.n4445 242.672
R5507 gnd.n5877 gnd.n4445 242.672
R5508 gnd.n4454 gnd.n4445 242.672
R5509 gnd.n4444 gnd.n4443 242.672
R5510 gnd.n4444 gnd.n857 242.672
R5511 gnd.n4444 gnd.n858 242.672
R5512 gnd.n4444 gnd.n859 242.672
R5513 gnd.n4444 gnd.n860 242.672
R5514 gnd.n4444 gnd.n861 242.672
R5515 gnd.n4444 gnd.n862 242.672
R5516 gnd.n4444 gnd.n863 242.672
R5517 gnd.n4444 gnd.n864 242.672
R5518 gnd.n4444 gnd.n865 242.672
R5519 gnd.n4444 gnd.n866 242.672
R5520 gnd.n4444 gnd.n867 242.672
R5521 gnd.n4444 gnd.n868 242.672
R5522 gnd.n4444 gnd.n869 242.672
R5523 gnd.n4444 gnd.n870 242.672
R5524 gnd.n4444 gnd.n871 242.672
R5525 gnd.n4444 gnd.n872 242.672
R5526 gnd.n4444 gnd.n873 242.672
R5527 gnd.n4444 gnd.n874 242.672
R5528 gnd.n2787 gnd.n2052 242.672
R5529 gnd.n2787 gnd.n2053 242.672
R5530 gnd.n2787 gnd.n2054 242.672
R5531 gnd.n2787 gnd.n2055 242.672
R5532 gnd.n2787 gnd.n2056 242.672
R5533 gnd.n2787 gnd.n2057 242.672
R5534 gnd.n2787 gnd.n2058 242.672
R5535 gnd.n2787 gnd.n2059 242.672
R5536 gnd.n2787 gnd.n2060 242.672
R5537 gnd.n2787 gnd.n2061 242.672
R5538 gnd.n2787 gnd.n2062 242.672
R5539 gnd.n2758 gnd.n2093 242.672
R5540 gnd.n2787 gnd.n2063 242.672
R5541 gnd.n2787 gnd.n2064 242.672
R5542 gnd.n2787 gnd.n2065 242.672
R5543 gnd.n2787 gnd.n2066 242.672
R5544 gnd.n2787 gnd.n2067 242.672
R5545 gnd.n2787 gnd.n2068 242.672
R5546 gnd.n2787 gnd.n2069 242.672
R5547 gnd.n2787 gnd.n2786 242.672
R5548 gnd.n3801 gnd.n1316 242.672
R5549 gnd.n3804 gnd.n1316 242.672
R5550 gnd.n3812 gnd.n1316 242.672
R5551 gnd.n3814 gnd.n1316 242.672
R5552 gnd.n3822 gnd.n1316 242.672
R5553 gnd.n3824 gnd.n1316 242.672
R5554 gnd.n3833 gnd.n1316 242.672
R5555 gnd.n3836 gnd.n1316 242.672
R5556 gnd.n3840 gnd.n3837 242.672
R5557 gnd.n3783 gnd.n1316 242.672
R5558 gnd.n3846 gnd.n1316 242.672
R5559 gnd.n3848 gnd.n1316 242.672
R5560 gnd.n3856 gnd.n1316 242.672
R5561 gnd.n3858 gnd.n1316 242.672
R5562 gnd.n3866 gnd.n1316 242.672
R5563 gnd.n3868 gnd.n1316 242.672
R5564 gnd.n3876 gnd.n1316 242.672
R5565 gnd.n3878 gnd.n1316 242.672
R5566 gnd.n3887 gnd.n1316 242.672
R5567 gnd.n3890 gnd.n1316 242.672
R5568 gnd.n172 gnd.n102 242.672
R5569 gnd.n6945 gnd.n102 242.672
R5570 gnd.n168 gnd.n102 242.672
R5571 gnd.n6952 gnd.n102 242.672
R5572 gnd.n161 gnd.n102 242.672
R5573 gnd.n6959 gnd.n102 242.672
R5574 gnd.n154 gnd.n102 242.672
R5575 gnd.n6966 gnd.n102 242.672
R5576 gnd.n147 gnd.n102 242.672
R5577 gnd.n6973 gnd.n102 242.672
R5578 gnd.n140 gnd.n102 242.672
R5579 gnd.n6983 gnd.n102 242.672
R5580 gnd.n133 gnd.n102 242.672
R5581 gnd.n6990 gnd.n102 242.672
R5582 gnd.n126 gnd.n102 242.672
R5583 gnd.n6997 gnd.n102 242.672
R5584 gnd.n119 gnd.n102 242.672
R5585 gnd.n7004 gnd.n102 242.672
R5586 gnd.n112 gnd.n102 242.672
R5587 gnd.n2837 gnd.n2836 242.672
R5588 gnd.n2837 gnd.n1967 242.672
R5589 gnd.n2837 gnd.n1968 242.672
R5590 gnd.n2837 gnd.n1969 242.672
R5591 gnd.n2837 gnd.n1970 242.672
R5592 gnd.n2837 gnd.n1971 242.672
R5593 gnd.n2837 gnd.n1972 242.672
R5594 gnd.n2837 gnd.n1973 242.672
R5595 gnd.n2837 gnd.n1974 242.672
R5596 gnd.n2837 gnd.n1975 242.672
R5597 gnd.n2837 gnd.n1976 242.672
R5598 gnd.n2837 gnd.n1977 242.672
R5599 gnd.n2837 gnd.n1978 242.672
R5600 gnd.n2837 gnd.n1979 242.672
R5601 gnd.n3562 gnd.n1315 242.672
R5602 gnd.n3551 gnd.n1315 242.672
R5603 gnd.n3549 gnd.n1315 242.672
R5604 gnd.n3541 gnd.n1315 242.672
R5605 gnd.n3539 gnd.n1315 242.672
R5606 gnd.n3521 gnd.n1315 242.672
R5607 gnd.n3519 gnd.n1315 242.672
R5608 gnd.n3413 gnd.n1315 242.672
R5609 gnd.n3500 gnd.n1315 242.672
R5610 gnd.n3422 gnd.n1315 242.672
R5611 gnd.n3481 gnd.n1315 242.672
R5612 gnd.n3431 gnd.n1315 242.672
R5613 gnd.n3462 gnd.n1315 242.672
R5614 gnd.n3440 gnd.n1315 242.672
R5615 gnd.n109 gnd.n105 240.244
R5616 gnd.n7006 gnd.n7005 240.244
R5617 gnd.n7003 gnd.n113 240.244
R5618 gnd.n6999 gnd.n6998 240.244
R5619 gnd.n6996 gnd.n120 240.244
R5620 gnd.n6992 gnd.n6991 240.244
R5621 gnd.n6989 gnd.n127 240.244
R5622 gnd.n6985 gnd.n6984 240.244
R5623 gnd.n6982 gnd.n134 240.244
R5624 gnd.n6975 gnd.n6974 240.244
R5625 gnd.n6972 gnd.n141 240.244
R5626 gnd.n6968 gnd.n6967 240.244
R5627 gnd.n6965 gnd.n148 240.244
R5628 gnd.n6961 gnd.n6960 240.244
R5629 gnd.n6958 gnd.n155 240.244
R5630 gnd.n6954 gnd.n6953 240.244
R5631 gnd.n6951 gnd.n162 240.244
R5632 gnd.n6947 gnd.n6946 240.244
R5633 gnd.n6944 gnd.n169 240.244
R5634 gnd.n3904 gnd.n1325 240.244
R5635 gnd.n3904 gnd.n1337 240.244
R5636 gnd.n3898 gnd.n1337 240.244
R5637 gnd.n3898 gnd.n1436 240.244
R5638 gnd.n1436 gnd.n1428 240.244
R5639 gnd.n3939 gnd.n1428 240.244
R5640 gnd.n3939 gnd.n1429 240.244
R5641 gnd.n1429 gnd.n1408 240.244
R5642 gnd.n3945 gnd.n1408 240.244
R5643 gnd.n3945 gnd.n1399 240.244
R5644 gnd.n1422 gnd.n1399 240.244
R5645 gnd.n3957 gnd.n1422 240.244
R5646 gnd.n3957 gnd.n1369 240.244
R5647 gnd.n3953 gnd.n1369 240.244
R5648 gnd.n3953 gnd.n1360 240.244
R5649 gnd.n3994 gnd.n1360 240.244
R5650 gnd.n3994 gnd.n324 240.244
R5651 gnd.n4009 gnd.n324 240.244
R5652 gnd.n4009 gnd.n314 240.244
R5653 gnd.n332 gnd.n314 240.244
R5654 gnd.n4004 gnd.n332 240.244
R5655 gnd.n4004 gnd.n270 240.244
R5656 gnd.n298 gnd.n270 240.244
R5657 gnd.n6681 gnd.n298 240.244
R5658 gnd.n6681 gnd.n299 240.244
R5659 gnd.n299 gnd.n293 240.244
R5660 gnd.n6748 gnd.n293 240.244
R5661 gnd.n6748 gnd.n294 240.244
R5662 gnd.n294 gnd.n286 240.244
R5663 gnd.n6743 gnd.n286 240.244
R5664 gnd.n6743 gnd.n256 240.244
R5665 gnd.n6740 gnd.n256 240.244
R5666 gnd.n6740 gnd.n250 240.244
R5667 gnd.n6737 gnd.n250 240.244
R5668 gnd.n6737 gnd.n243 240.244
R5669 gnd.n6734 gnd.n243 240.244
R5670 gnd.n6734 gnd.n233 240.244
R5671 gnd.n6731 gnd.n233 240.244
R5672 gnd.n6731 gnd.n226 240.244
R5673 gnd.n6728 gnd.n226 240.244
R5674 gnd.n6728 gnd.n220 240.244
R5675 gnd.n6725 gnd.n220 240.244
R5676 gnd.n6725 gnd.n213 240.244
R5677 gnd.n6722 gnd.n213 240.244
R5678 gnd.n6722 gnd.n204 240.244
R5679 gnd.n6719 gnd.n204 240.244
R5680 gnd.n6719 gnd.n197 240.244
R5681 gnd.n6714 gnd.n197 240.244
R5682 gnd.n6714 gnd.n189 240.244
R5683 gnd.n189 gnd.n179 240.244
R5684 gnd.n6935 gnd.n179 240.244
R5685 gnd.n6936 gnd.n6935 240.244
R5686 gnd.n6936 gnd.n101 240.244
R5687 gnd.n3803 gnd.n3802 240.244
R5688 gnd.n3805 gnd.n3803 240.244
R5689 gnd.n3811 gnd.n3793 240.244
R5690 gnd.n3815 gnd.n3813 240.244
R5691 gnd.n3821 gnd.n3789 240.244
R5692 gnd.n3825 gnd.n3823 240.244
R5693 gnd.n3832 gnd.n3785 240.244
R5694 gnd.n3835 gnd.n3834 240.244
R5695 gnd.n3845 gnd.n1484 240.244
R5696 gnd.n3849 gnd.n3847 240.244
R5697 gnd.n3855 gnd.n1480 240.244
R5698 gnd.n3859 gnd.n3857 240.244
R5699 gnd.n3865 gnd.n1476 240.244
R5700 gnd.n3869 gnd.n3867 240.244
R5701 gnd.n3875 gnd.n1472 240.244
R5702 gnd.n3879 gnd.n3877 240.244
R5703 gnd.n3886 gnd.n1468 240.244
R5704 gnd.n3889 gnd.n3888 240.244
R5705 gnd.n4058 gnd.n1330 240.244
R5706 gnd.n4054 gnd.n1330 240.244
R5707 gnd.n4054 gnd.n1335 240.244
R5708 gnd.n3931 gnd.n1335 240.244
R5709 gnd.n3931 gnd.n1432 240.244
R5710 gnd.n3937 gnd.n1432 240.244
R5711 gnd.n3937 gnd.n1406 240.244
R5712 gnd.n3968 gnd.n1406 240.244
R5713 gnd.n3968 gnd.n1401 240.244
R5714 gnd.n3976 gnd.n1401 240.244
R5715 gnd.n3976 gnd.n1402 240.244
R5716 gnd.n1402 gnd.n1367 240.244
R5717 gnd.n4021 gnd.n1367 240.244
R5718 gnd.n4021 gnd.n1363 240.244
R5719 gnd.n4027 gnd.n1363 240.244
R5720 gnd.n4027 gnd.n322 240.244
R5721 gnd.n6653 gnd.n322 240.244
R5722 gnd.n6653 gnd.n317 240.244
R5723 gnd.n6661 gnd.n317 240.244
R5724 gnd.n6661 gnd.n318 240.244
R5725 gnd.n318 gnd.n267 240.244
R5726 gnd.n6773 gnd.n267 240.244
R5727 gnd.n6773 gnd.n268 240.244
R5728 gnd.n6679 gnd.n268 240.244
R5729 gnd.n6679 gnd.n6678 240.244
R5730 gnd.n6678 gnd.n289 240.244
R5731 gnd.n6751 gnd.n289 240.244
R5732 gnd.n6752 gnd.n6751 240.244
R5733 gnd.n6755 gnd.n6752 240.244
R5734 gnd.n6755 gnd.n257 240.244
R5735 gnd.n6778 gnd.n257 240.244
R5736 gnd.n6778 gnd.n248 240.244
R5737 gnd.n6788 gnd.n248 240.244
R5738 gnd.n6788 gnd.n244 240.244
R5739 gnd.n6794 gnd.n244 240.244
R5740 gnd.n6794 gnd.n231 240.244
R5741 gnd.n6804 gnd.n231 240.244
R5742 gnd.n6804 gnd.n227 240.244
R5743 gnd.n6810 gnd.n227 240.244
R5744 gnd.n6810 gnd.n218 240.244
R5745 gnd.n6820 gnd.n218 240.244
R5746 gnd.n6820 gnd.n214 240.244
R5747 gnd.n6826 gnd.n214 240.244
R5748 gnd.n6826 gnd.n202 240.244
R5749 gnd.n6836 gnd.n202 240.244
R5750 gnd.n6836 gnd.n198 240.244
R5751 gnd.n6842 gnd.n198 240.244
R5752 gnd.n6842 gnd.n187 240.244
R5753 gnd.n6927 gnd.n187 240.244
R5754 gnd.n6927 gnd.n183 240.244
R5755 gnd.n6933 gnd.n183 240.244
R5756 gnd.n6933 gnd.n104 240.244
R5757 gnd.n7013 gnd.n104 240.244
R5758 gnd.n2070 gnd.n1190 240.244
R5759 gnd.n2785 gnd.n2071 240.244
R5760 gnd.n2781 gnd.n2780 240.244
R5761 gnd.n2777 gnd.n2776 240.244
R5762 gnd.n2773 gnd.n2772 240.244
R5763 gnd.n2769 gnd.n2768 240.244
R5764 gnd.n2765 gnd.n2764 240.244
R5765 gnd.n2761 gnd.n2760 240.244
R5766 gnd.n2624 gnd.n2623 240.244
R5767 gnd.n2621 gnd.n2620 240.244
R5768 gnd.n2617 gnd.n2616 240.244
R5769 gnd.n2613 gnd.n2612 240.244
R5770 gnd.n2609 gnd.n2608 240.244
R5771 gnd.n2605 gnd.n2604 240.244
R5772 gnd.n2601 gnd.n2600 240.244
R5773 gnd.n2597 gnd.n2596 240.244
R5774 gnd.n2593 gnd.n2592 240.244
R5775 gnd.n2589 gnd.n2588 240.244
R5776 gnd.n4365 gnd.n933 240.244
R5777 gnd.n937 gnd.n933 240.244
R5778 gnd.n4358 gnd.n937 240.244
R5779 gnd.n4358 gnd.n938 240.244
R5780 gnd.n951 gnd.n938 240.244
R5781 gnd.n2204 gnd.n951 240.244
R5782 gnd.n2204 gnd.n962 240.244
R5783 gnd.n2209 gnd.n962 240.244
R5784 gnd.n2209 gnd.n972 240.244
R5785 gnd.n2212 gnd.n972 240.244
R5786 gnd.n2212 gnd.n982 240.244
R5787 gnd.n2217 gnd.n982 240.244
R5788 gnd.n2217 gnd.n992 240.244
R5789 gnd.n2220 gnd.n992 240.244
R5790 gnd.n2220 gnd.n1002 240.244
R5791 gnd.n2225 gnd.n1002 240.244
R5792 gnd.n2225 gnd.n1012 240.244
R5793 gnd.n2228 gnd.n1012 240.244
R5794 gnd.n2228 gnd.n1022 240.244
R5795 gnd.n2233 gnd.n1022 240.244
R5796 gnd.n2233 gnd.n1032 240.244
R5797 gnd.n2236 gnd.n1032 240.244
R5798 gnd.n2236 gnd.n1042 240.244
R5799 gnd.n2241 gnd.n1042 240.244
R5800 gnd.n2241 gnd.n1050 240.244
R5801 gnd.n2244 gnd.n1050 240.244
R5802 gnd.n2244 gnd.n1060 240.244
R5803 gnd.n2256 gnd.n1060 240.244
R5804 gnd.n2256 gnd.n1067 240.244
R5805 gnd.n2252 gnd.n1067 240.244
R5806 gnd.n2252 gnd.n1077 240.244
R5807 gnd.n2418 gnd.n1077 240.244
R5808 gnd.n2418 gnd.n1087 240.244
R5809 gnd.n2425 gnd.n1087 240.244
R5810 gnd.n2425 gnd.n1097 240.244
R5811 gnd.n2435 gnd.n1097 240.244
R5812 gnd.n2435 gnd.n1108 240.244
R5813 gnd.n2139 gnd.n1108 240.244
R5814 gnd.n2139 gnd.n1118 240.244
R5815 gnd.n2443 gnd.n1118 240.244
R5816 gnd.n2443 gnd.n1129 240.244
R5817 gnd.n2448 gnd.n1129 240.244
R5818 gnd.n2448 gnd.n1139 240.244
R5819 gnd.n2458 gnd.n1139 240.244
R5820 gnd.n2458 gnd.n1150 240.244
R5821 gnd.n2127 gnd.n1150 240.244
R5822 gnd.n2127 gnd.n1160 240.244
R5823 gnd.n2528 gnd.n1160 240.244
R5824 gnd.n2528 gnd.n1171 240.244
R5825 gnd.n2535 gnd.n1171 240.244
R5826 gnd.n2535 gnd.n1182 240.244
R5827 gnd.n2581 gnd.n1182 240.244
R5828 gnd.n2581 gnd.n1192 240.244
R5829 gnd.n887 gnd.n886 240.244
R5830 gnd.n4437 gnd.n886 240.244
R5831 gnd.n4435 gnd.n4434 240.244
R5832 gnd.n4431 gnd.n4430 240.244
R5833 gnd.n4427 gnd.n4426 240.244
R5834 gnd.n4423 gnd.n4422 240.244
R5835 gnd.n4419 gnd.n4418 240.244
R5836 gnd.n4415 gnd.n4414 240.244
R5837 gnd.n4411 gnd.n4410 240.244
R5838 gnd.n4406 gnd.n4405 240.244
R5839 gnd.n4402 gnd.n4401 240.244
R5840 gnd.n4398 gnd.n4397 240.244
R5841 gnd.n4394 gnd.n4393 240.244
R5842 gnd.n4390 gnd.n4389 240.244
R5843 gnd.n4386 gnd.n4385 240.244
R5844 gnd.n4382 gnd.n4381 240.244
R5845 gnd.n4378 gnd.n4377 240.244
R5846 gnd.n4374 gnd.n4373 240.244
R5847 gnd.n928 gnd.n927 240.244
R5848 gnd.n2351 gnd.n888 240.244
R5849 gnd.n2351 gnd.n943 240.244
R5850 gnd.n4356 gnd.n943 240.244
R5851 gnd.n4356 gnd.n944 240.244
R5852 gnd.n4352 gnd.n944 240.244
R5853 gnd.n4352 gnd.n950 240.244
R5854 gnd.n4344 gnd.n950 240.244
R5855 gnd.n4344 gnd.n965 240.244
R5856 gnd.n4340 gnd.n965 240.244
R5857 gnd.n4340 gnd.n971 240.244
R5858 gnd.n4332 gnd.n971 240.244
R5859 gnd.n4332 gnd.n984 240.244
R5860 gnd.n4328 gnd.n984 240.244
R5861 gnd.n4328 gnd.n990 240.244
R5862 gnd.n4320 gnd.n990 240.244
R5863 gnd.n4320 gnd.n1005 240.244
R5864 gnd.n4316 gnd.n1005 240.244
R5865 gnd.n4316 gnd.n1011 240.244
R5866 gnd.n4308 gnd.n1011 240.244
R5867 gnd.n4308 gnd.n1024 240.244
R5868 gnd.n4304 gnd.n1024 240.244
R5869 gnd.n4304 gnd.n1030 240.244
R5870 gnd.n4296 gnd.n1030 240.244
R5871 gnd.n4296 gnd.n1045 240.244
R5872 gnd.n4292 gnd.n1045 240.244
R5873 gnd.n4292 gnd.n1049 240.244
R5874 gnd.n4284 gnd.n1049 240.244
R5875 gnd.n4284 gnd.n1062 240.244
R5876 gnd.n4279 gnd.n1062 240.244
R5877 gnd.n4279 gnd.n1065 240.244
R5878 gnd.n4271 gnd.n1065 240.244
R5879 gnd.n4271 gnd.n1080 240.244
R5880 gnd.n4267 gnd.n1080 240.244
R5881 gnd.n4267 gnd.n1085 240.244
R5882 gnd.n4259 gnd.n1085 240.244
R5883 gnd.n4259 gnd.n1100 240.244
R5884 gnd.n4255 gnd.n1100 240.244
R5885 gnd.n4255 gnd.n1106 240.244
R5886 gnd.n4247 gnd.n1106 240.244
R5887 gnd.n4247 gnd.n1121 240.244
R5888 gnd.n4243 gnd.n1121 240.244
R5889 gnd.n4243 gnd.n1127 240.244
R5890 gnd.n4235 gnd.n1127 240.244
R5891 gnd.n4235 gnd.n1142 240.244
R5892 gnd.n4231 gnd.n1142 240.244
R5893 gnd.n4231 gnd.n1148 240.244
R5894 gnd.n4223 gnd.n1148 240.244
R5895 gnd.n4223 gnd.n1163 240.244
R5896 gnd.n4219 gnd.n1163 240.244
R5897 gnd.n4219 gnd.n1169 240.244
R5898 gnd.n4211 gnd.n1169 240.244
R5899 gnd.n4211 gnd.n1185 240.244
R5900 gnd.n4207 gnd.n1185 240.244
R5901 gnd.n4451 gnd.n4447 240.244
R5902 gnd.n5879 gnd.n5878 240.244
R5903 gnd.n5876 gnd.n4455 240.244
R5904 gnd.n5872 gnd.n5871 240.244
R5905 gnd.n5869 gnd.n4462 240.244
R5906 gnd.n5865 gnd.n5864 240.244
R5907 gnd.n5862 gnd.n4469 240.244
R5908 gnd.n5858 gnd.n5857 240.244
R5909 gnd.n5446 gnd.n5054 240.244
R5910 gnd.n5054 gnd.n5045 240.244
R5911 gnd.n5467 gnd.n5045 240.244
R5912 gnd.n5467 gnd.n5038 240.244
R5913 gnd.n5477 gnd.n5038 240.244
R5914 gnd.n5477 gnd.n5029 240.244
R5915 gnd.n5029 gnd.n5018 240.244
R5916 gnd.n5498 gnd.n5018 240.244
R5917 gnd.n5498 gnd.n5012 240.244
R5918 gnd.n5508 gnd.n5012 240.244
R5919 gnd.n5508 gnd.n5003 240.244
R5920 gnd.n5003 gnd.n4992 240.244
R5921 gnd.n5529 gnd.n4992 240.244
R5922 gnd.n5529 gnd.n4986 240.244
R5923 gnd.n5539 gnd.n4986 240.244
R5924 gnd.n5539 gnd.n4977 240.244
R5925 gnd.n4977 gnd.n4967 240.244
R5926 gnd.n5560 gnd.n4967 240.244
R5927 gnd.n5560 gnd.n4960 240.244
R5928 gnd.n5570 gnd.n4960 240.244
R5929 gnd.n5570 gnd.n4951 240.244
R5930 gnd.n4951 gnd.n4942 240.244
R5931 gnd.n5591 gnd.n4942 240.244
R5932 gnd.n5591 gnd.n4935 240.244
R5933 gnd.n5601 gnd.n4935 240.244
R5934 gnd.n5601 gnd.n4926 240.244
R5935 gnd.n4926 gnd.n4917 240.244
R5936 gnd.n5622 gnd.n4917 240.244
R5937 gnd.n5622 gnd.n4910 240.244
R5938 gnd.n5632 gnd.n4910 240.244
R5939 gnd.n5632 gnd.n4902 240.244
R5940 gnd.n4902 gnd.n4893 240.244
R5941 gnd.n5652 gnd.n4893 240.244
R5942 gnd.n5652 gnd.n4880 240.244
R5943 gnd.n5673 gnd.n4880 240.244
R5944 gnd.n5673 gnd.n4869 240.244
R5945 gnd.n4869 gnd.n4860 240.244
R5946 gnd.n5696 gnd.n4860 240.244
R5947 gnd.n5697 gnd.n5696 240.244
R5948 gnd.n5698 gnd.n5697 240.244
R5949 gnd.n5698 gnd.n4840 240.244
R5950 gnd.n5726 gnd.n4840 240.244
R5951 gnd.n5726 gnd.n4831 240.244
R5952 gnd.n5742 gnd.n4831 240.244
R5953 gnd.n5743 gnd.n5742 240.244
R5954 gnd.n5743 gnd.n4813 240.244
R5955 gnd.n5770 gnd.n4813 240.244
R5956 gnd.n5770 gnd.n4797 240.244
R5957 gnd.n5785 gnd.n4797 240.244
R5958 gnd.n5785 gnd.n5784 240.244
R5959 gnd.n5784 gnd.n4804 240.244
R5960 gnd.n4804 gnd.n4798 240.244
R5961 gnd.n4798 gnd.n856 240.244
R5962 gnd.n5383 gnd.n5382 240.244
R5963 gnd.n5427 gnd.n5382 240.244
R5964 gnd.n5425 gnd.n5424 240.244
R5965 gnd.n5421 gnd.n5420 240.244
R5966 gnd.n5417 gnd.n5416 240.244
R5967 gnd.n5413 gnd.n5412 240.244
R5968 gnd.n5409 gnd.n5408 240.244
R5969 gnd.n5405 gnd.n5404 240.244
R5970 gnd.n5457 gnd.n5052 240.244
R5971 gnd.n5457 gnd.n5047 240.244
R5972 gnd.n5465 gnd.n5047 240.244
R5973 gnd.n5465 gnd.n5048 240.244
R5974 gnd.n5048 gnd.n5027 240.244
R5975 gnd.n5488 gnd.n5027 240.244
R5976 gnd.n5488 gnd.n5021 240.244
R5977 gnd.n5496 gnd.n5021 240.244
R5978 gnd.n5496 gnd.n5023 240.244
R5979 gnd.n5023 gnd.n5001 240.244
R5980 gnd.n5519 gnd.n5001 240.244
R5981 gnd.n5519 gnd.n4995 240.244
R5982 gnd.n5527 gnd.n4995 240.244
R5983 gnd.n5527 gnd.n4997 240.244
R5984 gnd.n4997 gnd.n4975 240.244
R5985 gnd.n5550 gnd.n4975 240.244
R5986 gnd.n5550 gnd.n4970 240.244
R5987 gnd.n5558 gnd.n4970 240.244
R5988 gnd.n5558 gnd.n4971 240.244
R5989 gnd.n4971 gnd.n4949 240.244
R5990 gnd.n5581 gnd.n4949 240.244
R5991 gnd.n5581 gnd.n4944 240.244
R5992 gnd.n5589 gnd.n4944 240.244
R5993 gnd.n5589 gnd.n4945 240.244
R5994 gnd.n4945 gnd.n4924 240.244
R5995 gnd.n5612 gnd.n4924 240.244
R5996 gnd.n5612 gnd.n4919 240.244
R5997 gnd.n5620 gnd.n4919 240.244
R5998 gnd.n5620 gnd.n4920 240.244
R5999 gnd.n4920 gnd.n4900 240.244
R6000 gnd.n5642 gnd.n4900 240.244
R6001 gnd.n5642 gnd.n4895 240.244
R6002 gnd.n5650 gnd.n4895 240.244
R6003 gnd.n5650 gnd.n4896 240.244
R6004 gnd.n4896 gnd.n4868 240.244
R6005 gnd.n5683 gnd.n4868 240.244
R6006 gnd.n5683 gnd.n4863 240.244
R6007 gnd.n5694 gnd.n4863 240.244
R6008 gnd.n5694 gnd.n4864 240.244
R6009 gnd.n5690 gnd.n4864 240.244
R6010 gnd.n5690 gnd.n4838 240.244
R6011 gnd.n5730 gnd.n4838 240.244
R6012 gnd.n5730 gnd.n4833 240.244
R6013 gnd.n5740 gnd.n4833 240.244
R6014 gnd.n5740 gnd.n4834 240.244
R6015 gnd.n4834 gnd.n4811 240.244
R6016 gnd.n5773 gnd.n4811 240.244
R6017 gnd.n5774 gnd.n5773 240.244
R6018 gnd.n5774 gnd.n4806 240.244
R6019 gnd.n5782 gnd.n4806 240.244
R6020 gnd.n5782 gnd.n4807 240.244
R6021 gnd.n4807 gnd.n4446 240.244
R6022 gnd.n5886 gnd.n4446 240.244
R6023 gnd.n4481 gnd.n853 240.244
R6024 gnd.n5847 gnd.n5846 240.244
R6025 gnd.n5844 gnd.n4485 240.244
R6026 gnd.n5840 gnd.n5839 240.244
R6027 gnd.n5837 gnd.n4492 240.244
R6028 gnd.n5833 gnd.n5832 240.244
R6029 gnd.n5830 gnd.n4499 240.244
R6030 gnd.n5826 gnd.n5825 240.244
R6031 gnd.n5823 gnd.n4506 240.244
R6032 gnd.n5819 gnd.n5818 240.244
R6033 gnd.n5816 gnd.n4513 240.244
R6034 gnd.n5812 gnd.n5811 240.244
R6035 gnd.n5809 gnd.n4523 240.244
R6036 gnd.n5201 gnd.n5097 240.244
R6037 gnd.n5207 gnd.n5097 240.244
R6038 gnd.n5207 gnd.n5089 240.244
R6039 gnd.n5217 gnd.n5089 240.244
R6040 gnd.n5217 gnd.n5085 240.244
R6041 gnd.n5223 gnd.n5085 240.244
R6042 gnd.n5223 gnd.n5076 240.244
R6043 gnd.n5233 gnd.n5076 240.244
R6044 gnd.n5233 gnd.n5071 240.244
R6045 gnd.n5374 gnd.n5071 240.244
R6046 gnd.n5374 gnd.n5072 240.244
R6047 gnd.n5072 gnd.n5064 240.244
R6048 gnd.n5369 gnd.n5064 240.244
R6049 gnd.n5369 gnd.n5055 240.244
R6050 gnd.n5366 gnd.n5055 240.244
R6051 gnd.n5366 gnd.n5365 240.244
R6052 gnd.n5365 gnd.n5040 240.244
R6053 gnd.n5360 gnd.n5040 240.244
R6054 gnd.n5360 gnd.n5030 240.244
R6055 gnd.n5357 gnd.n5030 240.244
R6056 gnd.n5357 gnd.n5356 240.244
R6057 gnd.n5356 gnd.n5013 240.244
R6058 gnd.n5352 gnd.n5013 240.244
R6059 gnd.n5352 gnd.n5004 240.244
R6060 gnd.n5349 gnd.n5004 240.244
R6061 gnd.n5349 gnd.n5348 240.244
R6062 gnd.n5348 gnd.n4987 240.244
R6063 gnd.n5344 gnd.n4987 240.244
R6064 gnd.n5344 gnd.n4978 240.244
R6065 gnd.n5289 gnd.n4978 240.244
R6066 gnd.n5290 gnd.n5289 240.244
R6067 gnd.n5290 gnd.n4962 240.244
R6068 gnd.n5286 gnd.n4962 240.244
R6069 gnd.n5286 gnd.n4952 240.244
R6070 gnd.n5282 gnd.n4952 240.244
R6071 gnd.n5282 gnd.n5281 240.244
R6072 gnd.n5281 gnd.n4937 240.244
R6073 gnd.n5276 gnd.n4937 240.244
R6074 gnd.n5276 gnd.n4927 240.244
R6075 gnd.n5273 gnd.n4927 240.244
R6076 gnd.n5273 gnd.n5271 240.244
R6077 gnd.n5271 gnd.n4912 240.244
R6078 gnd.n5267 gnd.n4912 240.244
R6079 gnd.n5267 gnd.n4903 240.244
R6080 gnd.n4903 gnd.n4886 240.244
R6081 gnd.n5662 gnd.n4886 240.244
R6082 gnd.n5662 gnd.n4882 240.244
R6083 gnd.n5670 gnd.n4882 240.244
R6084 gnd.n5670 gnd.n4870 240.244
R6085 gnd.n4870 gnd.n4851 240.244
R6086 gnd.n5706 gnd.n4851 240.244
R6087 gnd.n5706 gnd.n4846 240.244
R6088 gnd.n5714 gnd.n4846 240.244
R6089 gnd.n5714 gnd.n4847 240.244
R6090 gnd.n4847 gnd.n4824 240.244
R6091 gnd.n5751 gnd.n4824 240.244
R6092 gnd.n5751 gnd.n4819 240.244
R6093 gnd.n5759 gnd.n4819 240.244
R6094 gnd.n5759 gnd.n4820 240.244
R6095 gnd.n4820 gnd.n4531 240.244
R6096 gnd.n5792 gnd.n4531 240.244
R6097 gnd.n5792 gnd.n4532 240.244
R6098 gnd.n4532 gnd.n845 240.244
R6099 gnd.n5799 gnd.n845 240.244
R6100 gnd.n5799 gnd.n855 240.244
R6101 gnd.n5193 gnd.n5191 240.244
R6102 gnd.n5191 gnd.n5190 240.244
R6103 gnd.n5187 gnd.n5186 240.244
R6104 gnd.n5184 gnd.n5110 240.244
R6105 gnd.n5180 gnd.n5178 240.244
R6106 gnd.n5176 gnd.n5116 240.244
R6107 gnd.n5172 gnd.n5170 240.244
R6108 gnd.n5168 gnd.n5122 240.244
R6109 gnd.n5164 gnd.n5162 240.244
R6110 gnd.n5160 gnd.n5128 240.244
R6111 gnd.n5156 gnd.n5154 240.244
R6112 gnd.n5152 gnd.n5134 240.244
R6113 gnd.n5147 gnd.n5145 240.244
R6114 gnd.n5199 gnd.n5095 240.244
R6115 gnd.n5209 gnd.n5095 240.244
R6116 gnd.n5209 gnd.n5091 240.244
R6117 gnd.n5215 gnd.n5091 240.244
R6118 gnd.n5215 gnd.n5083 240.244
R6119 gnd.n5225 gnd.n5083 240.244
R6120 gnd.n5225 gnd.n5079 240.244
R6121 gnd.n5231 gnd.n5079 240.244
R6122 gnd.n5231 gnd.n5070 240.244
R6123 gnd.n5436 gnd.n5070 240.244
R6124 gnd.n5436 gnd.n5065 240.244
R6125 gnd.n5443 gnd.n5065 240.244
R6126 gnd.n5443 gnd.n5057 240.244
R6127 gnd.n5454 gnd.n5057 240.244
R6128 gnd.n5454 gnd.n5058 240.244
R6129 gnd.n5058 gnd.n5041 240.244
R6130 gnd.n5474 gnd.n5041 240.244
R6131 gnd.n5474 gnd.n5032 240.244
R6132 gnd.n5485 gnd.n5032 240.244
R6133 gnd.n5485 gnd.n5033 240.244
R6134 gnd.n5033 gnd.n5014 240.244
R6135 gnd.n5505 gnd.n5014 240.244
R6136 gnd.n5505 gnd.n5006 240.244
R6137 gnd.n5516 gnd.n5006 240.244
R6138 gnd.n5516 gnd.n5007 240.244
R6139 gnd.n5007 gnd.n4988 240.244
R6140 gnd.n5536 gnd.n4988 240.244
R6141 gnd.n5536 gnd.n4980 240.244
R6142 gnd.n5547 gnd.n4980 240.244
R6143 gnd.n5547 gnd.n4981 240.244
R6144 gnd.n4981 gnd.n4963 240.244
R6145 gnd.n5567 gnd.n4963 240.244
R6146 gnd.n5567 gnd.n4954 240.244
R6147 gnd.n5578 gnd.n4954 240.244
R6148 gnd.n5578 gnd.n4955 240.244
R6149 gnd.n4955 gnd.n4938 240.244
R6150 gnd.n5598 gnd.n4938 240.244
R6151 gnd.n5598 gnd.n4929 240.244
R6152 gnd.n5609 gnd.n4929 240.244
R6153 gnd.n5609 gnd.n4930 240.244
R6154 gnd.n4930 gnd.n4913 240.244
R6155 gnd.n5629 gnd.n4913 240.244
R6156 gnd.n5629 gnd.n4905 240.244
R6157 gnd.n5639 gnd.n4905 240.244
R6158 gnd.n5639 gnd.n4888 240.244
R6159 gnd.n5660 gnd.n4888 240.244
R6160 gnd.n5660 gnd.n4889 240.244
R6161 gnd.n4889 gnd.n4872 240.244
R6162 gnd.n5680 gnd.n4872 240.244
R6163 gnd.n5680 gnd.n4854 240.244
R6164 gnd.n5704 gnd.n4854 240.244
R6165 gnd.n5704 gnd.n4844 240.244
R6166 gnd.n5717 gnd.n4844 240.244
R6167 gnd.n5718 gnd.n5717 240.244
R6168 gnd.n5718 gnd.n4825 240.244
R6169 gnd.n5749 gnd.n4825 240.244
R6170 gnd.n5749 gnd.n4817 240.244
R6171 gnd.n5762 gnd.n4817 240.244
R6172 gnd.n5763 gnd.n5762 240.244
R6173 gnd.n5763 gnd.n4535 240.244
R6174 gnd.n5790 gnd.n4535 240.244
R6175 gnd.n5790 gnd.n847 240.244
R6176 gnd.n5893 gnd.n847 240.244
R6177 gnd.n5893 gnd.n848 240.244
R6178 gnd.n5889 gnd.n848 240.244
R6179 gnd.n6852 gnd.n6851 240.244
R6180 gnd.n6857 gnd.n6854 240.244
R6181 gnd.n6860 gnd.n6859 240.244
R6182 gnd.n6865 gnd.n6862 240.244
R6183 gnd.n6868 gnd.n6867 240.244
R6184 gnd.n6873 gnd.n6870 240.244
R6185 gnd.n6876 gnd.n6875 240.244
R6186 gnd.n6881 gnd.n6878 240.244
R6187 gnd.n6887 gnd.n6883 240.244
R6188 gnd.n3906 gnd.n1326 240.244
R6189 gnd.n3906 gnd.n1338 240.244
R6190 gnd.n1458 gnd.n1338 240.244
R6191 gnd.n1458 gnd.n1437 240.244
R6192 gnd.n3913 gnd.n1437 240.244
R6193 gnd.n3913 gnd.n1431 240.244
R6194 gnd.n3920 gnd.n1431 240.244
R6195 gnd.n3920 gnd.n1409 240.244
R6196 gnd.n1409 gnd.n1396 240.244
R6197 gnd.n3978 gnd.n1396 240.244
R6198 gnd.n3978 gnd.n1397 240.244
R6199 gnd.n1397 gnd.n1393 240.244
R6200 gnd.n1393 gnd.n1370 240.244
R6201 gnd.n3985 gnd.n1370 240.244
R6202 gnd.n3985 gnd.n1361 240.244
R6203 gnd.n3992 gnd.n1361 240.244
R6204 gnd.n3992 gnd.n325 240.244
R6205 gnd.n325 gnd.n311 240.244
R6206 gnd.n6663 gnd.n311 240.244
R6207 gnd.n6663 gnd.n312 240.244
R6208 gnd.n312 gnd.n308 240.244
R6209 gnd.n308 gnd.n271 240.244
R6210 gnd.n6670 gnd.n271 240.244
R6211 gnd.n6670 gnd.n301 240.244
R6212 gnd.n6676 gnd.n301 240.244
R6213 gnd.n6676 gnd.n304 240.244
R6214 gnd.n304 gnd.n66 240.244
R6215 gnd.n67 gnd.n66 240.244
R6216 gnd.n68 gnd.n67 240.244
R6217 gnd.n287 gnd.n68 240.244
R6218 gnd.n287 gnd.n71 240.244
R6219 gnd.n72 gnd.n71 240.244
R6220 gnd.n73 gnd.n72 240.244
R6221 gnd.n241 gnd.n73 240.244
R6222 gnd.n241 gnd.n76 240.244
R6223 gnd.n77 gnd.n76 240.244
R6224 gnd.n78 gnd.n77 240.244
R6225 gnd.n234 gnd.n78 240.244
R6226 gnd.n234 gnd.n81 240.244
R6227 gnd.n82 gnd.n81 240.244
R6228 gnd.n83 gnd.n82 240.244
R6229 gnd.n211 gnd.n83 240.244
R6230 gnd.n211 gnd.n86 240.244
R6231 gnd.n87 gnd.n86 240.244
R6232 gnd.n88 gnd.n87 240.244
R6233 gnd.n6717 gnd.n88 240.244
R6234 gnd.n6717 gnd.n91 240.244
R6235 gnd.n92 gnd.n91 240.244
R6236 gnd.n93 gnd.n92 240.244
R6237 gnd.n180 gnd.n93 240.244
R6238 gnd.n180 gnd.n96 240.244
R6239 gnd.n97 gnd.n96 240.244
R6240 gnd.n7015 gnd.n97 240.244
R6241 gnd.n3454 gnd.n3452 240.244
R6242 gnd.n3469 gnd.n3435 240.244
R6243 gnd.n3473 gnd.n3471 240.244
R6244 gnd.n3488 gnd.n3426 240.244
R6245 gnd.n3492 gnd.n3490 240.244
R6246 gnd.n3507 gnd.n3417 240.244
R6247 gnd.n3511 gnd.n3509 240.244
R6248 gnd.n3528 gnd.n3408 240.244
R6249 gnd.n3531 gnd.n3530 240.244
R6250 gnd.n1340 gnd.n1328 240.244
R6251 gnd.n4052 gnd.n1340 240.244
R6252 gnd.n4052 gnd.n1341 240.244
R6253 gnd.n1346 gnd.n1341 240.244
R6254 gnd.n1347 gnd.n1346 240.244
R6255 gnd.n1348 gnd.n1347 240.244
R6256 gnd.n3921 gnd.n1348 240.244
R6257 gnd.n3921 gnd.n1351 240.244
R6258 gnd.n1352 gnd.n1351 240.244
R6259 gnd.n1353 gnd.n1352 240.244
R6260 gnd.n1420 gnd.n1353 240.244
R6261 gnd.n1420 gnd.n1356 240.244
R6262 gnd.n1357 gnd.n1356 240.244
R6263 gnd.n1358 gnd.n1357 240.244
R6264 gnd.n4029 gnd.n1358 240.244
R6265 gnd.n4029 gnd.n326 240.244
R6266 gnd.n6651 gnd.n326 240.244
R6267 gnd.n6651 gnd.n327 240.244
R6268 gnd.n327 gnd.n316 240.244
R6269 gnd.n6644 gnd.n316 240.244
R6270 gnd.n6644 gnd.n272 240.244
R6271 gnd.n6771 gnd.n272 240.244
R6272 gnd.n6771 gnd.n273 240.244
R6273 gnd.n278 gnd.n273 240.244
R6274 gnd.n279 gnd.n278 240.244
R6275 gnd.n280 gnd.n279 240.244
R6276 gnd.n6749 gnd.n280 240.244
R6277 gnd.n6749 gnd.n284 240.244
R6278 gnd.n6757 gnd.n284 240.244
R6279 gnd.n6757 gnd.n255 240.244
R6280 gnd.n6780 gnd.n255 240.244
R6281 gnd.n6780 gnd.n251 240.244
R6282 gnd.n6786 gnd.n251 240.244
R6283 gnd.n6786 gnd.n240 240.244
R6284 gnd.n6796 gnd.n240 240.244
R6285 gnd.n6796 gnd.n236 240.244
R6286 gnd.n6802 gnd.n236 240.244
R6287 gnd.n6802 gnd.n225 240.244
R6288 gnd.n6812 gnd.n225 240.244
R6289 gnd.n6812 gnd.n221 240.244
R6290 gnd.n6818 gnd.n221 240.244
R6291 gnd.n6818 gnd.n210 240.244
R6292 gnd.n6828 gnd.n210 240.244
R6293 gnd.n6828 gnd.n206 240.244
R6294 gnd.n6834 gnd.n206 240.244
R6295 gnd.n6834 gnd.n196 240.244
R6296 gnd.n6844 gnd.n196 240.244
R6297 gnd.n6844 gnd.n190 240.244
R6298 gnd.n6925 gnd.n190 240.244
R6299 gnd.n6925 gnd.n191 240.244
R6300 gnd.n191 gnd.n182 240.244
R6301 gnd.n6849 gnd.n182 240.244
R6302 gnd.n6849 gnd.n103 240.244
R6303 gnd.n2037 gnd.n1195 240.244
R6304 gnd.n2038 gnd.n1987 240.244
R6305 gnd.n2041 gnd.n1988 240.244
R6306 gnd.n1997 gnd.n1996 240.244
R6307 gnd.n2043 gnd.n2004 240.244
R6308 gnd.n2046 gnd.n2005 240.244
R6309 gnd.n2015 gnd.n2014 240.244
R6310 gnd.n2048 gnd.n2022 240.244
R6311 gnd.n2034 gnd.n2023 240.244
R6312 gnd.n2353 gnd.n2273 240.244
R6313 gnd.n2354 gnd.n2353 240.244
R6314 gnd.n2354 gnd.n940 240.244
R6315 gnd.n2359 gnd.n940 240.244
R6316 gnd.n2359 gnd.n952 240.244
R6317 gnd.n2362 gnd.n952 240.244
R6318 gnd.n2362 gnd.n963 240.244
R6319 gnd.n2367 gnd.n963 240.244
R6320 gnd.n2367 gnd.n973 240.244
R6321 gnd.n2370 gnd.n973 240.244
R6322 gnd.n2370 gnd.n983 240.244
R6323 gnd.n2375 gnd.n983 240.244
R6324 gnd.n2375 gnd.n993 240.244
R6325 gnd.n2378 gnd.n993 240.244
R6326 gnd.n2378 gnd.n1003 240.244
R6327 gnd.n2383 gnd.n1003 240.244
R6328 gnd.n2383 gnd.n1013 240.244
R6329 gnd.n2386 gnd.n1013 240.244
R6330 gnd.n2386 gnd.n1023 240.244
R6331 gnd.n2391 gnd.n1023 240.244
R6332 gnd.n2391 gnd.n1033 240.244
R6333 gnd.n2394 gnd.n1033 240.244
R6334 gnd.n2394 gnd.n1043 240.244
R6335 gnd.n2399 gnd.n1043 240.244
R6336 gnd.n2399 gnd.n1051 240.244
R6337 gnd.n2402 gnd.n1051 240.244
R6338 gnd.n2402 gnd.n1061 240.244
R6339 gnd.n2258 gnd.n1061 240.244
R6340 gnd.n2258 gnd.n1068 240.244
R6341 gnd.n2410 gnd.n1068 240.244
R6342 gnd.n2410 gnd.n1078 240.244
R6343 gnd.n2416 gnd.n1078 240.244
R6344 gnd.n2416 gnd.n1088 240.244
R6345 gnd.n2427 gnd.n1088 240.244
R6346 gnd.n2427 gnd.n1098 240.244
R6347 gnd.n2433 gnd.n1098 240.244
R6348 gnd.n2433 gnd.n1109 240.244
R6349 gnd.n2472 gnd.n1109 240.244
R6350 gnd.n2472 gnd.n1119 240.244
R6351 gnd.n2144 gnd.n1119 240.244
R6352 gnd.n2144 gnd.n1130 240.244
R6353 gnd.n2145 gnd.n1130 240.244
R6354 gnd.n2145 gnd.n1140 240.244
R6355 gnd.n2460 gnd.n1140 240.244
R6356 gnd.n2460 gnd.n1151 240.244
R6357 gnd.n2520 gnd.n1151 240.244
R6358 gnd.n2520 gnd.n1161 240.244
R6359 gnd.n2526 gnd.n1161 240.244
R6360 gnd.n2526 gnd.n1172 240.244
R6361 gnd.n2537 gnd.n1172 240.244
R6362 gnd.n2537 gnd.n1183 240.244
R6363 gnd.n2579 gnd.n1183 240.244
R6364 gnd.n2579 gnd.n1193 240.244
R6365 gnd.n2333 gnd.n2332 240.244
R6366 gnd.n2329 gnd.n2328 240.244
R6367 gnd.n2325 gnd.n2324 240.244
R6368 gnd.n2321 gnd.n2320 240.244
R6369 gnd.n2317 gnd.n2316 240.244
R6370 gnd.n2313 gnd.n2312 240.244
R6371 gnd.n2309 gnd.n2308 240.244
R6372 gnd.n2305 gnd.n2304 240.244
R6373 gnd.n2293 gnd.n884 240.244
R6374 gnd.n2345 gnd.n2274 240.244
R6375 gnd.n2345 gnd.n2275 240.244
R6376 gnd.n2275 gnd.n942 240.244
R6377 gnd.n954 gnd.n942 240.244
R6378 gnd.n4350 gnd.n954 240.244
R6379 gnd.n4350 gnd.n955 240.244
R6380 gnd.n4346 gnd.n955 240.244
R6381 gnd.n4346 gnd.n961 240.244
R6382 gnd.n4338 gnd.n961 240.244
R6383 gnd.n4338 gnd.n974 240.244
R6384 gnd.n4334 gnd.n974 240.244
R6385 gnd.n4334 gnd.n980 240.244
R6386 gnd.n4326 gnd.n980 240.244
R6387 gnd.n4326 gnd.n995 240.244
R6388 gnd.n4322 gnd.n995 240.244
R6389 gnd.n4322 gnd.n1001 240.244
R6390 gnd.n4314 gnd.n1001 240.244
R6391 gnd.n4314 gnd.n1014 240.244
R6392 gnd.n4310 gnd.n1014 240.244
R6393 gnd.n4310 gnd.n1020 240.244
R6394 gnd.n4302 gnd.n1020 240.244
R6395 gnd.n4302 gnd.n1035 240.244
R6396 gnd.n4298 gnd.n1035 240.244
R6397 gnd.n4298 gnd.n1041 240.244
R6398 gnd.n4290 gnd.n1041 240.244
R6399 gnd.n4290 gnd.n1052 240.244
R6400 gnd.n4286 gnd.n1052 240.244
R6401 gnd.n4286 gnd.n1058 240.244
R6402 gnd.n4277 gnd.n1058 240.244
R6403 gnd.n4277 gnd.n1070 240.244
R6404 gnd.n4273 gnd.n1070 240.244
R6405 gnd.n4273 gnd.n1076 240.244
R6406 gnd.n4265 gnd.n1076 240.244
R6407 gnd.n4265 gnd.n1089 240.244
R6408 gnd.n4261 gnd.n1089 240.244
R6409 gnd.n4261 gnd.n1095 240.244
R6410 gnd.n4253 gnd.n1095 240.244
R6411 gnd.n4253 gnd.n1111 240.244
R6412 gnd.n4249 gnd.n1111 240.244
R6413 gnd.n4249 gnd.n1117 240.244
R6414 gnd.n4241 gnd.n1117 240.244
R6415 gnd.n4241 gnd.n1131 240.244
R6416 gnd.n4237 gnd.n1131 240.244
R6417 gnd.n4237 gnd.n1137 240.244
R6418 gnd.n4229 gnd.n1137 240.244
R6419 gnd.n4229 gnd.n1153 240.244
R6420 gnd.n4225 gnd.n1153 240.244
R6421 gnd.n4225 gnd.n1159 240.244
R6422 gnd.n4217 gnd.n1159 240.244
R6423 gnd.n4217 gnd.n1174 240.244
R6424 gnd.n4213 gnd.n1174 240.244
R6425 gnd.n4213 gnd.n1180 240.244
R6426 gnd.n4205 gnd.n1180 240.244
R6427 gnd.n6065 gnd.n673 240.244
R6428 gnd.n6071 gnd.n673 240.244
R6429 gnd.n6071 gnd.n671 240.244
R6430 gnd.n6075 gnd.n671 240.244
R6431 gnd.n6075 gnd.n667 240.244
R6432 gnd.n6081 gnd.n667 240.244
R6433 gnd.n6081 gnd.n665 240.244
R6434 gnd.n6085 gnd.n665 240.244
R6435 gnd.n6085 gnd.n661 240.244
R6436 gnd.n6091 gnd.n661 240.244
R6437 gnd.n6091 gnd.n659 240.244
R6438 gnd.n6095 gnd.n659 240.244
R6439 gnd.n6095 gnd.n655 240.244
R6440 gnd.n6101 gnd.n655 240.244
R6441 gnd.n6101 gnd.n653 240.244
R6442 gnd.n6105 gnd.n653 240.244
R6443 gnd.n6105 gnd.n649 240.244
R6444 gnd.n6111 gnd.n649 240.244
R6445 gnd.n6111 gnd.n647 240.244
R6446 gnd.n6115 gnd.n647 240.244
R6447 gnd.n6115 gnd.n643 240.244
R6448 gnd.n6121 gnd.n643 240.244
R6449 gnd.n6121 gnd.n641 240.244
R6450 gnd.n6125 gnd.n641 240.244
R6451 gnd.n6125 gnd.n637 240.244
R6452 gnd.n6131 gnd.n637 240.244
R6453 gnd.n6131 gnd.n635 240.244
R6454 gnd.n6135 gnd.n635 240.244
R6455 gnd.n6135 gnd.n631 240.244
R6456 gnd.n6141 gnd.n631 240.244
R6457 gnd.n6141 gnd.n629 240.244
R6458 gnd.n6145 gnd.n629 240.244
R6459 gnd.n6145 gnd.n625 240.244
R6460 gnd.n6151 gnd.n625 240.244
R6461 gnd.n6151 gnd.n623 240.244
R6462 gnd.n6155 gnd.n623 240.244
R6463 gnd.n6155 gnd.n619 240.244
R6464 gnd.n6161 gnd.n619 240.244
R6465 gnd.n6161 gnd.n617 240.244
R6466 gnd.n6165 gnd.n617 240.244
R6467 gnd.n6165 gnd.n613 240.244
R6468 gnd.n6171 gnd.n613 240.244
R6469 gnd.n6171 gnd.n611 240.244
R6470 gnd.n6175 gnd.n611 240.244
R6471 gnd.n6175 gnd.n607 240.244
R6472 gnd.n6181 gnd.n607 240.244
R6473 gnd.n6181 gnd.n605 240.244
R6474 gnd.n6185 gnd.n605 240.244
R6475 gnd.n6185 gnd.n601 240.244
R6476 gnd.n6191 gnd.n601 240.244
R6477 gnd.n6191 gnd.n599 240.244
R6478 gnd.n6195 gnd.n599 240.244
R6479 gnd.n6195 gnd.n595 240.244
R6480 gnd.n6201 gnd.n595 240.244
R6481 gnd.n6201 gnd.n593 240.244
R6482 gnd.n6205 gnd.n593 240.244
R6483 gnd.n6205 gnd.n589 240.244
R6484 gnd.n6211 gnd.n589 240.244
R6485 gnd.n6211 gnd.n587 240.244
R6486 gnd.n6215 gnd.n587 240.244
R6487 gnd.n6215 gnd.n583 240.244
R6488 gnd.n6221 gnd.n583 240.244
R6489 gnd.n6221 gnd.n581 240.244
R6490 gnd.n6225 gnd.n581 240.244
R6491 gnd.n6225 gnd.n577 240.244
R6492 gnd.n6231 gnd.n577 240.244
R6493 gnd.n6231 gnd.n575 240.244
R6494 gnd.n6235 gnd.n575 240.244
R6495 gnd.n6235 gnd.n571 240.244
R6496 gnd.n6241 gnd.n571 240.244
R6497 gnd.n6241 gnd.n569 240.244
R6498 gnd.n6245 gnd.n569 240.244
R6499 gnd.n6245 gnd.n565 240.244
R6500 gnd.n6251 gnd.n565 240.244
R6501 gnd.n6251 gnd.n563 240.244
R6502 gnd.n6255 gnd.n563 240.244
R6503 gnd.n6255 gnd.n559 240.244
R6504 gnd.n6261 gnd.n559 240.244
R6505 gnd.n6261 gnd.n557 240.244
R6506 gnd.n6265 gnd.n557 240.244
R6507 gnd.n6265 gnd.n553 240.244
R6508 gnd.n6271 gnd.n553 240.244
R6509 gnd.n6271 gnd.n551 240.244
R6510 gnd.n6275 gnd.n551 240.244
R6511 gnd.n6275 gnd.n547 240.244
R6512 gnd.n6281 gnd.n547 240.244
R6513 gnd.n6281 gnd.n545 240.244
R6514 gnd.n6285 gnd.n545 240.244
R6515 gnd.n6285 gnd.n541 240.244
R6516 gnd.n6291 gnd.n541 240.244
R6517 gnd.n6291 gnd.n539 240.244
R6518 gnd.n6295 gnd.n539 240.244
R6519 gnd.n6295 gnd.n535 240.244
R6520 gnd.n6301 gnd.n535 240.244
R6521 gnd.n6301 gnd.n533 240.244
R6522 gnd.n6305 gnd.n533 240.244
R6523 gnd.n6305 gnd.n529 240.244
R6524 gnd.n6311 gnd.n529 240.244
R6525 gnd.n6311 gnd.n527 240.244
R6526 gnd.n6315 gnd.n527 240.244
R6527 gnd.n6315 gnd.n523 240.244
R6528 gnd.n6321 gnd.n523 240.244
R6529 gnd.n6321 gnd.n521 240.244
R6530 gnd.n6325 gnd.n521 240.244
R6531 gnd.n6325 gnd.n517 240.244
R6532 gnd.n6331 gnd.n517 240.244
R6533 gnd.n6331 gnd.n515 240.244
R6534 gnd.n6335 gnd.n515 240.244
R6535 gnd.n6335 gnd.n511 240.244
R6536 gnd.n6341 gnd.n511 240.244
R6537 gnd.n6341 gnd.n509 240.244
R6538 gnd.n6345 gnd.n509 240.244
R6539 gnd.n6345 gnd.n505 240.244
R6540 gnd.n6351 gnd.n505 240.244
R6541 gnd.n6351 gnd.n503 240.244
R6542 gnd.n6355 gnd.n503 240.244
R6543 gnd.n6355 gnd.n499 240.244
R6544 gnd.n6361 gnd.n499 240.244
R6545 gnd.n6361 gnd.n497 240.244
R6546 gnd.n6365 gnd.n497 240.244
R6547 gnd.n6365 gnd.n493 240.244
R6548 gnd.n6371 gnd.n493 240.244
R6549 gnd.n6371 gnd.n491 240.244
R6550 gnd.n6375 gnd.n491 240.244
R6551 gnd.n6375 gnd.n487 240.244
R6552 gnd.n6381 gnd.n487 240.244
R6553 gnd.n6381 gnd.n485 240.244
R6554 gnd.n6385 gnd.n485 240.244
R6555 gnd.n6385 gnd.n481 240.244
R6556 gnd.n6391 gnd.n481 240.244
R6557 gnd.n6391 gnd.n479 240.244
R6558 gnd.n6395 gnd.n479 240.244
R6559 gnd.n6395 gnd.n475 240.244
R6560 gnd.n6401 gnd.n475 240.244
R6561 gnd.n6401 gnd.n473 240.244
R6562 gnd.n6405 gnd.n473 240.244
R6563 gnd.n6405 gnd.n469 240.244
R6564 gnd.n6412 gnd.n469 240.244
R6565 gnd.n6412 gnd.n467 240.244
R6566 gnd.n6416 gnd.n467 240.244
R6567 gnd.n6416 gnd.n464 240.244
R6568 gnd.n6422 gnd.n462 240.244
R6569 gnd.n6426 gnd.n462 240.244
R6570 gnd.n6426 gnd.n458 240.244
R6571 gnd.n6432 gnd.n458 240.244
R6572 gnd.n6432 gnd.n456 240.244
R6573 gnd.n6436 gnd.n456 240.244
R6574 gnd.n6436 gnd.n452 240.244
R6575 gnd.n6442 gnd.n452 240.244
R6576 gnd.n6442 gnd.n450 240.244
R6577 gnd.n6446 gnd.n450 240.244
R6578 gnd.n6446 gnd.n446 240.244
R6579 gnd.n6452 gnd.n446 240.244
R6580 gnd.n6452 gnd.n444 240.244
R6581 gnd.n6456 gnd.n444 240.244
R6582 gnd.n6456 gnd.n440 240.244
R6583 gnd.n6462 gnd.n440 240.244
R6584 gnd.n6462 gnd.n438 240.244
R6585 gnd.n6466 gnd.n438 240.244
R6586 gnd.n6466 gnd.n434 240.244
R6587 gnd.n6472 gnd.n434 240.244
R6588 gnd.n6472 gnd.n432 240.244
R6589 gnd.n6476 gnd.n432 240.244
R6590 gnd.n6476 gnd.n428 240.244
R6591 gnd.n6482 gnd.n428 240.244
R6592 gnd.n6482 gnd.n426 240.244
R6593 gnd.n6486 gnd.n426 240.244
R6594 gnd.n6486 gnd.n422 240.244
R6595 gnd.n6492 gnd.n422 240.244
R6596 gnd.n6492 gnd.n420 240.244
R6597 gnd.n6496 gnd.n420 240.244
R6598 gnd.n6496 gnd.n416 240.244
R6599 gnd.n6502 gnd.n416 240.244
R6600 gnd.n6502 gnd.n414 240.244
R6601 gnd.n6506 gnd.n414 240.244
R6602 gnd.n6506 gnd.n410 240.244
R6603 gnd.n6512 gnd.n410 240.244
R6604 gnd.n6512 gnd.n408 240.244
R6605 gnd.n6516 gnd.n408 240.244
R6606 gnd.n6516 gnd.n404 240.244
R6607 gnd.n6522 gnd.n404 240.244
R6608 gnd.n6522 gnd.n402 240.244
R6609 gnd.n6526 gnd.n402 240.244
R6610 gnd.n6526 gnd.n398 240.244
R6611 gnd.n6532 gnd.n398 240.244
R6612 gnd.n6532 gnd.n396 240.244
R6613 gnd.n6536 gnd.n396 240.244
R6614 gnd.n6536 gnd.n392 240.244
R6615 gnd.n6542 gnd.n392 240.244
R6616 gnd.n6542 gnd.n390 240.244
R6617 gnd.n6546 gnd.n390 240.244
R6618 gnd.n6546 gnd.n386 240.244
R6619 gnd.n6552 gnd.n386 240.244
R6620 gnd.n6552 gnd.n384 240.244
R6621 gnd.n6556 gnd.n384 240.244
R6622 gnd.n6556 gnd.n380 240.244
R6623 gnd.n6562 gnd.n380 240.244
R6624 gnd.n6562 gnd.n378 240.244
R6625 gnd.n6566 gnd.n378 240.244
R6626 gnd.n6566 gnd.n374 240.244
R6627 gnd.n6572 gnd.n374 240.244
R6628 gnd.n6572 gnd.n372 240.244
R6629 gnd.n6576 gnd.n372 240.244
R6630 gnd.n6576 gnd.n368 240.244
R6631 gnd.n6582 gnd.n368 240.244
R6632 gnd.n6582 gnd.n366 240.244
R6633 gnd.n6586 gnd.n366 240.244
R6634 gnd.n6586 gnd.n362 240.244
R6635 gnd.n6592 gnd.n362 240.244
R6636 gnd.n6592 gnd.n360 240.244
R6637 gnd.n6596 gnd.n360 240.244
R6638 gnd.n6596 gnd.n356 240.244
R6639 gnd.n6602 gnd.n356 240.244
R6640 gnd.n6602 gnd.n354 240.244
R6641 gnd.n6606 gnd.n354 240.244
R6642 gnd.n6606 gnd.n350 240.244
R6643 gnd.n6612 gnd.n350 240.244
R6644 gnd.n6612 gnd.n348 240.244
R6645 gnd.n6616 gnd.n348 240.244
R6646 gnd.n6616 gnd.n344 240.244
R6647 gnd.n6622 gnd.n344 240.244
R6648 gnd.n6622 gnd.n342 240.244
R6649 gnd.n6627 gnd.n342 240.244
R6650 gnd.n6627 gnd.n338 240.244
R6651 gnd.n6633 gnd.n338 240.244
R6652 gnd.n2165 gnd.n2164 240.244
R6653 gnd.n2165 gnd.n2156 240.244
R6654 gnd.n2182 gnd.n2156 240.244
R6655 gnd.n2182 gnd.n2157 240.244
R6656 gnd.n2178 gnd.n2157 240.244
R6657 gnd.n2178 gnd.n2177 240.244
R6658 gnd.n2177 gnd.n2137 240.244
R6659 gnd.n2475 gnd.n2137 240.244
R6660 gnd.n2476 gnd.n2475 240.244
R6661 gnd.n2477 gnd.n2476 240.244
R6662 gnd.n2477 gnd.n2133 240.244
R6663 gnd.n2483 gnd.n2133 240.244
R6664 gnd.n2484 gnd.n2483 240.244
R6665 gnd.n2485 gnd.n2484 240.244
R6666 gnd.n2485 gnd.n2128 240.244
R6667 gnd.n2517 gnd.n2128 240.244
R6668 gnd.n2517 gnd.n2129 240.244
R6669 gnd.n2513 gnd.n2129 240.244
R6670 gnd.n2513 gnd.n2512 240.244
R6671 gnd.n2512 gnd.n2511 240.244
R6672 gnd.n2511 gnd.n2493 240.244
R6673 gnd.n2507 gnd.n2493 240.244
R6674 gnd.n2507 gnd.n2506 240.244
R6675 gnd.n2506 gnd.n2505 240.244
R6676 gnd.n2505 gnd.n2499 240.244
R6677 gnd.n2499 gnd.n1965 240.244
R6678 gnd.n2839 gnd.n1965 240.244
R6679 gnd.n2839 gnd.n1961 240.244
R6680 gnd.n2845 gnd.n1961 240.244
R6681 gnd.n2845 gnd.n1954 240.244
R6682 gnd.n2859 gnd.n1954 240.244
R6683 gnd.n2859 gnd.n1950 240.244
R6684 gnd.n2865 gnd.n1950 240.244
R6685 gnd.n2865 gnd.n1941 240.244
R6686 gnd.n2879 gnd.n1941 240.244
R6687 gnd.n2879 gnd.n1937 240.244
R6688 gnd.n2885 gnd.n1937 240.244
R6689 gnd.n2885 gnd.n1928 240.244
R6690 gnd.n2899 gnd.n1928 240.244
R6691 gnd.n2899 gnd.n1924 240.244
R6692 gnd.n2905 gnd.n1924 240.244
R6693 gnd.n2905 gnd.n1915 240.244
R6694 gnd.n2919 gnd.n1915 240.244
R6695 gnd.n2919 gnd.n1911 240.244
R6696 gnd.n2925 gnd.n1911 240.244
R6697 gnd.n2925 gnd.n1900 240.244
R6698 gnd.n2957 gnd.n1900 240.244
R6699 gnd.n2957 gnd.n1896 240.244
R6700 gnd.n2963 gnd.n1896 240.244
R6701 gnd.n2963 gnd.n1825 240.244
R6702 gnd.n2984 gnd.n1825 240.244
R6703 gnd.n2984 gnd.n1820 240.244
R6704 gnd.n2995 gnd.n1820 240.244
R6705 gnd.n2995 gnd.n1821 240.244
R6706 gnd.n2991 gnd.n1821 240.244
R6707 gnd.n2991 gnd.n1788 240.244
R6708 gnd.n3045 gnd.n1788 240.244
R6709 gnd.n3045 gnd.n1784 240.244
R6710 gnd.n3051 gnd.n1784 240.244
R6711 gnd.n3051 gnd.n1768 240.244
R6712 gnd.n3112 gnd.n1768 240.244
R6713 gnd.n3112 gnd.n1763 240.244
R6714 gnd.n3120 gnd.n1763 240.244
R6715 gnd.n3120 gnd.n1764 240.244
R6716 gnd.n1764 gnd.n1739 240.244
R6717 gnd.n3148 gnd.n1739 240.244
R6718 gnd.n3148 gnd.n1735 240.244
R6719 gnd.n3154 gnd.n1735 240.244
R6720 gnd.n3154 gnd.n1718 240.244
R6721 gnd.n3176 gnd.n1718 240.244
R6722 gnd.n3176 gnd.n1713 240.244
R6723 gnd.n3184 gnd.n1713 240.244
R6724 gnd.n3184 gnd.n1714 240.244
R6725 gnd.n1714 gnd.n1690 240.244
R6726 gnd.n3215 gnd.n1690 240.244
R6727 gnd.n3215 gnd.n1685 240.244
R6728 gnd.n3229 gnd.n1685 240.244
R6729 gnd.n3229 gnd.n1686 240.244
R6730 gnd.n3225 gnd.n1686 240.244
R6731 gnd.n3225 gnd.n1658 240.244
R6732 gnd.n3282 gnd.n1658 240.244
R6733 gnd.n3282 gnd.n1654 240.244
R6734 gnd.n3288 gnd.n1654 240.244
R6735 gnd.n3288 gnd.n1635 240.244
R6736 gnd.n3311 gnd.n1635 240.244
R6737 gnd.n3311 gnd.n1629 240.244
R6738 gnd.n3320 gnd.n1629 240.244
R6739 gnd.n3320 gnd.n1631 240.244
R6740 gnd.n1631 gnd.n1537 240.244
R6741 gnd.n3620 gnd.n1537 240.244
R6742 gnd.n3620 gnd.n1538 240.244
R6743 gnd.n3616 gnd.n1538 240.244
R6744 gnd.n3616 gnd.n3615 240.244
R6745 gnd.n3615 gnd.n1544 240.244
R6746 gnd.n3609 gnd.n1544 240.244
R6747 gnd.n3609 gnd.n1550 240.244
R6748 gnd.n3605 gnd.n1550 240.244
R6749 gnd.n3605 gnd.n1558 240.244
R6750 gnd.n3599 gnd.n1558 240.244
R6751 gnd.n3599 gnd.n1565 240.244
R6752 gnd.n3595 gnd.n1565 240.244
R6753 gnd.n3595 gnd.n1571 240.244
R6754 gnd.n3589 gnd.n1571 240.244
R6755 gnd.n3589 gnd.n1575 240.244
R6756 gnd.n3585 gnd.n1575 240.244
R6757 gnd.n3585 gnd.n1581 240.244
R6758 gnd.n3579 gnd.n1581 240.244
R6759 gnd.n3579 gnd.n1588 240.244
R6760 gnd.n3575 gnd.n1588 240.244
R6761 gnd.n3575 gnd.n1596 240.244
R6762 gnd.n1596 gnd.n1307 240.244
R6763 gnd.n4073 gnd.n1307 240.244
R6764 gnd.n4073 gnd.n1308 240.244
R6765 gnd.n4069 gnd.n1308 240.244
R6766 gnd.n4069 gnd.n1314 240.244
R6767 gnd.n4065 gnd.n1314 240.244
R6768 gnd.n4065 gnd.n1317 240.244
R6769 gnd.n4061 gnd.n1317 240.244
R6770 gnd.n4061 gnd.n1323 240.244
R6771 gnd.n1445 gnd.n1323 240.244
R6772 gnd.n1446 gnd.n1445 240.244
R6773 gnd.n1446 gnd.n1439 240.244
R6774 gnd.n3928 gnd.n1439 240.244
R6775 gnd.n3928 gnd.n1440 240.244
R6776 gnd.n3924 gnd.n1440 240.244
R6777 gnd.n3924 gnd.n1411 240.244
R6778 gnd.n3965 gnd.n1411 240.244
R6779 gnd.n3965 gnd.n1412 240.244
R6780 gnd.n3961 gnd.n1412 240.244
R6781 gnd.n3961 gnd.n3960 240.244
R6782 gnd.n3960 gnd.n1372 240.244
R6783 gnd.n4018 gnd.n1372 240.244
R6784 gnd.n4018 gnd.n1373 240.244
R6785 gnd.n4014 gnd.n1373 240.244
R6786 gnd.n4014 gnd.n4013 240.244
R6787 gnd.n4013 gnd.n4012 240.244
R6788 gnd.n4012 gnd.n1379 240.244
R6789 gnd.n1379 gnd.n334 240.244
R6790 gnd.n6641 gnd.n334 240.244
R6791 gnd.n6641 gnd.n335 240.244
R6792 gnd.n6635 gnd.n335 240.244
R6793 gnd.n6061 gnd.n676 240.244
R6794 gnd.n6061 gnd.n678 240.244
R6795 gnd.n6057 gnd.n678 240.244
R6796 gnd.n6057 gnd.n684 240.244
R6797 gnd.n6053 gnd.n684 240.244
R6798 gnd.n6053 gnd.n686 240.244
R6799 gnd.n6049 gnd.n686 240.244
R6800 gnd.n6049 gnd.n692 240.244
R6801 gnd.n6045 gnd.n692 240.244
R6802 gnd.n6045 gnd.n694 240.244
R6803 gnd.n6041 gnd.n694 240.244
R6804 gnd.n6041 gnd.n700 240.244
R6805 gnd.n6037 gnd.n700 240.244
R6806 gnd.n6037 gnd.n702 240.244
R6807 gnd.n6033 gnd.n702 240.244
R6808 gnd.n6033 gnd.n708 240.244
R6809 gnd.n6029 gnd.n708 240.244
R6810 gnd.n6029 gnd.n710 240.244
R6811 gnd.n6025 gnd.n710 240.244
R6812 gnd.n6025 gnd.n716 240.244
R6813 gnd.n6021 gnd.n716 240.244
R6814 gnd.n6021 gnd.n718 240.244
R6815 gnd.n6017 gnd.n718 240.244
R6816 gnd.n6017 gnd.n724 240.244
R6817 gnd.n6013 gnd.n724 240.244
R6818 gnd.n6013 gnd.n726 240.244
R6819 gnd.n6009 gnd.n726 240.244
R6820 gnd.n6009 gnd.n732 240.244
R6821 gnd.n6005 gnd.n732 240.244
R6822 gnd.n6005 gnd.n734 240.244
R6823 gnd.n6001 gnd.n734 240.244
R6824 gnd.n6001 gnd.n740 240.244
R6825 gnd.n5997 gnd.n740 240.244
R6826 gnd.n5997 gnd.n742 240.244
R6827 gnd.n5993 gnd.n742 240.244
R6828 gnd.n5993 gnd.n748 240.244
R6829 gnd.n5989 gnd.n748 240.244
R6830 gnd.n5989 gnd.n750 240.244
R6831 gnd.n5985 gnd.n750 240.244
R6832 gnd.n5985 gnd.n756 240.244
R6833 gnd.n5981 gnd.n756 240.244
R6834 gnd.n5981 gnd.n758 240.244
R6835 gnd.n5977 gnd.n758 240.244
R6836 gnd.n5977 gnd.n764 240.244
R6837 gnd.n5973 gnd.n764 240.244
R6838 gnd.n5973 gnd.n766 240.244
R6839 gnd.n5969 gnd.n766 240.244
R6840 gnd.n5969 gnd.n772 240.244
R6841 gnd.n5965 gnd.n772 240.244
R6842 gnd.n5965 gnd.n774 240.244
R6843 gnd.n5961 gnd.n774 240.244
R6844 gnd.n5961 gnd.n780 240.244
R6845 gnd.n5957 gnd.n780 240.244
R6846 gnd.n5957 gnd.n782 240.244
R6847 gnd.n5953 gnd.n782 240.244
R6848 gnd.n5953 gnd.n788 240.244
R6849 gnd.n5949 gnd.n788 240.244
R6850 gnd.n5949 gnd.n790 240.244
R6851 gnd.n5945 gnd.n790 240.244
R6852 gnd.n5945 gnd.n796 240.244
R6853 gnd.n5941 gnd.n796 240.244
R6854 gnd.n5941 gnd.n798 240.244
R6855 gnd.n5937 gnd.n798 240.244
R6856 gnd.n5937 gnd.n804 240.244
R6857 gnd.n5933 gnd.n804 240.244
R6858 gnd.n5933 gnd.n806 240.244
R6859 gnd.n5929 gnd.n806 240.244
R6860 gnd.n5929 gnd.n812 240.244
R6861 gnd.n5925 gnd.n812 240.244
R6862 gnd.n5925 gnd.n814 240.244
R6863 gnd.n5921 gnd.n814 240.244
R6864 gnd.n5921 gnd.n820 240.244
R6865 gnd.n5917 gnd.n820 240.244
R6866 gnd.n5917 gnd.n822 240.244
R6867 gnd.n5913 gnd.n822 240.244
R6868 gnd.n5913 gnd.n828 240.244
R6869 gnd.n5909 gnd.n828 240.244
R6870 gnd.n5909 gnd.n830 240.244
R6871 gnd.n5905 gnd.n830 240.244
R6872 gnd.n5905 gnd.n836 240.244
R6873 gnd.n5901 gnd.n836 240.244
R6874 gnd.n5901 gnd.n838 240.244
R6875 gnd.n5897 gnd.n838 240.244
R6876 gnd.n5897 gnd.n844 240.244
R6877 gnd.n1201 gnd.n1200 240.244
R6878 gnd.n1202 gnd.n1201 240.244
R6879 gnd.n1948 gnd.n1202 240.244
R6880 gnd.n1948 gnd.n1205 240.244
R6881 gnd.n1206 gnd.n1205 240.244
R6882 gnd.n1207 gnd.n1206 240.244
R6883 gnd.n1935 gnd.n1207 240.244
R6884 gnd.n1935 gnd.n1210 240.244
R6885 gnd.n1211 gnd.n1210 240.244
R6886 gnd.n1212 gnd.n1211 240.244
R6887 gnd.n1922 gnd.n1212 240.244
R6888 gnd.n1922 gnd.n1215 240.244
R6889 gnd.n1216 gnd.n1215 240.244
R6890 gnd.n1217 gnd.n1216 240.244
R6891 gnd.n1909 gnd.n1217 240.244
R6892 gnd.n1909 gnd.n1220 240.244
R6893 gnd.n1221 gnd.n1220 240.244
R6894 gnd.n1222 gnd.n1221 240.244
R6895 gnd.n1861 gnd.n1222 240.244
R6896 gnd.n1861 gnd.n1225 240.244
R6897 gnd.n1226 gnd.n1225 240.244
R6898 gnd.n1227 gnd.n1226 240.244
R6899 gnd.n1817 gnd.n1227 240.244
R6900 gnd.n1817 gnd.n1230 240.244
R6901 gnd.n1231 gnd.n1230 240.244
R6902 gnd.n1232 gnd.n1231 240.244
R6903 gnd.n3034 gnd.n1232 240.244
R6904 gnd.n3034 gnd.n1235 240.244
R6905 gnd.n1236 gnd.n1235 240.244
R6906 gnd.n1237 gnd.n1236 240.244
R6907 gnd.n1774 gnd.n1237 240.244
R6908 gnd.n1774 gnd.n1240 240.244
R6909 gnd.n1241 gnd.n1240 240.244
R6910 gnd.n1242 gnd.n1241 240.244
R6911 gnd.n3098 gnd.n1242 240.244
R6912 gnd.n3098 gnd.n1245 240.244
R6913 gnd.n1246 gnd.n1245 240.244
R6914 gnd.n1247 gnd.n1246 240.244
R6915 gnd.n3165 gnd.n1247 240.244
R6916 gnd.n3165 gnd.n1250 240.244
R6917 gnd.n1251 gnd.n1250 240.244
R6918 gnd.n1252 gnd.n1251 240.244
R6919 gnd.n3195 gnd.n1252 240.244
R6920 gnd.n3195 gnd.n1255 240.244
R6921 gnd.n1256 gnd.n1255 240.244
R6922 gnd.n1257 gnd.n1256 240.244
R6923 gnd.n1681 gnd.n1257 240.244
R6924 gnd.n1681 gnd.n1260 240.244
R6925 gnd.n1261 gnd.n1260 240.244
R6926 gnd.n1262 gnd.n1261 240.244
R6927 gnd.n3272 gnd.n1262 240.244
R6928 gnd.n3272 gnd.n1265 240.244
R6929 gnd.n1266 gnd.n1265 240.244
R6930 gnd.n1267 gnd.n1266 240.244
R6931 gnd.n1646 gnd.n1267 240.244
R6932 gnd.n1646 gnd.n1270 240.244
R6933 gnd.n1271 gnd.n1270 240.244
R6934 gnd.n1272 gnd.n1271 240.244
R6935 gnd.n3341 gnd.n1272 240.244
R6936 gnd.n3341 gnd.n1275 240.244
R6937 gnd.n1276 gnd.n1275 240.244
R6938 gnd.n1277 gnd.n1276 240.244
R6939 gnd.n1545 gnd.n1277 240.244
R6940 gnd.n1545 gnd.n1280 240.244
R6941 gnd.n1281 gnd.n1280 240.244
R6942 gnd.n1282 gnd.n1281 240.244
R6943 gnd.n1560 gnd.n1282 240.244
R6944 gnd.n1560 gnd.n1285 240.244
R6945 gnd.n1286 gnd.n1285 240.244
R6946 gnd.n1287 gnd.n1286 240.244
R6947 gnd.n3370 gnd.n1287 240.244
R6948 gnd.n3370 gnd.n1290 240.244
R6949 gnd.n1291 gnd.n1290 240.244
R6950 gnd.n1292 gnd.n1291 240.244
R6951 gnd.n1583 gnd.n1292 240.244
R6952 gnd.n1583 gnd.n1295 240.244
R6953 gnd.n1296 gnd.n1295 240.244
R6954 gnd.n1297 gnd.n1296 240.244
R6955 gnd.n1598 gnd.n1297 240.244
R6956 gnd.n1598 gnd.n1300 240.244
R6957 gnd.n1301 gnd.n1300 240.244
R6958 gnd.n4076 gnd.n1301 240.244
R6959 gnd.n1981 gnd.n1980 240.244
R6960 gnd.n1991 gnd.n1980 240.244
R6961 gnd.n1993 gnd.n1992 240.244
R6962 gnd.n2001 gnd.n2000 240.244
R6963 gnd.n2009 gnd.n2008 240.244
R6964 gnd.n2011 gnd.n2010 240.244
R6965 gnd.n2019 gnd.n2018 240.244
R6966 gnd.n2029 gnd.n2028 240.244
R6967 gnd.n2031 gnd.n2030 240.244
R6968 gnd.n2543 gnd.n2542 240.244
R6969 gnd.n2545 gnd.n2544 240.244
R6970 gnd.n2549 gnd.n2548 240.244
R6971 gnd.n2555 gnd.n2550 240.244
R6972 gnd.n2557 gnd.n2556 240.244
R6973 gnd.n2849 gnd.n1956 240.244
R6974 gnd.n2855 gnd.n1956 240.244
R6975 gnd.n2855 gnd.n1947 240.244
R6976 gnd.n2869 gnd.n1947 240.244
R6977 gnd.n2869 gnd.n1943 240.244
R6978 gnd.n2875 gnd.n1943 240.244
R6979 gnd.n2875 gnd.n1934 240.244
R6980 gnd.n2889 gnd.n1934 240.244
R6981 gnd.n2889 gnd.n1930 240.244
R6982 gnd.n2895 gnd.n1930 240.244
R6983 gnd.n2895 gnd.n1921 240.244
R6984 gnd.n2909 gnd.n1921 240.244
R6985 gnd.n2909 gnd.n1917 240.244
R6986 gnd.n2915 gnd.n1917 240.244
R6987 gnd.n2915 gnd.n1908 240.244
R6988 gnd.n2929 gnd.n1908 240.244
R6989 gnd.n2929 gnd.n1902 240.244
R6990 gnd.n2953 gnd.n1902 240.244
R6991 gnd.n2953 gnd.n1903 240.244
R6992 gnd.n2934 gnd.n1903 240.244
R6993 gnd.n2935 gnd.n2934 240.244
R6994 gnd.n2936 gnd.n2935 240.244
R6995 gnd.n2939 gnd.n2936 240.244
R6996 gnd.n2941 gnd.n2939 240.244
R6997 gnd.n2941 gnd.n1805 240.244
R6998 gnd.n3012 gnd.n1805 240.244
R6999 gnd.n3012 gnd.n1797 240.244
R7000 gnd.n1797 gnd.n1789 240.244
R7001 gnd.n3025 gnd.n1789 240.244
R7002 gnd.n3025 gnd.n1800 240.244
R7003 gnd.n3018 gnd.n1800 240.244
R7004 gnd.n3018 gnd.n1770 240.244
R7005 gnd.n1770 gnd.n1754 240.244
R7006 gnd.n3131 gnd.n1754 240.244
R7007 gnd.n3131 gnd.n1748 240.244
R7008 gnd.n3138 gnd.n1748 240.244
R7009 gnd.n3138 gnd.n1749 240.244
R7010 gnd.n1749 gnd.n1725 240.244
R7011 gnd.n3167 gnd.n1725 240.244
R7012 gnd.n3167 gnd.n1721 240.244
R7013 gnd.n3173 gnd.n1721 240.244
R7014 gnd.n3173 gnd.n1705 240.244
R7015 gnd.n3197 gnd.n1705 240.244
R7016 gnd.n3197 gnd.n1699 240.244
R7017 gnd.n3204 gnd.n1699 240.244
R7018 gnd.n3204 gnd.n1700 240.244
R7019 gnd.n1700 gnd.n1674 240.244
R7020 gnd.n3240 gnd.n1674 240.244
R7021 gnd.n3240 gnd.n1669 240.244
R7022 gnd.n3250 gnd.n1669 240.244
R7023 gnd.n3250 gnd.n1666 240.244
R7024 gnd.n3244 gnd.n1666 240.244
R7025 gnd.n3244 gnd.n1643 240.244
R7026 gnd.n3300 gnd.n1643 240.244
R7027 gnd.n3300 gnd.n1638 240.244
R7028 gnd.n3307 gnd.n1638 240.244
R7029 gnd.n3307 gnd.n1628 240.244
R7030 gnd.n1628 gnd.n1617 240.244
R7031 gnd.n3343 gnd.n1617 240.244
R7032 gnd.n3343 gnd.n1613 240.244
R7033 gnd.n3350 gnd.n1613 240.244
R7034 gnd.n3352 gnd.n3350 240.244
R7035 gnd.n3353 gnd.n3352 240.244
R7036 gnd.n3353 gnd.n1547 240.244
R7037 gnd.n1548 gnd.n1547 240.244
R7038 gnd.n3360 gnd.n1548 240.244
R7039 gnd.n3361 gnd.n3360 240.244
R7040 gnd.n3361 gnd.n1562 240.244
R7041 gnd.n1563 gnd.n1562 240.244
R7042 gnd.n3368 gnd.n1563 240.244
R7043 gnd.n3372 gnd.n3368 240.244
R7044 gnd.n3372 gnd.n1572 240.244
R7045 gnd.n1573 gnd.n1572 240.244
R7046 gnd.n3379 gnd.n1573 240.244
R7047 gnd.n3380 gnd.n3379 240.244
R7048 gnd.n3380 gnd.n1585 240.244
R7049 gnd.n1586 gnd.n1585 240.244
R7050 gnd.n3387 gnd.n1586 240.244
R7051 gnd.n3388 gnd.n3387 240.244
R7052 gnd.n3388 gnd.n1600 240.244
R7053 gnd.n3570 gnd.n1600 240.244
R7054 gnd.n3570 gnd.n1305 240.244
R7055 gnd.n3461 gnd.n3460 240.244
R7056 gnd.n3464 gnd.n3463 240.244
R7057 gnd.n3480 gnd.n3479 240.244
R7058 gnd.n3483 gnd.n3482 240.244
R7059 gnd.n3499 gnd.n3498 240.244
R7060 gnd.n3502 gnd.n3501 240.244
R7061 gnd.n3518 gnd.n3517 240.244
R7062 gnd.n3522 gnd.n3520 240.244
R7063 gnd.n3538 gnd.n3402 240.244
R7064 gnd.n3542 gnd.n3540 240.244
R7065 gnd.n3548 gnd.n3398 240.244
R7066 gnd.n3552 gnd.n3550 240.244
R7067 gnd.n3561 gnd.n3394 240.244
R7068 gnd.n3564 gnd.n3563 240.244
R7069 gnd.n1845 gnd.n1844 240.132
R7070 gnd.n3637 gnd.n3636 240.132
R7071 gnd.n6064 gnd.n672 225.874
R7072 gnd.n6072 gnd.n672 225.874
R7073 gnd.n6073 gnd.n6072 225.874
R7074 gnd.n6074 gnd.n6073 225.874
R7075 gnd.n6074 gnd.n666 225.874
R7076 gnd.n6082 gnd.n666 225.874
R7077 gnd.n6083 gnd.n6082 225.874
R7078 gnd.n6084 gnd.n6083 225.874
R7079 gnd.n6084 gnd.n660 225.874
R7080 gnd.n6092 gnd.n660 225.874
R7081 gnd.n6093 gnd.n6092 225.874
R7082 gnd.n6094 gnd.n6093 225.874
R7083 gnd.n6094 gnd.n654 225.874
R7084 gnd.n6102 gnd.n654 225.874
R7085 gnd.n6103 gnd.n6102 225.874
R7086 gnd.n6104 gnd.n6103 225.874
R7087 gnd.n6104 gnd.n648 225.874
R7088 gnd.n6112 gnd.n648 225.874
R7089 gnd.n6113 gnd.n6112 225.874
R7090 gnd.n6114 gnd.n6113 225.874
R7091 gnd.n6114 gnd.n642 225.874
R7092 gnd.n6122 gnd.n642 225.874
R7093 gnd.n6123 gnd.n6122 225.874
R7094 gnd.n6124 gnd.n6123 225.874
R7095 gnd.n6124 gnd.n636 225.874
R7096 gnd.n6132 gnd.n636 225.874
R7097 gnd.n6133 gnd.n6132 225.874
R7098 gnd.n6134 gnd.n6133 225.874
R7099 gnd.n6134 gnd.n630 225.874
R7100 gnd.n6142 gnd.n630 225.874
R7101 gnd.n6143 gnd.n6142 225.874
R7102 gnd.n6144 gnd.n6143 225.874
R7103 gnd.n6144 gnd.n624 225.874
R7104 gnd.n6152 gnd.n624 225.874
R7105 gnd.n6153 gnd.n6152 225.874
R7106 gnd.n6154 gnd.n6153 225.874
R7107 gnd.n6154 gnd.n618 225.874
R7108 gnd.n6162 gnd.n618 225.874
R7109 gnd.n6163 gnd.n6162 225.874
R7110 gnd.n6164 gnd.n6163 225.874
R7111 gnd.n6164 gnd.n612 225.874
R7112 gnd.n6172 gnd.n612 225.874
R7113 gnd.n6173 gnd.n6172 225.874
R7114 gnd.n6174 gnd.n6173 225.874
R7115 gnd.n6174 gnd.n606 225.874
R7116 gnd.n6182 gnd.n606 225.874
R7117 gnd.n6183 gnd.n6182 225.874
R7118 gnd.n6184 gnd.n6183 225.874
R7119 gnd.n6184 gnd.n600 225.874
R7120 gnd.n6192 gnd.n600 225.874
R7121 gnd.n6193 gnd.n6192 225.874
R7122 gnd.n6194 gnd.n6193 225.874
R7123 gnd.n6194 gnd.n594 225.874
R7124 gnd.n6202 gnd.n594 225.874
R7125 gnd.n6203 gnd.n6202 225.874
R7126 gnd.n6204 gnd.n6203 225.874
R7127 gnd.n6204 gnd.n588 225.874
R7128 gnd.n6212 gnd.n588 225.874
R7129 gnd.n6213 gnd.n6212 225.874
R7130 gnd.n6214 gnd.n6213 225.874
R7131 gnd.n6214 gnd.n582 225.874
R7132 gnd.n6222 gnd.n582 225.874
R7133 gnd.n6223 gnd.n6222 225.874
R7134 gnd.n6224 gnd.n6223 225.874
R7135 gnd.n6224 gnd.n576 225.874
R7136 gnd.n6232 gnd.n576 225.874
R7137 gnd.n6233 gnd.n6232 225.874
R7138 gnd.n6234 gnd.n6233 225.874
R7139 gnd.n6234 gnd.n570 225.874
R7140 gnd.n6242 gnd.n570 225.874
R7141 gnd.n6243 gnd.n6242 225.874
R7142 gnd.n6244 gnd.n6243 225.874
R7143 gnd.n6244 gnd.n564 225.874
R7144 gnd.n6252 gnd.n564 225.874
R7145 gnd.n6253 gnd.n6252 225.874
R7146 gnd.n6254 gnd.n6253 225.874
R7147 gnd.n6254 gnd.n558 225.874
R7148 gnd.n6262 gnd.n558 225.874
R7149 gnd.n6263 gnd.n6262 225.874
R7150 gnd.n6264 gnd.n6263 225.874
R7151 gnd.n6264 gnd.n552 225.874
R7152 gnd.n6272 gnd.n552 225.874
R7153 gnd.n6273 gnd.n6272 225.874
R7154 gnd.n6274 gnd.n6273 225.874
R7155 gnd.n6274 gnd.n546 225.874
R7156 gnd.n6282 gnd.n546 225.874
R7157 gnd.n6283 gnd.n6282 225.874
R7158 gnd.n6284 gnd.n6283 225.874
R7159 gnd.n6284 gnd.n540 225.874
R7160 gnd.n6292 gnd.n540 225.874
R7161 gnd.n6293 gnd.n6292 225.874
R7162 gnd.n6294 gnd.n6293 225.874
R7163 gnd.n6294 gnd.n534 225.874
R7164 gnd.n6302 gnd.n534 225.874
R7165 gnd.n6303 gnd.n6302 225.874
R7166 gnd.n6304 gnd.n6303 225.874
R7167 gnd.n6304 gnd.n528 225.874
R7168 gnd.n6312 gnd.n528 225.874
R7169 gnd.n6313 gnd.n6312 225.874
R7170 gnd.n6314 gnd.n6313 225.874
R7171 gnd.n6314 gnd.n522 225.874
R7172 gnd.n6322 gnd.n522 225.874
R7173 gnd.n6323 gnd.n6322 225.874
R7174 gnd.n6324 gnd.n6323 225.874
R7175 gnd.n6324 gnd.n516 225.874
R7176 gnd.n6332 gnd.n516 225.874
R7177 gnd.n6333 gnd.n6332 225.874
R7178 gnd.n6334 gnd.n6333 225.874
R7179 gnd.n6334 gnd.n510 225.874
R7180 gnd.n6342 gnd.n510 225.874
R7181 gnd.n6343 gnd.n6342 225.874
R7182 gnd.n6344 gnd.n6343 225.874
R7183 gnd.n6344 gnd.n504 225.874
R7184 gnd.n6352 gnd.n504 225.874
R7185 gnd.n6353 gnd.n6352 225.874
R7186 gnd.n6354 gnd.n6353 225.874
R7187 gnd.n6354 gnd.n498 225.874
R7188 gnd.n6362 gnd.n498 225.874
R7189 gnd.n6363 gnd.n6362 225.874
R7190 gnd.n6364 gnd.n6363 225.874
R7191 gnd.n6364 gnd.n492 225.874
R7192 gnd.n6372 gnd.n492 225.874
R7193 gnd.n6373 gnd.n6372 225.874
R7194 gnd.n6374 gnd.n6373 225.874
R7195 gnd.n6374 gnd.n486 225.874
R7196 gnd.n6382 gnd.n486 225.874
R7197 gnd.n6383 gnd.n6382 225.874
R7198 gnd.n6384 gnd.n6383 225.874
R7199 gnd.n6384 gnd.n480 225.874
R7200 gnd.n6392 gnd.n480 225.874
R7201 gnd.n6393 gnd.n6392 225.874
R7202 gnd.n6394 gnd.n6393 225.874
R7203 gnd.n6394 gnd.n474 225.874
R7204 gnd.n6402 gnd.n474 225.874
R7205 gnd.n6403 gnd.n6402 225.874
R7206 gnd.n6404 gnd.n6403 225.874
R7207 gnd.n6404 gnd.n468 225.874
R7208 gnd.n6413 gnd.n468 225.874
R7209 gnd.n6414 gnd.n6413 225.874
R7210 gnd.n6415 gnd.n6414 225.874
R7211 gnd.n6415 gnd.n463 225.874
R7212 gnd.n5137 gnd.t79 224.174
R7213 gnd.n4518 gnd.t125 224.174
R7214 gnd.n3837 gnd.n3836 199.319
R7215 gnd.n3837 gnd.n3783 199.319
R7216 gnd.n2093 gnd.n2063 199.319
R7217 gnd.n2093 gnd.n2062 199.319
R7218 gnd.n1846 gnd.n1843 186.49
R7219 gnd.n3638 gnd.n3635 186.49
R7220 gnd.n4786 gnd.n4785 185
R7221 gnd.n4784 gnd.n4783 185
R7222 gnd.n4763 gnd.n4762 185
R7223 gnd.n4778 gnd.n4777 185
R7224 gnd.n4776 gnd.n4775 185
R7225 gnd.n4767 gnd.n4766 185
R7226 gnd.n4770 gnd.n4769 185
R7227 gnd.n4754 gnd.n4753 185
R7228 gnd.n4752 gnd.n4751 185
R7229 gnd.n4731 gnd.n4730 185
R7230 gnd.n4746 gnd.n4745 185
R7231 gnd.n4744 gnd.n4743 185
R7232 gnd.n4735 gnd.n4734 185
R7233 gnd.n4738 gnd.n4737 185
R7234 gnd.n4722 gnd.n4721 185
R7235 gnd.n4720 gnd.n4719 185
R7236 gnd.n4699 gnd.n4698 185
R7237 gnd.n4714 gnd.n4713 185
R7238 gnd.n4712 gnd.n4711 185
R7239 gnd.n4703 gnd.n4702 185
R7240 gnd.n4706 gnd.n4705 185
R7241 gnd.n4691 gnd.n4690 185
R7242 gnd.n4689 gnd.n4688 185
R7243 gnd.n4668 gnd.n4667 185
R7244 gnd.n4683 gnd.n4682 185
R7245 gnd.n4681 gnd.n4680 185
R7246 gnd.n4672 gnd.n4671 185
R7247 gnd.n4675 gnd.n4674 185
R7248 gnd.n4659 gnd.n4658 185
R7249 gnd.n4657 gnd.n4656 185
R7250 gnd.n4636 gnd.n4635 185
R7251 gnd.n4651 gnd.n4650 185
R7252 gnd.n4649 gnd.n4648 185
R7253 gnd.n4640 gnd.n4639 185
R7254 gnd.n4643 gnd.n4642 185
R7255 gnd.n4627 gnd.n4626 185
R7256 gnd.n4625 gnd.n4624 185
R7257 gnd.n4604 gnd.n4603 185
R7258 gnd.n4619 gnd.n4618 185
R7259 gnd.n4617 gnd.n4616 185
R7260 gnd.n4608 gnd.n4607 185
R7261 gnd.n4611 gnd.n4610 185
R7262 gnd.n4595 gnd.n4594 185
R7263 gnd.n4593 gnd.n4592 185
R7264 gnd.n4572 gnd.n4571 185
R7265 gnd.n4587 gnd.n4586 185
R7266 gnd.n4585 gnd.n4584 185
R7267 gnd.n4576 gnd.n4575 185
R7268 gnd.n4579 gnd.n4578 185
R7269 gnd.n4564 gnd.n4563 185
R7270 gnd.n4562 gnd.n4561 185
R7271 gnd.n4541 gnd.n4540 185
R7272 gnd.n4556 gnd.n4555 185
R7273 gnd.n4554 gnd.n4553 185
R7274 gnd.n4545 gnd.n4544 185
R7275 gnd.n4548 gnd.n4547 185
R7276 gnd.n5138 gnd.t78 178.987
R7277 gnd.n4519 gnd.t126 178.987
R7278 gnd.n1 gnd.t146 170.774
R7279 gnd.n7 gnd.t5 170.103
R7280 gnd.n6 gnd.t21 170.103
R7281 gnd.n5 gnd.t23 170.103
R7282 gnd.n4 gnd.t150 170.103
R7283 gnd.n3 gnd.t7 170.103
R7284 gnd.n2 gnd.t28 170.103
R7285 gnd.n1 gnd.t308 170.103
R7286 gnd.n3706 gnd.n3705 163.367
R7287 gnd.n3702 gnd.n3701 163.367
R7288 gnd.n3698 gnd.n3697 163.367
R7289 gnd.n3694 gnd.n3693 163.367
R7290 gnd.n3690 gnd.n3689 163.367
R7291 gnd.n3686 gnd.n3685 163.367
R7292 gnd.n3682 gnd.n3681 163.367
R7293 gnd.n3678 gnd.n3677 163.367
R7294 gnd.n3674 gnd.n3673 163.367
R7295 gnd.n3670 gnd.n3669 163.367
R7296 gnd.n3666 gnd.n3665 163.367
R7297 gnd.n3662 gnd.n3661 163.367
R7298 gnd.n3658 gnd.n3657 163.367
R7299 gnd.n3654 gnd.n3653 163.367
R7300 gnd.n3649 gnd.n3648 163.367
R7301 gnd.n3781 gnd.n1491 163.367
R7302 gnd.n3778 gnd.n3777 163.367
R7303 gnd.n3775 gnd.n1524 163.367
R7304 gnd.n3770 gnd.n3769 163.367
R7305 gnd.n3766 gnd.n3765 163.367
R7306 gnd.n3762 gnd.n3761 163.367
R7307 gnd.n3758 gnd.n3757 163.367
R7308 gnd.n3754 gnd.n3753 163.367
R7309 gnd.n3750 gnd.n3749 163.367
R7310 gnd.n3746 gnd.n3745 163.367
R7311 gnd.n3742 gnd.n3741 163.367
R7312 gnd.n3738 gnd.n3737 163.367
R7313 gnd.n3734 gnd.n3733 163.367
R7314 gnd.n3730 gnd.n3729 163.367
R7315 gnd.n3726 gnd.n3725 163.367
R7316 gnd.n3722 gnd.n3721 163.367
R7317 gnd.n3718 gnd.n3717 163.367
R7318 gnd.n2976 gnd.n1829 163.367
R7319 gnd.n2982 gnd.n1829 163.367
R7320 gnd.n2982 gnd.n1832 163.367
R7321 gnd.n1832 gnd.n1819 163.367
R7322 gnd.n1819 gnd.n1809 163.367
R7323 gnd.n3005 gnd.n1809 163.367
R7324 gnd.n3005 gnd.n1807 163.367
R7325 gnd.n3009 gnd.n1807 163.367
R7326 gnd.n3009 gnd.n1796 163.367
R7327 gnd.n3032 gnd.n1796 163.367
R7328 gnd.n3032 gnd.n1790 163.367
R7329 gnd.n3028 gnd.n1790 163.367
R7330 gnd.n3028 gnd.n1780 163.367
R7331 gnd.n1780 gnd.n1773 163.367
R7332 gnd.n3061 gnd.n1773 163.367
R7333 gnd.n3061 gnd.n1771 163.367
R7334 gnd.n3108 gnd.n1771 163.367
R7335 gnd.n3108 gnd.n1762 163.367
R7336 gnd.n3104 gnd.n1762 163.367
R7337 gnd.n3104 gnd.n1756 163.367
R7338 gnd.n3101 gnd.n1756 163.367
R7339 gnd.n3101 gnd.n1747 163.367
R7340 gnd.n3095 gnd.n1747 163.367
R7341 gnd.n3095 gnd.n1741 163.367
R7342 gnd.n3092 gnd.n1741 163.367
R7343 gnd.n3092 gnd.n1734 163.367
R7344 gnd.n3087 gnd.n1734 163.367
R7345 gnd.n3087 gnd.n1727 163.367
R7346 gnd.n3084 gnd.n1727 163.367
R7347 gnd.n3084 gnd.n1720 163.367
R7348 gnd.n1720 gnd.n1711 163.367
R7349 gnd.n1712 gnd.n1711 163.367
R7350 gnd.n1712 gnd.n1706 163.367
R7351 gnd.n3078 gnd.n1706 163.367
R7352 gnd.n3078 gnd.n1698 163.367
R7353 gnd.n3073 gnd.n1698 163.367
R7354 gnd.n3073 gnd.n1692 163.367
R7355 gnd.n3070 gnd.n1692 163.367
R7356 gnd.n3070 gnd.n1683 163.367
R7357 gnd.n3065 gnd.n1683 163.367
R7358 gnd.n3065 gnd.n1675 163.367
R7359 gnd.n1675 gnd.n1668 163.367
R7360 gnd.n3253 gnd.n1668 163.367
R7361 gnd.n3253 gnd.n1665 163.367
R7362 gnd.n3270 gnd.n1665 163.367
R7363 gnd.n3270 gnd.n1659 163.367
R7364 gnd.n3266 gnd.n1659 163.367
R7365 gnd.n3266 gnd.n1653 163.367
R7366 gnd.n3261 gnd.n1653 163.367
R7367 gnd.n3261 gnd.n1645 163.367
R7368 gnd.n3258 gnd.n1645 163.367
R7369 gnd.n3258 gnd.n1637 163.367
R7370 gnd.n1637 gnd.n1627 163.367
R7371 gnd.n1627 gnd.n1621 163.367
R7372 gnd.n3332 gnd.n1621 163.367
R7373 gnd.n3332 gnd.n1619 163.367
R7374 gnd.n3338 gnd.n1619 163.367
R7375 gnd.n3338 gnd.n1535 163.367
R7376 gnd.n1535 gnd.n1528 163.367
R7377 gnd.n3713 gnd.n1528 163.367
R7378 gnd.n2967 gnd.n1860 163.367
R7379 gnd.n2696 gnd.n1860 163.367
R7380 gnd.n2700 gnd.n2699 163.367
R7381 gnd.n2704 gnd.n2703 163.367
R7382 gnd.n2708 gnd.n2707 163.367
R7383 gnd.n2712 gnd.n2711 163.367
R7384 gnd.n2716 gnd.n2715 163.367
R7385 gnd.n2720 gnd.n2719 163.367
R7386 gnd.n2724 gnd.n2723 163.367
R7387 gnd.n2728 gnd.n2727 163.367
R7388 gnd.n2732 gnd.n2731 163.367
R7389 gnd.n2736 gnd.n2735 163.367
R7390 gnd.n2740 gnd.n2739 163.367
R7391 gnd.n2744 gnd.n2743 163.367
R7392 gnd.n2748 gnd.n2747 163.367
R7393 gnd.n2752 gnd.n2751 163.367
R7394 gnd.n2756 gnd.n2755 163.367
R7395 gnd.n2690 gnd.n2689 163.367
R7396 gnd.n2685 gnd.n2684 163.367
R7397 gnd.n2681 gnd.n2680 163.367
R7398 gnd.n2677 gnd.n2676 163.367
R7399 gnd.n2673 gnd.n2672 163.367
R7400 gnd.n2669 gnd.n2668 163.367
R7401 gnd.n2665 gnd.n2664 163.367
R7402 gnd.n2661 gnd.n2660 163.367
R7403 gnd.n2657 gnd.n2656 163.367
R7404 gnd.n2653 gnd.n2652 163.367
R7405 gnd.n2649 gnd.n2648 163.367
R7406 gnd.n2645 gnd.n2644 163.367
R7407 gnd.n2641 gnd.n2640 163.367
R7408 gnd.n2637 gnd.n2636 163.367
R7409 gnd.n2633 gnd.n2632 163.367
R7410 gnd.n2974 gnd.n1838 163.367
R7411 gnd.n1838 gnd.n1827 163.367
R7412 gnd.n1827 gnd.n1816 163.367
R7413 gnd.n2998 gnd.n1816 163.367
R7414 gnd.n2998 gnd.n1811 163.367
R7415 gnd.n3003 gnd.n1811 163.367
R7416 gnd.n3003 gnd.n1814 163.367
R7417 gnd.n1814 gnd.n1794 163.367
R7418 gnd.n3037 gnd.n1794 163.367
R7419 gnd.n3037 gnd.n1792 163.367
R7420 gnd.n3041 gnd.n1792 163.367
R7421 gnd.n3041 gnd.n1779 163.367
R7422 gnd.n3054 gnd.n1779 163.367
R7423 gnd.n3054 gnd.n1776 163.367
R7424 gnd.n3059 gnd.n1776 163.367
R7425 gnd.n3059 gnd.n1777 163.367
R7426 gnd.n1777 gnd.n1760 163.367
R7427 gnd.n3124 gnd.n1760 163.367
R7428 gnd.n3124 gnd.n1758 163.367
R7429 gnd.n3128 gnd.n1758 163.367
R7430 gnd.n3128 gnd.n1745 163.367
R7431 gnd.n3141 gnd.n1745 163.367
R7432 gnd.n3141 gnd.n1743 163.367
R7433 gnd.n3145 gnd.n1743 163.367
R7434 gnd.n3145 gnd.n1732 163.367
R7435 gnd.n3157 gnd.n1732 163.367
R7436 gnd.n3157 gnd.n1729 163.367
R7437 gnd.n3162 gnd.n1729 163.367
R7438 gnd.n3162 gnd.n1730 163.367
R7439 gnd.n1730 gnd.n1709 163.367
R7440 gnd.n3189 gnd.n1709 163.367
R7441 gnd.n3189 gnd.n1707 163.367
R7442 gnd.n3193 gnd.n1707 163.367
R7443 gnd.n3193 gnd.n1696 163.367
R7444 gnd.n3208 gnd.n1696 163.367
R7445 gnd.n3208 gnd.n1694 163.367
R7446 gnd.n3212 gnd.n1694 163.367
R7447 gnd.n3212 gnd.n1680 163.367
R7448 gnd.n3232 gnd.n1680 163.367
R7449 gnd.n3232 gnd.n1677 163.367
R7450 gnd.n3237 gnd.n1677 163.367
R7451 gnd.n3237 gnd.n1678 163.367
R7452 gnd.n1678 gnd.n1663 163.367
R7453 gnd.n3275 gnd.n1663 163.367
R7454 gnd.n3275 gnd.n1661 163.367
R7455 gnd.n3279 gnd.n1661 163.367
R7456 gnd.n3279 gnd.n1651 163.367
R7457 gnd.n3291 gnd.n1651 163.367
R7458 gnd.n3291 gnd.n1648 163.367
R7459 gnd.n3296 gnd.n1648 163.367
R7460 gnd.n3296 gnd.n1649 163.367
R7461 gnd.n1649 gnd.n1625 163.367
R7462 gnd.n3325 gnd.n1625 163.367
R7463 gnd.n3325 gnd.n1622 163.367
R7464 gnd.n3330 gnd.n1622 163.367
R7465 gnd.n3330 gnd.n1623 163.367
R7466 gnd.n1623 gnd.n1533 163.367
R7467 gnd.n3623 gnd.n1533 163.367
R7468 gnd.n3623 gnd.n1530 163.367
R7469 gnd.n3711 gnd.n1530 163.367
R7470 gnd.n3644 gnd.n3643 156.462
R7471 gnd.n3840 gnd.n3782 154.689
R7472 gnd.n2758 gnd.n2757 154.689
R7473 gnd.n4726 gnd.n4694 153.042
R7474 gnd.n4790 gnd.n4789 152.079
R7475 gnd.n4758 gnd.n4757 152.079
R7476 gnd.n4726 gnd.n4725 152.079
R7477 gnd.n1851 gnd.n1850 152
R7478 gnd.n1852 gnd.n1841 152
R7479 gnd.n1854 gnd.n1853 152
R7480 gnd.n1856 gnd.n1839 152
R7481 gnd.n1858 gnd.n1857 152
R7482 gnd.n3642 gnd.n3626 152
R7483 gnd.n3634 gnd.n3627 152
R7484 gnd.n3633 gnd.n3632 152
R7485 gnd.n3631 gnd.n3628 152
R7486 gnd.n3629 gnd.t103 150.546
R7487 gnd.t19 gnd.n4768 147.661
R7488 gnd.t314 gnd.n4736 147.661
R7489 gnd.t156 gnd.n4704 147.661
R7490 gnd.t148 gnd.n4673 147.661
R7491 gnd.t16 gnd.n4641 147.661
R7492 gnd.t306 gnd.n4609 147.661
R7493 gnd.t310 gnd.n4577 147.661
R7494 gnd.t32 gnd.n4546 147.661
R7495 gnd.n3780 gnd.n1490 143.351
R7496 gnd.n2754 gnd.n1877 143.351
R7497 gnd.n2754 gnd.n1878 143.351
R7498 gnd.n1848 gnd.t136 130.484
R7499 gnd.n1857 gnd.t133 126.766
R7500 gnd.n1855 gnd.t120 126.766
R7501 gnd.n1841 gnd.t41 126.766
R7502 gnd.n1849 gnd.t100 126.766
R7503 gnd.n3630 gnd.t38 126.766
R7504 gnd.n3632 gnd.t117 126.766
R7505 gnd.n3641 gnd.t130 126.766
R7506 gnd.n3643 gnd.t88 126.766
R7507 gnd.n4785 gnd.n4784 104.615
R7508 gnd.n4784 gnd.n4762 104.615
R7509 gnd.n4777 gnd.n4762 104.615
R7510 gnd.n4777 gnd.n4776 104.615
R7511 gnd.n4776 gnd.n4766 104.615
R7512 gnd.n4769 gnd.n4766 104.615
R7513 gnd.n4753 gnd.n4752 104.615
R7514 gnd.n4752 gnd.n4730 104.615
R7515 gnd.n4745 gnd.n4730 104.615
R7516 gnd.n4745 gnd.n4744 104.615
R7517 gnd.n4744 gnd.n4734 104.615
R7518 gnd.n4737 gnd.n4734 104.615
R7519 gnd.n4721 gnd.n4720 104.615
R7520 gnd.n4720 gnd.n4698 104.615
R7521 gnd.n4713 gnd.n4698 104.615
R7522 gnd.n4713 gnd.n4712 104.615
R7523 gnd.n4712 gnd.n4702 104.615
R7524 gnd.n4705 gnd.n4702 104.615
R7525 gnd.n4690 gnd.n4689 104.615
R7526 gnd.n4689 gnd.n4667 104.615
R7527 gnd.n4682 gnd.n4667 104.615
R7528 gnd.n4682 gnd.n4681 104.615
R7529 gnd.n4681 gnd.n4671 104.615
R7530 gnd.n4674 gnd.n4671 104.615
R7531 gnd.n4658 gnd.n4657 104.615
R7532 gnd.n4657 gnd.n4635 104.615
R7533 gnd.n4650 gnd.n4635 104.615
R7534 gnd.n4650 gnd.n4649 104.615
R7535 gnd.n4649 gnd.n4639 104.615
R7536 gnd.n4642 gnd.n4639 104.615
R7537 gnd.n4626 gnd.n4625 104.615
R7538 gnd.n4625 gnd.n4603 104.615
R7539 gnd.n4618 gnd.n4603 104.615
R7540 gnd.n4618 gnd.n4617 104.615
R7541 gnd.n4617 gnd.n4607 104.615
R7542 gnd.n4610 gnd.n4607 104.615
R7543 gnd.n4594 gnd.n4593 104.615
R7544 gnd.n4593 gnd.n4571 104.615
R7545 gnd.n4586 gnd.n4571 104.615
R7546 gnd.n4586 gnd.n4585 104.615
R7547 gnd.n4585 gnd.n4575 104.615
R7548 gnd.n4578 gnd.n4575 104.615
R7549 gnd.n4563 gnd.n4562 104.615
R7550 gnd.n4562 gnd.n4540 104.615
R7551 gnd.n4555 gnd.n4540 104.615
R7552 gnd.n4555 gnd.n4554 104.615
R7553 gnd.n4554 gnd.n4544 104.615
R7554 gnd.n4547 gnd.n4544 104.615
R7555 gnd.n5400 gnd.t69 100.632
R7556 gnd.n4474 gnd.t111 100.632
R7557 gnd.n7006 gnd.n112 99.6594
R7558 gnd.n7004 gnd.n7003 99.6594
R7559 gnd.n6999 gnd.n119 99.6594
R7560 gnd.n6997 gnd.n6996 99.6594
R7561 gnd.n6992 gnd.n126 99.6594
R7562 gnd.n6990 gnd.n6989 99.6594
R7563 gnd.n6985 gnd.n133 99.6594
R7564 gnd.n6983 gnd.n6982 99.6594
R7565 gnd.n6975 gnd.n140 99.6594
R7566 gnd.n6973 gnd.n6972 99.6594
R7567 gnd.n6968 gnd.n147 99.6594
R7568 gnd.n6966 gnd.n6965 99.6594
R7569 gnd.n6961 gnd.n154 99.6594
R7570 gnd.n6959 gnd.n6958 99.6594
R7571 gnd.n6954 gnd.n161 99.6594
R7572 gnd.n6952 gnd.n6951 99.6594
R7573 gnd.n6947 gnd.n168 99.6594
R7574 gnd.n6945 gnd.n6944 99.6594
R7575 gnd.n173 gnd.n172 99.6594
R7576 gnd.n3801 gnd.n1329 99.6594
R7577 gnd.n3805 gnd.n3804 99.6594
R7578 gnd.n3812 gnd.n3811 99.6594
R7579 gnd.n3815 gnd.n3814 99.6594
R7580 gnd.n3822 gnd.n3821 99.6594
R7581 gnd.n3825 gnd.n3824 99.6594
R7582 gnd.n3833 gnd.n3832 99.6594
R7583 gnd.n3836 gnd.n3835 99.6594
R7584 gnd.n3846 gnd.n3845 99.6594
R7585 gnd.n3849 gnd.n3848 99.6594
R7586 gnd.n3856 gnd.n3855 99.6594
R7587 gnd.n3859 gnd.n3858 99.6594
R7588 gnd.n3866 gnd.n3865 99.6594
R7589 gnd.n3869 gnd.n3868 99.6594
R7590 gnd.n3876 gnd.n3875 99.6594
R7591 gnd.n3879 gnd.n3878 99.6594
R7592 gnd.n3887 gnd.n3886 99.6594
R7593 gnd.n3890 gnd.n3889 99.6594
R7594 gnd.n2786 gnd.n2785 99.6594
R7595 gnd.n2781 gnd.n2069 99.6594
R7596 gnd.n2777 gnd.n2068 99.6594
R7597 gnd.n2773 gnd.n2067 99.6594
R7598 gnd.n2769 gnd.n2066 99.6594
R7599 gnd.n2765 gnd.n2065 99.6594
R7600 gnd.n2761 gnd.n2064 99.6594
R7601 gnd.n2623 gnd.n2062 99.6594
R7602 gnd.n2621 gnd.n2061 99.6594
R7603 gnd.n2617 gnd.n2060 99.6594
R7604 gnd.n2613 gnd.n2059 99.6594
R7605 gnd.n2609 gnd.n2058 99.6594
R7606 gnd.n2605 gnd.n2057 99.6594
R7607 gnd.n2601 gnd.n2056 99.6594
R7608 gnd.n2597 gnd.n2055 99.6594
R7609 gnd.n2593 gnd.n2054 99.6594
R7610 gnd.n2589 gnd.n2053 99.6594
R7611 gnd.n2111 gnd.n2052 99.6594
R7612 gnd.n4443 gnd.n4442 99.6594
R7613 gnd.n4437 gnd.n857 99.6594
R7614 gnd.n4434 gnd.n858 99.6594
R7615 gnd.n4430 gnd.n859 99.6594
R7616 gnd.n4426 gnd.n860 99.6594
R7617 gnd.n4422 gnd.n861 99.6594
R7618 gnd.n4418 gnd.n862 99.6594
R7619 gnd.n4414 gnd.n863 99.6594
R7620 gnd.n4410 gnd.n864 99.6594
R7621 gnd.n4405 gnd.n865 99.6594
R7622 gnd.n4401 gnd.n866 99.6594
R7623 gnd.n4397 gnd.n867 99.6594
R7624 gnd.n4393 gnd.n868 99.6594
R7625 gnd.n4389 gnd.n869 99.6594
R7626 gnd.n4385 gnd.n870 99.6594
R7627 gnd.n4381 gnd.n871 99.6594
R7628 gnd.n4377 gnd.n872 99.6594
R7629 gnd.n4373 gnd.n873 99.6594
R7630 gnd.n928 gnd.n874 99.6594
R7631 gnd.n5879 gnd.n4454 99.6594
R7632 gnd.n5877 gnd.n5876 99.6594
R7633 gnd.n5872 gnd.n4461 99.6594
R7634 gnd.n5870 gnd.n5869 99.6594
R7635 gnd.n5865 gnd.n4468 99.6594
R7636 gnd.n5863 gnd.n5862 99.6594
R7637 gnd.n5858 gnd.n4477 99.6594
R7638 gnd.n5856 gnd.n5855 99.6594
R7639 gnd.n5433 gnd.n5432 99.6594
R7640 gnd.n5427 gnd.n5375 99.6594
R7641 gnd.n5424 gnd.n5376 99.6594
R7642 gnd.n5420 gnd.n5377 99.6594
R7643 gnd.n5416 gnd.n5378 99.6594
R7644 gnd.n5412 gnd.n5379 99.6594
R7645 gnd.n5408 gnd.n5380 99.6594
R7646 gnd.n5404 gnd.n5381 99.6594
R7647 gnd.n5847 gnd.n4484 99.6594
R7648 gnd.n5845 gnd.n5844 99.6594
R7649 gnd.n5840 gnd.n4491 99.6594
R7650 gnd.n5838 gnd.n5837 99.6594
R7651 gnd.n5833 gnd.n4498 99.6594
R7652 gnd.n5831 gnd.n5830 99.6594
R7653 gnd.n5826 gnd.n4505 99.6594
R7654 gnd.n5824 gnd.n5823 99.6594
R7655 gnd.n5819 gnd.n4512 99.6594
R7656 gnd.n5817 gnd.n5816 99.6594
R7657 gnd.n5812 gnd.n4521 99.6594
R7658 gnd.n5810 gnd.n5809 99.6594
R7659 gnd.n5805 gnd.n5804 99.6594
R7660 gnd.n5192 gnd.n5102 99.6594
R7661 gnd.n5190 gnd.n5105 99.6594
R7662 gnd.n5186 gnd.n5185 99.6594
R7663 gnd.n5179 gnd.n5110 99.6594
R7664 gnd.n5178 gnd.n5177 99.6594
R7665 gnd.n5171 gnd.n5116 99.6594
R7666 gnd.n5170 gnd.n5169 99.6594
R7667 gnd.n5163 gnd.n5122 99.6594
R7668 gnd.n5162 gnd.n5161 99.6594
R7669 gnd.n5155 gnd.n5128 99.6594
R7670 gnd.n5154 gnd.n5153 99.6594
R7671 gnd.n5146 gnd.n5134 99.6594
R7672 gnd.n5145 gnd.n5144 99.6594
R7673 gnd.n6854 gnd.n6853 99.6594
R7674 gnd.n6859 gnd.n6858 99.6594
R7675 gnd.n6862 gnd.n6861 99.6594
R7676 gnd.n6867 gnd.n6866 99.6594
R7677 gnd.n6870 gnd.n6869 99.6594
R7678 gnd.n6875 gnd.n6874 99.6594
R7679 gnd.n6878 gnd.n6877 99.6594
R7680 gnd.n6883 gnd.n6882 99.6594
R7681 gnd.n6886 gnd.n99 99.6594
R7682 gnd.n3451 gnd.n3450 99.6594
R7683 gnd.n3454 gnd.n3453 99.6594
R7684 gnd.n3470 gnd.n3469 99.6594
R7685 gnd.n3473 gnd.n3472 99.6594
R7686 gnd.n3489 gnd.n3488 99.6594
R7687 gnd.n3492 gnd.n3491 99.6594
R7688 gnd.n3508 gnd.n3507 99.6594
R7689 gnd.n3511 gnd.n3510 99.6594
R7690 gnd.n3529 gnd.n3528 99.6594
R7691 gnd.n2039 gnd.n2038 99.6594
R7692 gnd.n2040 gnd.n1988 99.6594
R7693 gnd.n2042 gnd.n1996 99.6594
R7694 gnd.n2044 gnd.n2043 99.6594
R7695 gnd.n2045 gnd.n2005 99.6594
R7696 gnd.n2047 gnd.n2014 99.6594
R7697 gnd.n2049 gnd.n2048 99.6594
R7698 gnd.n2050 gnd.n2023 99.6594
R7699 gnd.n2789 gnd.n2788 99.6594
R7700 gnd.n2335 gnd.n875 99.6594
R7701 gnd.n2332 gnd.n876 99.6594
R7702 gnd.n2328 gnd.n877 99.6594
R7703 gnd.n2324 gnd.n878 99.6594
R7704 gnd.n2320 gnd.n879 99.6594
R7705 gnd.n2316 gnd.n880 99.6594
R7706 gnd.n2312 gnd.n881 99.6594
R7707 gnd.n2308 gnd.n882 99.6594
R7708 gnd.n2304 gnd.n883 99.6594
R7709 gnd.n2333 gnd.n875 99.6594
R7710 gnd.n2329 gnd.n876 99.6594
R7711 gnd.n2325 gnd.n877 99.6594
R7712 gnd.n2321 gnd.n878 99.6594
R7713 gnd.n2317 gnd.n879 99.6594
R7714 gnd.n2313 gnd.n880 99.6594
R7715 gnd.n2309 gnd.n881 99.6594
R7716 gnd.n2305 gnd.n882 99.6594
R7717 gnd.n2293 gnd.n883 99.6594
R7718 gnd.n2788 gnd.n2034 99.6594
R7719 gnd.n2050 gnd.n2022 99.6594
R7720 gnd.n2049 gnd.n2015 99.6594
R7721 gnd.n2047 gnd.n2046 99.6594
R7722 gnd.n2045 gnd.n2004 99.6594
R7723 gnd.n2044 gnd.n1997 99.6594
R7724 gnd.n2042 gnd.n2041 99.6594
R7725 gnd.n2040 gnd.n1987 99.6594
R7726 gnd.n2039 gnd.n2037 99.6594
R7727 gnd.n3452 gnd.n3451 99.6594
R7728 gnd.n3453 gnd.n3435 99.6594
R7729 gnd.n3471 gnd.n3470 99.6594
R7730 gnd.n3472 gnd.n3426 99.6594
R7731 gnd.n3490 gnd.n3489 99.6594
R7732 gnd.n3491 gnd.n3417 99.6594
R7733 gnd.n3509 gnd.n3508 99.6594
R7734 gnd.n3510 gnd.n3408 99.6594
R7735 gnd.n3530 gnd.n3529 99.6594
R7736 gnd.n6887 gnd.n6886 99.6594
R7737 gnd.n6882 gnd.n6881 99.6594
R7738 gnd.n6877 gnd.n6876 99.6594
R7739 gnd.n6874 gnd.n6873 99.6594
R7740 gnd.n6869 gnd.n6868 99.6594
R7741 gnd.n6866 gnd.n6865 99.6594
R7742 gnd.n6861 gnd.n6860 99.6594
R7743 gnd.n6858 gnd.n6857 99.6594
R7744 gnd.n6853 gnd.n6852 99.6594
R7745 gnd.n5193 gnd.n5192 99.6594
R7746 gnd.n5187 gnd.n5105 99.6594
R7747 gnd.n5185 gnd.n5184 99.6594
R7748 gnd.n5180 gnd.n5179 99.6594
R7749 gnd.n5177 gnd.n5176 99.6594
R7750 gnd.n5172 gnd.n5171 99.6594
R7751 gnd.n5169 gnd.n5168 99.6594
R7752 gnd.n5164 gnd.n5163 99.6594
R7753 gnd.n5161 gnd.n5160 99.6594
R7754 gnd.n5156 gnd.n5155 99.6594
R7755 gnd.n5153 gnd.n5152 99.6594
R7756 gnd.n5147 gnd.n5146 99.6594
R7757 gnd.n5144 gnd.n5100 99.6594
R7758 gnd.n5804 gnd.n4523 99.6594
R7759 gnd.n5811 gnd.n5810 99.6594
R7760 gnd.n4521 gnd.n4513 99.6594
R7761 gnd.n5818 gnd.n5817 99.6594
R7762 gnd.n4512 gnd.n4506 99.6594
R7763 gnd.n5825 gnd.n5824 99.6594
R7764 gnd.n4505 gnd.n4499 99.6594
R7765 gnd.n5832 gnd.n5831 99.6594
R7766 gnd.n4498 gnd.n4492 99.6594
R7767 gnd.n5839 gnd.n5838 99.6594
R7768 gnd.n4491 gnd.n4485 99.6594
R7769 gnd.n5846 gnd.n5845 99.6594
R7770 gnd.n4484 gnd.n4481 99.6594
R7771 gnd.n5433 gnd.n5383 99.6594
R7772 gnd.n5425 gnd.n5375 99.6594
R7773 gnd.n5421 gnd.n5376 99.6594
R7774 gnd.n5417 gnd.n5377 99.6594
R7775 gnd.n5413 gnd.n5378 99.6594
R7776 gnd.n5409 gnd.n5379 99.6594
R7777 gnd.n5405 gnd.n5380 99.6594
R7778 gnd.n5381 gnd.n5062 99.6594
R7779 gnd.n5857 gnd.n5856 99.6594
R7780 gnd.n4477 gnd.n4469 99.6594
R7781 gnd.n5864 gnd.n5863 99.6594
R7782 gnd.n4468 gnd.n4462 99.6594
R7783 gnd.n5871 gnd.n5870 99.6594
R7784 gnd.n4461 gnd.n4455 99.6594
R7785 gnd.n5878 gnd.n5877 99.6594
R7786 gnd.n4454 gnd.n4451 99.6594
R7787 gnd.n4443 gnd.n887 99.6594
R7788 gnd.n4435 gnd.n857 99.6594
R7789 gnd.n4431 gnd.n858 99.6594
R7790 gnd.n4427 gnd.n859 99.6594
R7791 gnd.n4423 gnd.n860 99.6594
R7792 gnd.n4419 gnd.n861 99.6594
R7793 gnd.n4415 gnd.n862 99.6594
R7794 gnd.n4411 gnd.n863 99.6594
R7795 gnd.n4406 gnd.n864 99.6594
R7796 gnd.n4402 gnd.n865 99.6594
R7797 gnd.n4398 gnd.n866 99.6594
R7798 gnd.n4394 gnd.n867 99.6594
R7799 gnd.n4390 gnd.n868 99.6594
R7800 gnd.n4386 gnd.n869 99.6594
R7801 gnd.n4382 gnd.n870 99.6594
R7802 gnd.n4378 gnd.n871 99.6594
R7803 gnd.n4374 gnd.n872 99.6594
R7804 gnd.n927 gnd.n873 99.6594
R7805 gnd.n4366 gnd.n874 99.6594
R7806 gnd.n2588 gnd.n2052 99.6594
R7807 gnd.n2592 gnd.n2053 99.6594
R7808 gnd.n2596 gnd.n2054 99.6594
R7809 gnd.n2600 gnd.n2055 99.6594
R7810 gnd.n2604 gnd.n2056 99.6594
R7811 gnd.n2608 gnd.n2057 99.6594
R7812 gnd.n2612 gnd.n2058 99.6594
R7813 gnd.n2616 gnd.n2059 99.6594
R7814 gnd.n2620 gnd.n2060 99.6594
R7815 gnd.n2624 gnd.n2061 99.6594
R7816 gnd.n2760 gnd.n2063 99.6594
R7817 gnd.n2764 gnd.n2064 99.6594
R7818 gnd.n2768 gnd.n2065 99.6594
R7819 gnd.n2772 gnd.n2066 99.6594
R7820 gnd.n2776 gnd.n2067 99.6594
R7821 gnd.n2780 gnd.n2068 99.6594
R7822 gnd.n2071 gnd.n2069 99.6594
R7823 gnd.n2786 gnd.n2070 99.6594
R7824 gnd.n3802 gnd.n3801 99.6594
R7825 gnd.n3804 gnd.n3793 99.6594
R7826 gnd.n3813 gnd.n3812 99.6594
R7827 gnd.n3814 gnd.n3789 99.6594
R7828 gnd.n3823 gnd.n3822 99.6594
R7829 gnd.n3824 gnd.n3785 99.6594
R7830 gnd.n3834 gnd.n3833 99.6594
R7831 gnd.n3783 gnd.n1484 99.6594
R7832 gnd.n3847 gnd.n3846 99.6594
R7833 gnd.n3848 gnd.n1480 99.6594
R7834 gnd.n3857 gnd.n3856 99.6594
R7835 gnd.n3858 gnd.n1476 99.6594
R7836 gnd.n3867 gnd.n3866 99.6594
R7837 gnd.n3868 gnd.n1472 99.6594
R7838 gnd.n3877 gnd.n3876 99.6594
R7839 gnd.n3878 gnd.n1468 99.6594
R7840 gnd.n3888 gnd.n3887 99.6594
R7841 gnd.n3891 gnd.n3890 99.6594
R7842 gnd.n172 gnd.n169 99.6594
R7843 gnd.n6946 gnd.n6945 99.6594
R7844 gnd.n168 gnd.n162 99.6594
R7845 gnd.n6953 gnd.n6952 99.6594
R7846 gnd.n161 gnd.n155 99.6594
R7847 gnd.n6960 gnd.n6959 99.6594
R7848 gnd.n154 gnd.n148 99.6594
R7849 gnd.n6967 gnd.n6966 99.6594
R7850 gnd.n147 gnd.n141 99.6594
R7851 gnd.n6974 gnd.n6973 99.6594
R7852 gnd.n140 gnd.n134 99.6594
R7853 gnd.n6984 gnd.n6983 99.6594
R7854 gnd.n133 gnd.n127 99.6594
R7855 gnd.n6991 gnd.n6990 99.6594
R7856 gnd.n126 gnd.n120 99.6594
R7857 gnd.n6998 gnd.n6997 99.6594
R7858 gnd.n119 gnd.n113 99.6594
R7859 gnd.n7005 gnd.n7004 99.6594
R7860 gnd.n112 gnd.n109 99.6594
R7861 gnd.n2836 gnd.n2835 99.6594
R7862 gnd.n1991 gnd.n1967 99.6594
R7863 gnd.n1993 gnd.n1968 99.6594
R7864 gnd.n2001 gnd.n1969 99.6594
R7865 gnd.n2009 gnd.n1970 99.6594
R7866 gnd.n2011 gnd.n1971 99.6594
R7867 gnd.n2019 gnd.n1972 99.6594
R7868 gnd.n2029 gnd.n1973 99.6594
R7869 gnd.n2031 gnd.n1974 99.6594
R7870 gnd.n2543 gnd.n1975 99.6594
R7871 gnd.n2545 gnd.n1976 99.6594
R7872 gnd.n2549 gnd.n1977 99.6594
R7873 gnd.n2555 gnd.n1978 99.6594
R7874 gnd.n2557 gnd.n1979 99.6594
R7875 gnd.n2836 gnd.n1981 99.6594
R7876 gnd.n1992 gnd.n1967 99.6594
R7877 gnd.n2000 gnd.n1968 99.6594
R7878 gnd.n2008 gnd.n1969 99.6594
R7879 gnd.n2010 gnd.n1970 99.6594
R7880 gnd.n2018 gnd.n1971 99.6594
R7881 gnd.n2028 gnd.n1972 99.6594
R7882 gnd.n2030 gnd.n1973 99.6594
R7883 gnd.n2542 gnd.n1974 99.6594
R7884 gnd.n2544 gnd.n1975 99.6594
R7885 gnd.n2548 gnd.n1976 99.6594
R7886 gnd.n2550 gnd.n1977 99.6594
R7887 gnd.n2556 gnd.n1978 99.6594
R7888 gnd.n1979 gnd.n1959 99.6594
R7889 gnd.n3460 gnd.n3440 99.6594
R7890 gnd.n3464 gnd.n3462 99.6594
R7891 gnd.n3479 gnd.n3431 99.6594
R7892 gnd.n3483 gnd.n3481 99.6594
R7893 gnd.n3498 gnd.n3422 99.6594
R7894 gnd.n3502 gnd.n3500 99.6594
R7895 gnd.n3517 gnd.n3413 99.6594
R7896 gnd.n3520 gnd.n3519 99.6594
R7897 gnd.n3521 gnd.n3402 99.6594
R7898 gnd.n3540 gnd.n3539 99.6594
R7899 gnd.n3541 gnd.n3398 99.6594
R7900 gnd.n3550 gnd.n3549 99.6594
R7901 gnd.n3551 gnd.n3394 99.6594
R7902 gnd.n3563 gnd.n3562 99.6594
R7903 gnd.n3562 gnd.n3561 99.6594
R7904 gnd.n3552 gnd.n3551 99.6594
R7905 gnd.n3549 gnd.n3548 99.6594
R7906 gnd.n3542 gnd.n3541 99.6594
R7907 gnd.n3539 gnd.n3538 99.6594
R7908 gnd.n3522 gnd.n3521 99.6594
R7909 gnd.n3519 gnd.n3518 99.6594
R7910 gnd.n3501 gnd.n3413 99.6594
R7911 gnd.n3500 gnd.n3499 99.6594
R7912 gnd.n3482 gnd.n3422 99.6594
R7913 gnd.n3481 gnd.n3480 99.6594
R7914 gnd.n3463 gnd.n3431 99.6594
R7915 gnd.n3462 gnd.n3461 99.6594
R7916 gnd.n3440 gnd.n1303 99.6594
R7917 gnd.n2551 gnd.t116 98.63
R7918 gnd.n6884 gnd.t53 98.63
R7919 gnd.n3405 gnd.t75 98.63
R7920 gnd.n2024 gnd.t107 98.63
R7921 gnd.n3838 gnd.t72 98.63
R7922 gnd.n1464 gnd.t58 98.63
R7923 gnd.n175 gnd.t143 98.63
R7924 gnd.n6977 gnd.t60 98.63
R7925 gnd.n907 gnd.t141 98.63
R7926 gnd.n929 gnd.t129 98.63
R7927 gnd.n2113 gnd.t64 98.63
R7928 gnd.n2091 gnd.t92 98.63
R7929 gnd.n2294 gnd.t83 98.63
R7930 gnd.n3553 gnd.t86 98.63
R7931 gnd.n6424 gnd.n6423 97.2811
R7932 gnd.n6425 gnd.n6424 97.2811
R7933 gnd.n6425 gnd.n457 97.2811
R7934 gnd.n6433 gnd.n457 97.2811
R7935 gnd.n6434 gnd.n6433 97.2811
R7936 gnd.n6435 gnd.n6434 97.2811
R7937 gnd.n6435 gnd.n451 97.2811
R7938 gnd.n6443 gnd.n451 97.2811
R7939 gnd.n6444 gnd.n6443 97.2811
R7940 gnd.n6445 gnd.n6444 97.2811
R7941 gnd.n6445 gnd.n445 97.2811
R7942 gnd.n6453 gnd.n445 97.2811
R7943 gnd.n6454 gnd.n6453 97.2811
R7944 gnd.n6455 gnd.n6454 97.2811
R7945 gnd.n6455 gnd.n439 97.2811
R7946 gnd.n6463 gnd.n439 97.2811
R7947 gnd.n6464 gnd.n6463 97.2811
R7948 gnd.n6465 gnd.n6464 97.2811
R7949 gnd.n6465 gnd.n433 97.2811
R7950 gnd.n6473 gnd.n433 97.2811
R7951 gnd.n6474 gnd.n6473 97.2811
R7952 gnd.n6475 gnd.n6474 97.2811
R7953 gnd.n6475 gnd.n427 97.2811
R7954 gnd.n6483 gnd.n427 97.2811
R7955 gnd.n6484 gnd.n6483 97.2811
R7956 gnd.n6485 gnd.n6484 97.2811
R7957 gnd.n6485 gnd.n421 97.2811
R7958 gnd.n6493 gnd.n421 97.2811
R7959 gnd.n6494 gnd.n6493 97.2811
R7960 gnd.n6495 gnd.n6494 97.2811
R7961 gnd.n6495 gnd.n415 97.2811
R7962 gnd.n6503 gnd.n415 97.2811
R7963 gnd.n6504 gnd.n6503 97.2811
R7964 gnd.n6505 gnd.n6504 97.2811
R7965 gnd.n6505 gnd.n409 97.2811
R7966 gnd.n6513 gnd.n409 97.2811
R7967 gnd.n6514 gnd.n6513 97.2811
R7968 gnd.n6515 gnd.n6514 97.2811
R7969 gnd.n6515 gnd.n403 97.2811
R7970 gnd.n6523 gnd.n403 97.2811
R7971 gnd.n6524 gnd.n6523 97.2811
R7972 gnd.n6525 gnd.n6524 97.2811
R7973 gnd.n6525 gnd.n397 97.2811
R7974 gnd.n6533 gnd.n397 97.2811
R7975 gnd.n6534 gnd.n6533 97.2811
R7976 gnd.n6535 gnd.n6534 97.2811
R7977 gnd.n6535 gnd.n391 97.2811
R7978 gnd.n6543 gnd.n391 97.2811
R7979 gnd.n6544 gnd.n6543 97.2811
R7980 gnd.n6545 gnd.n6544 97.2811
R7981 gnd.n6545 gnd.n385 97.2811
R7982 gnd.n6553 gnd.n385 97.2811
R7983 gnd.n6554 gnd.n6553 97.2811
R7984 gnd.n6555 gnd.n6554 97.2811
R7985 gnd.n6555 gnd.n379 97.2811
R7986 gnd.n6563 gnd.n379 97.2811
R7987 gnd.n6564 gnd.n6563 97.2811
R7988 gnd.n6565 gnd.n6564 97.2811
R7989 gnd.n6565 gnd.n373 97.2811
R7990 gnd.n6573 gnd.n373 97.2811
R7991 gnd.n6574 gnd.n6573 97.2811
R7992 gnd.n6575 gnd.n6574 97.2811
R7993 gnd.n6575 gnd.n367 97.2811
R7994 gnd.n6583 gnd.n367 97.2811
R7995 gnd.n6584 gnd.n6583 97.2811
R7996 gnd.n6585 gnd.n6584 97.2811
R7997 gnd.n6585 gnd.n361 97.2811
R7998 gnd.n6593 gnd.n361 97.2811
R7999 gnd.n6594 gnd.n6593 97.2811
R8000 gnd.n6595 gnd.n6594 97.2811
R8001 gnd.n6595 gnd.n355 97.2811
R8002 gnd.n6603 gnd.n355 97.2811
R8003 gnd.n6604 gnd.n6603 97.2811
R8004 gnd.n6605 gnd.n6604 97.2811
R8005 gnd.n6605 gnd.n349 97.2811
R8006 gnd.n6613 gnd.n349 97.2811
R8007 gnd.n6614 gnd.n6613 97.2811
R8008 gnd.n6615 gnd.n6614 97.2811
R8009 gnd.n6615 gnd.n343 97.2811
R8010 gnd.n6623 gnd.n343 97.2811
R8011 gnd.n6624 gnd.n6623 97.2811
R8012 gnd.n6626 gnd.n6624 97.2811
R8013 gnd.n6626 gnd.n6625 97.2811
R8014 gnd.n2629 gnd.t46 88.9408
R8015 gnd.n1525 gnd.t49 88.9408
R8016 gnd.n2693 gnd.t96 88.933
R8017 gnd.n3645 gnd.t98 88.933
R8018 gnd.n1848 gnd.n1847 81.8399
R8019 gnd.n5401 gnd.t68 74.8376
R8020 gnd.n4475 gnd.t112 74.8376
R8021 gnd.n2630 gnd.t45 72.8438
R8022 gnd.n1526 gnd.t50 72.8438
R8023 gnd.n1849 gnd.n1842 72.8411
R8024 gnd.n1855 gnd.n1840 72.8411
R8025 gnd.n3641 gnd.n3640 72.8411
R8026 gnd.n2552 gnd.t115 72.836
R8027 gnd.n2694 gnd.t95 72.836
R8028 gnd.n3646 gnd.t99 72.836
R8029 gnd.n6885 gnd.t54 72.836
R8030 gnd.n3406 gnd.t74 72.836
R8031 gnd.n2025 gnd.t108 72.836
R8032 gnd.n3839 gnd.t71 72.836
R8033 gnd.n1465 gnd.t57 72.836
R8034 gnd.n176 gnd.t144 72.836
R8035 gnd.n6978 gnd.t61 72.836
R8036 gnd.n908 gnd.t140 72.836
R8037 gnd.n930 gnd.t128 72.836
R8038 gnd.n2114 gnd.t65 72.836
R8039 gnd.n2092 gnd.t93 72.836
R8040 gnd.n2295 gnd.t82 72.836
R8041 gnd.n3554 gnd.t87 72.836
R8042 gnd.n3706 gnd.n1493 71.676
R8043 gnd.n3702 gnd.n1494 71.676
R8044 gnd.n3698 gnd.n1495 71.676
R8045 gnd.n3694 gnd.n1496 71.676
R8046 gnd.n3690 gnd.n1497 71.676
R8047 gnd.n3686 gnd.n1498 71.676
R8048 gnd.n3682 gnd.n1499 71.676
R8049 gnd.n3678 gnd.n1500 71.676
R8050 gnd.n3674 gnd.n1501 71.676
R8051 gnd.n3670 gnd.n1502 71.676
R8052 gnd.n3666 gnd.n1503 71.676
R8053 gnd.n3662 gnd.n1504 71.676
R8054 gnd.n3658 gnd.n1505 71.676
R8055 gnd.n3654 gnd.n1506 71.676
R8056 gnd.n3649 gnd.n1507 71.676
R8057 gnd.n1508 gnd.n1491 71.676
R8058 gnd.n3778 gnd.n1490 71.676
R8059 gnd.n3776 gnd.n3775 71.676
R8060 gnd.n3770 gnd.n1523 71.676
R8061 gnd.n3766 gnd.n1522 71.676
R8062 gnd.n3762 gnd.n1521 71.676
R8063 gnd.n3758 gnd.n1520 71.676
R8064 gnd.n3754 gnd.n1519 71.676
R8065 gnd.n3750 gnd.n1518 71.676
R8066 gnd.n3746 gnd.n1517 71.676
R8067 gnd.n3742 gnd.n1516 71.676
R8068 gnd.n3738 gnd.n1515 71.676
R8069 gnd.n3734 gnd.n1514 71.676
R8070 gnd.n3730 gnd.n1513 71.676
R8071 gnd.n3726 gnd.n1512 71.676
R8072 gnd.n3722 gnd.n1511 71.676
R8073 gnd.n3718 gnd.n1510 71.676
R8074 gnd.n3714 gnd.n1509 71.676
R8075 gnd.n2966 gnd.n1837 71.676
R8076 gnd.n2696 gnd.n1863 71.676
R8077 gnd.n2700 gnd.n1864 71.676
R8078 gnd.n2704 gnd.n1865 71.676
R8079 gnd.n2708 gnd.n1866 71.676
R8080 gnd.n2712 gnd.n1867 71.676
R8081 gnd.n2716 gnd.n1868 71.676
R8082 gnd.n2720 gnd.n1869 71.676
R8083 gnd.n2724 gnd.n1870 71.676
R8084 gnd.n2728 gnd.n1871 71.676
R8085 gnd.n2732 gnd.n1872 71.676
R8086 gnd.n2736 gnd.n1873 71.676
R8087 gnd.n2740 gnd.n1874 71.676
R8088 gnd.n2744 gnd.n1875 71.676
R8089 gnd.n2748 gnd.n1876 71.676
R8090 gnd.n2752 gnd.n1877 71.676
R8091 gnd.n2755 gnd.n1879 71.676
R8092 gnd.n2689 gnd.n1880 71.676
R8093 gnd.n2684 gnd.n1881 71.676
R8094 gnd.n2680 gnd.n1882 71.676
R8095 gnd.n2676 gnd.n1883 71.676
R8096 gnd.n2672 gnd.n1884 71.676
R8097 gnd.n2668 gnd.n1885 71.676
R8098 gnd.n2664 gnd.n1886 71.676
R8099 gnd.n2660 gnd.n1887 71.676
R8100 gnd.n2656 gnd.n1888 71.676
R8101 gnd.n2652 gnd.n1889 71.676
R8102 gnd.n2648 gnd.n1890 71.676
R8103 gnd.n2644 gnd.n1891 71.676
R8104 gnd.n2640 gnd.n1892 71.676
R8105 gnd.n2636 gnd.n1893 71.676
R8106 gnd.n2632 gnd.n1894 71.676
R8107 gnd.n2967 gnd.n2966 71.676
R8108 gnd.n2699 gnd.n1863 71.676
R8109 gnd.n2703 gnd.n1864 71.676
R8110 gnd.n2707 gnd.n1865 71.676
R8111 gnd.n2711 gnd.n1866 71.676
R8112 gnd.n2715 gnd.n1867 71.676
R8113 gnd.n2719 gnd.n1868 71.676
R8114 gnd.n2723 gnd.n1869 71.676
R8115 gnd.n2727 gnd.n1870 71.676
R8116 gnd.n2731 gnd.n1871 71.676
R8117 gnd.n2735 gnd.n1872 71.676
R8118 gnd.n2739 gnd.n1873 71.676
R8119 gnd.n2743 gnd.n1874 71.676
R8120 gnd.n2747 gnd.n1875 71.676
R8121 gnd.n2751 gnd.n1876 71.676
R8122 gnd.n2756 gnd.n1878 71.676
R8123 gnd.n2690 gnd.n1879 71.676
R8124 gnd.n2685 gnd.n1880 71.676
R8125 gnd.n2681 gnd.n1881 71.676
R8126 gnd.n2677 gnd.n1882 71.676
R8127 gnd.n2673 gnd.n1883 71.676
R8128 gnd.n2669 gnd.n1884 71.676
R8129 gnd.n2665 gnd.n1885 71.676
R8130 gnd.n2661 gnd.n1886 71.676
R8131 gnd.n2657 gnd.n1887 71.676
R8132 gnd.n2653 gnd.n1888 71.676
R8133 gnd.n2649 gnd.n1889 71.676
R8134 gnd.n2645 gnd.n1890 71.676
R8135 gnd.n2641 gnd.n1891 71.676
R8136 gnd.n2637 gnd.n1892 71.676
R8137 gnd.n2633 gnd.n1893 71.676
R8138 gnd.n1894 gnd.n1834 71.676
R8139 gnd.n3717 gnd.n1509 71.676
R8140 gnd.n3721 gnd.n1510 71.676
R8141 gnd.n3725 gnd.n1511 71.676
R8142 gnd.n3729 gnd.n1512 71.676
R8143 gnd.n3733 gnd.n1513 71.676
R8144 gnd.n3737 gnd.n1514 71.676
R8145 gnd.n3741 gnd.n1515 71.676
R8146 gnd.n3745 gnd.n1516 71.676
R8147 gnd.n3749 gnd.n1517 71.676
R8148 gnd.n3753 gnd.n1518 71.676
R8149 gnd.n3757 gnd.n1519 71.676
R8150 gnd.n3761 gnd.n1520 71.676
R8151 gnd.n3765 gnd.n1521 71.676
R8152 gnd.n3769 gnd.n1522 71.676
R8153 gnd.n1524 gnd.n1523 71.676
R8154 gnd.n3777 gnd.n3776 71.676
R8155 gnd.n3781 gnd.n3780 71.676
R8156 gnd.n3648 gnd.n1508 71.676
R8157 gnd.n3653 gnd.n1507 71.676
R8158 gnd.n3657 gnd.n1506 71.676
R8159 gnd.n3661 gnd.n1505 71.676
R8160 gnd.n3665 gnd.n1504 71.676
R8161 gnd.n3669 gnd.n1503 71.676
R8162 gnd.n3673 gnd.n1502 71.676
R8163 gnd.n3677 gnd.n1501 71.676
R8164 gnd.n3681 gnd.n1500 71.676
R8165 gnd.n3685 gnd.n1499 71.676
R8166 gnd.n3689 gnd.n1498 71.676
R8167 gnd.n3693 gnd.n1497 71.676
R8168 gnd.n3697 gnd.n1496 71.676
R8169 gnd.n3701 gnd.n1495 71.676
R8170 gnd.n3705 gnd.n1494 71.676
R8171 gnd.n1531 gnd.n1493 71.676
R8172 gnd.n8 gnd.t312 69.1507
R8173 gnd.n14 gnd.t11 68.4792
R8174 gnd.n13 gnd.t153 68.4792
R8175 gnd.n12 gnd.t1 68.4792
R8176 gnd.n11 gnd.t34 68.4792
R8177 gnd.n10 gnd.t9 68.4792
R8178 gnd.n9 gnd.t30 68.4792
R8179 gnd.n8 gnd.t3 68.4792
R8180 gnd.n5200 gnd.n5101 64.369
R8181 gnd.n2687 gnd.n2630 59.5399
R8182 gnd.n3772 gnd.n1526 59.5399
R8183 gnd.n2695 gnd.n2694 59.5399
R8184 gnd.n3651 gnd.n3646 59.5399
R8185 gnd.n2970 gnd.n1858 59.1804
R8186 gnd.n6625 gnd.n205 58.3688
R8187 gnd.n5887 gnd.n4445 57.3586
R8188 gnd.n4444 gnd.n885 57.3586
R8189 gnd.n7014 gnd.n102 57.3586
R8190 gnd.n5325 gnd.t160 56.607
R8191 gnd.n48 gnd.t261 56.607
R8192 gnd.n5294 gnd.t224 56.407
R8193 gnd.n5309 gnd.t201 56.407
R8194 gnd.n17 gnd.t256 56.407
R8195 gnd.n32 gnd.t232 56.407
R8196 gnd.n5338 gnd.t273 55.8337
R8197 gnd.n5307 gnd.t230 55.8337
R8198 gnd.n5322 gnd.t211 55.8337
R8199 gnd.n61 gnd.t239 55.8337
R8200 gnd.n30 gnd.t263 55.8337
R8201 gnd.n45 gnd.t242 55.8337
R8202 gnd.n1846 gnd.n1845 54.358
R8203 gnd.n3638 gnd.n3637 54.358
R8204 gnd.n5325 gnd.n5324 53.0052
R8205 gnd.n5327 gnd.n5326 53.0052
R8206 gnd.n5329 gnd.n5328 53.0052
R8207 gnd.n5331 gnd.n5330 53.0052
R8208 gnd.n5333 gnd.n5332 53.0052
R8209 gnd.n5335 gnd.n5334 53.0052
R8210 gnd.n5337 gnd.n5336 53.0052
R8211 gnd.n5294 gnd.n5293 53.0052
R8212 gnd.n5296 gnd.n5295 53.0052
R8213 gnd.n5298 gnd.n5297 53.0052
R8214 gnd.n5300 gnd.n5299 53.0052
R8215 gnd.n5302 gnd.n5301 53.0052
R8216 gnd.n5304 gnd.n5303 53.0052
R8217 gnd.n5306 gnd.n5305 53.0052
R8218 gnd.n5309 gnd.n5308 53.0052
R8219 gnd.n5311 gnd.n5310 53.0052
R8220 gnd.n5313 gnd.n5312 53.0052
R8221 gnd.n5315 gnd.n5314 53.0052
R8222 gnd.n5317 gnd.n5316 53.0052
R8223 gnd.n5319 gnd.n5318 53.0052
R8224 gnd.n5321 gnd.n5320 53.0052
R8225 gnd.n60 gnd.n59 53.0052
R8226 gnd.n58 gnd.n57 53.0052
R8227 gnd.n56 gnd.n55 53.0052
R8228 gnd.n54 gnd.n53 53.0052
R8229 gnd.n52 gnd.n51 53.0052
R8230 gnd.n50 gnd.n49 53.0052
R8231 gnd.n48 gnd.n47 53.0052
R8232 gnd.n29 gnd.n28 53.0052
R8233 gnd.n27 gnd.n26 53.0052
R8234 gnd.n25 gnd.n24 53.0052
R8235 gnd.n23 gnd.n22 53.0052
R8236 gnd.n21 gnd.n20 53.0052
R8237 gnd.n19 gnd.n18 53.0052
R8238 gnd.n17 gnd.n16 53.0052
R8239 gnd.n44 gnd.n43 53.0052
R8240 gnd.n42 gnd.n41 53.0052
R8241 gnd.n40 gnd.n39 53.0052
R8242 gnd.n38 gnd.n37 53.0052
R8243 gnd.n36 gnd.n35 53.0052
R8244 gnd.n34 gnd.n33 53.0052
R8245 gnd.n32 gnd.n31 53.0052
R8246 gnd.n3629 gnd.n3628 52.4801
R8247 gnd.n4769 gnd.t19 52.3082
R8248 gnd.n4737 gnd.t314 52.3082
R8249 gnd.n4705 gnd.t156 52.3082
R8250 gnd.n4674 gnd.t148 52.3082
R8251 gnd.n4642 gnd.t16 52.3082
R8252 gnd.n4610 gnd.t306 52.3082
R8253 gnd.n4578 gnd.t310 52.3082
R8254 gnd.n4547 gnd.t32 52.3082
R8255 gnd.n4599 gnd.n4567 51.4173
R8256 gnd.n4663 gnd.n4662 50.455
R8257 gnd.n4631 gnd.n4630 50.455
R8258 gnd.n4599 gnd.n4598 50.455
R8259 gnd.n5138 gnd.n5137 45.1884
R8260 gnd.n4519 gnd.n4518 45.1884
R8261 gnd.n3709 gnd.n3644 44.3322
R8262 gnd.n1849 gnd.n1848 44.3189
R8263 gnd.n2553 gnd.n2552 42.2793
R8264 gnd.n5150 gnd.n5138 42.2793
R8265 gnd.n4520 gnd.n4519 42.2793
R8266 gnd.n5403 gnd.n5401 42.2793
R8267 gnd.n4476 gnd.n4475 42.2793
R8268 gnd.n6890 gnd.n6885 42.2793
R8269 gnd.n3407 gnd.n3406 42.2793
R8270 gnd.n2026 gnd.n2025 42.2793
R8271 gnd.n1466 gnd.n1465 42.2793
R8272 gnd.n6942 gnd.n176 42.2793
R8273 gnd.n6979 gnd.n6978 42.2793
R8274 gnd.n4408 gnd.n908 42.2793
R8275 gnd.n931 gnd.n930 42.2793
R8276 gnd.n2587 gnd.n2114 42.2793
R8277 gnd.n2296 gnd.n2295 42.2793
R8278 gnd.n3555 gnd.n3554 42.2793
R8279 gnd.n1847 gnd.n1846 41.6274
R8280 gnd.n3639 gnd.n3638 41.6274
R8281 gnd.n1856 gnd.n1855 40.8975
R8282 gnd.n3642 gnd.n3641 40.8975
R8283 gnd.n3840 gnd.n3839 36.9518
R8284 gnd.n2758 gnd.n2092 36.9518
R8285 gnd.n1855 gnd.n1854 35.055
R8286 gnd.n1850 gnd.n1849 35.055
R8287 gnd.n3631 gnd.n3630 35.055
R8288 gnd.n3641 gnd.n3627 35.055
R8289 gnd.n6063 gnd.n6062 33.6139
R8290 gnd.n6062 gnd.n677 33.6139
R8291 gnd.n6056 gnd.n677 33.6139
R8292 gnd.n6056 gnd.n6055 33.6139
R8293 gnd.n6055 gnd.n6054 33.6139
R8294 gnd.n6054 gnd.n685 33.6139
R8295 gnd.n6048 gnd.n685 33.6139
R8296 gnd.n6048 gnd.n6047 33.6139
R8297 gnd.n6047 gnd.n6046 33.6139
R8298 gnd.n6046 gnd.n693 33.6139
R8299 gnd.n6040 gnd.n693 33.6139
R8300 gnd.n6040 gnd.n6039 33.6139
R8301 gnd.n6039 gnd.n6038 33.6139
R8302 gnd.n6038 gnd.n701 33.6139
R8303 gnd.n6032 gnd.n701 33.6139
R8304 gnd.n6032 gnd.n6031 33.6139
R8305 gnd.n6031 gnd.n6030 33.6139
R8306 gnd.n6030 gnd.n709 33.6139
R8307 gnd.n6024 gnd.n709 33.6139
R8308 gnd.n6024 gnd.n6023 33.6139
R8309 gnd.n6023 gnd.n6022 33.6139
R8310 gnd.n6022 gnd.n717 33.6139
R8311 gnd.n6016 gnd.n717 33.6139
R8312 gnd.n6016 gnd.n6015 33.6139
R8313 gnd.n6015 gnd.n6014 33.6139
R8314 gnd.n6014 gnd.n725 33.6139
R8315 gnd.n6008 gnd.n725 33.6139
R8316 gnd.n6008 gnd.n6007 33.6139
R8317 gnd.n6007 gnd.n6006 33.6139
R8318 gnd.n6006 gnd.n733 33.6139
R8319 gnd.n6000 gnd.n733 33.6139
R8320 gnd.n6000 gnd.n5999 33.6139
R8321 gnd.n5999 gnd.n5998 33.6139
R8322 gnd.n5998 gnd.n741 33.6139
R8323 gnd.n5992 gnd.n741 33.6139
R8324 gnd.n5992 gnd.n5991 33.6139
R8325 gnd.n5991 gnd.n5990 33.6139
R8326 gnd.n5990 gnd.n749 33.6139
R8327 gnd.n5984 gnd.n749 33.6139
R8328 gnd.n5984 gnd.n5983 33.6139
R8329 gnd.n5983 gnd.n5982 33.6139
R8330 gnd.n5982 gnd.n757 33.6139
R8331 gnd.n5976 gnd.n757 33.6139
R8332 gnd.n5976 gnd.n5975 33.6139
R8333 gnd.n5975 gnd.n5974 33.6139
R8334 gnd.n5974 gnd.n765 33.6139
R8335 gnd.n5968 gnd.n765 33.6139
R8336 gnd.n5968 gnd.n5967 33.6139
R8337 gnd.n5967 gnd.n5966 33.6139
R8338 gnd.n5966 gnd.n773 33.6139
R8339 gnd.n5960 gnd.n773 33.6139
R8340 gnd.n5960 gnd.n5959 33.6139
R8341 gnd.n5959 gnd.n5958 33.6139
R8342 gnd.n5958 gnd.n781 33.6139
R8343 gnd.n5952 gnd.n781 33.6139
R8344 gnd.n5952 gnd.n5951 33.6139
R8345 gnd.n5951 gnd.n5950 33.6139
R8346 gnd.n5950 gnd.n789 33.6139
R8347 gnd.n5944 gnd.n789 33.6139
R8348 gnd.n5944 gnd.n5943 33.6139
R8349 gnd.n5943 gnd.n5942 33.6139
R8350 gnd.n5942 gnd.n797 33.6139
R8351 gnd.n5936 gnd.n797 33.6139
R8352 gnd.n5936 gnd.n5935 33.6139
R8353 gnd.n5935 gnd.n5934 33.6139
R8354 gnd.n5934 gnd.n805 33.6139
R8355 gnd.n5928 gnd.n805 33.6139
R8356 gnd.n5928 gnd.n5927 33.6139
R8357 gnd.n5927 gnd.n5926 33.6139
R8358 gnd.n5926 gnd.n813 33.6139
R8359 gnd.n5920 gnd.n813 33.6139
R8360 gnd.n5920 gnd.n5919 33.6139
R8361 gnd.n5919 gnd.n5918 33.6139
R8362 gnd.n5918 gnd.n821 33.6139
R8363 gnd.n5912 gnd.n821 33.6139
R8364 gnd.n5912 gnd.n5911 33.6139
R8365 gnd.n5911 gnd.n5910 33.6139
R8366 gnd.n5910 gnd.n829 33.6139
R8367 gnd.n5904 gnd.n829 33.6139
R8368 gnd.n5904 gnd.n5903 33.6139
R8369 gnd.n5903 gnd.n5902 33.6139
R8370 gnd.n5902 gnd.n837 33.6139
R8371 gnd.n5896 gnd.n837 33.6139
R8372 gnd.n3715 gnd.n1527 32.3127
R8373 gnd.n2977 gnd.n1833 32.3127
R8374 gnd.n5200 gnd.n5096 31.8661
R8375 gnd.n5208 gnd.n5096 31.8661
R8376 gnd.n5216 gnd.n5090 31.8661
R8377 gnd.n5216 gnd.n5084 31.8661
R8378 gnd.n5224 gnd.n5084 31.8661
R8379 gnd.n5224 gnd.n5077 31.8661
R8380 gnd.n5232 gnd.n5077 31.8661
R8381 gnd.n5232 gnd.n5078 31.8661
R8382 gnd.n5444 gnd.n5063 31.8661
R8383 gnd.n2352 gnd.n885 31.8661
R8384 gnd.n4357 gnd.n939 31.8661
R8385 gnd.n4357 gnd.n941 31.8661
R8386 gnd.n4351 gnd.n941 31.8661
R8387 gnd.n4351 gnd.n953 31.8661
R8388 gnd.n4345 gnd.n964 31.8661
R8389 gnd.n4339 gnd.n964 31.8661
R8390 gnd.n4333 gnd.n981 31.8661
R8391 gnd.n4327 gnd.n991 31.8661
R8392 gnd.n4327 gnd.n994 31.8661
R8393 gnd.n4321 gnd.n1004 31.8661
R8394 gnd.n4315 gnd.n1004 31.8661
R8395 gnd.n4309 gnd.n1021 31.8661
R8396 gnd.n4303 gnd.n1031 31.8661
R8397 gnd.n4303 gnd.n1034 31.8661
R8398 gnd.n4297 gnd.n1044 31.8661
R8399 gnd.n4291 gnd.n1044 31.8661
R8400 gnd.n4285 gnd.n1059 31.8661
R8401 gnd.n4278 gnd.n1069 31.8661
R8402 gnd.n2035 gnd.n1194 31.8661
R8403 gnd.n2051 gnd.n1966 31.8661
R8404 gnd.n2838 gnd.n1966 31.8661
R8405 gnd.n2846 gnd.n1960 31.8661
R8406 gnd.n4074 gnd.n1306 31.8661
R8407 gnd.n4068 gnd.n4067 31.8661
R8408 gnd.n4067 gnd.n4066 31.8661
R8409 gnd.n4060 gnd.n1324 31.8661
R8410 gnd.n6680 gnd.n300 31.8661
R8411 gnd.n6750 gnd.n292 31.8661
R8412 gnd.n6756 gnd.n285 31.8661
R8413 gnd.n6756 gnd.n288 31.8661
R8414 gnd.n6779 gnd.n249 31.8661
R8415 gnd.n6787 gnd.n249 31.8661
R8416 gnd.n6795 gnd.n242 31.8661
R8417 gnd.n6803 gnd.n232 31.8661
R8418 gnd.n6803 gnd.n235 31.8661
R8419 gnd.n6811 gnd.n219 31.8661
R8420 gnd.n6819 gnd.n219 31.8661
R8421 gnd.n6827 gnd.n212 31.8661
R8422 gnd.n6835 gnd.n203 31.8661
R8423 gnd.n6843 gnd.n188 31.8661
R8424 gnd.n6926 gnd.n188 31.8661
R8425 gnd.n6926 gnd.n181 31.8661
R8426 gnd.n6934 gnd.n181 31.8661
R8427 gnd.n7014 gnd.n100 31.8661
R8428 gnd.n4333 gnd.t171 27.7236
R8429 gnd.t204 gnd.n212 27.7236
R8430 gnd.n4309 gnd.t167 27.0862
R8431 gnd.t246 gnd.n242 27.0862
R8432 gnd.n2417 gnd.n1079 26.7676
R8433 gnd.n4266 gnd.n1086 26.7676
R8434 gnd.n2426 gnd.n2183 26.7676
R8435 gnd.n4260 gnd.n1096 26.7676
R8436 gnd.n4254 gnd.n1107 26.7676
R8437 gnd.n2473 gnd.n1110 26.7676
R8438 gnd.n2442 gnd.n1120 26.7676
R8439 gnd.n4242 gnd.n1128 26.7676
R8440 gnd.n2447 gnd.n2446 26.7676
R8441 gnd.n4236 gnd.n1138 26.7676
R8442 gnd.n4230 gnd.n1149 26.7676
R8443 gnd.n2519 gnd.n1152 26.7676
R8444 gnd.n2527 gnd.n1162 26.7676
R8445 gnd.n4218 gnd.n1170 26.7676
R8446 gnd.n2536 gnd.n1173 26.7676
R8447 gnd.n4212 gnd.n1181 26.7676
R8448 gnd.n4206 gnd.n1191 26.7676
R8449 gnd.n4059 gnd.n1327 26.7676
R8450 gnd.n4053 gnd.n1339 26.7676
R8451 gnd.n3897 gnd.n1435 26.7676
R8452 gnd.n3930 gnd.n3929 26.7676
R8453 gnd.n1438 gnd.n1430 26.7676
R8454 gnd.n3922 gnd.n1407 26.7676
R8455 gnd.n3967 gnd.n3966 26.7676
R8456 gnd.n3977 gnd.n1400 26.7676
R8457 gnd.n3959 gnd.n1421 26.7676
R8458 gnd.n3958 gnd.n1368 26.7676
R8459 gnd.n4020 gnd.n4019 26.7676
R8460 gnd.n4028 gnd.n1362 26.7676
R8461 gnd.n3993 gnd.n323 26.7676
R8462 gnd.n4010 gnd.n313 26.7676
R8463 gnd.n6662 gnd.n315 26.7676
R8464 gnd.n6643 gnd.n6642 26.7676
R8465 gnd.n333 gnd.n269 26.7676
R8466 gnd.n1059 gnd.t161 26.4489
R8467 gnd.n4285 gnd.t202 26.4489
R8468 gnd.t234 gnd.n292 26.4489
R8469 gnd.n6750 gnd.t240 26.4489
R8470 gnd.n1021 gnd.t169 25.8116
R8471 gnd.n6795 gnd.t253 25.8116
R8472 gnd.n2552 gnd.n2551 25.7944
R8473 gnd.n5401 gnd.n5400 25.7944
R8474 gnd.n4475 gnd.n4474 25.7944
R8475 gnd.n6885 gnd.n6884 25.7944
R8476 gnd.n3406 gnd.n3405 25.7944
R8477 gnd.n2025 gnd.n2024 25.7944
R8478 gnd.n3839 gnd.n3838 25.7944
R8479 gnd.n1465 gnd.n1464 25.7944
R8480 gnd.n176 gnd.n175 25.7944
R8481 gnd.n6978 gnd.n6977 25.7944
R8482 gnd.n908 gnd.n907 25.7944
R8483 gnd.n930 gnd.n929 25.7944
R8484 gnd.n2114 gnd.n2113 25.7944
R8485 gnd.n2092 gnd.n2091 25.7944
R8486 gnd.n2295 gnd.n2294 25.7944
R8487 gnd.n3554 gnd.n3553 25.7944
R8488 gnd.n981 gnd.t227 25.1743
R8489 gnd.n6827 gnd.t192 25.1743
R8490 gnd.n5445 gnd.n5053 24.8557
R8491 gnd.n5056 gnd.n5046 24.8557
R8492 gnd.n5475 gnd.n5039 24.8557
R8493 gnd.n5476 gnd.n5028 24.8557
R8494 gnd.n5031 gnd.n5019 24.8557
R8495 gnd.n5497 gnd.n5020 24.8557
R8496 gnd.n5518 gnd.n5517 24.8557
R8497 gnd.n5005 gnd.n4993 24.8557
R8498 gnd.n5528 gnd.n4994 24.8557
R8499 gnd.n5538 gnd.n4976 24.8557
R8500 gnd.n5549 gnd.n5548 24.8557
R8501 gnd.n5559 gnd.n4969 24.8557
R8502 gnd.n5568 gnd.n4961 24.8557
R8503 gnd.n5569 gnd.n4950 24.8557
R8504 gnd.n5580 gnd.n5579 24.8557
R8505 gnd.n5599 gnd.n4936 24.8557
R8506 gnd.n5611 gnd.n5610 24.8557
R8507 gnd.n5272 gnd.n4928 24.8557
R8508 gnd.n5621 gnd.n4918 24.8557
R8509 gnd.n5630 gnd.n4911 24.8557
R8510 gnd.n5641 gnd.n5640 24.8557
R8511 gnd.n4904 gnd.n4894 24.8557
R8512 gnd.n4887 gnd.n4881 24.8557
R8513 gnd.n5672 gnd.n5671 24.8557
R8514 gnd.n5682 gnd.n5681 24.8557
R8515 gnd.n4871 gnd.n4862 24.8557
R8516 gnd.n4853 gnd.n4852 24.8557
R8517 gnd.n5716 gnd.n4845 24.8557
R8518 gnd.n5729 gnd.n5728 24.8557
R8519 gnd.n5741 gnd.n4832 24.8557
R8520 gnd.n5761 gnd.n4818 24.8557
R8521 gnd.n5772 gnd.n5771 24.8557
R8522 gnd.n5791 gnd.n4533 24.8557
R8523 gnd.n4805 gnd.n4534 24.8557
R8524 gnd.n5888 gnd.n854 24.8557
R8525 gnd.n5466 gnd.t31 23.2624
R8526 gnd.n6835 gnd.n205 22.9437
R8527 gnd.n5456 gnd.t67 22.6251
R8528 gnd.n2352 gnd.t81 22.6251
R8529 gnd.n2580 gnd.t63 22.6251
R8530 gnd.n3905 gnd.t56 22.6251
R8531 gnd.t52 gnd.n100 22.6251
R8532 gnd.n5435 gnd.t147 21.3504
R8533 gnd.t291 gnd.n4839 20.7131
R8534 gnd.t190 gnd.n1099 20.7131
R8535 gnd.n4011 gnd.t214 20.7131
R8536 gnd.n2787 gnd.n2035 20.3945
R8537 gnd.n1324 gnd.n1316 20.3945
R8538 gnd.n5896 gnd.n5895 20.1686
R8539 gnd.n2973 gnd.n2970 20.1371
R8540 gnd.n3710 gnd.n3709 20.1371
R8541 gnd.n5661 gnd.t293 20.0758
R8542 gnd.t178 gnd.n1141 20.0758
R8543 gnd.t188 gnd.n1398 20.0758
R8544 gnd.n1843 gnd.t102 19.8005
R8545 gnd.n1843 gnd.t138 19.8005
R8546 gnd.n1844 gnd.t122 19.8005
R8547 gnd.n1844 gnd.t43 19.8005
R8548 gnd.n3635 gnd.t132 19.8005
R8549 gnd.n3635 gnd.t90 19.8005
R8550 gnd.n3636 gnd.t40 19.8005
R8551 gnd.n3636 gnd.t119 19.8005
R8552 gnd.n1840 gnd.n1839 19.5087
R8553 gnd.n1853 gnd.n1840 19.5087
R8554 gnd.n1851 gnd.n1842 19.5087
R8555 gnd.n3640 gnd.n3634 19.5087
R8556 gnd.t299 gnd.n4925 19.4385
R8557 gnd.n2850 gnd.n1957 19.3944
R8558 gnd.n2854 gnd.n1957 19.3944
R8559 gnd.n2854 gnd.n1946 19.3944
R8560 gnd.n2870 gnd.n1946 19.3944
R8561 gnd.n2870 gnd.n1944 19.3944
R8562 gnd.n2874 gnd.n1944 19.3944
R8563 gnd.n2874 gnd.n1933 19.3944
R8564 gnd.n2890 gnd.n1933 19.3944
R8565 gnd.n2890 gnd.n1931 19.3944
R8566 gnd.n2894 gnd.n1931 19.3944
R8567 gnd.n2894 gnd.n1920 19.3944
R8568 gnd.n2910 gnd.n1920 19.3944
R8569 gnd.n2910 gnd.n1918 19.3944
R8570 gnd.n2914 gnd.n1918 19.3944
R8571 gnd.n2914 gnd.n1907 19.3944
R8572 gnd.n2930 gnd.n1907 19.3944
R8573 gnd.n2930 gnd.n1904 19.3944
R8574 gnd.n2952 gnd.n1904 19.3944
R8575 gnd.n2952 gnd.n1905 19.3944
R8576 gnd.n2948 gnd.n1905 19.3944
R8577 gnd.n2948 gnd.n2947 19.3944
R8578 gnd.n2947 gnd.n2946 19.3944
R8579 gnd.n2946 gnd.n2937 19.3944
R8580 gnd.n2942 gnd.n2937 19.3944
R8581 gnd.n2942 gnd.n1804 19.3944
R8582 gnd.n3013 gnd.n1804 19.3944
R8583 gnd.n3014 gnd.n3013 19.3944
R8584 gnd.n3014 gnd.n1801 19.3944
R8585 gnd.n3024 gnd.n1801 19.3944
R8586 gnd.n3024 gnd.n1802 19.3944
R8587 gnd.n3020 gnd.n1802 19.3944
R8588 gnd.n3020 gnd.n3019 19.3944
R8589 gnd.n3019 gnd.n1753 19.3944
R8590 gnd.n3132 gnd.n1753 19.3944
R8591 gnd.n3132 gnd.n1750 19.3944
R8592 gnd.n3137 gnd.n1750 19.3944
R8593 gnd.n3137 gnd.n1751 19.3944
R8594 gnd.n1751 gnd.n1724 19.3944
R8595 gnd.n3168 gnd.n1724 19.3944
R8596 gnd.n3168 gnd.n1722 19.3944
R8597 gnd.n3172 gnd.n1722 19.3944
R8598 gnd.n3172 gnd.n1704 19.3944
R8599 gnd.n3198 gnd.n1704 19.3944
R8600 gnd.n3198 gnd.n1701 19.3944
R8601 gnd.n3203 gnd.n1701 19.3944
R8602 gnd.n3203 gnd.n1702 19.3944
R8603 gnd.n1702 gnd.n1673 19.3944
R8604 gnd.n3241 gnd.n1673 19.3944
R8605 gnd.n3241 gnd.n1670 19.3944
R8606 gnd.n3249 gnd.n1670 19.3944
R8607 gnd.n3249 gnd.n1671 19.3944
R8608 gnd.n3245 gnd.n1671 19.3944
R8609 gnd.n3245 gnd.n1642 19.3944
R8610 gnd.n3301 gnd.n1642 19.3944
R8611 gnd.n3301 gnd.n1639 19.3944
R8612 gnd.n3306 gnd.n1639 19.3944
R8613 gnd.n3306 gnd.n1640 19.3944
R8614 gnd.n1640 gnd.n1616 19.3944
R8615 gnd.n3344 gnd.n1616 19.3944
R8616 gnd.n3344 gnd.n1614 19.3944
R8617 gnd.n3348 gnd.n1614 19.3944
R8618 gnd.n3348 gnd.n1612 19.3944
R8619 gnd.n3354 gnd.n1612 19.3944
R8620 gnd.n3354 gnd.n1610 19.3944
R8621 gnd.n3358 gnd.n1610 19.3944
R8622 gnd.n3359 gnd.n3358 19.3944
R8623 gnd.n3362 gnd.n3359 19.3944
R8624 gnd.n3362 gnd.n1608 19.3944
R8625 gnd.n3366 gnd.n1608 19.3944
R8626 gnd.n3367 gnd.n3366 19.3944
R8627 gnd.n3373 gnd.n3367 19.3944
R8628 gnd.n3373 gnd.n1606 19.3944
R8629 gnd.n3377 gnd.n1606 19.3944
R8630 gnd.n3378 gnd.n3377 19.3944
R8631 gnd.n3381 gnd.n3378 19.3944
R8632 gnd.n3381 gnd.n1604 19.3944
R8633 gnd.n3385 gnd.n1604 19.3944
R8634 gnd.n3386 gnd.n3385 19.3944
R8635 gnd.n3389 gnd.n3386 19.3944
R8636 gnd.n3389 gnd.n1601 19.3944
R8637 gnd.n3569 gnd.n1601 19.3944
R8638 gnd.n3569 gnd.n1602 19.3944
R8639 gnd.n2562 gnd.n2561 19.3944
R8640 gnd.n2561 gnd.n2560 19.3944
R8641 gnd.n2560 gnd.n2558 19.3944
R8642 gnd.n2834 gnd.n2833 19.3944
R8643 gnd.n2833 gnd.n1983 19.3944
R8644 gnd.n2826 gnd.n1983 19.3944
R8645 gnd.n2826 gnd.n2825 19.3944
R8646 gnd.n2825 gnd.n1994 19.3944
R8647 gnd.n2818 gnd.n1994 19.3944
R8648 gnd.n2818 gnd.n2817 19.3944
R8649 gnd.n2817 gnd.n2002 19.3944
R8650 gnd.n2810 gnd.n2002 19.3944
R8651 gnd.n2810 gnd.n2809 19.3944
R8652 gnd.n2809 gnd.n2012 19.3944
R8653 gnd.n2802 gnd.n2012 19.3944
R8654 gnd.n2802 gnd.n2801 19.3944
R8655 gnd.n2801 gnd.n2020 19.3944
R8656 gnd.n2794 gnd.n2020 19.3944
R8657 gnd.n2794 gnd.n2793 19.3944
R8658 gnd.n2793 gnd.n2032 19.3944
R8659 gnd.n2573 gnd.n2032 19.3944
R8660 gnd.n2573 gnd.n2572 19.3944
R8661 gnd.n2572 gnd.n2571 19.3944
R8662 gnd.n2571 gnd.n2546 19.3944
R8663 gnd.n2567 gnd.n2546 19.3944
R8664 gnd.n2567 gnd.n2566 19.3944
R8665 gnd.n2566 gnd.n2565 19.3944
R8666 gnd.n5195 gnd.n5194 19.3944
R8667 gnd.n5194 gnd.n5104 19.3944
R8668 gnd.n5189 gnd.n5104 19.3944
R8669 gnd.n5189 gnd.n5188 19.3944
R8670 gnd.n5188 gnd.n5109 19.3944
R8671 gnd.n5183 gnd.n5109 19.3944
R8672 gnd.n5183 gnd.n5182 19.3944
R8673 gnd.n5182 gnd.n5181 19.3944
R8674 gnd.n5181 gnd.n5115 19.3944
R8675 gnd.n5175 gnd.n5115 19.3944
R8676 gnd.n5175 gnd.n5174 19.3944
R8677 gnd.n5174 gnd.n5173 19.3944
R8678 gnd.n5173 gnd.n5121 19.3944
R8679 gnd.n5167 gnd.n5121 19.3944
R8680 gnd.n5167 gnd.n5166 19.3944
R8681 gnd.n5166 gnd.n5165 19.3944
R8682 gnd.n5165 gnd.n5127 19.3944
R8683 gnd.n5159 gnd.n5127 19.3944
R8684 gnd.n5159 gnd.n5158 19.3944
R8685 gnd.n5158 gnd.n5157 19.3944
R8686 gnd.n5157 gnd.n5133 19.3944
R8687 gnd.n5151 gnd.n5133 19.3944
R8688 gnd.n5149 gnd.n5148 19.3944
R8689 gnd.n5148 gnd.n5143 19.3944
R8690 gnd.n5143 gnd.n5141 19.3944
R8691 gnd.n5808 gnd.n4522 19.3944
R8692 gnd.n5808 gnd.n5807 19.3944
R8693 gnd.n5807 gnd.n5806 19.3944
R8694 gnd.n5850 gnd.n5849 19.3944
R8695 gnd.n5849 gnd.n5848 19.3944
R8696 gnd.n5848 gnd.n4483 19.3944
R8697 gnd.n5843 gnd.n4483 19.3944
R8698 gnd.n5843 gnd.n5842 19.3944
R8699 gnd.n5842 gnd.n5841 19.3944
R8700 gnd.n5841 gnd.n4490 19.3944
R8701 gnd.n5836 gnd.n4490 19.3944
R8702 gnd.n5836 gnd.n5835 19.3944
R8703 gnd.n5835 gnd.n5834 19.3944
R8704 gnd.n5834 gnd.n4497 19.3944
R8705 gnd.n5829 gnd.n4497 19.3944
R8706 gnd.n5829 gnd.n5828 19.3944
R8707 gnd.n5828 gnd.n5827 19.3944
R8708 gnd.n5827 gnd.n4504 19.3944
R8709 gnd.n5822 gnd.n4504 19.3944
R8710 gnd.n5822 gnd.n5821 19.3944
R8711 gnd.n5821 gnd.n5820 19.3944
R8712 gnd.n5820 gnd.n4511 19.3944
R8713 gnd.n5815 gnd.n4511 19.3944
R8714 gnd.n5815 gnd.n5814 19.3944
R8715 gnd.n5814 gnd.n5813 19.3944
R8716 gnd.n5448 gnd.n5447 19.3944
R8717 gnd.n5448 gnd.n5044 19.3944
R8718 gnd.n5468 gnd.n5044 19.3944
R8719 gnd.n5468 gnd.n5036 19.3944
R8720 gnd.n5478 gnd.n5036 19.3944
R8721 gnd.n5479 gnd.n5478 19.3944
R8722 gnd.n5479 gnd.n5017 19.3944
R8723 gnd.n5499 gnd.n5017 19.3944
R8724 gnd.n5499 gnd.n5010 19.3944
R8725 gnd.n5509 gnd.n5010 19.3944
R8726 gnd.n5510 gnd.n5509 19.3944
R8727 gnd.n5510 gnd.n4991 19.3944
R8728 gnd.n5530 gnd.n4991 19.3944
R8729 gnd.n5530 gnd.n4984 19.3944
R8730 gnd.n5540 gnd.n4984 19.3944
R8731 gnd.n5541 gnd.n5540 19.3944
R8732 gnd.n5541 gnd.n4966 19.3944
R8733 gnd.n5561 gnd.n4966 19.3944
R8734 gnd.n5561 gnd.n4958 19.3944
R8735 gnd.n5571 gnd.n4958 19.3944
R8736 gnd.n5572 gnd.n5571 19.3944
R8737 gnd.n5572 gnd.n4941 19.3944
R8738 gnd.n5592 gnd.n4941 19.3944
R8739 gnd.n5592 gnd.n4933 19.3944
R8740 gnd.n5602 gnd.n4933 19.3944
R8741 gnd.n5603 gnd.n5602 19.3944
R8742 gnd.n5603 gnd.n4916 19.3944
R8743 gnd.n5623 gnd.n4916 19.3944
R8744 gnd.n5623 gnd.n4908 19.3944
R8745 gnd.n5633 gnd.n4908 19.3944
R8746 gnd.n5634 gnd.n5633 19.3944
R8747 gnd.n5634 gnd.n4892 19.3944
R8748 gnd.n5653 gnd.n4892 19.3944
R8749 gnd.n5653 gnd.n4877 19.3944
R8750 gnd.n5674 gnd.n4877 19.3944
R8751 gnd.n5675 gnd.n5674 19.3944
R8752 gnd.n5676 gnd.n5675 19.3944
R8753 gnd.n5676 gnd.n4861 19.3944
R8754 gnd.n4861 gnd.n4859 19.3944
R8755 gnd.n5699 gnd.n4859 19.3944
R8756 gnd.n5699 gnd.n4841 19.3944
R8757 gnd.n5725 gnd.n4841 19.3944
R8758 gnd.n5725 gnd.n5724 19.3944
R8759 gnd.n5724 gnd.n4830 19.3944
R8760 gnd.n5744 gnd.n4830 19.3944
R8761 gnd.n5744 gnd.n4814 19.3944
R8762 gnd.n5769 gnd.n4814 19.3944
R8763 gnd.n5769 gnd.n4794 19.3944
R8764 gnd.n5786 gnd.n4794 19.3944
R8765 gnd.n5786 gnd.n4796 19.3944
R8766 gnd.n4803 gnd.n4796 19.3944
R8767 gnd.n4803 gnd.n4802 19.3944
R8768 gnd.n4802 gnd.n4801 19.3944
R8769 gnd.n5431 gnd.n5430 19.3944
R8770 gnd.n5430 gnd.n5429 19.3944
R8771 gnd.n5429 gnd.n5428 19.3944
R8772 gnd.n5428 gnd.n5426 19.3944
R8773 gnd.n5426 gnd.n5423 19.3944
R8774 gnd.n5423 gnd.n5422 19.3944
R8775 gnd.n5422 gnd.n5419 19.3944
R8776 gnd.n5419 gnd.n5418 19.3944
R8777 gnd.n5418 gnd.n5415 19.3944
R8778 gnd.n5415 gnd.n5414 19.3944
R8779 gnd.n5414 gnd.n5411 19.3944
R8780 gnd.n5411 gnd.n5410 19.3944
R8781 gnd.n5410 gnd.n5407 19.3944
R8782 gnd.n5407 gnd.n5406 19.3944
R8783 gnd.n5458 gnd.n5051 19.3944
R8784 gnd.n5458 gnd.n5049 19.3944
R8785 gnd.n5464 gnd.n5049 19.3944
R8786 gnd.n5464 gnd.n5463 19.3944
R8787 gnd.n5463 gnd.n5026 19.3944
R8788 gnd.n5489 gnd.n5026 19.3944
R8789 gnd.n5489 gnd.n5024 19.3944
R8790 gnd.n5495 gnd.n5024 19.3944
R8791 gnd.n5495 gnd.n5494 19.3944
R8792 gnd.n5494 gnd.n5000 19.3944
R8793 gnd.n5520 gnd.n5000 19.3944
R8794 gnd.n5520 gnd.n4998 19.3944
R8795 gnd.n5526 gnd.n4998 19.3944
R8796 gnd.n5526 gnd.n5525 19.3944
R8797 gnd.n5525 gnd.n4974 19.3944
R8798 gnd.n5551 gnd.n4974 19.3944
R8799 gnd.n5551 gnd.n4972 19.3944
R8800 gnd.n5557 gnd.n4972 19.3944
R8801 gnd.n5557 gnd.n5556 19.3944
R8802 gnd.n5556 gnd.n4948 19.3944
R8803 gnd.n5582 gnd.n4948 19.3944
R8804 gnd.n5582 gnd.n4946 19.3944
R8805 gnd.n5588 gnd.n4946 19.3944
R8806 gnd.n5588 gnd.n5587 19.3944
R8807 gnd.n5587 gnd.n4923 19.3944
R8808 gnd.n5613 gnd.n4923 19.3944
R8809 gnd.n5613 gnd.n4921 19.3944
R8810 gnd.n5619 gnd.n4921 19.3944
R8811 gnd.n5619 gnd.n5618 19.3944
R8812 gnd.n5618 gnd.n4899 19.3944
R8813 gnd.n5643 gnd.n4899 19.3944
R8814 gnd.n5643 gnd.n4897 19.3944
R8815 gnd.n5649 gnd.n4897 19.3944
R8816 gnd.n5649 gnd.n5648 19.3944
R8817 gnd.n5648 gnd.n4867 19.3944
R8818 gnd.n5684 gnd.n4867 19.3944
R8819 gnd.n5684 gnd.n4865 19.3944
R8820 gnd.n5693 gnd.n4865 19.3944
R8821 gnd.n5693 gnd.n5692 19.3944
R8822 gnd.n5692 gnd.n5691 19.3944
R8823 gnd.n5691 gnd.n4837 19.3944
R8824 gnd.n5731 gnd.n4837 19.3944
R8825 gnd.n5731 gnd.n4835 19.3944
R8826 gnd.n5739 gnd.n4835 19.3944
R8827 gnd.n5739 gnd.n5738 19.3944
R8828 gnd.n5738 gnd.n5737 19.3944
R8829 gnd.n5737 gnd.n4810 19.3944
R8830 gnd.n5775 gnd.n4810 19.3944
R8831 gnd.n5775 gnd.n4808 19.3944
R8832 gnd.n5781 gnd.n4808 19.3944
R8833 gnd.n5781 gnd.n5780 19.3944
R8834 gnd.n5780 gnd.n4448 19.3944
R8835 gnd.n5885 gnd.n4448 19.3944
R8836 gnd.n5882 gnd.n5881 19.3944
R8837 gnd.n5881 gnd.n5880 19.3944
R8838 gnd.n5880 gnd.n4453 19.3944
R8839 gnd.n5875 gnd.n4453 19.3944
R8840 gnd.n5875 gnd.n5874 19.3944
R8841 gnd.n5874 gnd.n5873 19.3944
R8842 gnd.n5873 gnd.n4460 19.3944
R8843 gnd.n5868 gnd.n4460 19.3944
R8844 gnd.n5868 gnd.n5867 19.3944
R8845 gnd.n5867 gnd.n5866 19.3944
R8846 gnd.n5866 gnd.n4467 19.3944
R8847 gnd.n5861 gnd.n4467 19.3944
R8848 gnd.n5861 gnd.n5860 19.3944
R8849 gnd.n5860 gnd.n5859 19.3944
R8850 gnd.n5202 gnd.n5098 19.3944
R8851 gnd.n5206 gnd.n5098 19.3944
R8852 gnd.n5206 gnd.n5088 19.3944
R8853 gnd.n5218 gnd.n5088 19.3944
R8854 gnd.n5218 gnd.n5086 19.3944
R8855 gnd.n5222 gnd.n5086 19.3944
R8856 gnd.n5222 gnd.n5075 19.3944
R8857 gnd.n5234 gnd.n5075 19.3944
R8858 gnd.n5234 gnd.n5073 19.3944
R8859 gnd.n5373 gnd.n5073 19.3944
R8860 gnd.n5373 gnd.n5372 19.3944
R8861 gnd.n5372 gnd.n5371 19.3944
R8862 gnd.n5371 gnd.n5370 19.3944
R8863 gnd.n5370 gnd.n5368 19.3944
R8864 gnd.n5368 gnd.n5367 19.3944
R8865 gnd.n5367 gnd.n5363 19.3944
R8866 gnd.n5363 gnd.n5362 19.3944
R8867 gnd.n5362 gnd.n5361 19.3944
R8868 gnd.n5361 gnd.n5359 19.3944
R8869 gnd.n5359 gnd.n5358 19.3944
R8870 gnd.n5358 gnd.n5355 19.3944
R8871 gnd.n5355 gnd.n5354 19.3944
R8872 gnd.n5354 gnd.n5353 19.3944
R8873 gnd.n5353 gnd.n5351 19.3944
R8874 gnd.n5351 gnd.n5350 19.3944
R8875 gnd.n5350 gnd.n5347 19.3944
R8876 gnd.n5347 gnd.n5346 19.3944
R8877 gnd.n5346 gnd.n5345 19.3944
R8878 gnd.n5345 gnd.n5343 19.3944
R8879 gnd.n5291 gnd.n5256 19.3944
R8880 gnd.n5288 gnd.n5287 19.3944
R8881 gnd.n5284 gnd.n5283 19.3944
R8882 gnd.n5279 gnd.n5278 19.3944
R8883 gnd.n5278 gnd.n5277 19.3944
R8884 gnd.n5277 gnd.n5275 19.3944
R8885 gnd.n5275 gnd.n5274 19.3944
R8886 gnd.n5274 gnd.n5270 19.3944
R8887 gnd.n5270 gnd.n5269 19.3944
R8888 gnd.n5269 gnd.n5268 19.3944
R8889 gnd.n5268 gnd.n5266 19.3944
R8890 gnd.n5266 gnd.n4885 19.3944
R8891 gnd.n5663 gnd.n4885 19.3944
R8892 gnd.n5663 gnd.n4883 19.3944
R8893 gnd.n5669 gnd.n4883 19.3944
R8894 gnd.n5669 gnd.n5668 19.3944
R8895 gnd.n5668 gnd.n4850 19.3944
R8896 gnd.n5707 gnd.n4850 19.3944
R8897 gnd.n5707 gnd.n4848 19.3944
R8898 gnd.n5713 gnd.n4848 19.3944
R8899 gnd.n5713 gnd.n5712 19.3944
R8900 gnd.n5712 gnd.n4823 19.3944
R8901 gnd.n5752 gnd.n4823 19.3944
R8902 gnd.n5752 gnd.n4821 19.3944
R8903 gnd.n5758 gnd.n4821 19.3944
R8904 gnd.n5758 gnd.n5757 19.3944
R8905 gnd.n5757 gnd.n4530 19.3944
R8906 gnd.n5793 gnd.n4530 19.3944
R8907 gnd.n5793 gnd.n4528 19.3944
R8908 gnd.n5797 gnd.n4528 19.3944
R8909 gnd.n5800 gnd.n5797 19.3944
R8910 gnd.n5801 gnd.n5800 19.3944
R8911 gnd.n5198 gnd.n5094 19.3944
R8912 gnd.n5210 gnd.n5094 19.3944
R8913 gnd.n5210 gnd.n5092 19.3944
R8914 gnd.n5214 gnd.n5092 19.3944
R8915 gnd.n5214 gnd.n5082 19.3944
R8916 gnd.n5226 gnd.n5082 19.3944
R8917 gnd.n5226 gnd.n5080 19.3944
R8918 gnd.n5230 gnd.n5080 19.3944
R8919 gnd.n5230 gnd.n5069 19.3944
R8920 gnd.n5437 gnd.n5069 19.3944
R8921 gnd.n5437 gnd.n5066 19.3944
R8922 gnd.n5442 gnd.n5066 19.3944
R8923 gnd.n5442 gnd.n5059 19.3944
R8924 gnd.n5453 gnd.n5059 19.3944
R8925 gnd.n5453 gnd.n5452 19.3944
R8926 gnd.n5452 gnd.n5042 19.3944
R8927 gnd.n5473 gnd.n5042 19.3944
R8928 gnd.n5473 gnd.n5034 19.3944
R8929 gnd.n5484 gnd.n5034 19.3944
R8930 gnd.n5484 gnd.n5483 19.3944
R8931 gnd.n5483 gnd.n5015 19.3944
R8932 gnd.n5504 gnd.n5015 19.3944
R8933 gnd.n5504 gnd.n5008 19.3944
R8934 gnd.n5515 gnd.n5008 19.3944
R8935 gnd.n5515 gnd.n5514 19.3944
R8936 gnd.n5514 gnd.n4989 19.3944
R8937 gnd.n5535 gnd.n4989 19.3944
R8938 gnd.n5535 gnd.n4982 19.3944
R8939 gnd.n5546 gnd.n4982 19.3944
R8940 gnd.n5546 gnd.n5545 19.3944
R8941 gnd.n5545 gnd.n4964 19.3944
R8942 gnd.n5566 gnd.n4964 19.3944
R8943 gnd.n5566 gnd.n4956 19.3944
R8944 gnd.n5577 gnd.n4956 19.3944
R8945 gnd.n5577 gnd.n5576 19.3944
R8946 gnd.n5576 gnd.n4939 19.3944
R8947 gnd.n5597 gnd.n4939 19.3944
R8948 gnd.n5597 gnd.n4931 19.3944
R8949 gnd.n5608 gnd.n4931 19.3944
R8950 gnd.n5608 gnd.n5607 19.3944
R8951 gnd.n5607 gnd.n4914 19.3944
R8952 gnd.n5628 gnd.n4914 19.3944
R8953 gnd.n5628 gnd.n4906 19.3944
R8954 gnd.n5638 gnd.n4906 19.3944
R8955 gnd.n5638 gnd.n4890 19.3944
R8956 gnd.n5659 gnd.n4890 19.3944
R8957 gnd.n5659 gnd.n5658 19.3944
R8958 gnd.n5658 gnd.n4873 19.3944
R8959 gnd.n5679 gnd.n4873 19.3944
R8960 gnd.n5679 gnd.n4855 19.3944
R8961 gnd.n5703 gnd.n4855 19.3944
R8962 gnd.n5703 gnd.n5702 19.3944
R8963 gnd.n5702 gnd.n4843 19.3944
R8964 gnd.n5719 gnd.n4843 19.3944
R8965 gnd.n5719 gnd.n4826 19.3944
R8966 gnd.n5748 gnd.n4826 19.3944
R8967 gnd.n5748 gnd.n5747 19.3944
R8968 gnd.n5747 gnd.n4816 19.3944
R8969 gnd.n5764 gnd.n4816 19.3944
R8970 gnd.n5764 gnd.n4536 19.3944
R8971 gnd.n5789 gnd.n4536 19.3944
R8972 gnd.n5789 gnd.n849 19.3944
R8973 gnd.n5892 gnd.n849 19.3944
R8974 gnd.n5892 gnd.n5891 19.3944
R8975 gnd.n5891 gnd.n5890 19.3944
R8976 gnd.n3907 gnd.n1460 19.3944
R8977 gnd.n3907 gnd.n1457 19.3944
R8978 gnd.n3911 gnd.n1457 19.3944
R8979 gnd.n3912 gnd.n3911 19.3944
R8980 gnd.n3914 gnd.n3912 19.3944
R8981 gnd.n3914 gnd.n1454 19.3944
R8982 gnd.n3919 gnd.n1454 19.3944
R8983 gnd.n3919 gnd.n1455 19.3944
R8984 gnd.n1455 gnd.n1395 19.3944
R8985 gnd.n3979 gnd.n1395 19.3944
R8986 gnd.n3979 gnd.n1392 19.3944
R8987 gnd.n3983 gnd.n1392 19.3944
R8988 gnd.n3984 gnd.n3983 19.3944
R8989 gnd.n3986 gnd.n3984 19.3944
R8990 gnd.n3986 gnd.n1389 19.3944
R8991 gnd.n3991 gnd.n1389 19.3944
R8992 gnd.n3991 gnd.n1390 19.3944
R8993 gnd.n1390 gnd.n310 19.3944
R8994 gnd.n6664 gnd.n310 19.3944
R8995 gnd.n6664 gnd.n307 19.3944
R8996 gnd.n6668 gnd.n307 19.3944
R8997 gnd.n6669 gnd.n6668 19.3944
R8998 gnd.n6671 gnd.n6669 19.3944
R8999 gnd.n6671 gnd.n305 19.3944
R9000 gnd.n6675 gnd.n305 19.3944
R9001 gnd.n6675 gnd.n65 19.3944
R9002 gnd.n7054 gnd.n65 19.3944
R9003 gnd.n7054 gnd.n7053 19.3944
R9004 gnd.n7053 gnd.n7052 19.3944
R9005 gnd.n7052 gnd.n69 19.3944
R9006 gnd.n7048 gnd.n69 19.3944
R9007 gnd.n7048 gnd.n7047 19.3944
R9008 gnd.n7047 gnd.n7046 19.3944
R9009 gnd.n7046 gnd.n74 19.3944
R9010 gnd.n7042 gnd.n74 19.3944
R9011 gnd.n7042 gnd.n7041 19.3944
R9012 gnd.n7041 gnd.n7040 19.3944
R9013 gnd.n7040 gnd.n79 19.3944
R9014 gnd.n7036 gnd.n79 19.3944
R9015 gnd.n7036 gnd.n7035 19.3944
R9016 gnd.n7035 gnd.n7034 19.3944
R9017 gnd.n7034 gnd.n84 19.3944
R9018 gnd.n7030 gnd.n84 19.3944
R9019 gnd.n7030 gnd.n7029 19.3944
R9020 gnd.n7029 gnd.n7028 19.3944
R9021 gnd.n7028 gnd.n89 19.3944
R9022 gnd.n7024 gnd.n89 19.3944
R9023 gnd.n7024 gnd.n7023 19.3944
R9024 gnd.n7023 gnd.n7022 19.3944
R9025 gnd.n7022 gnd.n94 19.3944
R9026 gnd.n7018 gnd.n94 19.3944
R9027 gnd.n7018 gnd.n7017 19.3944
R9028 gnd.n7017 gnd.n7016 19.3944
R9029 gnd.n6915 gnd.n6914 19.3944
R9030 gnd.n6914 gnd.n6913 19.3944
R9031 gnd.n6913 gnd.n6855 19.3944
R9032 gnd.n6909 gnd.n6855 19.3944
R9033 gnd.n6909 gnd.n6908 19.3944
R9034 gnd.n6908 gnd.n6907 19.3944
R9035 gnd.n6907 gnd.n6863 19.3944
R9036 gnd.n6903 gnd.n6863 19.3944
R9037 gnd.n6903 gnd.n6902 19.3944
R9038 gnd.n6902 gnd.n6901 19.3944
R9039 gnd.n6901 gnd.n6871 19.3944
R9040 gnd.n6897 gnd.n6871 19.3944
R9041 gnd.n6897 gnd.n6896 19.3944
R9042 gnd.n6896 gnd.n6895 19.3944
R9043 gnd.n6895 gnd.n6879 19.3944
R9044 gnd.n6891 gnd.n6879 19.3944
R9045 gnd.n3449 gnd.n3443 19.3944
R9046 gnd.n3455 gnd.n3443 19.3944
R9047 gnd.n3455 gnd.n3436 19.3944
R9048 gnd.n3468 gnd.n3436 19.3944
R9049 gnd.n3468 gnd.n3434 19.3944
R9050 gnd.n3474 gnd.n3434 19.3944
R9051 gnd.n3474 gnd.n3427 19.3944
R9052 gnd.n3487 gnd.n3427 19.3944
R9053 gnd.n3487 gnd.n3425 19.3944
R9054 gnd.n3493 gnd.n3425 19.3944
R9055 gnd.n3493 gnd.n3418 19.3944
R9056 gnd.n3506 gnd.n3418 19.3944
R9057 gnd.n3506 gnd.n3416 19.3944
R9058 gnd.n3512 gnd.n3416 19.3944
R9059 gnd.n3512 gnd.n3409 19.3944
R9060 gnd.n3527 gnd.n3409 19.3944
R9061 gnd.n3446 gnd.n1342 19.3944
R9062 gnd.n4051 gnd.n1342 19.3944
R9063 gnd.n4051 gnd.n1343 19.3944
R9064 gnd.n4047 gnd.n1343 19.3944
R9065 gnd.n4047 gnd.n4046 19.3944
R9066 gnd.n4046 gnd.n4045 19.3944
R9067 gnd.n4045 gnd.n1349 19.3944
R9068 gnd.n4041 gnd.n1349 19.3944
R9069 gnd.n4041 gnd.n4040 19.3944
R9070 gnd.n4040 gnd.n4039 19.3944
R9071 gnd.n4039 gnd.n1354 19.3944
R9072 gnd.n4035 gnd.n1354 19.3944
R9073 gnd.n4035 gnd.n4034 19.3944
R9074 gnd.n4034 gnd.n4033 19.3944
R9075 gnd.n4033 gnd.n4030 19.3944
R9076 gnd.n4030 gnd.n328 19.3944
R9077 gnd.n6650 gnd.n328 19.3944
R9078 gnd.n6650 gnd.n329 19.3944
R9079 gnd.n6646 gnd.n329 19.3944
R9080 gnd.n6646 gnd.n6645 19.3944
R9081 gnd.n6645 gnd.n274 19.3944
R9082 gnd.n6770 gnd.n274 19.3944
R9083 gnd.n6770 gnd.n275 19.3944
R9084 gnd.n6766 gnd.n275 19.3944
R9085 gnd.n6766 gnd.n6765 19.3944
R9086 gnd.n6765 gnd.n6764 19.3944
R9087 gnd.n6764 gnd.n281 19.3944
R9088 gnd.n6759 gnd.n281 19.3944
R9089 gnd.n6759 gnd.n6758 19.3944
R9090 gnd.n6758 gnd.n254 19.3944
R9091 gnd.n6781 gnd.n254 19.3944
R9092 gnd.n6781 gnd.n252 19.3944
R9093 gnd.n6785 gnd.n252 19.3944
R9094 gnd.n6785 gnd.n239 19.3944
R9095 gnd.n6797 gnd.n239 19.3944
R9096 gnd.n6797 gnd.n237 19.3944
R9097 gnd.n6801 gnd.n237 19.3944
R9098 gnd.n6801 gnd.n224 19.3944
R9099 gnd.n6813 gnd.n224 19.3944
R9100 gnd.n6813 gnd.n222 19.3944
R9101 gnd.n6817 gnd.n222 19.3944
R9102 gnd.n6817 gnd.n209 19.3944
R9103 gnd.n6829 gnd.n209 19.3944
R9104 gnd.n6829 gnd.n207 19.3944
R9105 gnd.n6833 gnd.n207 19.3944
R9106 gnd.n6833 gnd.n195 19.3944
R9107 gnd.n6845 gnd.n195 19.3944
R9108 gnd.n6845 gnd.n192 19.3944
R9109 gnd.n6924 gnd.n192 19.3944
R9110 gnd.n6924 gnd.n193 19.3944
R9111 gnd.n6920 gnd.n193 19.3944
R9112 gnd.n6920 gnd.n6919 19.3944
R9113 gnd.n6919 gnd.n6918 19.3944
R9114 gnd.n2036 gnd.n1197 19.3944
R9115 gnd.n2036 gnd.n1986 19.3944
R9116 gnd.n2830 gnd.n1986 19.3944
R9117 gnd.n2830 gnd.n2829 19.3944
R9118 gnd.n2829 gnd.n1989 19.3944
R9119 gnd.n2822 gnd.n1989 19.3944
R9120 gnd.n2822 gnd.n2821 19.3944
R9121 gnd.n2821 gnd.n1998 19.3944
R9122 gnd.n2814 gnd.n1998 19.3944
R9123 gnd.n2814 gnd.n2813 19.3944
R9124 gnd.n2813 gnd.n2006 19.3944
R9125 gnd.n2806 gnd.n2006 19.3944
R9126 gnd.n2806 gnd.n2805 19.3944
R9127 gnd.n2805 gnd.n2016 19.3944
R9128 gnd.n2798 gnd.n2016 19.3944
R9129 gnd.n2798 gnd.n2797 19.3944
R9130 gnd.n2166 gnd.n2162 19.3944
R9131 gnd.n2166 gnd.n2158 19.3944
R9132 gnd.n2181 gnd.n2158 19.3944
R9133 gnd.n2181 gnd.n2180 19.3944
R9134 gnd.n2180 gnd.n2179 19.3944
R9135 gnd.n2179 gnd.n2176 19.3944
R9136 gnd.n2176 gnd.n2175 19.3944
R9137 gnd.n2175 gnd.n2138 19.3944
R9138 gnd.n2138 gnd.n2136 19.3944
R9139 gnd.n2478 gnd.n2136 19.3944
R9140 gnd.n2478 gnd.n2134 19.3944
R9141 gnd.n2482 gnd.n2134 19.3944
R9142 gnd.n2482 gnd.n2132 19.3944
R9143 gnd.n2486 gnd.n2132 19.3944
R9144 gnd.n2486 gnd.n2130 19.3944
R9145 gnd.n2516 gnd.n2130 19.3944
R9146 gnd.n2516 gnd.n2515 19.3944
R9147 gnd.n2515 gnd.n2514 19.3944
R9148 gnd.n2514 gnd.n2492 19.3944
R9149 gnd.n2510 gnd.n2492 19.3944
R9150 gnd.n2510 gnd.n2509 19.3944
R9151 gnd.n2509 gnd.n2508 19.3944
R9152 gnd.n2508 gnd.n2498 19.3944
R9153 gnd.n2504 gnd.n2498 19.3944
R9154 gnd.n2504 gnd.n2503 19.3944
R9155 gnd.n2503 gnd.n1964 19.3944
R9156 gnd.n2840 gnd.n1964 19.3944
R9157 gnd.n2840 gnd.n1962 19.3944
R9158 gnd.n2844 gnd.n1962 19.3944
R9159 gnd.n2844 gnd.n1953 19.3944
R9160 gnd.n2860 gnd.n1953 19.3944
R9161 gnd.n2860 gnd.n1951 19.3944
R9162 gnd.n2864 gnd.n1951 19.3944
R9163 gnd.n2864 gnd.n1940 19.3944
R9164 gnd.n2880 gnd.n1940 19.3944
R9165 gnd.n2880 gnd.n1938 19.3944
R9166 gnd.n2884 gnd.n1938 19.3944
R9167 gnd.n2884 gnd.n1927 19.3944
R9168 gnd.n2900 gnd.n1927 19.3944
R9169 gnd.n2900 gnd.n1925 19.3944
R9170 gnd.n2904 gnd.n1925 19.3944
R9171 gnd.n2904 gnd.n1914 19.3944
R9172 gnd.n2920 gnd.n1914 19.3944
R9173 gnd.n2920 gnd.n1912 19.3944
R9174 gnd.n2924 gnd.n1912 19.3944
R9175 gnd.n2924 gnd.n1899 19.3944
R9176 gnd.n2958 gnd.n1899 19.3944
R9177 gnd.n2958 gnd.n1897 19.3944
R9178 gnd.n2962 gnd.n1897 19.3944
R9179 gnd.n2962 gnd.n1824 19.3944
R9180 gnd.n2985 gnd.n1824 19.3944
R9181 gnd.n2985 gnd.n1822 19.3944
R9182 gnd.n2994 gnd.n1822 19.3944
R9183 gnd.n2994 gnd.n2993 19.3944
R9184 gnd.n2993 gnd.n2992 19.3944
R9185 gnd.n2992 gnd.n1787 19.3944
R9186 gnd.n3046 gnd.n1787 19.3944
R9187 gnd.n3046 gnd.n1785 19.3944
R9188 gnd.n3050 gnd.n1785 19.3944
R9189 gnd.n3050 gnd.n1767 19.3944
R9190 gnd.n3113 gnd.n1767 19.3944
R9191 gnd.n3113 gnd.n1765 19.3944
R9192 gnd.n3119 gnd.n1765 19.3944
R9193 gnd.n3119 gnd.n3118 19.3944
R9194 gnd.n3118 gnd.n1738 19.3944
R9195 gnd.n3149 gnd.n1738 19.3944
R9196 gnd.n3149 gnd.n1736 19.3944
R9197 gnd.n3153 gnd.n1736 19.3944
R9198 gnd.n3153 gnd.n1717 19.3944
R9199 gnd.n3177 gnd.n1717 19.3944
R9200 gnd.n3177 gnd.n1715 19.3944
R9201 gnd.n3183 gnd.n1715 19.3944
R9202 gnd.n3183 gnd.n3182 19.3944
R9203 gnd.n3182 gnd.n1689 19.3944
R9204 gnd.n3216 gnd.n1689 19.3944
R9205 gnd.n3216 gnd.n1687 19.3944
R9206 gnd.n3228 gnd.n1687 19.3944
R9207 gnd.n3228 gnd.n3227 19.3944
R9208 gnd.n3227 gnd.n3226 19.3944
R9209 gnd.n3226 gnd.n1657 19.3944
R9210 gnd.n3283 gnd.n1657 19.3944
R9211 gnd.n3283 gnd.n1655 19.3944
R9212 gnd.n3287 gnd.n1655 19.3944
R9213 gnd.n3287 gnd.n1634 19.3944
R9214 gnd.n3312 gnd.n1634 19.3944
R9215 gnd.n3312 gnd.n1632 19.3944
R9216 gnd.n3319 gnd.n1632 19.3944
R9217 gnd.n3319 gnd.n3318 19.3944
R9218 gnd.n3318 gnd.n1539 19.3944
R9219 gnd.n3619 gnd.n1539 19.3944
R9220 gnd.n3619 gnd.n3618 19.3944
R9221 gnd.n3618 gnd.n3617 19.3944
R9222 gnd.n3617 gnd.n1543 19.3944
R9223 gnd.n1551 gnd.n1543 19.3944
R9224 gnd.n3608 gnd.n1551 19.3944
R9225 gnd.n3608 gnd.n3607 19.3944
R9226 gnd.n3607 gnd.n3606 19.3944
R9227 gnd.n3606 gnd.n1557 19.3944
R9228 gnd.n3598 gnd.n1557 19.3944
R9229 gnd.n3598 gnd.n3597 19.3944
R9230 gnd.n3597 gnd.n3596 19.3944
R9231 gnd.n3596 gnd.n1570 19.3944
R9232 gnd.n3588 gnd.n1570 19.3944
R9233 gnd.n3588 gnd.n3587 19.3944
R9234 gnd.n3587 gnd.n3586 19.3944
R9235 gnd.n3586 gnd.n1580 19.3944
R9236 gnd.n3578 gnd.n1580 19.3944
R9237 gnd.n3578 gnd.n3577 19.3944
R9238 gnd.n3577 gnd.n3576 19.3944
R9239 gnd.n3576 gnd.n1595 19.3944
R9240 gnd.n1595 gnd.n1309 19.3944
R9241 gnd.n4072 gnd.n1309 19.3944
R9242 gnd.n4072 gnd.n4071 19.3944
R9243 gnd.n4071 gnd.n4070 19.3944
R9244 gnd.n4070 gnd.n1313 19.3944
R9245 gnd.n4064 gnd.n1313 19.3944
R9246 gnd.n4064 gnd.n4063 19.3944
R9247 gnd.n4063 gnd.n4062 19.3944
R9248 gnd.n4062 gnd.n1322 19.3944
R9249 gnd.n1444 gnd.n1322 19.3944
R9250 gnd.n1447 gnd.n1444 19.3944
R9251 gnd.n1447 gnd.n1441 19.3944
R9252 gnd.n3927 gnd.n1441 19.3944
R9253 gnd.n3927 gnd.n3926 19.3944
R9254 gnd.n3926 gnd.n3925 19.3944
R9255 gnd.n3925 gnd.n1413 19.3944
R9256 gnd.n3964 gnd.n1413 19.3944
R9257 gnd.n3964 gnd.n3963 19.3944
R9258 gnd.n3963 gnd.n3962 19.3944
R9259 gnd.n3962 gnd.n1419 19.3944
R9260 gnd.n1419 gnd.n1374 19.3944
R9261 gnd.n4017 gnd.n1374 19.3944
R9262 gnd.n4017 gnd.n4016 19.3944
R9263 gnd.n4016 gnd.n4015 19.3944
R9264 gnd.n4015 gnd.n1378 19.3944
R9265 gnd.n1385 gnd.n1378 19.3944
R9266 gnd.n1385 gnd.n1384 19.3944
R9267 gnd.n1384 gnd.n336 19.3944
R9268 gnd.n6640 gnd.n336 19.3944
R9269 gnd.n6640 gnd.n6639 19.3944
R9270 gnd.n6639 gnd.n6636 19.3944
R9271 gnd.n6421 gnd.n461 19.3944
R9272 gnd.n6427 gnd.n461 19.3944
R9273 gnd.n6427 gnd.n459 19.3944
R9274 gnd.n6431 gnd.n459 19.3944
R9275 gnd.n6431 gnd.n455 19.3944
R9276 gnd.n6437 gnd.n455 19.3944
R9277 gnd.n6437 gnd.n453 19.3944
R9278 gnd.n6441 gnd.n453 19.3944
R9279 gnd.n6441 gnd.n449 19.3944
R9280 gnd.n6447 gnd.n449 19.3944
R9281 gnd.n6447 gnd.n447 19.3944
R9282 gnd.n6451 gnd.n447 19.3944
R9283 gnd.n6451 gnd.n443 19.3944
R9284 gnd.n6457 gnd.n443 19.3944
R9285 gnd.n6457 gnd.n441 19.3944
R9286 gnd.n6461 gnd.n441 19.3944
R9287 gnd.n6461 gnd.n437 19.3944
R9288 gnd.n6467 gnd.n437 19.3944
R9289 gnd.n6467 gnd.n435 19.3944
R9290 gnd.n6471 gnd.n435 19.3944
R9291 gnd.n6471 gnd.n431 19.3944
R9292 gnd.n6477 gnd.n431 19.3944
R9293 gnd.n6477 gnd.n429 19.3944
R9294 gnd.n6481 gnd.n429 19.3944
R9295 gnd.n6481 gnd.n425 19.3944
R9296 gnd.n6487 gnd.n425 19.3944
R9297 gnd.n6487 gnd.n423 19.3944
R9298 gnd.n6491 gnd.n423 19.3944
R9299 gnd.n6491 gnd.n419 19.3944
R9300 gnd.n6497 gnd.n419 19.3944
R9301 gnd.n6497 gnd.n417 19.3944
R9302 gnd.n6501 gnd.n417 19.3944
R9303 gnd.n6501 gnd.n413 19.3944
R9304 gnd.n6507 gnd.n413 19.3944
R9305 gnd.n6507 gnd.n411 19.3944
R9306 gnd.n6511 gnd.n411 19.3944
R9307 gnd.n6511 gnd.n407 19.3944
R9308 gnd.n6517 gnd.n407 19.3944
R9309 gnd.n6517 gnd.n405 19.3944
R9310 gnd.n6521 gnd.n405 19.3944
R9311 gnd.n6521 gnd.n401 19.3944
R9312 gnd.n6527 gnd.n401 19.3944
R9313 gnd.n6527 gnd.n399 19.3944
R9314 gnd.n6531 gnd.n399 19.3944
R9315 gnd.n6531 gnd.n395 19.3944
R9316 gnd.n6537 gnd.n395 19.3944
R9317 gnd.n6537 gnd.n393 19.3944
R9318 gnd.n6541 gnd.n393 19.3944
R9319 gnd.n6541 gnd.n389 19.3944
R9320 gnd.n6547 gnd.n389 19.3944
R9321 gnd.n6547 gnd.n387 19.3944
R9322 gnd.n6551 gnd.n387 19.3944
R9323 gnd.n6551 gnd.n383 19.3944
R9324 gnd.n6557 gnd.n383 19.3944
R9325 gnd.n6557 gnd.n381 19.3944
R9326 gnd.n6561 gnd.n381 19.3944
R9327 gnd.n6561 gnd.n377 19.3944
R9328 gnd.n6567 gnd.n377 19.3944
R9329 gnd.n6567 gnd.n375 19.3944
R9330 gnd.n6571 gnd.n375 19.3944
R9331 gnd.n6571 gnd.n371 19.3944
R9332 gnd.n6577 gnd.n371 19.3944
R9333 gnd.n6577 gnd.n369 19.3944
R9334 gnd.n6581 gnd.n369 19.3944
R9335 gnd.n6581 gnd.n365 19.3944
R9336 gnd.n6587 gnd.n365 19.3944
R9337 gnd.n6587 gnd.n363 19.3944
R9338 gnd.n6591 gnd.n363 19.3944
R9339 gnd.n6591 gnd.n359 19.3944
R9340 gnd.n6597 gnd.n359 19.3944
R9341 gnd.n6597 gnd.n357 19.3944
R9342 gnd.n6601 gnd.n357 19.3944
R9343 gnd.n6601 gnd.n353 19.3944
R9344 gnd.n6607 gnd.n353 19.3944
R9345 gnd.n6607 gnd.n351 19.3944
R9346 gnd.n6611 gnd.n351 19.3944
R9347 gnd.n6611 gnd.n347 19.3944
R9348 gnd.n6617 gnd.n347 19.3944
R9349 gnd.n6617 gnd.n345 19.3944
R9350 gnd.n6621 gnd.n345 19.3944
R9351 gnd.n6621 gnd.n341 19.3944
R9352 gnd.n6628 gnd.n341 19.3944
R9353 gnd.n6628 gnd.n339 19.3944
R9354 gnd.n6632 gnd.n339 19.3944
R9355 gnd.n6066 gnd.n674 19.3944
R9356 gnd.n6070 gnd.n674 19.3944
R9357 gnd.n6070 gnd.n670 19.3944
R9358 gnd.n6076 gnd.n670 19.3944
R9359 gnd.n6076 gnd.n668 19.3944
R9360 gnd.n6080 gnd.n668 19.3944
R9361 gnd.n6080 gnd.n664 19.3944
R9362 gnd.n6086 gnd.n664 19.3944
R9363 gnd.n6086 gnd.n662 19.3944
R9364 gnd.n6090 gnd.n662 19.3944
R9365 gnd.n6090 gnd.n658 19.3944
R9366 gnd.n6096 gnd.n658 19.3944
R9367 gnd.n6096 gnd.n656 19.3944
R9368 gnd.n6100 gnd.n656 19.3944
R9369 gnd.n6100 gnd.n652 19.3944
R9370 gnd.n6106 gnd.n652 19.3944
R9371 gnd.n6106 gnd.n650 19.3944
R9372 gnd.n6110 gnd.n650 19.3944
R9373 gnd.n6110 gnd.n646 19.3944
R9374 gnd.n6116 gnd.n646 19.3944
R9375 gnd.n6116 gnd.n644 19.3944
R9376 gnd.n6120 gnd.n644 19.3944
R9377 gnd.n6120 gnd.n640 19.3944
R9378 gnd.n6126 gnd.n640 19.3944
R9379 gnd.n6126 gnd.n638 19.3944
R9380 gnd.n6130 gnd.n638 19.3944
R9381 gnd.n6130 gnd.n634 19.3944
R9382 gnd.n6136 gnd.n634 19.3944
R9383 gnd.n6136 gnd.n632 19.3944
R9384 gnd.n6140 gnd.n632 19.3944
R9385 gnd.n6140 gnd.n628 19.3944
R9386 gnd.n6146 gnd.n628 19.3944
R9387 gnd.n6146 gnd.n626 19.3944
R9388 gnd.n6150 gnd.n626 19.3944
R9389 gnd.n6150 gnd.n622 19.3944
R9390 gnd.n6156 gnd.n622 19.3944
R9391 gnd.n6156 gnd.n620 19.3944
R9392 gnd.n6160 gnd.n620 19.3944
R9393 gnd.n6160 gnd.n616 19.3944
R9394 gnd.n6166 gnd.n616 19.3944
R9395 gnd.n6166 gnd.n614 19.3944
R9396 gnd.n6170 gnd.n614 19.3944
R9397 gnd.n6170 gnd.n610 19.3944
R9398 gnd.n6176 gnd.n610 19.3944
R9399 gnd.n6176 gnd.n608 19.3944
R9400 gnd.n6180 gnd.n608 19.3944
R9401 gnd.n6180 gnd.n604 19.3944
R9402 gnd.n6186 gnd.n604 19.3944
R9403 gnd.n6186 gnd.n602 19.3944
R9404 gnd.n6190 gnd.n602 19.3944
R9405 gnd.n6190 gnd.n598 19.3944
R9406 gnd.n6196 gnd.n598 19.3944
R9407 gnd.n6196 gnd.n596 19.3944
R9408 gnd.n6200 gnd.n596 19.3944
R9409 gnd.n6200 gnd.n592 19.3944
R9410 gnd.n6206 gnd.n592 19.3944
R9411 gnd.n6206 gnd.n590 19.3944
R9412 gnd.n6210 gnd.n590 19.3944
R9413 gnd.n6210 gnd.n586 19.3944
R9414 gnd.n6216 gnd.n586 19.3944
R9415 gnd.n6216 gnd.n584 19.3944
R9416 gnd.n6220 gnd.n584 19.3944
R9417 gnd.n6220 gnd.n580 19.3944
R9418 gnd.n6226 gnd.n580 19.3944
R9419 gnd.n6226 gnd.n578 19.3944
R9420 gnd.n6230 gnd.n578 19.3944
R9421 gnd.n6230 gnd.n574 19.3944
R9422 gnd.n6236 gnd.n574 19.3944
R9423 gnd.n6236 gnd.n572 19.3944
R9424 gnd.n6240 gnd.n572 19.3944
R9425 gnd.n6240 gnd.n568 19.3944
R9426 gnd.n6246 gnd.n568 19.3944
R9427 gnd.n6246 gnd.n566 19.3944
R9428 gnd.n6250 gnd.n566 19.3944
R9429 gnd.n6250 gnd.n562 19.3944
R9430 gnd.n6256 gnd.n562 19.3944
R9431 gnd.n6256 gnd.n560 19.3944
R9432 gnd.n6260 gnd.n560 19.3944
R9433 gnd.n6260 gnd.n556 19.3944
R9434 gnd.n6266 gnd.n556 19.3944
R9435 gnd.n6266 gnd.n554 19.3944
R9436 gnd.n6270 gnd.n554 19.3944
R9437 gnd.n6270 gnd.n550 19.3944
R9438 gnd.n6276 gnd.n550 19.3944
R9439 gnd.n6276 gnd.n548 19.3944
R9440 gnd.n6280 gnd.n548 19.3944
R9441 gnd.n6280 gnd.n544 19.3944
R9442 gnd.n6286 gnd.n544 19.3944
R9443 gnd.n6286 gnd.n542 19.3944
R9444 gnd.n6290 gnd.n542 19.3944
R9445 gnd.n6290 gnd.n538 19.3944
R9446 gnd.n6296 gnd.n538 19.3944
R9447 gnd.n6296 gnd.n536 19.3944
R9448 gnd.n6300 gnd.n536 19.3944
R9449 gnd.n6300 gnd.n532 19.3944
R9450 gnd.n6306 gnd.n532 19.3944
R9451 gnd.n6306 gnd.n530 19.3944
R9452 gnd.n6310 gnd.n530 19.3944
R9453 gnd.n6310 gnd.n526 19.3944
R9454 gnd.n6316 gnd.n526 19.3944
R9455 gnd.n6316 gnd.n524 19.3944
R9456 gnd.n6320 gnd.n524 19.3944
R9457 gnd.n6320 gnd.n520 19.3944
R9458 gnd.n6326 gnd.n520 19.3944
R9459 gnd.n6326 gnd.n518 19.3944
R9460 gnd.n6330 gnd.n518 19.3944
R9461 gnd.n6330 gnd.n514 19.3944
R9462 gnd.n6336 gnd.n514 19.3944
R9463 gnd.n6336 gnd.n512 19.3944
R9464 gnd.n6340 gnd.n512 19.3944
R9465 gnd.n6340 gnd.n508 19.3944
R9466 gnd.n6346 gnd.n508 19.3944
R9467 gnd.n6346 gnd.n506 19.3944
R9468 gnd.n6350 gnd.n506 19.3944
R9469 gnd.n6350 gnd.n502 19.3944
R9470 gnd.n6356 gnd.n502 19.3944
R9471 gnd.n6356 gnd.n500 19.3944
R9472 gnd.n6360 gnd.n500 19.3944
R9473 gnd.n6360 gnd.n496 19.3944
R9474 gnd.n6366 gnd.n496 19.3944
R9475 gnd.n6366 gnd.n494 19.3944
R9476 gnd.n6370 gnd.n494 19.3944
R9477 gnd.n6370 gnd.n490 19.3944
R9478 gnd.n6376 gnd.n490 19.3944
R9479 gnd.n6376 gnd.n488 19.3944
R9480 gnd.n6380 gnd.n488 19.3944
R9481 gnd.n6380 gnd.n484 19.3944
R9482 gnd.n6386 gnd.n484 19.3944
R9483 gnd.n6386 gnd.n482 19.3944
R9484 gnd.n6390 gnd.n482 19.3944
R9485 gnd.n6390 gnd.n478 19.3944
R9486 gnd.n6396 gnd.n478 19.3944
R9487 gnd.n6396 gnd.n476 19.3944
R9488 gnd.n6400 gnd.n476 19.3944
R9489 gnd.n6400 gnd.n472 19.3944
R9490 gnd.n6406 gnd.n472 19.3944
R9491 gnd.n6406 gnd.n470 19.3944
R9492 gnd.n6411 gnd.n470 19.3944
R9493 gnd.n6411 gnd.n466 19.3944
R9494 gnd.n6417 gnd.n466 19.3944
R9495 gnd.n6418 gnd.n6417 19.3944
R9496 gnd.n3800 gnd.n3797 19.3944
R9497 gnd.n3800 gnd.n3796 19.3944
R9498 gnd.n3806 gnd.n3796 19.3944
R9499 gnd.n3806 gnd.n3794 19.3944
R9500 gnd.n3810 gnd.n3794 19.3944
R9501 gnd.n3810 gnd.n3792 19.3944
R9502 gnd.n3816 gnd.n3792 19.3944
R9503 gnd.n3816 gnd.n3790 19.3944
R9504 gnd.n3820 gnd.n3790 19.3944
R9505 gnd.n3820 gnd.n3788 19.3944
R9506 gnd.n3826 gnd.n3788 19.3944
R9507 gnd.n3826 gnd.n3786 19.3944
R9508 gnd.n3831 gnd.n3786 19.3944
R9509 gnd.n3831 gnd.n3784 19.3944
R9510 gnd.n3784 gnd.n1487 19.3944
R9511 gnd.n3844 gnd.n1485 19.3944
R9512 gnd.n3844 gnd.n1483 19.3944
R9513 gnd.n3850 gnd.n1483 19.3944
R9514 gnd.n3850 gnd.n1481 19.3944
R9515 gnd.n3854 gnd.n1481 19.3944
R9516 gnd.n3854 gnd.n1479 19.3944
R9517 gnd.n3860 gnd.n1479 19.3944
R9518 gnd.n3860 gnd.n1477 19.3944
R9519 gnd.n3864 gnd.n1477 19.3944
R9520 gnd.n3864 gnd.n1475 19.3944
R9521 gnd.n3870 gnd.n1475 19.3944
R9522 gnd.n3870 gnd.n1473 19.3944
R9523 gnd.n3874 gnd.n1473 19.3944
R9524 gnd.n3874 gnd.n1471 19.3944
R9525 gnd.n3880 gnd.n1471 19.3944
R9526 gnd.n3880 gnd.n1469 19.3944
R9527 gnd.n3885 gnd.n1469 19.3944
R9528 gnd.n3885 gnd.n1467 19.3944
R9529 gnd.n3903 gnd.n1461 19.3944
R9530 gnd.n3903 gnd.n1462 19.3944
R9531 gnd.n3899 gnd.n1462 19.3944
R9532 gnd.n3899 gnd.n3896 19.3944
R9533 gnd.n3896 gnd.n1427 19.3944
R9534 gnd.n3940 gnd.n1427 19.3944
R9535 gnd.n3940 gnd.n1425 19.3944
R9536 gnd.n3944 gnd.n1425 19.3944
R9537 gnd.n3946 gnd.n3944 19.3944
R9538 gnd.n3947 gnd.n3946 19.3944
R9539 gnd.n3947 gnd.n1423 19.3944
R9540 gnd.n3956 gnd.n1423 19.3944
R9541 gnd.n3956 gnd.n3955 19.3944
R9542 gnd.n3955 gnd.n3954 19.3944
R9543 gnd.n3954 gnd.n1388 19.3944
R9544 gnd.n3995 gnd.n1388 19.3944
R9545 gnd.n3995 gnd.n1386 19.3944
R9546 gnd.n4008 gnd.n1386 19.3944
R9547 gnd.n4008 gnd.n4007 19.3944
R9548 gnd.n4007 gnd.n4006 19.3944
R9549 gnd.n4006 gnd.n4005 19.3944
R9550 gnd.n4005 gnd.n4003 19.3944
R9551 gnd.n4003 gnd.n297 19.3944
R9552 gnd.n6682 gnd.n297 19.3944
R9553 gnd.n6682 gnd.n295 19.3944
R9554 gnd.n6686 gnd.n295 19.3944
R9555 gnd.n6747 gnd.n6686 19.3944
R9556 gnd.n6747 gnd.n6746 19.3944
R9557 gnd.n6746 gnd.n6745 19.3944
R9558 gnd.n6745 gnd.n6744 19.3944
R9559 gnd.n6744 gnd.n6742 19.3944
R9560 gnd.n6742 gnd.n6741 19.3944
R9561 gnd.n6741 gnd.n6739 19.3944
R9562 gnd.n6739 gnd.n6738 19.3944
R9563 gnd.n6738 gnd.n6736 19.3944
R9564 gnd.n6736 gnd.n6735 19.3944
R9565 gnd.n6735 gnd.n6733 19.3944
R9566 gnd.n6733 gnd.n6732 19.3944
R9567 gnd.n6732 gnd.n6730 19.3944
R9568 gnd.n6730 gnd.n6729 19.3944
R9569 gnd.n6729 gnd.n6727 19.3944
R9570 gnd.n6727 gnd.n6726 19.3944
R9571 gnd.n6726 gnd.n6724 19.3944
R9572 gnd.n6724 gnd.n6723 19.3944
R9573 gnd.n6723 gnd.n6721 19.3944
R9574 gnd.n6721 gnd.n6720 19.3944
R9575 gnd.n6720 gnd.n6716 19.3944
R9576 gnd.n6716 gnd.n6715 19.3944
R9577 gnd.n6715 gnd.n6713 19.3944
R9578 gnd.n6713 gnd.n6712 19.3944
R9579 gnd.n6712 gnd.n178 19.3944
R9580 gnd.n6937 gnd.n178 19.3944
R9581 gnd.n6938 gnd.n6937 19.3944
R9582 gnd.n6976 gnd.n139 19.3944
R9583 gnd.n6971 gnd.n139 19.3944
R9584 gnd.n6971 gnd.n6970 19.3944
R9585 gnd.n6970 gnd.n6969 19.3944
R9586 gnd.n6969 gnd.n146 19.3944
R9587 gnd.n6964 gnd.n146 19.3944
R9588 gnd.n6964 gnd.n6963 19.3944
R9589 gnd.n6963 gnd.n6962 19.3944
R9590 gnd.n6962 gnd.n153 19.3944
R9591 gnd.n6957 gnd.n153 19.3944
R9592 gnd.n6957 gnd.n6956 19.3944
R9593 gnd.n6956 gnd.n6955 19.3944
R9594 gnd.n6955 gnd.n160 19.3944
R9595 gnd.n6950 gnd.n160 19.3944
R9596 gnd.n6950 gnd.n6949 19.3944
R9597 gnd.n6949 gnd.n6948 19.3944
R9598 gnd.n6948 gnd.n167 19.3944
R9599 gnd.n6943 gnd.n167 19.3944
R9600 gnd.n7009 gnd.n7008 19.3944
R9601 gnd.n7008 gnd.n7007 19.3944
R9602 gnd.n7007 gnd.n111 19.3944
R9603 gnd.n7002 gnd.n111 19.3944
R9604 gnd.n7002 gnd.n7001 19.3944
R9605 gnd.n7001 gnd.n7000 19.3944
R9606 gnd.n7000 gnd.n118 19.3944
R9607 gnd.n6995 gnd.n118 19.3944
R9608 gnd.n6995 gnd.n6994 19.3944
R9609 gnd.n6994 gnd.n6993 19.3944
R9610 gnd.n6993 gnd.n125 19.3944
R9611 gnd.n6988 gnd.n125 19.3944
R9612 gnd.n6988 gnd.n6987 19.3944
R9613 gnd.n6987 gnd.n6986 19.3944
R9614 gnd.n6986 gnd.n132 19.3944
R9615 gnd.n6981 gnd.n132 19.3944
R9616 gnd.n6981 gnd.n6980 19.3944
R9617 gnd.n4057 gnd.n4056 19.3944
R9618 gnd.n4056 gnd.n4055 19.3944
R9619 gnd.n4055 gnd.n1334 19.3944
R9620 gnd.n3932 gnd.n1334 19.3944
R9621 gnd.n3932 gnd.n1433 19.3944
R9622 gnd.n3936 gnd.n1433 19.3944
R9623 gnd.n3936 gnd.n1405 19.3944
R9624 gnd.n3969 gnd.n1405 19.3944
R9625 gnd.n3969 gnd.n1403 19.3944
R9626 gnd.n3975 gnd.n1403 19.3944
R9627 gnd.n3975 gnd.n3974 19.3944
R9628 gnd.n3974 gnd.n1366 19.3944
R9629 gnd.n4022 gnd.n1366 19.3944
R9630 gnd.n4022 gnd.n1364 19.3944
R9631 gnd.n4026 gnd.n1364 19.3944
R9632 gnd.n4026 gnd.n321 19.3944
R9633 gnd.n6654 gnd.n321 19.3944
R9634 gnd.n6654 gnd.n319 19.3944
R9635 gnd.n6660 gnd.n319 19.3944
R9636 gnd.n6660 gnd.n6659 19.3944
R9637 gnd.n6659 gnd.n266 19.3944
R9638 gnd.n6774 gnd.n266 19.3944
R9639 gnd.n265 gnd.n264 19.3944
R9640 gnd.n303 gnd.n264 19.3944
R9641 gnd.n291 gnd.n290 19.3944
R9642 gnd.n6754 gnd.n6753 19.3944
R9643 gnd.n6777 gnd.n258 19.3944
R9644 gnd.n6777 gnd.n247 19.3944
R9645 gnd.n6789 gnd.n247 19.3944
R9646 gnd.n6789 gnd.n245 19.3944
R9647 gnd.n6793 gnd.n245 19.3944
R9648 gnd.n6793 gnd.n230 19.3944
R9649 gnd.n6805 gnd.n230 19.3944
R9650 gnd.n6805 gnd.n228 19.3944
R9651 gnd.n6809 gnd.n228 19.3944
R9652 gnd.n6809 gnd.n217 19.3944
R9653 gnd.n6821 gnd.n217 19.3944
R9654 gnd.n6821 gnd.n215 19.3944
R9655 gnd.n6825 gnd.n215 19.3944
R9656 gnd.n6825 gnd.n201 19.3944
R9657 gnd.n6837 gnd.n201 19.3944
R9658 gnd.n6837 gnd.n199 19.3944
R9659 gnd.n6841 gnd.n199 19.3944
R9660 gnd.n6841 gnd.n186 19.3944
R9661 gnd.n6928 gnd.n186 19.3944
R9662 gnd.n6928 gnd.n184 19.3944
R9663 gnd.n6932 gnd.n184 19.3944
R9664 gnd.n6932 gnd.n106 19.3944
R9665 gnd.n7012 gnd.n106 19.3944
R9666 gnd.n4441 gnd.n4440 19.3944
R9667 gnd.n4440 gnd.n4439 19.3944
R9668 gnd.n4439 gnd.n4438 19.3944
R9669 gnd.n4438 gnd.n4436 19.3944
R9670 gnd.n4436 gnd.n4433 19.3944
R9671 gnd.n4433 gnd.n4432 19.3944
R9672 gnd.n4432 gnd.n4429 19.3944
R9673 gnd.n4429 gnd.n4428 19.3944
R9674 gnd.n4428 gnd.n4425 19.3944
R9675 gnd.n4425 gnd.n4424 19.3944
R9676 gnd.n4424 gnd.n4421 19.3944
R9677 gnd.n4421 gnd.n4420 19.3944
R9678 gnd.n4420 gnd.n4417 19.3944
R9679 gnd.n4417 gnd.n4416 19.3944
R9680 gnd.n4416 gnd.n4413 19.3944
R9681 gnd.n4413 gnd.n4412 19.3944
R9682 gnd.n4412 gnd.n4409 19.3944
R9683 gnd.n4407 gnd.n4404 19.3944
R9684 gnd.n4404 gnd.n4403 19.3944
R9685 gnd.n4403 gnd.n4400 19.3944
R9686 gnd.n4400 gnd.n4399 19.3944
R9687 gnd.n4399 gnd.n4396 19.3944
R9688 gnd.n4396 gnd.n4395 19.3944
R9689 gnd.n4395 gnd.n4392 19.3944
R9690 gnd.n4392 gnd.n4391 19.3944
R9691 gnd.n4391 gnd.n4388 19.3944
R9692 gnd.n4388 gnd.n4387 19.3944
R9693 gnd.n4387 gnd.n4384 19.3944
R9694 gnd.n4384 gnd.n4383 19.3944
R9695 gnd.n4383 gnd.n4380 19.3944
R9696 gnd.n4380 gnd.n4379 19.3944
R9697 gnd.n4379 gnd.n4376 19.3944
R9698 gnd.n4376 gnd.n4375 19.3944
R9699 gnd.n4375 gnd.n4372 19.3944
R9700 gnd.n4372 gnd.n4371 19.3944
R9701 gnd.n4364 gnd.n4363 19.3944
R9702 gnd.n4363 gnd.n934 19.3944
R9703 gnd.n4359 gnd.n934 19.3944
R9704 gnd.n4359 gnd.n936 19.3944
R9705 gnd.n2203 gnd.n936 19.3944
R9706 gnd.n2205 gnd.n2203 19.3944
R9707 gnd.n2205 gnd.n2201 19.3944
R9708 gnd.n2210 gnd.n2201 19.3944
R9709 gnd.n2211 gnd.n2210 19.3944
R9710 gnd.n2213 gnd.n2211 19.3944
R9711 gnd.n2213 gnd.n2199 19.3944
R9712 gnd.n2218 gnd.n2199 19.3944
R9713 gnd.n2219 gnd.n2218 19.3944
R9714 gnd.n2221 gnd.n2219 19.3944
R9715 gnd.n2221 gnd.n2197 19.3944
R9716 gnd.n2226 gnd.n2197 19.3944
R9717 gnd.n2227 gnd.n2226 19.3944
R9718 gnd.n2229 gnd.n2227 19.3944
R9719 gnd.n2229 gnd.n2195 19.3944
R9720 gnd.n2234 gnd.n2195 19.3944
R9721 gnd.n2235 gnd.n2234 19.3944
R9722 gnd.n2237 gnd.n2235 19.3944
R9723 gnd.n2237 gnd.n2193 19.3944
R9724 gnd.n2242 gnd.n2193 19.3944
R9725 gnd.n2243 gnd.n2242 19.3944
R9726 gnd.n2245 gnd.n2243 19.3944
R9727 gnd.n2245 gnd.n2190 19.3944
R9728 gnd.n2255 gnd.n2190 19.3944
R9729 gnd.n2255 gnd.n2254 19.3944
R9730 gnd.n2254 gnd.n2253 19.3944
R9731 gnd.n2253 gnd.n2186 19.3944
R9732 gnd.n2419 gnd.n2186 19.3944
R9733 gnd.n2419 gnd.n2184 19.3944
R9734 gnd.n2424 gnd.n2184 19.3944
R9735 gnd.n2424 gnd.n2151 19.3944
R9736 gnd.n2436 gnd.n2151 19.3944
R9737 gnd.n2437 gnd.n2436 19.3944
R9738 gnd.n2438 gnd.n2437 19.3944
R9739 gnd.n2438 gnd.n2149 19.3944
R9740 gnd.n2444 gnd.n2149 19.3944
R9741 gnd.n2445 gnd.n2444 19.3944
R9742 gnd.n2449 gnd.n2445 19.3944
R9743 gnd.n2449 gnd.n2147 19.3944
R9744 gnd.n2457 gnd.n2147 19.3944
R9745 gnd.n2457 gnd.n2456 19.3944
R9746 gnd.n2456 gnd.n2455 19.3944
R9747 gnd.n2455 gnd.n2123 19.3944
R9748 gnd.n2529 gnd.n2123 19.3944
R9749 gnd.n2529 gnd.n2121 19.3944
R9750 gnd.n2534 gnd.n2121 19.3944
R9751 gnd.n2534 gnd.n2116 19.3944
R9752 gnd.n2582 gnd.n2116 19.3944
R9753 gnd.n2583 gnd.n2582 19.3944
R9754 gnd.n2625 gnd.n2090 19.3944
R9755 gnd.n2625 gnd.n2622 19.3944
R9756 gnd.n2622 gnd.n2619 19.3944
R9757 gnd.n2619 gnd.n2618 19.3944
R9758 gnd.n2618 gnd.n2615 19.3944
R9759 gnd.n2615 gnd.n2614 19.3944
R9760 gnd.n2614 gnd.n2611 19.3944
R9761 gnd.n2611 gnd.n2610 19.3944
R9762 gnd.n2610 gnd.n2607 19.3944
R9763 gnd.n2607 gnd.n2606 19.3944
R9764 gnd.n2606 gnd.n2603 19.3944
R9765 gnd.n2603 gnd.n2602 19.3944
R9766 gnd.n2602 gnd.n2599 19.3944
R9767 gnd.n2599 gnd.n2598 19.3944
R9768 gnd.n2598 gnd.n2595 19.3944
R9769 gnd.n2595 gnd.n2594 19.3944
R9770 gnd.n2594 gnd.n2591 19.3944
R9771 gnd.n2591 gnd.n2590 19.3944
R9772 gnd.n2073 gnd.n2072 19.3944
R9773 gnd.n2784 gnd.n2072 19.3944
R9774 gnd.n2784 gnd.n2783 19.3944
R9775 gnd.n2783 gnd.n2782 19.3944
R9776 gnd.n2782 gnd.n2779 19.3944
R9777 gnd.n2779 gnd.n2778 19.3944
R9778 gnd.n2778 gnd.n2775 19.3944
R9779 gnd.n2775 gnd.n2774 19.3944
R9780 gnd.n2774 gnd.n2771 19.3944
R9781 gnd.n2771 gnd.n2770 19.3944
R9782 gnd.n2770 gnd.n2767 19.3944
R9783 gnd.n2767 gnd.n2766 19.3944
R9784 gnd.n2766 gnd.n2763 19.3944
R9785 gnd.n2763 gnd.n2762 19.3944
R9786 gnd.n2762 gnd.n2759 19.3944
R9787 gnd.n2344 gnd.n2276 19.3944
R9788 gnd.n2344 gnd.n2277 19.3944
R9789 gnd.n2340 gnd.n2277 19.3944
R9790 gnd.n2340 gnd.n956 19.3944
R9791 gnd.n4349 gnd.n956 19.3944
R9792 gnd.n4349 gnd.n4348 19.3944
R9793 gnd.n4348 gnd.n4347 19.3944
R9794 gnd.n4347 gnd.n960 19.3944
R9795 gnd.n4337 gnd.n960 19.3944
R9796 gnd.n4337 gnd.n4336 19.3944
R9797 gnd.n4336 gnd.n4335 19.3944
R9798 gnd.n4335 gnd.n979 19.3944
R9799 gnd.n4325 gnd.n979 19.3944
R9800 gnd.n4325 gnd.n4324 19.3944
R9801 gnd.n4324 gnd.n4323 19.3944
R9802 gnd.n4323 gnd.n1000 19.3944
R9803 gnd.n4313 gnd.n1000 19.3944
R9804 gnd.n4313 gnd.n4312 19.3944
R9805 gnd.n4312 gnd.n4311 19.3944
R9806 gnd.n4311 gnd.n1019 19.3944
R9807 gnd.n4301 gnd.n1019 19.3944
R9808 gnd.n4301 gnd.n4300 19.3944
R9809 gnd.n4300 gnd.n4299 19.3944
R9810 gnd.n4299 gnd.n1040 19.3944
R9811 gnd.n4289 gnd.n1040 19.3944
R9812 gnd.n4289 gnd.n4288 19.3944
R9813 gnd.n4288 gnd.n4287 19.3944
R9814 gnd.n4287 gnd.n1057 19.3944
R9815 gnd.n4276 gnd.n1057 19.3944
R9816 gnd.n4276 gnd.n4275 19.3944
R9817 gnd.n4275 gnd.n4274 19.3944
R9818 gnd.n4274 gnd.n1075 19.3944
R9819 gnd.n4264 gnd.n1075 19.3944
R9820 gnd.n4264 gnd.n4263 19.3944
R9821 gnd.n4263 gnd.n4262 19.3944
R9822 gnd.n4262 gnd.n1094 19.3944
R9823 gnd.n4252 gnd.n1094 19.3944
R9824 gnd.n4252 gnd.n4251 19.3944
R9825 gnd.n4251 gnd.n4250 19.3944
R9826 gnd.n4250 gnd.n1116 19.3944
R9827 gnd.n4240 gnd.n1116 19.3944
R9828 gnd.n4240 gnd.n4239 19.3944
R9829 gnd.n4239 gnd.n4238 19.3944
R9830 gnd.n4238 gnd.n1136 19.3944
R9831 gnd.n4228 gnd.n1136 19.3944
R9832 gnd.n4228 gnd.n4227 19.3944
R9833 gnd.n4227 gnd.n4226 19.3944
R9834 gnd.n4226 gnd.n1158 19.3944
R9835 gnd.n4216 gnd.n1158 19.3944
R9836 gnd.n4216 gnd.n4215 19.3944
R9837 gnd.n4215 gnd.n4214 19.3944
R9838 gnd.n4214 gnd.n1179 19.3944
R9839 gnd.n4204 gnd.n1179 19.3944
R9840 gnd.n2336 gnd.n2334 19.3944
R9841 gnd.n2334 gnd.n2331 19.3944
R9842 gnd.n2331 gnd.n2330 19.3944
R9843 gnd.n2330 gnd.n2327 19.3944
R9844 gnd.n2327 gnd.n2326 19.3944
R9845 gnd.n2326 gnd.n2323 19.3944
R9846 gnd.n2323 gnd.n2322 19.3944
R9847 gnd.n2322 gnd.n2319 19.3944
R9848 gnd.n2319 gnd.n2318 19.3944
R9849 gnd.n2318 gnd.n2315 19.3944
R9850 gnd.n2315 gnd.n2314 19.3944
R9851 gnd.n2314 gnd.n2311 19.3944
R9852 gnd.n2311 gnd.n2310 19.3944
R9853 gnd.n2310 gnd.n2307 19.3944
R9854 gnd.n2307 gnd.n2306 19.3944
R9855 gnd.n2306 gnd.n2303 19.3944
R9856 gnd.n2297 gnd.n2272 19.3944
R9857 gnd.n2355 gnd.n2272 19.3944
R9858 gnd.n2355 gnd.n2270 19.3944
R9859 gnd.n2360 gnd.n2270 19.3944
R9860 gnd.n2361 gnd.n2360 19.3944
R9861 gnd.n2363 gnd.n2361 19.3944
R9862 gnd.n2363 gnd.n2268 19.3944
R9863 gnd.n2368 gnd.n2268 19.3944
R9864 gnd.n2369 gnd.n2368 19.3944
R9865 gnd.n2371 gnd.n2369 19.3944
R9866 gnd.n2371 gnd.n2266 19.3944
R9867 gnd.n2376 gnd.n2266 19.3944
R9868 gnd.n2377 gnd.n2376 19.3944
R9869 gnd.n2379 gnd.n2377 19.3944
R9870 gnd.n2379 gnd.n2264 19.3944
R9871 gnd.n2384 gnd.n2264 19.3944
R9872 gnd.n2385 gnd.n2384 19.3944
R9873 gnd.n2387 gnd.n2385 19.3944
R9874 gnd.n2387 gnd.n2262 19.3944
R9875 gnd.n2392 gnd.n2262 19.3944
R9876 gnd.n2393 gnd.n2392 19.3944
R9877 gnd.n2395 gnd.n2393 19.3944
R9878 gnd.n2395 gnd.n2260 19.3944
R9879 gnd.n2400 gnd.n2260 19.3944
R9880 gnd.n2401 gnd.n2400 19.3944
R9881 gnd.n2403 gnd.n2401 19.3944
R9882 gnd.n2403 gnd.n2189 19.3944
R9883 gnd.n2408 gnd.n2189 19.3944
R9884 gnd.n2409 gnd.n2408 19.3944
R9885 gnd.n2411 gnd.n2409 19.3944
R9886 gnd.n2411 gnd.n2187 19.3944
R9887 gnd.n2415 gnd.n2187 19.3944
R9888 gnd.n2415 gnd.n2155 19.3944
R9889 gnd.n2428 gnd.n2155 19.3944
R9890 gnd.n2428 gnd.n2153 19.3944
R9891 gnd.n2432 gnd.n2153 19.3944
R9892 gnd.n2432 gnd.n2140 19.3944
R9893 gnd.n2471 gnd.n2140 19.3944
R9894 gnd.n2471 gnd.n2141 19.3944
R9895 gnd.n2467 gnd.n2141 19.3944
R9896 gnd.n2467 gnd.n2466 19.3944
R9897 gnd.n2466 gnd.n2465 19.3944
R9898 gnd.n2465 gnd.n2146 19.3944
R9899 gnd.n2461 gnd.n2146 19.3944
R9900 gnd.n2461 gnd.n2126 19.3944
R9901 gnd.n2521 gnd.n2126 19.3944
R9902 gnd.n2521 gnd.n2124 19.3944
R9903 gnd.n2525 gnd.n2124 19.3944
R9904 gnd.n2525 gnd.n2120 19.3944
R9905 gnd.n2538 gnd.n2120 19.3944
R9906 gnd.n2538 gnd.n2117 19.3944
R9907 gnd.n2578 gnd.n2117 19.3944
R9908 gnd.n2578 gnd.n2118 19.3944
R9909 gnd.n2350 gnd.n2346 19.3944
R9910 gnd.n2350 gnd.n945 19.3944
R9911 gnd.n4355 gnd.n945 19.3944
R9912 gnd.n4355 gnd.n4354 19.3944
R9913 gnd.n4354 gnd.n4353 19.3944
R9914 gnd.n4353 gnd.n949 19.3944
R9915 gnd.n4343 gnd.n949 19.3944
R9916 gnd.n4343 gnd.n4342 19.3944
R9917 gnd.n4342 gnd.n4341 19.3944
R9918 gnd.n4341 gnd.n970 19.3944
R9919 gnd.n4331 gnd.n970 19.3944
R9920 gnd.n4331 gnd.n4330 19.3944
R9921 gnd.n4330 gnd.n4329 19.3944
R9922 gnd.n4329 gnd.n989 19.3944
R9923 gnd.n4319 gnd.n989 19.3944
R9924 gnd.n4319 gnd.n4318 19.3944
R9925 gnd.n4318 gnd.n4317 19.3944
R9926 gnd.n4317 gnd.n1010 19.3944
R9927 gnd.n4307 gnd.n1010 19.3944
R9928 gnd.n4307 gnd.n4306 19.3944
R9929 gnd.n4306 gnd.n4305 19.3944
R9930 gnd.n4305 gnd.n1029 19.3944
R9931 gnd.n4295 gnd.n4294 19.3944
R9932 gnd.n4294 gnd.n4293 19.3944
R9933 gnd.n4283 gnd.n1063 19.3944
R9934 gnd.n4281 gnd.n4280 19.3944
R9935 gnd.n4270 gnd.n1081 19.3944
R9936 gnd.n4270 gnd.n4269 19.3944
R9937 gnd.n4269 gnd.n4268 19.3944
R9938 gnd.n4268 gnd.n1084 19.3944
R9939 gnd.n4258 gnd.n1084 19.3944
R9940 gnd.n4258 gnd.n4257 19.3944
R9941 gnd.n4257 gnd.n4256 19.3944
R9942 gnd.n4256 gnd.n1105 19.3944
R9943 gnd.n4246 gnd.n1105 19.3944
R9944 gnd.n4246 gnd.n4245 19.3944
R9945 gnd.n4245 gnd.n4244 19.3944
R9946 gnd.n4244 gnd.n1126 19.3944
R9947 gnd.n4234 gnd.n1126 19.3944
R9948 gnd.n4234 gnd.n4233 19.3944
R9949 gnd.n4233 gnd.n4232 19.3944
R9950 gnd.n4232 gnd.n1147 19.3944
R9951 gnd.n4222 gnd.n1147 19.3944
R9952 gnd.n4222 gnd.n4221 19.3944
R9953 gnd.n4221 gnd.n4220 19.3944
R9954 gnd.n4220 gnd.n1168 19.3944
R9955 gnd.n4210 gnd.n1168 19.3944
R9956 gnd.n4210 gnd.n4209 19.3944
R9957 gnd.n4209 gnd.n4208 19.3944
R9958 gnd.n6060 gnd.n679 19.3944
R9959 gnd.n6060 gnd.n6059 19.3944
R9960 gnd.n6059 gnd.n6058 19.3944
R9961 gnd.n6058 gnd.n683 19.3944
R9962 gnd.n6052 gnd.n683 19.3944
R9963 gnd.n6052 gnd.n6051 19.3944
R9964 gnd.n6051 gnd.n6050 19.3944
R9965 gnd.n6050 gnd.n691 19.3944
R9966 gnd.n6044 gnd.n691 19.3944
R9967 gnd.n6044 gnd.n6043 19.3944
R9968 gnd.n6043 gnd.n6042 19.3944
R9969 gnd.n6042 gnd.n699 19.3944
R9970 gnd.n6036 gnd.n699 19.3944
R9971 gnd.n6036 gnd.n6035 19.3944
R9972 gnd.n6035 gnd.n6034 19.3944
R9973 gnd.n6034 gnd.n707 19.3944
R9974 gnd.n6028 gnd.n707 19.3944
R9975 gnd.n6028 gnd.n6027 19.3944
R9976 gnd.n6027 gnd.n6026 19.3944
R9977 gnd.n6026 gnd.n715 19.3944
R9978 gnd.n6020 gnd.n715 19.3944
R9979 gnd.n6020 gnd.n6019 19.3944
R9980 gnd.n6019 gnd.n6018 19.3944
R9981 gnd.n6018 gnd.n723 19.3944
R9982 gnd.n6012 gnd.n723 19.3944
R9983 gnd.n6012 gnd.n6011 19.3944
R9984 gnd.n6011 gnd.n6010 19.3944
R9985 gnd.n6010 gnd.n731 19.3944
R9986 gnd.n6004 gnd.n731 19.3944
R9987 gnd.n6004 gnd.n6003 19.3944
R9988 gnd.n6003 gnd.n6002 19.3944
R9989 gnd.n6002 gnd.n739 19.3944
R9990 gnd.n5996 gnd.n739 19.3944
R9991 gnd.n5996 gnd.n5995 19.3944
R9992 gnd.n5995 gnd.n5994 19.3944
R9993 gnd.n5994 gnd.n747 19.3944
R9994 gnd.n5988 gnd.n747 19.3944
R9995 gnd.n5988 gnd.n5987 19.3944
R9996 gnd.n5987 gnd.n5986 19.3944
R9997 gnd.n5986 gnd.n755 19.3944
R9998 gnd.n5980 gnd.n755 19.3944
R9999 gnd.n5980 gnd.n5979 19.3944
R10000 gnd.n5979 gnd.n5978 19.3944
R10001 gnd.n5978 gnd.n763 19.3944
R10002 gnd.n5972 gnd.n763 19.3944
R10003 gnd.n5972 gnd.n5971 19.3944
R10004 gnd.n5971 gnd.n5970 19.3944
R10005 gnd.n5970 gnd.n771 19.3944
R10006 gnd.n5964 gnd.n771 19.3944
R10007 gnd.n5964 gnd.n5963 19.3944
R10008 gnd.n5963 gnd.n5962 19.3944
R10009 gnd.n5962 gnd.n779 19.3944
R10010 gnd.n5956 gnd.n779 19.3944
R10011 gnd.n5956 gnd.n5955 19.3944
R10012 gnd.n5955 gnd.n5954 19.3944
R10013 gnd.n5954 gnd.n787 19.3944
R10014 gnd.n5948 gnd.n787 19.3944
R10015 gnd.n5948 gnd.n5947 19.3944
R10016 gnd.n5947 gnd.n5946 19.3944
R10017 gnd.n5946 gnd.n795 19.3944
R10018 gnd.n5940 gnd.n795 19.3944
R10019 gnd.n5940 gnd.n5939 19.3944
R10020 gnd.n5939 gnd.n5938 19.3944
R10021 gnd.n5938 gnd.n803 19.3944
R10022 gnd.n5932 gnd.n803 19.3944
R10023 gnd.n5932 gnd.n5931 19.3944
R10024 gnd.n5931 gnd.n5930 19.3944
R10025 gnd.n5930 gnd.n811 19.3944
R10026 gnd.n5924 gnd.n811 19.3944
R10027 gnd.n5924 gnd.n5923 19.3944
R10028 gnd.n5923 gnd.n5922 19.3944
R10029 gnd.n5922 gnd.n819 19.3944
R10030 gnd.n5916 gnd.n819 19.3944
R10031 gnd.n5916 gnd.n5915 19.3944
R10032 gnd.n5915 gnd.n5914 19.3944
R10033 gnd.n5914 gnd.n827 19.3944
R10034 gnd.n5908 gnd.n827 19.3944
R10035 gnd.n5908 gnd.n5907 19.3944
R10036 gnd.n5907 gnd.n5906 19.3944
R10037 gnd.n5906 gnd.n835 19.3944
R10038 gnd.n5900 gnd.n835 19.3944
R10039 gnd.n5900 gnd.n5899 19.3944
R10040 gnd.n5899 gnd.n5898 19.3944
R10041 gnd.n5898 gnd.n843 19.3944
R10042 gnd.n4199 gnd.n4198 19.3944
R10043 gnd.n4198 gnd.n4197 19.3944
R10044 gnd.n4197 gnd.n1203 19.3944
R10045 gnd.n4193 gnd.n1203 19.3944
R10046 gnd.n4193 gnd.n4192 19.3944
R10047 gnd.n4192 gnd.n4191 19.3944
R10048 gnd.n4191 gnd.n1208 19.3944
R10049 gnd.n4187 gnd.n1208 19.3944
R10050 gnd.n4187 gnd.n4186 19.3944
R10051 gnd.n4186 gnd.n4185 19.3944
R10052 gnd.n4185 gnd.n1213 19.3944
R10053 gnd.n4181 gnd.n1213 19.3944
R10054 gnd.n4181 gnd.n4180 19.3944
R10055 gnd.n4180 gnd.n4179 19.3944
R10056 gnd.n4179 gnd.n1218 19.3944
R10057 gnd.n4175 gnd.n1218 19.3944
R10058 gnd.n4175 gnd.n4174 19.3944
R10059 gnd.n4174 gnd.n4173 19.3944
R10060 gnd.n4173 gnd.n1223 19.3944
R10061 gnd.n4169 gnd.n1223 19.3944
R10062 gnd.n4169 gnd.n4168 19.3944
R10063 gnd.n4168 gnd.n4167 19.3944
R10064 gnd.n4167 gnd.n1228 19.3944
R10065 gnd.n4163 gnd.n1228 19.3944
R10066 gnd.n4163 gnd.n4162 19.3944
R10067 gnd.n4162 gnd.n4161 19.3944
R10068 gnd.n4161 gnd.n1233 19.3944
R10069 gnd.n4157 gnd.n1233 19.3944
R10070 gnd.n4157 gnd.n4156 19.3944
R10071 gnd.n4156 gnd.n4155 19.3944
R10072 gnd.n4155 gnd.n1238 19.3944
R10073 gnd.n4151 gnd.n1238 19.3944
R10074 gnd.n4151 gnd.n4150 19.3944
R10075 gnd.n4150 gnd.n4149 19.3944
R10076 gnd.n4149 gnd.n1243 19.3944
R10077 gnd.n4145 gnd.n1243 19.3944
R10078 gnd.n4145 gnd.n4144 19.3944
R10079 gnd.n4144 gnd.n4143 19.3944
R10080 gnd.n4143 gnd.n1248 19.3944
R10081 gnd.n4139 gnd.n1248 19.3944
R10082 gnd.n4139 gnd.n4138 19.3944
R10083 gnd.n4138 gnd.n4137 19.3944
R10084 gnd.n4137 gnd.n1253 19.3944
R10085 gnd.n4133 gnd.n1253 19.3944
R10086 gnd.n4133 gnd.n4132 19.3944
R10087 gnd.n4132 gnd.n4131 19.3944
R10088 gnd.n4131 gnd.n1258 19.3944
R10089 gnd.n4127 gnd.n1258 19.3944
R10090 gnd.n4127 gnd.n4126 19.3944
R10091 gnd.n4126 gnd.n4125 19.3944
R10092 gnd.n4125 gnd.n1263 19.3944
R10093 gnd.n4121 gnd.n1263 19.3944
R10094 gnd.n4121 gnd.n4120 19.3944
R10095 gnd.n4120 gnd.n4119 19.3944
R10096 gnd.n4119 gnd.n1268 19.3944
R10097 gnd.n4115 gnd.n1268 19.3944
R10098 gnd.n4115 gnd.n4114 19.3944
R10099 gnd.n4114 gnd.n4113 19.3944
R10100 gnd.n4113 gnd.n1273 19.3944
R10101 gnd.n4109 gnd.n1273 19.3944
R10102 gnd.n4109 gnd.n4108 19.3944
R10103 gnd.n4108 gnd.n4107 19.3944
R10104 gnd.n4107 gnd.n1278 19.3944
R10105 gnd.n4103 gnd.n1278 19.3944
R10106 gnd.n4103 gnd.n4102 19.3944
R10107 gnd.n4102 gnd.n4101 19.3944
R10108 gnd.n4101 gnd.n1283 19.3944
R10109 gnd.n4097 gnd.n1283 19.3944
R10110 gnd.n4097 gnd.n4096 19.3944
R10111 gnd.n4096 gnd.n4095 19.3944
R10112 gnd.n4095 gnd.n1288 19.3944
R10113 gnd.n4091 gnd.n1288 19.3944
R10114 gnd.n4091 gnd.n4090 19.3944
R10115 gnd.n4090 gnd.n4089 19.3944
R10116 gnd.n4089 gnd.n1293 19.3944
R10117 gnd.n4085 gnd.n1293 19.3944
R10118 gnd.n4085 gnd.n4084 19.3944
R10119 gnd.n4084 gnd.n4083 19.3944
R10120 gnd.n4083 gnd.n1298 19.3944
R10121 gnd.n4079 gnd.n1298 19.3944
R10122 gnd.n4079 gnd.n4078 19.3944
R10123 gnd.n4078 gnd.n4077 19.3944
R10124 gnd.n3560 gnd.n3395 19.3944
R10125 gnd.n3560 gnd.n3393 19.3944
R10126 gnd.n3565 gnd.n3393 19.3944
R10127 gnd.n3459 gnd.n3441 19.3944
R10128 gnd.n3459 gnd.n3439 19.3944
R10129 gnd.n3465 gnd.n3439 19.3944
R10130 gnd.n3465 gnd.n3432 19.3944
R10131 gnd.n3478 gnd.n3432 19.3944
R10132 gnd.n3478 gnd.n3430 19.3944
R10133 gnd.n3484 gnd.n3430 19.3944
R10134 gnd.n3484 gnd.n3423 19.3944
R10135 gnd.n3497 gnd.n3423 19.3944
R10136 gnd.n3497 gnd.n3421 19.3944
R10137 gnd.n3503 gnd.n3421 19.3944
R10138 gnd.n3503 gnd.n3414 19.3944
R10139 gnd.n3516 gnd.n3414 19.3944
R10140 gnd.n3516 gnd.n3412 19.3944
R10141 gnd.n3524 gnd.n3412 19.3944
R10142 gnd.n3524 gnd.n3523 19.3944
R10143 gnd.n3523 gnd.n3403 19.3944
R10144 gnd.n3537 gnd.n3403 19.3944
R10145 gnd.n3537 gnd.n3401 19.3944
R10146 gnd.n3543 gnd.n3401 19.3944
R10147 gnd.n3543 gnd.n3399 19.3944
R10148 gnd.n3547 gnd.n3399 19.3944
R10149 gnd.n3547 gnd.n3397 19.3944
R10150 gnd.n3556 gnd.n3397 19.3944
R10151 gnd.t289 gnd.n4968 18.8012
R10152 gnd.n5590 gnd.t313 18.8012
R10153 gnd.n5434 gnd.n5063 18.4825
R10154 gnd.n3840 gnd.n1487 18.4247
R10155 gnd.n2759 gnd.n2758 18.4247
R10156 gnd.n6891 gnd.n6890 18.2308
R10157 gnd.n3527 gnd.n3407 18.2308
R10158 gnd.n2797 gnd.n2026 18.2308
R10159 gnd.n2303 gnd.n2296 18.2308
R10160 gnd.n5506 gnd.t290 18.1639
R10161 gnd.n5487 gnd.t303 17.5266
R10162 gnd.t210 gnd.n953 17.5266
R10163 gnd.n4224 gnd.t159 17.5266
R10164 gnd.n3938 gnd.t231 17.5266
R10165 gnd.n6843 gnd.t238 17.5266
R10166 gnd.n4996 gnd.t298 16.8893
R10167 gnd.t198 gnd.n994 16.8893
R10168 gnd.n4248 gnd.t157 16.8893
R10169 gnd.n1371 gnd.t165 16.8893
R10170 gnd.n6811 gnd.t207 16.8893
R10171 gnd.t77 gnd.n5090 16.2519
R10172 gnd.n4953 gnd.t297 16.2519
R10173 gnd.t185 gnd.n1034 16.2519
R10174 gnd.n4278 gnd.n1066 16.2519
R10175 gnd.n4272 gnd.t173 16.2519
R10176 gnd.n6772 gnd.t183 16.2519
R10177 gnd.n6680 gnd.n302 16.2519
R10178 gnd.n6779 gnd.t180 16.2519
R10179 gnd.n2630 gnd.n2629 16.0975
R10180 gnd.n1526 gnd.n1525 16.0975
R10181 gnd.n2694 gnd.n2693 16.0975
R10182 gnd.n3646 gnd.n3645 16.0975
R10183 gnd.n2838 gnd.n2837 15.9333
R10184 gnd.n2837 gnd.n1960 15.9333
R10185 gnd.n2848 gnd.n2846 15.9333
R10186 gnd.n2848 gnd.n2847 15.9333
R10187 gnd.n2847 gnd.n1955 15.9333
R10188 gnd.n2858 gnd.n1955 15.9333
R10189 gnd.n2857 gnd.n2856 15.9333
R10190 gnd.n2856 gnd.n1949 15.9333
R10191 gnd.n2866 gnd.n1949 15.9333
R10192 gnd.n2868 gnd.n2866 15.9333
R10193 gnd.n2868 gnd.n2867 15.9333
R10194 gnd.n2867 gnd.n1942 15.9333
R10195 gnd.n2878 gnd.n1942 15.9333
R10196 gnd.n2878 gnd.n2877 15.9333
R10197 gnd.n2876 gnd.n1936 15.9333
R10198 gnd.n2886 gnd.n1936 15.9333
R10199 gnd.n2888 gnd.n2886 15.9333
R10200 gnd.n2888 gnd.n2887 15.9333
R10201 gnd.n2887 gnd.n1929 15.9333
R10202 gnd.n2898 gnd.n1929 15.9333
R10203 gnd.n2898 gnd.n2897 15.9333
R10204 gnd.n2897 gnd.n2896 15.9333
R10205 gnd.n2906 gnd.n1923 15.9333
R10206 gnd.n2908 gnd.n2906 15.9333
R10207 gnd.n2908 gnd.n2907 15.9333
R10208 gnd.n2907 gnd.n1916 15.9333
R10209 gnd.n2918 gnd.n1916 15.9333
R10210 gnd.n2918 gnd.n2917 15.9333
R10211 gnd.n2917 gnd.n2916 15.9333
R10212 gnd.n2916 gnd.n1910 15.9333
R10213 gnd.n2926 gnd.n1910 15.9333
R10214 gnd.n2928 gnd.n2927 15.9333
R10215 gnd.n2927 gnd.n1901 15.9333
R10216 gnd.n2956 gnd.n1901 15.9333
R10217 gnd.n2956 gnd.n2955 15.9333
R10218 gnd.n2955 gnd.n2954 15.9333
R10219 gnd.n2954 gnd.n1862 15.9333
R10220 gnd.n2964 gnd.n1895 15.9333
R10221 gnd.n1830 gnd.n1828 15.9333
R10222 gnd.n2940 gnd.n1810 15.9333
R10223 gnd.n3011 gnd.n1806 15.9333
R10224 gnd.n3044 gnd.n3043 15.9333
R10225 gnd.n3052 gnd.n1783 15.9333
R10226 gnd.n3111 gnd.n3110 15.9333
R10227 gnd.n3122 gnd.n3121 15.9333
R10228 gnd.n3099 gnd.n1746 15.9333
R10229 gnd.n3175 gnd.n3174 15.9333
R10230 gnd.n3174 gnd.n1710 15.9333
R10231 gnd.n3068 gnd.n1682 15.9333
R10232 gnd.n3222 gnd.n1676 15.9333
R10233 gnd.n3251 gnd.n1664 15.9333
R10234 gnd.n3264 gnd.n1660 15.9333
R10235 gnd.n3299 gnd.n3298 15.9333
R10236 gnd.n3351 gnd.n1492 15.9333
R10237 gnd.n3614 gnd.n1546 15.9333
R10238 gnd.n3614 gnd.n3613 15.9333
R10239 gnd.n3613 gnd.n3612 15.9333
R10240 gnd.n3612 gnd.n3611 15.9333
R10241 gnd.n3611 gnd.n3610 15.9333
R10242 gnd.n3610 gnd.n1549 15.9333
R10243 gnd.n1561 gnd.n1559 15.9333
R10244 gnd.n3604 gnd.n1561 15.9333
R10245 gnd.n3604 gnd.n3603 15.9333
R10246 gnd.n3603 gnd.n3602 15.9333
R10247 gnd.n3602 gnd.n3601 15.9333
R10248 gnd.n3601 gnd.n3600 15.9333
R10249 gnd.n3600 gnd.n1564 15.9333
R10250 gnd.n3369 gnd.n1564 15.9333
R10251 gnd.n3371 gnd.n3369 15.9333
R10252 gnd.n3594 gnd.n3593 15.9333
R10253 gnd.n3593 gnd.n3592 15.9333
R10254 gnd.n3592 gnd.n3591 15.9333
R10255 gnd.n3591 gnd.n3590 15.9333
R10256 gnd.n3590 gnd.n1574 15.9333
R10257 gnd.n1582 gnd.n1574 15.9333
R10258 gnd.n1584 gnd.n1582 15.9333
R10259 gnd.n3584 gnd.n1584 15.9333
R10260 gnd.n3583 gnd.n3582 15.9333
R10261 gnd.n3582 gnd.n3581 15.9333
R10262 gnd.n3581 gnd.n3580 15.9333
R10263 gnd.n3580 gnd.n1587 15.9333
R10264 gnd.n1597 gnd.n1587 15.9333
R10265 gnd.n1599 gnd.n1597 15.9333
R10266 gnd.n3574 gnd.n1599 15.9333
R10267 gnd.n3574 gnd.n3573 15.9333
R10268 gnd.n3572 gnd.n3571 15.9333
R10269 gnd.n3571 gnd.n1304 15.9333
R10270 gnd.n4075 gnd.n1304 15.9333
R10271 gnd.n4075 gnd.n4074 15.9333
R10272 gnd.n1315 gnd.n1306 15.9333
R10273 gnd.n4068 gnd.n1315 15.9333
R10274 gnd.n4770 gnd.n4768 15.6674
R10275 gnd.n4738 gnd.n4736 15.6674
R10276 gnd.n4706 gnd.n4704 15.6674
R10277 gnd.n4675 gnd.n4673 15.6674
R10278 gnd.n4643 gnd.n4641 15.6674
R10279 gnd.n4611 gnd.n4609 15.6674
R10280 gnd.n4579 gnd.n4577 15.6674
R10281 gnd.n4548 gnd.n4546 15.6674
R10282 gnd.n5208 gnd.t77 15.6146
R10283 gnd.n5798 gnd.t110 15.6146
R10284 gnd.n4297 gnd.t185 15.6146
R10285 gnd.n2257 gnd.n1066 15.6146
R10286 gnd.t114 gnd.n2857 15.6146
R10287 gnd.n3573 gnd.t85 15.6146
R10288 gnd.n6677 gnd.n302 15.6146
R10289 gnd.n288 gnd.t180 15.6146
R10290 gnd.n1775 gnd.n1769 15.296
R10291 gnd.n3130 gnd.n1755 15.296
R10292 gnd.n3239 gnd.n3238 15.296
R10293 gnd.n3274 gnd.n3273 15.296
R10294 gnd.t118 gnd.n1534 15.296
R10295 gnd.n3630 gnd.n3629 15.0827
R10296 gnd.n1847 gnd.n1842 15.0481
R10297 gnd.n3640 gnd.n3639 15.0481
R10298 gnd.n5695 gnd.t292 14.9773
R10299 gnd.n4321 gnd.t198 14.9773
R10300 gnd.n2896 gnd.t311 14.9773
R10301 gnd.n3594 gnd.t4 14.9773
R10302 gnd.n235 gnd.t207 14.9773
R10303 gnd.n2983 gnd.t121 14.6587
R10304 gnd.n3010 gnd.n1795 14.6587
R10305 gnd.n3310 gnd.n3309 14.6587
R10306 gnd.n3622 gnd.n3621 14.6587
R10307 gnd.n5727 gnd.t15 14.34
R10308 gnd.n5760 gnd.t302 14.34
R10309 gnd.n4345 gnd.t210 14.34
R10310 gnd.n6718 gnd.t238 14.34
R10311 gnd.t155 gnd.n5002 13.7027
R10312 gnd.n5403 gnd.n5399 13.5763
R10313 gnd.n5854 gnd.n4476 13.5763
R10314 gnd.n1467 gnd.n1466 13.5763
R10315 gnd.n6943 gnd.n6942 13.5763
R10316 gnd.n4371 gnd.n931 13.5763
R10317 gnd.n2590 gnd.n2587 13.5763
R10318 gnd.n5435 gnd.n5434 13.384
R10319 gnd.n3042 gnd.n1791 13.384
R10320 gnd.n3147 gnd.n3146 13.384
R10321 gnd.t13 gnd.n1742 13.384
R10322 gnd.t24 gnd.n3164 13.384
R10323 gnd.n3185 gnd.t287 13.384
R10324 gnd.t17 gnd.n3205 13.384
R10325 gnd.n3214 gnd.n1691 13.384
R10326 gnd.n3289 gnd.n1644 13.384
R10327 gnd.n1858 gnd.n1839 13.1884
R10328 gnd.n1853 gnd.n1852 13.1884
R10329 gnd.n1852 gnd.n1851 13.1884
R10330 gnd.n3633 gnd.n3628 13.1884
R10331 gnd.n3634 gnd.n3633 13.1884
R10332 gnd.n1854 gnd.n1841 13.146
R10333 gnd.n1850 gnd.n1841 13.146
R10334 gnd.n3632 gnd.n3631 13.146
R10335 gnd.n3632 gnd.n3627 13.146
R10336 gnd.n2928 gnd.t307 13.0654
R10337 gnd.t152 gnd.n1549 13.0654
R10338 gnd.n4771 gnd.n4767 12.8005
R10339 gnd.n4739 gnd.n4735 12.8005
R10340 gnd.n4707 gnd.n4703 12.8005
R10341 gnd.n4676 gnd.n4672 12.8005
R10342 gnd.n4644 gnd.n4640 12.8005
R10343 gnd.n4612 gnd.n4608 12.8005
R10344 gnd.n4580 gnd.n4576 12.8005
R10345 gnd.n4549 gnd.n4545 12.8005
R10346 gnd.n2975 gnd.n1836 12.7467
R10347 gnd.n3035 gnd.n3033 12.7467
R10348 gnd.n3091 gnd.n1733 12.7467
R10349 gnd.n3207 gnd.n1697 12.7467
R10350 gnd.n3297 gnd.n1647 12.7467
R10351 gnd.n5406 gnd.n5403 12.4126
R10352 gnd.n5859 gnd.n4476 12.4126
R10353 gnd.n3892 gnd.n1466 12.4126
R10354 gnd.n6942 gnd.n174 12.4126
R10355 gnd.n4367 gnd.n931 12.4126
R10356 gnd.n2587 gnd.n2112 12.4126
R10357 gnd.n2970 gnd.n2969 12.1761
R10358 gnd.n3709 gnd.n3708 12.1761
R10359 gnd.n2940 gnd.t42 12.1094
R10360 gnd.n1782 gnd.n1781 12.1094
R10361 gnd.n3100 gnd.n1757 12.1094
R10362 gnd.n3231 gnd.n3230 12.1094
R10363 gnd.n3281 gnd.n3280 12.1094
R10364 gnd.n3331 gnd.t48 12.1094
R10365 gnd.n4775 gnd.n4774 12.0247
R10366 gnd.n4743 gnd.n4742 12.0247
R10367 gnd.n4711 gnd.n4710 12.0247
R10368 gnd.n4680 gnd.n4679 12.0247
R10369 gnd.n4648 gnd.n4647 12.0247
R10370 gnd.n4616 gnd.n4615 12.0247
R10371 gnd.n4584 gnd.n4583 12.0247
R10372 gnd.n4553 gnd.n4552 12.0247
R10373 gnd.n2787 gnd.n2051 11.4721
R10374 gnd.n1831 gnd.n1818 11.4721
R10375 gnd.n3163 gnd.n1728 11.4721
R10376 gnd.n3187 gnd.n3186 11.4721
R10377 gnd.n3324 gnd.n3323 11.4721
R10378 gnd.n3321 gnd.t39 11.4721
R10379 gnd.n3342 gnd.n3340 11.4721
R10380 gnd.n4066 gnd.n1316 11.4721
R10381 gnd.n4778 gnd.n4765 11.249
R10382 gnd.n4746 gnd.n4733 11.249
R10383 gnd.n4714 gnd.n4701 11.249
R10384 gnd.n4683 gnd.n4670 11.249
R10385 gnd.n4651 gnd.n4638 11.249
R10386 gnd.n4619 gnd.n4606 11.249
R10387 gnd.n4587 gnd.n4574 11.249
R10388 gnd.n4556 gnd.n4543 11.249
R10389 gnd.n5507 gnd.t155 11.1535
R10390 gnd.n2877 gnd.t145 11.1535
R10391 gnd.t10 gnd.n3583 11.1535
R10392 gnd.n3123 gnd.n1761 10.8348
R10393 gnd.n3224 gnd.n3223 10.8348
R10394 gnd.n3774 gnd.n1488 10.6151
R10395 gnd.n3774 gnd.n3773 10.6151
R10396 gnd.n3771 gnd.n3768 10.6151
R10397 gnd.n3768 gnd.n3767 10.6151
R10398 gnd.n3767 gnd.n3764 10.6151
R10399 gnd.n3764 gnd.n3763 10.6151
R10400 gnd.n3763 gnd.n3760 10.6151
R10401 gnd.n3760 gnd.n3759 10.6151
R10402 gnd.n3759 gnd.n3756 10.6151
R10403 gnd.n3756 gnd.n3755 10.6151
R10404 gnd.n3755 gnd.n3752 10.6151
R10405 gnd.n3752 gnd.n3751 10.6151
R10406 gnd.n3751 gnd.n3748 10.6151
R10407 gnd.n3748 gnd.n3747 10.6151
R10408 gnd.n3747 gnd.n3744 10.6151
R10409 gnd.n3744 gnd.n3743 10.6151
R10410 gnd.n3743 gnd.n3740 10.6151
R10411 gnd.n3740 gnd.n3739 10.6151
R10412 gnd.n3739 gnd.n3736 10.6151
R10413 gnd.n3736 gnd.n3735 10.6151
R10414 gnd.n3735 gnd.n3732 10.6151
R10415 gnd.n3732 gnd.n3731 10.6151
R10416 gnd.n3731 gnd.n3728 10.6151
R10417 gnd.n3728 gnd.n3727 10.6151
R10418 gnd.n3727 gnd.n3724 10.6151
R10419 gnd.n3724 gnd.n3723 10.6151
R10420 gnd.n3723 gnd.n3720 10.6151
R10421 gnd.n3720 gnd.n3719 10.6151
R10422 gnd.n3719 gnd.n3716 10.6151
R10423 gnd.n3716 gnd.n3715 10.6151
R10424 gnd.n2978 gnd.n2977 10.6151
R10425 gnd.n2981 gnd.n2978 10.6151
R10426 gnd.n2981 gnd.n2980 10.6151
R10427 gnd.n2980 gnd.n2979 10.6151
R10428 gnd.n2979 gnd.n1808 10.6151
R10429 gnd.n3006 gnd.n1808 10.6151
R10430 gnd.n3007 gnd.n3006 10.6151
R10431 gnd.n3008 gnd.n3007 10.6151
R10432 gnd.n3008 gnd.n1798 10.6151
R10433 gnd.n3031 gnd.n1798 10.6151
R10434 gnd.n3031 gnd.n3030 10.6151
R10435 gnd.n3030 gnd.n3029 10.6151
R10436 gnd.n3029 gnd.n1799 10.6151
R10437 gnd.n1799 gnd.n1772 10.6151
R10438 gnd.n3062 gnd.n1772 10.6151
R10439 gnd.n3063 gnd.n3062 10.6151
R10440 gnd.n3107 gnd.n3063 10.6151
R10441 gnd.n3107 gnd.n3106 10.6151
R10442 gnd.n3106 gnd.n3105 10.6151
R10443 gnd.n3105 gnd.n3103 10.6151
R10444 gnd.n3103 gnd.n3102 10.6151
R10445 gnd.n3102 gnd.n3097 10.6151
R10446 gnd.n3097 gnd.n3096 10.6151
R10447 gnd.n3096 gnd.n3094 10.6151
R10448 gnd.n3094 gnd.n3093 10.6151
R10449 gnd.n3093 gnd.n3089 10.6151
R10450 gnd.n3089 gnd.n3088 10.6151
R10451 gnd.n3088 gnd.n3086 10.6151
R10452 gnd.n3086 gnd.n3085 10.6151
R10453 gnd.n3085 gnd.n3083 10.6151
R10454 gnd.n3083 gnd.n3082 10.6151
R10455 gnd.n3082 gnd.n3081 10.6151
R10456 gnd.n3081 gnd.n3080 10.6151
R10457 gnd.n3080 gnd.n3079 10.6151
R10458 gnd.n3079 gnd.n3075 10.6151
R10459 gnd.n3075 gnd.n3074 10.6151
R10460 gnd.n3074 gnd.n3072 10.6151
R10461 gnd.n3072 gnd.n3071 10.6151
R10462 gnd.n3071 gnd.n3067 10.6151
R10463 gnd.n3067 gnd.n3066 10.6151
R10464 gnd.n3066 gnd.n3064 10.6151
R10465 gnd.n3064 gnd.n1667 10.6151
R10466 gnd.n3254 gnd.n1667 10.6151
R10467 gnd.n3255 gnd.n3254 10.6151
R10468 gnd.n3269 gnd.n3255 10.6151
R10469 gnd.n3269 gnd.n3268 10.6151
R10470 gnd.n3268 gnd.n3267 10.6151
R10471 gnd.n3267 gnd.n3263 10.6151
R10472 gnd.n3263 gnd.n3262 10.6151
R10473 gnd.n3262 gnd.n3260 10.6151
R10474 gnd.n3260 gnd.n3259 10.6151
R10475 gnd.n3259 gnd.n3257 10.6151
R10476 gnd.n3257 gnd.n3256 10.6151
R10477 gnd.n3256 gnd.n1620 10.6151
R10478 gnd.n3333 gnd.n1620 10.6151
R10479 gnd.n3334 gnd.n3333 10.6151
R10480 gnd.n3337 gnd.n3334 10.6151
R10481 gnd.n3337 gnd.n3336 10.6151
R10482 gnd.n3336 gnd.n3335 10.6151
R10483 gnd.n3335 gnd.n1527 10.6151
R10484 gnd.n2692 gnd.n2691 10.6151
R10485 gnd.n2691 gnd.n2688 10.6151
R10486 gnd.n2686 gnd.n2683 10.6151
R10487 gnd.n2683 gnd.n2682 10.6151
R10488 gnd.n2682 gnd.n2679 10.6151
R10489 gnd.n2679 gnd.n2678 10.6151
R10490 gnd.n2678 gnd.n2675 10.6151
R10491 gnd.n2675 gnd.n2674 10.6151
R10492 gnd.n2674 gnd.n2671 10.6151
R10493 gnd.n2671 gnd.n2670 10.6151
R10494 gnd.n2670 gnd.n2667 10.6151
R10495 gnd.n2667 gnd.n2666 10.6151
R10496 gnd.n2666 gnd.n2663 10.6151
R10497 gnd.n2663 gnd.n2662 10.6151
R10498 gnd.n2662 gnd.n2659 10.6151
R10499 gnd.n2659 gnd.n2658 10.6151
R10500 gnd.n2658 gnd.n2655 10.6151
R10501 gnd.n2655 gnd.n2654 10.6151
R10502 gnd.n2654 gnd.n2651 10.6151
R10503 gnd.n2651 gnd.n2650 10.6151
R10504 gnd.n2650 gnd.n2647 10.6151
R10505 gnd.n2647 gnd.n2646 10.6151
R10506 gnd.n2646 gnd.n2643 10.6151
R10507 gnd.n2643 gnd.n2642 10.6151
R10508 gnd.n2642 gnd.n2639 10.6151
R10509 gnd.n2639 gnd.n2638 10.6151
R10510 gnd.n2638 gnd.n2635 10.6151
R10511 gnd.n2635 gnd.n2634 10.6151
R10512 gnd.n2634 gnd.n2631 10.6151
R10513 gnd.n2631 gnd.n1833 10.6151
R10514 gnd.n2969 gnd.n2968 10.6151
R10515 gnd.n2968 gnd.n1859 10.6151
R10516 gnd.n2697 gnd.n1859 10.6151
R10517 gnd.n2698 gnd.n2697 10.6151
R10518 gnd.n2701 gnd.n2698 10.6151
R10519 gnd.n2702 gnd.n2701 10.6151
R10520 gnd.n2705 gnd.n2702 10.6151
R10521 gnd.n2706 gnd.n2705 10.6151
R10522 gnd.n2709 gnd.n2706 10.6151
R10523 gnd.n2710 gnd.n2709 10.6151
R10524 gnd.n2713 gnd.n2710 10.6151
R10525 gnd.n2714 gnd.n2713 10.6151
R10526 gnd.n2717 gnd.n2714 10.6151
R10527 gnd.n2718 gnd.n2717 10.6151
R10528 gnd.n2721 gnd.n2718 10.6151
R10529 gnd.n2722 gnd.n2721 10.6151
R10530 gnd.n2725 gnd.n2722 10.6151
R10531 gnd.n2726 gnd.n2725 10.6151
R10532 gnd.n2729 gnd.n2726 10.6151
R10533 gnd.n2730 gnd.n2729 10.6151
R10534 gnd.n2733 gnd.n2730 10.6151
R10535 gnd.n2734 gnd.n2733 10.6151
R10536 gnd.n2737 gnd.n2734 10.6151
R10537 gnd.n2738 gnd.n2737 10.6151
R10538 gnd.n2741 gnd.n2738 10.6151
R10539 gnd.n2742 gnd.n2741 10.6151
R10540 gnd.n2745 gnd.n2742 10.6151
R10541 gnd.n2746 gnd.n2745 10.6151
R10542 gnd.n2750 gnd.n2749 10.6151
R10543 gnd.n2753 gnd.n2750 10.6151
R10544 gnd.n3708 gnd.n3707 10.6151
R10545 gnd.n3707 gnd.n3704 10.6151
R10546 gnd.n3704 gnd.n3703 10.6151
R10547 gnd.n3703 gnd.n3700 10.6151
R10548 gnd.n3700 gnd.n3699 10.6151
R10549 gnd.n3699 gnd.n3696 10.6151
R10550 gnd.n3696 gnd.n3695 10.6151
R10551 gnd.n3695 gnd.n3692 10.6151
R10552 gnd.n3692 gnd.n3691 10.6151
R10553 gnd.n3691 gnd.n3688 10.6151
R10554 gnd.n3688 gnd.n3687 10.6151
R10555 gnd.n3687 gnd.n3684 10.6151
R10556 gnd.n3684 gnd.n3683 10.6151
R10557 gnd.n3683 gnd.n3680 10.6151
R10558 gnd.n3680 gnd.n3679 10.6151
R10559 gnd.n3679 gnd.n3676 10.6151
R10560 gnd.n3676 gnd.n3675 10.6151
R10561 gnd.n3675 gnd.n3672 10.6151
R10562 gnd.n3672 gnd.n3671 10.6151
R10563 gnd.n3671 gnd.n3668 10.6151
R10564 gnd.n3668 gnd.n3667 10.6151
R10565 gnd.n3667 gnd.n3664 10.6151
R10566 gnd.n3664 gnd.n3663 10.6151
R10567 gnd.n3663 gnd.n3660 10.6151
R10568 gnd.n3660 gnd.n3659 10.6151
R10569 gnd.n3659 gnd.n3656 10.6151
R10570 gnd.n3656 gnd.n3655 10.6151
R10571 gnd.n3655 gnd.n3652 10.6151
R10572 gnd.n3650 gnd.n3647 10.6151
R10573 gnd.n3647 gnd.n1489 10.6151
R10574 gnd.n2973 gnd.n2972 10.6151
R10575 gnd.n2972 gnd.n2971 10.6151
R10576 gnd.n2971 gnd.n1815 10.6151
R10577 gnd.n2999 gnd.n1815 10.6151
R10578 gnd.n3000 gnd.n2999 10.6151
R10579 gnd.n3002 gnd.n3000 10.6151
R10580 gnd.n3002 gnd.n3001 10.6151
R10581 gnd.n3001 gnd.n1793 10.6151
R10582 gnd.n3038 gnd.n1793 10.6151
R10583 gnd.n3039 gnd.n3038 10.6151
R10584 gnd.n3040 gnd.n3039 10.6151
R10585 gnd.n3040 gnd.n1778 10.6151
R10586 gnd.n3055 gnd.n1778 10.6151
R10587 gnd.n3056 gnd.n3055 10.6151
R10588 gnd.n3058 gnd.n3056 10.6151
R10589 gnd.n3058 gnd.n3057 10.6151
R10590 gnd.n3057 gnd.n1759 10.6151
R10591 gnd.n3125 gnd.n1759 10.6151
R10592 gnd.n3126 gnd.n3125 10.6151
R10593 gnd.n3127 gnd.n3126 10.6151
R10594 gnd.n3127 gnd.n1744 10.6151
R10595 gnd.n3142 gnd.n1744 10.6151
R10596 gnd.n3143 gnd.n3142 10.6151
R10597 gnd.n3144 gnd.n3143 10.6151
R10598 gnd.n3144 gnd.n1731 10.6151
R10599 gnd.n3158 gnd.n1731 10.6151
R10600 gnd.n3159 gnd.n3158 10.6151
R10601 gnd.n3161 gnd.n3159 10.6151
R10602 gnd.n3161 gnd.n3160 10.6151
R10603 gnd.n3160 gnd.n1708 10.6151
R10604 gnd.n3190 gnd.n1708 10.6151
R10605 gnd.n3191 gnd.n3190 10.6151
R10606 gnd.n3192 gnd.n3191 10.6151
R10607 gnd.n3192 gnd.n1695 10.6151
R10608 gnd.n3209 gnd.n1695 10.6151
R10609 gnd.n3210 gnd.n3209 10.6151
R10610 gnd.n3211 gnd.n3210 10.6151
R10611 gnd.n3211 gnd.n1679 10.6151
R10612 gnd.n3233 gnd.n1679 10.6151
R10613 gnd.n3234 gnd.n3233 10.6151
R10614 gnd.n3236 gnd.n3234 10.6151
R10615 gnd.n3236 gnd.n3235 10.6151
R10616 gnd.n3235 gnd.n1662 10.6151
R10617 gnd.n3276 gnd.n1662 10.6151
R10618 gnd.n3277 gnd.n3276 10.6151
R10619 gnd.n3278 gnd.n3277 10.6151
R10620 gnd.n3278 gnd.n1650 10.6151
R10621 gnd.n3292 gnd.n1650 10.6151
R10622 gnd.n3293 gnd.n3292 10.6151
R10623 gnd.n3295 gnd.n3293 10.6151
R10624 gnd.n3295 gnd.n3294 10.6151
R10625 gnd.n3294 gnd.n1624 10.6151
R10626 gnd.n3326 gnd.n1624 10.6151
R10627 gnd.n3327 gnd.n3326 10.6151
R10628 gnd.n3329 gnd.n3327 10.6151
R10629 gnd.n3329 gnd.n3328 10.6151
R10630 gnd.n3328 gnd.n1532 10.6151
R10631 gnd.n3624 gnd.n1532 10.6151
R10632 gnd.n3625 gnd.n3624 10.6151
R10633 gnd.n3710 gnd.n3625 10.6151
R10634 gnd.n5078 gnd.t147 10.5161
R10635 gnd.n5750 gnd.t15 10.5161
R10636 gnd.t302 gnd.n4812 10.5161
R10637 gnd.n2163 gnd.t173 10.5161
R10638 gnd.n6634 gnd.t183 10.5161
R10639 gnd.n4779 gnd.n4763 10.4732
R10640 gnd.n4747 gnd.n4731 10.4732
R10641 gnd.n4715 gnd.n4699 10.4732
R10642 gnd.n4684 gnd.n4668 10.4732
R10643 gnd.n4652 gnd.n4636 10.4732
R10644 gnd.n4620 gnd.n4604 10.4732
R10645 gnd.n4588 gnd.n4572 10.4732
R10646 gnd.n4557 gnd.n4541 10.4732
R10647 gnd.n2997 gnd.n1818 10.1975
R10648 gnd.n3053 gnd.t37 10.1975
R10649 gnd.n1728 gnd.n1719 10.1975
R10650 gnd.n3188 gnd.n3187 10.1975
R10651 gnd.n3265 gnd.t35 10.1975
R10652 gnd.n3342 gnd.n1618 10.1975
R10653 gnd.n5705 gnd.t292 9.87883
R10654 gnd.n2474 gnd.t157 9.87883
R10655 gnd.n2965 gnd.n1862 9.87883
R10656 gnd.t165 gnd.n1359 9.87883
R10657 gnd.n7057 gnd.n62 9.73455
R10658 gnd.n4783 gnd.n4782 9.69747
R10659 gnd.n4751 gnd.n4750 9.69747
R10660 gnd.n4719 gnd.n4718 9.69747
R10661 gnd.n4688 gnd.n4687 9.69747
R10662 gnd.n4656 gnd.n4655 9.69747
R10663 gnd.n4624 gnd.n4623 9.69747
R10664 gnd.n4592 gnd.n4591 9.69747
R10665 gnd.n4561 gnd.n4560 9.69747
R10666 gnd.n3129 gnd.n1757 9.56018
R10667 gnd.n3230 gnd.n1684 9.56018
R10668 gnd.t104 gnd.n1626 9.56018
R10669 gnd.n4202 gnd.n1197 9.45599
R10670 gnd.n3449 gnd.n3448 9.45599
R10671 gnd.n4789 gnd.n4788 9.45567
R10672 gnd.n4757 gnd.n4756 9.45567
R10673 gnd.n4725 gnd.n4724 9.45567
R10674 gnd.n4694 gnd.n4693 9.45567
R10675 gnd.n4662 gnd.n4661 9.45567
R10676 gnd.n4630 gnd.n4629 9.45567
R10677 gnd.n4598 gnd.n4597 9.45567
R10678 gnd.n4567 gnd.n4566 9.45567
R10679 gnd.n5340 gnd.n5339 9.39724
R10680 gnd.n4788 gnd.n4787 9.3005
R10681 gnd.n4761 gnd.n4760 9.3005
R10682 gnd.n4782 gnd.n4781 9.3005
R10683 gnd.n4780 gnd.n4779 9.3005
R10684 gnd.n4765 gnd.n4764 9.3005
R10685 gnd.n4774 gnd.n4773 9.3005
R10686 gnd.n4772 gnd.n4771 9.3005
R10687 gnd.n4756 gnd.n4755 9.3005
R10688 gnd.n4729 gnd.n4728 9.3005
R10689 gnd.n4750 gnd.n4749 9.3005
R10690 gnd.n4748 gnd.n4747 9.3005
R10691 gnd.n4733 gnd.n4732 9.3005
R10692 gnd.n4742 gnd.n4741 9.3005
R10693 gnd.n4740 gnd.n4739 9.3005
R10694 gnd.n4724 gnd.n4723 9.3005
R10695 gnd.n4697 gnd.n4696 9.3005
R10696 gnd.n4718 gnd.n4717 9.3005
R10697 gnd.n4716 gnd.n4715 9.3005
R10698 gnd.n4701 gnd.n4700 9.3005
R10699 gnd.n4710 gnd.n4709 9.3005
R10700 gnd.n4708 gnd.n4707 9.3005
R10701 gnd.n4693 gnd.n4692 9.3005
R10702 gnd.n4666 gnd.n4665 9.3005
R10703 gnd.n4687 gnd.n4686 9.3005
R10704 gnd.n4685 gnd.n4684 9.3005
R10705 gnd.n4670 gnd.n4669 9.3005
R10706 gnd.n4679 gnd.n4678 9.3005
R10707 gnd.n4677 gnd.n4676 9.3005
R10708 gnd.n4661 gnd.n4660 9.3005
R10709 gnd.n4634 gnd.n4633 9.3005
R10710 gnd.n4655 gnd.n4654 9.3005
R10711 gnd.n4653 gnd.n4652 9.3005
R10712 gnd.n4638 gnd.n4637 9.3005
R10713 gnd.n4647 gnd.n4646 9.3005
R10714 gnd.n4645 gnd.n4644 9.3005
R10715 gnd.n4629 gnd.n4628 9.3005
R10716 gnd.n4602 gnd.n4601 9.3005
R10717 gnd.n4623 gnd.n4622 9.3005
R10718 gnd.n4621 gnd.n4620 9.3005
R10719 gnd.n4606 gnd.n4605 9.3005
R10720 gnd.n4615 gnd.n4614 9.3005
R10721 gnd.n4613 gnd.n4612 9.3005
R10722 gnd.n4597 gnd.n4596 9.3005
R10723 gnd.n4570 gnd.n4569 9.3005
R10724 gnd.n4591 gnd.n4590 9.3005
R10725 gnd.n4589 gnd.n4588 9.3005
R10726 gnd.n4574 gnd.n4573 9.3005
R10727 gnd.n4583 gnd.n4582 9.3005
R10728 gnd.n4581 gnd.n4580 9.3005
R10729 gnd.n4566 gnd.n4565 9.3005
R10730 gnd.n4539 gnd.n4538 9.3005
R10731 gnd.n4560 gnd.n4559 9.3005
R10732 gnd.n4558 gnd.n4557 9.3005
R10733 gnd.n4543 gnd.n4542 9.3005
R10734 gnd.n4552 gnd.n4551 9.3005
R10735 gnd.n4550 gnd.n4549 9.3005
R10736 gnd.n5881 gnd.n4450 9.3005
R10737 gnd.n5880 gnd.n4452 9.3005
R10738 gnd.n4456 gnd.n4453 9.3005
R10739 gnd.n5875 gnd.n4457 9.3005
R10740 gnd.n5874 gnd.n4458 9.3005
R10741 gnd.n5873 gnd.n4459 9.3005
R10742 gnd.n4463 gnd.n4460 9.3005
R10743 gnd.n5868 gnd.n4464 9.3005
R10744 gnd.n5867 gnd.n4465 9.3005
R10745 gnd.n5866 gnd.n4466 9.3005
R10746 gnd.n4470 gnd.n4467 9.3005
R10747 gnd.n5861 gnd.n4471 9.3005
R10748 gnd.n5860 gnd.n4472 9.3005
R10749 gnd.n5859 gnd.n4473 9.3005
R10750 gnd.n4478 gnd.n4476 9.3005
R10751 gnd.n5854 gnd.n5853 9.3005
R10752 gnd.n5883 gnd.n5882 9.3005
R10753 gnd.n5459 gnd.n5458 9.3005
R10754 gnd.n5460 gnd.n5049 9.3005
R10755 gnd.n5464 gnd.n5461 9.3005
R10756 gnd.n5463 gnd.n5462 9.3005
R10757 gnd.n5026 gnd.n5025 9.3005
R10758 gnd.n5490 gnd.n5489 9.3005
R10759 gnd.n5491 gnd.n5024 9.3005
R10760 gnd.n5495 gnd.n5492 9.3005
R10761 gnd.n5494 gnd.n5493 9.3005
R10762 gnd.n5000 gnd.n4999 9.3005
R10763 gnd.n5521 gnd.n5520 9.3005
R10764 gnd.n5522 gnd.n4998 9.3005
R10765 gnd.n5526 gnd.n5523 9.3005
R10766 gnd.n5525 gnd.n5524 9.3005
R10767 gnd.n4974 gnd.n4973 9.3005
R10768 gnd.n5552 gnd.n5551 9.3005
R10769 gnd.n5553 gnd.n4972 9.3005
R10770 gnd.n5557 gnd.n5554 9.3005
R10771 gnd.n5556 gnd.n5555 9.3005
R10772 gnd.n4948 gnd.n4947 9.3005
R10773 gnd.n5583 gnd.n5582 9.3005
R10774 gnd.n5584 gnd.n4946 9.3005
R10775 gnd.n5588 gnd.n5585 9.3005
R10776 gnd.n5587 gnd.n5586 9.3005
R10777 gnd.n4923 gnd.n4922 9.3005
R10778 gnd.n5614 gnd.n5613 9.3005
R10779 gnd.n5615 gnd.n4921 9.3005
R10780 gnd.n5619 gnd.n5616 9.3005
R10781 gnd.n5618 gnd.n5617 9.3005
R10782 gnd.n4899 gnd.n4898 9.3005
R10783 gnd.n5644 gnd.n5643 9.3005
R10784 gnd.n5645 gnd.n4897 9.3005
R10785 gnd.n5649 gnd.n5646 9.3005
R10786 gnd.n5648 gnd.n5647 9.3005
R10787 gnd.n4867 gnd.n4866 9.3005
R10788 gnd.n5685 gnd.n5684 9.3005
R10789 gnd.n5686 gnd.n4865 9.3005
R10790 gnd.n5693 gnd.n5687 9.3005
R10791 gnd.n5692 gnd.n5688 9.3005
R10792 gnd.n5691 gnd.n5689 9.3005
R10793 gnd.n4837 gnd.n4836 9.3005
R10794 gnd.n5732 gnd.n5731 9.3005
R10795 gnd.n5733 gnd.n4835 9.3005
R10796 gnd.n5739 gnd.n5734 9.3005
R10797 gnd.n5738 gnd.n5735 9.3005
R10798 gnd.n5737 gnd.n5736 9.3005
R10799 gnd.n4810 gnd.n4809 9.3005
R10800 gnd.n5776 gnd.n5775 9.3005
R10801 gnd.n5777 gnd.n4808 9.3005
R10802 gnd.n5781 gnd.n5778 9.3005
R10803 gnd.n5780 gnd.n5779 9.3005
R10804 gnd.n4449 gnd.n4448 9.3005
R10805 gnd.n5885 gnd.n5884 9.3005
R10806 gnd.n5051 gnd.n5050 9.3005
R10807 gnd.n5403 gnd.n5402 9.3005
R10808 gnd.n5406 gnd.n5398 9.3005
R10809 gnd.n5407 gnd.n5397 9.3005
R10810 gnd.n5410 gnd.n5396 9.3005
R10811 gnd.n5411 gnd.n5395 9.3005
R10812 gnd.n5414 gnd.n5394 9.3005
R10813 gnd.n5415 gnd.n5393 9.3005
R10814 gnd.n5418 gnd.n5392 9.3005
R10815 gnd.n5419 gnd.n5391 9.3005
R10816 gnd.n5422 gnd.n5390 9.3005
R10817 gnd.n5423 gnd.n5389 9.3005
R10818 gnd.n5426 gnd.n5388 9.3005
R10819 gnd.n5428 gnd.n5387 9.3005
R10820 gnd.n5429 gnd.n5386 9.3005
R10821 gnd.n5430 gnd.n5385 9.3005
R10822 gnd.n5431 gnd.n5384 9.3005
R10823 gnd.n5399 gnd.n5067 9.3005
R10824 gnd.n5449 gnd.n5448 9.3005
R10825 gnd.n5450 gnd.n5044 9.3005
R10826 gnd.n5469 gnd.n5468 9.3005
R10827 gnd.n5471 gnd.n5036 9.3005
R10828 gnd.n5478 gnd.n5037 9.3005
R10829 gnd.n5480 gnd.n5479 9.3005
R10830 gnd.n5481 gnd.n5017 9.3005
R10831 gnd.n5500 gnd.n5499 9.3005
R10832 gnd.n5502 gnd.n5010 9.3005
R10833 gnd.n5509 gnd.n5011 9.3005
R10834 gnd.n5511 gnd.n5510 9.3005
R10835 gnd.n5512 gnd.n4991 9.3005
R10836 gnd.n5531 gnd.n5530 9.3005
R10837 gnd.n5533 gnd.n4984 9.3005
R10838 gnd.n5540 gnd.n4985 9.3005
R10839 gnd.n5542 gnd.n5541 9.3005
R10840 gnd.n5543 gnd.n4966 9.3005
R10841 gnd.n5562 gnd.n5561 9.3005
R10842 gnd.n5564 gnd.n4958 9.3005
R10843 gnd.n5571 gnd.n4959 9.3005
R10844 gnd.n5573 gnd.n5572 9.3005
R10845 gnd.n5574 gnd.n4941 9.3005
R10846 gnd.n5593 gnd.n5592 9.3005
R10847 gnd.n5595 gnd.n4933 9.3005
R10848 gnd.n5602 gnd.n4934 9.3005
R10849 gnd.n5604 gnd.n5603 9.3005
R10850 gnd.n5605 gnd.n4916 9.3005
R10851 gnd.n5624 gnd.n5623 9.3005
R10852 gnd.n5626 gnd.n4908 9.3005
R10853 gnd.n5633 gnd.n4909 9.3005
R10854 gnd.n5635 gnd.n5634 9.3005
R10855 gnd.n5636 gnd.n4892 9.3005
R10856 gnd.n5654 gnd.n5653 9.3005
R10857 gnd.n5656 gnd.n4877 9.3005
R10858 gnd.n5674 gnd.n4879 9.3005
R10859 gnd.n5675 gnd.n4874 9.3005
R10860 gnd.n5677 gnd.n5676 9.3005
R10861 gnd.n4875 gnd.n4861 9.3005
R10862 gnd.n4859 gnd.n4857 9.3005
R10863 gnd.n5700 gnd.n5699 9.3005
R10864 gnd.n4842 gnd.n4841 9.3005
R10865 gnd.n5725 gnd.n5721 9.3005
R10866 gnd.n5724 gnd.n5723 9.3005
R10867 gnd.n4830 gnd.n4828 9.3005
R10868 gnd.n5745 gnd.n5744 9.3005
R10869 gnd.n4815 gnd.n4814 9.3005
R10870 gnd.n5769 gnd.n5768 9.3005
R10871 gnd.n5766 gnd.n4794 9.3005
R10872 gnd.n5787 gnd.n5786 9.3005
R10873 gnd.n4796 gnd.n4795 9.3005
R10874 gnd.n4803 gnd.n4799 9.3005
R10875 gnd.n4802 gnd.n4800 9.3005
R10876 gnd.n4801 gnd.n4479 9.3005
R10877 gnd.n5447 gnd.n5061 9.3005
R10878 gnd.n5849 gnd.n4480 9.3005
R10879 gnd.n5848 gnd.n4482 9.3005
R10880 gnd.n4486 gnd.n4483 9.3005
R10881 gnd.n5843 gnd.n4487 9.3005
R10882 gnd.n5842 gnd.n4488 9.3005
R10883 gnd.n5841 gnd.n4489 9.3005
R10884 gnd.n4493 gnd.n4490 9.3005
R10885 gnd.n5836 gnd.n4494 9.3005
R10886 gnd.n5835 gnd.n4495 9.3005
R10887 gnd.n5834 gnd.n4496 9.3005
R10888 gnd.n4500 gnd.n4497 9.3005
R10889 gnd.n5829 gnd.n4501 9.3005
R10890 gnd.n5828 gnd.n4502 9.3005
R10891 gnd.n5827 gnd.n4503 9.3005
R10892 gnd.n4507 gnd.n4504 9.3005
R10893 gnd.n5822 gnd.n4508 9.3005
R10894 gnd.n5821 gnd.n4509 9.3005
R10895 gnd.n5820 gnd.n4510 9.3005
R10896 gnd.n4514 gnd.n4511 9.3005
R10897 gnd.n5815 gnd.n4515 9.3005
R10898 gnd.n5814 gnd.n4516 9.3005
R10899 gnd.n5813 gnd.n4517 9.3005
R10900 gnd.n4524 gnd.n4522 9.3005
R10901 gnd.n5808 gnd.n4525 9.3005
R10902 gnd.n5807 gnd.n4526 9.3005
R10903 gnd.n5806 gnd.n5803 9.3005
R10904 gnd.n5851 gnd.n5850 9.3005
R10905 gnd.n5278 gnd.n5257 9.3005
R10906 gnd.n5277 gnd.n5259 9.3005
R10907 gnd.n5275 gnd.n5260 9.3005
R10908 gnd.n5274 gnd.n5261 9.3005
R10909 gnd.n5270 gnd.n5262 9.3005
R10910 gnd.n5269 gnd.n5263 9.3005
R10911 gnd.n5268 gnd.n5264 9.3005
R10912 gnd.n5266 gnd.n5265 9.3005
R10913 gnd.n4885 gnd.n4884 9.3005
R10914 gnd.n5664 gnd.n5663 9.3005
R10915 gnd.n5665 gnd.n4883 9.3005
R10916 gnd.n5669 gnd.n5666 9.3005
R10917 gnd.n5668 gnd.n5667 9.3005
R10918 gnd.n4850 gnd.n4849 9.3005
R10919 gnd.n5708 gnd.n5707 9.3005
R10920 gnd.n5709 gnd.n4848 9.3005
R10921 gnd.n5713 gnd.n5710 9.3005
R10922 gnd.n5712 gnd.n5711 9.3005
R10923 gnd.n4823 gnd.n4822 9.3005
R10924 gnd.n5753 gnd.n5752 9.3005
R10925 gnd.n5754 gnd.n4821 9.3005
R10926 gnd.n5758 gnd.n5755 9.3005
R10927 gnd.n5757 gnd.n5756 9.3005
R10928 gnd.n4530 gnd.n4529 9.3005
R10929 gnd.n5794 gnd.n5793 9.3005
R10930 gnd.n5795 gnd.n4528 9.3005
R10931 gnd.n5797 gnd.n5796 9.3005
R10932 gnd.n5800 gnd.n4527 9.3005
R10933 gnd.n5802 gnd.n5801 9.3005
R10934 gnd.n5204 gnd.n5098 9.3005
R10935 gnd.n5206 gnd.n5205 9.3005
R10936 gnd.n5088 gnd.n5087 9.3005
R10937 gnd.n5219 gnd.n5218 9.3005
R10938 gnd.n5220 gnd.n5086 9.3005
R10939 gnd.n5222 gnd.n5221 9.3005
R10940 gnd.n5075 gnd.n5074 9.3005
R10941 gnd.n5235 gnd.n5234 9.3005
R10942 gnd.n5236 gnd.n5073 9.3005
R10943 gnd.n5373 gnd.n5237 9.3005
R10944 gnd.n5372 gnd.n5238 9.3005
R10945 gnd.n5371 gnd.n5239 9.3005
R10946 gnd.n5370 gnd.n5240 9.3005
R10947 gnd.n5368 gnd.n5241 9.3005
R10948 gnd.n5367 gnd.n5242 9.3005
R10949 gnd.n5363 gnd.n5243 9.3005
R10950 gnd.n5362 gnd.n5244 9.3005
R10951 gnd.n5361 gnd.n5245 9.3005
R10952 gnd.n5359 gnd.n5246 9.3005
R10953 gnd.n5358 gnd.n5247 9.3005
R10954 gnd.n5355 gnd.n5248 9.3005
R10955 gnd.n5354 gnd.n5249 9.3005
R10956 gnd.n5353 gnd.n5250 9.3005
R10957 gnd.n5351 gnd.n5251 9.3005
R10958 gnd.n5350 gnd.n5252 9.3005
R10959 gnd.n5347 gnd.n5253 9.3005
R10960 gnd.n5346 gnd.n5254 9.3005
R10961 gnd.n5345 gnd.n5255 9.3005
R10962 gnd.n5203 gnd.n5202 9.3005
R10963 gnd.n5143 gnd.n5142 9.3005
R10964 gnd.n5148 gnd.n5140 9.3005
R10965 gnd.n5149 gnd.n5139 9.3005
R10966 gnd.n5151 gnd.n5136 9.3005
R10967 gnd.n5135 gnd.n5133 9.3005
R10968 gnd.n5157 gnd.n5132 9.3005
R10969 gnd.n5158 gnd.n5131 9.3005
R10970 gnd.n5159 gnd.n5130 9.3005
R10971 gnd.n5129 gnd.n5127 9.3005
R10972 gnd.n5165 gnd.n5126 9.3005
R10973 gnd.n5166 gnd.n5125 9.3005
R10974 gnd.n5167 gnd.n5124 9.3005
R10975 gnd.n5123 gnd.n5121 9.3005
R10976 gnd.n5173 gnd.n5120 9.3005
R10977 gnd.n5174 gnd.n5119 9.3005
R10978 gnd.n5175 gnd.n5118 9.3005
R10979 gnd.n5117 gnd.n5115 9.3005
R10980 gnd.n5181 gnd.n5114 9.3005
R10981 gnd.n5182 gnd.n5113 9.3005
R10982 gnd.n5183 gnd.n5112 9.3005
R10983 gnd.n5111 gnd.n5109 9.3005
R10984 gnd.n5188 gnd.n5108 9.3005
R10985 gnd.n5189 gnd.n5107 9.3005
R10986 gnd.n5106 gnd.n5104 9.3005
R10987 gnd.n5194 gnd.n5103 9.3005
R10988 gnd.n5196 gnd.n5195 9.3005
R10989 gnd.n5141 gnd.n5099 9.3005
R10990 gnd.n5094 gnd.n5093 9.3005
R10991 gnd.n5211 gnd.n5210 9.3005
R10992 gnd.n5212 gnd.n5092 9.3005
R10993 gnd.n5214 gnd.n5213 9.3005
R10994 gnd.n5082 gnd.n5081 9.3005
R10995 gnd.n5227 gnd.n5226 9.3005
R10996 gnd.n5228 gnd.n5080 9.3005
R10997 gnd.n5230 gnd.n5229 9.3005
R10998 gnd.n5069 gnd.n5068 9.3005
R10999 gnd.n5438 gnd.n5437 9.3005
R11000 gnd.n5440 gnd.n5066 9.3005
R11001 gnd.n5442 gnd.n5441 9.3005
R11002 gnd.n5060 gnd.n5059 9.3005
R11003 gnd.n5453 gnd.n5451 9.3005
R11004 gnd.n5452 gnd.n5043 9.3005
R11005 gnd.n5470 gnd.n5042 9.3005
R11006 gnd.n5473 gnd.n5472 9.3005
R11007 gnd.n5035 gnd.n5034 9.3005
R11008 gnd.n5484 gnd.n5482 9.3005
R11009 gnd.n5483 gnd.n5016 9.3005
R11010 gnd.n5501 gnd.n5015 9.3005
R11011 gnd.n5504 gnd.n5503 9.3005
R11012 gnd.n5009 gnd.n5008 9.3005
R11013 gnd.n5515 gnd.n5513 9.3005
R11014 gnd.n5514 gnd.n4990 9.3005
R11015 gnd.n5532 gnd.n4989 9.3005
R11016 gnd.n5535 gnd.n5534 9.3005
R11017 gnd.n4983 gnd.n4982 9.3005
R11018 gnd.n5546 gnd.n5544 9.3005
R11019 gnd.n5545 gnd.n4965 9.3005
R11020 gnd.n5563 gnd.n4964 9.3005
R11021 gnd.n5566 gnd.n5565 9.3005
R11022 gnd.n4957 gnd.n4956 9.3005
R11023 gnd.n5577 gnd.n5575 9.3005
R11024 gnd.n5576 gnd.n4940 9.3005
R11025 gnd.n5594 gnd.n4939 9.3005
R11026 gnd.n5597 gnd.n5596 9.3005
R11027 gnd.n4932 gnd.n4931 9.3005
R11028 gnd.n5608 gnd.n5606 9.3005
R11029 gnd.n5607 gnd.n4915 9.3005
R11030 gnd.n5625 gnd.n4914 9.3005
R11031 gnd.n5628 gnd.n5627 9.3005
R11032 gnd.n4907 gnd.n4906 9.3005
R11033 gnd.n5638 gnd.n5637 9.3005
R11034 gnd.n4891 gnd.n4890 9.3005
R11035 gnd.n5659 gnd.n5655 9.3005
R11036 gnd.n5658 gnd.n5657 9.3005
R11037 gnd.n4878 gnd.n4873 9.3005
R11038 gnd.n5679 gnd.n5678 9.3005
R11039 gnd.n4876 gnd.n4855 9.3005
R11040 gnd.n5703 gnd.n4856 9.3005
R11041 gnd.n5702 gnd.n5701 9.3005
R11042 gnd.n4858 gnd.n4843 9.3005
R11043 gnd.n5720 gnd.n5719 9.3005
R11044 gnd.n5722 gnd.n4826 9.3005
R11045 gnd.n5748 gnd.n4827 9.3005
R11046 gnd.n5747 gnd.n5746 9.3005
R11047 gnd.n4829 gnd.n4816 9.3005
R11048 gnd.n5765 gnd.n5764 9.3005
R11049 gnd.n5767 gnd.n4536 9.3005
R11050 gnd.n5789 gnd.n5788 9.3005
R11051 gnd.n4793 gnd.n849 9.3005
R11052 gnd.n5892 gnd.n850 9.3005
R11053 gnd.n5891 gnd.n851 9.3005
R11054 gnd.n5890 gnd.n852 9.3005
R11055 gnd.n5198 gnd.n5197 9.3005
R11056 gnd.n6067 gnd.n6066 9.3005
R11057 gnd.n6068 gnd.n674 9.3005
R11058 gnd.n6070 gnd.n6069 9.3005
R11059 gnd.n670 gnd.n669 9.3005
R11060 gnd.n6077 gnd.n6076 9.3005
R11061 gnd.n6078 gnd.n668 9.3005
R11062 gnd.n6080 gnd.n6079 9.3005
R11063 gnd.n664 gnd.n663 9.3005
R11064 gnd.n6087 gnd.n6086 9.3005
R11065 gnd.n6088 gnd.n662 9.3005
R11066 gnd.n6090 gnd.n6089 9.3005
R11067 gnd.n658 gnd.n657 9.3005
R11068 gnd.n6097 gnd.n6096 9.3005
R11069 gnd.n6098 gnd.n656 9.3005
R11070 gnd.n6100 gnd.n6099 9.3005
R11071 gnd.n652 gnd.n651 9.3005
R11072 gnd.n6107 gnd.n6106 9.3005
R11073 gnd.n6108 gnd.n650 9.3005
R11074 gnd.n6110 gnd.n6109 9.3005
R11075 gnd.n646 gnd.n645 9.3005
R11076 gnd.n6117 gnd.n6116 9.3005
R11077 gnd.n6118 gnd.n644 9.3005
R11078 gnd.n6120 gnd.n6119 9.3005
R11079 gnd.n640 gnd.n639 9.3005
R11080 gnd.n6127 gnd.n6126 9.3005
R11081 gnd.n6128 gnd.n638 9.3005
R11082 gnd.n6130 gnd.n6129 9.3005
R11083 gnd.n634 gnd.n633 9.3005
R11084 gnd.n6137 gnd.n6136 9.3005
R11085 gnd.n6138 gnd.n632 9.3005
R11086 gnd.n6140 gnd.n6139 9.3005
R11087 gnd.n628 gnd.n627 9.3005
R11088 gnd.n6147 gnd.n6146 9.3005
R11089 gnd.n6148 gnd.n626 9.3005
R11090 gnd.n6150 gnd.n6149 9.3005
R11091 gnd.n622 gnd.n621 9.3005
R11092 gnd.n6157 gnd.n6156 9.3005
R11093 gnd.n6158 gnd.n620 9.3005
R11094 gnd.n6160 gnd.n6159 9.3005
R11095 gnd.n616 gnd.n615 9.3005
R11096 gnd.n6167 gnd.n6166 9.3005
R11097 gnd.n6168 gnd.n614 9.3005
R11098 gnd.n6170 gnd.n6169 9.3005
R11099 gnd.n610 gnd.n609 9.3005
R11100 gnd.n6177 gnd.n6176 9.3005
R11101 gnd.n6178 gnd.n608 9.3005
R11102 gnd.n6180 gnd.n6179 9.3005
R11103 gnd.n604 gnd.n603 9.3005
R11104 gnd.n6187 gnd.n6186 9.3005
R11105 gnd.n6188 gnd.n602 9.3005
R11106 gnd.n6190 gnd.n6189 9.3005
R11107 gnd.n598 gnd.n597 9.3005
R11108 gnd.n6197 gnd.n6196 9.3005
R11109 gnd.n6198 gnd.n596 9.3005
R11110 gnd.n6200 gnd.n6199 9.3005
R11111 gnd.n592 gnd.n591 9.3005
R11112 gnd.n6207 gnd.n6206 9.3005
R11113 gnd.n6208 gnd.n590 9.3005
R11114 gnd.n6210 gnd.n6209 9.3005
R11115 gnd.n586 gnd.n585 9.3005
R11116 gnd.n6217 gnd.n6216 9.3005
R11117 gnd.n6218 gnd.n584 9.3005
R11118 gnd.n6220 gnd.n6219 9.3005
R11119 gnd.n580 gnd.n579 9.3005
R11120 gnd.n6227 gnd.n6226 9.3005
R11121 gnd.n6228 gnd.n578 9.3005
R11122 gnd.n6230 gnd.n6229 9.3005
R11123 gnd.n574 gnd.n573 9.3005
R11124 gnd.n6237 gnd.n6236 9.3005
R11125 gnd.n6238 gnd.n572 9.3005
R11126 gnd.n6240 gnd.n6239 9.3005
R11127 gnd.n568 gnd.n567 9.3005
R11128 gnd.n6247 gnd.n6246 9.3005
R11129 gnd.n6248 gnd.n566 9.3005
R11130 gnd.n6250 gnd.n6249 9.3005
R11131 gnd.n562 gnd.n561 9.3005
R11132 gnd.n6257 gnd.n6256 9.3005
R11133 gnd.n6258 gnd.n560 9.3005
R11134 gnd.n6260 gnd.n6259 9.3005
R11135 gnd.n556 gnd.n555 9.3005
R11136 gnd.n6267 gnd.n6266 9.3005
R11137 gnd.n6268 gnd.n554 9.3005
R11138 gnd.n6270 gnd.n6269 9.3005
R11139 gnd.n550 gnd.n549 9.3005
R11140 gnd.n6277 gnd.n6276 9.3005
R11141 gnd.n6278 gnd.n548 9.3005
R11142 gnd.n6280 gnd.n6279 9.3005
R11143 gnd.n544 gnd.n543 9.3005
R11144 gnd.n6287 gnd.n6286 9.3005
R11145 gnd.n6288 gnd.n542 9.3005
R11146 gnd.n6290 gnd.n6289 9.3005
R11147 gnd.n538 gnd.n537 9.3005
R11148 gnd.n6297 gnd.n6296 9.3005
R11149 gnd.n6298 gnd.n536 9.3005
R11150 gnd.n6300 gnd.n6299 9.3005
R11151 gnd.n532 gnd.n531 9.3005
R11152 gnd.n6307 gnd.n6306 9.3005
R11153 gnd.n6308 gnd.n530 9.3005
R11154 gnd.n6310 gnd.n6309 9.3005
R11155 gnd.n526 gnd.n525 9.3005
R11156 gnd.n6317 gnd.n6316 9.3005
R11157 gnd.n6318 gnd.n524 9.3005
R11158 gnd.n6320 gnd.n6319 9.3005
R11159 gnd.n520 gnd.n519 9.3005
R11160 gnd.n6327 gnd.n6326 9.3005
R11161 gnd.n6328 gnd.n518 9.3005
R11162 gnd.n6330 gnd.n6329 9.3005
R11163 gnd.n514 gnd.n513 9.3005
R11164 gnd.n6337 gnd.n6336 9.3005
R11165 gnd.n6338 gnd.n512 9.3005
R11166 gnd.n6340 gnd.n6339 9.3005
R11167 gnd.n508 gnd.n507 9.3005
R11168 gnd.n6347 gnd.n6346 9.3005
R11169 gnd.n6348 gnd.n506 9.3005
R11170 gnd.n6350 gnd.n6349 9.3005
R11171 gnd.n502 gnd.n501 9.3005
R11172 gnd.n6357 gnd.n6356 9.3005
R11173 gnd.n6358 gnd.n500 9.3005
R11174 gnd.n6360 gnd.n6359 9.3005
R11175 gnd.n496 gnd.n495 9.3005
R11176 gnd.n6367 gnd.n6366 9.3005
R11177 gnd.n6368 gnd.n494 9.3005
R11178 gnd.n6370 gnd.n6369 9.3005
R11179 gnd.n490 gnd.n489 9.3005
R11180 gnd.n6377 gnd.n6376 9.3005
R11181 gnd.n6378 gnd.n488 9.3005
R11182 gnd.n6380 gnd.n6379 9.3005
R11183 gnd.n484 gnd.n483 9.3005
R11184 gnd.n6387 gnd.n6386 9.3005
R11185 gnd.n6388 gnd.n482 9.3005
R11186 gnd.n6390 gnd.n6389 9.3005
R11187 gnd.n478 gnd.n477 9.3005
R11188 gnd.n6397 gnd.n6396 9.3005
R11189 gnd.n6398 gnd.n476 9.3005
R11190 gnd.n6400 gnd.n6399 9.3005
R11191 gnd.n472 gnd.n471 9.3005
R11192 gnd.n6407 gnd.n6406 9.3005
R11193 gnd.n6408 gnd.n470 9.3005
R11194 gnd.n6411 gnd.n6410 9.3005
R11195 gnd.n6409 gnd.n466 9.3005
R11196 gnd.n6417 gnd.n465 9.3005
R11197 gnd.n6419 gnd.n6418 9.3005
R11198 gnd.n461 gnd.n460 9.3005
R11199 gnd.n6428 gnd.n6427 9.3005
R11200 gnd.n6429 gnd.n459 9.3005
R11201 gnd.n6431 gnd.n6430 9.3005
R11202 gnd.n455 gnd.n454 9.3005
R11203 gnd.n6438 gnd.n6437 9.3005
R11204 gnd.n6439 gnd.n453 9.3005
R11205 gnd.n6441 gnd.n6440 9.3005
R11206 gnd.n449 gnd.n448 9.3005
R11207 gnd.n6448 gnd.n6447 9.3005
R11208 gnd.n6449 gnd.n447 9.3005
R11209 gnd.n6451 gnd.n6450 9.3005
R11210 gnd.n443 gnd.n442 9.3005
R11211 gnd.n6458 gnd.n6457 9.3005
R11212 gnd.n6459 gnd.n441 9.3005
R11213 gnd.n6461 gnd.n6460 9.3005
R11214 gnd.n437 gnd.n436 9.3005
R11215 gnd.n6468 gnd.n6467 9.3005
R11216 gnd.n6469 gnd.n435 9.3005
R11217 gnd.n6471 gnd.n6470 9.3005
R11218 gnd.n431 gnd.n430 9.3005
R11219 gnd.n6478 gnd.n6477 9.3005
R11220 gnd.n6479 gnd.n429 9.3005
R11221 gnd.n6481 gnd.n6480 9.3005
R11222 gnd.n425 gnd.n424 9.3005
R11223 gnd.n6488 gnd.n6487 9.3005
R11224 gnd.n6489 gnd.n423 9.3005
R11225 gnd.n6491 gnd.n6490 9.3005
R11226 gnd.n419 gnd.n418 9.3005
R11227 gnd.n6498 gnd.n6497 9.3005
R11228 gnd.n6499 gnd.n417 9.3005
R11229 gnd.n6501 gnd.n6500 9.3005
R11230 gnd.n413 gnd.n412 9.3005
R11231 gnd.n6508 gnd.n6507 9.3005
R11232 gnd.n6509 gnd.n411 9.3005
R11233 gnd.n6511 gnd.n6510 9.3005
R11234 gnd.n407 gnd.n406 9.3005
R11235 gnd.n6518 gnd.n6517 9.3005
R11236 gnd.n6519 gnd.n405 9.3005
R11237 gnd.n6521 gnd.n6520 9.3005
R11238 gnd.n401 gnd.n400 9.3005
R11239 gnd.n6528 gnd.n6527 9.3005
R11240 gnd.n6529 gnd.n399 9.3005
R11241 gnd.n6531 gnd.n6530 9.3005
R11242 gnd.n395 gnd.n394 9.3005
R11243 gnd.n6538 gnd.n6537 9.3005
R11244 gnd.n6539 gnd.n393 9.3005
R11245 gnd.n6541 gnd.n6540 9.3005
R11246 gnd.n389 gnd.n388 9.3005
R11247 gnd.n6548 gnd.n6547 9.3005
R11248 gnd.n6549 gnd.n387 9.3005
R11249 gnd.n6551 gnd.n6550 9.3005
R11250 gnd.n383 gnd.n382 9.3005
R11251 gnd.n6558 gnd.n6557 9.3005
R11252 gnd.n6559 gnd.n381 9.3005
R11253 gnd.n6561 gnd.n6560 9.3005
R11254 gnd.n377 gnd.n376 9.3005
R11255 gnd.n6568 gnd.n6567 9.3005
R11256 gnd.n6569 gnd.n375 9.3005
R11257 gnd.n6571 gnd.n6570 9.3005
R11258 gnd.n371 gnd.n370 9.3005
R11259 gnd.n6578 gnd.n6577 9.3005
R11260 gnd.n6579 gnd.n369 9.3005
R11261 gnd.n6581 gnd.n6580 9.3005
R11262 gnd.n365 gnd.n364 9.3005
R11263 gnd.n6588 gnd.n6587 9.3005
R11264 gnd.n6589 gnd.n363 9.3005
R11265 gnd.n6591 gnd.n6590 9.3005
R11266 gnd.n359 gnd.n358 9.3005
R11267 gnd.n6598 gnd.n6597 9.3005
R11268 gnd.n6599 gnd.n357 9.3005
R11269 gnd.n6601 gnd.n6600 9.3005
R11270 gnd.n353 gnd.n352 9.3005
R11271 gnd.n6608 gnd.n6607 9.3005
R11272 gnd.n6609 gnd.n351 9.3005
R11273 gnd.n6611 gnd.n6610 9.3005
R11274 gnd.n347 gnd.n346 9.3005
R11275 gnd.n6618 gnd.n6617 9.3005
R11276 gnd.n6619 gnd.n345 9.3005
R11277 gnd.n6621 gnd.n6620 9.3005
R11278 gnd.n341 gnd.n340 9.3005
R11279 gnd.n6629 gnd.n6628 9.3005
R11280 gnd.n6630 gnd.n339 9.3005
R11281 gnd.n6632 gnd.n6631 9.3005
R11282 gnd.n6421 gnd.n6420 9.3005
R11283 gnd.n7008 gnd.n108 9.3005
R11284 gnd.n7007 gnd.n110 9.3005
R11285 gnd.n114 gnd.n111 9.3005
R11286 gnd.n7002 gnd.n115 9.3005
R11287 gnd.n7001 gnd.n116 9.3005
R11288 gnd.n7000 gnd.n117 9.3005
R11289 gnd.n121 gnd.n118 9.3005
R11290 gnd.n6995 gnd.n122 9.3005
R11291 gnd.n6994 gnd.n123 9.3005
R11292 gnd.n6993 gnd.n124 9.3005
R11293 gnd.n128 gnd.n125 9.3005
R11294 gnd.n6988 gnd.n129 9.3005
R11295 gnd.n6987 gnd.n130 9.3005
R11296 gnd.n6986 gnd.n131 9.3005
R11297 gnd.n135 gnd.n132 9.3005
R11298 gnd.n6981 gnd.n136 9.3005
R11299 gnd.n6980 gnd.n137 9.3005
R11300 gnd.n6976 gnd.n138 9.3005
R11301 gnd.n142 gnd.n139 9.3005
R11302 gnd.n6971 gnd.n143 9.3005
R11303 gnd.n6970 gnd.n144 9.3005
R11304 gnd.n6969 gnd.n145 9.3005
R11305 gnd.n149 gnd.n146 9.3005
R11306 gnd.n6964 gnd.n150 9.3005
R11307 gnd.n6963 gnd.n151 9.3005
R11308 gnd.n6962 gnd.n152 9.3005
R11309 gnd.n156 gnd.n153 9.3005
R11310 gnd.n6957 gnd.n157 9.3005
R11311 gnd.n6956 gnd.n158 9.3005
R11312 gnd.n6955 gnd.n159 9.3005
R11313 gnd.n163 gnd.n160 9.3005
R11314 gnd.n6950 gnd.n164 9.3005
R11315 gnd.n6949 gnd.n165 9.3005
R11316 gnd.n6948 gnd.n166 9.3005
R11317 gnd.n170 gnd.n167 9.3005
R11318 gnd.n6943 gnd.n171 9.3005
R11319 gnd.n6942 gnd.n6941 9.3005
R11320 gnd.n6940 gnd.n174 9.3005
R11321 gnd.n7010 gnd.n7009 9.3005
R11322 gnd.n3903 gnd.n3902 9.3005
R11323 gnd.n3901 gnd.n1462 9.3005
R11324 gnd.n3900 gnd.n3899 9.3005
R11325 gnd.n3896 gnd.n3895 9.3005
R11326 gnd.n1427 gnd.n1426 9.3005
R11327 gnd.n3941 gnd.n3940 9.3005
R11328 gnd.n3942 gnd.n1425 9.3005
R11329 gnd.n3944 gnd.n3943 9.3005
R11330 gnd.n3946 gnd.n1424 9.3005
R11331 gnd.n3948 gnd.n3947 9.3005
R11332 gnd.n3949 gnd.n1423 9.3005
R11333 gnd.n3956 gnd.n3950 9.3005
R11334 gnd.n3955 gnd.n3951 9.3005
R11335 gnd.n3954 gnd.n3952 9.3005
R11336 gnd.n1388 gnd.n1387 9.3005
R11337 gnd.n3996 gnd.n3995 9.3005
R11338 gnd.n3997 gnd.n1386 9.3005
R11339 gnd.n4008 gnd.n3998 9.3005
R11340 gnd.n4007 gnd.n3999 9.3005
R11341 gnd.n4006 gnd.n4000 9.3005
R11342 gnd.n4005 gnd.n4001 9.3005
R11343 gnd.n4003 gnd.n4002 9.3005
R11344 gnd.n297 gnd.n296 9.3005
R11345 gnd.n6683 gnd.n6682 9.3005
R11346 gnd.n6684 gnd.n295 9.3005
R11347 gnd.n6686 gnd.n6685 9.3005
R11348 gnd.n6747 gnd.n6687 9.3005
R11349 gnd.n6746 gnd.n6688 9.3005
R11350 gnd.n6745 gnd.n6689 9.3005
R11351 gnd.n6744 gnd.n6690 9.3005
R11352 gnd.n6742 gnd.n6691 9.3005
R11353 gnd.n6741 gnd.n6692 9.3005
R11354 gnd.n6739 gnd.n6693 9.3005
R11355 gnd.n6738 gnd.n6694 9.3005
R11356 gnd.n6736 gnd.n6695 9.3005
R11357 gnd.n6735 gnd.n6696 9.3005
R11358 gnd.n6733 gnd.n6697 9.3005
R11359 gnd.n6732 gnd.n6698 9.3005
R11360 gnd.n6730 gnd.n6699 9.3005
R11361 gnd.n6729 gnd.n6700 9.3005
R11362 gnd.n6727 gnd.n6701 9.3005
R11363 gnd.n6726 gnd.n6702 9.3005
R11364 gnd.n6724 gnd.n6703 9.3005
R11365 gnd.n6723 gnd.n6704 9.3005
R11366 gnd.n6721 gnd.n6705 9.3005
R11367 gnd.n6720 gnd.n6706 9.3005
R11368 gnd.n6716 gnd.n6707 9.3005
R11369 gnd.n6715 gnd.n6708 9.3005
R11370 gnd.n6713 gnd.n6709 9.3005
R11371 gnd.n6712 gnd.n6711 9.3005
R11372 gnd.n6710 gnd.n178 9.3005
R11373 gnd.n6937 gnd.n177 9.3005
R11374 gnd.n6939 gnd.n6938 9.3005
R11375 gnd.n3894 gnd.n1461 9.3005
R11376 gnd.n3883 gnd.n1467 9.3005
R11377 gnd.n3885 gnd.n3884 9.3005
R11378 gnd.n3882 gnd.n1469 9.3005
R11379 gnd.n3881 gnd.n3880 9.3005
R11380 gnd.n1471 gnd.n1470 9.3005
R11381 gnd.n3874 gnd.n3873 9.3005
R11382 gnd.n3872 gnd.n1473 9.3005
R11383 gnd.n3871 gnd.n3870 9.3005
R11384 gnd.n1475 gnd.n1474 9.3005
R11385 gnd.n3864 gnd.n3863 9.3005
R11386 gnd.n3862 gnd.n1477 9.3005
R11387 gnd.n3861 gnd.n3860 9.3005
R11388 gnd.n1479 gnd.n1478 9.3005
R11389 gnd.n3854 gnd.n3853 9.3005
R11390 gnd.n3852 gnd.n1481 9.3005
R11391 gnd.n3851 gnd.n3850 9.3005
R11392 gnd.n1483 gnd.n1482 9.3005
R11393 gnd.n3844 gnd.n3843 9.3005
R11394 gnd.n3842 gnd.n1485 9.3005
R11395 gnd.n1487 gnd.n1486 9.3005
R11396 gnd.n3829 gnd.n3784 9.3005
R11397 gnd.n3831 gnd.n3830 9.3005
R11398 gnd.n3828 gnd.n3786 9.3005
R11399 gnd.n3827 gnd.n3826 9.3005
R11400 gnd.n3788 gnd.n3787 9.3005
R11401 gnd.n3820 gnd.n3819 9.3005
R11402 gnd.n3818 gnd.n3790 9.3005
R11403 gnd.n3817 gnd.n3816 9.3005
R11404 gnd.n3792 gnd.n3791 9.3005
R11405 gnd.n3810 gnd.n3809 9.3005
R11406 gnd.n3808 gnd.n3794 9.3005
R11407 gnd.n3807 gnd.n3806 9.3005
R11408 gnd.n3796 gnd.n3795 9.3005
R11409 gnd.n3800 gnd.n3799 9.3005
R11410 gnd.n3798 gnd.n3797 9.3005
R11411 gnd.n1466 gnd.n1463 9.3005
R11412 gnd.n3893 gnd.n3892 9.3005
R11413 gnd.n4056 gnd.n1332 9.3005
R11414 gnd.n4055 gnd.n1333 9.3005
R11415 gnd.n1434 gnd.n1334 9.3005
R11416 gnd.n3933 gnd.n3932 9.3005
R11417 gnd.n3934 gnd.n1433 9.3005
R11418 gnd.n3936 gnd.n3935 9.3005
R11419 gnd.n1405 gnd.n1404 9.3005
R11420 gnd.n3970 gnd.n3969 9.3005
R11421 gnd.n3971 gnd.n1403 9.3005
R11422 gnd.n3975 gnd.n3972 9.3005
R11423 gnd.n3974 gnd.n3973 9.3005
R11424 gnd.n1366 gnd.n1365 9.3005
R11425 gnd.n4023 gnd.n4022 9.3005
R11426 gnd.n4024 gnd.n1364 9.3005
R11427 gnd.n4026 gnd.n4025 9.3005
R11428 gnd.n321 gnd.n320 9.3005
R11429 gnd.n6655 gnd.n6654 9.3005
R11430 gnd.n6656 gnd.n319 9.3005
R11431 gnd.n6660 gnd.n6657 9.3005
R11432 gnd.n6659 gnd.n6658 9.3005
R11433 gnd.n266 gnd.n259 9.3005
R11434 gnd.n247 gnd.n246 9.3005
R11435 gnd.n6790 gnd.n6789 9.3005
R11436 gnd.n6791 gnd.n245 9.3005
R11437 gnd.n6793 gnd.n6792 9.3005
R11438 gnd.n230 gnd.n229 9.3005
R11439 gnd.n6806 gnd.n6805 9.3005
R11440 gnd.n6807 gnd.n228 9.3005
R11441 gnd.n6809 gnd.n6808 9.3005
R11442 gnd.n217 gnd.n216 9.3005
R11443 gnd.n6822 gnd.n6821 9.3005
R11444 gnd.n6823 gnd.n215 9.3005
R11445 gnd.n6825 gnd.n6824 9.3005
R11446 gnd.n201 gnd.n200 9.3005
R11447 gnd.n6838 gnd.n6837 9.3005
R11448 gnd.n6839 gnd.n199 9.3005
R11449 gnd.n6841 gnd.n6840 9.3005
R11450 gnd.n186 gnd.n185 9.3005
R11451 gnd.n6929 gnd.n6928 9.3005
R11452 gnd.n6930 gnd.n184 9.3005
R11453 gnd.n6932 gnd.n6931 9.3005
R11454 gnd.n107 gnd.n106 9.3005
R11455 gnd.n7012 gnd.n7011 9.3005
R11456 gnd.n4057 gnd.n1331 9.3005
R11457 gnd.n6776 gnd.n264 9.3005
R11458 gnd.n6777 gnd.n6776 9.3005
R11459 gnd.n6639 gnd.n6638 9.3005
R11460 gnd.n6637 gnd.n6636 9.3005
R11461 gnd.n2168 gnd.n2158 9.3005
R11462 gnd.n2181 gnd.n2169 9.3005
R11463 gnd.n2180 gnd.n2170 9.3005
R11464 gnd.n2179 gnd.n2171 9.3005
R11465 gnd.n2176 gnd.n2172 9.3005
R11466 gnd.n2175 gnd.n2174 9.3005
R11467 gnd.n2173 gnd.n2138 9.3005
R11468 gnd.n2136 gnd.n2135 9.3005
R11469 gnd.n2479 gnd.n2478 9.3005
R11470 gnd.n2480 gnd.n2134 9.3005
R11471 gnd.n2482 gnd.n2481 9.3005
R11472 gnd.n2132 gnd.n2131 9.3005
R11473 gnd.n2487 gnd.n2486 9.3005
R11474 gnd.n2488 gnd.n2130 9.3005
R11475 gnd.n2516 gnd.n2489 9.3005
R11476 gnd.n2515 gnd.n2490 9.3005
R11477 gnd.n2514 gnd.n2491 9.3005
R11478 gnd.n2494 gnd.n2492 9.3005
R11479 gnd.n2510 gnd.n2495 9.3005
R11480 gnd.n2509 gnd.n2496 9.3005
R11481 gnd.n2508 gnd.n2497 9.3005
R11482 gnd.n2500 gnd.n2498 9.3005
R11483 gnd.n2504 gnd.n2501 9.3005
R11484 gnd.n2503 gnd.n2502 9.3005
R11485 gnd.n1964 gnd.n1963 9.3005
R11486 gnd.n2841 gnd.n2840 9.3005
R11487 gnd.n2842 gnd.n1962 9.3005
R11488 gnd.n2844 gnd.n2843 9.3005
R11489 gnd.n1953 gnd.n1952 9.3005
R11490 gnd.n2861 gnd.n2860 9.3005
R11491 gnd.n2862 gnd.n1951 9.3005
R11492 gnd.n2864 gnd.n2863 9.3005
R11493 gnd.n1940 gnd.n1939 9.3005
R11494 gnd.n2881 gnd.n2880 9.3005
R11495 gnd.n2882 gnd.n1938 9.3005
R11496 gnd.n2884 gnd.n2883 9.3005
R11497 gnd.n1927 gnd.n1926 9.3005
R11498 gnd.n2901 gnd.n2900 9.3005
R11499 gnd.n2902 gnd.n1925 9.3005
R11500 gnd.n2904 gnd.n2903 9.3005
R11501 gnd.n1914 gnd.n1913 9.3005
R11502 gnd.n2921 gnd.n2920 9.3005
R11503 gnd.n2922 gnd.n1912 9.3005
R11504 gnd.n2924 gnd.n2923 9.3005
R11505 gnd.n1899 gnd.n1898 9.3005
R11506 gnd.n2959 gnd.n2958 9.3005
R11507 gnd.n2960 gnd.n1897 9.3005
R11508 gnd.n2962 gnd.n2961 9.3005
R11509 gnd.n1824 gnd.n1823 9.3005
R11510 gnd.n2986 gnd.n2985 9.3005
R11511 gnd.n2987 gnd.n1822 9.3005
R11512 gnd.n2994 gnd.n2988 9.3005
R11513 gnd.n2993 gnd.n2989 9.3005
R11514 gnd.n2992 gnd.n2990 9.3005
R11515 gnd.n1787 gnd.n1786 9.3005
R11516 gnd.n3047 gnd.n3046 9.3005
R11517 gnd.n3048 gnd.n1785 9.3005
R11518 gnd.n3050 gnd.n3049 9.3005
R11519 gnd.n1767 gnd.n1766 9.3005
R11520 gnd.n3114 gnd.n3113 9.3005
R11521 gnd.n3115 gnd.n1765 9.3005
R11522 gnd.n3119 gnd.n3116 9.3005
R11523 gnd.n3118 gnd.n3117 9.3005
R11524 gnd.n1738 gnd.n1737 9.3005
R11525 gnd.n3150 gnd.n3149 9.3005
R11526 gnd.n3151 gnd.n1736 9.3005
R11527 gnd.n3153 gnd.n3152 9.3005
R11528 gnd.n1717 gnd.n1716 9.3005
R11529 gnd.n3178 gnd.n3177 9.3005
R11530 gnd.n3179 gnd.n1715 9.3005
R11531 gnd.n3183 gnd.n3180 9.3005
R11532 gnd.n3182 gnd.n3181 9.3005
R11533 gnd.n1689 gnd.n1688 9.3005
R11534 gnd.n3217 gnd.n3216 9.3005
R11535 gnd.n3218 gnd.n1687 9.3005
R11536 gnd.n3228 gnd.n3219 9.3005
R11537 gnd.n3227 gnd.n3220 9.3005
R11538 gnd.n3226 gnd.n3221 9.3005
R11539 gnd.n1657 gnd.n1656 9.3005
R11540 gnd.n3284 gnd.n3283 9.3005
R11541 gnd.n3285 gnd.n1655 9.3005
R11542 gnd.n3287 gnd.n3286 9.3005
R11543 gnd.n1634 gnd.n1633 9.3005
R11544 gnd.n3313 gnd.n3312 9.3005
R11545 gnd.n3314 gnd.n1632 9.3005
R11546 gnd.n3319 gnd.n3315 9.3005
R11547 gnd.n3318 gnd.n3317 9.3005
R11548 gnd.n3316 gnd.n1539 9.3005
R11549 gnd.n3619 gnd.n1540 9.3005
R11550 gnd.n3618 gnd.n1541 9.3005
R11551 gnd.n3617 gnd.n1542 9.3005
R11552 gnd.n1552 gnd.n1543 9.3005
R11553 gnd.n1553 gnd.n1551 9.3005
R11554 gnd.n3608 gnd.n1554 9.3005
R11555 gnd.n3607 gnd.n1555 9.3005
R11556 gnd.n3606 gnd.n1556 9.3005
R11557 gnd.n1566 gnd.n1557 9.3005
R11558 gnd.n3598 gnd.n1567 9.3005
R11559 gnd.n3597 gnd.n1568 9.3005
R11560 gnd.n3596 gnd.n1569 9.3005
R11561 gnd.n1576 gnd.n1570 9.3005
R11562 gnd.n3588 gnd.n1577 9.3005
R11563 gnd.n3587 gnd.n1578 9.3005
R11564 gnd.n3586 gnd.n1579 9.3005
R11565 gnd.n1589 gnd.n1580 9.3005
R11566 gnd.n3578 gnd.n1590 9.3005
R11567 gnd.n3577 gnd.n1591 9.3005
R11568 gnd.n3576 gnd.n1592 9.3005
R11569 gnd.n1595 gnd.n1594 9.3005
R11570 gnd.n1593 gnd.n1309 9.3005
R11571 gnd.n4072 gnd.n1310 9.3005
R11572 gnd.n4071 gnd.n1311 9.3005
R11573 gnd.n4070 gnd.n1312 9.3005
R11574 gnd.n1318 gnd.n1313 9.3005
R11575 gnd.n4064 gnd.n1319 9.3005
R11576 gnd.n4063 gnd.n1320 9.3005
R11577 gnd.n4062 gnd.n1321 9.3005
R11578 gnd.n1442 gnd.n1322 9.3005
R11579 gnd.n1444 gnd.n1443 9.3005
R11580 gnd.n1448 gnd.n1447 9.3005
R11581 gnd.n1449 gnd.n1441 9.3005
R11582 gnd.n3927 gnd.n1450 9.3005
R11583 gnd.n3926 gnd.n1451 9.3005
R11584 gnd.n3925 gnd.n1453 9.3005
R11585 gnd.n1452 gnd.n1413 9.3005
R11586 gnd.n3964 gnd.n1414 9.3005
R11587 gnd.n3963 gnd.n1415 9.3005
R11588 gnd.n3962 gnd.n1416 9.3005
R11589 gnd.n1419 gnd.n1418 9.3005
R11590 gnd.n1417 gnd.n1374 9.3005
R11591 gnd.n4017 gnd.n1375 9.3005
R11592 gnd.n4016 gnd.n1376 9.3005
R11593 gnd.n4015 gnd.n1377 9.3005
R11594 gnd.n1380 gnd.n1378 9.3005
R11595 gnd.n1385 gnd.n1381 9.3005
R11596 gnd.n1384 gnd.n1383 9.3005
R11597 gnd.n1382 gnd.n336 9.3005
R11598 gnd.n6640 gnd.n337 9.3005
R11599 gnd.n2759 gnd.n2089 9.3005
R11600 gnd.n2762 gnd.n2088 9.3005
R11601 gnd.n2763 gnd.n2087 9.3005
R11602 gnd.n2766 gnd.n2086 9.3005
R11603 gnd.n2767 gnd.n2085 9.3005
R11604 gnd.n2770 gnd.n2084 9.3005
R11605 gnd.n2771 gnd.n2083 9.3005
R11606 gnd.n2774 gnd.n2082 9.3005
R11607 gnd.n2775 gnd.n2081 9.3005
R11608 gnd.n2778 gnd.n2080 9.3005
R11609 gnd.n2779 gnd.n2079 9.3005
R11610 gnd.n2782 gnd.n2078 9.3005
R11611 gnd.n2783 gnd.n2077 9.3005
R11612 gnd.n2784 gnd.n2076 9.3005
R11613 gnd.n2075 gnd.n2072 9.3005
R11614 gnd.n2074 gnd.n2073 9.3005
R11615 gnd.n2626 gnd.n2625 9.3005
R11616 gnd.n2622 gnd.n2094 9.3005
R11617 gnd.n2619 gnd.n2095 9.3005
R11618 gnd.n2618 gnd.n2096 9.3005
R11619 gnd.n2615 gnd.n2097 9.3005
R11620 gnd.n2614 gnd.n2098 9.3005
R11621 gnd.n2611 gnd.n2099 9.3005
R11622 gnd.n2610 gnd.n2100 9.3005
R11623 gnd.n2607 gnd.n2101 9.3005
R11624 gnd.n2606 gnd.n2102 9.3005
R11625 gnd.n2603 gnd.n2103 9.3005
R11626 gnd.n2602 gnd.n2104 9.3005
R11627 gnd.n2599 gnd.n2105 9.3005
R11628 gnd.n2598 gnd.n2106 9.3005
R11629 gnd.n2595 gnd.n2107 9.3005
R11630 gnd.n2594 gnd.n2108 9.3005
R11631 gnd.n2591 gnd.n2109 9.3005
R11632 gnd.n2590 gnd.n2110 9.3005
R11633 gnd.n2587 gnd.n2586 9.3005
R11634 gnd.n2585 gnd.n2112 9.3005
R11635 gnd.n2627 gnd.n2090 9.3005
R11636 gnd.n2272 gnd.n2271 9.3005
R11637 gnd.n2356 gnd.n2355 9.3005
R11638 gnd.n2357 gnd.n2270 9.3005
R11639 gnd.n2360 gnd.n2358 9.3005
R11640 gnd.n2361 gnd.n2269 9.3005
R11641 gnd.n2364 gnd.n2363 9.3005
R11642 gnd.n2365 gnd.n2268 9.3005
R11643 gnd.n2368 gnd.n2366 9.3005
R11644 gnd.n2369 gnd.n2267 9.3005
R11645 gnd.n2372 gnd.n2371 9.3005
R11646 gnd.n2373 gnd.n2266 9.3005
R11647 gnd.n2376 gnd.n2374 9.3005
R11648 gnd.n2377 gnd.n2265 9.3005
R11649 gnd.n2380 gnd.n2379 9.3005
R11650 gnd.n2381 gnd.n2264 9.3005
R11651 gnd.n2384 gnd.n2382 9.3005
R11652 gnd.n2385 gnd.n2263 9.3005
R11653 gnd.n2388 gnd.n2387 9.3005
R11654 gnd.n2389 gnd.n2262 9.3005
R11655 gnd.n2392 gnd.n2390 9.3005
R11656 gnd.n2393 gnd.n2261 9.3005
R11657 gnd.n2396 gnd.n2395 9.3005
R11658 gnd.n2397 gnd.n2260 9.3005
R11659 gnd.n2400 gnd.n2398 9.3005
R11660 gnd.n2401 gnd.n2259 9.3005
R11661 gnd.n2404 gnd.n2403 9.3005
R11662 gnd.n2298 gnd.n2297 9.3005
R11663 gnd.n2303 gnd.n2302 9.3005
R11664 gnd.n2306 gnd.n2292 9.3005
R11665 gnd.n2307 gnd.n2291 9.3005
R11666 gnd.n2310 gnd.n2290 9.3005
R11667 gnd.n2311 gnd.n2289 9.3005
R11668 gnd.n2314 gnd.n2288 9.3005
R11669 gnd.n2315 gnd.n2287 9.3005
R11670 gnd.n2318 gnd.n2286 9.3005
R11671 gnd.n2319 gnd.n2285 9.3005
R11672 gnd.n2322 gnd.n2284 9.3005
R11673 gnd.n2323 gnd.n2283 9.3005
R11674 gnd.n2326 gnd.n2282 9.3005
R11675 gnd.n2327 gnd.n2281 9.3005
R11676 gnd.n2330 gnd.n2280 9.3005
R11677 gnd.n2331 gnd.n2279 9.3005
R11678 gnd.n2334 gnd.n2278 9.3005
R11679 gnd.n2337 gnd.n2336 9.3005
R11680 gnd.n2301 gnd.n2296 9.3005
R11681 gnd.n2300 gnd.n2299 9.3005
R11682 gnd.n2344 gnd.n2343 9.3005
R11683 gnd.n2342 gnd.n2277 9.3005
R11684 gnd.n2341 gnd.n2340 9.3005
R11685 gnd.n2339 gnd.n956 9.3005
R11686 gnd.n4349 gnd.n957 9.3005
R11687 gnd.n4348 gnd.n958 9.3005
R11688 gnd.n4347 gnd.n959 9.3005
R11689 gnd.n975 gnd.n960 9.3005
R11690 gnd.n4337 gnd.n976 9.3005
R11691 gnd.n4336 gnd.n977 9.3005
R11692 gnd.n4335 gnd.n978 9.3005
R11693 gnd.n996 gnd.n979 9.3005
R11694 gnd.n4325 gnd.n997 9.3005
R11695 gnd.n4324 gnd.n998 9.3005
R11696 gnd.n4323 gnd.n999 9.3005
R11697 gnd.n1015 gnd.n1000 9.3005
R11698 gnd.n4313 gnd.n1016 9.3005
R11699 gnd.n4312 gnd.n1017 9.3005
R11700 gnd.n4311 gnd.n1018 9.3005
R11701 gnd.n1036 gnd.n1019 9.3005
R11702 gnd.n4301 gnd.n1037 9.3005
R11703 gnd.n4300 gnd.n1038 9.3005
R11704 gnd.n4299 gnd.n1039 9.3005
R11705 gnd.n1053 gnd.n1040 9.3005
R11706 gnd.n4289 gnd.n1054 9.3005
R11707 gnd.n4288 gnd.n1055 9.3005
R11708 gnd.n4287 gnd.n1056 9.3005
R11709 gnd.n1071 gnd.n1057 9.3005
R11710 gnd.n4276 gnd.n1072 9.3005
R11711 gnd.n4275 gnd.n1073 9.3005
R11712 gnd.n4274 gnd.n1074 9.3005
R11713 gnd.n1090 gnd.n1075 9.3005
R11714 gnd.n4264 gnd.n1091 9.3005
R11715 gnd.n4263 gnd.n1092 9.3005
R11716 gnd.n4262 gnd.n1093 9.3005
R11717 gnd.n1112 gnd.n1094 9.3005
R11718 gnd.n4252 gnd.n1113 9.3005
R11719 gnd.n4251 gnd.n1114 9.3005
R11720 gnd.n4250 gnd.n1115 9.3005
R11721 gnd.n1132 gnd.n1116 9.3005
R11722 gnd.n4240 gnd.n1133 9.3005
R11723 gnd.n4239 gnd.n1134 9.3005
R11724 gnd.n4238 gnd.n1135 9.3005
R11725 gnd.n1154 gnd.n1136 9.3005
R11726 gnd.n4228 gnd.n1155 9.3005
R11727 gnd.n4227 gnd.n1156 9.3005
R11728 gnd.n4226 gnd.n1157 9.3005
R11729 gnd.n1175 gnd.n1158 9.3005
R11730 gnd.n4216 gnd.n1176 9.3005
R11731 gnd.n4215 gnd.n1177 9.3005
R11732 gnd.n4214 gnd.n1178 9.3005
R11733 gnd.n1196 gnd.n1179 9.3005
R11734 gnd.n4204 gnd.n4203 9.3005
R11735 gnd.n2338 gnd.n2276 9.3005
R11736 gnd.n4363 gnd.n4362 9.3005
R11737 gnd.n4361 gnd.n934 9.3005
R11738 gnd.n4360 gnd.n4359 9.3005
R11739 gnd.n936 gnd.n935 9.3005
R11740 gnd.n2203 gnd.n2202 9.3005
R11741 gnd.n2206 gnd.n2205 9.3005
R11742 gnd.n2207 gnd.n2201 9.3005
R11743 gnd.n2210 gnd.n2208 9.3005
R11744 gnd.n2211 gnd.n2200 9.3005
R11745 gnd.n2214 gnd.n2213 9.3005
R11746 gnd.n2215 gnd.n2199 9.3005
R11747 gnd.n2218 gnd.n2216 9.3005
R11748 gnd.n2219 gnd.n2198 9.3005
R11749 gnd.n2222 gnd.n2221 9.3005
R11750 gnd.n2223 gnd.n2197 9.3005
R11751 gnd.n2226 gnd.n2224 9.3005
R11752 gnd.n2227 gnd.n2196 9.3005
R11753 gnd.n2230 gnd.n2229 9.3005
R11754 gnd.n2231 gnd.n2195 9.3005
R11755 gnd.n2234 gnd.n2232 9.3005
R11756 gnd.n2235 gnd.n2194 9.3005
R11757 gnd.n2238 gnd.n2237 9.3005
R11758 gnd.n2239 gnd.n2193 9.3005
R11759 gnd.n2242 gnd.n2240 9.3005
R11760 gnd.n2243 gnd.n2192 9.3005
R11761 gnd.n2246 gnd.n2245 9.3005
R11762 gnd.n2248 gnd.n2190 9.3005
R11763 gnd.n2255 gnd.n2249 9.3005
R11764 gnd.n2254 gnd.n2250 9.3005
R11765 gnd.n2253 gnd.n2251 9.3005
R11766 gnd.n2186 gnd.n2185 9.3005
R11767 gnd.n2420 gnd.n2419 9.3005
R11768 gnd.n2421 gnd.n2184 9.3005
R11769 gnd.n2424 gnd.n2423 9.3005
R11770 gnd.n2422 gnd.n2151 9.3005
R11771 gnd.n2436 gnd.n2152 9.3005
R11772 gnd.n2437 gnd.n2150 9.3005
R11773 gnd.n2439 gnd.n2438 9.3005
R11774 gnd.n2440 gnd.n2149 9.3005
R11775 gnd.n2444 gnd.n2441 9.3005
R11776 gnd.n2445 gnd.n2148 9.3005
R11777 gnd.n2450 gnd.n2449 9.3005
R11778 gnd.n2451 gnd.n2147 9.3005
R11779 gnd.n2457 gnd.n2452 9.3005
R11780 gnd.n2456 gnd.n2453 9.3005
R11781 gnd.n2455 gnd.n2454 9.3005
R11782 gnd.n2123 gnd.n2122 9.3005
R11783 gnd.n2530 gnd.n2529 9.3005
R11784 gnd.n2531 gnd.n2121 9.3005
R11785 gnd.n2534 gnd.n2533 9.3005
R11786 gnd.n2532 gnd.n2116 9.3005
R11787 gnd.n2582 gnd.n2115 9.3005
R11788 gnd.n2584 gnd.n2583 9.3005
R11789 gnd.n4364 gnd.n932 9.3005
R11790 gnd.n4371 gnd.n4370 9.3005
R11791 gnd.n4372 gnd.n926 9.3005
R11792 gnd.n4375 gnd.n925 9.3005
R11793 gnd.n4376 gnd.n924 9.3005
R11794 gnd.n4379 gnd.n923 9.3005
R11795 gnd.n4380 gnd.n922 9.3005
R11796 gnd.n4383 gnd.n921 9.3005
R11797 gnd.n4384 gnd.n920 9.3005
R11798 gnd.n4387 gnd.n919 9.3005
R11799 gnd.n4388 gnd.n918 9.3005
R11800 gnd.n4391 gnd.n917 9.3005
R11801 gnd.n4392 gnd.n916 9.3005
R11802 gnd.n4395 gnd.n915 9.3005
R11803 gnd.n4396 gnd.n914 9.3005
R11804 gnd.n4399 gnd.n913 9.3005
R11805 gnd.n4400 gnd.n912 9.3005
R11806 gnd.n4403 gnd.n911 9.3005
R11807 gnd.n4404 gnd.n910 9.3005
R11808 gnd.n4407 gnd.n909 9.3005
R11809 gnd.n4409 gnd.n906 9.3005
R11810 gnd.n4412 gnd.n905 9.3005
R11811 gnd.n4413 gnd.n904 9.3005
R11812 gnd.n4416 gnd.n903 9.3005
R11813 gnd.n4417 gnd.n902 9.3005
R11814 gnd.n4420 gnd.n901 9.3005
R11815 gnd.n4421 gnd.n900 9.3005
R11816 gnd.n4424 gnd.n899 9.3005
R11817 gnd.n4425 gnd.n898 9.3005
R11818 gnd.n4428 gnd.n897 9.3005
R11819 gnd.n4429 gnd.n896 9.3005
R11820 gnd.n4432 gnd.n895 9.3005
R11821 gnd.n4433 gnd.n894 9.3005
R11822 gnd.n4436 gnd.n893 9.3005
R11823 gnd.n4438 gnd.n892 9.3005
R11824 gnd.n4439 gnd.n891 9.3005
R11825 gnd.n4440 gnd.n890 9.3005
R11826 gnd.n4441 gnd.n889 9.3005
R11827 gnd.n4369 gnd.n931 9.3005
R11828 gnd.n4368 gnd.n4367 9.3005
R11829 gnd.n2350 gnd.n2349 9.3005
R11830 gnd.n2348 gnd.n945 9.3005
R11831 gnd.n4355 gnd.n946 9.3005
R11832 gnd.n4354 gnd.n947 9.3005
R11833 gnd.n4353 gnd.n948 9.3005
R11834 gnd.n966 gnd.n949 9.3005
R11835 gnd.n4343 gnd.n967 9.3005
R11836 gnd.n4342 gnd.n968 9.3005
R11837 gnd.n4341 gnd.n969 9.3005
R11838 gnd.n985 gnd.n970 9.3005
R11839 gnd.n4331 gnd.n986 9.3005
R11840 gnd.n4330 gnd.n987 9.3005
R11841 gnd.n4329 gnd.n988 9.3005
R11842 gnd.n1006 gnd.n989 9.3005
R11843 gnd.n4319 gnd.n1007 9.3005
R11844 gnd.n4318 gnd.n1008 9.3005
R11845 gnd.n4317 gnd.n1009 9.3005
R11846 gnd.n1025 gnd.n1010 9.3005
R11847 gnd.n4307 gnd.n1026 9.3005
R11848 gnd.n4306 gnd.n1027 9.3005
R11849 gnd.n4305 gnd.n1028 9.3005
R11850 gnd.n4269 gnd.n1082 9.3005
R11851 gnd.n4268 gnd.n1083 9.3005
R11852 gnd.n1101 gnd.n1084 9.3005
R11853 gnd.n4258 gnd.n1102 9.3005
R11854 gnd.n4257 gnd.n1103 9.3005
R11855 gnd.n4256 gnd.n1104 9.3005
R11856 gnd.n1122 gnd.n1105 9.3005
R11857 gnd.n4246 gnd.n1123 9.3005
R11858 gnd.n4245 gnd.n1124 9.3005
R11859 gnd.n4244 gnd.n1125 9.3005
R11860 gnd.n1143 gnd.n1126 9.3005
R11861 gnd.n4234 gnd.n1144 9.3005
R11862 gnd.n4233 gnd.n1145 9.3005
R11863 gnd.n4232 gnd.n1146 9.3005
R11864 gnd.n1164 gnd.n1147 9.3005
R11865 gnd.n4222 gnd.n1165 9.3005
R11866 gnd.n4221 gnd.n1166 9.3005
R11867 gnd.n4220 gnd.n1167 9.3005
R11868 gnd.n1186 gnd.n1168 9.3005
R11869 gnd.n4210 gnd.n1187 9.3005
R11870 gnd.n4209 gnd.n1188 9.3005
R11871 gnd.n4208 gnd.n1189 9.3005
R11872 gnd.n2347 gnd.n2346 9.3005
R11873 gnd.n4294 gnd.n1047 9.3005
R11874 gnd.n4270 gnd.n1047 9.3005
R11875 gnd.n2167 gnd.n2166 9.3005
R11876 gnd.n2162 gnd.n2161 9.3005
R11877 gnd.n5898 gnd.n842 9.3005
R11878 gnd.n5899 gnd.n841 9.3005
R11879 gnd.n5900 gnd.n840 9.3005
R11880 gnd.n839 gnd.n835 9.3005
R11881 gnd.n5906 gnd.n834 9.3005
R11882 gnd.n5907 gnd.n833 9.3005
R11883 gnd.n5908 gnd.n832 9.3005
R11884 gnd.n831 gnd.n827 9.3005
R11885 gnd.n5914 gnd.n826 9.3005
R11886 gnd.n5915 gnd.n825 9.3005
R11887 gnd.n5916 gnd.n824 9.3005
R11888 gnd.n823 gnd.n819 9.3005
R11889 gnd.n5922 gnd.n818 9.3005
R11890 gnd.n5923 gnd.n817 9.3005
R11891 gnd.n5924 gnd.n816 9.3005
R11892 gnd.n815 gnd.n811 9.3005
R11893 gnd.n5930 gnd.n810 9.3005
R11894 gnd.n5931 gnd.n809 9.3005
R11895 gnd.n5932 gnd.n808 9.3005
R11896 gnd.n807 gnd.n803 9.3005
R11897 gnd.n5938 gnd.n802 9.3005
R11898 gnd.n5939 gnd.n801 9.3005
R11899 gnd.n5940 gnd.n800 9.3005
R11900 gnd.n799 gnd.n795 9.3005
R11901 gnd.n5946 gnd.n794 9.3005
R11902 gnd.n5947 gnd.n793 9.3005
R11903 gnd.n5948 gnd.n792 9.3005
R11904 gnd.n791 gnd.n787 9.3005
R11905 gnd.n5954 gnd.n786 9.3005
R11906 gnd.n5955 gnd.n785 9.3005
R11907 gnd.n5956 gnd.n784 9.3005
R11908 gnd.n783 gnd.n779 9.3005
R11909 gnd.n5962 gnd.n778 9.3005
R11910 gnd.n5963 gnd.n777 9.3005
R11911 gnd.n5964 gnd.n776 9.3005
R11912 gnd.n775 gnd.n771 9.3005
R11913 gnd.n5970 gnd.n770 9.3005
R11914 gnd.n5971 gnd.n769 9.3005
R11915 gnd.n5972 gnd.n768 9.3005
R11916 gnd.n767 gnd.n763 9.3005
R11917 gnd.n5978 gnd.n762 9.3005
R11918 gnd.n5979 gnd.n761 9.3005
R11919 gnd.n5980 gnd.n760 9.3005
R11920 gnd.n759 gnd.n755 9.3005
R11921 gnd.n5986 gnd.n754 9.3005
R11922 gnd.n5987 gnd.n753 9.3005
R11923 gnd.n5988 gnd.n752 9.3005
R11924 gnd.n751 gnd.n747 9.3005
R11925 gnd.n5994 gnd.n746 9.3005
R11926 gnd.n5995 gnd.n745 9.3005
R11927 gnd.n5996 gnd.n744 9.3005
R11928 gnd.n743 gnd.n739 9.3005
R11929 gnd.n6002 gnd.n738 9.3005
R11930 gnd.n6003 gnd.n737 9.3005
R11931 gnd.n6004 gnd.n736 9.3005
R11932 gnd.n735 gnd.n731 9.3005
R11933 gnd.n6010 gnd.n730 9.3005
R11934 gnd.n6011 gnd.n729 9.3005
R11935 gnd.n6012 gnd.n728 9.3005
R11936 gnd.n727 gnd.n723 9.3005
R11937 gnd.n6018 gnd.n722 9.3005
R11938 gnd.n6019 gnd.n721 9.3005
R11939 gnd.n6020 gnd.n720 9.3005
R11940 gnd.n719 gnd.n715 9.3005
R11941 gnd.n6026 gnd.n714 9.3005
R11942 gnd.n6027 gnd.n713 9.3005
R11943 gnd.n6028 gnd.n712 9.3005
R11944 gnd.n711 gnd.n707 9.3005
R11945 gnd.n6034 gnd.n706 9.3005
R11946 gnd.n6035 gnd.n705 9.3005
R11947 gnd.n6036 gnd.n704 9.3005
R11948 gnd.n703 gnd.n699 9.3005
R11949 gnd.n6042 gnd.n698 9.3005
R11950 gnd.n6043 gnd.n697 9.3005
R11951 gnd.n6044 gnd.n696 9.3005
R11952 gnd.n695 gnd.n691 9.3005
R11953 gnd.n6050 gnd.n690 9.3005
R11954 gnd.n6051 gnd.n689 9.3005
R11955 gnd.n6052 gnd.n688 9.3005
R11956 gnd.n687 gnd.n683 9.3005
R11957 gnd.n6058 gnd.n682 9.3005
R11958 gnd.n6059 gnd.n681 9.3005
R11959 gnd.n6060 gnd.n680 9.3005
R11960 gnd.n679 gnd.n675 9.3005
R11961 gnd.n2159 gnd.n843 9.3005
R11962 gnd.n3459 gnd.n3458 9.3005
R11963 gnd.n3439 gnd.n3437 9.3005
R11964 gnd.n3466 gnd.n3465 9.3005
R11965 gnd.n3433 gnd.n3432 9.3005
R11966 gnd.n3478 gnd.n3477 9.3005
R11967 gnd.n3430 gnd.n3428 9.3005
R11968 gnd.n3485 gnd.n3484 9.3005
R11969 gnd.n3424 gnd.n3423 9.3005
R11970 gnd.n3497 gnd.n3496 9.3005
R11971 gnd.n3421 gnd.n3419 9.3005
R11972 gnd.n3504 gnd.n3503 9.3005
R11973 gnd.n3415 gnd.n3414 9.3005
R11974 gnd.n3516 gnd.n3515 9.3005
R11975 gnd.n3412 gnd.n3410 9.3005
R11976 gnd.n3525 gnd.n3524 9.3005
R11977 gnd.n3523 gnd.n3404 9.3005
R11978 gnd.n3534 gnd.n3403 9.3005
R11979 gnd.n3537 gnd.n3536 9.3005
R11980 gnd.n3442 gnd.n3441 9.3005
R11981 gnd.n3527 gnd.n3526 9.3005
R11982 gnd.n3514 gnd.n3409 9.3005
R11983 gnd.n3513 gnd.n3512 9.3005
R11984 gnd.n3420 gnd.n3416 9.3005
R11985 gnd.n3506 gnd.n3505 9.3005
R11986 gnd.n3495 gnd.n3418 9.3005
R11987 gnd.n3494 gnd.n3493 9.3005
R11988 gnd.n3429 gnd.n3425 9.3005
R11989 gnd.n3487 gnd.n3486 9.3005
R11990 gnd.n3476 gnd.n3427 9.3005
R11991 gnd.n3475 gnd.n3474 9.3005
R11992 gnd.n3438 gnd.n3434 9.3005
R11993 gnd.n3468 gnd.n3467 9.3005
R11994 gnd.n3457 gnd.n3436 9.3005
R11995 gnd.n3456 gnd.n3455 9.3005
R11996 gnd.n3444 gnd.n3443 9.3005
R11997 gnd.n3411 gnd.n3407 9.3005
R11998 gnd.n3533 gnd.n3532 9.3005
R11999 gnd.n3401 gnd.n3400 9.3005
R12000 gnd.n3544 gnd.n3543 9.3005
R12001 gnd.n3545 gnd.n3399 9.3005
R12002 gnd.n3547 gnd.n3546 9.3005
R12003 gnd.n3397 gnd.n3396 9.3005
R12004 gnd.n3557 gnd.n3556 9.3005
R12005 gnd.n3558 gnd.n3395 9.3005
R12006 gnd.n3560 gnd.n3559 9.3005
R12007 gnd.n3393 gnd.n3392 9.3005
R12008 gnd.n3566 gnd.n3565 9.3005
R12009 gnd.n2852 gnd.n1957 9.3005
R12010 gnd.n2854 gnd.n2853 9.3005
R12011 gnd.n1946 gnd.n1945 9.3005
R12012 gnd.n2871 gnd.n2870 9.3005
R12013 gnd.n2872 gnd.n1944 9.3005
R12014 gnd.n2874 gnd.n2873 9.3005
R12015 gnd.n1933 gnd.n1932 9.3005
R12016 gnd.n2891 gnd.n2890 9.3005
R12017 gnd.n2892 gnd.n1931 9.3005
R12018 gnd.n2894 gnd.n2893 9.3005
R12019 gnd.n1920 gnd.n1919 9.3005
R12020 gnd.n2911 gnd.n2910 9.3005
R12021 gnd.n2912 gnd.n1918 9.3005
R12022 gnd.n2914 gnd.n2913 9.3005
R12023 gnd.n1907 gnd.n1906 9.3005
R12024 gnd.n2931 gnd.n2930 9.3005
R12025 gnd.n2932 gnd.n1904 9.3005
R12026 gnd.n2952 gnd.n2951 9.3005
R12027 gnd.n2950 gnd.n1905 9.3005
R12028 gnd.n2949 gnd.n2948 9.3005
R12029 gnd.n2947 gnd.n2933 9.3005
R12030 gnd.n2946 gnd.n2945 9.3005
R12031 gnd.n2944 gnd.n2937 9.3005
R12032 gnd.n2943 gnd.n2942 9.3005
R12033 gnd.n2938 gnd.n1804 9.3005
R12034 gnd.n3013 gnd.n1803 9.3005
R12035 gnd.n3015 gnd.n3014 9.3005
R12036 gnd.n3016 gnd.n1801 9.3005
R12037 gnd.n3024 gnd.n3023 9.3005
R12038 gnd.n3022 gnd.n1802 9.3005
R12039 gnd.n3021 gnd.n3020 9.3005
R12040 gnd.n3019 gnd.n3017 9.3005
R12041 gnd.n1753 gnd.n1752 9.3005
R12042 gnd.n3133 gnd.n3132 9.3005
R12043 gnd.n3134 gnd.n1750 9.3005
R12044 gnd.n3137 gnd.n3136 9.3005
R12045 gnd.n3135 gnd.n1751 9.3005
R12046 gnd.n1724 gnd.n1723 9.3005
R12047 gnd.n3169 gnd.n3168 9.3005
R12048 gnd.n3170 gnd.n1722 9.3005
R12049 gnd.n3172 gnd.n3171 9.3005
R12050 gnd.n1704 gnd.n1703 9.3005
R12051 gnd.n3199 gnd.n3198 9.3005
R12052 gnd.n3200 gnd.n1701 9.3005
R12053 gnd.n3203 gnd.n3202 9.3005
R12054 gnd.n3201 gnd.n1702 9.3005
R12055 gnd.n1673 gnd.n1672 9.3005
R12056 gnd.n3242 gnd.n3241 9.3005
R12057 gnd.n3243 gnd.n1670 9.3005
R12058 gnd.n3249 gnd.n3248 9.3005
R12059 gnd.n3247 gnd.n1671 9.3005
R12060 gnd.n3246 gnd.n3245 9.3005
R12061 gnd.n1642 gnd.n1641 9.3005
R12062 gnd.n3302 gnd.n3301 9.3005
R12063 gnd.n3303 gnd.n1639 9.3005
R12064 gnd.n3306 gnd.n3305 9.3005
R12065 gnd.n3304 gnd.n1640 9.3005
R12066 gnd.n1616 gnd.n1615 9.3005
R12067 gnd.n3345 gnd.n3344 9.3005
R12068 gnd.n3346 gnd.n1614 9.3005
R12069 gnd.n3348 gnd.n3347 9.3005
R12070 gnd.n1612 gnd.n1611 9.3005
R12071 gnd.n3355 gnd.n3354 9.3005
R12072 gnd.n3356 gnd.n1610 9.3005
R12073 gnd.n3358 gnd.n3357 9.3005
R12074 gnd.n3359 gnd.n1609 9.3005
R12075 gnd.n3363 gnd.n3362 9.3005
R12076 gnd.n3364 gnd.n1608 9.3005
R12077 gnd.n3366 gnd.n3365 9.3005
R12078 gnd.n3367 gnd.n1607 9.3005
R12079 gnd.n3374 gnd.n3373 9.3005
R12080 gnd.n3375 gnd.n1606 9.3005
R12081 gnd.n3377 gnd.n3376 9.3005
R12082 gnd.n3378 gnd.n1605 9.3005
R12083 gnd.n3382 gnd.n3381 9.3005
R12084 gnd.n3383 gnd.n1604 9.3005
R12085 gnd.n3385 gnd.n3384 9.3005
R12086 gnd.n3386 gnd.n1603 9.3005
R12087 gnd.n3390 gnd.n3389 9.3005
R12088 gnd.n3391 gnd.n1601 9.3005
R12089 gnd.n3569 gnd.n3568 9.3005
R12090 gnd.n3567 gnd.n1602 9.3005
R12091 gnd.n2851 gnd.n2850 9.3005
R12092 gnd.n2560 gnd.n2559 9.3005
R12093 gnd.n2561 gnd.n2554 9.3005
R12094 gnd.n2563 gnd.n2562 9.3005
R12095 gnd.n2565 gnd.n2564 9.3005
R12096 gnd.n2566 gnd.n2547 9.3005
R12097 gnd.n2568 gnd.n2567 9.3005
R12098 gnd.n2569 gnd.n2546 9.3005
R12099 gnd.n2571 gnd.n2570 9.3005
R12100 gnd.n2572 gnd.n2541 9.3005
R12101 gnd.n2558 gnd.n1958 9.3005
R12102 gnd.n2406 gnd.n2189 9.3005
R12103 gnd.n2408 gnd.n2407 9.3005
R12104 gnd.n2409 gnd.n2188 9.3005
R12105 gnd.n2412 gnd.n2411 9.3005
R12106 gnd.n2413 gnd.n2187 9.3005
R12107 gnd.n2415 gnd.n2414 9.3005
R12108 gnd.n2155 gnd.n2154 9.3005
R12109 gnd.n2429 gnd.n2428 9.3005
R12110 gnd.n2430 gnd.n2153 9.3005
R12111 gnd.n2432 gnd.n2431 9.3005
R12112 gnd.n2142 gnd.n2140 9.3005
R12113 gnd.n2471 gnd.n2470 9.3005
R12114 gnd.n2469 gnd.n2141 9.3005
R12115 gnd.n2468 gnd.n2467 9.3005
R12116 gnd.n2466 gnd.n2143 9.3005
R12117 gnd.n2465 gnd.n2464 9.3005
R12118 gnd.n2463 gnd.n2146 9.3005
R12119 gnd.n2462 gnd.n2461 9.3005
R12120 gnd.n2126 gnd.n2125 9.3005
R12121 gnd.n2522 gnd.n2521 9.3005
R12122 gnd.n2523 gnd.n2124 9.3005
R12123 gnd.n2525 gnd.n2524 9.3005
R12124 gnd.n2120 gnd.n2119 9.3005
R12125 gnd.n2539 gnd.n2538 9.3005
R12126 gnd.n2540 gnd.n2117 9.3005
R12127 gnd.n2578 gnd.n2577 9.3005
R12128 gnd.n2576 gnd.n2118 9.3005
R12129 gnd.n2574 gnd.n2573 9.3005
R12130 gnd.n2033 gnd.n2032 9.3005
R12131 gnd.n2793 gnd.n2792 9.3005
R12132 gnd.n2795 gnd.n2794 9.3005
R12133 gnd.n2021 gnd.n2020 9.3005
R12134 gnd.n2801 gnd.n2800 9.3005
R12135 gnd.n2803 gnd.n2802 9.3005
R12136 gnd.n2013 gnd.n2012 9.3005
R12137 gnd.n2809 gnd.n2808 9.3005
R12138 gnd.n2811 gnd.n2810 9.3005
R12139 gnd.n2003 gnd.n2002 9.3005
R12140 gnd.n2817 gnd.n2816 9.3005
R12141 gnd.n2819 gnd.n2818 9.3005
R12142 gnd.n1995 gnd.n1994 9.3005
R12143 gnd.n2825 gnd.n2824 9.3005
R12144 gnd.n2827 gnd.n2826 9.3005
R12145 gnd.n1985 gnd.n1983 9.3005
R12146 gnd.n2833 gnd.n2832 9.3005
R12147 gnd.n2834 gnd.n1982 9.3005
R12148 gnd.n2036 gnd.n1198 9.3005
R12149 gnd.n1986 gnd.n1984 9.3005
R12150 gnd.n2831 gnd.n2830 9.3005
R12151 gnd.n2829 gnd.n2828 9.3005
R12152 gnd.n1990 gnd.n1989 9.3005
R12153 gnd.n2823 gnd.n2822 9.3005
R12154 gnd.n2821 gnd.n2820 9.3005
R12155 gnd.n1999 gnd.n1998 9.3005
R12156 gnd.n2815 gnd.n2814 9.3005
R12157 gnd.n2813 gnd.n2812 9.3005
R12158 gnd.n2007 gnd.n2006 9.3005
R12159 gnd.n2807 gnd.n2806 9.3005
R12160 gnd.n2805 gnd.n2804 9.3005
R12161 gnd.n2017 gnd.n2016 9.3005
R12162 gnd.n2799 gnd.n2798 9.3005
R12163 gnd.n2797 gnd.n2796 9.3005
R12164 gnd.n2027 gnd.n2026 9.3005
R12165 gnd.n2791 gnd.n2790 9.3005
R12166 gnd.n4198 gnd.n1199 9.3005
R12167 gnd.n4197 gnd.n4196 9.3005
R12168 gnd.n4195 gnd.n1203 9.3005
R12169 gnd.n4194 gnd.n4193 9.3005
R12170 gnd.n4192 gnd.n1204 9.3005
R12171 gnd.n4191 gnd.n4190 9.3005
R12172 gnd.n4189 gnd.n1208 9.3005
R12173 gnd.n4188 gnd.n4187 9.3005
R12174 gnd.n4186 gnd.n1209 9.3005
R12175 gnd.n4185 gnd.n4184 9.3005
R12176 gnd.n4183 gnd.n1213 9.3005
R12177 gnd.n4182 gnd.n4181 9.3005
R12178 gnd.n4180 gnd.n1214 9.3005
R12179 gnd.n4179 gnd.n4178 9.3005
R12180 gnd.n4177 gnd.n1218 9.3005
R12181 gnd.n4176 gnd.n4175 9.3005
R12182 gnd.n4174 gnd.n1219 9.3005
R12183 gnd.n4173 gnd.n4172 9.3005
R12184 gnd.n4171 gnd.n1223 9.3005
R12185 gnd.n4170 gnd.n4169 9.3005
R12186 gnd.n4168 gnd.n1224 9.3005
R12187 gnd.n4167 gnd.n4166 9.3005
R12188 gnd.n4165 gnd.n1228 9.3005
R12189 gnd.n4164 gnd.n4163 9.3005
R12190 gnd.n4162 gnd.n1229 9.3005
R12191 gnd.n4161 gnd.n4160 9.3005
R12192 gnd.n4159 gnd.n1233 9.3005
R12193 gnd.n4158 gnd.n4157 9.3005
R12194 gnd.n4156 gnd.n1234 9.3005
R12195 gnd.n4155 gnd.n4154 9.3005
R12196 gnd.n4153 gnd.n1238 9.3005
R12197 gnd.n4152 gnd.n4151 9.3005
R12198 gnd.n4150 gnd.n1239 9.3005
R12199 gnd.n4149 gnd.n4148 9.3005
R12200 gnd.n4147 gnd.n1243 9.3005
R12201 gnd.n4146 gnd.n4145 9.3005
R12202 gnd.n4144 gnd.n1244 9.3005
R12203 gnd.n4143 gnd.n4142 9.3005
R12204 gnd.n4141 gnd.n1248 9.3005
R12205 gnd.n4140 gnd.n4139 9.3005
R12206 gnd.n4138 gnd.n1249 9.3005
R12207 gnd.n4137 gnd.n4136 9.3005
R12208 gnd.n4135 gnd.n1253 9.3005
R12209 gnd.n4134 gnd.n4133 9.3005
R12210 gnd.n4132 gnd.n1254 9.3005
R12211 gnd.n4131 gnd.n4130 9.3005
R12212 gnd.n4129 gnd.n1258 9.3005
R12213 gnd.n4128 gnd.n4127 9.3005
R12214 gnd.n4126 gnd.n1259 9.3005
R12215 gnd.n4125 gnd.n4124 9.3005
R12216 gnd.n4123 gnd.n1263 9.3005
R12217 gnd.n4122 gnd.n4121 9.3005
R12218 gnd.n4120 gnd.n1264 9.3005
R12219 gnd.n4119 gnd.n4118 9.3005
R12220 gnd.n4117 gnd.n1268 9.3005
R12221 gnd.n4116 gnd.n4115 9.3005
R12222 gnd.n4114 gnd.n1269 9.3005
R12223 gnd.n4113 gnd.n4112 9.3005
R12224 gnd.n4111 gnd.n1273 9.3005
R12225 gnd.n4110 gnd.n4109 9.3005
R12226 gnd.n4108 gnd.n1274 9.3005
R12227 gnd.n4107 gnd.n4106 9.3005
R12228 gnd.n4105 gnd.n1278 9.3005
R12229 gnd.n4104 gnd.n4103 9.3005
R12230 gnd.n4102 gnd.n1279 9.3005
R12231 gnd.n4101 gnd.n4100 9.3005
R12232 gnd.n4099 gnd.n1283 9.3005
R12233 gnd.n4098 gnd.n4097 9.3005
R12234 gnd.n4096 gnd.n1284 9.3005
R12235 gnd.n4095 gnd.n4094 9.3005
R12236 gnd.n4093 gnd.n1288 9.3005
R12237 gnd.n4092 gnd.n4091 9.3005
R12238 gnd.n4090 gnd.n1289 9.3005
R12239 gnd.n4089 gnd.n4088 9.3005
R12240 gnd.n4087 gnd.n1293 9.3005
R12241 gnd.n4086 gnd.n4085 9.3005
R12242 gnd.n4084 gnd.n1294 9.3005
R12243 gnd.n4083 gnd.n4082 9.3005
R12244 gnd.n4081 gnd.n1298 9.3005
R12245 gnd.n4080 gnd.n4079 9.3005
R12246 gnd.n4078 gnd.n1299 9.3005
R12247 gnd.n4077 gnd.n1302 9.3005
R12248 gnd.n4200 gnd.n4199 9.3005
R12249 gnd.n1344 gnd.n1342 9.3005
R12250 gnd.n4051 gnd.n4050 9.3005
R12251 gnd.n4049 gnd.n1343 9.3005
R12252 gnd.n4048 gnd.n4047 9.3005
R12253 gnd.n4046 gnd.n1345 9.3005
R12254 gnd.n4045 gnd.n4044 9.3005
R12255 gnd.n4043 gnd.n1349 9.3005
R12256 gnd.n4042 gnd.n4041 9.3005
R12257 gnd.n4040 gnd.n1350 9.3005
R12258 gnd.n4039 gnd.n4038 9.3005
R12259 gnd.n4037 gnd.n1354 9.3005
R12260 gnd.n4036 gnd.n4035 9.3005
R12261 gnd.n4034 gnd.n1355 9.3005
R12262 gnd.n4033 gnd.n4032 9.3005
R12263 gnd.n4031 gnd.n4030 9.3005
R12264 gnd.n330 gnd.n328 9.3005
R12265 gnd.n6650 gnd.n6649 9.3005
R12266 gnd.n6648 gnd.n329 9.3005
R12267 gnd.n6647 gnd.n6646 9.3005
R12268 gnd.n6645 gnd.n331 9.3005
R12269 gnd.n276 gnd.n274 9.3005
R12270 gnd.n6770 gnd.n6769 9.3005
R12271 gnd.n6768 gnd.n275 9.3005
R12272 gnd.n6767 gnd.n6766 9.3005
R12273 gnd.n6765 gnd.n277 9.3005
R12274 gnd.n6764 gnd.n6763 9.3005
R12275 gnd.n6761 gnd.n281 9.3005
R12276 gnd.n6760 gnd.n6759 9.3005
R12277 gnd.n6758 gnd.n283 9.3005
R12278 gnd.n254 gnd.n253 9.3005
R12279 gnd.n6782 gnd.n6781 9.3005
R12280 gnd.n6783 gnd.n252 9.3005
R12281 gnd.n6785 gnd.n6784 9.3005
R12282 gnd.n239 gnd.n238 9.3005
R12283 gnd.n6798 gnd.n6797 9.3005
R12284 gnd.n6799 gnd.n237 9.3005
R12285 gnd.n6801 gnd.n6800 9.3005
R12286 gnd.n224 gnd.n223 9.3005
R12287 gnd.n6814 gnd.n6813 9.3005
R12288 gnd.n6815 gnd.n222 9.3005
R12289 gnd.n6817 gnd.n6816 9.3005
R12290 gnd.n209 gnd.n208 9.3005
R12291 gnd.n6830 gnd.n6829 9.3005
R12292 gnd.n6831 gnd.n207 9.3005
R12293 gnd.n6833 gnd.n6832 9.3005
R12294 gnd.n195 gnd.n194 9.3005
R12295 gnd.n6846 gnd.n6845 9.3005
R12296 gnd.n6847 gnd.n192 9.3005
R12297 gnd.n6924 gnd.n6923 9.3005
R12298 gnd.n6922 gnd.n193 9.3005
R12299 gnd.n6921 gnd.n6920 9.3005
R12300 gnd.n6919 gnd.n6848 9.3005
R12301 gnd.n6918 gnd.n6917 9.3005
R12302 gnd.n3447 gnd.n3446 9.3005
R12303 gnd.n6914 gnd.n6850 9.3005
R12304 gnd.n6913 gnd.n6912 9.3005
R12305 gnd.n6911 gnd.n6855 9.3005
R12306 gnd.n6910 gnd.n6909 9.3005
R12307 gnd.n6908 gnd.n6856 9.3005
R12308 gnd.n6907 gnd.n6906 9.3005
R12309 gnd.n6905 gnd.n6863 9.3005
R12310 gnd.n6904 gnd.n6903 9.3005
R12311 gnd.n6902 gnd.n6864 9.3005
R12312 gnd.n6901 gnd.n6900 9.3005
R12313 gnd.n6899 gnd.n6871 9.3005
R12314 gnd.n6898 gnd.n6897 9.3005
R12315 gnd.n6896 gnd.n6872 9.3005
R12316 gnd.n6895 gnd.n6894 9.3005
R12317 gnd.n6893 gnd.n6879 9.3005
R12318 gnd.n6892 gnd.n6891 9.3005
R12319 gnd.n6890 gnd.n6880 9.3005
R12320 gnd.n6889 gnd.n6888 9.3005
R12321 gnd.n6916 gnd.n6915 9.3005
R12322 gnd.n3908 gnd.n3907 9.3005
R12323 gnd.n3909 gnd.n1457 9.3005
R12324 gnd.n3911 gnd.n3910 9.3005
R12325 gnd.n3912 gnd.n1456 9.3005
R12326 gnd.n3915 gnd.n3914 9.3005
R12327 gnd.n3916 gnd.n1454 9.3005
R12328 gnd.n3919 gnd.n3918 9.3005
R12329 gnd.n3917 gnd.n1455 9.3005
R12330 gnd.n1395 gnd.n1394 9.3005
R12331 gnd.n3980 gnd.n3979 9.3005
R12332 gnd.n3981 gnd.n1392 9.3005
R12333 gnd.n3983 gnd.n3982 9.3005
R12334 gnd.n3984 gnd.n1391 9.3005
R12335 gnd.n3987 gnd.n3986 9.3005
R12336 gnd.n3988 gnd.n1389 9.3005
R12337 gnd.n3991 gnd.n3990 9.3005
R12338 gnd.n3989 gnd.n1390 9.3005
R12339 gnd.n310 gnd.n309 9.3005
R12340 gnd.n6665 gnd.n6664 9.3005
R12341 gnd.n6666 gnd.n307 9.3005
R12342 gnd.n6668 gnd.n6667 9.3005
R12343 gnd.n6669 gnd.n306 9.3005
R12344 gnd.n6672 gnd.n6671 9.3005
R12345 gnd.n6673 gnd.n305 9.3005
R12346 gnd.n6675 gnd.n6674 9.3005
R12347 gnd.n65 gnd.n63 9.3005
R12348 gnd.n7055 gnd.n7054 9.3005
R12349 gnd.n7053 gnd.n64 9.3005
R12350 gnd.n7052 gnd.n7051 9.3005
R12351 gnd.n7050 gnd.n69 9.3005
R12352 gnd.n7049 gnd.n7048 9.3005
R12353 gnd.n7047 gnd.n70 9.3005
R12354 gnd.n7046 gnd.n7045 9.3005
R12355 gnd.n7044 gnd.n74 9.3005
R12356 gnd.n7043 gnd.n7042 9.3005
R12357 gnd.n7041 gnd.n75 9.3005
R12358 gnd.n7040 gnd.n7039 9.3005
R12359 gnd.n7038 gnd.n79 9.3005
R12360 gnd.n7037 gnd.n7036 9.3005
R12361 gnd.n7035 gnd.n80 9.3005
R12362 gnd.n7034 gnd.n7033 9.3005
R12363 gnd.n7032 gnd.n84 9.3005
R12364 gnd.n7031 gnd.n7030 9.3005
R12365 gnd.n7029 gnd.n85 9.3005
R12366 gnd.n7028 gnd.n7027 9.3005
R12367 gnd.n7026 gnd.n89 9.3005
R12368 gnd.n7025 gnd.n7024 9.3005
R12369 gnd.n7023 gnd.n90 9.3005
R12370 gnd.n7022 gnd.n7021 9.3005
R12371 gnd.n7020 gnd.n94 9.3005
R12372 gnd.n7019 gnd.n7018 9.3005
R12373 gnd.n7017 gnd.n95 9.3005
R12374 gnd.n7016 gnd.n98 9.3005
R12375 gnd.n1460 gnd.n1459 9.3005
R12376 gnd.t295 gnd.n4901 9.24152
R12377 gnd.n5783 gnd.t124 9.24152
R12378 gnd.t110 gnd.n846 9.24152
R12379 gnd.t81 gnd.n939 9.24152
R12380 gnd.n2518 gnd.t159 9.24152
R12381 gnd.t20 gnd.n1529 9.24152
R12382 gnd.n3923 gnd.t231 9.24152
R12383 gnd.n6934 gnd.t52 9.24152
R12384 gnd.t305 gnd.t295 8.92286
R12385 gnd.n1836 gnd.n1826 8.92286
R12386 gnd.t101 gnd.n1812 8.92286
R12387 gnd.n1781 gnd.t36 8.92286
R12388 gnd.n3109 gnd.t154 8.92286
R12389 gnd.n3156 gnd.n1733 8.92286
R12390 gnd.n3077 gnd.n1697 8.92286
R12391 gnd.n3252 gnd.t288 8.92286
R12392 gnd.n3281 gnd.t151 8.92286
R12393 gnd.n1647 gnd.n1636 8.92286
R12394 gnd.n3349 gnd.n1536 8.92286
R12395 gnd.n6718 gnd.n205 8.92286
R12396 gnd.n4786 gnd.n4761 8.92171
R12397 gnd.n4754 gnd.n4729 8.92171
R12398 gnd.n4722 gnd.n4697 8.92171
R12399 gnd.n4691 gnd.n4666 8.92171
R12400 gnd.n4659 gnd.n4634 8.92171
R12401 gnd.n4627 gnd.n4602 8.92171
R12402 gnd.n4595 gnd.n4570 8.92171
R12403 gnd.n4564 gnd.n4539 8.92171
R12404 gnd.n3644 gnd.n3626 8.72777
R12405 gnd.t297 gnd.n4943 8.60421
R12406 gnd.t8 gnd.n1726 8.60421
R12407 gnd.n3194 gnd.t149 8.60421
R12408 gnd.n5323 gnd.n5307 8.43467
R12409 gnd.n46 gnd.n30 8.43467
R12410 gnd.n2405 gnd.n0 8.41456
R12411 gnd.n7057 gnd.n7056 8.41456
R12412 gnd.n3027 gnd.n1791 8.28555
R12413 gnd.n3147 gnd.n1740 8.28555
R12414 gnd.n3214 gnd.n3213 8.28555
R12415 gnd.n3290 gnd.n3289 8.28555
R12416 gnd.n4787 gnd.n4759 8.14595
R12417 gnd.n4755 gnd.n4727 8.14595
R12418 gnd.n4723 gnd.n4695 8.14595
R12419 gnd.n4692 gnd.n4664 8.14595
R12420 gnd.n4660 gnd.n4632 8.14595
R12421 gnd.n4628 gnd.n4600 8.14595
R12422 gnd.n4596 gnd.n4568 8.14595
R12423 gnd.n4565 gnd.n4537 8.14595
R12424 gnd.n4792 gnd.n4791 7.97301
R12425 gnd.n5537 gnd.t298 7.9669
R12426 gnd.n5895 gnd.t124 7.9669
R12427 gnd.n6890 gnd.n6889 7.75808
R12428 gnd.n3532 gnd.n3407 7.75808
R12429 gnd.n2790 gnd.n2026 7.75808
R12430 gnd.n2299 gnd.n2296 7.75808
R12431 gnd.n5895 gnd.n5894 7.64824
R12432 gnd.n3027 gnd.n3026 7.64824
R12433 gnd.t25 gnd.n3139 7.64824
R12434 gnd.n3139 gnd.n1740 7.64824
R12435 gnd.n3213 gnd.n1693 7.64824
R12436 gnd.t26 gnd.n1693 7.64824
R12437 gnd.n3290 gnd.n1652 7.64824
R12438 gnd.t303 gnd.n5486 7.32958
R12439 gnd.n1857 gnd.n1856 7.30353
R12440 gnd.n3643 gnd.n3642 7.30353
R12441 gnd.n5445 gnd.n5444 7.01093
R12442 gnd.n5456 gnd.n5053 7.01093
R12443 gnd.n5455 gnd.n5056 7.01093
R12444 gnd.n5466 gnd.n5046 7.01093
R12445 gnd.n5364 gnd.n5039 7.01093
R12446 gnd.n5476 gnd.n5475 7.01093
R12447 gnd.n5487 gnd.n5028 7.01093
R12448 gnd.n5486 gnd.n5031 7.01093
R12449 gnd.n5497 gnd.n5019 7.01093
R12450 gnd.n5022 gnd.n5020 7.01093
R12451 gnd.n5507 gnd.n5506 7.01093
R12452 gnd.n5518 gnd.n5002 7.01093
R12453 gnd.n5528 gnd.n4993 7.01093
R12454 gnd.n4996 gnd.n4994 7.01093
R12455 gnd.n5538 gnd.n5537 7.01093
R12456 gnd.n5549 gnd.n4976 7.01093
R12457 gnd.n5559 gnd.n4968 7.01093
R12458 gnd.n4969 gnd.n4961 7.01093
R12459 gnd.n5580 gnd.n4950 7.01093
R12460 gnd.n5579 gnd.n4953 7.01093
R12461 gnd.n5590 gnd.n4943 7.01093
R12462 gnd.n5280 gnd.n4936 7.01093
R12463 gnd.n5600 gnd.n5599 7.01093
R12464 gnd.n5611 gnd.n4925 7.01093
R12465 gnd.n5610 gnd.n4928 7.01093
R12466 gnd.n4918 gnd.n4911 7.01093
R12467 gnd.n5631 gnd.n5630 7.01093
R12468 gnd.n5641 gnd.n4901 7.01093
R12469 gnd.n5640 gnd.n4904 7.01093
R12470 gnd.n5651 gnd.n4894 7.01093
R12471 gnd.n5661 gnd.n4887 7.01093
R12472 gnd.n5672 gnd.n4881 7.01093
R12473 gnd.n5695 gnd.n4862 7.01093
R12474 gnd.n5705 gnd.n4853 7.01093
R12475 gnd.n4852 gnd.n4845 7.01093
R12476 gnd.n5716 gnd.n5715 7.01093
R12477 gnd.n5729 gnd.n4839 7.01093
R12478 gnd.n5728 gnd.n5727 7.01093
R12479 gnd.n4832 gnd.n4818 7.01093
R12480 gnd.n5761 gnd.n5760 7.01093
R12481 gnd.n5772 gnd.n4812 7.01093
R12482 gnd.n5771 gnd.n4533 7.01093
R12483 gnd.n5791 gnd.n4534 7.01093
R12484 gnd.n5783 gnd.n4805 7.01093
R12485 gnd.n5894 gnd.n846 7.01093
R12486 gnd.n5798 gnd.n854 7.01093
R12487 gnd.n5888 gnd.n5887 7.01093
R12488 gnd.n2983 gnd.n1826 7.01093
R12489 gnd.n3036 gnd.n1795 7.01093
R12490 gnd.n3036 gnd.t137 7.01093
R12491 gnd.n3156 gnd.n3155 7.01093
R12492 gnd.n3077 gnd.n3076 7.01093
R12493 gnd.n3310 gnd.n1636 7.01093
R12494 gnd.n3621 gnd.n1536 7.01093
R12495 gnd.n3712 gnd.t131 7.01093
R12496 gnd.n5022 gnd.t290 6.69227
R12497 gnd.n5631 gnd.t305 6.69227
R12498 gnd.n5741 gnd.t296 6.69227
R12499 gnd.n4339 gnd.t227 6.69227
R12500 gnd.n2459 gnd.t178 6.69227
R12501 gnd.n1895 gnd.t2 6.69227
R12502 gnd.n3351 gnd.t20 6.69227
R12503 gnd.n1410 gnd.t188 6.69227
R12504 gnd.t192 gnd.n203 6.69227
R12505 gnd.n3773 gnd.n3772 6.5566
R12506 gnd.n2688 gnd.n2687 6.5566
R12507 gnd.n2749 gnd.n2695 6.5566
R12508 gnd.n3651 gnd.n3650 6.5566
R12509 gnd.t134 gnd.n1835 6.37362
R12510 gnd.n3060 gnd.n1775 6.37362
R12511 gnd.n3140 gnd.t25 6.37362
R12512 gnd.n3069 gnd.t26 6.37362
R12513 gnd.n3273 gnd.n3271 6.37362
R12514 gnd.n3308 gnd.t104 6.37362
R12515 gnd.n2562 gnd.n2553 6.20656
R12516 gnd.n6979 gnd.n6976 6.20656
R12517 gnd.n4408 gnd.n4407 6.20656
R12518 gnd.n3555 gnd.n3395 6.20656
R12519 gnd.n5548 gnd.t309 6.05496
R12520 gnd.n4979 gnd.t289 6.05496
R12521 gnd.n5280 gnd.t313 6.05496
R12522 gnd.n5682 gnd.t300 6.05496
R12523 gnd.n4315 gnd.t169 6.05496
R12524 gnd.n2434 gnd.t190 6.05496
R12525 gnd.n2965 gnd.n2964 6.05496
R12526 gnd.n3155 gnd.t8 6.05496
R12527 gnd.n3076 gnd.t149 6.05496
R12528 gnd.n3779 gnd.n1492 6.05496
R12529 gnd.n6652 gnd.t214 6.05496
R12530 gnd.t253 gnd.n232 6.05496
R12531 gnd.n4789 gnd.n4759 5.81868
R12532 gnd.n4757 gnd.n4727 5.81868
R12533 gnd.n4725 gnd.n4695 5.81868
R12534 gnd.n4694 gnd.n4664 5.81868
R12535 gnd.n4662 gnd.n4632 5.81868
R12536 gnd.n4630 gnd.n4600 5.81868
R12537 gnd.n4598 gnd.n4568 5.81868
R12538 gnd.n4567 gnd.n4537 5.81868
R12539 gnd.n2997 gnd.n2996 5.73631
R12540 gnd.n3004 gnd.n1810 5.73631
R12541 gnd.n3175 gnd.n1719 5.73631
R12542 gnd.n3188 gnd.n1710 5.73631
R12543 gnd.n3322 gnd.n3321 5.73631
R12544 gnd.n1630 gnd.n1618 5.73631
R12545 gnd.n3349 gnd.t131 5.73631
R12546 gnd.n3782 gnd.n1488 5.62001
R12547 gnd.n2757 gnd.n2692 5.62001
R12548 gnd.n2757 gnd.n2753 5.62001
R12549 gnd.n3782 gnd.n1489 5.62001
R12550 gnd.n5150 gnd.n5149 5.4308
R12551 gnd.n4522 gnd.n4520 5.4308
R12552 gnd.n5600 gnd.t299 5.41765
R12553 gnd.n5621 gnd.t301 5.41765
R12554 gnd.t18 gnd.n4871 5.41765
R12555 gnd.n4291 gnd.t161 5.41765
R12556 gnd.n2257 gnd.t202 5.41765
R12557 gnd.n1812 gnd.t27 5.41765
R12558 gnd.n3323 gnd.t0 5.41765
R12559 gnd.n6677 gnd.t234 5.41765
R12560 gnd.t240 gnd.n285 5.41765
R12561 gnd.n2163 gnd.n1069 5.09899
R12562 gnd.n4272 gnd.n1079 5.09899
R12563 gnd.n2417 gnd.n1086 5.09899
R12564 gnd.n2426 gnd.n1096 5.09899
R12565 gnd.n4260 gnd.n1099 5.09899
R12566 gnd.n2434 gnd.n1107 5.09899
R12567 gnd.n4254 gnd.n1110 5.09899
R12568 gnd.n2474 gnd.n2473 5.09899
R12569 gnd.n4248 gnd.n1120 5.09899
R12570 gnd.n2442 gnd.n1128 5.09899
R12571 gnd.n2447 gnd.n1138 5.09899
R12572 gnd.n4236 gnd.n1141 5.09899
R12573 gnd.n2459 gnd.n1149 5.09899
R12574 gnd.n4230 gnd.n1152 5.09899
R12575 gnd.n2519 gnd.n2518 5.09899
R12576 gnd.n4224 gnd.n1162 5.09899
R12577 gnd.n2527 gnd.n1170 5.09899
R12578 gnd.n4218 gnd.n1173 5.09899
R12579 gnd.n2536 gnd.n1181 5.09899
R12580 gnd.n4212 gnd.n1184 5.09899
R12581 gnd.n2580 gnd.n1191 5.09899
R12582 gnd.n4206 gnd.n1194 5.09899
R12583 gnd.n3110 gnd.n3109 5.09899
R12584 gnd.n3123 gnd.n3122 5.09899
R12585 gnd.n3223 gnd.n3222 5.09899
R12586 gnd.n3252 gnd.n3251 5.09899
R12587 gnd.n1546 gnd.t89 5.09899
R12588 gnd.n4060 gnd.n4059 5.09899
R12589 gnd.n3905 gnd.n1327 5.09899
R12590 gnd.n4053 gnd.n1336 5.09899
R12591 gnd.n3897 gnd.n1339 5.09899
R12592 gnd.n3930 gnd.n1435 5.09899
R12593 gnd.n3929 gnd.n1438 5.09899
R12594 gnd.n3938 gnd.n1430 5.09899
R12595 gnd.n3923 gnd.n3922 5.09899
R12596 gnd.n3967 gnd.n1407 5.09899
R12597 gnd.n3966 gnd.n1410 5.09899
R12598 gnd.n3977 gnd.n1398 5.09899
R12599 gnd.n1421 gnd.n1400 5.09899
R12600 gnd.n4020 gnd.n1368 5.09899
R12601 gnd.n4019 gnd.n1371 5.09899
R12602 gnd.n4028 gnd.n1359 5.09899
R12603 gnd.n3993 gnd.n1362 5.09899
R12604 gnd.n6652 gnd.n323 5.09899
R12605 gnd.n4011 gnd.n4010 5.09899
R12606 gnd.n6662 gnd.n313 5.09899
R12607 gnd.n6642 gnd.n333 5.09899
R12608 gnd.n6772 gnd.n269 5.09899
R12609 gnd.n6634 gnd.n300 5.09899
R12610 gnd.n4787 gnd.n4786 5.04292
R12611 gnd.n4755 gnd.n4754 5.04292
R12612 gnd.n4723 gnd.n4722 5.04292
R12613 gnd.n4692 gnd.n4691 5.04292
R12614 gnd.n4660 gnd.n4659 5.04292
R12615 gnd.n4628 gnd.n4627 5.04292
R12616 gnd.n4596 gnd.n4595 5.04292
R12617 gnd.n4565 gnd.n4564 5.04292
R12618 gnd.n5339 gnd.n5338 4.82753
R12619 gnd.n62 gnd.n61 4.82753
R12620 gnd.n5569 gnd.t304 4.78034
R12621 gnd.n5651 gnd.t293 4.78034
R12622 gnd.n1031 gnd.t167 4.78034
R12623 gnd.n4266 gnd.t163 4.78034
R12624 gnd.t145 gnd.n2876 4.78034
R12625 gnd.n3004 gnd.t27 4.78034
R12626 gnd.t0 gnd.n3322 4.78034
R12627 gnd.n3779 gnd.t89 4.78034
R12628 gnd.n3584 gnd.t10 4.78034
R12629 gnd.n6643 gnd.t196 4.78034
R12630 gnd.n6787 gnd.t246 4.78034
R12631 gnd.n5343 gnd.n5342 4.74817
R12632 gnd.n5292 gnd.n5288 4.74817
R12633 gnd.n5285 gnd.n5284 4.74817
R12634 gnd.n5279 gnd.n5258 4.74817
R12635 gnd.n5342 gnd.n5256 4.74817
R12636 gnd.n5292 gnd.n5291 4.74817
R12637 gnd.n5287 gnd.n5285 4.74817
R12638 gnd.n5283 gnd.n5258 4.74817
R12639 gnd.n6775 gnd.n6774 4.74817
R12640 gnd.n290 gnd.n263 4.74817
R12641 gnd.n6753 gnd.n262 4.74817
R12642 gnd.n261 gnd.n258 4.74817
R12643 gnd.n6775 gnd.n265 4.74817
R12644 gnd.n303 gnd.n263 4.74817
R12645 gnd.n291 gnd.n262 4.74817
R12646 gnd.n6754 gnd.n261 4.74817
R12647 gnd.n1046 gnd.n1029 4.74817
R12648 gnd.n1063 gnd.n1048 4.74817
R12649 gnd.n4282 gnd.n4281 4.74817
R12650 gnd.n1081 gnd.n1064 4.74817
R12651 gnd.n4295 gnd.n1046 4.74817
R12652 gnd.n4293 gnd.n1048 4.74817
R12653 gnd.n4283 gnd.n4282 4.74817
R12654 gnd.n4280 gnd.n1064 4.74817
R12655 gnd.n5323 gnd.n5322 4.7074
R12656 gnd.n46 gnd.n45 4.7074
R12657 gnd.n5339 gnd.n5323 4.65959
R12658 gnd.n62 gnd.n46 4.65959
R12659 gnd.n3841 gnd.n3840 4.6132
R12660 gnd.n2758 gnd.n2628 4.6132
R12661 gnd.n1831 gnd.n1830 4.46168
R12662 gnd.n1813 gnd.n1806 4.46168
R12663 gnd.n3164 gnd.n3163 4.46168
R12664 gnd.n3186 gnd.n3185 4.46168
R12665 gnd.n3324 gnd.n1626 4.46168
R12666 gnd.n3331 gnd.t39 4.46168
R12667 gnd.n3340 gnd.n3339 4.46168
R12668 gnd.n3639 gnd.n3626 4.46111
R12669 gnd.n4772 gnd.n4768 4.38594
R12670 gnd.n4740 gnd.n4736 4.38594
R12671 gnd.n4708 gnd.n4704 4.38594
R12672 gnd.n4677 gnd.n4673 4.38594
R12673 gnd.n4645 gnd.n4641 4.38594
R12674 gnd.n4613 gnd.n4609 4.38594
R12675 gnd.n4581 gnd.n4577 4.38594
R12676 gnd.n4550 gnd.n4546 4.38594
R12677 gnd.n4783 gnd.n4761 4.26717
R12678 gnd.n4751 gnd.n4729 4.26717
R12679 gnd.n4719 gnd.n4697 4.26717
R12680 gnd.n4688 gnd.n4666 4.26717
R12681 gnd.n4656 gnd.n4634 4.26717
R12682 gnd.n4624 gnd.n4602 4.26717
R12683 gnd.n4592 gnd.n4570 4.26717
R12684 gnd.n4561 gnd.n4539 4.26717
R12685 gnd.t294 gnd.n5005 4.14303
R12686 gnd.n5715 gnd.t291 4.14303
R12687 gnd.n991 gnd.t171 4.14303
R12688 gnd.n4242 gnd.t176 4.14303
R12689 gnd.t63 gnd.n1184 4.14303
R12690 gnd.t56 gnd.n1336 4.14303
R12691 gnd.t249 gnd.n3958 4.14303
R12692 gnd.n6819 gnd.t204 4.14303
R12693 gnd.n4791 gnd.n4790 4.08274
R12694 gnd.n3772 gnd.n3771 4.05904
R12695 gnd.n2687 gnd.n2686 4.05904
R12696 gnd.n2746 gnd.n2695 4.05904
R12697 gnd.n3652 gnd.n3651 4.05904
R12698 gnd.n15 gnd.n7 3.99943
R12699 gnd.n2996 gnd.t42 3.82437
R12700 gnd.n3026 gnd.t37 3.82437
R12701 gnd.n1783 gnd.n1782 3.82437
R12702 gnd.n3100 gnd.n3099 3.82437
R12703 gnd.n3231 gnd.n1682 3.82437
R12704 gnd.n3280 gnd.n1660 3.82437
R12705 gnd.t35 gnd.n1652 3.82437
R12706 gnd.n1630 gnd.t48 3.82437
R12707 gnd.n4791 gnd.n4663 3.70378
R12708 gnd.n5341 gnd.n5340 3.65935
R12709 gnd.n15 gnd.n14 3.60163
R12710 gnd.n4782 gnd.n4763 3.49141
R12711 gnd.n4750 gnd.n4731 3.49141
R12712 gnd.n4718 gnd.n4699 3.49141
R12713 gnd.n4687 gnd.n4668 3.49141
R12714 gnd.n4655 gnd.n4636 3.49141
R12715 gnd.n4623 gnd.n4604 3.49141
R12716 gnd.n4591 gnd.n4572 3.49141
R12717 gnd.n4560 gnd.n4541 3.49141
R12718 gnd.n2975 gnd.n1835 3.18706
R12719 gnd.t14 gnd.n3129 3.18706
R12720 gnd.n3091 gnd.n3090 3.18706
R12721 gnd.n3207 gnd.n3206 3.18706
R12722 gnd.n1684 gnd.t12 3.18706
R12723 gnd.n3712 gnd.n1529 3.18706
R12724 gnd.n5517 gnd.t294 2.8684
R12725 gnd.t307 gnd.n2926 2.8684
R12726 gnd.t2 gnd.t134 2.8684
R12727 gnd.n1559 gnd.t152 2.8684
R12728 gnd.n5324 gnd.t268 2.82907
R12729 gnd.n5324 gnd.t222 2.82907
R12730 gnd.n5326 gnd.t255 2.82907
R12731 gnd.n5326 gnd.t158 2.82907
R12732 gnd.n5328 gnd.t182 2.82907
R12733 gnd.n5328 gnd.t164 2.82907
R12734 gnd.n5330 gnd.t162 2.82907
R12735 gnd.n5330 gnd.t278 2.82907
R12736 gnd.n5332 gnd.t168 2.82907
R12737 gnd.n5332 gnd.t216 2.82907
R12738 gnd.n5334 gnd.t244 2.82907
R12739 gnd.n5334 gnd.t170 2.82907
R12740 gnd.n5336 gnd.t228 2.82907
R12741 gnd.n5336 gnd.t172 2.82907
R12742 gnd.n5293 gnd.t177 2.82907
R12743 gnd.n5293 gnd.t200 2.82907
R12744 gnd.n5295 gnd.t213 2.82907
R12745 gnd.n5295 gnd.t270 2.82907
R12746 gnd.n5297 gnd.t195 2.82907
R12747 gnd.n5297 gnd.t187 2.82907
R12748 gnd.n5299 gnd.t233 2.82907
R12749 gnd.n5299 gnd.t223 2.82907
R12750 gnd.n5301 gnd.t275 2.82907
R12751 gnd.n5301 gnd.t206 2.82907
R12752 gnd.n5303 gnd.t219 2.82907
R12753 gnd.n5303 gnd.t245 2.82907
R12754 gnd.n5305 gnd.t258 2.82907
R12755 gnd.n5305 gnd.t194 2.82907
R12756 gnd.n5308 gnd.t277 2.82907
R12757 gnd.n5308 gnd.t179 2.82907
R12758 gnd.n5310 gnd.t191 2.82907
R12759 gnd.n5310 gnd.t248 2.82907
R12760 gnd.n5312 gnd.t174 2.82907
R12761 gnd.n5312 gnd.t283 2.82907
R12762 gnd.n5314 gnd.t212 2.82907
R12763 gnd.n5314 gnd.t203 2.82907
R12764 gnd.n5316 gnd.t259 2.82907
R12765 gnd.n5316 gnd.t186 2.82907
R12766 gnd.n5318 gnd.t199 2.82907
R12767 gnd.n5318 gnd.t221 2.82907
R12768 gnd.n5320 gnd.t236 2.82907
R12769 gnd.n5320 gnd.t175 2.82907
R12770 gnd.n59 gnd.t266 2.82907
R12771 gnd.n59 gnd.t193 2.82907
R12772 gnd.n57 gnd.t284 2.82907
R12773 gnd.n57 gnd.t208 2.82907
R12774 gnd.n55 gnd.t181 2.82907
R12775 gnd.n55 gnd.t276 2.82907
R12776 gnd.n53 gnd.t251 2.82907
R12777 gnd.n53 gnd.t262 2.82907
R12778 gnd.n51 gnd.t264 2.82907
R12779 gnd.n51 gnd.t281 2.82907
R12780 gnd.n49 gnd.t260 2.82907
R12781 gnd.n49 gnd.t215 2.82907
R12782 gnd.n47 gnd.t189 2.82907
R12783 gnd.n47 gnd.t250 2.82907
R12784 gnd.n28 gnd.t225 2.82907
R12785 gnd.n28 gnd.t279 2.82907
R12786 gnd.n26 gnd.t272 2.82907
R12787 gnd.n26 gnd.t252 2.82907
R12788 gnd.n24 gnd.t237 2.82907
R12789 gnd.n24 gnd.t269 2.82907
R12790 gnd.n22 gnd.t257 2.82907
R12791 gnd.n22 gnd.t265 2.82907
R12792 gnd.n20 gnd.t218 2.82907
R12793 gnd.n20 gnd.t184 2.82907
R12794 gnd.n18 gnd.t166 2.82907
R12795 gnd.n18 gnd.t243 2.82907
R12796 gnd.n16 gnd.t229 2.82907
R12797 gnd.n16 gnd.t282 2.82907
R12798 gnd.n43 gnd.t205 2.82907
R12799 gnd.n43 gnd.t267 2.82907
R12800 gnd.n41 gnd.t254 2.82907
R12801 gnd.n41 gnd.t226 2.82907
R12802 gnd.n39 gnd.t217 2.82907
R12803 gnd.n39 gnd.t247 2.82907
R12804 gnd.n37 gnd.t235 2.82907
R12805 gnd.n37 gnd.t241 2.82907
R12806 gnd.n35 gnd.t197 2.82907
R12807 gnd.n35 gnd.t280 2.82907
R12808 gnd.n33 gnd.t274 2.82907
R12809 gnd.n33 gnd.t220 2.82907
R12810 gnd.n31 gnd.t209 2.82907
R12811 gnd.n31 gnd.t271 2.82907
R12812 gnd.n4779 gnd.n4778 2.71565
R12813 gnd.n4747 gnd.n4746 2.71565
R12814 gnd.n4715 gnd.n4714 2.71565
R12815 gnd.n4684 gnd.n4683 2.71565
R12816 gnd.n4652 gnd.n4651 2.71565
R12817 gnd.n4620 gnd.n4619 2.71565
R12818 gnd.n4588 gnd.n4587 2.71565
R12819 gnd.n4557 gnd.n4556 2.71565
R12820 gnd.n1813 gnd.t101 2.54975
R12821 gnd.n3043 gnd.n3042 2.54975
R12822 gnd.n3146 gnd.n1742 2.54975
R12823 gnd.n3090 gnd.t13 2.54975
R12824 gnd.n3166 gnd.t24 2.54975
R12825 gnd.n3196 gnd.t287 2.54975
R12826 gnd.n3206 gnd.t17 2.54975
R12827 gnd.n3205 gnd.n1691 2.54975
R12828 gnd.n3299 gnd.n1644 2.54975
R12829 gnd.n5342 gnd.n5341 2.27742
R12830 gnd.n5341 gnd.n5292 2.27742
R12831 gnd.n5341 gnd.n5285 2.27742
R12832 gnd.n5341 gnd.n5258 2.27742
R12833 gnd.n6776 gnd.n6775 2.27742
R12834 gnd.n6776 gnd.n263 2.27742
R12835 gnd.n6776 gnd.n262 2.27742
R12836 gnd.n6776 gnd.n261 2.27742
R12837 gnd.n1047 gnd.n1046 2.27742
R12838 gnd.n1048 gnd.n1047 2.27742
R12839 gnd.n4282 gnd.n1047 2.27742
R12840 gnd.n1064 gnd.n1047 2.27742
R12841 gnd.t67 gnd.n5455 2.23109
R12842 gnd.t304 gnd.n5568 2.23109
R12843 gnd.n3130 gnd.t6 2.23109
R12844 gnd.n3239 gnd.t33 2.23109
R12845 gnd.n4775 gnd.n4765 1.93989
R12846 gnd.n4743 gnd.n4733 1.93989
R12847 gnd.n4711 gnd.n4701 1.93989
R12848 gnd.n4680 gnd.n4670 1.93989
R12849 gnd.n4648 gnd.n4638 1.93989
R12850 gnd.n4616 gnd.n4606 1.93989
R12851 gnd.n4584 gnd.n4574 1.93989
R12852 gnd.n4553 gnd.n4543 1.93989
R12853 gnd.t137 gnd.n3035 1.91244
R12854 gnd.n3033 gnd.t286 1.91244
R12855 gnd.t154 gnd.n1761 1.91244
R12856 gnd.n3140 gnd.n1746 1.91244
R12857 gnd.n3069 gnd.n3068 1.91244
R12858 gnd.n3224 gnd.t288 1.91244
R12859 gnd.t285 gnd.n3297 1.91244
R12860 gnd.n5364 gnd.t31 1.59378
R12861 gnd.n5272 gnd.t301 1.59378
R12862 gnd.n5681 gnd.t18 1.59378
R12863 gnd.t29 gnd.n3052 1.59378
R12864 gnd.t22 gnd.n3264 1.59378
R12865 gnd.t121 gnd.n1828 1.27512
R12866 gnd.n3011 gnd.n3010 1.27512
R12867 gnd.n3044 gnd.t286 1.27512
R12868 gnd.n3166 gnd.n1726 1.27512
R12869 gnd.n3196 gnd.n3194 1.27512
R12870 gnd.n3298 gnd.t285 1.27512
R12871 gnd.n3309 gnd.n3308 1.27512
R12872 gnd.n3622 gnd.n1534 1.27512
R12873 gnd.n5151 gnd.n5150 1.16414
R12874 gnd.n5813 gnd.n4520 1.16414
R12875 gnd.n4774 gnd.n4767 1.16414
R12876 gnd.n4742 gnd.n4735 1.16414
R12877 gnd.n4710 gnd.n4703 1.16414
R12878 gnd.n4679 gnd.n4672 1.16414
R12879 gnd.n4647 gnd.n4640 1.16414
R12880 gnd.n4615 gnd.n4608 1.16414
R12881 gnd.n4583 gnd.n4576 1.16414
R12882 gnd.n4552 gnd.n4545 1.16414
R12883 gnd.n3840 gnd.n1485 0.970197
R12884 gnd.n2758 gnd.n2090 0.970197
R12885 gnd.n4758 gnd.n4726 0.962709
R12886 gnd.n4790 gnd.n4758 0.962709
R12887 gnd.n4631 gnd.n4599 0.962709
R12888 gnd.n4663 gnd.n4631 0.962709
R12889 gnd.t309 gnd.n4979 0.956468
R12890 gnd.n5671 gnd.t300 0.956468
R12891 gnd.n2446 gnd.t176 0.956468
R12892 gnd.t311 gnd.n1923 0.956468
R12893 gnd.t6 gnd.t14 0.956468
R12894 gnd.t12 gnd.t33 0.956468
R12895 gnd.n3371 gnd.t4 0.956468
R12896 gnd.n3959 gnd.t249 0.956468
R12897 gnd.n5333 gnd.n5331 0.773756
R12898 gnd.n56 gnd.n54 0.773756
R12899 gnd.n5338 gnd.n5337 0.773756
R12900 gnd.n5337 gnd.n5335 0.773756
R12901 gnd.n5335 gnd.n5333 0.773756
R12902 gnd.n5331 gnd.n5329 0.773756
R12903 gnd.n5329 gnd.n5327 0.773756
R12904 gnd.n5327 gnd.n5325 0.773756
R12905 gnd.n50 gnd.n48 0.773756
R12906 gnd.n52 gnd.n50 0.773756
R12907 gnd.n54 gnd.n52 0.773756
R12908 gnd.n58 gnd.n56 0.773756
R12909 gnd.n60 gnd.n58 0.773756
R12910 gnd.n61 gnd.n60 0.773756
R12911 gnd.n2 gnd.n1 0.672012
R12912 gnd.n3 gnd.n2 0.672012
R12913 gnd.n4 gnd.n3 0.672012
R12914 gnd.n5 gnd.n4 0.672012
R12915 gnd.n6 gnd.n5 0.672012
R12916 gnd.n7 gnd.n6 0.672012
R12917 gnd.n9 gnd.n8 0.672012
R12918 gnd.n10 gnd.n9 0.672012
R12919 gnd.n11 gnd.n10 0.672012
R12920 gnd.n12 gnd.n11 0.672012
R12921 gnd.n13 gnd.n12 0.672012
R12922 gnd.n14 gnd.n13 0.672012
R12923 gnd.n3060 gnd.t36 0.637812
R12924 gnd.n3111 gnd.n1769 0.637812
R12925 gnd.n3121 gnd.n1755 0.637812
R12926 gnd.n3238 gnd.n1676 0.637812
R12927 gnd.n3274 gnd.n1664 0.637812
R12928 gnd.n3271 gnd.t151 0.637812
R12929 gnd.n3339 gnd.t118 0.637812
R12930 gnd gnd.n0 0.59317
R12931 gnd.n5307 gnd.n5306 0.573776
R12932 gnd.n5306 gnd.n5304 0.573776
R12933 gnd.n5304 gnd.n5302 0.573776
R12934 gnd.n5302 gnd.n5300 0.573776
R12935 gnd.n5300 gnd.n5298 0.573776
R12936 gnd.n5298 gnd.n5296 0.573776
R12937 gnd.n5296 gnd.n5294 0.573776
R12938 gnd.n5322 gnd.n5321 0.573776
R12939 gnd.n5321 gnd.n5319 0.573776
R12940 gnd.n5319 gnd.n5317 0.573776
R12941 gnd.n5317 gnd.n5315 0.573776
R12942 gnd.n5315 gnd.n5313 0.573776
R12943 gnd.n5313 gnd.n5311 0.573776
R12944 gnd.n5311 gnd.n5309 0.573776
R12945 gnd.n19 gnd.n17 0.573776
R12946 gnd.n21 gnd.n19 0.573776
R12947 gnd.n23 gnd.n21 0.573776
R12948 gnd.n25 gnd.n23 0.573776
R12949 gnd.n27 gnd.n25 0.573776
R12950 gnd.n29 gnd.n27 0.573776
R12951 gnd.n30 gnd.n29 0.573776
R12952 gnd.n34 gnd.n32 0.573776
R12953 gnd.n36 gnd.n34 0.573776
R12954 gnd.n38 gnd.n36 0.573776
R12955 gnd.n40 gnd.n38 0.573776
R12956 gnd.n42 gnd.n40 0.573776
R12957 gnd.n44 gnd.n42 0.573776
R12958 gnd.n45 gnd.n44 0.573776
R12959 gnd.n7058 gnd.n7057 0.553533
R12960 gnd.n6776 gnd.n260 0.5435
R12961 gnd.n2160 gnd.n1047 0.5435
R12962 gnd.n4201 gnd.n4200 0.523366
R12963 gnd.n3445 gnd.n1302 0.523366
R12964 gnd.n2300 gnd.n2298 0.505073
R12965 gnd.n2338 gnd.n2337 0.505073
R12966 gnd.n6917 gnd.n6916 0.505073
R12967 gnd.n6888 gnd.n98 0.505073
R12968 gnd.n7011 gnd.n7010 0.492878
R12969 gnd.n6940 gnd.n6939 0.492878
R12970 gnd.n3894 gnd.n3893 0.492878
R12971 gnd.n3798 gnd.n1331 0.492878
R12972 gnd.n2074 gnd.n1189 0.492878
R12973 gnd.n2585 gnd.n2584 0.492878
R12974 gnd.n4368 gnd.n932 0.492878
R12975 gnd.n2347 gnd.n889 0.492878
R12976 gnd.n3567 gnd.n3566 0.489829
R12977 gnd.n2851 gnd.n1958 0.489829
R12978 gnd.n5803 gnd.n5802 0.486781
R12979 gnd.n5203 gnd.n5099 0.48678
R12980 gnd.n5884 gnd.n5883 0.480683
R12981 gnd.n5384 gnd.n5050 0.480683
R12982 gnd.n6067 gnd.n675 0.438
R12983 gnd.n6420 gnd.n6419 0.438
R12984 gnd.n4203 gnd.n4202 0.404992
R12985 gnd.n3448 gnd.n3447 0.404992
R12986 gnd.n2565 gnd.n2553 0.388379
R12987 gnd.n4771 gnd.n4770 0.388379
R12988 gnd.n4739 gnd.n4738 0.388379
R12989 gnd.n4707 gnd.n4706 0.388379
R12990 gnd.n4676 gnd.n4675 0.388379
R12991 gnd.n4644 gnd.n4643 0.388379
R12992 gnd.n4612 gnd.n4611 0.388379
R12993 gnd.n4580 gnd.n4579 0.388379
R12994 gnd.n4549 gnd.n4548 0.388379
R12995 gnd.n6980 gnd.n6979 0.388379
R12996 gnd.n4409 gnd.n4408 0.388379
R12997 gnd.n3556 gnd.n3555 0.388379
R12998 gnd.n6631 gnd.n260 0.381598
R12999 gnd.n2160 gnd.n2159 0.381598
R13000 gnd.n7058 gnd.n15 0.374463
R13001 gnd.n5750 gnd.t296 0.319156
R13002 gnd.n2183 gnd.t163 0.319156
R13003 gnd.n2858 gnd.t114 0.319156
R13004 gnd.n3053 gnd.t29 0.319156
R13005 gnd.n3265 gnd.t22 0.319156
R13006 gnd.t85 gnd.n3572 0.319156
R13007 gnd.t196 gnd.n315 0.319156
R13008 gnd.n5197 gnd.n5196 0.311721
R13009 gnd gnd.n7058 0.295112
R13010 gnd.n2576 gnd.n2575 0.27489
R13011 gnd.n3535 gnd.n1459 0.27489
R13012 gnd.n5853 gnd.n5852 0.268793
R13013 gnd.n5852 gnd.n5851 0.241354
R13014 gnd.n3841 gnd.n1486 0.229039
R13015 gnd.n3842 gnd.n3841 0.229039
R13016 gnd.n2628 gnd.n2089 0.229039
R13017 gnd.n2628 gnd.n2627 0.229039
R13018 gnd.n5439 gnd.n5067 0.206293
R13019 gnd.n5340 gnd.n0 0.169152
R13020 gnd.n4788 gnd.n4760 0.155672
R13021 gnd.n4781 gnd.n4760 0.155672
R13022 gnd.n4781 gnd.n4780 0.155672
R13023 gnd.n4780 gnd.n4764 0.155672
R13024 gnd.n4773 gnd.n4764 0.155672
R13025 gnd.n4773 gnd.n4772 0.155672
R13026 gnd.n4756 gnd.n4728 0.155672
R13027 gnd.n4749 gnd.n4728 0.155672
R13028 gnd.n4749 gnd.n4748 0.155672
R13029 gnd.n4748 gnd.n4732 0.155672
R13030 gnd.n4741 gnd.n4732 0.155672
R13031 gnd.n4741 gnd.n4740 0.155672
R13032 gnd.n4724 gnd.n4696 0.155672
R13033 gnd.n4717 gnd.n4696 0.155672
R13034 gnd.n4717 gnd.n4716 0.155672
R13035 gnd.n4716 gnd.n4700 0.155672
R13036 gnd.n4709 gnd.n4700 0.155672
R13037 gnd.n4709 gnd.n4708 0.155672
R13038 gnd.n4693 gnd.n4665 0.155672
R13039 gnd.n4686 gnd.n4665 0.155672
R13040 gnd.n4686 gnd.n4685 0.155672
R13041 gnd.n4685 gnd.n4669 0.155672
R13042 gnd.n4678 gnd.n4669 0.155672
R13043 gnd.n4678 gnd.n4677 0.155672
R13044 gnd.n4661 gnd.n4633 0.155672
R13045 gnd.n4654 gnd.n4633 0.155672
R13046 gnd.n4654 gnd.n4653 0.155672
R13047 gnd.n4653 gnd.n4637 0.155672
R13048 gnd.n4646 gnd.n4637 0.155672
R13049 gnd.n4646 gnd.n4645 0.155672
R13050 gnd.n4629 gnd.n4601 0.155672
R13051 gnd.n4622 gnd.n4601 0.155672
R13052 gnd.n4622 gnd.n4621 0.155672
R13053 gnd.n4621 gnd.n4605 0.155672
R13054 gnd.n4614 gnd.n4605 0.155672
R13055 gnd.n4614 gnd.n4613 0.155672
R13056 gnd.n4597 gnd.n4569 0.155672
R13057 gnd.n4590 gnd.n4569 0.155672
R13058 gnd.n4590 gnd.n4589 0.155672
R13059 gnd.n4589 gnd.n4573 0.155672
R13060 gnd.n4582 gnd.n4573 0.155672
R13061 gnd.n4582 gnd.n4581 0.155672
R13062 gnd.n4566 gnd.n4538 0.155672
R13063 gnd.n4559 gnd.n4538 0.155672
R13064 gnd.n4559 gnd.n4558 0.155672
R13065 gnd.n4558 gnd.n4542 0.155672
R13066 gnd.n4551 gnd.n4542 0.155672
R13067 gnd.n4551 gnd.n4550 0.155672
R13068 gnd.n5883 gnd.n4450 0.152939
R13069 gnd.n4452 gnd.n4450 0.152939
R13070 gnd.n4456 gnd.n4452 0.152939
R13071 gnd.n4457 gnd.n4456 0.152939
R13072 gnd.n4458 gnd.n4457 0.152939
R13073 gnd.n4459 gnd.n4458 0.152939
R13074 gnd.n4463 gnd.n4459 0.152939
R13075 gnd.n4464 gnd.n4463 0.152939
R13076 gnd.n4465 gnd.n4464 0.152939
R13077 gnd.n4466 gnd.n4465 0.152939
R13078 gnd.n4470 gnd.n4466 0.152939
R13079 gnd.n4471 gnd.n4470 0.152939
R13080 gnd.n4472 gnd.n4471 0.152939
R13081 gnd.n4473 gnd.n4472 0.152939
R13082 gnd.n4478 gnd.n4473 0.152939
R13083 gnd.n5853 gnd.n4478 0.152939
R13084 gnd.n5459 gnd.n5050 0.152939
R13085 gnd.n5460 gnd.n5459 0.152939
R13086 gnd.n5461 gnd.n5460 0.152939
R13087 gnd.n5462 gnd.n5461 0.152939
R13088 gnd.n5462 gnd.n5025 0.152939
R13089 gnd.n5490 gnd.n5025 0.152939
R13090 gnd.n5491 gnd.n5490 0.152939
R13091 gnd.n5492 gnd.n5491 0.152939
R13092 gnd.n5493 gnd.n5492 0.152939
R13093 gnd.n5493 gnd.n4999 0.152939
R13094 gnd.n5521 gnd.n4999 0.152939
R13095 gnd.n5522 gnd.n5521 0.152939
R13096 gnd.n5523 gnd.n5522 0.152939
R13097 gnd.n5524 gnd.n5523 0.152939
R13098 gnd.n5524 gnd.n4973 0.152939
R13099 gnd.n5552 gnd.n4973 0.152939
R13100 gnd.n5553 gnd.n5552 0.152939
R13101 gnd.n5554 gnd.n5553 0.152939
R13102 gnd.n5555 gnd.n5554 0.152939
R13103 gnd.n5555 gnd.n4947 0.152939
R13104 gnd.n5583 gnd.n4947 0.152939
R13105 gnd.n5584 gnd.n5583 0.152939
R13106 gnd.n5585 gnd.n5584 0.152939
R13107 gnd.n5586 gnd.n5585 0.152939
R13108 gnd.n5586 gnd.n4922 0.152939
R13109 gnd.n5614 gnd.n4922 0.152939
R13110 gnd.n5615 gnd.n5614 0.152939
R13111 gnd.n5616 gnd.n5615 0.152939
R13112 gnd.n5617 gnd.n5616 0.152939
R13113 gnd.n5617 gnd.n4898 0.152939
R13114 gnd.n5644 gnd.n4898 0.152939
R13115 gnd.n5645 gnd.n5644 0.152939
R13116 gnd.n5646 gnd.n5645 0.152939
R13117 gnd.n5647 gnd.n5646 0.152939
R13118 gnd.n5647 gnd.n4866 0.152939
R13119 gnd.n5685 gnd.n4866 0.152939
R13120 gnd.n5686 gnd.n5685 0.152939
R13121 gnd.n5687 gnd.n5686 0.152939
R13122 gnd.n5688 gnd.n5687 0.152939
R13123 gnd.n5689 gnd.n5688 0.152939
R13124 gnd.n5689 gnd.n4836 0.152939
R13125 gnd.n5732 gnd.n4836 0.152939
R13126 gnd.n5733 gnd.n5732 0.152939
R13127 gnd.n5734 gnd.n5733 0.152939
R13128 gnd.n5735 gnd.n5734 0.152939
R13129 gnd.n5736 gnd.n5735 0.152939
R13130 gnd.n5736 gnd.n4809 0.152939
R13131 gnd.n5776 gnd.n4809 0.152939
R13132 gnd.n5777 gnd.n5776 0.152939
R13133 gnd.n5778 gnd.n5777 0.152939
R13134 gnd.n5779 gnd.n5778 0.152939
R13135 gnd.n5779 gnd.n4449 0.152939
R13136 gnd.n5884 gnd.n4449 0.152939
R13137 gnd.n5385 gnd.n5384 0.152939
R13138 gnd.n5386 gnd.n5385 0.152939
R13139 gnd.n5387 gnd.n5386 0.152939
R13140 gnd.n5388 gnd.n5387 0.152939
R13141 gnd.n5389 gnd.n5388 0.152939
R13142 gnd.n5390 gnd.n5389 0.152939
R13143 gnd.n5391 gnd.n5390 0.152939
R13144 gnd.n5392 gnd.n5391 0.152939
R13145 gnd.n5393 gnd.n5392 0.152939
R13146 gnd.n5394 gnd.n5393 0.152939
R13147 gnd.n5395 gnd.n5394 0.152939
R13148 gnd.n5396 gnd.n5395 0.152939
R13149 gnd.n5397 gnd.n5396 0.152939
R13150 gnd.n5398 gnd.n5397 0.152939
R13151 gnd.n5402 gnd.n5398 0.152939
R13152 gnd.n5402 gnd.n5067 0.152939
R13153 gnd.n5851 gnd.n4480 0.152939
R13154 gnd.n4482 gnd.n4480 0.152939
R13155 gnd.n4486 gnd.n4482 0.152939
R13156 gnd.n4487 gnd.n4486 0.152939
R13157 gnd.n4488 gnd.n4487 0.152939
R13158 gnd.n4489 gnd.n4488 0.152939
R13159 gnd.n4493 gnd.n4489 0.152939
R13160 gnd.n4494 gnd.n4493 0.152939
R13161 gnd.n4495 gnd.n4494 0.152939
R13162 gnd.n4496 gnd.n4495 0.152939
R13163 gnd.n4500 gnd.n4496 0.152939
R13164 gnd.n4501 gnd.n4500 0.152939
R13165 gnd.n4502 gnd.n4501 0.152939
R13166 gnd.n4503 gnd.n4502 0.152939
R13167 gnd.n4507 gnd.n4503 0.152939
R13168 gnd.n4508 gnd.n4507 0.152939
R13169 gnd.n4509 gnd.n4508 0.152939
R13170 gnd.n4510 gnd.n4509 0.152939
R13171 gnd.n4514 gnd.n4510 0.152939
R13172 gnd.n4515 gnd.n4514 0.152939
R13173 gnd.n4516 gnd.n4515 0.152939
R13174 gnd.n4517 gnd.n4516 0.152939
R13175 gnd.n4524 gnd.n4517 0.152939
R13176 gnd.n4525 gnd.n4524 0.152939
R13177 gnd.n4526 gnd.n4525 0.152939
R13178 gnd.n5803 gnd.n4526 0.152939
R13179 gnd.n5259 gnd.n5257 0.152939
R13180 gnd.n5260 gnd.n5259 0.152939
R13181 gnd.n5261 gnd.n5260 0.152939
R13182 gnd.n5262 gnd.n5261 0.152939
R13183 gnd.n5263 gnd.n5262 0.152939
R13184 gnd.n5264 gnd.n5263 0.152939
R13185 gnd.n5265 gnd.n5264 0.152939
R13186 gnd.n5265 gnd.n4884 0.152939
R13187 gnd.n5664 gnd.n4884 0.152939
R13188 gnd.n5665 gnd.n5664 0.152939
R13189 gnd.n5666 gnd.n5665 0.152939
R13190 gnd.n5667 gnd.n5666 0.152939
R13191 gnd.n5667 gnd.n4849 0.152939
R13192 gnd.n5708 gnd.n4849 0.152939
R13193 gnd.n5709 gnd.n5708 0.152939
R13194 gnd.n5710 gnd.n5709 0.152939
R13195 gnd.n5711 gnd.n5710 0.152939
R13196 gnd.n5711 gnd.n4822 0.152939
R13197 gnd.n5753 gnd.n4822 0.152939
R13198 gnd.n5754 gnd.n5753 0.152939
R13199 gnd.n5755 gnd.n5754 0.152939
R13200 gnd.n5756 gnd.n5755 0.152939
R13201 gnd.n5756 gnd.n4529 0.152939
R13202 gnd.n5794 gnd.n4529 0.152939
R13203 gnd.n5795 gnd.n5794 0.152939
R13204 gnd.n5796 gnd.n5795 0.152939
R13205 gnd.n5796 gnd.n4527 0.152939
R13206 gnd.n5802 gnd.n4527 0.152939
R13207 gnd.n5204 gnd.n5203 0.152939
R13208 gnd.n5205 gnd.n5204 0.152939
R13209 gnd.n5205 gnd.n5087 0.152939
R13210 gnd.n5219 gnd.n5087 0.152939
R13211 gnd.n5220 gnd.n5219 0.152939
R13212 gnd.n5221 gnd.n5220 0.152939
R13213 gnd.n5221 gnd.n5074 0.152939
R13214 gnd.n5235 gnd.n5074 0.152939
R13215 gnd.n5236 gnd.n5235 0.152939
R13216 gnd.n5237 gnd.n5236 0.152939
R13217 gnd.n5238 gnd.n5237 0.152939
R13218 gnd.n5239 gnd.n5238 0.152939
R13219 gnd.n5240 gnd.n5239 0.152939
R13220 gnd.n5241 gnd.n5240 0.152939
R13221 gnd.n5242 gnd.n5241 0.152939
R13222 gnd.n5243 gnd.n5242 0.152939
R13223 gnd.n5244 gnd.n5243 0.152939
R13224 gnd.n5245 gnd.n5244 0.152939
R13225 gnd.n5246 gnd.n5245 0.152939
R13226 gnd.n5247 gnd.n5246 0.152939
R13227 gnd.n5248 gnd.n5247 0.152939
R13228 gnd.n5249 gnd.n5248 0.152939
R13229 gnd.n5250 gnd.n5249 0.152939
R13230 gnd.n5251 gnd.n5250 0.152939
R13231 gnd.n5252 gnd.n5251 0.152939
R13232 gnd.n5253 gnd.n5252 0.152939
R13233 gnd.n5254 gnd.n5253 0.152939
R13234 gnd.n5255 gnd.n5254 0.152939
R13235 gnd.n5196 gnd.n5103 0.152939
R13236 gnd.n5106 gnd.n5103 0.152939
R13237 gnd.n5107 gnd.n5106 0.152939
R13238 gnd.n5108 gnd.n5107 0.152939
R13239 gnd.n5111 gnd.n5108 0.152939
R13240 gnd.n5112 gnd.n5111 0.152939
R13241 gnd.n5113 gnd.n5112 0.152939
R13242 gnd.n5114 gnd.n5113 0.152939
R13243 gnd.n5117 gnd.n5114 0.152939
R13244 gnd.n5118 gnd.n5117 0.152939
R13245 gnd.n5119 gnd.n5118 0.152939
R13246 gnd.n5120 gnd.n5119 0.152939
R13247 gnd.n5123 gnd.n5120 0.152939
R13248 gnd.n5124 gnd.n5123 0.152939
R13249 gnd.n5125 gnd.n5124 0.152939
R13250 gnd.n5126 gnd.n5125 0.152939
R13251 gnd.n5129 gnd.n5126 0.152939
R13252 gnd.n5130 gnd.n5129 0.152939
R13253 gnd.n5131 gnd.n5130 0.152939
R13254 gnd.n5132 gnd.n5131 0.152939
R13255 gnd.n5135 gnd.n5132 0.152939
R13256 gnd.n5136 gnd.n5135 0.152939
R13257 gnd.n5139 gnd.n5136 0.152939
R13258 gnd.n5140 gnd.n5139 0.152939
R13259 gnd.n5142 gnd.n5140 0.152939
R13260 gnd.n5142 gnd.n5099 0.152939
R13261 gnd.n6068 gnd.n6067 0.152939
R13262 gnd.n6069 gnd.n6068 0.152939
R13263 gnd.n6069 gnd.n669 0.152939
R13264 gnd.n6077 gnd.n669 0.152939
R13265 gnd.n6078 gnd.n6077 0.152939
R13266 gnd.n6079 gnd.n6078 0.152939
R13267 gnd.n6079 gnd.n663 0.152939
R13268 gnd.n6087 gnd.n663 0.152939
R13269 gnd.n6088 gnd.n6087 0.152939
R13270 gnd.n6089 gnd.n6088 0.152939
R13271 gnd.n6089 gnd.n657 0.152939
R13272 gnd.n6097 gnd.n657 0.152939
R13273 gnd.n6098 gnd.n6097 0.152939
R13274 gnd.n6099 gnd.n6098 0.152939
R13275 gnd.n6099 gnd.n651 0.152939
R13276 gnd.n6107 gnd.n651 0.152939
R13277 gnd.n6108 gnd.n6107 0.152939
R13278 gnd.n6109 gnd.n6108 0.152939
R13279 gnd.n6109 gnd.n645 0.152939
R13280 gnd.n6117 gnd.n645 0.152939
R13281 gnd.n6118 gnd.n6117 0.152939
R13282 gnd.n6119 gnd.n6118 0.152939
R13283 gnd.n6119 gnd.n639 0.152939
R13284 gnd.n6127 gnd.n639 0.152939
R13285 gnd.n6128 gnd.n6127 0.152939
R13286 gnd.n6129 gnd.n6128 0.152939
R13287 gnd.n6129 gnd.n633 0.152939
R13288 gnd.n6137 gnd.n633 0.152939
R13289 gnd.n6138 gnd.n6137 0.152939
R13290 gnd.n6139 gnd.n6138 0.152939
R13291 gnd.n6139 gnd.n627 0.152939
R13292 gnd.n6147 gnd.n627 0.152939
R13293 gnd.n6148 gnd.n6147 0.152939
R13294 gnd.n6149 gnd.n6148 0.152939
R13295 gnd.n6149 gnd.n621 0.152939
R13296 gnd.n6157 gnd.n621 0.152939
R13297 gnd.n6158 gnd.n6157 0.152939
R13298 gnd.n6159 gnd.n6158 0.152939
R13299 gnd.n6159 gnd.n615 0.152939
R13300 gnd.n6167 gnd.n615 0.152939
R13301 gnd.n6168 gnd.n6167 0.152939
R13302 gnd.n6169 gnd.n6168 0.152939
R13303 gnd.n6169 gnd.n609 0.152939
R13304 gnd.n6177 gnd.n609 0.152939
R13305 gnd.n6178 gnd.n6177 0.152939
R13306 gnd.n6179 gnd.n6178 0.152939
R13307 gnd.n6179 gnd.n603 0.152939
R13308 gnd.n6187 gnd.n603 0.152939
R13309 gnd.n6188 gnd.n6187 0.152939
R13310 gnd.n6189 gnd.n6188 0.152939
R13311 gnd.n6189 gnd.n597 0.152939
R13312 gnd.n6197 gnd.n597 0.152939
R13313 gnd.n6198 gnd.n6197 0.152939
R13314 gnd.n6199 gnd.n6198 0.152939
R13315 gnd.n6199 gnd.n591 0.152939
R13316 gnd.n6207 gnd.n591 0.152939
R13317 gnd.n6208 gnd.n6207 0.152939
R13318 gnd.n6209 gnd.n6208 0.152939
R13319 gnd.n6209 gnd.n585 0.152939
R13320 gnd.n6217 gnd.n585 0.152939
R13321 gnd.n6218 gnd.n6217 0.152939
R13322 gnd.n6219 gnd.n6218 0.152939
R13323 gnd.n6219 gnd.n579 0.152939
R13324 gnd.n6227 gnd.n579 0.152939
R13325 gnd.n6228 gnd.n6227 0.152939
R13326 gnd.n6229 gnd.n6228 0.152939
R13327 gnd.n6229 gnd.n573 0.152939
R13328 gnd.n6237 gnd.n573 0.152939
R13329 gnd.n6238 gnd.n6237 0.152939
R13330 gnd.n6239 gnd.n6238 0.152939
R13331 gnd.n6239 gnd.n567 0.152939
R13332 gnd.n6247 gnd.n567 0.152939
R13333 gnd.n6248 gnd.n6247 0.152939
R13334 gnd.n6249 gnd.n6248 0.152939
R13335 gnd.n6249 gnd.n561 0.152939
R13336 gnd.n6257 gnd.n561 0.152939
R13337 gnd.n6258 gnd.n6257 0.152939
R13338 gnd.n6259 gnd.n6258 0.152939
R13339 gnd.n6259 gnd.n555 0.152939
R13340 gnd.n6267 gnd.n555 0.152939
R13341 gnd.n6268 gnd.n6267 0.152939
R13342 gnd.n6269 gnd.n6268 0.152939
R13343 gnd.n6269 gnd.n549 0.152939
R13344 gnd.n6277 gnd.n549 0.152939
R13345 gnd.n6278 gnd.n6277 0.152939
R13346 gnd.n6279 gnd.n6278 0.152939
R13347 gnd.n6279 gnd.n543 0.152939
R13348 gnd.n6287 gnd.n543 0.152939
R13349 gnd.n6288 gnd.n6287 0.152939
R13350 gnd.n6289 gnd.n6288 0.152939
R13351 gnd.n6289 gnd.n537 0.152939
R13352 gnd.n6297 gnd.n537 0.152939
R13353 gnd.n6298 gnd.n6297 0.152939
R13354 gnd.n6299 gnd.n6298 0.152939
R13355 gnd.n6299 gnd.n531 0.152939
R13356 gnd.n6307 gnd.n531 0.152939
R13357 gnd.n6308 gnd.n6307 0.152939
R13358 gnd.n6309 gnd.n6308 0.152939
R13359 gnd.n6309 gnd.n525 0.152939
R13360 gnd.n6317 gnd.n525 0.152939
R13361 gnd.n6318 gnd.n6317 0.152939
R13362 gnd.n6319 gnd.n6318 0.152939
R13363 gnd.n6319 gnd.n519 0.152939
R13364 gnd.n6327 gnd.n519 0.152939
R13365 gnd.n6328 gnd.n6327 0.152939
R13366 gnd.n6329 gnd.n6328 0.152939
R13367 gnd.n6329 gnd.n513 0.152939
R13368 gnd.n6337 gnd.n513 0.152939
R13369 gnd.n6338 gnd.n6337 0.152939
R13370 gnd.n6339 gnd.n6338 0.152939
R13371 gnd.n6339 gnd.n507 0.152939
R13372 gnd.n6347 gnd.n507 0.152939
R13373 gnd.n6348 gnd.n6347 0.152939
R13374 gnd.n6349 gnd.n6348 0.152939
R13375 gnd.n6349 gnd.n501 0.152939
R13376 gnd.n6357 gnd.n501 0.152939
R13377 gnd.n6358 gnd.n6357 0.152939
R13378 gnd.n6359 gnd.n6358 0.152939
R13379 gnd.n6359 gnd.n495 0.152939
R13380 gnd.n6367 gnd.n495 0.152939
R13381 gnd.n6368 gnd.n6367 0.152939
R13382 gnd.n6369 gnd.n6368 0.152939
R13383 gnd.n6369 gnd.n489 0.152939
R13384 gnd.n6377 gnd.n489 0.152939
R13385 gnd.n6378 gnd.n6377 0.152939
R13386 gnd.n6379 gnd.n6378 0.152939
R13387 gnd.n6379 gnd.n483 0.152939
R13388 gnd.n6387 gnd.n483 0.152939
R13389 gnd.n6388 gnd.n6387 0.152939
R13390 gnd.n6389 gnd.n6388 0.152939
R13391 gnd.n6389 gnd.n477 0.152939
R13392 gnd.n6397 gnd.n477 0.152939
R13393 gnd.n6398 gnd.n6397 0.152939
R13394 gnd.n6399 gnd.n6398 0.152939
R13395 gnd.n6399 gnd.n471 0.152939
R13396 gnd.n6407 gnd.n471 0.152939
R13397 gnd.n6408 gnd.n6407 0.152939
R13398 gnd.n6410 gnd.n6408 0.152939
R13399 gnd.n6410 gnd.n6409 0.152939
R13400 gnd.n6409 gnd.n465 0.152939
R13401 gnd.n6419 gnd.n465 0.152939
R13402 gnd.n6420 gnd.n460 0.152939
R13403 gnd.n6428 gnd.n460 0.152939
R13404 gnd.n6429 gnd.n6428 0.152939
R13405 gnd.n6430 gnd.n6429 0.152939
R13406 gnd.n6430 gnd.n454 0.152939
R13407 gnd.n6438 gnd.n454 0.152939
R13408 gnd.n6439 gnd.n6438 0.152939
R13409 gnd.n6440 gnd.n6439 0.152939
R13410 gnd.n6440 gnd.n448 0.152939
R13411 gnd.n6448 gnd.n448 0.152939
R13412 gnd.n6449 gnd.n6448 0.152939
R13413 gnd.n6450 gnd.n6449 0.152939
R13414 gnd.n6450 gnd.n442 0.152939
R13415 gnd.n6458 gnd.n442 0.152939
R13416 gnd.n6459 gnd.n6458 0.152939
R13417 gnd.n6460 gnd.n6459 0.152939
R13418 gnd.n6460 gnd.n436 0.152939
R13419 gnd.n6468 gnd.n436 0.152939
R13420 gnd.n6469 gnd.n6468 0.152939
R13421 gnd.n6470 gnd.n6469 0.152939
R13422 gnd.n6470 gnd.n430 0.152939
R13423 gnd.n6478 gnd.n430 0.152939
R13424 gnd.n6479 gnd.n6478 0.152939
R13425 gnd.n6480 gnd.n6479 0.152939
R13426 gnd.n6480 gnd.n424 0.152939
R13427 gnd.n6488 gnd.n424 0.152939
R13428 gnd.n6489 gnd.n6488 0.152939
R13429 gnd.n6490 gnd.n6489 0.152939
R13430 gnd.n6490 gnd.n418 0.152939
R13431 gnd.n6498 gnd.n418 0.152939
R13432 gnd.n6499 gnd.n6498 0.152939
R13433 gnd.n6500 gnd.n6499 0.152939
R13434 gnd.n6500 gnd.n412 0.152939
R13435 gnd.n6508 gnd.n412 0.152939
R13436 gnd.n6509 gnd.n6508 0.152939
R13437 gnd.n6510 gnd.n6509 0.152939
R13438 gnd.n6510 gnd.n406 0.152939
R13439 gnd.n6518 gnd.n406 0.152939
R13440 gnd.n6519 gnd.n6518 0.152939
R13441 gnd.n6520 gnd.n6519 0.152939
R13442 gnd.n6520 gnd.n400 0.152939
R13443 gnd.n6528 gnd.n400 0.152939
R13444 gnd.n6529 gnd.n6528 0.152939
R13445 gnd.n6530 gnd.n6529 0.152939
R13446 gnd.n6530 gnd.n394 0.152939
R13447 gnd.n6538 gnd.n394 0.152939
R13448 gnd.n6539 gnd.n6538 0.152939
R13449 gnd.n6540 gnd.n6539 0.152939
R13450 gnd.n6540 gnd.n388 0.152939
R13451 gnd.n6548 gnd.n388 0.152939
R13452 gnd.n6549 gnd.n6548 0.152939
R13453 gnd.n6550 gnd.n6549 0.152939
R13454 gnd.n6550 gnd.n382 0.152939
R13455 gnd.n6558 gnd.n382 0.152939
R13456 gnd.n6559 gnd.n6558 0.152939
R13457 gnd.n6560 gnd.n6559 0.152939
R13458 gnd.n6560 gnd.n376 0.152939
R13459 gnd.n6568 gnd.n376 0.152939
R13460 gnd.n6569 gnd.n6568 0.152939
R13461 gnd.n6570 gnd.n6569 0.152939
R13462 gnd.n6570 gnd.n370 0.152939
R13463 gnd.n6578 gnd.n370 0.152939
R13464 gnd.n6579 gnd.n6578 0.152939
R13465 gnd.n6580 gnd.n6579 0.152939
R13466 gnd.n6580 gnd.n364 0.152939
R13467 gnd.n6588 gnd.n364 0.152939
R13468 gnd.n6589 gnd.n6588 0.152939
R13469 gnd.n6590 gnd.n6589 0.152939
R13470 gnd.n6590 gnd.n358 0.152939
R13471 gnd.n6598 gnd.n358 0.152939
R13472 gnd.n6599 gnd.n6598 0.152939
R13473 gnd.n6600 gnd.n6599 0.152939
R13474 gnd.n6600 gnd.n352 0.152939
R13475 gnd.n6608 gnd.n352 0.152939
R13476 gnd.n6609 gnd.n6608 0.152939
R13477 gnd.n6610 gnd.n6609 0.152939
R13478 gnd.n6610 gnd.n346 0.152939
R13479 gnd.n6618 gnd.n346 0.152939
R13480 gnd.n6619 gnd.n6618 0.152939
R13481 gnd.n6620 gnd.n6619 0.152939
R13482 gnd.n6620 gnd.n340 0.152939
R13483 gnd.n6629 gnd.n340 0.152939
R13484 gnd.n6630 gnd.n6629 0.152939
R13485 gnd.n6631 gnd.n6630 0.152939
R13486 gnd.n6790 gnd.n246 0.152939
R13487 gnd.n6791 gnd.n6790 0.152939
R13488 gnd.n6792 gnd.n6791 0.152939
R13489 gnd.n6792 gnd.n229 0.152939
R13490 gnd.n6806 gnd.n229 0.152939
R13491 gnd.n6807 gnd.n6806 0.152939
R13492 gnd.n6808 gnd.n6807 0.152939
R13493 gnd.n6808 gnd.n216 0.152939
R13494 gnd.n6822 gnd.n216 0.152939
R13495 gnd.n6823 gnd.n6822 0.152939
R13496 gnd.n6824 gnd.n6823 0.152939
R13497 gnd.n6824 gnd.n200 0.152939
R13498 gnd.n6838 gnd.n200 0.152939
R13499 gnd.n6839 gnd.n6838 0.152939
R13500 gnd.n6840 gnd.n6839 0.152939
R13501 gnd.n6840 gnd.n185 0.152939
R13502 gnd.n6929 gnd.n185 0.152939
R13503 gnd.n6930 gnd.n6929 0.152939
R13504 gnd.n6931 gnd.n6930 0.152939
R13505 gnd.n6931 gnd.n107 0.152939
R13506 gnd.n7011 gnd.n107 0.152939
R13507 gnd.n7010 gnd.n108 0.152939
R13508 gnd.n110 gnd.n108 0.152939
R13509 gnd.n114 gnd.n110 0.152939
R13510 gnd.n115 gnd.n114 0.152939
R13511 gnd.n116 gnd.n115 0.152939
R13512 gnd.n117 gnd.n116 0.152939
R13513 gnd.n121 gnd.n117 0.152939
R13514 gnd.n122 gnd.n121 0.152939
R13515 gnd.n123 gnd.n122 0.152939
R13516 gnd.n124 gnd.n123 0.152939
R13517 gnd.n128 gnd.n124 0.152939
R13518 gnd.n129 gnd.n128 0.152939
R13519 gnd.n130 gnd.n129 0.152939
R13520 gnd.n131 gnd.n130 0.152939
R13521 gnd.n135 gnd.n131 0.152939
R13522 gnd.n136 gnd.n135 0.152939
R13523 gnd.n137 gnd.n136 0.152939
R13524 gnd.n138 gnd.n137 0.152939
R13525 gnd.n142 gnd.n138 0.152939
R13526 gnd.n143 gnd.n142 0.152939
R13527 gnd.n144 gnd.n143 0.152939
R13528 gnd.n145 gnd.n144 0.152939
R13529 gnd.n149 gnd.n145 0.152939
R13530 gnd.n150 gnd.n149 0.152939
R13531 gnd.n151 gnd.n150 0.152939
R13532 gnd.n152 gnd.n151 0.152939
R13533 gnd.n156 gnd.n152 0.152939
R13534 gnd.n157 gnd.n156 0.152939
R13535 gnd.n158 gnd.n157 0.152939
R13536 gnd.n159 gnd.n158 0.152939
R13537 gnd.n163 gnd.n159 0.152939
R13538 gnd.n164 gnd.n163 0.152939
R13539 gnd.n165 gnd.n164 0.152939
R13540 gnd.n166 gnd.n165 0.152939
R13541 gnd.n170 gnd.n166 0.152939
R13542 gnd.n171 gnd.n170 0.152939
R13543 gnd.n6941 gnd.n171 0.152939
R13544 gnd.n6941 gnd.n6940 0.152939
R13545 gnd.n3902 gnd.n3894 0.152939
R13546 gnd.n3902 gnd.n3901 0.152939
R13547 gnd.n3901 gnd.n3900 0.152939
R13548 gnd.n3900 gnd.n3895 0.152939
R13549 gnd.n3895 gnd.n1426 0.152939
R13550 gnd.n3941 gnd.n1426 0.152939
R13551 gnd.n3942 gnd.n3941 0.152939
R13552 gnd.n3943 gnd.n3942 0.152939
R13553 gnd.n3943 gnd.n1424 0.152939
R13554 gnd.n3948 gnd.n1424 0.152939
R13555 gnd.n3949 gnd.n3948 0.152939
R13556 gnd.n3950 gnd.n3949 0.152939
R13557 gnd.n3951 gnd.n3950 0.152939
R13558 gnd.n3952 gnd.n3951 0.152939
R13559 gnd.n3952 gnd.n1387 0.152939
R13560 gnd.n3996 gnd.n1387 0.152939
R13561 gnd.n3997 gnd.n3996 0.152939
R13562 gnd.n3998 gnd.n3997 0.152939
R13563 gnd.n3999 gnd.n3998 0.152939
R13564 gnd.n4000 gnd.n3999 0.152939
R13565 gnd.n4001 gnd.n4000 0.152939
R13566 gnd.n4002 gnd.n4001 0.152939
R13567 gnd.n4002 gnd.n296 0.152939
R13568 gnd.n6683 gnd.n296 0.152939
R13569 gnd.n6684 gnd.n6683 0.152939
R13570 gnd.n6685 gnd.n6684 0.152939
R13571 gnd.n6688 gnd.n6687 0.152939
R13572 gnd.n6689 gnd.n6688 0.152939
R13573 gnd.n6690 gnd.n6689 0.152939
R13574 gnd.n6691 gnd.n6690 0.152939
R13575 gnd.n6692 gnd.n6691 0.152939
R13576 gnd.n6693 gnd.n6692 0.152939
R13577 gnd.n6694 gnd.n6693 0.152939
R13578 gnd.n6695 gnd.n6694 0.152939
R13579 gnd.n6696 gnd.n6695 0.152939
R13580 gnd.n6697 gnd.n6696 0.152939
R13581 gnd.n6698 gnd.n6697 0.152939
R13582 gnd.n6699 gnd.n6698 0.152939
R13583 gnd.n6700 gnd.n6699 0.152939
R13584 gnd.n6701 gnd.n6700 0.152939
R13585 gnd.n6702 gnd.n6701 0.152939
R13586 gnd.n6703 gnd.n6702 0.152939
R13587 gnd.n6704 gnd.n6703 0.152939
R13588 gnd.n6705 gnd.n6704 0.152939
R13589 gnd.n6706 gnd.n6705 0.152939
R13590 gnd.n6707 gnd.n6706 0.152939
R13591 gnd.n6708 gnd.n6707 0.152939
R13592 gnd.n6709 gnd.n6708 0.152939
R13593 gnd.n6711 gnd.n6709 0.152939
R13594 gnd.n6711 gnd.n6710 0.152939
R13595 gnd.n6710 gnd.n177 0.152939
R13596 gnd.n6939 gnd.n177 0.152939
R13597 gnd.n3799 gnd.n3798 0.152939
R13598 gnd.n3799 gnd.n3795 0.152939
R13599 gnd.n3807 gnd.n3795 0.152939
R13600 gnd.n3808 gnd.n3807 0.152939
R13601 gnd.n3809 gnd.n3808 0.152939
R13602 gnd.n3809 gnd.n3791 0.152939
R13603 gnd.n3817 gnd.n3791 0.152939
R13604 gnd.n3818 gnd.n3817 0.152939
R13605 gnd.n3819 gnd.n3818 0.152939
R13606 gnd.n3819 gnd.n3787 0.152939
R13607 gnd.n3827 gnd.n3787 0.152939
R13608 gnd.n3828 gnd.n3827 0.152939
R13609 gnd.n3830 gnd.n3828 0.152939
R13610 gnd.n3830 gnd.n3829 0.152939
R13611 gnd.n3829 gnd.n1486 0.152939
R13612 gnd.n3843 gnd.n3842 0.152939
R13613 gnd.n3843 gnd.n1482 0.152939
R13614 gnd.n3851 gnd.n1482 0.152939
R13615 gnd.n3852 gnd.n3851 0.152939
R13616 gnd.n3853 gnd.n3852 0.152939
R13617 gnd.n3853 gnd.n1478 0.152939
R13618 gnd.n3861 gnd.n1478 0.152939
R13619 gnd.n3862 gnd.n3861 0.152939
R13620 gnd.n3863 gnd.n3862 0.152939
R13621 gnd.n3863 gnd.n1474 0.152939
R13622 gnd.n3871 gnd.n1474 0.152939
R13623 gnd.n3872 gnd.n3871 0.152939
R13624 gnd.n3873 gnd.n3872 0.152939
R13625 gnd.n3873 gnd.n1470 0.152939
R13626 gnd.n3881 gnd.n1470 0.152939
R13627 gnd.n3882 gnd.n3881 0.152939
R13628 gnd.n3884 gnd.n3882 0.152939
R13629 gnd.n3884 gnd.n3883 0.152939
R13630 gnd.n3883 gnd.n1463 0.152939
R13631 gnd.n3893 gnd.n1463 0.152939
R13632 gnd.n1332 gnd.n1331 0.152939
R13633 gnd.n1333 gnd.n1332 0.152939
R13634 gnd.n1434 gnd.n1333 0.152939
R13635 gnd.n3933 gnd.n1434 0.152939
R13636 gnd.n3934 gnd.n3933 0.152939
R13637 gnd.n3935 gnd.n3934 0.152939
R13638 gnd.n3935 gnd.n1404 0.152939
R13639 gnd.n3970 gnd.n1404 0.152939
R13640 gnd.n3971 gnd.n3970 0.152939
R13641 gnd.n3972 gnd.n3971 0.152939
R13642 gnd.n3973 gnd.n3972 0.152939
R13643 gnd.n3973 gnd.n1365 0.152939
R13644 gnd.n4023 gnd.n1365 0.152939
R13645 gnd.n4024 gnd.n4023 0.152939
R13646 gnd.n4025 gnd.n4024 0.152939
R13647 gnd.n4025 gnd.n320 0.152939
R13648 gnd.n6655 gnd.n320 0.152939
R13649 gnd.n6656 gnd.n6655 0.152939
R13650 gnd.n6657 gnd.n6656 0.152939
R13651 gnd.n6658 gnd.n6657 0.152939
R13652 gnd.n6658 gnd.n259 0.152939
R13653 gnd.n6638 gnd.n337 0.152939
R13654 gnd.n6638 gnd.n6637 0.152939
R13655 gnd.n2168 gnd.n2167 0.152939
R13656 gnd.n2169 gnd.n2168 0.152939
R13657 gnd.n2170 gnd.n2169 0.152939
R13658 gnd.n2171 gnd.n2170 0.152939
R13659 gnd.n2172 gnd.n2171 0.152939
R13660 gnd.n2174 gnd.n2172 0.152939
R13661 gnd.n2174 gnd.n2173 0.152939
R13662 gnd.n2173 gnd.n2135 0.152939
R13663 gnd.n2479 gnd.n2135 0.152939
R13664 gnd.n2480 gnd.n2479 0.152939
R13665 gnd.n2481 gnd.n2480 0.152939
R13666 gnd.n2481 gnd.n2131 0.152939
R13667 gnd.n2487 gnd.n2131 0.152939
R13668 gnd.n2488 gnd.n2487 0.152939
R13669 gnd.n2489 gnd.n2488 0.152939
R13670 gnd.n2490 gnd.n2489 0.152939
R13671 gnd.n2491 gnd.n2490 0.152939
R13672 gnd.n2494 gnd.n2491 0.152939
R13673 gnd.n2495 gnd.n2494 0.152939
R13674 gnd.n2496 gnd.n2495 0.152939
R13675 gnd.n2497 gnd.n2496 0.152939
R13676 gnd.n2500 gnd.n2497 0.152939
R13677 gnd.n2501 gnd.n2500 0.152939
R13678 gnd.n2502 gnd.n2501 0.152939
R13679 gnd.n2502 gnd.n1963 0.152939
R13680 gnd.n2841 gnd.n1963 0.152939
R13681 gnd.n2842 gnd.n2841 0.152939
R13682 gnd.n2843 gnd.n2842 0.152939
R13683 gnd.n2843 gnd.n1952 0.152939
R13684 gnd.n2861 gnd.n1952 0.152939
R13685 gnd.n2862 gnd.n2861 0.152939
R13686 gnd.n2863 gnd.n2862 0.152939
R13687 gnd.n2863 gnd.n1939 0.152939
R13688 gnd.n2881 gnd.n1939 0.152939
R13689 gnd.n2882 gnd.n2881 0.152939
R13690 gnd.n2883 gnd.n2882 0.152939
R13691 gnd.n2883 gnd.n1926 0.152939
R13692 gnd.n2901 gnd.n1926 0.152939
R13693 gnd.n2902 gnd.n2901 0.152939
R13694 gnd.n2903 gnd.n2902 0.152939
R13695 gnd.n2903 gnd.n1913 0.152939
R13696 gnd.n2921 gnd.n1913 0.152939
R13697 gnd.n2922 gnd.n2921 0.152939
R13698 gnd.n2923 gnd.n2922 0.152939
R13699 gnd.n2923 gnd.n1898 0.152939
R13700 gnd.n2959 gnd.n1898 0.152939
R13701 gnd.n2960 gnd.n2959 0.152939
R13702 gnd.n2961 gnd.n2960 0.152939
R13703 gnd.n2961 gnd.n1823 0.152939
R13704 gnd.n2986 gnd.n1823 0.152939
R13705 gnd.n2987 gnd.n2986 0.152939
R13706 gnd.n2988 gnd.n2987 0.152939
R13707 gnd.n2989 gnd.n2988 0.152939
R13708 gnd.n2990 gnd.n2989 0.152939
R13709 gnd.n2990 gnd.n1786 0.152939
R13710 gnd.n3047 gnd.n1786 0.152939
R13711 gnd.n3048 gnd.n3047 0.152939
R13712 gnd.n3049 gnd.n3048 0.152939
R13713 gnd.n3049 gnd.n1766 0.152939
R13714 gnd.n3114 gnd.n1766 0.152939
R13715 gnd.n3115 gnd.n3114 0.152939
R13716 gnd.n3116 gnd.n3115 0.152939
R13717 gnd.n3117 gnd.n3116 0.152939
R13718 gnd.n3117 gnd.n1737 0.152939
R13719 gnd.n3150 gnd.n1737 0.152939
R13720 gnd.n3151 gnd.n3150 0.152939
R13721 gnd.n3152 gnd.n3151 0.152939
R13722 gnd.n3152 gnd.n1716 0.152939
R13723 gnd.n3178 gnd.n1716 0.152939
R13724 gnd.n3179 gnd.n3178 0.152939
R13725 gnd.n3180 gnd.n3179 0.152939
R13726 gnd.n3181 gnd.n3180 0.152939
R13727 gnd.n3181 gnd.n1688 0.152939
R13728 gnd.n3217 gnd.n1688 0.152939
R13729 gnd.n3218 gnd.n3217 0.152939
R13730 gnd.n3219 gnd.n3218 0.152939
R13731 gnd.n3220 gnd.n3219 0.152939
R13732 gnd.n3221 gnd.n3220 0.152939
R13733 gnd.n3221 gnd.n1656 0.152939
R13734 gnd.n3284 gnd.n1656 0.152939
R13735 gnd.n3285 gnd.n3284 0.152939
R13736 gnd.n3286 gnd.n3285 0.152939
R13737 gnd.n3286 gnd.n1633 0.152939
R13738 gnd.n3313 gnd.n1633 0.152939
R13739 gnd.n3314 gnd.n3313 0.152939
R13740 gnd.n3315 gnd.n3314 0.152939
R13741 gnd.n3317 gnd.n3315 0.152939
R13742 gnd.n3317 gnd.n3316 0.152939
R13743 gnd.n3316 gnd.n1540 0.152939
R13744 gnd.n1541 gnd.n1540 0.152939
R13745 gnd.n1542 gnd.n1541 0.152939
R13746 gnd.n1552 gnd.n1542 0.152939
R13747 gnd.n1553 gnd.n1552 0.152939
R13748 gnd.n1554 gnd.n1553 0.152939
R13749 gnd.n1555 gnd.n1554 0.152939
R13750 gnd.n1556 gnd.n1555 0.152939
R13751 gnd.n1566 gnd.n1556 0.152939
R13752 gnd.n1567 gnd.n1566 0.152939
R13753 gnd.n1568 gnd.n1567 0.152939
R13754 gnd.n1569 gnd.n1568 0.152939
R13755 gnd.n1576 gnd.n1569 0.152939
R13756 gnd.n1577 gnd.n1576 0.152939
R13757 gnd.n1578 gnd.n1577 0.152939
R13758 gnd.n1579 gnd.n1578 0.152939
R13759 gnd.n1589 gnd.n1579 0.152939
R13760 gnd.n1590 gnd.n1589 0.152939
R13761 gnd.n1591 gnd.n1590 0.152939
R13762 gnd.n1592 gnd.n1591 0.152939
R13763 gnd.n1594 gnd.n1592 0.152939
R13764 gnd.n1594 gnd.n1593 0.152939
R13765 gnd.n1593 gnd.n1310 0.152939
R13766 gnd.n1311 gnd.n1310 0.152939
R13767 gnd.n1312 gnd.n1311 0.152939
R13768 gnd.n1318 gnd.n1312 0.152939
R13769 gnd.n1319 gnd.n1318 0.152939
R13770 gnd.n1320 gnd.n1319 0.152939
R13771 gnd.n1321 gnd.n1320 0.152939
R13772 gnd.n1442 gnd.n1321 0.152939
R13773 gnd.n1443 gnd.n1442 0.152939
R13774 gnd.n1448 gnd.n1443 0.152939
R13775 gnd.n1449 gnd.n1448 0.152939
R13776 gnd.n1450 gnd.n1449 0.152939
R13777 gnd.n1451 gnd.n1450 0.152939
R13778 gnd.n1453 gnd.n1451 0.152939
R13779 gnd.n1453 gnd.n1452 0.152939
R13780 gnd.n1452 gnd.n1414 0.152939
R13781 gnd.n1415 gnd.n1414 0.152939
R13782 gnd.n1416 gnd.n1415 0.152939
R13783 gnd.n1418 gnd.n1416 0.152939
R13784 gnd.n1418 gnd.n1417 0.152939
R13785 gnd.n1417 gnd.n1375 0.152939
R13786 gnd.n1376 gnd.n1375 0.152939
R13787 gnd.n1377 gnd.n1376 0.152939
R13788 gnd.n1380 gnd.n1377 0.152939
R13789 gnd.n1381 gnd.n1380 0.152939
R13790 gnd.n1383 gnd.n1381 0.152939
R13791 gnd.n1383 gnd.n1382 0.152939
R13792 gnd.n1382 gnd.n337 0.152939
R13793 gnd.n1083 gnd.n1082 0.152939
R13794 gnd.n1101 gnd.n1083 0.152939
R13795 gnd.n1102 gnd.n1101 0.152939
R13796 gnd.n1103 gnd.n1102 0.152939
R13797 gnd.n1104 gnd.n1103 0.152939
R13798 gnd.n1122 gnd.n1104 0.152939
R13799 gnd.n1123 gnd.n1122 0.152939
R13800 gnd.n1124 gnd.n1123 0.152939
R13801 gnd.n1125 gnd.n1124 0.152939
R13802 gnd.n1143 gnd.n1125 0.152939
R13803 gnd.n1144 gnd.n1143 0.152939
R13804 gnd.n1145 gnd.n1144 0.152939
R13805 gnd.n1146 gnd.n1145 0.152939
R13806 gnd.n1164 gnd.n1146 0.152939
R13807 gnd.n1165 gnd.n1164 0.152939
R13808 gnd.n1166 gnd.n1165 0.152939
R13809 gnd.n1167 gnd.n1166 0.152939
R13810 gnd.n1186 gnd.n1167 0.152939
R13811 gnd.n1187 gnd.n1186 0.152939
R13812 gnd.n1188 gnd.n1187 0.152939
R13813 gnd.n1189 gnd.n1188 0.152939
R13814 gnd.n2075 gnd.n2074 0.152939
R13815 gnd.n2076 gnd.n2075 0.152939
R13816 gnd.n2077 gnd.n2076 0.152939
R13817 gnd.n2078 gnd.n2077 0.152939
R13818 gnd.n2079 gnd.n2078 0.152939
R13819 gnd.n2080 gnd.n2079 0.152939
R13820 gnd.n2081 gnd.n2080 0.152939
R13821 gnd.n2082 gnd.n2081 0.152939
R13822 gnd.n2083 gnd.n2082 0.152939
R13823 gnd.n2084 gnd.n2083 0.152939
R13824 gnd.n2085 gnd.n2084 0.152939
R13825 gnd.n2086 gnd.n2085 0.152939
R13826 gnd.n2087 gnd.n2086 0.152939
R13827 gnd.n2088 gnd.n2087 0.152939
R13828 gnd.n2089 gnd.n2088 0.152939
R13829 gnd.n2627 gnd.n2626 0.152939
R13830 gnd.n2626 gnd.n2094 0.152939
R13831 gnd.n2095 gnd.n2094 0.152939
R13832 gnd.n2096 gnd.n2095 0.152939
R13833 gnd.n2097 gnd.n2096 0.152939
R13834 gnd.n2098 gnd.n2097 0.152939
R13835 gnd.n2099 gnd.n2098 0.152939
R13836 gnd.n2100 gnd.n2099 0.152939
R13837 gnd.n2101 gnd.n2100 0.152939
R13838 gnd.n2102 gnd.n2101 0.152939
R13839 gnd.n2103 gnd.n2102 0.152939
R13840 gnd.n2104 gnd.n2103 0.152939
R13841 gnd.n2105 gnd.n2104 0.152939
R13842 gnd.n2106 gnd.n2105 0.152939
R13843 gnd.n2107 gnd.n2106 0.152939
R13844 gnd.n2108 gnd.n2107 0.152939
R13845 gnd.n2109 gnd.n2108 0.152939
R13846 gnd.n2110 gnd.n2109 0.152939
R13847 gnd.n2586 gnd.n2110 0.152939
R13848 gnd.n2586 gnd.n2585 0.152939
R13849 gnd.n2298 gnd.n2271 0.152939
R13850 gnd.n2356 gnd.n2271 0.152939
R13851 gnd.n2357 gnd.n2356 0.152939
R13852 gnd.n2358 gnd.n2357 0.152939
R13853 gnd.n2358 gnd.n2269 0.152939
R13854 gnd.n2364 gnd.n2269 0.152939
R13855 gnd.n2365 gnd.n2364 0.152939
R13856 gnd.n2366 gnd.n2365 0.152939
R13857 gnd.n2366 gnd.n2267 0.152939
R13858 gnd.n2372 gnd.n2267 0.152939
R13859 gnd.n2373 gnd.n2372 0.152939
R13860 gnd.n2374 gnd.n2373 0.152939
R13861 gnd.n2374 gnd.n2265 0.152939
R13862 gnd.n2380 gnd.n2265 0.152939
R13863 gnd.n2381 gnd.n2380 0.152939
R13864 gnd.n2382 gnd.n2381 0.152939
R13865 gnd.n2382 gnd.n2263 0.152939
R13866 gnd.n2388 gnd.n2263 0.152939
R13867 gnd.n2389 gnd.n2388 0.152939
R13868 gnd.n2390 gnd.n2389 0.152939
R13869 gnd.n2390 gnd.n2261 0.152939
R13870 gnd.n2396 gnd.n2261 0.152939
R13871 gnd.n2397 gnd.n2396 0.152939
R13872 gnd.n2398 gnd.n2397 0.152939
R13873 gnd.n2398 gnd.n2259 0.152939
R13874 gnd.n2404 gnd.n2259 0.152939
R13875 gnd.n2337 gnd.n2278 0.152939
R13876 gnd.n2279 gnd.n2278 0.152939
R13877 gnd.n2280 gnd.n2279 0.152939
R13878 gnd.n2281 gnd.n2280 0.152939
R13879 gnd.n2282 gnd.n2281 0.152939
R13880 gnd.n2283 gnd.n2282 0.152939
R13881 gnd.n2284 gnd.n2283 0.152939
R13882 gnd.n2285 gnd.n2284 0.152939
R13883 gnd.n2286 gnd.n2285 0.152939
R13884 gnd.n2287 gnd.n2286 0.152939
R13885 gnd.n2288 gnd.n2287 0.152939
R13886 gnd.n2289 gnd.n2288 0.152939
R13887 gnd.n2290 gnd.n2289 0.152939
R13888 gnd.n2291 gnd.n2290 0.152939
R13889 gnd.n2292 gnd.n2291 0.152939
R13890 gnd.n2302 gnd.n2292 0.152939
R13891 gnd.n2302 gnd.n2301 0.152939
R13892 gnd.n2301 gnd.n2300 0.152939
R13893 gnd.n2343 gnd.n2338 0.152939
R13894 gnd.n2343 gnd.n2342 0.152939
R13895 gnd.n2342 gnd.n2341 0.152939
R13896 gnd.n2341 gnd.n2339 0.152939
R13897 gnd.n2339 gnd.n957 0.152939
R13898 gnd.n958 gnd.n957 0.152939
R13899 gnd.n959 gnd.n958 0.152939
R13900 gnd.n975 gnd.n959 0.152939
R13901 gnd.n976 gnd.n975 0.152939
R13902 gnd.n977 gnd.n976 0.152939
R13903 gnd.n978 gnd.n977 0.152939
R13904 gnd.n996 gnd.n978 0.152939
R13905 gnd.n997 gnd.n996 0.152939
R13906 gnd.n998 gnd.n997 0.152939
R13907 gnd.n999 gnd.n998 0.152939
R13908 gnd.n1015 gnd.n999 0.152939
R13909 gnd.n1016 gnd.n1015 0.152939
R13910 gnd.n1017 gnd.n1016 0.152939
R13911 gnd.n1018 gnd.n1017 0.152939
R13912 gnd.n1036 gnd.n1018 0.152939
R13913 gnd.n1037 gnd.n1036 0.152939
R13914 gnd.n1038 gnd.n1037 0.152939
R13915 gnd.n1039 gnd.n1038 0.152939
R13916 gnd.n1053 gnd.n1039 0.152939
R13917 gnd.n1054 gnd.n1053 0.152939
R13918 gnd.n1055 gnd.n1054 0.152939
R13919 gnd.n1071 gnd.n1056 0.152939
R13920 gnd.n1072 gnd.n1071 0.152939
R13921 gnd.n1073 gnd.n1072 0.152939
R13922 gnd.n1074 gnd.n1073 0.152939
R13923 gnd.n1090 gnd.n1074 0.152939
R13924 gnd.n1091 gnd.n1090 0.152939
R13925 gnd.n1092 gnd.n1091 0.152939
R13926 gnd.n1093 gnd.n1092 0.152939
R13927 gnd.n1112 gnd.n1093 0.152939
R13928 gnd.n1113 gnd.n1112 0.152939
R13929 gnd.n1114 gnd.n1113 0.152939
R13930 gnd.n1115 gnd.n1114 0.152939
R13931 gnd.n1132 gnd.n1115 0.152939
R13932 gnd.n1133 gnd.n1132 0.152939
R13933 gnd.n1134 gnd.n1133 0.152939
R13934 gnd.n1135 gnd.n1134 0.152939
R13935 gnd.n1154 gnd.n1135 0.152939
R13936 gnd.n1155 gnd.n1154 0.152939
R13937 gnd.n1156 gnd.n1155 0.152939
R13938 gnd.n1157 gnd.n1156 0.152939
R13939 gnd.n1175 gnd.n1157 0.152939
R13940 gnd.n1176 gnd.n1175 0.152939
R13941 gnd.n1177 gnd.n1176 0.152939
R13942 gnd.n1178 gnd.n1177 0.152939
R13943 gnd.n1196 gnd.n1178 0.152939
R13944 gnd.n4203 gnd.n1196 0.152939
R13945 gnd.n4362 gnd.n932 0.152939
R13946 gnd.n4362 gnd.n4361 0.152939
R13947 gnd.n4361 gnd.n4360 0.152939
R13948 gnd.n4360 gnd.n935 0.152939
R13949 gnd.n2202 gnd.n935 0.152939
R13950 gnd.n2206 gnd.n2202 0.152939
R13951 gnd.n2207 gnd.n2206 0.152939
R13952 gnd.n2208 gnd.n2207 0.152939
R13953 gnd.n2208 gnd.n2200 0.152939
R13954 gnd.n2214 gnd.n2200 0.152939
R13955 gnd.n2215 gnd.n2214 0.152939
R13956 gnd.n2216 gnd.n2215 0.152939
R13957 gnd.n2216 gnd.n2198 0.152939
R13958 gnd.n2222 gnd.n2198 0.152939
R13959 gnd.n2223 gnd.n2222 0.152939
R13960 gnd.n2224 gnd.n2223 0.152939
R13961 gnd.n2224 gnd.n2196 0.152939
R13962 gnd.n2230 gnd.n2196 0.152939
R13963 gnd.n2231 gnd.n2230 0.152939
R13964 gnd.n2232 gnd.n2231 0.152939
R13965 gnd.n2232 gnd.n2194 0.152939
R13966 gnd.n2238 gnd.n2194 0.152939
R13967 gnd.n2239 gnd.n2238 0.152939
R13968 gnd.n2240 gnd.n2239 0.152939
R13969 gnd.n2240 gnd.n2192 0.152939
R13970 gnd.n2246 gnd.n2192 0.152939
R13971 gnd.n2249 gnd.n2248 0.152939
R13972 gnd.n2250 gnd.n2249 0.152939
R13973 gnd.n2251 gnd.n2250 0.152939
R13974 gnd.n2251 gnd.n2185 0.152939
R13975 gnd.n2420 gnd.n2185 0.152939
R13976 gnd.n2421 gnd.n2420 0.152939
R13977 gnd.n2423 gnd.n2421 0.152939
R13978 gnd.n2423 gnd.n2422 0.152939
R13979 gnd.n2422 gnd.n2152 0.152939
R13980 gnd.n2152 gnd.n2150 0.152939
R13981 gnd.n2439 gnd.n2150 0.152939
R13982 gnd.n2440 gnd.n2439 0.152939
R13983 gnd.n2441 gnd.n2440 0.152939
R13984 gnd.n2441 gnd.n2148 0.152939
R13985 gnd.n2450 gnd.n2148 0.152939
R13986 gnd.n2451 gnd.n2450 0.152939
R13987 gnd.n2452 gnd.n2451 0.152939
R13988 gnd.n2453 gnd.n2452 0.152939
R13989 gnd.n2454 gnd.n2453 0.152939
R13990 gnd.n2454 gnd.n2122 0.152939
R13991 gnd.n2530 gnd.n2122 0.152939
R13992 gnd.n2531 gnd.n2530 0.152939
R13993 gnd.n2533 gnd.n2531 0.152939
R13994 gnd.n2533 gnd.n2532 0.152939
R13995 gnd.n2532 gnd.n2115 0.152939
R13996 gnd.n2584 gnd.n2115 0.152939
R13997 gnd.n890 gnd.n889 0.152939
R13998 gnd.n891 gnd.n890 0.152939
R13999 gnd.n892 gnd.n891 0.152939
R14000 gnd.n893 gnd.n892 0.152939
R14001 gnd.n894 gnd.n893 0.152939
R14002 gnd.n895 gnd.n894 0.152939
R14003 gnd.n896 gnd.n895 0.152939
R14004 gnd.n897 gnd.n896 0.152939
R14005 gnd.n898 gnd.n897 0.152939
R14006 gnd.n899 gnd.n898 0.152939
R14007 gnd.n900 gnd.n899 0.152939
R14008 gnd.n901 gnd.n900 0.152939
R14009 gnd.n902 gnd.n901 0.152939
R14010 gnd.n903 gnd.n902 0.152939
R14011 gnd.n904 gnd.n903 0.152939
R14012 gnd.n905 gnd.n904 0.152939
R14013 gnd.n906 gnd.n905 0.152939
R14014 gnd.n909 gnd.n906 0.152939
R14015 gnd.n910 gnd.n909 0.152939
R14016 gnd.n911 gnd.n910 0.152939
R14017 gnd.n912 gnd.n911 0.152939
R14018 gnd.n913 gnd.n912 0.152939
R14019 gnd.n914 gnd.n913 0.152939
R14020 gnd.n915 gnd.n914 0.152939
R14021 gnd.n916 gnd.n915 0.152939
R14022 gnd.n917 gnd.n916 0.152939
R14023 gnd.n918 gnd.n917 0.152939
R14024 gnd.n919 gnd.n918 0.152939
R14025 gnd.n920 gnd.n919 0.152939
R14026 gnd.n921 gnd.n920 0.152939
R14027 gnd.n922 gnd.n921 0.152939
R14028 gnd.n923 gnd.n922 0.152939
R14029 gnd.n924 gnd.n923 0.152939
R14030 gnd.n925 gnd.n924 0.152939
R14031 gnd.n926 gnd.n925 0.152939
R14032 gnd.n4370 gnd.n926 0.152939
R14033 gnd.n4370 gnd.n4369 0.152939
R14034 gnd.n4369 gnd.n4368 0.152939
R14035 gnd.n2349 gnd.n2347 0.152939
R14036 gnd.n2349 gnd.n2348 0.152939
R14037 gnd.n2348 gnd.n946 0.152939
R14038 gnd.n947 gnd.n946 0.152939
R14039 gnd.n948 gnd.n947 0.152939
R14040 gnd.n966 gnd.n948 0.152939
R14041 gnd.n967 gnd.n966 0.152939
R14042 gnd.n968 gnd.n967 0.152939
R14043 gnd.n969 gnd.n968 0.152939
R14044 gnd.n985 gnd.n969 0.152939
R14045 gnd.n986 gnd.n985 0.152939
R14046 gnd.n987 gnd.n986 0.152939
R14047 gnd.n988 gnd.n987 0.152939
R14048 gnd.n1006 gnd.n988 0.152939
R14049 gnd.n1007 gnd.n1006 0.152939
R14050 gnd.n1008 gnd.n1007 0.152939
R14051 gnd.n1009 gnd.n1008 0.152939
R14052 gnd.n1025 gnd.n1009 0.152939
R14053 gnd.n1026 gnd.n1025 0.152939
R14054 gnd.n1027 gnd.n1026 0.152939
R14055 gnd.n1028 gnd.n1027 0.152939
R14056 gnd.n2167 gnd.n2161 0.152939
R14057 gnd.n680 gnd.n675 0.152939
R14058 gnd.n681 gnd.n680 0.152939
R14059 gnd.n682 gnd.n681 0.152939
R14060 gnd.n687 gnd.n682 0.152939
R14061 gnd.n688 gnd.n687 0.152939
R14062 gnd.n689 gnd.n688 0.152939
R14063 gnd.n690 gnd.n689 0.152939
R14064 gnd.n695 gnd.n690 0.152939
R14065 gnd.n696 gnd.n695 0.152939
R14066 gnd.n697 gnd.n696 0.152939
R14067 gnd.n698 gnd.n697 0.152939
R14068 gnd.n703 gnd.n698 0.152939
R14069 gnd.n704 gnd.n703 0.152939
R14070 gnd.n705 gnd.n704 0.152939
R14071 gnd.n706 gnd.n705 0.152939
R14072 gnd.n711 gnd.n706 0.152939
R14073 gnd.n712 gnd.n711 0.152939
R14074 gnd.n713 gnd.n712 0.152939
R14075 gnd.n714 gnd.n713 0.152939
R14076 gnd.n719 gnd.n714 0.152939
R14077 gnd.n720 gnd.n719 0.152939
R14078 gnd.n721 gnd.n720 0.152939
R14079 gnd.n722 gnd.n721 0.152939
R14080 gnd.n727 gnd.n722 0.152939
R14081 gnd.n728 gnd.n727 0.152939
R14082 gnd.n729 gnd.n728 0.152939
R14083 gnd.n730 gnd.n729 0.152939
R14084 gnd.n735 gnd.n730 0.152939
R14085 gnd.n736 gnd.n735 0.152939
R14086 gnd.n737 gnd.n736 0.152939
R14087 gnd.n738 gnd.n737 0.152939
R14088 gnd.n743 gnd.n738 0.152939
R14089 gnd.n744 gnd.n743 0.152939
R14090 gnd.n745 gnd.n744 0.152939
R14091 gnd.n746 gnd.n745 0.152939
R14092 gnd.n751 gnd.n746 0.152939
R14093 gnd.n752 gnd.n751 0.152939
R14094 gnd.n753 gnd.n752 0.152939
R14095 gnd.n754 gnd.n753 0.152939
R14096 gnd.n759 gnd.n754 0.152939
R14097 gnd.n760 gnd.n759 0.152939
R14098 gnd.n761 gnd.n760 0.152939
R14099 gnd.n762 gnd.n761 0.152939
R14100 gnd.n767 gnd.n762 0.152939
R14101 gnd.n768 gnd.n767 0.152939
R14102 gnd.n769 gnd.n768 0.152939
R14103 gnd.n770 gnd.n769 0.152939
R14104 gnd.n775 gnd.n770 0.152939
R14105 gnd.n776 gnd.n775 0.152939
R14106 gnd.n777 gnd.n776 0.152939
R14107 gnd.n778 gnd.n777 0.152939
R14108 gnd.n783 gnd.n778 0.152939
R14109 gnd.n784 gnd.n783 0.152939
R14110 gnd.n785 gnd.n784 0.152939
R14111 gnd.n786 gnd.n785 0.152939
R14112 gnd.n791 gnd.n786 0.152939
R14113 gnd.n792 gnd.n791 0.152939
R14114 gnd.n793 gnd.n792 0.152939
R14115 gnd.n794 gnd.n793 0.152939
R14116 gnd.n799 gnd.n794 0.152939
R14117 gnd.n800 gnd.n799 0.152939
R14118 gnd.n801 gnd.n800 0.152939
R14119 gnd.n802 gnd.n801 0.152939
R14120 gnd.n807 gnd.n802 0.152939
R14121 gnd.n808 gnd.n807 0.152939
R14122 gnd.n809 gnd.n808 0.152939
R14123 gnd.n810 gnd.n809 0.152939
R14124 gnd.n815 gnd.n810 0.152939
R14125 gnd.n816 gnd.n815 0.152939
R14126 gnd.n817 gnd.n816 0.152939
R14127 gnd.n818 gnd.n817 0.152939
R14128 gnd.n823 gnd.n818 0.152939
R14129 gnd.n824 gnd.n823 0.152939
R14130 gnd.n825 gnd.n824 0.152939
R14131 gnd.n826 gnd.n825 0.152939
R14132 gnd.n831 gnd.n826 0.152939
R14133 gnd.n832 gnd.n831 0.152939
R14134 gnd.n833 gnd.n832 0.152939
R14135 gnd.n834 gnd.n833 0.152939
R14136 gnd.n839 gnd.n834 0.152939
R14137 gnd.n840 gnd.n839 0.152939
R14138 gnd.n841 gnd.n840 0.152939
R14139 gnd.n842 gnd.n841 0.152939
R14140 gnd.n2159 gnd.n842 0.152939
R14141 gnd.n3544 gnd.n3400 0.152939
R14142 gnd.n3545 gnd.n3544 0.152939
R14143 gnd.n3546 gnd.n3545 0.152939
R14144 gnd.n3546 gnd.n3396 0.152939
R14145 gnd.n3557 gnd.n3396 0.152939
R14146 gnd.n3558 gnd.n3557 0.152939
R14147 gnd.n3559 gnd.n3558 0.152939
R14148 gnd.n3559 gnd.n3392 0.152939
R14149 gnd.n3566 gnd.n3392 0.152939
R14150 gnd.n2852 gnd.n2851 0.152939
R14151 gnd.n2853 gnd.n2852 0.152939
R14152 gnd.n2853 gnd.n1945 0.152939
R14153 gnd.n2871 gnd.n1945 0.152939
R14154 gnd.n2872 gnd.n2871 0.152939
R14155 gnd.n2873 gnd.n2872 0.152939
R14156 gnd.n2873 gnd.n1932 0.152939
R14157 gnd.n2891 gnd.n1932 0.152939
R14158 gnd.n2892 gnd.n2891 0.152939
R14159 gnd.n2893 gnd.n2892 0.152939
R14160 gnd.n2893 gnd.n1919 0.152939
R14161 gnd.n2911 gnd.n1919 0.152939
R14162 gnd.n2912 gnd.n2911 0.152939
R14163 gnd.n2913 gnd.n2912 0.152939
R14164 gnd.n2913 gnd.n1906 0.152939
R14165 gnd.n2931 gnd.n1906 0.152939
R14166 gnd.n2932 gnd.n2931 0.152939
R14167 gnd.n2951 gnd.n2932 0.152939
R14168 gnd.n2951 gnd.n2950 0.152939
R14169 gnd.n2950 gnd.n2949 0.152939
R14170 gnd.n2949 gnd.n2933 0.152939
R14171 gnd.n2945 gnd.n2933 0.152939
R14172 gnd.n2945 gnd.n2944 0.152939
R14173 gnd.n2944 gnd.n2943 0.152939
R14174 gnd.n2943 gnd.n2938 0.152939
R14175 gnd.n2938 gnd.n1803 0.152939
R14176 gnd.n3015 gnd.n1803 0.152939
R14177 gnd.n3016 gnd.n3015 0.152939
R14178 gnd.n3023 gnd.n3016 0.152939
R14179 gnd.n3023 gnd.n3022 0.152939
R14180 gnd.n3022 gnd.n3021 0.152939
R14181 gnd.n3021 gnd.n3017 0.152939
R14182 gnd.n3017 gnd.n1752 0.152939
R14183 gnd.n3133 gnd.n1752 0.152939
R14184 gnd.n3134 gnd.n3133 0.152939
R14185 gnd.n3136 gnd.n3134 0.152939
R14186 gnd.n3136 gnd.n3135 0.152939
R14187 gnd.n3135 gnd.n1723 0.152939
R14188 gnd.n3169 gnd.n1723 0.152939
R14189 gnd.n3170 gnd.n3169 0.152939
R14190 gnd.n3171 gnd.n3170 0.152939
R14191 gnd.n3171 gnd.n1703 0.152939
R14192 gnd.n3199 gnd.n1703 0.152939
R14193 gnd.n3200 gnd.n3199 0.152939
R14194 gnd.n3202 gnd.n3200 0.152939
R14195 gnd.n3202 gnd.n3201 0.152939
R14196 gnd.n3201 gnd.n1672 0.152939
R14197 gnd.n3242 gnd.n1672 0.152939
R14198 gnd.n3243 gnd.n3242 0.152939
R14199 gnd.n3248 gnd.n3243 0.152939
R14200 gnd.n3248 gnd.n3247 0.152939
R14201 gnd.n3247 gnd.n3246 0.152939
R14202 gnd.n3246 gnd.n1641 0.152939
R14203 gnd.n3302 gnd.n1641 0.152939
R14204 gnd.n3303 gnd.n3302 0.152939
R14205 gnd.n3305 gnd.n3303 0.152939
R14206 gnd.n3305 gnd.n3304 0.152939
R14207 gnd.n3304 gnd.n1615 0.152939
R14208 gnd.n3345 gnd.n1615 0.152939
R14209 gnd.n3346 gnd.n3345 0.152939
R14210 gnd.n3347 gnd.n3346 0.152939
R14211 gnd.n3347 gnd.n1611 0.152939
R14212 gnd.n3355 gnd.n1611 0.152939
R14213 gnd.n3356 gnd.n3355 0.152939
R14214 gnd.n3357 gnd.n3356 0.152939
R14215 gnd.n3357 gnd.n1609 0.152939
R14216 gnd.n3363 gnd.n1609 0.152939
R14217 gnd.n3364 gnd.n3363 0.152939
R14218 gnd.n3365 gnd.n3364 0.152939
R14219 gnd.n3365 gnd.n1607 0.152939
R14220 gnd.n3374 gnd.n1607 0.152939
R14221 gnd.n3375 gnd.n3374 0.152939
R14222 gnd.n3376 gnd.n3375 0.152939
R14223 gnd.n3376 gnd.n1605 0.152939
R14224 gnd.n3382 gnd.n1605 0.152939
R14225 gnd.n3383 gnd.n3382 0.152939
R14226 gnd.n3384 gnd.n3383 0.152939
R14227 gnd.n3384 gnd.n1603 0.152939
R14228 gnd.n3390 gnd.n1603 0.152939
R14229 gnd.n3391 gnd.n3390 0.152939
R14230 gnd.n3568 gnd.n3391 0.152939
R14231 gnd.n3568 gnd.n3567 0.152939
R14232 gnd.n2570 gnd.n2541 0.152939
R14233 gnd.n2570 gnd.n2569 0.152939
R14234 gnd.n2569 gnd.n2568 0.152939
R14235 gnd.n2568 gnd.n2547 0.152939
R14236 gnd.n2564 gnd.n2547 0.152939
R14237 gnd.n2564 gnd.n2563 0.152939
R14238 gnd.n2563 gnd.n2554 0.152939
R14239 gnd.n2559 gnd.n2554 0.152939
R14240 gnd.n2559 gnd.n1958 0.152939
R14241 gnd.n2407 gnd.n2406 0.152939
R14242 gnd.n2407 gnd.n2188 0.152939
R14243 gnd.n2412 gnd.n2188 0.152939
R14244 gnd.n2413 gnd.n2412 0.152939
R14245 gnd.n2414 gnd.n2413 0.152939
R14246 gnd.n2414 gnd.n2154 0.152939
R14247 gnd.n2429 gnd.n2154 0.152939
R14248 gnd.n2430 gnd.n2429 0.152939
R14249 gnd.n2431 gnd.n2430 0.152939
R14250 gnd.n2431 gnd.n2142 0.152939
R14251 gnd.n2470 gnd.n2142 0.152939
R14252 gnd.n2470 gnd.n2469 0.152939
R14253 gnd.n2469 gnd.n2468 0.152939
R14254 gnd.n2468 gnd.n2143 0.152939
R14255 gnd.n2464 gnd.n2143 0.152939
R14256 gnd.n2464 gnd.n2463 0.152939
R14257 gnd.n2463 gnd.n2462 0.152939
R14258 gnd.n2462 gnd.n2125 0.152939
R14259 gnd.n2522 gnd.n2125 0.152939
R14260 gnd.n2523 gnd.n2522 0.152939
R14261 gnd.n2524 gnd.n2523 0.152939
R14262 gnd.n2524 gnd.n2119 0.152939
R14263 gnd.n2539 gnd.n2119 0.152939
R14264 gnd.n2540 gnd.n2539 0.152939
R14265 gnd.n2577 gnd.n2540 0.152939
R14266 gnd.n2577 gnd.n2576 0.152939
R14267 gnd.n4200 gnd.n1199 0.152939
R14268 gnd.n4196 gnd.n1199 0.152939
R14269 gnd.n4196 gnd.n4195 0.152939
R14270 gnd.n4195 gnd.n4194 0.152939
R14271 gnd.n4194 gnd.n1204 0.152939
R14272 gnd.n4190 gnd.n1204 0.152939
R14273 gnd.n4190 gnd.n4189 0.152939
R14274 gnd.n4189 gnd.n4188 0.152939
R14275 gnd.n4188 gnd.n1209 0.152939
R14276 gnd.n4184 gnd.n1209 0.152939
R14277 gnd.n4184 gnd.n4183 0.152939
R14278 gnd.n4183 gnd.n4182 0.152939
R14279 gnd.n4182 gnd.n1214 0.152939
R14280 gnd.n4178 gnd.n1214 0.152939
R14281 gnd.n4178 gnd.n4177 0.152939
R14282 gnd.n4177 gnd.n4176 0.152939
R14283 gnd.n4176 gnd.n1219 0.152939
R14284 gnd.n4172 gnd.n1219 0.152939
R14285 gnd.n4172 gnd.n4171 0.152939
R14286 gnd.n4171 gnd.n4170 0.152939
R14287 gnd.n4170 gnd.n1224 0.152939
R14288 gnd.n4166 gnd.n1224 0.152939
R14289 gnd.n4166 gnd.n4165 0.152939
R14290 gnd.n4165 gnd.n4164 0.152939
R14291 gnd.n4164 gnd.n1229 0.152939
R14292 gnd.n4160 gnd.n1229 0.152939
R14293 gnd.n4160 gnd.n4159 0.152939
R14294 gnd.n4159 gnd.n4158 0.152939
R14295 gnd.n4158 gnd.n1234 0.152939
R14296 gnd.n4154 gnd.n1234 0.152939
R14297 gnd.n4154 gnd.n4153 0.152939
R14298 gnd.n4153 gnd.n4152 0.152939
R14299 gnd.n4152 gnd.n1239 0.152939
R14300 gnd.n4148 gnd.n1239 0.152939
R14301 gnd.n4148 gnd.n4147 0.152939
R14302 gnd.n4147 gnd.n4146 0.152939
R14303 gnd.n4146 gnd.n1244 0.152939
R14304 gnd.n4142 gnd.n1244 0.152939
R14305 gnd.n4142 gnd.n4141 0.152939
R14306 gnd.n4141 gnd.n4140 0.152939
R14307 gnd.n4140 gnd.n1249 0.152939
R14308 gnd.n4136 gnd.n1249 0.152939
R14309 gnd.n4136 gnd.n4135 0.152939
R14310 gnd.n4135 gnd.n4134 0.152939
R14311 gnd.n4134 gnd.n1254 0.152939
R14312 gnd.n4130 gnd.n1254 0.152939
R14313 gnd.n4130 gnd.n4129 0.152939
R14314 gnd.n4129 gnd.n4128 0.152939
R14315 gnd.n4128 gnd.n1259 0.152939
R14316 gnd.n4124 gnd.n1259 0.152939
R14317 gnd.n4124 gnd.n4123 0.152939
R14318 gnd.n4123 gnd.n4122 0.152939
R14319 gnd.n4122 gnd.n1264 0.152939
R14320 gnd.n4118 gnd.n1264 0.152939
R14321 gnd.n4118 gnd.n4117 0.152939
R14322 gnd.n4117 gnd.n4116 0.152939
R14323 gnd.n4116 gnd.n1269 0.152939
R14324 gnd.n4112 gnd.n1269 0.152939
R14325 gnd.n4112 gnd.n4111 0.152939
R14326 gnd.n4111 gnd.n4110 0.152939
R14327 gnd.n4110 gnd.n1274 0.152939
R14328 gnd.n4106 gnd.n1274 0.152939
R14329 gnd.n4106 gnd.n4105 0.152939
R14330 gnd.n4105 gnd.n4104 0.152939
R14331 gnd.n4104 gnd.n1279 0.152939
R14332 gnd.n4100 gnd.n1279 0.152939
R14333 gnd.n4100 gnd.n4099 0.152939
R14334 gnd.n4099 gnd.n4098 0.152939
R14335 gnd.n4098 gnd.n1284 0.152939
R14336 gnd.n4094 gnd.n1284 0.152939
R14337 gnd.n4094 gnd.n4093 0.152939
R14338 gnd.n4093 gnd.n4092 0.152939
R14339 gnd.n4092 gnd.n1289 0.152939
R14340 gnd.n4088 gnd.n1289 0.152939
R14341 gnd.n4088 gnd.n4087 0.152939
R14342 gnd.n4087 gnd.n4086 0.152939
R14343 gnd.n4086 gnd.n1294 0.152939
R14344 gnd.n4082 gnd.n1294 0.152939
R14345 gnd.n4082 gnd.n4081 0.152939
R14346 gnd.n4081 gnd.n4080 0.152939
R14347 gnd.n4080 gnd.n1299 0.152939
R14348 gnd.n1302 gnd.n1299 0.152939
R14349 gnd.n3447 gnd.n1344 0.152939
R14350 gnd.n4050 gnd.n1344 0.152939
R14351 gnd.n4050 gnd.n4049 0.152939
R14352 gnd.n4049 gnd.n4048 0.152939
R14353 gnd.n4048 gnd.n1345 0.152939
R14354 gnd.n4044 gnd.n1345 0.152939
R14355 gnd.n4044 gnd.n4043 0.152939
R14356 gnd.n4043 gnd.n4042 0.152939
R14357 gnd.n4042 gnd.n1350 0.152939
R14358 gnd.n4038 gnd.n1350 0.152939
R14359 gnd.n4038 gnd.n4037 0.152939
R14360 gnd.n4037 gnd.n4036 0.152939
R14361 gnd.n4036 gnd.n1355 0.152939
R14362 gnd.n4032 gnd.n1355 0.152939
R14363 gnd.n4032 gnd.n4031 0.152939
R14364 gnd.n4031 gnd.n330 0.152939
R14365 gnd.n6649 gnd.n330 0.152939
R14366 gnd.n6649 gnd.n6648 0.152939
R14367 gnd.n6648 gnd.n6647 0.152939
R14368 gnd.n6647 gnd.n331 0.152939
R14369 gnd.n331 gnd.n276 0.152939
R14370 gnd.n6769 gnd.n276 0.152939
R14371 gnd.n6769 gnd.n6768 0.152939
R14372 gnd.n6768 gnd.n6767 0.152939
R14373 gnd.n6767 gnd.n277 0.152939
R14374 gnd.n6763 gnd.n277 0.152939
R14375 gnd.n6761 gnd.n6760 0.152939
R14376 gnd.n6760 gnd.n283 0.152939
R14377 gnd.n283 gnd.n253 0.152939
R14378 gnd.n6782 gnd.n253 0.152939
R14379 gnd.n6783 gnd.n6782 0.152939
R14380 gnd.n6784 gnd.n6783 0.152939
R14381 gnd.n6784 gnd.n238 0.152939
R14382 gnd.n6798 gnd.n238 0.152939
R14383 gnd.n6799 gnd.n6798 0.152939
R14384 gnd.n6800 gnd.n6799 0.152939
R14385 gnd.n6800 gnd.n223 0.152939
R14386 gnd.n6814 gnd.n223 0.152939
R14387 gnd.n6815 gnd.n6814 0.152939
R14388 gnd.n6816 gnd.n6815 0.152939
R14389 gnd.n6816 gnd.n208 0.152939
R14390 gnd.n6830 gnd.n208 0.152939
R14391 gnd.n6831 gnd.n6830 0.152939
R14392 gnd.n6832 gnd.n6831 0.152939
R14393 gnd.n6832 gnd.n194 0.152939
R14394 gnd.n6846 gnd.n194 0.152939
R14395 gnd.n6847 gnd.n6846 0.152939
R14396 gnd.n6923 gnd.n6847 0.152939
R14397 gnd.n6923 gnd.n6922 0.152939
R14398 gnd.n6922 gnd.n6921 0.152939
R14399 gnd.n6921 gnd.n6848 0.152939
R14400 gnd.n6917 gnd.n6848 0.152939
R14401 gnd.n6916 gnd.n6850 0.152939
R14402 gnd.n6912 gnd.n6850 0.152939
R14403 gnd.n6912 gnd.n6911 0.152939
R14404 gnd.n6911 gnd.n6910 0.152939
R14405 gnd.n6910 gnd.n6856 0.152939
R14406 gnd.n6906 gnd.n6856 0.152939
R14407 gnd.n6906 gnd.n6905 0.152939
R14408 gnd.n6905 gnd.n6904 0.152939
R14409 gnd.n6904 gnd.n6864 0.152939
R14410 gnd.n6900 gnd.n6864 0.152939
R14411 gnd.n6900 gnd.n6899 0.152939
R14412 gnd.n6899 gnd.n6898 0.152939
R14413 gnd.n6898 gnd.n6872 0.152939
R14414 gnd.n6894 gnd.n6872 0.152939
R14415 gnd.n6894 gnd.n6893 0.152939
R14416 gnd.n6893 gnd.n6892 0.152939
R14417 gnd.n6892 gnd.n6880 0.152939
R14418 gnd.n6888 gnd.n6880 0.152939
R14419 gnd.n3908 gnd.n1459 0.152939
R14420 gnd.n3909 gnd.n3908 0.152939
R14421 gnd.n3910 gnd.n3909 0.152939
R14422 gnd.n3910 gnd.n1456 0.152939
R14423 gnd.n3915 gnd.n1456 0.152939
R14424 gnd.n3916 gnd.n3915 0.152939
R14425 gnd.n3918 gnd.n3916 0.152939
R14426 gnd.n3918 gnd.n3917 0.152939
R14427 gnd.n3917 gnd.n1394 0.152939
R14428 gnd.n3980 gnd.n1394 0.152939
R14429 gnd.n3981 gnd.n3980 0.152939
R14430 gnd.n3982 gnd.n3981 0.152939
R14431 gnd.n3982 gnd.n1391 0.152939
R14432 gnd.n3987 gnd.n1391 0.152939
R14433 gnd.n3988 gnd.n3987 0.152939
R14434 gnd.n3990 gnd.n3988 0.152939
R14435 gnd.n3990 gnd.n3989 0.152939
R14436 gnd.n3989 gnd.n309 0.152939
R14437 gnd.n6665 gnd.n309 0.152939
R14438 gnd.n6666 gnd.n6665 0.152939
R14439 gnd.n6667 gnd.n6666 0.152939
R14440 gnd.n6667 gnd.n306 0.152939
R14441 gnd.n6672 gnd.n306 0.152939
R14442 gnd.n6673 gnd.n6672 0.152939
R14443 gnd.n6674 gnd.n6673 0.152939
R14444 gnd.n6674 gnd.n63 0.152939
R14445 gnd.n7055 gnd.n64 0.152939
R14446 gnd.n7051 gnd.n64 0.152939
R14447 gnd.n7051 gnd.n7050 0.152939
R14448 gnd.n7050 gnd.n7049 0.152939
R14449 gnd.n7049 gnd.n70 0.152939
R14450 gnd.n7045 gnd.n70 0.152939
R14451 gnd.n7045 gnd.n7044 0.152939
R14452 gnd.n7044 gnd.n7043 0.152939
R14453 gnd.n7043 gnd.n75 0.152939
R14454 gnd.n7039 gnd.n75 0.152939
R14455 gnd.n7039 gnd.n7038 0.152939
R14456 gnd.n7038 gnd.n7037 0.152939
R14457 gnd.n7037 gnd.n80 0.152939
R14458 gnd.n7033 gnd.n80 0.152939
R14459 gnd.n7033 gnd.n7032 0.152939
R14460 gnd.n7032 gnd.n7031 0.152939
R14461 gnd.n7031 gnd.n85 0.152939
R14462 gnd.n7027 gnd.n85 0.152939
R14463 gnd.n7027 gnd.n7026 0.152939
R14464 gnd.n7026 gnd.n7025 0.152939
R14465 gnd.n7025 gnd.n90 0.152939
R14466 gnd.n7021 gnd.n90 0.152939
R14467 gnd.n7021 gnd.n7020 0.152939
R14468 gnd.n7020 gnd.n7019 0.152939
R14469 gnd.n7019 gnd.n95 0.152939
R14470 gnd.n98 gnd.n95 0.152939
R14471 gnd.n3535 gnd.n3400 0.151415
R14472 gnd.n2575 gnd.n2541 0.151415
R14473 gnd.n5341 gnd.n5257 0.0767195
R14474 gnd.n5341 gnd.n5255 0.0767195
R14475 gnd.n6776 gnd.n246 0.0767195
R14476 gnd.n6685 gnd.n282 0.0767195
R14477 gnd.n6687 gnd.n282 0.0767195
R14478 gnd.n6776 gnd.n259 0.0767195
R14479 gnd.n1082 gnd.n1047 0.0767195
R14480 gnd.n2191 gnd.n1055 0.0767195
R14481 gnd.n2191 gnd.n1056 0.0767195
R14482 gnd.n2247 gnd.n2246 0.0767195
R14483 gnd.n2248 gnd.n2247 0.0767195
R14484 gnd.n1047 gnd.n1028 0.0767195
R14485 gnd.n6763 gnd.n6762 0.0767195
R14486 gnd.n6762 gnd.n6761 0.0767195
R14487 gnd.n7056 gnd.n63 0.0767195
R14488 gnd.n7056 gnd.n7055 0.0767195
R14489 gnd.n2405 gnd.n2404 0.0695946
R14490 gnd.n2406 gnd.n2405 0.0695946
R14491 gnd.n4202 gnd.n4201 0.063
R14492 gnd.n3448 gnd.n3445 0.063
R14493 gnd.n6637 gnd.n260 0.0569024
R14494 gnd.n2161 gnd.n2160 0.0569024
R14495 gnd.n5852 gnd.n4479 0.0477147
R14496 gnd.n5197 gnd.n5093 0.0442063
R14497 gnd.n5211 gnd.n5093 0.0442063
R14498 gnd.n5212 gnd.n5211 0.0442063
R14499 gnd.n5213 gnd.n5212 0.0442063
R14500 gnd.n5213 gnd.n5081 0.0442063
R14501 gnd.n5227 gnd.n5081 0.0442063
R14502 gnd.n5228 gnd.n5227 0.0442063
R14503 gnd.n5229 gnd.n5228 0.0442063
R14504 gnd.n5229 gnd.n5068 0.0442063
R14505 gnd.n5438 gnd.n5068 0.0442063
R14506 gnd.n5441 gnd.n5440 0.0344674
R14507 gnd.n3536 gnd.n3534 0.0344674
R14508 gnd.n2574 gnd.n2033 0.0344674
R14509 gnd.n5061 gnd.n5060 0.0269946
R14510 gnd.n5451 gnd.n5449 0.0269946
R14511 gnd.n5450 gnd.n5043 0.0269946
R14512 gnd.n5470 gnd.n5469 0.0269946
R14513 gnd.n5472 gnd.n5471 0.0269946
R14514 gnd.n5037 gnd.n5035 0.0269946
R14515 gnd.n5482 gnd.n5480 0.0269946
R14516 gnd.n5481 gnd.n5016 0.0269946
R14517 gnd.n5501 gnd.n5500 0.0269946
R14518 gnd.n5503 gnd.n5502 0.0269946
R14519 gnd.n5011 gnd.n5009 0.0269946
R14520 gnd.n5513 gnd.n5511 0.0269946
R14521 gnd.n5512 gnd.n4990 0.0269946
R14522 gnd.n5532 gnd.n5531 0.0269946
R14523 gnd.n5534 gnd.n5533 0.0269946
R14524 gnd.n4985 gnd.n4983 0.0269946
R14525 gnd.n5544 gnd.n5542 0.0269946
R14526 gnd.n5543 gnd.n4965 0.0269946
R14527 gnd.n5563 gnd.n5562 0.0269946
R14528 gnd.n5565 gnd.n5564 0.0269946
R14529 gnd.n4959 gnd.n4957 0.0269946
R14530 gnd.n5575 gnd.n5573 0.0269946
R14531 gnd.n5574 gnd.n4940 0.0269946
R14532 gnd.n5594 gnd.n5593 0.0269946
R14533 gnd.n5596 gnd.n5595 0.0269946
R14534 gnd.n4934 gnd.n4932 0.0269946
R14535 gnd.n5606 gnd.n5604 0.0269946
R14536 gnd.n5605 gnd.n4915 0.0269946
R14537 gnd.n5625 gnd.n5624 0.0269946
R14538 gnd.n5627 gnd.n5626 0.0269946
R14539 gnd.n4909 gnd.n4907 0.0269946
R14540 gnd.n5637 gnd.n5635 0.0269946
R14541 gnd.n5636 gnd.n4891 0.0269946
R14542 gnd.n5655 gnd.n5654 0.0269946
R14543 gnd.n5657 gnd.n5656 0.0269946
R14544 gnd.n4879 gnd.n4878 0.0269946
R14545 gnd.n5678 gnd.n4874 0.0269946
R14546 gnd.n5677 gnd.n4876 0.0269946
R14547 gnd.n4875 gnd.n4856 0.0269946
R14548 gnd.n5701 gnd.n4857 0.0269946
R14549 gnd.n5700 gnd.n4858 0.0269946
R14550 gnd.n5720 gnd.n4842 0.0269946
R14551 gnd.n5722 gnd.n5721 0.0269946
R14552 gnd.n5723 gnd.n4827 0.0269946
R14553 gnd.n5746 gnd.n4828 0.0269946
R14554 gnd.n5745 gnd.n4829 0.0269946
R14555 gnd.n5765 gnd.n4815 0.0269946
R14556 gnd.n5768 gnd.n5767 0.0269946
R14557 gnd.n5787 gnd.n4793 0.0269946
R14558 gnd.n4795 gnd.n850 0.0269946
R14559 gnd.n4799 gnd.n851 0.0269946
R14560 gnd.n4800 gnd.n852 0.0269946
R14561 gnd.n3445 gnd.n3444 0.0246168
R14562 gnd.n4201 gnd.n1198 0.0246168
R14563 gnd.n5440 gnd.n5439 0.0202011
R14564 gnd.n3444 gnd.n3442 0.0174837
R14565 gnd.n3456 gnd.n3442 0.0174837
R14566 gnd.n3458 gnd.n3456 0.0174837
R14567 gnd.n3458 gnd.n3457 0.0174837
R14568 gnd.n3457 gnd.n3437 0.0174837
R14569 gnd.n3467 gnd.n3437 0.0174837
R14570 gnd.n3467 gnd.n3466 0.0174837
R14571 gnd.n3466 gnd.n3438 0.0174837
R14572 gnd.n3438 gnd.n3433 0.0174837
R14573 gnd.n3475 gnd.n3433 0.0174837
R14574 gnd.n3477 gnd.n3475 0.0174837
R14575 gnd.n3477 gnd.n3476 0.0174837
R14576 gnd.n3476 gnd.n3428 0.0174837
R14577 gnd.n3486 gnd.n3428 0.0174837
R14578 gnd.n3486 gnd.n3485 0.0174837
R14579 gnd.n3485 gnd.n3429 0.0174837
R14580 gnd.n3429 gnd.n3424 0.0174837
R14581 gnd.n3494 gnd.n3424 0.0174837
R14582 gnd.n3496 gnd.n3494 0.0174837
R14583 gnd.n3496 gnd.n3495 0.0174837
R14584 gnd.n3495 gnd.n3419 0.0174837
R14585 gnd.n3505 gnd.n3419 0.0174837
R14586 gnd.n3505 gnd.n3504 0.0174837
R14587 gnd.n3504 gnd.n3420 0.0174837
R14588 gnd.n3420 gnd.n3415 0.0174837
R14589 gnd.n3513 gnd.n3415 0.0174837
R14590 gnd.n3515 gnd.n3513 0.0174837
R14591 gnd.n3515 gnd.n3514 0.0174837
R14592 gnd.n3514 gnd.n3410 0.0174837
R14593 gnd.n3526 gnd.n3410 0.0174837
R14594 gnd.n3526 gnd.n3525 0.0174837
R14595 gnd.n3525 gnd.n3411 0.0174837
R14596 gnd.n3411 gnd.n3404 0.0174837
R14597 gnd.n3533 gnd.n3404 0.0174837
R14598 gnd.n3534 gnd.n3533 0.0174837
R14599 gnd.n1982 gnd.n1198 0.0174837
R14600 gnd.n1984 gnd.n1982 0.0174837
R14601 gnd.n2832 gnd.n1984 0.0174837
R14602 gnd.n2832 gnd.n2831 0.0174837
R14603 gnd.n2831 gnd.n1985 0.0174837
R14604 gnd.n2828 gnd.n1985 0.0174837
R14605 gnd.n2828 gnd.n2827 0.0174837
R14606 gnd.n2827 gnd.n1990 0.0174837
R14607 gnd.n2824 gnd.n1990 0.0174837
R14608 gnd.n2824 gnd.n2823 0.0174837
R14609 gnd.n2823 gnd.n1995 0.0174837
R14610 gnd.n2820 gnd.n1995 0.0174837
R14611 gnd.n2820 gnd.n2819 0.0174837
R14612 gnd.n2819 gnd.n1999 0.0174837
R14613 gnd.n2816 gnd.n1999 0.0174837
R14614 gnd.n2816 gnd.n2815 0.0174837
R14615 gnd.n2815 gnd.n2003 0.0174837
R14616 gnd.n2812 gnd.n2003 0.0174837
R14617 gnd.n2812 gnd.n2811 0.0174837
R14618 gnd.n2811 gnd.n2007 0.0174837
R14619 gnd.n2808 gnd.n2007 0.0174837
R14620 gnd.n2808 gnd.n2807 0.0174837
R14621 gnd.n2807 gnd.n2013 0.0174837
R14622 gnd.n2804 gnd.n2013 0.0174837
R14623 gnd.n2804 gnd.n2803 0.0174837
R14624 gnd.n2803 gnd.n2017 0.0174837
R14625 gnd.n2800 gnd.n2017 0.0174837
R14626 gnd.n2800 gnd.n2799 0.0174837
R14627 gnd.n2799 gnd.n2021 0.0174837
R14628 gnd.n2796 gnd.n2021 0.0174837
R14629 gnd.n2796 gnd.n2795 0.0174837
R14630 gnd.n2795 gnd.n2027 0.0174837
R14631 gnd.n2792 gnd.n2027 0.0174837
R14632 gnd.n2792 gnd.n2791 0.0174837
R14633 gnd.n2791 gnd.n2033 0.0174837
R14634 gnd.n5439 gnd.n5438 0.0148637
R14635 gnd.n5766 gnd.n4792 0.0144266
R14636 gnd.n5788 gnd.n4792 0.0130679
R14637 gnd.n5441 gnd.n5061 0.00797283
R14638 gnd.n5449 gnd.n5060 0.00797283
R14639 gnd.n5451 gnd.n5450 0.00797283
R14640 gnd.n5469 gnd.n5043 0.00797283
R14641 gnd.n5471 gnd.n5470 0.00797283
R14642 gnd.n5472 gnd.n5037 0.00797283
R14643 gnd.n5480 gnd.n5035 0.00797283
R14644 gnd.n5482 gnd.n5481 0.00797283
R14645 gnd.n5500 gnd.n5016 0.00797283
R14646 gnd.n5502 gnd.n5501 0.00797283
R14647 gnd.n5503 gnd.n5011 0.00797283
R14648 gnd.n5511 gnd.n5009 0.00797283
R14649 gnd.n5513 gnd.n5512 0.00797283
R14650 gnd.n5531 gnd.n4990 0.00797283
R14651 gnd.n5533 gnd.n5532 0.00797283
R14652 gnd.n5534 gnd.n4985 0.00797283
R14653 gnd.n5542 gnd.n4983 0.00797283
R14654 gnd.n5544 gnd.n5543 0.00797283
R14655 gnd.n5562 gnd.n4965 0.00797283
R14656 gnd.n5564 gnd.n5563 0.00797283
R14657 gnd.n5565 gnd.n4959 0.00797283
R14658 gnd.n5573 gnd.n4957 0.00797283
R14659 gnd.n5575 gnd.n5574 0.00797283
R14660 gnd.n5593 gnd.n4940 0.00797283
R14661 gnd.n5595 gnd.n5594 0.00797283
R14662 gnd.n5596 gnd.n4934 0.00797283
R14663 gnd.n5604 gnd.n4932 0.00797283
R14664 gnd.n5606 gnd.n5605 0.00797283
R14665 gnd.n5624 gnd.n4915 0.00797283
R14666 gnd.n5626 gnd.n5625 0.00797283
R14667 gnd.n5627 gnd.n4909 0.00797283
R14668 gnd.n5635 gnd.n4907 0.00797283
R14669 gnd.n5637 gnd.n5636 0.00797283
R14670 gnd.n5654 gnd.n4891 0.00797283
R14671 gnd.n5656 gnd.n5655 0.00797283
R14672 gnd.n5657 gnd.n4879 0.00797283
R14673 gnd.n4878 gnd.n4874 0.00797283
R14674 gnd.n5678 gnd.n5677 0.00797283
R14675 gnd.n4876 gnd.n4875 0.00797283
R14676 gnd.n4857 gnd.n4856 0.00797283
R14677 gnd.n5701 gnd.n5700 0.00797283
R14678 gnd.n4858 gnd.n4842 0.00797283
R14679 gnd.n5721 gnd.n5720 0.00797283
R14680 gnd.n5723 gnd.n5722 0.00797283
R14681 gnd.n4828 gnd.n4827 0.00797283
R14682 gnd.n5746 gnd.n5745 0.00797283
R14683 gnd.n4829 gnd.n4815 0.00797283
R14684 gnd.n5768 gnd.n5765 0.00797283
R14685 gnd.n5767 gnd.n5766 0.00797283
R14686 gnd.n5788 gnd.n5787 0.00797283
R14687 gnd.n4795 gnd.n4793 0.00797283
R14688 gnd.n4799 gnd.n850 0.00797283
R14689 gnd.n4800 gnd.n851 0.00797283
R14690 gnd.n4479 gnd.n852 0.00797283
R14691 gnd.n6762 gnd.n282 0.00507153
R14692 gnd.n2247 gnd.n2191 0.00507153
R14693 gnd.n3536 gnd.n3535 0.000839674
R14694 gnd.n2575 gnd.n2574 0.000839674
R14695 vdd.n303 vdd.n267 756.745
R14696 vdd.n252 vdd.n216 756.745
R14697 vdd.n209 vdd.n173 756.745
R14698 vdd.n158 vdd.n122 756.745
R14699 vdd.n116 vdd.n80 756.745
R14700 vdd.n65 vdd.n29 756.745
R14701 vdd.n1498 vdd.n1462 756.745
R14702 vdd.n1549 vdd.n1513 756.745
R14703 vdd.n1404 vdd.n1368 756.745
R14704 vdd.n1455 vdd.n1419 756.745
R14705 vdd.n1311 vdd.n1275 756.745
R14706 vdd.n1362 vdd.n1326 756.745
R14707 vdd.n1889 vdd.t119 640.208
R14708 vdd.n793 vdd.t104 640.208
R14709 vdd.n1863 vdd.t146 640.208
R14710 vdd.n785 vdd.t130 640.208
R14711 vdd.n2634 vdd.t91 640.208
R14712 vdd.n2354 vdd.t127 640.208
R14713 vdd.n661 vdd.t108 640.208
R14714 vdd.n2351 vdd.t112 640.208
R14715 vdd.n625 vdd.t116 640.208
R14716 vdd.n855 vdd.t123 640.208
R14717 vdd.n1110 vdd.t140 592.009
R14718 vdd.n1147 vdd.t87 592.009
R14719 vdd.n1021 vdd.t98 592.009
R14720 vdd.n2045 vdd.t83 592.009
R14721 vdd.n1682 vdd.t95 592.009
R14722 vdd.n1642 vdd.t101 592.009
R14723 vdd.n3021 vdd.t143 592.009
R14724 vdd.n427 vdd.t136 592.009
R14725 vdd.n387 vdd.t149 592.009
R14726 vdd.n580 vdd.t76 592.009
R14727 vdd.n543 vdd.t80 592.009
R14728 vdd.n2808 vdd.t133 592.009
R14729 vdd.n304 vdd.n303 585
R14730 vdd.n302 vdd.n269 585
R14731 vdd.n301 vdd.n300 585
R14732 vdd.n272 vdd.n270 585
R14733 vdd.n295 vdd.n294 585
R14734 vdd.n293 vdd.n292 585
R14735 vdd.n276 vdd.n275 585
R14736 vdd.n287 vdd.n286 585
R14737 vdd.n285 vdd.n284 585
R14738 vdd.n280 vdd.n279 585
R14739 vdd.n253 vdd.n252 585
R14740 vdd.n251 vdd.n218 585
R14741 vdd.n250 vdd.n249 585
R14742 vdd.n221 vdd.n219 585
R14743 vdd.n244 vdd.n243 585
R14744 vdd.n242 vdd.n241 585
R14745 vdd.n225 vdd.n224 585
R14746 vdd.n236 vdd.n235 585
R14747 vdd.n234 vdd.n233 585
R14748 vdd.n229 vdd.n228 585
R14749 vdd.n210 vdd.n209 585
R14750 vdd.n208 vdd.n175 585
R14751 vdd.n207 vdd.n206 585
R14752 vdd.n178 vdd.n176 585
R14753 vdd.n201 vdd.n200 585
R14754 vdd.n199 vdd.n198 585
R14755 vdd.n182 vdd.n181 585
R14756 vdd.n193 vdd.n192 585
R14757 vdd.n191 vdd.n190 585
R14758 vdd.n186 vdd.n185 585
R14759 vdd.n159 vdd.n158 585
R14760 vdd.n157 vdd.n124 585
R14761 vdd.n156 vdd.n155 585
R14762 vdd.n127 vdd.n125 585
R14763 vdd.n150 vdd.n149 585
R14764 vdd.n148 vdd.n147 585
R14765 vdd.n131 vdd.n130 585
R14766 vdd.n142 vdd.n141 585
R14767 vdd.n140 vdd.n139 585
R14768 vdd.n135 vdd.n134 585
R14769 vdd.n117 vdd.n116 585
R14770 vdd.n115 vdd.n82 585
R14771 vdd.n114 vdd.n113 585
R14772 vdd.n85 vdd.n83 585
R14773 vdd.n108 vdd.n107 585
R14774 vdd.n106 vdd.n105 585
R14775 vdd.n89 vdd.n88 585
R14776 vdd.n100 vdd.n99 585
R14777 vdd.n98 vdd.n97 585
R14778 vdd.n93 vdd.n92 585
R14779 vdd.n66 vdd.n65 585
R14780 vdd.n64 vdd.n31 585
R14781 vdd.n63 vdd.n62 585
R14782 vdd.n34 vdd.n32 585
R14783 vdd.n57 vdd.n56 585
R14784 vdd.n55 vdd.n54 585
R14785 vdd.n38 vdd.n37 585
R14786 vdd.n49 vdd.n48 585
R14787 vdd.n47 vdd.n46 585
R14788 vdd.n42 vdd.n41 585
R14789 vdd.n1499 vdd.n1498 585
R14790 vdd.n1497 vdd.n1464 585
R14791 vdd.n1496 vdd.n1495 585
R14792 vdd.n1467 vdd.n1465 585
R14793 vdd.n1490 vdd.n1489 585
R14794 vdd.n1488 vdd.n1487 585
R14795 vdd.n1471 vdd.n1470 585
R14796 vdd.n1482 vdd.n1481 585
R14797 vdd.n1480 vdd.n1479 585
R14798 vdd.n1475 vdd.n1474 585
R14799 vdd.n1550 vdd.n1549 585
R14800 vdd.n1548 vdd.n1515 585
R14801 vdd.n1547 vdd.n1546 585
R14802 vdd.n1518 vdd.n1516 585
R14803 vdd.n1541 vdd.n1540 585
R14804 vdd.n1539 vdd.n1538 585
R14805 vdd.n1522 vdd.n1521 585
R14806 vdd.n1533 vdd.n1532 585
R14807 vdd.n1531 vdd.n1530 585
R14808 vdd.n1526 vdd.n1525 585
R14809 vdd.n1405 vdd.n1404 585
R14810 vdd.n1403 vdd.n1370 585
R14811 vdd.n1402 vdd.n1401 585
R14812 vdd.n1373 vdd.n1371 585
R14813 vdd.n1396 vdd.n1395 585
R14814 vdd.n1394 vdd.n1393 585
R14815 vdd.n1377 vdd.n1376 585
R14816 vdd.n1388 vdd.n1387 585
R14817 vdd.n1386 vdd.n1385 585
R14818 vdd.n1381 vdd.n1380 585
R14819 vdd.n1456 vdd.n1455 585
R14820 vdd.n1454 vdd.n1421 585
R14821 vdd.n1453 vdd.n1452 585
R14822 vdd.n1424 vdd.n1422 585
R14823 vdd.n1447 vdd.n1446 585
R14824 vdd.n1445 vdd.n1444 585
R14825 vdd.n1428 vdd.n1427 585
R14826 vdd.n1439 vdd.n1438 585
R14827 vdd.n1437 vdd.n1436 585
R14828 vdd.n1432 vdd.n1431 585
R14829 vdd.n1312 vdd.n1311 585
R14830 vdd.n1310 vdd.n1277 585
R14831 vdd.n1309 vdd.n1308 585
R14832 vdd.n1280 vdd.n1278 585
R14833 vdd.n1303 vdd.n1302 585
R14834 vdd.n1301 vdd.n1300 585
R14835 vdd.n1284 vdd.n1283 585
R14836 vdd.n1295 vdd.n1294 585
R14837 vdd.n1293 vdd.n1292 585
R14838 vdd.n1288 vdd.n1287 585
R14839 vdd.n1363 vdd.n1362 585
R14840 vdd.n1361 vdd.n1328 585
R14841 vdd.n1360 vdd.n1359 585
R14842 vdd.n1331 vdd.n1329 585
R14843 vdd.n1354 vdd.n1353 585
R14844 vdd.n1352 vdd.n1351 585
R14845 vdd.n1335 vdd.n1334 585
R14846 vdd.n1346 vdd.n1345 585
R14847 vdd.n1344 vdd.n1343 585
R14848 vdd.n1339 vdd.n1338 585
R14849 vdd.n3137 vdd.n352 488.781
R14850 vdd.n3019 vdd.n350 488.781
R14851 vdd.n2941 vdd.n515 488.781
R14852 vdd.n2939 vdd.n517 488.781
R14853 vdd.n2040 vdd.n903 488.781
R14854 vdd.n2043 vdd.n2042 488.781
R14855 vdd.n1216 vdd.n981 488.781
R14856 vdd.n1214 vdd.n984 488.781
R14857 vdd.n281 vdd.t207 329.043
R14858 vdd.n230 vdd.t42 329.043
R14859 vdd.n187 vdd.t11 329.043
R14860 vdd.n136 vdd.t72 329.043
R14861 vdd.n94 vdd.t38 329.043
R14862 vdd.n43 vdd.t16 329.043
R14863 vdd.n1476 vdd.t208 329.043
R14864 vdd.n1527 vdd.t200 329.043
R14865 vdd.n1382 vdd.t54 329.043
R14866 vdd.n1433 vdd.t188 329.043
R14867 vdd.n1289 vdd.t18 329.043
R14868 vdd.n1340 vdd.t63 329.043
R14869 vdd.n1110 vdd.t142 319.788
R14870 vdd.n1147 vdd.t90 319.788
R14871 vdd.n1021 vdd.t100 319.788
R14872 vdd.n2045 vdd.t85 319.788
R14873 vdd.n1682 vdd.t96 319.788
R14874 vdd.n1642 vdd.t102 319.788
R14875 vdd.n3021 vdd.t144 319.788
R14876 vdd.n427 vdd.t138 319.788
R14877 vdd.n387 vdd.t150 319.788
R14878 vdd.n580 vdd.t79 319.788
R14879 vdd.n543 vdd.t82 319.788
R14880 vdd.n2808 vdd.t135 319.788
R14881 vdd.n1111 vdd.t141 303.69
R14882 vdd.n1148 vdd.t89 303.69
R14883 vdd.n1022 vdd.t99 303.69
R14884 vdd.n2046 vdd.t86 303.69
R14885 vdd.n1683 vdd.t97 303.69
R14886 vdd.n1643 vdd.t103 303.69
R14887 vdd.n3022 vdd.t145 303.69
R14888 vdd.n428 vdd.t139 303.69
R14889 vdd.n388 vdd.t151 303.69
R14890 vdd.n581 vdd.t78 303.69
R14891 vdd.n544 vdd.t81 303.69
R14892 vdd.n2809 vdd.t134 303.69
R14893 vdd.n2577 vdd.n741 297.074
R14894 vdd.n2770 vdd.n635 297.074
R14895 vdd.n2707 vdd.n632 297.074
R14896 vdd.n2500 vdd.n742 297.074
R14897 vdd.n2315 vdd.n782 297.074
R14898 vdd.n2246 vdd.n2245 297.074
R14899 vdd.n1992 vdd.n878 297.074
R14900 vdd.n2088 vdd.n876 297.074
R14901 vdd.n2686 vdd.n633 297.074
R14902 vdd.n2773 vdd.n2772 297.074
R14903 vdd.n2349 vdd.n743 297.074
R14904 vdd.n2575 vdd.n744 297.074
R14905 vdd.n2243 vdd.n791 297.074
R14906 vdd.n789 vdd.n764 297.074
R14907 vdd.n1929 vdd.n879 297.074
R14908 vdd.n2086 vdd.n880 297.074
R14909 vdd.n2688 vdd.n633 185
R14910 vdd.n2771 vdd.n633 185
R14911 vdd.n2690 vdd.n2689 185
R14912 vdd.n2689 vdd.n631 185
R14913 vdd.n2691 vdd.n667 185
R14914 vdd.n2701 vdd.n667 185
R14915 vdd.n2692 vdd.n676 185
R14916 vdd.n676 vdd.n674 185
R14917 vdd.n2694 vdd.n2693 185
R14918 vdd.n2695 vdd.n2694 185
R14919 vdd.n2647 vdd.n675 185
R14920 vdd.n675 vdd.n671 185
R14921 vdd.n2646 vdd.n2645 185
R14922 vdd.n2645 vdd.n2644 185
R14923 vdd.n678 vdd.n677 185
R14924 vdd.n679 vdd.n678 185
R14925 vdd.n2637 vdd.n2636 185
R14926 vdd.n2638 vdd.n2637 185
R14927 vdd.n2633 vdd.n688 185
R14928 vdd.n688 vdd.n685 185
R14929 vdd.n2632 vdd.n2631 185
R14930 vdd.n2631 vdd.n2630 185
R14931 vdd.n690 vdd.n689 185
R14932 vdd.n698 vdd.n690 185
R14933 vdd.n2623 vdd.n2622 185
R14934 vdd.n2624 vdd.n2623 185
R14935 vdd.n2621 vdd.n699 185
R14936 vdd.n2472 vdd.n699 185
R14937 vdd.n2620 vdd.n2619 185
R14938 vdd.n2619 vdd.n2618 185
R14939 vdd.n701 vdd.n700 185
R14940 vdd.n702 vdd.n701 185
R14941 vdd.n2611 vdd.n2610 185
R14942 vdd.n2612 vdd.n2611 185
R14943 vdd.n2609 vdd.n711 185
R14944 vdd.n711 vdd.n708 185
R14945 vdd.n2608 vdd.n2607 185
R14946 vdd.n2607 vdd.n2606 185
R14947 vdd.n713 vdd.n712 185
R14948 vdd.n721 vdd.n713 185
R14949 vdd.n2599 vdd.n2598 185
R14950 vdd.n2600 vdd.n2599 185
R14951 vdd.n2597 vdd.n722 185
R14952 vdd.n728 vdd.n722 185
R14953 vdd.n2596 vdd.n2595 185
R14954 vdd.n2595 vdd.n2594 185
R14955 vdd.n724 vdd.n723 185
R14956 vdd.n725 vdd.n724 185
R14957 vdd.n2587 vdd.n2586 185
R14958 vdd.n2588 vdd.n2587 185
R14959 vdd.n2585 vdd.n734 185
R14960 vdd.n2493 vdd.n734 185
R14961 vdd.n2584 vdd.n2583 185
R14962 vdd.n2583 vdd.n2582 185
R14963 vdd.n736 vdd.n735 185
R14964 vdd.t66 vdd.n736 185
R14965 vdd.n2575 vdd.n2574 185
R14966 vdd.n2576 vdd.n2575 185
R14967 vdd.n2573 vdd.n744 185
R14968 vdd.n2572 vdd.n2571 185
R14969 vdd.n746 vdd.n745 185
R14970 vdd.n2358 vdd.n2357 185
R14971 vdd.n2360 vdd.n2359 185
R14972 vdd.n2362 vdd.n2361 185
R14973 vdd.n2364 vdd.n2363 185
R14974 vdd.n2366 vdd.n2365 185
R14975 vdd.n2368 vdd.n2367 185
R14976 vdd.n2370 vdd.n2369 185
R14977 vdd.n2372 vdd.n2371 185
R14978 vdd.n2374 vdd.n2373 185
R14979 vdd.n2376 vdd.n2375 185
R14980 vdd.n2378 vdd.n2377 185
R14981 vdd.n2380 vdd.n2379 185
R14982 vdd.n2382 vdd.n2381 185
R14983 vdd.n2384 vdd.n2383 185
R14984 vdd.n2386 vdd.n2385 185
R14985 vdd.n2388 vdd.n2387 185
R14986 vdd.n2390 vdd.n2389 185
R14987 vdd.n2392 vdd.n2391 185
R14988 vdd.n2394 vdd.n2393 185
R14989 vdd.n2396 vdd.n2395 185
R14990 vdd.n2398 vdd.n2397 185
R14991 vdd.n2400 vdd.n2399 185
R14992 vdd.n2402 vdd.n2401 185
R14993 vdd.n2404 vdd.n2403 185
R14994 vdd.n2406 vdd.n2405 185
R14995 vdd.n2408 vdd.n2407 185
R14996 vdd.n2410 vdd.n2409 185
R14997 vdd.n2412 vdd.n2411 185
R14998 vdd.n2414 vdd.n2413 185
R14999 vdd.n2416 vdd.n2415 185
R15000 vdd.n2418 vdd.n2417 185
R15001 vdd.n2419 vdd.n2349 185
R15002 vdd.n2569 vdd.n2349 185
R15003 vdd.n2774 vdd.n2773 185
R15004 vdd.n2775 vdd.n624 185
R15005 vdd.n2777 vdd.n2776 185
R15006 vdd.n2779 vdd.n622 185
R15007 vdd.n2781 vdd.n2780 185
R15008 vdd.n2782 vdd.n621 185
R15009 vdd.n2784 vdd.n2783 185
R15010 vdd.n2786 vdd.n619 185
R15011 vdd.n2788 vdd.n2787 185
R15012 vdd.n2789 vdd.n618 185
R15013 vdd.n2791 vdd.n2790 185
R15014 vdd.n2793 vdd.n616 185
R15015 vdd.n2795 vdd.n2794 185
R15016 vdd.n2796 vdd.n615 185
R15017 vdd.n2798 vdd.n2797 185
R15018 vdd.n2800 vdd.n614 185
R15019 vdd.n2801 vdd.n611 185
R15020 vdd.n2804 vdd.n2803 185
R15021 vdd.n612 vdd.n610 185
R15022 vdd.n2660 vdd.n2659 185
R15023 vdd.n2662 vdd.n2661 185
R15024 vdd.n2664 vdd.n2656 185
R15025 vdd.n2666 vdd.n2665 185
R15026 vdd.n2667 vdd.n2655 185
R15027 vdd.n2669 vdd.n2668 185
R15028 vdd.n2671 vdd.n2653 185
R15029 vdd.n2673 vdd.n2672 185
R15030 vdd.n2674 vdd.n2652 185
R15031 vdd.n2676 vdd.n2675 185
R15032 vdd.n2678 vdd.n2650 185
R15033 vdd.n2680 vdd.n2679 185
R15034 vdd.n2681 vdd.n2649 185
R15035 vdd.n2683 vdd.n2682 185
R15036 vdd.n2685 vdd.n2648 185
R15037 vdd.n2687 vdd.n2686 185
R15038 vdd.n2686 vdd.n613 185
R15039 vdd.n2772 vdd.n628 185
R15040 vdd.n2772 vdd.n2771 185
R15041 vdd.n2424 vdd.n630 185
R15042 vdd.n631 vdd.n630 185
R15043 vdd.n2425 vdd.n666 185
R15044 vdd.n2701 vdd.n666 185
R15045 vdd.n2427 vdd.n2426 185
R15046 vdd.n2426 vdd.n674 185
R15047 vdd.n2428 vdd.n673 185
R15048 vdd.n2695 vdd.n673 185
R15049 vdd.n2430 vdd.n2429 185
R15050 vdd.n2429 vdd.n671 185
R15051 vdd.n2431 vdd.n681 185
R15052 vdd.n2644 vdd.n681 185
R15053 vdd.n2433 vdd.n2432 185
R15054 vdd.n2432 vdd.n679 185
R15055 vdd.n2434 vdd.n687 185
R15056 vdd.n2638 vdd.n687 185
R15057 vdd.n2436 vdd.n2435 185
R15058 vdd.n2435 vdd.n685 185
R15059 vdd.n2437 vdd.n692 185
R15060 vdd.n2630 vdd.n692 185
R15061 vdd.n2439 vdd.n2438 185
R15062 vdd.n2438 vdd.n698 185
R15063 vdd.n2440 vdd.n697 185
R15064 vdd.n2624 vdd.n697 185
R15065 vdd.n2474 vdd.n2473 185
R15066 vdd.n2473 vdd.n2472 185
R15067 vdd.n2475 vdd.n704 185
R15068 vdd.n2618 vdd.n704 185
R15069 vdd.n2477 vdd.n2476 185
R15070 vdd.n2476 vdd.n702 185
R15071 vdd.n2478 vdd.n710 185
R15072 vdd.n2612 vdd.n710 185
R15073 vdd.n2480 vdd.n2479 185
R15074 vdd.n2479 vdd.n708 185
R15075 vdd.n2481 vdd.n715 185
R15076 vdd.n2606 vdd.n715 185
R15077 vdd.n2483 vdd.n2482 185
R15078 vdd.n2482 vdd.n721 185
R15079 vdd.n2484 vdd.n720 185
R15080 vdd.n2600 vdd.n720 185
R15081 vdd.n2486 vdd.n2485 185
R15082 vdd.n2485 vdd.n728 185
R15083 vdd.n2487 vdd.n727 185
R15084 vdd.n2594 vdd.n727 185
R15085 vdd.n2489 vdd.n2488 185
R15086 vdd.n2488 vdd.n725 185
R15087 vdd.n2490 vdd.n733 185
R15088 vdd.n2588 vdd.n733 185
R15089 vdd.n2492 vdd.n2491 185
R15090 vdd.n2493 vdd.n2492 185
R15091 vdd.n2423 vdd.n738 185
R15092 vdd.n2582 vdd.n738 185
R15093 vdd.n2422 vdd.n2421 185
R15094 vdd.n2421 vdd.t66 185
R15095 vdd.n2420 vdd.n743 185
R15096 vdd.n2576 vdd.n743 185
R15097 vdd.n2040 vdd.n2039 185
R15098 vdd.n2041 vdd.n2040 185
R15099 vdd.n904 vdd.n902 185
R15100 vdd.n1606 vdd.n902 185
R15101 vdd.n1609 vdd.n1608 185
R15102 vdd.n1608 vdd.n1607 185
R15103 vdd.n907 vdd.n906 185
R15104 vdd.n908 vdd.n907 185
R15105 vdd.n1595 vdd.n1594 185
R15106 vdd.n1596 vdd.n1595 185
R15107 vdd.n916 vdd.n915 185
R15108 vdd.n1587 vdd.n915 185
R15109 vdd.n1590 vdd.n1589 185
R15110 vdd.n1589 vdd.n1588 185
R15111 vdd.n919 vdd.n918 185
R15112 vdd.n925 vdd.n919 185
R15113 vdd.n1578 vdd.n1577 185
R15114 vdd.n1579 vdd.n1578 185
R15115 vdd.n927 vdd.n926 185
R15116 vdd.n1570 vdd.n926 185
R15117 vdd.n1573 vdd.n1572 185
R15118 vdd.n1572 vdd.n1571 185
R15119 vdd.n930 vdd.n929 185
R15120 vdd.n931 vdd.n930 185
R15121 vdd.n1561 vdd.n1560 185
R15122 vdd.n1562 vdd.n1561 185
R15123 vdd.n939 vdd.n938 185
R15124 vdd.n938 vdd.n937 185
R15125 vdd.n1274 vdd.n1273 185
R15126 vdd.n1273 vdd.n1272 185
R15127 vdd.n942 vdd.n941 185
R15128 vdd.n948 vdd.n942 185
R15129 vdd.n1263 vdd.n1262 185
R15130 vdd.n1264 vdd.n1263 185
R15131 vdd.n950 vdd.n949 185
R15132 vdd.n1255 vdd.n949 185
R15133 vdd.n1258 vdd.n1257 185
R15134 vdd.n1257 vdd.n1256 185
R15135 vdd.n953 vdd.n952 185
R15136 vdd.n960 vdd.n953 185
R15137 vdd.n1246 vdd.n1245 185
R15138 vdd.n1247 vdd.n1246 185
R15139 vdd.n962 vdd.n961 185
R15140 vdd.n961 vdd.n959 185
R15141 vdd.n1241 vdd.n1240 185
R15142 vdd.n1240 vdd.n1239 185
R15143 vdd.n965 vdd.n964 185
R15144 vdd.n966 vdd.n965 185
R15145 vdd.n1230 vdd.n1229 185
R15146 vdd.n1231 vdd.n1230 185
R15147 vdd.n974 vdd.n973 185
R15148 vdd.n973 vdd.n972 185
R15149 vdd.n1225 vdd.n1224 185
R15150 vdd.n1224 vdd.n1223 185
R15151 vdd.n977 vdd.n976 185
R15152 vdd.n983 vdd.n977 185
R15153 vdd.n1214 vdd.n1213 185
R15154 vdd.n1215 vdd.n1214 185
R15155 vdd.n1210 vdd.n984 185
R15156 vdd.n1209 vdd.n987 185
R15157 vdd.n1208 vdd.n988 185
R15158 vdd.n988 vdd.n982 185
R15159 vdd.n991 vdd.n989 185
R15160 vdd.n1204 vdd.n993 185
R15161 vdd.n1203 vdd.n994 185
R15162 vdd.n1202 vdd.n996 185
R15163 vdd.n999 vdd.n997 185
R15164 vdd.n1198 vdd.n1001 185
R15165 vdd.n1197 vdd.n1002 185
R15166 vdd.n1196 vdd.n1004 185
R15167 vdd.n1007 vdd.n1005 185
R15168 vdd.n1192 vdd.n1009 185
R15169 vdd.n1191 vdd.n1010 185
R15170 vdd.n1190 vdd.n1012 185
R15171 vdd.n1015 vdd.n1013 185
R15172 vdd.n1186 vdd.n1017 185
R15173 vdd.n1185 vdd.n1018 185
R15174 vdd.n1184 vdd.n1020 185
R15175 vdd.n1025 vdd.n1023 185
R15176 vdd.n1180 vdd.n1027 185
R15177 vdd.n1179 vdd.n1028 185
R15178 vdd.n1178 vdd.n1030 185
R15179 vdd.n1033 vdd.n1031 185
R15180 vdd.n1174 vdd.n1035 185
R15181 vdd.n1173 vdd.n1036 185
R15182 vdd.n1172 vdd.n1038 185
R15183 vdd.n1041 vdd.n1039 185
R15184 vdd.n1168 vdd.n1043 185
R15185 vdd.n1167 vdd.n1044 185
R15186 vdd.n1166 vdd.n1046 185
R15187 vdd.n1049 vdd.n1047 185
R15188 vdd.n1162 vdd.n1051 185
R15189 vdd.n1161 vdd.n1052 185
R15190 vdd.n1160 vdd.n1054 185
R15191 vdd.n1057 vdd.n1055 185
R15192 vdd.n1156 vdd.n1059 185
R15193 vdd.n1155 vdd.n1060 185
R15194 vdd.n1154 vdd.n1062 185
R15195 vdd.n1065 vdd.n1063 185
R15196 vdd.n1150 vdd.n1067 185
R15197 vdd.n1149 vdd.n1146 185
R15198 vdd.n1144 vdd.n1068 185
R15199 vdd.n1143 vdd.n1142 185
R15200 vdd.n1073 vdd.n1070 185
R15201 vdd.n1138 vdd.n1074 185
R15202 vdd.n1137 vdd.n1076 185
R15203 vdd.n1136 vdd.n1077 185
R15204 vdd.n1081 vdd.n1078 185
R15205 vdd.n1132 vdd.n1082 185
R15206 vdd.n1131 vdd.n1084 185
R15207 vdd.n1130 vdd.n1085 185
R15208 vdd.n1089 vdd.n1086 185
R15209 vdd.n1126 vdd.n1090 185
R15210 vdd.n1125 vdd.n1092 185
R15211 vdd.n1124 vdd.n1093 185
R15212 vdd.n1097 vdd.n1094 185
R15213 vdd.n1120 vdd.n1098 185
R15214 vdd.n1119 vdd.n1100 185
R15215 vdd.n1118 vdd.n1101 185
R15216 vdd.n1105 vdd.n1102 185
R15217 vdd.n1114 vdd.n1106 185
R15218 vdd.n1113 vdd.n1108 185
R15219 vdd.n1109 vdd.n981 185
R15220 vdd.n982 vdd.n981 185
R15221 vdd.n2044 vdd.n2043 185
R15222 vdd.n2048 vdd.n897 185
R15223 vdd.n1711 vdd.n896 185
R15224 vdd.n1714 vdd.n1713 185
R15225 vdd.n1716 vdd.n1715 185
R15226 vdd.n1719 vdd.n1718 185
R15227 vdd.n1721 vdd.n1720 185
R15228 vdd.n1723 vdd.n1709 185
R15229 vdd.n1725 vdd.n1724 185
R15230 vdd.n1726 vdd.n1703 185
R15231 vdd.n1728 vdd.n1727 185
R15232 vdd.n1730 vdd.n1701 185
R15233 vdd.n1732 vdd.n1731 185
R15234 vdd.n1733 vdd.n1696 185
R15235 vdd.n1735 vdd.n1734 185
R15236 vdd.n1737 vdd.n1694 185
R15237 vdd.n1739 vdd.n1738 185
R15238 vdd.n1740 vdd.n1690 185
R15239 vdd.n1742 vdd.n1741 185
R15240 vdd.n1744 vdd.n1687 185
R15241 vdd.n1746 vdd.n1745 185
R15242 vdd.n1688 vdd.n1681 185
R15243 vdd.n1750 vdd.n1685 185
R15244 vdd.n1751 vdd.n1677 185
R15245 vdd.n1753 vdd.n1752 185
R15246 vdd.n1755 vdd.n1675 185
R15247 vdd.n1757 vdd.n1756 185
R15248 vdd.n1758 vdd.n1670 185
R15249 vdd.n1760 vdd.n1759 185
R15250 vdd.n1762 vdd.n1668 185
R15251 vdd.n1764 vdd.n1763 185
R15252 vdd.n1765 vdd.n1663 185
R15253 vdd.n1767 vdd.n1766 185
R15254 vdd.n1769 vdd.n1661 185
R15255 vdd.n1771 vdd.n1770 185
R15256 vdd.n1772 vdd.n1656 185
R15257 vdd.n1774 vdd.n1773 185
R15258 vdd.n1776 vdd.n1654 185
R15259 vdd.n1778 vdd.n1777 185
R15260 vdd.n1779 vdd.n1650 185
R15261 vdd.n1781 vdd.n1780 185
R15262 vdd.n1783 vdd.n1647 185
R15263 vdd.n1785 vdd.n1784 185
R15264 vdd.n1648 vdd.n1641 185
R15265 vdd.n1789 vdd.n1645 185
R15266 vdd.n1790 vdd.n1637 185
R15267 vdd.n1792 vdd.n1791 185
R15268 vdd.n1794 vdd.n1635 185
R15269 vdd.n1796 vdd.n1795 185
R15270 vdd.n1797 vdd.n1630 185
R15271 vdd.n1799 vdd.n1798 185
R15272 vdd.n1801 vdd.n1628 185
R15273 vdd.n1803 vdd.n1802 185
R15274 vdd.n1804 vdd.n1623 185
R15275 vdd.n1806 vdd.n1805 185
R15276 vdd.n1808 vdd.n1622 185
R15277 vdd.n1809 vdd.n1619 185
R15278 vdd.n1812 vdd.n1811 185
R15279 vdd.n1621 vdd.n1617 185
R15280 vdd.n2029 vdd.n1615 185
R15281 vdd.n2031 vdd.n2030 185
R15282 vdd.n2033 vdd.n1613 185
R15283 vdd.n2035 vdd.n2034 185
R15284 vdd.n2036 vdd.n903 185
R15285 vdd.n2042 vdd.n900 185
R15286 vdd.n2042 vdd.n2041 185
R15287 vdd.n911 vdd.n899 185
R15288 vdd.n1606 vdd.n899 185
R15289 vdd.n1605 vdd.n1604 185
R15290 vdd.n1607 vdd.n1605 185
R15291 vdd.n910 vdd.n909 185
R15292 vdd.n909 vdd.n908 185
R15293 vdd.n1598 vdd.n1597 185
R15294 vdd.n1597 vdd.n1596 185
R15295 vdd.n914 vdd.n913 185
R15296 vdd.n1587 vdd.n914 185
R15297 vdd.n1586 vdd.n1585 185
R15298 vdd.n1588 vdd.n1586 185
R15299 vdd.n921 vdd.n920 185
R15300 vdd.n925 vdd.n920 185
R15301 vdd.n1581 vdd.n1580 185
R15302 vdd.n1580 vdd.n1579 185
R15303 vdd.n924 vdd.n923 185
R15304 vdd.n1570 vdd.n924 185
R15305 vdd.n1569 vdd.n1568 185
R15306 vdd.n1571 vdd.n1569 185
R15307 vdd.n933 vdd.n932 185
R15308 vdd.n932 vdd.n931 185
R15309 vdd.n1564 vdd.n1563 185
R15310 vdd.n1563 vdd.n1562 185
R15311 vdd.n936 vdd.n935 185
R15312 vdd.n937 vdd.n936 185
R15313 vdd.n1271 vdd.n1270 185
R15314 vdd.n1272 vdd.n1271 185
R15315 vdd.n944 vdd.n943 185
R15316 vdd.n948 vdd.n943 185
R15317 vdd.n1266 vdd.n1265 185
R15318 vdd.n1265 vdd.n1264 185
R15319 vdd.n947 vdd.n946 185
R15320 vdd.n1255 vdd.n947 185
R15321 vdd.n1254 vdd.n1253 185
R15322 vdd.n1256 vdd.n1254 185
R15323 vdd.n955 vdd.n954 185
R15324 vdd.n960 vdd.n954 185
R15325 vdd.n1249 vdd.n1248 185
R15326 vdd.n1248 vdd.n1247 185
R15327 vdd.n958 vdd.n957 185
R15328 vdd.n959 vdd.n958 185
R15329 vdd.n1238 vdd.n1237 185
R15330 vdd.n1239 vdd.n1238 185
R15331 vdd.n968 vdd.n967 185
R15332 vdd.n967 vdd.n966 185
R15333 vdd.n1233 vdd.n1232 185
R15334 vdd.n1232 vdd.n1231 185
R15335 vdd.n971 vdd.n970 185
R15336 vdd.n972 vdd.n971 185
R15337 vdd.n1222 vdd.n1221 185
R15338 vdd.n1223 vdd.n1222 185
R15339 vdd.n979 vdd.n978 185
R15340 vdd.n983 vdd.n978 185
R15341 vdd.n1217 vdd.n1216 185
R15342 vdd.n1216 vdd.n1215 185
R15343 vdd.n784 vdd.n782 185
R15344 vdd.n2244 vdd.n782 185
R15345 vdd.n2166 vdd.n801 185
R15346 vdd.n801 vdd.t159 185
R15347 vdd.n2168 vdd.n2167 185
R15348 vdd.n2169 vdd.n2168 185
R15349 vdd.n2165 vdd.n800 185
R15350 vdd.n1868 vdd.n800 185
R15351 vdd.n2164 vdd.n2163 185
R15352 vdd.n2163 vdd.n2162 185
R15353 vdd.n803 vdd.n802 185
R15354 vdd.n804 vdd.n803 185
R15355 vdd.n2153 vdd.n2152 185
R15356 vdd.n2154 vdd.n2153 185
R15357 vdd.n2151 vdd.n814 185
R15358 vdd.n814 vdd.n811 185
R15359 vdd.n2150 vdd.n2149 185
R15360 vdd.n2149 vdd.n2148 185
R15361 vdd.n816 vdd.n815 185
R15362 vdd.n817 vdd.n816 185
R15363 vdd.n2141 vdd.n2140 185
R15364 vdd.n2142 vdd.n2141 185
R15365 vdd.n2139 vdd.n825 185
R15366 vdd.n830 vdd.n825 185
R15367 vdd.n2138 vdd.n2137 185
R15368 vdd.n2137 vdd.n2136 185
R15369 vdd.n827 vdd.n826 185
R15370 vdd.n836 vdd.n827 185
R15371 vdd.n2129 vdd.n2128 185
R15372 vdd.n2130 vdd.n2129 185
R15373 vdd.n2127 vdd.n837 185
R15374 vdd.n1969 vdd.n837 185
R15375 vdd.n2126 vdd.n2125 185
R15376 vdd.n2125 vdd.n2124 185
R15377 vdd.n839 vdd.n838 185
R15378 vdd.n840 vdd.n839 185
R15379 vdd.n2117 vdd.n2116 185
R15380 vdd.n2118 vdd.n2117 185
R15381 vdd.n2115 vdd.n849 185
R15382 vdd.n849 vdd.n846 185
R15383 vdd.n2114 vdd.n2113 185
R15384 vdd.n2113 vdd.n2112 185
R15385 vdd.n851 vdd.n850 185
R15386 vdd.n861 vdd.n851 185
R15387 vdd.n2104 vdd.n2103 185
R15388 vdd.n2105 vdd.n2104 185
R15389 vdd.n2102 vdd.n862 185
R15390 vdd.n862 vdd.n858 185
R15391 vdd.n2101 vdd.n2100 185
R15392 vdd.n2100 vdd.n2099 185
R15393 vdd.n864 vdd.n863 185
R15394 vdd.n865 vdd.n864 185
R15395 vdd.n2092 vdd.n2091 185
R15396 vdd.n2093 vdd.n2092 185
R15397 vdd.n2090 vdd.n874 185
R15398 vdd.n874 vdd.n871 185
R15399 vdd.n2089 vdd.n2088 185
R15400 vdd.n2088 vdd.n2087 185
R15401 vdd.n876 vdd.n875 185
R15402 vdd.n1824 vdd.n1823 185
R15403 vdd.n1825 vdd.n1821 185
R15404 vdd.n1821 vdd.n877 185
R15405 vdd.n1827 vdd.n1826 185
R15406 vdd.n1829 vdd.n1820 185
R15407 vdd.n1832 vdd.n1831 185
R15408 vdd.n1833 vdd.n1819 185
R15409 vdd.n1835 vdd.n1834 185
R15410 vdd.n1837 vdd.n1818 185
R15411 vdd.n1840 vdd.n1839 185
R15412 vdd.n1841 vdd.n1817 185
R15413 vdd.n1843 vdd.n1842 185
R15414 vdd.n1845 vdd.n1816 185
R15415 vdd.n1848 vdd.n1847 185
R15416 vdd.n1849 vdd.n1815 185
R15417 vdd.n1851 vdd.n1850 185
R15418 vdd.n1853 vdd.n1814 185
R15419 vdd.n2026 vdd.n1854 185
R15420 vdd.n2025 vdd.n2024 185
R15421 vdd.n2022 vdd.n1855 185
R15422 vdd.n2020 vdd.n2019 185
R15423 vdd.n2018 vdd.n1856 185
R15424 vdd.n2017 vdd.n2016 185
R15425 vdd.n2014 vdd.n1857 185
R15426 vdd.n2012 vdd.n2011 185
R15427 vdd.n2010 vdd.n1858 185
R15428 vdd.n2009 vdd.n2008 185
R15429 vdd.n2006 vdd.n1859 185
R15430 vdd.n2004 vdd.n2003 185
R15431 vdd.n2002 vdd.n1860 185
R15432 vdd.n2001 vdd.n2000 185
R15433 vdd.n1998 vdd.n1861 185
R15434 vdd.n1996 vdd.n1995 185
R15435 vdd.n1994 vdd.n1862 185
R15436 vdd.n1993 vdd.n1992 185
R15437 vdd.n2247 vdd.n2246 185
R15438 vdd.n2249 vdd.n2248 185
R15439 vdd.n2251 vdd.n2250 185
R15440 vdd.n2254 vdd.n2253 185
R15441 vdd.n2256 vdd.n2255 185
R15442 vdd.n2258 vdd.n2257 185
R15443 vdd.n2260 vdd.n2259 185
R15444 vdd.n2262 vdd.n2261 185
R15445 vdd.n2264 vdd.n2263 185
R15446 vdd.n2266 vdd.n2265 185
R15447 vdd.n2268 vdd.n2267 185
R15448 vdd.n2270 vdd.n2269 185
R15449 vdd.n2272 vdd.n2271 185
R15450 vdd.n2274 vdd.n2273 185
R15451 vdd.n2276 vdd.n2275 185
R15452 vdd.n2278 vdd.n2277 185
R15453 vdd.n2280 vdd.n2279 185
R15454 vdd.n2282 vdd.n2281 185
R15455 vdd.n2284 vdd.n2283 185
R15456 vdd.n2286 vdd.n2285 185
R15457 vdd.n2288 vdd.n2287 185
R15458 vdd.n2290 vdd.n2289 185
R15459 vdd.n2292 vdd.n2291 185
R15460 vdd.n2294 vdd.n2293 185
R15461 vdd.n2296 vdd.n2295 185
R15462 vdd.n2298 vdd.n2297 185
R15463 vdd.n2300 vdd.n2299 185
R15464 vdd.n2302 vdd.n2301 185
R15465 vdd.n2304 vdd.n2303 185
R15466 vdd.n2306 vdd.n2305 185
R15467 vdd.n2308 vdd.n2307 185
R15468 vdd.n2310 vdd.n2309 185
R15469 vdd.n2312 vdd.n2311 185
R15470 vdd.n2313 vdd.n783 185
R15471 vdd.n2315 vdd.n2314 185
R15472 vdd.n2316 vdd.n2315 185
R15473 vdd.n2245 vdd.n787 185
R15474 vdd.n2245 vdd.n2244 185
R15475 vdd.n1866 vdd.n788 185
R15476 vdd.t159 vdd.n788 185
R15477 vdd.n1867 vdd.n798 185
R15478 vdd.n2169 vdd.n798 185
R15479 vdd.n1870 vdd.n1869 185
R15480 vdd.n1869 vdd.n1868 185
R15481 vdd.n1871 vdd.n805 185
R15482 vdd.n2162 vdd.n805 185
R15483 vdd.n1873 vdd.n1872 185
R15484 vdd.n1872 vdd.n804 185
R15485 vdd.n1874 vdd.n812 185
R15486 vdd.n2154 vdd.n812 185
R15487 vdd.n1876 vdd.n1875 185
R15488 vdd.n1875 vdd.n811 185
R15489 vdd.n1877 vdd.n818 185
R15490 vdd.n2148 vdd.n818 185
R15491 vdd.n1879 vdd.n1878 185
R15492 vdd.n1878 vdd.n817 185
R15493 vdd.n1880 vdd.n823 185
R15494 vdd.n2142 vdd.n823 185
R15495 vdd.n1882 vdd.n1881 185
R15496 vdd.n1881 vdd.n830 185
R15497 vdd.n1883 vdd.n828 185
R15498 vdd.n2136 vdd.n828 185
R15499 vdd.n1885 vdd.n1884 185
R15500 vdd.n1884 vdd.n836 185
R15501 vdd.n1886 vdd.n834 185
R15502 vdd.n2130 vdd.n834 185
R15503 vdd.n1971 vdd.n1970 185
R15504 vdd.n1970 vdd.n1969 185
R15505 vdd.n1972 vdd.n841 185
R15506 vdd.n2124 vdd.n841 185
R15507 vdd.n1974 vdd.n1973 185
R15508 vdd.n1973 vdd.n840 185
R15509 vdd.n1975 vdd.n847 185
R15510 vdd.n2118 vdd.n847 185
R15511 vdd.n1977 vdd.n1976 185
R15512 vdd.n1976 vdd.n846 185
R15513 vdd.n1978 vdd.n852 185
R15514 vdd.n2112 vdd.n852 185
R15515 vdd.n1980 vdd.n1979 185
R15516 vdd.n1979 vdd.n861 185
R15517 vdd.n1981 vdd.n859 185
R15518 vdd.n2105 vdd.n859 185
R15519 vdd.n1983 vdd.n1982 185
R15520 vdd.n1982 vdd.n858 185
R15521 vdd.n1984 vdd.n866 185
R15522 vdd.n2099 vdd.n866 185
R15523 vdd.n1986 vdd.n1985 185
R15524 vdd.n1985 vdd.n865 185
R15525 vdd.n1987 vdd.n872 185
R15526 vdd.n2093 vdd.n872 185
R15527 vdd.n1989 vdd.n1988 185
R15528 vdd.n1988 vdd.n871 185
R15529 vdd.n1990 vdd.n878 185
R15530 vdd.n2087 vdd.n878 185
R15531 vdd.n3137 vdd.n3136 185
R15532 vdd.n3138 vdd.n3137 185
R15533 vdd.n347 vdd.n346 185
R15534 vdd.n3139 vdd.n347 185
R15535 vdd.n3142 vdd.n3141 185
R15536 vdd.n3141 vdd.n3140 185
R15537 vdd.n3143 vdd.n341 185
R15538 vdd.n341 vdd.n340 185
R15539 vdd.n3145 vdd.n3144 185
R15540 vdd.n3146 vdd.n3145 185
R15541 vdd.n336 vdd.n335 185
R15542 vdd.n3147 vdd.n336 185
R15543 vdd.n3150 vdd.n3149 185
R15544 vdd.n3149 vdd.n3148 185
R15545 vdd.n3151 vdd.n330 185
R15546 vdd.n330 vdd.n329 185
R15547 vdd.n3153 vdd.n3152 185
R15548 vdd.n3154 vdd.n3153 185
R15549 vdd.n324 vdd.n323 185
R15550 vdd.n3155 vdd.n324 185
R15551 vdd.n3158 vdd.n3157 185
R15552 vdd.n3157 vdd.n3156 185
R15553 vdd.n3159 vdd.n319 185
R15554 vdd.n325 vdd.n319 185
R15555 vdd.n3161 vdd.n3160 185
R15556 vdd.n3162 vdd.n3161 185
R15557 vdd.n315 vdd.n313 185
R15558 vdd.n3163 vdd.n315 185
R15559 vdd.n3166 vdd.n3165 185
R15560 vdd.n3165 vdd.n3164 185
R15561 vdd.n314 vdd.n312 185
R15562 vdd.n481 vdd.n314 185
R15563 vdd.n2988 vdd.n2987 185
R15564 vdd.n2989 vdd.n2988 185
R15565 vdd.n483 vdd.n482 185
R15566 vdd.n2980 vdd.n482 185
R15567 vdd.n2983 vdd.n2982 185
R15568 vdd.n2982 vdd.n2981 185
R15569 vdd.n486 vdd.n485 185
R15570 vdd.n493 vdd.n486 185
R15571 vdd.n2971 vdd.n2970 185
R15572 vdd.n2972 vdd.n2971 185
R15573 vdd.n495 vdd.n494 185
R15574 vdd.n494 vdd.n492 185
R15575 vdd.n2966 vdd.n2965 185
R15576 vdd.n2965 vdd.n2964 185
R15577 vdd.n498 vdd.n497 185
R15578 vdd.n499 vdd.n498 185
R15579 vdd.n2955 vdd.n2954 185
R15580 vdd.n2956 vdd.n2955 185
R15581 vdd.n507 vdd.n506 185
R15582 vdd.n506 vdd.n505 185
R15583 vdd.n2950 vdd.n2949 185
R15584 vdd.n2949 vdd.n2948 185
R15585 vdd.n510 vdd.n509 185
R15586 vdd.n511 vdd.n510 185
R15587 vdd.n2939 vdd.n2938 185
R15588 vdd.n2940 vdd.n2939 185
R15589 vdd.n2935 vdd.n517 185
R15590 vdd.n2934 vdd.n2933 185
R15591 vdd.n2931 vdd.n519 185
R15592 vdd.n2931 vdd.n516 185
R15593 vdd.n2930 vdd.n2929 185
R15594 vdd.n2928 vdd.n2927 185
R15595 vdd.n2926 vdd.n2925 185
R15596 vdd.n2924 vdd.n2923 185
R15597 vdd.n2922 vdd.n525 185
R15598 vdd.n2920 vdd.n2919 185
R15599 vdd.n2918 vdd.n526 185
R15600 vdd.n2917 vdd.n2916 185
R15601 vdd.n2914 vdd.n531 185
R15602 vdd.n2912 vdd.n2911 185
R15603 vdd.n2910 vdd.n532 185
R15604 vdd.n2909 vdd.n2908 185
R15605 vdd.n2906 vdd.n537 185
R15606 vdd.n2904 vdd.n2903 185
R15607 vdd.n2902 vdd.n538 185
R15608 vdd.n2901 vdd.n2900 185
R15609 vdd.n2898 vdd.n545 185
R15610 vdd.n2896 vdd.n2895 185
R15611 vdd.n2894 vdd.n546 185
R15612 vdd.n2893 vdd.n2892 185
R15613 vdd.n2890 vdd.n551 185
R15614 vdd.n2888 vdd.n2887 185
R15615 vdd.n2886 vdd.n552 185
R15616 vdd.n2885 vdd.n2884 185
R15617 vdd.n2882 vdd.n557 185
R15618 vdd.n2880 vdd.n2879 185
R15619 vdd.n2878 vdd.n558 185
R15620 vdd.n2877 vdd.n2876 185
R15621 vdd.n2874 vdd.n563 185
R15622 vdd.n2872 vdd.n2871 185
R15623 vdd.n2870 vdd.n564 185
R15624 vdd.n2869 vdd.n2868 185
R15625 vdd.n2866 vdd.n569 185
R15626 vdd.n2864 vdd.n2863 185
R15627 vdd.n2862 vdd.n570 185
R15628 vdd.n2861 vdd.n2860 185
R15629 vdd.n2858 vdd.n575 185
R15630 vdd.n2856 vdd.n2855 185
R15631 vdd.n2854 vdd.n576 185
R15632 vdd.n585 vdd.n579 185
R15633 vdd.n2850 vdd.n2849 185
R15634 vdd.n2847 vdd.n583 185
R15635 vdd.n2846 vdd.n2845 185
R15636 vdd.n2844 vdd.n2843 185
R15637 vdd.n2842 vdd.n589 185
R15638 vdd.n2840 vdd.n2839 185
R15639 vdd.n2838 vdd.n590 185
R15640 vdd.n2837 vdd.n2836 185
R15641 vdd.n2834 vdd.n595 185
R15642 vdd.n2832 vdd.n2831 185
R15643 vdd.n2830 vdd.n596 185
R15644 vdd.n2829 vdd.n2828 185
R15645 vdd.n2826 vdd.n601 185
R15646 vdd.n2824 vdd.n2823 185
R15647 vdd.n2822 vdd.n602 185
R15648 vdd.n2821 vdd.n2820 185
R15649 vdd.n2818 vdd.n2817 185
R15650 vdd.n2816 vdd.n2815 185
R15651 vdd.n2814 vdd.n2813 185
R15652 vdd.n2812 vdd.n2811 185
R15653 vdd.n2807 vdd.n515 185
R15654 vdd.n516 vdd.n515 185
R15655 vdd.n3020 vdd.n3019 185
R15656 vdd.n3024 vdd.n462 185
R15657 vdd.n3026 vdd.n3025 185
R15658 vdd.n3028 vdd.n460 185
R15659 vdd.n3030 vdd.n3029 185
R15660 vdd.n3031 vdd.n455 185
R15661 vdd.n3033 vdd.n3032 185
R15662 vdd.n3035 vdd.n453 185
R15663 vdd.n3037 vdd.n3036 185
R15664 vdd.n3038 vdd.n448 185
R15665 vdd.n3040 vdd.n3039 185
R15666 vdd.n3042 vdd.n446 185
R15667 vdd.n3044 vdd.n3043 185
R15668 vdd.n3045 vdd.n441 185
R15669 vdd.n3047 vdd.n3046 185
R15670 vdd.n3049 vdd.n439 185
R15671 vdd.n3051 vdd.n3050 185
R15672 vdd.n3052 vdd.n435 185
R15673 vdd.n3054 vdd.n3053 185
R15674 vdd.n3056 vdd.n432 185
R15675 vdd.n3058 vdd.n3057 185
R15676 vdd.n433 vdd.n426 185
R15677 vdd.n3062 vdd.n430 185
R15678 vdd.n3063 vdd.n422 185
R15679 vdd.n3065 vdd.n3064 185
R15680 vdd.n3067 vdd.n420 185
R15681 vdd.n3069 vdd.n3068 185
R15682 vdd.n3070 vdd.n415 185
R15683 vdd.n3072 vdd.n3071 185
R15684 vdd.n3074 vdd.n413 185
R15685 vdd.n3076 vdd.n3075 185
R15686 vdd.n3077 vdd.n408 185
R15687 vdd.n3079 vdd.n3078 185
R15688 vdd.n3081 vdd.n406 185
R15689 vdd.n3083 vdd.n3082 185
R15690 vdd.n3084 vdd.n401 185
R15691 vdd.n3086 vdd.n3085 185
R15692 vdd.n3088 vdd.n399 185
R15693 vdd.n3090 vdd.n3089 185
R15694 vdd.n3091 vdd.n395 185
R15695 vdd.n3093 vdd.n3092 185
R15696 vdd.n3095 vdd.n392 185
R15697 vdd.n3097 vdd.n3096 185
R15698 vdd.n393 vdd.n386 185
R15699 vdd.n3101 vdd.n390 185
R15700 vdd.n3102 vdd.n382 185
R15701 vdd.n3104 vdd.n3103 185
R15702 vdd.n3106 vdd.n380 185
R15703 vdd.n3108 vdd.n3107 185
R15704 vdd.n3109 vdd.n375 185
R15705 vdd.n3111 vdd.n3110 185
R15706 vdd.n3113 vdd.n373 185
R15707 vdd.n3115 vdd.n3114 185
R15708 vdd.n3116 vdd.n368 185
R15709 vdd.n3118 vdd.n3117 185
R15710 vdd.n3120 vdd.n366 185
R15711 vdd.n3122 vdd.n3121 185
R15712 vdd.n3123 vdd.n360 185
R15713 vdd.n3125 vdd.n3124 185
R15714 vdd.n3127 vdd.n359 185
R15715 vdd.n3128 vdd.n358 185
R15716 vdd.n3131 vdd.n3130 185
R15717 vdd.n3132 vdd.n356 185
R15718 vdd.n3133 vdd.n352 185
R15719 vdd.n3015 vdd.n350 185
R15720 vdd.n3138 vdd.n350 185
R15721 vdd.n3014 vdd.n349 185
R15722 vdd.n3139 vdd.n349 185
R15723 vdd.n3013 vdd.n348 185
R15724 vdd.n3140 vdd.n348 185
R15725 vdd.n468 vdd.n467 185
R15726 vdd.n467 vdd.n340 185
R15727 vdd.n3009 vdd.n339 185
R15728 vdd.n3146 vdd.n339 185
R15729 vdd.n3008 vdd.n338 185
R15730 vdd.n3147 vdd.n338 185
R15731 vdd.n3007 vdd.n337 185
R15732 vdd.n3148 vdd.n337 185
R15733 vdd.n471 vdd.n470 185
R15734 vdd.n470 vdd.n329 185
R15735 vdd.n3003 vdd.n328 185
R15736 vdd.n3154 vdd.n328 185
R15737 vdd.n3002 vdd.n327 185
R15738 vdd.n3155 vdd.n327 185
R15739 vdd.n3001 vdd.n326 185
R15740 vdd.n3156 vdd.n326 185
R15741 vdd.n474 vdd.n473 185
R15742 vdd.n473 vdd.n325 185
R15743 vdd.n2997 vdd.n318 185
R15744 vdd.n3162 vdd.n318 185
R15745 vdd.n2996 vdd.n317 185
R15746 vdd.n3163 vdd.n317 185
R15747 vdd.n2995 vdd.n316 185
R15748 vdd.n3164 vdd.n316 185
R15749 vdd.n480 vdd.n476 185
R15750 vdd.n481 vdd.n480 185
R15751 vdd.n2991 vdd.n2990 185
R15752 vdd.n2990 vdd.n2989 185
R15753 vdd.n479 vdd.n478 185
R15754 vdd.n2980 vdd.n479 185
R15755 vdd.n2979 vdd.n2978 185
R15756 vdd.n2981 vdd.n2979 185
R15757 vdd.n488 vdd.n487 185
R15758 vdd.n493 vdd.n487 185
R15759 vdd.n2974 vdd.n2973 185
R15760 vdd.n2973 vdd.n2972 185
R15761 vdd.n491 vdd.n490 185
R15762 vdd.n492 vdd.n491 185
R15763 vdd.n2963 vdd.n2962 185
R15764 vdd.n2964 vdd.n2963 185
R15765 vdd.n501 vdd.n500 185
R15766 vdd.n500 vdd.n499 185
R15767 vdd.n2958 vdd.n2957 185
R15768 vdd.n2957 vdd.n2956 185
R15769 vdd.n504 vdd.n503 185
R15770 vdd.n505 vdd.n504 185
R15771 vdd.n2947 vdd.n2946 185
R15772 vdd.n2948 vdd.n2947 185
R15773 vdd.n513 vdd.n512 185
R15774 vdd.n512 vdd.n511 185
R15775 vdd.n2942 vdd.n2941 185
R15776 vdd.n2941 vdd.n2940 185
R15777 vdd.n741 vdd.n740 185
R15778 vdd.n2567 vdd.n2566 185
R15779 vdd.n2565 vdd.n2350 185
R15780 vdd.n2569 vdd.n2350 185
R15781 vdd.n2564 vdd.n2563 185
R15782 vdd.n2562 vdd.n2561 185
R15783 vdd.n2560 vdd.n2559 185
R15784 vdd.n2558 vdd.n2557 185
R15785 vdd.n2556 vdd.n2555 185
R15786 vdd.n2554 vdd.n2553 185
R15787 vdd.n2552 vdd.n2551 185
R15788 vdd.n2550 vdd.n2549 185
R15789 vdd.n2548 vdd.n2547 185
R15790 vdd.n2546 vdd.n2545 185
R15791 vdd.n2544 vdd.n2543 185
R15792 vdd.n2542 vdd.n2541 185
R15793 vdd.n2540 vdd.n2539 185
R15794 vdd.n2538 vdd.n2537 185
R15795 vdd.n2536 vdd.n2535 185
R15796 vdd.n2534 vdd.n2533 185
R15797 vdd.n2532 vdd.n2531 185
R15798 vdd.n2530 vdd.n2529 185
R15799 vdd.n2528 vdd.n2527 185
R15800 vdd.n2526 vdd.n2525 185
R15801 vdd.n2524 vdd.n2523 185
R15802 vdd.n2522 vdd.n2521 185
R15803 vdd.n2520 vdd.n2519 185
R15804 vdd.n2518 vdd.n2517 185
R15805 vdd.n2516 vdd.n2515 185
R15806 vdd.n2514 vdd.n2513 185
R15807 vdd.n2512 vdd.n2511 185
R15808 vdd.n2510 vdd.n2509 185
R15809 vdd.n2508 vdd.n2507 185
R15810 vdd.n2505 vdd.n2504 185
R15811 vdd.n2503 vdd.n2502 185
R15812 vdd.n2501 vdd.n2500 185
R15813 vdd.n2708 vdd.n2707 185
R15814 vdd.n2709 vdd.n660 185
R15815 vdd.n2711 vdd.n2710 185
R15816 vdd.n2713 vdd.n658 185
R15817 vdd.n2715 vdd.n2714 185
R15818 vdd.n2716 vdd.n657 185
R15819 vdd.n2718 vdd.n2717 185
R15820 vdd.n2720 vdd.n655 185
R15821 vdd.n2722 vdd.n2721 185
R15822 vdd.n2723 vdd.n654 185
R15823 vdd.n2725 vdd.n2724 185
R15824 vdd.n2727 vdd.n652 185
R15825 vdd.n2729 vdd.n2728 185
R15826 vdd.n2730 vdd.n651 185
R15827 vdd.n2732 vdd.n2731 185
R15828 vdd.n2734 vdd.n649 185
R15829 vdd.n2736 vdd.n2735 185
R15830 vdd.n2738 vdd.n648 185
R15831 vdd.n2740 vdd.n2739 185
R15832 vdd.n2742 vdd.n646 185
R15833 vdd.n2744 vdd.n2743 185
R15834 vdd.n2745 vdd.n645 185
R15835 vdd.n2747 vdd.n2746 185
R15836 vdd.n2749 vdd.n643 185
R15837 vdd.n2751 vdd.n2750 185
R15838 vdd.n2752 vdd.n642 185
R15839 vdd.n2754 vdd.n2753 185
R15840 vdd.n2756 vdd.n640 185
R15841 vdd.n2758 vdd.n2757 185
R15842 vdd.n2759 vdd.n639 185
R15843 vdd.n2761 vdd.n2760 185
R15844 vdd.n2763 vdd.n638 185
R15845 vdd.n2764 vdd.n637 185
R15846 vdd.n2767 vdd.n2766 185
R15847 vdd.n2768 vdd.n635 185
R15848 vdd.n635 vdd.n613 185
R15849 vdd.n2705 vdd.n632 185
R15850 vdd.n2771 vdd.n632 185
R15851 vdd.n2704 vdd.n2703 185
R15852 vdd.n2703 vdd.n631 185
R15853 vdd.n2702 vdd.n664 185
R15854 vdd.n2702 vdd.n2701 185
R15855 vdd.n2456 vdd.n665 185
R15856 vdd.n674 vdd.n665 185
R15857 vdd.n2457 vdd.n672 185
R15858 vdd.n2695 vdd.n672 185
R15859 vdd.n2459 vdd.n2458 185
R15860 vdd.n2458 vdd.n671 185
R15861 vdd.n2460 vdd.n680 185
R15862 vdd.n2644 vdd.n680 185
R15863 vdd.n2462 vdd.n2461 185
R15864 vdd.n2461 vdd.n679 185
R15865 vdd.n2463 vdd.n686 185
R15866 vdd.n2638 vdd.n686 185
R15867 vdd.n2465 vdd.n2464 185
R15868 vdd.n2464 vdd.n685 185
R15869 vdd.n2466 vdd.n691 185
R15870 vdd.n2630 vdd.n691 185
R15871 vdd.n2468 vdd.n2467 185
R15872 vdd.n2467 vdd.n698 185
R15873 vdd.n2469 vdd.n696 185
R15874 vdd.n2624 vdd.n696 185
R15875 vdd.n2471 vdd.n2470 185
R15876 vdd.n2472 vdd.n2471 185
R15877 vdd.n2455 vdd.n703 185
R15878 vdd.n2618 vdd.n703 185
R15879 vdd.n2454 vdd.n2453 185
R15880 vdd.n2453 vdd.n702 185
R15881 vdd.n2452 vdd.n709 185
R15882 vdd.n2612 vdd.n709 185
R15883 vdd.n2451 vdd.n2450 185
R15884 vdd.n2450 vdd.n708 185
R15885 vdd.n2449 vdd.n714 185
R15886 vdd.n2606 vdd.n714 185
R15887 vdd.n2448 vdd.n2447 185
R15888 vdd.n2447 vdd.n721 185
R15889 vdd.n2446 vdd.n719 185
R15890 vdd.n2600 vdd.n719 185
R15891 vdd.n2445 vdd.n2444 185
R15892 vdd.n2444 vdd.n728 185
R15893 vdd.n2443 vdd.n726 185
R15894 vdd.n2594 vdd.n726 185
R15895 vdd.n2442 vdd.n2441 185
R15896 vdd.n2441 vdd.n725 185
R15897 vdd.n2353 vdd.n732 185
R15898 vdd.n2588 vdd.n732 185
R15899 vdd.n2495 vdd.n2494 185
R15900 vdd.n2494 vdd.n2493 185
R15901 vdd.n2496 vdd.n737 185
R15902 vdd.n2582 vdd.n737 185
R15903 vdd.n2498 vdd.n2497 185
R15904 vdd.n2497 vdd.t66 185
R15905 vdd.n2499 vdd.n742 185
R15906 vdd.n2576 vdd.n742 185
R15907 vdd.n2578 vdd.n2577 185
R15908 vdd.n2577 vdd.n2576 185
R15909 vdd.n2579 vdd.n739 185
R15910 vdd.n739 vdd.t66 185
R15911 vdd.n2581 vdd.n2580 185
R15912 vdd.n2582 vdd.n2581 185
R15913 vdd.n731 vdd.n730 185
R15914 vdd.n2493 vdd.n731 185
R15915 vdd.n2590 vdd.n2589 185
R15916 vdd.n2589 vdd.n2588 185
R15917 vdd.n2591 vdd.n729 185
R15918 vdd.n729 vdd.n725 185
R15919 vdd.n2593 vdd.n2592 185
R15920 vdd.n2594 vdd.n2593 185
R15921 vdd.n718 vdd.n717 185
R15922 vdd.n728 vdd.n718 185
R15923 vdd.n2602 vdd.n2601 185
R15924 vdd.n2601 vdd.n2600 185
R15925 vdd.n2603 vdd.n716 185
R15926 vdd.n721 vdd.n716 185
R15927 vdd.n2605 vdd.n2604 185
R15928 vdd.n2606 vdd.n2605 185
R15929 vdd.n707 vdd.n706 185
R15930 vdd.n708 vdd.n707 185
R15931 vdd.n2614 vdd.n2613 185
R15932 vdd.n2613 vdd.n2612 185
R15933 vdd.n2615 vdd.n705 185
R15934 vdd.n705 vdd.n702 185
R15935 vdd.n2617 vdd.n2616 185
R15936 vdd.n2618 vdd.n2617 185
R15937 vdd.n695 vdd.n694 185
R15938 vdd.n2472 vdd.n695 185
R15939 vdd.n2626 vdd.n2625 185
R15940 vdd.n2625 vdd.n2624 185
R15941 vdd.n2627 vdd.n693 185
R15942 vdd.n698 vdd.n693 185
R15943 vdd.n2629 vdd.n2628 185
R15944 vdd.n2630 vdd.n2629 185
R15945 vdd.n684 vdd.n683 185
R15946 vdd.n685 vdd.n684 185
R15947 vdd.n2640 vdd.n2639 185
R15948 vdd.n2639 vdd.n2638 185
R15949 vdd.n2641 vdd.n682 185
R15950 vdd.n682 vdd.n679 185
R15951 vdd.n2643 vdd.n2642 185
R15952 vdd.n2644 vdd.n2643 185
R15953 vdd.n670 vdd.n669 185
R15954 vdd.n671 vdd.n670 185
R15955 vdd.n2697 vdd.n2696 185
R15956 vdd.n2696 vdd.n2695 185
R15957 vdd.n2698 vdd.n668 185
R15958 vdd.n674 vdd.n668 185
R15959 vdd.n2700 vdd.n2699 185
R15960 vdd.n2701 vdd.n2700 185
R15961 vdd.n636 vdd.n634 185
R15962 vdd.n634 vdd.n631 185
R15963 vdd.n2770 vdd.n2769 185
R15964 vdd.n2771 vdd.n2770 185
R15965 vdd.n2243 vdd.n2242 185
R15966 vdd.n2244 vdd.n2243 185
R15967 vdd.n792 vdd.n790 185
R15968 vdd.n790 vdd.t159 185
R15969 vdd.n2158 vdd.n799 185
R15970 vdd.n2169 vdd.n799 185
R15971 vdd.n2159 vdd.n808 185
R15972 vdd.n1868 vdd.n808 185
R15973 vdd.n2161 vdd.n2160 185
R15974 vdd.n2162 vdd.n2161 185
R15975 vdd.n2157 vdd.n807 185
R15976 vdd.n807 vdd.n804 185
R15977 vdd.n2156 vdd.n2155 185
R15978 vdd.n2155 vdd.n2154 185
R15979 vdd.n810 vdd.n809 185
R15980 vdd.n811 vdd.n810 185
R15981 vdd.n2147 vdd.n2146 185
R15982 vdd.n2148 vdd.n2147 185
R15983 vdd.n2145 vdd.n820 185
R15984 vdd.n820 vdd.n817 185
R15985 vdd.n2144 vdd.n2143 185
R15986 vdd.n2143 vdd.n2142 185
R15987 vdd.n822 vdd.n821 185
R15988 vdd.n830 vdd.n822 185
R15989 vdd.n2135 vdd.n2134 185
R15990 vdd.n2136 vdd.n2135 185
R15991 vdd.n2133 vdd.n831 185
R15992 vdd.n836 vdd.n831 185
R15993 vdd.n2132 vdd.n2131 185
R15994 vdd.n2131 vdd.n2130 185
R15995 vdd.n833 vdd.n832 185
R15996 vdd.n1969 vdd.n833 185
R15997 vdd.n2123 vdd.n2122 185
R15998 vdd.n2124 vdd.n2123 185
R15999 vdd.n2121 vdd.n843 185
R16000 vdd.n843 vdd.n840 185
R16001 vdd.n2120 vdd.n2119 185
R16002 vdd.n2119 vdd.n2118 185
R16003 vdd.n845 vdd.n844 185
R16004 vdd.n846 vdd.n845 185
R16005 vdd.n2111 vdd.n2110 185
R16006 vdd.n2112 vdd.n2111 185
R16007 vdd.n2108 vdd.n854 185
R16008 vdd.n861 vdd.n854 185
R16009 vdd.n2107 vdd.n2106 185
R16010 vdd.n2106 vdd.n2105 185
R16011 vdd.n857 vdd.n856 185
R16012 vdd.n858 vdd.n857 185
R16013 vdd.n2098 vdd.n2097 185
R16014 vdd.n2099 vdd.n2098 185
R16015 vdd.n2096 vdd.n868 185
R16016 vdd.n868 vdd.n865 185
R16017 vdd.n2095 vdd.n2094 185
R16018 vdd.n2094 vdd.n2093 185
R16019 vdd.n870 vdd.n869 185
R16020 vdd.n871 vdd.n870 185
R16021 vdd.n2086 vdd.n2085 185
R16022 vdd.n2087 vdd.n2086 185
R16023 vdd.n2174 vdd.n764 185
R16024 vdd.n2316 vdd.n764 185
R16025 vdd.n2176 vdd.n2175 185
R16026 vdd.n2178 vdd.n2177 185
R16027 vdd.n2180 vdd.n2179 185
R16028 vdd.n2182 vdd.n2181 185
R16029 vdd.n2184 vdd.n2183 185
R16030 vdd.n2186 vdd.n2185 185
R16031 vdd.n2188 vdd.n2187 185
R16032 vdd.n2190 vdd.n2189 185
R16033 vdd.n2192 vdd.n2191 185
R16034 vdd.n2194 vdd.n2193 185
R16035 vdd.n2196 vdd.n2195 185
R16036 vdd.n2198 vdd.n2197 185
R16037 vdd.n2200 vdd.n2199 185
R16038 vdd.n2202 vdd.n2201 185
R16039 vdd.n2204 vdd.n2203 185
R16040 vdd.n2206 vdd.n2205 185
R16041 vdd.n2208 vdd.n2207 185
R16042 vdd.n2210 vdd.n2209 185
R16043 vdd.n2212 vdd.n2211 185
R16044 vdd.n2214 vdd.n2213 185
R16045 vdd.n2216 vdd.n2215 185
R16046 vdd.n2218 vdd.n2217 185
R16047 vdd.n2220 vdd.n2219 185
R16048 vdd.n2222 vdd.n2221 185
R16049 vdd.n2224 vdd.n2223 185
R16050 vdd.n2226 vdd.n2225 185
R16051 vdd.n2228 vdd.n2227 185
R16052 vdd.n2230 vdd.n2229 185
R16053 vdd.n2232 vdd.n2231 185
R16054 vdd.n2234 vdd.n2233 185
R16055 vdd.n2236 vdd.n2235 185
R16056 vdd.n2238 vdd.n2237 185
R16057 vdd.n2240 vdd.n2239 185
R16058 vdd.n2241 vdd.n791 185
R16059 vdd.n2173 vdd.n789 185
R16060 vdd.n2244 vdd.n789 185
R16061 vdd.n2172 vdd.n2171 185
R16062 vdd.n2171 vdd.t159 185
R16063 vdd.n2170 vdd.n796 185
R16064 vdd.n2170 vdd.n2169 185
R16065 vdd.n1950 vdd.n797 185
R16066 vdd.n1868 vdd.n797 185
R16067 vdd.n1951 vdd.n806 185
R16068 vdd.n2162 vdd.n806 185
R16069 vdd.n1953 vdd.n1952 185
R16070 vdd.n1952 vdd.n804 185
R16071 vdd.n1954 vdd.n813 185
R16072 vdd.n2154 vdd.n813 185
R16073 vdd.n1956 vdd.n1955 185
R16074 vdd.n1955 vdd.n811 185
R16075 vdd.n1957 vdd.n819 185
R16076 vdd.n2148 vdd.n819 185
R16077 vdd.n1959 vdd.n1958 185
R16078 vdd.n1958 vdd.n817 185
R16079 vdd.n1960 vdd.n824 185
R16080 vdd.n2142 vdd.n824 185
R16081 vdd.n1962 vdd.n1961 185
R16082 vdd.n1961 vdd.n830 185
R16083 vdd.n1963 vdd.n829 185
R16084 vdd.n2136 vdd.n829 185
R16085 vdd.n1965 vdd.n1964 185
R16086 vdd.n1964 vdd.n836 185
R16087 vdd.n1966 vdd.n835 185
R16088 vdd.n2130 vdd.n835 185
R16089 vdd.n1968 vdd.n1967 185
R16090 vdd.n1969 vdd.n1968 185
R16091 vdd.n1949 vdd.n842 185
R16092 vdd.n2124 vdd.n842 185
R16093 vdd.n1948 vdd.n1947 185
R16094 vdd.n1947 vdd.n840 185
R16095 vdd.n1946 vdd.n848 185
R16096 vdd.n2118 vdd.n848 185
R16097 vdd.n1945 vdd.n1944 185
R16098 vdd.n1944 vdd.n846 185
R16099 vdd.n1943 vdd.n853 185
R16100 vdd.n2112 vdd.n853 185
R16101 vdd.n1942 vdd.n1941 185
R16102 vdd.n1941 vdd.n861 185
R16103 vdd.n1940 vdd.n860 185
R16104 vdd.n2105 vdd.n860 185
R16105 vdd.n1939 vdd.n1938 185
R16106 vdd.n1938 vdd.n858 185
R16107 vdd.n1937 vdd.n867 185
R16108 vdd.n2099 vdd.n867 185
R16109 vdd.n1936 vdd.n1935 185
R16110 vdd.n1935 vdd.n865 185
R16111 vdd.n1934 vdd.n873 185
R16112 vdd.n2093 vdd.n873 185
R16113 vdd.n1933 vdd.n1932 185
R16114 vdd.n1932 vdd.n871 185
R16115 vdd.n1931 vdd.n879 185
R16116 vdd.n2087 vdd.n879 185
R16117 vdd.n2084 vdd.n880 185
R16118 vdd.n2083 vdd.n2082 185
R16119 vdd.n2080 vdd.n881 185
R16120 vdd.n2078 vdd.n2077 185
R16121 vdd.n2076 vdd.n882 185
R16122 vdd.n2075 vdd.n2074 185
R16123 vdd.n2072 vdd.n883 185
R16124 vdd.n2070 vdd.n2069 185
R16125 vdd.n2068 vdd.n884 185
R16126 vdd.n2067 vdd.n2066 185
R16127 vdd.n2064 vdd.n885 185
R16128 vdd.n2062 vdd.n2061 185
R16129 vdd.n2060 vdd.n886 185
R16130 vdd.n2059 vdd.n2058 185
R16131 vdd.n2056 vdd.n887 185
R16132 vdd.n2054 vdd.n2053 185
R16133 vdd.n2052 vdd.n888 185
R16134 vdd.n2051 vdd.n890 185
R16135 vdd.n1896 vdd.n891 185
R16136 vdd.n1899 vdd.n1898 185
R16137 vdd.n1901 vdd.n1900 185
R16138 vdd.n1903 vdd.n1895 185
R16139 vdd.n1906 vdd.n1905 185
R16140 vdd.n1907 vdd.n1894 185
R16141 vdd.n1909 vdd.n1908 185
R16142 vdd.n1911 vdd.n1893 185
R16143 vdd.n1914 vdd.n1913 185
R16144 vdd.n1915 vdd.n1892 185
R16145 vdd.n1917 vdd.n1916 185
R16146 vdd.n1919 vdd.n1891 185
R16147 vdd.n1922 vdd.n1921 185
R16148 vdd.n1923 vdd.n1888 185
R16149 vdd.n1926 vdd.n1925 185
R16150 vdd.n1928 vdd.n1887 185
R16151 vdd.n1930 vdd.n1929 185
R16152 vdd.n1929 vdd.n877 185
R16153 vdd.n303 vdd.n302 171.744
R16154 vdd.n302 vdd.n301 171.744
R16155 vdd.n301 vdd.n270 171.744
R16156 vdd.n294 vdd.n270 171.744
R16157 vdd.n294 vdd.n293 171.744
R16158 vdd.n293 vdd.n275 171.744
R16159 vdd.n286 vdd.n275 171.744
R16160 vdd.n286 vdd.n285 171.744
R16161 vdd.n285 vdd.n279 171.744
R16162 vdd.n252 vdd.n251 171.744
R16163 vdd.n251 vdd.n250 171.744
R16164 vdd.n250 vdd.n219 171.744
R16165 vdd.n243 vdd.n219 171.744
R16166 vdd.n243 vdd.n242 171.744
R16167 vdd.n242 vdd.n224 171.744
R16168 vdd.n235 vdd.n224 171.744
R16169 vdd.n235 vdd.n234 171.744
R16170 vdd.n234 vdd.n228 171.744
R16171 vdd.n209 vdd.n208 171.744
R16172 vdd.n208 vdd.n207 171.744
R16173 vdd.n207 vdd.n176 171.744
R16174 vdd.n200 vdd.n176 171.744
R16175 vdd.n200 vdd.n199 171.744
R16176 vdd.n199 vdd.n181 171.744
R16177 vdd.n192 vdd.n181 171.744
R16178 vdd.n192 vdd.n191 171.744
R16179 vdd.n191 vdd.n185 171.744
R16180 vdd.n158 vdd.n157 171.744
R16181 vdd.n157 vdd.n156 171.744
R16182 vdd.n156 vdd.n125 171.744
R16183 vdd.n149 vdd.n125 171.744
R16184 vdd.n149 vdd.n148 171.744
R16185 vdd.n148 vdd.n130 171.744
R16186 vdd.n141 vdd.n130 171.744
R16187 vdd.n141 vdd.n140 171.744
R16188 vdd.n140 vdd.n134 171.744
R16189 vdd.n116 vdd.n115 171.744
R16190 vdd.n115 vdd.n114 171.744
R16191 vdd.n114 vdd.n83 171.744
R16192 vdd.n107 vdd.n83 171.744
R16193 vdd.n107 vdd.n106 171.744
R16194 vdd.n106 vdd.n88 171.744
R16195 vdd.n99 vdd.n88 171.744
R16196 vdd.n99 vdd.n98 171.744
R16197 vdd.n98 vdd.n92 171.744
R16198 vdd.n65 vdd.n64 171.744
R16199 vdd.n64 vdd.n63 171.744
R16200 vdd.n63 vdd.n32 171.744
R16201 vdd.n56 vdd.n32 171.744
R16202 vdd.n56 vdd.n55 171.744
R16203 vdd.n55 vdd.n37 171.744
R16204 vdd.n48 vdd.n37 171.744
R16205 vdd.n48 vdd.n47 171.744
R16206 vdd.n47 vdd.n41 171.744
R16207 vdd.n1498 vdd.n1497 171.744
R16208 vdd.n1497 vdd.n1496 171.744
R16209 vdd.n1496 vdd.n1465 171.744
R16210 vdd.n1489 vdd.n1465 171.744
R16211 vdd.n1489 vdd.n1488 171.744
R16212 vdd.n1488 vdd.n1470 171.744
R16213 vdd.n1481 vdd.n1470 171.744
R16214 vdd.n1481 vdd.n1480 171.744
R16215 vdd.n1480 vdd.n1474 171.744
R16216 vdd.n1549 vdd.n1548 171.744
R16217 vdd.n1548 vdd.n1547 171.744
R16218 vdd.n1547 vdd.n1516 171.744
R16219 vdd.n1540 vdd.n1516 171.744
R16220 vdd.n1540 vdd.n1539 171.744
R16221 vdd.n1539 vdd.n1521 171.744
R16222 vdd.n1532 vdd.n1521 171.744
R16223 vdd.n1532 vdd.n1531 171.744
R16224 vdd.n1531 vdd.n1525 171.744
R16225 vdd.n1404 vdd.n1403 171.744
R16226 vdd.n1403 vdd.n1402 171.744
R16227 vdd.n1402 vdd.n1371 171.744
R16228 vdd.n1395 vdd.n1371 171.744
R16229 vdd.n1395 vdd.n1394 171.744
R16230 vdd.n1394 vdd.n1376 171.744
R16231 vdd.n1387 vdd.n1376 171.744
R16232 vdd.n1387 vdd.n1386 171.744
R16233 vdd.n1386 vdd.n1380 171.744
R16234 vdd.n1455 vdd.n1454 171.744
R16235 vdd.n1454 vdd.n1453 171.744
R16236 vdd.n1453 vdd.n1422 171.744
R16237 vdd.n1446 vdd.n1422 171.744
R16238 vdd.n1446 vdd.n1445 171.744
R16239 vdd.n1445 vdd.n1427 171.744
R16240 vdd.n1438 vdd.n1427 171.744
R16241 vdd.n1438 vdd.n1437 171.744
R16242 vdd.n1437 vdd.n1431 171.744
R16243 vdd.n1311 vdd.n1310 171.744
R16244 vdd.n1310 vdd.n1309 171.744
R16245 vdd.n1309 vdd.n1278 171.744
R16246 vdd.n1302 vdd.n1278 171.744
R16247 vdd.n1302 vdd.n1301 171.744
R16248 vdd.n1301 vdd.n1283 171.744
R16249 vdd.n1294 vdd.n1283 171.744
R16250 vdd.n1294 vdd.n1293 171.744
R16251 vdd.n1293 vdd.n1287 171.744
R16252 vdd.n1362 vdd.n1361 171.744
R16253 vdd.n1361 vdd.n1360 171.744
R16254 vdd.n1360 vdd.n1329 171.744
R16255 vdd.n1353 vdd.n1329 171.744
R16256 vdd.n1353 vdd.n1352 171.744
R16257 vdd.n1352 vdd.n1334 171.744
R16258 vdd.n1345 vdd.n1334 171.744
R16259 vdd.n1345 vdd.n1344 171.744
R16260 vdd.n1344 vdd.n1338 171.744
R16261 vdd.n3130 vdd.n356 146.341
R16262 vdd.n3128 vdd.n3127 146.341
R16263 vdd.n3125 vdd.n360 146.341
R16264 vdd.n3121 vdd.n3120 146.341
R16265 vdd.n3118 vdd.n368 146.341
R16266 vdd.n3114 vdd.n3113 146.341
R16267 vdd.n3111 vdd.n375 146.341
R16268 vdd.n3107 vdd.n3106 146.341
R16269 vdd.n3104 vdd.n382 146.341
R16270 vdd.n393 vdd.n390 146.341
R16271 vdd.n3096 vdd.n3095 146.341
R16272 vdd.n3093 vdd.n395 146.341
R16273 vdd.n3089 vdd.n3088 146.341
R16274 vdd.n3086 vdd.n401 146.341
R16275 vdd.n3082 vdd.n3081 146.341
R16276 vdd.n3079 vdd.n408 146.341
R16277 vdd.n3075 vdd.n3074 146.341
R16278 vdd.n3072 vdd.n415 146.341
R16279 vdd.n3068 vdd.n3067 146.341
R16280 vdd.n3065 vdd.n422 146.341
R16281 vdd.n433 vdd.n430 146.341
R16282 vdd.n3057 vdd.n3056 146.341
R16283 vdd.n3054 vdd.n435 146.341
R16284 vdd.n3050 vdd.n3049 146.341
R16285 vdd.n3047 vdd.n441 146.341
R16286 vdd.n3043 vdd.n3042 146.341
R16287 vdd.n3040 vdd.n448 146.341
R16288 vdd.n3036 vdd.n3035 146.341
R16289 vdd.n3033 vdd.n455 146.341
R16290 vdd.n3029 vdd.n3028 146.341
R16291 vdd.n3026 vdd.n462 146.341
R16292 vdd.n2941 vdd.n512 146.341
R16293 vdd.n2947 vdd.n512 146.341
R16294 vdd.n2947 vdd.n504 146.341
R16295 vdd.n2957 vdd.n504 146.341
R16296 vdd.n2957 vdd.n500 146.341
R16297 vdd.n2963 vdd.n500 146.341
R16298 vdd.n2963 vdd.n491 146.341
R16299 vdd.n2973 vdd.n491 146.341
R16300 vdd.n2973 vdd.n487 146.341
R16301 vdd.n2979 vdd.n487 146.341
R16302 vdd.n2979 vdd.n479 146.341
R16303 vdd.n2990 vdd.n479 146.341
R16304 vdd.n2990 vdd.n480 146.341
R16305 vdd.n480 vdd.n316 146.341
R16306 vdd.n317 vdd.n316 146.341
R16307 vdd.n318 vdd.n317 146.341
R16308 vdd.n473 vdd.n318 146.341
R16309 vdd.n473 vdd.n326 146.341
R16310 vdd.n327 vdd.n326 146.341
R16311 vdd.n328 vdd.n327 146.341
R16312 vdd.n470 vdd.n328 146.341
R16313 vdd.n470 vdd.n337 146.341
R16314 vdd.n338 vdd.n337 146.341
R16315 vdd.n339 vdd.n338 146.341
R16316 vdd.n467 vdd.n339 146.341
R16317 vdd.n467 vdd.n348 146.341
R16318 vdd.n349 vdd.n348 146.341
R16319 vdd.n350 vdd.n349 146.341
R16320 vdd.n2933 vdd.n2931 146.341
R16321 vdd.n2931 vdd.n2930 146.341
R16322 vdd.n2927 vdd.n2926 146.341
R16323 vdd.n2923 vdd.n2922 146.341
R16324 vdd.n2920 vdd.n526 146.341
R16325 vdd.n2916 vdd.n2914 146.341
R16326 vdd.n2912 vdd.n532 146.341
R16327 vdd.n2908 vdd.n2906 146.341
R16328 vdd.n2904 vdd.n538 146.341
R16329 vdd.n2900 vdd.n2898 146.341
R16330 vdd.n2896 vdd.n546 146.341
R16331 vdd.n2892 vdd.n2890 146.341
R16332 vdd.n2888 vdd.n552 146.341
R16333 vdd.n2884 vdd.n2882 146.341
R16334 vdd.n2880 vdd.n558 146.341
R16335 vdd.n2876 vdd.n2874 146.341
R16336 vdd.n2872 vdd.n564 146.341
R16337 vdd.n2868 vdd.n2866 146.341
R16338 vdd.n2864 vdd.n570 146.341
R16339 vdd.n2860 vdd.n2858 146.341
R16340 vdd.n2856 vdd.n576 146.341
R16341 vdd.n2849 vdd.n585 146.341
R16342 vdd.n2847 vdd.n2846 146.341
R16343 vdd.n2843 vdd.n2842 146.341
R16344 vdd.n2840 vdd.n590 146.341
R16345 vdd.n2836 vdd.n2834 146.341
R16346 vdd.n2832 vdd.n596 146.341
R16347 vdd.n2828 vdd.n2826 146.341
R16348 vdd.n2824 vdd.n602 146.341
R16349 vdd.n2820 vdd.n2818 146.341
R16350 vdd.n2815 vdd.n2814 146.341
R16351 vdd.n2811 vdd.n515 146.341
R16352 vdd.n2939 vdd.n510 146.341
R16353 vdd.n2949 vdd.n510 146.341
R16354 vdd.n2949 vdd.n506 146.341
R16355 vdd.n2955 vdd.n506 146.341
R16356 vdd.n2955 vdd.n498 146.341
R16357 vdd.n2965 vdd.n498 146.341
R16358 vdd.n2965 vdd.n494 146.341
R16359 vdd.n2971 vdd.n494 146.341
R16360 vdd.n2971 vdd.n486 146.341
R16361 vdd.n2982 vdd.n486 146.341
R16362 vdd.n2982 vdd.n482 146.341
R16363 vdd.n2988 vdd.n482 146.341
R16364 vdd.n2988 vdd.n314 146.341
R16365 vdd.n3165 vdd.n314 146.341
R16366 vdd.n3165 vdd.n315 146.341
R16367 vdd.n3161 vdd.n315 146.341
R16368 vdd.n3161 vdd.n319 146.341
R16369 vdd.n3157 vdd.n319 146.341
R16370 vdd.n3157 vdd.n324 146.341
R16371 vdd.n3153 vdd.n324 146.341
R16372 vdd.n3153 vdd.n330 146.341
R16373 vdd.n3149 vdd.n330 146.341
R16374 vdd.n3149 vdd.n336 146.341
R16375 vdd.n3145 vdd.n336 146.341
R16376 vdd.n3145 vdd.n341 146.341
R16377 vdd.n3141 vdd.n341 146.341
R16378 vdd.n3141 vdd.n347 146.341
R16379 vdd.n3137 vdd.n347 146.341
R16380 vdd.n2034 vdd.n2033 146.341
R16381 vdd.n2031 vdd.n1615 146.341
R16382 vdd.n1811 vdd.n1621 146.341
R16383 vdd.n1809 vdd.n1808 146.341
R16384 vdd.n1806 vdd.n1623 146.341
R16385 vdd.n1802 vdd.n1801 146.341
R16386 vdd.n1799 vdd.n1630 146.341
R16387 vdd.n1795 vdd.n1794 146.341
R16388 vdd.n1792 vdd.n1637 146.341
R16389 vdd.n1648 vdd.n1645 146.341
R16390 vdd.n1784 vdd.n1783 146.341
R16391 vdd.n1781 vdd.n1650 146.341
R16392 vdd.n1777 vdd.n1776 146.341
R16393 vdd.n1774 vdd.n1656 146.341
R16394 vdd.n1770 vdd.n1769 146.341
R16395 vdd.n1767 vdd.n1663 146.341
R16396 vdd.n1763 vdd.n1762 146.341
R16397 vdd.n1760 vdd.n1670 146.341
R16398 vdd.n1756 vdd.n1755 146.341
R16399 vdd.n1753 vdd.n1677 146.341
R16400 vdd.n1688 vdd.n1685 146.341
R16401 vdd.n1745 vdd.n1744 146.341
R16402 vdd.n1742 vdd.n1690 146.341
R16403 vdd.n1738 vdd.n1737 146.341
R16404 vdd.n1735 vdd.n1696 146.341
R16405 vdd.n1731 vdd.n1730 146.341
R16406 vdd.n1728 vdd.n1703 146.341
R16407 vdd.n1724 vdd.n1723 146.341
R16408 vdd.n1721 vdd.n1718 146.341
R16409 vdd.n1716 vdd.n1713 146.341
R16410 vdd.n1711 vdd.n897 146.341
R16411 vdd.n1216 vdd.n978 146.341
R16412 vdd.n1222 vdd.n978 146.341
R16413 vdd.n1222 vdd.n971 146.341
R16414 vdd.n1232 vdd.n971 146.341
R16415 vdd.n1232 vdd.n967 146.341
R16416 vdd.n1238 vdd.n967 146.341
R16417 vdd.n1238 vdd.n958 146.341
R16418 vdd.n1248 vdd.n958 146.341
R16419 vdd.n1248 vdd.n954 146.341
R16420 vdd.n1254 vdd.n954 146.341
R16421 vdd.n1254 vdd.n947 146.341
R16422 vdd.n1265 vdd.n947 146.341
R16423 vdd.n1265 vdd.n943 146.341
R16424 vdd.n1271 vdd.n943 146.341
R16425 vdd.n1271 vdd.n936 146.341
R16426 vdd.n1563 vdd.n936 146.341
R16427 vdd.n1563 vdd.n932 146.341
R16428 vdd.n1569 vdd.n932 146.341
R16429 vdd.n1569 vdd.n924 146.341
R16430 vdd.n1580 vdd.n924 146.341
R16431 vdd.n1580 vdd.n920 146.341
R16432 vdd.n1586 vdd.n920 146.341
R16433 vdd.n1586 vdd.n914 146.341
R16434 vdd.n1597 vdd.n914 146.341
R16435 vdd.n1597 vdd.n909 146.341
R16436 vdd.n1605 vdd.n909 146.341
R16437 vdd.n1605 vdd.n899 146.341
R16438 vdd.n2042 vdd.n899 146.341
R16439 vdd.n988 vdd.n987 146.341
R16440 vdd.n991 vdd.n988 146.341
R16441 vdd.n994 vdd.n993 146.341
R16442 vdd.n999 vdd.n996 146.341
R16443 vdd.n1002 vdd.n1001 146.341
R16444 vdd.n1007 vdd.n1004 146.341
R16445 vdd.n1010 vdd.n1009 146.341
R16446 vdd.n1015 vdd.n1012 146.341
R16447 vdd.n1018 vdd.n1017 146.341
R16448 vdd.n1025 vdd.n1020 146.341
R16449 vdd.n1028 vdd.n1027 146.341
R16450 vdd.n1033 vdd.n1030 146.341
R16451 vdd.n1036 vdd.n1035 146.341
R16452 vdd.n1041 vdd.n1038 146.341
R16453 vdd.n1044 vdd.n1043 146.341
R16454 vdd.n1049 vdd.n1046 146.341
R16455 vdd.n1052 vdd.n1051 146.341
R16456 vdd.n1057 vdd.n1054 146.341
R16457 vdd.n1060 vdd.n1059 146.341
R16458 vdd.n1065 vdd.n1062 146.341
R16459 vdd.n1146 vdd.n1067 146.341
R16460 vdd.n1144 vdd.n1143 146.341
R16461 vdd.n1074 vdd.n1073 146.341
R16462 vdd.n1077 vdd.n1076 146.341
R16463 vdd.n1082 vdd.n1081 146.341
R16464 vdd.n1085 vdd.n1084 146.341
R16465 vdd.n1090 vdd.n1089 146.341
R16466 vdd.n1093 vdd.n1092 146.341
R16467 vdd.n1098 vdd.n1097 146.341
R16468 vdd.n1101 vdd.n1100 146.341
R16469 vdd.n1106 vdd.n1105 146.341
R16470 vdd.n1108 vdd.n981 146.341
R16471 vdd.n1214 vdd.n977 146.341
R16472 vdd.n1224 vdd.n977 146.341
R16473 vdd.n1224 vdd.n973 146.341
R16474 vdd.n1230 vdd.n973 146.341
R16475 vdd.n1230 vdd.n965 146.341
R16476 vdd.n1240 vdd.n965 146.341
R16477 vdd.n1240 vdd.n961 146.341
R16478 vdd.n1246 vdd.n961 146.341
R16479 vdd.n1246 vdd.n953 146.341
R16480 vdd.n1257 vdd.n953 146.341
R16481 vdd.n1257 vdd.n949 146.341
R16482 vdd.n1263 vdd.n949 146.341
R16483 vdd.n1263 vdd.n942 146.341
R16484 vdd.n1273 vdd.n942 146.341
R16485 vdd.n1273 vdd.n938 146.341
R16486 vdd.n1561 vdd.n938 146.341
R16487 vdd.n1561 vdd.n930 146.341
R16488 vdd.n1572 vdd.n930 146.341
R16489 vdd.n1572 vdd.n926 146.341
R16490 vdd.n1578 vdd.n926 146.341
R16491 vdd.n1578 vdd.n919 146.341
R16492 vdd.n1589 vdd.n919 146.341
R16493 vdd.n1589 vdd.n915 146.341
R16494 vdd.n1595 vdd.n915 146.341
R16495 vdd.n1595 vdd.n907 146.341
R16496 vdd.n1608 vdd.n907 146.341
R16497 vdd.n1608 vdd.n902 146.341
R16498 vdd.n2040 vdd.n902 146.341
R16499 vdd.n901 vdd.n877 141.707
R16500 vdd.n613 vdd.n516 141.707
R16501 vdd.n1889 vdd.t122 127.284
R16502 vdd.n793 vdd.t106 127.284
R16503 vdd.n1863 vdd.t148 127.284
R16504 vdd.n785 vdd.t131 127.284
R16505 vdd.n2634 vdd.t93 127.284
R16506 vdd.n2634 vdd.t94 127.284
R16507 vdd.n2354 vdd.t129 127.284
R16508 vdd.n661 vdd.t110 127.284
R16509 vdd.n2351 vdd.t115 127.284
R16510 vdd.n625 vdd.t117 127.284
R16511 vdd.n855 vdd.t125 127.284
R16512 vdd.n855 vdd.t126 127.284
R16513 vdd.n22 vdd.n20 117.314
R16514 vdd.n17 vdd.n15 117.314
R16515 vdd.n27 vdd.n26 116.927
R16516 vdd.n24 vdd.n23 116.927
R16517 vdd.n22 vdd.n21 116.927
R16518 vdd.n17 vdd.n16 116.927
R16519 vdd.n19 vdd.n18 116.927
R16520 vdd.n27 vdd.n25 116.927
R16521 vdd.n1890 vdd.t121 111.188
R16522 vdd.n794 vdd.t107 111.188
R16523 vdd.n1864 vdd.t147 111.188
R16524 vdd.n786 vdd.t132 111.188
R16525 vdd.n2355 vdd.t128 111.188
R16526 vdd.n662 vdd.t111 111.188
R16527 vdd.n2352 vdd.t114 111.188
R16528 vdd.n626 vdd.t118 111.188
R16529 vdd.n2577 vdd.n739 99.5127
R16530 vdd.n2581 vdd.n739 99.5127
R16531 vdd.n2581 vdd.n731 99.5127
R16532 vdd.n2589 vdd.n731 99.5127
R16533 vdd.n2589 vdd.n729 99.5127
R16534 vdd.n2593 vdd.n729 99.5127
R16535 vdd.n2593 vdd.n718 99.5127
R16536 vdd.n2601 vdd.n718 99.5127
R16537 vdd.n2601 vdd.n716 99.5127
R16538 vdd.n2605 vdd.n716 99.5127
R16539 vdd.n2605 vdd.n707 99.5127
R16540 vdd.n2613 vdd.n707 99.5127
R16541 vdd.n2613 vdd.n705 99.5127
R16542 vdd.n2617 vdd.n705 99.5127
R16543 vdd.n2617 vdd.n695 99.5127
R16544 vdd.n2625 vdd.n695 99.5127
R16545 vdd.n2625 vdd.n693 99.5127
R16546 vdd.n2629 vdd.n693 99.5127
R16547 vdd.n2629 vdd.n684 99.5127
R16548 vdd.n2639 vdd.n684 99.5127
R16549 vdd.n2639 vdd.n682 99.5127
R16550 vdd.n2643 vdd.n682 99.5127
R16551 vdd.n2643 vdd.n670 99.5127
R16552 vdd.n2696 vdd.n670 99.5127
R16553 vdd.n2696 vdd.n668 99.5127
R16554 vdd.n2700 vdd.n668 99.5127
R16555 vdd.n2700 vdd.n634 99.5127
R16556 vdd.n2770 vdd.n634 99.5127
R16557 vdd.n2766 vdd.n635 99.5127
R16558 vdd.n2764 vdd.n2763 99.5127
R16559 vdd.n2761 vdd.n639 99.5127
R16560 vdd.n2757 vdd.n2756 99.5127
R16561 vdd.n2754 vdd.n642 99.5127
R16562 vdd.n2750 vdd.n2749 99.5127
R16563 vdd.n2747 vdd.n645 99.5127
R16564 vdd.n2743 vdd.n2742 99.5127
R16565 vdd.n2740 vdd.n648 99.5127
R16566 vdd.n2735 vdd.n2734 99.5127
R16567 vdd.n2732 vdd.n651 99.5127
R16568 vdd.n2728 vdd.n2727 99.5127
R16569 vdd.n2725 vdd.n654 99.5127
R16570 vdd.n2721 vdd.n2720 99.5127
R16571 vdd.n2718 vdd.n657 99.5127
R16572 vdd.n2714 vdd.n2713 99.5127
R16573 vdd.n2711 vdd.n660 99.5127
R16574 vdd.n2497 vdd.n742 99.5127
R16575 vdd.n2497 vdd.n737 99.5127
R16576 vdd.n2494 vdd.n737 99.5127
R16577 vdd.n2494 vdd.n732 99.5127
R16578 vdd.n2441 vdd.n732 99.5127
R16579 vdd.n2441 vdd.n726 99.5127
R16580 vdd.n2444 vdd.n726 99.5127
R16581 vdd.n2444 vdd.n719 99.5127
R16582 vdd.n2447 vdd.n719 99.5127
R16583 vdd.n2447 vdd.n714 99.5127
R16584 vdd.n2450 vdd.n714 99.5127
R16585 vdd.n2450 vdd.n709 99.5127
R16586 vdd.n2453 vdd.n709 99.5127
R16587 vdd.n2453 vdd.n703 99.5127
R16588 vdd.n2471 vdd.n703 99.5127
R16589 vdd.n2471 vdd.n696 99.5127
R16590 vdd.n2467 vdd.n696 99.5127
R16591 vdd.n2467 vdd.n691 99.5127
R16592 vdd.n2464 vdd.n691 99.5127
R16593 vdd.n2464 vdd.n686 99.5127
R16594 vdd.n2461 vdd.n686 99.5127
R16595 vdd.n2461 vdd.n680 99.5127
R16596 vdd.n2458 vdd.n680 99.5127
R16597 vdd.n2458 vdd.n672 99.5127
R16598 vdd.n672 vdd.n665 99.5127
R16599 vdd.n2702 vdd.n665 99.5127
R16600 vdd.n2703 vdd.n2702 99.5127
R16601 vdd.n2703 vdd.n632 99.5127
R16602 vdd.n2567 vdd.n2350 99.5127
R16603 vdd.n2563 vdd.n2350 99.5127
R16604 vdd.n2561 vdd.n2560 99.5127
R16605 vdd.n2557 vdd.n2556 99.5127
R16606 vdd.n2553 vdd.n2552 99.5127
R16607 vdd.n2549 vdd.n2548 99.5127
R16608 vdd.n2545 vdd.n2544 99.5127
R16609 vdd.n2541 vdd.n2540 99.5127
R16610 vdd.n2537 vdd.n2536 99.5127
R16611 vdd.n2533 vdd.n2532 99.5127
R16612 vdd.n2529 vdd.n2528 99.5127
R16613 vdd.n2525 vdd.n2524 99.5127
R16614 vdd.n2521 vdd.n2520 99.5127
R16615 vdd.n2517 vdd.n2516 99.5127
R16616 vdd.n2513 vdd.n2512 99.5127
R16617 vdd.n2509 vdd.n2508 99.5127
R16618 vdd.n2504 vdd.n2503 99.5127
R16619 vdd.n2315 vdd.n783 99.5127
R16620 vdd.n2311 vdd.n2310 99.5127
R16621 vdd.n2307 vdd.n2306 99.5127
R16622 vdd.n2303 vdd.n2302 99.5127
R16623 vdd.n2299 vdd.n2298 99.5127
R16624 vdd.n2295 vdd.n2294 99.5127
R16625 vdd.n2291 vdd.n2290 99.5127
R16626 vdd.n2287 vdd.n2286 99.5127
R16627 vdd.n2283 vdd.n2282 99.5127
R16628 vdd.n2279 vdd.n2278 99.5127
R16629 vdd.n2275 vdd.n2274 99.5127
R16630 vdd.n2271 vdd.n2270 99.5127
R16631 vdd.n2267 vdd.n2266 99.5127
R16632 vdd.n2263 vdd.n2262 99.5127
R16633 vdd.n2259 vdd.n2258 99.5127
R16634 vdd.n2255 vdd.n2254 99.5127
R16635 vdd.n2250 vdd.n2249 99.5127
R16636 vdd.n1988 vdd.n878 99.5127
R16637 vdd.n1988 vdd.n872 99.5127
R16638 vdd.n1985 vdd.n872 99.5127
R16639 vdd.n1985 vdd.n866 99.5127
R16640 vdd.n1982 vdd.n866 99.5127
R16641 vdd.n1982 vdd.n859 99.5127
R16642 vdd.n1979 vdd.n859 99.5127
R16643 vdd.n1979 vdd.n852 99.5127
R16644 vdd.n1976 vdd.n852 99.5127
R16645 vdd.n1976 vdd.n847 99.5127
R16646 vdd.n1973 vdd.n847 99.5127
R16647 vdd.n1973 vdd.n841 99.5127
R16648 vdd.n1970 vdd.n841 99.5127
R16649 vdd.n1970 vdd.n834 99.5127
R16650 vdd.n1884 vdd.n834 99.5127
R16651 vdd.n1884 vdd.n828 99.5127
R16652 vdd.n1881 vdd.n828 99.5127
R16653 vdd.n1881 vdd.n823 99.5127
R16654 vdd.n1878 vdd.n823 99.5127
R16655 vdd.n1878 vdd.n818 99.5127
R16656 vdd.n1875 vdd.n818 99.5127
R16657 vdd.n1875 vdd.n812 99.5127
R16658 vdd.n1872 vdd.n812 99.5127
R16659 vdd.n1872 vdd.n805 99.5127
R16660 vdd.n1869 vdd.n805 99.5127
R16661 vdd.n1869 vdd.n798 99.5127
R16662 vdd.n798 vdd.n788 99.5127
R16663 vdd.n2245 vdd.n788 99.5127
R16664 vdd.n1823 vdd.n1821 99.5127
R16665 vdd.n1827 vdd.n1821 99.5127
R16666 vdd.n1831 vdd.n1829 99.5127
R16667 vdd.n1835 vdd.n1819 99.5127
R16668 vdd.n1839 vdd.n1837 99.5127
R16669 vdd.n1843 vdd.n1817 99.5127
R16670 vdd.n1847 vdd.n1845 99.5127
R16671 vdd.n1851 vdd.n1815 99.5127
R16672 vdd.n1854 vdd.n1853 99.5127
R16673 vdd.n2024 vdd.n2022 99.5127
R16674 vdd.n2020 vdd.n1856 99.5127
R16675 vdd.n2016 vdd.n2014 99.5127
R16676 vdd.n2012 vdd.n1858 99.5127
R16677 vdd.n2008 vdd.n2006 99.5127
R16678 vdd.n2004 vdd.n1860 99.5127
R16679 vdd.n2000 vdd.n1998 99.5127
R16680 vdd.n1996 vdd.n1862 99.5127
R16681 vdd.n2088 vdd.n874 99.5127
R16682 vdd.n2092 vdd.n874 99.5127
R16683 vdd.n2092 vdd.n864 99.5127
R16684 vdd.n2100 vdd.n864 99.5127
R16685 vdd.n2100 vdd.n862 99.5127
R16686 vdd.n2104 vdd.n862 99.5127
R16687 vdd.n2104 vdd.n851 99.5127
R16688 vdd.n2113 vdd.n851 99.5127
R16689 vdd.n2113 vdd.n849 99.5127
R16690 vdd.n2117 vdd.n849 99.5127
R16691 vdd.n2117 vdd.n839 99.5127
R16692 vdd.n2125 vdd.n839 99.5127
R16693 vdd.n2125 vdd.n837 99.5127
R16694 vdd.n2129 vdd.n837 99.5127
R16695 vdd.n2129 vdd.n827 99.5127
R16696 vdd.n2137 vdd.n827 99.5127
R16697 vdd.n2137 vdd.n825 99.5127
R16698 vdd.n2141 vdd.n825 99.5127
R16699 vdd.n2141 vdd.n816 99.5127
R16700 vdd.n2149 vdd.n816 99.5127
R16701 vdd.n2149 vdd.n814 99.5127
R16702 vdd.n2153 vdd.n814 99.5127
R16703 vdd.n2153 vdd.n803 99.5127
R16704 vdd.n2163 vdd.n803 99.5127
R16705 vdd.n2163 vdd.n800 99.5127
R16706 vdd.n2168 vdd.n800 99.5127
R16707 vdd.n2168 vdd.n801 99.5127
R16708 vdd.n801 vdd.n782 99.5127
R16709 vdd.n2686 vdd.n2685 99.5127
R16710 vdd.n2683 vdd.n2649 99.5127
R16711 vdd.n2679 vdd.n2678 99.5127
R16712 vdd.n2676 vdd.n2652 99.5127
R16713 vdd.n2672 vdd.n2671 99.5127
R16714 vdd.n2669 vdd.n2655 99.5127
R16715 vdd.n2665 vdd.n2664 99.5127
R16716 vdd.n2662 vdd.n2659 99.5127
R16717 vdd.n2803 vdd.n612 99.5127
R16718 vdd.n2801 vdd.n2800 99.5127
R16719 vdd.n2798 vdd.n615 99.5127
R16720 vdd.n2794 vdd.n2793 99.5127
R16721 vdd.n2791 vdd.n618 99.5127
R16722 vdd.n2787 vdd.n2786 99.5127
R16723 vdd.n2784 vdd.n621 99.5127
R16724 vdd.n2780 vdd.n2779 99.5127
R16725 vdd.n2777 vdd.n624 99.5127
R16726 vdd.n2421 vdd.n743 99.5127
R16727 vdd.n2421 vdd.n738 99.5127
R16728 vdd.n2492 vdd.n738 99.5127
R16729 vdd.n2492 vdd.n733 99.5127
R16730 vdd.n2488 vdd.n733 99.5127
R16731 vdd.n2488 vdd.n727 99.5127
R16732 vdd.n2485 vdd.n727 99.5127
R16733 vdd.n2485 vdd.n720 99.5127
R16734 vdd.n2482 vdd.n720 99.5127
R16735 vdd.n2482 vdd.n715 99.5127
R16736 vdd.n2479 vdd.n715 99.5127
R16737 vdd.n2479 vdd.n710 99.5127
R16738 vdd.n2476 vdd.n710 99.5127
R16739 vdd.n2476 vdd.n704 99.5127
R16740 vdd.n2473 vdd.n704 99.5127
R16741 vdd.n2473 vdd.n697 99.5127
R16742 vdd.n2438 vdd.n697 99.5127
R16743 vdd.n2438 vdd.n692 99.5127
R16744 vdd.n2435 vdd.n692 99.5127
R16745 vdd.n2435 vdd.n687 99.5127
R16746 vdd.n2432 vdd.n687 99.5127
R16747 vdd.n2432 vdd.n681 99.5127
R16748 vdd.n2429 vdd.n681 99.5127
R16749 vdd.n2429 vdd.n673 99.5127
R16750 vdd.n2426 vdd.n673 99.5127
R16751 vdd.n2426 vdd.n666 99.5127
R16752 vdd.n666 vdd.n630 99.5127
R16753 vdd.n2772 vdd.n630 99.5127
R16754 vdd.n2571 vdd.n746 99.5127
R16755 vdd.n2359 vdd.n2358 99.5127
R16756 vdd.n2363 vdd.n2362 99.5127
R16757 vdd.n2367 vdd.n2366 99.5127
R16758 vdd.n2371 vdd.n2370 99.5127
R16759 vdd.n2375 vdd.n2374 99.5127
R16760 vdd.n2379 vdd.n2378 99.5127
R16761 vdd.n2383 vdd.n2382 99.5127
R16762 vdd.n2387 vdd.n2386 99.5127
R16763 vdd.n2391 vdd.n2390 99.5127
R16764 vdd.n2395 vdd.n2394 99.5127
R16765 vdd.n2399 vdd.n2398 99.5127
R16766 vdd.n2403 vdd.n2402 99.5127
R16767 vdd.n2407 vdd.n2406 99.5127
R16768 vdd.n2411 vdd.n2410 99.5127
R16769 vdd.n2415 vdd.n2414 99.5127
R16770 vdd.n2417 vdd.n2349 99.5127
R16771 vdd.n2575 vdd.n736 99.5127
R16772 vdd.n2583 vdd.n736 99.5127
R16773 vdd.n2583 vdd.n734 99.5127
R16774 vdd.n2587 vdd.n734 99.5127
R16775 vdd.n2587 vdd.n724 99.5127
R16776 vdd.n2595 vdd.n724 99.5127
R16777 vdd.n2595 vdd.n722 99.5127
R16778 vdd.n2599 vdd.n722 99.5127
R16779 vdd.n2599 vdd.n713 99.5127
R16780 vdd.n2607 vdd.n713 99.5127
R16781 vdd.n2607 vdd.n711 99.5127
R16782 vdd.n2611 vdd.n711 99.5127
R16783 vdd.n2611 vdd.n701 99.5127
R16784 vdd.n2619 vdd.n701 99.5127
R16785 vdd.n2619 vdd.n699 99.5127
R16786 vdd.n2623 vdd.n699 99.5127
R16787 vdd.n2623 vdd.n690 99.5127
R16788 vdd.n2631 vdd.n690 99.5127
R16789 vdd.n2631 vdd.n688 99.5127
R16790 vdd.n2637 vdd.n688 99.5127
R16791 vdd.n2637 vdd.n678 99.5127
R16792 vdd.n2645 vdd.n678 99.5127
R16793 vdd.n2645 vdd.n675 99.5127
R16794 vdd.n2694 vdd.n675 99.5127
R16795 vdd.n2694 vdd.n676 99.5127
R16796 vdd.n676 vdd.n667 99.5127
R16797 vdd.n2689 vdd.n667 99.5127
R16798 vdd.n2689 vdd.n633 99.5127
R16799 vdd.n2239 vdd.n2238 99.5127
R16800 vdd.n2235 vdd.n2234 99.5127
R16801 vdd.n2231 vdd.n2230 99.5127
R16802 vdd.n2227 vdd.n2226 99.5127
R16803 vdd.n2223 vdd.n2222 99.5127
R16804 vdd.n2219 vdd.n2218 99.5127
R16805 vdd.n2215 vdd.n2214 99.5127
R16806 vdd.n2211 vdd.n2210 99.5127
R16807 vdd.n2207 vdd.n2206 99.5127
R16808 vdd.n2203 vdd.n2202 99.5127
R16809 vdd.n2199 vdd.n2198 99.5127
R16810 vdd.n2195 vdd.n2194 99.5127
R16811 vdd.n2191 vdd.n2190 99.5127
R16812 vdd.n2187 vdd.n2186 99.5127
R16813 vdd.n2183 vdd.n2182 99.5127
R16814 vdd.n2179 vdd.n2178 99.5127
R16815 vdd.n2175 vdd.n764 99.5127
R16816 vdd.n1932 vdd.n879 99.5127
R16817 vdd.n1932 vdd.n873 99.5127
R16818 vdd.n1935 vdd.n873 99.5127
R16819 vdd.n1935 vdd.n867 99.5127
R16820 vdd.n1938 vdd.n867 99.5127
R16821 vdd.n1938 vdd.n860 99.5127
R16822 vdd.n1941 vdd.n860 99.5127
R16823 vdd.n1941 vdd.n853 99.5127
R16824 vdd.n1944 vdd.n853 99.5127
R16825 vdd.n1944 vdd.n848 99.5127
R16826 vdd.n1947 vdd.n848 99.5127
R16827 vdd.n1947 vdd.n842 99.5127
R16828 vdd.n1968 vdd.n842 99.5127
R16829 vdd.n1968 vdd.n835 99.5127
R16830 vdd.n1964 vdd.n835 99.5127
R16831 vdd.n1964 vdd.n829 99.5127
R16832 vdd.n1961 vdd.n829 99.5127
R16833 vdd.n1961 vdd.n824 99.5127
R16834 vdd.n1958 vdd.n824 99.5127
R16835 vdd.n1958 vdd.n819 99.5127
R16836 vdd.n1955 vdd.n819 99.5127
R16837 vdd.n1955 vdd.n813 99.5127
R16838 vdd.n1952 vdd.n813 99.5127
R16839 vdd.n1952 vdd.n806 99.5127
R16840 vdd.n806 vdd.n797 99.5127
R16841 vdd.n2170 vdd.n797 99.5127
R16842 vdd.n2171 vdd.n2170 99.5127
R16843 vdd.n2171 vdd.n789 99.5127
R16844 vdd.n2082 vdd.n2080 99.5127
R16845 vdd.n2078 vdd.n882 99.5127
R16846 vdd.n2074 vdd.n2072 99.5127
R16847 vdd.n2070 vdd.n884 99.5127
R16848 vdd.n2066 vdd.n2064 99.5127
R16849 vdd.n2062 vdd.n886 99.5127
R16850 vdd.n2058 vdd.n2056 99.5127
R16851 vdd.n2054 vdd.n888 99.5127
R16852 vdd.n1896 vdd.n890 99.5127
R16853 vdd.n1901 vdd.n1898 99.5127
R16854 vdd.n1905 vdd.n1903 99.5127
R16855 vdd.n1909 vdd.n1894 99.5127
R16856 vdd.n1913 vdd.n1911 99.5127
R16857 vdd.n1917 vdd.n1892 99.5127
R16858 vdd.n1921 vdd.n1919 99.5127
R16859 vdd.n1926 vdd.n1888 99.5127
R16860 vdd.n1929 vdd.n1928 99.5127
R16861 vdd.n2086 vdd.n870 99.5127
R16862 vdd.n2094 vdd.n870 99.5127
R16863 vdd.n2094 vdd.n868 99.5127
R16864 vdd.n2098 vdd.n868 99.5127
R16865 vdd.n2098 vdd.n857 99.5127
R16866 vdd.n2106 vdd.n857 99.5127
R16867 vdd.n2106 vdd.n854 99.5127
R16868 vdd.n2111 vdd.n854 99.5127
R16869 vdd.n2111 vdd.n845 99.5127
R16870 vdd.n2119 vdd.n845 99.5127
R16871 vdd.n2119 vdd.n843 99.5127
R16872 vdd.n2123 vdd.n843 99.5127
R16873 vdd.n2123 vdd.n833 99.5127
R16874 vdd.n2131 vdd.n833 99.5127
R16875 vdd.n2131 vdd.n831 99.5127
R16876 vdd.n2135 vdd.n831 99.5127
R16877 vdd.n2135 vdd.n822 99.5127
R16878 vdd.n2143 vdd.n822 99.5127
R16879 vdd.n2143 vdd.n820 99.5127
R16880 vdd.n2147 vdd.n820 99.5127
R16881 vdd.n2147 vdd.n810 99.5127
R16882 vdd.n2155 vdd.n810 99.5127
R16883 vdd.n2155 vdd.n807 99.5127
R16884 vdd.n2161 vdd.n807 99.5127
R16885 vdd.n2161 vdd.n808 99.5127
R16886 vdd.n808 vdd.n799 99.5127
R16887 vdd.n799 vdd.n790 99.5127
R16888 vdd.n2243 vdd.n790 99.5127
R16889 vdd.n9 vdd.n7 98.9633
R16890 vdd.n2 vdd.n0 98.9633
R16891 vdd.n9 vdd.n8 98.6055
R16892 vdd.n11 vdd.n10 98.6055
R16893 vdd.n13 vdd.n12 98.6055
R16894 vdd.n6 vdd.n5 98.6055
R16895 vdd.n4 vdd.n3 98.6055
R16896 vdd.n2 vdd.n1 98.6055
R16897 vdd.t207 vdd.n279 85.8723
R16898 vdd.t42 vdd.n228 85.8723
R16899 vdd.t11 vdd.n185 85.8723
R16900 vdd.t72 vdd.n134 85.8723
R16901 vdd.t38 vdd.n92 85.8723
R16902 vdd.t16 vdd.n41 85.8723
R16903 vdd.t208 vdd.n1474 85.8723
R16904 vdd.t200 vdd.n1525 85.8723
R16905 vdd.t54 vdd.n1380 85.8723
R16906 vdd.t188 vdd.n1431 85.8723
R16907 vdd.t18 vdd.n1287 85.8723
R16908 vdd.t63 vdd.n1338 85.8723
R16909 vdd.n2635 vdd.n2634 78.546
R16910 vdd.n2109 vdd.n855 78.546
R16911 vdd.n266 vdd.n265 75.1835
R16912 vdd.n264 vdd.n263 75.1835
R16913 vdd.n262 vdd.n261 75.1835
R16914 vdd.n260 vdd.n259 75.1835
R16915 vdd.n258 vdd.n257 75.1835
R16916 vdd.n172 vdd.n171 75.1835
R16917 vdd.n170 vdd.n169 75.1835
R16918 vdd.n168 vdd.n167 75.1835
R16919 vdd.n166 vdd.n165 75.1835
R16920 vdd.n164 vdd.n163 75.1835
R16921 vdd.n79 vdd.n78 75.1835
R16922 vdd.n77 vdd.n76 75.1835
R16923 vdd.n75 vdd.n74 75.1835
R16924 vdd.n73 vdd.n72 75.1835
R16925 vdd.n71 vdd.n70 75.1835
R16926 vdd.n1504 vdd.n1503 75.1835
R16927 vdd.n1506 vdd.n1505 75.1835
R16928 vdd.n1508 vdd.n1507 75.1835
R16929 vdd.n1510 vdd.n1509 75.1835
R16930 vdd.n1512 vdd.n1511 75.1835
R16931 vdd.n1410 vdd.n1409 75.1835
R16932 vdd.n1412 vdd.n1411 75.1835
R16933 vdd.n1414 vdd.n1413 75.1835
R16934 vdd.n1416 vdd.n1415 75.1835
R16935 vdd.n1418 vdd.n1417 75.1835
R16936 vdd.n1317 vdd.n1316 75.1835
R16937 vdd.n1319 vdd.n1318 75.1835
R16938 vdd.n1321 vdd.n1320 75.1835
R16939 vdd.n1323 vdd.n1322 75.1835
R16940 vdd.n1325 vdd.n1324 75.1835
R16941 vdd.n2570 vdd.n2569 72.8958
R16942 vdd.n2569 vdd.n2333 72.8958
R16943 vdd.n2569 vdd.n2334 72.8958
R16944 vdd.n2569 vdd.n2335 72.8958
R16945 vdd.n2569 vdd.n2336 72.8958
R16946 vdd.n2569 vdd.n2337 72.8958
R16947 vdd.n2569 vdd.n2338 72.8958
R16948 vdd.n2569 vdd.n2339 72.8958
R16949 vdd.n2569 vdd.n2340 72.8958
R16950 vdd.n2569 vdd.n2341 72.8958
R16951 vdd.n2569 vdd.n2342 72.8958
R16952 vdd.n2569 vdd.n2343 72.8958
R16953 vdd.n2569 vdd.n2344 72.8958
R16954 vdd.n2569 vdd.n2345 72.8958
R16955 vdd.n2569 vdd.n2346 72.8958
R16956 vdd.n2569 vdd.n2347 72.8958
R16957 vdd.n2569 vdd.n2348 72.8958
R16958 vdd.n629 vdd.n613 72.8958
R16959 vdd.n2778 vdd.n613 72.8958
R16960 vdd.n623 vdd.n613 72.8958
R16961 vdd.n2785 vdd.n613 72.8958
R16962 vdd.n620 vdd.n613 72.8958
R16963 vdd.n2792 vdd.n613 72.8958
R16964 vdd.n617 vdd.n613 72.8958
R16965 vdd.n2799 vdd.n613 72.8958
R16966 vdd.n2802 vdd.n613 72.8958
R16967 vdd.n2658 vdd.n613 72.8958
R16968 vdd.n2663 vdd.n613 72.8958
R16969 vdd.n2657 vdd.n613 72.8958
R16970 vdd.n2670 vdd.n613 72.8958
R16971 vdd.n2654 vdd.n613 72.8958
R16972 vdd.n2677 vdd.n613 72.8958
R16973 vdd.n2651 vdd.n613 72.8958
R16974 vdd.n2684 vdd.n613 72.8958
R16975 vdd.n1822 vdd.n877 72.8958
R16976 vdd.n1828 vdd.n877 72.8958
R16977 vdd.n1830 vdd.n877 72.8958
R16978 vdd.n1836 vdd.n877 72.8958
R16979 vdd.n1838 vdd.n877 72.8958
R16980 vdd.n1844 vdd.n877 72.8958
R16981 vdd.n1846 vdd.n877 72.8958
R16982 vdd.n1852 vdd.n877 72.8958
R16983 vdd.n2023 vdd.n877 72.8958
R16984 vdd.n2021 vdd.n877 72.8958
R16985 vdd.n2015 vdd.n877 72.8958
R16986 vdd.n2013 vdd.n877 72.8958
R16987 vdd.n2007 vdd.n877 72.8958
R16988 vdd.n2005 vdd.n877 72.8958
R16989 vdd.n1999 vdd.n877 72.8958
R16990 vdd.n1997 vdd.n877 72.8958
R16991 vdd.n1991 vdd.n877 72.8958
R16992 vdd.n2316 vdd.n765 72.8958
R16993 vdd.n2316 vdd.n766 72.8958
R16994 vdd.n2316 vdd.n767 72.8958
R16995 vdd.n2316 vdd.n768 72.8958
R16996 vdd.n2316 vdd.n769 72.8958
R16997 vdd.n2316 vdd.n770 72.8958
R16998 vdd.n2316 vdd.n771 72.8958
R16999 vdd.n2316 vdd.n772 72.8958
R17000 vdd.n2316 vdd.n773 72.8958
R17001 vdd.n2316 vdd.n774 72.8958
R17002 vdd.n2316 vdd.n775 72.8958
R17003 vdd.n2316 vdd.n776 72.8958
R17004 vdd.n2316 vdd.n777 72.8958
R17005 vdd.n2316 vdd.n778 72.8958
R17006 vdd.n2316 vdd.n779 72.8958
R17007 vdd.n2316 vdd.n780 72.8958
R17008 vdd.n2316 vdd.n781 72.8958
R17009 vdd.n2569 vdd.n2568 72.8958
R17010 vdd.n2569 vdd.n2317 72.8958
R17011 vdd.n2569 vdd.n2318 72.8958
R17012 vdd.n2569 vdd.n2319 72.8958
R17013 vdd.n2569 vdd.n2320 72.8958
R17014 vdd.n2569 vdd.n2321 72.8958
R17015 vdd.n2569 vdd.n2322 72.8958
R17016 vdd.n2569 vdd.n2323 72.8958
R17017 vdd.n2569 vdd.n2324 72.8958
R17018 vdd.n2569 vdd.n2325 72.8958
R17019 vdd.n2569 vdd.n2326 72.8958
R17020 vdd.n2569 vdd.n2327 72.8958
R17021 vdd.n2569 vdd.n2328 72.8958
R17022 vdd.n2569 vdd.n2329 72.8958
R17023 vdd.n2569 vdd.n2330 72.8958
R17024 vdd.n2569 vdd.n2331 72.8958
R17025 vdd.n2569 vdd.n2332 72.8958
R17026 vdd.n2706 vdd.n613 72.8958
R17027 vdd.n2712 vdd.n613 72.8958
R17028 vdd.n659 vdd.n613 72.8958
R17029 vdd.n2719 vdd.n613 72.8958
R17030 vdd.n656 vdd.n613 72.8958
R17031 vdd.n2726 vdd.n613 72.8958
R17032 vdd.n653 vdd.n613 72.8958
R17033 vdd.n2733 vdd.n613 72.8958
R17034 vdd.n650 vdd.n613 72.8958
R17035 vdd.n2741 vdd.n613 72.8958
R17036 vdd.n647 vdd.n613 72.8958
R17037 vdd.n2748 vdd.n613 72.8958
R17038 vdd.n644 vdd.n613 72.8958
R17039 vdd.n2755 vdd.n613 72.8958
R17040 vdd.n641 vdd.n613 72.8958
R17041 vdd.n2762 vdd.n613 72.8958
R17042 vdd.n2765 vdd.n613 72.8958
R17043 vdd.n2316 vdd.n763 72.8958
R17044 vdd.n2316 vdd.n762 72.8958
R17045 vdd.n2316 vdd.n761 72.8958
R17046 vdd.n2316 vdd.n760 72.8958
R17047 vdd.n2316 vdd.n759 72.8958
R17048 vdd.n2316 vdd.n758 72.8958
R17049 vdd.n2316 vdd.n757 72.8958
R17050 vdd.n2316 vdd.n756 72.8958
R17051 vdd.n2316 vdd.n755 72.8958
R17052 vdd.n2316 vdd.n754 72.8958
R17053 vdd.n2316 vdd.n753 72.8958
R17054 vdd.n2316 vdd.n752 72.8958
R17055 vdd.n2316 vdd.n751 72.8958
R17056 vdd.n2316 vdd.n750 72.8958
R17057 vdd.n2316 vdd.n749 72.8958
R17058 vdd.n2316 vdd.n748 72.8958
R17059 vdd.n2316 vdd.n747 72.8958
R17060 vdd.n2081 vdd.n877 72.8958
R17061 vdd.n2079 vdd.n877 72.8958
R17062 vdd.n2073 vdd.n877 72.8958
R17063 vdd.n2071 vdd.n877 72.8958
R17064 vdd.n2065 vdd.n877 72.8958
R17065 vdd.n2063 vdd.n877 72.8958
R17066 vdd.n2057 vdd.n877 72.8958
R17067 vdd.n2055 vdd.n877 72.8958
R17068 vdd.n889 vdd.n877 72.8958
R17069 vdd.n1897 vdd.n877 72.8958
R17070 vdd.n1902 vdd.n877 72.8958
R17071 vdd.n1904 vdd.n877 72.8958
R17072 vdd.n1910 vdd.n877 72.8958
R17073 vdd.n1912 vdd.n877 72.8958
R17074 vdd.n1918 vdd.n877 72.8958
R17075 vdd.n1920 vdd.n877 72.8958
R17076 vdd.n1927 vdd.n877 72.8958
R17077 vdd.n986 vdd.n982 66.2847
R17078 vdd.n992 vdd.n982 66.2847
R17079 vdd.n995 vdd.n982 66.2847
R17080 vdd.n1000 vdd.n982 66.2847
R17081 vdd.n1003 vdd.n982 66.2847
R17082 vdd.n1008 vdd.n982 66.2847
R17083 vdd.n1011 vdd.n982 66.2847
R17084 vdd.n1016 vdd.n982 66.2847
R17085 vdd.n1019 vdd.n982 66.2847
R17086 vdd.n1026 vdd.n982 66.2847
R17087 vdd.n1029 vdd.n982 66.2847
R17088 vdd.n1034 vdd.n982 66.2847
R17089 vdd.n1037 vdd.n982 66.2847
R17090 vdd.n1042 vdd.n982 66.2847
R17091 vdd.n1045 vdd.n982 66.2847
R17092 vdd.n1050 vdd.n982 66.2847
R17093 vdd.n1053 vdd.n982 66.2847
R17094 vdd.n1058 vdd.n982 66.2847
R17095 vdd.n1061 vdd.n982 66.2847
R17096 vdd.n1066 vdd.n982 66.2847
R17097 vdd.n1145 vdd.n982 66.2847
R17098 vdd.n1069 vdd.n982 66.2847
R17099 vdd.n1075 vdd.n982 66.2847
R17100 vdd.n1080 vdd.n982 66.2847
R17101 vdd.n1083 vdd.n982 66.2847
R17102 vdd.n1088 vdd.n982 66.2847
R17103 vdd.n1091 vdd.n982 66.2847
R17104 vdd.n1096 vdd.n982 66.2847
R17105 vdd.n1099 vdd.n982 66.2847
R17106 vdd.n1104 vdd.n982 66.2847
R17107 vdd.n1107 vdd.n982 66.2847
R17108 vdd.n901 vdd.n898 66.2847
R17109 vdd.n1712 vdd.n901 66.2847
R17110 vdd.n1717 vdd.n901 66.2847
R17111 vdd.n1722 vdd.n901 66.2847
R17112 vdd.n1710 vdd.n901 66.2847
R17113 vdd.n1729 vdd.n901 66.2847
R17114 vdd.n1702 vdd.n901 66.2847
R17115 vdd.n1736 vdd.n901 66.2847
R17116 vdd.n1695 vdd.n901 66.2847
R17117 vdd.n1743 vdd.n901 66.2847
R17118 vdd.n1689 vdd.n901 66.2847
R17119 vdd.n1684 vdd.n901 66.2847
R17120 vdd.n1754 vdd.n901 66.2847
R17121 vdd.n1676 vdd.n901 66.2847
R17122 vdd.n1761 vdd.n901 66.2847
R17123 vdd.n1669 vdd.n901 66.2847
R17124 vdd.n1768 vdd.n901 66.2847
R17125 vdd.n1662 vdd.n901 66.2847
R17126 vdd.n1775 vdd.n901 66.2847
R17127 vdd.n1655 vdd.n901 66.2847
R17128 vdd.n1782 vdd.n901 66.2847
R17129 vdd.n1649 vdd.n901 66.2847
R17130 vdd.n1644 vdd.n901 66.2847
R17131 vdd.n1793 vdd.n901 66.2847
R17132 vdd.n1636 vdd.n901 66.2847
R17133 vdd.n1800 vdd.n901 66.2847
R17134 vdd.n1629 vdd.n901 66.2847
R17135 vdd.n1807 vdd.n901 66.2847
R17136 vdd.n1810 vdd.n901 66.2847
R17137 vdd.n1620 vdd.n901 66.2847
R17138 vdd.n2032 vdd.n901 66.2847
R17139 vdd.n1614 vdd.n901 66.2847
R17140 vdd.n2932 vdd.n516 66.2847
R17141 vdd.n520 vdd.n516 66.2847
R17142 vdd.n523 vdd.n516 66.2847
R17143 vdd.n2921 vdd.n516 66.2847
R17144 vdd.n2915 vdd.n516 66.2847
R17145 vdd.n2913 vdd.n516 66.2847
R17146 vdd.n2907 vdd.n516 66.2847
R17147 vdd.n2905 vdd.n516 66.2847
R17148 vdd.n2899 vdd.n516 66.2847
R17149 vdd.n2897 vdd.n516 66.2847
R17150 vdd.n2891 vdd.n516 66.2847
R17151 vdd.n2889 vdd.n516 66.2847
R17152 vdd.n2883 vdd.n516 66.2847
R17153 vdd.n2881 vdd.n516 66.2847
R17154 vdd.n2875 vdd.n516 66.2847
R17155 vdd.n2873 vdd.n516 66.2847
R17156 vdd.n2867 vdd.n516 66.2847
R17157 vdd.n2865 vdd.n516 66.2847
R17158 vdd.n2859 vdd.n516 66.2847
R17159 vdd.n2857 vdd.n516 66.2847
R17160 vdd.n584 vdd.n516 66.2847
R17161 vdd.n2848 vdd.n516 66.2847
R17162 vdd.n586 vdd.n516 66.2847
R17163 vdd.n2841 vdd.n516 66.2847
R17164 vdd.n2835 vdd.n516 66.2847
R17165 vdd.n2833 vdd.n516 66.2847
R17166 vdd.n2827 vdd.n516 66.2847
R17167 vdd.n2825 vdd.n516 66.2847
R17168 vdd.n2819 vdd.n516 66.2847
R17169 vdd.n607 vdd.n516 66.2847
R17170 vdd.n609 vdd.n516 66.2847
R17171 vdd.n3018 vdd.n351 66.2847
R17172 vdd.n3027 vdd.n351 66.2847
R17173 vdd.n461 vdd.n351 66.2847
R17174 vdd.n3034 vdd.n351 66.2847
R17175 vdd.n454 vdd.n351 66.2847
R17176 vdd.n3041 vdd.n351 66.2847
R17177 vdd.n447 vdd.n351 66.2847
R17178 vdd.n3048 vdd.n351 66.2847
R17179 vdd.n440 vdd.n351 66.2847
R17180 vdd.n3055 vdd.n351 66.2847
R17181 vdd.n434 vdd.n351 66.2847
R17182 vdd.n429 vdd.n351 66.2847
R17183 vdd.n3066 vdd.n351 66.2847
R17184 vdd.n421 vdd.n351 66.2847
R17185 vdd.n3073 vdd.n351 66.2847
R17186 vdd.n414 vdd.n351 66.2847
R17187 vdd.n3080 vdd.n351 66.2847
R17188 vdd.n407 vdd.n351 66.2847
R17189 vdd.n3087 vdd.n351 66.2847
R17190 vdd.n400 vdd.n351 66.2847
R17191 vdd.n3094 vdd.n351 66.2847
R17192 vdd.n394 vdd.n351 66.2847
R17193 vdd.n389 vdd.n351 66.2847
R17194 vdd.n3105 vdd.n351 66.2847
R17195 vdd.n381 vdd.n351 66.2847
R17196 vdd.n3112 vdd.n351 66.2847
R17197 vdd.n374 vdd.n351 66.2847
R17198 vdd.n3119 vdd.n351 66.2847
R17199 vdd.n367 vdd.n351 66.2847
R17200 vdd.n3126 vdd.n351 66.2847
R17201 vdd.n3129 vdd.n351 66.2847
R17202 vdd.n355 vdd.n351 66.2847
R17203 vdd.n356 vdd.n355 52.4337
R17204 vdd.n3129 vdd.n3128 52.4337
R17205 vdd.n3126 vdd.n3125 52.4337
R17206 vdd.n3121 vdd.n367 52.4337
R17207 vdd.n3119 vdd.n3118 52.4337
R17208 vdd.n3114 vdd.n374 52.4337
R17209 vdd.n3112 vdd.n3111 52.4337
R17210 vdd.n3107 vdd.n381 52.4337
R17211 vdd.n3105 vdd.n3104 52.4337
R17212 vdd.n390 vdd.n389 52.4337
R17213 vdd.n3096 vdd.n394 52.4337
R17214 vdd.n3094 vdd.n3093 52.4337
R17215 vdd.n3089 vdd.n400 52.4337
R17216 vdd.n3087 vdd.n3086 52.4337
R17217 vdd.n3082 vdd.n407 52.4337
R17218 vdd.n3080 vdd.n3079 52.4337
R17219 vdd.n3075 vdd.n414 52.4337
R17220 vdd.n3073 vdd.n3072 52.4337
R17221 vdd.n3068 vdd.n421 52.4337
R17222 vdd.n3066 vdd.n3065 52.4337
R17223 vdd.n430 vdd.n429 52.4337
R17224 vdd.n3057 vdd.n434 52.4337
R17225 vdd.n3055 vdd.n3054 52.4337
R17226 vdd.n3050 vdd.n440 52.4337
R17227 vdd.n3048 vdd.n3047 52.4337
R17228 vdd.n3043 vdd.n447 52.4337
R17229 vdd.n3041 vdd.n3040 52.4337
R17230 vdd.n3036 vdd.n454 52.4337
R17231 vdd.n3034 vdd.n3033 52.4337
R17232 vdd.n3029 vdd.n461 52.4337
R17233 vdd.n3027 vdd.n3026 52.4337
R17234 vdd.n3019 vdd.n3018 52.4337
R17235 vdd.n2932 vdd.n517 52.4337
R17236 vdd.n2930 vdd.n520 52.4337
R17237 vdd.n2926 vdd.n523 52.4337
R17238 vdd.n2922 vdd.n2921 52.4337
R17239 vdd.n2915 vdd.n526 52.4337
R17240 vdd.n2914 vdd.n2913 52.4337
R17241 vdd.n2907 vdd.n532 52.4337
R17242 vdd.n2906 vdd.n2905 52.4337
R17243 vdd.n2899 vdd.n538 52.4337
R17244 vdd.n2898 vdd.n2897 52.4337
R17245 vdd.n2891 vdd.n546 52.4337
R17246 vdd.n2890 vdd.n2889 52.4337
R17247 vdd.n2883 vdd.n552 52.4337
R17248 vdd.n2882 vdd.n2881 52.4337
R17249 vdd.n2875 vdd.n558 52.4337
R17250 vdd.n2874 vdd.n2873 52.4337
R17251 vdd.n2867 vdd.n564 52.4337
R17252 vdd.n2866 vdd.n2865 52.4337
R17253 vdd.n2859 vdd.n570 52.4337
R17254 vdd.n2858 vdd.n2857 52.4337
R17255 vdd.n584 vdd.n576 52.4337
R17256 vdd.n2849 vdd.n2848 52.4337
R17257 vdd.n2846 vdd.n586 52.4337
R17258 vdd.n2842 vdd.n2841 52.4337
R17259 vdd.n2835 vdd.n590 52.4337
R17260 vdd.n2834 vdd.n2833 52.4337
R17261 vdd.n2827 vdd.n596 52.4337
R17262 vdd.n2826 vdd.n2825 52.4337
R17263 vdd.n2819 vdd.n602 52.4337
R17264 vdd.n2818 vdd.n607 52.4337
R17265 vdd.n2814 vdd.n609 52.4337
R17266 vdd.n2034 vdd.n1614 52.4337
R17267 vdd.n2032 vdd.n2031 52.4337
R17268 vdd.n1621 vdd.n1620 52.4337
R17269 vdd.n1810 vdd.n1809 52.4337
R17270 vdd.n1807 vdd.n1806 52.4337
R17271 vdd.n1802 vdd.n1629 52.4337
R17272 vdd.n1800 vdd.n1799 52.4337
R17273 vdd.n1795 vdd.n1636 52.4337
R17274 vdd.n1793 vdd.n1792 52.4337
R17275 vdd.n1645 vdd.n1644 52.4337
R17276 vdd.n1784 vdd.n1649 52.4337
R17277 vdd.n1782 vdd.n1781 52.4337
R17278 vdd.n1777 vdd.n1655 52.4337
R17279 vdd.n1775 vdd.n1774 52.4337
R17280 vdd.n1770 vdd.n1662 52.4337
R17281 vdd.n1768 vdd.n1767 52.4337
R17282 vdd.n1763 vdd.n1669 52.4337
R17283 vdd.n1761 vdd.n1760 52.4337
R17284 vdd.n1756 vdd.n1676 52.4337
R17285 vdd.n1754 vdd.n1753 52.4337
R17286 vdd.n1685 vdd.n1684 52.4337
R17287 vdd.n1745 vdd.n1689 52.4337
R17288 vdd.n1743 vdd.n1742 52.4337
R17289 vdd.n1738 vdd.n1695 52.4337
R17290 vdd.n1736 vdd.n1735 52.4337
R17291 vdd.n1731 vdd.n1702 52.4337
R17292 vdd.n1729 vdd.n1728 52.4337
R17293 vdd.n1724 vdd.n1710 52.4337
R17294 vdd.n1722 vdd.n1721 52.4337
R17295 vdd.n1717 vdd.n1716 52.4337
R17296 vdd.n1712 vdd.n1711 52.4337
R17297 vdd.n2043 vdd.n898 52.4337
R17298 vdd.n986 vdd.n984 52.4337
R17299 vdd.n992 vdd.n991 52.4337
R17300 vdd.n995 vdd.n994 52.4337
R17301 vdd.n1000 vdd.n999 52.4337
R17302 vdd.n1003 vdd.n1002 52.4337
R17303 vdd.n1008 vdd.n1007 52.4337
R17304 vdd.n1011 vdd.n1010 52.4337
R17305 vdd.n1016 vdd.n1015 52.4337
R17306 vdd.n1019 vdd.n1018 52.4337
R17307 vdd.n1026 vdd.n1025 52.4337
R17308 vdd.n1029 vdd.n1028 52.4337
R17309 vdd.n1034 vdd.n1033 52.4337
R17310 vdd.n1037 vdd.n1036 52.4337
R17311 vdd.n1042 vdd.n1041 52.4337
R17312 vdd.n1045 vdd.n1044 52.4337
R17313 vdd.n1050 vdd.n1049 52.4337
R17314 vdd.n1053 vdd.n1052 52.4337
R17315 vdd.n1058 vdd.n1057 52.4337
R17316 vdd.n1061 vdd.n1060 52.4337
R17317 vdd.n1066 vdd.n1065 52.4337
R17318 vdd.n1146 vdd.n1145 52.4337
R17319 vdd.n1143 vdd.n1069 52.4337
R17320 vdd.n1075 vdd.n1074 52.4337
R17321 vdd.n1080 vdd.n1077 52.4337
R17322 vdd.n1083 vdd.n1082 52.4337
R17323 vdd.n1088 vdd.n1085 52.4337
R17324 vdd.n1091 vdd.n1090 52.4337
R17325 vdd.n1096 vdd.n1093 52.4337
R17326 vdd.n1099 vdd.n1098 52.4337
R17327 vdd.n1104 vdd.n1101 52.4337
R17328 vdd.n1107 vdd.n1106 52.4337
R17329 vdd.n987 vdd.n986 52.4337
R17330 vdd.n993 vdd.n992 52.4337
R17331 vdd.n996 vdd.n995 52.4337
R17332 vdd.n1001 vdd.n1000 52.4337
R17333 vdd.n1004 vdd.n1003 52.4337
R17334 vdd.n1009 vdd.n1008 52.4337
R17335 vdd.n1012 vdd.n1011 52.4337
R17336 vdd.n1017 vdd.n1016 52.4337
R17337 vdd.n1020 vdd.n1019 52.4337
R17338 vdd.n1027 vdd.n1026 52.4337
R17339 vdd.n1030 vdd.n1029 52.4337
R17340 vdd.n1035 vdd.n1034 52.4337
R17341 vdd.n1038 vdd.n1037 52.4337
R17342 vdd.n1043 vdd.n1042 52.4337
R17343 vdd.n1046 vdd.n1045 52.4337
R17344 vdd.n1051 vdd.n1050 52.4337
R17345 vdd.n1054 vdd.n1053 52.4337
R17346 vdd.n1059 vdd.n1058 52.4337
R17347 vdd.n1062 vdd.n1061 52.4337
R17348 vdd.n1067 vdd.n1066 52.4337
R17349 vdd.n1145 vdd.n1144 52.4337
R17350 vdd.n1073 vdd.n1069 52.4337
R17351 vdd.n1076 vdd.n1075 52.4337
R17352 vdd.n1081 vdd.n1080 52.4337
R17353 vdd.n1084 vdd.n1083 52.4337
R17354 vdd.n1089 vdd.n1088 52.4337
R17355 vdd.n1092 vdd.n1091 52.4337
R17356 vdd.n1097 vdd.n1096 52.4337
R17357 vdd.n1100 vdd.n1099 52.4337
R17358 vdd.n1105 vdd.n1104 52.4337
R17359 vdd.n1108 vdd.n1107 52.4337
R17360 vdd.n898 vdd.n897 52.4337
R17361 vdd.n1713 vdd.n1712 52.4337
R17362 vdd.n1718 vdd.n1717 52.4337
R17363 vdd.n1723 vdd.n1722 52.4337
R17364 vdd.n1710 vdd.n1703 52.4337
R17365 vdd.n1730 vdd.n1729 52.4337
R17366 vdd.n1702 vdd.n1696 52.4337
R17367 vdd.n1737 vdd.n1736 52.4337
R17368 vdd.n1695 vdd.n1690 52.4337
R17369 vdd.n1744 vdd.n1743 52.4337
R17370 vdd.n1689 vdd.n1688 52.4337
R17371 vdd.n1684 vdd.n1677 52.4337
R17372 vdd.n1755 vdd.n1754 52.4337
R17373 vdd.n1676 vdd.n1670 52.4337
R17374 vdd.n1762 vdd.n1761 52.4337
R17375 vdd.n1669 vdd.n1663 52.4337
R17376 vdd.n1769 vdd.n1768 52.4337
R17377 vdd.n1662 vdd.n1656 52.4337
R17378 vdd.n1776 vdd.n1775 52.4337
R17379 vdd.n1655 vdd.n1650 52.4337
R17380 vdd.n1783 vdd.n1782 52.4337
R17381 vdd.n1649 vdd.n1648 52.4337
R17382 vdd.n1644 vdd.n1637 52.4337
R17383 vdd.n1794 vdd.n1793 52.4337
R17384 vdd.n1636 vdd.n1630 52.4337
R17385 vdd.n1801 vdd.n1800 52.4337
R17386 vdd.n1629 vdd.n1623 52.4337
R17387 vdd.n1808 vdd.n1807 52.4337
R17388 vdd.n1811 vdd.n1810 52.4337
R17389 vdd.n1620 vdd.n1615 52.4337
R17390 vdd.n2033 vdd.n2032 52.4337
R17391 vdd.n1614 vdd.n903 52.4337
R17392 vdd.n2933 vdd.n2932 52.4337
R17393 vdd.n2927 vdd.n520 52.4337
R17394 vdd.n2923 vdd.n523 52.4337
R17395 vdd.n2921 vdd.n2920 52.4337
R17396 vdd.n2916 vdd.n2915 52.4337
R17397 vdd.n2913 vdd.n2912 52.4337
R17398 vdd.n2908 vdd.n2907 52.4337
R17399 vdd.n2905 vdd.n2904 52.4337
R17400 vdd.n2900 vdd.n2899 52.4337
R17401 vdd.n2897 vdd.n2896 52.4337
R17402 vdd.n2892 vdd.n2891 52.4337
R17403 vdd.n2889 vdd.n2888 52.4337
R17404 vdd.n2884 vdd.n2883 52.4337
R17405 vdd.n2881 vdd.n2880 52.4337
R17406 vdd.n2876 vdd.n2875 52.4337
R17407 vdd.n2873 vdd.n2872 52.4337
R17408 vdd.n2868 vdd.n2867 52.4337
R17409 vdd.n2865 vdd.n2864 52.4337
R17410 vdd.n2860 vdd.n2859 52.4337
R17411 vdd.n2857 vdd.n2856 52.4337
R17412 vdd.n585 vdd.n584 52.4337
R17413 vdd.n2848 vdd.n2847 52.4337
R17414 vdd.n2843 vdd.n586 52.4337
R17415 vdd.n2841 vdd.n2840 52.4337
R17416 vdd.n2836 vdd.n2835 52.4337
R17417 vdd.n2833 vdd.n2832 52.4337
R17418 vdd.n2828 vdd.n2827 52.4337
R17419 vdd.n2825 vdd.n2824 52.4337
R17420 vdd.n2820 vdd.n2819 52.4337
R17421 vdd.n2815 vdd.n607 52.4337
R17422 vdd.n2811 vdd.n609 52.4337
R17423 vdd.n3018 vdd.n462 52.4337
R17424 vdd.n3028 vdd.n3027 52.4337
R17425 vdd.n461 vdd.n455 52.4337
R17426 vdd.n3035 vdd.n3034 52.4337
R17427 vdd.n454 vdd.n448 52.4337
R17428 vdd.n3042 vdd.n3041 52.4337
R17429 vdd.n447 vdd.n441 52.4337
R17430 vdd.n3049 vdd.n3048 52.4337
R17431 vdd.n440 vdd.n435 52.4337
R17432 vdd.n3056 vdd.n3055 52.4337
R17433 vdd.n434 vdd.n433 52.4337
R17434 vdd.n429 vdd.n422 52.4337
R17435 vdd.n3067 vdd.n3066 52.4337
R17436 vdd.n421 vdd.n415 52.4337
R17437 vdd.n3074 vdd.n3073 52.4337
R17438 vdd.n414 vdd.n408 52.4337
R17439 vdd.n3081 vdd.n3080 52.4337
R17440 vdd.n407 vdd.n401 52.4337
R17441 vdd.n3088 vdd.n3087 52.4337
R17442 vdd.n400 vdd.n395 52.4337
R17443 vdd.n3095 vdd.n3094 52.4337
R17444 vdd.n394 vdd.n393 52.4337
R17445 vdd.n389 vdd.n382 52.4337
R17446 vdd.n3106 vdd.n3105 52.4337
R17447 vdd.n381 vdd.n375 52.4337
R17448 vdd.n3113 vdd.n3112 52.4337
R17449 vdd.n374 vdd.n368 52.4337
R17450 vdd.n3120 vdd.n3119 52.4337
R17451 vdd.n367 vdd.n360 52.4337
R17452 vdd.n3127 vdd.n3126 52.4337
R17453 vdd.n3130 vdd.n3129 52.4337
R17454 vdd.n355 vdd.n352 52.4337
R17455 vdd.t156 vdd.t204 51.4683
R17456 vdd.n258 vdd.n256 42.0461
R17457 vdd.n164 vdd.n162 42.0461
R17458 vdd.n71 vdd.n69 42.0461
R17459 vdd.n1504 vdd.n1502 42.0461
R17460 vdd.n1410 vdd.n1408 42.0461
R17461 vdd.n1317 vdd.n1315 42.0461
R17462 vdd.n308 vdd.n307 41.6884
R17463 vdd.n214 vdd.n213 41.6884
R17464 vdd.n121 vdd.n120 41.6884
R17465 vdd.n1554 vdd.n1553 41.6884
R17466 vdd.n1460 vdd.n1459 41.6884
R17467 vdd.n1367 vdd.n1366 41.6884
R17468 vdd.n1112 vdd.n1111 41.1157
R17469 vdd.n1149 vdd.n1148 41.1157
R17470 vdd.n1023 vdd.n1022 41.1157
R17471 vdd.n3023 vdd.n3022 41.1157
R17472 vdd.n3062 vdd.n428 41.1157
R17473 vdd.n3101 vdd.n388 41.1157
R17474 vdd.n2765 vdd.n2764 39.2114
R17475 vdd.n2762 vdd.n2761 39.2114
R17476 vdd.n2757 vdd.n641 39.2114
R17477 vdd.n2755 vdd.n2754 39.2114
R17478 vdd.n2750 vdd.n644 39.2114
R17479 vdd.n2748 vdd.n2747 39.2114
R17480 vdd.n2743 vdd.n647 39.2114
R17481 vdd.n2741 vdd.n2740 39.2114
R17482 vdd.n2735 vdd.n650 39.2114
R17483 vdd.n2733 vdd.n2732 39.2114
R17484 vdd.n2728 vdd.n653 39.2114
R17485 vdd.n2726 vdd.n2725 39.2114
R17486 vdd.n2721 vdd.n656 39.2114
R17487 vdd.n2719 vdd.n2718 39.2114
R17488 vdd.n2714 vdd.n659 39.2114
R17489 vdd.n2712 vdd.n2711 39.2114
R17490 vdd.n2707 vdd.n2706 39.2114
R17491 vdd.n2568 vdd.n741 39.2114
R17492 vdd.n2563 vdd.n2317 39.2114
R17493 vdd.n2560 vdd.n2318 39.2114
R17494 vdd.n2556 vdd.n2319 39.2114
R17495 vdd.n2552 vdd.n2320 39.2114
R17496 vdd.n2548 vdd.n2321 39.2114
R17497 vdd.n2544 vdd.n2322 39.2114
R17498 vdd.n2540 vdd.n2323 39.2114
R17499 vdd.n2536 vdd.n2324 39.2114
R17500 vdd.n2532 vdd.n2325 39.2114
R17501 vdd.n2528 vdd.n2326 39.2114
R17502 vdd.n2524 vdd.n2327 39.2114
R17503 vdd.n2520 vdd.n2328 39.2114
R17504 vdd.n2516 vdd.n2329 39.2114
R17505 vdd.n2512 vdd.n2330 39.2114
R17506 vdd.n2508 vdd.n2331 39.2114
R17507 vdd.n2503 vdd.n2332 39.2114
R17508 vdd.n2311 vdd.n781 39.2114
R17509 vdd.n2307 vdd.n780 39.2114
R17510 vdd.n2303 vdd.n779 39.2114
R17511 vdd.n2299 vdd.n778 39.2114
R17512 vdd.n2295 vdd.n777 39.2114
R17513 vdd.n2291 vdd.n776 39.2114
R17514 vdd.n2287 vdd.n775 39.2114
R17515 vdd.n2283 vdd.n774 39.2114
R17516 vdd.n2279 vdd.n773 39.2114
R17517 vdd.n2275 vdd.n772 39.2114
R17518 vdd.n2271 vdd.n771 39.2114
R17519 vdd.n2267 vdd.n770 39.2114
R17520 vdd.n2263 vdd.n769 39.2114
R17521 vdd.n2259 vdd.n768 39.2114
R17522 vdd.n2255 vdd.n767 39.2114
R17523 vdd.n2250 vdd.n766 39.2114
R17524 vdd.n2246 vdd.n765 39.2114
R17525 vdd.n1822 vdd.n876 39.2114
R17526 vdd.n1828 vdd.n1827 39.2114
R17527 vdd.n1831 vdd.n1830 39.2114
R17528 vdd.n1836 vdd.n1835 39.2114
R17529 vdd.n1839 vdd.n1838 39.2114
R17530 vdd.n1844 vdd.n1843 39.2114
R17531 vdd.n1847 vdd.n1846 39.2114
R17532 vdd.n1852 vdd.n1851 39.2114
R17533 vdd.n2023 vdd.n1854 39.2114
R17534 vdd.n2022 vdd.n2021 39.2114
R17535 vdd.n2015 vdd.n1856 39.2114
R17536 vdd.n2014 vdd.n2013 39.2114
R17537 vdd.n2007 vdd.n1858 39.2114
R17538 vdd.n2006 vdd.n2005 39.2114
R17539 vdd.n1999 vdd.n1860 39.2114
R17540 vdd.n1998 vdd.n1997 39.2114
R17541 vdd.n1991 vdd.n1862 39.2114
R17542 vdd.n2684 vdd.n2683 39.2114
R17543 vdd.n2679 vdd.n2651 39.2114
R17544 vdd.n2677 vdd.n2676 39.2114
R17545 vdd.n2672 vdd.n2654 39.2114
R17546 vdd.n2670 vdd.n2669 39.2114
R17547 vdd.n2665 vdd.n2657 39.2114
R17548 vdd.n2663 vdd.n2662 39.2114
R17549 vdd.n2658 vdd.n612 39.2114
R17550 vdd.n2802 vdd.n2801 39.2114
R17551 vdd.n2799 vdd.n2798 39.2114
R17552 vdd.n2794 vdd.n617 39.2114
R17553 vdd.n2792 vdd.n2791 39.2114
R17554 vdd.n2787 vdd.n620 39.2114
R17555 vdd.n2785 vdd.n2784 39.2114
R17556 vdd.n2780 vdd.n623 39.2114
R17557 vdd.n2778 vdd.n2777 39.2114
R17558 vdd.n2773 vdd.n629 39.2114
R17559 vdd.n2570 vdd.n744 39.2114
R17560 vdd.n2333 vdd.n746 39.2114
R17561 vdd.n2359 vdd.n2334 39.2114
R17562 vdd.n2363 vdd.n2335 39.2114
R17563 vdd.n2367 vdd.n2336 39.2114
R17564 vdd.n2371 vdd.n2337 39.2114
R17565 vdd.n2375 vdd.n2338 39.2114
R17566 vdd.n2379 vdd.n2339 39.2114
R17567 vdd.n2383 vdd.n2340 39.2114
R17568 vdd.n2387 vdd.n2341 39.2114
R17569 vdd.n2391 vdd.n2342 39.2114
R17570 vdd.n2395 vdd.n2343 39.2114
R17571 vdd.n2399 vdd.n2344 39.2114
R17572 vdd.n2403 vdd.n2345 39.2114
R17573 vdd.n2407 vdd.n2346 39.2114
R17574 vdd.n2411 vdd.n2347 39.2114
R17575 vdd.n2415 vdd.n2348 39.2114
R17576 vdd.n2571 vdd.n2570 39.2114
R17577 vdd.n2358 vdd.n2333 39.2114
R17578 vdd.n2362 vdd.n2334 39.2114
R17579 vdd.n2366 vdd.n2335 39.2114
R17580 vdd.n2370 vdd.n2336 39.2114
R17581 vdd.n2374 vdd.n2337 39.2114
R17582 vdd.n2378 vdd.n2338 39.2114
R17583 vdd.n2382 vdd.n2339 39.2114
R17584 vdd.n2386 vdd.n2340 39.2114
R17585 vdd.n2390 vdd.n2341 39.2114
R17586 vdd.n2394 vdd.n2342 39.2114
R17587 vdd.n2398 vdd.n2343 39.2114
R17588 vdd.n2402 vdd.n2344 39.2114
R17589 vdd.n2406 vdd.n2345 39.2114
R17590 vdd.n2410 vdd.n2346 39.2114
R17591 vdd.n2414 vdd.n2347 39.2114
R17592 vdd.n2417 vdd.n2348 39.2114
R17593 vdd.n629 vdd.n624 39.2114
R17594 vdd.n2779 vdd.n2778 39.2114
R17595 vdd.n623 vdd.n621 39.2114
R17596 vdd.n2786 vdd.n2785 39.2114
R17597 vdd.n620 vdd.n618 39.2114
R17598 vdd.n2793 vdd.n2792 39.2114
R17599 vdd.n617 vdd.n615 39.2114
R17600 vdd.n2800 vdd.n2799 39.2114
R17601 vdd.n2803 vdd.n2802 39.2114
R17602 vdd.n2659 vdd.n2658 39.2114
R17603 vdd.n2664 vdd.n2663 39.2114
R17604 vdd.n2657 vdd.n2655 39.2114
R17605 vdd.n2671 vdd.n2670 39.2114
R17606 vdd.n2654 vdd.n2652 39.2114
R17607 vdd.n2678 vdd.n2677 39.2114
R17608 vdd.n2651 vdd.n2649 39.2114
R17609 vdd.n2685 vdd.n2684 39.2114
R17610 vdd.n1823 vdd.n1822 39.2114
R17611 vdd.n1829 vdd.n1828 39.2114
R17612 vdd.n1830 vdd.n1819 39.2114
R17613 vdd.n1837 vdd.n1836 39.2114
R17614 vdd.n1838 vdd.n1817 39.2114
R17615 vdd.n1845 vdd.n1844 39.2114
R17616 vdd.n1846 vdd.n1815 39.2114
R17617 vdd.n1853 vdd.n1852 39.2114
R17618 vdd.n2024 vdd.n2023 39.2114
R17619 vdd.n2021 vdd.n2020 39.2114
R17620 vdd.n2016 vdd.n2015 39.2114
R17621 vdd.n2013 vdd.n2012 39.2114
R17622 vdd.n2008 vdd.n2007 39.2114
R17623 vdd.n2005 vdd.n2004 39.2114
R17624 vdd.n2000 vdd.n1999 39.2114
R17625 vdd.n1997 vdd.n1996 39.2114
R17626 vdd.n1992 vdd.n1991 39.2114
R17627 vdd.n2249 vdd.n765 39.2114
R17628 vdd.n2254 vdd.n766 39.2114
R17629 vdd.n2258 vdd.n767 39.2114
R17630 vdd.n2262 vdd.n768 39.2114
R17631 vdd.n2266 vdd.n769 39.2114
R17632 vdd.n2270 vdd.n770 39.2114
R17633 vdd.n2274 vdd.n771 39.2114
R17634 vdd.n2278 vdd.n772 39.2114
R17635 vdd.n2282 vdd.n773 39.2114
R17636 vdd.n2286 vdd.n774 39.2114
R17637 vdd.n2290 vdd.n775 39.2114
R17638 vdd.n2294 vdd.n776 39.2114
R17639 vdd.n2298 vdd.n777 39.2114
R17640 vdd.n2302 vdd.n778 39.2114
R17641 vdd.n2306 vdd.n779 39.2114
R17642 vdd.n2310 vdd.n780 39.2114
R17643 vdd.n783 vdd.n781 39.2114
R17644 vdd.n2568 vdd.n2567 39.2114
R17645 vdd.n2561 vdd.n2317 39.2114
R17646 vdd.n2557 vdd.n2318 39.2114
R17647 vdd.n2553 vdd.n2319 39.2114
R17648 vdd.n2549 vdd.n2320 39.2114
R17649 vdd.n2545 vdd.n2321 39.2114
R17650 vdd.n2541 vdd.n2322 39.2114
R17651 vdd.n2537 vdd.n2323 39.2114
R17652 vdd.n2533 vdd.n2324 39.2114
R17653 vdd.n2529 vdd.n2325 39.2114
R17654 vdd.n2525 vdd.n2326 39.2114
R17655 vdd.n2521 vdd.n2327 39.2114
R17656 vdd.n2517 vdd.n2328 39.2114
R17657 vdd.n2513 vdd.n2329 39.2114
R17658 vdd.n2509 vdd.n2330 39.2114
R17659 vdd.n2504 vdd.n2331 39.2114
R17660 vdd.n2500 vdd.n2332 39.2114
R17661 vdd.n2706 vdd.n660 39.2114
R17662 vdd.n2713 vdd.n2712 39.2114
R17663 vdd.n659 vdd.n657 39.2114
R17664 vdd.n2720 vdd.n2719 39.2114
R17665 vdd.n656 vdd.n654 39.2114
R17666 vdd.n2727 vdd.n2726 39.2114
R17667 vdd.n653 vdd.n651 39.2114
R17668 vdd.n2734 vdd.n2733 39.2114
R17669 vdd.n650 vdd.n648 39.2114
R17670 vdd.n2742 vdd.n2741 39.2114
R17671 vdd.n647 vdd.n645 39.2114
R17672 vdd.n2749 vdd.n2748 39.2114
R17673 vdd.n644 vdd.n642 39.2114
R17674 vdd.n2756 vdd.n2755 39.2114
R17675 vdd.n641 vdd.n639 39.2114
R17676 vdd.n2763 vdd.n2762 39.2114
R17677 vdd.n2766 vdd.n2765 39.2114
R17678 vdd.n791 vdd.n747 39.2114
R17679 vdd.n2238 vdd.n748 39.2114
R17680 vdd.n2234 vdd.n749 39.2114
R17681 vdd.n2230 vdd.n750 39.2114
R17682 vdd.n2226 vdd.n751 39.2114
R17683 vdd.n2222 vdd.n752 39.2114
R17684 vdd.n2218 vdd.n753 39.2114
R17685 vdd.n2214 vdd.n754 39.2114
R17686 vdd.n2210 vdd.n755 39.2114
R17687 vdd.n2206 vdd.n756 39.2114
R17688 vdd.n2202 vdd.n757 39.2114
R17689 vdd.n2198 vdd.n758 39.2114
R17690 vdd.n2194 vdd.n759 39.2114
R17691 vdd.n2190 vdd.n760 39.2114
R17692 vdd.n2186 vdd.n761 39.2114
R17693 vdd.n2182 vdd.n762 39.2114
R17694 vdd.n2178 vdd.n763 39.2114
R17695 vdd.n2081 vdd.n880 39.2114
R17696 vdd.n2080 vdd.n2079 39.2114
R17697 vdd.n2073 vdd.n882 39.2114
R17698 vdd.n2072 vdd.n2071 39.2114
R17699 vdd.n2065 vdd.n884 39.2114
R17700 vdd.n2064 vdd.n2063 39.2114
R17701 vdd.n2057 vdd.n886 39.2114
R17702 vdd.n2056 vdd.n2055 39.2114
R17703 vdd.n889 vdd.n888 39.2114
R17704 vdd.n1897 vdd.n1896 39.2114
R17705 vdd.n1902 vdd.n1901 39.2114
R17706 vdd.n1905 vdd.n1904 39.2114
R17707 vdd.n1910 vdd.n1909 39.2114
R17708 vdd.n1913 vdd.n1912 39.2114
R17709 vdd.n1918 vdd.n1917 39.2114
R17710 vdd.n1921 vdd.n1920 39.2114
R17711 vdd.n1927 vdd.n1926 39.2114
R17712 vdd.n2175 vdd.n763 39.2114
R17713 vdd.n2179 vdd.n762 39.2114
R17714 vdd.n2183 vdd.n761 39.2114
R17715 vdd.n2187 vdd.n760 39.2114
R17716 vdd.n2191 vdd.n759 39.2114
R17717 vdd.n2195 vdd.n758 39.2114
R17718 vdd.n2199 vdd.n757 39.2114
R17719 vdd.n2203 vdd.n756 39.2114
R17720 vdd.n2207 vdd.n755 39.2114
R17721 vdd.n2211 vdd.n754 39.2114
R17722 vdd.n2215 vdd.n753 39.2114
R17723 vdd.n2219 vdd.n752 39.2114
R17724 vdd.n2223 vdd.n751 39.2114
R17725 vdd.n2227 vdd.n750 39.2114
R17726 vdd.n2231 vdd.n749 39.2114
R17727 vdd.n2235 vdd.n748 39.2114
R17728 vdd.n2239 vdd.n747 39.2114
R17729 vdd.n2082 vdd.n2081 39.2114
R17730 vdd.n2079 vdd.n2078 39.2114
R17731 vdd.n2074 vdd.n2073 39.2114
R17732 vdd.n2071 vdd.n2070 39.2114
R17733 vdd.n2066 vdd.n2065 39.2114
R17734 vdd.n2063 vdd.n2062 39.2114
R17735 vdd.n2058 vdd.n2057 39.2114
R17736 vdd.n2055 vdd.n2054 39.2114
R17737 vdd.n890 vdd.n889 39.2114
R17738 vdd.n1898 vdd.n1897 39.2114
R17739 vdd.n1903 vdd.n1902 39.2114
R17740 vdd.n1904 vdd.n1894 39.2114
R17741 vdd.n1911 vdd.n1910 39.2114
R17742 vdd.n1912 vdd.n1892 39.2114
R17743 vdd.n1919 vdd.n1918 39.2114
R17744 vdd.n1920 vdd.n1888 39.2114
R17745 vdd.n1928 vdd.n1927 39.2114
R17746 vdd.n2047 vdd.n2046 37.2369
R17747 vdd.n1750 vdd.n1683 37.2369
R17748 vdd.n1789 vdd.n1643 37.2369
R17749 vdd.n2854 vdd.n581 37.2369
R17750 vdd.n545 vdd.n544 37.2369
R17751 vdd.n2810 vdd.n2809 37.2369
R17752 vdd.n2089 vdd.n875 31.6883
R17753 vdd.n2314 vdd.n784 31.6883
R17754 vdd.n2247 vdd.n787 31.6883
R17755 vdd.n1993 vdd.n1990 31.6883
R17756 vdd.n2501 vdd.n2499 31.6883
R17757 vdd.n2708 vdd.n2705 31.6883
R17758 vdd.n2578 vdd.n740 31.6883
R17759 vdd.n2769 vdd.n2768 31.6883
R17760 vdd.n2688 vdd.n2687 31.6883
R17761 vdd.n2774 vdd.n628 31.6883
R17762 vdd.n2420 vdd.n2419 31.6883
R17763 vdd.n2574 vdd.n2573 31.6883
R17764 vdd.n2085 vdd.n2084 31.6883
R17765 vdd.n2242 vdd.n2241 31.6883
R17766 vdd.n2174 vdd.n2173 31.6883
R17767 vdd.n1931 vdd.n1930 31.6883
R17768 vdd.n1924 vdd.n1890 30.449
R17769 vdd.n795 vdd.n794 30.449
R17770 vdd.n1865 vdd.n1864 30.449
R17771 vdd.n2252 vdd.n786 30.449
R17772 vdd.n2356 vdd.n2355 30.449
R17773 vdd.n663 vdd.n662 30.449
R17774 vdd.n2506 vdd.n2352 30.449
R17775 vdd.n627 vdd.n626 30.449
R17776 vdd.n1215 vdd.n982 20.633
R17777 vdd.n2041 vdd.n901 20.633
R17778 vdd.n2940 vdd.n516 20.633
R17779 vdd.n3138 vdd.n351 20.633
R17780 vdd.n1217 vdd.n979 19.3944
R17781 vdd.n1221 vdd.n979 19.3944
R17782 vdd.n1221 vdd.n970 19.3944
R17783 vdd.n1233 vdd.n970 19.3944
R17784 vdd.n1233 vdd.n968 19.3944
R17785 vdd.n1237 vdd.n968 19.3944
R17786 vdd.n1237 vdd.n957 19.3944
R17787 vdd.n1249 vdd.n957 19.3944
R17788 vdd.n1249 vdd.n955 19.3944
R17789 vdd.n1253 vdd.n955 19.3944
R17790 vdd.n1253 vdd.n946 19.3944
R17791 vdd.n1266 vdd.n946 19.3944
R17792 vdd.n1266 vdd.n944 19.3944
R17793 vdd.n1270 vdd.n944 19.3944
R17794 vdd.n1270 vdd.n935 19.3944
R17795 vdd.n1564 vdd.n935 19.3944
R17796 vdd.n1564 vdd.n933 19.3944
R17797 vdd.n1568 vdd.n933 19.3944
R17798 vdd.n1568 vdd.n923 19.3944
R17799 vdd.n1581 vdd.n923 19.3944
R17800 vdd.n1581 vdd.n921 19.3944
R17801 vdd.n1585 vdd.n921 19.3944
R17802 vdd.n1585 vdd.n913 19.3944
R17803 vdd.n1598 vdd.n913 19.3944
R17804 vdd.n1598 vdd.n910 19.3944
R17805 vdd.n1604 vdd.n910 19.3944
R17806 vdd.n1604 vdd.n911 19.3944
R17807 vdd.n911 vdd.n900 19.3944
R17808 vdd.n1142 vdd.n1068 19.3944
R17809 vdd.n1142 vdd.n1070 19.3944
R17810 vdd.n1138 vdd.n1070 19.3944
R17811 vdd.n1138 vdd.n1137 19.3944
R17812 vdd.n1137 vdd.n1136 19.3944
R17813 vdd.n1136 vdd.n1078 19.3944
R17814 vdd.n1132 vdd.n1078 19.3944
R17815 vdd.n1132 vdd.n1131 19.3944
R17816 vdd.n1131 vdd.n1130 19.3944
R17817 vdd.n1130 vdd.n1086 19.3944
R17818 vdd.n1126 vdd.n1086 19.3944
R17819 vdd.n1126 vdd.n1125 19.3944
R17820 vdd.n1125 vdd.n1124 19.3944
R17821 vdd.n1124 vdd.n1094 19.3944
R17822 vdd.n1120 vdd.n1094 19.3944
R17823 vdd.n1120 vdd.n1119 19.3944
R17824 vdd.n1119 vdd.n1118 19.3944
R17825 vdd.n1118 vdd.n1102 19.3944
R17826 vdd.n1114 vdd.n1102 19.3944
R17827 vdd.n1114 vdd.n1113 19.3944
R17828 vdd.n1180 vdd.n1179 19.3944
R17829 vdd.n1179 vdd.n1178 19.3944
R17830 vdd.n1178 vdd.n1031 19.3944
R17831 vdd.n1174 vdd.n1031 19.3944
R17832 vdd.n1174 vdd.n1173 19.3944
R17833 vdd.n1173 vdd.n1172 19.3944
R17834 vdd.n1172 vdd.n1039 19.3944
R17835 vdd.n1168 vdd.n1039 19.3944
R17836 vdd.n1168 vdd.n1167 19.3944
R17837 vdd.n1167 vdd.n1166 19.3944
R17838 vdd.n1166 vdd.n1047 19.3944
R17839 vdd.n1162 vdd.n1047 19.3944
R17840 vdd.n1162 vdd.n1161 19.3944
R17841 vdd.n1161 vdd.n1160 19.3944
R17842 vdd.n1160 vdd.n1055 19.3944
R17843 vdd.n1156 vdd.n1055 19.3944
R17844 vdd.n1156 vdd.n1155 19.3944
R17845 vdd.n1155 vdd.n1154 19.3944
R17846 vdd.n1154 vdd.n1063 19.3944
R17847 vdd.n1150 vdd.n1063 19.3944
R17848 vdd.n1210 vdd.n1209 19.3944
R17849 vdd.n1209 vdd.n1208 19.3944
R17850 vdd.n1208 vdd.n989 19.3944
R17851 vdd.n1204 vdd.n989 19.3944
R17852 vdd.n1204 vdd.n1203 19.3944
R17853 vdd.n1203 vdd.n1202 19.3944
R17854 vdd.n1202 vdd.n997 19.3944
R17855 vdd.n1198 vdd.n997 19.3944
R17856 vdd.n1198 vdd.n1197 19.3944
R17857 vdd.n1197 vdd.n1196 19.3944
R17858 vdd.n1196 vdd.n1005 19.3944
R17859 vdd.n1192 vdd.n1005 19.3944
R17860 vdd.n1192 vdd.n1191 19.3944
R17861 vdd.n1191 vdd.n1190 19.3944
R17862 vdd.n1190 vdd.n1013 19.3944
R17863 vdd.n1186 vdd.n1013 19.3944
R17864 vdd.n1186 vdd.n1185 19.3944
R17865 vdd.n1185 vdd.n1184 19.3944
R17866 vdd.n1746 vdd.n1681 19.3944
R17867 vdd.n1746 vdd.n1687 19.3944
R17868 vdd.n1741 vdd.n1687 19.3944
R17869 vdd.n1741 vdd.n1740 19.3944
R17870 vdd.n1740 vdd.n1739 19.3944
R17871 vdd.n1739 vdd.n1694 19.3944
R17872 vdd.n1734 vdd.n1694 19.3944
R17873 vdd.n1734 vdd.n1733 19.3944
R17874 vdd.n1733 vdd.n1732 19.3944
R17875 vdd.n1732 vdd.n1701 19.3944
R17876 vdd.n1727 vdd.n1701 19.3944
R17877 vdd.n1727 vdd.n1726 19.3944
R17878 vdd.n1726 vdd.n1725 19.3944
R17879 vdd.n1725 vdd.n1709 19.3944
R17880 vdd.n1720 vdd.n1709 19.3944
R17881 vdd.n1720 vdd.n1719 19.3944
R17882 vdd.n1715 vdd.n1714 19.3944
R17883 vdd.n2048 vdd.n896 19.3944
R17884 vdd.n1785 vdd.n1641 19.3944
R17885 vdd.n1785 vdd.n1647 19.3944
R17886 vdd.n1780 vdd.n1647 19.3944
R17887 vdd.n1780 vdd.n1779 19.3944
R17888 vdd.n1779 vdd.n1778 19.3944
R17889 vdd.n1778 vdd.n1654 19.3944
R17890 vdd.n1773 vdd.n1654 19.3944
R17891 vdd.n1773 vdd.n1772 19.3944
R17892 vdd.n1772 vdd.n1771 19.3944
R17893 vdd.n1771 vdd.n1661 19.3944
R17894 vdd.n1766 vdd.n1661 19.3944
R17895 vdd.n1766 vdd.n1765 19.3944
R17896 vdd.n1765 vdd.n1764 19.3944
R17897 vdd.n1764 vdd.n1668 19.3944
R17898 vdd.n1759 vdd.n1668 19.3944
R17899 vdd.n1759 vdd.n1758 19.3944
R17900 vdd.n1758 vdd.n1757 19.3944
R17901 vdd.n1757 vdd.n1675 19.3944
R17902 vdd.n1752 vdd.n1675 19.3944
R17903 vdd.n1752 vdd.n1751 19.3944
R17904 vdd.n2036 vdd.n2035 19.3944
R17905 vdd.n2035 vdd.n1613 19.3944
R17906 vdd.n2030 vdd.n2029 19.3944
R17907 vdd.n1812 vdd.n1617 19.3944
R17908 vdd.n1812 vdd.n1619 19.3944
R17909 vdd.n1622 vdd.n1619 19.3944
R17910 vdd.n1805 vdd.n1622 19.3944
R17911 vdd.n1805 vdd.n1804 19.3944
R17912 vdd.n1804 vdd.n1803 19.3944
R17913 vdd.n1803 vdd.n1628 19.3944
R17914 vdd.n1798 vdd.n1628 19.3944
R17915 vdd.n1798 vdd.n1797 19.3944
R17916 vdd.n1797 vdd.n1796 19.3944
R17917 vdd.n1796 vdd.n1635 19.3944
R17918 vdd.n1791 vdd.n1635 19.3944
R17919 vdd.n1791 vdd.n1790 19.3944
R17920 vdd.n1213 vdd.n976 19.3944
R17921 vdd.n1225 vdd.n976 19.3944
R17922 vdd.n1225 vdd.n974 19.3944
R17923 vdd.n1229 vdd.n974 19.3944
R17924 vdd.n1229 vdd.n964 19.3944
R17925 vdd.n1241 vdd.n964 19.3944
R17926 vdd.n1241 vdd.n962 19.3944
R17927 vdd.n1245 vdd.n962 19.3944
R17928 vdd.n1245 vdd.n952 19.3944
R17929 vdd.n1258 vdd.n952 19.3944
R17930 vdd.n1258 vdd.n950 19.3944
R17931 vdd.n1262 vdd.n950 19.3944
R17932 vdd.n1262 vdd.n941 19.3944
R17933 vdd.n1274 vdd.n941 19.3944
R17934 vdd.n1274 vdd.n939 19.3944
R17935 vdd.n1560 vdd.n939 19.3944
R17936 vdd.n1560 vdd.n929 19.3944
R17937 vdd.n1573 vdd.n929 19.3944
R17938 vdd.n1573 vdd.n927 19.3944
R17939 vdd.n1577 vdd.n927 19.3944
R17940 vdd.n1577 vdd.n918 19.3944
R17941 vdd.n1590 vdd.n918 19.3944
R17942 vdd.n1590 vdd.n916 19.3944
R17943 vdd.n1594 vdd.n916 19.3944
R17944 vdd.n1594 vdd.n906 19.3944
R17945 vdd.n1609 vdd.n906 19.3944
R17946 vdd.n1609 vdd.n904 19.3944
R17947 vdd.n2039 vdd.n904 19.3944
R17948 vdd.n2942 vdd.n513 19.3944
R17949 vdd.n2946 vdd.n513 19.3944
R17950 vdd.n2946 vdd.n503 19.3944
R17951 vdd.n2958 vdd.n503 19.3944
R17952 vdd.n2958 vdd.n501 19.3944
R17953 vdd.n2962 vdd.n501 19.3944
R17954 vdd.n2962 vdd.n490 19.3944
R17955 vdd.n2974 vdd.n490 19.3944
R17956 vdd.n2974 vdd.n488 19.3944
R17957 vdd.n2978 vdd.n488 19.3944
R17958 vdd.n2978 vdd.n478 19.3944
R17959 vdd.n2991 vdd.n478 19.3944
R17960 vdd.n2991 vdd.n476 19.3944
R17961 vdd.n2995 vdd.n476 19.3944
R17962 vdd.n2996 vdd.n2995 19.3944
R17963 vdd.n2997 vdd.n2996 19.3944
R17964 vdd.n2997 vdd.n474 19.3944
R17965 vdd.n3001 vdd.n474 19.3944
R17966 vdd.n3002 vdd.n3001 19.3944
R17967 vdd.n3003 vdd.n3002 19.3944
R17968 vdd.n3003 vdd.n471 19.3944
R17969 vdd.n3007 vdd.n471 19.3944
R17970 vdd.n3008 vdd.n3007 19.3944
R17971 vdd.n3009 vdd.n3008 19.3944
R17972 vdd.n3009 vdd.n468 19.3944
R17973 vdd.n3013 vdd.n468 19.3944
R17974 vdd.n3014 vdd.n3013 19.3944
R17975 vdd.n3015 vdd.n3014 19.3944
R17976 vdd.n3058 vdd.n426 19.3944
R17977 vdd.n3058 vdd.n432 19.3944
R17978 vdd.n3053 vdd.n432 19.3944
R17979 vdd.n3053 vdd.n3052 19.3944
R17980 vdd.n3052 vdd.n3051 19.3944
R17981 vdd.n3051 vdd.n439 19.3944
R17982 vdd.n3046 vdd.n439 19.3944
R17983 vdd.n3046 vdd.n3045 19.3944
R17984 vdd.n3045 vdd.n3044 19.3944
R17985 vdd.n3044 vdd.n446 19.3944
R17986 vdd.n3039 vdd.n446 19.3944
R17987 vdd.n3039 vdd.n3038 19.3944
R17988 vdd.n3038 vdd.n3037 19.3944
R17989 vdd.n3037 vdd.n453 19.3944
R17990 vdd.n3032 vdd.n453 19.3944
R17991 vdd.n3032 vdd.n3031 19.3944
R17992 vdd.n3031 vdd.n3030 19.3944
R17993 vdd.n3030 vdd.n460 19.3944
R17994 vdd.n3025 vdd.n460 19.3944
R17995 vdd.n3025 vdd.n3024 19.3944
R17996 vdd.n3097 vdd.n386 19.3944
R17997 vdd.n3097 vdd.n392 19.3944
R17998 vdd.n3092 vdd.n392 19.3944
R17999 vdd.n3092 vdd.n3091 19.3944
R18000 vdd.n3091 vdd.n3090 19.3944
R18001 vdd.n3090 vdd.n399 19.3944
R18002 vdd.n3085 vdd.n399 19.3944
R18003 vdd.n3085 vdd.n3084 19.3944
R18004 vdd.n3084 vdd.n3083 19.3944
R18005 vdd.n3083 vdd.n406 19.3944
R18006 vdd.n3078 vdd.n406 19.3944
R18007 vdd.n3078 vdd.n3077 19.3944
R18008 vdd.n3077 vdd.n3076 19.3944
R18009 vdd.n3076 vdd.n413 19.3944
R18010 vdd.n3071 vdd.n413 19.3944
R18011 vdd.n3071 vdd.n3070 19.3944
R18012 vdd.n3070 vdd.n3069 19.3944
R18013 vdd.n3069 vdd.n420 19.3944
R18014 vdd.n3064 vdd.n420 19.3944
R18015 vdd.n3064 vdd.n3063 19.3944
R18016 vdd.n3133 vdd.n3132 19.3944
R18017 vdd.n3132 vdd.n3131 19.3944
R18018 vdd.n3131 vdd.n358 19.3944
R18019 vdd.n359 vdd.n358 19.3944
R18020 vdd.n3124 vdd.n359 19.3944
R18021 vdd.n3124 vdd.n3123 19.3944
R18022 vdd.n3123 vdd.n3122 19.3944
R18023 vdd.n3122 vdd.n366 19.3944
R18024 vdd.n3117 vdd.n366 19.3944
R18025 vdd.n3117 vdd.n3116 19.3944
R18026 vdd.n3116 vdd.n3115 19.3944
R18027 vdd.n3115 vdd.n373 19.3944
R18028 vdd.n3110 vdd.n373 19.3944
R18029 vdd.n3110 vdd.n3109 19.3944
R18030 vdd.n3109 vdd.n3108 19.3944
R18031 vdd.n3108 vdd.n380 19.3944
R18032 vdd.n3103 vdd.n380 19.3944
R18033 vdd.n3103 vdd.n3102 19.3944
R18034 vdd.n2938 vdd.n509 19.3944
R18035 vdd.n2950 vdd.n509 19.3944
R18036 vdd.n2950 vdd.n507 19.3944
R18037 vdd.n2954 vdd.n507 19.3944
R18038 vdd.n2954 vdd.n497 19.3944
R18039 vdd.n2966 vdd.n497 19.3944
R18040 vdd.n2966 vdd.n495 19.3944
R18041 vdd.n2970 vdd.n495 19.3944
R18042 vdd.n2970 vdd.n485 19.3944
R18043 vdd.n2983 vdd.n485 19.3944
R18044 vdd.n2983 vdd.n483 19.3944
R18045 vdd.n2987 vdd.n483 19.3944
R18046 vdd.n2987 vdd.n312 19.3944
R18047 vdd.n3166 vdd.n312 19.3944
R18048 vdd.n3166 vdd.n313 19.3944
R18049 vdd.n3160 vdd.n313 19.3944
R18050 vdd.n3160 vdd.n3159 19.3944
R18051 vdd.n3159 vdd.n3158 19.3944
R18052 vdd.n3158 vdd.n323 19.3944
R18053 vdd.n3152 vdd.n323 19.3944
R18054 vdd.n3152 vdd.n3151 19.3944
R18055 vdd.n3151 vdd.n3150 19.3944
R18056 vdd.n3150 vdd.n335 19.3944
R18057 vdd.n3144 vdd.n335 19.3944
R18058 vdd.n3144 vdd.n3143 19.3944
R18059 vdd.n3143 vdd.n3142 19.3944
R18060 vdd.n3142 vdd.n346 19.3944
R18061 vdd.n3136 vdd.n346 19.3944
R18062 vdd.n2895 vdd.n2894 19.3944
R18063 vdd.n2894 vdd.n2893 19.3944
R18064 vdd.n2893 vdd.n551 19.3944
R18065 vdd.n2887 vdd.n551 19.3944
R18066 vdd.n2887 vdd.n2886 19.3944
R18067 vdd.n2886 vdd.n2885 19.3944
R18068 vdd.n2885 vdd.n557 19.3944
R18069 vdd.n2879 vdd.n557 19.3944
R18070 vdd.n2879 vdd.n2878 19.3944
R18071 vdd.n2878 vdd.n2877 19.3944
R18072 vdd.n2877 vdd.n563 19.3944
R18073 vdd.n2871 vdd.n563 19.3944
R18074 vdd.n2871 vdd.n2870 19.3944
R18075 vdd.n2870 vdd.n2869 19.3944
R18076 vdd.n2869 vdd.n569 19.3944
R18077 vdd.n2863 vdd.n569 19.3944
R18078 vdd.n2863 vdd.n2862 19.3944
R18079 vdd.n2862 vdd.n2861 19.3944
R18080 vdd.n2861 vdd.n575 19.3944
R18081 vdd.n2855 vdd.n575 19.3944
R18082 vdd.n2935 vdd.n2934 19.3944
R18083 vdd.n2934 vdd.n519 19.3944
R18084 vdd.n2929 vdd.n2928 19.3944
R18085 vdd.n2925 vdd.n2924 19.3944
R18086 vdd.n2924 vdd.n525 19.3944
R18087 vdd.n2919 vdd.n525 19.3944
R18088 vdd.n2919 vdd.n2918 19.3944
R18089 vdd.n2918 vdd.n2917 19.3944
R18090 vdd.n2917 vdd.n531 19.3944
R18091 vdd.n2911 vdd.n531 19.3944
R18092 vdd.n2911 vdd.n2910 19.3944
R18093 vdd.n2910 vdd.n2909 19.3944
R18094 vdd.n2909 vdd.n537 19.3944
R18095 vdd.n2903 vdd.n537 19.3944
R18096 vdd.n2903 vdd.n2902 19.3944
R18097 vdd.n2902 vdd.n2901 19.3944
R18098 vdd.n2850 vdd.n579 19.3944
R18099 vdd.n2850 vdd.n583 19.3944
R18100 vdd.n2845 vdd.n583 19.3944
R18101 vdd.n2845 vdd.n2844 19.3944
R18102 vdd.n2844 vdd.n589 19.3944
R18103 vdd.n2839 vdd.n589 19.3944
R18104 vdd.n2839 vdd.n2838 19.3944
R18105 vdd.n2838 vdd.n2837 19.3944
R18106 vdd.n2837 vdd.n595 19.3944
R18107 vdd.n2831 vdd.n595 19.3944
R18108 vdd.n2831 vdd.n2830 19.3944
R18109 vdd.n2830 vdd.n2829 19.3944
R18110 vdd.n2829 vdd.n601 19.3944
R18111 vdd.n2823 vdd.n601 19.3944
R18112 vdd.n2823 vdd.n2822 19.3944
R18113 vdd.n2822 vdd.n2821 19.3944
R18114 vdd.n2817 vdd.n2816 19.3944
R18115 vdd.n2813 vdd.n2812 19.3944
R18116 vdd.n1149 vdd.n1068 19.0066
R18117 vdd.n1750 vdd.n1681 19.0066
R18118 vdd.n3062 vdd.n426 19.0066
R18119 vdd.n2854 vdd.n579 19.0066
R18120 vdd.n1890 vdd.n1889 16.0975
R18121 vdd.n794 vdd.n793 16.0975
R18122 vdd.n1111 vdd.n1110 16.0975
R18123 vdd.n1148 vdd.n1147 16.0975
R18124 vdd.n1022 vdd.n1021 16.0975
R18125 vdd.n2046 vdd.n2045 16.0975
R18126 vdd.n1683 vdd.n1682 16.0975
R18127 vdd.n1643 vdd.n1642 16.0975
R18128 vdd.n1864 vdd.n1863 16.0975
R18129 vdd.n786 vdd.n785 16.0975
R18130 vdd.n2355 vdd.n2354 16.0975
R18131 vdd.n3022 vdd.n3021 16.0975
R18132 vdd.n428 vdd.n427 16.0975
R18133 vdd.n388 vdd.n387 16.0975
R18134 vdd.n581 vdd.n580 16.0975
R18135 vdd.n544 vdd.n543 16.0975
R18136 vdd.n662 vdd.n661 16.0975
R18137 vdd.n2352 vdd.n2351 16.0975
R18138 vdd.n2809 vdd.n2808 16.0975
R18139 vdd.n626 vdd.n625 16.0975
R18140 vdd.t204 vdd.n2316 15.4182
R18141 vdd.n2569 vdd.t156 15.4182
R18142 vdd.n28 vdd.n27 14.6905
R18143 vdd.n2087 vdd.n877 14.5112
R18144 vdd.n2771 vdd.n613 14.5112
R18145 vdd.n304 vdd.n269 13.1884
R18146 vdd.n253 vdd.n218 13.1884
R18147 vdd.n210 vdd.n175 13.1884
R18148 vdd.n159 vdd.n124 13.1884
R18149 vdd.n117 vdd.n82 13.1884
R18150 vdd.n66 vdd.n31 13.1884
R18151 vdd.n1499 vdd.n1464 13.1884
R18152 vdd.n1550 vdd.n1515 13.1884
R18153 vdd.n1405 vdd.n1370 13.1884
R18154 vdd.n1456 vdd.n1421 13.1884
R18155 vdd.n1312 vdd.n1277 13.1884
R18156 vdd.n1363 vdd.n1328 13.1884
R18157 vdd.n1180 vdd.n1023 12.9944
R18158 vdd.n1184 vdd.n1023 12.9944
R18159 vdd.n1789 vdd.n1641 12.9944
R18160 vdd.n1790 vdd.n1789 12.9944
R18161 vdd.n3101 vdd.n386 12.9944
R18162 vdd.n3102 vdd.n3101 12.9944
R18163 vdd.n2895 vdd.n545 12.9944
R18164 vdd.n2901 vdd.n545 12.9944
R18165 vdd.n305 vdd.n267 12.8005
R18166 vdd.n300 vdd.n271 12.8005
R18167 vdd.n254 vdd.n216 12.8005
R18168 vdd.n249 vdd.n220 12.8005
R18169 vdd.n211 vdd.n173 12.8005
R18170 vdd.n206 vdd.n177 12.8005
R18171 vdd.n160 vdd.n122 12.8005
R18172 vdd.n155 vdd.n126 12.8005
R18173 vdd.n118 vdd.n80 12.8005
R18174 vdd.n113 vdd.n84 12.8005
R18175 vdd.n67 vdd.n29 12.8005
R18176 vdd.n62 vdd.n33 12.8005
R18177 vdd.n1500 vdd.n1462 12.8005
R18178 vdd.n1495 vdd.n1466 12.8005
R18179 vdd.n1551 vdd.n1513 12.8005
R18180 vdd.n1546 vdd.n1517 12.8005
R18181 vdd.n1406 vdd.n1368 12.8005
R18182 vdd.n1401 vdd.n1372 12.8005
R18183 vdd.n1457 vdd.n1419 12.8005
R18184 vdd.n1452 vdd.n1423 12.8005
R18185 vdd.n1313 vdd.n1275 12.8005
R18186 vdd.n1308 vdd.n1279 12.8005
R18187 vdd.n1364 vdd.n1326 12.8005
R18188 vdd.n1359 vdd.n1330 12.8005
R18189 vdd.n299 vdd.n272 12.0247
R18190 vdd.n248 vdd.n221 12.0247
R18191 vdd.n205 vdd.n178 12.0247
R18192 vdd.n154 vdd.n127 12.0247
R18193 vdd.n112 vdd.n85 12.0247
R18194 vdd.n61 vdd.n34 12.0247
R18195 vdd.n1494 vdd.n1467 12.0247
R18196 vdd.n1545 vdd.n1518 12.0247
R18197 vdd.n1400 vdd.n1373 12.0247
R18198 vdd.n1451 vdd.n1424 12.0247
R18199 vdd.n1307 vdd.n1280 12.0247
R18200 vdd.n1358 vdd.n1331 12.0247
R18201 vdd.n1215 vdd.n983 11.337
R18202 vdd.n1223 vdd.n972 11.337
R18203 vdd.n1231 vdd.n972 11.337
R18204 vdd.n1239 vdd.n966 11.337
R18205 vdd.n1247 vdd.n959 11.337
R18206 vdd.n1256 vdd.n1255 11.337
R18207 vdd.n1264 vdd.n948 11.337
R18208 vdd.n1562 vdd.n937 11.337
R18209 vdd.n1571 vdd.n931 11.337
R18210 vdd.n1579 vdd.n925 11.337
R18211 vdd.n1588 vdd.n1587 11.337
R18212 vdd.n1596 vdd.n908 11.337
R18213 vdd.n1607 vdd.n908 11.337
R18214 vdd.n1607 vdd.n1606 11.337
R18215 vdd.n2948 vdd.n511 11.337
R18216 vdd.n2948 vdd.n505 11.337
R18217 vdd.n2956 vdd.n505 11.337
R18218 vdd.n2964 vdd.n499 11.337
R18219 vdd.n2972 vdd.n492 11.337
R18220 vdd.n2981 vdd.n2980 11.337
R18221 vdd.n2989 vdd.n481 11.337
R18222 vdd.n3163 vdd.n3162 11.337
R18223 vdd.n3156 vdd.n325 11.337
R18224 vdd.n3154 vdd.n329 11.337
R18225 vdd.n3148 vdd.n3147 11.337
R18226 vdd.n3146 vdd.n340 11.337
R18227 vdd.n3140 vdd.n340 11.337
R18228 vdd.n3139 vdd.n3138 11.337
R18229 vdd.n296 vdd.n295 11.249
R18230 vdd.n245 vdd.n244 11.249
R18231 vdd.n202 vdd.n201 11.249
R18232 vdd.n151 vdd.n150 11.249
R18233 vdd.n109 vdd.n108 11.249
R18234 vdd.n58 vdd.n57 11.249
R18235 vdd.n1491 vdd.n1490 11.249
R18236 vdd.n1542 vdd.n1541 11.249
R18237 vdd.n1397 vdd.n1396 11.249
R18238 vdd.n1448 vdd.n1447 11.249
R18239 vdd.n1304 vdd.n1303 11.249
R18240 vdd.n1355 vdd.n1354 11.249
R18241 vdd.n2244 vdd.t154 11.1103
R18242 vdd.n2576 vdd.t23 11.1103
R18243 vdd.n1231 vdd.t62 10.9969
R18244 vdd.t10 vdd.n3146 10.9969
R18245 vdd.n960 vdd.t50 10.7702
R18246 vdd.t19 vdd.n3155 10.7702
R18247 vdd.n281 vdd.n280 10.7238
R18248 vdd.n230 vdd.n229 10.7238
R18249 vdd.n187 vdd.n186 10.7238
R18250 vdd.n136 vdd.n135 10.7238
R18251 vdd.n94 vdd.n93 10.7238
R18252 vdd.n43 vdd.n42 10.7238
R18253 vdd.n1476 vdd.n1475 10.7238
R18254 vdd.n1527 vdd.n1526 10.7238
R18255 vdd.n1382 vdd.n1381 10.7238
R18256 vdd.n1433 vdd.n1432 10.7238
R18257 vdd.n1289 vdd.n1288 10.7238
R18258 vdd.n1340 vdd.n1339 10.7238
R18259 vdd.n2090 vdd.n2089 10.6151
R18260 vdd.n2091 vdd.n2090 10.6151
R18261 vdd.n2091 vdd.n863 10.6151
R18262 vdd.n2101 vdd.n863 10.6151
R18263 vdd.n2102 vdd.n2101 10.6151
R18264 vdd.n2103 vdd.n2102 10.6151
R18265 vdd.n2103 vdd.n850 10.6151
R18266 vdd.n2114 vdd.n850 10.6151
R18267 vdd.n2115 vdd.n2114 10.6151
R18268 vdd.n2116 vdd.n2115 10.6151
R18269 vdd.n2116 vdd.n838 10.6151
R18270 vdd.n2126 vdd.n838 10.6151
R18271 vdd.n2127 vdd.n2126 10.6151
R18272 vdd.n2128 vdd.n2127 10.6151
R18273 vdd.n2128 vdd.n826 10.6151
R18274 vdd.n2138 vdd.n826 10.6151
R18275 vdd.n2139 vdd.n2138 10.6151
R18276 vdd.n2140 vdd.n2139 10.6151
R18277 vdd.n2140 vdd.n815 10.6151
R18278 vdd.n2150 vdd.n815 10.6151
R18279 vdd.n2151 vdd.n2150 10.6151
R18280 vdd.n2152 vdd.n2151 10.6151
R18281 vdd.n2152 vdd.n802 10.6151
R18282 vdd.n2164 vdd.n802 10.6151
R18283 vdd.n2165 vdd.n2164 10.6151
R18284 vdd.n2167 vdd.n2165 10.6151
R18285 vdd.n2167 vdd.n2166 10.6151
R18286 vdd.n2166 vdd.n784 10.6151
R18287 vdd.n2314 vdd.n2313 10.6151
R18288 vdd.n2313 vdd.n2312 10.6151
R18289 vdd.n2312 vdd.n2309 10.6151
R18290 vdd.n2309 vdd.n2308 10.6151
R18291 vdd.n2308 vdd.n2305 10.6151
R18292 vdd.n2305 vdd.n2304 10.6151
R18293 vdd.n2304 vdd.n2301 10.6151
R18294 vdd.n2301 vdd.n2300 10.6151
R18295 vdd.n2300 vdd.n2297 10.6151
R18296 vdd.n2297 vdd.n2296 10.6151
R18297 vdd.n2296 vdd.n2293 10.6151
R18298 vdd.n2293 vdd.n2292 10.6151
R18299 vdd.n2292 vdd.n2289 10.6151
R18300 vdd.n2289 vdd.n2288 10.6151
R18301 vdd.n2288 vdd.n2285 10.6151
R18302 vdd.n2285 vdd.n2284 10.6151
R18303 vdd.n2284 vdd.n2281 10.6151
R18304 vdd.n2281 vdd.n2280 10.6151
R18305 vdd.n2280 vdd.n2277 10.6151
R18306 vdd.n2277 vdd.n2276 10.6151
R18307 vdd.n2276 vdd.n2273 10.6151
R18308 vdd.n2273 vdd.n2272 10.6151
R18309 vdd.n2272 vdd.n2269 10.6151
R18310 vdd.n2269 vdd.n2268 10.6151
R18311 vdd.n2268 vdd.n2265 10.6151
R18312 vdd.n2265 vdd.n2264 10.6151
R18313 vdd.n2264 vdd.n2261 10.6151
R18314 vdd.n2261 vdd.n2260 10.6151
R18315 vdd.n2260 vdd.n2257 10.6151
R18316 vdd.n2257 vdd.n2256 10.6151
R18317 vdd.n2256 vdd.n2253 10.6151
R18318 vdd.n2251 vdd.n2248 10.6151
R18319 vdd.n2248 vdd.n2247 10.6151
R18320 vdd.n1990 vdd.n1989 10.6151
R18321 vdd.n1989 vdd.n1987 10.6151
R18322 vdd.n1987 vdd.n1986 10.6151
R18323 vdd.n1986 vdd.n1984 10.6151
R18324 vdd.n1984 vdd.n1983 10.6151
R18325 vdd.n1983 vdd.n1981 10.6151
R18326 vdd.n1981 vdd.n1980 10.6151
R18327 vdd.n1980 vdd.n1978 10.6151
R18328 vdd.n1978 vdd.n1977 10.6151
R18329 vdd.n1977 vdd.n1975 10.6151
R18330 vdd.n1975 vdd.n1974 10.6151
R18331 vdd.n1974 vdd.n1972 10.6151
R18332 vdd.n1972 vdd.n1971 10.6151
R18333 vdd.n1971 vdd.n1886 10.6151
R18334 vdd.n1886 vdd.n1885 10.6151
R18335 vdd.n1885 vdd.n1883 10.6151
R18336 vdd.n1883 vdd.n1882 10.6151
R18337 vdd.n1882 vdd.n1880 10.6151
R18338 vdd.n1880 vdd.n1879 10.6151
R18339 vdd.n1879 vdd.n1877 10.6151
R18340 vdd.n1877 vdd.n1876 10.6151
R18341 vdd.n1876 vdd.n1874 10.6151
R18342 vdd.n1874 vdd.n1873 10.6151
R18343 vdd.n1873 vdd.n1871 10.6151
R18344 vdd.n1871 vdd.n1870 10.6151
R18345 vdd.n1870 vdd.n1867 10.6151
R18346 vdd.n1867 vdd.n1866 10.6151
R18347 vdd.n1866 vdd.n787 10.6151
R18348 vdd.n1824 vdd.n875 10.6151
R18349 vdd.n1825 vdd.n1824 10.6151
R18350 vdd.n1826 vdd.n1825 10.6151
R18351 vdd.n1826 vdd.n1820 10.6151
R18352 vdd.n1832 vdd.n1820 10.6151
R18353 vdd.n1833 vdd.n1832 10.6151
R18354 vdd.n1834 vdd.n1833 10.6151
R18355 vdd.n1834 vdd.n1818 10.6151
R18356 vdd.n1840 vdd.n1818 10.6151
R18357 vdd.n1841 vdd.n1840 10.6151
R18358 vdd.n1842 vdd.n1841 10.6151
R18359 vdd.n1842 vdd.n1816 10.6151
R18360 vdd.n1848 vdd.n1816 10.6151
R18361 vdd.n1849 vdd.n1848 10.6151
R18362 vdd.n1850 vdd.n1849 10.6151
R18363 vdd.n1850 vdd.n1814 10.6151
R18364 vdd.n2026 vdd.n1814 10.6151
R18365 vdd.n2026 vdd.n2025 10.6151
R18366 vdd.n2025 vdd.n1855 10.6151
R18367 vdd.n2019 vdd.n1855 10.6151
R18368 vdd.n2019 vdd.n2018 10.6151
R18369 vdd.n2018 vdd.n2017 10.6151
R18370 vdd.n2017 vdd.n1857 10.6151
R18371 vdd.n2011 vdd.n1857 10.6151
R18372 vdd.n2011 vdd.n2010 10.6151
R18373 vdd.n2010 vdd.n2009 10.6151
R18374 vdd.n2009 vdd.n1859 10.6151
R18375 vdd.n2003 vdd.n1859 10.6151
R18376 vdd.n2003 vdd.n2002 10.6151
R18377 vdd.n2002 vdd.n2001 10.6151
R18378 vdd.n2001 vdd.n1861 10.6151
R18379 vdd.n1995 vdd.n1994 10.6151
R18380 vdd.n1994 vdd.n1993 10.6151
R18381 vdd.n2499 vdd.n2498 10.6151
R18382 vdd.n2498 vdd.n2496 10.6151
R18383 vdd.n2496 vdd.n2495 10.6151
R18384 vdd.n2495 vdd.n2353 10.6151
R18385 vdd.n2442 vdd.n2353 10.6151
R18386 vdd.n2443 vdd.n2442 10.6151
R18387 vdd.n2445 vdd.n2443 10.6151
R18388 vdd.n2446 vdd.n2445 10.6151
R18389 vdd.n2448 vdd.n2446 10.6151
R18390 vdd.n2449 vdd.n2448 10.6151
R18391 vdd.n2451 vdd.n2449 10.6151
R18392 vdd.n2452 vdd.n2451 10.6151
R18393 vdd.n2454 vdd.n2452 10.6151
R18394 vdd.n2455 vdd.n2454 10.6151
R18395 vdd.n2470 vdd.n2455 10.6151
R18396 vdd.n2470 vdd.n2469 10.6151
R18397 vdd.n2469 vdd.n2468 10.6151
R18398 vdd.n2468 vdd.n2466 10.6151
R18399 vdd.n2466 vdd.n2465 10.6151
R18400 vdd.n2465 vdd.n2463 10.6151
R18401 vdd.n2463 vdd.n2462 10.6151
R18402 vdd.n2462 vdd.n2460 10.6151
R18403 vdd.n2460 vdd.n2459 10.6151
R18404 vdd.n2459 vdd.n2457 10.6151
R18405 vdd.n2457 vdd.n2456 10.6151
R18406 vdd.n2456 vdd.n664 10.6151
R18407 vdd.n2704 vdd.n664 10.6151
R18408 vdd.n2705 vdd.n2704 10.6151
R18409 vdd.n2566 vdd.n740 10.6151
R18410 vdd.n2566 vdd.n2565 10.6151
R18411 vdd.n2565 vdd.n2564 10.6151
R18412 vdd.n2564 vdd.n2562 10.6151
R18413 vdd.n2562 vdd.n2559 10.6151
R18414 vdd.n2559 vdd.n2558 10.6151
R18415 vdd.n2558 vdd.n2555 10.6151
R18416 vdd.n2555 vdd.n2554 10.6151
R18417 vdd.n2554 vdd.n2551 10.6151
R18418 vdd.n2551 vdd.n2550 10.6151
R18419 vdd.n2550 vdd.n2547 10.6151
R18420 vdd.n2547 vdd.n2546 10.6151
R18421 vdd.n2546 vdd.n2543 10.6151
R18422 vdd.n2543 vdd.n2542 10.6151
R18423 vdd.n2542 vdd.n2539 10.6151
R18424 vdd.n2539 vdd.n2538 10.6151
R18425 vdd.n2538 vdd.n2535 10.6151
R18426 vdd.n2535 vdd.n2534 10.6151
R18427 vdd.n2534 vdd.n2531 10.6151
R18428 vdd.n2531 vdd.n2530 10.6151
R18429 vdd.n2530 vdd.n2527 10.6151
R18430 vdd.n2527 vdd.n2526 10.6151
R18431 vdd.n2526 vdd.n2523 10.6151
R18432 vdd.n2523 vdd.n2522 10.6151
R18433 vdd.n2522 vdd.n2519 10.6151
R18434 vdd.n2519 vdd.n2518 10.6151
R18435 vdd.n2518 vdd.n2515 10.6151
R18436 vdd.n2515 vdd.n2514 10.6151
R18437 vdd.n2514 vdd.n2511 10.6151
R18438 vdd.n2511 vdd.n2510 10.6151
R18439 vdd.n2510 vdd.n2507 10.6151
R18440 vdd.n2505 vdd.n2502 10.6151
R18441 vdd.n2502 vdd.n2501 10.6151
R18442 vdd.n2579 vdd.n2578 10.6151
R18443 vdd.n2580 vdd.n2579 10.6151
R18444 vdd.n2580 vdd.n730 10.6151
R18445 vdd.n2590 vdd.n730 10.6151
R18446 vdd.n2591 vdd.n2590 10.6151
R18447 vdd.n2592 vdd.n2591 10.6151
R18448 vdd.n2592 vdd.n717 10.6151
R18449 vdd.n2602 vdd.n717 10.6151
R18450 vdd.n2603 vdd.n2602 10.6151
R18451 vdd.n2604 vdd.n2603 10.6151
R18452 vdd.n2604 vdd.n706 10.6151
R18453 vdd.n2614 vdd.n706 10.6151
R18454 vdd.n2615 vdd.n2614 10.6151
R18455 vdd.n2616 vdd.n2615 10.6151
R18456 vdd.n2616 vdd.n694 10.6151
R18457 vdd.n2626 vdd.n694 10.6151
R18458 vdd.n2627 vdd.n2626 10.6151
R18459 vdd.n2628 vdd.n2627 10.6151
R18460 vdd.n2628 vdd.n683 10.6151
R18461 vdd.n2640 vdd.n683 10.6151
R18462 vdd.n2641 vdd.n2640 10.6151
R18463 vdd.n2642 vdd.n2641 10.6151
R18464 vdd.n2642 vdd.n669 10.6151
R18465 vdd.n2697 vdd.n669 10.6151
R18466 vdd.n2698 vdd.n2697 10.6151
R18467 vdd.n2699 vdd.n2698 10.6151
R18468 vdd.n2699 vdd.n636 10.6151
R18469 vdd.n2769 vdd.n636 10.6151
R18470 vdd.n2768 vdd.n2767 10.6151
R18471 vdd.n2767 vdd.n637 10.6151
R18472 vdd.n638 vdd.n637 10.6151
R18473 vdd.n2760 vdd.n638 10.6151
R18474 vdd.n2760 vdd.n2759 10.6151
R18475 vdd.n2759 vdd.n2758 10.6151
R18476 vdd.n2758 vdd.n640 10.6151
R18477 vdd.n2753 vdd.n640 10.6151
R18478 vdd.n2753 vdd.n2752 10.6151
R18479 vdd.n2752 vdd.n2751 10.6151
R18480 vdd.n2751 vdd.n643 10.6151
R18481 vdd.n2746 vdd.n643 10.6151
R18482 vdd.n2746 vdd.n2745 10.6151
R18483 vdd.n2745 vdd.n2744 10.6151
R18484 vdd.n2744 vdd.n646 10.6151
R18485 vdd.n2739 vdd.n646 10.6151
R18486 vdd.n2739 vdd.n2738 10.6151
R18487 vdd.n2738 vdd.n2736 10.6151
R18488 vdd.n2736 vdd.n649 10.6151
R18489 vdd.n2731 vdd.n649 10.6151
R18490 vdd.n2731 vdd.n2730 10.6151
R18491 vdd.n2730 vdd.n2729 10.6151
R18492 vdd.n2729 vdd.n652 10.6151
R18493 vdd.n2724 vdd.n652 10.6151
R18494 vdd.n2724 vdd.n2723 10.6151
R18495 vdd.n2723 vdd.n2722 10.6151
R18496 vdd.n2722 vdd.n655 10.6151
R18497 vdd.n2717 vdd.n655 10.6151
R18498 vdd.n2717 vdd.n2716 10.6151
R18499 vdd.n2716 vdd.n2715 10.6151
R18500 vdd.n2715 vdd.n658 10.6151
R18501 vdd.n2710 vdd.n2709 10.6151
R18502 vdd.n2709 vdd.n2708 10.6151
R18503 vdd.n2687 vdd.n2648 10.6151
R18504 vdd.n2682 vdd.n2648 10.6151
R18505 vdd.n2682 vdd.n2681 10.6151
R18506 vdd.n2681 vdd.n2680 10.6151
R18507 vdd.n2680 vdd.n2650 10.6151
R18508 vdd.n2675 vdd.n2650 10.6151
R18509 vdd.n2675 vdd.n2674 10.6151
R18510 vdd.n2674 vdd.n2673 10.6151
R18511 vdd.n2673 vdd.n2653 10.6151
R18512 vdd.n2668 vdd.n2653 10.6151
R18513 vdd.n2668 vdd.n2667 10.6151
R18514 vdd.n2667 vdd.n2666 10.6151
R18515 vdd.n2666 vdd.n2656 10.6151
R18516 vdd.n2661 vdd.n2656 10.6151
R18517 vdd.n2661 vdd.n2660 10.6151
R18518 vdd.n2660 vdd.n610 10.6151
R18519 vdd.n2804 vdd.n610 10.6151
R18520 vdd.n2804 vdd.n611 10.6151
R18521 vdd.n614 vdd.n611 10.6151
R18522 vdd.n2797 vdd.n614 10.6151
R18523 vdd.n2797 vdd.n2796 10.6151
R18524 vdd.n2796 vdd.n2795 10.6151
R18525 vdd.n2795 vdd.n616 10.6151
R18526 vdd.n2790 vdd.n616 10.6151
R18527 vdd.n2790 vdd.n2789 10.6151
R18528 vdd.n2789 vdd.n2788 10.6151
R18529 vdd.n2788 vdd.n619 10.6151
R18530 vdd.n2783 vdd.n619 10.6151
R18531 vdd.n2783 vdd.n2782 10.6151
R18532 vdd.n2782 vdd.n2781 10.6151
R18533 vdd.n2781 vdd.n622 10.6151
R18534 vdd.n2776 vdd.n2775 10.6151
R18535 vdd.n2775 vdd.n2774 10.6151
R18536 vdd.n2422 vdd.n2420 10.6151
R18537 vdd.n2423 vdd.n2422 10.6151
R18538 vdd.n2491 vdd.n2423 10.6151
R18539 vdd.n2491 vdd.n2490 10.6151
R18540 vdd.n2490 vdd.n2489 10.6151
R18541 vdd.n2489 vdd.n2487 10.6151
R18542 vdd.n2487 vdd.n2486 10.6151
R18543 vdd.n2486 vdd.n2484 10.6151
R18544 vdd.n2484 vdd.n2483 10.6151
R18545 vdd.n2483 vdd.n2481 10.6151
R18546 vdd.n2481 vdd.n2480 10.6151
R18547 vdd.n2480 vdd.n2478 10.6151
R18548 vdd.n2478 vdd.n2477 10.6151
R18549 vdd.n2477 vdd.n2475 10.6151
R18550 vdd.n2475 vdd.n2474 10.6151
R18551 vdd.n2474 vdd.n2440 10.6151
R18552 vdd.n2440 vdd.n2439 10.6151
R18553 vdd.n2439 vdd.n2437 10.6151
R18554 vdd.n2437 vdd.n2436 10.6151
R18555 vdd.n2436 vdd.n2434 10.6151
R18556 vdd.n2434 vdd.n2433 10.6151
R18557 vdd.n2433 vdd.n2431 10.6151
R18558 vdd.n2431 vdd.n2430 10.6151
R18559 vdd.n2430 vdd.n2428 10.6151
R18560 vdd.n2428 vdd.n2427 10.6151
R18561 vdd.n2427 vdd.n2425 10.6151
R18562 vdd.n2425 vdd.n2424 10.6151
R18563 vdd.n2424 vdd.n628 10.6151
R18564 vdd.n2573 vdd.n2572 10.6151
R18565 vdd.n2572 vdd.n745 10.6151
R18566 vdd.n2357 vdd.n745 10.6151
R18567 vdd.n2360 vdd.n2357 10.6151
R18568 vdd.n2361 vdd.n2360 10.6151
R18569 vdd.n2364 vdd.n2361 10.6151
R18570 vdd.n2365 vdd.n2364 10.6151
R18571 vdd.n2368 vdd.n2365 10.6151
R18572 vdd.n2369 vdd.n2368 10.6151
R18573 vdd.n2372 vdd.n2369 10.6151
R18574 vdd.n2373 vdd.n2372 10.6151
R18575 vdd.n2376 vdd.n2373 10.6151
R18576 vdd.n2377 vdd.n2376 10.6151
R18577 vdd.n2380 vdd.n2377 10.6151
R18578 vdd.n2381 vdd.n2380 10.6151
R18579 vdd.n2384 vdd.n2381 10.6151
R18580 vdd.n2385 vdd.n2384 10.6151
R18581 vdd.n2388 vdd.n2385 10.6151
R18582 vdd.n2389 vdd.n2388 10.6151
R18583 vdd.n2392 vdd.n2389 10.6151
R18584 vdd.n2393 vdd.n2392 10.6151
R18585 vdd.n2396 vdd.n2393 10.6151
R18586 vdd.n2397 vdd.n2396 10.6151
R18587 vdd.n2400 vdd.n2397 10.6151
R18588 vdd.n2401 vdd.n2400 10.6151
R18589 vdd.n2404 vdd.n2401 10.6151
R18590 vdd.n2405 vdd.n2404 10.6151
R18591 vdd.n2408 vdd.n2405 10.6151
R18592 vdd.n2409 vdd.n2408 10.6151
R18593 vdd.n2412 vdd.n2409 10.6151
R18594 vdd.n2413 vdd.n2412 10.6151
R18595 vdd.n2418 vdd.n2416 10.6151
R18596 vdd.n2419 vdd.n2418 10.6151
R18597 vdd.n2574 vdd.n735 10.6151
R18598 vdd.n2584 vdd.n735 10.6151
R18599 vdd.n2585 vdd.n2584 10.6151
R18600 vdd.n2586 vdd.n2585 10.6151
R18601 vdd.n2586 vdd.n723 10.6151
R18602 vdd.n2596 vdd.n723 10.6151
R18603 vdd.n2597 vdd.n2596 10.6151
R18604 vdd.n2598 vdd.n2597 10.6151
R18605 vdd.n2598 vdd.n712 10.6151
R18606 vdd.n2608 vdd.n712 10.6151
R18607 vdd.n2609 vdd.n2608 10.6151
R18608 vdd.n2610 vdd.n2609 10.6151
R18609 vdd.n2610 vdd.n700 10.6151
R18610 vdd.n2620 vdd.n700 10.6151
R18611 vdd.n2621 vdd.n2620 10.6151
R18612 vdd.n2622 vdd.n2621 10.6151
R18613 vdd.n2622 vdd.n689 10.6151
R18614 vdd.n2632 vdd.n689 10.6151
R18615 vdd.n2633 vdd.n2632 10.6151
R18616 vdd.n2636 vdd.n2633 10.6151
R18617 vdd.n2646 vdd.n677 10.6151
R18618 vdd.n2647 vdd.n2646 10.6151
R18619 vdd.n2693 vdd.n2647 10.6151
R18620 vdd.n2693 vdd.n2692 10.6151
R18621 vdd.n2692 vdd.n2691 10.6151
R18622 vdd.n2691 vdd.n2690 10.6151
R18623 vdd.n2690 vdd.n2688 10.6151
R18624 vdd.n2085 vdd.n869 10.6151
R18625 vdd.n2095 vdd.n869 10.6151
R18626 vdd.n2096 vdd.n2095 10.6151
R18627 vdd.n2097 vdd.n2096 10.6151
R18628 vdd.n2097 vdd.n856 10.6151
R18629 vdd.n2107 vdd.n856 10.6151
R18630 vdd.n2108 vdd.n2107 10.6151
R18631 vdd.n2110 vdd.n844 10.6151
R18632 vdd.n2120 vdd.n844 10.6151
R18633 vdd.n2121 vdd.n2120 10.6151
R18634 vdd.n2122 vdd.n2121 10.6151
R18635 vdd.n2122 vdd.n832 10.6151
R18636 vdd.n2132 vdd.n832 10.6151
R18637 vdd.n2133 vdd.n2132 10.6151
R18638 vdd.n2134 vdd.n2133 10.6151
R18639 vdd.n2134 vdd.n821 10.6151
R18640 vdd.n2144 vdd.n821 10.6151
R18641 vdd.n2145 vdd.n2144 10.6151
R18642 vdd.n2146 vdd.n2145 10.6151
R18643 vdd.n2146 vdd.n809 10.6151
R18644 vdd.n2156 vdd.n809 10.6151
R18645 vdd.n2157 vdd.n2156 10.6151
R18646 vdd.n2160 vdd.n2157 10.6151
R18647 vdd.n2160 vdd.n2159 10.6151
R18648 vdd.n2159 vdd.n2158 10.6151
R18649 vdd.n2158 vdd.n792 10.6151
R18650 vdd.n2242 vdd.n792 10.6151
R18651 vdd.n2241 vdd.n2240 10.6151
R18652 vdd.n2240 vdd.n2237 10.6151
R18653 vdd.n2237 vdd.n2236 10.6151
R18654 vdd.n2236 vdd.n2233 10.6151
R18655 vdd.n2233 vdd.n2232 10.6151
R18656 vdd.n2232 vdd.n2229 10.6151
R18657 vdd.n2229 vdd.n2228 10.6151
R18658 vdd.n2228 vdd.n2225 10.6151
R18659 vdd.n2225 vdd.n2224 10.6151
R18660 vdd.n2224 vdd.n2221 10.6151
R18661 vdd.n2221 vdd.n2220 10.6151
R18662 vdd.n2220 vdd.n2217 10.6151
R18663 vdd.n2217 vdd.n2216 10.6151
R18664 vdd.n2216 vdd.n2213 10.6151
R18665 vdd.n2213 vdd.n2212 10.6151
R18666 vdd.n2212 vdd.n2209 10.6151
R18667 vdd.n2209 vdd.n2208 10.6151
R18668 vdd.n2208 vdd.n2205 10.6151
R18669 vdd.n2205 vdd.n2204 10.6151
R18670 vdd.n2204 vdd.n2201 10.6151
R18671 vdd.n2201 vdd.n2200 10.6151
R18672 vdd.n2200 vdd.n2197 10.6151
R18673 vdd.n2197 vdd.n2196 10.6151
R18674 vdd.n2196 vdd.n2193 10.6151
R18675 vdd.n2193 vdd.n2192 10.6151
R18676 vdd.n2192 vdd.n2189 10.6151
R18677 vdd.n2189 vdd.n2188 10.6151
R18678 vdd.n2188 vdd.n2185 10.6151
R18679 vdd.n2185 vdd.n2184 10.6151
R18680 vdd.n2184 vdd.n2181 10.6151
R18681 vdd.n2181 vdd.n2180 10.6151
R18682 vdd.n2177 vdd.n2176 10.6151
R18683 vdd.n2176 vdd.n2174 10.6151
R18684 vdd.n1933 vdd.n1931 10.6151
R18685 vdd.n1934 vdd.n1933 10.6151
R18686 vdd.n1936 vdd.n1934 10.6151
R18687 vdd.n1937 vdd.n1936 10.6151
R18688 vdd.n1939 vdd.n1937 10.6151
R18689 vdd.n1940 vdd.n1939 10.6151
R18690 vdd.n1942 vdd.n1940 10.6151
R18691 vdd.n1943 vdd.n1942 10.6151
R18692 vdd.n1945 vdd.n1943 10.6151
R18693 vdd.n1946 vdd.n1945 10.6151
R18694 vdd.n1948 vdd.n1946 10.6151
R18695 vdd.n1949 vdd.n1948 10.6151
R18696 vdd.n1967 vdd.n1949 10.6151
R18697 vdd.n1967 vdd.n1966 10.6151
R18698 vdd.n1966 vdd.n1965 10.6151
R18699 vdd.n1965 vdd.n1963 10.6151
R18700 vdd.n1963 vdd.n1962 10.6151
R18701 vdd.n1962 vdd.n1960 10.6151
R18702 vdd.n1960 vdd.n1959 10.6151
R18703 vdd.n1959 vdd.n1957 10.6151
R18704 vdd.n1957 vdd.n1956 10.6151
R18705 vdd.n1956 vdd.n1954 10.6151
R18706 vdd.n1954 vdd.n1953 10.6151
R18707 vdd.n1953 vdd.n1951 10.6151
R18708 vdd.n1951 vdd.n1950 10.6151
R18709 vdd.n1950 vdd.n796 10.6151
R18710 vdd.n2172 vdd.n796 10.6151
R18711 vdd.n2173 vdd.n2172 10.6151
R18712 vdd.n2084 vdd.n2083 10.6151
R18713 vdd.n2083 vdd.n881 10.6151
R18714 vdd.n2077 vdd.n881 10.6151
R18715 vdd.n2077 vdd.n2076 10.6151
R18716 vdd.n2076 vdd.n2075 10.6151
R18717 vdd.n2075 vdd.n883 10.6151
R18718 vdd.n2069 vdd.n883 10.6151
R18719 vdd.n2069 vdd.n2068 10.6151
R18720 vdd.n2068 vdd.n2067 10.6151
R18721 vdd.n2067 vdd.n885 10.6151
R18722 vdd.n2061 vdd.n885 10.6151
R18723 vdd.n2061 vdd.n2060 10.6151
R18724 vdd.n2060 vdd.n2059 10.6151
R18725 vdd.n2059 vdd.n887 10.6151
R18726 vdd.n2053 vdd.n887 10.6151
R18727 vdd.n2053 vdd.n2052 10.6151
R18728 vdd.n2052 vdd.n2051 10.6151
R18729 vdd.n2051 vdd.n891 10.6151
R18730 vdd.n1899 vdd.n891 10.6151
R18731 vdd.n1900 vdd.n1899 10.6151
R18732 vdd.n1900 vdd.n1895 10.6151
R18733 vdd.n1906 vdd.n1895 10.6151
R18734 vdd.n1907 vdd.n1906 10.6151
R18735 vdd.n1908 vdd.n1907 10.6151
R18736 vdd.n1908 vdd.n1893 10.6151
R18737 vdd.n1914 vdd.n1893 10.6151
R18738 vdd.n1915 vdd.n1914 10.6151
R18739 vdd.n1916 vdd.n1915 10.6151
R18740 vdd.n1916 vdd.n1891 10.6151
R18741 vdd.n1922 vdd.n1891 10.6151
R18742 vdd.n1923 vdd.n1922 10.6151
R18743 vdd.n1925 vdd.n1887 10.6151
R18744 vdd.n1930 vdd.n1887 10.6151
R18745 vdd.n1272 vdd.t8 10.5435
R18746 vdd.n2041 vdd.t84 10.5435
R18747 vdd.n2940 vdd.t77 10.5435
R18748 vdd.n3164 vdd.t191 10.5435
R18749 vdd.n292 vdd.n274 10.4732
R18750 vdd.n241 vdd.n223 10.4732
R18751 vdd.n198 vdd.n180 10.4732
R18752 vdd.n147 vdd.n129 10.4732
R18753 vdd.n105 vdd.n87 10.4732
R18754 vdd.n54 vdd.n36 10.4732
R18755 vdd.n1487 vdd.n1469 10.4732
R18756 vdd.n1538 vdd.n1520 10.4732
R18757 vdd.n1393 vdd.n1375 10.4732
R18758 vdd.n1444 vdd.n1426 10.4732
R18759 vdd.n1300 vdd.n1282 10.4732
R18760 vdd.n1351 vdd.n1333 10.4732
R18761 vdd.n1570 vdd.t30 10.3167
R18762 vdd.t52 vdd.n493 10.3167
R18763 vdd.n1223 vdd.t88 9.86327
R18764 vdd.n3140 vdd.t137 9.86327
R18765 vdd.n291 vdd.n276 9.69747
R18766 vdd.n240 vdd.n225 9.69747
R18767 vdd.n197 vdd.n182 9.69747
R18768 vdd.n146 vdd.n131 9.69747
R18769 vdd.n104 vdd.n89 9.69747
R18770 vdd.n53 vdd.n38 9.69747
R18771 vdd.n1486 vdd.n1471 9.69747
R18772 vdd.n1537 vdd.n1522 9.69747
R18773 vdd.n1392 vdd.n1377 9.69747
R18774 vdd.n1443 vdd.n1428 9.69747
R18775 vdd.n1299 vdd.n1284 9.69747
R18776 vdd.n1350 vdd.n1335 9.69747
R18777 vdd.n2027 vdd.n2026 9.67831
R18778 vdd.n2738 vdd.n2737 9.67831
R18779 vdd.n2805 vdd.n2804 9.67831
R18780 vdd.n2051 vdd.n2050 9.67831
R18781 vdd.n307 vdd.n306 9.45567
R18782 vdd.n256 vdd.n255 9.45567
R18783 vdd.n213 vdd.n212 9.45567
R18784 vdd.n162 vdd.n161 9.45567
R18785 vdd.n120 vdd.n119 9.45567
R18786 vdd.n69 vdd.n68 9.45567
R18787 vdd.n1502 vdd.n1501 9.45567
R18788 vdd.n1553 vdd.n1552 9.45567
R18789 vdd.n1408 vdd.n1407 9.45567
R18790 vdd.n1459 vdd.n1458 9.45567
R18791 vdd.n1315 vdd.n1314 9.45567
R18792 vdd.n1366 vdd.n1365 9.45567
R18793 vdd.n1787 vdd.n1641 9.3005
R18794 vdd.n1786 vdd.n1785 9.3005
R18795 vdd.n1647 vdd.n1646 9.3005
R18796 vdd.n1780 vdd.n1651 9.3005
R18797 vdd.n1779 vdd.n1652 9.3005
R18798 vdd.n1778 vdd.n1653 9.3005
R18799 vdd.n1657 vdd.n1654 9.3005
R18800 vdd.n1773 vdd.n1658 9.3005
R18801 vdd.n1772 vdd.n1659 9.3005
R18802 vdd.n1771 vdd.n1660 9.3005
R18803 vdd.n1664 vdd.n1661 9.3005
R18804 vdd.n1766 vdd.n1665 9.3005
R18805 vdd.n1765 vdd.n1666 9.3005
R18806 vdd.n1764 vdd.n1667 9.3005
R18807 vdd.n1671 vdd.n1668 9.3005
R18808 vdd.n1759 vdd.n1672 9.3005
R18809 vdd.n1758 vdd.n1673 9.3005
R18810 vdd.n1757 vdd.n1674 9.3005
R18811 vdd.n1678 vdd.n1675 9.3005
R18812 vdd.n1752 vdd.n1679 9.3005
R18813 vdd.n1751 vdd.n1680 9.3005
R18814 vdd.n1750 vdd.n1749 9.3005
R18815 vdd.n1748 vdd.n1681 9.3005
R18816 vdd.n1747 vdd.n1746 9.3005
R18817 vdd.n1687 vdd.n1686 9.3005
R18818 vdd.n1741 vdd.n1691 9.3005
R18819 vdd.n1740 vdd.n1692 9.3005
R18820 vdd.n1739 vdd.n1693 9.3005
R18821 vdd.n1697 vdd.n1694 9.3005
R18822 vdd.n1734 vdd.n1698 9.3005
R18823 vdd.n1733 vdd.n1699 9.3005
R18824 vdd.n1732 vdd.n1700 9.3005
R18825 vdd.n1704 vdd.n1701 9.3005
R18826 vdd.n1727 vdd.n1705 9.3005
R18827 vdd.n1726 vdd.n1706 9.3005
R18828 vdd.n1725 vdd.n1707 9.3005
R18829 vdd.n1709 vdd.n1708 9.3005
R18830 vdd.n1720 vdd.n892 9.3005
R18831 vdd.n1789 vdd.n1788 9.3005
R18832 vdd.n1813 vdd.n1812 9.3005
R18833 vdd.n1619 vdd.n1618 9.3005
R18834 vdd.n1624 vdd.n1622 9.3005
R18835 vdd.n1805 vdd.n1625 9.3005
R18836 vdd.n1804 vdd.n1626 9.3005
R18837 vdd.n1803 vdd.n1627 9.3005
R18838 vdd.n1631 vdd.n1628 9.3005
R18839 vdd.n1798 vdd.n1632 9.3005
R18840 vdd.n1797 vdd.n1633 9.3005
R18841 vdd.n1796 vdd.n1634 9.3005
R18842 vdd.n1638 vdd.n1635 9.3005
R18843 vdd.n1791 vdd.n1639 9.3005
R18844 vdd.n1790 vdd.n1640 9.3005
R18845 vdd.n2035 vdd.n1612 9.3005
R18846 vdd.n2037 vdd.n2036 9.3005
R18847 vdd.n1558 vdd.n939 9.3005
R18848 vdd.n1560 vdd.n1559 9.3005
R18849 vdd.n929 vdd.n928 9.3005
R18850 vdd.n1574 vdd.n1573 9.3005
R18851 vdd.n1575 vdd.n927 9.3005
R18852 vdd.n1577 vdd.n1576 9.3005
R18853 vdd.n918 vdd.n917 9.3005
R18854 vdd.n1591 vdd.n1590 9.3005
R18855 vdd.n1592 vdd.n916 9.3005
R18856 vdd.n1594 vdd.n1593 9.3005
R18857 vdd.n906 vdd.n905 9.3005
R18858 vdd.n1610 vdd.n1609 9.3005
R18859 vdd.n1611 vdd.n904 9.3005
R18860 vdd.n2039 vdd.n2038 9.3005
R18861 vdd.n283 vdd.n282 9.3005
R18862 vdd.n278 vdd.n277 9.3005
R18863 vdd.n289 vdd.n288 9.3005
R18864 vdd.n291 vdd.n290 9.3005
R18865 vdd.n274 vdd.n273 9.3005
R18866 vdd.n297 vdd.n296 9.3005
R18867 vdd.n299 vdd.n298 9.3005
R18868 vdd.n271 vdd.n268 9.3005
R18869 vdd.n306 vdd.n305 9.3005
R18870 vdd.n232 vdd.n231 9.3005
R18871 vdd.n227 vdd.n226 9.3005
R18872 vdd.n238 vdd.n237 9.3005
R18873 vdd.n240 vdd.n239 9.3005
R18874 vdd.n223 vdd.n222 9.3005
R18875 vdd.n246 vdd.n245 9.3005
R18876 vdd.n248 vdd.n247 9.3005
R18877 vdd.n220 vdd.n217 9.3005
R18878 vdd.n255 vdd.n254 9.3005
R18879 vdd.n189 vdd.n188 9.3005
R18880 vdd.n184 vdd.n183 9.3005
R18881 vdd.n195 vdd.n194 9.3005
R18882 vdd.n197 vdd.n196 9.3005
R18883 vdd.n180 vdd.n179 9.3005
R18884 vdd.n203 vdd.n202 9.3005
R18885 vdd.n205 vdd.n204 9.3005
R18886 vdd.n177 vdd.n174 9.3005
R18887 vdd.n212 vdd.n211 9.3005
R18888 vdd.n138 vdd.n137 9.3005
R18889 vdd.n133 vdd.n132 9.3005
R18890 vdd.n144 vdd.n143 9.3005
R18891 vdd.n146 vdd.n145 9.3005
R18892 vdd.n129 vdd.n128 9.3005
R18893 vdd.n152 vdd.n151 9.3005
R18894 vdd.n154 vdd.n153 9.3005
R18895 vdd.n126 vdd.n123 9.3005
R18896 vdd.n161 vdd.n160 9.3005
R18897 vdd.n96 vdd.n95 9.3005
R18898 vdd.n91 vdd.n90 9.3005
R18899 vdd.n102 vdd.n101 9.3005
R18900 vdd.n104 vdd.n103 9.3005
R18901 vdd.n87 vdd.n86 9.3005
R18902 vdd.n110 vdd.n109 9.3005
R18903 vdd.n112 vdd.n111 9.3005
R18904 vdd.n84 vdd.n81 9.3005
R18905 vdd.n119 vdd.n118 9.3005
R18906 vdd.n45 vdd.n44 9.3005
R18907 vdd.n40 vdd.n39 9.3005
R18908 vdd.n51 vdd.n50 9.3005
R18909 vdd.n53 vdd.n52 9.3005
R18910 vdd.n36 vdd.n35 9.3005
R18911 vdd.n59 vdd.n58 9.3005
R18912 vdd.n61 vdd.n60 9.3005
R18913 vdd.n33 vdd.n30 9.3005
R18914 vdd.n68 vdd.n67 9.3005
R18915 vdd.n2854 vdd.n2853 9.3005
R18916 vdd.n2855 vdd.n578 9.3005
R18917 vdd.n577 vdd.n575 9.3005
R18918 vdd.n2861 vdd.n574 9.3005
R18919 vdd.n2862 vdd.n573 9.3005
R18920 vdd.n2863 vdd.n572 9.3005
R18921 vdd.n571 vdd.n569 9.3005
R18922 vdd.n2869 vdd.n568 9.3005
R18923 vdd.n2870 vdd.n567 9.3005
R18924 vdd.n2871 vdd.n566 9.3005
R18925 vdd.n565 vdd.n563 9.3005
R18926 vdd.n2877 vdd.n562 9.3005
R18927 vdd.n2878 vdd.n561 9.3005
R18928 vdd.n2879 vdd.n560 9.3005
R18929 vdd.n559 vdd.n557 9.3005
R18930 vdd.n2885 vdd.n556 9.3005
R18931 vdd.n2886 vdd.n555 9.3005
R18932 vdd.n2887 vdd.n554 9.3005
R18933 vdd.n553 vdd.n551 9.3005
R18934 vdd.n2893 vdd.n550 9.3005
R18935 vdd.n2894 vdd.n549 9.3005
R18936 vdd.n2895 vdd.n548 9.3005
R18937 vdd.n547 vdd.n545 9.3005
R18938 vdd.n2901 vdd.n542 9.3005
R18939 vdd.n2902 vdd.n541 9.3005
R18940 vdd.n2903 vdd.n540 9.3005
R18941 vdd.n539 vdd.n537 9.3005
R18942 vdd.n2909 vdd.n536 9.3005
R18943 vdd.n2910 vdd.n535 9.3005
R18944 vdd.n2911 vdd.n534 9.3005
R18945 vdd.n533 vdd.n531 9.3005
R18946 vdd.n2917 vdd.n530 9.3005
R18947 vdd.n2918 vdd.n529 9.3005
R18948 vdd.n2919 vdd.n528 9.3005
R18949 vdd.n527 vdd.n525 9.3005
R18950 vdd.n2924 vdd.n524 9.3005
R18951 vdd.n2934 vdd.n518 9.3005
R18952 vdd.n2936 vdd.n2935 9.3005
R18953 vdd.n509 vdd.n508 9.3005
R18954 vdd.n2951 vdd.n2950 9.3005
R18955 vdd.n2952 vdd.n507 9.3005
R18956 vdd.n2954 vdd.n2953 9.3005
R18957 vdd.n497 vdd.n496 9.3005
R18958 vdd.n2967 vdd.n2966 9.3005
R18959 vdd.n2968 vdd.n495 9.3005
R18960 vdd.n2970 vdd.n2969 9.3005
R18961 vdd.n485 vdd.n484 9.3005
R18962 vdd.n2984 vdd.n2983 9.3005
R18963 vdd.n2985 vdd.n483 9.3005
R18964 vdd.n2987 vdd.n2986 9.3005
R18965 vdd.n312 vdd.n310 9.3005
R18966 vdd.n2938 vdd.n2937 9.3005
R18967 vdd.n3167 vdd.n3166 9.3005
R18968 vdd.n313 vdd.n311 9.3005
R18969 vdd.n3160 vdd.n320 9.3005
R18970 vdd.n3159 vdd.n321 9.3005
R18971 vdd.n3158 vdd.n322 9.3005
R18972 vdd.n331 vdd.n323 9.3005
R18973 vdd.n3152 vdd.n332 9.3005
R18974 vdd.n3151 vdd.n333 9.3005
R18975 vdd.n3150 vdd.n334 9.3005
R18976 vdd.n342 vdd.n335 9.3005
R18977 vdd.n3144 vdd.n343 9.3005
R18978 vdd.n3143 vdd.n344 9.3005
R18979 vdd.n3142 vdd.n345 9.3005
R18980 vdd.n353 vdd.n346 9.3005
R18981 vdd.n3136 vdd.n3135 9.3005
R18982 vdd.n3132 vdd.n354 9.3005
R18983 vdd.n3131 vdd.n357 9.3005
R18984 vdd.n361 vdd.n358 9.3005
R18985 vdd.n362 vdd.n359 9.3005
R18986 vdd.n3124 vdd.n363 9.3005
R18987 vdd.n3123 vdd.n364 9.3005
R18988 vdd.n3122 vdd.n365 9.3005
R18989 vdd.n369 vdd.n366 9.3005
R18990 vdd.n3117 vdd.n370 9.3005
R18991 vdd.n3116 vdd.n371 9.3005
R18992 vdd.n3115 vdd.n372 9.3005
R18993 vdd.n376 vdd.n373 9.3005
R18994 vdd.n3110 vdd.n377 9.3005
R18995 vdd.n3109 vdd.n378 9.3005
R18996 vdd.n3108 vdd.n379 9.3005
R18997 vdd.n383 vdd.n380 9.3005
R18998 vdd.n3103 vdd.n384 9.3005
R18999 vdd.n3102 vdd.n385 9.3005
R19000 vdd.n3101 vdd.n3100 9.3005
R19001 vdd.n3099 vdd.n386 9.3005
R19002 vdd.n3098 vdd.n3097 9.3005
R19003 vdd.n392 vdd.n391 9.3005
R19004 vdd.n3092 vdd.n396 9.3005
R19005 vdd.n3091 vdd.n397 9.3005
R19006 vdd.n3090 vdd.n398 9.3005
R19007 vdd.n402 vdd.n399 9.3005
R19008 vdd.n3085 vdd.n403 9.3005
R19009 vdd.n3084 vdd.n404 9.3005
R19010 vdd.n3083 vdd.n405 9.3005
R19011 vdd.n409 vdd.n406 9.3005
R19012 vdd.n3078 vdd.n410 9.3005
R19013 vdd.n3077 vdd.n411 9.3005
R19014 vdd.n3076 vdd.n412 9.3005
R19015 vdd.n416 vdd.n413 9.3005
R19016 vdd.n3071 vdd.n417 9.3005
R19017 vdd.n3070 vdd.n418 9.3005
R19018 vdd.n3069 vdd.n419 9.3005
R19019 vdd.n423 vdd.n420 9.3005
R19020 vdd.n3064 vdd.n424 9.3005
R19021 vdd.n3063 vdd.n425 9.3005
R19022 vdd.n3062 vdd.n3061 9.3005
R19023 vdd.n3060 vdd.n426 9.3005
R19024 vdd.n3059 vdd.n3058 9.3005
R19025 vdd.n432 vdd.n431 9.3005
R19026 vdd.n3053 vdd.n436 9.3005
R19027 vdd.n3052 vdd.n437 9.3005
R19028 vdd.n3051 vdd.n438 9.3005
R19029 vdd.n442 vdd.n439 9.3005
R19030 vdd.n3046 vdd.n443 9.3005
R19031 vdd.n3045 vdd.n444 9.3005
R19032 vdd.n3044 vdd.n445 9.3005
R19033 vdd.n449 vdd.n446 9.3005
R19034 vdd.n3039 vdd.n450 9.3005
R19035 vdd.n3038 vdd.n451 9.3005
R19036 vdd.n3037 vdd.n452 9.3005
R19037 vdd.n456 vdd.n453 9.3005
R19038 vdd.n3032 vdd.n457 9.3005
R19039 vdd.n3031 vdd.n458 9.3005
R19040 vdd.n3030 vdd.n459 9.3005
R19041 vdd.n463 vdd.n460 9.3005
R19042 vdd.n3025 vdd.n464 9.3005
R19043 vdd.n3024 vdd.n465 9.3005
R19044 vdd.n3020 vdd.n3017 9.3005
R19045 vdd.n3134 vdd.n3133 9.3005
R19046 vdd.n2944 vdd.n513 9.3005
R19047 vdd.n2946 vdd.n2945 9.3005
R19048 vdd.n503 vdd.n502 9.3005
R19049 vdd.n2959 vdd.n2958 9.3005
R19050 vdd.n2960 vdd.n501 9.3005
R19051 vdd.n2962 vdd.n2961 9.3005
R19052 vdd.n490 vdd.n489 9.3005
R19053 vdd.n2975 vdd.n2974 9.3005
R19054 vdd.n2976 vdd.n488 9.3005
R19055 vdd.n2978 vdd.n2977 9.3005
R19056 vdd.n478 vdd.n477 9.3005
R19057 vdd.n2992 vdd.n2991 9.3005
R19058 vdd.n2993 vdd.n476 9.3005
R19059 vdd.n2995 vdd.n2994 9.3005
R19060 vdd.n2996 vdd.n475 9.3005
R19061 vdd.n2998 vdd.n2997 9.3005
R19062 vdd.n2999 vdd.n474 9.3005
R19063 vdd.n3001 vdd.n3000 9.3005
R19064 vdd.n3002 vdd.n472 9.3005
R19065 vdd.n3004 vdd.n3003 9.3005
R19066 vdd.n3005 vdd.n471 9.3005
R19067 vdd.n3007 vdd.n3006 9.3005
R19068 vdd.n3008 vdd.n469 9.3005
R19069 vdd.n3010 vdd.n3009 9.3005
R19070 vdd.n3011 vdd.n468 9.3005
R19071 vdd.n3013 vdd.n3012 9.3005
R19072 vdd.n3014 vdd.n466 9.3005
R19073 vdd.n3016 vdd.n3015 9.3005
R19074 vdd.n2943 vdd.n2942 9.3005
R19075 vdd.n2807 vdd.n514 9.3005
R19076 vdd.n2812 vdd.n2806 9.3005
R19077 vdd.n2822 vdd.n605 9.3005
R19078 vdd.n2823 vdd.n604 9.3005
R19079 vdd.n603 vdd.n601 9.3005
R19080 vdd.n2829 vdd.n600 9.3005
R19081 vdd.n2830 vdd.n599 9.3005
R19082 vdd.n2831 vdd.n598 9.3005
R19083 vdd.n597 vdd.n595 9.3005
R19084 vdd.n2837 vdd.n594 9.3005
R19085 vdd.n2838 vdd.n593 9.3005
R19086 vdd.n2839 vdd.n592 9.3005
R19087 vdd.n591 vdd.n589 9.3005
R19088 vdd.n2844 vdd.n588 9.3005
R19089 vdd.n2845 vdd.n587 9.3005
R19090 vdd.n583 vdd.n582 9.3005
R19091 vdd.n2851 vdd.n2850 9.3005
R19092 vdd.n2852 vdd.n579 9.3005
R19093 vdd.n2049 vdd.n2048 9.3005
R19094 vdd.n2044 vdd.n895 9.3005
R19095 vdd.n1219 vdd.n979 9.3005
R19096 vdd.n1221 vdd.n1220 9.3005
R19097 vdd.n970 vdd.n969 9.3005
R19098 vdd.n1234 vdd.n1233 9.3005
R19099 vdd.n1235 vdd.n968 9.3005
R19100 vdd.n1237 vdd.n1236 9.3005
R19101 vdd.n957 vdd.n956 9.3005
R19102 vdd.n1250 vdd.n1249 9.3005
R19103 vdd.n1251 vdd.n955 9.3005
R19104 vdd.n1253 vdd.n1252 9.3005
R19105 vdd.n946 vdd.n945 9.3005
R19106 vdd.n1267 vdd.n1266 9.3005
R19107 vdd.n1268 vdd.n944 9.3005
R19108 vdd.n1270 vdd.n1269 9.3005
R19109 vdd.n935 vdd.n934 9.3005
R19110 vdd.n1565 vdd.n1564 9.3005
R19111 vdd.n1566 vdd.n933 9.3005
R19112 vdd.n1568 vdd.n1567 9.3005
R19113 vdd.n923 vdd.n922 9.3005
R19114 vdd.n1582 vdd.n1581 9.3005
R19115 vdd.n1583 vdd.n921 9.3005
R19116 vdd.n1585 vdd.n1584 9.3005
R19117 vdd.n913 vdd.n912 9.3005
R19118 vdd.n1599 vdd.n1598 9.3005
R19119 vdd.n1600 vdd.n910 9.3005
R19120 vdd.n1604 vdd.n1603 9.3005
R19121 vdd.n1602 vdd.n911 9.3005
R19122 vdd.n1601 vdd.n900 9.3005
R19123 vdd.n1218 vdd.n1217 9.3005
R19124 vdd.n1113 vdd.n1103 9.3005
R19125 vdd.n1115 vdd.n1114 9.3005
R19126 vdd.n1116 vdd.n1102 9.3005
R19127 vdd.n1118 vdd.n1117 9.3005
R19128 vdd.n1119 vdd.n1095 9.3005
R19129 vdd.n1121 vdd.n1120 9.3005
R19130 vdd.n1122 vdd.n1094 9.3005
R19131 vdd.n1124 vdd.n1123 9.3005
R19132 vdd.n1125 vdd.n1087 9.3005
R19133 vdd.n1127 vdd.n1126 9.3005
R19134 vdd.n1128 vdd.n1086 9.3005
R19135 vdd.n1130 vdd.n1129 9.3005
R19136 vdd.n1131 vdd.n1079 9.3005
R19137 vdd.n1133 vdd.n1132 9.3005
R19138 vdd.n1134 vdd.n1078 9.3005
R19139 vdd.n1136 vdd.n1135 9.3005
R19140 vdd.n1137 vdd.n1072 9.3005
R19141 vdd.n1139 vdd.n1138 9.3005
R19142 vdd.n1140 vdd.n1070 9.3005
R19143 vdd.n1142 vdd.n1141 9.3005
R19144 vdd.n1071 vdd.n1068 9.3005
R19145 vdd.n1149 vdd.n1064 9.3005
R19146 vdd.n1151 vdd.n1150 9.3005
R19147 vdd.n1152 vdd.n1063 9.3005
R19148 vdd.n1154 vdd.n1153 9.3005
R19149 vdd.n1155 vdd.n1056 9.3005
R19150 vdd.n1157 vdd.n1156 9.3005
R19151 vdd.n1158 vdd.n1055 9.3005
R19152 vdd.n1160 vdd.n1159 9.3005
R19153 vdd.n1161 vdd.n1048 9.3005
R19154 vdd.n1163 vdd.n1162 9.3005
R19155 vdd.n1164 vdd.n1047 9.3005
R19156 vdd.n1166 vdd.n1165 9.3005
R19157 vdd.n1167 vdd.n1040 9.3005
R19158 vdd.n1169 vdd.n1168 9.3005
R19159 vdd.n1170 vdd.n1039 9.3005
R19160 vdd.n1172 vdd.n1171 9.3005
R19161 vdd.n1173 vdd.n1032 9.3005
R19162 vdd.n1175 vdd.n1174 9.3005
R19163 vdd.n1176 vdd.n1031 9.3005
R19164 vdd.n1178 vdd.n1177 9.3005
R19165 vdd.n1179 vdd.n1024 9.3005
R19166 vdd.n1181 vdd.n1180 9.3005
R19167 vdd.n1182 vdd.n1023 9.3005
R19168 vdd.n1184 vdd.n1183 9.3005
R19169 vdd.n1185 vdd.n1014 9.3005
R19170 vdd.n1187 vdd.n1186 9.3005
R19171 vdd.n1188 vdd.n1013 9.3005
R19172 vdd.n1190 vdd.n1189 9.3005
R19173 vdd.n1191 vdd.n1006 9.3005
R19174 vdd.n1193 vdd.n1192 9.3005
R19175 vdd.n1194 vdd.n1005 9.3005
R19176 vdd.n1196 vdd.n1195 9.3005
R19177 vdd.n1197 vdd.n998 9.3005
R19178 vdd.n1199 vdd.n1198 9.3005
R19179 vdd.n1200 vdd.n997 9.3005
R19180 vdd.n1202 vdd.n1201 9.3005
R19181 vdd.n1203 vdd.n990 9.3005
R19182 vdd.n1205 vdd.n1204 9.3005
R19183 vdd.n1206 vdd.n989 9.3005
R19184 vdd.n1208 vdd.n1207 9.3005
R19185 vdd.n1209 vdd.n985 9.3005
R19186 vdd.n1211 vdd.n1210 9.3005
R19187 vdd.n1109 vdd.n980 9.3005
R19188 vdd.n976 vdd.n975 9.3005
R19189 vdd.n1226 vdd.n1225 9.3005
R19190 vdd.n1227 vdd.n974 9.3005
R19191 vdd.n1229 vdd.n1228 9.3005
R19192 vdd.n964 vdd.n963 9.3005
R19193 vdd.n1242 vdd.n1241 9.3005
R19194 vdd.n1243 vdd.n962 9.3005
R19195 vdd.n1245 vdd.n1244 9.3005
R19196 vdd.n952 vdd.n951 9.3005
R19197 vdd.n1259 vdd.n1258 9.3005
R19198 vdd.n1260 vdd.n950 9.3005
R19199 vdd.n1262 vdd.n1261 9.3005
R19200 vdd.n941 vdd.n940 9.3005
R19201 vdd.n1213 vdd.n1212 9.3005
R19202 vdd.n1557 vdd.n1274 9.3005
R19203 vdd.n1478 vdd.n1477 9.3005
R19204 vdd.n1473 vdd.n1472 9.3005
R19205 vdd.n1484 vdd.n1483 9.3005
R19206 vdd.n1486 vdd.n1485 9.3005
R19207 vdd.n1469 vdd.n1468 9.3005
R19208 vdd.n1492 vdd.n1491 9.3005
R19209 vdd.n1494 vdd.n1493 9.3005
R19210 vdd.n1466 vdd.n1463 9.3005
R19211 vdd.n1501 vdd.n1500 9.3005
R19212 vdd.n1529 vdd.n1528 9.3005
R19213 vdd.n1524 vdd.n1523 9.3005
R19214 vdd.n1535 vdd.n1534 9.3005
R19215 vdd.n1537 vdd.n1536 9.3005
R19216 vdd.n1520 vdd.n1519 9.3005
R19217 vdd.n1543 vdd.n1542 9.3005
R19218 vdd.n1545 vdd.n1544 9.3005
R19219 vdd.n1517 vdd.n1514 9.3005
R19220 vdd.n1552 vdd.n1551 9.3005
R19221 vdd.n1384 vdd.n1383 9.3005
R19222 vdd.n1379 vdd.n1378 9.3005
R19223 vdd.n1390 vdd.n1389 9.3005
R19224 vdd.n1392 vdd.n1391 9.3005
R19225 vdd.n1375 vdd.n1374 9.3005
R19226 vdd.n1398 vdd.n1397 9.3005
R19227 vdd.n1400 vdd.n1399 9.3005
R19228 vdd.n1372 vdd.n1369 9.3005
R19229 vdd.n1407 vdd.n1406 9.3005
R19230 vdd.n1435 vdd.n1434 9.3005
R19231 vdd.n1430 vdd.n1429 9.3005
R19232 vdd.n1441 vdd.n1440 9.3005
R19233 vdd.n1443 vdd.n1442 9.3005
R19234 vdd.n1426 vdd.n1425 9.3005
R19235 vdd.n1449 vdd.n1448 9.3005
R19236 vdd.n1451 vdd.n1450 9.3005
R19237 vdd.n1423 vdd.n1420 9.3005
R19238 vdd.n1458 vdd.n1457 9.3005
R19239 vdd.n1291 vdd.n1290 9.3005
R19240 vdd.n1286 vdd.n1285 9.3005
R19241 vdd.n1297 vdd.n1296 9.3005
R19242 vdd.n1299 vdd.n1298 9.3005
R19243 vdd.n1282 vdd.n1281 9.3005
R19244 vdd.n1305 vdd.n1304 9.3005
R19245 vdd.n1307 vdd.n1306 9.3005
R19246 vdd.n1279 vdd.n1276 9.3005
R19247 vdd.n1314 vdd.n1313 9.3005
R19248 vdd.n1342 vdd.n1341 9.3005
R19249 vdd.n1337 vdd.n1336 9.3005
R19250 vdd.n1348 vdd.n1347 9.3005
R19251 vdd.n1350 vdd.n1349 9.3005
R19252 vdd.n1333 vdd.n1332 9.3005
R19253 vdd.n1356 vdd.n1355 9.3005
R19254 vdd.n1358 vdd.n1357 9.3005
R19255 vdd.n1330 vdd.n1327 9.3005
R19256 vdd.n1365 vdd.n1364 9.3005
R19257 vdd.n288 vdd.n287 8.92171
R19258 vdd.n237 vdd.n236 8.92171
R19259 vdd.n194 vdd.n193 8.92171
R19260 vdd.n143 vdd.n142 8.92171
R19261 vdd.n101 vdd.n100 8.92171
R19262 vdd.n50 vdd.n49 8.92171
R19263 vdd.n1483 vdd.n1482 8.92171
R19264 vdd.n1534 vdd.n1533 8.92171
R19265 vdd.n1389 vdd.n1388 8.92171
R19266 vdd.n1440 vdd.n1439 8.92171
R19267 vdd.n1296 vdd.n1295 8.92171
R19268 vdd.n1347 vdd.n1346 8.92171
R19269 vdd.n215 vdd.n121 8.81535
R19270 vdd.n1461 vdd.n1367 8.81535
R19271 vdd.n1596 vdd.t17 8.72962
R19272 vdd.n2956 vdd.t15 8.72962
R19273 vdd.t21 vdd.n1570 8.50289
R19274 vdd.n493 vdd.t6 8.50289
R19275 vdd.n28 vdd.n14 8.42249
R19276 vdd.n1272 vdd.t162 8.27616
R19277 vdd.n3164 vdd.t60 8.27616
R19278 vdd.n3168 vdd.n3167 8.16225
R19279 vdd.n1557 vdd.n1556 8.16225
R19280 vdd.n284 vdd.n278 8.14595
R19281 vdd.n233 vdd.n227 8.14595
R19282 vdd.n190 vdd.n184 8.14595
R19283 vdd.n139 vdd.n133 8.14595
R19284 vdd.n97 vdd.n91 8.14595
R19285 vdd.n46 vdd.n40 8.14595
R19286 vdd.n1479 vdd.n1473 8.14595
R19287 vdd.n1530 vdd.n1524 8.14595
R19288 vdd.n1385 vdd.n1379 8.14595
R19289 vdd.n1436 vdd.n1430 8.14595
R19290 vdd.n1292 vdd.n1286 8.14595
R19291 vdd.n1343 vdd.n1337 8.14595
R19292 vdd.n2635 vdd.n677 8.11757
R19293 vdd.n2109 vdd.n2108 8.11757
R19294 vdd.t36 vdd.n960 8.04943
R19295 vdd.n3155 vdd.t34 8.04943
R19296 vdd.n2087 vdd.n871 7.70933
R19297 vdd.n2093 vdd.n871 7.70933
R19298 vdd.n2099 vdd.n865 7.70933
R19299 vdd.n2099 vdd.n858 7.70933
R19300 vdd.n2105 vdd.n858 7.70933
R19301 vdd.n2105 vdd.n861 7.70933
R19302 vdd.n2112 vdd.n846 7.70933
R19303 vdd.n2118 vdd.n846 7.70933
R19304 vdd.n2124 vdd.n840 7.70933
R19305 vdd.n2130 vdd.n836 7.70933
R19306 vdd.n2136 vdd.n830 7.70933
R19307 vdd.n2148 vdd.n817 7.70933
R19308 vdd.n2154 vdd.n811 7.70933
R19309 vdd.n2154 vdd.n804 7.70933
R19310 vdd.n2162 vdd.n804 7.70933
R19311 vdd.n2169 vdd.t159 7.70933
R19312 vdd.n2244 vdd.t159 7.70933
R19313 vdd.n2576 vdd.t66 7.70933
R19314 vdd.n2582 vdd.t66 7.70933
R19315 vdd.n2588 vdd.n725 7.70933
R19316 vdd.n2594 vdd.n725 7.70933
R19317 vdd.n2594 vdd.n728 7.70933
R19318 vdd.n2600 vdd.n721 7.70933
R19319 vdd.n2612 vdd.n708 7.70933
R19320 vdd.n2618 vdd.n702 7.70933
R19321 vdd.n2624 vdd.n698 7.70933
R19322 vdd.n2630 vdd.n685 7.70933
R19323 vdd.n2638 vdd.n685 7.70933
R19324 vdd.n2644 vdd.n679 7.70933
R19325 vdd.n2644 vdd.n671 7.70933
R19326 vdd.n2695 vdd.n671 7.70933
R19327 vdd.n2695 vdd.n674 7.70933
R19328 vdd.n2701 vdd.n631 7.70933
R19329 vdd.n2771 vdd.n631 7.70933
R19330 vdd.n283 vdd.n280 7.3702
R19331 vdd.n232 vdd.n229 7.3702
R19332 vdd.n189 vdd.n186 7.3702
R19333 vdd.n138 vdd.n135 7.3702
R19334 vdd.n96 vdd.n93 7.3702
R19335 vdd.n45 vdd.n42 7.3702
R19336 vdd.n1478 vdd.n1475 7.3702
R19337 vdd.n1529 vdd.n1526 7.3702
R19338 vdd.n1384 vdd.n1381 7.3702
R19339 vdd.n1435 vdd.n1432 7.3702
R19340 vdd.n1291 vdd.n1288 7.3702
R19341 vdd.n1342 vdd.n1339 7.3702
R19342 vdd.n1239 vdd.t186 7.1425
R19343 vdd.n3148 vdd.t12 7.1425
R19344 vdd.n1150 vdd.n1149 6.98232
R19345 vdd.n1751 vdd.n1750 6.98232
R19346 vdd.n3063 vdd.n3062 6.98232
R19347 vdd.n2855 vdd.n2854 6.98232
R19348 vdd.n1255 vdd.t26 6.91577
R19349 vdd.n325 vdd.t164 6.91577
R19350 vdd.n1562 vdd.t46 6.68904
R19351 vdd.n2989 vdd.t32 6.68904
R19352 vdd.n925 vdd.t168 6.46231
R19353 vdd.t40 vdd.n492 6.46231
R19354 vdd.n3168 vdd.n309 6.27748
R19355 vdd.n1556 vdd.n1555 6.27748
R19356 vdd.n2124 vdd.t181 6.00885
R19357 vdd.n2624 vdd.t199 6.00885
R19358 vdd.n861 vdd.t124 5.89549
R19359 vdd.t92 vdd.n679 5.89549
R19360 vdd.n284 vdd.n283 5.81868
R19361 vdd.n233 vdd.n232 5.81868
R19362 vdd.n190 vdd.n189 5.81868
R19363 vdd.n139 vdd.n138 5.81868
R19364 vdd.n97 vdd.n96 5.81868
R19365 vdd.n46 vdd.n45 5.81868
R19366 vdd.n1479 vdd.n1478 5.81868
R19367 vdd.n1530 vdd.n1529 5.81868
R19368 vdd.n1385 vdd.n1384 5.81868
R19369 vdd.n1436 vdd.n1435 5.81868
R19370 vdd.n1292 vdd.n1291 5.81868
R19371 vdd.n1343 vdd.n1342 5.81868
R19372 vdd.t120 vdd.n865 5.78212
R19373 vdd.n1868 vdd.t105 5.78212
R19374 vdd.n2493 vdd.t113 5.78212
R19375 vdd.n674 vdd.t109 5.78212
R19376 vdd.n2252 vdd.n2251 5.77611
R19377 vdd.n1995 vdd.n1865 5.77611
R19378 vdd.n2506 vdd.n2505 5.77611
R19379 vdd.n2710 vdd.n663 5.77611
R19380 vdd.n2776 vdd.n627 5.77611
R19381 vdd.n2416 vdd.n2356 5.77611
R19382 vdd.n2177 vdd.n795 5.77611
R19383 vdd.n1925 vdd.n1924 5.77611
R19384 vdd.n1112 vdd.n1109 5.62474
R19385 vdd.n2047 vdd.n2044 5.62474
R19386 vdd.n3023 vdd.n3020 5.62474
R19387 vdd.n2810 vdd.n2807 5.62474
R19388 vdd.t28 vdd.n817 5.44203
R19389 vdd.n721 vdd.t226 5.44203
R19390 vdd.t68 vdd.n840 5.10193
R19391 vdd.n830 vdd.t71 5.10193
R19392 vdd.t59 vdd.n708 5.10193
R19393 vdd.n698 vdd.t45 5.10193
R19394 vdd.n287 vdd.n278 5.04292
R19395 vdd.n236 vdd.n227 5.04292
R19396 vdd.n193 vdd.n184 5.04292
R19397 vdd.n142 vdd.n133 5.04292
R19398 vdd.n100 vdd.n91 5.04292
R19399 vdd.n49 vdd.n40 5.04292
R19400 vdd.n1482 vdd.n1473 5.04292
R19401 vdd.n1533 vdd.n1524 5.04292
R19402 vdd.n1388 vdd.n1379 5.04292
R19403 vdd.n1439 vdd.n1430 5.04292
R19404 vdd.n1295 vdd.n1286 5.04292
R19405 vdd.n1346 vdd.n1337 5.04292
R19406 vdd.n1588 vdd.t168 4.8752
R19407 vdd.t0 vdd.t57 4.8752
R19408 vdd.t182 vdd.t43 4.8752
R19409 vdd.t55 vdd.t5 4.8752
R19410 vdd.t152 vdd.t158 4.8752
R19411 vdd.n2964 vdd.t40 4.8752
R19412 vdd.n2253 vdd.n2252 4.83952
R19413 vdd.n1865 vdd.n1861 4.83952
R19414 vdd.n2507 vdd.n2506 4.83952
R19415 vdd.n663 vdd.n658 4.83952
R19416 vdd.n627 vdd.n622 4.83952
R19417 vdd.n2413 vdd.n2356 4.83952
R19418 vdd.n2180 vdd.n795 4.83952
R19419 vdd.n1924 vdd.n1923 4.83952
R19420 vdd.n1719 vdd.n893 4.74817
R19421 vdd.n1714 vdd.n894 4.74817
R19422 vdd.n1616 vdd.n1613 4.74817
R19423 vdd.n2028 vdd.n1617 4.74817
R19424 vdd.n2030 vdd.n1616 4.74817
R19425 vdd.n2029 vdd.n2028 4.74817
R19426 vdd.n521 vdd.n519 4.74817
R19427 vdd.n2925 vdd.n522 4.74817
R19428 vdd.n2928 vdd.n522 4.74817
R19429 vdd.n2929 vdd.n521 4.74817
R19430 vdd.n2817 vdd.n606 4.74817
R19431 vdd.n2813 vdd.n608 4.74817
R19432 vdd.n2816 vdd.n608 4.74817
R19433 vdd.n2821 vdd.n606 4.74817
R19434 vdd.n1715 vdd.n893 4.74817
R19435 vdd.n896 vdd.n894 4.74817
R19436 vdd.n309 vdd.n308 4.7074
R19437 vdd.n215 vdd.n214 4.7074
R19438 vdd.n1555 vdd.n1554 4.7074
R19439 vdd.n1461 vdd.n1460 4.7074
R19440 vdd.t46 vdd.n931 4.64847
R19441 vdd.n2980 vdd.t32 4.64847
R19442 vdd.n2130 vdd.t1 4.53511
R19443 vdd.n2618 vdd.t3 4.53511
R19444 vdd.n1264 vdd.t26 4.42174
R19445 vdd.n3162 vdd.t164 4.42174
R19446 vdd.n2162 vdd.t197 4.30838
R19447 vdd.n2588 vdd.t69 4.30838
R19448 vdd.n288 vdd.n276 4.26717
R19449 vdd.n237 vdd.n225 4.26717
R19450 vdd.n194 vdd.n182 4.26717
R19451 vdd.n143 vdd.n131 4.26717
R19452 vdd.n101 vdd.n89 4.26717
R19453 vdd.n50 vdd.n38 4.26717
R19454 vdd.n1483 vdd.n1471 4.26717
R19455 vdd.n1534 vdd.n1522 4.26717
R19456 vdd.n1389 vdd.n1377 4.26717
R19457 vdd.n1440 vdd.n1428 4.26717
R19458 vdd.n1296 vdd.n1284 4.26717
R19459 vdd.n1347 vdd.n1335 4.26717
R19460 vdd.t186 vdd.n959 4.19501
R19461 vdd.t12 vdd.n329 4.19501
R19462 vdd.n309 vdd.n215 4.10845
R19463 vdd.n1555 vdd.n1461 4.10845
R19464 vdd.n265 vdd.t173 4.06363
R19465 vdd.n265 vdd.t64 4.06363
R19466 vdd.n263 vdd.t165 4.06363
R19467 vdd.n263 vdd.t161 4.06363
R19468 vdd.n261 vdd.t203 4.06363
R19469 vdd.n261 vdd.t61 4.06363
R19470 vdd.n259 vdd.t183 4.06363
R19471 vdd.n259 vdd.t49 4.06363
R19472 vdd.n257 vdd.t41 4.06363
R19473 vdd.n257 vdd.t53 4.06363
R19474 vdd.n171 vdd.t167 4.06363
R19475 vdd.n171 vdd.t13 4.06363
R19476 vdd.n169 vdd.t229 4.06363
R19477 vdd.n169 vdd.t228 4.06363
R19478 vdd.n167 vdd.t192 4.06363
R19479 vdd.n167 vdd.t174 4.06363
R19480 vdd.n165 vdd.t7 4.06363
R19481 vdd.n165 vdd.t33 4.06363
R19482 vdd.n163 vdd.t231 4.06363
R19483 vdd.n163 vdd.t190 4.06363
R19484 vdd.n78 vdd.t35 4.06363
R19485 vdd.n78 vdd.t185 4.06363
R19486 vdd.n76 vdd.t170 4.06363
R19487 vdd.n76 vdd.t20 4.06363
R19488 vdd.n74 vdd.t202 4.06363
R19489 vdd.n74 vdd.t166 4.06363
R19490 vdd.n72 vdd.t172 4.06363
R19491 vdd.n72 vdd.t180 4.06363
R19492 vdd.n70 vdd.t176 4.06363
R19493 vdd.n70 vdd.t73 4.06363
R19494 vdd.n1503 vdd.t48 4.06363
R19495 vdd.n1503 vdd.t209 4.06363
R19496 vdd.n1505 vdd.t195 4.06363
R19497 vdd.n1505 vdd.t25 4.06363
R19498 vdd.n1507 vdd.t230 4.06363
R19499 vdd.n1507 vdd.t184 4.06363
R19500 vdd.n1509 vdd.t175 4.06363
R19501 vdd.n1509 vdd.t27 4.06363
R19502 vdd.n1511 vdd.t201 4.06363
R19503 vdd.n1511 vdd.t65 4.06363
R19504 vdd.n1409 vdd.t39 4.06363
R19505 vdd.n1409 vdd.t177 4.06363
R19506 vdd.n1411 vdd.t194 4.06363
R19507 vdd.n1411 vdd.t74 4.06363
R19508 vdd.n1413 vdd.t163 4.06363
R19509 vdd.n1413 vdd.t9 4.06363
R19510 vdd.n1415 vdd.t196 4.06363
R19511 vdd.n1415 vdd.t75 4.06363
R19512 vdd.n1417 vdd.t189 4.06363
R19513 vdd.n1417 vdd.t179 4.06363
R19514 vdd.n1316 vdd.t31 4.06363
R19515 vdd.n1316 vdd.t169 4.06363
R19516 vdd.n1318 vdd.t47 4.06363
R19517 vdd.n1318 vdd.t22 4.06363
R19518 vdd.n1320 vdd.t206 4.06363
R19519 vdd.n1320 vdd.t193 4.06363
R19520 vdd.n1322 vdd.t51 4.06363
R19521 vdd.n1322 vdd.t171 4.06363
R19522 vdd.n1324 vdd.t187 4.06363
R19523 vdd.n1324 vdd.t37 4.06363
R19524 vdd.n26 vdd.t221 3.9605
R19525 vdd.n26 vdd.t220 3.9605
R19526 vdd.n23 vdd.t214 3.9605
R19527 vdd.n23 vdd.t213 3.9605
R19528 vdd.n21 vdd.t218 3.9605
R19529 vdd.n21 vdd.t222 3.9605
R19530 vdd.n20 vdd.t210 3.9605
R19531 vdd.n20 vdd.t212 3.9605
R19532 vdd.n15 vdd.t215 3.9605
R19533 vdd.n15 vdd.t223 3.9605
R19534 vdd.n16 vdd.t217 3.9605
R19535 vdd.n16 vdd.t211 3.9605
R19536 vdd.n18 vdd.t225 3.9605
R19537 vdd.n18 vdd.t219 3.9605
R19538 vdd.n25 vdd.t216 3.9605
R19539 vdd.n25 vdd.t224 3.9605
R19540 vdd.n7 vdd.t153 3.61217
R19541 vdd.n7 vdd.t4 3.61217
R19542 vdd.n8 vdd.t56 3.61217
R19543 vdd.n8 vdd.t227 3.61217
R19544 vdd.n10 vdd.t67 3.61217
R19545 vdd.n10 vdd.t70 3.61217
R19546 vdd.n12 vdd.t157 3.61217
R19547 vdd.n12 vdd.t24 3.61217
R19548 vdd.n5 vdd.t155 3.61217
R19549 vdd.n5 vdd.t205 3.61217
R19550 vdd.n3 vdd.t198 3.61217
R19551 vdd.n3 vdd.t160 3.61217
R19552 vdd.n1 vdd.t29 3.61217
R19553 vdd.n1 vdd.t44 3.61217
R19554 vdd.n0 vdd.t2 3.61217
R19555 vdd.n0 vdd.t58 3.61217
R19556 vdd.n292 vdd.n291 3.49141
R19557 vdd.n241 vdd.n240 3.49141
R19558 vdd.n198 vdd.n197 3.49141
R19559 vdd.n147 vdd.n146 3.49141
R19560 vdd.n105 vdd.n104 3.49141
R19561 vdd.n54 vdd.n53 3.49141
R19562 vdd.n1487 vdd.n1486 3.49141
R19563 vdd.n1538 vdd.n1537 3.49141
R19564 vdd.n1393 vdd.n1392 3.49141
R19565 vdd.n1444 vdd.n1443 3.49141
R19566 vdd.n1300 vdd.n1299 3.49141
R19567 vdd.n1351 vdd.n1350 3.49141
R19568 vdd.n1868 vdd.t197 3.40145
R19569 vdd.n2316 vdd.t154 3.40145
R19570 vdd.n2569 vdd.t23 3.40145
R19571 vdd.n2493 vdd.t69 3.40145
R19572 vdd.n1247 vdd.t36 3.28809
R19573 vdd.t34 vdd.n3154 3.28809
R19574 vdd.n1969 vdd.t1 3.17472
R19575 vdd.n2472 vdd.t3 3.17472
R19576 vdd.n948 vdd.t162 3.06136
R19577 vdd.t60 vdd.n3163 3.06136
R19578 vdd.n1571 vdd.t21 2.83463
R19579 vdd.n2981 vdd.t6 2.83463
R19580 vdd.n295 vdd.n274 2.71565
R19581 vdd.n244 vdd.n223 2.71565
R19582 vdd.n201 vdd.n180 2.71565
R19583 vdd.n150 vdd.n129 2.71565
R19584 vdd.n108 vdd.n87 2.71565
R19585 vdd.n57 vdd.n36 2.71565
R19586 vdd.n1490 vdd.n1469 2.71565
R19587 vdd.n1541 vdd.n1520 2.71565
R19588 vdd.n1396 vdd.n1375 2.71565
R19589 vdd.n1447 vdd.n1426 2.71565
R19590 vdd.n1303 vdd.n1282 2.71565
R19591 vdd.n1354 vdd.n1333 2.71565
R19592 vdd.n1587 vdd.t17 2.6079
R19593 vdd.n2118 vdd.t68 2.6079
R19594 vdd.n2142 vdd.t71 2.6079
R19595 vdd.n2606 vdd.t59 2.6079
R19596 vdd.n2630 vdd.t45 2.6079
R19597 vdd.t15 vdd.n499 2.6079
R19598 vdd.n2636 vdd.n2635 2.49806
R19599 vdd.n2110 vdd.n2109 2.49806
R19600 vdd.n282 vdd.n281 2.4129
R19601 vdd.n231 vdd.n230 2.4129
R19602 vdd.n188 vdd.n187 2.4129
R19603 vdd.n137 vdd.n136 2.4129
R19604 vdd.n95 vdd.n94 2.4129
R19605 vdd.n44 vdd.n43 2.4129
R19606 vdd.n1477 vdd.n1476 2.4129
R19607 vdd.n1528 vdd.n1527 2.4129
R19608 vdd.n1383 vdd.n1382 2.4129
R19609 vdd.n1434 vdd.n1433 2.4129
R19610 vdd.n1290 vdd.n1289 2.4129
R19611 vdd.n1341 vdd.n1340 2.4129
R19612 vdd.n2027 vdd.n1616 2.27742
R19613 vdd.n2028 vdd.n2027 2.27742
R19614 vdd.n2737 vdd.n522 2.27742
R19615 vdd.n2737 vdd.n521 2.27742
R19616 vdd.n2805 vdd.n608 2.27742
R19617 vdd.n2805 vdd.n606 2.27742
R19618 vdd.n2050 vdd.n893 2.27742
R19619 vdd.n2050 vdd.n894 2.27742
R19620 vdd.n2142 vdd.t28 2.2678
R19621 vdd.n2606 vdd.t226 2.2678
R19622 vdd.t43 vdd.n811 2.04107
R19623 vdd.n728 vdd.t55 2.04107
R19624 vdd.n296 vdd.n272 1.93989
R19625 vdd.n245 vdd.n221 1.93989
R19626 vdd.n202 vdd.n178 1.93989
R19627 vdd.n151 vdd.n127 1.93989
R19628 vdd.n109 vdd.n85 1.93989
R19629 vdd.n58 vdd.n34 1.93989
R19630 vdd.n1491 vdd.n1467 1.93989
R19631 vdd.n1542 vdd.n1518 1.93989
R19632 vdd.n1397 vdd.n1373 1.93989
R19633 vdd.n1448 vdd.n1424 1.93989
R19634 vdd.n1304 vdd.n1280 1.93989
R19635 vdd.n1355 vdd.n1331 1.93989
R19636 vdd.n2093 vdd.t120 1.92771
R19637 vdd.n2169 vdd.t105 1.92771
R19638 vdd.n2582 vdd.t113 1.92771
R19639 vdd.n2701 vdd.t109 1.92771
R19640 vdd.n1969 vdd.t181 1.70098
R19641 vdd.n836 vdd.t0 1.70098
R19642 vdd.t158 vdd.n702 1.70098
R19643 vdd.n2472 vdd.t199 1.70098
R19644 vdd.n983 vdd.t88 1.47425
R19645 vdd.t137 vdd.n3139 1.47425
R19646 vdd.n307 vdd.n267 1.16414
R19647 vdd.n300 vdd.n299 1.16414
R19648 vdd.n256 vdd.n216 1.16414
R19649 vdd.n249 vdd.n248 1.16414
R19650 vdd.n213 vdd.n173 1.16414
R19651 vdd.n206 vdd.n205 1.16414
R19652 vdd.n162 vdd.n122 1.16414
R19653 vdd.n155 vdd.n154 1.16414
R19654 vdd.n120 vdd.n80 1.16414
R19655 vdd.n113 vdd.n112 1.16414
R19656 vdd.n69 vdd.n29 1.16414
R19657 vdd.n62 vdd.n61 1.16414
R19658 vdd.n1502 vdd.n1462 1.16414
R19659 vdd.n1495 vdd.n1494 1.16414
R19660 vdd.n1553 vdd.n1513 1.16414
R19661 vdd.n1546 vdd.n1545 1.16414
R19662 vdd.n1408 vdd.n1368 1.16414
R19663 vdd.n1401 vdd.n1400 1.16414
R19664 vdd.n1459 vdd.n1419 1.16414
R19665 vdd.n1452 vdd.n1451 1.16414
R19666 vdd.n1315 vdd.n1275 1.16414
R19667 vdd.n1308 vdd.n1307 1.16414
R19668 vdd.n1366 vdd.n1326 1.16414
R19669 vdd.n1359 vdd.n1358 1.16414
R19670 vdd.n2136 vdd.t57 1.13415
R19671 vdd.n2612 vdd.t152 1.13415
R19672 vdd.n1579 vdd.t30 1.02079
R19673 vdd.t124 vdd.t14 1.02079
R19674 vdd.t178 vdd.t92 1.02079
R19675 vdd.n2972 vdd.t52 1.02079
R19676 vdd.n1113 vdd.n1112 0.970197
R19677 vdd.n2048 vdd.n2047 0.970197
R19678 vdd.n3024 vdd.n3023 0.970197
R19679 vdd.n2812 vdd.n2810 0.970197
R19680 vdd.n1556 vdd.n28 0.800283
R19681 vdd.t8 vdd.n937 0.794056
R19682 vdd.n1606 vdd.t84 0.794056
R19683 vdd.n2112 vdd.t14 0.794056
R19684 vdd.n2148 vdd.t182 0.794056
R19685 vdd.n2600 vdd.t5 0.794056
R19686 vdd.n2638 vdd.t178 0.794056
R19687 vdd.t77 vdd.n511 0.794056
R19688 vdd.n481 vdd.t191 0.794056
R19689 vdd vdd.n3168 0.79245
R19690 vdd.n1256 vdd.t50 0.567326
R19691 vdd.n3156 vdd.t19 0.567326
R19692 vdd.n2038 vdd.n2037 0.509646
R19693 vdd.n2937 vdd.n2936 0.509646
R19694 vdd.n3135 vdd.n3134 0.509646
R19695 vdd.n3017 vdd.n3016 0.509646
R19696 vdd.n2943 vdd.n514 0.509646
R19697 vdd.n1601 vdd.n895 0.509646
R19698 vdd.n1218 vdd.n980 0.509646
R19699 vdd.n1212 vdd.n1211 0.509646
R19700 vdd.n4 vdd.n2 0.459552
R19701 vdd.n11 vdd.n9 0.459552
R19702 vdd.n305 vdd.n304 0.388379
R19703 vdd.n271 vdd.n269 0.388379
R19704 vdd.n254 vdd.n253 0.388379
R19705 vdd.n220 vdd.n218 0.388379
R19706 vdd.n211 vdd.n210 0.388379
R19707 vdd.n177 vdd.n175 0.388379
R19708 vdd.n160 vdd.n159 0.388379
R19709 vdd.n126 vdd.n124 0.388379
R19710 vdd.n118 vdd.n117 0.388379
R19711 vdd.n84 vdd.n82 0.388379
R19712 vdd.n67 vdd.n66 0.388379
R19713 vdd.n33 vdd.n31 0.388379
R19714 vdd.n1500 vdd.n1499 0.388379
R19715 vdd.n1466 vdd.n1464 0.388379
R19716 vdd.n1551 vdd.n1550 0.388379
R19717 vdd.n1517 vdd.n1515 0.388379
R19718 vdd.n1406 vdd.n1405 0.388379
R19719 vdd.n1372 vdd.n1370 0.388379
R19720 vdd.n1457 vdd.n1456 0.388379
R19721 vdd.n1423 vdd.n1421 0.388379
R19722 vdd.n1313 vdd.n1312 0.388379
R19723 vdd.n1279 vdd.n1277 0.388379
R19724 vdd.n1364 vdd.n1363 0.388379
R19725 vdd.n1330 vdd.n1328 0.388379
R19726 vdd.n19 vdd.n17 0.387128
R19727 vdd.n24 vdd.n22 0.387128
R19728 vdd.n6 vdd.n4 0.358259
R19729 vdd.n13 vdd.n11 0.358259
R19730 vdd.n260 vdd.n258 0.358259
R19731 vdd.n262 vdd.n260 0.358259
R19732 vdd.n264 vdd.n262 0.358259
R19733 vdd.n266 vdd.n264 0.358259
R19734 vdd.n308 vdd.n266 0.358259
R19735 vdd.n166 vdd.n164 0.358259
R19736 vdd.n168 vdd.n166 0.358259
R19737 vdd.n170 vdd.n168 0.358259
R19738 vdd.n172 vdd.n170 0.358259
R19739 vdd.n214 vdd.n172 0.358259
R19740 vdd.n73 vdd.n71 0.358259
R19741 vdd.n75 vdd.n73 0.358259
R19742 vdd.n77 vdd.n75 0.358259
R19743 vdd.n79 vdd.n77 0.358259
R19744 vdd.n121 vdd.n79 0.358259
R19745 vdd.n1554 vdd.n1512 0.358259
R19746 vdd.n1512 vdd.n1510 0.358259
R19747 vdd.n1510 vdd.n1508 0.358259
R19748 vdd.n1508 vdd.n1506 0.358259
R19749 vdd.n1506 vdd.n1504 0.358259
R19750 vdd.n1460 vdd.n1418 0.358259
R19751 vdd.n1418 vdd.n1416 0.358259
R19752 vdd.n1416 vdd.n1414 0.358259
R19753 vdd.n1414 vdd.n1412 0.358259
R19754 vdd.n1412 vdd.n1410 0.358259
R19755 vdd.n1367 vdd.n1325 0.358259
R19756 vdd.n1325 vdd.n1323 0.358259
R19757 vdd.n1323 vdd.n1321 0.358259
R19758 vdd.n1321 vdd.n1319 0.358259
R19759 vdd.n1319 vdd.n1317 0.358259
R19760 vdd.t62 vdd.n966 0.340595
R19761 vdd.n3147 vdd.t10 0.340595
R19762 vdd.n14 vdd.n6 0.334552
R19763 vdd.n14 vdd.n13 0.334552
R19764 vdd.n27 vdd.n19 0.21707
R19765 vdd.n27 vdd.n24 0.21707
R19766 vdd.n306 vdd.n268 0.155672
R19767 vdd.n298 vdd.n268 0.155672
R19768 vdd.n298 vdd.n297 0.155672
R19769 vdd.n297 vdd.n273 0.155672
R19770 vdd.n290 vdd.n273 0.155672
R19771 vdd.n290 vdd.n289 0.155672
R19772 vdd.n289 vdd.n277 0.155672
R19773 vdd.n282 vdd.n277 0.155672
R19774 vdd.n255 vdd.n217 0.155672
R19775 vdd.n247 vdd.n217 0.155672
R19776 vdd.n247 vdd.n246 0.155672
R19777 vdd.n246 vdd.n222 0.155672
R19778 vdd.n239 vdd.n222 0.155672
R19779 vdd.n239 vdd.n238 0.155672
R19780 vdd.n238 vdd.n226 0.155672
R19781 vdd.n231 vdd.n226 0.155672
R19782 vdd.n212 vdd.n174 0.155672
R19783 vdd.n204 vdd.n174 0.155672
R19784 vdd.n204 vdd.n203 0.155672
R19785 vdd.n203 vdd.n179 0.155672
R19786 vdd.n196 vdd.n179 0.155672
R19787 vdd.n196 vdd.n195 0.155672
R19788 vdd.n195 vdd.n183 0.155672
R19789 vdd.n188 vdd.n183 0.155672
R19790 vdd.n161 vdd.n123 0.155672
R19791 vdd.n153 vdd.n123 0.155672
R19792 vdd.n153 vdd.n152 0.155672
R19793 vdd.n152 vdd.n128 0.155672
R19794 vdd.n145 vdd.n128 0.155672
R19795 vdd.n145 vdd.n144 0.155672
R19796 vdd.n144 vdd.n132 0.155672
R19797 vdd.n137 vdd.n132 0.155672
R19798 vdd.n119 vdd.n81 0.155672
R19799 vdd.n111 vdd.n81 0.155672
R19800 vdd.n111 vdd.n110 0.155672
R19801 vdd.n110 vdd.n86 0.155672
R19802 vdd.n103 vdd.n86 0.155672
R19803 vdd.n103 vdd.n102 0.155672
R19804 vdd.n102 vdd.n90 0.155672
R19805 vdd.n95 vdd.n90 0.155672
R19806 vdd.n68 vdd.n30 0.155672
R19807 vdd.n60 vdd.n30 0.155672
R19808 vdd.n60 vdd.n59 0.155672
R19809 vdd.n59 vdd.n35 0.155672
R19810 vdd.n52 vdd.n35 0.155672
R19811 vdd.n52 vdd.n51 0.155672
R19812 vdd.n51 vdd.n39 0.155672
R19813 vdd.n44 vdd.n39 0.155672
R19814 vdd.n1501 vdd.n1463 0.155672
R19815 vdd.n1493 vdd.n1463 0.155672
R19816 vdd.n1493 vdd.n1492 0.155672
R19817 vdd.n1492 vdd.n1468 0.155672
R19818 vdd.n1485 vdd.n1468 0.155672
R19819 vdd.n1485 vdd.n1484 0.155672
R19820 vdd.n1484 vdd.n1472 0.155672
R19821 vdd.n1477 vdd.n1472 0.155672
R19822 vdd.n1552 vdd.n1514 0.155672
R19823 vdd.n1544 vdd.n1514 0.155672
R19824 vdd.n1544 vdd.n1543 0.155672
R19825 vdd.n1543 vdd.n1519 0.155672
R19826 vdd.n1536 vdd.n1519 0.155672
R19827 vdd.n1536 vdd.n1535 0.155672
R19828 vdd.n1535 vdd.n1523 0.155672
R19829 vdd.n1528 vdd.n1523 0.155672
R19830 vdd.n1407 vdd.n1369 0.155672
R19831 vdd.n1399 vdd.n1369 0.155672
R19832 vdd.n1399 vdd.n1398 0.155672
R19833 vdd.n1398 vdd.n1374 0.155672
R19834 vdd.n1391 vdd.n1374 0.155672
R19835 vdd.n1391 vdd.n1390 0.155672
R19836 vdd.n1390 vdd.n1378 0.155672
R19837 vdd.n1383 vdd.n1378 0.155672
R19838 vdd.n1458 vdd.n1420 0.155672
R19839 vdd.n1450 vdd.n1420 0.155672
R19840 vdd.n1450 vdd.n1449 0.155672
R19841 vdd.n1449 vdd.n1425 0.155672
R19842 vdd.n1442 vdd.n1425 0.155672
R19843 vdd.n1442 vdd.n1441 0.155672
R19844 vdd.n1441 vdd.n1429 0.155672
R19845 vdd.n1434 vdd.n1429 0.155672
R19846 vdd.n1314 vdd.n1276 0.155672
R19847 vdd.n1306 vdd.n1276 0.155672
R19848 vdd.n1306 vdd.n1305 0.155672
R19849 vdd.n1305 vdd.n1281 0.155672
R19850 vdd.n1298 vdd.n1281 0.155672
R19851 vdd.n1298 vdd.n1297 0.155672
R19852 vdd.n1297 vdd.n1285 0.155672
R19853 vdd.n1290 vdd.n1285 0.155672
R19854 vdd.n1365 vdd.n1327 0.155672
R19855 vdd.n1357 vdd.n1327 0.155672
R19856 vdd.n1357 vdd.n1356 0.155672
R19857 vdd.n1356 vdd.n1332 0.155672
R19858 vdd.n1349 vdd.n1332 0.155672
R19859 vdd.n1349 vdd.n1348 0.155672
R19860 vdd.n1348 vdd.n1336 0.155672
R19861 vdd.n1341 vdd.n1336 0.155672
R19862 vdd.n1813 vdd.n1618 0.152939
R19863 vdd.n1624 vdd.n1618 0.152939
R19864 vdd.n1625 vdd.n1624 0.152939
R19865 vdd.n1626 vdd.n1625 0.152939
R19866 vdd.n1627 vdd.n1626 0.152939
R19867 vdd.n1631 vdd.n1627 0.152939
R19868 vdd.n1632 vdd.n1631 0.152939
R19869 vdd.n1633 vdd.n1632 0.152939
R19870 vdd.n1634 vdd.n1633 0.152939
R19871 vdd.n1638 vdd.n1634 0.152939
R19872 vdd.n1639 vdd.n1638 0.152939
R19873 vdd.n1640 vdd.n1639 0.152939
R19874 vdd.n1788 vdd.n1640 0.152939
R19875 vdd.n1788 vdd.n1787 0.152939
R19876 vdd.n1787 vdd.n1786 0.152939
R19877 vdd.n1786 vdd.n1646 0.152939
R19878 vdd.n1651 vdd.n1646 0.152939
R19879 vdd.n1652 vdd.n1651 0.152939
R19880 vdd.n1653 vdd.n1652 0.152939
R19881 vdd.n1657 vdd.n1653 0.152939
R19882 vdd.n1658 vdd.n1657 0.152939
R19883 vdd.n1659 vdd.n1658 0.152939
R19884 vdd.n1660 vdd.n1659 0.152939
R19885 vdd.n1664 vdd.n1660 0.152939
R19886 vdd.n1665 vdd.n1664 0.152939
R19887 vdd.n1666 vdd.n1665 0.152939
R19888 vdd.n1667 vdd.n1666 0.152939
R19889 vdd.n1671 vdd.n1667 0.152939
R19890 vdd.n1672 vdd.n1671 0.152939
R19891 vdd.n1673 vdd.n1672 0.152939
R19892 vdd.n1674 vdd.n1673 0.152939
R19893 vdd.n1678 vdd.n1674 0.152939
R19894 vdd.n1679 vdd.n1678 0.152939
R19895 vdd.n1680 vdd.n1679 0.152939
R19896 vdd.n1749 vdd.n1680 0.152939
R19897 vdd.n1749 vdd.n1748 0.152939
R19898 vdd.n1748 vdd.n1747 0.152939
R19899 vdd.n1747 vdd.n1686 0.152939
R19900 vdd.n1691 vdd.n1686 0.152939
R19901 vdd.n1692 vdd.n1691 0.152939
R19902 vdd.n1693 vdd.n1692 0.152939
R19903 vdd.n1697 vdd.n1693 0.152939
R19904 vdd.n1698 vdd.n1697 0.152939
R19905 vdd.n1699 vdd.n1698 0.152939
R19906 vdd.n1700 vdd.n1699 0.152939
R19907 vdd.n1704 vdd.n1700 0.152939
R19908 vdd.n1705 vdd.n1704 0.152939
R19909 vdd.n1706 vdd.n1705 0.152939
R19910 vdd.n1707 vdd.n1706 0.152939
R19911 vdd.n1708 vdd.n1707 0.152939
R19912 vdd.n1708 vdd.n892 0.152939
R19913 vdd.n2037 vdd.n1612 0.152939
R19914 vdd.n1559 vdd.n1558 0.152939
R19915 vdd.n1559 vdd.n928 0.152939
R19916 vdd.n1574 vdd.n928 0.152939
R19917 vdd.n1575 vdd.n1574 0.152939
R19918 vdd.n1576 vdd.n1575 0.152939
R19919 vdd.n1576 vdd.n917 0.152939
R19920 vdd.n1591 vdd.n917 0.152939
R19921 vdd.n1592 vdd.n1591 0.152939
R19922 vdd.n1593 vdd.n1592 0.152939
R19923 vdd.n1593 vdd.n905 0.152939
R19924 vdd.n1610 vdd.n905 0.152939
R19925 vdd.n1611 vdd.n1610 0.152939
R19926 vdd.n2038 vdd.n1611 0.152939
R19927 vdd.n527 vdd.n524 0.152939
R19928 vdd.n528 vdd.n527 0.152939
R19929 vdd.n529 vdd.n528 0.152939
R19930 vdd.n530 vdd.n529 0.152939
R19931 vdd.n533 vdd.n530 0.152939
R19932 vdd.n534 vdd.n533 0.152939
R19933 vdd.n535 vdd.n534 0.152939
R19934 vdd.n536 vdd.n535 0.152939
R19935 vdd.n539 vdd.n536 0.152939
R19936 vdd.n540 vdd.n539 0.152939
R19937 vdd.n541 vdd.n540 0.152939
R19938 vdd.n542 vdd.n541 0.152939
R19939 vdd.n547 vdd.n542 0.152939
R19940 vdd.n548 vdd.n547 0.152939
R19941 vdd.n549 vdd.n548 0.152939
R19942 vdd.n550 vdd.n549 0.152939
R19943 vdd.n553 vdd.n550 0.152939
R19944 vdd.n554 vdd.n553 0.152939
R19945 vdd.n555 vdd.n554 0.152939
R19946 vdd.n556 vdd.n555 0.152939
R19947 vdd.n559 vdd.n556 0.152939
R19948 vdd.n560 vdd.n559 0.152939
R19949 vdd.n561 vdd.n560 0.152939
R19950 vdd.n562 vdd.n561 0.152939
R19951 vdd.n565 vdd.n562 0.152939
R19952 vdd.n566 vdd.n565 0.152939
R19953 vdd.n567 vdd.n566 0.152939
R19954 vdd.n568 vdd.n567 0.152939
R19955 vdd.n571 vdd.n568 0.152939
R19956 vdd.n572 vdd.n571 0.152939
R19957 vdd.n573 vdd.n572 0.152939
R19958 vdd.n574 vdd.n573 0.152939
R19959 vdd.n577 vdd.n574 0.152939
R19960 vdd.n578 vdd.n577 0.152939
R19961 vdd.n2853 vdd.n578 0.152939
R19962 vdd.n2853 vdd.n2852 0.152939
R19963 vdd.n2852 vdd.n2851 0.152939
R19964 vdd.n2851 vdd.n582 0.152939
R19965 vdd.n587 vdd.n582 0.152939
R19966 vdd.n588 vdd.n587 0.152939
R19967 vdd.n591 vdd.n588 0.152939
R19968 vdd.n592 vdd.n591 0.152939
R19969 vdd.n593 vdd.n592 0.152939
R19970 vdd.n594 vdd.n593 0.152939
R19971 vdd.n597 vdd.n594 0.152939
R19972 vdd.n598 vdd.n597 0.152939
R19973 vdd.n599 vdd.n598 0.152939
R19974 vdd.n600 vdd.n599 0.152939
R19975 vdd.n603 vdd.n600 0.152939
R19976 vdd.n604 vdd.n603 0.152939
R19977 vdd.n605 vdd.n604 0.152939
R19978 vdd.n2936 vdd.n518 0.152939
R19979 vdd.n2937 vdd.n508 0.152939
R19980 vdd.n2951 vdd.n508 0.152939
R19981 vdd.n2952 vdd.n2951 0.152939
R19982 vdd.n2953 vdd.n2952 0.152939
R19983 vdd.n2953 vdd.n496 0.152939
R19984 vdd.n2967 vdd.n496 0.152939
R19985 vdd.n2968 vdd.n2967 0.152939
R19986 vdd.n2969 vdd.n2968 0.152939
R19987 vdd.n2969 vdd.n484 0.152939
R19988 vdd.n2984 vdd.n484 0.152939
R19989 vdd.n2985 vdd.n2984 0.152939
R19990 vdd.n2986 vdd.n2985 0.152939
R19991 vdd.n2986 vdd.n310 0.152939
R19992 vdd.n320 vdd.n311 0.152939
R19993 vdd.n321 vdd.n320 0.152939
R19994 vdd.n322 vdd.n321 0.152939
R19995 vdd.n331 vdd.n322 0.152939
R19996 vdd.n332 vdd.n331 0.152939
R19997 vdd.n333 vdd.n332 0.152939
R19998 vdd.n334 vdd.n333 0.152939
R19999 vdd.n342 vdd.n334 0.152939
R20000 vdd.n343 vdd.n342 0.152939
R20001 vdd.n344 vdd.n343 0.152939
R20002 vdd.n345 vdd.n344 0.152939
R20003 vdd.n353 vdd.n345 0.152939
R20004 vdd.n3135 vdd.n353 0.152939
R20005 vdd.n3134 vdd.n354 0.152939
R20006 vdd.n357 vdd.n354 0.152939
R20007 vdd.n361 vdd.n357 0.152939
R20008 vdd.n362 vdd.n361 0.152939
R20009 vdd.n363 vdd.n362 0.152939
R20010 vdd.n364 vdd.n363 0.152939
R20011 vdd.n365 vdd.n364 0.152939
R20012 vdd.n369 vdd.n365 0.152939
R20013 vdd.n370 vdd.n369 0.152939
R20014 vdd.n371 vdd.n370 0.152939
R20015 vdd.n372 vdd.n371 0.152939
R20016 vdd.n376 vdd.n372 0.152939
R20017 vdd.n377 vdd.n376 0.152939
R20018 vdd.n378 vdd.n377 0.152939
R20019 vdd.n379 vdd.n378 0.152939
R20020 vdd.n383 vdd.n379 0.152939
R20021 vdd.n384 vdd.n383 0.152939
R20022 vdd.n385 vdd.n384 0.152939
R20023 vdd.n3100 vdd.n385 0.152939
R20024 vdd.n3100 vdd.n3099 0.152939
R20025 vdd.n3099 vdd.n3098 0.152939
R20026 vdd.n3098 vdd.n391 0.152939
R20027 vdd.n396 vdd.n391 0.152939
R20028 vdd.n397 vdd.n396 0.152939
R20029 vdd.n398 vdd.n397 0.152939
R20030 vdd.n402 vdd.n398 0.152939
R20031 vdd.n403 vdd.n402 0.152939
R20032 vdd.n404 vdd.n403 0.152939
R20033 vdd.n405 vdd.n404 0.152939
R20034 vdd.n409 vdd.n405 0.152939
R20035 vdd.n410 vdd.n409 0.152939
R20036 vdd.n411 vdd.n410 0.152939
R20037 vdd.n412 vdd.n411 0.152939
R20038 vdd.n416 vdd.n412 0.152939
R20039 vdd.n417 vdd.n416 0.152939
R20040 vdd.n418 vdd.n417 0.152939
R20041 vdd.n419 vdd.n418 0.152939
R20042 vdd.n423 vdd.n419 0.152939
R20043 vdd.n424 vdd.n423 0.152939
R20044 vdd.n425 vdd.n424 0.152939
R20045 vdd.n3061 vdd.n425 0.152939
R20046 vdd.n3061 vdd.n3060 0.152939
R20047 vdd.n3060 vdd.n3059 0.152939
R20048 vdd.n3059 vdd.n431 0.152939
R20049 vdd.n436 vdd.n431 0.152939
R20050 vdd.n437 vdd.n436 0.152939
R20051 vdd.n438 vdd.n437 0.152939
R20052 vdd.n442 vdd.n438 0.152939
R20053 vdd.n443 vdd.n442 0.152939
R20054 vdd.n444 vdd.n443 0.152939
R20055 vdd.n445 vdd.n444 0.152939
R20056 vdd.n449 vdd.n445 0.152939
R20057 vdd.n450 vdd.n449 0.152939
R20058 vdd.n451 vdd.n450 0.152939
R20059 vdd.n452 vdd.n451 0.152939
R20060 vdd.n456 vdd.n452 0.152939
R20061 vdd.n457 vdd.n456 0.152939
R20062 vdd.n458 vdd.n457 0.152939
R20063 vdd.n459 vdd.n458 0.152939
R20064 vdd.n463 vdd.n459 0.152939
R20065 vdd.n464 vdd.n463 0.152939
R20066 vdd.n465 vdd.n464 0.152939
R20067 vdd.n3017 vdd.n465 0.152939
R20068 vdd.n2944 vdd.n2943 0.152939
R20069 vdd.n2945 vdd.n2944 0.152939
R20070 vdd.n2945 vdd.n502 0.152939
R20071 vdd.n2959 vdd.n502 0.152939
R20072 vdd.n2960 vdd.n2959 0.152939
R20073 vdd.n2961 vdd.n2960 0.152939
R20074 vdd.n2961 vdd.n489 0.152939
R20075 vdd.n2975 vdd.n489 0.152939
R20076 vdd.n2976 vdd.n2975 0.152939
R20077 vdd.n2977 vdd.n2976 0.152939
R20078 vdd.n2977 vdd.n477 0.152939
R20079 vdd.n2992 vdd.n477 0.152939
R20080 vdd.n2993 vdd.n2992 0.152939
R20081 vdd.n2994 vdd.n2993 0.152939
R20082 vdd.n2994 vdd.n475 0.152939
R20083 vdd.n2998 vdd.n475 0.152939
R20084 vdd.n2999 vdd.n2998 0.152939
R20085 vdd.n3000 vdd.n2999 0.152939
R20086 vdd.n3000 vdd.n472 0.152939
R20087 vdd.n3004 vdd.n472 0.152939
R20088 vdd.n3005 vdd.n3004 0.152939
R20089 vdd.n3006 vdd.n3005 0.152939
R20090 vdd.n3006 vdd.n469 0.152939
R20091 vdd.n3010 vdd.n469 0.152939
R20092 vdd.n3011 vdd.n3010 0.152939
R20093 vdd.n3012 vdd.n3011 0.152939
R20094 vdd.n3012 vdd.n466 0.152939
R20095 vdd.n3016 vdd.n466 0.152939
R20096 vdd.n2806 vdd.n514 0.152939
R20097 vdd.n2049 vdd.n895 0.152939
R20098 vdd.n1219 vdd.n1218 0.152939
R20099 vdd.n1220 vdd.n1219 0.152939
R20100 vdd.n1220 vdd.n969 0.152939
R20101 vdd.n1234 vdd.n969 0.152939
R20102 vdd.n1235 vdd.n1234 0.152939
R20103 vdd.n1236 vdd.n1235 0.152939
R20104 vdd.n1236 vdd.n956 0.152939
R20105 vdd.n1250 vdd.n956 0.152939
R20106 vdd.n1251 vdd.n1250 0.152939
R20107 vdd.n1252 vdd.n1251 0.152939
R20108 vdd.n1252 vdd.n945 0.152939
R20109 vdd.n1267 vdd.n945 0.152939
R20110 vdd.n1268 vdd.n1267 0.152939
R20111 vdd.n1269 vdd.n1268 0.152939
R20112 vdd.n1269 vdd.n934 0.152939
R20113 vdd.n1565 vdd.n934 0.152939
R20114 vdd.n1566 vdd.n1565 0.152939
R20115 vdd.n1567 vdd.n1566 0.152939
R20116 vdd.n1567 vdd.n922 0.152939
R20117 vdd.n1582 vdd.n922 0.152939
R20118 vdd.n1583 vdd.n1582 0.152939
R20119 vdd.n1584 vdd.n1583 0.152939
R20120 vdd.n1584 vdd.n912 0.152939
R20121 vdd.n1599 vdd.n912 0.152939
R20122 vdd.n1600 vdd.n1599 0.152939
R20123 vdd.n1603 vdd.n1600 0.152939
R20124 vdd.n1603 vdd.n1602 0.152939
R20125 vdd.n1602 vdd.n1601 0.152939
R20126 vdd.n1211 vdd.n985 0.152939
R20127 vdd.n1207 vdd.n985 0.152939
R20128 vdd.n1207 vdd.n1206 0.152939
R20129 vdd.n1206 vdd.n1205 0.152939
R20130 vdd.n1205 vdd.n990 0.152939
R20131 vdd.n1201 vdd.n990 0.152939
R20132 vdd.n1201 vdd.n1200 0.152939
R20133 vdd.n1200 vdd.n1199 0.152939
R20134 vdd.n1199 vdd.n998 0.152939
R20135 vdd.n1195 vdd.n998 0.152939
R20136 vdd.n1195 vdd.n1194 0.152939
R20137 vdd.n1194 vdd.n1193 0.152939
R20138 vdd.n1193 vdd.n1006 0.152939
R20139 vdd.n1189 vdd.n1006 0.152939
R20140 vdd.n1189 vdd.n1188 0.152939
R20141 vdd.n1188 vdd.n1187 0.152939
R20142 vdd.n1187 vdd.n1014 0.152939
R20143 vdd.n1183 vdd.n1014 0.152939
R20144 vdd.n1183 vdd.n1182 0.152939
R20145 vdd.n1182 vdd.n1181 0.152939
R20146 vdd.n1181 vdd.n1024 0.152939
R20147 vdd.n1177 vdd.n1024 0.152939
R20148 vdd.n1177 vdd.n1176 0.152939
R20149 vdd.n1176 vdd.n1175 0.152939
R20150 vdd.n1175 vdd.n1032 0.152939
R20151 vdd.n1171 vdd.n1032 0.152939
R20152 vdd.n1171 vdd.n1170 0.152939
R20153 vdd.n1170 vdd.n1169 0.152939
R20154 vdd.n1169 vdd.n1040 0.152939
R20155 vdd.n1165 vdd.n1040 0.152939
R20156 vdd.n1165 vdd.n1164 0.152939
R20157 vdd.n1164 vdd.n1163 0.152939
R20158 vdd.n1163 vdd.n1048 0.152939
R20159 vdd.n1159 vdd.n1048 0.152939
R20160 vdd.n1159 vdd.n1158 0.152939
R20161 vdd.n1158 vdd.n1157 0.152939
R20162 vdd.n1157 vdd.n1056 0.152939
R20163 vdd.n1153 vdd.n1056 0.152939
R20164 vdd.n1153 vdd.n1152 0.152939
R20165 vdd.n1152 vdd.n1151 0.152939
R20166 vdd.n1151 vdd.n1064 0.152939
R20167 vdd.n1071 vdd.n1064 0.152939
R20168 vdd.n1141 vdd.n1071 0.152939
R20169 vdd.n1141 vdd.n1140 0.152939
R20170 vdd.n1140 vdd.n1139 0.152939
R20171 vdd.n1139 vdd.n1072 0.152939
R20172 vdd.n1135 vdd.n1072 0.152939
R20173 vdd.n1135 vdd.n1134 0.152939
R20174 vdd.n1134 vdd.n1133 0.152939
R20175 vdd.n1133 vdd.n1079 0.152939
R20176 vdd.n1129 vdd.n1079 0.152939
R20177 vdd.n1129 vdd.n1128 0.152939
R20178 vdd.n1128 vdd.n1127 0.152939
R20179 vdd.n1127 vdd.n1087 0.152939
R20180 vdd.n1123 vdd.n1087 0.152939
R20181 vdd.n1123 vdd.n1122 0.152939
R20182 vdd.n1122 vdd.n1121 0.152939
R20183 vdd.n1121 vdd.n1095 0.152939
R20184 vdd.n1117 vdd.n1095 0.152939
R20185 vdd.n1117 vdd.n1116 0.152939
R20186 vdd.n1116 vdd.n1115 0.152939
R20187 vdd.n1115 vdd.n1103 0.152939
R20188 vdd.n1103 vdd.n980 0.152939
R20189 vdd.n1212 vdd.n975 0.152939
R20190 vdd.n1226 vdd.n975 0.152939
R20191 vdd.n1227 vdd.n1226 0.152939
R20192 vdd.n1228 vdd.n1227 0.152939
R20193 vdd.n1228 vdd.n963 0.152939
R20194 vdd.n1242 vdd.n963 0.152939
R20195 vdd.n1243 vdd.n1242 0.152939
R20196 vdd.n1244 vdd.n1243 0.152939
R20197 vdd.n1244 vdd.n951 0.152939
R20198 vdd.n1259 vdd.n951 0.152939
R20199 vdd.n1260 vdd.n1259 0.152939
R20200 vdd.n1261 vdd.n1260 0.152939
R20201 vdd.n1261 vdd.n940 0.152939
R20202 vdd.n1558 vdd.n1557 0.145814
R20203 vdd.n3167 vdd.n310 0.145814
R20204 vdd.n3167 vdd.n311 0.145814
R20205 vdd.n1557 vdd.n940 0.145814
R20206 vdd.n2027 vdd.n1612 0.110256
R20207 vdd.n2737 vdd.n518 0.110256
R20208 vdd.n2806 vdd.n2805 0.110256
R20209 vdd.n2050 vdd.n2049 0.110256
R20210 vdd.n2027 vdd.n1813 0.0431829
R20211 vdd.n2050 vdd.n892 0.0431829
R20212 vdd.n2737 vdd.n524 0.0431829
R20213 vdd.n2805 vdd.n605 0.0431829
R20214 vdd vdd.n28 0.00833333
R20215 a_n6308_8799.n133 a_n6308_8799.t75 490.524
R20216 a_n6308_8799.n144 a_n6308_8799.t82 490.524
R20217 a_n6308_8799.n156 a_n6308_8799.t92 490.524
R20218 a_n6308_8799.n99 a_n6308_8799.t52 490.524
R20219 a_n6308_8799.n110 a_n6308_8799.t58 490.524
R20220 a_n6308_8799.n122 a_n6308_8799.t91 490.524
R20221 a_n6308_8799.n29 a_n6308_8799.t61 484.3
R20222 a_n6308_8799.n139 a_n6308_8799.t60 464.166
R20223 a_n6308_8799.n138 a_n6308_8799.t42 464.166
R20224 a_n6308_8799.n129 a_n6308_8799.t88 464.166
R20225 a_n6308_8799.n137 a_n6308_8799.t62 464.166
R20226 a_n6308_8799.n136 a_n6308_8799.t47 464.166
R20227 a_n6308_8799.n130 a_n6308_8799.t90 464.166
R20228 a_n6308_8799.n135 a_n6308_8799.t72 464.166
R20229 a_n6308_8799.n134 a_n6308_8799.t70 464.166
R20230 a_n6308_8799.n131 a_n6308_8799.t31 464.166
R20231 a_n6308_8799.n132 a_n6308_8799.t76 464.166
R20232 a_n6308_8799.n38 a_n6308_8799.t66 484.3
R20233 a_n6308_8799.n150 a_n6308_8799.t65 464.166
R20234 a_n6308_8799.n149 a_n6308_8799.t54 464.166
R20235 a_n6308_8799.n140 a_n6308_8799.t96 464.166
R20236 a_n6308_8799.n148 a_n6308_8799.t69 464.166
R20237 a_n6308_8799.n147 a_n6308_8799.t55 464.166
R20238 a_n6308_8799.n141 a_n6308_8799.t28 464.166
R20239 a_n6308_8799.n146 a_n6308_8799.t81 464.166
R20240 a_n6308_8799.n145 a_n6308_8799.t80 464.166
R20241 a_n6308_8799.n142 a_n6308_8799.t38 464.166
R20242 a_n6308_8799.n143 a_n6308_8799.t83 464.166
R20243 a_n6308_8799.n47 a_n6308_8799.t98 484.3
R20244 a_n6308_8799.n162 a_n6308_8799.t40 464.166
R20245 a_n6308_8799.n161 a_n6308_8799.t67 464.166
R20246 a_n6308_8799.n152 a_n6308_8799.t30 464.166
R20247 a_n6308_8799.n160 a_n6308_8799.t85 464.166
R20248 a_n6308_8799.n159 a_n6308_8799.t46 464.166
R20249 a_n6308_8799.n153 a_n6308_8799.t73 464.166
R20250 a_n6308_8799.n158 a_n6308_8799.t32 464.166
R20251 a_n6308_8799.n157 a_n6308_8799.t50 464.166
R20252 a_n6308_8799.n154 a_n6308_8799.t94 464.166
R20253 a_n6308_8799.n155 a_n6308_8799.t78 464.166
R20254 a_n6308_8799.n98 a_n6308_8799.t53 464.166
R20255 a_n6308_8799.n97 a_n6308_8799.t77 464.166
R20256 a_n6308_8799.n100 a_n6308_8799.t29 464.166
R20257 a_n6308_8799.n96 a_n6308_8799.t49 464.166
R20258 a_n6308_8799.n101 a_n6308_8799.t64 464.166
R20259 a_n6308_8799.n102 a_n6308_8799.t89 464.166
R20260 a_n6308_8799.n95 a_n6308_8799.t36 464.166
R20261 a_n6308_8799.n103 a_n6308_8799.t48 464.166
R20262 a_n6308_8799.n94 a_n6308_8799.t87 464.166
R20263 a_n6308_8799.n104 a_n6308_8799.t35 464.166
R20264 a_n6308_8799.n109 a_n6308_8799.t59 464.166
R20265 a_n6308_8799.n108 a_n6308_8799.t84 464.166
R20266 a_n6308_8799.n111 a_n6308_8799.t37 464.166
R20267 a_n6308_8799.n107 a_n6308_8799.t57 464.166
R20268 a_n6308_8799.n112 a_n6308_8799.t71 464.166
R20269 a_n6308_8799.n113 a_n6308_8799.t97 464.166
R20270 a_n6308_8799.n106 a_n6308_8799.t45 464.166
R20271 a_n6308_8799.n114 a_n6308_8799.t56 464.166
R20272 a_n6308_8799.n105 a_n6308_8799.t93 464.166
R20273 a_n6308_8799.n115 a_n6308_8799.t41 464.166
R20274 a_n6308_8799.n121 a_n6308_8799.t79 464.166
R20275 a_n6308_8799.n120 a_n6308_8799.t95 464.166
R20276 a_n6308_8799.n123 a_n6308_8799.t63 464.166
R20277 a_n6308_8799.n119 a_n6308_8799.t33 464.166
R20278 a_n6308_8799.n124 a_n6308_8799.t74 464.166
R20279 a_n6308_8799.n125 a_n6308_8799.t44 464.166
R20280 a_n6308_8799.n118 a_n6308_8799.t86 464.166
R20281 a_n6308_8799.n126 a_n6308_8799.t51 464.166
R20282 a_n6308_8799.n117 a_n6308_8799.t68 464.166
R20283 a_n6308_8799.n127 a_n6308_8799.t39 464.166
R20284 a_n6308_8799.n37 a_n6308_8799.n36 75.3623
R20285 a_n6308_8799.n35 a_n6308_8799.n20 70.3058
R20286 a_n6308_8799.n20 a_n6308_8799.n34 70.1674
R20287 a_n6308_8799.n34 a_n6308_8799.n130 20.9683
R20288 a_n6308_8799.n33 a_n6308_8799.n21 75.0448
R20289 a_n6308_8799.n136 a_n6308_8799.n33 11.2134
R20290 a_n6308_8799.n32 a_n6308_8799.n21 80.4688
R20291 a_n6308_8799.n23 a_n6308_8799.n31 74.73
R20292 a_n6308_8799.n30 a_n6308_8799.n23 70.1674
R20293 a_n6308_8799.n139 a_n6308_8799.n30 20.9683
R20294 a_n6308_8799.n22 a_n6308_8799.n29 70.5844
R20295 a_n6308_8799.n46 a_n6308_8799.n45 75.3623
R20296 a_n6308_8799.n44 a_n6308_8799.n16 70.3058
R20297 a_n6308_8799.n16 a_n6308_8799.n43 70.1674
R20298 a_n6308_8799.n43 a_n6308_8799.n141 20.9683
R20299 a_n6308_8799.n42 a_n6308_8799.n17 75.0448
R20300 a_n6308_8799.n147 a_n6308_8799.n42 11.2134
R20301 a_n6308_8799.n41 a_n6308_8799.n17 80.4688
R20302 a_n6308_8799.n19 a_n6308_8799.n40 74.73
R20303 a_n6308_8799.n39 a_n6308_8799.n19 70.1674
R20304 a_n6308_8799.n150 a_n6308_8799.n39 20.9683
R20305 a_n6308_8799.n18 a_n6308_8799.n38 70.5844
R20306 a_n6308_8799.n55 a_n6308_8799.n54 75.3623
R20307 a_n6308_8799.n53 a_n6308_8799.n12 70.3058
R20308 a_n6308_8799.n12 a_n6308_8799.n52 70.1674
R20309 a_n6308_8799.n52 a_n6308_8799.n153 20.9683
R20310 a_n6308_8799.n51 a_n6308_8799.n13 75.0448
R20311 a_n6308_8799.n159 a_n6308_8799.n51 11.2134
R20312 a_n6308_8799.n50 a_n6308_8799.n13 80.4688
R20313 a_n6308_8799.n15 a_n6308_8799.n49 74.73
R20314 a_n6308_8799.n48 a_n6308_8799.n15 70.1674
R20315 a_n6308_8799.n162 a_n6308_8799.n48 20.9683
R20316 a_n6308_8799.n14 a_n6308_8799.n47 70.5844
R20317 a_n6308_8799.n8 a_n6308_8799.n64 70.5844
R20318 a_n6308_8799.n63 a_n6308_8799.n9 70.1674
R20319 a_n6308_8799.n63 a_n6308_8799.n94 20.9683
R20320 a_n6308_8799.n9 a_n6308_8799.n62 74.73
R20321 a_n6308_8799.n103 a_n6308_8799.n62 11.843
R20322 a_n6308_8799.n61 a_n6308_8799.n10 80.4688
R20323 a_n6308_8799.n61 a_n6308_8799.n95 0.365327
R20324 a_n6308_8799.n10 a_n6308_8799.n60 75.0448
R20325 a_n6308_8799.n59 a_n6308_8799.n11 70.1674
R20326 a_n6308_8799.n59 a_n6308_8799.n96 20.9683
R20327 a_n6308_8799.n11 a_n6308_8799.n58 70.3058
R20328 a_n6308_8799.n100 a_n6308_8799.n58 20.6913
R20329 a_n6308_8799.n57 a_n6308_8799.n56 75.3623
R20330 a_n6308_8799.n4 a_n6308_8799.n73 70.5844
R20331 a_n6308_8799.n72 a_n6308_8799.n5 70.1674
R20332 a_n6308_8799.n72 a_n6308_8799.n105 20.9683
R20333 a_n6308_8799.n5 a_n6308_8799.n71 74.73
R20334 a_n6308_8799.n114 a_n6308_8799.n71 11.843
R20335 a_n6308_8799.n70 a_n6308_8799.n6 80.4688
R20336 a_n6308_8799.n70 a_n6308_8799.n106 0.365327
R20337 a_n6308_8799.n6 a_n6308_8799.n69 75.0448
R20338 a_n6308_8799.n68 a_n6308_8799.n7 70.1674
R20339 a_n6308_8799.n68 a_n6308_8799.n107 20.9683
R20340 a_n6308_8799.n7 a_n6308_8799.n67 70.3058
R20341 a_n6308_8799.n111 a_n6308_8799.n67 20.6913
R20342 a_n6308_8799.n66 a_n6308_8799.n65 75.3623
R20343 a_n6308_8799.n0 a_n6308_8799.n82 70.5844
R20344 a_n6308_8799.n81 a_n6308_8799.n1 70.1674
R20345 a_n6308_8799.n81 a_n6308_8799.n117 20.9683
R20346 a_n6308_8799.n1 a_n6308_8799.n80 74.73
R20347 a_n6308_8799.n126 a_n6308_8799.n80 11.843
R20348 a_n6308_8799.n79 a_n6308_8799.n2 80.4688
R20349 a_n6308_8799.n79 a_n6308_8799.n118 0.365327
R20350 a_n6308_8799.n2 a_n6308_8799.n78 75.0448
R20351 a_n6308_8799.n77 a_n6308_8799.n3 70.1674
R20352 a_n6308_8799.n77 a_n6308_8799.n119 20.9683
R20353 a_n6308_8799.n3 a_n6308_8799.n76 70.3058
R20354 a_n6308_8799.n123 a_n6308_8799.n76 20.6913
R20355 a_n6308_8799.n75 a_n6308_8799.n74 75.3623
R20356 a_n6308_8799.n24 a_n6308_8799.n83 98.9633
R20357 a_n6308_8799.n25 a_n6308_8799.n168 98.9631
R20358 a_n6308_8799.n25 a_n6308_8799.n167 98.6055
R20359 a_n6308_8799.n24 a_n6308_8799.n85 98.6055
R20360 a_n6308_8799.n24 a_n6308_8799.n84 98.6055
R20361 a_n6308_8799.n169 a_n6308_8799.n25 98.6054
R20362 a_n6308_8799.n27 a_n6308_8799.n86 81.2902
R20363 a_n6308_8799.n28 a_n6308_8799.n90 81.2902
R20364 a_n6308_8799.n28 a_n6308_8799.n88 81.2902
R20365 a_n6308_8799.n26 a_n6308_8799.n92 80.9324
R20366 a_n6308_8799.n27 a_n6308_8799.n93 80.9324
R20367 a_n6308_8799.n27 a_n6308_8799.n87 80.9324
R20368 a_n6308_8799.n28 a_n6308_8799.n91 80.9324
R20369 a_n6308_8799.n28 a_n6308_8799.n89 80.9324
R20370 a_n6308_8799.n30 a_n6308_8799.n138 20.9683
R20371 a_n6308_8799.n137 a_n6308_8799.n136 48.2005
R20372 a_n6308_8799.n135 a_n6308_8799.n34 20.9683
R20373 a_n6308_8799.n132 a_n6308_8799.n131 48.2005
R20374 a_n6308_8799.n39 a_n6308_8799.n149 20.9683
R20375 a_n6308_8799.n148 a_n6308_8799.n147 48.2005
R20376 a_n6308_8799.n146 a_n6308_8799.n43 20.9683
R20377 a_n6308_8799.n143 a_n6308_8799.n142 48.2005
R20378 a_n6308_8799.n48 a_n6308_8799.n161 20.9683
R20379 a_n6308_8799.n160 a_n6308_8799.n159 48.2005
R20380 a_n6308_8799.n158 a_n6308_8799.n52 20.9683
R20381 a_n6308_8799.n155 a_n6308_8799.n154 48.2005
R20382 a_n6308_8799.n98 a_n6308_8799.n97 48.2005
R20383 a_n6308_8799.n101 a_n6308_8799.n59 20.9683
R20384 a_n6308_8799.n102 a_n6308_8799.n95 48.2005
R20385 a_n6308_8799.n104 a_n6308_8799.n63 20.9683
R20386 a_n6308_8799.n109 a_n6308_8799.n108 48.2005
R20387 a_n6308_8799.n112 a_n6308_8799.n68 20.9683
R20388 a_n6308_8799.n113 a_n6308_8799.n106 48.2005
R20389 a_n6308_8799.n115 a_n6308_8799.n72 20.9683
R20390 a_n6308_8799.n121 a_n6308_8799.n120 48.2005
R20391 a_n6308_8799.n124 a_n6308_8799.n77 20.9683
R20392 a_n6308_8799.n125 a_n6308_8799.n118 48.2005
R20393 a_n6308_8799.n127 a_n6308_8799.n81 20.9683
R20394 a_n6308_8799.n32 a_n6308_8799.n129 47.835
R20395 a_n6308_8799.n35 a_n6308_8799.n134 20.6913
R20396 a_n6308_8799.n41 a_n6308_8799.n140 47.835
R20397 a_n6308_8799.n44 a_n6308_8799.n145 20.6913
R20398 a_n6308_8799.n50 a_n6308_8799.n152 47.835
R20399 a_n6308_8799.n53 a_n6308_8799.n157 20.6913
R20400 a_n6308_8799.n96 a_n6308_8799.n58 21.4216
R20401 a_n6308_8799.n107 a_n6308_8799.n67 21.4216
R20402 a_n6308_8799.n119 a_n6308_8799.n76 21.4216
R20403 a_n6308_8799.t34 a_n6308_8799.n64 484.3
R20404 a_n6308_8799.t43 a_n6308_8799.n73 484.3
R20405 a_n6308_8799.t99 a_n6308_8799.n82 484.3
R20406 a_n6308_8799.n57 a_n6308_8799.n99 45.0871
R20407 a_n6308_8799.n66 a_n6308_8799.n110 45.0871
R20408 a_n6308_8799.n75 a_n6308_8799.n122 45.0871
R20409 a_n6308_8799.n37 a_n6308_8799.n133 45.0871
R20410 a_n6308_8799.n46 a_n6308_8799.n144 45.0871
R20411 a_n6308_8799.n55 a_n6308_8799.n156 45.0871
R20412 a_n6308_8799.n31 a_n6308_8799.n129 11.843
R20413 a_n6308_8799.n134 a_n6308_8799.n36 36.139
R20414 a_n6308_8799.n40 a_n6308_8799.n140 11.843
R20415 a_n6308_8799.n145 a_n6308_8799.n45 36.139
R20416 a_n6308_8799.n49 a_n6308_8799.n152 11.843
R20417 a_n6308_8799.n157 a_n6308_8799.n54 36.139
R20418 a_n6308_8799.n100 a_n6308_8799.n56 36.139
R20419 a_n6308_8799.n94 a_n6308_8799.n62 34.4824
R20420 a_n6308_8799.n111 a_n6308_8799.n65 36.139
R20421 a_n6308_8799.n105 a_n6308_8799.n71 34.4824
R20422 a_n6308_8799.n123 a_n6308_8799.n74 36.139
R20423 a_n6308_8799.n117 a_n6308_8799.n80 34.4824
R20424 a_n6308_8799.n33 a_n6308_8799.n130 35.3134
R20425 a_n6308_8799.n42 a_n6308_8799.n141 35.3134
R20426 a_n6308_8799.n51 a_n6308_8799.n153 35.3134
R20427 a_n6308_8799.n60 a_n6308_8799.n101 35.3134
R20428 a_n6308_8799.n102 a_n6308_8799.n60 11.2134
R20429 a_n6308_8799.n69 a_n6308_8799.n112 35.3134
R20430 a_n6308_8799.n113 a_n6308_8799.n69 11.2134
R20431 a_n6308_8799.n78 a_n6308_8799.n124 35.3134
R20432 a_n6308_8799.n125 a_n6308_8799.n78 11.2134
R20433 a_n6308_8799.n138 a_n6308_8799.n31 34.4824
R20434 a_n6308_8799.n36 a_n6308_8799.n131 10.5784
R20435 a_n6308_8799.n149 a_n6308_8799.n40 34.4824
R20436 a_n6308_8799.n45 a_n6308_8799.n142 10.5784
R20437 a_n6308_8799.n161 a_n6308_8799.n49 34.4824
R20438 a_n6308_8799.n54 a_n6308_8799.n154 10.5784
R20439 a_n6308_8799.n56 a_n6308_8799.n97 10.5784
R20440 a_n6308_8799.n65 a_n6308_8799.n108 10.5784
R20441 a_n6308_8799.n74 a_n6308_8799.n120 10.5784
R20442 a_n6308_8799.n133 a_n6308_8799.n132 14.1472
R20443 a_n6308_8799.n144 a_n6308_8799.n143 14.1472
R20444 a_n6308_8799.n156 a_n6308_8799.n155 14.1472
R20445 a_n6308_8799.n99 a_n6308_8799.n98 14.1472
R20446 a_n6308_8799.n110 a_n6308_8799.n109 14.1472
R20447 a_n6308_8799.n122 a_n6308_8799.n121 14.1472
R20448 a_n6308_8799.n165 a_n6308_8799.n27 12.3339
R20449 a_n6308_8799.n166 a_n6308_8799.n165 11.4887
R20450 a_n6308_8799.n151 a_n6308_8799.n22 9.01755
R20451 a_n6308_8799.n116 a_n6308_8799.n8 9.01755
R20452 a_n6308_8799.n164 a_n6308_8799.n128 6.81251
R20453 a_n6308_8799.n164 a_n6308_8799.n163 6.5703
R20454 a_n6308_8799.n151 a_n6308_8799.n18 4.90959
R20455 a_n6308_8799.n163 a_n6308_8799.n14 4.90959
R20456 a_n6308_8799.n116 a_n6308_8799.n4 4.90959
R20457 a_n6308_8799.n128 a_n6308_8799.n0 4.90959
R20458 a_n6308_8799.n163 a_n6308_8799.n151 4.10845
R20459 a_n6308_8799.n128 a_n6308_8799.n116 4.10845
R20460 a_n6308_8799.n168 a_n6308_8799.t12 3.61217
R20461 a_n6308_8799.n168 a_n6308_8799.t18 3.61217
R20462 a_n6308_8799.n167 a_n6308_8799.t19 3.61217
R20463 a_n6308_8799.n167 a_n6308_8799.t10 3.61217
R20464 a_n6308_8799.n85 a_n6308_8799.t11 3.61217
R20465 a_n6308_8799.n85 a_n6308_8799.t22 3.61217
R20466 a_n6308_8799.n84 a_n6308_8799.t16 3.61217
R20467 a_n6308_8799.n84 a_n6308_8799.t25 3.61217
R20468 a_n6308_8799.n83 a_n6308_8799.t1 3.61217
R20469 a_n6308_8799.n83 a_n6308_8799.t7 3.61217
R20470 a_n6308_8799.n169 a_n6308_8799.t17 3.61217
R20471 a_n6308_8799.t0 a_n6308_8799.n169 3.61217
R20472 a_n6308_8799.n165 a_n6308_8799.n164 3.4105
R20473 a_n6308_8799.n92 a_n6308_8799.t13 2.82907
R20474 a_n6308_8799.n92 a_n6308_8799.t27 2.82907
R20475 a_n6308_8799.n93 a_n6308_8799.t24 2.82907
R20476 a_n6308_8799.n93 a_n6308_8799.t20 2.82907
R20477 a_n6308_8799.n87 a_n6308_8799.t9 2.82907
R20478 a_n6308_8799.n87 a_n6308_8799.t2 2.82907
R20479 a_n6308_8799.n86 a_n6308_8799.t23 2.82907
R20480 a_n6308_8799.n86 a_n6308_8799.t5 2.82907
R20481 a_n6308_8799.n90 a_n6308_8799.t3 2.82907
R20482 a_n6308_8799.n90 a_n6308_8799.t6 2.82907
R20483 a_n6308_8799.n91 a_n6308_8799.t4 2.82907
R20484 a_n6308_8799.n91 a_n6308_8799.t8 2.82907
R20485 a_n6308_8799.n89 a_n6308_8799.t14 2.82907
R20486 a_n6308_8799.n89 a_n6308_8799.t21 2.82907
R20487 a_n6308_8799.n88 a_n6308_8799.t26 2.82907
R20488 a_n6308_8799.n88 a_n6308_8799.t15 2.82907
R20489 a_n6308_8799.n29 a_n6308_8799.n139 22.3251
R20490 a_n6308_8799.n38 a_n6308_8799.n150 22.3251
R20491 a_n6308_8799.n47 a_n6308_8799.n162 22.3251
R20492 a_n6308_8799.n64 a_n6308_8799.n104 22.3251
R20493 a_n6308_8799.n73 a_n6308_8799.n115 22.3251
R20494 a_n6308_8799.n82 a_n6308_8799.n127 22.3251
R20495 a_n6308_8799.n32 a_n6308_8799.n137 0.365327
R20496 a_n6308_8799.n135 a_n6308_8799.n35 21.4216
R20497 a_n6308_8799.n41 a_n6308_8799.n148 0.365327
R20498 a_n6308_8799.n146 a_n6308_8799.n44 21.4216
R20499 a_n6308_8799.n50 a_n6308_8799.n160 0.365327
R20500 a_n6308_8799.n158 a_n6308_8799.n53 21.4216
R20501 a_n6308_8799.n103 a_n6308_8799.n61 47.835
R20502 a_n6308_8799.n114 a_n6308_8799.n70 47.835
R20503 a_n6308_8799.n126 a_n6308_8799.n79 47.835
R20504 a_n6308_8799.n26 a_n6308_8799.n28 31.7978
R20505 a_n6308_8799.n25 a_n6308_8799.n166 30.6769
R20506 a_n6308_8799.n166 a_n6308_8799.n24 18.4882
R20507 a_n6308_8799.n23 a_n6308_8799.n21 0.758076
R20508 a_n6308_8799.n21 a_n6308_8799.n20 0.758076
R20509 a_n6308_8799.n37 a_n6308_8799.n20 0.758076
R20510 a_n6308_8799.n19 a_n6308_8799.n17 0.758076
R20511 a_n6308_8799.n17 a_n6308_8799.n16 0.758076
R20512 a_n6308_8799.n46 a_n6308_8799.n16 0.758076
R20513 a_n6308_8799.n15 a_n6308_8799.n13 0.758076
R20514 a_n6308_8799.n13 a_n6308_8799.n12 0.758076
R20515 a_n6308_8799.n55 a_n6308_8799.n12 0.758076
R20516 a_n6308_8799.n11 a_n6308_8799.n10 0.758076
R20517 a_n6308_8799.n10 a_n6308_8799.n9 0.758076
R20518 a_n6308_8799.n9 a_n6308_8799.n8 0.758076
R20519 a_n6308_8799.n7 a_n6308_8799.n6 0.758076
R20520 a_n6308_8799.n6 a_n6308_8799.n5 0.758076
R20521 a_n6308_8799.n5 a_n6308_8799.n4 0.758076
R20522 a_n6308_8799.n3 a_n6308_8799.n2 0.758076
R20523 a_n6308_8799.n2 a_n6308_8799.n1 0.758076
R20524 a_n6308_8799.n1 a_n6308_8799.n0 0.758076
R20525 a_n6308_8799.n27 a_n6308_8799.n26 0.716017
R20526 a_n6308_8799.n75 a_n6308_8799.n3 0.568682
R20527 a_n6308_8799.n66 a_n6308_8799.n7 0.568682
R20528 a_n6308_8799.n57 a_n6308_8799.n11 0.568682
R20529 a_n6308_8799.n15 a_n6308_8799.n14 0.568682
R20530 a_n6308_8799.n19 a_n6308_8799.n18 0.568682
R20531 a_n6308_8799.n23 a_n6308_8799.n22 0.568682
R20532 a_n1986_13878.n3 a_n1986_13878.t20 539.01
R20533 a_n1986_13878.n91 a_n1986_13878.t2 512.366
R20534 a_n1986_13878.n90 a_n1986_13878.t12 512.366
R20535 a_n1986_13878.n52 a_n1986_13878.t18 512.366
R20536 a_n1986_13878.n89 a_n1986_13878.t8 512.366
R20537 a_n1986_13878.n7 a_n1986_13878.t67 539.01
R20538 a_n1986_13878.n80 a_n1986_13878.t50 512.366
R20539 a_n1986_13878.n79 a_n1986_13878.t54 512.366
R20540 a_n1986_13878.n53 a_n1986_13878.t44 512.366
R20541 a_n1986_13878.n78 a_n1986_13878.t59 512.366
R20542 a_n1986_13878.n20 a_n1986_13878.t22 539.01
R20543 a_n1986_13878.n61 a_n1986_13878.t16 512.366
R20544 a_n1986_13878.n62 a_n1986_13878.t6 512.366
R20545 a_n1986_13878.n56 a_n1986_13878.t4 512.366
R20546 a_n1986_13878.n63 a_n1986_13878.t14 512.366
R20547 a_n1986_13878.n24 a_n1986_13878.t62 539.01
R20548 a_n1986_13878.n58 a_n1986_13878.t63 512.366
R20549 a_n1986_13878.n59 a_n1986_13878.t42 512.366
R20550 a_n1986_13878.n57 a_n1986_13878.t48 512.366
R20551 a_n1986_13878.n60 a_n1986_13878.t57 512.366
R20552 a_n1986_13878.n75 a_n1986_13878.t56 512.366
R20553 a_n1986_13878.n65 a_n1986_13878.t47 512.366
R20554 a_n1986_13878.n76 a_n1986_13878.t41 512.366
R20555 a_n1986_13878.n73 a_n1986_13878.t64 512.366
R20556 a_n1986_13878.n66 a_n1986_13878.t53 512.366
R20557 a_n1986_13878.n74 a_n1986_13878.t52 512.366
R20558 a_n1986_13878.n71 a_n1986_13878.t60 512.366
R20559 a_n1986_13878.n67 a_n1986_13878.t45 512.366
R20560 a_n1986_13878.n72 a_n1986_13878.t46 512.366
R20561 a_n1986_13878.n69 a_n1986_13878.t49 512.366
R20562 a_n1986_13878.n68 a_n1986_13878.t58 512.366
R20563 a_n1986_13878.n70 a_n1986_13878.t40 512.366
R20564 a_n1986_13878.n51 a_n1986_13878.n0 70.3058
R20565 a_n1986_13878.n48 a_n1986_13878.n5 70.3058
R20566 a_n1986_13878.n17 a_n1986_13878.n37 70.3058
R20567 a_n1986_13878.n21 a_n1986_13878.n34 70.3058
R20568 a_n1986_13878.n33 a_n1986_13878.n22 70.1674
R20569 a_n1986_13878.n33 a_n1986_13878.n57 20.9683
R20570 a_n1986_13878.n22 a_n1986_13878.n32 75.0448
R20571 a_n1986_13878.n59 a_n1986_13878.n32 11.2134
R20572 a_n1986_13878.n23 a_n1986_13878.n24 44.8194
R20573 a_n1986_13878.n36 a_n1986_13878.n18 70.1674
R20574 a_n1986_13878.n36 a_n1986_13878.n56 20.9683
R20575 a_n1986_13878.n18 a_n1986_13878.n35 75.0448
R20576 a_n1986_13878.n62 a_n1986_13878.n35 11.2134
R20577 a_n1986_13878.n19 a_n1986_13878.n20 44.8194
R20578 a_n1986_13878.n8 a_n1986_13878.n45 70.1674
R20579 a_n1986_13878.n10 a_n1986_13878.n43 70.1674
R20580 a_n1986_13878.n12 a_n1986_13878.n41 70.1674
R20581 a_n1986_13878.n15 a_n1986_13878.n39 70.1674
R20582 a_n1986_13878.n70 a_n1986_13878.n39 20.9683
R20583 a_n1986_13878.n38 a_n1986_13878.n16 75.0448
R20584 a_n1986_13878.n38 a_n1986_13878.n68 11.2134
R20585 a_n1986_13878.n16 a_n1986_13878.n69 161.3
R20586 a_n1986_13878.n72 a_n1986_13878.n41 20.9683
R20587 a_n1986_13878.n40 a_n1986_13878.n13 75.0448
R20588 a_n1986_13878.n40 a_n1986_13878.n67 11.2134
R20589 a_n1986_13878.n13 a_n1986_13878.n71 161.3
R20590 a_n1986_13878.n74 a_n1986_13878.n43 20.9683
R20591 a_n1986_13878.n42 a_n1986_13878.n11 75.0448
R20592 a_n1986_13878.n42 a_n1986_13878.n66 11.2134
R20593 a_n1986_13878.n11 a_n1986_13878.n73 161.3
R20594 a_n1986_13878.n76 a_n1986_13878.n45 20.9683
R20595 a_n1986_13878.n44 a_n1986_13878.n9 75.0448
R20596 a_n1986_13878.n44 a_n1986_13878.n65 11.2134
R20597 a_n1986_13878.n9 a_n1986_13878.n75 161.3
R20598 a_n1986_13878.n6 a_n1986_13878.n47 70.1674
R20599 a_n1986_13878.n47 a_n1986_13878.n53 20.9683
R20600 a_n1986_13878.n46 a_n1986_13878.n6 75.0448
R20601 a_n1986_13878.n79 a_n1986_13878.n46 11.2134
R20602 a_n1986_13878.n4 a_n1986_13878.n7 44.8194
R20603 a_n1986_13878.n2 a_n1986_13878.n50 70.1674
R20604 a_n1986_13878.n50 a_n1986_13878.n52 20.9683
R20605 a_n1986_13878.n49 a_n1986_13878.n2 75.0448
R20606 a_n1986_13878.n90 a_n1986_13878.n49 11.2134
R20607 a_n1986_13878.n1 a_n1986_13878.n3 44.8194
R20608 a_n1986_13878.n30 a_n1986_13878.n87 81.2902
R20609 a_n1986_13878.n31 a_n1986_13878.n83 81.2902
R20610 a_n1986_13878.n31 a_n1986_13878.n81 81.2902
R20611 a_n1986_13878.n30 a_n1986_13878.n88 80.9324
R20612 a_n1986_13878.n30 a_n1986_13878.n86 80.9324
R20613 a_n1986_13878.n29 a_n1986_13878.n85 80.9324
R20614 a_n1986_13878.n31 a_n1986_13878.n84 80.9324
R20615 a_n1986_13878.n31 a_n1986_13878.n82 80.9324
R20616 a_n1986_13878.n25 a_n1986_13878.t23 74.6477
R20617 a_n1986_13878.t1 a_n1986_13878.n28 74.6477
R20618 a_n1986_13878.n27 a_n1986_13878.t21 74.2899
R20619 a_n1986_13878.n26 a_n1986_13878.t11 74.2897
R20620 a_n1986_13878.n28 a_n1986_13878.n94 70.6783
R20621 a_n1986_13878.n28 a_n1986_13878.n93 70.6783
R20622 a_n1986_13878.n26 a_n1986_13878.n55 70.6783
R20623 a_n1986_13878.n25 a_n1986_13878.n54 70.6783
R20624 a_n1986_13878.n91 a_n1986_13878.n90 48.2005
R20625 a_n1986_13878.n89 a_n1986_13878.n50 20.9683
R20626 a_n1986_13878.n80 a_n1986_13878.n79 48.2005
R20627 a_n1986_13878.n78 a_n1986_13878.n47 20.9683
R20628 a_n1986_13878.n62 a_n1986_13878.n61 48.2005
R20629 a_n1986_13878.n63 a_n1986_13878.n36 20.9683
R20630 a_n1986_13878.n59 a_n1986_13878.n58 48.2005
R20631 a_n1986_13878.n60 a_n1986_13878.n33 20.9683
R20632 a_n1986_13878.n75 a_n1986_13878.n65 48.2005
R20633 a_n1986_13878.t61 a_n1986_13878.n45 533.335
R20634 a_n1986_13878.n73 a_n1986_13878.n66 48.2005
R20635 a_n1986_13878.t66 a_n1986_13878.n43 533.335
R20636 a_n1986_13878.n71 a_n1986_13878.n67 48.2005
R20637 a_n1986_13878.t55 a_n1986_13878.n41 533.335
R20638 a_n1986_13878.n69 a_n1986_13878.n68 48.2005
R20639 a_n1986_13878.t51 a_n1986_13878.n39 533.335
R20640 a_n1986_13878.n51 a_n1986_13878.t0 533.058
R20641 a_n1986_13878.n48 a_n1986_13878.t65 533.058
R20642 a_n1986_13878.t10 a_n1986_13878.n37 533.058
R20643 a_n1986_13878.t43 a_n1986_13878.n34 533.058
R20644 a_n1986_13878.n49 a_n1986_13878.n52 35.3134
R20645 a_n1986_13878.n46 a_n1986_13878.n53 35.3134
R20646 a_n1986_13878.n56 a_n1986_13878.n35 35.3134
R20647 a_n1986_13878.n57 a_n1986_13878.n32 35.3134
R20648 a_n1986_13878.n76 a_n1986_13878.n44 35.3134
R20649 a_n1986_13878.n74 a_n1986_13878.n42 35.3134
R20650 a_n1986_13878.n72 a_n1986_13878.n40 35.3134
R20651 a_n1986_13878.n70 a_n1986_13878.n38 35.3134
R20652 a_n1986_13878.n29 a_n1986_13878.n31 31.0592
R20653 a_n1986_13878.n0 a_n1986_13878.n30 23.891
R20654 a_n1986_13878.n23 a_n1986_13878.n14 12.046
R20655 a_n1986_13878.n5 a_n1986_13878.n77 11.8414
R20656 a_n1986_13878.n92 a_n1986_13878.n1 10.5365
R20657 a_n1986_13878.n64 a_n1986_13878.n26 9.50122
R20658 a_n1986_13878.n16 a_n1986_13878.n14 7.47588
R20659 a_n1986_13878.n77 a_n1986_13878.n8 7.47588
R20660 a_n1986_13878.n64 a_n1986_13878.n17 6.70126
R20661 a_n1986_13878.n27 a_n1986_13878.n92 5.65783
R20662 a_n1986_13878.n77 a_n1986_13878.n64 5.3452
R20663 a_n1986_13878.n19 a_n1986_13878.n21 3.95126
R20664 a_n1986_13878.n94 a_n1986_13878.t19 3.61217
R20665 a_n1986_13878.n94 a_n1986_13878.t9 3.61217
R20666 a_n1986_13878.n93 a_n1986_13878.t3 3.61217
R20667 a_n1986_13878.n93 a_n1986_13878.t13 3.61217
R20668 a_n1986_13878.n55 a_n1986_13878.t5 3.61217
R20669 a_n1986_13878.n55 a_n1986_13878.t15 3.61217
R20670 a_n1986_13878.n54 a_n1986_13878.t17 3.61217
R20671 a_n1986_13878.n54 a_n1986_13878.t7 3.61217
R20672 a_n1986_13878.n0 a_n1986_13878.n4 3.42095
R20673 a_n1986_13878.n87 a_n1986_13878.t39 2.82907
R20674 a_n1986_13878.n87 a_n1986_13878.t37 2.82907
R20675 a_n1986_13878.n88 a_n1986_13878.t25 2.82907
R20676 a_n1986_13878.n88 a_n1986_13878.t38 2.82907
R20677 a_n1986_13878.n86 a_n1986_13878.t27 2.82907
R20678 a_n1986_13878.n86 a_n1986_13878.t33 2.82907
R20679 a_n1986_13878.n85 a_n1986_13878.t29 2.82907
R20680 a_n1986_13878.n85 a_n1986_13878.t28 2.82907
R20681 a_n1986_13878.n83 a_n1986_13878.t30 2.82907
R20682 a_n1986_13878.n83 a_n1986_13878.t26 2.82907
R20683 a_n1986_13878.n84 a_n1986_13878.t36 2.82907
R20684 a_n1986_13878.n84 a_n1986_13878.t31 2.82907
R20685 a_n1986_13878.n82 a_n1986_13878.t24 2.82907
R20686 a_n1986_13878.n82 a_n1986_13878.t34 2.82907
R20687 a_n1986_13878.n81 a_n1986_13878.t35 2.82907
R20688 a_n1986_13878.n81 a_n1986_13878.t32 2.82907
R20689 a_n1986_13878.n92 a_n1986_13878.n14 1.30542
R20690 a_n1986_13878.n11 a_n1986_13878.n12 1.04595
R20691 a_n1986_13878.n3 a_n1986_13878.n91 13.657
R20692 a_n1986_13878.n89 a_n1986_13878.n51 21.4216
R20693 a_n1986_13878.n7 a_n1986_13878.n80 13.657
R20694 a_n1986_13878.n78 a_n1986_13878.n48 21.4216
R20695 a_n1986_13878.n61 a_n1986_13878.n20 13.657
R20696 a_n1986_13878.n37 a_n1986_13878.n63 21.4216
R20697 a_n1986_13878.n58 a_n1986_13878.n24 13.657
R20698 a_n1986_13878.n34 a_n1986_13878.n60 21.4216
R20699 a_n1986_13878.n2 a_n1986_13878.n0 1.2505
R20700 a_n1986_13878.n23 a_n1986_13878.n22 0.758076
R20701 a_n1986_13878.n22 a_n1986_13878.n21 0.758076
R20702 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R20703 a_n1986_13878.n18 a_n1986_13878.n17 0.758076
R20704 a_n1986_13878.n16 a_n1986_13878.n15 0.758076
R20705 a_n1986_13878.n13 a_n1986_13878.n12 0.758076
R20706 a_n1986_13878.n11 a_n1986_13878.n10 0.758076
R20707 a_n1986_13878.n9 a_n1986_13878.n8 0.758076
R20708 a_n1986_13878.n6 a_n1986_13878.n4 0.758076
R20709 a_n1986_13878.n6 a_n1986_13878.n5 0.758076
R20710 a_n1986_13878.n2 a_n1986_13878.n1 0.758076
R20711 a_n1986_13878.n30 a_n1986_13878.n29 0.716017
R20712 a_n1986_13878.n28 a_n1986_13878.n27 0.716017
R20713 a_n1986_13878.n26 a_n1986_13878.n25 0.716017
R20714 a_n1986_13878.n13 a_n1986_13878.n15 0.67853
R20715 a_n1986_13878.n9 a_n1986_13878.n10 0.67853
R20716 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R20717 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R20718 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R20719 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20720 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20721 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R20722 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R20723 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R20724 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R20725 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R20726 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R20727 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R20728 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R20729 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R20730 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R20731 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R20732 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R20733 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R20734 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R20735 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R20736 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R20737 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R20738 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R20739 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R20740 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R20741 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R20742 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R20743 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R20744 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R20745 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R20746 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R20747 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R20748 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R20749 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R20750 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R20751 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R20752 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R20753 output.n41 output.n15 289.615
R20754 output.n72 output.n46 289.615
R20755 output.n104 output.n78 289.615
R20756 output.n136 output.n110 289.615
R20757 output.n77 output.n45 197.26
R20758 output.n77 output.n76 196.298
R20759 output.n109 output.n108 196.298
R20760 output.n141 output.n140 196.298
R20761 output.n42 output.n41 185
R20762 output.n40 output.n39 185
R20763 output.n19 output.n18 185
R20764 output.n34 output.n33 185
R20765 output.n32 output.n31 185
R20766 output.n23 output.n22 185
R20767 output.n26 output.n25 185
R20768 output.n73 output.n72 185
R20769 output.n71 output.n70 185
R20770 output.n50 output.n49 185
R20771 output.n65 output.n64 185
R20772 output.n63 output.n62 185
R20773 output.n54 output.n53 185
R20774 output.n57 output.n56 185
R20775 output.n105 output.n104 185
R20776 output.n103 output.n102 185
R20777 output.n82 output.n81 185
R20778 output.n97 output.n96 185
R20779 output.n95 output.n94 185
R20780 output.n86 output.n85 185
R20781 output.n89 output.n88 185
R20782 output.n137 output.n136 185
R20783 output.n135 output.n134 185
R20784 output.n114 output.n113 185
R20785 output.n129 output.n128 185
R20786 output.n127 output.n126 185
R20787 output.n118 output.n117 185
R20788 output.n121 output.n120 185
R20789 output.t0 output.n24 147.661
R20790 output.t19 output.n55 147.661
R20791 output.t2 output.n87 147.661
R20792 output.t1 output.n119 147.661
R20793 output.n41 output.n40 104.615
R20794 output.n40 output.n18 104.615
R20795 output.n33 output.n18 104.615
R20796 output.n33 output.n32 104.615
R20797 output.n32 output.n22 104.615
R20798 output.n25 output.n22 104.615
R20799 output.n72 output.n71 104.615
R20800 output.n71 output.n49 104.615
R20801 output.n64 output.n49 104.615
R20802 output.n64 output.n63 104.615
R20803 output.n63 output.n53 104.615
R20804 output.n56 output.n53 104.615
R20805 output.n104 output.n103 104.615
R20806 output.n103 output.n81 104.615
R20807 output.n96 output.n81 104.615
R20808 output.n96 output.n95 104.615
R20809 output.n95 output.n85 104.615
R20810 output.n88 output.n85 104.615
R20811 output.n136 output.n135 104.615
R20812 output.n135 output.n113 104.615
R20813 output.n128 output.n113 104.615
R20814 output.n128 output.n127 104.615
R20815 output.n127 output.n117 104.615
R20816 output.n120 output.n117 104.615
R20817 output.n1 output.t16 77.056
R20818 output.n14 output.t17 76.6694
R20819 output.n1 output.n0 72.7095
R20820 output.n3 output.n2 72.7095
R20821 output.n5 output.n4 72.7095
R20822 output.n7 output.n6 72.7095
R20823 output.n9 output.n8 72.7095
R20824 output.n11 output.n10 72.7095
R20825 output.n13 output.n12 72.7095
R20826 output.n25 output.t0 52.3082
R20827 output.n56 output.t19 52.3082
R20828 output.n88 output.t2 52.3082
R20829 output.n120 output.t1 52.3082
R20830 output.n26 output.n24 15.6674
R20831 output.n57 output.n55 15.6674
R20832 output.n89 output.n87 15.6674
R20833 output.n121 output.n119 15.6674
R20834 output.n27 output.n23 12.8005
R20835 output.n58 output.n54 12.8005
R20836 output.n90 output.n86 12.8005
R20837 output.n122 output.n118 12.8005
R20838 output.n31 output.n30 12.0247
R20839 output.n62 output.n61 12.0247
R20840 output.n94 output.n93 12.0247
R20841 output.n126 output.n125 12.0247
R20842 output.n34 output.n21 11.249
R20843 output.n65 output.n52 11.249
R20844 output.n97 output.n84 11.249
R20845 output.n129 output.n116 11.249
R20846 output.n35 output.n19 10.4732
R20847 output.n66 output.n50 10.4732
R20848 output.n98 output.n82 10.4732
R20849 output.n130 output.n114 10.4732
R20850 output.n39 output.n38 9.69747
R20851 output.n70 output.n69 9.69747
R20852 output.n102 output.n101 9.69747
R20853 output.n134 output.n133 9.69747
R20854 output.n45 output.n44 9.45567
R20855 output.n76 output.n75 9.45567
R20856 output.n108 output.n107 9.45567
R20857 output.n140 output.n139 9.45567
R20858 output.n44 output.n43 9.3005
R20859 output.n17 output.n16 9.3005
R20860 output.n38 output.n37 9.3005
R20861 output.n36 output.n35 9.3005
R20862 output.n21 output.n20 9.3005
R20863 output.n30 output.n29 9.3005
R20864 output.n28 output.n27 9.3005
R20865 output.n75 output.n74 9.3005
R20866 output.n48 output.n47 9.3005
R20867 output.n69 output.n68 9.3005
R20868 output.n67 output.n66 9.3005
R20869 output.n52 output.n51 9.3005
R20870 output.n61 output.n60 9.3005
R20871 output.n59 output.n58 9.3005
R20872 output.n107 output.n106 9.3005
R20873 output.n80 output.n79 9.3005
R20874 output.n101 output.n100 9.3005
R20875 output.n99 output.n98 9.3005
R20876 output.n84 output.n83 9.3005
R20877 output.n93 output.n92 9.3005
R20878 output.n91 output.n90 9.3005
R20879 output.n139 output.n138 9.3005
R20880 output.n112 output.n111 9.3005
R20881 output.n133 output.n132 9.3005
R20882 output.n131 output.n130 9.3005
R20883 output.n116 output.n115 9.3005
R20884 output.n125 output.n124 9.3005
R20885 output.n123 output.n122 9.3005
R20886 output.n42 output.n17 8.92171
R20887 output.n73 output.n48 8.92171
R20888 output.n105 output.n80 8.92171
R20889 output.n137 output.n112 8.92171
R20890 output output.n141 8.15037
R20891 output.n43 output.n15 8.14595
R20892 output.n74 output.n46 8.14595
R20893 output.n106 output.n78 8.14595
R20894 output.n138 output.n110 8.14595
R20895 output.n45 output.n15 5.81868
R20896 output.n76 output.n46 5.81868
R20897 output.n108 output.n78 5.81868
R20898 output.n140 output.n110 5.81868
R20899 output.n43 output.n42 5.04292
R20900 output.n74 output.n73 5.04292
R20901 output.n106 output.n105 5.04292
R20902 output.n138 output.n137 5.04292
R20903 output.n28 output.n24 4.38594
R20904 output.n59 output.n55 4.38594
R20905 output.n91 output.n87 4.38594
R20906 output.n123 output.n119 4.38594
R20907 output.n39 output.n17 4.26717
R20908 output.n70 output.n48 4.26717
R20909 output.n102 output.n80 4.26717
R20910 output.n134 output.n112 4.26717
R20911 output.n0 output.t5 3.9605
R20912 output.n0 output.t10 3.9605
R20913 output.n2 output.t14 3.9605
R20914 output.n2 output.t6 3.9605
R20915 output.n4 output.t9 3.9605
R20916 output.n4 output.t7 3.9605
R20917 output.n6 output.t13 3.9605
R20918 output.n6 output.t15 3.9605
R20919 output.n8 output.t18 3.9605
R20920 output.n8 output.t11 3.9605
R20921 output.n10 output.t12 3.9605
R20922 output.n10 output.t3 3.9605
R20923 output.n12 output.t4 3.9605
R20924 output.n12 output.t8 3.9605
R20925 output.n38 output.n19 3.49141
R20926 output.n69 output.n50 3.49141
R20927 output.n101 output.n82 3.49141
R20928 output.n133 output.n114 3.49141
R20929 output.n35 output.n34 2.71565
R20930 output.n66 output.n65 2.71565
R20931 output.n98 output.n97 2.71565
R20932 output.n130 output.n129 2.71565
R20933 output.n31 output.n21 1.93989
R20934 output.n62 output.n52 1.93989
R20935 output.n94 output.n84 1.93989
R20936 output.n126 output.n116 1.93989
R20937 output.n30 output.n23 1.16414
R20938 output.n61 output.n54 1.16414
R20939 output.n93 output.n86 1.16414
R20940 output.n125 output.n118 1.16414
R20941 output.n141 output.n109 0.962709
R20942 output.n109 output.n77 0.962709
R20943 output.n27 output.n26 0.388379
R20944 output.n58 output.n57 0.388379
R20945 output.n90 output.n89 0.388379
R20946 output.n122 output.n121 0.388379
R20947 output.n14 output.n13 0.387128
R20948 output.n13 output.n11 0.387128
R20949 output.n11 output.n9 0.387128
R20950 output.n9 output.n7 0.387128
R20951 output.n7 output.n5 0.387128
R20952 output.n5 output.n3 0.387128
R20953 output.n3 output.n1 0.387128
R20954 output.n44 output.n16 0.155672
R20955 output.n37 output.n16 0.155672
R20956 output.n37 output.n36 0.155672
R20957 output.n36 output.n20 0.155672
R20958 output.n29 output.n20 0.155672
R20959 output.n29 output.n28 0.155672
R20960 output.n75 output.n47 0.155672
R20961 output.n68 output.n47 0.155672
R20962 output.n68 output.n67 0.155672
R20963 output.n67 output.n51 0.155672
R20964 output.n60 output.n51 0.155672
R20965 output.n60 output.n59 0.155672
R20966 output.n107 output.n79 0.155672
R20967 output.n100 output.n79 0.155672
R20968 output.n100 output.n99 0.155672
R20969 output.n99 output.n83 0.155672
R20970 output.n92 output.n83 0.155672
R20971 output.n92 output.n91 0.155672
R20972 output.n139 output.n111 0.155672
R20973 output.n132 output.n111 0.155672
R20974 output.n132 output.n131 0.155672
R20975 output.n131 output.n115 0.155672
R20976 output.n124 output.n115 0.155672
R20977 output.n124 output.n123 0.155672
R20978 output output.n14 0.126227
R20979 plus.n27 plus.t19 436.949
R20980 plus.n5 plus.t11 436.949
R20981 plus.n28 plus.t5 415.966
R20982 plus.n30 plus.t17 415.966
R20983 plus.n34 plus.t20 415.966
R20984 plus.n35 plus.t10 415.966
R20985 plus.n23 plus.t6 415.966
R20986 plus.n41 plus.t9 415.966
R20987 plus.n42 plus.t16 415.966
R20988 plus.n20 plus.t7 415.966
R20989 plus.n19 plus.t15 415.966
R20990 plus.n1 plus.t12 415.966
R20991 plus.n13 plus.t18 415.966
R20992 plus.n12 plus.t14 415.966
R20993 plus.n4 plus.t8 415.966
R20994 plus.n6 plus.t13 415.966
R20995 plus.n46 plus.t4 243.97
R20996 plus.n46 plus.n45 223.454
R20997 plus.n48 plus.n47 223.454
R20998 plus.n43 plus.n42 161.3
R20999 plus.n41 plus.n22 161.3
R21000 plus.n40 plus.n39 161.3
R21001 plus.n38 plus.n23 161.3
R21002 plus.n37 plus.n36 161.3
R21003 plus.n35 plus.n24 161.3
R21004 plus.n34 plus.n33 161.3
R21005 plus.n32 plus.n25 161.3
R21006 plus.n31 plus.n30 161.3
R21007 plus.n29 plus.n26 161.3
R21008 plus.n8 plus.n7 161.3
R21009 plus.n9 plus.n4 161.3
R21010 plus.n11 plus.n10 161.3
R21011 plus.n12 plus.n3 161.3
R21012 plus.n13 plus.n2 161.3
R21013 plus.n15 plus.n14 161.3
R21014 plus.n16 plus.n1 161.3
R21015 plus.n18 plus.n17 161.3
R21016 plus.n19 plus.n0 161.3
R21017 plus.n21 plus.n20 161.3
R21018 plus.n27 plus.n26 70.4033
R21019 plus.n8 plus.n5 70.4033
R21020 plus.n35 plus.n34 48.2005
R21021 plus.n42 plus.n41 48.2005
R21022 plus.n20 plus.n19 48.2005
R21023 plus.n13 plus.n12 48.2005
R21024 plus.n30 plus.n29 37.246
R21025 plus.n40 plus.n23 37.246
R21026 plus.n18 plus.n1 37.246
R21027 plus.n7 plus.n4 37.246
R21028 plus.n30 plus.n25 35.7853
R21029 plus.n36 plus.n23 35.7853
R21030 plus.n14 plus.n1 35.7853
R21031 plus.n11 plus.n4 35.7853
R21032 plus.n44 plus.n43 28.5744
R21033 plus.n28 plus.n27 20.9576
R21034 plus.n6 plus.n5 20.9576
R21035 plus.n45 plus.t0 19.8005
R21036 plus.n45 plus.t1 19.8005
R21037 plus.n47 plus.t3 19.8005
R21038 plus.n47 plus.t2 19.8005
R21039 plus plus.n49 14.2034
R21040 plus.n34 plus.n25 12.4157
R21041 plus.n36 plus.n35 12.4157
R21042 plus.n14 plus.n13 12.4157
R21043 plus.n12 plus.n11 12.4157
R21044 plus.n44 plus.n21 11.76
R21045 plus.n29 plus.n28 10.955
R21046 plus.n41 plus.n40 10.955
R21047 plus.n19 plus.n18 10.955
R21048 plus.n7 plus.n6 10.955
R21049 plus.n49 plus.n48 5.40567
R21050 plus.n49 plus.n44 1.188
R21051 plus.n48 plus.n46 0.716017
R21052 plus.n31 plus.n26 0.189894
R21053 plus.n32 plus.n31 0.189894
R21054 plus.n33 plus.n32 0.189894
R21055 plus.n33 plus.n24 0.189894
R21056 plus.n37 plus.n24 0.189894
R21057 plus.n38 plus.n37 0.189894
R21058 plus.n39 plus.n38 0.189894
R21059 plus.n39 plus.n22 0.189894
R21060 plus.n43 plus.n22 0.189894
R21061 plus.n21 plus.n0 0.189894
R21062 plus.n17 plus.n0 0.189894
R21063 plus.n17 plus.n16 0.189894
R21064 plus.n16 plus.n15 0.189894
R21065 plus.n15 plus.n2 0.189894
R21066 plus.n3 plus.n2 0.189894
R21067 plus.n10 plus.n3 0.189894
R21068 plus.n10 plus.n9 0.189894
R21069 plus.n9 plus.n8 0.189894
R21070 a_n2903_n3924.n10 a_n2903_n3924.t21 214.994
R21071 a_n2903_n3924.n0 a_n2903_n3924.t16 214.975
R21072 a_n2903_n3924.n0 a_n2903_n3924.t18 214.321
R21073 a_n2903_n3924.n11 a_n2903_n3924.t19 214.321
R21074 a_n2903_n3924.n12 a_n2903_n3924.t22 214.321
R21075 a_n2903_n3924.n13 a_n2903_n3924.t17 214.321
R21076 a_n2903_n3924.n14 a_n2903_n3924.t20 214.321
R21077 a_n2903_n3924.n10 a_n2903_n3924.t39 214.321
R21078 a_n2903_n3924.n1 a_n2903_n3924.t1 55.8337
R21079 a_n2903_n3924.n2 a_n2903_n3924.t36 55.8337
R21080 a_n2903_n3924.n9 a_n2903_n3924.t28 55.8337
R21081 a_n2903_n3924.n34 a_n2903_n3924.t4 55.8335
R21082 a_n2903_n3924.n32 a_n2903_n3924.t25 55.8335
R21083 a_n2903_n3924.n25 a_n2903_n3924.t34 55.8335
R21084 a_n2903_n3924.n24 a_n2903_n3924.t9 55.8335
R21085 a_n2903_n3924.n17 a_n2903_n3924.t13 55.8335
R21086 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R21087 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R21088 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R21089 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R21090 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R21091 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R21092 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R21093 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R21094 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R21095 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R21096 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R21097 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R21098 a_n2903_n3924.n16 a_n2903_n3924.n9 12.1555
R21099 a_n2903_n3924.n34 a_n2903_n3924.n33 12.1555
R21100 a_n2903_n3924.n17 a_n2903_n3924.n16 5.07593
R21101 a_n2903_n3924.n33 a_n2903_n3924.n32 5.07593
R21102 a_n2903_n3924.n35 a_n2903_n3924.t14 2.82907
R21103 a_n2903_n3924.n35 a_n2903_n3924.t11 2.82907
R21104 a_n2903_n3924.n37 a_n2903_n3924.t0 2.82907
R21105 a_n2903_n3924.n37 a_n2903_n3924.t10 2.82907
R21106 a_n2903_n3924.n3 a_n2903_n3924.t37 2.82907
R21107 a_n2903_n3924.n3 a_n2903_n3924.t38 2.82907
R21108 a_n2903_n3924.n5 a_n2903_n3924.t32 2.82907
R21109 a_n2903_n3924.n5 a_n2903_n3924.t24 2.82907
R21110 a_n2903_n3924.n7 a_n2903_n3924.t27 2.82907
R21111 a_n2903_n3924.n7 a_n2903_n3924.t26 2.82907
R21112 a_n2903_n3924.n30 a_n2903_n3924.t30 2.82907
R21113 a_n2903_n3924.n30 a_n2903_n3924.t29 2.82907
R21114 a_n2903_n3924.n28 a_n2903_n3924.t33 2.82907
R21115 a_n2903_n3924.n28 a_n2903_n3924.t35 2.82907
R21116 a_n2903_n3924.n26 a_n2903_n3924.t31 2.82907
R21117 a_n2903_n3924.n26 a_n2903_n3924.t23 2.82907
R21118 a_n2903_n3924.n22 a_n2903_n3924.t12 2.82907
R21119 a_n2903_n3924.n22 a_n2903_n3924.t7 2.82907
R21120 a_n2903_n3924.n20 a_n2903_n3924.t2 2.82907
R21121 a_n2903_n3924.n20 a_n2903_n3924.t6 2.82907
R21122 a_n2903_n3924.n18 a_n2903_n3924.t5 2.82907
R21123 a_n2903_n3924.n18 a_n2903_n3924.t8 2.82907
R21124 a_n2903_n3924.t15 a_n2903_n3924.n40 2.82907
R21125 a_n2903_n3924.n40 a_n2903_n3924.t3 2.82907
R21126 a_n2903_n3924.n33 a_n2903_n3924.n0 1.95694
R21127 a_n2903_n3924.n16 a_n2903_n3924.n15 1.95694
R21128 a_n2903_n3924.n11 a_n2903_n3924.n0 0.69018
R21129 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R21130 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R21131 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R21132 a_n2903_n3924.n15 a_n2903_n3924.n10 0.511401
R21133 a_n2903_n3924.n19 a_n2903_n3924.n17 0.358259
R21134 a_n2903_n3924.n21 a_n2903_n3924.n19 0.358259
R21135 a_n2903_n3924.n23 a_n2903_n3924.n21 0.358259
R21136 a_n2903_n3924.n24 a_n2903_n3924.n23 0.358259
R21137 a_n2903_n3924.n27 a_n2903_n3924.n25 0.358259
R21138 a_n2903_n3924.n29 a_n2903_n3924.n27 0.358259
R21139 a_n2903_n3924.n31 a_n2903_n3924.n29 0.358259
R21140 a_n2903_n3924.n32 a_n2903_n3924.n31 0.358259
R21141 a_n2903_n3924.n9 a_n2903_n3924.n8 0.358259
R21142 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R21143 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R21144 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R21145 a_n2903_n3924.n39 a_n2903_n3924.n1 0.358259
R21146 a_n2903_n3924.n39 a_n2903_n3924.n38 0.358259
R21147 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R21148 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R21149 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R21150 a_n2903_n3924.n2 a_n2903_n3924.n1 0.235414
R21151 a_n2903_n3924.n15 a_n2903_n3924.n14 0.16111
R21152 outputibias.n27 outputibias.n1 289.615
R21153 outputibias.n58 outputibias.n32 289.615
R21154 outputibias.n90 outputibias.n64 289.615
R21155 outputibias.n122 outputibias.n96 289.615
R21156 outputibias.n28 outputibias.n27 185
R21157 outputibias.n26 outputibias.n25 185
R21158 outputibias.n5 outputibias.n4 185
R21159 outputibias.n20 outputibias.n19 185
R21160 outputibias.n18 outputibias.n17 185
R21161 outputibias.n9 outputibias.n8 185
R21162 outputibias.n12 outputibias.n11 185
R21163 outputibias.n59 outputibias.n58 185
R21164 outputibias.n57 outputibias.n56 185
R21165 outputibias.n36 outputibias.n35 185
R21166 outputibias.n51 outputibias.n50 185
R21167 outputibias.n49 outputibias.n48 185
R21168 outputibias.n40 outputibias.n39 185
R21169 outputibias.n43 outputibias.n42 185
R21170 outputibias.n91 outputibias.n90 185
R21171 outputibias.n89 outputibias.n88 185
R21172 outputibias.n68 outputibias.n67 185
R21173 outputibias.n83 outputibias.n82 185
R21174 outputibias.n81 outputibias.n80 185
R21175 outputibias.n72 outputibias.n71 185
R21176 outputibias.n75 outputibias.n74 185
R21177 outputibias.n123 outputibias.n122 185
R21178 outputibias.n121 outputibias.n120 185
R21179 outputibias.n100 outputibias.n99 185
R21180 outputibias.n115 outputibias.n114 185
R21181 outputibias.n113 outputibias.n112 185
R21182 outputibias.n104 outputibias.n103 185
R21183 outputibias.n107 outputibias.n106 185
R21184 outputibias.n0 outputibias.t8 178.945
R21185 outputibias.n133 outputibias.t9 177.018
R21186 outputibias.n132 outputibias.t10 177.018
R21187 outputibias.n0 outputibias.t11 177.018
R21188 outputibias.t7 outputibias.n10 147.661
R21189 outputibias.t5 outputibias.n41 147.661
R21190 outputibias.t1 outputibias.n73 147.661
R21191 outputibias.t3 outputibias.n105 147.661
R21192 outputibias.n128 outputibias.t6 132.363
R21193 outputibias.n128 outputibias.t4 130.436
R21194 outputibias.n129 outputibias.t0 130.436
R21195 outputibias.n130 outputibias.t2 130.436
R21196 outputibias.n27 outputibias.n26 104.615
R21197 outputibias.n26 outputibias.n4 104.615
R21198 outputibias.n19 outputibias.n4 104.615
R21199 outputibias.n19 outputibias.n18 104.615
R21200 outputibias.n18 outputibias.n8 104.615
R21201 outputibias.n11 outputibias.n8 104.615
R21202 outputibias.n58 outputibias.n57 104.615
R21203 outputibias.n57 outputibias.n35 104.615
R21204 outputibias.n50 outputibias.n35 104.615
R21205 outputibias.n50 outputibias.n49 104.615
R21206 outputibias.n49 outputibias.n39 104.615
R21207 outputibias.n42 outputibias.n39 104.615
R21208 outputibias.n90 outputibias.n89 104.615
R21209 outputibias.n89 outputibias.n67 104.615
R21210 outputibias.n82 outputibias.n67 104.615
R21211 outputibias.n82 outputibias.n81 104.615
R21212 outputibias.n81 outputibias.n71 104.615
R21213 outputibias.n74 outputibias.n71 104.615
R21214 outputibias.n122 outputibias.n121 104.615
R21215 outputibias.n121 outputibias.n99 104.615
R21216 outputibias.n114 outputibias.n99 104.615
R21217 outputibias.n114 outputibias.n113 104.615
R21218 outputibias.n113 outputibias.n103 104.615
R21219 outputibias.n106 outputibias.n103 104.615
R21220 outputibias.n63 outputibias.n31 95.6354
R21221 outputibias.n63 outputibias.n62 94.6732
R21222 outputibias.n95 outputibias.n94 94.6732
R21223 outputibias.n127 outputibias.n126 94.6732
R21224 outputibias.n11 outputibias.t7 52.3082
R21225 outputibias.n42 outputibias.t5 52.3082
R21226 outputibias.n74 outputibias.t1 52.3082
R21227 outputibias.n106 outputibias.t3 52.3082
R21228 outputibias.n12 outputibias.n10 15.6674
R21229 outputibias.n43 outputibias.n41 15.6674
R21230 outputibias.n75 outputibias.n73 15.6674
R21231 outputibias.n107 outputibias.n105 15.6674
R21232 outputibias.n13 outputibias.n9 12.8005
R21233 outputibias.n44 outputibias.n40 12.8005
R21234 outputibias.n76 outputibias.n72 12.8005
R21235 outputibias.n108 outputibias.n104 12.8005
R21236 outputibias.n17 outputibias.n16 12.0247
R21237 outputibias.n48 outputibias.n47 12.0247
R21238 outputibias.n80 outputibias.n79 12.0247
R21239 outputibias.n112 outputibias.n111 12.0247
R21240 outputibias.n20 outputibias.n7 11.249
R21241 outputibias.n51 outputibias.n38 11.249
R21242 outputibias.n83 outputibias.n70 11.249
R21243 outputibias.n115 outputibias.n102 11.249
R21244 outputibias.n21 outputibias.n5 10.4732
R21245 outputibias.n52 outputibias.n36 10.4732
R21246 outputibias.n84 outputibias.n68 10.4732
R21247 outputibias.n116 outputibias.n100 10.4732
R21248 outputibias.n25 outputibias.n24 9.69747
R21249 outputibias.n56 outputibias.n55 9.69747
R21250 outputibias.n88 outputibias.n87 9.69747
R21251 outputibias.n120 outputibias.n119 9.69747
R21252 outputibias.n31 outputibias.n30 9.45567
R21253 outputibias.n62 outputibias.n61 9.45567
R21254 outputibias.n94 outputibias.n93 9.45567
R21255 outputibias.n126 outputibias.n125 9.45567
R21256 outputibias.n30 outputibias.n29 9.3005
R21257 outputibias.n3 outputibias.n2 9.3005
R21258 outputibias.n24 outputibias.n23 9.3005
R21259 outputibias.n22 outputibias.n21 9.3005
R21260 outputibias.n7 outputibias.n6 9.3005
R21261 outputibias.n16 outputibias.n15 9.3005
R21262 outputibias.n14 outputibias.n13 9.3005
R21263 outputibias.n61 outputibias.n60 9.3005
R21264 outputibias.n34 outputibias.n33 9.3005
R21265 outputibias.n55 outputibias.n54 9.3005
R21266 outputibias.n53 outputibias.n52 9.3005
R21267 outputibias.n38 outputibias.n37 9.3005
R21268 outputibias.n47 outputibias.n46 9.3005
R21269 outputibias.n45 outputibias.n44 9.3005
R21270 outputibias.n93 outputibias.n92 9.3005
R21271 outputibias.n66 outputibias.n65 9.3005
R21272 outputibias.n87 outputibias.n86 9.3005
R21273 outputibias.n85 outputibias.n84 9.3005
R21274 outputibias.n70 outputibias.n69 9.3005
R21275 outputibias.n79 outputibias.n78 9.3005
R21276 outputibias.n77 outputibias.n76 9.3005
R21277 outputibias.n125 outputibias.n124 9.3005
R21278 outputibias.n98 outputibias.n97 9.3005
R21279 outputibias.n119 outputibias.n118 9.3005
R21280 outputibias.n117 outputibias.n116 9.3005
R21281 outputibias.n102 outputibias.n101 9.3005
R21282 outputibias.n111 outputibias.n110 9.3005
R21283 outputibias.n109 outputibias.n108 9.3005
R21284 outputibias.n28 outputibias.n3 8.92171
R21285 outputibias.n59 outputibias.n34 8.92171
R21286 outputibias.n91 outputibias.n66 8.92171
R21287 outputibias.n123 outputibias.n98 8.92171
R21288 outputibias.n29 outputibias.n1 8.14595
R21289 outputibias.n60 outputibias.n32 8.14595
R21290 outputibias.n92 outputibias.n64 8.14595
R21291 outputibias.n124 outputibias.n96 8.14595
R21292 outputibias.n31 outputibias.n1 5.81868
R21293 outputibias.n62 outputibias.n32 5.81868
R21294 outputibias.n94 outputibias.n64 5.81868
R21295 outputibias.n126 outputibias.n96 5.81868
R21296 outputibias.n131 outputibias.n130 5.20947
R21297 outputibias.n29 outputibias.n28 5.04292
R21298 outputibias.n60 outputibias.n59 5.04292
R21299 outputibias.n92 outputibias.n91 5.04292
R21300 outputibias.n124 outputibias.n123 5.04292
R21301 outputibias.n131 outputibias.n127 4.42209
R21302 outputibias.n14 outputibias.n10 4.38594
R21303 outputibias.n45 outputibias.n41 4.38594
R21304 outputibias.n77 outputibias.n73 4.38594
R21305 outputibias.n109 outputibias.n105 4.38594
R21306 outputibias.n132 outputibias.n131 4.28454
R21307 outputibias.n25 outputibias.n3 4.26717
R21308 outputibias.n56 outputibias.n34 4.26717
R21309 outputibias.n88 outputibias.n66 4.26717
R21310 outputibias.n120 outputibias.n98 4.26717
R21311 outputibias.n24 outputibias.n5 3.49141
R21312 outputibias.n55 outputibias.n36 3.49141
R21313 outputibias.n87 outputibias.n68 3.49141
R21314 outputibias.n119 outputibias.n100 3.49141
R21315 outputibias.n21 outputibias.n20 2.71565
R21316 outputibias.n52 outputibias.n51 2.71565
R21317 outputibias.n84 outputibias.n83 2.71565
R21318 outputibias.n116 outputibias.n115 2.71565
R21319 outputibias.n17 outputibias.n7 1.93989
R21320 outputibias.n48 outputibias.n38 1.93989
R21321 outputibias.n80 outputibias.n70 1.93989
R21322 outputibias.n112 outputibias.n102 1.93989
R21323 outputibias.n130 outputibias.n129 1.9266
R21324 outputibias.n129 outputibias.n128 1.9266
R21325 outputibias.n133 outputibias.n132 1.92658
R21326 outputibias.n134 outputibias.n133 1.29913
R21327 outputibias.n16 outputibias.n9 1.16414
R21328 outputibias.n47 outputibias.n40 1.16414
R21329 outputibias.n79 outputibias.n72 1.16414
R21330 outputibias.n111 outputibias.n104 1.16414
R21331 outputibias.n127 outputibias.n95 0.962709
R21332 outputibias.n95 outputibias.n63 0.962709
R21333 outputibias.n13 outputibias.n12 0.388379
R21334 outputibias.n44 outputibias.n43 0.388379
R21335 outputibias.n76 outputibias.n75 0.388379
R21336 outputibias.n108 outputibias.n107 0.388379
R21337 outputibias.n134 outputibias.n0 0.337251
R21338 outputibias outputibias.n134 0.302375
R21339 outputibias.n30 outputibias.n2 0.155672
R21340 outputibias.n23 outputibias.n2 0.155672
R21341 outputibias.n23 outputibias.n22 0.155672
R21342 outputibias.n22 outputibias.n6 0.155672
R21343 outputibias.n15 outputibias.n6 0.155672
R21344 outputibias.n15 outputibias.n14 0.155672
R21345 outputibias.n61 outputibias.n33 0.155672
R21346 outputibias.n54 outputibias.n33 0.155672
R21347 outputibias.n54 outputibias.n53 0.155672
R21348 outputibias.n53 outputibias.n37 0.155672
R21349 outputibias.n46 outputibias.n37 0.155672
R21350 outputibias.n46 outputibias.n45 0.155672
R21351 outputibias.n93 outputibias.n65 0.155672
R21352 outputibias.n86 outputibias.n65 0.155672
R21353 outputibias.n86 outputibias.n85 0.155672
R21354 outputibias.n85 outputibias.n69 0.155672
R21355 outputibias.n78 outputibias.n69 0.155672
R21356 outputibias.n78 outputibias.n77 0.155672
R21357 outputibias.n125 outputibias.n97 0.155672
R21358 outputibias.n118 outputibias.n97 0.155672
R21359 outputibias.n118 outputibias.n117 0.155672
R21360 outputibias.n117 outputibias.n101 0.155672
R21361 outputibias.n110 outputibias.n101 0.155672
R21362 outputibias.n110 outputibias.n109 0.155672
R21363 minus.n27 minus.t20 436.949
R21364 minus.n5 minus.t11 436.949
R21365 minus.n42 minus.t17 415.966
R21366 minus.n41 minus.t10 415.966
R21367 minus.n23 minus.t5 415.966
R21368 minus.n35 minus.t13 415.966
R21369 minus.n34 minus.t9 415.966
R21370 minus.n26 minus.t19 415.966
R21371 minus.n28 minus.t7 415.966
R21372 minus.n6 minus.t14 415.966
R21373 minus.n8 minus.t8 415.966
R21374 minus.n12 minus.t12 415.966
R21375 minus.n13 minus.t18 415.966
R21376 minus.n1 minus.t15 415.966
R21377 minus.n19 minus.t16 415.966
R21378 minus.n20 minus.t6 415.966
R21379 minus.n48 minus.t1 243.255
R21380 minus.n47 minus.n45 224.169
R21381 minus.n47 minus.n46 223.454
R21382 minus.n30 minus.n29 161.3
R21383 minus.n31 minus.n26 161.3
R21384 minus.n33 minus.n32 161.3
R21385 minus.n34 minus.n25 161.3
R21386 minus.n35 minus.n24 161.3
R21387 minus.n37 minus.n36 161.3
R21388 minus.n38 minus.n23 161.3
R21389 minus.n40 minus.n39 161.3
R21390 minus.n41 minus.n22 161.3
R21391 minus.n43 minus.n42 161.3
R21392 minus.n21 minus.n20 161.3
R21393 minus.n19 minus.n0 161.3
R21394 minus.n18 minus.n17 161.3
R21395 minus.n16 minus.n1 161.3
R21396 minus.n15 minus.n14 161.3
R21397 minus.n13 minus.n2 161.3
R21398 minus.n12 minus.n11 161.3
R21399 minus.n10 minus.n3 161.3
R21400 minus.n9 minus.n8 161.3
R21401 minus.n7 minus.n4 161.3
R21402 minus.n30 minus.n27 70.4033
R21403 minus.n5 minus.n4 70.4033
R21404 minus.n42 minus.n41 48.2005
R21405 minus.n35 minus.n34 48.2005
R21406 minus.n13 minus.n12 48.2005
R21407 minus.n20 minus.n19 48.2005
R21408 minus.n40 minus.n23 37.246
R21409 minus.n29 minus.n26 37.246
R21410 minus.n8 minus.n7 37.246
R21411 minus.n18 minus.n1 37.246
R21412 minus.n36 minus.n23 35.7853
R21413 minus.n33 minus.n26 35.7853
R21414 minus.n8 minus.n3 35.7853
R21415 minus.n14 minus.n1 35.7853
R21416 minus.n44 minus.n43 28.7903
R21417 minus.n28 minus.n27 20.9576
R21418 minus.n6 minus.n5 20.9576
R21419 minus.n46 minus.t3 19.8005
R21420 minus.n46 minus.t4 19.8005
R21421 minus.n45 minus.t2 19.8005
R21422 minus.n45 minus.t0 19.8005
R21423 minus.n36 minus.n35 12.4157
R21424 minus.n34 minus.n33 12.4157
R21425 minus.n12 minus.n3 12.4157
R21426 minus.n14 minus.n13 12.4157
R21427 minus.n44 minus.n21 11.9759
R21428 minus minus.n49 11.7812
R21429 minus.n41 minus.n40 10.955
R21430 minus.n29 minus.n28 10.955
R21431 minus.n7 minus.n6 10.955
R21432 minus.n19 minus.n18 10.955
R21433 minus.n49 minus.n48 4.80222
R21434 minus.n49 minus.n44 0.972091
R21435 minus.n48 minus.n47 0.716017
R21436 minus.n43 minus.n22 0.189894
R21437 minus.n39 minus.n22 0.189894
R21438 minus.n39 minus.n38 0.189894
R21439 minus.n38 minus.n37 0.189894
R21440 minus.n37 minus.n24 0.189894
R21441 minus.n25 minus.n24 0.189894
R21442 minus.n32 minus.n25 0.189894
R21443 minus.n32 minus.n31 0.189894
R21444 minus.n31 minus.n30 0.189894
R21445 minus.n9 minus.n4 0.189894
R21446 minus.n10 minus.n9 0.189894
R21447 minus.n11 minus.n10 0.189894
R21448 minus.n11 minus.n2 0.189894
R21449 minus.n15 minus.n2 0.189894
R21450 minus.n16 minus.n15 0.189894
R21451 minus.n17 minus.n16 0.189894
R21452 minus.n17 minus.n0 0.189894
R21453 minus.n21 minus.n0 0.189894
R21454 diffpairibias.n0 diffpairibias.t18 436.822
R21455 diffpairibias.n21 diffpairibias.t19 435.479
R21456 diffpairibias.n20 diffpairibias.t16 435.479
R21457 diffpairibias.n19 diffpairibias.t17 435.479
R21458 diffpairibias.n18 diffpairibias.t21 435.479
R21459 diffpairibias.n0 diffpairibias.t22 435.479
R21460 diffpairibias.n1 diffpairibias.t20 435.479
R21461 diffpairibias.n2 diffpairibias.t23 435.479
R21462 diffpairibias.n10 diffpairibias.t0 377.536
R21463 diffpairibias.n10 diffpairibias.t8 376.193
R21464 diffpairibias.n11 diffpairibias.t10 376.193
R21465 diffpairibias.n12 diffpairibias.t6 376.193
R21466 diffpairibias.n13 diffpairibias.t2 376.193
R21467 diffpairibias.n14 diffpairibias.t12 376.193
R21468 diffpairibias.n15 diffpairibias.t4 376.193
R21469 diffpairibias.n16 diffpairibias.t14 376.193
R21470 diffpairibias.n3 diffpairibias.t1 113.368
R21471 diffpairibias.n3 diffpairibias.t9 112.698
R21472 diffpairibias.n4 diffpairibias.t11 112.698
R21473 diffpairibias.n5 diffpairibias.t7 112.698
R21474 diffpairibias.n6 diffpairibias.t3 112.698
R21475 diffpairibias.n7 diffpairibias.t13 112.698
R21476 diffpairibias.n8 diffpairibias.t5 112.698
R21477 diffpairibias.n9 diffpairibias.t15 112.698
R21478 diffpairibias.n17 diffpairibias.n16 4.77242
R21479 diffpairibias.n17 diffpairibias.n9 4.30807
R21480 diffpairibias.n18 diffpairibias.n17 4.13945
R21481 diffpairibias.n16 diffpairibias.n15 1.34352
R21482 diffpairibias.n15 diffpairibias.n14 1.34352
R21483 diffpairibias.n14 diffpairibias.n13 1.34352
R21484 diffpairibias.n13 diffpairibias.n12 1.34352
R21485 diffpairibias.n12 diffpairibias.n11 1.34352
R21486 diffpairibias.n11 diffpairibias.n10 1.34352
R21487 diffpairibias.n2 diffpairibias.n1 1.34352
R21488 diffpairibias.n1 diffpairibias.n0 1.34352
R21489 diffpairibias.n19 diffpairibias.n18 1.34352
R21490 diffpairibias.n20 diffpairibias.n19 1.34352
R21491 diffpairibias.n21 diffpairibias.n20 1.34352
R21492 diffpairibias.n22 diffpairibias.n21 0.862419
R21493 diffpairibias diffpairibias.n22 0.684875
R21494 diffpairibias.n9 diffpairibias.n8 0.672012
R21495 diffpairibias.n8 diffpairibias.n7 0.672012
R21496 diffpairibias.n7 diffpairibias.n6 0.672012
R21497 diffpairibias.n6 diffpairibias.n5 0.672012
R21498 diffpairibias.n5 diffpairibias.n4 0.672012
R21499 diffpairibias.n4 diffpairibias.n3 0.672012
R21500 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus commonsourceibias 0.314643f
C1 plus commonsourceibias 0.268404f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13571f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 91.981f
C7 minus diffpairibias 1.62e-19
C8 commonsourceibias output 0.006808f
C9 vdd plus 0.069331f
C10 CSoutput minus 2.95655f
C11 plus diffpairibias 2.39e-19
C12 commonsourceibias outputibias 0.003832f
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.829163f
C15 commonsourceibias diffpairibias 0.052851f
C16 CSoutput commonsourceibias 36.982002f
C17 minus plus 8.5425f
C18 diffpairibias gnd 48.96824f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150147p
C22 plus gnd 28.85172f
C23 minus gnd 25.2504f
C24 CSoutput gnd 0.101655p
C25 vdd gnd 0.377288p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031083f
C74 minus.t15 gnd 0.314031f
C75 minus.n1 gnd 0.145186f
C76 minus.n2 gnd 0.031083f
C77 minus.n3 gnd 0.007053f
C78 minus.n4 gnd 0.098964f
C79 minus.t11 gnd 0.320848f
C80 minus.n5 gnd 0.135338f
C81 minus.t14 gnd 0.314031f
C82 minus.n6 gnd 0.143366f
C83 minus.n7 gnd 0.007053f
C84 minus.t8 gnd 0.314031f
C85 minus.n8 gnd 0.145186f
C86 minus.n9 gnd 0.031083f
C87 minus.n10 gnd 0.031083f
C88 minus.n11 gnd 0.031083f
C89 minus.t12 gnd 0.314031f
C90 minus.n12 gnd 0.143557f
C91 minus.t18 gnd 0.314031f
C92 minus.n13 gnd 0.143557f
C93 minus.n14 gnd 0.007053f
C94 minus.n15 gnd 0.031083f
C95 minus.n16 gnd 0.031083f
C96 minus.n17 gnd 0.031083f
C97 minus.n18 gnd 0.007053f
C98 minus.t16 gnd 0.314031f
C99 minus.n19 gnd 0.143366f
C100 minus.t6 gnd 0.314031f
C101 minus.n20 gnd 0.141928f
C102 minus.n21 gnd 0.351353f
C103 minus.n22 gnd 0.031083f
C104 minus.t17 gnd 0.314031f
C105 minus.t10 gnd 0.314031f
C106 minus.t5 gnd 0.314031f
C107 minus.n23 gnd 0.145186f
C108 minus.n24 gnd 0.031083f
C109 minus.t13 gnd 0.314031f
C110 minus.t9 gnd 0.314031f
C111 minus.n25 gnd 0.031083f
C112 minus.t19 gnd 0.314031f
C113 minus.n26 gnd 0.145186f
C114 minus.t20 gnd 0.320848f
C115 minus.n27 gnd 0.135338f
C116 minus.t7 gnd 0.314031f
C117 minus.n28 gnd 0.143366f
C118 minus.n29 gnd 0.007053f
C119 minus.n30 gnd 0.098964f
C120 minus.n31 gnd 0.031083f
C121 minus.n32 gnd 0.031083f
C122 minus.n33 gnd 0.007053f
C123 minus.n34 gnd 0.143557f
C124 minus.n35 gnd 0.143557f
C125 minus.n36 gnd 0.007053f
C126 minus.n37 gnd 0.031083f
C127 minus.n38 gnd 0.031083f
C128 minus.n39 gnd 0.031083f
C129 minus.n40 gnd 0.007053f
C130 minus.n41 gnd 0.143366f
C131 minus.n42 gnd 0.141928f
C132 minus.n43 gnd 0.836604f
C133 minus.n44 gnd 1.28731f
C134 minus.t2 gnd 0.009582f
C135 minus.t0 gnd 0.009582f
C136 minus.n45 gnd 0.031508f
C137 minus.t3 gnd 0.009582f
C138 minus.t4 gnd 0.009582f
C139 minus.n46 gnd 0.031076f
C140 minus.n47 gnd 0.265222f
C141 minus.t1 gnd 0.053333f
C142 minus.n48 gnd 0.144729f
C143 minus.n49 gnd 2.11885f
C144 outputibias.t11 gnd 0.11477f
C145 outputibias.t8 gnd 0.115567f
C146 outputibias.n0 gnd 0.130108f
C147 outputibias.n1 gnd 0.001372f
C148 outputibias.n2 gnd 9.76e-19
C149 outputibias.n3 gnd 5.24e-19
C150 outputibias.n4 gnd 0.001239f
C151 outputibias.n5 gnd 5.55e-19
C152 outputibias.n6 gnd 9.76e-19
C153 outputibias.n7 gnd 5.24e-19
C154 outputibias.n8 gnd 0.001239f
C155 outputibias.n9 gnd 5.55e-19
C156 outputibias.n10 gnd 0.004176f
C157 outputibias.t7 gnd 0.00202f
C158 outputibias.n11 gnd 9.3e-19
C159 outputibias.n12 gnd 7.32e-19
C160 outputibias.n13 gnd 5.24e-19
C161 outputibias.n14 gnd 0.02322f
C162 outputibias.n15 gnd 9.76e-19
C163 outputibias.n16 gnd 5.24e-19
C164 outputibias.n17 gnd 5.55e-19
C165 outputibias.n18 gnd 0.001239f
C166 outputibias.n19 gnd 0.001239f
C167 outputibias.n20 gnd 5.55e-19
C168 outputibias.n21 gnd 5.24e-19
C169 outputibias.n22 gnd 9.76e-19
C170 outputibias.n23 gnd 9.76e-19
C171 outputibias.n24 gnd 5.24e-19
C172 outputibias.n25 gnd 5.55e-19
C173 outputibias.n26 gnd 0.001239f
C174 outputibias.n27 gnd 0.002683f
C175 outputibias.n28 gnd 5.55e-19
C176 outputibias.n29 gnd 5.24e-19
C177 outputibias.n30 gnd 0.002256f
C178 outputibias.n31 gnd 0.005781f
C179 outputibias.n32 gnd 0.001372f
C180 outputibias.n33 gnd 9.76e-19
C181 outputibias.n34 gnd 5.24e-19
C182 outputibias.n35 gnd 0.001239f
C183 outputibias.n36 gnd 5.55e-19
C184 outputibias.n37 gnd 9.76e-19
C185 outputibias.n38 gnd 5.24e-19
C186 outputibias.n39 gnd 0.001239f
C187 outputibias.n40 gnd 5.55e-19
C188 outputibias.n41 gnd 0.004176f
C189 outputibias.t5 gnd 0.00202f
C190 outputibias.n42 gnd 9.3e-19
C191 outputibias.n43 gnd 7.32e-19
C192 outputibias.n44 gnd 5.24e-19
C193 outputibias.n45 gnd 0.02322f
C194 outputibias.n46 gnd 9.76e-19
C195 outputibias.n47 gnd 5.24e-19
C196 outputibias.n48 gnd 5.55e-19
C197 outputibias.n49 gnd 0.001239f
C198 outputibias.n50 gnd 0.001239f
C199 outputibias.n51 gnd 5.55e-19
C200 outputibias.n52 gnd 5.24e-19
C201 outputibias.n53 gnd 9.76e-19
C202 outputibias.n54 gnd 9.76e-19
C203 outputibias.n55 gnd 5.24e-19
C204 outputibias.n56 gnd 5.55e-19
C205 outputibias.n57 gnd 0.001239f
C206 outputibias.n58 gnd 0.002683f
C207 outputibias.n59 gnd 5.55e-19
C208 outputibias.n60 gnd 5.24e-19
C209 outputibias.n61 gnd 0.002256f
C210 outputibias.n62 gnd 0.005197f
C211 outputibias.n63 gnd 0.121892f
C212 outputibias.n64 gnd 0.001372f
C213 outputibias.n65 gnd 9.76e-19
C214 outputibias.n66 gnd 5.24e-19
C215 outputibias.n67 gnd 0.001239f
C216 outputibias.n68 gnd 5.55e-19
C217 outputibias.n69 gnd 9.76e-19
C218 outputibias.n70 gnd 5.24e-19
C219 outputibias.n71 gnd 0.001239f
C220 outputibias.n72 gnd 5.55e-19
C221 outputibias.n73 gnd 0.004176f
C222 outputibias.t1 gnd 0.00202f
C223 outputibias.n74 gnd 9.3e-19
C224 outputibias.n75 gnd 7.32e-19
C225 outputibias.n76 gnd 5.24e-19
C226 outputibias.n77 gnd 0.02322f
C227 outputibias.n78 gnd 9.76e-19
C228 outputibias.n79 gnd 5.24e-19
C229 outputibias.n80 gnd 5.55e-19
C230 outputibias.n81 gnd 0.001239f
C231 outputibias.n82 gnd 0.001239f
C232 outputibias.n83 gnd 5.55e-19
C233 outputibias.n84 gnd 5.24e-19
C234 outputibias.n85 gnd 9.76e-19
C235 outputibias.n86 gnd 9.76e-19
C236 outputibias.n87 gnd 5.24e-19
C237 outputibias.n88 gnd 5.55e-19
C238 outputibias.n89 gnd 0.001239f
C239 outputibias.n90 gnd 0.002683f
C240 outputibias.n91 gnd 5.55e-19
C241 outputibias.n92 gnd 5.24e-19
C242 outputibias.n93 gnd 0.002256f
C243 outputibias.n94 gnd 0.005197f
C244 outputibias.n95 gnd 0.064513f
C245 outputibias.n96 gnd 0.001372f
C246 outputibias.n97 gnd 9.76e-19
C247 outputibias.n98 gnd 5.24e-19
C248 outputibias.n99 gnd 0.001239f
C249 outputibias.n100 gnd 5.55e-19
C250 outputibias.n101 gnd 9.76e-19
C251 outputibias.n102 gnd 5.24e-19
C252 outputibias.n103 gnd 0.001239f
C253 outputibias.n104 gnd 5.55e-19
C254 outputibias.n105 gnd 0.004176f
C255 outputibias.t3 gnd 0.00202f
C256 outputibias.n106 gnd 9.3e-19
C257 outputibias.n107 gnd 7.32e-19
C258 outputibias.n108 gnd 5.24e-19
C259 outputibias.n109 gnd 0.02322f
C260 outputibias.n110 gnd 9.76e-19
C261 outputibias.n111 gnd 5.24e-19
C262 outputibias.n112 gnd 5.55e-19
C263 outputibias.n113 gnd 0.001239f
C264 outputibias.n114 gnd 0.001239f
C265 outputibias.n115 gnd 5.55e-19
C266 outputibias.n116 gnd 5.24e-19
C267 outputibias.n117 gnd 9.76e-19
C268 outputibias.n118 gnd 9.76e-19
C269 outputibias.n119 gnd 5.24e-19
C270 outputibias.n120 gnd 5.55e-19
C271 outputibias.n121 gnd 0.001239f
C272 outputibias.n122 gnd 0.002683f
C273 outputibias.n123 gnd 5.55e-19
C274 outputibias.n124 gnd 5.24e-19
C275 outputibias.n125 gnd 0.002256f
C276 outputibias.n126 gnd 0.005197f
C277 outputibias.n127 gnd 0.084814f
C278 outputibias.t2 gnd 0.108319f
C279 outputibias.t0 gnd 0.108319f
C280 outputibias.t4 gnd 0.108319f
C281 outputibias.t6 gnd 0.109238f
C282 outputibias.n128 gnd 0.134674f
C283 outputibias.n129 gnd 0.07244f
C284 outputibias.n130 gnd 0.079818f
C285 outputibias.n131 gnd 0.164901f
C286 outputibias.t10 gnd 0.11477f
C287 outputibias.n132 gnd 0.067481f
C288 outputibias.t9 gnd 0.11477f
C289 outputibias.n133 gnd 0.065115f
C290 outputibias.n134 gnd 0.029159f
C291 a_n2903_n3924.n0 gnd 2.07284f
C292 a_n2903_n3924.t3 gnd 0.094832f
C293 a_n2903_n3924.t1 gnd 0.985605f
C294 a_n2903_n3924.n1 gnd 0.334506f
C295 a_n2903_n3924.t16 gnd 1.22783f
C296 a_n2903_n3924.t36 gnd 0.985605f
C297 a_n2903_n3924.n2 gnd 0.334506f
C298 a_n2903_n3924.t37 gnd 0.094832f
C299 a_n2903_n3924.t38 gnd 0.094832f
C300 a_n2903_n3924.n3 gnd 0.774508f
C301 a_n2903_n3924.n4 gnd 0.314114f
C302 a_n2903_n3924.t32 gnd 0.094832f
C303 a_n2903_n3924.t24 gnd 0.094832f
C304 a_n2903_n3924.n5 gnd 0.774508f
C305 a_n2903_n3924.n6 gnd 0.314114f
C306 a_n2903_n3924.t27 gnd 0.094832f
C307 a_n2903_n3924.t26 gnd 0.094832f
C308 a_n2903_n3924.n7 gnd 0.774508f
C309 a_n2903_n3924.n8 gnd 0.314114f
C310 a_n2903_n3924.t28 gnd 0.985605f
C311 a_n2903_n3924.n9 gnd 0.850542f
C312 a_n2903_n3924.t21 gnd 1.22634f
C313 a_n2903_n3924.t39 gnd 1.22459f
C314 a_n2903_n3924.n10 gnd 1.34231f
C315 a_n2903_n3924.t18 gnd 1.22459f
C316 a_n2903_n3924.t19 gnd 1.22459f
C317 a_n2903_n3924.n11 gnd 0.8625f
C318 a_n2903_n3924.t22 gnd 1.22459f
C319 a_n2903_n3924.n12 gnd 0.8625f
C320 a_n2903_n3924.t17 gnd 1.22459f
C321 a_n2903_n3924.n13 gnd 0.8625f
C322 a_n2903_n3924.t20 gnd 1.22459f
C323 a_n2903_n3924.n14 gnd 0.614303f
C324 a_n2903_n3924.n15 gnd 0.466167f
C325 a_n2903_n3924.n16 gnd 0.885261f
C326 a_n2903_n3924.t13 gnd 0.985601f
C327 a_n2903_n3924.n17 gnd 0.54064f
C328 a_n2903_n3924.t5 gnd 0.094832f
C329 a_n2903_n3924.t8 gnd 0.094832f
C330 a_n2903_n3924.n18 gnd 0.774507f
C331 a_n2903_n3924.n19 gnd 0.314115f
C332 a_n2903_n3924.t2 gnd 0.094832f
C333 a_n2903_n3924.t6 gnd 0.094832f
C334 a_n2903_n3924.n20 gnd 0.774507f
C335 a_n2903_n3924.n21 gnd 0.314115f
C336 a_n2903_n3924.t12 gnd 0.094832f
C337 a_n2903_n3924.t7 gnd 0.094832f
C338 a_n2903_n3924.n22 gnd 0.774507f
C339 a_n2903_n3924.n23 gnd 0.314115f
C340 a_n2903_n3924.t9 gnd 0.985601f
C341 a_n2903_n3924.n24 gnd 0.334509f
C342 a_n2903_n3924.t34 gnd 0.985601f
C343 a_n2903_n3924.n25 gnd 0.334509f
C344 a_n2903_n3924.t31 gnd 0.094832f
C345 a_n2903_n3924.t23 gnd 0.094832f
C346 a_n2903_n3924.n26 gnd 0.774507f
C347 a_n2903_n3924.n27 gnd 0.314115f
C348 a_n2903_n3924.t33 gnd 0.094832f
C349 a_n2903_n3924.t35 gnd 0.094832f
C350 a_n2903_n3924.n28 gnd 0.774507f
C351 a_n2903_n3924.n29 gnd 0.314115f
C352 a_n2903_n3924.t30 gnd 0.094832f
C353 a_n2903_n3924.t29 gnd 0.094832f
C354 a_n2903_n3924.n30 gnd 0.774507f
C355 a_n2903_n3924.n31 gnd 0.314115f
C356 a_n2903_n3924.t25 gnd 0.985601f
C357 a_n2903_n3924.n32 gnd 0.54064f
C358 a_n2903_n3924.n33 gnd 0.885261f
C359 a_n2903_n3924.t4 gnd 0.985601f
C360 a_n2903_n3924.n34 gnd 0.850545f
C361 a_n2903_n3924.t14 gnd 0.094832f
C362 a_n2903_n3924.t11 gnd 0.094832f
C363 a_n2903_n3924.n35 gnd 0.774508f
C364 a_n2903_n3924.n36 gnd 0.314114f
C365 a_n2903_n3924.t0 gnd 0.094832f
C366 a_n2903_n3924.t10 gnd 0.094832f
C367 a_n2903_n3924.n37 gnd 0.774508f
C368 a_n2903_n3924.n38 gnd 0.314114f
C369 a_n2903_n3924.n39 gnd 0.314113f
C370 a_n2903_n3924.n40 gnd 0.774509f
C371 a_n2903_n3924.t15 gnd 0.094832f
C372 plus.n0 gnd 0.022128f
C373 plus.t7 gnd 0.223557f
C374 plus.t15 gnd 0.223557f
C375 plus.t12 gnd 0.223557f
C376 plus.n1 gnd 0.103357f
C377 plus.n2 gnd 0.022128f
C378 plus.t18 gnd 0.223557f
C379 plus.n3 gnd 0.022128f
C380 plus.t14 gnd 0.223557f
C381 plus.t8 gnd 0.223557f
C382 plus.n4 gnd 0.103357f
C383 plus.t11 gnd 0.22841f
C384 plus.n5 gnd 0.096346f
C385 plus.t13 gnd 0.223557f
C386 plus.n6 gnd 0.102061f
C387 plus.n7 gnd 0.005021f
C388 plus.n8 gnd 0.070452f
C389 plus.n9 gnd 0.022128f
C390 plus.n10 gnd 0.022128f
C391 plus.n11 gnd 0.005021f
C392 plus.n12 gnd 0.102198f
C393 plus.n13 gnd 0.102198f
C394 plus.n14 gnd 0.005021f
C395 plus.n15 gnd 0.022128f
C396 plus.n16 gnd 0.022128f
C397 plus.n17 gnd 0.022128f
C398 plus.n18 gnd 0.005021f
C399 plus.n19 gnd 0.102061f
C400 plus.n20 gnd 0.101038f
C401 plus.n21 gnd 0.244413f
C402 plus.n22 gnd 0.022128f
C403 plus.t6 gnd 0.223557f
C404 plus.n23 gnd 0.103357f
C405 plus.n24 gnd 0.022128f
C406 plus.n25 gnd 0.005021f
C407 plus.t20 gnd 0.223557f
C408 plus.n26 gnd 0.070452f
C409 plus.t5 gnd 0.223557f
C410 plus.t19 gnd 0.22841f
C411 plus.n27 gnd 0.096346f
C412 plus.n28 gnd 0.102061f
C413 plus.n29 gnd 0.005021f
C414 plus.t17 gnd 0.223557f
C415 plus.n30 gnd 0.103357f
C416 plus.n31 gnd 0.022128f
C417 plus.n32 gnd 0.022128f
C418 plus.n33 gnd 0.022128f
C419 plus.n34 gnd 0.102198f
C420 plus.t10 gnd 0.223557f
C421 plus.n35 gnd 0.102198f
C422 plus.n36 gnd 0.005021f
C423 plus.n37 gnd 0.022128f
C424 plus.n38 gnd 0.022128f
C425 plus.n39 gnd 0.022128f
C426 plus.n40 gnd 0.005021f
C427 plus.t9 gnd 0.223557f
C428 plus.n41 gnd 0.102061f
C429 plus.t16 gnd 0.223557f
C430 plus.n42 gnd 0.101038f
C431 plus.n43 gnd 0.58668f
C432 plus.n44 gnd 0.907705f
C433 plus.t4 gnd 0.038199f
C434 plus.t0 gnd 0.006821f
C435 plus.t1 gnd 0.006821f
C436 plus.n45 gnd 0.022123f
C437 plus.n46 gnd 0.171743f
C438 plus.t3 gnd 0.006821f
C439 plus.t2 gnd 0.006821f
C440 plus.n47 gnd 0.022123f
C441 plus.n48 gnd 0.128914f
C442 plus.n49 gnd 2.34093f
C443 output.t16 gnd 0.464308f
C444 output.t5 gnd 0.044422f
C445 output.t10 gnd 0.044422f
C446 output.n0 gnd 0.364624f
C447 output.n1 gnd 0.614102f
C448 output.t14 gnd 0.044422f
C449 output.t6 gnd 0.044422f
C450 output.n2 gnd 0.364624f
C451 output.n3 gnd 0.350265f
C452 output.t9 gnd 0.044422f
C453 output.t7 gnd 0.044422f
C454 output.n4 gnd 0.364624f
C455 output.n5 gnd 0.350265f
C456 output.t13 gnd 0.044422f
C457 output.t15 gnd 0.044422f
C458 output.n6 gnd 0.364624f
C459 output.n7 gnd 0.350265f
C460 output.t18 gnd 0.044422f
C461 output.t11 gnd 0.044422f
C462 output.n8 gnd 0.364624f
C463 output.n9 gnd 0.350265f
C464 output.t12 gnd 0.044422f
C465 output.t3 gnd 0.044422f
C466 output.n10 gnd 0.364624f
C467 output.n11 gnd 0.350265f
C468 output.t4 gnd 0.044422f
C469 output.t8 gnd 0.044422f
C470 output.n12 gnd 0.364624f
C471 output.n13 gnd 0.350265f
C472 output.t17 gnd 0.462979f
C473 output.n14 gnd 0.28994f
C474 output.n15 gnd 0.015803f
C475 output.n16 gnd 0.011243f
C476 output.n17 gnd 0.006041f
C477 output.n18 gnd 0.01428f
C478 output.n19 gnd 0.006397f
C479 output.n20 gnd 0.011243f
C480 output.n21 gnd 0.006041f
C481 output.n22 gnd 0.01428f
C482 output.n23 gnd 0.006397f
C483 output.n24 gnd 0.048111f
C484 output.t0 gnd 0.023274f
C485 output.n25 gnd 0.01071f
C486 output.n26 gnd 0.008435f
C487 output.n27 gnd 0.006041f
C488 output.n28 gnd 0.267512f
C489 output.n29 gnd 0.011243f
C490 output.n30 gnd 0.006041f
C491 output.n31 gnd 0.006397f
C492 output.n32 gnd 0.01428f
C493 output.n33 gnd 0.01428f
C494 output.n34 gnd 0.006397f
C495 output.n35 gnd 0.006041f
C496 output.n36 gnd 0.011243f
C497 output.n37 gnd 0.011243f
C498 output.n38 gnd 0.006041f
C499 output.n39 gnd 0.006397f
C500 output.n40 gnd 0.01428f
C501 output.n41 gnd 0.030913f
C502 output.n42 gnd 0.006397f
C503 output.n43 gnd 0.006041f
C504 output.n44 gnd 0.025987f
C505 output.n45 gnd 0.097665f
C506 output.n46 gnd 0.015803f
C507 output.n47 gnd 0.011243f
C508 output.n48 gnd 0.006041f
C509 output.n49 gnd 0.01428f
C510 output.n50 gnd 0.006397f
C511 output.n51 gnd 0.011243f
C512 output.n52 gnd 0.006041f
C513 output.n53 gnd 0.01428f
C514 output.n54 gnd 0.006397f
C515 output.n55 gnd 0.048111f
C516 output.t19 gnd 0.023274f
C517 output.n56 gnd 0.01071f
C518 output.n57 gnd 0.008435f
C519 output.n58 gnd 0.006041f
C520 output.n59 gnd 0.267512f
C521 output.n60 gnd 0.011243f
C522 output.n61 gnd 0.006041f
C523 output.n62 gnd 0.006397f
C524 output.n63 gnd 0.01428f
C525 output.n64 gnd 0.01428f
C526 output.n65 gnd 0.006397f
C527 output.n66 gnd 0.006041f
C528 output.n67 gnd 0.011243f
C529 output.n68 gnd 0.011243f
C530 output.n69 gnd 0.006041f
C531 output.n70 gnd 0.006397f
C532 output.n71 gnd 0.01428f
C533 output.n72 gnd 0.030913f
C534 output.n73 gnd 0.006397f
C535 output.n74 gnd 0.006041f
C536 output.n75 gnd 0.025987f
C537 output.n76 gnd 0.09306f
C538 output.n77 gnd 1.65264f
C539 output.n78 gnd 0.015803f
C540 output.n79 gnd 0.011243f
C541 output.n80 gnd 0.006041f
C542 output.n81 gnd 0.01428f
C543 output.n82 gnd 0.006397f
C544 output.n83 gnd 0.011243f
C545 output.n84 gnd 0.006041f
C546 output.n85 gnd 0.01428f
C547 output.n86 gnd 0.006397f
C548 output.n87 gnd 0.048111f
C549 output.t2 gnd 0.023274f
C550 output.n88 gnd 0.01071f
C551 output.n89 gnd 0.008435f
C552 output.n90 gnd 0.006041f
C553 output.n91 gnd 0.267512f
C554 output.n92 gnd 0.011243f
C555 output.n93 gnd 0.006041f
C556 output.n94 gnd 0.006397f
C557 output.n95 gnd 0.01428f
C558 output.n96 gnd 0.01428f
C559 output.n97 gnd 0.006397f
C560 output.n98 gnd 0.006041f
C561 output.n99 gnd 0.011243f
C562 output.n100 gnd 0.011243f
C563 output.n101 gnd 0.006041f
C564 output.n102 gnd 0.006397f
C565 output.n103 gnd 0.01428f
C566 output.n104 gnd 0.030913f
C567 output.n105 gnd 0.006397f
C568 output.n106 gnd 0.006041f
C569 output.n107 gnd 0.025987f
C570 output.n108 gnd 0.09306f
C571 output.n109 gnd 0.713089f
C572 output.n110 gnd 0.015803f
C573 output.n111 gnd 0.011243f
C574 output.n112 gnd 0.006041f
C575 output.n113 gnd 0.01428f
C576 output.n114 gnd 0.006397f
C577 output.n115 gnd 0.011243f
C578 output.n116 gnd 0.006041f
C579 output.n117 gnd 0.01428f
C580 output.n118 gnd 0.006397f
C581 output.n119 gnd 0.048111f
C582 output.t1 gnd 0.023274f
C583 output.n120 gnd 0.01071f
C584 output.n121 gnd 0.008435f
C585 output.n122 gnd 0.006041f
C586 output.n123 gnd 0.267512f
C587 output.n124 gnd 0.011243f
C588 output.n125 gnd 0.006041f
C589 output.n126 gnd 0.006397f
C590 output.n127 gnd 0.01428f
C591 output.n128 gnd 0.01428f
C592 output.n129 gnd 0.006397f
C593 output.n130 gnd 0.006041f
C594 output.n131 gnd 0.011243f
C595 output.n132 gnd 0.011243f
C596 output.n133 gnd 0.006041f
C597 output.n134 gnd 0.006397f
C598 output.n135 gnd 0.01428f
C599 output.n136 gnd 0.030913f
C600 output.n137 gnd 0.006397f
C601 output.n138 gnd 0.006041f
C602 output.n139 gnd 0.025987f
C603 output.n140 gnd 0.09306f
C604 output.n141 gnd 1.67353f
C605 a_n1808_13878.t4 gnd 0.185195f
C606 a_n1808_13878.t0 gnd 0.185195f
C607 a_n1808_13878.t2 gnd 0.185195f
C608 a_n1808_13878.n0 gnd 1.4598f
C609 a_n1808_13878.t6 gnd 0.185195f
C610 a_n1808_13878.t1 gnd 0.185195f
C611 a_n1808_13878.n1 gnd 1.45825f
C612 a_n1808_13878.n2 gnd 2.03762f
C613 a_n1808_13878.t5 gnd 0.185195f
C614 a_n1808_13878.t9 gnd 0.185195f
C615 a_n1808_13878.n3 gnd 1.46067f
C616 a_n1808_13878.t10 gnd 0.185195f
C617 a_n1808_13878.t3 gnd 0.185195f
C618 a_n1808_13878.n4 gnd 1.45825f
C619 a_n1808_13878.n5 gnd 1.31079f
C620 a_n1808_13878.t7 gnd 0.185195f
C621 a_n1808_13878.t8 gnd 0.185195f
C622 a_n1808_13878.n6 gnd 1.45825f
C623 a_n1808_13878.n7 gnd 1.80025f
C624 a_n1808_13878.t13 gnd 1.73408f
C625 a_n1808_13878.t16 gnd 0.185195f
C626 a_n1808_13878.t17 gnd 0.185195f
C627 a_n1808_13878.n8 gnd 1.30452f
C628 a_n1808_13878.n9 gnd 1.4576f
C629 a_n1808_13878.t12 gnd 1.73062f
C630 a_n1808_13878.n10 gnd 0.733487f
C631 a_n1808_13878.t15 gnd 1.73062f
C632 a_n1808_13878.n11 gnd 0.733487f
C633 a_n1808_13878.t18 gnd 0.185195f
C634 a_n1808_13878.t19 gnd 0.185195f
C635 a_n1808_13878.n12 gnd 1.30452f
C636 a_n1808_13878.n13 gnd 0.74059f
C637 a_n1808_13878.t14 gnd 1.73062f
C638 a_n1808_13878.n14 gnd 1.7272f
C639 a_n1808_13878.n15 gnd 2.51438f
C640 a_n1808_13878.n16 gnd 3.69301f
C641 a_n1808_13878.n17 gnd 1.45826f
C642 a_n1808_13878.t11 gnd 0.185195f
C643 a_n1986_13878.n0 gnd 3.20192f
C644 a_n1986_13878.n1 gnd 0.64915f
C645 a_n1986_13878.n2 gnd 0.219304f
C646 a_n1986_13878.n3 gnd 0.286909f
C647 a_n1986_13878.n4 gnd 0.452885f
C648 a_n1986_13878.n5 gnd 0.674778f
C649 a_n1986_13878.n6 gnd 0.219304f
C650 a_n1986_13878.n7 gnd 0.286909f
C651 a_n1986_13878.n8 gnd 0.534226f
C652 a_n1986_13878.n9 gnd 0.208083f
C653 a_n1986_13878.n10 gnd 0.153257f
C654 a_n1986_13878.n11 gnd 0.240872f
C655 a_n1986_13878.n12 gnd 0.186046f
C656 a_n1986_13878.n13 gnd 0.208083f
C657 a_n1986_13878.n14 gnd 1.02197f
C658 a_n1986_13878.n15 gnd 0.153257f
C659 a_n1986_13878.n16 gnd 0.589052f
C660 a_n1986_13878.n17 gnd 0.439018f
C661 a_n1986_13878.n18 gnd 0.219304f
C662 a_n1986_13878.n19 gnd 0.500138f
C663 a_n1986_13878.n20 gnd 0.286909f
C664 a_n1986_13878.n21 gnd 0.445312f
C665 a_n1986_13878.n22 gnd 0.219304f
C666 a_n1986_13878.n23 gnd 0.742922f
C667 a_n1986_13878.n24 gnd 0.286909f
C668 a_n1986_13878.n25 gnd 1.19721f
C669 a_n1986_13878.n26 gnd 1.9455f
C670 a_n1986_13878.n27 gnd 1.1624f
C671 a_n1986_13878.n28 gnd 1.8055f
C672 a_n1986_13878.n29 gnd 2.46475f
C673 a_n1986_13878.n30 gnd 3.82161f
C674 a_n1986_13878.n31 gnd 3.20861f
C675 a_n1986_13878.n32 gnd 0.008491f
C676 a_n1986_13878.n34 gnd 0.290112f
C677 a_n1986_13878.n35 gnd 0.008491f
C678 a_n1986_13878.n37 gnd 0.290112f
C679 a_n1986_13878.n38 gnd 0.008491f
C680 a_n1986_13878.n39 gnd 0.2897f
C681 a_n1986_13878.n40 gnd 0.008491f
C682 a_n1986_13878.n41 gnd 0.2897f
C683 a_n1986_13878.n42 gnd 0.008491f
C684 a_n1986_13878.n43 gnd 0.2897f
C685 a_n1986_13878.n44 gnd 0.008491f
C686 a_n1986_13878.n45 gnd 0.2897f
C687 a_n1986_13878.n46 gnd 0.008491f
C688 a_n1986_13878.n48 gnd 0.290112f
C689 a_n1986_13878.n49 gnd 0.008491f
C690 a_n1986_13878.n51 gnd 0.290112f
C691 a_n1986_13878.t20 gnd 0.722451f
C692 a_n1986_13878.t2 gnd 0.707549f
C693 a_n1986_13878.t12 gnd 0.707549f
C694 a_n1986_13878.t18 gnd 0.707549f
C695 a_n1986_13878.n52 gnd 0.311083f
C696 a_n1986_13878.t8 gnd 0.707549f
C697 a_n1986_13878.t0 gnd 0.719248f
C698 a_n1986_13878.t67 gnd 0.722451f
C699 a_n1986_13878.t50 gnd 0.707549f
C700 a_n1986_13878.t54 gnd 0.707549f
C701 a_n1986_13878.t44 gnd 0.707549f
C702 a_n1986_13878.n53 gnd 0.311083f
C703 a_n1986_13878.t59 gnd 0.707549f
C704 a_n1986_13878.t65 gnd 0.719248f
C705 a_n1986_13878.t23 gnd 1.4243f
C706 a_n1986_13878.t17 gnd 0.152112f
C707 a_n1986_13878.t7 gnd 0.152112f
C708 a_n1986_13878.n54 gnd 1.07147f
C709 a_n1986_13878.t5 gnd 0.152112f
C710 a_n1986_13878.t15 gnd 0.152112f
C711 a_n1986_13878.n55 gnd 1.07147f
C712 a_n1986_13878.t11 gnd 1.42146f
C713 a_n1986_13878.t4 gnd 0.707549f
C714 a_n1986_13878.n56 gnd 0.311083f
C715 a_n1986_13878.t14 gnd 0.707549f
C716 a_n1986_13878.t16 gnd 0.707549f
C717 a_n1986_13878.t48 gnd 0.707549f
C718 a_n1986_13878.n57 gnd 0.311083f
C719 a_n1986_13878.t57 gnd 0.707549f
C720 a_n1986_13878.t63 gnd 0.707549f
C721 a_n1986_13878.t62 gnd 0.722451f
C722 a_n1986_13878.n58 gnd 0.313741f
C723 a_n1986_13878.t42 gnd 0.707549f
C724 a_n1986_13878.n59 gnd 0.307133f
C725 a_n1986_13878.n60 gnd 0.313742f
C726 a_n1986_13878.t43 gnd 0.719248f
C727 a_n1986_13878.t22 gnd 0.722451f
C728 a_n1986_13878.n61 gnd 0.313741f
C729 a_n1986_13878.t6 gnd 0.707549f
C730 a_n1986_13878.n62 gnd 0.307133f
C731 a_n1986_13878.n63 gnd 0.313742f
C732 a_n1986_13878.t10 gnd 0.719248f
C733 a_n1986_13878.n64 gnd 1.14966f
C734 a_n1986_13878.t47 gnd 0.707549f
C735 a_n1986_13878.n65 gnd 0.307133f
C736 a_n1986_13878.t53 gnd 0.707549f
C737 a_n1986_13878.n66 gnd 0.307133f
C738 a_n1986_13878.t45 gnd 0.707549f
C739 a_n1986_13878.n67 gnd 0.307133f
C740 a_n1986_13878.t58 gnd 0.707549f
C741 a_n1986_13878.n68 gnd 0.307133f
C742 a_n1986_13878.t49 gnd 0.707549f
C743 a_n1986_13878.n69 gnd 0.301556f
C744 a_n1986_13878.t40 gnd 0.707549f
C745 a_n1986_13878.n70 gnd 0.311083f
C746 a_n1986_13878.t51 gnd 0.719405f
C747 a_n1986_13878.t60 gnd 0.707549f
C748 a_n1986_13878.n71 gnd 0.301556f
C749 a_n1986_13878.t46 gnd 0.707549f
C750 a_n1986_13878.n72 gnd 0.311083f
C751 a_n1986_13878.t55 gnd 0.719405f
C752 a_n1986_13878.t64 gnd 0.707549f
C753 a_n1986_13878.n73 gnd 0.301556f
C754 a_n1986_13878.t52 gnd 0.707549f
C755 a_n1986_13878.n74 gnd 0.311083f
C756 a_n1986_13878.t66 gnd 0.719405f
C757 a_n1986_13878.t56 gnd 0.707549f
C758 a_n1986_13878.n75 gnd 0.301556f
C759 a_n1986_13878.t41 gnd 0.707549f
C760 a_n1986_13878.n76 gnd 0.311083f
C761 a_n1986_13878.t61 gnd 0.719405f
C762 a_n1986_13878.n77 gnd 1.35928f
C763 a_n1986_13878.n78 gnd 0.313742f
C764 a_n1986_13878.n79 gnd 0.307133f
C765 a_n1986_13878.n80 gnd 0.313741f
C766 a_n1986_13878.t35 gnd 0.118309f
C767 a_n1986_13878.t32 gnd 0.118309f
C768 a_n1986_13878.n81 gnd 1.04709f
C769 a_n1986_13878.t24 gnd 0.118309f
C770 a_n1986_13878.t34 gnd 0.118309f
C771 a_n1986_13878.n82 gnd 1.04542f
C772 a_n1986_13878.t30 gnd 0.118309f
C773 a_n1986_13878.t26 gnd 0.118309f
C774 a_n1986_13878.n83 gnd 1.04709f
C775 a_n1986_13878.t36 gnd 0.118309f
C776 a_n1986_13878.t31 gnd 0.118309f
C777 a_n1986_13878.n84 gnd 1.04542f
C778 a_n1986_13878.t29 gnd 0.118309f
C779 a_n1986_13878.t28 gnd 0.118309f
C780 a_n1986_13878.n85 gnd 1.04542f
C781 a_n1986_13878.t27 gnd 0.118309f
C782 a_n1986_13878.t33 gnd 0.118309f
C783 a_n1986_13878.n86 gnd 1.04542f
C784 a_n1986_13878.t39 gnd 0.118309f
C785 a_n1986_13878.t37 gnd 0.118309f
C786 a_n1986_13878.n87 gnd 1.04709f
C787 a_n1986_13878.t25 gnd 0.118309f
C788 a_n1986_13878.t38 gnd 0.118309f
C789 a_n1986_13878.n88 gnd 1.04542f
C790 a_n1986_13878.n89 gnd 0.313742f
C791 a_n1986_13878.n90 gnd 0.307133f
C792 a_n1986_13878.n91 gnd 0.313741f
C793 a_n1986_13878.n92 gnd 0.799185f
C794 a_n1986_13878.t21 gnd 1.42146f
C795 a_n1986_13878.t3 gnd 0.152112f
C796 a_n1986_13878.t13 gnd 0.152112f
C797 a_n1986_13878.n93 gnd 1.07147f
C798 a_n1986_13878.t19 gnd 0.152112f
C799 a_n1986_13878.t9 gnd 0.152112f
C800 a_n1986_13878.n94 gnd 1.07147f
C801 a_n1986_13878.t1 gnd 1.4243f
C802 a_n6308_8799.n0 gnd 0.178004f
C803 a_n6308_8799.n1 gnd 0.208454f
C804 a_n6308_8799.n2 gnd 0.208454f
C805 a_n6308_8799.n3 gnd 0.208454f
C806 a_n6308_8799.n4 gnd 0.178004f
C807 a_n6308_8799.n5 gnd 0.208454f
C808 a_n6308_8799.n6 gnd 0.208454f
C809 a_n6308_8799.n7 gnd 0.208454f
C810 a_n6308_8799.n8 gnd 0.343842f
C811 a_n6308_8799.n9 gnd 0.208454f
C812 a_n6308_8799.n10 gnd 0.208454f
C813 a_n6308_8799.n11 gnd 0.208454f
C814 a_n6308_8799.n12 gnd 0.208454f
C815 a_n6308_8799.n13 gnd 0.208454f
C816 a_n6308_8799.n14 gnd 0.178004f
C817 a_n6308_8799.n15 gnd 0.208454f
C818 a_n6308_8799.n16 gnd 0.208454f
C819 a_n6308_8799.n17 gnd 0.208454f
C820 a_n6308_8799.n18 gnd 0.178004f
C821 a_n6308_8799.n19 gnd 0.208454f
C822 a_n6308_8799.n20 gnd 0.208454f
C823 a_n6308_8799.n21 gnd 0.208454f
C824 a_n6308_8799.n22 gnd 0.343842f
C825 a_n6308_8799.n23 gnd 0.208454f
C826 a_n6308_8799.n24 gnd 2.87873f
C827 a_n6308_8799.n25 gnd 3.94079f
C828 a_n6308_8799.n26 gnd 2.3968f
C829 a_n6308_8799.n27 gnd 1.40084f
C830 a_n6308_8799.n28 gnd 3.10097f
C831 a_n6308_8799.n29 gnd 0.25209f
C832 a_n6308_8799.n31 gnd 0.007764f
C833 a_n6308_8799.n32 gnd 0.011735f
C834 a_n6308_8799.n33 gnd 0.008071f
C835 a_n6308_8799.n35 gnd 4.03e-19
C836 a_n6308_8799.n36 gnd 0.008364f
C837 a_n6308_8799.n37 gnd 0.263716f
C838 a_n6308_8799.n38 gnd 0.25209f
C839 a_n6308_8799.n40 gnd 0.007764f
C840 a_n6308_8799.n41 gnd 0.011735f
C841 a_n6308_8799.n42 gnd 0.008071f
C842 a_n6308_8799.n44 gnd 4.03e-19
C843 a_n6308_8799.n45 gnd 0.008364f
C844 a_n6308_8799.n46 gnd 0.263716f
C845 a_n6308_8799.n47 gnd 0.25209f
C846 a_n6308_8799.n49 gnd 0.007764f
C847 a_n6308_8799.n50 gnd 0.011735f
C848 a_n6308_8799.n51 gnd 0.008071f
C849 a_n6308_8799.n53 gnd 4.03e-19
C850 a_n6308_8799.n54 gnd 0.008364f
C851 a_n6308_8799.n55 gnd 0.263716f
C852 a_n6308_8799.n56 gnd 0.008364f
C853 a_n6308_8799.n57 gnd 0.263716f
C854 a_n6308_8799.n58 gnd 4.03e-19
C855 a_n6308_8799.n60 gnd 0.008071f
C856 a_n6308_8799.n61 gnd 0.011735f
C857 a_n6308_8799.n62 gnd 0.007764f
C858 a_n6308_8799.n64 gnd 0.25209f
C859 a_n6308_8799.n65 gnd 0.008364f
C860 a_n6308_8799.n66 gnd 0.263716f
C861 a_n6308_8799.n67 gnd 4.03e-19
C862 a_n6308_8799.n69 gnd 0.008071f
C863 a_n6308_8799.n70 gnd 0.011735f
C864 a_n6308_8799.n71 gnd 0.007764f
C865 a_n6308_8799.n73 gnd 0.25209f
C866 a_n6308_8799.n74 gnd 0.008364f
C867 a_n6308_8799.n75 gnd 0.263716f
C868 a_n6308_8799.n76 gnd 4.03e-19
C869 a_n6308_8799.n78 gnd 0.008071f
C870 a_n6308_8799.n79 gnd 0.011735f
C871 a_n6308_8799.n80 gnd 0.007764f
C872 a_n6308_8799.n82 gnd 0.25209f
C873 a_n6308_8799.t17 gnd 0.144586f
C874 a_n6308_8799.t1 gnd 0.144586f
C875 a_n6308_8799.t7 gnd 0.144586f
C876 a_n6308_8799.n83 gnd 1.14038f
C877 a_n6308_8799.t16 gnd 0.144586f
C878 a_n6308_8799.t25 gnd 0.144586f
C879 a_n6308_8799.n84 gnd 1.13849f
C880 a_n6308_8799.t11 gnd 0.144586f
C881 a_n6308_8799.t22 gnd 0.144586f
C882 a_n6308_8799.n85 gnd 1.13849f
C883 a_n6308_8799.t23 gnd 0.112456f
C884 a_n6308_8799.t5 gnd 0.112456f
C885 a_n6308_8799.n86 gnd 0.995285f
C886 a_n6308_8799.t9 gnd 0.112456f
C887 a_n6308_8799.t2 gnd 0.112456f
C888 a_n6308_8799.n87 gnd 0.993701f
C889 a_n6308_8799.t26 gnd 0.112456f
C890 a_n6308_8799.t15 gnd 0.112456f
C891 a_n6308_8799.n88 gnd 0.995284f
C892 a_n6308_8799.t14 gnd 0.112456f
C893 a_n6308_8799.t21 gnd 0.112456f
C894 a_n6308_8799.n89 gnd 0.9937f
C895 a_n6308_8799.t3 gnd 0.112456f
C896 a_n6308_8799.t6 gnd 0.112456f
C897 a_n6308_8799.n90 gnd 0.995284f
C898 a_n6308_8799.t4 gnd 0.112456f
C899 a_n6308_8799.t8 gnd 0.112456f
C900 a_n6308_8799.n91 gnd 0.9937f
C901 a_n6308_8799.t13 gnd 0.112456f
C902 a_n6308_8799.t27 gnd 0.112456f
C903 a_n6308_8799.n92 gnd 0.993701f
C904 a_n6308_8799.t24 gnd 0.112456f
C905 a_n6308_8799.t20 gnd 0.112456f
C906 a_n6308_8799.n93 gnd 0.993701f
C907 a_n6308_8799.t87 gnd 0.599522f
C908 a_n6308_8799.n94 gnd 0.271337f
C909 a_n6308_8799.t35 gnd 0.599522f
C910 a_n6308_8799.t36 gnd 0.599522f
C911 a_n6308_8799.n95 gnd 0.262457f
C912 a_n6308_8799.t49 gnd 0.599522f
C913 a_n6308_8799.n96 gnd 0.273879f
C914 a_n6308_8799.t64 gnd 0.599522f
C915 a_n6308_8799.t77 gnd 0.599522f
C916 a_n6308_8799.n97 gnd 0.267276f
C917 a_n6308_8799.t52 gnd 0.613613f
C918 a_n6308_8799.t53 gnd 0.599522f
C919 a_n6308_8799.n98 gnd 0.273442f
C920 a_n6308_8799.n99 gnd 0.249913f
C921 a_n6308_8799.t29 gnd 0.599522f
C922 a_n6308_8799.n100 gnd 0.271219f
C923 a_n6308_8799.n101 gnd 0.271352f
C924 a_n6308_8799.t89 gnd 0.599522f
C925 a_n6308_8799.n102 gnd 0.267597f
C926 a_n6308_8799.t48 gnd 0.599522f
C927 a_n6308_8799.n103 gnd 0.267848f
C928 a_n6308_8799.n104 gnd 0.273443f
C929 a_n6308_8799.t34 gnd 0.610406f
C930 a_n6308_8799.t93 gnd 0.599522f
C931 a_n6308_8799.n105 gnd 0.271337f
C932 a_n6308_8799.t41 gnd 0.599522f
C933 a_n6308_8799.t45 gnd 0.599522f
C934 a_n6308_8799.n106 gnd 0.262457f
C935 a_n6308_8799.t57 gnd 0.599522f
C936 a_n6308_8799.n107 gnd 0.273879f
C937 a_n6308_8799.t71 gnd 0.599522f
C938 a_n6308_8799.t84 gnd 0.599522f
C939 a_n6308_8799.n108 gnd 0.267276f
C940 a_n6308_8799.t58 gnd 0.613613f
C941 a_n6308_8799.t59 gnd 0.599522f
C942 a_n6308_8799.n109 gnd 0.273442f
C943 a_n6308_8799.n110 gnd 0.249913f
C944 a_n6308_8799.t37 gnd 0.599522f
C945 a_n6308_8799.n111 gnd 0.271219f
C946 a_n6308_8799.n112 gnd 0.271352f
C947 a_n6308_8799.t97 gnd 0.599522f
C948 a_n6308_8799.n113 gnd 0.267597f
C949 a_n6308_8799.t56 gnd 0.599522f
C950 a_n6308_8799.n114 gnd 0.267848f
C951 a_n6308_8799.n115 gnd 0.273443f
C952 a_n6308_8799.t43 gnd 0.610406f
C953 a_n6308_8799.n116 gnd 0.900047f
C954 a_n6308_8799.t68 gnd 0.599522f
C955 a_n6308_8799.n117 gnd 0.271337f
C956 a_n6308_8799.t39 gnd 0.599522f
C957 a_n6308_8799.t86 gnd 0.599522f
C958 a_n6308_8799.n118 gnd 0.262457f
C959 a_n6308_8799.t33 gnd 0.599522f
C960 a_n6308_8799.n119 gnd 0.273879f
C961 a_n6308_8799.t74 gnd 0.599522f
C962 a_n6308_8799.t95 gnd 0.599522f
C963 a_n6308_8799.n120 gnd 0.267276f
C964 a_n6308_8799.t91 gnd 0.613613f
C965 a_n6308_8799.t79 gnd 0.599522f
C966 a_n6308_8799.n121 gnd 0.273442f
C967 a_n6308_8799.n122 gnd 0.249913f
C968 a_n6308_8799.t63 gnd 0.599522f
C969 a_n6308_8799.n123 gnd 0.271219f
C970 a_n6308_8799.n124 gnd 0.271352f
C971 a_n6308_8799.t44 gnd 0.599522f
C972 a_n6308_8799.n125 gnd 0.267597f
C973 a_n6308_8799.t51 gnd 0.599522f
C974 a_n6308_8799.n126 gnd 0.267848f
C975 a_n6308_8799.n127 gnd 0.273443f
C976 a_n6308_8799.t99 gnd 0.610406f
C977 a_n6308_8799.n128 gnd 1.40092f
C978 a_n6308_8799.t61 gnd 0.610406f
C979 a_n6308_8799.t60 gnd 0.599522f
C980 a_n6308_8799.t42 gnd 0.599522f
C981 a_n6308_8799.t88 gnd 0.599522f
C982 a_n6308_8799.n129 gnd 0.267848f
C983 a_n6308_8799.t62 gnd 0.599522f
C984 a_n6308_8799.t47 gnd 0.599522f
C985 a_n6308_8799.t90 gnd 0.599522f
C986 a_n6308_8799.n130 gnd 0.271352f
C987 a_n6308_8799.t72 gnd 0.599522f
C988 a_n6308_8799.t70 gnd 0.599522f
C989 a_n6308_8799.t31 gnd 0.599522f
C990 a_n6308_8799.n131 gnd 0.267276f
C991 a_n6308_8799.t75 gnd 0.613613f
C992 a_n6308_8799.t76 gnd 0.599522f
C993 a_n6308_8799.n132 gnd 0.273442f
C994 a_n6308_8799.n133 gnd 0.249913f
C995 a_n6308_8799.n134 gnd 0.271219f
C996 a_n6308_8799.n135 gnd 0.273879f
C997 a_n6308_8799.n136 gnd 0.267597f
C998 a_n6308_8799.n137 gnd 0.262457f
C999 a_n6308_8799.n138 gnd 0.271337f
C1000 a_n6308_8799.n139 gnd 0.273443f
C1001 a_n6308_8799.t66 gnd 0.610406f
C1002 a_n6308_8799.t65 gnd 0.599522f
C1003 a_n6308_8799.t54 gnd 0.599522f
C1004 a_n6308_8799.t96 gnd 0.599522f
C1005 a_n6308_8799.n140 gnd 0.267848f
C1006 a_n6308_8799.t69 gnd 0.599522f
C1007 a_n6308_8799.t55 gnd 0.599522f
C1008 a_n6308_8799.t28 gnd 0.599522f
C1009 a_n6308_8799.n141 gnd 0.271352f
C1010 a_n6308_8799.t81 gnd 0.599522f
C1011 a_n6308_8799.t80 gnd 0.599522f
C1012 a_n6308_8799.t38 gnd 0.599522f
C1013 a_n6308_8799.n142 gnd 0.267276f
C1014 a_n6308_8799.t82 gnd 0.613613f
C1015 a_n6308_8799.t83 gnd 0.599522f
C1016 a_n6308_8799.n143 gnd 0.273442f
C1017 a_n6308_8799.n144 gnd 0.249913f
C1018 a_n6308_8799.n145 gnd 0.271219f
C1019 a_n6308_8799.n146 gnd 0.273879f
C1020 a_n6308_8799.n147 gnd 0.267597f
C1021 a_n6308_8799.n148 gnd 0.262457f
C1022 a_n6308_8799.n149 gnd 0.271337f
C1023 a_n6308_8799.n150 gnd 0.273443f
C1024 a_n6308_8799.n151 gnd 0.900047f
C1025 a_n6308_8799.t98 gnd 0.610406f
C1026 a_n6308_8799.t40 gnd 0.599522f
C1027 a_n6308_8799.t67 gnd 0.599522f
C1028 a_n6308_8799.t30 gnd 0.599522f
C1029 a_n6308_8799.n152 gnd 0.267848f
C1030 a_n6308_8799.t85 gnd 0.599522f
C1031 a_n6308_8799.t46 gnd 0.599522f
C1032 a_n6308_8799.t73 gnd 0.599522f
C1033 a_n6308_8799.n153 gnd 0.271352f
C1034 a_n6308_8799.t32 gnd 0.599522f
C1035 a_n6308_8799.t50 gnd 0.599522f
C1036 a_n6308_8799.t94 gnd 0.599522f
C1037 a_n6308_8799.n154 gnd 0.267276f
C1038 a_n6308_8799.t92 gnd 0.613613f
C1039 a_n6308_8799.t78 gnd 0.599522f
C1040 a_n6308_8799.n155 gnd 0.273442f
C1041 a_n6308_8799.n156 gnd 0.249913f
C1042 a_n6308_8799.n157 gnd 0.271219f
C1043 a_n6308_8799.n158 gnd 0.273879f
C1044 a_n6308_8799.n159 gnd 0.267597f
C1045 a_n6308_8799.n160 gnd 0.262457f
C1046 a_n6308_8799.n161 gnd 0.271337f
C1047 a_n6308_8799.n162 gnd 0.273443f
C1048 a_n6308_8799.n163 gnd 1.17834f
C1049 a_n6308_8799.n164 gnd 12.2976f
C1050 a_n6308_8799.n165 gnd 4.38763f
C1051 a_n6308_8799.n166 gnd 5.71511f
C1052 a_n6308_8799.t19 gnd 0.144586f
C1053 a_n6308_8799.t10 gnd 0.144586f
C1054 a_n6308_8799.n167 gnd 1.13849f
C1055 a_n6308_8799.t12 gnd 0.144586f
C1056 a_n6308_8799.t18 gnd 0.144586f
C1057 a_n6308_8799.n168 gnd 1.14037f
C1058 a_n6308_8799.n169 gnd 1.13849f
C1059 a_n6308_8799.t0 gnd 0.144586f
C1060 vdd.t2 gnd 0.035814f
C1061 vdd.t58 gnd 0.035814f
C1062 vdd.n0 gnd 0.282475f
C1063 vdd.t29 gnd 0.035814f
C1064 vdd.t44 gnd 0.035814f
C1065 vdd.n1 gnd 0.282008f
C1066 vdd.n2 gnd 0.260066f
C1067 vdd.t198 gnd 0.035814f
C1068 vdd.t160 gnd 0.035814f
C1069 vdd.n3 gnd 0.282008f
C1070 vdd.n4 gnd 0.131525f
C1071 vdd.t155 gnd 0.035814f
C1072 vdd.t205 gnd 0.035814f
C1073 vdd.n5 gnd 0.282008f
C1074 vdd.n6 gnd 0.123412f
C1075 vdd.t153 gnd 0.035814f
C1076 vdd.t4 gnd 0.035814f
C1077 vdd.n7 gnd 0.282475f
C1078 vdd.t56 gnd 0.035814f
C1079 vdd.t227 gnd 0.035814f
C1080 vdd.n8 gnd 0.282008f
C1081 vdd.n9 gnd 0.260066f
C1082 vdd.t67 gnd 0.035814f
C1083 vdd.t70 gnd 0.035814f
C1084 vdd.n10 gnd 0.282008f
C1085 vdd.n11 gnd 0.131525f
C1086 vdd.t157 gnd 0.035814f
C1087 vdd.t24 gnd 0.035814f
C1088 vdd.n12 gnd 0.282008f
C1089 vdd.n13 gnd 0.123412f
C1090 vdd.n14 gnd 0.08725f
C1091 vdd.t215 gnd 0.019897f
C1092 vdd.t223 gnd 0.019897f
C1093 vdd.n15 gnd 0.183143f
C1094 vdd.t217 gnd 0.019897f
C1095 vdd.t211 gnd 0.019897f
C1096 vdd.n16 gnd 0.182607f
C1097 vdd.n17 gnd 0.317793f
C1098 vdd.t225 gnd 0.019897f
C1099 vdd.t219 gnd 0.019897f
C1100 vdd.n18 gnd 0.182607f
C1101 vdd.n19 gnd 0.131475f
C1102 vdd.t210 gnd 0.019897f
C1103 vdd.t212 gnd 0.019897f
C1104 vdd.n20 gnd 0.183143f
C1105 vdd.t218 gnd 0.019897f
C1106 vdd.t222 gnd 0.019897f
C1107 vdd.n21 gnd 0.182607f
C1108 vdd.n22 gnd 0.317793f
C1109 vdd.t214 gnd 0.019897f
C1110 vdd.t213 gnd 0.019897f
C1111 vdd.n23 gnd 0.182607f
C1112 vdd.n24 gnd 0.131475f
C1113 vdd.t216 gnd 0.019897f
C1114 vdd.t224 gnd 0.019897f
C1115 vdd.n25 gnd 0.182607f
C1116 vdd.t221 gnd 0.019897f
C1117 vdd.t220 gnd 0.019897f
C1118 vdd.n26 gnd 0.182607f
C1119 vdd.n27 gnd 21.037899f
C1120 vdd.n28 gnd 7.7082f
C1121 vdd.n29 gnd 0.005427f
C1122 vdd.n30 gnd 0.005036f
C1123 vdd.n31 gnd 0.002786f
C1124 vdd.n32 gnd 0.006396f
C1125 vdd.n33 gnd 0.002706f
C1126 vdd.n34 gnd 0.002865f
C1127 vdd.n35 gnd 0.005036f
C1128 vdd.n36 gnd 0.002706f
C1129 vdd.n37 gnd 0.006396f
C1130 vdd.n38 gnd 0.002865f
C1131 vdd.n39 gnd 0.005036f
C1132 vdd.n40 gnd 0.002706f
C1133 vdd.n41 gnd 0.004797f
C1134 vdd.n42 gnd 0.004811f
C1135 vdd.t16 gnd 0.013741f
C1136 vdd.n43 gnd 0.030574f
C1137 vdd.n44 gnd 0.159114f
C1138 vdd.n45 gnd 0.002706f
C1139 vdd.n46 gnd 0.002865f
C1140 vdd.n47 gnd 0.006396f
C1141 vdd.n48 gnd 0.006396f
C1142 vdd.n49 gnd 0.002865f
C1143 vdd.n50 gnd 0.002706f
C1144 vdd.n51 gnd 0.005036f
C1145 vdd.n52 gnd 0.005036f
C1146 vdd.n53 gnd 0.002706f
C1147 vdd.n54 gnd 0.002865f
C1148 vdd.n55 gnd 0.006396f
C1149 vdd.n56 gnd 0.006396f
C1150 vdd.n57 gnd 0.002865f
C1151 vdd.n58 gnd 0.002706f
C1152 vdd.n59 gnd 0.005036f
C1153 vdd.n60 gnd 0.005036f
C1154 vdd.n61 gnd 0.002706f
C1155 vdd.n62 gnd 0.002865f
C1156 vdd.n63 gnd 0.006396f
C1157 vdd.n64 gnd 0.006396f
C1158 vdd.n65 gnd 0.015121f
C1159 vdd.n66 gnd 0.002786f
C1160 vdd.n67 gnd 0.002706f
C1161 vdd.n68 gnd 0.013016f
C1162 vdd.n69 gnd 0.009087f
C1163 vdd.t176 gnd 0.031835f
C1164 vdd.t73 gnd 0.031835f
C1165 vdd.n70 gnd 0.218793f
C1166 vdd.n71 gnd 0.172047f
C1167 vdd.t172 gnd 0.031835f
C1168 vdd.t180 gnd 0.031835f
C1169 vdd.n72 gnd 0.218793f
C1170 vdd.n73 gnd 0.138841f
C1171 vdd.t202 gnd 0.031835f
C1172 vdd.t166 gnd 0.031835f
C1173 vdd.n74 gnd 0.218793f
C1174 vdd.n75 gnd 0.138841f
C1175 vdd.t170 gnd 0.031835f
C1176 vdd.t20 gnd 0.031835f
C1177 vdd.n76 gnd 0.218793f
C1178 vdd.n77 gnd 0.138841f
C1179 vdd.t35 gnd 0.031835f
C1180 vdd.t185 gnd 0.031835f
C1181 vdd.n78 gnd 0.218793f
C1182 vdd.n79 gnd 0.138841f
C1183 vdd.n80 gnd 0.005427f
C1184 vdd.n81 gnd 0.005036f
C1185 vdd.n82 gnd 0.002786f
C1186 vdd.n83 gnd 0.006396f
C1187 vdd.n84 gnd 0.002706f
C1188 vdd.n85 gnd 0.002865f
C1189 vdd.n86 gnd 0.005036f
C1190 vdd.n87 gnd 0.002706f
C1191 vdd.n88 gnd 0.006396f
C1192 vdd.n89 gnd 0.002865f
C1193 vdd.n90 gnd 0.005036f
C1194 vdd.n91 gnd 0.002706f
C1195 vdd.n92 gnd 0.004797f
C1196 vdd.n93 gnd 0.004811f
C1197 vdd.t38 gnd 0.013741f
C1198 vdd.n94 gnd 0.030574f
C1199 vdd.n95 gnd 0.159114f
C1200 vdd.n96 gnd 0.002706f
C1201 vdd.n97 gnd 0.002865f
C1202 vdd.n98 gnd 0.006396f
C1203 vdd.n99 gnd 0.006396f
C1204 vdd.n100 gnd 0.002865f
C1205 vdd.n101 gnd 0.002706f
C1206 vdd.n102 gnd 0.005036f
C1207 vdd.n103 gnd 0.005036f
C1208 vdd.n104 gnd 0.002706f
C1209 vdd.n105 gnd 0.002865f
C1210 vdd.n106 gnd 0.006396f
C1211 vdd.n107 gnd 0.006396f
C1212 vdd.n108 gnd 0.002865f
C1213 vdd.n109 gnd 0.002706f
C1214 vdd.n110 gnd 0.005036f
C1215 vdd.n111 gnd 0.005036f
C1216 vdd.n112 gnd 0.002706f
C1217 vdd.n113 gnd 0.002865f
C1218 vdd.n114 gnd 0.006396f
C1219 vdd.n115 gnd 0.006396f
C1220 vdd.n116 gnd 0.015121f
C1221 vdd.n117 gnd 0.002786f
C1222 vdd.n118 gnd 0.002706f
C1223 vdd.n119 gnd 0.013016f
C1224 vdd.n120 gnd 0.008802f
C1225 vdd.n121 gnd 0.103298f
C1226 vdd.n122 gnd 0.005427f
C1227 vdd.n123 gnd 0.005036f
C1228 vdd.n124 gnd 0.002786f
C1229 vdd.n125 gnd 0.006396f
C1230 vdd.n126 gnd 0.002706f
C1231 vdd.n127 gnd 0.002865f
C1232 vdd.n128 gnd 0.005036f
C1233 vdd.n129 gnd 0.002706f
C1234 vdd.n130 gnd 0.006396f
C1235 vdd.n131 gnd 0.002865f
C1236 vdd.n132 gnd 0.005036f
C1237 vdd.n133 gnd 0.002706f
C1238 vdd.n134 gnd 0.004797f
C1239 vdd.n135 gnd 0.004811f
C1240 vdd.t72 gnd 0.013741f
C1241 vdd.n136 gnd 0.030574f
C1242 vdd.n137 gnd 0.159114f
C1243 vdd.n138 gnd 0.002706f
C1244 vdd.n139 gnd 0.002865f
C1245 vdd.n140 gnd 0.006396f
C1246 vdd.n141 gnd 0.006396f
C1247 vdd.n142 gnd 0.002865f
C1248 vdd.n143 gnd 0.002706f
C1249 vdd.n144 gnd 0.005036f
C1250 vdd.n145 gnd 0.005036f
C1251 vdd.n146 gnd 0.002706f
C1252 vdd.n147 gnd 0.002865f
C1253 vdd.n148 gnd 0.006396f
C1254 vdd.n149 gnd 0.006396f
C1255 vdd.n150 gnd 0.002865f
C1256 vdd.n151 gnd 0.002706f
C1257 vdd.n152 gnd 0.005036f
C1258 vdd.n153 gnd 0.005036f
C1259 vdd.n154 gnd 0.002706f
C1260 vdd.n155 gnd 0.002865f
C1261 vdd.n156 gnd 0.006396f
C1262 vdd.n157 gnd 0.006396f
C1263 vdd.n158 gnd 0.015121f
C1264 vdd.n159 gnd 0.002786f
C1265 vdd.n160 gnd 0.002706f
C1266 vdd.n161 gnd 0.013016f
C1267 vdd.n162 gnd 0.009087f
C1268 vdd.t231 gnd 0.031835f
C1269 vdd.t190 gnd 0.031835f
C1270 vdd.n163 gnd 0.218793f
C1271 vdd.n164 gnd 0.172047f
C1272 vdd.t7 gnd 0.031835f
C1273 vdd.t33 gnd 0.031835f
C1274 vdd.n165 gnd 0.218793f
C1275 vdd.n166 gnd 0.138841f
C1276 vdd.t192 gnd 0.031835f
C1277 vdd.t174 gnd 0.031835f
C1278 vdd.n167 gnd 0.218793f
C1279 vdd.n168 gnd 0.138841f
C1280 vdd.t229 gnd 0.031835f
C1281 vdd.t228 gnd 0.031835f
C1282 vdd.n169 gnd 0.218793f
C1283 vdd.n170 gnd 0.138841f
C1284 vdd.t167 gnd 0.031835f
C1285 vdd.t13 gnd 0.031835f
C1286 vdd.n171 gnd 0.218793f
C1287 vdd.n172 gnd 0.138841f
C1288 vdd.n173 gnd 0.005427f
C1289 vdd.n174 gnd 0.005036f
C1290 vdd.n175 gnd 0.002786f
C1291 vdd.n176 gnd 0.006396f
C1292 vdd.n177 gnd 0.002706f
C1293 vdd.n178 gnd 0.002865f
C1294 vdd.n179 gnd 0.005036f
C1295 vdd.n180 gnd 0.002706f
C1296 vdd.n181 gnd 0.006396f
C1297 vdd.n182 gnd 0.002865f
C1298 vdd.n183 gnd 0.005036f
C1299 vdd.n184 gnd 0.002706f
C1300 vdd.n185 gnd 0.004797f
C1301 vdd.n186 gnd 0.004811f
C1302 vdd.t11 gnd 0.013741f
C1303 vdd.n187 gnd 0.030574f
C1304 vdd.n188 gnd 0.159114f
C1305 vdd.n189 gnd 0.002706f
C1306 vdd.n190 gnd 0.002865f
C1307 vdd.n191 gnd 0.006396f
C1308 vdd.n192 gnd 0.006396f
C1309 vdd.n193 gnd 0.002865f
C1310 vdd.n194 gnd 0.002706f
C1311 vdd.n195 gnd 0.005036f
C1312 vdd.n196 gnd 0.005036f
C1313 vdd.n197 gnd 0.002706f
C1314 vdd.n198 gnd 0.002865f
C1315 vdd.n199 gnd 0.006396f
C1316 vdd.n200 gnd 0.006396f
C1317 vdd.n201 gnd 0.002865f
C1318 vdd.n202 gnd 0.002706f
C1319 vdd.n203 gnd 0.005036f
C1320 vdd.n204 gnd 0.005036f
C1321 vdd.n205 gnd 0.002706f
C1322 vdd.n206 gnd 0.002865f
C1323 vdd.n207 gnd 0.006396f
C1324 vdd.n208 gnd 0.006396f
C1325 vdd.n209 gnd 0.015121f
C1326 vdd.n210 gnd 0.002786f
C1327 vdd.n211 gnd 0.002706f
C1328 vdd.n212 gnd 0.013016f
C1329 vdd.n213 gnd 0.008802f
C1330 vdd.n214 gnd 0.061452f
C1331 vdd.n215 gnd 0.221428f
C1332 vdd.n216 gnd 0.005427f
C1333 vdd.n217 gnd 0.005036f
C1334 vdd.n218 gnd 0.002786f
C1335 vdd.n219 gnd 0.006396f
C1336 vdd.n220 gnd 0.002706f
C1337 vdd.n221 gnd 0.002865f
C1338 vdd.n222 gnd 0.005036f
C1339 vdd.n223 gnd 0.002706f
C1340 vdd.n224 gnd 0.006396f
C1341 vdd.n225 gnd 0.002865f
C1342 vdd.n226 gnd 0.005036f
C1343 vdd.n227 gnd 0.002706f
C1344 vdd.n228 gnd 0.004797f
C1345 vdd.n229 gnd 0.004811f
C1346 vdd.t42 gnd 0.013741f
C1347 vdd.n230 gnd 0.030574f
C1348 vdd.n231 gnd 0.159114f
C1349 vdd.n232 gnd 0.002706f
C1350 vdd.n233 gnd 0.002865f
C1351 vdd.n234 gnd 0.006396f
C1352 vdd.n235 gnd 0.006396f
C1353 vdd.n236 gnd 0.002865f
C1354 vdd.n237 gnd 0.002706f
C1355 vdd.n238 gnd 0.005036f
C1356 vdd.n239 gnd 0.005036f
C1357 vdd.n240 gnd 0.002706f
C1358 vdd.n241 gnd 0.002865f
C1359 vdd.n242 gnd 0.006396f
C1360 vdd.n243 gnd 0.006396f
C1361 vdd.n244 gnd 0.002865f
C1362 vdd.n245 gnd 0.002706f
C1363 vdd.n246 gnd 0.005036f
C1364 vdd.n247 gnd 0.005036f
C1365 vdd.n248 gnd 0.002706f
C1366 vdd.n249 gnd 0.002865f
C1367 vdd.n250 gnd 0.006396f
C1368 vdd.n251 gnd 0.006396f
C1369 vdd.n252 gnd 0.015121f
C1370 vdd.n253 gnd 0.002786f
C1371 vdd.n254 gnd 0.002706f
C1372 vdd.n255 gnd 0.013016f
C1373 vdd.n256 gnd 0.009087f
C1374 vdd.t41 gnd 0.031835f
C1375 vdd.t53 gnd 0.031835f
C1376 vdd.n257 gnd 0.218793f
C1377 vdd.n258 gnd 0.172047f
C1378 vdd.t183 gnd 0.031835f
C1379 vdd.t49 gnd 0.031835f
C1380 vdd.n259 gnd 0.218793f
C1381 vdd.n260 gnd 0.138841f
C1382 vdd.t203 gnd 0.031835f
C1383 vdd.t61 gnd 0.031835f
C1384 vdd.n261 gnd 0.218793f
C1385 vdd.n262 gnd 0.138841f
C1386 vdd.t165 gnd 0.031835f
C1387 vdd.t161 gnd 0.031835f
C1388 vdd.n263 gnd 0.218793f
C1389 vdd.n264 gnd 0.138841f
C1390 vdd.t173 gnd 0.031835f
C1391 vdd.t64 gnd 0.031835f
C1392 vdd.n265 gnd 0.218793f
C1393 vdd.n266 gnd 0.138841f
C1394 vdd.n267 gnd 0.005427f
C1395 vdd.n268 gnd 0.005036f
C1396 vdd.n269 gnd 0.002786f
C1397 vdd.n270 gnd 0.006396f
C1398 vdd.n271 gnd 0.002706f
C1399 vdd.n272 gnd 0.002865f
C1400 vdd.n273 gnd 0.005036f
C1401 vdd.n274 gnd 0.002706f
C1402 vdd.n275 gnd 0.006396f
C1403 vdd.n276 gnd 0.002865f
C1404 vdd.n277 gnd 0.005036f
C1405 vdd.n278 gnd 0.002706f
C1406 vdd.n279 gnd 0.004797f
C1407 vdd.n280 gnd 0.004811f
C1408 vdd.t207 gnd 0.013741f
C1409 vdd.n281 gnd 0.030574f
C1410 vdd.n282 gnd 0.159114f
C1411 vdd.n283 gnd 0.002706f
C1412 vdd.n284 gnd 0.002865f
C1413 vdd.n285 gnd 0.006396f
C1414 vdd.n286 gnd 0.006396f
C1415 vdd.n287 gnd 0.002865f
C1416 vdd.n288 gnd 0.002706f
C1417 vdd.n289 gnd 0.005036f
C1418 vdd.n290 gnd 0.005036f
C1419 vdd.n291 gnd 0.002706f
C1420 vdd.n292 gnd 0.002865f
C1421 vdd.n293 gnd 0.006396f
C1422 vdd.n294 gnd 0.006396f
C1423 vdd.n295 gnd 0.002865f
C1424 vdd.n296 gnd 0.002706f
C1425 vdd.n297 gnd 0.005036f
C1426 vdd.n298 gnd 0.005036f
C1427 vdd.n299 gnd 0.002706f
C1428 vdd.n300 gnd 0.002865f
C1429 vdd.n301 gnd 0.006396f
C1430 vdd.n302 gnd 0.006396f
C1431 vdd.n303 gnd 0.015121f
C1432 vdd.n304 gnd 0.002786f
C1433 vdd.n305 gnd 0.002706f
C1434 vdd.n306 gnd 0.013016f
C1435 vdd.n307 gnd 0.008802f
C1436 vdd.n308 gnd 0.061452f
C1437 vdd.n309 gnd 0.243357f
C1438 vdd.n310 gnd 0.009854f
C1439 vdd.n311 gnd 0.009854f
C1440 vdd.n312 gnd 0.007959f
C1441 vdd.n313 gnd 0.007959f
C1442 vdd.n314 gnd 0.009888f
C1443 vdd.n315 gnd 0.009888f
C1444 vdd.t191 gnd 0.505262f
C1445 vdd.n316 gnd 0.009888f
C1446 vdd.n317 gnd 0.009888f
C1447 vdd.n318 gnd 0.009888f
C1448 vdd.t164 gnd 0.505262f
C1449 vdd.n319 gnd 0.009888f
C1450 vdd.n320 gnd 0.009888f
C1451 vdd.n321 gnd 0.009888f
C1452 vdd.n322 gnd 0.009888f
C1453 vdd.n323 gnd 0.007959f
C1454 vdd.n324 gnd 0.009888f
C1455 vdd.n325 gnd 0.813471f
C1456 vdd.n326 gnd 0.009888f
C1457 vdd.n327 gnd 0.009888f
C1458 vdd.n328 gnd 0.009888f
C1459 vdd.n329 gnd 0.692209f
C1460 vdd.n330 gnd 0.009888f
C1461 vdd.n331 gnd 0.009888f
C1462 vdd.n332 gnd 0.009888f
C1463 vdd.n333 gnd 0.009888f
C1464 vdd.n334 gnd 0.009888f
C1465 vdd.n335 gnd 0.007959f
C1466 vdd.n336 gnd 0.009888f
C1467 vdd.t12 gnd 0.505262f
C1468 vdd.n337 gnd 0.009888f
C1469 vdd.n338 gnd 0.009888f
C1470 vdd.n339 gnd 0.009888f
C1471 vdd.n340 gnd 1.01052f
C1472 vdd.n341 gnd 0.009888f
C1473 vdd.n342 gnd 0.009888f
C1474 vdd.n343 gnd 0.009888f
C1475 vdd.n344 gnd 0.009888f
C1476 vdd.n345 gnd 0.009888f
C1477 vdd.n346 gnd 0.007959f
C1478 vdd.n347 gnd 0.009888f
C1479 vdd.n348 gnd 0.009888f
C1480 vdd.n349 gnd 0.009888f
C1481 vdd.n350 gnd 0.023302f
C1482 vdd.n351 gnd 2.3242f
C1483 vdd.n352 gnd 0.023667f
C1484 vdd.n353 gnd 0.009888f
C1485 vdd.n354 gnd 0.009888f
C1486 vdd.n356 gnd 0.009888f
C1487 vdd.n357 gnd 0.009888f
C1488 vdd.n358 gnd 0.007959f
C1489 vdd.n359 gnd 0.007959f
C1490 vdd.n360 gnd 0.009888f
C1491 vdd.n361 gnd 0.009888f
C1492 vdd.n362 gnd 0.009888f
C1493 vdd.n363 gnd 0.009888f
C1494 vdd.n364 gnd 0.009888f
C1495 vdd.n365 gnd 0.009888f
C1496 vdd.n366 gnd 0.007959f
C1497 vdd.n368 gnd 0.009888f
C1498 vdd.n369 gnd 0.009888f
C1499 vdd.n370 gnd 0.009888f
C1500 vdd.n371 gnd 0.009888f
C1501 vdd.n372 gnd 0.009888f
C1502 vdd.n373 gnd 0.007959f
C1503 vdd.n375 gnd 0.009888f
C1504 vdd.n376 gnd 0.009888f
C1505 vdd.n377 gnd 0.009888f
C1506 vdd.n378 gnd 0.009888f
C1507 vdd.n379 gnd 0.009888f
C1508 vdd.n380 gnd 0.007959f
C1509 vdd.n382 gnd 0.009888f
C1510 vdd.n383 gnd 0.009888f
C1511 vdd.n384 gnd 0.009888f
C1512 vdd.n385 gnd 0.009888f
C1513 vdd.n386 gnd 0.006646f
C1514 vdd.t151 gnd 0.12165f
C1515 vdd.t150 gnd 0.130011f
C1516 vdd.t149 gnd 0.158874f
C1517 vdd.n387 gnd 0.203654f
C1518 vdd.n388 gnd 0.171902f
C1519 vdd.n390 gnd 0.009888f
C1520 vdd.n391 gnd 0.009888f
C1521 vdd.n392 gnd 0.007959f
C1522 vdd.n393 gnd 0.009888f
C1523 vdd.n395 gnd 0.009888f
C1524 vdd.n396 gnd 0.009888f
C1525 vdd.n397 gnd 0.009888f
C1526 vdd.n398 gnd 0.009888f
C1527 vdd.n399 gnd 0.007959f
C1528 vdd.n401 gnd 0.009888f
C1529 vdd.n402 gnd 0.009888f
C1530 vdd.n403 gnd 0.009888f
C1531 vdd.n404 gnd 0.009888f
C1532 vdd.n405 gnd 0.009888f
C1533 vdd.n406 gnd 0.007959f
C1534 vdd.n408 gnd 0.009888f
C1535 vdd.n409 gnd 0.009888f
C1536 vdd.n410 gnd 0.009888f
C1537 vdd.n411 gnd 0.009888f
C1538 vdd.n412 gnd 0.009888f
C1539 vdd.n413 gnd 0.007959f
C1540 vdd.n415 gnd 0.009888f
C1541 vdd.n416 gnd 0.009888f
C1542 vdd.n417 gnd 0.009888f
C1543 vdd.n418 gnd 0.009888f
C1544 vdd.n419 gnd 0.009888f
C1545 vdd.n420 gnd 0.007959f
C1546 vdd.n422 gnd 0.009888f
C1547 vdd.n423 gnd 0.009888f
C1548 vdd.n424 gnd 0.009888f
C1549 vdd.n425 gnd 0.009888f
C1550 vdd.n426 gnd 0.007879f
C1551 vdd.t139 gnd 0.12165f
C1552 vdd.t138 gnd 0.130011f
C1553 vdd.t136 gnd 0.158874f
C1554 vdd.n427 gnd 0.203654f
C1555 vdd.n428 gnd 0.171902f
C1556 vdd.n430 gnd 0.009888f
C1557 vdd.n431 gnd 0.009888f
C1558 vdd.n432 gnd 0.007959f
C1559 vdd.n433 gnd 0.009888f
C1560 vdd.n435 gnd 0.009888f
C1561 vdd.n436 gnd 0.009888f
C1562 vdd.n437 gnd 0.009888f
C1563 vdd.n438 gnd 0.009888f
C1564 vdd.n439 gnd 0.007959f
C1565 vdd.n441 gnd 0.009888f
C1566 vdd.n442 gnd 0.009888f
C1567 vdd.n443 gnd 0.009888f
C1568 vdd.n444 gnd 0.009888f
C1569 vdd.n445 gnd 0.009888f
C1570 vdd.n446 gnd 0.007959f
C1571 vdd.n448 gnd 0.009888f
C1572 vdd.n449 gnd 0.009888f
C1573 vdd.n450 gnd 0.009888f
C1574 vdd.n451 gnd 0.009888f
C1575 vdd.n452 gnd 0.009888f
C1576 vdd.n453 gnd 0.007959f
C1577 vdd.n455 gnd 0.009888f
C1578 vdd.n456 gnd 0.009888f
C1579 vdd.n457 gnd 0.009888f
C1580 vdd.n458 gnd 0.009888f
C1581 vdd.n459 gnd 0.009888f
C1582 vdd.n460 gnd 0.007959f
C1583 vdd.n462 gnd 0.009888f
C1584 vdd.n463 gnd 0.009888f
C1585 vdd.n464 gnd 0.009888f
C1586 vdd.n465 gnd 0.009888f
C1587 vdd.n466 gnd 0.009888f
C1588 vdd.n467 gnd 0.009888f
C1589 vdd.n468 gnd 0.007959f
C1590 vdd.n469 gnd 0.009888f
C1591 vdd.n470 gnd 0.009888f
C1592 vdd.n471 gnd 0.007959f
C1593 vdd.n472 gnd 0.009888f
C1594 vdd.n473 gnd 0.009888f
C1595 vdd.n474 gnd 0.007959f
C1596 vdd.n475 gnd 0.009888f
C1597 vdd.n476 gnd 0.007959f
C1598 vdd.n477 gnd 0.009888f
C1599 vdd.n478 gnd 0.007959f
C1600 vdd.n479 gnd 0.009888f
C1601 vdd.n480 gnd 0.009888f
C1602 vdd.t32 gnd 0.505262f
C1603 vdd.n481 gnd 0.54063f
C1604 vdd.n482 gnd 0.009888f
C1605 vdd.n483 gnd 0.007959f
C1606 vdd.n484 gnd 0.009888f
C1607 vdd.n485 gnd 0.007959f
C1608 vdd.n486 gnd 0.009888f
C1609 vdd.t6 gnd 0.505262f
C1610 vdd.n487 gnd 0.009888f
C1611 vdd.n488 gnd 0.007959f
C1612 vdd.n489 gnd 0.009888f
C1613 vdd.n490 gnd 0.007959f
C1614 vdd.n491 gnd 0.009888f
C1615 vdd.n492 gnd 0.793261f
C1616 vdd.n493 gnd 0.838735f
C1617 vdd.t52 gnd 0.505262f
C1618 vdd.n494 gnd 0.009888f
C1619 vdd.n495 gnd 0.007959f
C1620 vdd.n496 gnd 0.009888f
C1621 vdd.n497 gnd 0.007959f
C1622 vdd.n498 gnd 0.009888f
C1623 vdd.n499 gnd 0.621472f
C1624 vdd.n500 gnd 0.009888f
C1625 vdd.n501 gnd 0.007959f
C1626 vdd.n502 gnd 0.009888f
C1627 vdd.n503 gnd 0.007959f
C1628 vdd.n504 gnd 0.009888f
C1629 vdd.n505 gnd 1.01052f
C1630 vdd.t15 gnd 0.505262f
C1631 vdd.n506 gnd 0.009888f
C1632 vdd.n507 gnd 0.007959f
C1633 vdd.n508 gnd 0.009888f
C1634 vdd.n509 gnd 0.007959f
C1635 vdd.n510 gnd 0.009888f
C1636 vdd.n511 gnd 0.54063f
C1637 vdd.n512 gnd 0.009888f
C1638 vdd.n513 gnd 0.007959f
C1639 vdd.n514 gnd 0.023667f
C1640 vdd.n515 gnd 0.023667f
C1641 vdd.n516 gnd 7.23535f
C1642 vdd.t77 gnd 0.505262f
C1643 vdd.n517 gnd 0.023667f
C1644 vdd.n518 gnd 0.008504f
C1645 vdd.n519 gnd 0.007959f
C1646 vdd.n524 gnd 0.006328f
C1647 vdd.n525 gnd 0.007959f
C1648 vdd.n526 gnd 0.009888f
C1649 vdd.n527 gnd 0.009888f
C1650 vdd.n528 gnd 0.009888f
C1651 vdd.n529 gnd 0.009888f
C1652 vdd.n530 gnd 0.009888f
C1653 vdd.n531 gnd 0.007959f
C1654 vdd.n532 gnd 0.009888f
C1655 vdd.n533 gnd 0.009888f
C1656 vdd.n534 gnd 0.009888f
C1657 vdd.n535 gnd 0.009888f
C1658 vdd.n536 gnd 0.009888f
C1659 vdd.n537 gnd 0.007959f
C1660 vdd.n538 gnd 0.009888f
C1661 vdd.n539 gnd 0.009888f
C1662 vdd.n540 gnd 0.009888f
C1663 vdd.n541 gnd 0.009888f
C1664 vdd.n542 gnd 0.009888f
C1665 vdd.t81 gnd 0.12165f
C1666 vdd.t82 gnd 0.130011f
C1667 vdd.t80 gnd 0.158874f
C1668 vdd.n543 gnd 0.203654f
C1669 vdd.n544 gnd 0.171106f
C1670 vdd.n545 gnd 0.016236f
C1671 vdd.n546 gnd 0.009888f
C1672 vdd.n547 gnd 0.009888f
C1673 vdd.n548 gnd 0.009888f
C1674 vdd.n549 gnd 0.009888f
C1675 vdd.n550 gnd 0.009888f
C1676 vdd.n551 gnd 0.007959f
C1677 vdd.n552 gnd 0.009888f
C1678 vdd.n553 gnd 0.009888f
C1679 vdd.n554 gnd 0.009888f
C1680 vdd.n555 gnd 0.009888f
C1681 vdd.n556 gnd 0.009888f
C1682 vdd.n557 gnd 0.007959f
C1683 vdd.n558 gnd 0.009888f
C1684 vdd.n559 gnd 0.009888f
C1685 vdd.n560 gnd 0.009888f
C1686 vdd.n561 gnd 0.009888f
C1687 vdd.n562 gnd 0.009888f
C1688 vdd.n563 gnd 0.007959f
C1689 vdd.n564 gnd 0.009888f
C1690 vdd.n565 gnd 0.009888f
C1691 vdd.n566 gnd 0.009888f
C1692 vdd.n567 gnd 0.009888f
C1693 vdd.n568 gnd 0.009888f
C1694 vdd.n569 gnd 0.007959f
C1695 vdd.n570 gnd 0.009888f
C1696 vdd.n571 gnd 0.009888f
C1697 vdd.n572 gnd 0.009888f
C1698 vdd.n573 gnd 0.009888f
C1699 vdd.n574 gnd 0.009888f
C1700 vdd.n575 gnd 0.007959f
C1701 vdd.n576 gnd 0.009888f
C1702 vdd.n577 gnd 0.009888f
C1703 vdd.n578 gnd 0.009888f
C1704 vdd.n579 gnd 0.007879f
C1705 vdd.t78 gnd 0.12165f
C1706 vdd.t79 gnd 0.130011f
C1707 vdd.t76 gnd 0.158874f
C1708 vdd.n580 gnd 0.203654f
C1709 vdd.n581 gnd 0.171106f
C1710 vdd.n582 gnd 0.009888f
C1711 vdd.n583 gnd 0.007959f
C1712 vdd.n585 gnd 0.009888f
C1713 vdd.n587 gnd 0.009888f
C1714 vdd.n588 gnd 0.009888f
C1715 vdd.n589 gnd 0.007959f
C1716 vdd.n590 gnd 0.009888f
C1717 vdd.n591 gnd 0.009888f
C1718 vdd.n592 gnd 0.009888f
C1719 vdd.n593 gnd 0.009888f
C1720 vdd.n594 gnd 0.009888f
C1721 vdd.n595 gnd 0.007959f
C1722 vdd.n596 gnd 0.009888f
C1723 vdd.n597 gnd 0.009888f
C1724 vdd.n598 gnd 0.009888f
C1725 vdd.n599 gnd 0.009888f
C1726 vdd.n600 gnd 0.009888f
C1727 vdd.n601 gnd 0.007959f
C1728 vdd.n602 gnd 0.009888f
C1729 vdd.n603 gnd 0.009888f
C1730 vdd.n604 gnd 0.009888f
C1731 vdd.n605 gnd 0.006328f
C1732 vdd.n610 gnd 0.006724f
C1733 vdd.n611 gnd 0.006724f
C1734 vdd.n612 gnd 0.006724f
C1735 vdd.n613 gnd 6.96251f
C1736 vdd.n614 gnd 0.006724f
C1737 vdd.n615 gnd 0.006724f
C1738 vdd.n616 gnd 0.006724f
C1739 vdd.n618 gnd 0.006724f
C1740 vdd.n619 gnd 0.006724f
C1741 vdd.n621 gnd 0.006724f
C1742 vdd.n622 gnd 0.004895f
C1743 vdd.n624 gnd 0.006724f
C1744 vdd.t118 gnd 0.271714f
C1745 vdd.t117 gnd 0.278133f
C1746 vdd.t116 gnd 0.177385f
C1747 vdd.n625 gnd 0.095867f
C1748 vdd.n626 gnd 0.054379f
C1749 vdd.n627 gnd 0.00961f
C1750 vdd.n628 gnd 0.015715f
C1751 vdd.n630 gnd 0.006724f
C1752 vdd.n631 gnd 0.687156f
C1753 vdd.n632 gnd 0.014896f
C1754 vdd.n633 gnd 0.014896f
C1755 vdd.n634 gnd 0.006724f
C1756 vdd.n635 gnd 0.015955f
C1757 vdd.n636 gnd 0.006724f
C1758 vdd.n637 gnd 0.006724f
C1759 vdd.n638 gnd 0.006724f
C1760 vdd.n639 gnd 0.006724f
C1761 vdd.n640 gnd 0.006724f
C1762 vdd.n642 gnd 0.006724f
C1763 vdd.n643 gnd 0.006724f
C1764 vdd.n645 gnd 0.006724f
C1765 vdd.n646 gnd 0.006724f
C1766 vdd.n648 gnd 0.006724f
C1767 vdd.n649 gnd 0.006724f
C1768 vdd.n651 gnd 0.006724f
C1769 vdd.n652 gnd 0.006724f
C1770 vdd.n654 gnd 0.006724f
C1771 vdd.n655 gnd 0.006724f
C1772 vdd.n657 gnd 0.006724f
C1773 vdd.n658 gnd 0.004895f
C1774 vdd.n660 gnd 0.006724f
C1775 vdd.t111 gnd 0.271714f
C1776 vdd.t110 gnd 0.278133f
C1777 vdd.t108 gnd 0.177385f
C1778 vdd.n661 gnd 0.095867f
C1779 vdd.n662 gnd 0.054379f
C1780 vdd.n663 gnd 0.00961f
C1781 vdd.n664 gnd 0.006724f
C1782 vdd.n665 gnd 0.006724f
C1783 vdd.t109 gnd 0.343578f
C1784 vdd.n666 gnd 0.006724f
C1785 vdd.n667 gnd 0.006724f
C1786 vdd.n668 gnd 0.006724f
C1787 vdd.n669 gnd 0.006724f
C1788 vdd.n670 gnd 0.006724f
C1789 vdd.n671 gnd 0.687156f
C1790 vdd.n672 gnd 0.006724f
C1791 vdd.n673 gnd 0.006724f
C1792 vdd.n674 gnd 0.601262f
C1793 vdd.n675 gnd 0.006724f
C1794 vdd.n676 gnd 0.006724f
C1795 vdd.n677 gnd 0.005933f
C1796 vdd.n678 gnd 0.006724f
C1797 vdd.n679 gnd 0.606314f
C1798 vdd.n680 gnd 0.006724f
C1799 vdd.n681 gnd 0.006724f
C1800 vdd.n682 gnd 0.006724f
C1801 vdd.n683 gnd 0.006724f
C1802 vdd.n684 gnd 0.006724f
C1803 vdd.n685 gnd 0.687156f
C1804 vdd.n686 gnd 0.006724f
C1805 vdd.n687 gnd 0.006724f
C1806 vdd.t92 gnd 0.30821f
C1807 vdd.t178 gnd 0.080842f
C1808 vdd.n688 gnd 0.006724f
C1809 vdd.n689 gnd 0.006724f
C1810 vdd.n690 gnd 0.006724f
C1811 vdd.t45 gnd 0.343578f
C1812 vdd.n691 gnd 0.006724f
C1813 vdd.n692 gnd 0.006724f
C1814 vdd.n693 gnd 0.006724f
C1815 vdd.n694 gnd 0.006724f
C1816 vdd.n695 gnd 0.006724f
C1817 vdd.t199 gnd 0.343578f
C1818 vdd.n696 gnd 0.006724f
C1819 vdd.n697 gnd 0.006724f
C1820 vdd.n698 gnd 0.570946f
C1821 vdd.n699 gnd 0.006724f
C1822 vdd.n700 gnd 0.006724f
C1823 vdd.n701 gnd 0.006724f
C1824 vdd.n702 gnd 0.419367f
C1825 vdd.n703 gnd 0.006724f
C1826 vdd.n704 gnd 0.006724f
C1827 vdd.t3 gnd 0.343578f
C1828 vdd.n705 gnd 0.006724f
C1829 vdd.n706 gnd 0.006724f
C1830 vdd.n707 gnd 0.006724f
C1831 vdd.n708 gnd 0.570946f
C1832 vdd.n709 gnd 0.006724f
C1833 vdd.n710 gnd 0.006724f
C1834 vdd.t158 gnd 0.293052f
C1835 vdd.t152 gnd 0.267789f
C1836 vdd.n711 gnd 0.006724f
C1837 vdd.n712 gnd 0.006724f
C1838 vdd.n713 gnd 0.006724f
C1839 vdd.t226 gnd 0.343578f
C1840 vdd.n714 gnd 0.006724f
C1841 vdd.n715 gnd 0.006724f
C1842 vdd.t59 gnd 0.343578f
C1843 vdd.n716 gnd 0.006724f
C1844 vdd.n717 gnd 0.006724f
C1845 vdd.n718 gnd 0.006724f
C1846 vdd.t5 gnd 0.252631f
C1847 vdd.n719 gnd 0.006724f
C1848 vdd.n720 gnd 0.006724f
C1849 vdd.n721 gnd 0.586104f
C1850 vdd.n722 gnd 0.006724f
C1851 vdd.n723 gnd 0.006724f
C1852 vdd.n724 gnd 0.006724f
C1853 vdd.n725 gnd 0.687156f
C1854 vdd.n726 gnd 0.006724f
C1855 vdd.n727 gnd 0.006724f
C1856 vdd.t55 gnd 0.30821f
C1857 vdd.n728 gnd 0.434525f
C1858 vdd.n729 gnd 0.006724f
C1859 vdd.n730 gnd 0.006724f
C1860 vdd.n731 gnd 0.006724f
C1861 vdd.t69 gnd 0.343578f
C1862 vdd.n732 gnd 0.006724f
C1863 vdd.n733 gnd 0.006724f
C1864 vdd.n734 gnd 0.006724f
C1865 vdd.n735 gnd 0.006724f
C1866 vdd.n736 gnd 0.006724f
C1867 vdd.t66 gnd 0.687156f
C1868 vdd.n737 gnd 0.006724f
C1869 vdd.n738 gnd 0.006724f
C1870 vdd.t113 gnd 0.343578f
C1871 vdd.n739 gnd 0.006724f
C1872 vdd.n740 gnd 0.015955f
C1873 vdd.n741 gnd 0.015955f
C1874 vdd.t23 gnd 0.646735f
C1875 vdd.n742 gnd 0.014896f
C1876 vdd.n743 gnd 0.014896f
C1877 vdd.n744 gnd 0.015955f
C1878 vdd.n745 gnd 0.006724f
C1879 vdd.n746 gnd 0.006724f
C1880 vdd.t154 gnd 0.646735f
C1881 vdd.n764 gnd 0.015955f
C1882 vdd.n782 gnd 0.014896f
C1883 vdd.n783 gnd 0.006724f
C1884 vdd.n784 gnd 0.014896f
C1885 vdd.t132 gnd 0.271714f
C1886 vdd.t131 gnd 0.278133f
C1887 vdd.t130 gnd 0.177385f
C1888 vdd.n785 gnd 0.095867f
C1889 vdd.n786 gnd 0.054379f
C1890 vdd.n787 gnd 0.015715f
C1891 vdd.n788 gnd 0.006724f
C1892 vdd.t159 gnd 0.687156f
C1893 vdd.n789 gnd 0.014896f
C1894 vdd.n790 gnd 0.006724f
C1895 vdd.n791 gnd 0.015955f
C1896 vdd.n792 gnd 0.006724f
C1897 vdd.t107 gnd 0.271714f
C1898 vdd.t106 gnd 0.278133f
C1899 vdd.t104 gnd 0.177385f
C1900 vdd.n793 gnd 0.095867f
C1901 vdd.n794 gnd 0.054379f
C1902 vdd.n795 gnd 0.00961f
C1903 vdd.n796 gnd 0.006724f
C1904 vdd.n797 gnd 0.006724f
C1905 vdd.t105 gnd 0.343578f
C1906 vdd.n798 gnd 0.006724f
C1907 vdd.n799 gnd 0.006724f
C1908 vdd.n800 gnd 0.006724f
C1909 vdd.n801 gnd 0.006724f
C1910 vdd.n802 gnd 0.006724f
C1911 vdd.n803 gnd 0.006724f
C1912 vdd.n804 gnd 0.687156f
C1913 vdd.n805 gnd 0.006724f
C1914 vdd.n806 gnd 0.006724f
C1915 vdd.t197 gnd 0.343578f
C1916 vdd.n807 gnd 0.006724f
C1917 vdd.n808 gnd 0.006724f
C1918 vdd.n809 gnd 0.006724f
C1919 vdd.n810 gnd 0.006724f
C1920 vdd.n811 gnd 0.434525f
C1921 vdd.n812 gnd 0.006724f
C1922 vdd.n813 gnd 0.006724f
C1923 vdd.n814 gnd 0.006724f
C1924 vdd.n815 gnd 0.006724f
C1925 vdd.n816 gnd 0.006724f
C1926 vdd.n817 gnd 0.586104f
C1927 vdd.n818 gnd 0.006724f
C1928 vdd.n819 gnd 0.006724f
C1929 vdd.t43 gnd 0.30821f
C1930 vdd.t182 gnd 0.252631f
C1931 vdd.n820 gnd 0.006724f
C1932 vdd.n821 gnd 0.006724f
C1933 vdd.n822 gnd 0.006724f
C1934 vdd.t71 gnd 0.343578f
C1935 vdd.n823 gnd 0.006724f
C1936 vdd.n824 gnd 0.006724f
C1937 vdd.t28 gnd 0.343578f
C1938 vdd.n825 gnd 0.006724f
C1939 vdd.n826 gnd 0.006724f
C1940 vdd.n827 gnd 0.006724f
C1941 vdd.t57 gnd 0.267789f
C1942 vdd.n828 gnd 0.006724f
C1943 vdd.n829 gnd 0.006724f
C1944 vdd.n830 gnd 0.570946f
C1945 vdd.n831 gnd 0.006724f
C1946 vdd.n832 gnd 0.006724f
C1947 vdd.n833 gnd 0.006724f
C1948 vdd.t1 gnd 0.343578f
C1949 vdd.n834 gnd 0.006724f
C1950 vdd.n835 gnd 0.006724f
C1951 vdd.t0 gnd 0.293052f
C1952 vdd.n836 gnd 0.419367f
C1953 vdd.n837 gnd 0.006724f
C1954 vdd.n838 gnd 0.006724f
C1955 vdd.n839 gnd 0.006724f
C1956 vdd.n840 gnd 0.570946f
C1957 vdd.n841 gnd 0.006724f
C1958 vdd.n842 gnd 0.006724f
C1959 vdd.t181 gnd 0.343578f
C1960 vdd.n843 gnd 0.006724f
C1961 vdd.n844 gnd 0.006724f
C1962 vdd.n845 gnd 0.006724f
C1963 vdd.n846 gnd 0.687156f
C1964 vdd.n847 gnd 0.006724f
C1965 vdd.n848 gnd 0.006724f
C1966 vdd.t68 gnd 0.343578f
C1967 vdd.n849 gnd 0.006724f
C1968 vdd.n850 gnd 0.006724f
C1969 vdd.n851 gnd 0.006724f
C1970 vdd.t14 gnd 0.080842f
C1971 vdd.n852 gnd 0.006724f
C1972 vdd.n853 gnd 0.006724f
C1973 vdd.n854 gnd 0.006724f
C1974 vdd.t125 gnd 0.278133f
C1975 vdd.t123 gnd 0.177385f
C1976 vdd.t126 gnd 0.278133f
C1977 vdd.n855 gnd 0.156322f
C1978 vdd.n856 gnd 0.006724f
C1979 vdd.n857 gnd 0.006724f
C1980 vdd.n858 gnd 0.687156f
C1981 vdd.n859 gnd 0.006724f
C1982 vdd.n860 gnd 0.006724f
C1983 vdd.t124 gnd 0.30821f
C1984 vdd.n861 gnd 0.606314f
C1985 vdd.n862 gnd 0.006724f
C1986 vdd.n863 gnd 0.006724f
C1987 vdd.n864 gnd 0.006724f
C1988 vdd.n865 gnd 0.601262f
C1989 vdd.n866 gnd 0.006724f
C1990 vdd.n867 gnd 0.006724f
C1991 vdd.n868 gnd 0.006724f
C1992 vdd.n869 gnd 0.006724f
C1993 vdd.n870 gnd 0.006724f
C1994 vdd.n871 gnd 0.687156f
C1995 vdd.n872 gnd 0.006724f
C1996 vdd.n873 gnd 0.006724f
C1997 vdd.t120 gnd 0.343578f
C1998 vdd.n874 gnd 0.006724f
C1999 vdd.n875 gnd 0.015955f
C2000 vdd.n876 gnd 0.015955f
C2001 vdd.n877 gnd 6.96251f
C2002 vdd.n878 gnd 0.014896f
C2003 vdd.n879 gnd 0.014896f
C2004 vdd.n880 gnd 0.015955f
C2005 vdd.n881 gnd 0.006724f
C2006 vdd.n882 gnd 0.006724f
C2007 vdd.n883 gnd 0.006724f
C2008 vdd.n884 gnd 0.006724f
C2009 vdd.n885 gnd 0.006724f
C2010 vdd.n886 gnd 0.006724f
C2011 vdd.n887 gnd 0.006724f
C2012 vdd.n888 gnd 0.006724f
C2013 vdd.n890 gnd 0.006724f
C2014 vdd.n891 gnd 0.006724f
C2015 vdd.n892 gnd 0.006328f
C2016 vdd.n895 gnd 0.023667f
C2017 vdd.n896 gnd 0.007959f
C2018 vdd.n897 gnd 0.009888f
C2019 vdd.n899 gnd 0.009888f
C2020 vdd.n900 gnd 0.006606f
C2021 vdd.t84 gnd 0.505262f
C2022 vdd.n901 gnd 7.23535f
C2023 vdd.n902 gnd 0.009888f
C2024 vdd.n903 gnd 0.023667f
C2025 vdd.n904 gnd 0.007959f
C2026 vdd.n905 gnd 0.009888f
C2027 vdd.n906 gnd 0.007959f
C2028 vdd.n907 gnd 0.009888f
C2029 vdd.n908 gnd 1.01052f
C2030 vdd.n909 gnd 0.009888f
C2031 vdd.n910 gnd 0.007959f
C2032 vdd.n911 gnd 0.007959f
C2033 vdd.n912 gnd 0.009888f
C2034 vdd.n913 gnd 0.007959f
C2035 vdd.n914 gnd 0.009888f
C2036 vdd.t17 gnd 0.505262f
C2037 vdd.n915 gnd 0.009888f
C2038 vdd.n916 gnd 0.007959f
C2039 vdd.n917 gnd 0.009888f
C2040 vdd.n918 gnd 0.007959f
C2041 vdd.n919 gnd 0.009888f
C2042 vdd.t168 gnd 0.505262f
C2043 vdd.n920 gnd 0.009888f
C2044 vdd.n921 gnd 0.007959f
C2045 vdd.n922 gnd 0.009888f
C2046 vdd.n923 gnd 0.007959f
C2047 vdd.n924 gnd 0.009888f
C2048 vdd.t30 gnd 0.505262f
C2049 vdd.n925 gnd 0.793261f
C2050 vdd.n926 gnd 0.009888f
C2051 vdd.n927 gnd 0.007959f
C2052 vdd.n928 gnd 0.009888f
C2053 vdd.n929 gnd 0.007959f
C2054 vdd.n930 gnd 0.009888f
C2055 vdd.n931 gnd 0.712419f
C2056 vdd.n932 gnd 0.009888f
C2057 vdd.n933 gnd 0.007959f
C2058 vdd.n934 gnd 0.009888f
C2059 vdd.n935 gnd 0.007959f
C2060 vdd.n936 gnd 0.009888f
C2061 vdd.n937 gnd 0.54063f
C2062 vdd.t46 gnd 0.505262f
C2063 vdd.n938 gnd 0.009888f
C2064 vdd.n939 gnd 0.007959f
C2065 vdd.n940 gnd 0.009854f
C2066 vdd.n941 gnd 0.007959f
C2067 vdd.n942 gnd 0.009888f
C2068 vdd.t162 gnd 0.505262f
C2069 vdd.n943 gnd 0.009888f
C2070 vdd.n944 gnd 0.007959f
C2071 vdd.n945 gnd 0.009888f
C2072 vdd.n946 gnd 0.007959f
C2073 vdd.n947 gnd 0.009888f
C2074 vdd.t26 gnd 0.505262f
C2075 vdd.n948 gnd 0.641682f
C2076 vdd.n949 gnd 0.009888f
C2077 vdd.n950 gnd 0.007959f
C2078 vdd.n951 gnd 0.009888f
C2079 vdd.n952 gnd 0.007959f
C2080 vdd.n953 gnd 0.009888f
C2081 vdd.t50 gnd 0.505262f
C2082 vdd.n954 gnd 0.009888f
C2083 vdd.n955 gnd 0.007959f
C2084 vdd.n956 gnd 0.009888f
C2085 vdd.n957 gnd 0.007959f
C2086 vdd.n958 gnd 0.009888f
C2087 vdd.n959 gnd 0.692209f
C2088 vdd.n960 gnd 0.838735f
C2089 vdd.t36 gnd 0.505262f
C2090 vdd.n961 gnd 0.009888f
C2091 vdd.n962 gnd 0.007959f
C2092 vdd.n963 gnd 0.009888f
C2093 vdd.n964 gnd 0.007959f
C2094 vdd.n965 gnd 0.009888f
C2095 vdd.n966 gnd 0.52042f
C2096 vdd.n967 gnd 0.009888f
C2097 vdd.n968 gnd 0.007959f
C2098 vdd.n969 gnd 0.009888f
C2099 vdd.n970 gnd 0.007959f
C2100 vdd.n971 gnd 0.009888f
C2101 vdd.n972 gnd 1.01052f
C2102 vdd.t62 gnd 0.505262f
C2103 vdd.n973 gnd 0.009888f
C2104 vdd.n974 gnd 0.007959f
C2105 vdd.n975 gnd 0.009888f
C2106 vdd.n976 gnd 0.007959f
C2107 vdd.n977 gnd 0.009888f
C2108 vdd.t88 gnd 0.505262f
C2109 vdd.n978 gnd 0.009888f
C2110 vdd.n979 gnd 0.007959f
C2111 vdd.n980 gnd 0.023667f
C2112 vdd.n981 gnd 0.023667f
C2113 vdd.n982 gnd 2.3242f
C2114 vdd.n983 gnd 0.570946f
C2115 vdd.n984 gnd 0.023667f
C2116 vdd.n985 gnd 0.009888f
C2117 vdd.n987 gnd 0.009888f
C2118 vdd.n988 gnd 0.009888f
C2119 vdd.n989 gnd 0.007959f
C2120 vdd.n990 gnd 0.009888f
C2121 vdd.n991 gnd 0.009888f
C2122 vdd.n993 gnd 0.009888f
C2123 vdd.n994 gnd 0.009888f
C2124 vdd.n996 gnd 0.009888f
C2125 vdd.n997 gnd 0.007959f
C2126 vdd.n998 gnd 0.009888f
C2127 vdd.n999 gnd 0.009888f
C2128 vdd.n1001 gnd 0.009888f
C2129 vdd.n1002 gnd 0.009888f
C2130 vdd.n1004 gnd 0.009888f
C2131 vdd.n1005 gnd 0.007959f
C2132 vdd.n1006 gnd 0.009888f
C2133 vdd.n1007 gnd 0.009888f
C2134 vdd.n1009 gnd 0.009888f
C2135 vdd.n1010 gnd 0.009888f
C2136 vdd.n1012 gnd 0.009888f
C2137 vdd.n1013 gnd 0.007959f
C2138 vdd.n1014 gnd 0.009888f
C2139 vdd.n1015 gnd 0.009888f
C2140 vdd.n1017 gnd 0.009888f
C2141 vdd.n1018 gnd 0.009888f
C2142 vdd.n1020 gnd 0.009888f
C2143 vdd.t99 gnd 0.12165f
C2144 vdd.t100 gnd 0.130011f
C2145 vdd.t98 gnd 0.158874f
C2146 vdd.n1021 gnd 0.203654f
C2147 vdd.n1022 gnd 0.171902f
C2148 vdd.n1023 gnd 0.017032f
C2149 vdd.n1024 gnd 0.009888f
C2150 vdd.n1025 gnd 0.009888f
C2151 vdd.n1027 gnd 0.009888f
C2152 vdd.n1028 gnd 0.009888f
C2153 vdd.n1030 gnd 0.009888f
C2154 vdd.n1031 gnd 0.007959f
C2155 vdd.n1032 gnd 0.009888f
C2156 vdd.n1033 gnd 0.009888f
C2157 vdd.n1035 gnd 0.009888f
C2158 vdd.n1036 gnd 0.009888f
C2159 vdd.n1038 gnd 0.009888f
C2160 vdd.n1039 gnd 0.007959f
C2161 vdd.n1040 gnd 0.009888f
C2162 vdd.n1041 gnd 0.009888f
C2163 vdd.n1043 gnd 0.009888f
C2164 vdd.n1044 gnd 0.009888f
C2165 vdd.n1046 gnd 0.009888f
C2166 vdd.n1047 gnd 0.007959f
C2167 vdd.n1048 gnd 0.009888f
C2168 vdd.n1049 gnd 0.009888f
C2169 vdd.n1051 gnd 0.009888f
C2170 vdd.n1052 gnd 0.009888f
C2171 vdd.n1054 gnd 0.009888f
C2172 vdd.n1055 gnd 0.007959f
C2173 vdd.n1056 gnd 0.009888f
C2174 vdd.n1057 gnd 0.009888f
C2175 vdd.n1059 gnd 0.009888f
C2176 vdd.n1060 gnd 0.009888f
C2177 vdd.n1062 gnd 0.009888f
C2178 vdd.n1063 gnd 0.007959f
C2179 vdd.n1064 gnd 0.009888f
C2180 vdd.n1065 gnd 0.009888f
C2181 vdd.n1067 gnd 0.009888f
C2182 vdd.n1068 gnd 0.007879f
C2183 vdd.n1070 gnd 0.007959f
C2184 vdd.n1071 gnd 0.009888f
C2185 vdd.n1072 gnd 0.009888f
C2186 vdd.n1073 gnd 0.009888f
C2187 vdd.n1074 gnd 0.009888f
C2188 vdd.n1076 gnd 0.009888f
C2189 vdd.n1077 gnd 0.009888f
C2190 vdd.n1078 gnd 0.007959f
C2191 vdd.n1079 gnd 0.009888f
C2192 vdd.n1081 gnd 0.009888f
C2193 vdd.n1082 gnd 0.009888f
C2194 vdd.n1084 gnd 0.009888f
C2195 vdd.n1085 gnd 0.009888f
C2196 vdd.n1086 gnd 0.007959f
C2197 vdd.n1087 gnd 0.009888f
C2198 vdd.n1089 gnd 0.009888f
C2199 vdd.n1090 gnd 0.009888f
C2200 vdd.n1092 gnd 0.009888f
C2201 vdd.n1093 gnd 0.009888f
C2202 vdd.n1094 gnd 0.007959f
C2203 vdd.n1095 gnd 0.009888f
C2204 vdd.n1097 gnd 0.009888f
C2205 vdd.n1098 gnd 0.009888f
C2206 vdd.n1100 gnd 0.009888f
C2207 vdd.n1101 gnd 0.009888f
C2208 vdd.n1102 gnd 0.007959f
C2209 vdd.n1103 gnd 0.009888f
C2210 vdd.n1105 gnd 0.009888f
C2211 vdd.n1106 gnd 0.009888f
C2212 vdd.n1108 gnd 0.009888f
C2213 vdd.n1109 gnd 0.00378f
C2214 vdd.t141 gnd 0.12165f
C2215 vdd.t142 gnd 0.130011f
C2216 vdd.t140 gnd 0.158874f
C2217 vdd.n1110 gnd 0.203654f
C2218 vdd.n1111 gnd 0.171902f
C2219 vdd.n1112 gnd 0.013052f
C2220 vdd.n1113 gnd 0.004178f
C2221 vdd.n1114 gnd 0.007959f
C2222 vdd.n1115 gnd 0.009888f
C2223 vdd.n1116 gnd 0.009888f
C2224 vdd.n1117 gnd 0.009888f
C2225 vdd.n1118 gnd 0.007959f
C2226 vdd.n1119 gnd 0.007959f
C2227 vdd.n1120 gnd 0.007959f
C2228 vdd.n1121 gnd 0.009888f
C2229 vdd.n1122 gnd 0.009888f
C2230 vdd.n1123 gnd 0.009888f
C2231 vdd.n1124 gnd 0.007959f
C2232 vdd.n1125 gnd 0.007959f
C2233 vdd.n1126 gnd 0.007959f
C2234 vdd.n1127 gnd 0.009888f
C2235 vdd.n1128 gnd 0.009888f
C2236 vdd.n1129 gnd 0.009888f
C2237 vdd.n1130 gnd 0.007959f
C2238 vdd.n1131 gnd 0.007959f
C2239 vdd.n1132 gnd 0.007959f
C2240 vdd.n1133 gnd 0.009888f
C2241 vdd.n1134 gnd 0.009888f
C2242 vdd.n1135 gnd 0.009888f
C2243 vdd.n1136 gnd 0.007959f
C2244 vdd.n1137 gnd 0.007959f
C2245 vdd.n1138 gnd 0.007959f
C2246 vdd.n1139 gnd 0.009888f
C2247 vdd.n1140 gnd 0.009888f
C2248 vdd.n1141 gnd 0.009888f
C2249 vdd.n1142 gnd 0.007959f
C2250 vdd.n1143 gnd 0.009888f
C2251 vdd.n1144 gnd 0.009888f
C2252 vdd.n1146 gnd 0.009888f
C2253 vdd.t89 gnd 0.12165f
C2254 vdd.t90 gnd 0.130011f
C2255 vdd.t87 gnd 0.158874f
C2256 vdd.n1147 gnd 0.203654f
C2257 vdd.n1148 gnd 0.171902f
C2258 vdd.n1149 gnd 0.017032f
C2259 vdd.n1150 gnd 0.005412f
C2260 vdd.n1151 gnd 0.009888f
C2261 vdd.n1152 gnd 0.009888f
C2262 vdd.n1153 gnd 0.009888f
C2263 vdd.n1154 gnd 0.007959f
C2264 vdd.n1155 gnd 0.007959f
C2265 vdd.n1156 gnd 0.007959f
C2266 vdd.n1157 gnd 0.009888f
C2267 vdd.n1158 gnd 0.009888f
C2268 vdd.n1159 gnd 0.009888f
C2269 vdd.n1160 gnd 0.007959f
C2270 vdd.n1161 gnd 0.007959f
C2271 vdd.n1162 gnd 0.007959f
C2272 vdd.n1163 gnd 0.009888f
C2273 vdd.n1164 gnd 0.009888f
C2274 vdd.n1165 gnd 0.009888f
C2275 vdd.n1166 gnd 0.007959f
C2276 vdd.n1167 gnd 0.007959f
C2277 vdd.n1168 gnd 0.007959f
C2278 vdd.n1169 gnd 0.009888f
C2279 vdd.n1170 gnd 0.009888f
C2280 vdd.n1171 gnd 0.009888f
C2281 vdd.n1172 gnd 0.007959f
C2282 vdd.n1173 gnd 0.007959f
C2283 vdd.n1174 gnd 0.007959f
C2284 vdd.n1175 gnd 0.009888f
C2285 vdd.n1176 gnd 0.009888f
C2286 vdd.n1177 gnd 0.009888f
C2287 vdd.n1178 gnd 0.007959f
C2288 vdd.n1179 gnd 0.007959f
C2289 vdd.n1180 gnd 0.006646f
C2290 vdd.n1181 gnd 0.009888f
C2291 vdd.n1182 gnd 0.009888f
C2292 vdd.n1183 gnd 0.009888f
C2293 vdd.n1184 gnd 0.006646f
C2294 vdd.n1185 gnd 0.007959f
C2295 vdd.n1186 gnd 0.007959f
C2296 vdd.n1187 gnd 0.009888f
C2297 vdd.n1188 gnd 0.009888f
C2298 vdd.n1189 gnd 0.009888f
C2299 vdd.n1190 gnd 0.007959f
C2300 vdd.n1191 gnd 0.007959f
C2301 vdd.n1192 gnd 0.007959f
C2302 vdd.n1193 gnd 0.009888f
C2303 vdd.n1194 gnd 0.009888f
C2304 vdd.n1195 gnd 0.009888f
C2305 vdd.n1196 gnd 0.007959f
C2306 vdd.n1197 gnd 0.007959f
C2307 vdd.n1198 gnd 0.007959f
C2308 vdd.n1199 gnd 0.009888f
C2309 vdd.n1200 gnd 0.009888f
C2310 vdd.n1201 gnd 0.009888f
C2311 vdd.n1202 gnd 0.007959f
C2312 vdd.n1203 gnd 0.007959f
C2313 vdd.n1204 gnd 0.007959f
C2314 vdd.n1205 gnd 0.009888f
C2315 vdd.n1206 gnd 0.009888f
C2316 vdd.n1207 gnd 0.009888f
C2317 vdd.n1208 gnd 0.007959f
C2318 vdd.n1209 gnd 0.007959f
C2319 vdd.n1210 gnd 0.006606f
C2320 vdd.n1211 gnd 0.023667f
C2321 vdd.n1212 gnd 0.023302f
C2322 vdd.n1213 gnd 0.006606f
C2323 vdd.n1214 gnd 0.023302f
C2324 vdd.n1215 gnd 1.42484f
C2325 vdd.n1216 gnd 0.023302f
C2326 vdd.n1217 gnd 0.006606f
C2327 vdd.n1218 gnd 0.023302f
C2328 vdd.n1219 gnd 0.009888f
C2329 vdd.n1220 gnd 0.009888f
C2330 vdd.n1221 gnd 0.007959f
C2331 vdd.n1222 gnd 0.009888f
C2332 vdd.n1223 gnd 0.94484f
C2333 vdd.n1224 gnd 0.009888f
C2334 vdd.n1225 gnd 0.007959f
C2335 vdd.n1226 gnd 0.009888f
C2336 vdd.n1227 gnd 0.009888f
C2337 vdd.n1228 gnd 0.009888f
C2338 vdd.n1229 gnd 0.007959f
C2339 vdd.n1230 gnd 0.009888f
C2340 vdd.n1231 gnd 0.995366f
C2341 vdd.n1232 gnd 0.009888f
C2342 vdd.n1233 gnd 0.007959f
C2343 vdd.n1234 gnd 0.009888f
C2344 vdd.n1235 gnd 0.009888f
C2345 vdd.n1236 gnd 0.009888f
C2346 vdd.n1237 gnd 0.007959f
C2347 vdd.n1238 gnd 0.009888f
C2348 vdd.t186 gnd 0.505262f
C2349 vdd.n1239 gnd 0.823577f
C2350 vdd.n1240 gnd 0.009888f
C2351 vdd.n1241 gnd 0.007959f
C2352 vdd.n1242 gnd 0.009888f
C2353 vdd.n1243 gnd 0.009888f
C2354 vdd.n1244 gnd 0.009888f
C2355 vdd.n1245 gnd 0.007959f
C2356 vdd.n1246 gnd 0.009888f
C2357 vdd.n1247 gnd 0.651788f
C2358 vdd.n1248 gnd 0.009888f
C2359 vdd.n1249 gnd 0.007959f
C2360 vdd.n1250 gnd 0.009888f
C2361 vdd.n1251 gnd 0.009888f
C2362 vdd.n1252 gnd 0.009888f
C2363 vdd.n1253 gnd 0.007959f
C2364 vdd.n1254 gnd 0.009888f
C2365 vdd.n1255 gnd 0.813471f
C2366 vdd.n1256 gnd 0.530525f
C2367 vdd.n1257 gnd 0.009888f
C2368 vdd.n1258 gnd 0.007959f
C2369 vdd.n1259 gnd 0.009888f
C2370 vdd.n1260 gnd 0.009888f
C2371 vdd.n1261 gnd 0.009888f
C2372 vdd.n1262 gnd 0.007959f
C2373 vdd.n1263 gnd 0.009888f
C2374 vdd.n1264 gnd 0.702314f
C2375 vdd.n1265 gnd 0.009888f
C2376 vdd.n1266 gnd 0.007959f
C2377 vdd.n1267 gnd 0.009888f
C2378 vdd.n1268 gnd 0.009888f
C2379 vdd.n1269 gnd 0.009888f
C2380 vdd.n1270 gnd 0.007959f
C2381 vdd.n1271 gnd 0.009888f
C2382 vdd.t8 gnd 0.505262f
C2383 vdd.n1272 gnd 0.838735f
C2384 vdd.n1273 gnd 0.009888f
C2385 vdd.n1274 gnd 0.007959f
C2386 vdd.n1275 gnd 0.005427f
C2387 vdd.n1276 gnd 0.005036f
C2388 vdd.n1277 gnd 0.002786f
C2389 vdd.n1278 gnd 0.006396f
C2390 vdd.n1279 gnd 0.002706f
C2391 vdd.n1280 gnd 0.002865f
C2392 vdd.n1281 gnd 0.005036f
C2393 vdd.n1282 gnd 0.002706f
C2394 vdd.n1283 gnd 0.006396f
C2395 vdd.n1284 gnd 0.002865f
C2396 vdd.n1285 gnd 0.005036f
C2397 vdd.n1286 gnd 0.002706f
C2398 vdd.n1287 gnd 0.004797f
C2399 vdd.n1288 gnd 0.004811f
C2400 vdd.t18 gnd 0.013741f
C2401 vdd.n1289 gnd 0.030574f
C2402 vdd.n1290 gnd 0.159114f
C2403 vdd.n1291 gnd 0.002706f
C2404 vdd.n1292 gnd 0.002865f
C2405 vdd.n1293 gnd 0.006396f
C2406 vdd.n1294 gnd 0.006396f
C2407 vdd.n1295 gnd 0.002865f
C2408 vdd.n1296 gnd 0.002706f
C2409 vdd.n1297 gnd 0.005036f
C2410 vdd.n1298 gnd 0.005036f
C2411 vdd.n1299 gnd 0.002706f
C2412 vdd.n1300 gnd 0.002865f
C2413 vdd.n1301 gnd 0.006396f
C2414 vdd.n1302 gnd 0.006396f
C2415 vdd.n1303 gnd 0.002865f
C2416 vdd.n1304 gnd 0.002706f
C2417 vdd.n1305 gnd 0.005036f
C2418 vdd.n1306 gnd 0.005036f
C2419 vdd.n1307 gnd 0.002706f
C2420 vdd.n1308 gnd 0.002865f
C2421 vdd.n1309 gnd 0.006396f
C2422 vdd.n1310 gnd 0.006396f
C2423 vdd.n1311 gnd 0.015121f
C2424 vdd.n1312 gnd 0.002786f
C2425 vdd.n1313 gnd 0.002706f
C2426 vdd.n1314 gnd 0.013016f
C2427 vdd.n1315 gnd 0.009087f
C2428 vdd.t31 gnd 0.031835f
C2429 vdd.t169 gnd 0.031835f
C2430 vdd.n1316 gnd 0.218793f
C2431 vdd.n1317 gnd 0.172047f
C2432 vdd.t47 gnd 0.031835f
C2433 vdd.t22 gnd 0.031835f
C2434 vdd.n1318 gnd 0.218793f
C2435 vdd.n1319 gnd 0.138841f
C2436 vdd.t206 gnd 0.031835f
C2437 vdd.t193 gnd 0.031835f
C2438 vdd.n1320 gnd 0.218793f
C2439 vdd.n1321 gnd 0.138841f
C2440 vdd.t51 gnd 0.031835f
C2441 vdd.t171 gnd 0.031835f
C2442 vdd.n1322 gnd 0.218793f
C2443 vdd.n1323 gnd 0.138841f
C2444 vdd.t187 gnd 0.031835f
C2445 vdd.t37 gnd 0.031835f
C2446 vdd.n1324 gnd 0.218793f
C2447 vdd.n1325 gnd 0.138841f
C2448 vdd.n1326 gnd 0.005427f
C2449 vdd.n1327 gnd 0.005036f
C2450 vdd.n1328 gnd 0.002786f
C2451 vdd.n1329 gnd 0.006396f
C2452 vdd.n1330 gnd 0.002706f
C2453 vdd.n1331 gnd 0.002865f
C2454 vdd.n1332 gnd 0.005036f
C2455 vdd.n1333 gnd 0.002706f
C2456 vdd.n1334 gnd 0.006396f
C2457 vdd.n1335 gnd 0.002865f
C2458 vdd.n1336 gnd 0.005036f
C2459 vdd.n1337 gnd 0.002706f
C2460 vdd.n1338 gnd 0.004797f
C2461 vdd.n1339 gnd 0.004811f
C2462 vdd.t63 gnd 0.013741f
C2463 vdd.n1340 gnd 0.030574f
C2464 vdd.n1341 gnd 0.159114f
C2465 vdd.n1342 gnd 0.002706f
C2466 vdd.n1343 gnd 0.002865f
C2467 vdd.n1344 gnd 0.006396f
C2468 vdd.n1345 gnd 0.006396f
C2469 vdd.n1346 gnd 0.002865f
C2470 vdd.n1347 gnd 0.002706f
C2471 vdd.n1348 gnd 0.005036f
C2472 vdd.n1349 gnd 0.005036f
C2473 vdd.n1350 gnd 0.002706f
C2474 vdd.n1351 gnd 0.002865f
C2475 vdd.n1352 gnd 0.006396f
C2476 vdd.n1353 gnd 0.006396f
C2477 vdd.n1354 gnd 0.002865f
C2478 vdd.n1355 gnd 0.002706f
C2479 vdd.n1356 gnd 0.005036f
C2480 vdd.n1357 gnd 0.005036f
C2481 vdd.n1358 gnd 0.002706f
C2482 vdd.n1359 gnd 0.002865f
C2483 vdd.n1360 gnd 0.006396f
C2484 vdd.n1361 gnd 0.006396f
C2485 vdd.n1362 gnd 0.015121f
C2486 vdd.n1363 gnd 0.002786f
C2487 vdd.n1364 gnd 0.002706f
C2488 vdd.n1365 gnd 0.013016f
C2489 vdd.n1366 gnd 0.008802f
C2490 vdd.n1367 gnd 0.103298f
C2491 vdd.n1368 gnd 0.005427f
C2492 vdd.n1369 gnd 0.005036f
C2493 vdd.n1370 gnd 0.002786f
C2494 vdd.n1371 gnd 0.006396f
C2495 vdd.n1372 gnd 0.002706f
C2496 vdd.n1373 gnd 0.002865f
C2497 vdd.n1374 gnd 0.005036f
C2498 vdd.n1375 gnd 0.002706f
C2499 vdd.n1376 gnd 0.006396f
C2500 vdd.n1377 gnd 0.002865f
C2501 vdd.n1378 gnd 0.005036f
C2502 vdd.n1379 gnd 0.002706f
C2503 vdd.n1380 gnd 0.004797f
C2504 vdd.n1381 gnd 0.004811f
C2505 vdd.t54 gnd 0.013741f
C2506 vdd.n1382 gnd 0.030574f
C2507 vdd.n1383 gnd 0.159114f
C2508 vdd.n1384 gnd 0.002706f
C2509 vdd.n1385 gnd 0.002865f
C2510 vdd.n1386 gnd 0.006396f
C2511 vdd.n1387 gnd 0.006396f
C2512 vdd.n1388 gnd 0.002865f
C2513 vdd.n1389 gnd 0.002706f
C2514 vdd.n1390 gnd 0.005036f
C2515 vdd.n1391 gnd 0.005036f
C2516 vdd.n1392 gnd 0.002706f
C2517 vdd.n1393 gnd 0.002865f
C2518 vdd.n1394 gnd 0.006396f
C2519 vdd.n1395 gnd 0.006396f
C2520 vdd.n1396 gnd 0.002865f
C2521 vdd.n1397 gnd 0.002706f
C2522 vdd.n1398 gnd 0.005036f
C2523 vdd.n1399 gnd 0.005036f
C2524 vdd.n1400 gnd 0.002706f
C2525 vdd.n1401 gnd 0.002865f
C2526 vdd.n1402 gnd 0.006396f
C2527 vdd.n1403 gnd 0.006396f
C2528 vdd.n1404 gnd 0.015121f
C2529 vdd.n1405 gnd 0.002786f
C2530 vdd.n1406 gnd 0.002706f
C2531 vdd.n1407 gnd 0.013016f
C2532 vdd.n1408 gnd 0.009087f
C2533 vdd.t39 gnd 0.031835f
C2534 vdd.t177 gnd 0.031835f
C2535 vdd.n1409 gnd 0.218793f
C2536 vdd.n1410 gnd 0.172047f
C2537 vdd.t194 gnd 0.031835f
C2538 vdd.t74 gnd 0.031835f
C2539 vdd.n1411 gnd 0.218793f
C2540 vdd.n1412 gnd 0.138841f
C2541 vdd.t163 gnd 0.031835f
C2542 vdd.t9 gnd 0.031835f
C2543 vdd.n1413 gnd 0.218793f
C2544 vdd.n1414 gnd 0.138841f
C2545 vdd.t196 gnd 0.031835f
C2546 vdd.t75 gnd 0.031835f
C2547 vdd.n1415 gnd 0.218793f
C2548 vdd.n1416 gnd 0.138841f
C2549 vdd.t189 gnd 0.031835f
C2550 vdd.t179 gnd 0.031835f
C2551 vdd.n1417 gnd 0.218793f
C2552 vdd.n1418 gnd 0.138841f
C2553 vdd.n1419 gnd 0.005427f
C2554 vdd.n1420 gnd 0.005036f
C2555 vdd.n1421 gnd 0.002786f
C2556 vdd.n1422 gnd 0.006396f
C2557 vdd.n1423 gnd 0.002706f
C2558 vdd.n1424 gnd 0.002865f
C2559 vdd.n1425 gnd 0.005036f
C2560 vdd.n1426 gnd 0.002706f
C2561 vdd.n1427 gnd 0.006396f
C2562 vdd.n1428 gnd 0.002865f
C2563 vdd.n1429 gnd 0.005036f
C2564 vdd.n1430 gnd 0.002706f
C2565 vdd.n1431 gnd 0.004797f
C2566 vdd.n1432 gnd 0.004811f
C2567 vdd.t188 gnd 0.013741f
C2568 vdd.n1433 gnd 0.030574f
C2569 vdd.n1434 gnd 0.159114f
C2570 vdd.n1435 gnd 0.002706f
C2571 vdd.n1436 gnd 0.002865f
C2572 vdd.n1437 gnd 0.006396f
C2573 vdd.n1438 gnd 0.006396f
C2574 vdd.n1439 gnd 0.002865f
C2575 vdd.n1440 gnd 0.002706f
C2576 vdd.n1441 gnd 0.005036f
C2577 vdd.n1442 gnd 0.005036f
C2578 vdd.n1443 gnd 0.002706f
C2579 vdd.n1444 gnd 0.002865f
C2580 vdd.n1445 gnd 0.006396f
C2581 vdd.n1446 gnd 0.006396f
C2582 vdd.n1447 gnd 0.002865f
C2583 vdd.n1448 gnd 0.002706f
C2584 vdd.n1449 gnd 0.005036f
C2585 vdd.n1450 gnd 0.005036f
C2586 vdd.n1451 gnd 0.002706f
C2587 vdd.n1452 gnd 0.002865f
C2588 vdd.n1453 gnd 0.006396f
C2589 vdd.n1454 gnd 0.006396f
C2590 vdd.n1455 gnd 0.015121f
C2591 vdd.n1456 gnd 0.002786f
C2592 vdd.n1457 gnd 0.002706f
C2593 vdd.n1458 gnd 0.013016f
C2594 vdd.n1459 gnd 0.008802f
C2595 vdd.n1460 gnd 0.061452f
C2596 vdd.n1461 gnd 0.221428f
C2597 vdd.n1462 gnd 0.005427f
C2598 vdd.n1463 gnd 0.005036f
C2599 vdd.n1464 gnd 0.002786f
C2600 vdd.n1465 gnd 0.006396f
C2601 vdd.n1466 gnd 0.002706f
C2602 vdd.n1467 gnd 0.002865f
C2603 vdd.n1468 gnd 0.005036f
C2604 vdd.n1469 gnd 0.002706f
C2605 vdd.n1470 gnd 0.006396f
C2606 vdd.n1471 gnd 0.002865f
C2607 vdd.n1472 gnd 0.005036f
C2608 vdd.n1473 gnd 0.002706f
C2609 vdd.n1474 gnd 0.004797f
C2610 vdd.n1475 gnd 0.004811f
C2611 vdd.t208 gnd 0.013741f
C2612 vdd.n1476 gnd 0.030574f
C2613 vdd.n1477 gnd 0.159114f
C2614 vdd.n1478 gnd 0.002706f
C2615 vdd.n1479 gnd 0.002865f
C2616 vdd.n1480 gnd 0.006396f
C2617 vdd.n1481 gnd 0.006396f
C2618 vdd.n1482 gnd 0.002865f
C2619 vdd.n1483 gnd 0.002706f
C2620 vdd.n1484 gnd 0.005036f
C2621 vdd.n1485 gnd 0.005036f
C2622 vdd.n1486 gnd 0.002706f
C2623 vdd.n1487 gnd 0.002865f
C2624 vdd.n1488 gnd 0.006396f
C2625 vdd.n1489 gnd 0.006396f
C2626 vdd.n1490 gnd 0.002865f
C2627 vdd.n1491 gnd 0.002706f
C2628 vdd.n1492 gnd 0.005036f
C2629 vdd.n1493 gnd 0.005036f
C2630 vdd.n1494 gnd 0.002706f
C2631 vdd.n1495 gnd 0.002865f
C2632 vdd.n1496 gnd 0.006396f
C2633 vdd.n1497 gnd 0.006396f
C2634 vdd.n1498 gnd 0.015121f
C2635 vdd.n1499 gnd 0.002786f
C2636 vdd.n1500 gnd 0.002706f
C2637 vdd.n1501 gnd 0.013016f
C2638 vdd.n1502 gnd 0.009087f
C2639 vdd.t48 gnd 0.031835f
C2640 vdd.t209 gnd 0.031835f
C2641 vdd.n1503 gnd 0.218793f
C2642 vdd.n1504 gnd 0.172047f
C2643 vdd.t195 gnd 0.031835f
C2644 vdd.t25 gnd 0.031835f
C2645 vdd.n1505 gnd 0.218793f
C2646 vdd.n1506 gnd 0.138841f
C2647 vdd.t230 gnd 0.031835f
C2648 vdd.t184 gnd 0.031835f
C2649 vdd.n1507 gnd 0.218793f
C2650 vdd.n1508 gnd 0.138841f
C2651 vdd.t175 gnd 0.031835f
C2652 vdd.t27 gnd 0.031835f
C2653 vdd.n1509 gnd 0.218793f
C2654 vdd.n1510 gnd 0.138841f
C2655 vdd.t201 gnd 0.031835f
C2656 vdd.t65 gnd 0.031835f
C2657 vdd.n1511 gnd 0.218793f
C2658 vdd.n1512 gnd 0.138841f
C2659 vdd.n1513 gnd 0.005427f
C2660 vdd.n1514 gnd 0.005036f
C2661 vdd.n1515 gnd 0.002786f
C2662 vdd.n1516 gnd 0.006396f
C2663 vdd.n1517 gnd 0.002706f
C2664 vdd.n1518 gnd 0.002865f
C2665 vdd.n1519 gnd 0.005036f
C2666 vdd.n1520 gnd 0.002706f
C2667 vdd.n1521 gnd 0.006396f
C2668 vdd.n1522 gnd 0.002865f
C2669 vdd.n1523 gnd 0.005036f
C2670 vdd.n1524 gnd 0.002706f
C2671 vdd.n1525 gnd 0.004797f
C2672 vdd.n1526 gnd 0.004811f
C2673 vdd.t200 gnd 0.013741f
C2674 vdd.n1527 gnd 0.030574f
C2675 vdd.n1528 gnd 0.159114f
C2676 vdd.n1529 gnd 0.002706f
C2677 vdd.n1530 gnd 0.002865f
C2678 vdd.n1531 gnd 0.006396f
C2679 vdd.n1532 gnd 0.006396f
C2680 vdd.n1533 gnd 0.002865f
C2681 vdd.n1534 gnd 0.002706f
C2682 vdd.n1535 gnd 0.005036f
C2683 vdd.n1536 gnd 0.005036f
C2684 vdd.n1537 gnd 0.002706f
C2685 vdd.n1538 gnd 0.002865f
C2686 vdd.n1539 gnd 0.006396f
C2687 vdd.n1540 gnd 0.006396f
C2688 vdd.n1541 gnd 0.002865f
C2689 vdd.n1542 gnd 0.002706f
C2690 vdd.n1543 gnd 0.005036f
C2691 vdd.n1544 gnd 0.005036f
C2692 vdd.n1545 gnd 0.002706f
C2693 vdd.n1546 gnd 0.002865f
C2694 vdd.n1547 gnd 0.006396f
C2695 vdd.n1548 gnd 0.006396f
C2696 vdd.n1549 gnd 0.015121f
C2697 vdd.n1550 gnd 0.002786f
C2698 vdd.n1551 gnd 0.002706f
C2699 vdd.n1552 gnd 0.013016f
C2700 vdd.n1553 gnd 0.008802f
C2701 vdd.n1554 gnd 0.061452f
C2702 vdd.n1555 gnd 0.243357f
C2703 vdd.n1556 gnd 2.19025f
C2704 vdd.n1557 gnd 0.588621f
C2705 vdd.n1558 gnd 0.009854f
C2706 vdd.n1559 gnd 0.009888f
C2707 vdd.n1560 gnd 0.007959f
C2708 vdd.n1561 gnd 0.009888f
C2709 vdd.n1562 gnd 0.803366f
C2710 vdd.n1563 gnd 0.009888f
C2711 vdd.n1564 gnd 0.007959f
C2712 vdd.n1565 gnd 0.009888f
C2713 vdd.n1566 gnd 0.009888f
C2714 vdd.n1567 gnd 0.009888f
C2715 vdd.n1568 gnd 0.007959f
C2716 vdd.n1569 gnd 0.009888f
C2717 vdd.n1570 gnd 0.838735f
C2718 vdd.t21 gnd 0.505262f
C2719 vdd.n1571 gnd 0.631577f
C2720 vdd.n1572 gnd 0.009888f
C2721 vdd.n1573 gnd 0.007959f
C2722 vdd.n1574 gnd 0.009888f
C2723 vdd.n1575 gnd 0.009888f
C2724 vdd.n1576 gnd 0.009888f
C2725 vdd.n1577 gnd 0.007959f
C2726 vdd.n1578 gnd 0.009888f
C2727 vdd.n1579 gnd 0.550735f
C2728 vdd.n1580 gnd 0.009888f
C2729 vdd.n1581 gnd 0.007959f
C2730 vdd.n1582 gnd 0.009888f
C2731 vdd.n1583 gnd 0.009888f
C2732 vdd.n1584 gnd 0.009888f
C2733 vdd.n1585 gnd 0.007959f
C2734 vdd.n1586 gnd 0.009888f
C2735 vdd.n1587 gnd 0.621472f
C2736 vdd.n1588 gnd 0.722524f
C2737 vdd.n1589 gnd 0.009888f
C2738 vdd.n1590 gnd 0.007959f
C2739 vdd.n1591 gnd 0.009888f
C2740 vdd.n1592 gnd 0.009888f
C2741 vdd.n1593 gnd 0.009888f
C2742 vdd.n1594 gnd 0.007959f
C2743 vdd.n1595 gnd 0.009888f
C2744 vdd.n1596 gnd 0.894313f
C2745 vdd.n1597 gnd 0.009888f
C2746 vdd.n1598 gnd 0.007959f
C2747 vdd.n1599 gnd 0.009888f
C2748 vdd.n1600 gnd 0.009888f
C2749 vdd.n1601 gnd 0.023302f
C2750 vdd.n1602 gnd 0.009888f
C2751 vdd.n1603 gnd 0.009888f
C2752 vdd.n1604 gnd 0.007959f
C2753 vdd.n1605 gnd 0.009888f
C2754 vdd.n1606 gnd 0.54063f
C2755 vdd.n1607 gnd 1.01052f
C2756 vdd.n1608 gnd 0.009888f
C2757 vdd.n1609 gnd 0.007959f
C2758 vdd.n1610 gnd 0.009888f
C2759 vdd.n1611 gnd 0.009888f
C2760 vdd.n1612 gnd 0.008504f
C2761 vdd.n1613 gnd 0.007959f
C2762 vdd.n1615 gnd 0.009888f
C2763 vdd.n1617 gnd 0.007959f
C2764 vdd.n1618 gnd 0.009888f
C2765 vdd.n1619 gnd 0.007959f
C2766 vdd.n1621 gnd 0.009888f
C2767 vdd.n1622 gnd 0.007959f
C2768 vdd.n1623 gnd 0.009888f
C2769 vdd.n1624 gnd 0.009888f
C2770 vdd.n1625 gnd 0.009888f
C2771 vdd.n1626 gnd 0.009888f
C2772 vdd.n1627 gnd 0.009888f
C2773 vdd.n1628 gnd 0.007959f
C2774 vdd.n1630 gnd 0.009888f
C2775 vdd.n1631 gnd 0.009888f
C2776 vdd.n1632 gnd 0.009888f
C2777 vdd.n1633 gnd 0.009888f
C2778 vdd.n1634 gnd 0.009888f
C2779 vdd.n1635 gnd 0.007959f
C2780 vdd.n1637 gnd 0.009888f
C2781 vdd.n1638 gnd 0.009888f
C2782 vdd.n1639 gnd 0.009888f
C2783 vdd.n1640 gnd 0.009888f
C2784 vdd.n1641 gnd 0.006646f
C2785 vdd.t103 gnd 0.12165f
C2786 vdd.t102 gnd 0.130011f
C2787 vdd.t101 gnd 0.158874f
C2788 vdd.n1642 gnd 0.203654f
C2789 vdd.n1643 gnd 0.171106f
C2790 vdd.n1645 gnd 0.009888f
C2791 vdd.n1646 gnd 0.009888f
C2792 vdd.n1647 gnd 0.007959f
C2793 vdd.n1648 gnd 0.009888f
C2794 vdd.n1650 gnd 0.009888f
C2795 vdd.n1651 gnd 0.009888f
C2796 vdd.n1652 gnd 0.009888f
C2797 vdd.n1653 gnd 0.009888f
C2798 vdd.n1654 gnd 0.007959f
C2799 vdd.n1656 gnd 0.009888f
C2800 vdd.n1657 gnd 0.009888f
C2801 vdd.n1658 gnd 0.009888f
C2802 vdd.n1659 gnd 0.009888f
C2803 vdd.n1660 gnd 0.009888f
C2804 vdd.n1661 gnd 0.007959f
C2805 vdd.n1663 gnd 0.009888f
C2806 vdd.n1664 gnd 0.009888f
C2807 vdd.n1665 gnd 0.009888f
C2808 vdd.n1666 gnd 0.009888f
C2809 vdd.n1667 gnd 0.009888f
C2810 vdd.n1668 gnd 0.007959f
C2811 vdd.n1670 gnd 0.009888f
C2812 vdd.n1671 gnd 0.009888f
C2813 vdd.n1672 gnd 0.009888f
C2814 vdd.n1673 gnd 0.009888f
C2815 vdd.n1674 gnd 0.009888f
C2816 vdd.n1675 gnd 0.007959f
C2817 vdd.n1677 gnd 0.009888f
C2818 vdd.n1678 gnd 0.009888f
C2819 vdd.n1679 gnd 0.009888f
C2820 vdd.n1680 gnd 0.009888f
C2821 vdd.n1681 gnd 0.007879f
C2822 vdd.t97 gnd 0.12165f
C2823 vdd.t96 gnd 0.130011f
C2824 vdd.t95 gnd 0.158874f
C2825 vdd.n1682 gnd 0.203654f
C2826 vdd.n1683 gnd 0.171106f
C2827 vdd.n1685 gnd 0.009888f
C2828 vdd.n1686 gnd 0.009888f
C2829 vdd.n1687 gnd 0.007959f
C2830 vdd.n1688 gnd 0.009888f
C2831 vdd.n1690 gnd 0.009888f
C2832 vdd.n1691 gnd 0.009888f
C2833 vdd.n1692 gnd 0.009888f
C2834 vdd.n1693 gnd 0.009888f
C2835 vdd.n1694 gnd 0.007959f
C2836 vdd.n1696 gnd 0.009888f
C2837 vdd.n1697 gnd 0.009888f
C2838 vdd.n1698 gnd 0.009888f
C2839 vdd.n1699 gnd 0.009888f
C2840 vdd.n1700 gnd 0.009888f
C2841 vdd.n1701 gnd 0.007959f
C2842 vdd.n1703 gnd 0.009888f
C2843 vdd.n1704 gnd 0.009888f
C2844 vdd.n1705 gnd 0.009888f
C2845 vdd.n1706 gnd 0.009888f
C2846 vdd.n1707 gnd 0.009888f
C2847 vdd.n1708 gnd 0.009888f
C2848 vdd.n1709 gnd 0.007959f
C2849 vdd.n1711 gnd 0.009888f
C2850 vdd.n1713 gnd 0.009888f
C2851 vdd.n1714 gnd 0.007959f
C2852 vdd.n1715 gnd 0.007959f
C2853 vdd.n1716 gnd 0.009888f
C2854 vdd.n1718 gnd 0.009888f
C2855 vdd.n1719 gnd 0.007959f
C2856 vdd.n1720 gnd 0.007959f
C2857 vdd.n1721 gnd 0.009888f
C2858 vdd.n1723 gnd 0.009888f
C2859 vdd.n1724 gnd 0.009888f
C2860 vdd.n1725 gnd 0.007959f
C2861 vdd.n1726 gnd 0.007959f
C2862 vdd.n1727 gnd 0.007959f
C2863 vdd.n1728 gnd 0.009888f
C2864 vdd.n1730 gnd 0.009888f
C2865 vdd.n1731 gnd 0.009888f
C2866 vdd.n1732 gnd 0.007959f
C2867 vdd.n1733 gnd 0.007959f
C2868 vdd.n1734 gnd 0.007959f
C2869 vdd.n1735 gnd 0.009888f
C2870 vdd.n1737 gnd 0.009888f
C2871 vdd.n1738 gnd 0.009888f
C2872 vdd.n1739 gnd 0.007959f
C2873 vdd.n1740 gnd 0.007959f
C2874 vdd.n1741 gnd 0.007959f
C2875 vdd.n1742 gnd 0.009888f
C2876 vdd.n1744 gnd 0.009888f
C2877 vdd.n1745 gnd 0.009888f
C2878 vdd.n1746 gnd 0.007959f
C2879 vdd.n1747 gnd 0.009888f
C2880 vdd.n1748 gnd 0.009888f
C2881 vdd.n1749 gnd 0.009888f
C2882 vdd.n1750 gnd 0.016236f
C2883 vdd.n1751 gnd 0.005412f
C2884 vdd.n1752 gnd 0.007959f
C2885 vdd.n1753 gnd 0.009888f
C2886 vdd.n1755 gnd 0.009888f
C2887 vdd.n1756 gnd 0.009888f
C2888 vdd.n1757 gnd 0.007959f
C2889 vdd.n1758 gnd 0.007959f
C2890 vdd.n1759 gnd 0.007959f
C2891 vdd.n1760 gnd 0.009888f
C2892 vdd.n1762 gnd 0.009888f
C2893 vdd.n1763 gnd 0.009888f
C2894 vdd.n1764 gnd 0.007959f
C2895 vdd.n1765 gnd 0.007959f
C2896 vdd.n1766 gnd 0.007959f
C2897 vdd.n1767 gnd 0.009888f
C2898 vdd.n1769 gnd 0.009888f
C2899 vdd.n1770 gnd 0.009888f
C2900 vdd.n1771 gnd 0.007959f
C2901 vdd.n1772 gnd 0.007959f
C2902 vdd.n1773 gnd 0.007959f
C2903 vdd.n1774 gnd 0.009888f
C2904 vdd.n1776 gnd 0.009888f
C2905 vdd.n1777 gnd 0.009888f
C2906 vdd.n1778 gnd 0.007959f
C2907 vdd.n1779 gnd 0.007959f
C2908 vdd.n1780 gnd 0.007959f
C2909 vdd.n1781 gnd 0.009888f
C2910 vdd.n1783 gnd 0.009888f
C2911 vdd.n1784 gnd 0.009888f
C2912 vdd.n1785 gnd 0.007959f
C2913 vdd.n1786 gnd 0.009888f
C2914 vdd.n1787 gnd 0.009888f
C2915 vdd.n1788 gnd 0.009888f
C2916 vdd.n1789 gnd 0.016236f
C2917 vdd.n1790 gnd 0.006646f
C2918 vdd.n1791 gnd 0.007959f
C2919 vdd.n1792 gnd 0.009888f
C2920 vdd.n1794 gnd 0.009888f
C2921 vdd.n1795 gnd 0.009888f
C2922 vdd.n1796 gnd 0.007959f
C2923 vdd.n1797 gnd 0.007959f
C2924 vdd.n1798 gnd 0.007959f
C2925 vdd.n1799 gnd 0.009888f
C2926 vdd.n1801 gnd 0.009888f
C2927 vdd.n1802 gnd 0.009888f
C2928 vdd.n1803 gnd 0.007959f
C2929 vdd.n1804 gnd 0.007959f
C2930 vdd.n1805 gnd 0.007959f
C2931 vdd.n1806 gnd 0.009888f
C2932 vdd.n1808 gnd 0.009888f
C2933 vdd.n1809 gnd 0.009888f
C2934 vdd.n1811 gnd 0.009888f
C2935 vdd.n1812 gnd 0.007959f
C2936 vdd.n1813 gnd 0.006328f
C2937 vdd.n1814 gnd 0.006724f
C2938 vdd.n1815 gnd 0.006724f
C2939 vdd.n1816 gnd 0.006724f
C2940 vdd.n1817 gnd 0.006724f
C2941 vdd.n1818 gnd 0.006724f
C2942 vdd.n1819 gnd 0.006724f
C2943 vdd.n1820 gnd 0.006724f
C2944 vdd.n1821 gnd 0.006724f
C2945 vdd.n1823 gnd 0.006724f
C2946 vdd.n1824 gnd 0.006724f
C2947 vdd.n1825 gnd 0.006724f
C2948 vdd.n1826 gnd 0.006724f
C2949 vdd.n1827 gnd 0.006724f
C2950 vdd.n1829 gnd 0.006724f
C2951 vdd.n1831 gnd 0.006724f
C2952 vdd.n1832 gnd 0.006724f
C2953 vdd.n1833 gnd 0.006724f
C2954 vdd.n1834 gnd 0.006724f
C2955 vdd.n1835 gnd 0.006724f
C2956 vdd.n1837 gnd 0.006724f
C2957 vdd.n1839 gnd 0.006724f
C2958 vdd.n1840 gnd 0.006724f
C2959 vdd.n1841 gnd 0.006724f
C2960 vdd.n1842 gnd 0.006724f
C2961 vdd.n1843 gnd 0.006724f
C2962 vdd.n1845 gnd 0.006724f
C2963 vdd.n1847 gnd 0.006724f
C2964 vdd.n1848 gnd 0.006724f
C2965 vdd.n1849 gnd 0.006724f
C2966 vdd.n1850 gnd 0.006724f
C2967 vdd.n1851 gnd 0.006724f
C2968 vdd.n1853 gnd 0.006724f
C2969 vdd.n1854 gnd 0.006724f
C2970 vdd.n1855 gnd 0.006724f
C2971 vdd.n1856 gnd 0.006724f
C2972 vdd.n1857 gnd 0.006724f
C2973 vdd.n1858 gnd 0.006724f
C2974 vdd.n1859 gnd 0.006724f
C2975 vdd.n1860 gnd 0.006724f
C2976 vdd.n1861 gnd 0.004895f
C2977 vdd.n1862 gnd 0.006724f
C2978 vdd.t147 gnd 0.271714f
C2979 vdd.t148 gnd 0.278133f
C2980 vdd.t146 gnd 0.177385f
C2981 vdd.n1863 gnd 0.095867f
C2982 vdd.n1864 gnd 0.054379f
C2983 vdd.n1865 gnd 0.00961f
C2984 vdd.n1866 gnd 0.006724f
C2985 vdd.n1867 gnd 0.006724f
C2986 vdd.n1868 gnd 0.409262f
C2987 vdd.n1869 gnd 0.006724f
C2988 vdd.n1870 gnd 0.006724f
C2989 vdd.n1871 gnd 0.006724f
C2990 vdd.n1872 gnd 0.006724f
C2991 vdd.n1873 gnd 0.006724f
C2992 vdd.n1874 gnd 0.006724f
C2993 vdd.n1875 gnd 0.006724f
C2994 vdd.n1876 gnd 0.006724f
C2995 vdd.n1877 gnd 0.006724f
C2996 vdd.n1878 gnd 0.006724f
C2997 vdd.n1879 gnd 0.006724f
C2998 vdd.n1880 gnd 0.006724f
C2999 vdd.n1881 gnd 0.006724f
C3000 vdd.n1882 gnd 0.006724f
C3001 vdd.n1883 gnd 0.006724f
C3002 vdd.n1884 gnd 0.006724f
C3003 vdd.n1885 gnd 0.006724f
C3004 vdd.n1886 gnd 0.006724f
C3005 vdd.n1887 gnd 0.006724f
C3006 vdd.n1888 gnd 0.006724f
C3007 vdd.t121 gnd 0.271714f
C3008 vdd.t122 gnd 0.278133f
C3009 vdd.t119 gnd 0.177385f
C3010 vdd.n1889 gnd 0.095867f
C3011 vdd.n1890 gnd 0.054379f
C3012 vdd.n1891 gnd 0.006724f
C3013 vdd.n1892 gnd 0.006724f
C3014 vdd.n1893 gnd 0.006724f
C3015 vdd.n1894 gnd 0.006724f
C3016 vdd.n1895 gnd 0.006724f
C3017 vdd.n1896 gnd 0.006724f
C3018 vdd.n1898 gnd 0.006724f
C3019 vdd.n1899 gnd 0.006724f
C3020 vdd.n1900 gnd 0.006724f
C3021 vdd.n1901 gnd 0.006724f
C3022 vdd.n1903 gnd 0.006724f
C3023 vdd.n1905 gnd 0.006724f
C3024 vdd.n1906 gnd 0.006724f
C3025 vdd.n1907 gnd 0.006724f
C3026 vdd.n1908 gnd 0.006724f
C3027 vdd.n1909 gnd 0.006724f
C3028 vdd.n1911 gnd 0.006724f
C3029 vdd.n1913 gnd 0.006724f
C3030 vdd.n1914 gnd 0.006724f
C3031 vdd.n1915 gnd 0.006724f
C3032 vdd.n1916 gnd 0.006724f
C3033 vdd.n1917 gnd 0.006724f
C3034 vdd.n1919 gnd 0.006724f
C3035 vdd.n1921 gnd 0.006724f
C3036 vdd.n1922 gnd 0.006724f
C3037 vdd.n1923 gnd 0.004895f
C3038 vdd.n1924 gnd 0.00961f
C3039 vdd.n1925 gnd 0.005191f
C3040 vdd.n1926 gnd 0.006724f
C3041 vdd.n1928 gnd 0.006724f
C3042 vdd.n1929 gnd 0.015955f
C3043 vdd.n1930 gnd 0.015955f
C3044 vdd.n1931 gnd 0.014896f
C3045 vdd.n1932 gnd 0.006724f
C3046 vdd.n1933 gnd 0.006724f
C3047 vdd.n1934 gnd 0.006724f
C3048 vdd.n1935 gnd 0.006724f
C3049 vdd.n1936 gnd 0.006724f
C3050 vdd.n1937 gnd 0.006724f
C3051 vdd.n1938 gnd 0.006724f
C3052 vdd.n1939 gnd 0.006724f
C3053 vdd.n1940 gnd 0.006724f
C3054 vdd.n1941 gnd 0.006724f
C3055 vdd.n1942 gnd 0.006724f
C3056 vdd.n1943 gnd 0.006724f
C3057 vdd.n1944 gnd 0.006724f
C3058 vdd.n1945 gnd 0.006724f
C3059 vdd.n1946 gnd 0.006724f
C3060 vdd.n1947 gnd 0.006724f
C3061 vdd.n1948 gnd 0.006724f
C3062 vdd.n1949 gnd 0.006724f
C3063 vdd.n1950 gnd 0.006724f
C3064 vdd.n1951 gnd 0.006724f
C3065 vdd.n1952 gnd 0.006724f
C3066 vdd.n1953 gnd 0.006724f
C3067 vdd.n1954 gnd 0.006724f
C3068 vdd.n1955 gnd 0.006724f
C3069 vdd.n1956 gnd 0.006724f
C3070 vdd.n1957 gnd 0.006724f
C3071 vdd.n1958 gnd 0.006724f
C3072 vdd.n1959 gnd 0.006724f
C3073 vdd.n1960 gnd 0.006724f
C3074 vdd.n1961 gnd 0.006724f
C3075 vdd.n1962 gnd 0.006724f
C3076 vdd.n1963 gnd 0.006724f
C3077 vdd.n1964 gnd 0.006724f
C3078 vdd.n1965 gnd 0.006724f
C3079 vdd.n1966 gnd 0.006724f
C3080 vdd.n1967 gnd 0.006724f
C3081 vdd.n1968 gnd 0.006724f
C3082 vdd.n1969 gnd 0.217263f
C3083 vdd.n1970 gnd 0.006724f
C3084 vdd.n1971 gnd 0.006724f
C3085 vdd.n1972 gnd 0.006724f
C3086 vdd.n1973 gnd 0.006724f
C3087 vdd.n1974 gnd 0.006724f
C3088 vdd.n1975 gnd 0.006724f
C3089 vdd.n1976 gnd 0.006724f
C3090 vdd.n1977 gnd 0.006724f
C3091 vdd.n1978 gnd 0.006724f
C3092 vdd.n1979 gnd 0.006724f
C3093 vdd.n1980 gnd 0.006724f
C3094 vdd.n1981 gnd 0.006724f
C3095 vdd.n1982 gnd 0.006724f
C3096 vdd.n1983 gnd 0.006724f
C3097 vdd.n1984 gnd 0.006724f
C3098 vdd.n1985 gnd 0.006724f
C3099 vdd.n1986 gnd 0.006724f
C3100 vdd.n1987 gnd 0.006724f
C3101 vdd.n1988 gnd 0.006724f
C3102 vdd.n1989 gnd 0.006724f
C3103 vdd.n1990 gnd 0.014896f
C3104 vdd.n1992 gnd 0.015955f
C3105 vdd.n1993 gnd 0.015955f
C3106 vdd.n1994 gnd 0.006724f
C3107 vdd.n1995 gnd 0.005191f
C3108 vdd.n1996 gnd 0.006724f
C3109 vdd.n1998 gnd 0.006724f
C3110 vdd.n2000 gnd 0.006724f
C3111 vdd.n2001 gnd 0.006724f
C3112 vdd.n2002 gnd 0.006724f
C3113 vdd.n2003 gnd 0.006724f
C3114 vdd.n2004 gnd 0.006724f
C3115 vdd.n2006 gnd 0.006724f
C3116 vdd.n2008 gnd 0.006724f
C3117 vdd.n2009 gnd 0.006724f
C3118 vdd.n2010 gnd 0.006724f
C3119 vdd.n2011 gnd 0.006724f
C3120 vdd.n2012 gnd 0.006724f
C3121 vdd.n2014 gnd 0.006724f
C3122 vdd.n2016 gnd 0.006724f
C3123 vdd.n2017 gnd 0.006724f
C3124 vdd.n2018 gnd 0.006724f
C3125 vdd.n2019 gnd 0.006724f
C3126 vdd.n2020 gnd 0.006724f
C3127 vdd.n2022 gnd 0.006724f
C3128 vdd.n2024 gnd 0.006724f
C3129 vdd.n2025 gnd 0.006724f
C3130 vdd.n2026 gnd 0.020056f
C3131 vdd.n2027 gnd 0.59455f
C3132 vdd.n2029 gnd 0.007959f
C3133 vdd.n2030 gnd 0.007959f
C3134 vdd.n2031 gnd 0.009888f
C3135 vdd.n2033 gnd 0.009888f
C3136 vdd.n2034 gnd 0.009888f
C3137 vdd.n2035 gnd 0.007959f
C3138 vdd.n2036 gnd 0.006606f
C3139 vdd.n2037 gnd 0.023667f
C3140 vdd.n2038 gnd 0.023302f
C3141 vdd.n2039 gnd 0.006606f
C3142 vdd.n2040 gnd 0.023302f
C3143 vdd.n2041 gnd 1.38947f
C3144 vdd.n2042 gnd 0.023302f
C3145 vdd.n2043 gnd 0.023667f
C3146 vdd.n2044 gnd 0.00378f
C3147 vdd.t86 gnd 0.12165f
C3148 vdd.t85 gnd 0.130011f
C3149 vdd.t83 gnd 0.158874f
C3150 vdd.n2045 gnd 0.203654f
C3151 vdd.n2046 gnd 0.171106f
C3152 vdd.n2047 gnd 0.012257f
C3153 vdd.n2048 gnd 0.004178f
C3154 vdd.n2049 gnd 0.008504f
C3155 vdd.n2050 gnd 0.59455f
C3156 vdd.n2051 gnd 0.020056f
C3157 vdd.n2052 gnd 0.006724f
C3158 vdd.n2053 gnd 0.006724f
C3159 vdd.n2054 gnd 0.006724f
C3160 vdd.n2056 gnd 0.006724f
C3161 vdd.n2058 gnd 0.006724f
C3162 vdd.n2059 gnd 0.006724f
C3163 vdd.n2060 gnd 0.006724f
C3164 vdd.n2061 gnd 0.006724f
C3165 vdd.n2062 gnd 0.006724f
C3166 vdd.n2064 gnd 0.006724f
C3167 vdd.n2066 gnd 0.006724f
C3168 vdd.n2067 gnd 0.006724f
C3169 vdd.n2068 gnd 0.006724f
C3170 vdd.n2069 gnd 0.006724f
C3171 vdd.n2070 gnd 0.006724f
C3172 vdd.n2072 gnd 0.006724f
C3173 vdd.n2074 gnd 0.006724f
C3174 vdd.n2075 gnd 0.006724f
C3175 vdd.n2076 gnd 0.006724f
C3176 vdd.n2077 gnd 0.006724f
C3177 vdd.n2078 gnd 0.006724f
C3178 vdd.n2080 gnd 0.006724f
C3179 vdd.n2082 gnd 0.006724f
C3180 vdd.n2083 gnd 0.006724f
C3181 vdd.n2084 gnd 0.015955f
C3182 vdd.n2085 gnd 0.014896f
C3183 vdd.n2086 gnd 0.014896f
C3184 vdd.n2087 gnd 0.990313f
C3185 vdd.n2088 gnd 0.014896f
C3186 vdd.n2089 gnd 0.014896f
C3187 vdd.n2090 gnd 0.006724f
C3188 vdd.n2091 gnd 0.006724f
C3189 vdd.n2092 gnd 0.006724f
C3190 vdd.n2093 gnd 0.429473f
C3191 vdd.n2094 gnd 0.006724f
C3192 vdd.n2095 gnd 0.006724f
C3193 vdd.n2096 gnd 0.006724f
C3194 vdd.n2097 gnd 0.006724f
C3195 vdd.n2098 gnd 0.006724f
C3196 vdd.n2099 gnd 0.687156f
C3197 vdd.n2100 gnd 0.006724f
C3198 vdd.n2101 gnd 0.006724f
C3199 vdd.n2102 gnd 0.006724f
C3200 vdd.n2103 gnd 0.006724f
C3201 vdd.n2104 gnd 0.006724f
C3202 vdd.n2105 gnd 0.687156f
C3203 vdd.n2106 gnd 0.006724f
C3204 vdd.n2107 gnd 0.006724f
C3205 vdd.n2108 gnd 0.005933f
C3206 vdd.n2109 gnd 0.019478f
C3207 vdd.n2110 gnd 0.004153f
C3208 vdd.n2111 gnd 0.006724f
C3209 vdd.n2112 gnd 0.378946f
C3210 vdd.n2113 gnd 0.006724f
C3211 vdd.n2114 gnd 0.006724f
C3212 vdd.n2115 gnd 0.006724f
C3213 vdd.n2116 gnd 0.006724f
C3214 vdd.n2117 gnd 0.006724f
C3215 vdd.n2118 gnd 0.459788f
C3216 vdd.n2119 gnd 0.006724f
C3217 vdd.n2120 gnd 0.006724f
C3218 vdd.n2121 gnd 0.006724f
C3219 vdd.n2122 gnd 0.006724f
C3220 vdd.n2123 gnd 0.006724f
C3221 vdd.n2124 gnd 0.611367f
C3222 vdd.n2125 gnd 0.006724f
C3223 vdd.n2126 gnd 0.006724f
C3224 vdd.n2127 gnd 0.006724f
C3225 vdd.n2128 gnd 0.006724f
C3226 vdd.n2129 gnd 0.006724f
C3227 vdd.n2130 gnd 0.545683f
C3228 vdd.n2131 gnd 0.006724f
C3229 vdd.n2132 gnd 0.006724f
C3230 vdd.n2133 gnd 0.006724f
C3231 vdd.n2134 gnd 0.006724f
C3232 vdd.n2135 gnd 0.006724f
C3233 vdd.n2136 gnd 0.394104f
C3234 vdd.n2137 gnd 0.006724f
C3235 vdd.n2138 gnd 0.006724f
C3236 vdd.n2139 gnd 0.006724f
C3237 vdd.n2140 gnd 0.006724f
C3238 vdd.n2141 gnd 0.006724f
C3239 vdd.n2142 gnd 0.217263f
C3240 vdd.n2143 gnd 0.006724f
C3241 vdd.n2144 gnd 0.006724f
C3242 vdd.n2145 gnd 0.006724f
C3243 vdd.n2146 gnd 0.006724f
C3244 vdd.n2147 gnd 0.006724f
C3245 vdd.n2148 gnd 0.378946f
C3246 vdd.n2149 gnd 0.006724f
C3247 vdd.n2150 gnd 0.006724f
C3248 vdd.n2151 gnd 0.006724f
C3249 vdd.n2152 gnd 0.006724f
C3250 vdd.n2153 gnd 0.006724f
C3251 vdd.n2154 gnd 0.687156f
C3252 vdd.n2155 gnd 0.006724f
C3253 vdd.n2156 gnd 0.006724f
C3254 vdd.n2157 gnd 0.006724f
C3255 vdd.n2158 gnd 0.006724f
C3256 vdd.n2159 gnd 0.006724f
C3257 vdd.n2160 gnd 0.006724f
C3258 vdd.n2161 gnd 0.006724f
C3259 vdd.n2162 gnd 0.535578f
C3260 vdd.n2163 gnd 0.006724f
C3261 vdd.n2164 gnd 0.006724f
C3262 vdd.n2165 gnd 0.006724f
C3263 vdd.n2166 gnd 0.006724f
C3264 vdd.n2167 gnd 0.006724f
C3265 vdd.n2168 gnd 0.006724f
C3266 vdd.n2169 gnd 0.429473f
C3267 vdd.n2170 gnd 0.006724f
C3268 vdd.n2171 gnd 0.006724f
C3269 vdd.n2172 gnd 0.006724f
C3270 vdd.n2173 gnd 0.015715f
C3271 vdd.n2174 gnd 0.015136f
C3272 vdd.n2175 gnd 0.006724f
C3273 vdd.n2176 gnd 0.006724f
C3274 vdd.n2177 gnd 0.005191f
C3275 vdd.n2178 gnd 0.006724f
C3276 vdd.n2179 gnd 0.006724f
C3277 vdd.n2180 gnd 0.004895f
C3278 vdd.n2181 gnd 0.006724f
C3279 vdd.n2182 gnd 0.006724f
C3280 vdd.n2183 gnd 0.006724f
C3281 vdd.n2184 gnd 0.006724f
C3282 vdd.n2185 gnd 0.006724f
C3283 vdd.n2186 gnd 0.006724f
C3284 vdd.n2187 gnd 0.006724f
C3285 vdd.n2188 gnd 0.006724f
C3286 vdd.n2189 gnd 0.006724f
C3287 vdd.n2190 gnd 0.006724f
C3288 vdd.n2191 gnd 0.006724f
C3289 vdd.n2192 gnd 0.006724f
C3290 vdd.n2193 gnd 0.006724f
C3291 vdd.n2194 gnd 0.006724f
C3292 vdd.n2195 gnd 0.006724f
C3293 vdd.n2196 gnd 0.006724f
C3294 vdd.n2197 gnd 0.006724f
C3295 vdd.n2198 gnd 0.006724f
C3296 vdd.n2199 gnd 0.006724f
C3297 vdd.n2200 gnd 0.006724f
C3298 vdd.n2201 gnd 0.006724f
C3299 vdd.n2202 gnd 0.006724f
C3300 vdd.n2203 gnd 0.006724f
C3301 vdd.n2204 gnd 0.006724f
C3302 vdd.n2205 gnd 0.006724f
C3303 vdd.n2206 gnd 0.006724f
C3304 vdd.n2207 gnd 0.006724f
C3305 vdd.n2208 gnd 0.006724f
C3306 vdd.n2209 gnd 0.006724f
C3307 vdd.n2210 gnd 0.006724f
C3308 vdd.n2211 gnd 0.006724f
C3309 vdd.n2212 gnd 0.006724f
C3310 vdd.n2213 gnd 0.006724f
C3311 vdd.n2214 gnd 0.006724f
C3312 vdd.n2215 gnd 0.006724f
C3313 vdd.n2216 gnd 0.006724f
C3314 vdd.n2217 gnd 0.006724f
C3315 vdd.n2218 gnd 0.006724f
C3316 vdd.n2219 gnd 0.006724f
C3317 vdd.n2220 gnd 0.006724f
C3318 vdd.n2221 gnd 0.006724f
C3319 vdd.n2222 gnd 0.006724f
C3320 vdd.n2223 gnd 0.006724f
C3321 vdd.n2224 gnd 0.006724f
C3322 vdd.n2225 gnd 0.006724f
C3323 vdd.n2226 gnd 0.006724f
C3324 vdd.n2227 gnd 0.006724f
C3325 vdd.n2228 gnd 0.006724f
C3326 vdd.n2229 gnd 0.006724f
C3327 vdd.n2230 gnd 0.006724f
C3328 vdd.n2231 gnd 0.006724f
C3329 vdd.n2232 gnd 0.006724f
C3330 vdd.n2233 gnd 0.006724f
C3331 vdd.n2234 gnd 0.006724f
C3332 vdd.n2235 gnd 0.006724f
C3333 vdd.n2236 gnd 0.006724f
C3334 vdd.n2237 gnd 0.006724f
C3335 vdd.n2238 gnd 0.006724f
C3336 vdd.n2239 gnd 0.006724f
C3337 vdd.n2240 gnd 0.006724f
C3338 vdd.n2241 gnd 0.015955f
C3339 vdd.n2242 gnd 0.014896f
C3340 vdd.n2243 gnd 0.014896f
C3341 vdd.n2244 gnd 0.838735f
C3342 vdd.n2245 gnd 0.014896f
C3343 vdd.n2246 gnd 0.015955f
C3344 vdd.n2247 gnd 0.015136f
C3345 vdd.n2248 gnd 0.006724f
C3346 vdd.n2249 gnd 0.006724f
C3347 vdd.n2250 gnd 0.006724f
C3348 vdd.n2251 gnd 0.005191f
C3349 vdd.n2252 gnd 0.00961f
C3350 vdd.n2253 gnd 0.004895f
C3351 vdd.n2254 gnd 0.006724f
C3352 vdd.n2255 gnd 0.006724f
C3353 vdd.n2256 gnd 0.006724f
C3354 vdd.n2257 gnd 0.006724f
C3355 vdd.n2258 gnd 0.006724f
C3356 vdd.n2259 gnd 0.006724f
C3357 vdd.n2260 gnd 0.006724f
C3358 vdd.n2261 gnd 0.006724f
C3359 vdd.n2262 gnd 0.006724f
C3360 vdd.n2263 gnd 0.006724f
C3361 vdd.n2264 gnd 0.006724f
C3362 vdd.n2265 gnd 0.006724f
C3363 vdd.n2266 gnd 0.006724f
C3364 vdd.n2267 gnd 0.006724f
C3365 vdd.n2268 gnd 0.006724f
C3366 vdd.n2269 gnd 0.006724f
C3367 vdd.n2270 gnd 0.006724f
C3368 vdd.n2271 gnd 0.006724f
C3369 vdd.n2272 gnd 0.006724f
C3370 vdd.n2273 gnd 0.006724f
C3371 vdd.n2274 gnd 0.006724f
C3372 vdd.n2275 gnd 0.006724f
C3373 vdd.n2276 gnd 0.006724f
C3374 vdd.n2277 gnd 0.006724f
C3375 vdd.n2278 gnd 0.006724f
C3376 vdd.n2279 gnd 0.006724f
C3377 vdd.n2280 gnd 0.006724f
C3378 vdd.n2281 gnd 0.006724f
C3379 vdd.n2282 gnd 0.006724f
C3380 vdd.n2283 gnd 0.006724f
C3381 vdd.n2284 gnd 0.006724f
C3382 vdd.n2285 gnd 0.006724f
C3383 vdd.n2286 gnd 0.006724f
C3384 vdd.n2287 gnd 0.006724f
C3385 vdd.n2288 gnd 0.006724f
C3386 vdd.n2289 gnd 0.006724f
C3387 vdd.n2290 gnd 0.006724f
C3388 vdd.n2291 gnd 0.006724f
C3389 vdd.n2292 gnd 0.006724f
C3390 vdd.n2293 gnd 0.006724f
C3391 vdd.n2294 gnd 0.006724f
C3392 vdd.n2295 gnd 0.006724f
C3393 vdd.n2296 gnd 0.006724f
C3394 vdd.n2297 gnd 0.006724f
C3395 vdd.n2298 gnd 0.006724f
C3396 vdd.n2299 gnd 0.006724f
C3397 vdd.n2300 gnd 0.006724f
C3398 vdd.n2301 gnd 0.006724f
C3399 vdd.n2302 gnd 0.006724f
C3400 vdd.n2303 gnd 0.006724f
C3401 vdd.n2304 gnd 0.006724f
C3402 vdd.n2305 gnd 0.006724f
C3403 vdd.n2306 gnd 0.006724f
C3404 vdd.n2307 gnd 0.006724f
C3405 vdd.n2308 gnd 0.006724f
C3406 vdd.n2309 gnd 0.006724f
C3407 vdd.n2310 gnd 0.006724f
C3408 vdd.n2311 gnd 0.006724f
C3409 vdd.n2312 gnd 0.006724f
C3410 vdd.n2313 gnd 0.006724f
C3411 vdd.n2314 gnd 0.015955f
C3412 vdd.n2315 gnd 0.015955f
C3413 vdd.n2316 gnd 0.838735f
C3414 vdd.t204 gnd 2.98104f
C3415 vdd.t156 gnd 2.98104f
C3416 vdd.n2349 gnd 0.015955f
C3417 vdd.n2350 gnd 0.006724f
C3418 vdd.t114 gnd 0.271714f
C3419 vdd.t115 gnd 0.278133f
C3420 vdd.t112 gnd 0.177385f
C3421 vdd.n2351 gnd 0.095867f
C3422 vdd.n2352 gnd 0.054379f
C3423 vdd.n2353 gnd 0.006724f
C3424 vdd.t128 gnd 0.271714f
C3425 vdd.t129 gnd 0.278133f
C3426 vdd.t127 gnd 0.177385f
C3427 vdd.n2354 gnd 0.095867f
C3428 vdd.n2355 gnd 0.054379f
C3429 vdd.n2356 gnd 0.00961f
C3430 vdd.n2357 gnd 0.006724f
C3431 vdd.n2358 gnd 0.006724f
C3432 vdd.n2359 gnd 0.006724f
C3433 vdd.n2360 gnd 0.006724f
C3434 vdd.n2361 gnd 0.006724f
C3435 vdd.n2362 gnd 0.006724f
C3436 vdd.n2363 gnd 0.006724f
C3437 vdd.n2364 gnd 0.006724f
C3438 vdd.n2365 gnd 0.006724f
C3439 vdd.n2366 gnd 0.006724f
C3440 vdd.n2367 gnd 0.006724f
C3441 vdd.n2368 gnd 0.006724f
C3442 vdd.n2369 gnd 0.006724f
C3443 vdd.n2370 gnd 0.006724f
C3444 vdd.n2371 gnd 0.006724f
C3445 vdd.n2372 gnd 0.006724f
C3446 vdd.n2373 gnd 0.006724f
C3447 vdd.n2374 gnd 0.006724f
C3448 vdd.n2375 gnd 0.006724f
C3449 vdd.n2376 gnd 0.006724f
C3450 vdd.n2377 gnd 0.006724f
C3451 vdd.n2378 gnd 0.006724f
C3452 vdd.n2379 gnd 0.006724f
C3453 vdd.n2380 gnd 0.006724f
C3454 vdd.n2381 gnd 0.006724f
C3455 vdd.n2382 gnd 0.006724f
C3456 vdd.n2383 gnd 0.006724f
C3457 vdd.n2384 gnd 0.006724f
C3458 vdd.n2385 gnd 0.006724f
C3459 vdd.n2386 gnd 0.006724f
C3460 vdd.n2387 gnd 0.006724f
C3461 vdd.n2388 gnd 0.006724f
C3462 vdd.n2389 gnd 0.006724f
C3463 vdd.n2390 gnd 0.006724f
C3464 vdd.n2391 gnd 0.006724f
C3465 vdd.n2392 gnd 0.006724f
C3466 vdd.n2393 gnd 0.006724f
C3467 vdd.n2394 gnd 0.006724f
C3468 vdd.n2395 gnd 0.006724f
C3469 vdd.n2396 gnd 0.006724f
C3470 vdd.n2397 gnd 0.006724f
C3471 vdd.n2398 gnd 0.006724f
C3472 vdd.n2399 gnd 0.006724f
C3473 vdd.n2400 gnd 0.006724f
C3474 vdd.n2401 gnd 0.006724f
C3475 vdd.n2402 gnd 0.006724f
C3476 vdd.n2403 gnd 0.006724f
C3477 vdd.n2404 gnd 0.006724f
C3478 vdd.n2405 gnd 0.006724f
C3479 vdd.n2406 gnd 0.006724f
C3480 vdd.n2407 gnd 0.006724f
C3481 vdd.n2408 gnd 0.006724f
C3482 vdd.n2409 gnd 0.006724f
C3483 vdd.n2410 gnd 0.006724f
C3484 vdd.n2411 gnd 0.006724f
C3485 vdd.n2412 gnd 0.006724f
C3486 vdd.n2413 gnd 0.004895f
C3487 vdd.n2414 gnd 0.006724f
C3488 vdd.n2415 gnd 0.006724f
C3489 vdd.n2416 gnd 0.005191f
C3490 vdd.n2417 gnd 0.006724f
C3491 vdd.n2418 gnd 0.006724f
C3492 vdd.n2419 gnd 0.015955f
C3493 vdd.n2420 gnd 0.014896f
C3494 vdd.n2421 gnd 0.006724f
C3495 vdd.n2422 gnd 0.006724f
C3496 vdd.n2423 gnd 0.006724f
C3497 vdd.n2424 gnd 0.006724f
C3498 vdd.n2425 gnd 0.006724f
C3499 vdd.n2426 gnd 0.006724f
C3500 vdd.n2427 gnd 0.006724f
C3501 vdd.n2428 gnd 0.006724f
C3502 vdd.n2429 gnd 0.006724f
C3503 vdd.n2430 gnd 0.006724f
C3504 vdd.n2431 gnd 0.006724f
C3505 vdd.n2432 gnd 0.006724f
C3506 vdd.n2433 gnd 0.006724f
C3507 vdd.n2434 gnd 0.006724f
C3508 vdd.n2435 gnd 0.006724f
C3509 vdd.n2436 gnd 0.006724f
C3510 vdd.n2437 gnd 0.006724f
C3511 vdd.n2438 gnd 0.006724f
C3512 vdd.n2439 gnd 0.006724f
C3513 vdd.n2440 gnd 0.006724f
C3514 vdd.n2441 gnd 0.006724f
C3515 vdd.n2442 gnd 0.006724f
C3516 vdd.n2443 gnd 0.006724f
C3517 vdd.n2444 gnd 0.006724f
C3518 vdd.n2445 gnd 0.006724f
C3519 vdd.n2446 gnd 0.006724f
C3520 vdd.n2447 gnd 0.006724f
C3521 vdd.n2448 gnd 0.006724f
C3522 vdd.n2449 gnd 0.006724f
C3523 vdd.n2450 gnd 0.006724f
C3524 vdd.n2451 gnd 0.006724f
C3525 vdd.n2452 gnd 0.006724f
C3526 vdd.n2453 gnd 0.006724f
C3527 vdd.n2454 gnd 0.006724f
C3528 vdd.n2455 gnd 0.006724f
C3529 vdd.n2456 gnd 0.006724f
C3530 vdd.n2457 gnd 0.006724f
C3531 vdd.n2458 gnd 0.006724f
C3532 vdd.n2459 gnd 0.006724f
C3533 vdd.n2460 gnd 0.006724f
C3534 vdd.n2461 gnd 0.006724f
C3535 vdd.n2462 gnd 0.006724f
C3536 vdd.n2463 gnd 0.006724f
C3537 vdd.n2464 gnd 0.006724f
C3538 vdd.n2465 gnd 0.006724f
C3539 vdd.n2466 gnd 0.006724f
C3540 vdd.n2467 gnd 0.006724f
C3541 vdd.n2468 gnd 0.006724f
C3542 vdd.n2469 gnd 0.006724f
C3543 vdd.n2470 gnd 0.006724f
C3544 vdd.n2471 gnd 0.006724f
C3545 vdd.n2472 gnd 0.217263f
C3546 vdd.n2473 gnd 0.006724f
C3547 vdd.n2474 gnd 0.006724f
C3548 vdd.n2475 gnd 0.006724f
C3549 vdd.n2476 gnd 0.006724f
C3550 vdd.n2477 gnd 0.006724f
C3551 vdd.n2478 gnd 0.006724f
C3552 vdd.n2479 gnd 0.006724f
C3553 vdd.n2480 gnd 0.006724f
C3554 vdd.n2481 gnd 0.006724f
C3555 vdd.n2482 gnd 0.006724f
C3556 vdd.n2483 gnd 0.006724f
C3557 vdd.n2484 gnd 0.006724f
C3558 vdd.n2485 gnd 0.006724f
C3559 vdd.n2486 gnd 0.006724f
C3560 vdd.n2487 gnd 0.006724f
C3561 vdd.n2488 gnd 0.006724f
C3562 vdd.n2489 gnd 0.006724f
C3563 vdd.n2490 gnd 0.006724f
C3564 vdd.n2491 gnd 0.006724f
C3565 vdd.n2492 gnd 0.006724f
C3566 vdd.n2493 gnd 0.409262f
C3567 vdd.n2494 gnd 0.006724f
C3568 vdd.n2495 gnd 0.006724f
C3569 vdd.n2496 gnd 0.006724f
C3570 vdd.n2497 gnd 0.006724f
C3571 vdd.n2498 gnd 0.006724f
C3572 vdd.n2499 gnd 0.014896f
C3573 vdd.n2500 gnd 0.015955f
C3574 vdd.n2501 gnd 0.015955f
C3575 vdd.n2502 gnd 0.006724f
C3576 vdd.n2503 gnd 0.006724f
C3577 vdd.n2504 gnd 0.006724f
C3578 vdd.n2505 gnd 0.005191f
C3579 vdd.n2506 gnd 0.00961f
C3580 vdd.n2507 gnd 0.004895f
C3581 vdd.n2508 gnd 0.006724f
C3582 vdd.n2509 gnd 0.006724f
C3583 vdd.n2510 gnd 0.006724f
C3584 vdd.n2511 gnd 0.006724f
C3585 vdd.n2512 gnd 0.006724f
C3586 vdd.n2513 gnd 0.006724f
C3587 vdd.n2514 gnd 0.006724f
C3588 vdd.n2515 gnd 0.006724f
C3589 vdd.n2516 gnd 0.006724f
C3590 vdd.n2517 gnd 0.006724f
C3591 vdd.n2518 gnd 0.006724f
C3592 vdd.n2519 gnd 0.006724f
C3593 vdd.n2520 gnd 0.006724f
C3594 vdd.n2521 gnd 0.006724f
C3595 vdd.n2522 gnd 0.006724f
C3596 vdd.n2523 gnd 0.006724f
C3597 vdd.n2524 gnd 0.006724f
C3598 vdd.n2525 gnd 0.006724f
C3599 vdd.n2526 gnd 0.006724f
C3600 vdd.n2527 gnd 0.006724f
C3601 vdd.n2528 gnd 0.006724f
C3602 vdd.n2529 gnd 0.006724f
C3603 vdd.n2530 gnd 0.006724f
C3604 vdd.n2531 gnd 0.006724f
C3605 vdd.n2532 gnd 0.006724f
C3606 vdd.n2533 gnd 0.006724f
C3607 vdd.n2534 gnd 0.006724f
C3608 vdd.n2535 gnd 0.006724f
C3609 vdd.n2536 gnd 0.006724f
C3610 vdd.n2537 gnd 0.006724f
C3611 vdd.n2538 gnd 0.006724f
C3612 vdd.n2539 gnd 0.006724f
C3613 vdd.n2540 gnd 0.006724f
C3614 vdd.n2541 gnd 0.006724f
C3615 vdd.n2542 gnd 0.006724f
C3616 vdd.n2543 gnd 0.006724f
C3617 vdd.n2544 gnd 0.006724f
C3618 vdd.n2545 gnd 0.006724f
C3619 vdd.n2546 gnd 0.006724f
C3620 vdd.n2547 gnd 0.006724f
C3621 vdd.n2548 gnd 0.006724f
C3622 vdd.n2549 gnd 0.006724f
C3623 vdd.n2550 gnd 0.006724f
C3624 vdd.n2551 gnd 0.006724f
C3625 vdd.n2552 gnd 0.006724f
C3626 vdd.n2553 gnd 0.006724f
C3627 vdd.n2554 gnd 0.006724f
C3628 vdd.n2555 gnd 0.006724f
C3629 vdd.n2556 gnd 0.006724f
C3630 vdd.n2557 gnd 0.006724f
C3631 vdd.n2558 gnd 0.006724f
C3632 vdd.n2559 gnd 0.006724f
C3633 vdd.n2560 gnd 0.006724f
C3634 vdd.n2561 gnd 0.006724f
C3635 vdd.n2562 gnd 0.006724f
C3636 vdd.n2563 gnd 0.006724f
C3637 vdd.n2564 gnd 0.006724f
C3638 vdd.n2565 gnd 0.006724f
C3639 vdd.n2566 gnd 0.006724f
C3640 vdd.n2567 gnd 0.006724f
C3641 vdd.n2569 gnd 0.838735f
C3642 vdd.n2571 gnd 0.006724f
C3643 vdd.n2572 gnd 0.006724f
C3644 vdd.n2573 gnd 0.015955f
C3645 vdd.n2574 gnd 0.014896f
C3646 vdd.n2575 gnd 0.014896f
C3647 vdd.n2576 gnd 0.838735f
C3648 vdd.n2577 gnd 0.014896f
C3649 vdd.n2578 gnd 0.014896f
C3650 vdd.n2579 gnd 0.006724f
C3651 vdd.n2580 gnd 0.006724f
C3652 vdd.n2581 gnd 0.006724f
C3653 vdd.n2582 gnd 0.429473f
C3654 vdd.n2583 gnd 0.006724f
C3655 vdd.n2584 gnd 0.006724f
C3656 vdd.n2585 gnd 0.006724f
C3657 vdd.n2586 gnd 0.006724f
C3658 vdd.n2587 gnd 0.006724f
C3659 vdd.n2588 gnd 0.535578f
C3660 vdd.n2589 gnd 0.006724f
C3661 vdd.n2590 gnd 0.006724f
C3662 vdd.n2591 gnd 0.006724f
C3663 vdd.n2592 gnd 0.006724f
C3664 vdd.n2593 gnd 0.006724f
C3665 vdd.n2594 gnd 0.687156f
C3666 vdd.n2595 gnd 0.006724f
C3667 vdd.n2596 gnd 0.006724f
C3668 vdd.n2597 gnd 0.006724f
C3669 vdd.n2598 gnd 0.006724f
C3670 vdd.n2599 gnd 0.006724f
C3671 vdd.n2600 gnd 0.378946f
C3672 vdd.n2601 gnd 0.006724f
C3673 vdd.n2602 gnd 0.006724f
C3674 vdd.n2603 gnd 0.006724f
C3675 vdd.n2604 gnd 0.006724f
C3676 vdd.n2605 gnd 0.006724f
C3677 vdd.n2606 gnd 0.217263f
C3678 vdd.n2607 gnd 0.006724f
C3679 vdd.n2608 gnd 0.006724f
C3680 vdd.n2609 gnd 0.006724f
C3681 vdd.n2610 gnd 0.006724f
C3682 vdd.n2611 gnd 0.006724f
C3683 vdd.n2612 gnd 0.394104f
C3684 vdd.n2613 gnd 0.006724f
C3685 vdd.n2614 gnd 0.006724f
C3686 vdd.n2615 gnd 0.006724f
C3687 vdd.n2616 gnd 0.006724f
C3688 vdd.n2617 gnd 0.006724f
C3689 vdd.n2618 gnd 0.545683f
C3690 vdd.n2619 gnd 0.006724f
C3691 vdd.n2620 gnd 0.006724f
C3692 vdd.n2621 gnd 0.006724f
C3693 vdd.n2622 gnd 0.006724f
C3694 vdd.n2623 gnd 0.006724f
C3695 vdd.n2624 gnd 0.611367f
C3696 vdd.n2625 gnd 0.006724f
C3697 vdd.n2626 gnd 0.006724f
C3698 vdd.n2627 gnd 0.006724f
C3699 vdd.n2628 gnd 0.006724f
C3700 vdd.n2629 gnd 0.006724f
C3701 vdd.n2630 gnd 0.459788f
C3702 vdd.n2631 gnd 0.006724f
C3703 vdd.n2632 gnd 0.006724f
C3704 vdd.n2633 gnd 0.006724f
C3705 vdd.t93 gnd 0.278133f
C3706 vdd.t91 gnd 0.177385f
C3707 vdd.t94 gnd 0.278133f
C3708 vdd.n2634 gnd 0.156322f
C3709 vdd.n2635 gnd 0.019478f
C3710 vdd.n2636 gnd 0.004153f
C3711 vdd.n2637 gnd 0.006724f
C3712 vdd.n2638 gnd 0.378946f
C3713 vdd.n2639 gnd 0.006724f
C3714 vdd.n2640 gnd 0.006724f
C3715 vdd.n2641 gnd 0.006724f
C3716 vdd.n2642 gnd 0.006724f
C3717 vdd.n2643 gnd 0.006724f
C3718 vdd.n2644 gnd 0.687156f
C3719 vdd.n2645 gnd 0.006724f
C3720 vdd.n2646 gnd 0.006724f
C3721 vdd.n2647 gnd 0.006724f
C3722 vdd.n2648 gnd 0.006724f
C3723 vdd.n2649 gnd 0.006724f
C3724 vdd.n2650 gnd 0.006724f
C3725 vdd.n2652 gnd 0.006724f
C3726 vdd.n2653 gnd 0.006724f
C3727 vdd.n2655 gnd 0.006724f
C3728 vdd.n2656 gnd 0.006724f
C3729 vdd.n2659 gnd 0.006724f
C3730 vdd.n2660 gnd 0.006724f
C3731 vdd.n2661 gnd 0.006724f
C3732 vdd.n2662 gnd 0.006724f
C3733 vdd.n2664 gnd 0.006724f
C3734 vdd.n2665 gnd 0.006724f
C3735 vdd.n2666 gnd 0.006724f
C3736 vdd.n2667 gnd 0.006724f
C3737 vdd.n2668 gnd 0.006724f
C3738 vdd.n2669 gnd 0.006724f
C3739 vdd.n2671 gnd 0.006724f
C3740 vdd.n2672 gnd 0.006724f
C3741 vdd.n2673 gnd 0.006724f
C3742 vdd.n2674 gnd 0.006724f
C3743 vdd.n2675 gnd 0.006724f
C3744 vdd.n2676 gnd 0.006724f
C3745 vdd.n2678 gnd 0.006724f
C3746 vdd.n2679 gnd 0.006724f
C3747 vdd.n2680 gnd 0.006724f
C3748 vdd.n2681 gnd 0.006724f
C3749 vdd.n2682 gnd 0.006724f
C3750 vdd.n2683 gnd 0.006724f
C3751 vdd.n2685 gnd 0.006724f
C3752 vdd.n2686 gnd 0.015955f
C3753 vdd.n2687 gnd 0.015955f
C3754 vdd.n2688 gnd 0.014896f
C3755 vdd.n2689 gnd 0.006724f
C3756 vdd.n2690 gnd 0.006724f
C3757 vdd.n2691 gnd 0.006724f
C3758 vdd.n2692 gnd 0.006724f
C3759 vdd.n2693 gnd 0.006724f
C3760 vdd.n2694 gnd 0.006724f
C3761 vdd.n2695 gnd 0.687156f
C3762 vdd.n2696 gnd 0.006724f
C3763 vdd.n2697 gnd 0.006724f
C3764 vdd.n2698 gnd 0.006724f
C3765 vdd.n2699 gnd 0.006724f
C3766 vdd.n2700 gnd 0.006724f
C3767 vdd.n2701 gnd 0.429473f
C3768 vdd.n2702 gnd 0.006724f
C3769 vdd.n2703 gnd 0.006724f
C3770 vdd.n2704 gnd 0.006724f
C3771 vdd.n2705 gnd 0.015715f
C3772 vdd.n2707 gnd 0.015955f
C3773 vdd.n2708 gnd 0.015136f
C3774 vdd.n2709 gnd 0.006724f
C3775 vdd.n2710 gnd 0.005191f
C3776 vdd.n2711 gnd 0.006724f
C3777 vdd.n2713 gnd 0.006724f
C3778 vdd.n2714 gnd 0.006724f
C3779 vdd.n2715 gnd 0.006724f
C3780 vdd.n2716 gnd 0.006724f
C3781 vdd.n2717 gnd 0.006724f
C3782 vdd.n2718 gnd 0.006724f
C3783 vdd.n2720 gnd 0.006724f
C3784 vdd.n2721 gnd 0.006724f
C3785 vdd.n2722 gnd 0.006724f
C3786 vdd.n2723 gnd 0.006724f
C3787 vdd.n2724 gnd 0.006724f
C3788 vdd.n2725 gnd 0.006724f
C3789 vdd.n2727 gnd 0.006724f
C3790 vdd.n2728 gnd 0.006724f
C3791 vdd.n2729 gnd 0.006724f
C3792 vdd.n2730 gnd 0.006724f
C3793 vdd.n2731 gnd 0.006724f
C3794 vdd.n2732 gnd 0.006724f
C3795 vdd.n2734 gnd 0.006724f
C3796 vdd.n2735 gnd 0.006724f
C3797 vdd.n2736 gnd 0.006724f
C3798 vdd.n2737 gnd 0.598448f
C3799 vdd.n2738 gnd 0.016158f
C3800 vdd.n2739 gnd 0.006724f
C3801 vdd.n2740 gnd 0.006724f
C3802 vdd.n2742 gnd 0.006724f
C3803 vdd.n2743 gnd 0.006724f
C3804 vdd.n2744 gnd 0.006724f
C3805 vdd.n2745 gnd 0.006724f
C3806 vdd.n2746 gnd 0.006724f
C3807 vdd.n2747 gnd 0.006724f
C3808 vdd.n2749 gnd 0.006724f
C3809 vdd.n2750 gnd 0.006724f
C3810 vdd.n2751 gnd 0.006724f
C3811 vdd.n2752 gnd 0.006724f
C3812 vdd.n2753 gnd 0.006724f
C3813 vdd.n2754 gnd 0.006724f
C3814 vdd.n2756 gnd 0.006724f
C3815 vdd.n2757 gnd 0.006724f
C3816 vdd.n2758 gnd 0.006724f
C3817 vdd.n2759 gnd 0.006724f
C3818 vdd.n2760 gnd 0.006724f
C3819 vdd.n2761 gnd 0.006724f
C3820 vdd.n2763 gnd 0.006724f
C3821 vdd.n2764 gnd 0.006724f
C3822 vdd.n2766 gnd 0.006724f
C3823 vdd.n2767 gnd 0.006724f
C3824 vdd.n2768 gnd 0.015955f
C3825 vdd.n2769 gnd 0.014896f
C3826 vdd.n2770 gnd 0.014896f
C3827 vdd.n2771 gnd 0.990313f
C3828 vdd.n2772 gnd 0.014896f
C3829 vdd.n2773 gnd 0.015955f
C3830 vdd.n2774 gnd 0.015136f
C3831 vdd.n2775 gnd 0.006724f
C3832 vdd.n2776 gnd 0.005191f
C3833 vdd.n2777 gnd 0.006724f
C3834 vdd.n2779 gnd 0.006724f
C3835 vdd.n2780 gnd 0.006724f
C3836 vdd.n2781 gnd 0.006724f
C3837 vdd.n2782 gnd 0.006724f
C3838 vdd.n2783 gnd 0.006724f
C3839 vdd.n2784 gnd 0.006724f
C3840 vdd.n2786 gnd 0.006724f
C3841 vdd.n2787 gnd 0.006724f
C3842 vdd.n2788 gnd 0.006724f
C3843 vdd.n2789 gnd 0.006724f
C3844 vdd.n2790 gnd 0.006724f
C3845 vdd.n2791 gnd 0.006724f
C3846 vdd.n2793 gnd 0.006724f
C3847 vdd.n2794 gnd 0.006724f
C3848 vdd.n2795 gnd 0.006724f
C3849 vdd.n2796 gnd 0.006724f
C3850 vdd.n2797 gnd 0.006724f
C3851 vdd.n2798 gnd 0.006724f
C3852 vdd.n2800 gnd 0.006724f
C3853 vdd.n2801 gnd 0.006724f
C3854 vdd.n2803 gnd 0.006724f
C3855 vdd.n2804 gnd 0.016158f
C3856 vdd.n2805 gnd 0.598448f
C3857 vdd.n2806 gnd 0.008504f
C3858 vdd.n2807 gnd 0.00378f
C3859 vdd.t134 gnd 0.12165f
C3860 vdd.t135 gnd 0.130011f
C3861 vdd.t133 gnd 0.158874f
C3862 vdd.n2808 gnd 0.203654f
C3863 vdd.n2809 gnd 0.171106f
C3864 vdd.n2810 gnd 0.012257f
C3865 vdd.n2811 gnd 0.009888f
C3866 vdd.n2812 gnd 0.004178f
C3867 vdd.n2813 gnd 0.007959f
C3868 vdd.n2814 gnd 0.009888f
C3869 vdd.n2815 gnd 0.009888f
C3870 vdd.n2816 gnd 0.007959f
C3871 vdd.n2817 gnd 0.007959f
C3872 vdd.n2818 gnd 0.009888f
C3873 vdd.n2820 gnd 0.009888f
C3874 vdd.n2821 gnd 0.007959f
C3875 vdd.n2822 gnd 0.007959f
C3876 vdd.n2823 gnd 0.007959f
C3877 vdd.n2824 gnd 0.009888f
C3878 vdd.n2826 gnd 0.009888f
C3879 vdd.n2828 gnd 0.009888f
C3880 vdd.n2829 gnd 0.007959f
C3881 vdd.n2830 gnd 0.007959f
C3882 vdd.n2831 gnd 0.007959f
C3883 vdd.n2832 gnd 0.009888f
C3884 vdd.n2834 gnd 0.009888f
C3885 vdd.n2836 gnd 0.009888f
C3886 vdd.n2837 gnd 0.007959f
C3887 vdd.n2838 gnd 0.007959f
C3888 vdd.n2839 gnd 0.007959f
C3889 vdd.n2840 gnd 0.009888f
C3890 vdd.n2842 gnd 0.009888f
C3891 vdd.n2843 gnd 0.009888f
C3892 vdd.n2844 gnd 0.007959f
C3893 vdd.n2845 gnd 0.007959f
C3894 vdd.n2846 gnd 0.009888f
C3895 vdd.n2847 gnd 0.009888f
C3896 vdd.n2849 gnd 0.009888f
C3897 vdd.n2850 gnd 0.007959f
C3898 vdd.n2851 gnd 0.009888f
C3899 vdd.n2852 gnd 0.009888f
C3900 vdd.n2853 gnd 0.009888f
C3901 vdd.n2854 gnd 0.016236f
C3902 vdd.n2855 gnd 0.005412f
C3903 vdd.n2856 gnd 0.009888f
C3904 vdd.n2858 gnd 0.009888f
C3905 vdd.n2860 gnd 0.009888f
C3906 vdd.n2861 gnd 0.007959f
C3907 vdd.n2862 gnd 0.007959f
C3908 vdd.n2863 gnd 0.007959f
C3909 vdd.n2864 gnd 0.009888f
C3910 vdd.n2866 gnd 0.009888f
C3911 vdd.n2868 gnd 0.009888f
C3912 vdd.n2869 gnd 0.007959f
C3913 vdd.n2870 gnd 0.007959f
C3914 vdd.n2871 gnd 0.007959f
C3915 vdd.n2872 gnd 0.009888f
C3916 vdd.n2874 gnd 0.009888f
C3917 vdd.n2876 gnd 0.009888f
C3918 vdd.n2877 gnd 0.007959f
C3919 vdd.n2878 gnd 0.007959f
C3920 vdd.n2879 gnd 0.007959f
C3921 vdd.n2880 gnd 0.009888f
C3922 vdd.n2882 gnd 0.009888f
C3923 vdd.n2884 gnd 0.009888f
C3924 vdd.n2885 gnd 0.007959f
C3925 vdd.n2886 gnd 0.007959f
C3926 vdd.n2887 gnd 0.007959f
C3927 vdd.n2888 gnd 0.009888f
C3928 vdd.n2890 gnd 0.009888f
C3929 vdd.n2892 gnd 0.009888f
C3930 vdd.n2893 gnd 0.007959f
C3931 vdd.n2894 gnd 0.007959f
C3932 vdd.n2895 gnd 0.006646f
C3933 vdd.n2896 gnd 0.009888f
C3934 vdd.n2898 gnd 0.009888f
C3935 vdd.n2900 gnd 0.009888f
C3936 vdd.n2901 gnd 0.006646f
C3937 vdd.n2902 gnd 0.007959f
C3938 vdd.n2903 gnd 0.007959f
C3939 vdd.n2904 gnd 0.009888f
C3940 vdd.n2906 gnd 0.009888f
C3941 vdd.n2908 gnd 0.009888f
C3942 vdd.n2909 gnd 0.007959f
C3943 vdd.n2910 gnd 0.007959f
C3944 vdd.n2911 gnd 0.007959f
C3945 vdd.n2912 gnd 0.009888f
C3946 vdd.n2914 gnd 0.009888f
C3947 vdd.n2916 gnd 0.009888f
C3948 vdd.n2917 gnd 0.007959f
C3949 vdd.n2918 gnd 0.007959f
C3950 vdd.n2919 gnd 0.007959f
C3951 vdd.n2920 gnd 0.009888f
C3952 vdd.n2922 gnd 0.009888f
C3953 vdd.n2923 gnd 0.009888f
C3954 vdd.n2924 gnd 0.007959f
C3955 vdd.n2925 gnd 0.007959f
C3956 vdd.n2926 gnd 0.009888f
C3957 vdd.n2927 gnd 0.009888f
C3958 vdd.n2928 gnd 0.007959f
C3959 vdd.n2929 gnd 0.007959f
C3960 vdd.n2930 gnd 0.009888f
C3961 vdd.n2931 gnd 0.009888f
C3962 vdd.n2933 gnd 0.009888f
C3963 vdd.n2934 gnd 0.007959f
C3964 vdd.n2935 gnd 0.006606f
C3965 vdd.n2936 gnd 0.023667f
C3966 vdd.n2937 gnd 0.023302f
C3967 vdd.n2938 gnd 0.006606f
C3968 vdd.n2939 gnd 0.023302f
C3969 vdd.n2940 gnd 1.38947f
C3970 vdd.n2941 gnd 0.023302f
C3971 vdd.n2942 gnd 0.006606f
C3972 vdd.n2943 gnd 0.023302f
C3973 vdd.n2944 gnd 0.009888f
C3974 vdd.n2945 gnd 0.009888f
C3975 vdd.n2946 gnd 0.007959f
C3976 vdd.n2947 gnd 0.009888f
C3977 vdd.n2948 gnd 1.01052f
C3978 vdd.n2949 gnd 0.009888f
C3979 vdd.n2950 gnd 0.007959f
C3980 vdd.n2951 gnd 0.009888f
C3981 vdd.n2952 gnd 0.009888f
C3982 vdd.n2953 gnd 0.009888f
C3983 vdd.n2954 gnd 0.007959f
C3984 vdd.n2955 gnd 0.009888f
C3985 vdd.n2956 gnd 0.894313f
C3986 vdd.n2957 gnd 0.009888f
C3987 vdd.n2958 gnd 0.007959f
C3988 vdd.n2959 gnd 0.009888f
C3989 vdd.n2960 gnd 0.009888f
C3990 vdd.n2961 gnd 0.009888f
C3991 vdd.n2962 gnd 0.007959f
C3992 vdd.n2963 gnd 0.009888f
C3993 vdd.t40 gnd 0.505262f
C3994 vdd.n2964 gnd 0.722524f
C3995 vdd.n2965 gnd 0.009888f
C3996 vdd.n2966 gnd 0.007959f
C3997 vdd.n2967 gnd 0.009888f
C3998 vdd.n2968 gnd 0.009888f
C3999 vdd.n2969 gnd 0.009888f
C4000 vdd.n2970 gnd 0.007959f
C4001 vdd.n2971 gnd 0.009888f
C4002 vdd.n2972 gnd 0.550735f
C4003 vdd.n2973 gnd 0.009888f
C4004 vdd.n2974 gnd 0.007959f
C4005 vdd.n2975 gnd 0.009888f
C4006 vdd.n2976 gnd 0.009888f
C4007 vdd.n2977 gnd 0.009888f
C4008 vdd.n2978 gnd 0.007959f
C4009 vdd.n2979 gnd 0.009888f
C4010 vdd.n2980 gnd 0.712419f
C4011 vdd.n2981 gnd 0.631577f
C4012 vdd.n2982 gnd 0.009888f
C4013 vdd.n2983 gnd 0.007959f
C4014 vdd.n2984 gnd 0.009888f
C4015 vdd.n2985 gnd 0.009888f
C4016 vdd.n2986 gnd 0.009888f
C4017 vdd.n2987 gnd 0.007959f
C4018 vdd.n2988 gnd 0.009888f
C4019 vdd.n2989 gnd 0.803366f
C4020 vdd.n2990 gnd 0.009888f
C4021 vdd.n2991 gnd 0.007959f
C4022 vdd.n2992 gnd 0.009888f
C4023 vdd.n2993 gnd 0.009888f
C4024 vdd.n2994 gnd 0.009888f
C4025 vdd.n2995 gnd 0.007959f
C4026 vdd.n2996 gnd 0.007959f
C4027 vdd.n2997 gnd 0.007959f
C4028 vdd.n2998 gnd 0.009888f
C4029 vdd.n2999 gnd 0.009888f
C4030 vdd.n3000 gnd 0.009888f
C4031 vdd.n3001 gnd 0.007959f
C4032 vdd.n3002 gnd 0.007959f
C4033 vdd.n3003 gnd 0.007959f
C4034 vdd.n3004 gnd 0.009888f
C4035 vdd.n3005 gnd 0.009888f
C4036 vdd.n3006 gnd 0.009888f
C4037 vdd.n3007 gnd 0.007959f
C4038 vdd.n3008 gnd 0.007959f
C4039 vdd.n3009 gnd 0.007959f
C4040 vdd.n3010 gnd 0.009888f
C4041 vdd.n3011 gnd 0.009888f
C4042 vdd.n3012 gnd 0.009888f
C4043 vdd.n3013 gnd 0.007959f
C4044 vdd.n3014 gnd 0.007959f
C4045 vdd.n3015 gnd 0.006606f
C4046 vdd.n3016 gnd 0.023302f
C4047 vdd.n3017 gnd 0.023667f
C4048 vdd.n3019 gnd 0.023667f
C4049 vdd.n3020 gnd 0.00378f
C4050 vdd.t145 gnd 0.12165f
C4051 vdd.t144 gnd 0.130011f
C4052 vdd.t143 gnd 0.158874f
C4053 vdd.n3021 gnd 0.203654f
C4054 vdd.n3022 gnd 0.171902f
C4055 vdd.n3023 gnd 0.013052f
C4056 vdd.n3024 gnd 0.004178f
C4057 vdd.n3025 gnd 0.007959f
C4058 vdd.n3026 gnd 0.009888f
C4059 vdd.n3028 gnd 0.009888f
C4060 vdd.n3029 gnd 0.009888f
C4061 vdd.n3030 gnd 0.007959f
C4062 vdd.n3031 gnd 0.007959f
C4063 vdd.n3032 gnd 0.007959f
C4064 vdd.n3033 gnd 0.009888f
C4065 vdd.n3035 gnd 0.009888f
C4066 vdd.n3036 gnd 0.009888f
C4067 vdd.n3037 gnd 0.007959f
C4068 vdd.n3038 gnd 0.007959f
C4069 vdd.n3039 gnd 0.007959f
C4070 vdd.n3040 gnd 0.009888f
C4071 vdd.n3042 gnd 0.009888f
C4072 vdd.n3043 gnd 0.009888f
C4073 vdd.n3044 gnd 0.007959f
C4074 vdd.n3045 gnd 0.007959f
C4075 vdd.n3046 gnd 0.007959f
C4076 vdd.n3047 gnd 0.009888f
C4077 vdd.n3049 gnd 0.009888f
C4078 vdd.n3050 gnd 0.009888f
C4079 vdd.n3051 gnd 0.007959f
C4080 vdd.n3052 gnd 0.007959f
C4081 vdd.n3053 gnd 0.007959f
C4082 vdd.n3054 gnd 0.009888f
C4083 vdd.n3056 gnd 0.009888f
C4084 vdd.n3057 gnd 0.009888f
C4085 vdd.n3058 gnd 0.007959f
C4086 vdd.n3059 gnd 0.009888f
C4087 vdd.n3060 gnd 0.009888f
C4088 vdd.n3061 gnd 0.009888f
C4089 vdd.n3062 gnd 0.017032f
C4090 vdd.n3063 gnd 0.005412f
C4091 vdd.n3064 gnd 0.007959f
C4092 vdd.n3065 gnd 0.009888f
C4093 vdd.n3067 gnd 0.009888f
C4094 vdd.n3068 gnd 0.009888f
C4095 vdd.n3069 gnd 0.007959f
C4096 vdd.n3070 gnd 0.007959f
C4097 vdd.n3071 gnd 0.007959f
C4098 vdd.n3072 gnd 0.009888f
C4099 vdd.n3074 gnd 0.009888f
C4100 vdd.n3075 gnd 0.009888f
C4101 vdd.n3076 gnd 0.007959f
C4102 vdd.n3077 gnd 0.007959f
C4103 vdd.n3078 gnd 0.007959f
C4104 vdd.n3079 gnd 0.009888f
C4105 vdd.n3081 gnd 0.009888f
C4106 vdd.n3082 gnd 0.009888f
C4107 vdd.n3083 gnd 0.007959f
C4108 vdd.n3084 gnd 0.007959f
C4109 vdd.n3085 gnd 0.007959f
C4110 vdd.n3086 gnd 0.009888f
C4111 vdd.n3088 gnd 0.009888f
C4112 vdd.n3089 gnd 0.009888f
C4113 vdd.n3090 gnd 0.007959f
C4114 vdd.n3091 gnd 0.007959f
C4115 vdd.n3092 gnd 0.007959f
C4116 vdd.n3093 gnd 0.009888f
C4117 vdd.n3095 gnd 0.009888f
C4118 vdd.n3096 gnd 0.009888f
C4119 vdd.n3097 gnd 0.007959f
C4120 vdd.n3098 gnd 0.009888f
C4121 vdd.n3099 gnd 0.009888f
C4122 vdd.n3100 gnd 0.009888f
C4123 vdd.n3101 gnd 0.017032f
C4124 vdd.n3102 gnd 0.006646f
C4125 vdd.n3103 gnd 0.007959f
C4126 vdd.n3104 gnd 0.009888f
C4127 vdd.n3106 gnd 0.009888f
C4128 vdd.n3107 gnd 0.009888f
C4129 vdd.n3108 gnd 0.007959f
C4130 vdd.n3109 gnd 0.007959f
C4131 vdd.n3110 gnd 0.007959f
C4132 vdd.n3111 gnd 0.009888f
C4133 vdd.n3113 gnd 0.009888f
C4134 vdd.n3114 gnd 0.009888f
C4135 vdd.n3115 gnd 0.007959f
C4136 vdd.n3116 gnd 0.007959f
C4137 vdd.n3117 gnd 0.007959f
C4138 vdd.n3118 gnd 0.009888f
C4139 vdd.n3120 gnd 0.009888f
C4140 vdd.n3121 gnd 0.009888f
C4141 vdd.n3122 gnd 0.007959f
C4142 vdd.n3123 gnd 0.007959f
C4143 vdd.n3124 gnd 0.007959f
C4144 vdd.n3125 gnd 0.009888f
C4145 vdd.n3127 gnd 0.009888f
C4146 vdd.n3128 gnd 0.009888f
C4147 vdd.n3130 gnd 0.009888f
C4148 vdd.n3131 gnd 0.007959f
C4149 vdd.n3132 gnd 0.007959f
C4150 vdd.n3133 gnd 0.006606f
C4151 vdd.n3134 gnd 0.023667f
C4152 vdd.n3135 gnd 0.023302f
C4153 vdd.n3136 gnd 0.006606f
C4154 vdd.n3137 gnd 0.023302f
C4155 vdd.n3138 gnd 1.42484f
C4156 vdd.n3139 gnd 0.570946f
C4157 vdd.t137 gnd 0.505262f
C4158 vdd.n3140 gnd 0.94484f
C4159 vdd.n3141 gnd 0.009888f
C4160 vdd.n3142 gnd 0.007959f
C4161 vdd.n3143 gnd 0.007959f
C4162 vdd.n3144 gnd 0.007959f
C4163 vdd.n3145 gnd 0.009888f
C4164 vdd.n3146 gnd 0.995366f
C4165 vdd.t10 gnd 0.505262f
C4166 vdd.n3147 gnd 0.52042f
C4167 vdd.n3148 gnd 0.823577f
C4168 vdd.n3149 gnd 0.009888f
C4169 vdd.n3150 gnd 0.007959f
C4170 vdd.n3151 gnd 0.007959f
C4171 vdd.n3152 gnd 0.007959f
C4172 vdd.n3153 gnd 0.009888f
C4173 vdd.n3154 gnd 0.651788f
C4174 vdd.t34 gnd 0.505262f
C4175 vdd.n3155 gnd 0.838735f
C4176 vdd.t19 gnd 0.505262f
C4177 vdd.n3156 gnd 0.530525f
C4178 vdd.n3157 gnd 0.009888f
C4179 vdd.n3158 gnd 0.007959f
C4180 vdd.n3159 gnd 0.007959f
C4181 vdd.n3160 gnd 0.007959f
C4182 vdd.n3161 gnd 0.009888f
C4183 vdd.n3162 gnd 0.702314f
C4184 vdd.n3163 gnd 0.641682f
C4185 vdd.t60 gnd 0.505262f
C4186 vdd.n3164 gnd 0.838735f
C4187 vdd.n3165 gnd 0.009888f
C4188 vdd.n3166 gnd 0.007959f
C4189 vdd.n3167 gnd 0.58862f
C4190 vdd.n3168 gnd 2.17886f
C4191 commonsourceibias.n0 gnd 0.010545f
C4192 commonsourceibias.t94 gnd 0.159685f
C4193 commonsourceibias.t109 gnd 0.147652f
C4194 commonsourceibias.n1 gnd 0.006423f
C4195 commonsourceibias.n2 gnd 0.007903f
C4196 commonsourceibias.t72 gnd 0.147652f
C4197 commonsourceibias.n3 gnd 0.008017f
C4198 commonsourceibias.n4 gnd 0.007903f
C4199 commonsourceibias.t70 gnd 0.147652f
C4200 commonsourceibias.n5 gnd 0.058913f
C4201 commonsourceibias.t102 gnd 0.147652f
C4202 commonsourceibias.n6 gnd 0.006393f
C4203 commonsourceibias.n7 gnd 0.007903f
C4204 commonsourceibias.t116 gnd 0.147652f
C4205 commonsourceibias.n8 gnd 0.00763f
C4206 commonsourceibias.n9 gnd 0.007903f
C4207 commonsourceibias.t66 gnd 0.147652f
C4208 commonsourceibias.n10 gnd 0.058913f
C4209 commonsourceibias.t92 gnd 0.147652f
C4210 commonsourceibias.n11 gnd 0.006383f
C4211 commonsourceibias.n12 gnd 0.010545f
C4212 commonsourceibias.t28 gnd 0.159685f
C4213 commonsourceibias.t48 gnd 0.147652f
C4214 commonsourceibias.n13 gnd 0.006423f
C4215 commonsourceibias.n14 gnd 0.007903f
C4216 commonsourceibias.t34 gnd 0.147652f
C4217 commonsourceibias.n15 gnd 0.008017f
C4218 commonsourceibias.n16 gnd 0.007903f
C4219 commonsourceibias.t26 gnd 0.147652f
C4220 commonsourceibias.n17 gnd 0.058913f
C4221 commonsourceibias.t44 gnd 0.147652f
C4222 commonsourceibias.n18 gnd 0.006393f
C4223 commonsourceibias.n19 gnd 0.007903f
C4224 commonsourceibias.t16 gnd 0.147652f
C4225 commonsourceibias.n20 gnd 0.00763f
C4226 commonsourceibias.n21 gnd 0.007903f
C4227 commonsourceibias.t12 gnd 0.147652f
C4228 commonsourceibias.n22 gnd 0.058913f
C4229 commonsourceibias.t36 gnd 0.147652f
C4230 commonsourceibias.n23 gnd 0.006383f
C4231 commonsourceibias.n24 gnd 0.007903f
C4232 commonsourceibias.t30 gnd 0.147652f
C4233 commonsourceibias.t4 gnd 0.147652f
C4234 commonsourceibias.n25 gnd 0.058913f
C4235 commonsourceibias.n26 gnd 0.007903f
C4236 commonsourceibias.t8 gnd 0.147652f
C4237 commonsourceibias.n27 gnd 0.058913f
C4238 commonsourceibias.n28 gnd 0.007903f
C4239 commonsourceibias.t14 gnd 0.147652f
C4240 commonsourceibias.n29 gnd 0.058913f
C4241 commonsourceibias.n30 gnd 0.007903f
C4242 commonsourceibias.t42 gnd 0.147652f
C4243 commonsourceibias.n31 gnd 0.008983f
C4244 commonsourceibias.n32 gnd 0.007903f
C4245 commonsourceibias.t18 gnd 0.147652f
C4246 commonsourceibias.n33 gnd 0.010623f
C4247 commonsourceibias.t0 gnd 0.164481f
C4248 commonsourceibias.t50 gnd 0.147652f
C4249 commonsourceibias.n34 gnd 0.065644f
C4250 commonsourceibias.n35 gnd 0.070328f
C4251 commonsourceibias.n36 gnd 0.033639f
C4252 commonsourceibias.n37 gnd 0.007903f
C4253 commonsourceibias.n38 gnd 0.006423f
C4254 commonsourceibias.n39 gnd 0.01089f
C4255 commonsourceibias.n40 gnd 0.058913f
C4256 commonsourceibias.n41 gnd 0.010937f
C4257 commonsourceibias.n42 gnd 0.007903f
C4258 commonsourceibias.n43 gnd 0.007903f
C4259 commonsourceibias.n44 gnd 0.007903f
C4260 commonsourceibias.n45 gnd 0.008017f
C4261 commonsourceibias.n46 gnd 0.058913f
C4262 commonsourceibias.n47 gnd 0.009741f
C4263 commonsourceibias.n48 gnd 0.010776f
C4264 commonsourceibias.n49 gnd 0.007903f
C4265 commonsourceibias.n50 gnd 0.007903f
C4266 commonsourceibias.n51 gnd 0.010705f
C4267 commonsourceibias.n52 gnd 0.006393f
C4268 commonsourceibias.n53 gnd 0.010838f
C4269 commonsourceibias.n54 gnd 0.007903f
C4270 commonsourceibias.n55 gnd 0.007903f
C4271 commonsourceibias.n56 gnd 0.010904f
C4272 commonsourceibias.n57 gnd 0.009403f
C4273 commonsourceibias.n58 gnd 0.00763f
C4274 commonsourceibias.n59 gnd 0.007903f
C4275 commonsourceibias.n60 gnd 0.007903f
C4276 commonsourceibias.n61 gnd 0.009667f
C4277 commonsourceibias.n62 gnd 0.01085f
C4278 commonsourceibias.n63 gnd 0.058913f
C4279 commonsourceibias.n64 gnd 0.010777f
C4280 commonsourceibias.n65 gnd 0.007903f
C4281 commonsourceibias.n66 gnd 0.007903f
C4282 commonsourceibias.n67 gnd 0.007903f
C4283 commonsourceibias.n68 gnd 0.010777f
C4284 commonsourceibias.n69 gnd 0.058913f
C4285 commonsourceibias.n70 gnd 0.01085f
C4286 commonsourceibias.n71 gnd 0.009667f
C4287 commonsourceibias.n72 gnd 0.007903f
C4288 commonsourceibias.n73 gnd 0.007903f
C4289 commonsourceibias.n74 gnd 0.007903f
C4290 commonsourceibias.n75 gnd 0.009403f
C4291 commonsourceibias.n76 gnd 0.010904f
C4292 commonsourceibias.n77 gnd 0.058913f
C4293 commonsourceibias.n78 gnd 0.010838f
C4294 commonsourceibias.n79 gnd 0.007903f
C4295 commonsourceibias.n80 gnd 0.007903f
C4296 commonsourceibias.n81 gnd 0.007903f
C4297 commonsourceibias.n82 gnd 0.010705f
C4298 commonsourceibias.n83 gnd 0.058913f
C4299 commonsourceibias.n84 gnd 0.010776f
C4300 commonsourceibias.n85 gnd 0.009741f
C4301 commonsourceibias.n86 gnd 0.007903f
C4302 commonsourceibias.n87 gnd 0.007903f
C4303 commonsourceibias.n88 gnd 0.007903f
C4304 commonsourceibias.n89 gnd 0.008983f
C4305 commonsourceibias.n90 gnd 0.010937f
C4306 commonsourceibias.n91 gnd 0.058913f
C4307 commonsourceibias.n92 gnd 0.01089f
C4308 commonsourceibias.n93 gnd 0.007903f
C4309 commonsourceibias.n94 gnd 0.007903f
C4310 commonsourceibias.n95 gnd 0.007903f
C4311 commonsourceibias.n96 gnd 0.010623f
C4312 commonsourceibias.n97 gnd 0.058913f
C4313 commonsourceibias.n98 gnd 0.010649f
C4314 commonsourceibias.n99 gnd 0.071041f
C4315 commonsourceibias.n100 gnd 0.079434f
C4316 commonsourceibias.t29 gnd 0.017054f
C4317 commonsourceibias.t49 gnd 0.017054f
C4318 commonsourceibias.n101 gnd 0.150693f
C4319 commonsourceibias.n102 gnd 0.130533f
C4320 commonsourceibias.t35 gnd 0.017054f
C4321 commonsourceibias.t27 gnd 0.017054f
C4322 commonsourceibias.n103 gnd 0.150693f
C4323 commonsourceibias.n104 gnd 0.069219f
C4324 commonsourceibias.t45 gnd 0.017054f
C4325 commonsourceibias.t17 gnd 0.017054f
C4326 commonsourceibias.n105 gnd 0.150693f
C4327 commonsourceibias.n106 gnd 0.069219f
C4328 commonsourceibias.t13 gnd 0.017054f
C4329 commonsourceibias.t37 gnd 0.017054f
C4330 commonsourceibias.n107 gnd 0.150693f
C4331 commonsourceibias.n108 gnd 0.057829f
C4332 commonsourceibias.t51 gnd 0.017054f
C4333 commonsourceibias.t1 gnd 0.017054f
C4334 commonsourceibias.n109 gnd 0.151197f
C4335 commonsourceibias.t43 gnd 0.017054f
C4336 commonsourceibias.t19 gnd 0.017054f
C4337 commonsourceibias.n110 gnd 0.150693f
C4338 commonsourceibias.n111 gnd 0.140418f
C4339 commonsourceibias.t9 gnd 0.017054f
C4340 commonsourceibias.t15 gnd 0.017054f
C4341 commonsourceibias.n112 gnd 0.150693f
C4342 commonsourceibias.n113 gnd 0.069219f
C4343 commonsourceibias.t31 gnd 0.017054f
C4344 commonsourceibias.t5 gnd 0.017054f
C4345 commonsourceibias.n114 gnd 0.150693f
C4346 commonsourceibias.n115 gnd 0.057829f
C4347 commonsourceibias.n116 gnd 0.070025f
C4348 commonsourceibias.n117 gnd 0.007903f
C4349 commonsourceibias.t89 gnd 0.147652f
C4350 commonsourceibias.t105 gnd 0.147652f
C4351 commonsourceibias.n118 gnd 0.058913f
C4352 commonsourceibias.n119 gnd 0.007903f
C4353 commonsourceibias.t85 gnd 0.147652f
C4354 commonsourceibias.n120 gnd 0.058913f
C4355 commonsourceibias.n121 gnd 0.007903f
C4356 commonsourceibias.t82 gnd 0.147652f
C4357 commonsourceibias.n122 gnd 0.058913f
C4358 commonsourceibias.n123 gnd 0.007903f
C4359 commonsourceibias.t97 gnd 0.147652f
C4360 commonsourceibias.n124 gnd 0.008983f
C4361 commonsourceibias.n125 gnd 0.007903f
C4362 commonsourceibias.t111 gnd 0.147652f
C4363 commonsourceibias.n126 gnd 0.010623f
C4364 commonsourceibias.t88 gnd 0.164481f
C4365 commonsourceibias.t75 gnd 0.147652f
C4366 commonsourceibias.n127 gnd 0.065644f
C4367 commonsourceibias.n128 gnd 0.070328f
C4368 commonsourceibias.n129 gnd 0.033639f
C4369 commonsourceibias.n130 gnd 0.007903f
C4370 commonsourceibias.n131 gnd 0.006423f
C4371 commonsourceibias.n132 gnd 0.01089f
C4372 commonsourceibias.n133 gnd 0.058913f
C4373 commonsourceibias.n134 gnd 0.010937f
C4374 commonsourceibias.n135 gnd 0.007903f
C4375 commonsourceibias.n136 gnd 0.007903f
C4376 commonsourceibias.n137 gnd 0.007903f
C4377 commonsourceibias.n138 gnd 0.008017f
C4378 commonsourceibias.n139 gnd 0.058913f
C4379 commonsourceibias.n140 gnd 0.009741f
C4380 commonsourceibias.n141 gnd 0.010776f
C4381 commonsourceibias.n142 gnd 0.007903f
C4382 commonsourceibias.n143 gnd 0.007903f
C4383 commonsourceibias.n144 gnd 0.010705f
C4384 commonsourceibias.n145 gnd 0.006393f
C4385 commonsourceibias.n146 gnd 0.010838f
C4386 commonsourceibias.n147 gnd 0.007903f
C4387 commonsourceibias.n148 gnd 0.007903f
C4388 commonsourceibias.n149 gnd 0.010904f
C4389 commonsourceibias.n150 gnd 0.009403f
C4390 commonsourceibias.n151 gnd 0.00763f
C4391 commonsourceibias.n152 gnd 0.007903f
C4392 commonsourceibias.n153 gnd 0.007903f
C4393 commonsourceibias.n154 gnd 0.009667f
C4394 commonsourceibias.n155 gnd 0.01085f
C4395 commonsourceibias.n156 gnd 0.058913f
C4396 commonsourceibias.n157 gnd 0.010777f
C4397 commonsourceibias.n158 gnd 0.007865f
C4398 commonsourceibias.n159 gnd 0.057129f
C4399 commonsourceibias.n160 gnd 0.007865f
C4400 commonsourceibias.n161 gnd 0.010777f
C4401 commonsourceibias.n162 gnd 0.058913f
C4402 commonsourceibias.n163 gnd 0.01085f
C4403 commonsourceibias.n164 gnd 0.009667f
C4404 commonsourceibias.n165 gnd 0.007903f
C4405 commonsourceibias.n166 gnd 0.007903f
C4406 commonsourceibias.n167 gnd 0.007903f
C4407 commonsourceibias.n168 gnd 0.009403f
C4408 commonsourceibias.n169 gnd 0.010904f
C4409 commonsourceibias.n170 gnd 0.058913f
C4410 commonsourceibias.n171 gnd 0.010838f
C4411 commonsourceibias.n172 gnd 0.007903f
C4412 commonsourceibias.n173 gnd 0.007903f
C4413 commonsourceibias.n174 gnd 0.007903f
C4414 commonsourceibias.n175 gnd 0.010705f
C4415 commonsourceibias.n176 gnd 0.058913f
C4416 commonsourceibias.n177 gnd 0.010776f
C4417 commonsourceibias.n178 gnd 0.009741f
C4418 commonsourceibias.n179 gnd 0.007903f
C4419 commonsourceibias.n180 gnd 0.007903f
C4420 commonsourceibias.n181 gnd 0.007903f
C4421 commonsourceibias.n182 gnd 0.008983f
C4422 commonsourceibias.n183 gnd 0.010937f
C4423 commonsourceibias.n184 gnd 0.058913f
C4424 commonsourceibias.n185 gnd 0.01089f
C4425 commonsourceibias.n186 gnd 0.007903f
C4426 commonsourceibias.n187 gnd 0.007903f
C4427 commonsourceibias.n188 gnd 0.007903f
C4428 commonsourceibias.n189 gnd 0.010623f
C4429 commonsourceibias.n190 gnd 0.058913f
C4430 commonsourceibias.n191 gnd 0.010649f
C4431 commonsourceibias.n192 gnd 0.071041f
C4432 commonsourceibias.n193 gnd 0.046914f
C4433 commonsourceibias.n194 gnd 0.010545f
C4434 commonsourceibias.t96 gnd 0.147652f
C4435 commonsourceibias.n195 gnd 0.006423f
C4436 commonsourceibias.n196 gnd 0.007903f
C4437 commonsourceibias.t65 gnd 0.147652f
C4438 commonsourceibias.n197 gnd 0.008017f
C4439 commonsourceibias.n198 gnd 0.007903f
C4440 commonsourceibias.t127 gnd 0.147652f
C4441 commonsourceibias.n199 gnd 0.058913f
C4442 commonsourceibias.t87 gnd 0.147652f
C4443 commonsourceibias.n200 gnd 0.006393f
C4444 commonsourceibias.n201 gnd 0.007903f
C4445 commonsourceibias.t104 gnd 0.147652f
C4446 commonsourceibias.n202 gnd 0.00763f
C4447 commonsourceibias.n203 gnd 0.007903f
C4448 commonsourceibias.t122 gnd 0.147652f
C4449 commonsourceibias.n204 gnd 0.058913f
C4450 commonsourceibias.t80 gnd 0.147652f
C4451 commonsourceibias.n205 gnd 0.006383f
C4452 commonsourceibias.n206 gnd 0.007903f
C4453 commonsourceibias.t76 gnd 0.147652f
C4454 commonsourceibias.t90 gnd 0.147652f
C4455 commonsourceibias.n207 gnd 0.058913f
C4456 commonsourceibias.n208 gnd 0.007903f
C4457 commonsourceibias.t74 gnd 0.147652f
C4458 commonsourceibias.n209 gnd 0.058913f
C4459 commonsourceibias.n210 gnd 0.007903f
C4460 commonsourceibias.t71 gnd 0.147652f
C4461 commonsourceibias.n211 gnd 0.058913f
C4462 commonsourceibias.n212 gnd 0.007903f
C4463 commonsourceibias.t83 gnd 0.147652f
C4464 commonsourceibias.n213 gnd 0.008983f
C4465 commonsourceibias.n214 gnd 0.007903f
C4466 commonsourceibias.t98 gnd 0.147652f
C4467 commonsourceibias.n215 gnd 0.010623f
C4468 commonsourceibias.t77 gnd 0.164481f
C4469 commonsourceibias.t67 gnd 0.147652f
C4470 commonsourceibias.n216 gnd 0.065644f
C4471 commonsourceibias.n217 gnd 0.070328f
C4472 commonsourceibias.n218 gnd 0.033639f
C4473 commonsourceibias.n219 gnd 0.007903f
C4474 commonsourceibias.n220 gnd 0.006423f
C4475 commonsourceibias.n221 gnd 0.01089f
C4476 commonsourceibias.n222 gnd 0.058913f
C4477 commonsourceibias.n223 gnd 0.010937f
C4478 commonsourceibias.n224 gnd 0.007903f
C4479 commonsourceibias.n225 gnd 0.007903f
C4480 commonsourceibias.n226 gnd 0.007903f
C4481 commonsourceibias.n227 gnd 0.008017f
C4482 commonsourceibias.n228 gnd 0.058913f
C4483 commonsourceibias.n229 gnd 0.009741f
C4484 commonsourceibias.n230 gnd 0.010776f
C4485 commonsourceibias.n231 gnd 0.007903f
C4486 commonsourceibias.n232 gnd 0.007903f
C4487 commonsourceibias.n233 gnd 0.010705f
C4488 commonsourceibias.n234 gnd 0.006393f
C4489 commonsourceibias.n235 gnd 0.010838f
C4490 commonsourceibias.n236 gnd 0.007903f
C4491 commonsourceibias.n237 gnd 0.007903f
C4492 commonsourceibias.n238 gnd 0.010904f
C4493 commonsourceibias.n239 gnd 0.009403f
C4494 commonsourceibias.n240 gnd 0.00763f
C4495 commonsourceibias.n241 gnd 0.007903f
C4496 commonsourceibias.n242 gnd 0.007903f
C4497 commonsourceibias.n243 gnd 0.009667f
C4498 commonsourceibias.n244 gnd 0.01085f
C4499 commonsourceibias.n245 gnd 0.058913f
C4500 commonsourceibias.n246 gnd 0.010777f
C4501 commonsourceibias.n247 gnd 0.007903f
C4502 commonsourceibias.n248 gnd 0.007903f
C4503 commonsourceibias.n249 gnd 0.007903f
C4504 commonsourceibias.n250 gnd 0.010777f
C4505 commonsourceibias.n251 gnd 0.058913f
C4506 commonsourceibias.n252 gnd 0.01085f
C4507 commonsourceibias.n253 gnd 0.009667f
C4508 commonsourceibias.n254 gnd 0.007903f
C4509 commonsourceibias.n255 gnd 0.007903f
C4510 commonsourceibias.n256 gnd 0.007903f
C4511 commonsourceibias.n257 gnd 0.009403f
C4512 commonsourceibias.n258 gnd 0.010904f
C4513 commonsourceibias.n259 gnd 0.058913f
C4514 commonsourceibias.n260 gnd 0.010838f
C4515 commonsourceibias.n261 gnd 0.007903f
C4516 commonsourceibias.n262 gnd 0.007903f
C4517 commonsourceibias.n263 gnd 0.007903f
C4518 commonsourceibias.n264 gnd 0.010705f
C4519 commonsourceibias.n265 gnd 0.058913f
C4520 commonsourceibias.n266 gnd 0.010776f
C4521 commonsourceibias.n267 gnd 0.009741f
C4522 commonsourceibias.n268 gnd 0.007903f
C4523 commonsourceibias.n269 gnd 0.007903f
C4524 commonsourceibias.n270 gnd 0.007903f
C4525 commonsourceibias.n271 gnd 0.008983f
C4526 commonsourceibias.n272 gnd 0.010937f
C4527 commonsourceibias.n273 gnd 0.058913f
C4528 commonsourceibias.n274 gnd 0.01089f
C4529 commonsourceibias.n275 gnd 0.007903f
C4530 commonsourceibias.n276 gnd 0.007903f
C4531 commonsourceibias.n277 gnd 0.007903f
C4532 commonsourceibias.n278 gnd 0.010623f
C4533 commonsourceibias.n279 gnd 0.058913f
C4534 commonsourceibias.n280 gnd 0.010649f
C4535 commonsourceibias.t81 gnd 0.159685f
C4536 commonsourceibias.n281 gnd 0.071041f
C4537 commonsourceibias.n282 gnd 0.02535f
C4538 commonsourceibias.n283 gnd 0.398385f
C4539 commonsourceibias.n284 gnd 0.010545f
C4540 commonsourceibias.t113 gnd 0.159685f
C4541 commonsourceibias.t123 gnd 0.147652f
C4542 commonsourceibias.n285 gnd 0.006423f
C4543 commonsourceibias.n286 gnd 0.007903f
C4544 commonsourceibias.t68 gnd 0.147652f
C4545 commonsourceibias.n287 gnd 0.008017f
C4546 commonsourceibias.n288 gnd 0.007903f
C4547 commonsourceibias.t119 gnd 0.147652f
C4548 commonsourceibias.n289 gnd 0.006393f
C4549 commonsourceibias.n290 gnd 0.007903f
C4550 commonsourceibias.t64 gnd 0.147652f
C4551 commonsourceibias.n291 gnd 0.00763f
C4552 commonsourceibias.n292 gnd 0.007903f
C4553 commonsourceibias.t112 gnd 0.147652f
C4554 commonsourceibias.n293 gnd 0.006383f
C4555 commonsourceibias.n294 gnd 0.007903f
C4556 commonsourceibias.t107 gnd 0.147652f
C4557 commonsourceibias.t121 gnd 0.147652f
C4558 commonsourceibias.n295 gnd 0.058913f
C4559 commonsourceibias.n296 gnd 0.007903f
C4560 commonsourceibias.t78 gnd 0.147652f
C4561 commonsourceibias.n297 gnd 0.058913f
C4562 commonsourceibias.n298 gnd 0.007903f
C4563 commonsourceibias.t101 gnd 0.147652f
C4564 commonsourceibias.n299 gnd 0.058913f
C4565 commonsourceibias.n300 gnd 0.007903f
C4566 commonsourceibias.t115 gnd 0.147652f
C4567 commonsourceibias.n301 gnd 0.008983f
C4568 commonsourceibias.n302 gnd 0.007903f
C4569 commonsourceibias.t125 gnd 0.147652f
C4570 commonsourceibias.n303 gnd 0.010623f
C4571 commonsourceibias.t108 gnd 0.164481f
C4572 commonsourceibias.t91 gnd 0.147652f
C4573 commonsourceibias.n304 gnd 0.065644f
C4574 commonsourceibias.n305 gnd 0.070328f
C4575 commonsourceibias.n306 gnd 0.033639f
C4576 commonsourceibias.n307 gnd 0.007903f
C4577 commonsourceibias.n308 gnd 0.006423f
C4578 commonsourceibias.n309 gnd 0.01089f
C4579 commonsourceibias.n310 gnd 0.058913f
C4580 commonsourceibias.n311 gnd 0.010937f
C4581 commonsourceibias.n312 gnd 0.007903f
C4582 commonsourceibias.n313 gnd 0.007903f
C4583 commonsourceibias.n314 gnd 0.007903f
C4584 commonsourceibias.n315 gnd 0.008017f
C4585 commonsourceibias.n316 gnd 0.058913f
C4586 commonsourceibias.n317 gnd 0.009741f
C4587 commonsourceibias.n318 gnd 0.010776f
C4588 commonsourceibias.n319 gnd 0.007903f
C4589 commonsourceibias.n320 gnd 0.007903f
C4590 commonsourceibias.n321 gnd 0.010705f
C4591 commonsourceibias.n322 gnd 0.006393f
C4592 commonsourceibias.n323 gnd 0.010838f
C4593 commonsourceibias.n324 gnd 0.007903f
C4594 commonsourceibias.n325 gnd 0.007903f
C4595 commonsourceibias.n326 gnd 0.010904f
C4596 commonsourceibias.n327 gnd 0.009403f
C4597 commonsourceibias.n328 gnd 0.00763f
C4598 commonsourceibias.n329 gnd 0.007903f
C4599 commonsourceibias.n330 gnd 0.007903f
C4600 commonsourceibias.n331 gnd 0.009667f
C4601 commonsourceibias.n332 gnd 0.01085f
C4602 commonsourceibias.n333 gnd 0.058913f
C4603 commonsourceibias.n334 gnd 0.010777f
C4604 commonsourceibias.n335 gnd 0.007865f
C4605 commonsourceibias.t23 gnd 0.017054f
C4606 commonsourceibias.t41 gnd 0.017054f
C4607 commonsourceibias.n336 gnd 0.151197f
C4608 commonsourceibias.t3 gnd 0.017054f
C4609 commonsourceibias.t33 gnd 0.017054f
C4610 commonsourceibias.n337 gnd 0.150693f
C4611 commonsourceibias.n338 gnd 0.140418f
C4612 commonsourceibias.t61 gnd 0.017054f
C4613 commonsourceibias.t59 gnd 0.017054f
C4614 commonsourceibias.n339 gnd 0.150693f
C4615 commonsourceibias.n340 gnd 0.069219f
C4616 commonsourceibias.t47 gnd 0.017054f
C4617 commonsourceibias.t55 gnd 0.017054f
C4618 commonsourceibias.n341 gnd 0.150693f
C4619 commonsourceibias.n342 gnd 0.057829f
C4620 commonsourceibias.n343 gnd 0.010545f
C4621 commonsourceibias.t38 gnd 0.147652f
C4622 commonsourceibias.n344 gnd 0.006423f
C4623 commonsourceibias.n345 gnd 0.007903f
C4624 commonsourceibias.t20 gnd 0.147652f
C4625 commonsourceibias.n346 gnd 0.008017f
C4626 commonsourceibias.n347 gnd 0.007903f
C4627 commonsourceibias.t24 gnd 0.147652f
C4628 commonsourceibias.n348 gnd 0.006393f
C4629 commonsourceibias.n349 gnd 0.007903f
C4630 commonsourceibias.t56 gnd 0.147652f
C4631 commonsourceibias.n350 gnd 0.00763f
C4632 commonsourceibias.n351 gnd 0.007903f
C4633 commonsourceibias.t10 gnd 0.147652f
C4634 commonsourceibias.n352 gnd 0.006383f
C4635 commonsourceibias.n353 gnd 0.007903f
C4636 commonsourceibias.t54 gnd 0.147652f
C4637 commonsourceibias.t46 gnd 0.147652f
C4638 commonsourceibias.n354 gnd 0.058913f
C4639 commonsourceibias.n355 gnd 0.007903f
C4640 commonsourceibias.t58 gnd 0.147652f
C4641 commonsourceibias.n356 gnd 0.058913f
C4642 commonsourceibias.n357 gnd 0.007903f
C4643 commonsourceibias.t60 gnd 0.147652f
C4644 commonsourceibias.n358 gnd 0.058913f
C4645 commonsourceibias.n359 gnd 0.007903f
C4646 commonsourceibias.t32 gnd 0.147652f
C4647 commonsourceibias.n360 gnd 0.008983f
C4648 commonsourceibias.n361 gnd 0.007903f
C4649 commonsourceibias.t2 gnd 0.147652f
C4650 commonsourceibias.n362 gnd 0.010623f
C4651 commonsourceibias.t22 gnd 0.164481f
C4652 commonsourceibias.t40 gnd 0.147652f
C4653 commonsourceibias.n363 gnd 0.065644f
C4654 commonsourceibias.n364 gnd 0.070328f
C4655 commonsourceibias.n365 gnd 0.033639f
C4656 commonsourceibias.n366 gnd 0.007903f
C4657 commonsourceibias.n367 gnd 0.006423f
C4658 commonsourceibias.n368 gnd 0.01089f
C4659 commonsourceibias.n369 gnd 0.058913f
C4660 commonsourceibias.n370 gnd 0.010937f
C4661 commonsourceibias.n371 gnd 0.007903f
C4662 commonsourceibias.n372 gnd 0.007903f
C4663 commonsourceibias.n373 gnd 0.007903f
C4664 commonsourceibias.n374 gnd 0.008017f
C4665 commonsourceibias.n375 gnd 0.058913f
C4666 commonsourceibias.n376 gnd 0.009741f
C4667 commonsourceibias.n377 gnd 0.010776f
C4668 commonsourceibias.n378 gnd 0.007903f
C4669 commonsourceibias.n379 gnd 0.007903f
C4670 commonsourceibias.n380 gnd 0.010705f
C4671 commonsourceibias.n381 gnd 0.006393f
C4672 commonsourceibias.n382 gnd 0.010838f
C4673 commonsourceibias.n383 gnd 0.007903f
C4674 commonsourceibias.n384 gnd 0.007903f
C4675 commonsourceibias.n385 gnd 0.010904f
C4676 commonsourceibias.n386 gnd 0.009403f
C4677 commonsourceibias.n387 gnd 0.00763f
C4678 commonsourceibias.n388 gnd 0.007903f
C4679 commonsourceibias.n389 gnd 0.007903f
C4680 commonsourceibias.n390 gnd 0.009667f
C4681 commonsourceibias.n391 gnd 0.01085f
C4682 commonsourceibias.n392 gnd 0.058913f
C4683 commonsourceibias.n393 gnd 0.010777f
C4684 commonsourceibias.n394 gnd 0.007903f
C4685 commonsourceibias.n395 gnd 0.007903f
C4686 commonsourceibias.n396 gnd 0.007903f
C4687 commonsourceibias.n397 gnd 0.010777f
C4688 commonsourceibias.n398 gnd 0.058913f
C4689 commonsourceibias.n399 gnd 0.01085f
C4690 commonsourceibias.t6 gnd 0.147652f
C4691 commonsourceibias.n400 gnd 0.058913f
C4692 commonsourceibias.n401 gnd 0.009667f
C4693 commonsourceibias.n402 gnd 0.007903f
C4694 commonsourceibias.n403 gnd 0.007903f
C4695 commonsourceibias.n404 gnd 0.007903f
C4696 commonsourceibias.n405 gnd 0.009403f
C4697 commonsourceibias.n406 gnd 0.010904f
C4698 commonsourceibias.n407 gnd 0.058913f
C4699 commonsourceibias.n408 gnd 0.010838f
C4700 commonsourceibias.n409 gnd 0.007903f
C4701 commonsourceibias.n410 gnd 0.007903f
C4702 commonsourceibias.n411 gnd 0.007903f
C4703 commonsourceibias.n412 gnd 0.010705f
C4704 commonsourceibias.n413 gnd 0.058913f
C4705 commonsourceibias.n414 gnd 0.010776f
C4706 commonsourceibias.t62 gnd 0.147652f
C4707 commonsourceibias.n415 gnd 0.058913f
C4708 commonsourceibias.n416 gnd 0.009741f
C4709 commonsourceibias.n417 gnd 0.007903f
C4710 commonsourceibias.n418 gnd 0.007903f
C4711 commonsourceibias.n419 gnd 0.007903f
C4712 commonsourceibias.n420 gnd 0.008983f
C4713 commonsourceibias.n421 gnd 0.010937f
C4714 commonsourceibias.n422 gnd 0.058913f
C4715 commonsourceibias.n423 gnd 0.01089f
C4716 commonsourceibias.n424 gnd 0.007903f
C4717 commonsourceibias.n425 gnd 0.007903f
C4718 commonsourceibias.n426 gnd 0.007903f
C4719 commonsourceibias.n427 gnd 0.010623f
C4720 commonsourceibias.n428 gnd 0.058913f
C4721 commonsourceibias.n429 gnd 0.010649f
C4722 commonsourceibias.t52 gnd 0.159685f
C4723 commonsourceibias.n430 gnd 0.071041f
C4724 commonsourceibias.n431 gnd 0.079434f
C4725 commonsourceibias.t39 gnd 0.017054f
C4726 commonsourceibias.t53 gnd 0.017054f
C4727 commonsourceibias.n432 gnd 0.150693f
C4728 commonsourceibias.n433 gnd 0.130533f
C4729 commonsourceibias.t63 gnd 0.017054f
C4730 commonsourceibias.t21 gnd 0.017054f
C4731 commonsourceibias.n434 gnd 0.150693f
C4732 commonsourceibias.n435 gnd 0.069219f
C4733 commonsourceibias.t57 gnd 0.017054f
C4734 commonsourceibias.t25 gnd 0.017054f
C4735 commonsourceibias.n436 gnd 0.150693f
C4736 commonsourceibias.n437 gnd 0.069219f
C4737 commonsourceibias.t11 gnd 0.017054f
C4738 commonsourceibias.t7 gnd 0.017054f
C4739 commonsourceibias.n438 gnd 0.150693f
C4740 commonsourceibias.n439 gnd 0.057829f
C4741 commonsourceibias.n440 gnd 0.070025f
C4742 commonsourceibias.n441 gnd 0.057129f
C4743 commonsourceibias.n442 gnd 0.007865f
C4744 commonsourceibias.n443 gnd 0.010777f
C4745 commonsourceibias.n444 gnd 0.058913f
C4746 commonsourceibias.n445 gnd 0.01085f
C4747 commonsourceibias.t126 gnd 0.147652f
C4748 commonsourceibias.n446 gnd 0.058913f
C4749 commonsourceibias.n447 gnd 0.009667f
C4750 commonsourceibias.n448 gnd 0.007903f
C4751 commonsourceibias.n449 gnd 0.007903f
C4752 commonsourceibias.n450 gnd 0.007903f
C4753 commonsourceibias.n451 gnd 0.009403f
C4754 commonsourceibias.n452 gnd 0.010904f
C4755 commonsourceibias.n453 gnd 0.058913f
C4756 commonsourceibias.n454 gnd 0.010838f
C4757 commonsourceibias.n455 gnd 0.007903f
C4758 commonsourceibias.n456 gnd 0.007903f
C4759 commonsourceibias.n457 gnd 0.007903f
C4760 commonsourceibias.n458 gnd 0.010705f
C4761 commonsourceibias.n459 gnd 0.058913f
C4762 commonsourceibias.n460 gnd 0.010776f
C4763 commonsourceibias.t84 gnd 0.147652f
C4764 commonsourceibias.n461 gnd 0.058913f
C4765 commonsourceibias.n462 gnd 0.009741f
C4766 commonsourceibias.n463 gnd 0.007903f
C4767 commonsourceibias.n464 gnd 0.007903f
C4768 commonsourceibias.n465 gnd 0.007903f
C4769 commonsourceibias.n466 gnd 0.008983f
C4770 commonsourceibias.n467 gnd 0.010937f
C4771 commonsourceibias.n468 gnd 0.058913f
C4772 commonsourceibias.n469 gnd 0.01089f
C4773 commonsourceibias.n470 gnd 0.007903f
C4774 commonsourceibias.n471 gnd 0.007903f
C4775 commonsourceibias.n472 gnd 0.007903f
C4776 commonsourceibias.n473 gnd 0.010623f
C4777 commonsourceibias.n474 gnd 0.058913f
C4778 commonsourceibias.n475 gnd 0.010649f
C4779 commonsourceibias.n476 gnd 0.071041f
C4780 commonsourceibias.n477 gnd 0.046914f
C4781 commonsourceibias.n478 gnd 0.010545f
C4782 commonsourceibias.t114 gnd 0.147652f
C4783 commonsourceibias.n479 gnd 0.006423f
C4784 commonsourceibias.n480 gnd 0.007903f
C4785 commonsourceibias.t124 gnd 0.147652f
C4786 commonsourceibias.n481 gnd 0.008017f
C4787 commonsourceibias.n482 gnd 0.007903f
C4788 commonsourceibias.t106 gnd 0.147652f
C4789 commonsourceibias.n483 gnd 0.006393f
C4790 commonsourceibias.n484 gnd 0.007903f
C4791 commonsourceibias.t120 gnd 0.147652f
C4792 commonsourceibias.n485 gnd 0.00763f
C4793 commonsourceibias.n486 gnd 0.007903f
C4794 commonsourceibias.t100 gnd 0.147652f
C4795 commonsourceibias.n487 gnd 0.006383f
C4796 commonsourceibias.n488 gnd 0.007903f
C4797 commonsourceibias.t93 gnd 0.147652f
C4798 commonsourceibias.t110 gnd 0.147652f
C4799 commonsourceibias.n489 gnd 0.058913f
C4800 commonsourceibias.n490 gnd 0.007903f
C4801 commonsourceibias.t69 gnd 0.147652f
C4802 commonsourceibias.n491 gnd 0.058913f
C4803 commonsourceibias.n492 gnd 0.007903f
C4804 commonsourceibias.t86 gnd 0.147652f
C4805 commonsourceibias.n493 gnd 0.058913f
C4806 commonsourceibias.n494 gnd 0.007903f
C4807 commonsourceibias.t103 gnd 0.147652f
C4808 commonsourceibias.n495 gnd 0.008983f
C4809 commonsourceibias.n496 gnd 0.007903f
C4810 commonsourceibias.t118 gnd 0.147652f
C4811 commonsourceibias.n497 gnd 0.010623f
C4812 commonsourceibias.t95 gnd 0.164481f
C4813 commonsourceibias.t79 gnd 0.147652f
C4814 commonsourceibias.n498 gnd 0.065644f
C4815 commonsourceibias.n499 gnd 0.070328f
C4816 commonsourceibias.n500 gnd 0.033639f
C4817 commonsourceibias.n501 gnd 0.007903f
C4818 commonsourceibias.n502 gnd 0.006423f
C4819 commonsourceibias.n503 gnd 0.01089f
C4820 commonsourceibias.n504 gnd 0.058913f
C4821 commonsourceibias.n505 gnd 0.010937f
C4822 commonsourceibias.n506 gnd 0.007903f
C4823 commonsourceibias.n507 gnd 0.007903f
C4824 commonsourceibias.n508 gnd 0.007903f
C4825 commonsourceibias.n509 gnd 0.008017f
C4826 commonsourceibias.n510 gnd 0.058913f
C4827 commonsourceibias.n511 gnd 0.009741f
C4828 commonsourceibias.n512 gnd 0.010776f
C4829 commonsourceibias.n513 gnd 0.007903f
C4830 commonsourceibias.n514 gnd 0.007903f
C4831 commonsourceibias.n515 gnd 0.010705f
C4832 commonsourceibias.n516 gnd 0.006393f
C4833 commonsourceibias.n517 gnd 0.010838f
C4834 commonsourceibias.n518 gnd 0.007903f
C4835 commonsourceibias.n519 gnd 0.007903f
C4836 commonsourceibias.n520 gnd 0.010904f
C4837 commonsourceibias.n521 gnd 0.009403f
C4838 commonsourceibias.n522 gnd 0.00763f
C4839 commonsourceibias.n523 gnd 0.007903f
C4840 commonsourceibias.n524 gnd 0.007903f
C4841 commonsourceibias.n525 gnd 0.009667f
C4842 commonsourceibias.n526 gnd 0.01085f
C4843 commonsourceibias.n527 gnd 0.058913f
C4844 commonsourceibias.n528 gnd 0.010777f
C4845 commonsourceibias.n529 gnd 0.007903f
C4846 commonsourceibias.n530 gnd 0.007903f
C4847 commonsourceibias.n531 gnd 0.007903f
C4848 commonsourceibias.n532 gnd 0.010777f
C4849 commonsourceibias.n533 gnd 0.058913f
C4850 commonsourceibias.n534 gnd 0.01085f
C4851 commonsourceibias.t117 gnd 0.147652f
C4852 commonsourceibias.n535 gnd 0.058913f
C4853 commonsourceibias.n536 gnd 0.009667f
C4854 commonsourceibias.n537 gnd 0.007903f
C4855 commonsourceibias.n538 gnd 0.007903f
C4856 commonsourceibias.n539 gnd 0.007903f
C4857 commonsourceibias.n540 gnd 0.009403f
C4858 commonsourceibias.n541 gnd 0.010904f
C4859 commonsourceibias.n542 gnd 0.058913f
C4860 commonsourceibias.n543 gnd 0.010838f
C4861 commonsourceibias.n544 gnd 0.007903f
C4862 commonsourceibias.n545 gnd 0.007903f
C4863 commonsourceibias.n546 gnd 0.007903f
C4864 commonsourceibias.n547 gnd 0.010705f
C4865 commonsourceibias.n548 gnd 0.058913f
C4866 commonsourceibias.n549 gnd 0.010776f
C4867 commonsourceibias.t73 gnd 0.147652f
C4868 commonsourceibias.n550 gnd 0.058913f
C4869 commonsourceibias.n551 gnd 0.009741f
C4870 commonsourceibias.n552 gnd 0.007903f
C4871 commonsourceibias.n553 gnd 0.007903f
C4872 commonsourceibias.n554 gnd 0.007903f
C4873 commonsourceibias.n555 gnd 0.008983f
C4874 commonsourceibias.n556 gnd 0.010937f
C4875 commonsourceibias.n557 gnd 0.058913f
C4876 commonsourceibias.n558 gnd 0.01089f
C4877 commonsourceibias.n559 gnd 0.007903f
C4878 commonsourceibias.n560 gnd 0.007903f
C4879 commonsourceibias.n561 gnd 0.007903f
C4880 commonsourceibias.n562 gnd 0.010623f
C4881 commonsourceibias.n563 gnd 0.058913f
C4882 commonsourceibias.n564 gnd 0.010649f
C4883 commonsourceibias.t99 gnd 0.159685f
C4884 commonsourceibias.n565 gnd 0.071041f
C4885 commonsourceibias.n566 gnd 0.02535f
C4886 commonsourceibias.n567 gnd 0.218509f
C4887 commonsourceibias.n568 gnd 4.2686f
C4888 a_n1986_8322.n0 gnd 1.477f
C4889 a_n1986_8322.n1 gnd 1.24631f
C4890 a_n1986_8322.n2 gnd 1.11016f
C4891 a_n1986_8322.n3 gnd 0.766493f
C4892 a_n1986_8322.n4 gnd 1.11016f
C4893 a_n1986_8322.t19 gnd 0.124841p
C4894 a_n1986_8322.t9 gnd 0.093529f
C4895 a_n1986_8322.t17 gnd 0.875761f
C4896 a_n1986_8322.t20 gnd 0.093529f
C4897 a_n1986_8322.t8 gnd 0.093529f
C4898 a_n1986_8322.n5 gnd 0.65882f
C4899 a_n1986_8322.t6 gnd 0.093529f
C4900 a_n1986_8322.t12 gnd 0.093529f
C4901 a_n1986_8322.n6 gnd 0.65882f
C4902 a_n1986_8322.t2 gnd 0.874017f
C4903 a_n1986_8322.n7 gnd 1.39891f
C4904 a_n1986_8322.t18 gnd 0.875761f
C4905 a_n1986_8322.t11 gnd 0.093529f
C4906 a_n1986_8322.t10 gnd 0.093529f
C4907 a_n1986_8322.n8 gnd 0.65882f
C4908 a_n1986_8322.t16 gnd 0.874017f
C4909 a_n1986_8322.t4 gnd 0.874017f
C4910 a_n1986_8322.t5 gnd 0.093529f
C4911 a_n1986_8322.t3 gnd 0.093529f
C4912 a_n1986_8322.n9 gnd 0.65882f
C4913 a_n1986_8322.t1 gnd 0.874017f
C4914 a_n1986_8322.n10 gnd 1.59065f
C4915 a_n1986_8322.n11 gnd 3.48702f
C4916 a_n1986_8322.t15 gnd 0.874017f
C4917 a_n1986_8322.t7 gnd 0.093529f
C4918 a_n1986_8322.t13 gnd 0.093529f
C4919 a_n1986_8322.n12 gnd 0.65882f
C4920 a_n1986_8322.t14 gnd 0.875759f
C4921 a_n1986_8322.n13 gnd 0.658822f
C4922 a_n1986_8322.t0 gnd 0.093529f
C4923 CSoutput.n0 gnd 0.040834f
C4924 CSoutput.t149 gnd 0.270108f
C4925 CSoutput.n1 gnd 0.121967f
C4926 CSoutput.n2 gnd 0.040834f
C4927 CSoutput.t154 gnd 0.270108f
C4928 CSoutput.n3 gnd 0.032364f
C4929 CSoutput.n4 gnd 0.040834f
C4930 CSoutput.t142 gnd 0.270108f
C4931 CSoutput.n5 gnd 0.027908f
C4932 CSoutput.n6 gnd 0.040834f
C4933 CSoutput.t152 gnd 0.270108f
C4934 CSoutput.t150 gnd 0.270108f
C4935 CSoutput.n7 gnd 0.120638f
C4936 CSoutput.n8 gnd 0.040834f
C4937 CSoutput.t141 gnd 0.270108f
C4938 CSoutput.n9 gnd 0.026609f
C4939 CSoutput.n10 gnd 0.040834f
C4940 CSoutput.t146 gnd 0.270108f
C4941 CSoutput.t148 gnd 0.270108f
C4942 CSoutput.n11 gnd 0.120638f
C4943 CSoutput.n12 gnd 0.040834f
C4944 CSoutput.t137 gnd 0.270108f
C4945 CSoutput.n13 gnd 0.027908f
C4946 CSoutput.n14 gnd 0.040834f
C4947 CSoutput.t157 gnd 0.270108f
C4948 CSoutput.t147 gnd 0.270108f
C4949 CSoutput.n15 gnd 0.120638f
C4950 CSoutput.n16 gnd 0.040834f
C4951 CSoutput.t151 gnd 0.270108f
C4952 CSoutput.n17 gnd 0.029807f
C4953 CSoutput.t138 gnd 0.322787f
C4954 CSoutput.t155 gnd 0.270108f
C4955 CSoutput.n18 gnd 0.154008f
C4956 CSoutput.n19 gnd 0.149441f
C4957 CSoutput.n20 gnd 0.17337f
C4958 CSoutput.n21 gnd 0.040834f
C4959 CSoutput.n22 gnd 0.034081f
C4960 CSoutput.n23 gnd 0.120638f
C4961 CSoutput.n24 gnd 0.032853f
C4962 CSoutput.n25 gnd 0.032364f
C4963 CSoutput.n26 gnd 0.040834f
C4964 CSoutput.n27 gnd 0.040834f
C4965 CSoutput.n28 gnd 0.033819f
C4966 CSoutput.n29 gnd 0.028713f
C4967 CSoutput.n30 gnd 0.123324f
C4968 CSoutput.n31 gnd 0.029108f
C4969 CSoutput.n32 gnd 0.040834f
C4970 CSoutput.n33 gnd 0.040834f
C4971 CSoutput.n34 gnd 0.040834f
C4972 CSoutput.n35 gnd 0.033458f
C4973 CSoutput.n36 gnd 0.120638f
C4974 CSoutput.n37 gnd 0.031998f
C4975 CSoutput.n38 gnd 0.033219f
C4976 CSoutput.n39 gnd 0.040834f
C4977 CSoutput.n40 gnd 0.040834f
C4978 CSoutput.n41 gnd 0.034074f
C4979 CSoutput.n42 gnd 0.031143f
C4980 CSoutput.n43 gnd 0.120638f
C4981 CSoutput.n44 gnd 0.031933f
C4982 CSoutput.n45 gnd 0.040834f
C4983 CSoutput.n46 gnd 0.040834f
C4984 CSoutput.n47 gnd 0.040834f
C4985 CSoutput.n48 gnd 0.031933f
C4986 CSoutput.n49 gnd 0.120638f
C4987 CSoutput.n50 gnd 0.031143f
C4988 CSoutput.n51 gnd 0.034074f
C4989 CSoutput.n52 gnd 0.040834f
C4990 CSoutput.n53 gnd 0.040834f
C4991 CSoutput.n54 gnd 0.033219f
C4992 CSoutput.n55 gnd 0.031998f
C4993 CSoutput.n56 gnd 0.120638f
C4994 CSoutput.n57 gnd 0.033458f
C4995 CSoutput.n58 gnd 0.040834f
C4996 CSoutput.n59 gnd 0.040834f
C4997 CSoutput.n60 gnd 0.040834f
C4998 CSoutput.n61 gnd 0.029108f
C4999 CSoutput.n62 gnd 0.123324f
C5000 CSoutput.n63 gnd 0.028713f
C5001 CSoutput.t153 gnd 0.270108f
C5002 CSoutput.n64 gnd 0.120638f
C5003 CSoutput.n65 gnd 0.033819f
C5004 CSoutput.n66 gnd 0.040834f
C5005 CSoutput.n67 gnd 0.040834f
C5006 CSoutput.n68 gnd 0.040834f
C5007 CSoutput.n69 gnd 0.032853f
C5008 CSoutput.n70 gnd 0.120638f
C5009 CSoutput.n71 gnd 0.034081f
C5010 CSoutput.n72 gnd 0.029807f
C5011 CSoutput.n73 gnd 0.040834f
C5012 CSoutput.n74 gnd 0.040834f
C5013 CSoutput.n75 gnd 0.030912f
C5014 CSoutput.n76 gnd 0.018359f
C5015 CSoutput.t140 gnd 0.303486f
C5016 CSoutput.n77 gnd 0.15076f
C5017 CSoutput.n78 gnd 0.645087f
C5018 CSoutput.t79 gnd 0.050935f
C5019 CSoutput.t13 gnd 0.050935f
C5020 CSoutput.n79 gnd 0.394354f
C5021 CSoutput.t22 gnd 0.050935f
C5022 CSoutput.t29 gnd 0.050935f
C5023 CSoutput.n80 gnd 0.393651f
C5024 CSoutput.n81 gnd 0.399555f
C5025 CSoutput.t102 gnd 0.050935f
C5026 CSoutput.t47 gnd 0.050935f
C5027 CSoutput.n82 gnd 0.393651f
C5028 CSoutput.n83 gnd 0.196884f
C5029 CSoutput.t81 gnd 0.050935f
C5030 CSoutput.t115 gnd 0.050935f
C5031 CSoutput.n84 gnd 0.393651f
C5032 CSoutput.n85 gnd 0.196884f
C5033 CSoutput.t33 gnd 0.050935f
C5034 CSoutput.t50 gnd 0.050935f
C5035 CSoutput.n86 gnd 0.393651f
C5036 CSoutput.n87 gnd 0.196884f
C5037 CSoutput.t61 gnd 0.050935f
C5038 CSoutput.t97 gnd 0.050935f
C5039 CSoutput.n88 gnd 0.393651f
C5040 CSoutput.n89 gnd 0.361039f
C5041 CSoutput.t87 gnd 0.050935f
C5042 CSoutput.t53 gnd 0.050935f
C5043 CSoutput.n90 gnd 0.394354f
C5044 CSoutput.t71 gnd 0.050935f
C5045 CSoutput.t35 gnd 0.050935f
C5046 CSoutput.n91 gnd 0.393651f
C5047 CSoutput.n92 gnd 0.399555f
C5048 CSoutput.t9 gnd 0.050935f
C5049 CSoutput.t103 gnd 0.050935f
C5050 CSoutput.n93 gnd 0.393651f
C5051 CSoutput.n94 gnd 0.196884f
C5052 CSoutput.t72 gnd 0.050935f
C5053 CSoutput.t74 gnd 0.050935f
C5054 CSoutput.n95 gnd 0.393651f
C5055 CSoutput.n96 gnd 0.196884f
C5056 CSoutput.t88 gnd 0.050935f
C5057 CSoutput.t105 gnd 0.050935f
C5058 CSoutput.n97 gnd 0.393651f
C5059 CSoutput.n98 gnd 0.196884f
C5060 CSoutput.t98 gnd 0.050935f
C5061 CSoutput.t99 gnd 0.050935f
C5062 CSoutput.n99 gnd 0.393651f
C5063 CSoutput.n100 gnd 0.293603f
C5064 CSoutput.n101 gnd 0.370232f
C5065 CSoutput.t126 gnd 0.050935f
C5066 CSoutput.t125 gnd 0.050935f
C5067 CSoutput.n102 gnd 0.394354f
C5068 CSoutput.t23 gnd 0.050935f
C5069 CSoutput.t48 gnd 0.050935f
C5070 CSoutput.n103 gnd 0.393651f
C5071 CSoutput.n104 gnd 0.399555f
C5072 CSoutput.t95 gnd 0.050935f
C5073 CSoutput.t104 gnd 0.050935f
C5074 CSoutput.n105 gnd 0.393651f
C5075 CSoutput.n106 gnd 0.196884f
C5076 CSoutput.t24 gnd 0.050935f
C5077 CSoutput.t134 gnd 0.050935f
C5078 CSoutput.n107 gnd 0.393651f
C5079 CSoutput.n108 gnd 0.196884f
C5080 CSoutput.t63 gnd 0.050935f
C5081 CSoutput.t85 gnd 0.050935f
C5082 CSoutput.n109 gnd 0.393651f
C5083 CSoutput.n110 gnd 0.196884f
C5084 CSoutput.t107 gnd 0.050935f
C5085 CSoutput.t108 gnd 0.050935f
C5086 CSoutput.n111 gnd 0.393651f
C5087 CSoutput.n112 gnd 0.293603f
C5088 CSoutput.n113 gnd 0.413824f
C5089 CSoutput.n114 gnd 7.535f
C5090 CSoutput.n116 gnd 0.722347f
C5091 CSoutput.n117 gnd 0.54176f
C5092 CSoutput.n118 gnd 0.722347f
C5093 CSoutput.n119 gnd 0.722347f
C5094 CSoutput.n120 gnd 1.94478f
C5095 CSoutput.n121 gnd 0.722347f
C5096 CSoutput.n122 gnd 0.722347f
C5097 CSoutput.t144 gnd 0.902934f
C5098 CSoutput.n123 gnd 0.722347f
C5099 CSoutput.n124 gnd 0.722347f
C5100 CSoutput.n128 gnd 0.722347f
C5101 CSoutput.n132 gnd 0.722347f
C5102 CSoutput.n133 gnd 0.722347f
C5103 CSoutput.n135 gnd 0.722347f
C5104 CSoutput.n140 gnd 0.722347f
C5105 CSoutput.n142 gnd 0.722347f
C5106 CSoutput.n143 gnd 0.722347f
C5107 CSoutput.n145 gnd 0.722347f
C5108 CSoutput.n146 gnd 0.722347f
C5109 CSoutput.n148 gnd 0.722347f
C5110 CSoutput.t139 gnd 12.0703f
C5111 CSoutput.n150 gnd 0.722347f
C5112 CSoutput.n151 gnd 0.54176f
C5113 CSoutput.n152 gnd 0.722347f
C5114 CSoutput.n153 gnd 0.722347f
C5115 CSoutput.n154 gnd 1.94478f
C5116 CSoutput.n155 gnd 0.722347f
C5117 CSoutput.n156 gnd 0.722347f
C5118 CSoutput.t156 gnd 0.902934f
C5119 CSoutput.n157 gnd 0.722347f
C5120 CSoutput.n158 gnd 0.722347f
C5121 CSoutput.n162 gnd 0.722347f
C5122 CSoutput.n166 gnd 0.722347f
C5123 CSoutput.n167 gnd 0.722347f
C5124 CSoutput.n169 gnd 0.722347f
C5125 CSoutput.n174 gnd 0.722347f
C5126 CSoutput.n176 gnd 0.722347f
C5127 CSoutput.n177 gnd 0.722347f
C5128 CSoutput.n179 gnd 0.722347f
C5129 CSoutput.n180 gnd 0.722347f
C5130 CSoutput.n182 gnd 0.722347f
C5131 CSoutput.n183 gnd 0.54176f
C5132 CSoutput.n185 gnd 0.722347f
C5133 CSoutput.n186 gnd 0.54176f
C5134 CSoutput.n187 gnd 0.722347f
C5135 CSoutput.n188 gnd 0.722347f
C5136 CSoutput.n189 gnd 1.94478f
C5137 CSoutput.n190 gnd 0.722347f
C5138 CSoutput.n191 gnd 0.722347f
C5139 CSoutput.t136 gnd 0.902934f
C5140 CSoutput.n192 gnd 0.722347f
C5141 CSoutput.n193 gnd 1.94478f
C5142 CSoutput.n195 gnd 0.722347f
C5143 CSoutput.n196 gnd 0.722347f
C5144 CSoutput.n198 gnd 0.722347f
C5145 CSoutput.n199 gnd 0.722347f
C5146 CSoutput.t145 gnd 11.873599f
C5147 CSoutput.t143 gnd 12.0703f
C5148 CSoutput.n205 gnd 2.26611f
C5149 CSoutput.n206 gnd 9.23131f
C5150 CSoutput.n207 gnd 9.617579f
C5151 CSoutput.n212 gnd 2.45481f
C5152 CSoutput.n218 gnd 0.722347f
C5153 CSoutput.n220 gnd 0.722347f
C5154 CSoutput.n222 gnd 0.722347f
C5155 CSoutput.n224 gnd 0.722347f
C5156 CSoutput.n226 gnd 0.722347f
C5157 CSoutput.n232 gnd 0.722347f
C5158 CSoutput.n239 gnd 1.32523f
C5159 CSoutput.n240 gnd 1.32523f
C5160 CSoutput.n241 gnd 0.722347f
C5161 CSoutput.n242 gnd 0.722347f
C5162 CSoutput.n244 gnd 0.54176f
C5163 CSoutput.n245 gnd 0.463969f
C5164 CSoutput.n247 gnd 0.54176f
C5165 CSoutput.n248 gnd 0.463969f
C5166 CSoutput.n249 gnd 0.54176f
C5167 CSoutput.n251 gnd 0.722347f
C5168 CSoutput.n253 gnd 1.94478f
C5169 CSoutput.n254 gnd 2.26611f
C5170 CSoutput.n255 gnd 8.49043f
C5171 CSoutput.n257 gnd 0.54176f
C5172 CSoutput.n258 gnd 1.39398f
C5173 CSoutput.n259 gnd 0.54176f
C5174 CSoutput.n261 gnd 0.722347f
C5175 CSoutput.n263 gnd 1.94478f
C5176 CSoutput.n264 gnd 4.23605f
C5177 CSoutput.t12 gnd 0.050935f
C5178 CSoutput.t86 gnd 0.050935f
C5179 CSoutput.n265 gnd 0.394354f
C5180 CSoutput.t70 gnd 0.050935f
C5181 CSoutput.t82 gnd 0.050935f
C5182 CSoutput.n266 gnd 0.393651f
C5183 CSoutput.n267 gnd 0.399555f
C5184 CSoutput.t89 gnd 0.050935f
C5185 CSoutput.t109 gnd 0.050935f
C5186 CSoutput.n268 gnd 0.393651f
C5187 CSoutput.n269 gnd 0.196884f
C5188 CSoutput.t76 gnd 0.050935f
C5189 CSoutput.t80 gnd 0.050935f
C5190 CSoutput.n270 gnd 0.393651f
C5191 CSoutput.n271 gnd 0.196884f
C5192 CSoutput.t21 gnd 0.050935f
C5193 CSoutput.t32 gnd 0.050935f
C5194 CSoutput.n272 gnd 0.393651f
C5195 CSoutput.n273 gnd 0.196884f
C5196 CSoutput.t96 gnd 0.050935f
C5197 CSoutput.t34 gnd 0.050935f
C5198 CSoutput.n274 gnd 0.393651f
C5199 CSoutput.n275 gnd 0.361039f
C5200 CSoutput.t69 gnd 0.050935f
C5201 CSoutput.t135 gnd 0.050935f
C5202 CSoutput.n276 gnd 0.394354f
C5203 CSoutput.t100 gnd 0.050935f
C5204 CSoutput.t8 gnd 0.050935f
C5205 CSoutput.n277 gnd 0.393651f
C5206 CSoutput.n278 gnd 0.399555f
C5207 CSoutput.t30 gnd 0.050935f
C5208 CSoutput.t101 gnd 0.050935f
C5209 CSoutput.n279 gnd 0.393651f
C5210 CSoutput.n280 gnd 0.196884f
C5211 CSoutput.t84 gnd 0.050935f
C5212 CSoutput.t133 gnd 0.050935f
C5213 CSoutput.n281 gnd 0.393651f
C5214 CSoutput.n282 gnd 0.196884f
C5215 CSoutput.t132 gnd 0.050935f
C5216 CSoutput.t78 gnd 0.050935f
C5217 CSoutput.n283 gnd 0.393651f
C5218 CSoutput.n284 gnd 0.196884f
C5219 CSoutput.t11 gnd 0.050935f
C5220 CSoutput.t10 gnd 0.050935f
C5221 CSoutput.n285 gnd 0.393651f
C5222 CSoutput.n286 gnd 0.293603f
C5223 CSoutput.n287 gnd 0.370232f
C5224 CSoutput.t37 gnd 0.050935f
C5225 CSoutput.t36 gnd 0.050935f
C5226 CSoutput.n288 gnd 0.394354f
C5227 CSoutput.t52 gnd 0.050935f
C5228 CSoutput.t94 gnd 0.050935f
C5229 CSoutput.n289 gnd 0.393651f
C5230 CSoutput.n290 gnd 0.399555f
C5231 CSoutput.t49 gnd 0.050935f
C5232 CSoutput.t110 gnd 0.050935f
C5233 CSoutput.n291 gnd 0.393651f
C5234 CSoutput.n292 gnd 0.196884f
C5235 CSoutput.t60 gnd 0.050935f
C5236 CSoutput.t75 gnd 0.050935f
C5237 CSoutput.n293 gnd 0.393651f
C5238 CSoutput.n294 gnd 0.196884f
C5239 CSoutput.t73 gnd 0.050935f
C5240 CSoutput.t83 gnd 0.050935f
C5241 CSoutput.n295 gnd 0.393651f
C5242 CSoutput.n296 gnd 0.196884f
C5243 CSoutput.t62 gnd 0.050935f
C5244 CSoutput.t116 gnd 0.050935f
C5245 CSoutput.n297 gnd 0.393649f
C5246 CSoutput.n298 gnd 0.293605f
C5247 CSoutput.n299 gnd 0.413824f
C5248 CSoutput.n300 gnd 10.7889f
C5249 CSoutput.t46 gnd 0.044568f
C5250 CSoutput.t38 gnd 0.044568f
C5251 CSoutput.n301 gnd 0.395136f
C5252 CSoutput.t111 gnd 0.044568f
C5253 CSoutput.t92 gnd 0.044568f
C5254 CSoutput.n302 gnd 0.393818f
C5255 CSoutput.n303 gnd 0.366964f
C5256 CSoutput.t0 gnd 0.044568f
C5257 CSoutput.t64 gnd 0.044568f
C5258 CSoutput.n304 gnd 0.393818f
C5259 CSoutput.n305 gnd 0.180896f
C5260 CSoutput.t27 gnd 0.044568f
C5261 CSoutput.t77 gnd 0.044568f
C5262 CSoutput.n306 gnd 0.393818f
C5263 CSoutput.n307 gnd 0.180896f
C5264 CSoutput.t45 gnd 0.044568f
C5265 CSoutput.t118 gnd 0.044568f
C5266 CSoutput.n308 gnd 0.393818f
C5267 CSoutput.n309 gnd 0.180896f
C5268 CSoutput.t122 gnd 0.044568f
C5269 CSoutput.t124 gnd 0.044568f
C5270 CSoutput.n310 gnd 0.393818f
C5271 CSoutput.n311 gnd 0.180896f
C5272 CSoutput.t117 gnd 0.044568f
C5273 CSoutput.t6 gnd 0.044568f
C5274 CSoutput.n312 gnd 0.393818f
C5275 CSoutput.n313 gnd 0.180896f
C5276 CSoutput.t58 gnd 0.044568f
C5277 CSoutput.t127 gnd 0.044568f
C5278 CSoutput.n314 gnd 0.393818f
C5279 CSoutput.n315 gnd 0.333609f
C5280 CSoutput.t57 gnd 0.044568f
C5281 CSoutput.t56 gnd 0.044568f
C5282 CSoutput.n316 gnd 0.395136f
C5283 CSoutput.t106 gnd 0.044568f
C5284 CSoutput.t7 gnd 0.044568f
C5285 CSoutput.n317 gnd 0.393818f
C5286 CSoutput.n318 gnd 0.366964f
C5287 CSoutput.t40 gnd 0.044568f
C5288 CSoutput.t14 gnd 0.044568f
C5289 CSoutput.n319 gnd 0.393818f
C5290 CSoutput.n320 gnd 0.180896f
C5291 CSoutput.t55 gnd 0.044568f
C5292 CSoutput.t20 gnd 0.044568f
C5293 CSoutput.n321 gnd 0.393818f
C5294 CSoutput.n322 gnd 0.180896f
C5295 CSoutput.t31 gnd 0.044568f
C5296 CSoutput.t44 gnd 0.044568f
C5297 CSoutput.n323 gnd 0.393818f
C5298 CSoutput.n324 gnd 0.180896f
C5299 CSoutput.t120 gnd 0.044568f
C5300 CSoutput.t119 gnd 0.044568f
C5301 CSoutput.n325 gnd 0.393818f
C5302 CSoutput.n326 gnd 0.180896f
C5303 CSoutput.t112 gnd 0.044568f
C5304 CSoutput.t123 gnd 0.044568f
C5305 CSoutput.n327 gnd 0.393818f
C5306 CSoutput.n328 gnd 0.180896f
C5307 CSoutput.t65 gnd 0.044568f
C5308 CSoutput.t2 gnd 0.044568f
C5309 CSoutput.n329 gnd 0.393818f
C5310 CSoutput.n330 gnd 0.274639f
C5311 CSoutput.n331 gnd 0.5103f
C5312 CSoutput.n332 gnd 11.4489f
C5313 CSoutput.t42 gnd 0.044568f
C5314 CSoutput.t67 gnd 0.044568f
C5315 CSoutput.n333 gnd 0.395136f
C5316 CSoutput.t4 gnd 0.044568f
C5317 CSoutput.t114 gnd 0.044568f
C5318 CSoutput.n334 gnd 0.393818f
C5319 CSoutput.n335 gnd 0.366964f
C5320 CSoutput.t19 gnd 0.044568f
C5321 CSoutput.t54 gnd 0.044568f
C5322 CSoutput.n336 gnd 0.393818f
C5323 CSoutput.n337 gnd 0.180896f
C5324 CSoutput.t121 gnd 0.044568f
C5325 CSoutput.t1 gnd 0.044568f
C5326 CSoutput.n338 gnd 0.393818f
C5327 CSoutput.n339 gnd 0.180896f
C5328 CSoutput.t130 gnd 0.044568f
C5329 CSoutput.t16 gnd 0.044568f
C5330 CSoutput.n340 gnd 0.393818f
C5331 CSoutput.n341 gnd 0.180896f
C5332 CSoutput.t91 gnd 0.044568f
C5333 CSoutput.t128 gnd 0.044568f
C5334 CSoutput.n342 gnd 0.393818f
C5335 CSoutput.n343 gnd 0.180896f
C5336 CSoutput.t5 gnd 0.044568f
C5337 CSoutput.t113 gnd 0.044568f
C5338 CSoutput.n344 gnd 0.393818f
C5339 CSoutput.n345 gnd 0.180896f
C5340 CSoutput.t39 gnd 0.044568f
C5341 CSoutput.t129 gnd 0.044568f
C5342 CSoutput.n346 gnd 0.393818f
C5343 CSoutput.n347 gnd 0.333609f
C5344 CSoutput.t28 gnd 0.044568f
C5345 CSoutput.t51 gnd 0.044568f
C5346 CSoutput.n348 gnd 0.395136f
C5347 CSoutput.t66 gnd 0.044568f
C5348 CSoutput.t43 gnd 0.044568f
C5349 CSoutput.n349 gnd 0.393818f
C5350 CSoutput.n350 gnd 0.366964f
C5351 CSoutput.t68 gnd 0.044568f
C5352 CSoutput.t25 gnd 0.044568f
C5353 CSoutput.n351 gnd 0.393818f
C5354 CSoutput.n352 gnd 0.180896f
C5355 CSoutput.t131 gnd 0.044568f
C5356 CSoutput.t59 gnd 0.044568f
C5357 CSoutput.n353 gnd 0.393818f
C5358 CSoutput.n354 gnd 0.180896f
C5359 CSoutput.t26 gnd 0.044568f
C5360 CSoutput.t17 gnd 0.044568f
C5361 CSoutput.n355 gnd 0.393818f
C5362 CSoutput.n356 gnd 0.180896f
C5363 CSoutput.t18 gnd 0.044568f
C5364 CSoutput.t41 gnd 0.044568f
C5365 CSoutput.n357 gnd 0.393818f
C5366 CSoutput.n358 gnd 0.180896f
C5367 CSoutput.t93 gnd 0.044568f
C5368 CSoutput.t90 gnd 0.044568f
C5369 CSoutput.n359 gnd 0.393818f
C5370 CSoutput.n360 gnd 0.180896f
C5371 CSoutput.t15 gnd 0.044568f
C5372 CSoutput.t3 gnd 0.044568f
C5373 CSoutput.n361 gnd 0.393818f
C5374 CSoutput.n362 gnd 0.274639f
C5375 CSoutput.n363 gnd 0.5103f
C5376 CSoutput.n364 gnd 6.55902f
C5377 CSoutput.n365 gnd 13.2435f
.ends

