* NGSPICE file created from opamp496.ext - technology: sky130A

.subckt opamp496 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n7636_8799.t44 plus.t5 a_n2903_n3924.t44 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t143 commonsourceibias.t64 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t7 a_n2982_13878.t72 vdd.t211 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2804_13878.t31 a_n2982_13878.t59 a_n2982_13878.t60 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 gnd.t248 gnd.t246 gnd.t247 gnd.t199 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 CSoutput.t144 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X6 vdd.t155 a_n7636_8799.t48 CSoutput.t7 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X7 gnd.t261 commonsourceibias.t65 CSoutput.t142 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t245 gnd.t243 minus.t4 gnd.t244 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X9 CSoutput.t141 commonsourceibias.t66 gnd.t63 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 CSoutput.t140 commonsourceibias.t67 gnd.t250 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 a_n2903_n3924.t28 plus.t6 a_n7636_8799.t43 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X12 vdd.t91 vdd.t89 vdd.t90 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X13 a_n2903_n3924.t51 minus.t5 a_n2982_13878.t68 gnd.t337 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X14 a_n2982_8322.t37 a_n2982_13878.t73 a_n7636_8799.t6 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 vdd.t4 CSoutput.t145 output.t15 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X16 CSoutput.t34 a_n7636_8799.t49 vdd.t154 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 CSoutput.t139 commonsourceibias.t68 gnd.t271 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t120 commonsourceibias.t69 CSoutput.t138 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t137 commonsourceibias.t70 gnd.t267 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t13 commonsourceibias.t71 CSoutput.t136 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t135 commonsourceibias.t72 gnd.t96 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 vdd.t153 a_n7636_8799.t50 CSoutput.t33 vdd.t126 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X23 CSoutput.t134 commonsourceibias.t73 gnd.t74 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 gnd.t275 commonsourceibias.t74 CSoutput.t133 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X25 a_n2982_13878.t65 minus.t6 a_n2903_n3924.t48 gnd.t336 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X26 commonsourceibias.t63 commonsourceibias.t62 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 CSoutput.t132 commonsourceibias.t75 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n7636_8799.t10 a_n2982_13878.t74 a_n2982_8322.t36 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 a_n2982_13878.t1 minus.t7 a_n2903_n3924.t2 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X30 vdd.t152 a_n7636_8799.t51 CSoutput.t32 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 CSoutput.t146 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X32 a_n7636_8799.t5 a_n2982_13878.t75 a_n2982_8322.t35 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t131 commonsourceibias.t76 gnd.t310 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 gnd.t353 commonsourceibias.t77 CSoutput.t130 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t242 gnd.t240 gnd.t241 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 CSoutput.t129 commonsourceibias.t78 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t128 commonsourceibias.t79 gnd.t316 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 a_n2903_n3924.t21 minus.t8 a_n2982_13878.t14 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X39 gnd.t239 gnd.t237 gnd.t238 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X40 CSoutput.t127 commonsourceibias.t80 gnd.t122 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n2903_n3924.t16 diffpairibias.t16 gnd.t293 gnd.t292 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 gnd.t324 commonsourceibias.t81 CSoutput.t126 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 CSoutput.t125 commonsourceibias.t82 gnd.t318 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X44 gnd.t259 commonsourceibias.t60 commonsourceibias.t61 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 CSoutput.t124 commonsourceibias.t83 gnd.t62 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 output.t18 outputibias.t8 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X47 gnd.t263 commonsourceibias.t84 CSoutput.t123 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 a_n2903_n3924.t46 plus.t7 a_n7636_8799.t42 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X49 CSoutput.t122 commonsourceibias.t85 gnd.t264 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 vdd.t88 vdd.t86 vdd.t87 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X51 a_n2804_13878.t30 a_n2982_13878.t51 a_n2982_13878.t52 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X52 gnd.t325 commonsourceibias.t86 CSoutput.t121 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 vdd.t5 CSoutput.t147 output.t14 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X54 a_n7636_8799.t41 plus.t8 a_n2903_n3924.t35 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X55 CSoutput.t120 commonsourceibias.t87 gnd.t326 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n2982_13878.t44 a_n2982_13878.t43 a_n2804_13878.t29 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 gnd.t300 commonsourceibias.t88 CSoutput.t119 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 a_n7636_8799.t40 plus.t9 a_n2903_n3924.t24 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X59 CSoutput.t39 a_n7636_8799.t52 vdd.t151 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 gnd.t367 commonsourceibias.t58 commonsourceibias.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 vdd.t85 vdd.t83 vdd.t84 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 CSoutput.t118 commonsourceibias.t89 gnd.t322 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 gnd.t236 gnd.t233 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X64 vdd.t150 a_n7636_8799.t53 CSoutput.t38 vdd.t126 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X65 gnd.t232 gnd.t230 gnd.t231 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X66 CSoutput.t117 commonsourceibias.t90 gnd.t102 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 diffpairibias.t15 diffpairibias.t14 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X68 a_n2903_n3924.t43 plus.t10 a_n7636_8799.t39 gnd.t340 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X69 a_n2982_13878.t0 minus.t9 a_n2903_n3924.t1 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X70 a_n2982_13878.t36 a_n2982_13878.t35 a_n2804_13878.t28 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X71 CSoutput.t116 commonsourceibias.t91 gnd.t350 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X72 CSoutput.t115 commonsourceibias.t92 gnd.t255 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 gnd.t14 commonsourceibias.t93 CSoutput.t114 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 gnd.t296 commonsourceibias.t94 CSoutput.t113 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 a_n7636_8799.t9 a_n2982_13878.t76 a_n2982_8322.t34 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X76 CSoutput.t37 a_n7636_8799.t54 vdd.t149 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 gnd.t71 commonsourceibias.t95 CSoutput.t112 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t229 gnd.t227 plus.t2 gnd.t228 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X79 a_n2982_13878.t40 a_n2982_13878.t39 a_n2804_13878.t27 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X80 vdd.t148 a_n7636_8799.t55 CSoutput.t28 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 vdd.t147 a_n7636_8799.t56 CSoutput.t27 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 a_n7636_8799.t15 a_n2982_13878.t77 a_n2982_8322.t33 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X83 CSoutput.t111 commonsourceibias.t96 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 diffpairibias.t13 diffpairibias.t12 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 CSoutput.t26 a_n7636_8799.t57 vdd.t146 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 gnd.t87 commonsourceibias.t56 commonsourceibias.t57 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd.t121 commonsourceibias.t97 CSoutput.t110 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t109 commonsourceibias.t98 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n7636_8799.t13 a_n2982_13878.t78 a_n2982_8322.t32 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 gnd.t36 commonsourceibias.t99 CSoutput.t108 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 gnd.t226 gnd.t224 gnd.t225 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X92 CSoutput.t107 commonsourceibias.t100 gnd.t314 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput.t106 commonsourceibias.t101 gnd.t25 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n2982_8322.t31 a_n2982_13878.t79 a_n7636_8799.t14 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 gnd.t117 commonsourceibias.t102 CSoutput.t105 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 CSoutput.t22 a_n7636_8799.t58 vdd.t145 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X97 CSoutput.t148 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X98 gnd.t279 commonsourceibias.t54 commonsourceibias.t55 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t223 gnd.t221 gnd.t222 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X100 gnd.t220 gnd.t218 plus.t1 gnd.t219 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X101 output.t13 CSoutput.t149 vdd.t2 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X102 a_n2903_n3924.t33 plus.t11 a_n7636_8799.t38 gnd.t339 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X103 gnd.t76 commonsourceibias.t103 CSoutput.t104 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 a_n2903_n3924.t0 diffpairibias.t17 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X105 vdd.t144 a_n7636_8799.t59 CSoutput.t21 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 gnd.t217 gnd.t215 gnd.t216 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X107 a_n2982_13878.t46 a_n2982_13878.t45 a_n2804_13878.t26 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X108 gnd.t303 commonsourceibias.t104 CSoutput.t103 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 a_n7636_8799.t4 a_n2982_13878.t80 a_n2982_8322.t30 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X110 a_n2982_13878.t18 a_n2982_13878.t17 a_n2804_13878.t25 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X111 gnd.t214 gnd.t212 gnd.t213 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X112 CSoutput.t102 commonsourceibias.t105 gnd.t86 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 gnd.t75 commonsourceibias.t106 CSoutput.t101 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n2982_13878.t3 minus.t10 a_n2903_n3924.t4 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X115 output.t12 CSoutput.t150 vdd.t0 gnd.t125 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X116 vdd.t82 vdd.t80 vdd.t81 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 gnd.t358 commonsourceibias.t52 commonsourceibias.t53 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 gnd.t302 commonsourceibias.t107 CSoutput.t100 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 CSoutput.t20 a_n7636_8799.t60 vdd.t143 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 output.t19 outputibias.t9 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X122 a_n2903_n3924.t49 minus.t11 a_n2982_13878.t66 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X123 a_n2804_13878.t24 a_n2982_13878.t23 a_n2982_13878.t24 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X124 CSoutput.t151 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X125 vdd.t207 a_n2982_13878.t81 a_n2982_8322.t13 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 a_n2982_13878.t22 a_n2982_13878.t21 a_n2804_13878.t23 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 a_n2982_8322.t12 a_n2982_13878.t82 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 gnd.t99 commonsourceibias.t108 CSoutput.t99 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X129 a_n2903_n3924.t14 diffpairibias.t18 gnd.t287 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 output.t11 CSoutput.t152 vdd.t14 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X131 CSoutput.t16 a_n7636_8799.t61 vdd.t142 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X132 vdd.t9 CSoutput.t153 output.t10 gnd.t106 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X133 gnd.t357 commonsourceibias.t109 CSoutput.t98 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 gnd.t252 commonsourceibias.t50 commonsourceibias.t51 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 CSoutput.t97 commonsourceibias.t110 gnd.t88 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 gnd.t49 commonsourceibias.t111 CSoutput.t96 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 CSoutput.t95 commonsourceibias.t112 gnd.t366 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X138 CSoutput.t94 commonsourceibias.t113 gnd.t89 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n2903_n3924.t52 minus.t12 a_n2982_13878.t69 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X140 a_n2903_n3924.t22 minus.t13 a_n2982_13878.t63 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X141 CSoutput.t154 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X142 vdd.t203 a_n2982_13878.t83 a_n2804_13878.t6 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 a_n2982_13878.t8 minus.t14 a_n2903_n3924.t10 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X144 a_n2903_n3924.t45 plus.t12 a_n7636_8799.t37 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X145 a_n2903_n3924.t25 plus.t13 a_n7636_8799.t36 gnd.t338 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X146 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X147 a_n2982_13878.t2 minus.t15 a_n2903_n3924.t3 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X148 gnd.t211 gnd.t209 gnd.t210 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X149 a_n2804_13878.t22 a_n2982_13878.t55 a_n2982_13878.t56 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 a_n2982_8322.t29 a_n2982_13878.t84 a_n7636_8799.t18 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 gnd.t208 gnd.t206 plus.t0 gnd.t207 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X152 a_n7636_8799.t35 plus.t14 a_n2903_n3924.t29 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X153 a_n7636_8799.t34 plus.t15 a_n2903_n3924.t30 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X154 vdd.t71 vdd.t69 vdd.t70 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X155 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X156 a_n2982_8322.t11 a_n2982_13878.t85 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X157 a_n7636_8799.t16 a_n2982_13878.t86 a_n2982_8322.t28 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 CSoutput.t15 a_n7636_8799.t62 vdd.t141 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 diffpairibias.t11 diffpairibias.t10 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X160 vdd.t140 a_n7636_8799.t63 CSoutput.t14 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 a_n2982_13878.t64 minus.t16 a_n2903_n3924.t23 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X162 a_n2982_13878.t32 a_n2982_13878.t31 a_n2804_13878.t21 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 CSoutput.t93 commonsourceibias.t114 gnd.t48 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 a_n7636_8799.t11 a_n2982_13878.t87 a_n2982_8322.t27 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 commonsourceibias.t49 commonsourceibias.t48 gnd.t359 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 output.t9 CSoutput.t155 vdd.t8 gnd.t107 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X167 gnd.t343 commonsourceibias.t115 CSoutput.t92 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 a_n2804_13878.t20 a_n2982_13878.t61 a_n2982_13878.t62 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X169 a_n2903_n3924.t8 minus.t17 a_n2982_13878.t7 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X170 gnd.t205 gnd.t202 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X171 CSoutput.t91 commonsourceibias.t116 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 vdd.t64 vdd.t62 vdd.t63 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X173 output.t8 CSoutput.t156 vdd.t15 gnd.t108 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 CSoutput.t43 a_n7636_8799.t64 vdd.t138 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 gnd.t201 gnd.t198 gnd.t200 gnd.t199 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X176 CSoutput.t90 commonsourceibias.t117 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 gnd.t197 gnd.t195 gnd.t196 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X178 vdd.t196 a_n2982_13878.t88 a_n2982_8322.t10 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X179 a_n2804_13878.t19 a_n2982_13878.t57 a_n2982_13878.t58 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 outputibias.t7 outputibias.t6 gnd.t298 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X181 vdd.t137 a_n7636_8799.t65 CSoutput.t42 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 gnd.t7 commonsourceibias.t118 CSoutput.t89 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t266 commonsourceibias.t119 CSoutput.t88 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n2982_13878.t20 a_n2982_13878.t19 a_n2804_13878.t18 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 commonsourceibias.t47 commonsourceibias.t46 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 minus.t3 gnd.t192 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X187 gnd.t317 commonsourceibias.t120 CSoutput.t87 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X188 outputibias.t5 outputibias.t4 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X189 a_n2903_n3924.t39 plus.t16 a_n7636_8799.t33 gnd.t337 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X190 vdd.t136 a_n7636_8799.t66 CSoutput.t4 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 CSoutput.t86 commonsourceibias.t121 gnd.t249 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 a_n2903_n3924.t9 diffpairibias.t19 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 gnd.t191 gnd.t188 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X194 a_n2903_n3924.t13 diffpairibias.t20 gnd.t285 gnd.t284 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X195 commonsourceibias.t45 commonsourceibias.t44 gnd.t319 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 vdd.t135 a_n7636_8799.t67 CSoutput.t3 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 a_n7636_8799.t32 plus.t17 a_n2903_n3924.t27 gnd.t336 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X198 gnd.t187 gnd.t185 gnd.t186 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X199 gnd.t184 gnd.t182 gnd.t183 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X200 vdd.t61 vdd.t59 vdd.t60 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 vdd.t7 CSoutput.t157 output.t7 gnd.t126 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X202 CSoutput.t85 commonsourceibias.t122 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 CSoutput.t84 commonsourceibias.t123 gnd.t299 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 a_n2804_13878.t17 a_n2982_13878.t33 a_n2982_13878.t34 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 a_n2982_8322.t26 a_n2982_13878.t89 a_n7636_8799.t3 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 CSoutput.t2 a_n7636_8799.t68 vdd.t134 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 commonsourceibias.t43 commonsourceibias.t42 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 gnd.t356 commonsourceibias.t40 commonsourceibias.t41 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 vdd.t12 CSoutput.t158 output.t6 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X210 diffpairibias.t9 diffpairibias.t8 gnd.t345 gnd.t344 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X211 a_n2804_13878.t5 a_n2982_13878.t90 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 vdd.t190 a_n2982_13878.t91 a_n2804_13878.t4 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X213 CSoutput.t83 commonsourceibias.t124 gnd.t118 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t82 commonsourceibias.t125 gnd.t64 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 vdd.t58 vdd.t56 vdd.t57 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X216 CSoutput.t11 a_n7636_8799.t69 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t274 commonsourceibias.t38 commonsourceibias.t39 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t131 a_n7636_8799.t70 CSoutput.t10 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t55 vdd.t53 vdd.t54 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X220 commonsourceibias.t37 commonsourceibias.t36 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 outputibias.t3 outputibias.t2 gnd.t273 gnd.t272 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X222 plus.t4 gnd.t179 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X223 a_n2804_13878.t16 a_n2982_13878.t53 a_n2982_13878.t54 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 a_n2903_n3924.t11 minus.t18 a_n2982_13878.t9 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X225 gnd.t294 commonsourceibias.t126 CSoutput.t81 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 commonsourceibias.t35 commonsourceibias.t34 gnd.t277 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X227 vdd.t129 a_n7636_8799.t71 CSoutput.t47 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 a_n2982_13878.t11 minus.t19 a_n2903_n3924.t18 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X229 gnd.t268 commonsourceibias.t32 commonsourceibias.t33 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 a_n2982_8322.t25 a_n2982_13878.t92 a_n7636_8799.t7 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X231 CSoutput.t80 commonsourceibias.t127 gnd.t251 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 CSoutput.t46 a_n7636_8799.t72 vdd.t128 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X233 a_n2982_13878.t30 a_n2982_13878.t29 a_n2804_13878.t15 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X234 diffpairibias.t7 diffpairibias.t6 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X235 vdd.t127 a_n7636_8799.t73 CSoutput.t36 vdd.t126 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X236 commonsourceibias.t31 commonsourceibias.t30 gnd.t348 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 a_n2982_13878.t10 minus.t20 a_n2903_n3924.t17 gnd.t304 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X238 a_n2804_13878.t14 a_n2982_13878.t49 a_n2982_13878.t50 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X239 a_n2982_13878.t6 minus.t21 a_n2903_n3924.t7 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X240 vdd.t185 a_n2982_13878.t93 a_n2982_8322.t9 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X241 vdd.t125 a_n7636_8799.t74 CSoutput.t35 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 a_n2903_n3924.t53 minus.t22 a_n2982_13878.t70 gnd.t340 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X243 a_n7636_8799.t31 plus.t18 a_n2903_n3924.t34 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X244 gnd.t66 commonsourceibias.t128 CSoutput.t79 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 a_n2903_n3924.t20 minus.t23 a_n2982_13878.t13 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X246 gnd.t315 commonsourceibias.t28 commonsourceibias.t29 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 CSoutput.t78 commonsourceibias.t129 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X248 a_n2804_13878.t3 a_n2982_13878.t94 vdd.t183 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X249 output.t5 CSoutput.t159 vdd.t3 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X250 gnd.t178 gnd.t176 minus.t2 gnd.t177 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X251 gnd.t5 commonsourceibias.t130 CSoutput.t77 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 vdd.t52 vdd.t49 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X253 gnd.t175 gnd.t172 gnd.t174 gnd.t173 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 vdd.t48 vdd.t46 vdd.t47 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X255 a_n2903_n3924.t12 diffpairibias.t21 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X256 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X257 vdd.t181 a_n2982_13878.t95 a_n2982_8322.t8 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X258 a_n2982_8322.t24 a_n2982_13878.t96 a_n7636_8799.t0 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 gnd.t73 commonsourceibias.t26 commonsourceibias.t27 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 a_n7636_8799.t30 plus.t19 a_n2903_n3924.t37 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X261 output.t16 outputibias.t10 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X262 gnd.t171 gnd.t169 gnd.t170 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X263 gnd.t24 commonsourceibias.t24 commonsourceibias.t25 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t41 vdd.t38 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X265 gnd.t168 gnd.t166 gnd.t167 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X266 CSoutput.t76 commonsourceibias.t131 gnd.t327 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 a_n2903_n3924.t41 plus.t20 a_n7636_8799.t29 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X268 vdd.t123 a_n7636_8799.t75 CSoutput.t30 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X269 vdd.t10 CSoutput.t160 output.t4 gnd.t109 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X270 CSoutput.t29 a_n7636_8799.t76 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X271 CSoutput.t75 commonsourceibias.t132 gnd.t328 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 output.t17 outputibias.t11 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X273 a_n2804_13878.t13 a_n2982_13878.t41 a_n2982_13878.t42 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X274 CSoutput.t25 a_n7636_8799.t77 vdd.t120 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X275 a_n2982_8322.t23 a_n2982_13878.t97 a_n7636_8799.t45 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 diffpairibias.t5 diffpairibias.t4 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X277 gnd.t165 gnd.t162 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X278 CSoutput.t24 a_n7636_8799.t78 vdd.t119 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 gnd.t57 commonsourceibias.t22 commonsourceibias.t23 gnd.t56 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X280 output.t3 CSoutput.t161 vdd.t6 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X281 vdd.t37 vdd.t34 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X282 CSoutput.t74 commonsourceibias.t133 gnd.t329 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 a_n2982_8322.t7 a_n2982_13878.t98 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X284 gnd.t330 commonsourceibias.t134 CSoutput.t73 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 vdd.t177 a_n2982_13878.t99 a_n2804_13878.t2 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X286 plus.t3 gnd.t159 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X287 CSoutput.t23 a_n7636_8799.t79 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 a_n2903_n3924.t26 plus.t21 a_n7636_8799.t28 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X289 gnd.t331 commonsourceibias.t135 CSoutput.t72 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t349 commonsourceibias.t136 CSoutput.t71 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 output.t2 CSoutput.t162 vdd.t13 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X292 a_n2903_n3924.t19 minus.t24 a_n2982_13878.t12 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X293 a_n2982_8322.t22 a_n2982_13878.t100 a_n7636_8799.t17 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X294 commonsourceibias.t21 commonsourceibias.t20 gnd.t352 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 vdd.t1 CSoutput.t163 output.t1 gnd.t112 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X296 a_n7636_8799.t12 a_n2982_13878.t101 a_n2982_8322.t21 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X297 a_n7636_8799.t27 plus.t22 a_n2903_n3924.t47 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X298 a_n2804_13878.t1 a_n2982_13878.t102 vdd.t167 vdd.t166 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X299 gnd.t333 commonsourceibias.t137 CSoutput.t70 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 vdd.t33 vdd.t31 vdd.t32 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X301 vdd.t116 a_n7636_8799.t80 CSoutput.t45 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 a_n2982_13878.t5 minus.t25 a_n2903_n3924.t6 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X303 CSoutput.t44 a_n7636_8799.t81 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X304 commonsourceibias.t19 commonsourceibias.t18 gnd.t332 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 a_n2982_13878.t38 a_n2982_13878.t37 a_n2804_13878.t12 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X306 a_n7636_8799.t1 a_n2982_13878.t103 a_n2982_8322.t20 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X307 gnd.t158 gnd.t155 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X308 a_n7636_8799.t2 a_n2982_13878.t104 a_n2982_8322.t19 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X309 gnd.t101 commonsourceibias.t138 CSoutput.t69 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 commonsourceibias.t17 commonsourceibias.t16 gnd.t301 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 a_n7636_8799.t26 plus.t23 a_n2903_n3924.t32 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X312 gnd.t154 gnd.t151 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X313 gnd.t150 gnd.t148 minus.t1 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X314 a_n2982_8322.t18 a_n2982_13878.t105 a_n7636_8799.t19 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X315 gnd.t119 commonsourceibias.t139 CSoutput.t68 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 CSoutput.t67 commonsourceibias.t140 gnd.t309 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X317 a_n2903_n3924.t50 minus.t26 a_n2982_13878.t67 gnd.t339 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X318 vdd.t113 a_n7636_8799.t82 CSoutput.t6 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t312 commonsourceibias.t14 commonsourceibias.t15 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 CSoutput.t5 a_n7636_8799.t83 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 CSoutput.t9 a_n7636_8799.t84 vdd.t109 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t8 a_n7636_8799.t85 vdd.t108 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 gnd.t147 gnd.t144 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X324 a_n2804_13878.t11 a_n2982_13878.t25 a_n2982_13878.t26 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X325 a_n2903_n3924.t38 plus.t24 a_n7636_8799.t25 gnd.t82 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X326 vdd.t107 a_n7636_8799.t86 CSoutput.t19 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 gnd.t256 commonsourceibias.t12 commonsourceibias.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X328 commonsourceibias.t11 commonsourceibias.t10 gnd.t276 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 gnd.t83 commonsourceibias.t141 CSoutput.t66 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n2903_n3924.t55 diffpairibias.t22 gnd.t361 gnd.t360 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X331 gnd.t351 commonsourceibias.t142 CSoutput.t65 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 CSoutput.t64 commonsourceibias.t143 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 vdd.t106 a_n7636_8799.t87 CSoutput.t18 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X334 gnd.t346 commonsourceibias.t144 CSoutput.t63 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 CSoutput.t17 a_n7636_8799.t88 vdd.t105 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 CSoutput.t62 commonsourceibias.t145 gnd.t100 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 a_n2982_13878.t48 a_n2982_13878.t47 a_n2804_13878.t10 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X338 gnd.t143 gnd.t140 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X339 a_n7636_8799.t46 a_n2982_13878.t106 a_n2982_8322.t17 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X340 vdd.t11 CSoutput.t164 output.t0 gnd.t113 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X341 vdd.t104 a_n7636_8799.t89 CSoutput.t41 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t40 a_n7636_8799.t90 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 a_n7636_8799.t24 plus.t25 a_n2903_n3924.t31 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X344 vdd.t30 vdd.t28 vdd.t29 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 CSoutput.t61 commonsourceibias.t146 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 gnd.t295 commonsourceibias.t147 CSoutput.t60 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X347 commonsourceibias.t9 commonsourceibias.t8 gnd.t45 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 diffpairibias.t3 diffpairibias.t2 gnd.t365 gnd.t364 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X349 CSoutput.t165 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X350 a_n2982_8322.t16 a_n2982_13878.t107 a_n7636_8799.t47 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X351 gnd.t98 commonsourceibias.t148 CSoutput.t59 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 a_n2903_n3924.t40 plus.t26 a_n7636_8799.t23 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X353 vdd.t101 a_n7636_8799.t91 CSoutput.t1 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 gnd.t139 gnd.t136 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X355 diffpairibias.t1 diffpairibias.t0 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X356 gnd.t42 commonsourceibias.t149 CSoutput.t58 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 commonsourceibias.t7 commonsourceibias.t6 gnd.t257 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 gnd.t61 commonsourceibias.t150 CSoutput.t57 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 a_n2903_n3924.t36 plus.t27 a_n7636_8799.t22 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X360 CSoutput.t56 commonsourceibias.t151 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X361 vdd.t163 a_n2982_13878.t108 a_n2804_13878.t0 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X362 a_n7636_8799.t21 plus.t28 a_n2903_n3924.t42 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X363 CSoutput.t0 a_n7636_8799.t92 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 a_n2903_n3924.t54 minus.t27 a_n2982_13878.t71 gnd.t338 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X365 vdd.t97 a_n7636_8799.t93 CSoutput.t13 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 gnd.t308 commonsourceibias.t4 commonsourceibias.t5 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 gnd.t311 commonsourceibias.t152 CSoutput.t55 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 a_n2982_8322.t15 a_n2982_13878.t109 a_n7636_8799.t20 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X369 a_n2982_13878.t4 minus.t28 a_n2903_n3924.t5 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X370 commonsourceibias.t3 commonsourceibias.t2 gnd.t265 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 gnd.t123 commonsourceibias.t153 CSoutput.t54 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 gnd.t135 gnd.t132 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X373 gnd.t347 commonsourceibias.t154 CSoutput.t53 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 a_n2982_8322.t14 a_n2982_13878.t110 a_n7636_8799.t8 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X375 vdd.t95 a_n7636_8799.t94 CSoutput.t12 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t31 a_n7636_8799.t95 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 gnd.t59 commonsourceibias.t155 CSoutput.t52 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 vdd.t27 vdd.t24 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X379 a_n2982_8322.t6 a_n2982_13878.t111 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X380 gnd.t342 commonsourceibias.t156 CSoutput.t51 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X381 a_n2804_13878.t9 a_n2982_13878.t15 a_n2982_13878.t16 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X382 gnd.t341 commonsourceibias.t157 CSoutput.t50 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 CSoutput.t49 commonsourceibias.t158 gnd.t323 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 commonsourceibias.t1 commonsourceibias.t0 gnd.t278 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X385 CSoutput.t48 commonsourceibias.t159 gnd.t97 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 minus.t0 gnd.t129 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X387 outputibias.t1 outputibias.t0 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X388 vdd.t23 vdd.t20 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X389 a_n2903_n3924.t15 diffpairibias.t23 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X390 vdd.t19 vdd.t16 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X391 a_n2982_13878.t28 a_n2982_13878.t27 a_n2804_13878.t8 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t0 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t1 19.8005
R93 plus.n85 plus.t4 19.8005
R94 plus.n87 plus.t2 19.8005
R95 plus.n87 plus.t3 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 14.5734
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n2903_n3924.n11 a_n2903_n3924.t12 214.643
R160 a_n2903_n3924.n7 a_n2903_n3924.t14 214.321
R161 a_n2903_n3924.n7 a_n2903_n3924.t55 214.321
R162 a_n2903_n3924.n5 a_n2903_n3924.t13 214.321
R163 a_n2903_n3924.n5 a_n2903_n3924.t15 214.321
R164 a_n2903_n3924.n6 a_n2903_n3924.t9 214.321
R165 a_n2903_n3924.n6 a_n2903_n3924.t16 214.321
R166 a_n2903_n3924.n11 a_n2903_n3924.t0 214.321
R167 a_n2903_n3924.n1 a_n2903_n3924.t41 55.8337
R168 a_n2903_n3924.n1 a_n2903_n3924.t5 55.8337
R169 a_n2903_n3924.n10 a_n2903_n3924.t22 55.8337
R170 a_n2903_n3924.n0 a_n2903_n3924.t35 55.8335
R171 a_n2903_n3924.n8 a_n2903_n3924.t18 55.8335
R172 a_n2903_n3924.n4 a_n2903_n3924.t21 55.8335
R173 a_n2903_n3924.n4 a_n2903_n3924.t30 55.8335
R174 a_n2903_n3924.n3 a_n2903_n3924.t26 55.8335
R175 a_n2903_n3924.n0 a_n2903_n3924.n28 53.0052
R176 a_n2903_n3924.n0 a_n2903_n3924.n29 53.0052
R177 a_n2903_n3924.n0 a_n2903_n3924.n30 53.0052
R178 a_n2903_n3924.n1 a_n2903_n3924.n31 53.0052
R179 a_n2903_n3924.n1 a_n2903_n3924.n32 53.0052
R180 a_n2903_n3924.n1 a_n2903_n3924.n12 53.0052
R181 a_n2903_n3924.n9 a_n2903_n3924.n13 53.0052
R182 a_n2903_n3924.n9 a_n2903_n3924.n14 53.0052
R183 a_n2903_n3924.n10 a_n2903_n3924.n15 53.0052
R184 a_n2903_n3924.n8 a_n2903_n3924.n26 53.0051
R185 a_n2903_n3924.n2 a_n2903_n3924.n25 53.0051
R186 a_n2903_n3924.n2 a_n2903_n3924.n24 53.0051
R187 a_n2903_n3924.n2 a_n2903_n3924.n23 53.0051
R188 a_n2903_n3924.n2 a_n2903_n3924.n22 53.0051
R189 a_n2903_n3924.n4 a_n2903_n3924.n21 53.0051
R190 a_n2903_n3924.n4 a_n2903_n3924.n20 53.0051
R191 a_n2903_n3924.n4 a_n2903_n3924.n19 53.0051
R192 a_n2903_n3924.n3 a_n2903_n3924.n18 53.0051
R193 a_n2903_n3924.n3 a_n2903_n3924.n17 53.0051
R194 a_n2903_n3924.n33 a_n2903_n3924.n1 53.0051
R195 a_n2903_n3924.n16 a_n2903_n3924.n10 12.1986
R196 a_n2903_n3924.n0 a_n2903_n3924.n27 12.1986
R197 a_n2903_n3924.n3 a_n2903_n3924.n16 5.11903
R198 a_n2903_n3924.n27 a_n2903_n3924.n8 5.11903
R199 a_n2903_n3924.n28 a_n2903_n3924.t42 2.82907
R200 a_n2903_n3924.n28 a_n2903_n3924.t43 2.82907
R201 a_n2903_n3924.n29 a_n2903_n3924.t29 2.82907
R202 a_n2903_n3924.n29 a_n2903_n3924.t45 2.82907
R203 a_n2903_n3924.n30 a_n2903_n3924.t24 2.82907
R204 a_n2903_n3924.n30 a_n2903_n3924.t46 2.82907
R205 a_n2903_n3924.n31 a_n2903_n3924.t31 2.82907
R206 a_n2903_n3924.n31 a_n2903_n3924.t36 2.82907
R207 a_n2903_n3924.n32 a_n2903_n3924.t37 2.82907
R208 a_n2903_n3924.n32 a_n2903_n3924.t40 2.82907
R209 a_n2903_n3924.n12 a_n2903_n3924.t23 2.82907
R210 a_n2903_n3924.n12 a_n2903_n3924.t8 2.82907
R211 a_n2903_n3924.n13 a_n2903_n3924.t7 2.82907
R212 a_n2903_n3924.n13 a_n2903_n3924.t20 2.82907
R213 a_n2903_n3924.n14 a_n2903_n3924.t48 2.82907
R214 a_n2903_n3924.n14 a_n2903_n3924.t50 2.82907
R215 a_n2903_n3924.n15 a_n2903_n3924.t3 2.82907
R216 a_n2903_n3924.n15 a_n2903_n3924.t51 2.82907
R217 a_n2903_n3924.n26 a_n2903_n3924.t10 2.82907
R218 a_n2903_n3924.n26 a_n2903_n3924.t53 2.82907
R219 a_n2903_n3924.n25 a_n2903_n3924.t6 2.82907
R220 a_n2903_n3924.n25 a_n2903_n3924.t19 2.82907
R221 a_n2903_n3924.n24 a_n2903_n3924.t17 2.82907
R222 a_n2903_n3924.n24 a_n2903_n3924.t11 2.82907
R223 a_n2903_n3924.n23 a_n2903_n3924.t4 2.82907
R224 a_n2903_n3924.n23 a_n2903_n3924.t52 2.82907
R225 a_n2903_n3924.n22 a_n2903_n3924.t2 2.82907
R226 a_n2903_n3924.n22 a_n2903_n3924.t49 2.82907
R227 a_n2903_n3924.n21 a_n2903_n3924.t34 2.82907
R228 a_n2903_n3924.n21 a_n2903_n3924.t25 2.82907
R229 a_n2903_n3924.n20 a_n2903_n3924.t32 2.82907
R230 a_n2903_n3924.n20 a_n2903_n3924.t38 2.82907
R231 a_n2903_n3924.n19 a_n2903_n3924.t44 2.82907
R232 a_n2903_n3924.n19 a_n2903_n3924.t28 2.82907
R233 a_n2903_n3924.n18 a_n2903_n3924.t27 2.82907
R234 a_n2903_n3924.n18 a_n2903_n3924.t33 2.82907
R235 a_n2903_n3924.n17 a_n2903_n3924.t47 2.82907
R236 a_n2903_n3924.n17 a_n2903_n3924.t39 2.82907
R237 a_n2903_n3924.t1 a_n2903_n3924.n33 2.82907
R238 a_n2903_n3924.n33 a_n2903_n3924.t54 2.82907
R239 a_n2903_n3924.n1 a_n2903_n3924.n0 2.66429
R240 a_n2903_n3924.n27 a_n2903_n3924.n7 2.16406
R241 a_n2903_n3924.n2 a_n2903_n3924.n4 2.01128
R242 a_n2903_n3924.n16 a_n2903_n3924.n11 1.95694
R243 a_n2903_n3924.n4 a_n2903_n3924.n3 1.77636
R244 a_n2903_n3924.n8 a_n2903_n3924.n2 1.77636
R245 a_n2903_n3924.n11 a_n2903_n3924.n6 1.69309
R246 a_n2903_n3924.n9 a_n2903_n3924.n1 1.56731
R247 a_n2903_n3924.n5 a_n2903_n3924.n7 1.34352
R248 a_n2903_n3924.n6 a_n2903_n3924.n5 1.34352
R249 a_n2903_n3924.n10 a_n2903_n3924.n9 1.3324
R250 a_n7636_8799.n99 a_n7636_8799.t58 485.149
R251 a_n7636_8799.n121 a_n7636_8799.t61 485.149
R252 a_n7636_8799.n144 a_n7636_8799.t76 485.149
R253 a_n7636_8799.n31 a_n7636_8799.t87 485.149
R254 a_n7636_8799.n53 a_n7636_8799.t94 485.149
R255 a_n7636_8799.n76 a_n7636_8799.t75 485.149
R256 a_n7636_8799.n114 a_n7636_8799.t50 464.166
R257 a_n7636_8799.n113 a_n7636_8799.t49 464.166
R258 a_n7636_8799.n95 a_n7636_8799.t80 464.166
R259 a_n7636_8799.n107 a_n7636_8799.t57 464.166
R260 a_n7636_8799.n106 a_n7636_8799.t51 464.166
R261 a_n7636_8799.n98 a_n7636_8799.t84 464.166
R262 a_n7636_8799.n100 a_n7636_8799.t67 464.166
R263 a_n7636_8799.n136 a_n7636_8799.t53 464.166
R264 a_n7636_8799.n135 a_n7636_8799.t52 464.166
R265 a_n7636_8799.n117 a_n7636_8799.t91 464.166
R266 a_n7636_8799.n129 a_n7636_8799.t60 464.166
R267 a_n7636_8799.n128 a_n7636_8799.t56 464.166
R268 a_n7636_8799.n120 a_n7636_8799.t92 464.166
R269 a_n7636_8799.n122 a_n7636_8799.t74 464.166
R270 a_n7636_8799.n159 a_n7636_8799.t73 464.166
R271 a_n7636_8799.n158 a_n7636_8799.t79 464.166
R272 a_n7636_8799.n140 a_n7636_8799.t55 464.166
R273 a_n7636_8799.n152 a_n7636_8799.t90 464.166
R274 a_n7636_8799.n151 a_n7636_8799.t63 464.166
R275 a_n7636_8799.n143 a_n7636_8799.t85 464.166
R276 a_n7636_8799.n145 a_n7636_8799.t59 464.166
R277 a_n7636_8799.n32 a_n7636_8799.t88 464.166
R278 a_n7636_8799.n34 a_n7636_8799.t66 464.166
R279 a_n7636_8799.n38 a_n7636_8799.t78 464.166
R280 a_n7636_8799.n39 a_n7636_8799.t86 464.166
R281 a_n7636_8799.n27 a_n7636_8799.t64 464.166
R282 a_n7636_8799.n45 a_n7636_8799.t65 464.166
R283 a_n7636_8799.n46 a_n7636_8799.t77 464.166
R284 a_n7636_8799.n54 a_n7636_8799.t95 464.166
R285 a_n7636_8799.n56 a_n7636_8799.t71 464.166
R286 a_n7636_8799.n60 a_n7636_8799.t83 464.166
R287 a_n7636_8799.n61 a_n7636_8799.t93 464.166
R288 a_n7636_8799.n49 a_n7636_8799.t69 464.166
R289 a_n7636_8799.n67 a_n7636_8799.t70 464.166
R290 a_n7636_8799.n68 a_n7636_8799.t81 464.166
R291 a_n7636_8799.n77 a_n7636_8799.t68 464.166
R292 a_n7636_8799.n79 a_n7636_8799.t82 464.166
R293 a_n7636_8799.n83 a_n7636_8799.t62 464.166
R294 a_n7636_8799.n84 a_n7636_8799.t89 464.166
R295 a_n7636_8799.n72 a_n7636_8799.t54 464.166
R296 a_n7636_8799.n90 a_n7636_8799.t48 464.166
R297 a_n7636_8799.n91 a_n7636_8799.t72 464.166
R298 a_n7636_8799.n102 a_n7636_8799.n101 161.3
R299 a_n7636_8799.n103 a_n7636_8799.n98 161.3
R300 a_n7636_8799.n105 a_n7636_8799.n104 161.3
R301 a_n7636_8799.n106 a_n7636_8799.n97 161.3
R302 a_n7636_8799.n107 a_n7636_8799.n96 161.3
R303 a_n7636_8799.n109 a_n7636_8799.n108 161.3
R304 a_n7636_8799.n110 a_n7636_8799.n95 161.3
R305 a_n7636_8799.n112 a_n7636_8799.n111 161.3
R306 a_n7636_8799.n113 a_n7636_8799.n94 161.3
R307 a_n7636_8799.n115 a_n7636_8799.n114 161.3
R308 a_n7636_8799.n124 a_n7636_8799.n123 161.3
R309 a_n7636_8799.n125 a_n7636_8799.n120 161.3
R310 a_n7636_8799.n127 a_n7636_8799.n126 161.3
R311 a_n7636_8799.n128 a_n7636_8799.n119 161.3
R312 a_n7636_8799.n129 a_n7636_8799.n118 161.3
R313 a_n7636_8799.n131 a_n7636_8799.n130 161.3
R314 a_n7636_8799.n132 a_n7636_8799.n117 161.3
R315 a_n7636_8799.n134 a_n7636_8799.n133 161.3
R316 a_n7636_8799.n135 a_n7636_8799.n116 161.3
R317 a_n7636_8799.n137 a_n7636_8799.n136 161.3
R318 a_n7636_8799.n147 a_n7636_8799.n146 161.3
R319 a_n7636_8799.n148 a_n7636_8799.n143 161.3
R320 a_n7636_8799.n150 a_n7636_8799.n149 161.3
R321 a_n7636_8799.n151 a_n7636_8799.n142 161.3
R322 a_n7636_8799.n152 a_n7636_8799.n141 161.3
R323 a_n7636_8799.n154 a_n7636_8799.n153 161.3
R324 a_n7636_8799.n155 a_n7636_8799.n140 161.3
R325 a_n7636_8799.n157 a_n7636_8799.n156 161.3
R326 a_n7636_8799.n158 a_n7636_8799.n139 161.3
R327 a_n7636_8799.n160 a_n7636_8799.n159 161.3
R328 a_n7636_8799.n47 a_n7636_8799.n46 161.3
R329 a_n7636_8799.n45 a_n7636_8799.n26 161.3
R330 a_n7636_8799.n44 a_n7636_8799.n43 161.3
R331 a_n7636_8799.n42 a_n7636_8799.n27 161.3
R332 a_n7636_8799.n41 a_n7636_8799.n40 161.3
R333 a_n7636_8799.n39 a_n7636_8799.n28 161.3
R334 a_n7636_8799.n38 a_n7636_8799.n37 161.3
R335 a_n7636_8799.n36 a_n7636_8799.n29 161.3
R336 a_n7636_8799.n35 a_n7636_8799.n34 161.3
R337 a_n7636_8799.n33 a_n7636_8799.n30 161.3
R338 a_n7636_8799.n69 a_n7636_8799.n68 161.3
R339 a_n7636_8799.n67 a_n7636_8799.n48 161.3
R340 a_n7636_8799.n66 a_n7636_8799.n65 161.3
R341 a_n7636_8799.n64 a_n7636_8799.n49 161.3
R342 a_n7636_8799.n63 a_n7636_8799.n62 161.3
R343 a_n7636_8799.n61 a_n7636_8799.n50 161.3
R344 a_n7636_8799.n60 a_n7636_8799.n59 161.3
R345 a_n7636_8799.n58 a_n7636_8799.n51 161.3
R346 a_n7636_8799.n57 a_n7636_8799.n56 161.3
R347 a_n7636_8799.n55 a_n7636_8799.n52 161.3
R348 a_n7636_8799.n92 a_n7636_8799.n91 161.3
R349 a_n7636_8799.n90 a_n7636_8799.n71 161.3
R350 a_n7636_8799.n89 a_n7636_8799.n88 161.3
R351 a_n7636_8799.n87 a_n7636_8799.n72 161.3
R352 a_n7636_8799.n86 a_n7636_8799.n85 161.3
R353 a_n7636_8799.n84 a_n7636_8799.n73 161.3
R354 a_n7636_8799.n83 a_n7636_8799.n82 161.3
R355 a_n7636_8799.n81 a_n7636_8799.n74 161.3
R356 a_n7636_8799.n80 a_n7636_8799.n79 161.3
R357 a_n7636_8799.n78 a_n7636_8799.n75 161.3
R358 a_n7636_8799.n16 a_n7636_8799.n14 98.9633
R359 a_n7636_8799.n5 a_n7636_8799.n3 98.9631
R360 a_n7636_8799.n24 a_n7636_8799.n23 98.6055
R361 a_n7636_8799.n22 a_n7636_8799.n21 98.6055
R362 a_n7636_8799.n20 a_n7636_8799.n19 98.6055
R363 a_n7636_8799.n18 a_n7636_8799.n17 98.6055
R364 a_n7636_8799.n16 a_n7636_8799.n15 98.6055
R365 a_n7636_8799.n5 a_n7636_8799.n4 98.6055
R366 a_n7636_8799.n7 a_n7636_8799.n6 98.6055
R367 a_n7636_8799.n9 a_n7636_8799.n8 98.6055
R368 a_n7636_8799.n11 a_n7636_8799.n10 98.6055
R369 a_n7636_8799.n13 a_n7636_8799.n12 98.6055
R370 a_n7636_8799.n166 a_n7636_8799.n164 81.3764
R371 a_n7636_8799.n178 a_n7636_8799.n176 81.3764
R372 a_n7636_8799.n2 a_n7636_8799.n0 81.3764
R373 a_n7636_8799.n183 a_n7636_8799.n182 80.9326
R374 a_n7636_8799.n175 a_n7636_8799.n174 80.9324
R375 a_n7636_8799.n173 a_n7636_8799.n172 80.9324
R376 a_n7636_8799.n171 a_n7636_8799.n170 80.9324
R377 a_n7636_8799.n168 a_n7636_8799.n167 80.9324
R378 a_n7636_8799.n166 a_n7636_8799.n165 80.9324
R379 a_n7636_8799.n178 a_n7636_8799.n177 80.9324
R380 a_n7636_8799.n180 a_n7636_8799.n179 80.9324
R381 a_n7636_8799.n2 a_n7636_8799.n1 80.9324
R382 a_n7636_8799.n102 a_n7636_8799.n99 70.4033
R383 a_n7636_8799.n124 a_n7636_8799.n121 70.4033
R384 a_n7636_8799.n147 a_n7636_8799.n144 70.4033
R385 a_n7636_8799.n31 a_n7636_8799.n30 70.4033
R386 a_n7636_8799.n53 a_n7636_8799.n52 70.4033
R387 a_n7636_8799.n76 a_n7636_8799.n75 70.4033
R388 a_n7636_8799.n114 a_n7636_8799.n113 48.2005
R389 a_n7636_8799.n107 a_n7636_8799.n106 48.2005
R390 a_n7636_8799.n136 a_n7636_8799.n135 48.2005
R391 a_n7636_8799.n129 a_n7636_8799.n128 48.2005
R392 a_n7636_8799.n159 a_n7636_8799.n158 48.2005
R393 a_n7636_8799.n152 a_n7636_8799.n151 48.2005
R394 a_n7636_8799.n39 a_n7636_8799.n38 48.2005
R395 a_n7636_8799.n46 a_n7636_8799.n45 48.2005
R396 a_n7636_8799.n61 a_n7636_8799.n60 48.2005
R397 a_n7636_8799.n68 a_n7636_8799.n67 48.2005
R398 a_n7636_8799.n84 a_n7636_8799.n83 48.2005
R399 a_n7636_8799.n91 a_n7636_8799.n90 48.2005
R400 a_n7636_8799.n112 a_n7636_8799.n95 37.246
R401 a_n7636_8799.n101 a_n7636_8799.n98 37.246
R402 a_n7636_8799.n134 a_n7636_8799.n117 37.246
R403 a_n7636_8799.n123 a_n7636_8799.n120 37.246
R404 a_n7636_8799.n157 a_n7636_8799.n140 37.246
R405 a_n7636_8799.n146 a_n7636_8799.n143 37.246
R406 a_n7636_8799.n34 a_n7636_8799.n33 37.246
R407 a_n7636_8799.n44 a_n7636_8799.n27 37.246
R408 a_n7636_8799.n56 a_n7636_8799.n55 37.246
R409 a_n7636_8799.n66 a_n7636_8799.n49 37.246
R410 a_n7636_8799.n79 a_n7636_8799.n78 37.246
R411 a_n7636_8799.n89 a_n7636_8799.n72 37.246
R412 a_n7636_8799.n108 a_n7636_8799.n95 35.7853
R413 a_n7636_8799.n105 a_n7636_8799.n98 35.7853
R414 a_n7636_8799.n130 a_n7636_8799.n117 35.7853
R415 a_n7636_8799.n127 a_n7636_8799.n120 35.7853
R416 a_n7636_8799.n153 a_n7636_8799.n140 35.7853
R417 a_n7636_8799.n150 a_n7636_8799.n143 35.7853
R418 a_n7636_8799.n34 a_n7636_8799.n29 35.7853
R419 a_n7636_8799.n40 a_n7636_8799.n27 35.7853
R420 a_n7636_8799.n56 a_n7636_8799.n51 35.7853
R421 a_n7636_8799.n62 a_n7636_8799.n49 35.7853
R422 a_n7636_8799.n79 a_n7636_8799.n74 35.7853
R423 a_n7636_8799.n85 a_n7636_8799.n72 35.7853
R424 a_n7636_8799.n25 a_n7636_8799.n13 34.1553
R425 a_n7636_8799.n181 a_n7636_8799.n175 33.4185
R426 a_n7636_8799.n100 a_n7636_8799.n99 20.9576
R427 a_n7636_8799.n122 a_n7636_8799.n121 20.9576
R428 a_n7636_8799.n145 a_n7636_8799.n144 20.9576
R429 a_n7636_8799.n32 a_n7636_8799.n31 20.9576
R430 a_n7636_8799.n54 a_n7636_8799.n53 20.9576
R431 a_n7636_8799.n77 a_n7636_8799.n76 20.9576
R432 a_n7636_8799.n25 a_n7636_8799.n24 20.7339
R433 a_n7636_8799.n108 a_n7636_8799.n107 12.4157
R434 a_n7636_8799.n106 a_n7636_8799.n105 12.4157
R435 a_n7636_8799.n130 a_n7636_8799.n129 12.4157
R436 a_n7636_8799.n128 a_n7636_8799.n127 12.4157
R437 a_n7636_8799.n153 a_n7636_8799.n152 12.4157
R438 a_n7636_8799.n151 a_n7636_8799.n150 12.4157
R439 a_n7636_8799.n38 a_n7636_8799.n29 12.4157
R440 a_n7636_8799.n40 a_n7636_8799.n39 12.4157
R441 a_n7636_8799.n60 a_n7636_8799.n51 12.4157
R442 a_n7636_8799.n62 a_n7636_8799.n61 12.4157
R443 a_n7636_8799.n83 a_n7636_8799.n74 12.4157
R444 a_n7636_8799.n85 a_n7636_8799.n84 12.4157
R445 a_n7636_8799.n169 a_n7636_8799.n163 12.3339
R446 a_n7636_8799.n163 a_n7636_8799.n25 11.4887
R447 a_n7636_8799.n113 a_n7636_8799.n112 10.955
R448 a_n7636_8799.n101 a_n7636_8799.n100 10.955
R449 a_n7636_8799.n135 a_n7636_8799.n134 10.955
R450 a_n7636_8799.n123 a_n7636_8799.n122 10.955
R451 a_n7636_8799.n158 a_n7636_8799.n157 10.955
R452 a_n7636_8799.n146 a_n7636_8799.n145 10.955
R453 a_n7636_8799.n33 a_n7636_8799.n32 10.955
R454 a_n7636_8799.n45 a_n7636_8799.n44 10.955
R455 a_n7636_8799.n55 a_n7636_8799.n54 10.955
R456 a_n7636_8799.n67 a_n7636_8799.n66 10.955
R457 a_n7636_8799.n78 a_n7636_8799.n77 10.955
R458 a_n7636_8799.n90 a_n7636_8799.n89 10.955
R459 a_n7636_8799.n138 a_n7636_8799.n115 9.05164
R460 a_n7636_8799.n70 a_n7636_8799.n47 9.05164
R461 a_n7636_8799.n162 a_n7636_8799.n93 7.2142
R462 a_n7636_8799.n162 a_n7636_8799.n161 6.79277
R463 a_n7636_8799.n138 a_n7636_8799.n137 4.94368
R464 a_n7636_8799.n161 a_n7636_8799.n160 4.94368
R465 a_n7636_8799.n70 a_n7636_8799.n69 4.94368
R466 a_n7636_8799.n93 a_n7636_8799.n92 4.94368
R467 a_n7636_8799.n161 a_n7636_8799.n138 4.10845
R468 a_n7636_8799.n93 a_n7636_8799.n70 4.10845
R469 a_n7636_8799.n23 a_n7636_8799.t18 3.61217
R470 a_n7636_8799.n23 a_n7636_8799.t1 3.61217
R471 a_n7636_8799.n21 a_n7636_8799.t3 3.61217
R472 a_n7636_8799.n21 a_n7636_8799.t15 3.61217
R473 a_n7636_8799.n19 a_n7636_8799.t47 3.61217
R474 a_n7636_8799.n19 a_n7636_8799.t10 3.61217
R475 a_n7636_8799.n17 a_n7636_8799.t45 3.61217
R476 a_n7636_8799.n17 a_n7636_8799.t46 3.61217
R477 a_n7636_8799.n15 a_n7636_8799.t7 3.61217
R478 a_n7636_8799.n15 a_n7636_8799.t4 3.61217
R479 a_n7636_8799.n14 a_n7636_8799.t8 3.61217
R480 a_n7636_8799.n14 a_n7636_8799.t11 3.61217
R481 a_n7636_8799.n3 a_n7636_8799.t0 3.61217
R482 a_n7636_8799.n3 a_n7636_8799.t5 3.61217
R483 a_n7636_8799.n4 a_n7636_8799.t6 3.61217
R484 a_n7636_8799.n4 a_n7636_8799.t16 3.61217
R485 a_n7636_8799.n6 a_n7636_8799.t17 3.61217
R486 a_n7636_8799.n6 a_n7636_8799.t12 3.61217
R487 a_n7636_8799.n8 a_n7636_8799.t19 3.61217
R488 a_n7636_8799.n8 a_n7636_8799.t9 3.61217
R489 a_n7636_8799.n10 a_n7636_8799.t14 3.61217
R490 a_n7636_8799.n10 a_n7636_8799.t2 3.61217
R491 a_n7636_8799.n12 a_n7636_8799.t20 3.61217
R492 a_n7636_8799.n12 a_n7636_8799.t13 3.61217
R493 a_n7636_8799.n163 a_n7636_8799.n162 3.4105
R494 a_n7636_8799.n176 a_n7636_8799.t36 2.82907
R495 a_n7636_8799.n176 a_n7636_8799.t34 2.82907
R496 a_n7636_8799.n177 a_n7636_8799.t25 2.82907
R497 a_n7636_8799.n177 a_n7636_8799.t31 2.82907
R498 a_n7636_8799.n179 a_n7636_8799.t43 2.82907
R499 a_n7636_8799.n179 a_n7636_8799.t26 2.82907
R500 a_n7636_8799.n1 a_n7636_8799.t33 2.82907
R501 a_n7636_8799.n1 a_n7636_8799.t32 2.82907
R502 a_n7636_8799.n0 a_n7636_8799.t28 2.82907
R503 a_n7636_8799.n0 a_n7636_8799.t27 2.82907
R504 a_n7636_8799.n174 a_n7636_8799.t39 2.82907
R505 a_n7636_8799.n174 a_n7636_8799.t41 2.82907
R506 a_n7636_8799.n172 a_n7636_8799.t37 2.82907
R507 a_n7636_8799.n172 a_n7636_8799.t21 2.82907
R508 a_n7636_8799.n170 a_n7636_8799.t42 2.82907
R509 a_n7636_8799.n170 a_n7636_8799.t35 2.82907
R510 a_n7636_8799.n167 a_n7636_8799.t22 2.82907
R511 a_n7636_8799.n167 a_n7636_8799.t40 2.82907
R512 a_n7636_8799.n165 a_n7636_8799.t23 2.82907
R513 a_n7636_8799.n165 a_n7636_8799.t24 2.82907
R514 a_n7636_8799.n164 a_n7636_8799.t29 2.82907
R515 a_n7636_8799.n164 a_n7636_8799.t30 2.82907
R516 a_n7636_8799.n183 a_n7636_8799.t38 2.82907
R517 a_n7636_8799.t44 a_n7636_8799.n183 2.82907
R518 a_n7636_8799.n168 a_n7636_8799.n166 0.444466
R519 a_n7636_8799.n173 a_n7636_8799.n171 0.444466
R520 a_n7636_8799.n175 a_n7636_8799.n173 0.444466
R521 a_n7636_8799.n182 a_n7636_8799.n2 0.444466
R522 a_n7636_8799.n180 a_n7636_8799.n178 0.444466
R523 a_n7636_8799.n18 a_n7636_8799.n16 0.358259
R524 a_n7636_8799.n20 a_n7636_8799.n18 0.358259
R525 a_n7636_8799.n22 a_n7636_8799.n20 0.358259
R526 a_n7636_8799.n24 a_n7636_8799.n22 0.358259
R527 a_n7636_8799.n13 a_n7636_8799.n11 0.358259
R528 a_n7636_8799.n11 a_n7636_8799.n9 0.358259
R529 a_n7636_8799.n9 a_n7636_8799.n7 0.358259
R530 a_n7636_8799.n7 a_n7636_8799.n5 0.358259
R531 a_n7636_8799.n169 a_n7636_8799.n168 0.222483
R532 a_n7636_8799.n171 a_n7636_8799.n169 0.222483
R533 a_n7636_8799.n182 a_n7636_8799.n181 0.222483
R534 a_n7636_8799.n181 a_n7636_8799.n180 0.222483
R535 a_n7636_8799.n115 a_n7636_8799.n94 0.189894
R536 a_n7636_8799.n111 a_n7636_8799.n94 0.189894
R537 a_n7636_8799.n111 a_n7636_8799.n110 0.189894
R538 a_n7636_8799.n110 a_n7636_8799.n109 0.189894
R539 a_n7636_8799.n109 a_n7636_8799.n96 0.189894
R540 a_n7636_8799.n97 a_n7636_8799.n96 0.189894
R541 a_n7636_8799.n104 a_n7636_8799.n97 0.189894
R542 a_n7636_8799.n104 a_n7636_8799.n103 0.189894
R543 a_n7636_8799.n103 a_n7636_8799.n102 0.189894
R544 a_n7636_8799.n137 a_n7636_8799.n116 0.189894
R545 a_n7636_8799.n133 a_n7636_8799.n116 0.189894
R546 a_n7636_8799.n133 a_n7636_8799.n132 0.189894
R547 a_n7636_8799.n132 a_n7636_8799.n131 0.189894
R548 a_n7636_8799.n131 a_n7636_8799.n118 0.189894
R549 a_n7636_8799.n119 a_n7636_8799.n118 0.189894
R550 a_n7636_8799.n126 a_n7636_8799.n119 0.189894
R551 a_n7636_8799.n126 a_n7636_8799.n125 0.189894
R552 a_n7636_8799.n125 a_n7636_8799.n124 0.189894
R553 a_n7636_8799.n160 a_n7636_8799.n139 0.189894
R554 a_n7636_8799.n156 a_n7636_8799.n139 0.189894
R555 a_n7636_8799.n156 a_n7636_8799.n155 0.189894
R556 a_n7636_8799.n155 a_n7636_8799.n154 0.189894
R557 a_n7636_8799.n154 a_n7636_8799.n141 0.189894
R558 a_n7636_8799.n142 a_n7636_8799.n141 0.189894
R559 a_n7636_8799.n149 a_n7636_8799.n142 0.189894
R560 a_n7636_8799.n149 a_n7636_8799.n148 0.189894
R561 a_n7636_8799.n148 a_n7636_8799.n147 0.189894
R562 a_n7636_8799.n35 a_n7636_8799.n30 0.189894
R563 a_n7636_8799.n36 a_n7636_8799.n35 0.189894
R564 a_n7636_8799.n37 a_n7636_8799.n36 0.189894
R565 a_n7636_8799.n37 a_n7636_8799.n28 0.189894
R566 a_n7636_8799.n41 a_n7636_8799.n28 0.189894
R567 a_n7636_8799.n42 a_n7636_8799.n41 0.189894
R568 a_n7636_8799.n43 a_n7636_8799.n42 0.189894
R569 a_n7636_8799.n43 a_n7636_8799.n26 0.189894
R570 a_n7636_8799.n47 a_n7636_8799.n26 0.189894
R571 a_n7636_8799.n57 a_n7636_8799.n52 0.189894
R572 a_n7636_8799.n58 a_n7636_8799.n57 0.189894
R573 a_n7636_8799.n59 a_n7636_8799.n58 0.189894
R574 a_n7636_8799.n59 a_n7636_8799.n50 0.189894
R575 a_n7636_8799.n63 a_n7636_8799.n50 0.189894
R576 a_n7636_8799.n64 a_n7636_8799.n63 0.189894
R577 a_n7636_8799.n65 a_n7636_8799.n64 0.189894
R578 a_n7636_8799.n65 a_n7636_8799.n48 0.189894
R579 a_n7636_8799.n69 a_n7636_8799.n48 0.189894
R580 a_n7636_8799.n80 a_n7636_8799.n75 0.189894
R581 a_n7636_8799.n81 a_n7636_8799.n80 0.189894
R582 a_n7636_8799.n82 a_n7636_8799.n81 0.189894
R583 a_n7636_8799.n82 a_n7636_8799.n73 0.189894
R584 a_n7636_8799.n86 a_n7636_8799.n73 0.189894
R585 a_n7636_8799.n87 a_n7636_8799.n86 0.189894
R586 a_n7636_8799.n88 a_n7636_8799.n87 0.189894
R587 a_n7636_8799.n88 a_n7636_8799.n71 0.189894
R588 a_n7636_8799.n92 a_n7636_8799.n71 0.189894
R589 gnd.n7066 gnd.n518 1490.86
R590 gnd.n4043 gnd.n3749 939.716
R591 gnd.n7565 gnd.n206 795.207
R592 gnd.n346 gnd.n209 795.207
R593 gnd.n5378 gnd.n1339 795.207
R594 gnd.n5446 gnd.n1341 795.207
R595 gnd.n6382 gnd.n1091 795.207
R596 gnd.n4665 gnd.n1094 795.207
R597 gnd.n3883 gnd.n3786 795.207
R598 gnd.n3922 gnd.n2262 795.207
R599 gnd.n4653 gnd.n2058 771.183
R600 gnd.n6139 gnd.n1316 771.183
R601 gnd.n4675 gnd.n2069 771.183
R602 gnd.n5534 gnd.n1318 771.183
R603 gnd.n3657 gnd.n2273 766.379
R604 gnd.n3660 gnd.n3659 766.379
R605 gnd.n2899 gnd.n2802 766.379
R606 gnd.n2895 gnd.n2800 766.379
R607 gnd.n3748 gnd.n2295 756.769
R608 gnd.n3651 gnd.n3650 756.769
R609 gnd.n2992 gnd.n2709 756.769
R610 gnd.n2990 gnd.n2712 756.769
R611 gnd.n6644 gnd.n770 756.769
R612 gnd.n7065 gnd.n519 756.769
R613 gnd.n7279 gnd.n7277 756.769
R614 gnd.n6468 gnd.n935 756.769
R615 gnd.n7563 gnd.n211 739.952
R616 gnd.n7454 gnd.n208 739.952
R617 gnd.n5898 gnd.n1338 739.952
R618 gnd.n6121 gnd.n1342 739.952
R619 gnd.n6380 gnd.n1096 739.952
R620 gnd.n4532 gnd.n1093 739.952
R621 gnd.n4046 gnd.n4045 739.952
R622 gnd.n4041 gnd.n2258 739.952
R623 gnd.n6640 gnd.n770 585
R624 gnd.n770 gnd.n769 585
R625 gnd.n6639 gnd.n6638 585
R626 gnd.n6638 gnd.n6637 585
R627 gnd.n773 gnd.n772 585
R628 gnd.n6636 gnd.n773 585
R629 gnd.n6634 gnd.n6633 585
R630 gnd.n6635 gnd.n6634 585
R631 gnd.n6632 gnd.n775 585
R632 gnd.n775 gnd.n774 585
R633 gnd.n6631 gnd.n6630 585
R634 gnd.n6630 gnd.n6629 585
R635 gnd.n781 gnd.n780 585
R636 gnd.n6628 gnd.n781 585
R637 gnd.n6626 gnd.n6625 585
R638 gnd.n6627 gnd.n6626 585
R639 gnd.n6624 gnd.n783 585
R640 gnd.n783 gnd.n782 585
R641 gnd.n6623 gnd.n6622 585
R642 gnd.n6622 gnd.n6621 585
R643 gnd.n789 gnd.n788 585
R644 gnd.n6620 gnd.n789 585
R645 gnd.n6618 gnd.n6617 585
R646 gnd.n6619 gnd.n6618 585
R647 gnd.n6616 gnd.n791 585
R648 gnd.n791 gnd.n790 585
R649 gnd.n6615 gnd.n6614 585
R650 gnd.n6614 gnd.n6613 585
R651 gnd.n797 gnd.n796 585
R652 gnd.n6612 gnd.n797 585
R653 gnd.n6610 gnd.n6609 585
R654 gnd.n6611 gnd.n6610 585
R655 gnd.n6608 gnd.n799 585
R656 gnd.n799 gnd.n798 585
R657 gnd.n6607 gnd.n6606 585
R658 gnd.n6606 gnd.n6605 585
R659 gnd.n805 gnd.n804 585
R660 gnd.n6604 gnd.n805 585
R661 gnd.n6602 gnd.n6601 585
R662 gnd.n6603 gnd.n6602 585
R663 gnd.n6600 gnd.n807 585
R664 gnd.n807 gnd.n806 585
R665 gnd.n6599 gnd.n6598 585
R666 gnd.n6598 gnd.n6597 585
R667 gnd.n813 gnd.n812 585
R668 gnd.n6596 gnd.n813 585
R669 gnd.n6594 gnd.n6593 585
R670 gnd.n6595 gnd.n6594 585
R671 gnd.n6592 gnd.n815 585
R672 gnd.n815 gnd.n814 585
R673 gnd.n6591 gnd.n6590 585
R674 gnd.n6590 gnd.n6589 585
R675 gnd.n821 gnd.n820 585
R676 gnd.n6588 gnd.n821 585
R677 gnd.n6586 gnd.n6585 585
R678 gnd.n6587 gnd.n6586 585
R679 gnd.n6584 gnd.n823 585
R680 gnd.n823 gnd.n822 585
R681 gnd.n6583 gnd.n6582 585
R682 gnd.n6582 gnd.n6581 585
R683 gnd.n829 gnd.n828 585
R684 gnd.n6580 gnd.n829 585
R685 gnd.n6578 gnd.n6577 585
R686 gnd.n6579 gnd.n6578 585
R687 gnd.n6576 gnd.n831 585
R688 gnd.n831 gnd.n830 585
R689 gnd.n6575 gnd.n6574 585
R690 gnd.n6574 gnd.n6573 585
R691 gnd.n837 gnd.n836 585
R692 gnd.n6572 gnd.n837 585
R693 gnd.n6570 gnd.n6569 585
R694 gnd.n6571 gnd.n6570 585
R695 gnd.n6568 gnd.n839 585
R696 gnd.n839 gnd.n838 585
R697 gnd.n6567 gnd.n6566 585
R698 gnd.n6566 gnd.n6565 585
R699 gnd.n845 gnd.n844 585
R700 gnd.n6564 gnd.n845 585
R701 gnd.n6562 gnd.n6561 585
R702 gnd.n6563 gnd.n6562 585
R703 gnd.n6560 gnd.n847 585
R704 gnd.n847 gnd.n846 585
R705 gnd.n6559 gnd.n6558 585
R706 gnd.n6558 gnd.n6557 585
R707 gnd.n853 gnd.n852 585
R708 gnd.n6556 gnd.n853 585
R709 gnd.n6554 gnd.n6553 585
R710 gnd.n6555 gnd.n6554 585
R711 gnd.n6552 gnd.n855 585
R712 gnd.n855 gnd.n854 585
R713 gnd.n6551 gnd.n6550 585
R714 gnd.n6550 gnd.n6549 585
R715 gnd.n861 gnd.n860 585
R716 gnd.n6548 gnd.n861 585
R717 gnd.n6546 gnd.n6545 585
R718 gnd.n6547 gnd.n6546 585
R719 gnd.n6544 gnd.n863 585
R720 gnd.n863 gnd.n862 585
R721 gnd.n6543 gnd.n6542 585
R722 gnd.n6542 gnd.n6541 585
R723 gnd.n869 gnd.n868 585
R724 gnd.n6540 gnd.n869 585
R725 gnd.n6538 gnd.n6537 585
R726 gnd.n6539 gnd.n6538 585
R727 gnd.n6536 gnd.n871 585
R728 gnd.n871 gnd.n870 585
R729 gnd.n6535 gnd.n6534 585
R730 gnd.n6534 gnd.n6533 585
R731 gnd.n877 gnd.n876 585
R732 gnd.n6532 gnd.n877 585
R733 gnd.n6530 gnd.n6529 585
R734 gnd.n6531 gnd.n6530 585
R735 gnd.n6528 gnd.n879 585
R736 gnd.n879 gnd.n878 585
R737 gnd.n6527 gnd.n6526 585
R738 gnd.n6526 gnd.n6525 585
R739 gnd.n885 gnd.n884 585
R740 gnd.n6524 gnd.n885 585
R741 gnd.n6522 gnd.n6521 585
R742 gnd.n6523 gnd.n6522 585
R743 gnd.n6520 gnd.n887 585
R744 gnd.n887 gnd.n886 585
R745 gnd.n6519 gnd.n6518 585
R746 gnd.n6518 gnd.n6517 585
R747 gnd.n893 gnd.n892 585
R748 gnd.n6516 gnd.n893 585
R749 gnd.n6514 gnd.n6513 585
R750 gnd.n6515 gnd.n6514 585
R751 gnd.n6512 gnd.n895 585
R752 gnd.n895 gnd.n894 585
R753 gnd.n6511 gnd.n6510 585
R754 gnd.n6510 gnd.n6509 585
R755 gnd.n901 gnd.n900 585
R756 gnd.n6508 gnd.n901 585
R757 gnd.n6506 gnd.n6505 585
R758 gnd.n6507 gnd.n6506 585
R759 gnd.n6504 gnd.n903 585
R760 gnd.n903 gnd.n902 585
R761 gnd.n6503 gnd.n6502 585
R762 gnd.n6502 gnd.n6501 585
R763 gnd.n909 gnd.n908 585
R764 gnd.n6500 gnd.n909 585
R765 gnd.n6498 gnd.n6497 585
R766 gnd.n6499 gnd.n6498 585
R767 gnd.n6496 gnd.n911 585
R768 gnd.n911 gnd.n910 585
R769 gnd.n6495 gnd.n6494 585
R770 gnd.n6494 gnd.n6493 585
R771 gnd.n917 gnd.n916 585
R772 gnd.n6492 gnd.n917 585
R773 gnd.n6490 gnd.n6489 585
R774 gnd.n6491 gnd.n6490 585
R775 gnd.n6488 gnd.n919 585
R776 gnd.n919 gnd.n918 585
R777 gnd.n6487 gnd.n6486 585
R778 gnd.n6486 gnd.n6485 585
R779 gnd.n925 gnd.n924 585
R780 gnd.n6484 gnd.n925 585
R781 gnd.n6482 gnd.n6481 585
R782 gnd.n6483 gnd.n6482 585
R783 gnd.n6480 gnd.n927 585
R784 gnd.n927 gnd.n926 585
R785 gnd.n6479 gnd.n6478 585
R786 gnd.n6478 gnd.n6477 585
R787 gnd.n933 gnd.n932 585
R788 gnd.n6476 gnd.n933 585
R789 gnd.n6474 gnd.n6473 585
R790 gnd.n6475 gnd.n6474 585
R791 gnd.n6644 gnd.n6643 585
R792 gnd.n6645 gnd.n6644 585
R793 gnd.n768 gnd.n767 585
R794 gnd.n6646 gnd.n768 585
R795 gnd.n6649 gnd.n6648 585
R796 gnd.n6648 gnd.n6647 585
R797 gnd.n765 gnd.n764 585
R798 gnd.n764 gnd.n763 585
R799 gnd.n6654 gnd.n6653 585
R800 gnd.n6655 gnd.n6654 585
R801 gnd.n762 gnd.n761 585
R802 gnd.n6656 gnd.n762 585
R803 gnd.n6659 gnd.n6658 585
R804 gnd.n6658 gnd.n6657 585
R805 gnd.n759 gnd.n758 585
R806 gnd.n758 gnd.n757 585
R807 gnd.n6664 gnd.n6663 585
R808 gnd.n6665 gnd.n6664 585
R809 gnd.n756 gnd.n755 585
R810 gnd.n6666 gnd.n756 585
R811 gnd.n6669 gnd.n6668 585
R812 gnd.n6668 gnd.n6667 585
R813 gnd.n753 gnd.n752 585
R814 gnd.n752 gnd.n751 585
R815 gnd.n6674 gnd.n6673 585
R816 gnd.n6675 gnd.n6674 585
R817 gnd.n750 gnd.n749 585
R818 gnd.n6676 gnd.n750 585
R819 gnd.n6679 gnd.n6678 585
R820 gnd.n6678 gnd.n6677 585
R821 gnd.n747 gnd.n746 585
R822 gnd.n746 gnd.n745 585
R823 gnd.n6684 gnd.n6683 585
R824 gnd.n6685 gnd.n6684 585
R825 gnd.n744 gnd.n743 585
R826 gnd.n6686 gnd.n744 585
R827 gnd.n6689 gnd.n6688 585
R828 gnd.n6688 gnd.n6687 585
R829 gnd.n741 gnd.n740 585
R830 gnd.n740 gnd.n739 585
R831 gnd.n6694 gnd.n6693 585
R832 gnd.n6695 gnd.n6694 585
R833 gnd.n738 gnd.n737 585
R834 gnd.n6696 gnd.n738 585
R835 gnd.n6699 gnd.n6698 585
R836 gnd.n6698 gnd.n6697 585
R837 gnd.n735 gnd.n734 585
R838 gnd.n734 gnd.n733 585
R839 gnd.n6704 gnd.n6703 585
R840 gnd.n6705 gnd.n6704 585
R841 gnd.n732 gnd.n731 585
R842 gnd.n6706 gnd.n732 585
R843 gnd.n6709 gnd.n6708 585
R844 gnd.n6708 gnd.n6707 585
R845 gnd.n729 gnd.n728 585
R846 gnd.n728 gnd.n727 585
R847 gnd.n6714 gnd.n6713 585
R848 gnd.n6715 gnd.n6714 585
R849 gnd.n726 gnd.n725 585
R850 gnd.n6716 gnd.n726 585
R851 gnd.n6719 gnd.n6718 585
R852 gnd.n6718 gnd.n6717 585
R853 gnd.n723 gnd.n722 585
R854 gnd.n722 gnd.n721 585
R855 gnd.n6724 gnd.n6723 585
R856 gnd.n6725 gnd.n6724 585
R857 gnd.n720 gnd.n719 585
R858 gnd.n6726 gnd.n720 585
R859 gnd.n6729 gnd.n6728 585
R860 gnd.n6728 gnd.n6727 585
R861 gnd.n717 gnd.n716 585
R862 gnd.n716 gnd.n715 585
R863 gnd.n6734 gnd.n6733 585
R864 gnd.n6735 gnd.n6734 585
R865 gnd.n714 gnd.n713 585
R866 gnd.n6736 gnd.n714 585
R867 gnd.n6739 gnd.n6738 585
R868 gnd.n6738 gnd.n6737 585
R869 gnd.n711 gnd.n710 585
R870 gnd.n710 gnd.n709 585
R871 gnd.n6744 gnd.n6743 585
R872 gnd.n6745 gnd.n6744 585
R873 gnd.n708 gnd.n707 585
R874 gnd.n6746 gnd.n708 585
R875 gnd.n6749 gnd.n6748 585
R876 gnd.n6748 gnd.n6747 585
R877 gnd.n705 gnd.n704 585
R878 gnd.n704 gnd.n703 585
R879 gnd.n6754 gnd.n6753 585
R880 gnd.n6755 gnd.n6754 585
R881 gnd.n702 gnd.n701 585
R882 gnd.n6756 gnd.n702 585
R883 gnd.n6759 gnd.n6758 585
R884 gnd.n6758 gnd.n6757 585
R885 gnd.n699 gnd.n698 585
R886 gnd.n698 gnd.n697 585
R887 gnd.n6764 gnd.n6763 585
R888 gnd.n6765 gnd.n6764 585
R889 gnd.n696 gnd.n695 585
R890 gnd.n6766 gnd.n696 585
R891 gnd.n6769 gnd.n6768 585
R892 gnd.n6768 gnd.n6767 585
R893 gnd.n693 gnd.n692 585
R894 gnd.n692 gnd.n691 585
R895 gnd.n6774 gnd.n6773 585
R896 gnd.n6775 gnd.n6774 585
R897 gnd.n690 gnd.n689 585
R898 gnd.n6776 gnd.n690 585
R899 gnd.n6779 gnd.n6778 585
R900 gnd.n6778 gnd.n6777 585
R901 gnd.n687 gnd.n686 585
R902 gnd.n686 gnd.n685 585
R903 gnd.n6784 gnd.n6783 585
R904 gnd.n6785 gnd.n6784 585
R905 gnd.n684 gnd.n683 585
R906 gnd.n6786 gnd.n684 585
R907 gnd.n6789 gnd.n6788 585
R908 gnd.n6788 gnd.n6787 585
R909 gnd.n681 gnd.n680 585
R910 gnd.n680 gnd.n679 585
R911 gnd.n6794 gnd.n6793 585
R912 gnd.n6795 gnd.n6794 585
R913 gnd.n678 gnd.n677 585
R914 gnd.n6796 gnd.n678 585
R915 gnd.n6799 gnd.n6798 585
R916 gnd.n6798 gnd.n6797 585
R917 gnd.n675 gnd.n674 585
R918 gnd.n674 gnd.n673 585
R919 gnd.n6804 gnd.n6803 585
R920 gnd.n6805 gnd.n6804 585
R921 gnd.n672 gnd.n671 585
R922 gnd.n6806 gnd.n672 585
R923 gnd.n6809 gnd.n6808 585
R924 gnd.n6808 gnd.n6807 585
R925 gnd.n669 gnd.n668 585
R926 gnd.n668 gnd.n667 585
R927 gnd.n6814 gnd.n6813 585
R928 gnd.n6815 gnd.n6814 585
R929 gnd.n666 gnd.n665 585
R930 gnd.n6816 gnd.n666 585
R931 gnd.n6819 gnd.n6818 585
R932 gnd.n6818 gnd.n6817 585
R933 gnd.n663 gnd.n662 585
R934 gnd.n662 gnd.n661 585
R935 gnd.n6824 gnd.n6823 585
R936 gnd.n6825 gnd.n6824 585
R937 gnd.n660 gnd.n659 585
R938 gnd.n6826 gnd.n660 585
R939 gnd.n6829 gnd.n6828 585
R940 gnd.n6828 gnd.n6827 585
R941 gnd.n657 gnd.n656 585
R942 gnd.n656 gnd.n655 585
R943 gnd.n6834 gnd.n6833 585
R944 gnd.n6835 gnd.n6834 585
R945 gnd.n654 gnd.n653 585
R946 gnd.n6836 gnd.n654 585
R947 gnd.n6839 gnd.n6838 585
R948 gnd.n6838 gnd.n6837 585
R949 gnd.n651 gnd.n650 585
R950 gnd.n650 gnd.n649 585
R951 gnd.n6844 gnd.n6843 585
R952 gnd.n6845 gnd.n6844 585
R953 gnd.n648 gnd.n647 585
R954 gnd.n6846 gnd.n648 585
R955 gnd.n6849 gnd.n6848 585
R956 gnd.n6848 gnd.n6847 585
R957 gnd.n645 gnd.n644 585
R958 gnd.n644 gnd.n643 585
R959 gnd.n6854 gnd.n6853 585
R960 gnd.n6855 gnd.n6854 585
R961 gnd.n642 gnd.n641 585
R962 gnd.n6856 gnd.n642 585
R963 gnd.n6859 gnd.n6858 585
R964 gnd.n6858 gnd.n6857 585
R965 gnd.n639 gnd.n638 585
R966 gnd.n638 gnd.n637 585
R967 gnd.n6864 gnd.n6863 585
R968 gnd.n6865 gnd.n6864 585
R969 gnd.n636 gnd.n635 585
R970 gnd.n6866 gnd.n636 585
R971 gnd.n6869 gnd.n6868 585
R972 gnd.n6868 gnd.n6867 585
R973 gnd.n633 gnd.n632 585
R974 gnd.n632 gnd.n631 585
R975 gnd.n6874 gnd.n6873 585
R976 gnd.n6875 gnd.n6874 585
R977 gnd.n630 gnd.n629 585
R978 gnd.n6876 gnd.n630 585
R979 gnd.n6879 gnd.n6878 585
R980 gnd.n6878 gnd.n6877 585
R981 gnd.n627 gnd.n626 585
R982 gnd.n626 gnd.n625 585
R983 gnd.n6884 gnd.n6883 585
R984 gnd.n6885 gnd.n6884 585
R985 gnd.n624 gnd.n623 585
R986 gnd.n6886 gnd.n624 585
R987 gnd.n6889 gnd.n6888 585
R988 gnd.n6888 gnd.n6887 585
R989 gnd.n621 gnd.n620 585
R990 gnd.n620 gnd.n619 585
R991 gnd.n6894 gnd.n6893 585
R992 gnd.n6895 gnd.n6894 585
R993 gnd.n618 gnd.n617 585
R994 gnd.n6896 gnd.n618 585
R995 gnd.n6899 gnd.n6898 585
R996 gnd.n6898 gnd.n6897 585
R997 gnd.n615 gnd.n614 585
R998 gnd.n614 gnd.n613 585
R999 gnd.n6904 gnd.n6903 585
R1000 gnd.n6905 gnd.n6904 585
R1001 gnd.n612 gnd.n611 585
R1002 gnd.n6906 gnd.n612 585
R1003 gnd.n6909 gnd.n6908 585
R1004 gnd.n6908 gnd.n6907 585
R1005 gnd.n609 gnd.n608 585
R1006 gnd.n608 gnd.n607 585
R1007 gnd.n6914 gnd.n6913 585
R1008 gnd.n6915 gnd.n6914 585
R1009 gnd.n606 gnd.n605 585
R1010 gnd.n6916 gnd.n606 585
R1011 gnd.n6919 gnd.n6918 585
R1012 gnd.n6918 gnd.n6917 585
R1013 gnd.n603 gnd.n602 585
R1014 gnd.n602 gnd.n601 585
R1015 gnd.n6924 gnd.n6923 585
R1016 gnd.n6925 gnd.n6924 585
R1017 gnd.n600 gnd.n599 585
R1018 gnd.n6926 gnd.n600 585
R1019 gnd.n6929 gnd.n6928 585
R1020 gnd.n6928 gnd.n6927 585
R1021 gnd.n597 gnd.n596 585
R1022 gnd.n596 gnd.n595 585
R1023 gnd.n6934 gnd.n6933 585
R1024 gnd.n6935 gnd.n6934 585
R1025 gnd.n594 gnd.n593 585
R1026 gnd.n6936 gnd.n594 585
R1027 gnd.n6939 gnd.n6938 585
R1028 gnd.n6938 gnd.n6937 585
R1029 gnd.n591 gnd.n590 585
R1030 gnd.n590 gnd.n589 585
R1031 gnd.n6944 gnd.n6943 585
R1032 gnd.n6945 gnd.n6944 585
R1033 gnd.n588 gnd.n587 585
R1034 gnd.n6946 gnd.n588 585
R1035 gnd.n6949 gnd.n6948 585
R1036 gnd.n6948 gnd.n6947 585
R1037 gnd.n585 gnd.n584 585
R1038 gnd.n584 gnd.n583 585
R1039 gnd.n6954 gnd.n6953 585
R1040 gnd.n6955 gnd.n6954 585
R1041 gnd.n582 gnd.n581 585
R1042 gnd.n6956 gnd.n582 585
R1043 gnd.n6959 gnd.n6958 585
R1044 gnd.n6958 gnd.n6957 585
R1045 gnd.n579 gnd.n578 585
R1046 gnd.n578 gnd.n577 585
R1047 gnd.n6964 gnd.n6963 585
R1048 gnd.n6965 gnd.n6964 585
R1049 gnd.n576 gnd.n575 585
R1050 gnd.n6966 gnd.n576 585
R1051 gnd.n6969 gnd.n6968 585
R1052 gnd.n6968 gnd.n6967 585
R1053 gnd.n573 gnd.n572 585
R1054 gnd.n572 gnd.n571 585
R1055 gnd.n6974 gnd.n6973 585
R1056 gnd.n6975 gnd.n6974 585
R1057 gnd.n570 gnd.n569 585
R1058 gnd.n6976 gnd.n570 585
R1059 gnd.n6979 gnd.n6978 585
R1060 gnd.n6978 gnd.n6977 585
R1061 gnd.n567 gnd.n566 585
R1062 gnd.n566 gnd.n565 585
R1063 gnd.n6984 gnd.n6983 585
R1064 gnd.n6985 gnd.n6984 585
R1065 gnd.n564 gnd.n563 585
R1066 gnd.n6986 gnd.n564 585
R1067 gnd.n6989 gnd.n6988 585
R1068 gnd.n6988 gnd.n6987 585
R1069 gnd.n561 gnd.n560 585
R1070 gnd.n560 gnd.n559 585
R1071 gnd.n6994 gnd.n6993 585
R1072 gnd.n6995 gnd.n6994 585
R1073 gnd.n558 gnd.n557 585
R1074 gnd.n6996 gnd.n558 585
R1075 gnd.n6999 gnd.n6998 585
R1076 gnd.n6998 gnd.n6997 585
R1077 gnd.n555 gnd.n554 585
R1078 gnd.n554 gnd.n553 585
R1079 gnd.n7004 gnd.n7003 585
R1080 gnd.n7005 gnd.n7004 585
R1081 gnd.n552 gnd.n551 585
R1082 gnd.n7006 gnd.n552 585
R1083 gnd.n7009 gnd.n7008 585
R1084 gnd.n7008 gnd.n7007 585
R1085 gnd.n549 gnd.n548 585
R1086 gnd.n548 gnd.n547 585
R1087 gnd.n7014 gnd.n7013 585
R1088 gnd.n7015 gnd.n7014 585
R1089 gnd.n546 gnd.n545 585
R1090 gnd.n7016 gnd.n546 585
R1091 gnd.n7019 gnd.n7018 585
R1092 gnd.n7018 gnd.n7017 585
R1093 gnd.n543 gnd.n542 585
R1094 gnd.n542 gnd.n541 585
R1095 gnd.n7024 gnd.n7023 585
R1096 gnd.n7025 gnd.n7024 585
R1097 gnd.n540 gnd.n539 585
R1098 gnd.n7026 gnd.n540 585
R1099 gnd.n7029 gnd.n7028 585
R1100 gnd.n7028 gnd.n7027 585
R1101 gnd.n537 gnd.n536 585
R1102 gnd.n536 gnd.n535 585
R1103 gnd.n7034 gnd.n7033 585
R1104 gnd.n7035 gnd.n7034 585
R1105 gnd.n534 gnd.n533 585
R1106 gnd.n7036 gnd.n534 585
R1107 gnd.n7039 gnd.n7038 585
R1108 gnd.n7038 gnd.n7037 585
R1109 gnd.n531 gnd.n530 585
R1110 gnd.n530 gnd.n529 585
R1111 gnd.n7044 gnd.n7043 585
R1112 gnd.n7045 gnd.n7044 585
R1113 gnd.n528 gnd.n527 585
R1114 gnd.n7046 gnd.n528 585
R1115 gnd.n7049 gnd.n7048 585
R1116 gnd.n7048 gnd.n7047 585
R1117 gnd.n525 gnd.n524 585
R1118 gnd.n524 gnd.n523 585
R1119 gnd.n7055 gnd.n7054 585
R1120 gnd.n7056 gnd.n7055 585
R1121 gnd.n522 gnd.n521 585
R1122 gnd.n7057 gnd.n522 585
R1123 gnd.n7060 gnd.n7059 585
R1124 gnd.n7059 gnd.n7058 585
R1125 gnd.n7061 gnd.n519 585
R1126 gnd.n519 gnd.n518 585
R1127 gnd.n394 gnd.n393 585
R1128 gnd.n7268 gnd.n393 585
R1129 gnd.n7271 gnd.n7270 585
R1130 gnd.n7270 gnd.n7269 585
R1131 gnd.n397 gnd.n396 585
R1132 gnd.n7267 gnd.n397 585
R1133 gnd.n7265 gnd.n7264 585
R1134 gnd.n7266 gnd.n7265 585
R1135 gnd.n400 gnd.n399 585
R1136 gnd.n399 gnd.n398 585
R1137 gnd.n7260 gnd.n7259 585
R1138 gnd.n7259 gnd.n7258 585
R1139 gnd.n403 gnd.n402 585
R1140 gnd.n7257 gnd.n403 585
R1141 gnd.n7255 gnd.n7254 585
R1142 gnd.n7256 gnd.n7255 585
R1143 gnd.n406 gnd.n405 585
R1144 gnd.n405 gnd.n404 585
R1145 gnd.n7250 gnd.n7249 585
R1146 gnd.n7249 gnd.n7248 585
R1147 gnd.n409 gnd.n408 585
R1148 gnd.n7247 gnd.n409 585
R1149 gnd.n7245 gnd.n7244 585
R1150 gnd.n7246 gnd.n7245 585
R1151 gnd.n412 gnd.n411 585
R1152 gnd.n411 gnd.n410 585
R1153 gnd.n7240 gnd.n7239 585
R1154 gnd.n7239 gnd.n7238 585
R1155 gnd.n415 gnd.n414 585
R1156 gnd.n7237 gnd.n415 585
R1157 gnd.n7235 gnd.n7234 585
R1158 gnd.n7236 gnd.n7235 585
R1159 gnd.n418 gnd.n417 585
R1160 gnd.n417 gnd.n416 585
R1161 gnd.n7230 gnd.n7229 585
R1162 gnd.n7229 gnd.n7228 585
R1163 gnd.n421 gnd.n420 585
R1164 gnd.n7227 gnd.n421 585
R1165 gnd.n7225 gnd.n7224 585
R1166 gnd.n7226 gnd.n7225 585
R1167 gnd.n424 gnd.n423 585
R1168 gnd.n423 gnd.n422 585
R1169 gnd.n7220 gnd.n7219 585
R1170 gnd.n7219 gnd.n7218 585
R1171 gnd.n427 gnd.n426 585
R1172 gnd.n7217 gnd.n427 585
R1173 gnd.n7215 gnd.n7214 585
R1174 gnd.n7216 gnd.n7215 585
R1175 gnd.n430 gnd.n429 585
R1176 gnd.n429 gnd.n428 585
R1177 gnd.n7210 gnd.n7209 585
R1178 gnd.n7209 gnd.n7208 585
R1179 gnd.n433 gnd.n432 585
R1180 gnd.n7207 gnd.n433 585
R1181 gnd.n7205 gnd.n7204 585
R1182 gnd.n7206 gnd.n7205 585
R1183 gnd.n436 gnd.n435 585
R1184 gnd.n435 gnd.n434 585
R1185 gnd.n7200 gnd.n7199 585
R1186 gnd.n7199 gnd.n7198 585
R1187 gnd.n439 gnd.n438 585
R1188 gnd.n7197 gnd.n439 585
R1189 gnd.n7195 gnd.n7194 585
R1190 gnd.n7196 gnd.n7195 585
R1191 gnd.n442 gnd.n441 585
R1192 gnd.n441 gnd.n440 585
R1193 gnd.n7190 gnd.n7189 585
R1194 gnd.n7189 gnd.n7188 585
R1195 gnd.n445 gnd.n444 585
R1196 gnd.n7187 gnd.n445 585
R1197 gnd.n7185 gnd.n7184 585
R1198 gnd.n7186 gnd.n7185 585
R1199 gnd.n448 gnd.n447 585
R1200 gnd.n447 gnd.n446 585
R1201 gnd.n7180 gnd.n7179 585
R1202 gnd.n7179 gnd.n7178 585
R1203 gnd.n451 gnd.n450 585
R1204 gnd.n7177 gnd.n451 585
R1205 gnd.n7175 gnd.n7174 585
R1206 gnd.n7176 gnd.n7175 585
R1207 gnd.n454 gnd.n453 585
R1208 gnd.n453 gnd.n452 585
R1209 gnd.n7170 gnd.n7169 585
R1210 gnd.n7169 gnd.n7168 585
R1211 gnd.n457 gnd.n456 585
R1212 gnd.n7167 gnd.n457 585
R1213 gnd.n7165 gnd.n7164 585
R1214 gnd.n7166 gnd.n7165 585
R1215 gnd.n460 gnd.n459 585
R1216 gnd.n459 gnd.n458 585
R1217 gnd.n7160 gnd.n7159 585
R1218 gnd.n7159 gnd.n7158 585
R1219 gnd.n463 gnd.n462 585
R1220 gnd.n7157 gnd.n463 585
R1221 gnd.n7155 gnd.n7154 585
R1222 gnd.n7156 gnd.n7155 585
R1223 gnd.n466 gnd.n465 585
R1224 gnd.n465 gnd.n464 585
R1225 gnd.n7150 gnd.n7149 585
R1226 gnd.n7149 gnd.n7148 585
R1227 gnd.n469 gnd.n468 585
R1228 gnd.n7147 gnd.n469 585
R1229 gnd.n7145 gnd.n7144 585
R1230 gnd.n7146 gnd.n7145 585
R1231 gnd.n472 gnd.n471 585
R1232 gnd.n471 gnd.n470 585
R1233 gnd.n7140 gnd.n7139 585
R1234 gnd.n7139 gnd.n7138 585
R1235 gnd.n475 gnd.n474 585
R1236 gnd.n7137 gnd.n475 585
R1237 gnd.n7135 gnd.n7134 585
R1238 gnd.n7136 gnd.n7135 585
R1239 gnd.n478 gnd.n477 585
R1240 gnd.n477 gnd.n476 585
R1241 gnd.n7130 gnd.n7129 585
R1242 gnd.n7129 gnd.n7128 585
R1243 gnd.n481 gnd.n480 585
R1244 gnd.n7127 gnd.n481 585
R1245 gnd.n7125 gnd.n7124 585
R1246 gnd.n7126 gnd.n7125 585
R1247 gnd.n484 gnd.n483 585
R1248 gnd.n483 gnd.n482 585
R1249 gnd.n7120 gnd.n7119 585
R1250 gnd.n7119 gnd.n7118 585
R1251 gnd.n487 gnd.n486 585
R1252 gnd.n7117 gnd.n487 585
R1253 gnd.n7115 gnd.n7114 585
R1254 gnd.n7116 gnd.n7115 585
R1255 gnd.n490 gnd.n489 585
R1256 gnd.n489 gnd.n488 585
R1257 gnd.n7110 gnd.n7109 585
R1258 gnd.n7109 gnd.n7108 585
R1259 gnd.n493 gnd.n492 585
R1260 gnd.n7107 gnd.n493 585
R1261 gnd.n7105 gnd.n7104 585
R1262 gnd.n7106 gnd.n7105 585
R1263 gnd.n496 gnd.n495 585
R1264 gnd.n495 gnd.n494 585
R1265 gnd.n7100 gnd.n7099 585
R1266 gnd.n7099 gnd.n7098 585
R1267 gnd.n499 gnd.n498 585
R1268 gnd.n7097 gnd.n499 585
R1269 gnd.n7095 gnd.n7094 585
R1270 gnd.n7096 gnd.n7095 585
R1271 gnd.n502 gnd.n501 585
R1272 gnd.n501 gnd.n500 585
R1273 gnd.n7090 gnd.n7089 585
R1274 gnd.n7089 gnd.n7088 585
R1275 gnd.n505 gnd.n504 585
R1276 gnd.n7087 gnd.n505 585
R1277 gnd.n7085 gnd.n7084 585
R1278 gnd.n7086 gnd.n7085 585
R1279 gnd.n508 gnd.n507 585
R1280 gnd.n507 gnd.n506 585
R1281 gnd.n7080 gnd.n7079 585
R1282 gnd.n7079 gnd.n7078 585
R1283 gnd.n511 gnd.n510 585
R1284 gnd.n7077 gnd.n511 585
R1285 gnd.n7075 gnd.n7074 585
R1286 gnd.n7076 gnd.n7075 585
R1287 gnd.n514 gnd.n513 585
R1288 gnd.n513 gnd.n512 585
R1289 gnd.n7070 gnd.n7069 585
R1290 gnd.n7069 gnd.n7068 585
R1291 gnd.n517 gnd.n516 585
R1292 gnd.n7067 gnd.n517 585
R1293 gnd.n7065 gnd.n7064 585
R1294 gnd.n7066 gnd.n7065 585
R1295 gnd.n6383 gnd.n6382 585
R1296 gnd.n6382 gnd.n6381 585
R1297 gnd.n6384 gnd.n1087 585
R1298 gnd.n4358 gnd.n1087 585
R1299 gnd.n6386 gnd.n6385 585
R1300 gnd.n6387 gnd.n6386 585
R1301 gnd.n1071 gnd.n1070 585
R1302 gnd.n4351 gnd.n1071 585
R1303 gnd.n6395 gnd.n6394 585
R1304 gnd.n6394 gnd.n6393 585
R1305 gnd.n6396 gnd.n1066 585
R1306 gnd.n4346 gnd.n1066 585
R1307 gnd.n6398 gnd.n6397 585
R1308 gnd.n6399 gnd.n6398 585
R1309 gnd.n1051 gnd.n1050 585
R1310 gnd.n4373 gnd.n1051 585
R1311 gnd.n6407 gnd.n6406 585
R1312 gnd.n6406 gnd.n6405 585
R1313 gnd.n6408 gnd.n1046 585
R1314 gnd.n4339 gnd.n1046 585
R1315 gnd.n6410 gnd.n6409 585
R1316 gnd.n6411 gnd.n6410 585
R1317 gnd.n1031 gnd.n1030 585
R1318 gnd.n4331 gnd.n1031 585
R1319 gnd.n6419 gnd.n6418 585
R1320 gnd.n6418 gnd.n6417 585
R1321 gnd.n6420 gnd.n1026 585
R1322 gnd.n4324 gnd.n1026 585
R1323 gnd.n6422 gnd.n6421 585
R1324 gnd.n6423 gnd.n6422 585
R1325 gnd.n1011 gnd.n1010 585
R1326 gnd.n4316 gnd.n1011 585
R1327 gnd.n6431 gnd.n6430 585
R1328 gnd.n6430 gnd.n6429 585
R1329 gnd.n6432 gnd.n1006 585
R1330 gnd.n4263 gnd.n1006 585
R1331 gnd.n6434 gnd.n6433 585
R1332 gnd.n6435 gnd.n6434 585
R1333 gnd.n992 gnd.n991 585
R1334 gnd.n4254 gnd.n992 585
R1335 gnd.n6443 gnd.n6442 585
R1336 gnd.n6442 gnd.n6441 585
R1337 gnd.n6444 gnd.n986 585
R1338 gnd.n4248 gnd.n986 585
R1339 gnd.n6446 gnd.n6445 585
R1340 gnd.n6447 gnd.n6446 585
R1341 gnd.n987 gnd.n985 585
R1342 gnd.n4277 gnd.n985 585
R1343 gnd.n4243 gnd.n4242 585
R1344 gnd.n4242 gnd.n4241 585
R1345 gnd.n2144 gnd.n2143 585
R1346 gnd.n4236 gnd.n2144 585
R1347 gnd.n4218 gnd.n4217 585
R1348 gnd.n4217 gnd.n4216 585
R1349 gnd.n4219 gnd.n2156 585
R1350 gnd.n4227 gnd.n2156 585
R1351 gnd.n4221 gnd.n4220 585
R1352 gnd.n4222 gnd.n4221 585
R1353 gnd.n2163 gnd.n2162 585
R1354 gnd.n4176 gnd.n2162 585
R1355 gnd.n964 gnd.n963 585
R1356 gnd.n4178 gnd.n964 585
R1357 gnd.n6456 gnd.n6455 585
R1358 gnd.n6455 gnd.n6454 585
R1359 gnd.n6457 gnd.n958 585
R1360 gnd.n4184 gnd.n958 585
R1361 gnd.n6459 gnd.n6458 585
R1362 gnd.n6460 gnd.n6459 585
R1363 gnd.n959 gnd.n957 585
R1364 gnd.n4190 gnd.n957 585
R1365 gnd.n4156 gnd.n945 585
R1366 gnd.n6466 gnd.n945 585
R1367 gnd.n4155 gnd.n4154 585
R1368 gnd.n4154 gnd.n941 585
R1369 gnd.n4153 gnd.n2181 585
R1370 gnd.n4153 gnd.n4152 585
R1371 gnd.n4140 gnd.n2182 585
R1372 gnd.n4136 gnd.n2182 585
R1373 gnd.n4142 gnd.n4141 585
R1374 gnd.n4143 gnd.n4142 585
R1375 gnd.n2195 gnd.n2194 585
R1376 gnd.n2194 gnd.n2191 585
R1377 gnd.n4109 gnd.n2207 585
R1378 gnd.n4121 gnd.n2207 585
R1379 gnd.n4110 gnd.n2217 585
R1380 gnd.n2217 gnd.n2215 585
R1381 gnd.n4112 gnd.n4111 585
R1382 gnd.n4113 gnd.n4112 585
R1383 gnd.n2218 gnd.n2216 585
R1384 gnd.n4099 gnd.n2216 585
R1385 gnd.n4072 gnd.n4071 585
R1386 gnd.n4071 gnd.n2225 585
R1387 gnd.n4073 gnd.n2232 585
R1388 gnd.n4087 gnd.n2232 585
R1389 gnd.n4074 gnd.n2244 585
R1390 gnd.n2244 gnd.n2242 585
R1391 gnd.n4076 gnd.n4075 585
R1392 gnd.n4077 gnd.n4076 585
R1393 gnd.n2245 gnd.n2243 585
R1394 gnd.n2243 gnd.n2239 585
R1395 gnd.n2267 gnd.n2253 585
R1396 gnd.n4061 gnd.n2253 585
R1397 gnd.n2265 gnd.n2263 585
R1398 gnd.n2263 gnd.n2251 585
R1399 gnd.n4052 gnd.n4051 585
R1400 gnd.n4053 gnd.n4052 585
R1401 gnd.n2264 gnd.n2262 585
R1402 gnd.n2262 gnd.n2259 585
R1403 gnd.n3923 gnd.n3922 585
R1404 gnd.n3921 gnd.n3920 585
R1405 gnd.n3919 gnd.n3918 585
R1406 gnd.n3917 gnd.n3916 585
R1407 gnd.n3915 gnd.n3914 585
R1408 gnd.n3913 gnd.n3912 585
R1409 gnd.n3911 gnd.n3910 585
R1410 gnd.n3909 gnd.n3908 585
R1411 gnd.n3907 gnd.n3906 585
R1412 gnd.n3905 gnd.n3904 585
R1413 gnd.n3903 gnd.n3902 585
R1414 gnd.n3901 gnd.n3900 585
R1415 gnd.n3899 gnd.n3898 585
R1416 gnd.n3897 gnd.n3896 585
R1417 gnd.n3895 gnd.n3894 585
R1418 gnd.n3893 gnd.n3892 585
R1419 gnd.n3891 gnd.n3890 585
R1420 gnd.n3870 gnd.n3867 585
R1421 gnd.n3886 gnd.n3786 585
R1422 gnd.n4043 gnd.n3786 585
R1423 gnd.n4666 gnd.n4665 585
R1424 gnd.n4663 gnd.n2077 585
R1425 gnd.n4662 gnd.n4661 585
R1426 gnd.n4593 gnd.n2079 585
R1427 gnd.n4602 gnd.n4594 585
R1428 gnd.n4603 gnd.n4591 585
R1429 gnd.n4590 gnd.n4583 585
R1430 gnd.n4610 gnd.n4582 585
R1431 gnd.n4611 gnd.n4581 585
R1432 gnd.n4579 gnd.n4571 585
R1433 gnd.n4618 gnd.n4570 585
R1434 gnd.n4619 gnd.n4568 585
R1435 gnd.n4567 gnd.n4560 585
R1436 gnd.n4626 gnd.n4559 585
R1437 gnd.n4627 gnd.n4558 585
R1438 gnd.n4556 gnd.n4548 585
R1439 gnd.n4634 gnd.n4547 585
R1440 gnd.n4635 gnd.n4545 585
R1441 gnd.n4544 gnd.n1091 585
R1442 gnd.n1100 gnd.n1091 585
R1443 gnd.n4360 gnd.n1094 585
R1444 gnd.n6381 gnd.n1094 585
R1445 gnd.n4361 gnd.n4359 585
R1446 gnd.n4359 gnd.n4358 585
R1447 gnd.n2108 gnd.n1085 585
R1448 gnd.n6387 gnd.n1085 585
R1449 gnd.n4365 gnd.n2107 585
R1450 gnd.n4351 gnd.n2107 585
R1451 gnd.n4366 gnd.n1074 585
R1452 gnd.n6393 gnd.n1074 585
R1453 gnd.n4367 gnd.n2106 585
R1454 gnd.n4346 gnd.n2106 585
R1455 gnd.n2103 gnd.n1064 585
R1456 gnd.n6399 gnd.n1064 585
R1457 gnd.n4372 gnd.n4371 585
R1458 gnd.n4373 gnd.n4372 585
R1459 gnd.n2102 gnd.n1054 585
R1460 gnd.n6405 gnd.n1054 585
R1461 gnd.n4338 gnd.n4337 585
R1462 gnd.n4339 gnd.n4338 585
R1463 gnd.n2111 gnd.n1044 585
R1464 gnd.n6411 gnd.n1044 585
R1465 gnd.n4333 gnd.n4332 585
R1466 gnd.n4332 gnd.n4331 585
R1467 gnd.n2113 gnd.n1034 585
R1468 gnd.n6417 gnd.n1034 585
R1469 gnd.n4323 gnd.n4322 585
R1470 gnd.n4324 gnd.n4323 585
R1471 gnd.n2116 gnd.n1024 585
R1472 gnd.n6423 gnd.n1024 585
R1473 gnd.n4318 gnd.n4317 585
R1474 gnd.n4317 gnd.n4316 585
R1475 gnd.n2118 gnd.n1014 585
R1476 gnd.n6429 gnd.n1014 585
R1477 gnd.n4265 gnd.n4264 585
R1478 gnd.n4264 gnd.n4263 585
R1479 gnd.n2140 gnd.n1004 585
R1480 gnd.n6435 gnd.n1004 585
R1481 gnd.n4269 gnd.n2139 585
R1482 gnd.n4254 gnd.n2139 585
R1483 gnd.n4270 gnd.n995 585
R1484 gnd.n6441 gnd.n995 585
R1485 gnd.n4271 gnd.n2138 585
R1486 gnd.n4248 gnd.n2138 585
R1487 gnd.n2135 gnd.n983 585
R1488 gnd.n6447 gnd.n983 585
R1489 gnd.n4276 gnd.n4275 585
R1490 gnd.n4277 gnd.n4276 585
R1491 gnd.n2134 gnd.n2133 585
R1492 gnd.n4241 gnd.n2133 585
R1493 gnd.n4235 gnd.n4234 585
R1494 gnd.n4236 gnd.n4235 585
R1495 gnd.n2150 gnd.n2149 585
R1496 gnd.n4216 gnd.n2149 585
R1497 gnd.n4229 gnd.n4228 585
R1498 gnd.n4228 gnd.n4227 585
R1499 gnd.n2153 gnd.n2152 585
R1500 gnd.n4222 gnd.n2153 585
R1501 gnd.n4175 gnd.n4174 585
R1502 gnd.n4176 gnd.n4175 585
R1503 gnd.n4170 gnd.n4169 585
R1504 gnd.n4178 gnd.n4169 585
R1505 gnd.n2178 gnd.n967 585
R1506 gnd.n6454 gnd.n967 585
R1507 gnd.n4186 gnd.n4185 585
R1508 gnd.n4185 gnd.n4184 585
R1509 gnd.n4187 gnd.n955 585
R1510 gnd.n6460 gnd.n955 585
R1511 gnd.n4189 gnd.n4188 585
R1512 gnd.n4190 gnd.n4189 585
R1513 gnd.n2174 gnd.n943 585
R1514 gnd.n6466 gnd.n943 585
R1515 gnd.n4132 gnd.n4131 585
R1516 gnd.n4131 gnd.n941 585
R1517 gnd.n4133 gnd.n2185 585
R1518 gnd.n4152 gnd.n2185 585
R1519 gnd.n4135 gnd.n4134 585
R1520 gnd.n4136 gnd.n4135 585
R1521 gnd.n2202 gnd.n2193 585
R1522 gnd.n4143 gnd.n2193 585
R1523 gnd.n4124 gnd.n4123 585
R1524 gnd.n4123 gnd.n2191 585
R1525 gnd.n4122 gnd.n2204 585
R1526 gnd.n4122 gnd.n4121 585
R1527 gnd.n4095 gnd.n2205 585
R1528 gnd.n2215 gnd.n2205 585
R1529 gnd.n4096 gnd.n2214 585
R1530 gnd.n4113 gnd.n2214 585
R1531 gnd.n4098 gnd.n4097 585
R1532 gnd.n4099 gnd.n4098 585
R1533 gnd.n2227 gnd.n2226 585
R1534 gnd.n2226 gnd.n2225 585
R1535 gnd.n4089 gnd.n4088 585
R1536 gnd.n4088 gnd.n4087 585
R1537 gnd.n2230 gnd.n2229 585
R1538 gnd.n2242 gnd.n2230 585
R1539 gnd.n3876 gnd.n2241 585
R1540 gnd.n4077 gnd.n2241 585
R1541 gnd.n3878 gnd.n3877 585
R1542 gnd.n3877 gnd.n2239 585
R1543 gnd.n3879 gnd.n2252 585
R1544 gnd.n4061 gnd.n2252 585
R1545 gnd.n3881 gnd.n3880 585
R1546 gnd.n3880 gnd.n2251 585
R1547 gnd.n3882 gnd.n2261 585
R1548 gnd.n4053 gnd.n2261 585
R1549 gnd.n3884 gnd.n3883 585
R1550 gnd.n3883 gnd.n2259 585
R1551 gnd.n3657 gnd.n3656 585
R1552 gnd.n3658 gnd.n3657 585
R1553 gnd.n2348 gnd.n2347 585
R1554 gnd.n2354 gnd.n2347 585
R1555 gnd.n3632 gnd.n2366 585
R1556 gnd.n2366 gnd.n2353 585
R1557 gnd.n3634 gnd.n3633 585
R1558 gnd.n3635 gnd.n3634 585
R1559 gnd.n2367 gnd.n2365 585
R1560 gnd.n2365 gnd.n2361 585
R1561 gnd.n3366 gnd.n3365 585
R1562 gnd.n3365 gnd.n3364 585
R1563 gnd.n2372 gnd.n2371 585
R1564 gnd.n3335 gnd.n2372 585
R1565 gnd.n3355 gnd.n3354 585
R1566 gnd.n3354 gnd.n3353 585
R1567 gnd.n2379 gnd.n2378 585
R1568 gnd.n3341 gnd.n2379 585
R1569 gnd.n3311 gnd.n2399 585
R1570 gnd.n2399 gnd.n2398 585
R1571 gnd.n3313 gnd.n3312 585
R1572 gnd.n3314 gnd.n3313 585
R1573 gnd.n2400 gnd.n2397 585
R1574 gnd.n2408 gnd.n2397 585
R1575 gnd.n3289 gnd.n2420 585
R1576 gnd.n2420 gnd.n2407 585
R1577 gnd.n3291 gnd.n3290 585
R1578 gnd.n3292 gnd.n3291 585
R1579 gnd.n2421 gnd.n2419 585
R1580 gnd.n2419 gnd.n2415 585
R1581 gnd.n3277 gnd.n3276 585
R1582 gnd.n3276 gnd.n3275 585
R1583 gnd.n2426 gnd.n2425 585
R1584 gnd.n2436 gnd.n2426 585
R1585 gnd.n3266 gnd.n3265 585
R1586 gnd.n3265 gnd.n3264 585
R1587 gnd.n2433 gnd.n2432 585
R1588 gnd.n3252 gnd.n2433 585
R1589 gnd.n3226 gnd.n2454 585
R1590 gnd.n2454 gnd.n2443 585
R1591 gnd.n3228 gnd.n3227 585
R1592 gnd.n3229 gnd.n3228 585
R1593 gnd.n2455 gnd.n2453 585
R1594 gnd.n2463 gnd.n2453 585
R1595 gnd.n3204 gnd.n2475 585
R1596 gnd.n2475 gnd.n2462 585
R1597 gnd.n3206 gnd.n3205 585
R1598 gnd.n3207 gnd.n3206 585
R1599 gnd.n2476 gnd.n2474 585
R1600 gnd.n2474 gnd.n2470 585
R1601 gnd.n3192 gnd.n3191 585
R1602 gnd.n3191 gnd.n3190 585
R1603 gnd.n2481 gnd.n2480 585
R1604 gnd.n2490 gnd.n2481 585
R1605 gnd.n3181 gnd.n3180 585
R1606 gnd.n3180 gnd.n3179 585
R1607 gnd.n2488 gnd.n2487 585
R1608 gnd.n3167 gnd.n2488 585
R1609 gnd.n2605 gnd.n2604 585
R1610 gnd.n2605 gnd.n2497 585
R1611 gnd.n3124 gnd.n3123 585
R1612 gnd.n3123 gnd.n3122 585
R1613 gnd.n3125 gnd.n2599 585
R1614 gnd.n2610 gnd.n2599 585
R1615 gnd.n3127 gnd.n3126 585
R1616 gnd.n3128 gnd.n3127 585
R1617 gnd.n2600 gnd.n2598 585
R1618 gnd.n2623 gnd.n2598 585
R1619 gnd.n2583 gnd.n2582 585
R1620 gnd.n2586 gnd.n2583 585
R1621 gnd.n3138 gnd.n3137 585
R1622 gnd.n3137 gnd.n3136 585
R1623 gnd.n3139 gnd.n2577 585
R1624 gnd.n3098 gnd.n2577 585
R1625 gnd.n3141 gnd.n3140 585
R1626 gnd.n3142 gnd.n3141 585
R1627 gnd.n2578 gnd.n2576 585
R1628 gnd.n2637 gnd.n2576 585
R1629 gnd.n3090 gnd.n3089 585
R1630 gnd.n3089 gnd.n3088 585
R1631 gnd.n2634 gnd.n2633 585
R1632 gnd.n3072 gnd.n2634 585
R1633 gnd.n3059 gnd.n2653 585
R1634 gnd.n2653 gnd.n2652 585
R1635 gnd.n3061 gnd.n3060 585
R1636 gnd.n3062 gnd.n3061 585
R1637 gnd.n2654 gnd.n2651 585
R1638 gnd.n2660 gnd.n2651 585
R1639 gnd.n3040 gnd.n3039 585
R1640 gnd.n3041 gnd.n3040 585
R1641 gnd.n2671 gnd.n2670 585
R1642 gnd.n2670 gnd.n2666 585
R1643 gnd.n3030 gnd.n3029 585
R1644 gnd.n3031 gnd.n3030 585
R1645 gnd.n2681 gnd.n2680 585
R1646 gnd.n2686 gnd.n2680 585
R1647 gnd.n3008 gnd.n2699 585
R1648 gnd.n2699 gnd.n2685 585
R1649 gnd.n3010 gnd.n3009 585
R1650 gnd.n3011 gnd.n3010 585
R1651 gnd.n2700 gnd.n2698 585
R1652 gnd.n2698 gnd.n2694 585
R1653 gnd.n2999 gnd.n2998 585
R1654 gnd.n3000 gnd.n2999 585
R1655 gnd.n2707 gnd.n2706 585
R1656 gnd.n2711 gnd.n2706 585
R1657 gnd.n2976 gnd.n2728 585
R1658 gnd.n2728 gnd.n2710 585
R1659 gnd.n2978 gnd.n2977 585
R1660 gnd.n2979 gnd.n2978 585
R1661 gnd.n2729 gnd.n2727 585
R1662 gnd.n2727 gnd.n2718 585
R1663 gnd.n2971 gnd.n2970 585
R1664 gnd.n2970 gnd.n2969 585
R1665 gnd.n2776 gnd.n2775 585
R1666 gnd.n2777 gnd.n2776 585
R1667 gnd.n2930 gnd.n2929 585
R1668 gnd.n2931 gnd.n2930 585
R1669 gnd.n2786 gnd.n2785 585
R1670 gnd.n2785 gnd.n2784 585
R1671 gnd.n2925 gnd.n2924 585
R1672 gnd.n2924 gnd.n2923 585
R1673 gnd.n2789 gnd.n2788 585
R1674 gnd.n2790 gnd.n2789 585
R1675 gnd.n2914 gnd.n2913 585
R1676 gnd.n2915 gnd.n2914 585
R1677 gnd.n2797 gnd.n2796 585
R1678 gnd.n2906 gnd.n2796 585
R1679 gnd.n2909 gnd.n2908 585
R1680 gnd.n2908 gnd.n2907 585
R1681 gnd.n2800 gnd.n2799 585
R1682 gnd.n2801 gnd.n2800 585
R1683 gnd.n2895 gnd.n2894 585
R1684 gnd.n2893 gnd.n2819 585
R1685 gnd.n2892 gnd.n2818 585
R1686 gnd.n2897 gnd.n2818 585
R1687 gnd.n2891 gnd.n2890 585
R1688 gnd.n2889 gnd.n2888 585
R1689 gnd.n2887 gnd.n2886 585
R1690 gnd.n2885 gnd.n2884 585
R1691 gnd.n2883 gnd.n2882 585
R1692 gnd.n2881 gnd.n2880 585
R1693 gnd.n2879 gnd.n2878 585
R1694 gnd.n2877 gnd.n2876 585
R1695 gnd.n2875 gnd.n2874 585
R1696 gnd.n2873 gnd.n2872 585
R1697 gnd.n2871 gnd.n2870 585
R1698 gnd.n2869 gnd.n2868 585
R1699 gnd.n2867 gnd.n2866 585
R1700 gnd.n2865 gnd.n2864 585
R1701 gnd.n2863 gnd.n2862 585
R1702 gnd.n2861 gnd.n2860 585
R1703 gnd.n2859 gnd.n2858 585
R1704 gnd.n2857 gnd.n2856 585
R1705 gnd.n2855 gnd.n2854 585
R1706 gnd.n2853 gnd.n2852 585
R1707 gnd.n2851 gnd.n2850 585
R1708 gnd.n2849 gnd.n2848 585
R1709 gnd.n2806 gnd.n2805 585
R1710 gnd.n2900 gnd.n2899 585
R1711 gnd.n3661 gnd.n3660 585
R1712 gnd.n3663 gnd.n3662 585
R1713 gnd.n3665 gnd.n3664 585
R1714 gnd.n3667 gnd.n3666 585
R1715 gnd.n3669 gnd.n3668 585
R1716 gnd.n3671 gnd.n3670 585
R1717 gnd.n3673 gnd.n3672 585
R1718 gnd.n3675 gnd.n3674 585
R1719 gnd.n3677 gnd.n3676 585
R1720 gnd.n3679 gnd.n3678 585
R1721 gnd.n3681 gnd.n3680 585
R1722 gnd.n3683 gnd.n3682 585
R1723 gnd.n3685 gnd.n3684 585
R1724 gnd.n3687 gnd.n3686 585
R1725 gnd.n3689 gnd.n3688 585
R1726 gnd.n3691 gnd.n3690 585
R1727 gnd.n3693 gnd.n3692 585
R1728 gnd.n3695 gnd.n3694 585
R1729 gnd.n3697 gnd.n3696 585
R1730 gnd.n3699 gnd.n3698 585
R1731 gnd.n3701 gnd.n3700 585
R1732 gnd.n3703 gnd.n3702 585
R1733 gnd.n3705 gnd.n3704 585
R1734 gnd.n3707 gnd.n3706 585
R1735 gnd.n3709 gnd.n3708 585
R1736 gnd.n3710 gnd.n2315 585
R1737 gnd.n3711 gnd.n2273 585
R1738 gnd.n3749 gnd.n2273 585
R1739 gnd.n3659 gnd.n2345 585
R1740 gnd.n3659 gnd.n3658 585
R1741 gnd.n3328 gnd.n2344 585
R1742 gnd.n2354 gnd.n2344 585
R1743 gnd.n3330 gnd.n3329 585
R1744 gnd.n3329 gnd.n2353 585
R1745 gnd.n3331 gnd.n2363 585
R1746 gnd.n3635 gnd.n2363 585
R1747 gnd.n3333 gnd.n3332 585
R1748 gnd.n3332 gnd.n2361 585
R1749 gnd.n3334 gnd.n2374 585
R1750 gnd.n3364 gnd.n2374 585
R1751 gnd.n3337 gnd.n3336 585
R1752 gnd.n3336 gnd.n3335 585
R1753 gnd.n3338 gnd.n2381 585
R1754 gnd.n3353 gnd.n2381 585
R1755 gnd.n3340 gnd.n3339 585
R1756 gnd.n3341 gnd.n3340 585
R1757 gnd.n2391 gnd.n2390 585
R1758 gnd.n2398 gnd.n2390 585
R1759 gnd.n3316 gnd.n3315 585
R1760 gnd.n3315 gnd.n3314 585
R1761 gnd.n2394 gnd.n2393 585
R1762 gnd.n2408 gnd.n2394 585
R1763 gnd.n3242 gnd.n3241 585
R1764 gnd.n3241 gnd.n2407 585
R1765 gnd.n3243 gnd.n2417 585
R1766 gnd.n3292 gnd.n2417 585
R1767 gnd.n3245 gnd.n3244 585
R1768 gnd.n3244 gnd.n2415 585
R1769 gnd.n3246 gnd.n2428 585
R1770 gnd.n3275 gnd.n2428 585
R1771 gnd.n3248 gnd.n3247 585
R1772 gnd.n3247 gnd.n2436 585
R1773 gnd.n3249 gnd.n2435 585
R1774 gnd.n3264 gnd.n2435 585
R1775 gnd.n3251 gnd.n3250 585
R1776 gnd.n3252 gnd.n3251 585
R1777 gnd.n2447 gnd.n2446 585
R1778 gnd.n2446 gnd.n2443 585
R1779 gnd.n3231 gnd.n3230 585
R1780 gnd.n3230 gnd.n3229 585
R1781 gnd.n2450 gnd.n2449 585
R1782 gnd.n2463 gnd.n2450 585
R1783 gnd.n3155 gnd.n3154 585
R1784 gnd.n3154 gnd.n2462 585
R1785 gnd.n3156 gnd.n2472 585
R1786 gnd.n3207 gnd.n2472 585
R1787 gnd.n3158 gnd.n3157 585
R1788 gnd.n3157 gnd.n2470 585
R1789 gnd.n3159 gnd.n2483 585
R1790 gnd.n3190 gnd.n2483 585
R1791 gnd.n3161 gnd.n3160 585
R1792 gnd.n3160 gnd.n2490 585
R1793 gnd.n3162 gnd.n2489 585
R1794 gnd.n3179 gnd.n2489 585
R1795 gnd.n3164 gnd.n3163 585
R1796 gnd.n3167 gnd.n3164 585
R1797 gnd.n2500 gnd.n2499 585
R1798 gnd.n2499 gnd.n2497 585
R1799 gnd.n2607 gnd.n2606 585
R1800 gnd.n3122 gnd.n2606 585
R1801 gnd.n2609 gnd.n2608 585
R1802 gnd.n2610 gnd.n2609 585
R1803 gnd.n2620 gnd.n2596 585
R1804 gnd.n3128 gnd.n2596 585
R1805 gnd.n2622 gnd.n2621 585
R1806 gnd.n2623 gnd.n2622 585
R1807 gnd.n2619 gnd.n2618 585
R1808 gnd.n2619 gnd.n2586 585
R1809 gnd.n2617 gnd.n2584 585
R1810 gnd.n3136 gnd.n2584 585
R1811 gnd.n2573 gnd.n2571 585
R1812 gnd.n3098 gnd.n2573 585
R1813 gnd.n3144 gnd.n3143 585
R1814 gnd.n3143 gnd.n3142 585
R1815 gnd.n2572 gnd.n2570 585
R1816 gnd.n2637 gnd.n2572 585
R1817 gnd.n3069 gnd.n2636 585
R1818 gnd.n3088 gnd.n2636 585
R1819 gnd.n3071 gnd.n3070 585
R1820 gnd.n3072 gnd.n3071 585
R1821 gnd.n2646 gnd.n2645 585
R1822 gnd.n2652 gnd.n2645 585
R1823 gnd.n3064 gnd.n3063 585
R1824 gnd.n3063 gnd.n3062 585
R1825 gnd.n2649 gnd.n2648 585
R1826 gnd.n2660 gnd.n2649 585
R1827 gnd.n2949 gnd.n2668 585
R1828 gnd.n3041 gnd.n2668 585
R1829 gnd.n2951 gnd.n2950 585
R1830 gnd.n2950 gnd.n2666 585
R1831 gnd.n2952 gnd.n2679 585
R1832 gnd.n3031 gnd.n2679 585
R1833 gnd.n2954 gnd.n2953 585
R1834 gnd.n2954 gnd.n2686 585
R1835 gnd.n2956 gnd.n2955 585
R1836 gnd.n2955 gnd.n2685 585
R1837 gnd.n2957 gnd.n2696 585
R1838 gnd.n3011 gnd.n2696 585
R1839 gnd.n2959 gnd.n2958 585
R1840 gnd.n2958 gnd.n2694 585
R1841 gnd.n2960 gnd.n2705 585
R1842 gnd.n3000 gnd.n2705 585
R1843 gnd.n2962 gnd.n2961 585
R1844 gnd.n2962 gnd.n2711 585
R1845 gnd.n2964 gnd.n2963 585
R1846 gnd.n2963 gnd.n2710 585
R1847 gnd.n2965 gnd.n2726 585
R1848 gnd.n2979 gnd.n2726 585
R1849 gnd.n2966 gnd.n2779 585
R1850 gnd.n2779 gnd.n2718 585
R1851 gnd.n2968 gnd.n2967 585
R1852 gnd.n2969 gnd.n2968 585
R1853 gnd.n2780 gnd.n2778 585
R1854 gnd.n2778 gnd.n2777 585
R1855 gnd.n2933 gnd.n2932 585
R1856 gnd.n2932 gnd.n2931 585
R1857 gnd.n2783 gnd.n2782 585
R1858 gnd.n2784 gnd.n2783 585
R1859 gnd.n2922 gnd.n2921 585
R1860 gnd.n2923 gnd.n2922 585
R1861 gnd.n2792 gnd.n2791 585
R1862 gnd.n2791 gnd.n2790 585
R1863 gnd.n2917 gnd.n2916 585
R1864 gnd.n2916 gnd.n2915 585
R1865 gnd.n2795 gnd.n2794 585
R1866 gnd.n2906 gnd.n2795 585
R1867 gnd.n2905 gnd.n2904 585
R1868 gnd.n2907 gnd.n2905 585
R1869 gnd.n2803 gnd.n2802 585
R1870 gnd.n2802 gnd.n2801 585
R1871 gnd.n7566 gnd.n7565 585
R1872 gnd.n7565 gnd.n7564 585
R1873 gnd.n7567 gnd.n202 585
R1874 gnd.n7413 gnd.n202 585
R1875 gnd.n7569 gnd.n7568 585
R1876 gnd.n7570 gnd.n7569 585
R1877 gnd.n189 gnd.n188 585
R1878 gnd.n192 gnd.n189 585
R1879 gnd.n7578 gnd.n7577 585
R1880 gnd.n7577 gnd.n7576 585
R1881 gnd.n7579 gnd.n184 585
R1882 gnd.n184 gnd.n183 585
R1883 gnd.n7581 gnd.n7580 585
R1884 gnd.n7582 gnd.n7581 585
R1885 gnd.n169 gnd.n168 585
R1886 gnd.n173 gnd.n169 585
R1887 gnd.n7590 gnd.n7589 585
R1888 gnd.n7589 gnd.n7588 585
R1889 gnd.n7591 gnd.n164 585
R1890 gnd.n170 gnd.n164 585
R1891 gnd.n7593 gnd.n7592 585
R1892 gnd.n7594 gnd.n7593 585
R1893 gnd.n151 gnd.n150 585
R1894 gnd.n161 gnd.n151 585
R1895 gnd.n7602 gnd.n7601 585
R1896 gnd.n7601 gnd.n7600 585
R1897 gnd.n7603 gnd.n146 585
R1898 gnd.n146 gnd.n145 585
R1899 gnd.n7605 gnd.n7604 585
R1900 gnd.n7606 gnd.n7605 585
R1901 gnd.n131 gnd.n130 585
R1902 gnd.n7385 gnd.n131 585
R1903 gnd.n7614 gnd.n7613 585
R1904 gnd.n7613 gnd.n7612 585
R1905 gnd.n7615 gnd.n126 585
R1906 gnd.n132 gnd.n126 585
R1907 gnd.n7617 gnd.n7616 585
R1908 gnd.n7618 gnd.n7617 585
R1909 gnd.n113 gnd.n112 585
R1910 gnd.n7343 gnd.n113 585
R1911 gnd.n7626 gnd.n7625 585
R1912 gnd.n7625 gnd.n7624 585
R1913 gnd.n7627 gnd.n107 585
R1914 gnd.n7333 gnd.n107 585
R1915 gnd.n7629 gnd.n7628 585
R1916 gnd.n7630 gnd.n7629 585
R1917 gnd.n108 gnd.n106 585
R1918 gnd.n7324 gnd.n106 585
R1919 gnd.n7319 gnd.n7318 585
R1920 gnd.n7318 gnd.n7317 585
R1921 gnd.n7316 gnd.n88 585
R1922 gnd.n7638 gnd.n88 585
R1923 gnd.n7315 gnd.n7314 585
R1924 gnd.n7314 gnd.n7313 585
R1925 gnd.n368 gnd.n366 585
R1926 gnd.n7300 gnd.n368 585
R1927 gnd.n7306 gnd.n7305 585
R1928 gnd.n7305 gnd.n7304 585
R1929 gnd.n374 gnd.n373 585
R1930 gnd.n1460 gnd.n374 585
R1931 gnd.n6053 gnd.n1453 585
R1932 gnd.n6049 gnd.n1453 585
R1933 gnd.n6055 gnd.n6054 585
R1934 gnd.n6056 gnd.n6055 585
R1935 gnd.n1441 gnd.n1440 585
R1936 gnd.n6021 gnd.n1441 585
R1937 gnd.n6064 gnd.n6063 585
R1938 gnd.n6063 gnd.n6062 585
R1939 gnd.n6065 gnd.n1436 585
R1940 gnd.n6037 gnd.n1436 585
R1941 gnd.n6067 gnd.n6066 585
R1942 gnd.n6068 gnd.n6067 585
R1943 gnd.n1420 gnd.n1419 585
R1944 gnd.n6012 gnd.n1420 585
R1945 gnd.n6076 gnd.n6075 585
R1946 gnd.n6075 gnd.n6074 585
R1947 gnd.n6077 gnd.n1415 585
R1948 gnd.n6004 gnd.n1415 585
R1949 gnd.n6079 gnd.n6078 585
R1950 gnd.n6080 gnd.n6079 585
R1951 gnd.n1401 gnd.n1400 585
R1952 gnd.n5998 gnd.n1401 585
R1953 gnd.n6088 gnd.n6087 585
R1954 gnd.n6087 gnd.n6086 585
R1955 gnd.n6089 gnd.n1396 585
R1956 gnd.n5990 gnd.n1396 585
R1957 gnd.n6091 gnd.n6090 585
R1958 gnd.n6092 gnd.n6091 585
R1959 gnd.n1380 gnd.n1379 585
R1960 gnd.n5928 gnd.n1380 585
R1961 gnd.n6100 gnd.n6099 585
R1962 gnd.n6099 gnd.n6098 585
R1963 gnd.n6101 gnd.n1375 585
R1964 gnd.n5936 gnd.n1375 585
R1965 gnd.n6103 gnd.n6102 585
R1966 gnd.n6104 gnd.n6103 585
R1967 gnd.n1360 gnd.n1359 585
R1968 gnd.n5917 gnd.n1360 585
R1969 gnd.n6112 gnd.n6111 585
R1970 gnd.n6111 gnd.n6110 585
R1971 gnd.n6113 gnd.n1354 585
R1972 gnd.n5909 gnd.n1354 585
R1973 gnd.n6115 gnd.n6114 585
R1974 gnd.n6116 gnd.n6115 585
R1975 gnd.n1355 gnd.n1353 585
R1976 gnd.n5361 gnd.n1353 585
R1977 gnd.n5902 gnd.n1341 585
R1978 gnd.n6122 gnd.n1341 585
R1979 gnd.n5447 gnd.n5446 585
R1980 gnd.n5411 gnd.n5410 585
R1981 gnd.n5461 gnd.n5460 585
R1982 gnd.n5463 gnd.n5409 585
R1983 gnd.n5466 gnd.n5465 585
R1984 gnd.n5402 gnd.n5401 585
R1985 gnd.n5480 gnd.n5479 585
R1986 gnd.n5482 gnd.n5400 585
R1987 gnd.n5485 gnd.n5484 585
R1988 gnd.n5393 gnd.n5392 585
R1989 gnd.n5499 gnd.n5498 585
R1990 gnd.n5501 gnd.n5391 585
R1991 gnd.n5504 gnd.n5503 585
R1992 gnd.n5384 gnd.n5383 585
R1993 gnd.n5519 gnd.n5518 585
R1994 gnd.n5521 gnd.n5382 585
R1995 gnd.n5524 gnd.n5523 585
R1996 gnd.n5525 gnd.n5379 585
R1997 gnd.n5378 gnd.n5377 585
R1998 gnd.n5378 gnd.n1329 585
R1999 gnd.n347 gnd.n346 585
R2000 gnd.n7420 gnd.n342 585
R2001 gnd.n7422 gnd.n7421 585
R2002 gnd.n7424 gnd.n340 585
R2003 gnd.n7426 gnd.n7425 585
R2004 gnd.n7427 gnd.n335 585
R2005 gnd.n7429 gnd.n7428 585
R2006 gnd.n7431 gnd.n333 585
R2007 gnd.n7433 gnd.n7432 585
R2008 gnd.n7434 gnd.n328 585
R2009 gnd.n7436 gnd.n7435 585
R2010 gnd.n7438 gnd.n326 585
R2011 gnd.n7440 gnd.n7439 585
R2012 gnd.n7441 gnd.n321 585
R2013 gnd.n7443 gnd.n7442 585
R2014 gnd.n7445 gnd.n319 585
R2015 gnd.n7447 gnd.n7446 585
R2016 gnd.n7448 gnd.n317 585
R2017 gnd.n7449 gnd.n206 585
R2018 gnd.n210 gnd.n206 585
R2019 gnd.n7416 gnd.n209 585
R2020 gnd.n7564 gnd.n209 585
R2021 gnd.n7415 gnd.n7414 585
R2022 gnd.n7414 gnd.n7413 585
R2023 gnd.n351 gnd.n201 585
R2024 gnd.n7570 gnd.n201 585
R2025 gnd.n7366 gnd.n7365 585
R2026 gnd.n7365 gnd.n192 585
R2027 gnd.n7367 gnd.n191 585
R2028 gnd.n7576 gnd.n191 585
R2029 gnd.n7369 gnd.n7368 585
R2030 gnd.n7368 gnd.n183 585
R2031 gnd.n7370 gnd.n182 585
R2032 gnd.n7582 gnd.n182 585
R2033 gnd.n7372 gnd.n7371 585
R2034 gnd.n7371 gnd.n173 585
R2035 gnd.n7373 gnd.n172 585
R2036 gnd.n7588 gnd.n172 585
R2037 gnd.n7375 gnd.n7374 585
R2038 gnd.n7374 gnd.n170 585
R2039 gnd.n7376 gnd.n163 585
R2040 gnd.n7594 gnd.n163 585
R2041 gnd.n7378 gnd.n7377 585
R2042 gnd.n7377 gnd.n161 585
R2043 gnd.n7379 gnd.n153 585
R2044 gnd.n7600 gnd.n153 585
R2045 gnd.n7381 gnd.n7380 585
R2046 gnd.n7380 gnd.n145 585
R2047 gnd.n7382 gnd.n144 585
R2048 gnd.n7606 gnd.n144 585
R2049 gnd.n7384 gnd.n7383 585
R2050 gnd.n7385 gnd.n7384 585
R2051 gnd.n354 gnd.n134 585
R2052 gnd.n7612 gnd.n134 585
R2053 gnd.n7348 gnd.n7347 585
R2054 gnd.n7347 gnd.n132 585
R2055 gnd.n7346 gnd.n125 585
R2056 gnd.n7618 gnd.n125 585
R2057 gnd.n7345 gnd.n7344 585
R2058 gnd.n7344 gnd.n7343 585
R2059 gnd.n356 gnd.n116 585
R2060 gnd.n7624 gnd.n116 585
R2061 gnd.n7332 gnd.n7331 585
R2062 gnd.n7333 gnd.n7332 585
R2063 gnd.n360 gnd.n104 585
R2064 gnd.n7630 gnd.n104 585
R2065 gnd.n7326 gnd.n7325 585
R2066 gnd.n7325 gnd.n7324 585
R2067 gnd.n84 gnd.n83 585
R2068 gnd.n7317 gnd.n84 585
R2069 gnd.n7640 gnd.n7639 585
R2070 gnd.n7639 gnd.n7638 585
R2071 gnd.n7641 gnd.n82 585
R2072 gnd.n7313 gnd.n82 585
R2073 gnd.n7299 gnd.n81 585
R2074 gnd.n7300 gnd.n7299 585
R2075 gnd.n6025 gnd.n377 585
R2076 gnd.n7304 gnd.n377 585
R2077 gnd.n6024 gnd.n6023 585
R2078 gnd.n6023 gnd.n1460 585
R2079 gnd.n6029 gnd.n1459 585
R2080 gnd.n6049 gnd.n1459 585
R2081 gnd.n6030 gnd.n1452 585
R2082 gnd.n6056 gnd.n1452 585
R2083 gnd.n6031 gnd.n6022 585
R2084 gnd.n6022 gnd.n6021 585
R2085 gnd.n1467 gnd.n1443 585
R2086 gnd.n6062 gnd.n1443 585
R2087 gnd.n6036 gnd.n6035 585
R2088 gnd.n6037 gnd.n6036 585
R2089 gnd.n1466 gnd.n1434 585
R2090 gnd.n6068 gnd.n1434 585
R2091 gnd.n6011 gnd.n6010 585
R2092 gnd.n6012 gnd.n6011 585
R2093 gnd.n1472 gnd.n1423 585
R2094 gnd.n6074 gnd.n1423 585
R2095 gnd.n6006 gnd.n6005 585
R2096 gnd.n6005 gnd.n6004 585
R2097 gnd.n1474 gnd.n1414 585
R2098 gnd.n6080 gnd.n1414 585
R2099 gnd.n5997 gnd.n5996 585
R2100 gnd.n5998 gnd.n5997 585
R2101 gnd.n1478 gnd.n1403 585
R2102 gnd.n6086 gnd.n1403 585
R2103 gnd.n5992 gnd.n5991 585
R2104 gnd.n5991 gnd.n5990 585
R2105 gnd.n1480 gnd.n1394 585
R2106 gnd.n6092 gnd.n1394 585
R2107 gnd.n5930 gnd.n5929 585
R2108 gnd.n5929 gnd.n5928 585
R2109 gnd.n1489 gnd.n1383 585
R2110 gnd.n6098 gnd.n1383 585
R2111 gnd.n5935 gnd.n5934 585
R2112 gnd.n5936 gnd.n5935 585
R2113 gnd.n1488 gnd.n1374 585
R2114 gnd.n6104 gnd.n1374 585
R2115 gnd.n5916 gnd.n5915 585
R2116 gnd.n5917 gnd.n5916 585
R2117 gnd.n1493 gnd.n1363 585
R2118 gnd.n6110 gnd.n1363 585
R2119 gnd.n5911 gnd.n5910 585
R2120 gnd.n5910 gnd.n5909 585
R2121 gnd.n1495 gnd.n1351 585
R2122 gnd.n6116 gnd.n1351 585
R2123 gnd.n5363 gnd.n5362 585
R2124 gnd.n5362 gnd.n5361 585
R2125 gnd.n5364 gnd.n1339 585
R2126 gnd.n6122 gnd.n1339 585
R2127 gnd.n3644 gnd.n2295 585
R2128 gnd.n2295 gnd.n2272 585
R2129 gnd.n3645 gnd.n2356 585
R2130 gnd.n2356 gnd.n2346 585
R2131 gnd.n3647 gnd.n3646 585
R2132 gnd.n3648 gnd.n3647 585
R2133 gnd.n2357 gnd.n2355 585
R2134 gnd.n2364 gnd.n2355 585
R2135 gnd.n3638 gnd.n3637 585
R2136 gnd.n3637 gnd.n3636 585
R2137 gnd.n2360 gnd.n2359 585
R2138 gnd.n3363 gnd.n2360 585
R2139 gnd.n3349 gnd.n2383 585
R2140 gnd.n2383 gnd.n2373 585
R2141 gnd.n3351 gnd.n3350 585
R2142 gnd.n3352 gnd.n3351 585
R2143 gnd.n2384 gnd.n2382 585
R2144 gnd.n2382 gnd.n2380 585
R2145 gnd.n3344 gnd.n3343 585
R2146 gnd.n3343 gnd.n3342 585
R2147 gnd.n2387 gnd.n2386 585
R2148 gnd.n2396 gnd.n2387 585
R2149 gnd.n3300 gnd.n2410 585
R2150 gnd.n2410 gnd.n2395 585
R2151 gnd.n3302 gnd.n3301 585
R2152 gnd.n3303 gnd.n3302 585
R2153 gnd.n2411 gnd.n2409 585
R2154 gnd.n2418 gnd.n2409 585
R2155 gnd.n3295 gnd.n3294 585
R2156 gnd.n3294 gnd.n3293 585
R2157 gnd.n2414 gnd.n2413 585
R2158 gnd.n3274 gnd.n2414 585
R2159 gnd.n3260 gnd.n2438 585
R2160 gnd.n2438 gnd.n2427 585
R2161 gnd.n3262 gnd.n3261 585
R2162 gnd.n3263 gnd.n3262 585
R2163 gnd.n2439 gnd.n2437 585
R2164 gnd.n2437 gnd.n2434 585
R2165 gnd.n3255 gnd.n3254 585
R2166 gnd.n3254 gnd.n3253 585
R2167 gnd.n2442 gnd.n2441 585
R2168 gnd.n2452 gnd.n2442 585
R2169 gnd.n3215 gnd.n2465 585
R2170 gnd.n2465 gnd.n2451 585
R2171 gnd.n3217 gnd.n3216 585
R2172 gnd.n3218 gnd.n3217 585
R2173 gnd.n2466 gnd.n2464 585
R2174 gnd.n2473 gnd.n2464 585
R2175 gnd.n3210 gnd.n3209 585
R2176 gnd.n3209 gnd.n3208 585
R2177 gnd.n2469 gnd.n2468 585
R2178 gnd.n3189 gnd.n2469 585
R2179 gnd.n3175 gnd.n2492 585
R2180 gnd.n2492 gnd.n2482 585
R2181 gnd.n3177 gnd.n3176 585
R2182 gnd.n3178 gnd.n3177 585
R2183 gnd.n2493 gnd.n2491 585
R2184 gnd.n3166 gnd.n2491 585
R2185 gnd.n3170 gnd.n3169 585
R2186 gnd.n3169 gnd.n3168 585
R2187 gnd.n2496 gnd.n2495 585
R2188 gnd.n3121 gnd.n2496 585
R2189 gnd.n2614 gnd.n2613 585
R2190 gnd.n2615 gnd.n2614 585
R2191 gnd.n2594 gnd.n2593 585
R2192 gnd.n2597 gnd.n2594 585
R2193 gnd.n3131 gnd.n3130 585
R2194 gnd.n3130 gnd.n3129 585
R2195 gnd.n3132 gnd.n2588 585
R2196 gnd.n2624 gnd.n2588 585
R2197 gnd.n3134 gnd.n3133 585
R2198 gnd.n3135 gnd.n3134 585
R2199 gnd.n2589 gnd.n2587 585
R2200 gnd.n3099 gnd.n2587 585
R2201 gnd.n3083 gnd.n3082 585
R2202 gnd.n3082 gnd.n2575 585
R2203 gnd.n3084 gnd.n2639 585
R2204 gnd.n2639 gnd.n2574 585
R2205 gnd.n3086 gnd.n3085 585
R2206 gnd.n3087 gnd.n3086 585
R2207 gnd.n2640 gnd.n2638 585
R2208 gnd.n2638 gnd.n2635 585
R2209 gnd.n3075 gnd.n3074 585
R2210 gnd.n3074 gnd.n3073 585
R2211 gnd.n2643 gnd.n2642 585
R2212 gnd.n2650 gnd.n2643 585
R2213 gnd.n3049 gnd.n3048 585
R2214 gnd.n3050 gnd.n3049 585
R2215 gnd.n2662 gnd.n2661 585
R2216 gnd.n2669 gnd.n2661 585
R2217 gnd.n3044 gnd.n3043 585
R2218 gnd.n3043 gnd.n3042 585
R2219 gnd.n2665 gnd.n2664 585
R2220 gnd.n3032 gnd.n2665 585
R2221 gnd.n3019 gnd.n2689 585
R2222 gnd.n2689 gnd.n2688 585
R2223 gnd.n3021 gnd.n3020 585
R2224 gnd.n3022 gnd.n3021 585
R2225 gnd.n2690 gnd.n2687 585
R2226 gnd.n2697 gnd.n2687 585
R2227 gnd.n3014 gnd.n3013 585
R2228 gnd.n3013 gnd.n3012 585
R2229 gnd.n2693 gnd.n2692 585
R2230 gnd.n3001 gnd.n2693 585
R2231 gnd.n2988 gnd.n2714 585
R2232 gnd.n2714 gnd.n2713 585
R2233 gnd.n2990 gnd.n2989 585
R2234 gnd.n2991 gnd.n2990 585
R2235 gnd.n2984 gnd.n2712 585
R2236 gnd.n2983 gnd.n2982 585
R2237 gnd.n2717 gnd.n2716 585
R2238 gnd.n2980 gnd.n2717 585
R2239 gnd.n2739 gnd.n2738 585
R2240 gnd.n2742 gnd.n2741 585
R2241 gnd.n2740 gnd.n2735 585
R2242 gnd.n2747 gnd.n2746 585
R2243 gnd.n2749 gnd.n2748 585
R2244 gnd.n2752 gnd.n2751 585
R2245 gnd.n2750 gnd.n2733 585
R2246 gnd.n2757 gnd.n2756 585
R2247 gnd.n2759 gnd.n2758 585
R2248 gnd.n2762 gnd.n2761 585
R2249 gnd.n2760 gnd.n2731 585
R2250 gnd.n2767 gnd.n2766 585
R2251 gnd.n2771 gnd.n2768 585
R2252 gnd.n2772 gnd.n2709 585
R2253 gnd.n3650 gnd.n2310 585
R2254 gnd.n3717 gnd.n3716 585
R2255 gnd.n3719 gnd.n3718 585
R2256 gnd.n3721 gnd.n3720 585
R2257 gnd.n3723 gnd.n3722 585
R2258 gnd.n3725 gnd.n3724 585
R2259 gnd.n3727 gnd.n3726 585
R2260 gnd.n3729 gnd.n3728 585
R2261 gnd.n3731 gnd.n3730 585
R2262 gnd.n3733 gnd.n3732 585
R2263 gnd.n3735 gnd.n3734 585
R2264 gnd.n3737 gnd.n3736 585
R2265 gnd.n3739 gnd.n3738 585
R2266 gnd.n3742 gnd.n3741 585
R2267 gnd.n3740 gnd.n2298 585
R2268 gnd.n3746 gnd.n2296 585
R2269 gnd.n3748 gnd.n3747 585
R2270 gnd.n3749 gnd.n3748 585
R2271 gnd.n3651 gnd.n2351 585
R2272 gnd.n3651 gnd.n2272 585
R2273 gnd.n3653 gnd.n3652 585
R2274 gnd.n3652 gnd.n2346 585
R2275 gnd.n3649 gnd.n2350 585
R2276 gnd.n3649 gnd.n3648 585
R2277 gnd.n3628 gnd.n2352 585
R2278 gnd.n2364 gnd.n2352 585
R2279 gnd.n3627 gnd.n2362 585
R2280 gnd.n3636 gnd.n2362 585
R2281 gnd.n3362 gnd.n2369 585
R2282 gnd.n3363 gnd.n3362 585
R2283 gnd.n3361 gnd.n3360 585
R2284 gnd.n3361 gnd.n2373 585
R2285 gnd.n3359 gnd.n2375 585
R2286 gnd.n3352 gnd.n2375 585
R2287 gnd.n2388 gnd.n2376 585
R2288 gnd.n2388 gnd.n2380 585
R2289 gnd.n3308 gnd.n2389 585
R2290 gnd.n3342 gnd.n2389 585
R2291 gnd.n3307 gnd.n3306 585
R2292 gnd.n3306 gnd.n2396 585
R2293 gnd.n3305 gnd.n2404 585
R2294 gnd.n3305 gnd.n2395 585
R2295 gnd.n3304 gnd.n2406 585
R2296 gnd.n3304 gnd.n3303 585
R2297 gnd.n3283 gnd.n2405 585
R2298 gnd.n2418 gnd.n2405 585
R2299 gnd.n3282 gnd.n2416 585
R2300 gnd.n3293 gnd.n2416 585
R2301 gnd.n3273 gnd.n2423 585
R2302 gnd.n3274 gnd.n3273 585
R2303 gnd.n3272 gnd.n3271 585
R2304 gnd.n3272 gnd.n2427 585
R2305 gnd.n3270 gnd.n2429 585
R2306 gnd.n3263 gnd.n2429 585
R2307 gnd.n2444 gnd.n2430 585
R2308 gnd.n2444 gnd.n2434 585
R2309 gnd.n3223 gnd.n2445 585
R2310 gnd.n3253 gnd.n2445 585
R2311 gnd.n3222 gnd.n3221 585
R2312 gnd.n3221 gnd.n2452 585
R2313 gnd.n3220 gnd.n2459 585
R2314 gnd.n3220 gnd.n2451 585
R2315 gnd.n3219 gnd.n2461 585
R2316 gnd.n3219 gnd.n3218 585
R2317 gnd.n3198 gnd.n2460 585
R2318 gnd.n2473 gnd.n2460 585
R2319 gnd.n3197 gnd.n2471 585
R2320 gnd.n3208 gnd.n2471 585
R2321 gnd.n3188 gnd.n2478 585
R2322 gnd.n3189 gnd.n3188 585
R2323 gnd.n3187 gnd.n3186 585
R2324 gnd.n3187 gnd.n2482 585
R2325 gnd.n3185 gnd.n2484 585
R2326 gnd.n3178 gnd.n2484 585
R2327 gnd.n3165 gnd.n2485 585
R2328 gnd.n3166 gnd.n3165 585
R2329 gnd.n3118 gnd.n2498 585
R2330 gnd.n3168 gnd.n2498 585
R2331 gnd.n3120 gnd.n3119 585
R2332 gnd.n3121 gnd.n3120 585
R2333 gnd.n3113 gnd.n2616 585
R2334 gnd.n2616 gnd.n2615 585
R2335 gnd.n3111 gnd.n3110 585
R2336 gnd.n3110 gnd.n2597 585
R2337 gnd.n3108 gnd.n2595 585
R2338 gnd.n3129 gnd.n2595 585
R2339 gnd.n2626 gnd.n2625 585
R2340 gnd.n2625 gnd.n2624 585
R2341 gnd.n3102 gnd.n2585 585
R2342 gnd.n3135 gnd.n2585 585
R2343 gnd.n3101 gnd.n3100 585
R2344 gnd.n3100 gnd.n3099 585
R2345 gnd.n3097 gnd.n2628 585
R2346 gnd.n3097 gnd.n2575 585
R2347 gnd.n3096 gnd.n3095 585
R2348 gnd.n3096 gnd.n2574 585
R2349 gnd.n2631 gnd.n2630 585
R2350 gnd.n3087 gnd.n2630 585
R2351 gnd.n3055 gnd.n3054 585
R2352 gnd.n3054 gnd.n2635 585
R2353 gnd.n3056 gnd.n2644 585
R2354 gnd.n3073 gnd.n2644 585
R2355 gnd.n3053 gnd.n3052 585
R2356 gnd.n3052 gnd.n2650 585
R2357 gnd.n3051 gnd.n2658 585
R2358 gnd.n3051 gnd.n3050 585
R2359 gnd.n3036 gnd.n2659 585
R2360 gnd.n2669 gnd.n2659 585
R2361 gnd.n3035 gnd.n2667 585
R2362 gnd.n3042 gnd.n2667 585
R2363 gnd.n3034 gnd.n3033 585
R2364 gnd.n3033 gnd.n3032 585
R2365 gnd.n2678 gnd.n2675 585
R2366 gnd.n2688 gnd.n2678 585
R2367 gnd.n3024 gnd.n3023 585
R2368 gnd.n3023 gnd.n3022 585
R2369 gnd.n2684 gnd.n2683 585
R2370 gnd.n2697 gnd.n2684 585
R2371 gnd.n3004 gnd.n2695 585
R2372 gnd.n3012 gnd.n2695 585
R2373 gnd.n3003 gnd.n3002 585
R2374 gnd.n3002 gnd.n3001 585
R2375 gnd.n2704 gnd.n2702 585
R2376 gnd.n2713 gnd.n2704 585
R2377 gnd.n2993 gnd.n2992 585
R2378 gnd.n2992 gnd.n2991 585
R2379 gnd.n5653 gnd.n5652 585
R2380 gnd.n5654 gnd.n5653 585
R2381 gnd.n5567 gnd.n1574 585
R2382 gnd.n1581 gnd.n1574 585
R2383 gnd.n5566 gnd.n5565 585
R2384 gnd.n5565 gnd.n5564 585
R2385 gnd.n1577 gnd.n1576 585
R2386 gnd.n5335 gnd.n1577 585
R2387 gnd.n5324 gnd.n1624 585
R2388 gnd.n1624 gnd.n1618 585
R2389 gnd.n5326 gnd.n5325 585
R2390 gnd.n5327 gnd.n5326 585
R2391 gnd.n5323 gnd.n1623 585
R2392 gnd.n5317 gnd.n1623 585
R2393 gnd.n5322 gnd.n5321 585
R2394 gnd.n5321 gnd.n5320 585
R2395 gnd.n1626 gnd.n1625 585
R2396 gnd.n5304 gnd.n1626 585
R2397 gnd.n5279 gnd.n5278 585
R2398 gnd.n5278 gnd.n1637 585
R2399 gnd.n5280 gnd.n1646 585
R2400 gnd.n5293 gnd.n1646 585
R2401 gnd.n5281 gnd.n1656 585
R2402 gnd.n1656 gnd.n1645 585
R2403 gnd.n5283 gnd.n5282 585
R2404 gnd.n5284 gnd.n5283 585
R2405 gnd.n5277 gnd.n1655 585
R2406 gnd.n5272 gnd.n1655 585
R2407 gnd.n5276 gnd.n5275 585
R2408 gnd.n5275 gnd.n5274 585
R2409 gnd.n1658 gnd.n1657 585
R2410 gnd.n5259 gnd.n1658 585
R2411 gnd.n5248 gnd.n1673 585
R2412 gnd.n1673 gnd.n1667 585
R2413 gnd.n5250 gnd.n5249 585
R2414 gnd.n5251 gnd.n5250 585
R2415 gnd.n5247 gnd.n1672 585
R2416 gnd.n1679 gnd.n1672 585
R2417 gnd.n5246 gnd.n5245 585
R2418 gnd.n5245 gnd.n5244 585
R2419 gnd.n1675 gnd.n1674 585
R2420 gnd.n5125 gnd.n1675 585
R2421 gnd.n5232 gnd.n5231 585
R2422 gnd.n5233 gnd.n5232 585
R2423 gnd.n5230 gnd.n1691 585
R2424 gnd.n1691 gnd.n1687 585
R2425 gnd.n5229 gnd.n5228 585
R2426 gnd.n5228 gnd.n5227 585
R2427 gnd.n1693 gnd.n1692 585
R2428 gnd.n5135 gnd.n1693 585
R2429 gnd.n5201 gnd.n5200 585
R2430 gnd.n5202 gnd.n5201 585
R2431 gnd.n5199 gnd.n1704 585
R2432 gnd.n1704 gnd.n1701 585
R2433 gnd.n5198 gnd.n5197 585
R2434 gnd.n5197 gnd.n5196 585
R2435 gnd.n1706 gnd.n1705 585
R2436 gnd.n5142 gnd.n1706 585
R2437 gnd.n5182 gnd.n5181 585
R2438 gnd.n5183 gnd.n5182 585
R2439 gnd.n5180 gnd.n1717 585
R2440 gnd.n5175 gnd.n1717 585
R2441 gnd.n5179 gnd.n5178 585
R2442 gnd.n5178 gnd.n5177 585
R2443 gnd.n1719 gnd.n1718 585
R2444 gnd.n1731 gnd.n1719 585
R2445 gnd.n5111 gnd.n5110 585
R2446 gnd.n5111 gnd.n1730 585
R2447 gnd.n5115 gnd.n5114 585
R2448 gnd.n5114 gnd.n5113 585
R2449 gnd.n5116 gnd.n1737 585
R2450 gnd.n5155 gnd.n1737 585
R2451 gnd.n5117 gnd.n1746 585
R2452 gnd.n5041 gnd.n1746 585
R2453 gnd.n5119 gnd.n5118 585
R2454 gnd.n5120 gnd.n5119 585
R2455 gnd.n5109 gnd.n1745 585
R2456 gnd.n5104 gnd.n1745 585
R2457 gnd.n5108 gnd.n5107 585
R2458 gnd.n5107 gnd.n5106 585
R2459 gnd.n1748 gnd.n1747 585
R2460 gnd.n5093 gnd.n1748 585
R2461 gnd.n5083 gnd.n1766 585
R2462 gnd.n1766 gnd.n1757 585
R2463 gnd.n5085 gnd.n5084 585
R2464 gnd.n5086 gnd.n5085 585
R2465 gnd.n5082 gnd.n1765 585
R2466 gnd.n1770 gnd.n1765 585
R2467 gnd.n5081 gnd.n5080 585
R2468 gnd.n5080 gnd.n5079 585
R2469 gnd.n1768 gnd.n1767 585
R2470 gnd.n5033 gnd.n1768 585
R2471 gnd.n5067 gnd.n5066 585
R2472 gnd.n5068 gnd.n5067 585
R2473 gnd.n5065 gnd.n1781 585
R2474 gnd.n1781 gnd.n1777 585
R2475 gnd.n5064 gnd.n5063 585
R2476 gnd.n5063 gnd.n5062 585
R2477 gnd.n1783 gnd.n1782 585
R2478 gnd.n5023 gnd.n1783 585
R2479 gnd.n5008 gnd.n5007 585
R2480 gnd.n5007 gnd.n1793 585
R2481 gnd.n5009 gnd.n1803 585
R2482 gnd.n4992 gnd.n1803 585
R2483 gnd.n5011 gnd.n5010 585
R2484 gnd.n5012 gnd.n5011 585
R2485 gnd.n5006 gnd.n1802 585
R2486 gnd.n1802 gnd.n1799 585
R2487 gnd.n5005 gnd.n5004 585
R2488 gnd.n5004 gnd.n5003 585
R2489 gnd.n1805 gnd.n1804 585
R2490 gnd.n4983 gnd.n1805 585
R2491 gnd.n4968 gnd.n4967 585
R2492 gnd.n4967 gnd.n1816 585
R2493 gnd.n4969 gnd.n1826 585
R2494 gnd.n4956 gnd.n1826 585
R2495 gnd.n4971 gnd.n4970 585
R2496 gnd.n4972 gnd.n4971 585
R2497 gnd.n4966 gnd.n1825 585
R2498 gnd.n1825 gnd.n1822 585
R2499 gnd.n4965 gnd.n4964 585
R2500 gnd.n4964 gnd.n4963 585
R2501 gnd.n1828 gnd.n1827 585
R2502 gnd.n1841 gnd.n1828 585
R2503 gnd.n4941 gnd.n4940 585
R2504 gnd.n4942 gnd.n4941 585
R2505 gnd.n4939 gnd.n1843 585
R2506 gnd.n4934 gnd.n1843 585
R2507 gnd.n4938 gnd.n4937 585
R2508 gnd.n4937 gnd.n4936 585
R2509 gnd.n1845 gnd.n1844 585
R2510 gnd.n4920 gnd.n1845 585
R2511 gnd.n4908 gnd.n1863 585
R2512 gnd.n1863 gnd.n1855 585
R2513 gnd.n4910 gnd.n4909 585
R2514 gnd.n4911 gnd.n4910 585
R2515 gnd.n4907 gnd.n1862 585
R2516 gnd.n4852 gnd.n1862 585
R2517 gnd.n4906 gnd.n4905 585
R2518 gnd.n4905 gnd.n4904 585
R2519 gnd.n1865 gnd.n1864 585
R2520 gnd.n4878 gnd.n1865 585
R2521 gnd.n4891 gnd.n4890 585
R2522 gnd.n4892 gnd.n4891 585
R2523 gnd.n4889 gnd.n1876 585
R2524 gnd.n4884 gnd.n1876 585
R2525 gnd.n4888 gnd.n4887 585
R2526 gnd.n4887 gnd.n4886 585
R2527 gnd.n1878 gnd.n1877 585
R2528 gnd.n4873 gnd.n1878 585
R2529 gnd.n4825 gnd.n4822 585
R2530 gnd.n4825 gnd.n4824 585
R2531 gnd.n4826 gnd.n4821 585
R2532 gnd.n4826 gnd.n1892 585
R2533 gnd.n4828 gnd.n4827 585
R2534 gnd.n4827 gnd.n1891 585
R2535 gnd.n4829 gnd.n1903 585
R2536 gnd.n4809 gnd.n1903 585
R2537 gnd.n4831 gnd.n4830 585
R2538 gnd.n4832 gnd.n4831 585
R2539 gnd.n4820 gnd.n1902 585
R2540 gnd.n4815 gnd.n1902 585
R2541 gnd.n4819 gnd.n4818 585
R2542 gnd.n4818 gnd.n4817 585
R2543 gnd.n1905 gnd.n1904 585
R2544 gnd.n4800 gnd.n1905 585
R2545 gnd.n1928 gnd.n1927 585
R2546 gnd.n4775 gnd.n1928 585
R2547 gnd.n4779 gnd.n4778 585
R2548 gnd.n4778 gnd.n4777 585
R2549 gnd.n4780 gnd.n1917 585
R2550 gnd.n4791 gnd.n1917 585
R2551 gnd.n4781 gnd.n1925 585
R2552 gnd.n1929 gnd.n1925 585
R2553 gnd.n4783 gnd.n4782 585
R2554 gnd.n4784 gnd.n4783 585
R2555 gnd.n1926 gnd.n1924 585
R2556 gnd.n4757 gnd.n1924 585
R2557 gnd.n4750 gnd.n4749 585
R2558 gnd.n4751 gnd.n4750 585
R2559 gnd.n4748 gnd.n1939 585
R2560 gnd.n1939 gnd.n1223 585
R2561 gnd.n4747 gnd.n4746 585
R2562 gnd.n4746 gnd.n1221 585
R2563 gnd.n4745 gnd.n1940 585
R2564 gnd.n4745 gnd.n4744 585
R2565 gnd.n1209 gnd.n1208 585
R2566 gnd.n2020 gnd.n1209 585
R2567 gnd.n6258 gnd.n6257 585
R2568 gnd.n6257 gnd.n6256 585
R2569 gnd.n6259 gnd.n1187 585
R2570 gnd.n2026 gnd.n1187 585
R2571 gnd.n6324 gnd.n6323 585
R2572 gnd.n6322 gnd.n1186 585
R2573 gnd.n6321 gnd.n1185 585
R2574 gnd.n6326 gnd.n1185 585
R2575 gnd.n6320 gnd.n6319 585
R2576 gnd.n6318 gnd.n6317 585
R2577 gnd.n6316 gnd.n6315 585
R2578 gnd.n6314 gnd.n6313 585
R2579 gnd.n6312 gnd.n6311 585
R2580 gnd.n6310 gnd.n6309 585
R2581 gnd.n6308 gnd.n6307 585
R2582 gnd.n6306 gnd.n6305 585
R2583 gnd.n6304 gnd.n6303 585
R2584 gnd.n6302 gnd.n6301 585
R2585 gnd.n6300 gnd.n6299 585
R2586 gnd.n6298 gnd.n6297 585
R2587 gnd.n6296 gnd.n6295 585
R2588 gnd.n6294 gnd.n6293 585
R2589 gnd.n6292 gnd.n6291 585
R2590 gnd.n6290 gnd.n6289 585
R2591 gnd.n6288 gnd.n6287 585
R2592 gnd.n6286 gnd.n6285 585
R2593 gnd.n6284 gnd.n6283 585
R2594 gnd.n6282 gnd.n6281 585
R2595 gnd.n6280 gnd.n6279 585
R2596 gnd.n6278 gnd.n6277 585
R2597 gnd.n6276 gnd.n6275 585
R2598 gnd.n6274 gnd.n6273 585
R2599 gnd.n6272 gnd.n6271 585
R2600 gnd.n6270 gnd.n6269 585
R2601 gnd.n6268 gnd.n6267 585
R2602 gnd.n6266 gnd.n6265 585
R2603 gnd.n6264 gnd.n1149 585
R2604 gnd.n6329 gnd.n6328 585
R2605 gnd.n1151 gnd.n1148 585
R2606 gnd.n1953 gnd.n1952 585
R2607 gnd.n1955 gnd.n1954 585
R2608 gnd.n1958 gnd.n1957 585
R2609 gnd.n1960 gnd.n1959 585
R2610 gnd.n1962 gnd.n1961 585
R2611 gnd.n1964 gnd.n1963 585
R2612 gnd.n1966 gnd.n1965 585
R2613 gnd.n1968 gnd.n1967 585
R2614 gnd.n1970 gnd.n1969 585
R2615 gnd.n1972 gnd.n1971 585
R2616 gnd.n1974 gnd.n1973 585
R2617 gnd.n1976 gnd.n1975 585
R2618 gnd.n1978 gnd.n1977 585
R2619 gnd.n1980 gnd.n1979 585
R2620 gnd.n1982 gnd.n1981 585
R2621 gnd.n1984 gnd.n1983 585
R2622 gnd.n1986 gnd.n1985 585
R2623 gnd.n1988 gnd.n1987 585
R2624 gnd.n1990 gnd.n1989 585
R2625 gnd.n1992 gnd.n1991 585
R2626 gnd.n1994 gnd.n1993 585
R2627 gnd.n1996 gnd.n1995 585
R2628 gnd.n1998 gnd.n1997 585
R2629 gnd.n2000 gnd.n1999 585
R2630 gnd.n2002 gnd.n2001 585
R2631 gnd.n2004 gnd.n2003 585
R2632 gnd.n2006 gnd.n2005 585
R2633 gnd.n2008 gnd.n2007 585
R2634 gnd.n2010 gnd.n2009 585
R2635 gnd.n2012 gnd.n2011 585
R2636 gnd.n2013 gnd.n1949 585
R2637 gnd.n5657 gnd.n5656 585
R2638 gnd.n5659 gnd.n5658 585
R2639 gnd.n5661 gnd.n5660 585
R2640 gnd.n5663 gnd.n5662 585
R2641 gnd.n5665 gnd.n5664 585
R2642 gnd.n5667 gnd.n5666 585
R2643 gnd.n5669 gnd.n5668 585
R2644 gnd.n5671 gnd.n5670 585
R2645 gnd.n5673 gnd.n5672 585
R2646 gnd.n5675 gnd.n5674 585
R2647 gnd.n5677 gnd.n5676 585
R2648 gnd.n5679 gnd.n5678 585
R2649 gnd.n5681 gnd.n5680 585
R2650 gnd.n5683 gnd.n5682 585
R2651 gnd.n5685 gnd.n5684 585
R2652 gnd.n5687 gnd.n5686 585
R2653 gnd.n5689 gnd.n5688 585
R2654 gnd.n5691 gnd.n5690 585
R2655 gnd.n5693 gnd.n5692 585
R2656 gnd.n5695 gnd.n5694 585
R2657 gnd.n5697 gnd.n5696 585
R2658 gnd.n5699 gnd.n5698 585
R2659 gnd.n5701 gnd.n5700 585
R2660 gnd.n5703 gnd.n5702 585
R2661 gnd.n5705 gnd.n5704 585
R2662 gnd.n5707 gnd.n5706 585
R2663 gnd.n5709 gnd.n5708 585
R2664 gnd.n5711 gnd.n5710 585
R2665 gnd.n5713 gnd.n5712 585
R2666 gnd.n5715 gnd.n1568 585
R2667 gnd.n5717 gnd.n5716 585
R2668 gnd.n5719 gnd.n1532 585
R2669 gnd.n5721 gnd.n5720 585
R2670 gnd.n5724 gnd.n5723 585
R2671 gnd.n1535 gnd.n1533 585
R2672 gnd.n5590 gnd.n5589 585
R2673 gnd.n5592 gnd.n5591 585
R2674 gnd.n5595 gnd.n5594 585
R2675 gnd.n5597 gnd.n5596 585
R2676 gnd.n5599 gnd.n5598 585
R2677 gnd.n5601 gnd.n5600 585
R2678 gnd.n5603 gnd.n5602 585
R2679 gnd.n5605 gnd.n5604 585
R2680 gnd.n5607 gnd.n5606 585
R2681 gnd.n5609 gnd.n5608 585
R2682 gnd.n5611 gnd.n5610 585
R2683 gnd.n5613 gnd.n5612 585
R2684 gnd.n5615 gnd.n5614 585
R2685 gnd.n5617 gnd.n5616 585
R2686 gnd.n5619 gnd.n5618 585
R2687 gnd.n5621 gnd.n5620 585
R2688 gnd.n5623 gnd.n5622 585
R2689 gnd.n5625 gnd.n5624 585
R2690 gnd.n5627 gnd.n5626 585
R2691 gnd.n5629 gnd.n5628 585
R2692 gnd.n5631 gnd.n5630 585
R2693 gnd.n5633 gnd.n5632 585
R2694 gnd.n5635 gnd.n5634 585
R2695 gnd.n5637 gnd.n5636 585
R2696 gnd.n5639 gnd.n5638 585
R2697 gnd.n5641 gnd.n5640 585
R2698 gnd.n5643 gnd.n5642 585
R2699 gnd.n5645 gnd.n5644 585
R2700 gnd.n5647 gnd.n5646 585
R2701 gnd.n5649 gnd.n5648 585
R2702 gnd.n5650 gnd.n1575 585
R2703 gnd.n5655 gnd.n1571 585
R2704 gnd.n5655 gnd.n5654 585
R2705 gnd.n5331 gnd.n1572 585
R2706 gnd.n1581 gnd.n1572 585
R2707 gnd.n5332 gnd.n1579 585
R2708 gnd.n5564 gnd.n1579 585
R2709 gnd.n5334 gnd.n5333 585
R2710 gnd.n5335 gnd.n5334 585
R2711 gnd.n5330 gnd.n1619 585
R2712 gnd.n1619 gnd.n1618 585
R2713 gnd.n5329 gnd.n5328 585
R2714 gnd.n5328 gnd.n5327 585
R2715 gnd.n1621 gnd.n1620 585
R2716 gnd.n5317 gnd.n1621 585
R2717 gnd.n5288 gnd.n1628 585
R2718 gnd.n5320 gnd.n1628 585
R2719 gnd.n5289 gnd.n1638 585
R2720 gnd.n5304 gnd.n1638 585
R2721 gnd.n5290 gnd.n1649 585
R2722 gnd.n1649 gnd.n1637 585
R2723 gnd.n5292 gnd.n5291 585
R2724 gnd.n5293 gnd.n5292 585
R2725 gnd.n5287 gnd.n1648 585
R2726 gnd.n1648 gnd.n1645 585
R2727 gnd.n5286 gnd.n5285 585
R2728 gnd.n5285 gnd.n5284 585
R2729 gnd.n1651 gnd.n1650 585
R2730 gnd.n5272 gnd.n1651 585
R2731 gnd.n5255 gnd.n1659 585
R2732 gnd.n5274 gnd.n1659 585
R2733 gnd.n5257 gnd.n5256 585
R2734 gnd.n5259 gnd.n5257 585
R2735 gnd.n5254 gnd.n1669 585
R2736 gnd.n1669 gnd.n1667 585
R2737 gnd.n5253 gnd.n5252 585
R2738 gnd.n5252 gnd.n5251 585
R2739 gnd.n1671 gnd.n1670 585
R2740 gnd.n1679 gnd.n1671 585
R2741 gnd.n5124 gnd.n1677 585
R2742 gnd.n5244 gnd.n1677 585
R2743 gnd.n5127 gnd.n5126 585
R2744 gnd.n5126 gnd.n5125 585
R2745 gnd.n5128 gnd.n1689 585
R2746 gnd.n5233 gnd.n1689 585
R2747 gnd.n5130 gnd.n5129 585
R2748 gnd.n5129 gnd.n1687 585
R2749 gnd.n5131 gnd.n1694 585
R2750 gnd.n5227 gnd.n1694 585
R2751 gnd.n5137 gnd.n5136 585
R2752 gnd.n5136 gnd.n5135 585
R2753 gnd.n5138 gnd.n1702 585
R2754 gnd.n5202 gnd.n1702 585
R2755 gnd.n5140 gnd.n5139 585
R2756 gnd.n5139 gnd.n1701 585
R2757 gnd.n5141 gnd.n1708 585
R2758 gnd.n5196 gnd.n1708 585
R2759 gnd.n5144 gnd.n5143 585
R2760 gnd.n5143 gnd.n5142 585
R2761 gnd.n5145 gnd.n1715 585
R2762 gnd.n5183 gnd.n1715 585
R2763 gnd.n5146 gnd.n1722 585
R2764 gnd.n5175 gnd.n1722 585
R2765 gnd.n5147 gnd.n1721 585
R2766 gnd.n5177 gnd.n1721 585
R2767 gnd.n5149 gnd.n5148 585
R2768 gnd.n5149 gnd.n1731 585
R2769 gnd.n5151 gnd.n5150 585
R2770 gnd.n5150 gnd.n1730 585
R2771 gnd.n5152 gnd.n1740 585
R2772 gnd.n5113 gnd.n1740 585
R2773 gnd.n5154 gnd.n5153 585
R2774 gnd.n5155 gnd.n5154 585
R2775 gnd.n5123 gnd.n1739 585
R2776 gnd.n5041 gnd.n1739 585
R2777 gnd.n5122 gnd.n5121 585
R2778 gnd.n5121 gnd.n5120 585
R2779 gnd.n1742 gnd.n1741 585
R2780 gnd.n5104 gnd.n1742 585
R2781 gnd.n5090 gnd.n1750 585
R2782 gnd.n5106 gnd.n1750 585
R2783 gnd.n5092 gnd.n5091 585
R2784 gnd.n5093 gnd.n5092 585
R2785 gnd.n5089 gnd.n1759 585
R2786 gnd.n1759 gnd.n1757 585
R2787 gnd.n5088 gnd.n5087 585
R2788 gnd.n5087 gnd.n5086 585
R2789 gnd.n1761 gnd.n1760 585
R2790 gnd.n1770 gnd.n1761 585
R2791 gnd.n5030 gnd.n1769 585
R2792 gnd.n5079 gnd.n1769 585
R2793 gnd.n5032 gnd.n5031 585
R2794 gnd.n5033 gnd.n5032 585
R2795 gnd.n5029 gnd.n1779 585
R2796 gnd.n5068 gnd.n1779 585
R2797 gnd.n5028 gnd.n5027 585
R2798 gnd.n5027 gnd.n1777 585
R2799 gnd.n5026 gnd.n1785 585
R2800 gnd.n5062 gnd.n1785 585
R2801 gnd.n5025 gnd.n5024 585
R2802 gnd.n5024 gnd.n5023 585
R2803 gnd.n1792 gnd.n1791 585
R2804 gnd.n1793 gnd.n1792 585
R2805 gnd.n4991 gnd.n4990 585
R2806 gnd.n4992 gnd.n4991 585
R2807 gnd.n4989 gnd.n1800 585
R2808 gnd.n5012 gnd.n1800 585
R2809 gnd.n4988 gnd.n4987 585
R2810 gnd.n4987 gnd.n1799 585
R2811 gnd.n4986 gnd.n1807 585
R2812 gnd.n5003 gnd.n1807 585
R2813 gnd.n4985 gnd.n4984 585
R2814 gnd.n4984 gnd.n4983 585
R2815 gnd.n1815 gnd.n1814 585
R2816 gnd.n1816 gnd.n1815 585
R2817 gnd.n4958 gnd.n4957 585
R2818 gnd.n4957 gnd.n4956 585
R2819 gnd.n4959 gnd.n1823 585
R2820 gnd.n4972 gnd.n1823 585
R2821 gnd.n4960 gnd.n1831 585
R2822 gnd.n1831 gnd.n1822 585
R2823 gnd.n4962 gnd.n4961 585
R2824 gnd.n4963 gnd.n4962 585
R2825 gnd.n1832 gnd.n1830 585
R2826 gnd.n1841 gnd.n1830 585
R2827 gnd.n4915 gnd.n1840 585
R2828 gnd.n4942 gnd.n1840 585
R2829 gnd.n4916 gnd.n1848 585
R2830 gnd.n4934 gnd.n1848 585
R2831 gnd.n4917 gnd.n1847 585
R2832 gnd.n4936 gnd.n1847 585
R2833 gnd.n4919 gnd.n4918 585
R2834 gnd.n4920 gnd.n4919 585
R2835 gnd.n4914 gnd.n1857 585
R2836 gnd.n1857 gnd.n1855 585
R2837 gnd.n4913 gnd.n4912 585
R2838 gnd.n4912 gnd.n4911 585
R2839 gnd.n1859 gnd.n1858 585
R2840 gnd.n4852 gnd.n1859 585
R2841 gnd.n4877 gnd.n1867 585
R2842 gnd.n4904 gnd.n1867 585
R2843 gnd.n4880 gnd.n4879 585
R2844 gnd.n4879 gnd.n4878 585
R2845 gnd.n4881 gnd.n1874 585
R2846 gnd.n4892 gnd.n1874 585
R2847 gnd.n4883 gnd.n4882 585
R2848 gnd.n4884 gnd.n4883 585
R2849 gnd.n4876 gnd.n1880 585
R2850 gnd.n4886 gnd.n1880 585
R2851 gnd.n4875 gnd.n4874 585
R2852 gnd.n4874 gnd.n4873 585
R2853 gnd.n1883 gnd.n1882 585
R2854 gnd.n4824 gnd.n1883 585
R2855 gnd.n4806 gnd.n4805 585
R2856 gnd.n4806 gnd.n1892 585
R2857 gnd.n4807 gnd.n4804 585
R2858 gnd.n4807 gnd.n1891 585
R2859 gnd.n4811 gnd.n4810 585
R2860 gnd.n4810 gnd.n4809 585
R2861 gnd.n4812 gnd.n1900 585
R2862 gnd.n4832 gnd.n1900 585
R2863 gnd.n4814 gnd.n4813 585
R2864 gnd.n4815 gnd.n4814 585
R2865 gnd.n4803 gnd.n1907 585
R2866 gnd.n4817 gnd.n1907 585
R2867 gnd.n4802 gnd.n4801 585
R2868 gnd.n4801 gnd.n4800 585
R2869 gnd.n1909 gnd.n1908 585
R2870 gnd.n4775 gnd.n1909 585
R2871 gnd.n4788 gnd.n1919 585
R2872 gnd.n4777 gnd.n1919 585
R2873 gnd.n4790 gnd.n4789 585
R2874 gnd.n4791 gnd.n4790 585
R2875 gnd.n4787 gnd.n1918 585
R2876 gnd.n1929 gnd.n1918 585
R2877 gnd.n4786 gnd.n4785 585
R2878 gnd.n4785 gnd.n4784 585
R2879 gnd.n1921 gnd.n1920 585
R2880 gnd.n4757 gnd.n1921 585
R2881 gnd.n2014 gnd.n1938 585
R2882 gnd.n4751 gnd.n1938 585
R2883 gnd.n2016 gnd.n2015 585
R2884 gnd.n2016 gnd.n1223 585
R2885 gnd.n2018 gnd.n2017 585
R2886 gnd.n2017 gnd.n1221 585
R2887 gnd.n2019 gnd.n1942 585
R2888 gnd.n4744 gnd.n1942 585
R2889 gnd.n2022 gnd.n2021 585
R2890 gnd.n2021 gnd.n2020 585
R2891 gnd.n2023 gnd.n1211 585
R2892 gnd.n6256 gnd.n1211 585
R2893 gnd.n2025 gnd.n2024 585
R2894 gnd.n2026 gnd.n2025 585
R2895 gnd.n6380 gnd.n6379 585
R2896 gnd.n6381 gnd.n6380 585
R2897 gnd.n1082 gnd.n1081 585
R2898 gnd.n4358 gnd.n1082 585
R2899 gnd.n6389 gnd.n6388 585
R2900 gnd.n6388 gnd.n6387 585
R2901 gnd.n6390 gnd.n1076 585
R2902 gnd.n4351 gnd.n1076 585
R2903 gnd.n6392 gnd.n6391 585
R2904 gnd.n6393 gnd.n6392 585
R2905 gnd.n1062 gnd.n1061 585
R2906 gnd.n4346 gnd.n1062 585
R2907 gnd.n6401 gnd.n6400 585
R2908 gnd.n6400 gnd.n6399 585
R2909 gnd.n6402 gnd.n1056 585
R2910 gnd.n4373 gnd.n1056 585
R2911 gnd.n6404 gnd.n6403 585
R2912 gnd.n6405 gnd.n6404 585
R2913 gnd.n1041 gnd.n1040 585
R2914 gnd.n4339 gnd.n1041 585
R2915 gnd.n6413 gnd.n6412 585
R2916 gnd.n6412 gnd.n6411 585
R2917 gnd.n6414 gnd.n1035 585
R2918 gnd.n4331 gnd.n1035 585
R2919 gnd.n6416 gnd.n6415 585
R2920 gnd.n6417 gnd.n6416 585
R2921 gnd.n1022 gnd.n1021 585
R2922 gnd.n4324 gnd.n1022 585
R2923 gnd.n6425 gnd.n6424 585
R2924 gnd.n6424 gnd.n6423 585
R2925 gnd.n6426 gnd.n1016 585
R2926 gnd.n4316 gnd.n1016 585
R2927 gnd.n6428 gnd.n6427 585
R2928 gnd.n6429 gnd.n6428 585
R2929 gnd.n1001 gnd.n1000 585
R2930 gnd.n4263 gnd.n1001 585
R2931 gnd.n6437 gnd.n6436 585
R2932 gnd.n6436 gnd.n6435 585
R2933 gnd.n6438 gnd.n996 585
R2934 gnd.n4254 gnd.n996 585
R2935 gnd.n6440 gnd.n6439 585
R2936 gnd.n6441 gnd.n6440 585
R2937 gnd.n981 gnd.n979 585
R2938 gnd.n4248 gnd.n981 585
R2939 gnd.n6449 gnd.n6448 585
R2940 gnd.n6448 gnd.n6447 585
R2941 gnd.n980 gnd.n978 585
R2942 gnd.n4277 gnd.n980 585
R2943 gnd.n4240 gnd.n4239 585
R2944 gnd.n4241 gnd.n4240 585
R2945 gnd.n4238 gnd.n4237 585
R2946 gnd.n4237 gnd.n4236 585
R2947 gnd.n4224 gnd.n2147 585
R2948 gnd.n4216 gnd.n2147 585
R2949 gnd.n4226 gnd.n4225 585
R2950 gnd.n4227 gnd.n4226 585
R2951 gnd.n4223 gnd.n2158 585
R2952 gnd.n4223 gnd.n4222 585
R2953 gnd.n2157 gnd.n977 585
R2954 gnd.n4176 gnd.n2157 585
R2955 gnd.n970 gnd.n969 585
R2956 gnd.n4178 gnd.n969 585
R2957 gnd.n6453 gnd.n6452 585
R2958 gnd.n6454 gnd.n6453 585
R2959 gnd.n953 gnd.n952 585
R2960 gnd.n4184 gnd.n953 585
R2961 gnd.n6462 gnd.n6461 585
R2962 gnd.n6461 gnd.n6460 585
R2963 gnd.n6463 gnd.n947 585
R2964 gnd.n4190 gnd.n947 585
R2965 gnd.n6465 gnd.n6464 585
R2966 gnd.n6466 gnd.n6465 585
R2967 gnd.n948 gnd.n946 585
R2968 gnd.n946 gnd.n941 585
R2969 gnd.n4151 gnd.n4150 585
R2970 gnd.n4152 gnd.n4151 585
R2971 gnd.n2187 gnd.n2186 585
R2972 gnd.n4136 gnd.n2186 585
R2973 gnd.n4145 gnd.n4144 585
R2974 gnd.n4144 gnd.n4143 585
R2975 gnd.n2190 gnd.n2189 585
R2976 gnd.n2191 gnd.n2190 585
R2977 gnd.n4120 gnd.n4119 585
R2978 gnd.n4121 gnd.n4120 585
R2979 gnd.n2209 gnd.n2208 585
R2980 gnd.n2215 gnd.n2208 585
R2981 gnd.n4115 gnd.n4114 585
R2982 gnd.n4114 gnd.n4113 585
R2983 gnd.n2212 gnd.n2211 585
R2984 gnd.n4099 gnd.n2212 585
R2985 gnd.n4084 gnd.n2234 585
R2986 gnd.n2234 gnd.n2225 585
R2987 gnd.n4086 gnd.n4085 585
R2988 gnd.n4087 gnd.n4086 585
R2989 gnd.n2235 gnd.n2233 585
R2990 gnd.n2242 gnd.n2233 585
R2991 gnd.n4079 gnd.n4078 585
R2992 gnd.n4078 gnd.n4077 585
R2993 gnd.n2238 gnd.n2237 585
R2994 gnd.n2239 gnd.n2238 585
R2995 gnd.n4060 gnd.n4059 585
R2996 gnd.n4061 gnd.n4060 585
R2997 gnd.n2255 gnd.n2254 585
R2998 gnd.n2254 gnd.n2251 585
R2999 gnd.n4055 gnd.n4054 585
R3000 gnd.n4054 gnd.n4053 585
R3001 gnd.n2258 gnd.n2257 585
R3002 gnd.n2259 gnd.n2258 585
R3003 gnd.n4041 gnd.n4040 585
R3004 gnd.n4039 gnd.n3788 585
R3005 gnd.n4038 gnd.n3787 585
R3006 gnd.n4043 gnd.n3787 585
R3007 gnd.n4037 gnd.n4036 585
R3008 gnd.n4035 gnd.n4034 585
R3009 gnd.n4033 gnd.n4032 585
R3010 gnd.n4031 gnd.n4030 585
R3011 gnd.n4029 gnd.n4028 585
R3012 gnd.n4027 gnd.n4026 585
R3013 gnd.n4025 gnd.n4024 585
R3014 gnd.n4023 gnd.n4022 585
R3015 gnd.n4021 gnd.n4020 585
R3016 gnd.n4019 gnd.n4018 585
R3017 gnd.n4017 gnd.n4016 585
R3018 gnd.n4015 gnd.n4014 585
R3019 gnd.n4013 gnd.n4012 585
R3020 gnd.n4011 gnd.n4010 585
R3021 gnd.n4009 gnd.n4008 585
R3022 gnd.n4006 gnd.n4005 585
R3023 gnd.n4004 gnd.n4003 585
R3024 gnd.n4002 gnd.n4001 585
R3025 gnd.n4000 gnd.n3999 585
R3026 gnd.n3998 gnd.n3997 585
R3027 gnd.n3996 gnd.n3995 585
R3028 gnd.n3994 gnd.n3993 585
R3029 gnd.n3992 gnd.n3991 585
R3030 gnd.n3990 gnd.n3989 585
R3031 gnd.n3988 gnd.n3987 585
R3032 gnd.n3986 gnd.n3985 585
R3033 gnd.n3984 gnd.n3983 585
R3034 gnd.n3982 gnd.n3981 585
R3035 gnd.n3980 gnd.n3979 585
R3036 gnd.n3978 gnd.n3977 585
R3037 gnd.n3976 gnd.n3975 585
R3038 gnd.n3974 gnd.n3973 585
R3039 gnd.n3972 gnd.n3971 585
R3040 gnd.n3970 gnd.n3969 585
R3041 gnd.n3968 gnd.n3967 585
R3042 gnd.n3966 gnd.n3965 585
R3043 gnd.n3964 gnd.n3963 585
R3044 gnd.n3962 gnd.n3961 585
R3045 gnd.n3960 gnd.n3959 585
R3046 gnd.n3958 gnd.n3957 585
R3047 gnd.n3956 gnd.n3955 585
R3048 gnd.n3954 gnd.n3953 585
R3049 gnd.n3952 gnd.n3951 585
R3050 gnd.n3950 gnd.n3949 585
R3051 gnd.n3948 gnd.n3947 585
R3052 gnd.n3946 gnd.n3945 585
R3053 gnd.n3944 gnd.n3943 585
R3054 gnd.n3942 gnd.n3941 585
R3055 gnd.n3940 gnd.n3939 585
R3056 gnd.n3938 gnd.n3937 585
R3057 gnd.n3936 gnd.n3935 585
R3058 gnd.n3934 gnd.n3933 585
R3059 gnd.n3932 gnd.n3931 585
R3060 gnd.n3930 gnd.n3929 585
R3061 gnd.n3928 gnd.n2271 585
R3062 gnd.n4045 gnd.n2270 585
R3063 gnd.n4533 gnd.n4532 585
R3064 gnd.n4530 gnd.n4426 585
R3065 gnd.n4529 gnd.n4528 585
R3066 gnd.n4522 gnd.n4428 585
R3067 gnd.n4524 gnd.n4523 585
R3068 gnd.n4520 gnd.n4430 585
R3069 gnd.n4519 gnd.n4518 585
R3070 gnd.n4512 gnd.n4432 585
R3071 gnd.n4514 gnd.n4513 585
R3072 gnd.n4510 gnd.n4434 585
R3073 gnd.n4509 gnd.n4508 585
R3074 gnd.n4502 gnd.n4436 585
R3075 gnd.n4504 gnd.n4503 585
R3076 gnd.n4500 gnd.n4438 585
R3077 gnd.n4499 gnd.n4498 585
R3078 gnd.n4492 gnd.n4440 585
R3079 gnd.n4494 gnd.n4493 585
R3080 gnd.n4490 gnd.n4442 585
R3081 gnd.n4489 gnd.n4488 585
R3082 gnd.n4482 gnd.n4444 585
R3083 gnd.n4484 gnd.n4483 585
R3084 gnd.n4480 gnd.n4448 585
R3085 gnd.n4479 gnd.n4478 585
R3086 gnd.n4472 gnd.n4450 585
R3087 gnd.n4474 gnd.n4473 585
R3088 gnd.n4470 gnd.n4452 585
R3089 gnd.n4469 gnd.n4468 585
R3090 gnd.n4462 gnd.n4454 585
R3091 gnd.n4464 gnd.n4463 585
R3092 gnd.n4460 gnd.n4457 585
R3093 gnd.n4459 gnd.n1144 585
R3094 gnd.n6331 gnd.n1140 585
R3095 gnd.n6333 gnd.n6332 585
R3096 gnd.n6335 gnd.n1138 585
R3097 gnd.n6337 gnd.n6336 585
R3098 gnd.n6338 gnd.n1133 585
R3099 gnd.n6340 gnd.n6339 585
R3100 gnd.n6342 gnd.n1131 585
R3101 gnd.n6344 gnd.n6343 585
R3102 gnd.n6346 gnd.n1124 585
R3103 gnd.n6348 gnd.n6347 585
R3104 gnd.n6350 gnd.n1122 585
R3105 gnd.n6352 gnd.n6351 585
R3106 gnd.n6353 gnd.n1117 585
R3107 gnd.n6355 gnd.n6354 585
R3108 gnd.n6357 gnd.n1115 585
R3109 gnd.n6359 gnd.n6358 585
R3110 gnd.n6360 gnd.n1110 585
R3111 gnd.n6362 gnd.n6361 585
R3112 gnd.n6364 gnd.n1108 585
R3113 gnd.n6366 gnd.n6365 585
R3114 gnd.n6367 gnd.n1102 585
R3115 gnd.n6369 gnd.n6368 585
R3116 gnd.n6371 gnd.n1101 585
R3117 gnd.n6372 gnd.n1099 585
R3118 gnd.n6375 gnd.n6374 585
R3119 gnd.n6376 gnd.n1096 585
R3120 gnd.n1100 gnd.n1096 585
R3121 gnd.n4355 gnd.n1093 585
R3122 gnd.n6381 gnd.n1093 585
R3123 gnd.n4357 gnd.n4356 585
R3124 gnd.n4358 gnd.n4357 585
R3125 gnd.n4354 gnd.n1084 585
R3126 gnd.n6387 gnd.n1084 585
R3127 gnd.n4353 gnd.n4352 585
R3128 gnd.n4352 gnd.n4351 585
R3129 gnd.n4349 gnd.n1073 585
R3130 gnd.n6393 gnd.n1073 585
R3131 gnd.n4348 gnd.n4347 585
R3132 gnd.n4347 gnd.n4346 585
R3133 gnd.n4345 gnd.n1063 585
R3134 gnd.n6399 gnd.n1063 585
R3135 gnd.n4344 gnd.n2101 585
R3136 gnd.n4373 gnd.n2101 585
R3137 gnd.n4342 gnd.n1053 585
R3138 gnd.n6405 gnd.n1053 585
R3139 gnd.n4341 gnd.n4340 585
R3140 gnd.n4340 gnd.n4339 585
R3141 gnd.n2110 gnd.n1043 585
R3142 gnd.n6411 gnd.n1043 585
R3143 gnd.n4330 gnd.n4329 585
R3144 gnd.n4331 gnd.n4330 585
R3145 gnd.n4327 gnd.n1033 585
R3146 gnd.n6417 gnd.n1033 585
R3147 gnd.n4326 gnd.n4325 585
R3148 gnd.n4325 gnd.n4324 585
R3149 gnd.n2115 gnd.n1023 585
R3150 gnd.n6423 gnd.n1023 585
R3151 gnd.n4259 gnd.n2119 585
R3152 gnd.n4316 gnd.n2119 585
R3153 gnd.n4260 gnd.n1013 585
R3154 gnd.n6429 gnd.n1013 585
R3155 gnd.n4262 gnd.n4261 585
R3156 gnd.n4263 gnd.n4262 585
R3157 gnd.n4257 gnd.n1003 585
R3158 gnd.n6435 gnd.n1003 585
R3159 gnd.n4256 gnd.n4255 585
R3160 gnd.n4255 gnd.n4254 585
R3161 gnd.n4251 gnd.n994 585
R3162 gnd.n6441 gnd.n994 585
R3163 gnd.n4250 gnd.n4249 585
R3164 gnd.n4249 gnd.n4248 585
R3165 gnd.n4247 gnd.n982 585
R3166 gnd.n6447 gnd.n982 585
R3167 gnd.n4246 gnd.n2132 585
R3168 gnd.n4277 gnd.n2132 585
R3169 gnd.n2146 gnd.n2141 585
R3170 gnd.n4241 gnd.n2146 585
R3171 gnd.n4163 gnd.n2148 585
R3172 gnd.n4236 gnd.n2148 585
R3173 gnd.n4164 gnd.n2167 585
R3174 gnd.n4216 gnd.n2167 585
R3175 gnd.n4165 gnd.n2154 585
R3176 gnd.n4227 gnd.n2154 585
R3177 gnd.n4166 gnd.n2160 585
R3178 gnd.n4222 gnd.n2160 585
R3179 gnd.n4168 gnd.n4167 585
R3180 gnd.n4176 gnd.n4168 585
R3181 gnd.n4180 gnd.n4179 585
R3182 gnd.n4179 gnd.n4178 585
R3183 gnd.n4181 gnd.n966 585
R3184 gnd.n6454 gnd.n966 585
R3185 gnd.n4183 gnd.n4182 585
R3186 gnd.n4184 gnd.n4183 585
R3187 gnd.n4160 gnd.n954 585
R3188 gnd.n6460 gnd.n954 585
R3189 gnd.n4159 gnd.n2173 585
R3190 gnd.n4190 gnd.n2173 585
R3191 gnd.n2179 gnd.n942 585
R3192 gnd.n6466 gnd.n942 585
R3193 gnd.n2200 gnd.n2199 585
R3194 gnd.n2199 gnd.n941 585
R3195 gnd.n2201 gnd.n2184 585
R3196 gnd.n4152 gnd.n2184 585
R3197 gnd.n4138 gnd.n4137 585
R3198 gnd.n4137 gnd.n4136 585
R3199 gnd.n2198 gnd.n2192 585
R3200 gnd.n4143 gnd.n2192 585
R3201 gnd.n4106 gnd.n4105 585
R3202 gnd.n4105 gnd.n2191 585
R3203 gnd.n4107 gnd.n2206 585
R3204 gnd.n4121 gnd.n2206 585
R3205 gnd.n4104 gnd.n4103 585
R3206 gnd.n4103 gnd.n2215 585
R3207 gnd.n4102 gnd.n2213 585
R3208 gnd.n4113 gnd.n2213 585
R3209 gnd.n4101 gnd.n4100 585
R3210 gnd.n4100 gnd.n4099 585
R3211 gnd.n2224 gnd.n2222 585
R3212 gnd.n2225 gnd.n2224 585
R3213 gnd.n4068 gnd.n2231 585
R3214 gnd.n4087 gnd.n2231 585
R3215 gnd.n4067 gnd.n4066 585
R3216 gnd.n4066 gnd.n2242 585
R3217 gnd.n4065 gnd.n2240 585
R3218 gnd.n4077 gnd.n2240 585
R3219 gnd.n4064 gnd.n4063 585
R3220 gnd.n4063 gnd.n2239 585
R3221 gnd.n4062 gnd.n2248 585
R3222 gnd.n4062 gnd.n4061 585
R3223 gnd.n4048 gnd.n2250 585
R3224 gnd.n2251 gnd.n2250 585
R3225 gnd.n4049 gnd.n2260 585
R3226 gnd.n4053 gnd.n2260 585
R3227 gnd.n4047 gnd.n4046 585
R3228 gnd.n4046 gnd.n2259 585
R3229 gnd.n7563 gnd.n7562 585
R3230 gnd.n7564 gnd.n7563 585
R3231 gnd.n199 gnd.n198 585
R3232 gnd.n7413 gnd.n199 585
R3233 gnd.n7572 gnd.n7571 585
R3234 gnd.n7571 gnd.n7570 585
R3235 gnd.n7573 gnd.n193 585
R3236 gnd.n193 gnd.n192 585
R3237 gnd.n7575 gnd.n7574 585
R3238 gnd.n7576 gnd.n7575 585
R3239 gnd.n180 gnd.n179 585
R3240 gnd.n183 gnd.n180 585
R3241 gnd.n7584 gnd.n7583 585
R3242 gnd.n7583 gnd.n7582 585
R3243 gnd.n7585 gnd.n174 585
R3244 gnd.n174 gnd.n173 585
R3245 gnd.n7587 gnd.n7586 585
R3246 gnd.n7588 gnd.n7587 585
R3247 gnd.n160 gnd.n159 585
R3248 gnd.n170 gnd.n160 585
R3249 gnd.n7596 gnd.n7595 585
R3250 gnd.n7595 gnd.n7594 585
R3251 gnd.n7597 gnd.n154 585
R3252 gnd.n161 gnd.n154 585
R3253 gnd.n7599 gnd.n7598 585
R3254 gnd.n7600 gnd.n7599 585
R3255 gnd.n142 gnd.n141 585
R3256 gnd.n145 gnd.n142 585
R3257 gnd.n7608 gnd.n7607 585
R3258 gnd.n7607 gnd.n7606 585
R3259 gnd.n7609 gnd.n136 585
R3260 gnd.n7385 gnd.n136 585
R3261 gnd.n7611 gnd.n7610 585
R3262 gnd.n7612 gnd.n7611 585
R3263 gnd.n122 gnd.n121 585
R3264 gnd.n132 gnd.n122 585
R3265 gnd.n7620 gnd.n7619 585
R3266 gnd.n7619 gnd.n7618 585
R3267 gnd.n7621 gnd.n117 585
R3268 gnd.n7343 gnd.n117 585
R3269 gnd.n7623 gnd.n7622 585
R3270 gnd.n7624 gnd.n7623 585
R3271 gnd.n101 gnd.n99 585
R3272 gnd.n7333 gnd.n101 585
R3273 gnd.n7632 gnd.n7631 585
R3274 gnd.n7631 gnd.n7630 585
R3275 gnd.n100 gnd.n92 585
R3276 gnd.n7324 gnd.n100 585
R3277 gnd.n7635 gnd.n90 585
R3278 gnd.n7317 gnd.n90 585
R3279 gnd.n7637 gnd.n7636 585
R3280 gnd.n7638 gnd.n7637 585
R3281 gnd.n379 gnd.n89 585
R3282 gnd.n7313 gnd.n89 585
R3283 gnd.n7301 gnd.n380 585
R3284 gnd.n7301 gnd.n7300 585
R3285 gnd.n7303 gnd.n7302 585
R3286 gnd.n7304 gnd.n7303 585
R3287 gnd.n378 gnd.n97 585
R3288 gnd.n1460 gnd.n378 585
R3289 gnd.n1449 gnd.n1448 585
R3290 gnd.n6049 gnd.n1449 585
R3291 gnd.n6058 gnd.n6057 585
R3292 gnd.n6057 gnd.n6056 585
R3293 gnd.n6059 gnd.n1445 585
R3294 gnd.n6021 gnd.n1445 585
R3295 gnd.n6061 gnd.n6060 585
R3296 gnd.n6062 gnd.n6061 585
R3297 gnd.n1431 gnd.n1430 585
R3298 gnd.n6037 gnd.n1431 585
R3299 gnd.n6070 gnd.n6069 585
R3300 gnd.n6069 gnd.n6068 585
R3301 gnd.n6071 gnd.n1425 585
R3302 gnd.n6012 gnd.n1425 585
R3303 gnd.n6073 gnd.n6072 585
R3304 gnd.n6074 gnd.n6073 585
R3305 gnd.n1411 gnd.n1410 585
R3306 gnd.n6004 gnd.n1411 585
R3307 gnd.n6082 gnd.n6081 585
R3308 gnd.n6081 gnd.n6080 585
R3309 gnd.n6083 gnd.n1405 585
R3310 gnd.n5998 gnd.n1405 585
R3311 gnd.n6085 gnd.n6084 585
R3312 gnd.n6086 gnd.n6085 585
R3313 gnd.n1391 gnd.n1390 585
R3314 gnd.n5990 gnd.n1391 585
R3315 gnd.n6094 gnd.n6093 585
R3316 gnd.n6093 gnd.n6092 585
R3317 gnd.n6095 gnd.n1385 585
R3318 gnd.n5928 gnd.n1385 585
R3319 gnd.n6097 gnd.n6096 585
R3320 gnd.n6098 gnd.n6097 585
R3321 gnd.n1371 gnd.n1370 585
R3322 gnd.n5936 gnd.n1371 585
R3323 gnd.n6106 gnd.n6105 585
R3324 gnd.n6105 gnd.n6104 585
R3325 gnd.n6107 gnd.n1365 585
R3326 gnd.n5917 gnd.n1365 585
R3327 gnd.n6109 gnd.n6108 585
R3328 gnd.n6110 gnd.n6109 585
R3329 gnd.n1348 gnd.n1347 585
R3330 gnd.n5909 gnd.n1348 585
R3331 gnd.n6118 gnd.n6117 585
R3332 gnd.n6117 gnd.n6116 585
R3333 gnd.n6119 gnd.n1343 585
R3334 gnd.n5361 gnd.n1343 585
R3335 gnd.n6121 gnd.n6120 585
R3336 gnd.n6122 gnd.n6121 585
R3337 gnd.n5750 gnd.n1342 585
R3338 gnd.n5755 gnd.n5753 585
R3339 gnd.n5756 gnd.n5749 585
R3340 gnd.n5756 gnd.n1329 585
R3341 gnd.n5759 gnd.n5758 585
R3342 gnd.n5747 gnd.n5746 585
R3343 gnd.n5764 gnd.n5763 585
R3344 gnd.n5766 gnd.n5745 585
R3345 gnd.n5769 gnd.n5768 585
R3346 gnd.n5743 gnd.n5742 585
R3347 gnd.n5774 gnd.n5773 585
R3348 gnd.n5776 gnd.n5741 585
R3349 gnd.n5779 gnd.n5778 585
R3350 gnd.n5739 gnd.n5738 585
R3351 gnd.n5784 gnd.n5783 585
R3352 gnd.n5786 gnd.n5737 585
R3353 gnd.n5789 gnd.n5788 585
R3354 gnd.n5735 gnd.n5734 585
R3355 gnd.n5797 gnd.n5796 585
R3356 gnd.n5799 gnd.n5733 585
R3357 gnd.n5802 gnd.n5801 585
R3358 gnd.n5731 gnd.n5730 585
R3359 gnd.n5807 gnd.n5806 585
R3360 gnd.n5809 gnd.n5729 585
R3361 gnd.n5812 gnd.n5811 585
R3362 gnd.n5727 gnd.n5726 585
R3363 gnd.n5818 gnd.n5817 585
R3364 gnd.n5822 gnd.n1531 585
R3365 gnd.n5825 gnd.n5824 585
R3366 gnd.n1529 gnd.n1528 585
R3367 gnd.n5830 gnd.n5829 585
R3368 gnd.n5832 gnd.n1527 585
R3369 gnd.n5835 gnd.n5834 585
R3370 gnd.n1525 gnd.n1524 585
R3371 gnd.n5840 gnd.n5839 585
R3372 gnd.n5842 gnd.n1523 585
R3373 gnd.n5847 gnd.n5844 585
R3374 gnd.n1521 gnd.n1520 585
R3375 gnd.n5852 gnd.n5851 585
R3376 gnd.n5854 gnd.n1519 585
R3377 gnd.n5857 gnd.n5856 585
R3378 gnd.n1517 gnd.n1516 585
R3379 gnd.n5862 gnd.n5861 585
R3380 gnd.n5864 gnd.n1515 585
R3381 gnd.n5867 gnd.n5866 585
R3382 gnd.n1513 gnd.n1512 585
R3383 gnd.n5872 gnd.n5871 585
R3384 gnd.n5874 gnd.n1511 585
R3385 gnd.n5877 gnd.n5876 585
R3386 gnd.n1509 gnd.n1508 585
R3387 gnd.n5882 gnd.n5881 585
R3388 gnd.n5884 gnd.n1507 585
R3389 gnd.n5887 gnd.n5886 585
R3390 gnd.n1505 gnd.n1504 585
R3391 gnd.n5893 gnd.n5892 585
R3392 gnd.n5895 gnd.n1503 585
R3393 gnd.n5896 gnd.n1502 585
R3394 gnd.n5899 gnd.n5898 585
R3395 gnd.n7454 gnd.n7453 585
R3396 gnd.n7456 gnd.n313 585
R3397 gnd.n7458 gnd.n7457 585
R3398 gnd.n7459 gnd.n306 585
R3399 gnd.n7461 gnd.n7460 585
R3400 gnd.n7463 gnd.n304 585
R3401 gnd.n7465 gnd.n7464 585
R3402 gnd.n7466 gnd.n299 585
R3403 gnd.n7468 gnd.n7467 585
R3404 gnd.n7470 gnd.n297 585
R3405 gnd.n7472 gnd.n7471 585
R3406 gnd.n7473 gnd.n292 585
R3407 gnd.n7475 gnd.n7474 585
R3408 gnd.n7477 gnd.n290 585
R3409 gnd.n7479 gnd.n7478 585
R3410 gnd.n7480 gnd.n285 585
R3411 gnd.n7482 gnd.n7481 585
R3412 gnd.n7484 gnd.n284 585
R3413 gnd.n7485 gnd.n281 585
R3414 gnd.n7488 gnd.n7487 585
R3415 gnd.n283 gnd.n277 585
R3416 gnd.n7492 gnd.n274 585
R3417 gnd.n7494 gnd.n7493 585
R3418 gnd.n7496 gnd.n272 585
R3419 gnd.n7498 gnd.n7497 585
R3420 gnd.n7499 gnd.n267 585
R3421 gnd.n7501 gnd.n7500 585
R3422 gnd.n7503 gnd.n265 585
R3423 gnd.n7505 gnd.n7504 585
R3424 gnd.n7506 gnd.n260 585
R3425 gnd.n7508 gnd.n7507 585
R3426 gnd.n7510 gnd.n258 585
R3427 gnd.n7512 gnd.n7511 585
R3428 gnd.n7513 gnd.n253 585
R3429 gnd.n7515 gnd.n7514 585
R3430 gnd.n7517 gnd.n251 585
R3431 gnd.n7519 gnd.n7518 585
R3432 gnd.n7520 gnd.n246 585
R3433 gnd.n7522 gnd.n7521 585
R3434 gnd.n7524 gnd.n244 585
R3435 gnd.n7526 gnd.n7525 585
R3436 gnd.n7530 gnd.n239 585
R3437 gnd.n7532 gnd.n7531 585
R3438 gnd.n7534 gnd.n237 585
R3439 gnd.n7536 gnd.n7535 585
R3440 gnd.n7537 gnd.n232 585
R3441 gnd.n7539 gnd.n7538 585
R3442 gnd.n7541 gnd.n230 585
R3443 gnd.n7543 gnd.n7542 585
R3444 gnd.n7544 gnd.n225 585
R3445 gnd.n7546 gnd.n7545 585
R3446 gnd.n7548 gnd.n223 585
R3447 gnd.n7550 gnd.n7549 585
R3448 gnd.n7551 gnd.n218 585
R3449 gnd.n7553 gnd.n7552 585
R3450 gnd.n7555 gnd.n216 585
R3451 gnd.n7557 gnd.n7556 585
R3452 gnd.n7558 gnd.n214 585
R3453 gnd.n7559 gnd.n211 585
R3454 gnd.n211 gnd.n210 585
R3455 gnd.n7410 gnd.n208 585
R3456 gnd.n7564 gnd.n208 585
R3457 gnd.n7412 gnd.n7411 585
R3458 gnd.n7413 gnd.n7412 585
R3459 gnd.n7409 gnd.n200 585
R3460 gnd.n7570 gnd.n200 585
R3461 gnd.n7408 gnd.n7407 585
R3462 gnd.n7407 gnd.n192 585
R3463 gnd.n7405 gnd.n190 585
R3464 gnd.n7576 gnd.n190 585
R3465 gnd.n7404 gnd.n7403 585
R3466 gnd.n7403 gnd.n183 585
R3467 gnd.n7402 gnd.n181 585
R3468 gnd.n7582 gnd.n181 585
R3469 gnd.n7401 gnd.n7400 585
R3470 gnd.n7400 gnd.n173 585
R3471 gnd.n7398 gnd.n171 585
R3472 gnd.n7588 gnd.n171 585
R3473 gnd.n7397 gnd.n7396 585
R3474 gnd.n7396 gnd.n170 585
R3475 gnd.n7395 gnd.n162 585
R3476 gnd.n7594 gnd.n162 585
R3477 gnd.n7394 gnd.n7393 585
R3478 gnd.n7393 gnd.n161 585
R3479 gnd.n7391 gnd.n152 585
R3480 gnd.n7600 gnd.n152 585
R3481 gnd.n7390 gnd.n7389 585
R3482 gnd.n7389 gnd.n145 585
R3483 gnd.n7388 gnd.n143 585
R3484 gnd.n7606 gnd.n143 585
R3485 gnd.n7387 gnd.n7386 585
R3486 gnd.n7386 gnd.n7385 585
R3487 gnd.n352 gnd.n133 585
R3488 gnd.n7612 gnd.n133 585
R3489 gnd.n7339 gnd.n7338 585
R3490 gnd.n7338 gnd.n132 585
R3491 gnd.n7340 gnd.n124 585
R3492 gnd.n7618 gnd.n124 585
R3493 gnd.n7342 gnd.n7341 585
R3494 gnd.n7343 gnd.n7342 585
R3495 gnd.n7336 gnd.n115 585
R3496 gnd.n7624 gnd.n115 585
R3497 gnd.n7335 gnd.n7334 585
R3498 gnd.n7334 gnd.n7333 585
R3499 gnd.n359 gnd.n103 585
R3500 gnd.n7630 gnd.n103 585
R3501 gnd.n7323 gnd.n7322 585
R3502 gnd.n7324 gnd.n7323 585
R3503 gnd.n364 gnd.n363 585
R3504 gnd.n7317 gnd.n363 585
R3505 gnd.n7310 gnd.n86 585
R3506 gnd.n7638 gnd.n86 585
R3507 gnd.n7312 gnd.n7311 585
R3508 gnd.n7313 gnd.n7312 585
R3509 gnd.n7309 gnd.n370 585
R3510 gnd.n7300 gnd.n370 585
R3511 gnd.n376 gnd.n371 585
R3512 gnd.n7304 gnd.n376 585
R3513 gnd.n1457 gnd.n1456 585
R3514 gnd.n1460 gnd.n1457 585
R3515 gnd.n6051 gnd.n6050 585
R3516 gnd.n6050 gnd.n6049 585
R3517 gnd.n1455 gnd.n1451 585
R3518 gnd.n6056 gnd.n1451 585
R3519 gnd.n6020 gnd.n6019 585
R3520 gnd.n6021 gnd.n6020 585
R3521 gnd.n6017 gnd.n1442 585
R3522 gnd.n6062 gnd.n1442 585
R3523 gnd.n6016 gnd.n1465 585
R3524 gnd.n6037 gnd.n1465 585
R3525 gnd.n6015 gnd.n1433 585
R3526 gnd.n6068 gnd.n1433 585
R3527 gnd.n6014 gnd.n6013 585
R3528 gnd.n6013 gnd.n6012 585
R3529 gnd.n1470 gnd.n1422 585
R3530 gnd.n6074 gnd.n1422 585
R3531 gnd.n6003 gnd.n6002 585
R3532 gnd.n6004 gnd.n6003 585
R3533 gnd.n6001 gnd.n1413 585
R3534 gnd.n6080 gnd.n1413 585
R3535 gnd.n6000 gnd.n5999 585
R3536 gnd.n5999 gnd.n5998 585
R3537 gnd.n1476 gnd.n1402 585
R3538 gnd.n6086 gnd.n1402 585
R3539 gnd.n5924 gnd.n1481 585
R3540 gnd.n5990 gnd.n1481 585
R3541 gnd.n5925 gnd.n1393 585
R3542 gnd.n6092 gnd.n1393 585
R3543 gnd.n5927 gnd.n5926 585
R3544 gnd.n5928 gnd.n5927 585
R3545 gnd.n5922 gnd.n1382 585
R3546 gnd.n6098 gnd.n1382 585
R3547 gnd.n5921 gnd.n1487 585
R3548 gnd.n5936 gnd.n1487 585
R3549 gnd.n5920 gnd.n1373 585
R3550 gnd.n6104 gnd.n1373 585
R3551 gnd.n5919 gnd.n5918 585
R3552 gnd.n5918 gnd.n5917 585
R3553 gnd.n1491 gnd.n1362 585
R3554 gnd.n6110 gnd.n1362 585
R3555 gnd.n5908 gnd.n5907 585
R3556 gnd.n5909 gnd.n5908 585
R3557 gnd.n5906 gnd.n1350 585
R3558 gnd.n6116 gnd.n1350 585
R3559 gnd.n5905 gnd.n1497 585
R3560 gnd.n5361 gnd.n1497 585
R3561 gnd.n1496 gnd.n1338 585
R3562 gnd.n6122 gnd.n1338 585
R3563 gnd.n6472 gnd.n935 585
R3564 gnd.n2183 gnd.n935 585
R3565 gnd.n7277 gnd.n7276 585
R3566 gnd.n7277 gnd.n135 585
R3567 gnd.n7279 gnd.n392 585
R3568 gnd.n7279 gnd.n7278 585
R3569 gnd.n7281 gnd.n7280 585
R3570 gnd.n7280 gnd.n123 585
R3571 gnd.n7282 gnd.n387 585
R3572 gnd.n387 gnd.n358 585
R3573 gnd.n7284 gnd.n7283 585
R3574 gnd.n7284 gnd.n114 585
R3575 gnd.n7285 gnd.n386 585
R3576 gnd.n7285 gnd.n105 585
R3577 gnd.n7287 gnd.n7286 585
R3578 gnd.n7286 gnd.n102 585
R3579 gnd.n7289 gnd.n385 585
R3580 gnd.n385 gnd.n362 585
R3581 gnd.n7291 gnd.n7290 585
R3582 gnd.n7291 gnd.n87 585
R3583 gnd.n7293 gnd.n7292 585
R3584 gnd.n7292 gnd.n85 585
R3585 gnd.n7294 gnd.n382 585
R3586 gnd.n382 gnd.n369 585
R3587 gnd.n7297 gnd.n7296 585
R3588 gnd.n7298 gnd.n7297 585
R3589 gnd.n383 gnd.n381 585
R3590 gnd.n381 gnd.n375 585
R3591 gnd.n6047 gnd.n6046 585
R3592 gnd.n6048 gnd.n6047 585
R3593 gnd.n6044 gnd.n1461 585
R3594 gnd.n1461 gnd.n1458 585
R3595 gnd.n6042 gnd.n6041 585
R3596 gnd.n6041 gnd.n1450 585
R3597 gnd.n6040 gnd.n1462 585
R3598 gnd.n6040 gnd.n1444 585
R3599 gnd.n6039 gnd.n1464 585
R3600 gnd.n6039 gnd.n6038 585
R3601 gnd.n5977 gnd.n1463 585
R3602 gnd.n1463 gnd.n1435 585
R3603 gnd.n5979 gnd.n5978 585
R3604 gnd.n5978 gnd.n1432 585
R3605 gnd.n5980 gnd.n5969 585
R3606 gnd.n5969 gnd.n1424 585
R3607 gnd.n5982 gnd.n5981 585
R3608 gnd.n5982 gnd.n1421 585
R3609 gnd.n5983 gnd.n5968 585
R3610 gnd.n5983 gnd.n1475 585
R3611 gnd.n5985 gnd.n5984 585
R3612 gnd.n5984 gnd.n1412 585
R3613 gnd.n5986 gnd.n1483 585
R3614 gnd.n1483 gnd.n1404 585
R3615 gnd.n5988 gnd.n5987 585
R3616 gnd.n5989 gnd.n5988 585
R3617 gnd.n1484 gnd.n1482 585
R3618 gnd.n1482 gnd.n1395 585
R3619 gnd.n5962 gnd.n5961 585
R3620 gnd.n5961 gnd.n1392 585
R3621 gnd.n5960 gnd.n1486 585
R3622 gnd.n5960 gnd.n1384 585
R3623 gnd.n5959 gnd.n5958 585
R3624 gnd.n5959 gnd.n1381 585
R3625 gnd.n5939 gnd.n5938 585
R3626 gnd.n5938 gnd.n5937 585
R3627 gnd.n5954 gnd.n5953 585
R3628 gnd.n5953 gnd.n1372 585
R3629 gnd.n5952 gnd.n5941 585
R3630 gnd.n5952 gnd.n1364 585
R3631 gnd.n5951 gnd.n5950 585
R3632 gnd.n5951 gnd.n1361 585
R3633 gnd.n5943 gnd.n5942 585
R3634 gnd.n5942 gnd.n1352 585
R3635 gnd.n5946 gnd.n5945 585
R3636 gnd.n5945 gnd.n1349 585
R3637 gnd.n1336 gnd.n1335 585
R3638 gnd.n1340 gnd.n1336 585
R3639 gnd.n6125 gnd.n6124 585
R3640 gnd.n6124 gnd.n6123 585
R3641 gnd.n6126 gnd.n1330 585
R3642 gnd.n1337 gnd.n1330 585
R3643 gnd.n6128 gnd.n6127 585
R3644 gnd.n6129 gnd.n6128 585
R3645 gnd.n1327 gnd.n1326 585
R3646 gnd.n6130 gnd.n1327 585
R3647 gnd.n6133 gnd.n6132 585
R3648 gnd.n6132 gnd.n6131 585
R3649 gnd.n6134 gnd.n1321 585
R3650 gnd.n1321 gnd.n1319 585
R3651 gnd.n6136 gnd.n6135 585
R3652 gnd.n6137 gnd.n6136 585
R3653 gnd.n1322 gnd.n1320 585
R3654 gnd.n1320 gnd.n1317 585
R3655 gnd.n1604 gnd.n1603 585
R3656 gnd.n5542 gnd.n1604 585
R3657 gnd.n5546 gnd.n5545 585
R3658 gnd.n5545 gnd.n5544 585
R3659 gnd.n5547 gnd.n1594 585
R3660 gnd.n1605 gnd.n1594 585
R3661 gnd.n5549 gnd.n5548 585
R3662 gnd.n5550 gnd.n5549 585
R3663 gnd.n1595 gnd.n1589 585
R3664 gnd.n5553 gnd.n1589 585
R3665 gnd.n5556 gnd.n1588 585
R3666 gnd.n5556 gnd.n5555 585
R3667 gnd.n5558 gnd.n5557 585
R3668 gnd.n5557 gnd.n1536 585
R3669 gnd.n5559 gnd.n1583 585
R3670 gnd.n1583 gnd.n1573 585
R3671 gnd.n5561 gnd.n5560 585
R3672 gnd.n5562 gnd.n5561 585
R3673 gnd.n1584 gnd.n1582 585
R3674 gnd.n1582 gnd.n1578 585
R3675 gnd.n5313 gnd.n1632 585
R3676 gnd.n1632 gnd.n1631 585
R3677 gnd.n5315 gnd.n5314 585
R3678 gnd.n5316 gnd.n5315 585
R3679 gnd.n1633 gnd.n1630 585
R3680 gnd.n1630 gnd.n1627 585
R3681 gnd.n5307 gnd.n5306 585
R3682 gnd.n5306 gnd.n5305 585
R3683 gnd.n1636 gnd.n1635 585
R3684 gnd.n5293 gnd.n1636 585
R3685 gnd.n5268 gnd.n1662 585
R3686 gnd.n1662 gnd.n1654 585
R3687 gnd.n5270 gnd.n5269 585
R3688 gnd.n5271 gnd.n5270 585
R3689 gnd.n1663 gnd.n1661 585
R3690 gnd.n5258 gnd.n1661 585
R3691 gnd.n5263 gnd.n5262 585
R3692 gnd.n5262 gnd.n5261 585
R3693 gnd.n1666 gnd.n1665 585
R3694 gnd.n1678 gnd.n1666 585
R3695 gnd.n5242 gnd.n5241 585
R3696 gnd.n5243 gnd.n5242 585
R3697 gnd.n1683 gnd.n1682 585
R3698 gnd.n1690 gnd.n1682 585
R3699 gnd.n5237 gnd.n5236 585
R3700 gnd.n5236 gnd.n5235 585
R3701 gnd.n1686 gnd.n1685 585
R3702 gnd.n5132 gnd.n1686 585
R3703 gnd.n5191 gnd.n1710 585
R3704 gnd.n1710 gnd.n1703 585
R3705 gnd.n5193 gnd.n5192 585
R3706 gnd.n5194 gnd.n5193 585
R3707 gnd.n1711 gnd.n1709 585
R3708 gnd.n1709 gnd.n1707 585
R3709 gnd.n5186 gnd.n5185 585
R3710 gnd.n5185 gnd.n5184 585
R3711 gnd.n1714 gnd.n1713 585
R3712 gnd.n5176 gnd.n1714 585
R3713 gnd.n5162 gnd.n5161 585
R3714 gnd.n5163 gnd.n5162 585
R3715 gnd.n1733 gnd.n1732 585
R3716 gnd.n5112 gnd.n1732 585
R3717 gnd.n5157 gnd.n5156 585
R3718 gnd.n5156 gnd.n5155 585
R3719 gnd.n1736 gnd.n1735 585
R3720 gnd.n1744 gnd.n1736 585
R3721 gnd.n5102 gnd.n5101 585
R3722 gnd.n5103 gnd.n5102 585
R3723 gnd.n1753 gnd.n1752 585
R3724 gnd.n1752 gnd.n1749 585
R3725 gnd.n5097 gnd.n5096 585
R3726 gnd.n5096 gnd.n5095 585
R3727 gnd.n1756 gnd.n1755 585
R3728 gnd.n1762 gnd.n1756 585
R3729 gnd.n5077 gnd.n5076 585
R3730 gnd.n5078 gnd.n5077 585
R3731 gnd.n1773 gnd.n1772 585
R3732 gnd.n1780 gnd.n1772 585
R3733 gnd.n5072 gnd.n5071 585
R3734 gnd.n5071 gnd.n5070 585
R3735 gnd.n1776 gnd.n1775 585
R3736 gnd.n1784 gnd.n1776 585
R3737 gnd.n5020 gnd.n5019 585
R3738 gnd.n5021 gnd.n5020 585
R3739 gnd.n1795 gnd.n1794 585
R3740 gnd.n1813 gnd.n1794 585
R3741 gnd.n5015 gnd.n5014 585
R3742 gnd.n5014 gnd.n5013 585
R3743 gnd.n1798 gnd.n1797 585
R3744 gnd.n1806 gnd.n1798 585
R3745 gnd.n4980 gnd.n4979 585
R3746 gnd.n4981 gnd.n4980 585
R3747 gnd.n1818 gnd.n1817 585
R3748 gnd.n1833 gnd.n1817 585
R3749 gnd.n4975 gnd.n4974 585
R3750 gnd.n4974 gnd.n4973 585
R3751 gnd.n1821 gnd.n1820 585
R3752 gnd.n4963 gnd.n1821 585
R3753 gnd.n4930 gnd.n1850 585
R3754 gnd.n1850 gnd.n1842 585
R3755 gnd.n4932 gnd.n4931 585
R3756 gnd.n4933 gnd.n4932 585
R3757 gnd.n1851 gnd.n1849 585
R3758 gnd.n1849 gnd.n1846 585
R3759 gnd.n4925 gnd.n4924 585
R3760 gnd.n4924 gnd.n4923 585
R3761 gnd.n1854 gnd.n1853 585
R3762 gnd.n1860 gnd.n1854 585
R3763 gnd.n4902 gnd.n4901 585
R3764 gnd.n4903 gnd.n4902 585
R3765 gnd.n1869 gnd.n1868 585
R3766 gnd.n1875 gnd.n1868 585
R3767 gnd.n4897 gnd.n4896 585
R3768 gnd.n4896 gnd.n4895 585
R3769 gnd.n1872 gnd.n1871 585
R3770 gnd.n1879 gnd.n1872 585
R3771 gnd.n4840 gnd.n1894 585
R3772 gnd.n1894 gnd.n1884 585
R3773 gnd.n4842 gnd.n4841 585
R3774 gnd.n4843 gnd.n4842 585
R3775 gnd.n1895 gnd.n1893 585
R3776 gnd.n4808 gnd.n1893 585
R3777 gnd.n4835 gnd.n4834 585
R3778 gnd.n4834 gnd.n4833 585
R3779 gnd.n1898 gnd.n1897 585
R3780 gnd.n4816 gnd.n1898 585
R3781 gnd.n4798 gnd.n4797 585
R3782 gnd.n4799 gnd.n4798 585
R3783 gnd.n1913 gnd.n1912 585
R3784 gnd.n4776 gnd.n1912 585
R3785 gnd.n4793 gnd.n4792 585
R3786 gnd.n4792 gnd.n4791 585
R3787 gnd.n1916 gnd.n1915 585
R3788 gnd.n1923 gnd.n1916 585
R3789 gnd.n4755 gnd.n4754 585
R3790 gnd.n4756 gnd.n4755 585
R3791 gnd.n1220 gnd.n1219 585
R3792 gnd.n1937 gnd.n1220 585
R3793 gnd.n6251 gnd.n6250 585
R3794 gnd.n6250 gnd.n6249 585
R3795 gnd.n6252 gnd.n1214 585
R3796 gnd.n1941 gnd.n1214 585
R3797 gnd.n6254 gnd.n6253 585
R3798 gnd.n6255 gnd.n6254 585
R3799 gnd.n1215 gnd.n1213 585
R3800 gnd.n2027 gnd.n1213 585
R3801 gnd.n4717 gnd.n2038 585
R3802 gnd.n2038 gnd.n1184 585
R3803 gnd.n4719 gnd.n4718 585
R3804 gnd.n4720 gnd.n4719 585
R3805 gnd.n2039 gnd.n2037 585
R3806 gnd.n2037 gnd.n2035 585
R3807 gnd.n4711 gnd.n4710 585
R3808 gnd.n4710 gnd.n4709 585
R3809 gnd.n2042 gnd.n2041 585
R3810 gnd.n2051 gnd.n2042 585
R3811 gnd.n4684 gnd.n2063 585
R3812 gnd.n2063 gnd.n2050 585
R3813 gnd.n4686 gnd.n4685 585
R3814 gnd.n4687 gnd.n4686 585
R3815 gnd.n2064 gnd.n2062 585
R3816 gnd.n2062 gnd.n2059 585
R3817 gnd.n4679 gnd.n4678 585
R3818 gnd.n4678 gnd.n4677 585
R3819 gnd.n2067 gnd.n2066 585
R3820 gnd.n2068 gnd.n2067 585
R3821 gnd.n4400 gnd.n4399 585
R3822 gnd.n4401 gnd.n4400 585
R3823 gnd.n2089 gnd.n2088 585
R3824 gnd.n2088 gnd.n2087 585
R3825 gnd.n4395 gnd.n4394 585
R3826 gnd.n4394 gnd.n4393 585
R3827 gnd.n4392 gnd.n2091 585
R3828 gnd.n4392 gnd.n4391 585
R3829 gnd.n4390 gnd.n4389 585
R3830 gnd.n4390 gnd.n1095 585
R3831 gnd.n2093 gnd.n2092 585
R3832 gnd.n2092 gnd.n1092 585
R3833 gnd.n4385 gnd.n4384 585
R3834 gnd.n4384 gnd.n1086 585
R3835 gnd.n4383 gnd.n2095 585
R3836 gnd.n4383 gnd.n1083 585
R3837 gnd.n4382 gnd.n4381 585
R3838 gnd.n4382 gnd.n1075 585
R3839 gnd.n2097 gnd.n2096 585
R3840 gnd.n2096 gnd.n1072 585
R3841 gnd.n4377 gnd.n4376 585
R3842 gnd.n4376 gnd.n1065 585
R3843 gnd.n4375 gnd.n2099 585
R3844 gnd.n4375 gnd.n4374 585
R3845 gnd.n4303 gnd.n2100 585
R3846 gnd.n2100 gnd.n1055 585
R3847 gnd.n4305 gnd.n4304 585
R3848 gnd.n4304 gnd.n1052 585
R3849 gnd.n4306 gnd.n4297 585
R3850 gnd.n4297 gnd.n1045 585
R3851 gnd.n4308 gnd.n4307 585
R3852 gnd.n4308 gnd.n1042 585
R3853 gnd.n4309 gnd.n4296 585
R3854 gnd.n4309 gnd.n2114 585
R3855 gnd.n4311 gnd.n4310 585
R3856 gnd.n4310 gnd.n1032 585
R3857 gnd.n4312 gnd.n2121 585
R3858 gnd.n2121 gnd.n1025 585
R3859 gnd.n4314 gnd.n4313 585
R3860 gnd.n4315 gnd.n4314 585
R3861 gnd.n2122 gnd.n2120 585
R3862 gnd.n2120 gnd.n1015 585
R3863 gnd.n4290 gnd.n4289 585
R3864 gnd.n4289 gnd.n1012 585
R3865 gnd.n4288 gnd.n2124 585
R3866 gnd.n4288 gnd.n1005 585
R3867 gnd.n4287 gnd.n4286 585
R3868 gnd.n4287 gnd.n1002 585
R3869 gnd.n2126 gnd.n2125 585
R3870 gnd.n4253 gnd.n2125 585
R3871 gnd.n4282 gnd.n4281 585
R3872 gnd.n4281 gnd.n993 585
R3873 gnd.n4280 gnd.n2127 585
R3874 gnd.n4280 gnd.n984 585
R3875 gnd.n4279 gnd.n2130 585
R3876 gnd.n4279 gnd.n4278 585
R3877 gnd.n4210 gnd.n2128 585
R3878 gnd.n2131 gnd.n2128 585
R3879 gnd.n4212 gnd.n2169 585
R3880 gnd.n2169 gnd.n2145 585
R3881 gnd.n4214 gnd.n4213 585
R3882 gnd.n4215 gnd.n4214 585
R3883 gnd.n4208 gnd.n2168 585
R3884 gnd.n2168 gnd.n2155 585
R3885 gnd.n4207 gnd.n4206 585
R3886 gnd.n4206 gnd.n2161 585
R3887 gnd.n4205 gnd.n4204 585
R3888 gnd.n4205 gnd.n2159 585
R3889 gnd.n4203 gnd.n2171 585
R3890 gnd.n4177 gnd.n2171 585
R3891 gnd.n4201 gnd.n4200 585
R3892 gnd.n4200 gnd.n968 585
R3893 gnd.n4199 gnd.n2172 585
R3894 gnd.n4199 gnd.n965 585
R3895 gnd.n4198 gnd.n4197 585
R3896 gnd.n4198 gnd.n956 585
R3897 gnd.n4193 gnd.n4192 585
R3898 gnd.n4192 gnd.n4191 585
R3899 gnd.n940 gnd.n939 585
R3900 gnd.n944 gnd.n940 585
R3901 gnd.n6469 gnd.n6468 585
R3902 gnd.n6468 gnd.n6467 585
R3903 gnd.n6140 gnd.n6139 585
R3904 gnd.n6139 gnd.n6138 585
R3905 gnd.n1315 gnd.n1313 585
R3906 gnd.n5541 gnd.n1315 585
R3907 gnd.n6144 gnd.n1312 585
R3908 gnd.n5543 gnd.n1312 585
R3909 gnd.n6145 gnd.n1311 585
R3910 gnd.n1606 gnd.n1311 585
R3911 gnd.n6146 gnd.n1310 585
R3912 gnd.n1593 gnd.n1310 585
R3913 gnd.n5551 gnd.n1308 585
R3914 gnd.n5552 gnd.n5551 585
R3915 gnd.n6150 gnd.n1307 585
R3916 gnd.n5554 gnd.n1307 585
R3917 gnd.n6151 gnd.n1306 585
R3918 gnd.n1590 gnd.n1306 585
R3919 gnd.n6152 gnd.n1305 585
R3920 gnd.n5346 gnd.n1305 585
R3921 gnd.n5343 gnd.n1303 585
R3922 gnd.n5344 gnd.n5343 585
R3923 gnd.n6156 gnd.n1302 585
R3924 gnd.n5563 gnd.n1302 585
R3925 gnd.n6157 gnd.n1301 585
R3926 gnd.n5336 gnd.n1301 585
R3927 gnd.n6158 gnd.n1300 585
R3928 gnd.n1622 gnd.n1300 585
R3929 gnd.n5318 gnd.n1298 585
R3930 gnd.n5319 gnd.n5318 585
R3931 gnd.n6162 gnd.n1297 585
R3932 gnd.n5303 gnd.n1297 585
R3933 gnd.n6163 gnd.n1296 585
R3934 gnd.n1647 gnd.n1296 585
R3935 gnd.n6164 gnd.n1295 585
R3936 gnd.n5294 gnd.n1295 585
R3937 gnd.n1652 gnd.n1293 585
R3938 gnd.n1653 gnd.n1652 585
R3939 gnd.n6168 gnd.n1292 585
R3940 gnd.n5273 gnd.n1292 585
R3941 gnd.n6169 gnd.n1291 585
R3942 gnd.n5260 gnd.n1291 585
R3943 gnd.n6170 gnd.n1290 585
R3944 gnd.n5211 gnd.n1290 585
R3945 gnd.n1680 gnd.n1288 585
R3946 gnd.n1681 gnd.n1680 585
R3947 gnd.n6174 gnd.n1287 585
R3948 gnd.n1676 gnd.n1287 585
R3949 gnd.n6175 gnd.n1286 585
R3950 gnd.n5234 gnd.n1286 585
R3951 gnd.n6176 gnd.n1285 585
R3952 gnd.n5226 gnd.n1285 585
R3953 gnd.n5133 gnd.n1283 585
R3954 gnd.n5134 gnd.n5133 585
R3955 gnd.n6180 gnd.n1282 585
R3956 gnd.n5203 gnd.n1282 585
R3957 gnd.n6181 gnd.n1281 585
R3958 gnd.n5195 gnd.n1281 585
R3959 gnd.n6182 gnd.n1280 585
R3960 gnd.n1716 gnd.n1280 585
R3961 gnd.n5173 gnd.n1278 585
R3962 gnd.n5174 gnd.n5173 585
R3963 gnd.n6186 gnd.n1277 585
R3964 gnd.n1720 gnd.n1277 585
R3965 gnd.n6187 gnd.n1276 585
R3966 gnd.n5164 gnd.n1276 585
R3967 gnd.n6188 gnd.n1275 585
R3968 gnd.n1738 gnd.n1275 585
R3969 gnd.n5042 gnd.n1273 585
R3970 gnd.n5043 gnd.n5042 585
R3971 gnd.n6192 gnd.n1272 585
R3972 gnd.n1743 gnd.n1272 585
R3973 gnd.n6193 gnd.n1271 585
R3974 gnd.n5105 gnd.n1271 585
R3975 gnd.n6194 gnd.n1270 585
R3976 gnd.n5094 gnd.n1270 585
R3977 gnd.n1763 gnd.n1268 585
R3978 gnd.n1764 gnd.n1763 585
R3979 gnd.n6198 gnd.n1267 585
R3980 gnd.n1771 gnd.n1267 585
R3981 gnd.n6199 gnd.n1266 585
R3982 gnd.n5034 gnd.n1266 585
R3983 gnd.n6200 gnd.n1265 585
R3984 gnd.n5069 gnd.n1265 585
R3985 gnd.n5060 gnd.n1263 585
R3986 gnd.n5061 gnd.n5060 585
R3987 gnd.n6204 gnd.n1262 585
R3988 gnd.n5022 gnd.n1262 585
R3989 gnd.n6205 gnd.n1261 585
R3990 gnd.n4993 gnd.n1261 585
R3991 gnd.n6206 gnd.n1260 585
R3992 gnd.n1801 gnd.n1260 585
R3993 gnd.n5001 gnd.n1258 585
R3994 gnd.n5002 gnd.n5001 585
R3995 gnd.n6210 gnd.n1257 585
R3996 gnd.n4982 gnd.n1257 585
R3997 gnd.n6211 gnd.n1256 585
R3998 gnd.n4955 gnd.n1256 585
R3999 gnd.n6212 gnd.n1255 585
R4000 gnd.n1824 gnd.n1255 585
R4001 gnd.n4946 gnd.n1253 585
R4002 gnd.n4947 gnd.n4946 585
R4003 gnd.n6216 gnd.n1252 585
R4004 gnd.n1829 gnd.n1252 585
R4005 gnd.n6217 gnd.n1251 585
R4006 gnd.n4943 gnd.n1251 585
R4007 gnd.n6218 gnd.n1250 585
R4008 gnd.n4935 gnd.n1250 585
R4009 gnd.n4921 gnd.n1248 585
R4010 gnd.n4922 gnd.n4921 585
R4011 gnd.n6222 gnd.n1247 585
R4012 gnd.n1861 gnd.n1247 585
R4013 gnd.n6223 gnd.n1246 585
R4014 gnd.n4853 gnd.n1246 585
R4015 gnd.n6224 gnd.n1245 585
R4016 gnd.n1866 gnd.n1245 585
R4017 gnd.n4893 gnd.n1243 585
R4018 gnd.n4894 gnd.n4893 585
R4019 gnd.n6228 gnd.n1242 585
R4020 gnd.n4885 gnd.n1242 585
R4021 gnd.n6229 gnd.n1241 585
R4022 gnd.n4872 gnd.n1241 585
R4023 gnd.n6230 gnd.n1240 585
R4024 gnd.n4823 gnd.n1240 585
R4025 gnd.n4844 gnd.n1238 585
R4026 gnd.n4845 gnd.n4844 585
R4027 gnd.n6234 gnd.n1237 585
R4028 gnd.n1901 gnd.n1237 585
R4029 gnd.n6235 gnd.n1236 585
R4030 gnd.n1899 gnd.n1236 585
R4031 gnd.n6236 gnd.n1235 585
R4032 gnd.n1906 gnd.n1235 585
R4033 gnd.n1910 gnd.n1233 585
R4034 gnd.n1911 gnd.n1910 585
R4035 gnd.n6240 gnd.n1232 585
R4036 gnd.n4774 gnd.n1232 585
R4037 gnd.n6241 gnd.n1231 585
R4038 gnd.n1930 gnd.n1231 585
R4039 gnd.n6242 gnd.n1230 585
R4040 gnd.n1922 gnd.n1230 585
R4041 gnd.n1227 gnd.n1225 585
R4042 gnd.n4758 gnd.n1225 585
R4043 gnd.n6247 gnd.n6246 585
R4044 gnd.n6248 gnd.n6247 585
R4045 gnd.n1226 gnd.n1224 585
R4046 gnd.n4743 gnd.n1224 585
R4047 gnd.n4727 gnd.n4726 585
R4048 gnd.n4726 gnd.n1212 585
R4049 gnd.n2031 gnd.n2029 585
R4050 gnd.n2029 gnd.n1210 585
R4051 gnd.n4732 gnd.n4731 585
R4052 gnd.n4733 gnd.n4732 585
R4053 gnd.n2030 gnd.n2028 585
R4054 gnd.n2028 gnd.n1152 585
R4055 gnd.n4723 gnd.n4722 585
R4056 gnd.n4722 gnd.n4721 585
R4057 gnd.n2034 gnd.n2033 585
R4058 gnd.n4708 gnd.n2034 585
R4059 gnd.n2055 gnd.n2053 585
R4060 gnd.n2053 gnd.n2043 585
R4061 gnd.n4696 gnd.n4695 585
R4062 gnd.n4697 gnd.n4696 585
R4063 gnd.n2054 gnd.n2052 585
R4064 gnd.n2061 gnd.n2052 585
R4065 gnd.n4690 gnd.n4689 585
R4066 gnd.n4689 gnd.n4688 585
R4067 gnd.n2058 gnd.n2057 585
R4068 gnd.n4676 gnd.n2058 585
R4069 gnd.n4653 gnd.n4652 585
R4070 gnd.n4651 gnd.n4415 585
R4071 gnd.n4417 gnd.n4414 585
R4072 gnd.n4655 gnd.n4414 585
R4073 gnd.n4647 gnd.n4419 585
R4074 gnd.n4646 gnd.n4420 585
R4075 gnd.n4645 gnd.n4421 585
R4076 gnd.n4537 gnd.n4422 585
R4077 gnd.n4640 gnd.n4538 585
R4078 gnd.n4639 gnd.n4539 585
R4079 gnd.n4638 gnd.n4540 585
R4080 gnd.n4550 gnd.n4541 585
R4081 gnd.n4631 gnd.n4551 585
R4082 gnd.n4630 gnd.n4552 585
R4083 gnd.n4554 gnd.n4553 585
R4084 gnd.n4623 gnd.n4562 585
R4085 gnd.n4622 gnd.n4563 585
R4086 gnd.n4573 gnd.n4564 585
R4087 gnd.n4615 gnd.n4574 585
R4088 gnd.n4614 gnd.n4575 585
R4089 gnd.n4577 gnd.n4576 585
R4090 gnd.n4607 gnd.n4585 585
R4091 gnd.n4606 gnd.n4586 585
R4092 gnd.n4596 gnd.n4587 585
R4093 gnd.n4599 gnd.n4597 585
R4094 gnd.n4598 gnd.n2085 585
R4095 gnd.n4658 gnd.n4657 585
R4096 gnd.n2086 gnd.n2072 585
R4097 gnd.n4669 gnd.n2073 585
R4098 gnd.n4670 gnd.n2069 585
R4099 gnd.n1609 gnd.n1318 585
R4100 gnd.n6138 gnd.n1318 585
R4101 gnd.n5540 gnd.n5539 585
R4102 gnd.n5541 gnd.n5540 585
R4103 gnd.n1608 gnd.n1607 585
R4104 gnd.n5543 gnd.n1607 585
R4105 gnd.n5357 gnd.n5356 585
R4106 gnd.n5356 gnd.n1606 585
R4107 gnd.n5355 gnd.n5354 585
R4108 gnd.n5355 gnd.n1593 585
R4109 gnd.n5353 gnd.n1592 585
R4110 gnd.n5552 gnd.n1592 585
R4111 gnd.n1611 gnd.n1591 585
R4112 gnd.n5554 gnd.n1591 585
R4113 gnd.n5349 gnd.n5348 585
R4114 gnd.n5348 gnd.n1590 585
R4115 gnd.n5347 gnd.n1613 585
R4116 gnd.n5347 gnd.n5346 585
R4117 gnd.n5345 gnd.n5342 585
R4118 gnd.n5345 gnd.n5344 585
R4119 gnd.n1614 gnd.n1580 585
R4120 gnd.n5563 gnd.n1580 585
R4121 gnd.n5338 gnd.n5337 585
R4122 gnd.n5337 gnd.n5336 585
R4123 gnd.n1617 gnd.n1616 585
R4124 gnd.n1622 gnd.n1617 585
R4125 gnd.n1641 gnd.n1629 585
R4126 gnd.n5319 gnd.n1629 585
R4127 gnd.n5302 gnd.n5301 585
R4128 gnd.n5303 gnd.n5302 585
R4129 gnd.n1640 gnd.n1639 585
R4130 gnd.n1647 gnd.n1639 585
R4131 gnd.n5296 gnd.n5295 585
R4132 gnd.n5295 gnd.n5294 585
R4133 gnd.n1644 gnd.n1643 585
R4134 gnd.n1653 gnd.n1644 585
R4135 gnd.n5214 gnd.n1660 585
R4136 gnd.n5273 gnd.n1660 585
R4137 gnd.n5213 gnd.n1668 585
R4138 gnd.n5260 gnd.n1668 585
R4139 gnd.n5218 gnd.n5212 585
R4140 gnd.n5212 gnd.n5211 585
R4141 gnd.n5219 gnd.n5210 585
R4142 gnd.n5210 gnd.n1681 585
R4143 gnd.n5220 gnd.n5209 585
R4144 gnd.n5209 gnd.n1676 585
R4145 gnd.n1697 gnd.n1688 585
R4146 gnd.n5234 gnd.n1688 585
R4147 gnd.n5225 gnd.n5224 585
R4148 gnd.n5226 gnd.n5225 585
R4149 gnd.n1696 gnd.n1695 585
R4150 gnd.n5134 gnd.n1695 585
R4151 gnd.n5205 gnd.n5204 585
R4152 gnd.n5204 gnd.n5203 585
R4153 gnd.n1700 gnd.n1699 585
R4154 gnd.n5195 gnd.n1700 585
R4155 gnd.n1726 gnd.n1724 585
R4156 gnd.n1724 gnd.n1716 585
R4157 gnd.n5172 gnd.n5171 585
R4158 gnd.n5174 gnd.n5172 585
R4159 gnd.n1725 gnd.n1723 585
R4160 gnd.n1723 gnd.n1720 585
R4161 gnd.n5166 gnd.n5165 585
R4162 gnd.n5165 gnd.n5164 585
R4163 gnd.n1729 gnd.n1728 585
R4164 gnd.n1738 gnd.n1729 585
R4165 gnd.n5046 gnd.n5044 585
R4166 gnd.n5044 gnd.n5043 585
R4167 gnd.n5047 gnd.n5040 585
R4168 gnd.n5040 gnd.n1743 585
R4169 gnd.n5048 gnd.n1751 585
R4170 gnd.n5105 gnd.n1751 585
R4171 gnd.n5038 gnd.n1758 585
R4172 gnd.n5094 gnd.n1758 585
R4173 gnd.n5052 gnd.n5037 585
R4174 gnd.n5037 gnd.n1764 585
R4175 gnd.n5053 gnd.n5036 585
R4176 gnd.n5036 gnd.n1771 585
R4177 gnd.n5054 gnd.n5035 585
R4178 gnd.n5035 gnd.n5034 585
R4179 gnd.n1788 gnd.n1778 585
R4180 gnd.n5069 gnd.n1778 585
R4181 gnd.n5059 gnd.n5058 585
R4182 gnd.n5061 gnd.n5059 585
R4183 gnd.n1787 gnd.n1786 585
R4184 gnd.n5022 gnd.n1786 585
R4185 gnd.n4995 gnd.n4994 585
R4186 gnd.n4994 gnd.n4993 585
R4187 gnd.n1811 gnd.n1809 585
R4188 gnd.n1809 gnd.n1801 585
R4189 gnd.n5000 gnd.n4999 585
R4190 gnd.n5002 gnd.n5000 585
R4191 gnd.n1810 gnd.n1808 585
R4192 gnd.n4982 gnd.n1808 585
R4193 gnd.n4954 gnd.n4953 585
R4194 gnd.n4955 gnd.n4954 585
R4195 gnd.n1835 gnd.n1834 585
R4196 gnd.n1834 gnd.n1824 585
R4197 gnd.n4949 gnd.n4948 585
R4198 gnd.n4948 gnd.n4947 585
R4199 gnd.n4945 gnd.n1837 585
R4200 gnd.n4945 gnd.n1829 585
R4201 gnd.n4944 gnd.n1839 585
R4202 gnd.n4944 gnd.n4943 585
R4203 gnd.n4859 gnd.n1838 585
R4204 gnd.n4935 gnd.n1838 585
R4205 gnd.n4860 gnd.n1856 585
R4206 gnd.n4922 gnd.n1856 585
R4207 gnd.n4856 gnd.n4855 585
R4208 gnd.n4855 gnd.n1861 585
R4209 gnd.n4864 gnd.n4854 585
R4210 gnd.n4854 gnd.n4853 585
R4211 gnd.n4865 gnd.n4851 585
R4212 gnd.n4851 gnd.n1866 585
R4213 gnd.n4866 gnd.n1873 585
R4214 gnd.n4894 gnd.n1873 585
R4215 gnd.n1887 gnd.n1881 585
R4216 gnd.n4885 gnd.n1881 585
R4217 gnd.n4871 gnd.n4870 585
R4218 gnd.n4872 gnd.n4871 585
R4219 gnd.n1886 gnd.n1885 585
R4220 gnd.n4823 gnd.n1885 585
R4221 gnd.n4847 gnd.n4846 585
R4222 gnd.n4846 gnd.n4845 585
R4223 gnd.n1890 gnd.n1889 585
R4224 gnd.n1901 gnd.n1890 585
R4225 gnd.n4767 gnd.n4766 585
R4226 gnd.n4766 gnd.n1899 585
R4227 gnd.n4768 gnd.n4765 585
R4228 gnd.n4765 gnd.n1906 585
R4229 gnd.n1934 gnd.n1932 585
R4230 gnd.n1932 gnd.n1911 585
R4231 gnd.n4773 gnd.n4772 585
R4232 gnd.n4774 gnd.n4773 585
R4233 gnd.n1933 gnd.n1931 585
R4234 gnd.n1931 gnd.n1930 585
R4235 gnd.n4761 gnd.n4760 585
R4236 gnd.n4760 gnd.n1922 585
R4237 gnd.n4759 gnd.n1936 585
R4238 gnd.n4759 gnd.n4758 585
R4239 gnd.n1945 gnd.n1222 585
R4240 gnd.n6248 gnd.n1222 585
R4241 gnd.n4742 gnd.n4741 585
R4242 gnd.n4743 gnd.n4742 585
R4243 gnd.n1944 gnd.n1943 585
R4244 gnd.n1943 gnd.n1212 585
R4245 gnd.n4736 gnd.n4735 585
R4246 gnd.n4735 gnd.n1210 585
R4247 gnd.n4734 gnd.n1947 585
R4248 gnd.n4734 gnd.n4733 585
R4249 gnd.n4702 gnd.n1948 585
R4250 gnd.n1948 gnd.n1152 585
R4251 gnd.n2046 gnd.n2036 585
R4252 gnd.n4721 gnd.n2036 585
R4253 gnd.n4707 gnd.n4706 585
R4254 gnd.n4708 gnd.n4707 585
R4255 gnd.n2045 gnd.n2044 585
R4256 gnd.n2044 gnd.n2043 585
R4257 gnd.n4699 gnd.n4698 585
R4258 gnd.n4698 gnd.n4697 585
R4259 gnd.n2049 gnd.n2048 585
R4260 gnd.n2061 gnd.n2049 585
R4261 gnd.n2070 gnd.n2060 585
R4262 gnd.n4688 gnd.n2060 585
R4263 gnd.n4675 gnd.n4674 585
R4264 gnd.n4676 gnd.n4675 585
R4265 gnd.n5514 gnd.n5369 585
R4266 gnd.n5369 gnd.n1328 585
R4267 gnd.n5515 gnd.n5512 585
R4268 gnd.n5510 gnd.n5387 585
R4269 gnd.n5509 gnd.n5508 585
R4270 gnd.n5493 gnd.n5389 585
R4271 gnd.n5495 gnd.n5494 585
R4272 gnd.n5491 gnd.n5396 585
R4273 gnd.n5490 gnd.n5489 585
R4274 gnd.n5474 gnd.n5398 585
R4275 gnd.n5476 gnd.n5475 585
R4276 gnd.n5472 gnd.n5405 585
R4277 gnd.n5471 gnd.n5470 585
R4278 gnd.n5455 gnd.n5407 585
R4279 gnd.n5457 gnd.n5456 585
R4280 gnd.n5453 gnd.n5414 585
R4281 gnd.n5452 gnd.n5451 585
R4282 gnd.n5440 gnd.n5416 585
R4283 gnd.n5442 gnd.n5441 585
R4284 gnd.n5438 gnd.n5417 585
R4285 gnd.n5437 gnd.n5436 585
R4286 gnd.n5429 gnd.n5419 585
R4287 gnd.n5431 gnd.n5430 585
R4288 gnd.n5427 gnd.n5421 585
R4289 gnd.n5426 gnd.n5425 585
R4290 gnd.n5423 gnd.n1316 585
R4291 gnd.n5535 gnd.n5534 585
R4292 gnd.n5532 gnd.n5367 585
R4293 gnd.n5531 gnd.n5368 585
R4294 gnd.n5529 gnd.n5528 585
R4295 gnd.n6645 gnd.n769 493.813
R4296 gnd.n5653 gnd.n1575 482.89
R4297 gnd.n5656 gnd.n5655 482.89
R4298 gnd.n2025 gnd.n1949 482.89
R4299 gnd.n6324 gnd.n1187 482.89
R4300 gnd.n1950 gnd.t198 443.966
R4301 gnd.n1569 gnd.t221 443.966
R4302 gnd.n6261 gnd.t246 443.966
R4303 gnd.n5587 gnd.t151 443.966
R4304 gnd.n2082 gnd.t188 371.625
R4305 gnd.n5380 gnd.t215 371.625
R4306 gnd.n2075 gnd.t240 371.625
R4307 gnd.n5793 gnd.t212 371.625
R4308 gnd.n5845 gnd.t209 371.625
R4309 gnd.n1500 gnd.t140 371.625
R4310 gnd.n311 gnd.t237 371.625
R4311 gnd.n278 gnd.t155 371.625
R4312 gnd.n7527 gnd.t195 371.625
R4313 gnd.n348 gnd.t182 371.625
R4314 gnd.n3807 gnd.t169 371.625
R4315 gnd.n3829 gnd.t166 371.625
R4316 gnd.n3850 gnd.t144 371.625
R4317 gnd.n3868 gnd.t224 371.625
R4318 gnd.n1128 gnd.t230 371.625
R4319 gnd.n4424 gnd.t162 371.625
R4320 gnd.n4446 gnd.t185 371.625
R4321 gnd.n5370 gnd.t172 371.625
R4322 gnd.n2769 gnd.t202 323.425
R4323 gnd.n2311 gnd.t233 323.425
R4324 gnd.n3617 gnd.n3591 289.615
R4325 gnd.n3585 gnd.n3559 289.615
R4326 gnd.n3553 gnd.n3527 289.615
R4327 gnd.n3522 gnd.n3496 289.615
R4328 gnd.n3490 gnd.n3464 289.615
R4329 gnd.n3458 gnd.n3432 289.615
R4330 gnd.n3426 gnd.n3400 289.615
R4331 gnd.n3395 gnd.n3369 289.615
R4332 gnd.n2843 gnd.t136 279.217
R4333 gnd.n2337 gnd.t132 279.217
R4334 gnd.n1194 gnd.t229 260.649
R4335 gnd.n5579 gnd.t150 260.649
R4336 gnd.n6326 gnd.n6325 256.663
R4337 gnd.n6326 gnd.n1153 256.663
R4338 gnd.n6326 gnd.n1154 256.663
R4339 gnd.n6326 gnd.n1155 256.663
R4340 gnd.n6326 gnd.n1156 256.663
R4341 gnd.n6326 gnd.n1157 256.663
R4342 gnd.n6326 gnd.n1158 256.663
R4343 gnd.n6326 gnd.n1159 256.663
R4344 gnd.n6326 gnd.n1160 256.663
R4345 gnd.n6326 gnd.n1161 256.663
R4346 gnd.n6326 gnd.n1162 256.663
R4347 gnd.n6326 gnd.n1163 256.663
R4348 gnd.n6326 gnd.n1164 256.663
R4349 gnd.n6326 gnd.n1165 256.663
R4350 gnd.n6326 gnd.n1166 256.663
R4351 gnd.n6326 gnd.n1167 256.663
R4352 gnd.n6329 gnd.n1150 256.663
R4353 gnd.n6327 gnd.n6326 256.663
R4354 gnd.n6326 gnd.n1168 256.663
R4355 gnd.n6326 gnd.n1169 256.663
R4356 gnd.n6326 gnd.n1170 256.663
R4357 gnd.n6326 gnd.n1171 256.663
R4358 gnd.n6326 gnd.n1172 256.663
R4359 gnd.n6326 gnd.n1173 256.663
R4360 gnd.n6326 gnd.n1174 256.663
R4361 gnd.n6326 gnd.n1175 256.663
R4362 gnd.n6326 gnd.n1176 256.663
R4363 gnd.n6326 gnd.n1177 256.663
R4364 gnd.n6326 gnd.n1178 256.663
R4365 gnd.n6326 gnd.n1179 256.663
R4366 gnd.n6326 gnd.n1180 256.663
R4367 gnd.n6326 gnd.n1181 256.663
R4368 gnd.n6326 gnd.n1182 256.663
R4369 gnd.n6326 gnd.n1183 256.663
R4370 gnd.n5721 gnd.n1553 256.663
R4371 gnd.n5721 gnd.n1554 256.663
R4372 gnd.n5721 gnd.n1555 256.663
R4373 gnd.n5721 gnd.n1556 256.663
R4374 gnd.n5721 gnd.n1557 256.663
R4375 gnd.n5721 gnd.n1558 256.663
R4376 gnd.n5721 gnd.n1559 256.663
R4377 gnd.n5721 gnd.n1560 256.663
R4378 gnd.n5721 gnd.n1561 256.663
R4379 gnd.n5721 gnd.n1562 256.663
R4380 gnd.n5721 gnd.n1563 256.663
R4381 gnd.n5721 gnd.n1564 256.663
R4382 gnd.n5721 gnd.n1565 256.663
R4383 gnd.n5721 gnd.n1566 256.663
R4384 gnd.n5721 gnd.n1567 256.663
R4385 gnd.n5721 gnd.n5718 256.663
R4386 gnd.n5724 gnd.n1534 256.663
R4387 gnd.n5722 gnd.n5721 256.663
R4388 gnd.n5721 gnd.n1552 256.663
R4389 gnd.n5721 gnd.n1551 256.663
R4390 gnd.n5721 gnd.n1550 256.663
R4391 gnd.n5721 gnd.n1549 256.663
R4392 gnd.n5721 gnd.n1548 256.663
R4393 gnd.n5721 gnd.n1547 256.663
R4394 gnd.n5721 gnd.n1546 256.663
R4395 gnd.n5721 gnd.n1545 256.663
R4396 gnd.n5721 gnd.n1544 256.663
R4397 gnd.n5721 gnd.n1543 256.663
R4398 gnd.n5721 gnd.n1542 256.663
R4399 gnd.n5721 gnd.n1541 256.663
R4400 gnd.n5721 gnd.n1540 256.663
R4401 gnd.n5721 gnd.n1539 256.663
R4402 gnd.n5721 gnd.n1538 256.663
R4403 gnd.n5721 gnd.n1537 256.663
R4404 gnd.n4043 gnd.n3777 242.672
R4405 gnd.n4043 gnd.n3778 242.672
R4406 gnd.n4043 gnd.n3779 242.672
R4407 gnd.n4043 gnd.n3780 242.672
R4408 gnd.n4043 gnd.n3781 242.672
R4409 gnd.n4043 gnd.n3782 242.672
R4410 gnd.n4043 gnd.n3783 242.672
R4411 gnd.n4043 gnd.n3784 242.672
R4412 gnd.n4043 gnd.n3785 242.672
R4413 gnd.n4664 gnd.n1100 242.672
R4414 gnd.n2078 gnd.n1100 242.672
R4415 gnd.n4592 gnd.n1100 242.672
R4416 gnd.n4589 gnd.n1100 242.672
R4417 gnd.n4580 gnd.n1100 242.672
R4418 gnd.n4569 gnd.n1100 242.672
R4419 gnd.n4566 gnd.n1100 242.672
R4420 gnd.n4557 gnd.n1100 242.672
R4421 gnd.n4546 gnd.n1100 242.672
R4422 gnd.n2897 gnd.n2896 242.672
R4423 gnd.n2897 gnd.n2807 242.672
R4424 gnd.n2897 gnd.n2808 242.672
R4425 gnd.n2897 gnd.n2809 242.672
R4426 gnd.n2897 gnd.n2810 242.672
R4427 gnd.n2897 gnd.n2811 242.672
R4428 gnd.n2897 gnd.n2812 242.672
R4429 gnd.n2897 gnd.n2813 242.672
R4430 gnd.n2897 gnd.n2814 242.672
R4431 gnd.n2897 gnd.n2815 242.672
R4432 gnd.n2897 gnd.n2816 242.672
R4433 gnd.n2897 gnd.n2817 242.672
R4434 gnd.n2898 gnd.n2897 242.672
R4435 gnd.n3749 gnd.n2286 242.672
R4436 gnd.n3749 gnd.n2285 242.672
R4437 gnd.n3749 gnd.n2284 242.672
R4438 gnd.n3749 gnd.n2283 242.672
R4439 gnd.n3749 gnd.n2282 242.672
R4440 gnd.n3749 gnd.n2281 242.672
R4441 gnd.n3749 gnd.n2280 242.672
R4442 gnd.n3749 gnd.n2279 242.672
R4443 gnd.n3749 gnd.n2278 242.672
R4444 gnd.n3749 gnd.n2277 242.672
R4445 gnd.n3749 gnd.n2276 242.672
R4446 gnd.n3749 gnd.n2275 242.672
R4447 gnd.n3749 gnd.n2274 242.672
R4448 gnd.n5445 gnd.n1329 242.672
R4449 gnd.n5462 gnd.n1329 242.672
R4450 gnd.n5464 gnd.n1329 242.672
R4451 gnd.n5481 gnd.n1329 242.672
R4452 gnd.n5483 gnd.n1329 242.672
R4453 gnd.n5500 gnd.n1329 242.672
R4454 gnd.n5502 gnd.n1329 242.672
R4455 gnd.n5520 gnd.n1329 242.672
R4456 gnd.n5522 gnd.n1329 242.672
R4457 gnd.n345 gnd.n210 242.672
R4458 gnd.n7423 gnd.n210 242.672
R4459 gnd.n341 gnd.n210 242.672
R4460 gnd.n7430 gnd.n210 242.672
R4461 gnd.n334 gnd.n210 242.672
R4462 gnd.n7437 gnd.n210 242.672
R4463 gnd.n327 gnd.n210 242.672
R4464 gnd.n7444 gnd.n210 242.672
R4465 gnd.n320 gnd.n210 242.672
R4466 gnd.n2981 gnd.n2980 242.672
R4467 gnd.n2980 gnd.n2719 242.672
R4468 gnd.n2980 gnd.n2720 242.672
R4469 gnd.n2980 gnd.n2721 242.672
R4470 gnd.n2980 gnd.n2722 242.672
R4471 gnd.n2980 gnd.n2723 242.672
R4472 gnd.n2980 gnd.n2724 242.672
R4473 gnd.n2980 gnd.n2725 242.672
R4474 gnd.n3749 gnd.n2287 242.672
R4475 gnd.n3749 gnd.n2288 242.672
R4476 gnd.n3749 gnd.n2289 242.672
R4477 gnd.n3749 gnd.n2290 242.672
R4478 gnd.n3749 gnd.n2291 242.672
R4479 gnd.n3749 gnd.n2292 242.672
R4480 gnd.n3749 gnd.n2293 242.672
R4481 gnd.n3749 gnd.n2294 242.672
R4482 gnd.n4043 gnd.n4042 242.672
R4483 gnd.n4043 gnd.n3750 242.672
R4484 gnd.n4043 gnd.n3751 242.672
R4485 gnd.n4043 gnd.n3752 242.672
R4486 gnd.n4043 gnd.n3753 242.672
R4487 gnd.n4043 gnd.n3754 242.672
R4488 gnd.n4043 gnd.n3755 242.672
R4489 gnd.n4043 gnd.n3756 242.672
R4490 gnd.n4043 gnd.n3757 242.672
R4491 gnd.n4043 gnd.n3758 242.672
R4492 gnd.n4043 gnd.n3759 242.672
R4493 gnd.n4043 gnd.n3760 242.672
R4494 gnd.n4043 gnd.n3761 242.672
R4495 gnd.n4043 gnd.n3762 242.672
R4496 gnd.n4043 gnd.n3763 242.672
R4497 gnd.n4043 gnd.n3764 242.672
R4498 gnd.n4043 gnd.n3765 242.672
R4499 gnd.n4043 gnd.n3766 242.672
R4500 gnd.n4043 gnd.n3767 242.672
R4501 gnd.n4043 gnd.n3768 242.672
R4502 gnd.n4043 gnd.n3769 242.672
R4503 gnd.n4043 gnd.n3770 242.672
R4504 gnd.n4043 gnd.n3771 242.672
R4505 gnd.n4043 gnd.n3772 242.672
R4506 gnd.n4043 gnd.n3773 242.672
R4507 gnd.n4043 gnd.n3774 242.672
R4508 gnd.n4043 gnd.n3775 242.672
R4509 gnd.n4043 gnd.n3776 242.672
R4510 gnd.n4044 gnd.n4043 242.672
R4511 gnd.n4531 gnd.n1100 242.672
R4512 gnd.n4427 gnd.n1100 242.672
R4513 gnd.n4521 gnd.n1100 242.672
R4514 gnd.n4431 gnd.n1100 242.672
R4515 gnd.n4511 gnd.n1100 242.672
R4516 gnd.n4435 gnd.n1100 242.672
R4517 gnd.n4501 gnd.n1100 242.672
R4518 gnd.n4439 gnd.n1100 242.672
R4519 gnd.n4491 gnd.n1100 242.672
R4520 gnd.n4443 gnd.n1100 242.672
R4521 gnd.n4481 gnd.n1100 242.672
R4522 gnd.n4449 gnd.n1100 242.672
R4523 gnd.n4471 gnd.n1100 242.672
R4524 gnd.n4453 gnd.n1100 242.672
R4525 gnd.n4461 gnd.n1100 242.672
R4526 gnd.n4458 gnd.n1100 242.672
R4527 gnd.n6330 gnd.n1146 242.672
R4528 gnd.n1145 gnd.n1100 242.672
R4529 gnd.n6334 gnd.n1100 242.672
R4530 gnd.n1139 gnd.n1100 242.672
R4531 gnd.n6341 gnd.n1100 242.672
R4532 gnd.n1132 gnd.n1100 242.672
R4533 gnd.n6349 gnd.n1100 242.672
R4534 gnd.n1123 gnd.n1100 242.672
R4535 gnd.n6356 gnd.n1100 242.672
R4536 gnd.n1116 gnd.n1100 242.672
R4537 gnd.n6363 gnd.n1100 242.672
R4538 gnd.n1109 gnd.n1100 242.672
R4539 gnd.n6370 gnd.n1100 242.672
R4540 gnd.n6373 gnd.n1100 242.672
R4541 gnd.n5754 gnd.n1329 242.672
R4542 gnd.n5757 gnd.n1329 242.672
R4543 gnd.n5765 gnd.n1329 242.672
R4544 gnd.n5767 gnd.n1329 242.672
R4545 gnd.n5775 gnd.n1329 242.672
R4546 gnd.n5777 gnd.n1329 242.672
R4547 gnd.n5785 gnd.n1329 242.672
R4548 gnd.n5787 gnd.n1329 242.672
R4549 gnd.n5798 gnd.n1329 242.672
R4550 gnd.n5800 gnd.n1329 242.672
R4551 gnd.n5808 gnd.n1329 242.672
R4552 gnd.n5810 gnd.n1329 242.672
R4553 gnd.n5819 gnd.n1329 242.672
R4554 gnd.n5820 gnd.n5725 242.672
R4555 gnd.n5821 gnd.n1329 242.672
R4556 gnd.n5823 gnd.n1329 242.672
R4557 gnd.n5831 gnd.n1329 242.672
R4558 gnd.n5833 gnd.n1329 242.672
R4559 gnd.n5841 gnd.n1329 242.672
R4560 gnd.n5843 gnd.n1329 242.672
R4561 gnd.n5853 gnd.n1329 242.672
R4562 gnd.n5855 gnd.n1329 242.672
R4563 gnd.n5863 gnd.n1329 242.672
R4564 gnd.n5865 gnd.n1329 242.672
R4565 gnd.n5873 gnd.n1329 242.672
R4566 gnd.n5875 gnd.n1329 242.672
R4567 gnd.n5883 gnd.n1329 242.672
R4568 gnd.n5885 gnd.n1329 242.672
R4569 gnd.n5894 gnd.n1329 242.672
R4570 gnd.n5897 gnd.n1329 242.672
R4571 gnd.n7455 gnd.n210 242.672
R4572 gnd.n314 gnd.n210 242.672
R4573 gnd.n7462 gnd.n210 242.672
R4574 gnd.n305 gnd.n210 242.672
R4575 gnd.n7469 gnd.n210 242.672
R4576 gnd.n298 gnd.n210 242.672
R4577 gnd.n7476 gnd.n210 242.672
R4578 gnd.n291 gnd.n210 242.672
R4579 gnd.n7483 gnd.n210 242.672
R4580 gnd.n7486 gnd.n210 242.672
R4581 gnd.n282 gnd.n210 242.672
R4582 gnd.n7495 gnd.n210 242.672
R4583 gnd.n273 gnd.n210 242.672
R4584 gnd.n7502 gnd.n210 242.672
R4585 gnd.n266 gnd.n210 242.672
R4586 gnd.n7509 gnd.n210 242.672
R4587 gnd.n259 gnd.n210 242.672
R4588 gnd.n7516 gnd.n210 242.672
R4589 gnd.n252 gnd.n210 242.672
R4590 gnd.n7523 gnd.n210 242.672
R4591 gnd.n245 gnd.n210 242.672
R4592 gnd.n7533 gnd.n210 242.672
R4593 gnd.n238 gnd.n210 242.672
R4594 gnd.n7540 gnd.n210 242.672
R4595 gnd.n231 gnd.n210 242.672
R4596 gnd.n7547 gnd.n210 242.672
R4597 gnd.n224 gnd.n210 242.672
R4598 gnd.n7554 gnd.n210 242.672
R4599 gnd.n217 gnd.n210 242.672
R4600 gnd.n4655 gnd.n4654 242.672
R4601 gnd.n4655 gnd.n4402 242.672
R4602 gnd.n4655 gnd.n4403 242.672
R4603 gnd.n4655 gnd.n4404 242.672
R4604 gnd.n4655 gnd.n4405 242.672
R4605 gnd.n4655 gnd.n4406 242.672
R4606 gnd.n4655 gnd.n4407 242.672
R4607 gnd.n4655 gnd.n4408 242.672
R4608 gnd.n4655 gnd.n4409 242.672
R4609 gnd.n4655 gnd.n4410 242.672
R4610 gnd.n4655 gnd.n4411 242.672
R4611 gnd.n4655 gnd.n4412 242.672
R4612 gnd.n4656 gnd.n4655 242.672
R4613 gnd.n4655 gnd.n4413 242.672
R4614 gnd.n5511 gnd.n1328 242.672
R4615 gnd.n5388 gnd.n1328 242.672
R4616 gnd.n5492 gnd.n1328 242.672
R4617 gnd.n5397 gnd.n1328 242.672
R4618 gnd.n5473 gnd.n1328 242.672
R4619 gnd.n5406 gnd.n1328 242.672
R4620 gnd.n5454 gnd.n1328 242.672
R4621 gnd.n5415 gnd.n1328 242.672
R4622 gnd.n5439 gnd.n1328 242.672
R4623 gnd.n5418 gnd.n1328 242.672
R4624 gnd.n5428 gnd.n1328 242.672
R4625 gnd.n5422 gnd.n1328 242.672
R4626 gnd.n5533 gnd.n1328 242.672
R4627 gnd.n5530 gnd.n1328 242.672
R4628 gnd.n214 gnd.n211 240.244
R4629 gnd.n7556 gnd.n7555 240.244
R4630 gnd.n7553 gnd.n218 240.244
R4631 gnd.n7549 gnd.n7548 240.244
R4632 gnd.n7546 gnd.n225 240.244
R4633 gnd.n7542 gnd.n7541 240.244
R4634 gnd.n7539 gnd.n232 240.244
R4635 gnd.n7535 gnd.n7534 240.244
R4636 gnd.n7532 gnd.n239 240.244
R4637 gnd.n7525 gnd.n7524 240.244
R4638 gnd.n7522 gnd.n246 240.244
R4639 gnd.n7518 gnd.n7517 240.244
R4640 gnd.n7515 gnd.n253 240.244
R4641 gnd.n7511 gnd.n7510 240.244
R4642 gnd.n7508 gnd.n260 240.244
R4643 gnd.n7504 gnd.n7503 240.244
R4644 gnd.n7501 gnd.n267 240.244
R4645 gnd.n7497 gnd.n7496 240.244
R4646 gnd.n7494 gnd.n274 240.244
R4647 gnd.n7487 gnd.n283 240.244
R4648 gnd.n7485 gnd.n7484 240.244
R4649 gnd.n7482 gnd.n285 240.244
R4650 gnd.n7478 gnd.n7477 240.244
R4651 gnd.n7475 gnd.n292 240.244
R4652 gnd.n7471 gnd.n7470 240.244
R4653 gnd.n7468 gnd.n299 240.244
R4654 gnd.n7464 gnd.n7463 240.244
R4655 gnd.n7461 gnd.n306 240.244
R4656 gnd.n7457 gnd.n7456 240.244
R4657 gnd.n1497 gnd.n1338 240.244
R4658 gnd.n1497 gnd.n1350 240.244
R4659 gnd.n5908 gnd.n1350 240.244
R4660 gnd.n5908 gnd.n1362 240.244
R4661 gnd.n5918 gnd.n1362 240.244
R4662 gnd.n5918 gnd.n1373 240.244
R4663 gnd.n1487 gnd.n1373 240.244
R4664 gnd.n1487 gnd.n1382 240.244
R4665 gnd.n5927 gnd.n1382 240.244
R4666 gnd.n5927 gnd.n1393 240.244
R4667 gnd.n1481 gnd.n1393 240.244
R4668 gnd.n1481 gnd.n1402 240.244
R4669 gnd.n5999 gnd.n1402 240.244
R4670 gnd.n5999 gnd.n1413 240.244
R4671 gnd.n6003 gnd.n1413 240.244
R4672 gnd.n6003 gnd.n1422 240.244
R4673 gnd.n6013 gnd.n1422 240.244
R4674 gnd.n6013 gnd.n1433 240.244
R4675 gnd.n1465 gnd.n1433 240.244
R4676 gnd.n1465 gnd.n1442 240.244
R4677 gnd.n6020 gnd.n1442 240.244
R4678 gnd.n6020 gnd.n1451 240.244
R4679 gnd.n6050 gnd.n1451 240.244
R4680 gnd.n6050 gnd.n1457 240.244
R4681 gnd.n1457 gnd.n376 240.244
R4682 gnd.n376 gnd.n370 240.244
R4683 gnd.n7312 gnd.n370 240.244
R4684 gnd.n7312 gnd.n86 240.244
R4685 gnd.n363 gnd.n86 240.244
R4686 gnd.n7323 gnd.n363 240.244
R4687 gnd.n7323 gnd.n103 240.244
R4688 gnd.n7334 gnd.n103 240.244
R4689 gnd.n7334 gnd.n115 240.244
R4690 gnd.n7342 gnd.n115 240.244
R4691 gnd.n7342 gnd.n124 240.244
R4692 gnd.n7338 gnd.n124 240.244
R4693 gnd.n7338 gnd.n133 240.244
R4694 gnd.n7386 gnd.n133 240.244
R4695 gnd.n7386 gnd.n143 240.244
R4696 gnd.n7389 gnd.n143 240.244
R4697 gnd.n7389 gnd.n152 240.244
R4698 gnd.n7393 gnd.n152 240.244
R4699 gnd.n7393 gnd.n162 240.244
R4700 gnd.n7396 gnd.n162 240.244
R4701 gnd.n7396 gnd.n171 240.244
R4702 gnd.n7400 gnd.n171 240.244
R4703 gnd.n7400 gnd.n181 240.244
R4704 gnd.n7403 gnd.n181 240.244
R4705 gnd.n7403 gnd.n190 240.244
R4706 gnd.n7407 gnd.n190 240.244
R4707 gnd.n7407 gnd.n200 240.244
R4708 gnd.n7412 gnd.n200 240.244
R4709 gnd.n7412 gnd.n208 240.244
R4710 gnd.n5756 gnd.n5755 240.244
R4711 gnd.n5758 gnd.n5756 240.244
R4712 gnd.n5764 gnd.n5746 240.244
R4713 gnd.n5768 gnd.n5766 240.244
R4714 gnd.n5774 gnd.n5742 240.244
R4715 gnd.n5778 gnd.n5776 240.244
R4716 gnd.n5784 gnd.n5738 240.244
R4717 gnd.n5788 gnd.n5786 240.244
R4718 gnd.n5797 gnd.n5734 240.244
R4719 gnd.n5801 gnd.n5799 240.244
R4720 gnd.n5807 gnd.n5730 240.244
R4721 gnd.n5811 gnd.n5809 240.244
R4722 gnd.n5818 gnd.n5726 240.244
R4723 gnd.n5824 gnd.n5822 240.244
R4724 gnd.n5830 gnd.n1528 240.244
R4725 gnd.n5834 gnd.n5832 240.244
R4726 gnd.n5840 gnd.n1524 240.244
R4727 gnd.n5844 gnd.n5842 240.244
R4728 gnd.n5852 gnd.n1520 240.244
R4729 gnd.n5856 gnd.n5854 240.244
R4730 gnd.n5862 gnd.n1516 240.244
R4731 gnd.n5866 gnd.n5864 240.244
R4732 gnd.n5872 gnd.n1512 240.244
R4733 gnd.n5876 gnd.n5874 240.244
R4734 gnd.n5882 gnd.n1508 240.244
R4735 gnd.n5886 gnd.n5884 240.244
R4736 gnd.n5893 gnd.n1504 240.244
R4737 gnd.n5896 gnd.n5895 240.244
R4738 gnd.n6121 gnd.n1343 240.244
R4739 gnd.n6117 gnd.n1343 240.244
R4740 gnd.n6117 gnd.n1348 240.244
R4741 gnd.n6109 gnd.n1348 240.244
R4742 gnd.n6109 gnd.n1365 240.244
R4743 gnd.n6105 gnd.n1365 240.244
R4744 gnd.n6105 gnd.n1371 240.244
R4745 gnd.n6097 gnd.n1371 240.244
R4746 gnd.n6097 gnd.n1385 240.244
R4747 gnd.n6093 gnd.n1385 240.244
R4748 gnd.n6093 gnd.n1391 240.244
R4749 gnd.n6085 gnd.n1391 240.244
R4750 gnd.n6085 gnd.n1405 240.244
R4751 gnd.n6081 gnd.n1405 240.244
R4752 gnd.n6081 gnd.n1411 240.244
R4753 gnd.n6073 gnd.n1411 240.244
R4754 gnd.n6073 gnd.n1425 240.244
R4755 gnd.n6069 gnd.n1425 240.244
R4756 gnd.n6069 gnd.n1431 240.244
R4757 gnd.n6061 gnd.n1431 240.244
R4758 gnd.n6061 gnd.n1445 240.244
R4759 gnd.n6057 gnd.n1445 240.244
R4760 gnd.n6057 gnd.n1449 240.244
R4761 gnd.n1449 gnd.n378 240.244
R4762 gnd.n7303 gnd.n378 240.244
R4763 gnd.n7303 gnd.n7301 240.244
R4764 gnd.n7301 gnd.n89 240.244
R4765 gnd.n7637 gnd.n89 240.244
R4766 gnd.n7637 gnd.n90 240.244
R4767 gnd.n100 gnd.n90 240.244
R4768 gnd.n7631 gnd.n100 240.244
R4769 gnd.n7631 gnd.n101 240.244
R4770 gnd.n7623 gnd.n101 240.244
R4771 gnd.n7623 gnd.n117 240.244
R4772 gnd.n7619 gnd.n117 240.244
R4773 gnd.n7619 gnd.n122 240.244
R4774 gnd.n7611 gnd.n122 240.244
R4775 gnd.n7611 gnd.n136 240.244
R4776 gnd.n7607 gnd.n136 240.244
R4777 gnd.n7607 gnd.n142 240.244
R4778 gnd.n7599 gnd.n142 240.244
R4779 gnd.n7599 gnd.n154 240.244
R4780 gnd.n7595 gnd.n154 240.244
R4781 gnd.n7595 gnd.n160 240.244
R4782 gnd.n7587 gnd.n160 240.244
R4783 gnd.n7587 gnd.n174 240.244
R4784 gnd.n7583 gnd.n174 240.244
R4785 gnd.n7583 gnd.n180 240.244
R4786 gnd.n7575 gnd.n180 240.244
R4787 gnd.n7575 gnd.n193 240.244
R4788 gnd.n7571 gnd.n193 240.244
R4789 gnd.n7571 gnd.n199 240.244
R4790 gnd.n7563 gnd.n199 240.244
R4791 gnd.n6374 gnd.n1096 240.244
R4792 gnd.n6372 gnd.n6371 240.244
R4793 gnd.n6369 gnd.n1102 240.244
R4794 gnd.n6365 gnd.n6364 240.244
R4795 gnd.n6362 gnd.n1110 240.244
R4796 gnd.n6358 gnd.n6357 240.244
R4797 gnd.n6355 gnd.n1117 240.244
R4798 gnd.n6351 gnd.n6350 240.244
R4799 gnd.n6348 gnd.n1124 240.244
R4800 gnd.n6343 gnd.n6342 240.244
R4801 gnd.n6340 gnd.n1133 240.244
R4802 gnd.n6336 gnd.n6335 240.244
R4803 gnd.n6333 gnd.n1140 240.244
R4804 gnd.n4460 gnd.n4459 240.244
R4805 gnd.n4463 gnd.n4462 240.244
R4806 gnd.n4470 gnd.n4469 240.244
R4807 gnd.n4473 gnd.n4472 240.244
R4808 gnd.n4480 gnd.n4479 240.244
R4809 gnd.n4483 gnd.n4482 240.244
R4810 gnd.n4490 gnd.n4489 240.244
R4811 gnd.n4493 gnd.n4492 240.244
R4812 gnd.n4500 gnd.n4499 240.244
R4813 gnd.n4503 gnd.n4502 240.244
R4814 gnd.n4510 gnd.n4509 240.244
R4815 gnd.n4513 gnd.n4512 240.244
R4816 gnd.n4520 gnd.n4519 240.244
R4817 gnd.n4523 gnd.n4522 240.244
R4818 gnd.n4530 gnd.n4529 240.244
R4819 gnd.n4046 gnd.n2260 240.244
R4820 gnd.n2260 gnd.n2250 240.244
R4821 gnd.n4062 gnd.n2250 240.244
R4822 gnd.n4063 gnd.n4062 240.244
R4823 gnd.n4063 gnd.n2240 240.244
R4824 gnd.n4066 gnd.n2240 240.244
R4825 gnd.n4066 gnd.n2231 240.244
R4826 gnd.n2231 gnd.n2224 240.244
R4827 gnd.n4100 gnd.n2224 240.244
R4828 gnd.n4100 gnd.n2213 240.244
R4829 gnd.n4103 gnd.n2213 240.244
R4830 gnd.n4103 gnd.n2206 240.244
R4831 gnd.n4105 gnd.n2206 240.244
R4832 gnd.n4105 gnd.n2192 240.244
R4833 gnd.n4137 gnd.n2192 240.244
R4834 gnd.n4137 gnd.n2184 240.244
R4835 gnd.n2199 gnd.n2184 240.244
R4836 gnd.n2199 gnd.n942 240.244
R4837 gnd.n2173 gnd.n942 240.244
R4838 gnd.n2173 gnd.n954 240.244
R4839 gnd.n4183 gnd.n954 240.244
R4840 gnd.n4183 gnd.n966 240.244
R4841 gnd.n4179 gnd.n966 240.244
R4842 gnd.n4179 gnd.n4168 240.244
R4843 gnd.n4168 gnd.n2160 240.244
R4844 gnd.n2160 gnd.n2154 240.244
R4845 gnd.n2167 gnd.n2154 240.244
R4846 gnd.n2167 gnd.n2148 240.244
R4847 gnd.n2148 gnd.n2146 240.244
R4848 gnd.n2146 gnd.n2132 240.244
R4849 gnd.n2132 gnd.n982 240.244
R4850 gnd.n4249 gnd.n982 240.244
R4851 gnd.n4249 gnd.n994 240.244
R4852 gnd.n4255 gnd.n994 240.244
R4853 gnd.n4255 gnd.n1003 240.244
R4854 gnd.n4262 gnd.n1003 240.244
R4855 gnd.n4262 gnd.n1013 240.244
R4856 gnd.n2119 gnd.n1013 240.244
R4857 gnd.n2119 gnd.n1023 240.244
R4858 gnd.n4325 gnd.n1023 240.244
R4859 gnd.n4325 gnd.n1033 240.244
R4860 gnd.n4330 gnd.n1033 240.244
R4861 gnd.n4330 gnd.n1043 240.244
R4862 gnd.n4340 gnd.n1043 240.244
R4863 gnd.n4340 gnd.n1053 240.244
R4864 gnd.n2101 gnd.n1053 240.244
R4865 gnd.n2101 gnd.n1063 240.244
R4866 gnd.n4347 gnd.n1063 240.244
R4867 gnd.n4347 gnd.n1073 240.244
R4868 gnd.n4352 gnd.n1073 240.244
R4869 gnd.n4352 gnd.n1084 240.244
R4870 gnd.n4357 gnd.n1084 240.244
R4871 gnd.n4357 gnd.n1093 240.244
R4872 gnd.n3788 gnd.n3787 240.244
R4873 gnd.n4036 gnd.n3787 240.244
R4874 gnd.n4034 gnd.n4033 240.244
R4875 gnd.n4030 gnd.n4029 240.244
R4876 gnd.n4026 gnd.n4025 240.244
R4877 gnd.n4022 gnd.n4021 240.244
R4878 gnd.n4018 gnd.n4017 240.244
R4879 gnd.n4014 gnd.n4013 240.244
R4880 gnd.n4010 gnd.n4009 240.244
R4881 gnd.n4005 gnd.n4004 240.244
R4882 gnd.n4001 gnd.n4000 240.244
R4883 gnd.n3997 gnd.n3996 240.244
R4884 gnd.n3993 gnd.n3992 240.244
R4885 gnd.n3989 gnd.n3988 240.244
R4886 gnd.n3985 gnd.n3984 240.244
R4887 gnd.n3981 gnd.n3980 240.244
R4888 gnd.n3977 gnd.n3976 240.244
R4889 gnd.n3973 gnd.n3972 240.244
R4890 gnd.n3969 gnd.n3968 240.244
R4891 gnd.n3965 gnd.n3964 240.244
R4892 gnd.n3961 gnd.n3960 240.244
R4893 gnd.n3957 gnd.n3956 240.244
R4894 gnd.n3953 gnd.n3952 240.244
R4895 gnd.n3949 gnd.n3948 240.244
R4896 gnd.n3945 gnd.n3944 240.244
R4897 gnd.n3941 gnd.n3940 240.244
R4898 gnd.n3937 gnd.n3936 240.244
R4899 gnd.n3933 gnd.n3932 240.244
R4900 gnd.n3929 gnd.n2271 240.244
R4901 gnd.n4054 gnd.n2258 240.244
R4902 gnd.n4054 gnd.n2254 240.244
R4903 gnd.n4060 gnd.n2254 240.244
R4904 gnd.n4060 gnd.n2238 240.244
R4905 gnd.n4078 gnd.n2238 240.244
R4906 gnd.n4078 gnd.n2233 240.244
R4907 gnd.n4086 gnd.n2233 240.244
R4908 gnd.n4086 gnd.n2234 240.244
R4909 gnd.n2234 gnd.n2212 240.244
R4910 gnd.n4114 gnd.n2212 240.244
R4911 gnd.n4114 gnd.n2208 240.244
R4912 gnd.n4120 gnd.n2208 240.244
R4913 gnd.n4120 gnd.n2190 240.244
R4914 gnd.n4144 gnd.n2190 240.244
R4915 gnd.n4144 gnd.n2186 240.244
R4916 gnd.n4151 gnd.n2186 240.244
R4917 gnd.n4151 gnd.n946 240.244
R4918 gnd.n6465 gnd.n946 240.244
R4919 gnd.n6465 gnd.n947 240.244
R4920 gnd.n6461 gnd.n947 240.244
R4921 gnd.n6461 gnd.n953 240.244
R4922 gnd.n6453 gnd.n953 240.244
R4923 gnd.n6453 gnd.n969 240.244
R4924 gnd.n2157 gnd.n969 240.244
R4925 gnd.n4223 gnd.n2157 240.244
R4926 gnd.n4226 gnd.n4223 240.244
R4927 gnd.n4226 gnd.n2147 240.244
R4928 gnd.n4237 gnd.n2147 240.244
R4929 gnd.n4240 gnd.n4237 240.244
R4930 gnd.n4240 gnd.n980 240.244
R4931 gnd.n6448 gnd.n980 240.244
R4932 gnd.n6448 gnd.n981 240.244
R4933 gnd.n6440 gnd.n981 240.244
R4934 gnd.n6440 gnd.n996 240.244
R4935 gnd.n6436 gnd.n996 240.244
R4936 gnd.n6436 gnd.n1001 240.244
R4937 gnd.n6428 gnd.n1001 240.244
R4938 gnd.n6428 gnd.n1016 240.244
R4939 gnd.n6424 gnd.n1016 240.244
R4940 gnd.n6424 gnd.n1022 240.244
R4941 gnd.n6416 gnd.n1022 240.244
R4942 gnd.n6416 gnd.n1035 240.244
R4943 gnd.n6412 gnd.n1035 240.244
R4944 gnd.n6412 gnd.n1041 240.244
R4945 gnd.n6404 gnd.n1041 240.244
R4946 gnd.n6404 gnd.n1056 240.244
R4947 gnd.n6400 gnd.n1056 240.244
R4948 gnd.n6400 gnd.n1062 240.244
R4949 gnd.n6392 gnd.n1062 240.244
R4950 gnd.n6392 gnd.n1076 240.244
R4951 gnd.n6388 gnd.n1076 240.244
R4952 gnd.n6388 gnd.n1082 240.244
R4953 gnd.n6380 gnd.n1082 240.244
R4954 gnd.n3748 gnd.n2296 240.244
R4955 gnd.n3741 gnd.n3740 240.244
R4956 gnd.n3738 gnd.n3737 240.244
R4957 gnd.n3734 gnd.n3733 240.244
R4958 gnd.n3730 gnd.n3729 240.244
R4959 gnd.n3726 gnd.n3725 240.244
R4960 gnd.n3722 gnd.n3721 240.244
R4961 gnd.n3718 gnd.n3717 240.244
R4962 gnd.n2992 gnd.n2704 240.244
R4963 gnd.n3002 gnd.n2704 240.244
R4964 gnd.n3002 gnd.n2695 240.244
R4965 gnd.n2695 gnd.n2684 240.244
R4966 gnd.n3023 gnd.n2684 240.244
R4967 gnd.n3023 gnd.n2678 240.244
R4968 gnd.n3033 gnd.n2678 240.244
R4969 gnd.n3033 gnd.n2667 240.244
R4970 gnd.n2667 gnd.n2659 240.244
R4971 gnd.n3051 gnd.n2659 240.244
R4972 gnd.n3052 gnd.n3051 240.244
R4973 gnd.n3052 gnd.n2644 240.244
R4974 gnd.n3054 gnd.n2644 240.244
R4975 gnd.n3054 gnd.n2630 240.244
R4976 gnd.n3096 gnd.n2630 240.244
R4977 gnd.n3097 gnd.n3096 240.244
R4978 gnd.n3100 gnd.n3097 240.244
R4979 gnd.n3100 gnd.n2585 240.244
R4980 gnd.n2625 gnd.n2585 240.244
R4981 gnd.n2625 gnd.n2595 240.244
R4982 gnd.n3110 gnd.n2595 240.244
R4983 gnd.n3110 gnd.n2616 240.244
R4984 gnd.n3120 gnd.n2616 240.244
R4985 gnd.n3120 gnd.n2498 240.244
R4986 gnd.n3165 gnd.n2498 240.244
R4987 gnd.n3165 gnd.n2484 240.244
R4988 gnd.n3187 gnd.n2484 240.244
R4989 gnd.n3188 gnd.n3187 240.244
R4990 gnd.n3188 gnd.n2471 240.244
R4991 gnd.n2471 gnd.n2460 240.244
R4992 gnd.n3219 gnd.n2460 240.244
R4993 gnd.n3220 gnd.n3219 240.244
R4994 gnd.n3221 gnd.n3220 240.244
R4995 gnd.n3221 gnd.n2445 240.244
R4996 gnd.n2445 gnd.n2444 240.244
R4997 gnd.n2444 gnd.n2429 240.244
R4998 gnd.n3272 gnd.n2429 240.244
R4999 gnd.n3273 gnd.n3272 240.244
R5000 gnd.n3273 gnd.n2416 240.244
R5001 gnd.n2416 gnd.n2405 240.244
R5002 gnd.n3304 gnd.n2405 240.244
R5003 gnd.n3305 gnd.n3304 240.244
R5004 gnd.n3306 gnd.n3305 240.244
R5005 gnd.n3306 gnd.n2389 240.244
R5006 gnd.n2389 gnd.n2388 240.244
R5007 gnd.n2388 gnd.n2375 240.244
R5008 gnd.n3361 gnd.n2375 240.244
R5009 gnd.n3362 gnd.n3361 240.244
R5010 gnd.n3362 gnd.n2362 240.244
R5011 gnd.n2362 gnd.n2352 240.244
R5012 gnd.n3649 gnd.n2352 240.244
R5013 gnd.n3652 gnd.n3649 240.244
R5014 gnd.n3652 gnd.n3651 240.244
R5015 gnd.n2982 gnd.n2717 240.244
R5016 gnd.n2738 gnd.n2717 240.244
R5017 gnd.n2741 gnd.n2740 240.244
R5018 gnd.n2748 gnd.n2747 240.244
R5019 gnd.n2751 gnd.n2750 240.244
R5020 gnd.n2758 gnd.n2757 240.244
R5021 gnd.n2761 gnd.n2760 240.244
R5022 gnd.n2768 gnd.n2767 240.244
R5023 gnd.n2990 gnd.n2714 240.244
R5024 gnd.n2714 gnd.n2693 240.244
R5025 gnd.n3013 gnd.n2693 240.244
R5026 gnd.n3013 gnd.n2687 240.244
R5027 gnd.n3021 gnd.n2687 240.244
R5028 gnd.n3021 gnd.n2689 240.244
R5029 gnd.n2689 gnd.n2665 240.244
R5030 gnd.n3043 gnd.n2665 240.244
R5031 gnd.n3043 gnd.n2661 240.244
R5032 gnd.n3049 gnd.n2661 240.244
R5033 gnd.n3049 gnd.n2643 240.244
R5034 gnd.n3074 gnd.n2643 240.244
R5035 gnd.n3074 gnd.n2638 240.244
R5036 gnd.n3086 gnd.n2638 240.244
R5037 gnd.n3086 gnd.n2639 240.244
R5038 gnd.n3082 gnd.n2639 240.244
R5039 gnd.n3082 gnd.n2587 240.244
R5040 gnd.n3134 gnd.n2587 240.244
R5041 gnd.n3134 gnd.n2588 240.244
R5042 gnd.n3130 gnd.n2588 240.244
R5043 gnd.n3130 gnd.n2594 240.244
R5044 gnd.n2614 gnd.n2594 240.244
R5045 gnd.n2614 gnd.n2496 240.244
R5046 gnd.n3169 gnd.n2496 240.244
R5047 gnd.n3169 gnd.n2491 240.244
R5048 gnd.n3177 gnd.n2491 240.244
R5049 gnd.n3177 gnd.n2492 240.244
R5050 gnd.n2492 gnd.n2469 240.244
R5051 gnd.n3209 gnd.n2469 240.244
R5052 gnd.n3209 gnd.n2464 240.244
R5053 gnd.n3217 gnd.n2464 240.244
R5054 gnd.n3217 gnd.n2465 240.244
R5055 gnd.n2465 gnd.n2442 240.244
R5056 gnd.n3254 gnd.n2442 240.244
R5057 gnd.n3254 gnd.n2437 240.244
R5058 gnd.n3262 gnd.n2437 240.244
R5059 gnd.n3262 gnd.n2438 240.244
R5060 gnd.n2438 gnd.n2414 240.244
R5061 gnd.n3294 gnd.n2414 240.244
R5062 gnd.n3294 gnd.n2409 240.244
R5063 gnd.n3302 gnd.n2409 240.244
R5064 gnd.n3302 gnd.n2410 240.244
R5065 gnd.n2410 gnd.n2387 240.244
R5066 gnd.n3343 gnd.n2387 240.244
R5067 gnd.n3343 gnd.n2382 240.244
R5068 gnd.n3351 gnd.n2382 240.244
R5069 gnd.n3351 gnd.n2383 240.244
R5070 gnd.n2383 gnd.n2360 240.244
R5071 gnd.n3637 gnd.n2360 240.244
R5072 gnd.n3637 gnd.n2355 240.244
R5073 gnd.n3647 gnd.n2355 240.244
R5074 gnd.n3647 gnd.n2356 240.244
R5075 gnd.n2356 gnd.n2295 240.244
R5076 gnd.n317 gnd.n206 240.244
R5077 gnd.n7446 gnd.n7445 240.244
R5078 gnd.n7443 gnd.n321 240.244
R5079 gnd.n7439 gnd.n7438 240.244
R5080 gnd.n7436 gnd.n328 240.244
R5081 gnd.n7432 gnd.n7431 240.244
R5082 gnd.n7429 gnd.n335 240.244
R5083 gnd.n7425 gnd.n7424 240.244
R5084 gnd.n7422 gnd.n342 240.244
R5085 gnd.n5362 gnd.n1339 240.244
R5086 gnd.n5362 gnd.n1351 240.244
R5087 gnd.n5910 gnd.n1351 240.244
R5088 gnd.n5910 gnd.n1363 240.244
R5089 gnd.n5916 gnd.n1363 240.244
R5090 gnd.n5916 gnd.n1374 240.244
R5091 gnd.n5935 gnd.n1374 240.244
R5092 gnd.n5935 gnd.n1383 240.244
R5093 gnd.n5929 gnd.n1383 240.244
R5094 gnd.n5929 gnd.n1394 240.244
R5095 gnd.n5991 gnd.n1394 240.244
R5096 gnd.n5991 gnd.n1403 240.244
R5097 gnd.n5997 gnd.n1403 240.244
R5098 gnd.n5997 gnd.n1414 240.244
R5099 gnd.n6005 gnd.n1414 240.244
R5100 gnd.n6005 gnd.n1423 240.244
R5101 gnd.n6011 gnd.n1423 240.244
R5102 gnd.n6011 gnd.n1434 240.244
R5103 gnd.n6036 gnd.n1434 240.244
R5104 gnd.n6036 gnd.n1443 240.244
R5105 gnd.n6022 gnd.n1443 240.244
R5106 gnd.n6022 gnd.n1452 240.244
R5107 gnd.n1459 gnd.n1452 240.244
R5108 gnd.n6023 gnd.n1459 240.244
R5109 gnd.n6023 gnd.n377 240.244
R5110 gnd.n7299 gnd.n377 240.244
R5111 gnd.n7299 gnd.n82 240.244
R5112 gnd.n7639 gnd.n82 240.244
R5113 gnd.n7639 gnd.n84 240.244
R5114 gnd.n7325 gnd.n84 240.244
R5115 gnd.n7325 gnd.n104 240.244
R5116 gnd.n7332 gnd.n104 240.244
R5117 gnd.n7332 gnd.n116 240.244
R5118 gnd.n7344 gnd.n116 240.244
R5119 gnd.n7344 gnd.n125 240.244
R5120 gnd.n7347 gnd.n125 240.244
R5121 gnd.n7347 gnd.n134 240.244
R5122 gnd.n7384 gnd.n134 240.244
R5123 gnd.n7384 gnd.n144 240.244
R5124 gnd.n7380 gnd.n144 240.244
R5125 gnd.n7380 gnd.n153 240.244
R5126 gnd.n7377 gnd.n153 240.244
R5127 gnd.n7377 gnd.n163 240.244
R5128 gnd.n7374 gnd.n163 240.244
R5129 gnd.n7374 gnd.n172 240.244
R5130 gnd.n7371 gnd.n172 240.244
R5131 gnd.n7371 gnd.n182 240.244
R5132 gnd.n7368 gnd.n182 240.244
R5133 gnd.n7368 gnd.n191 240.244
R5134 gnd.n7365 gnd.n191 240.244
R5135 gnd.n7365 gnd.n201 240.244
R5136 gnd.n7414 gnd.n201 240.244
R5137 gnd.n7414 gnd.n209 240.244
R5138 gnd.n5461 gnd.n5410 240.244
R5139 gnd.n5465 gnd.n5463 240.244
R5140 gnd.n5480 gnd.n5401 240.244
R5141 gnd.n5484 gnd.n5482 240.244
R5142 gnd.n5499 gnd.n5392 240.244
R5143 gnd.n5503 gnd.n5501 240.244
R5144 gnd.n5519 gnd.n5383 240.244
R5145 gnd.n5523 gnd.n5521 240.244
R5146 gnd.n5379 gnd.n5378 240.244
R5147 gnd.n1353 gnd.n1341 240.244
R5148 gnd.n6115 gnd.n1353 240.244
R5149 gnd.n6115 gnd.n1354 240.244
R5150 gnd.n6111 gnd.n1354 240.244
R5151 gnd.n6111 gnd.n1360 240.244
R5152 gnd.n6103 gnd.n1360 240.244
R5153 gnd.n6103 gnd.n1375 240.244
R5154 gnd.n6099 gnd.n1375 240.244
R5155 gnd.n6099 gnd.n1380 240.244
R5156 gnd.n6091 gnd.n1380 240.244
R5157 gnd.n6091 gnd.n1396 240.244
R5158 gnd.n6087 gnd.n1396 240.244
R5159 gnd.n6087 gnd.n1401 240.244
R5160 gnd.n6079 gnd.n1401 240.244
R5161 gnd.n6079 gnd.n1415 240.244
R5162 gnd.n6075 gnd.n1415 240.244
R5163 gnd.n6075 gnd.n1420 240.244
R5164 gnd.n6067 gnd.n1420 240.244
R5165 gnd.n6067 gnd.n1436 240.244
R5166 gnd.n6063 gnd.n1436 240.244
R5167 gnd.n6063 gnd.n1441 240.244
R5168 gnd.n6055 gnd.n1441 240.244
R5169 gnd.n6055 gnd.n1453 240.244
R5170 gnd.n1453 gnd.n374 240.244
R5171 gnd.n7305 gnd.n374 240.244
R5172 gnd.n7305 gnd.n368 240.244
R5173 gnd.n7314 gnd.n368 240.244
R5174 gnd.n7314 gnd.n88 240.244
R5175 gnd.n7318 gnd.n88 240.244
R5176 gnd.n7318 gnd.n106 240.244
R5177 gnd.n7629 gnd.n106 240.244
R5178 gnd.n7629 gnd.n107 240.244
R5179 gnd.n7625 gnd.n107 240.244
R5180 gnd.n7625 gnd.n113 240.244
R5181 gnd.n7617 gnd.n113 240.244
R5182 gnd.n7617 gnd.n126 240.244
R5183 gnd.n7613 gnd.n126 240.244
R5184 gnd.n7613 gnd.n131 240.244
R5185 gnd.n7605 gnd.n131 240.244
R5186 gnd.n7605 gnd.n146 240.244
R5187 gnd.n7601 gnd.n146 240.244
R5188 gnd.n7601 gnd.n151 240.244
R5189 gnd.n7593 gnd.n151 240.244
R5190 gnd.n7593 gnd.n164 240.244
R5191 gnd.n7589 gnd.n164 240.244
R5192 gnd.n7589 gnd.n169 240.244
R5193 gnd.n7581 gnd.n169 240.244
R5194 gnd.n7581 gnd.n184 240.244
R5195 gnd.n7577 gnd.n184 240.244
R5196 gnd.n7577 gnd.n189 240.244
R5197 gnd.n7569 gnd.n189 240.244
R5198 gnd.n7569 gnd.n202 240.244
R5199 gnd.n7565 gnd.n202 240.244
R5200 gnd.n2315 gnd.n2273 240.244
R5201 gnd.n3708 gnd.n3707 240.244
R5202 gnd.n3704 gnd.n3703 240.244
R5203 gnd.n3700 gnd.n3699 240.244
R5204 gnd.n3696 gnd.n3695 240.244
R5205 gnd.n3692 gnd.n3691 240.244
R5206 gnd.n3688 gnd.n3687 240.244
R5207 gnd.n3684 gnd.n3683 240.244
R5208 gnd.n3680 gnd.n3679 240.244
R5209 gnd.n3676 gnd.n3675 240.244
R5210 gnd.n3672 gnd.n3671 240.244
R5211 gnd.n3668 gnd.n3667 240.244
R5212 gnd.n3664 gnd.n3663 240.244
R5213 gnd.n2905 gnd.n2802 240.244
R5214 gnd.n2905 gnd.n2795 240.244
R5215 gnd.n2916 gnd.n2795 240.244
R5216 gnd.n2916 gnd.n2791 240.244
R5217 gnd.n2922 gnd.n2791 240.244
R5218 gnd.n2922 gnd.n2783 240.244
R5219 gnd.n2932 gnd.n2783 240.244
R5220 gnd.n2932 gnd.n2778 240.244
R5221 gnd.n2968 gnd.n2778 240.244
R5222 gnd.n2968 gnd.n2779 240.244
R5223 gnd.n2779 gnd.n2726 240.244
R5224 gnd.n2963 gnd.n2726 240.244
R5225 gnd.n2963 gnd.n2962 240.244
R5226 gnd.n2962 gnd.n2705 240.244
R5227 gnd.n2958 gnd.n2705 240.244
R5228 gnd.n2958 gnd.n2696 240.244
R5229 gnd.n2955 gnd.n2696 240.244
R5230 gnd.n2955 gnd.n2954 240.244
R5231 gnd.n2954 gnd.n2679 240.244
R5232 gnd.n2950 gnd.n2679 240.244
R5233 gnd.n2950 gnd.n2668 240.244
R5234 gnd.n2668 gnd.n2649 240.244
R5235 gnd.n3063 gnd.n2649 240.244
R5236 gnd.n3063 gnd.n2645 240.244
R5237 gnd.n3071 gnd.n2645 240.244
R5238 gnd.n3071 gnd.n2636 240.244
R5239 gnd.n2636 gnd.n2572 240.244
R5240 gnd.n3143 gnd.n2572 240.244
R5241 gnd.n3143 gnd.n2573 240.244
R5242 gnd.n2584 gnd.n2573 240.244
R5243 gnd.n2619 gnd.n2584 240.244
R5244 gnd.n2622 gnd.n2619 240.244
R5245 gnd.n2622 gnd.n2596 240.244
R5246 gnd.n2609 gnd.n2596 240.244
R5247 gnd.n2609 gnd.n2606 240.244
R5248 gnd.n2606 gnd.n2499 240.244
R5249 gnd.n3164 gnd.n2499 240.244
R5250 gnd.n3164 gnd.n2489 240.244
R5251 gnd.n3160 gnd.n2489 240.244
R5252 gnd.n3160 gnd.n2483 240.244
R5253 gnd.n3157 gnd.n2483 240.244
R5254 gnd.n3157 gnd.n2472 240.244
R5255 gnd.n3154 gnd.n2472 240.244
R5256 gnd.n3154 gnd.n2450 240.244
R5257 gnd.n3230 gnd.n2450 240.244
R5258 gnd.n3230 gnd.n2446 240.244
R5259 gnd.n3251 gnd.n2446 240.244
R5260 gnd.n3251 gnd.n2435 240.244
R5261 gnd.n3247 gnd.n2435 240.244
R5262 gnd.n3247 gnd.n2428 240.244
R5263 gnd.n3244 gnd.n2428 240.244
R5264 gnd.n3244 gnd.n2417 240.244
R5265 gnd.n3241 gnd.n2417 240.244
R5266 gnd.n3241 gnd.n2394 240.244
R5267 gnd.n3315 gnd.n2394 240.244
R5268 gnd.n3315 gnd.n2390 240.244
R5269 gnd.n3340 gnd.n2390 240.244
R5270 gnd.n3340 gnd.n2381 240.244
R5271 gnd.n3336 gnd.n2381 240.244
R5272 gnd.n3336 gnd.n2374 240.244
R5273 gnd.n3332 gnd.n2374 240.244
R5274 gnd.n3332 gnd.n2363 240.244
R5275 gnd.n3329 gnd.n2363 240.244
R5276 gnd.n3329 gnd.n2344 240.244
R5277 gnd.n3659 gnd.n2344 240.244
R5278 gnd.n2819 gnd.n2818 240.244
R5279 gnd.n2890 gnd.n2818 240.244
R5280 gnd.n2888 gnd.n2887 240.244
R5281 gnd.n2884 gnd.n2883 240.244
R5282 gnd.n2880 gnd.n2879 240.244
R5283 gnd.n2876 gnd.n2875 240.244
R5284 gnd.n2872 gnd.n2871 240.244
R5285 gnd.n2868 gnd.n2867 240.244
R5286 gnd.n2864 gnd.n2863 240.244
R5287 gnd.n2860 gnd.n2859 240.244
R5288 gnd.n2856 gnd.n2855 240.244
R5289 gnd.n2852 gnd.n2851 240.244
R5290 gnd.n2848 gnd.n2806 240.244
R5291 gnd.n2908 gnd.n2800 240.244
R5292 gnd.n2908 gnd.n2796 240.244
R5293 gnd.n2914 gnd.n2796 240.244
R5294 gnd.n2914 gnd.n2789 240.244
R5295 gnd.n2924 gnd.n2789 240.244
R5296 gnd.n2924 gnd.n2785 240.244
R5297 gnd.n2930 gnd.n2785 240.244
R5298 gnd.n2930 gnd.n2776 240.244
R5299 gnd.n2970 gnd.n2776 240.244
R5300 gnd.n2970 gnd.n2727 240.244
R5301 gnd.n2978 gnd.n2727 240.244
R5302 gnd.n2978 gnd.n2728 240.244
R5303 gnd.n2728 gnd.n2706 240.244
R5304 gnd.n2999 gnd.n2706 240.244
R5305 gnd.n2999 gnd.n2698 240.244
R5306 gnd.n3010 gnd.n2698 240.244
R5307 gnd.n3010 gnd.n2699 240.244
R5308 gnd.n2699 gnd.n2680 240.244
R5309 gnd.n3030 gnd.n2680 240.244
R5310 gnd.n3030 gnd.n2670 240.244
R5311 gnd.n3040 gnd.n2670 240.244
R5312 gnd.n3040 gnd.n2651 240.244
R5313 gnd.n3061 gnd.n2651 240.244
R5314 gnd.n3061 gnd.n2653 240.244
R5315 gnd.n2653 gnd.n2634 240.244
R5316 gnd.n3089 gnd.n2634 240.244
R5317 gnd.n3089 gnd.n2576 240.244
R5318 gnd.n3141 gnd.n2576 240.244
R5319 gnd.n3141 gnd.n2577 240.244
R5320 gnd.n3137 gnd.n2577 240.244
R5321 gnd.n3137 gnd.n2583 240.244
R5322 gnd.n2598 gnd.n2583 240.244
R5323 gnd.n3127 gnd.n2598 240.244
R5324 gnd.n3127 gnd.n2599 240.244
R5325 gnd.n3123 gnd.n2599 240.244
R5326 gnd.n3123 gnd.n2605 240.244
R5327 gnd.n2605 gnd.n2488 240.244
R5328 gnd.n3180 gnd.n2488 240.244
R5329 gnd.n3180 gnd.n2481 240.244
R5330 gnd.n3191 gnd.n2481 240.244
R5331 gnd.n3191 gnd.n2474 240.244
R5332 gnd.n3206 gnd.n2474 240.244
R5333 gnd.n3206 gnd.n2475 240.244
R5334 gnd.n2475 gnd.n2453 240.244
R5335 gnd.n3228 gnd.n2453 240.244
R5336 gnd.n3228 gnd.n2454 240.244
R5337 gnd.n2454 gnd.n2433 240.244
R5338 gnd.n3265 gnd.n2433 240.244
R5339 gnd.n3265 gnd.n2426 240.244
R5340 gnd.n3276 gnd.n2426 240.244
R5341 gnd.n3276 gnd.n2419 240.244
R5342 gnd.n3291 gnd.n2419 240.244
R5343 gnd.n3291 gnd.n2420 240.244
R5344 gnd.n2420 gnd.n2397 240.244
R5345 gnd.n3313 gnd.n2397 240.244
R5346 gnd.n3313 gnd.n2399 240.244
R5347 gnd.n2399 gnd.n2379 240.244
R5348 gnd.n3354 gnd.n2379 240.244
R5349 gnd.n3354 gnd.n2372 240.244
R5350 gnd.n3365 gnd.n2372 240.244
R5351 gnd.n3365 gnd.n2365 240.244
R5352 gnd.n3634 gnd.n2365 240.244
R5353 gnd.n3634 gnd.n2366 240.244
R5354 gnd.n2366 gnd.n2347 240.244
R5355 gnd.n3657 gnd.n2347 240.244
R5356 gnd.n4545 gnd.n1091 240.244
R5357 gnd.n4556 gnd.n4547 240.244
R5358 gnd.n4559 gnd.n4558 240.244
R5359 gnd.n4568 gnd.n4567 240.244
R5360 gnd.n4579 gnd.n4570 240.244
R5361 gnd.n4582 gnd.n4581 240.244
R5362 gnd.n4591 gnd.n4590 240.244
R5363 gnd.n4594 gnd.n4593 240.244
R5364 gnd.n4663 gnd.n4662 240.244
R5365 gnd.n3883 gnd.n2261 240.244
R5366 gnd.n3880 gnd.n2261 240.244
R5367 gnd.n3880 gnd.n2252 240.244
R5368 gnd.n3877 gnd.n2252 240.244
R5369 gnd.n3877 gnd.n2241 240.244
R5370 gnd.n2241 gnd.n2230 240.244
R5371 gnd.n4088 gnd.n2230 240.244
R5372 gnd.n4088 gnd.n2226 240.244
R5373 gnd.n4098 gnd.n2226 240.244
R5374 gnd.n4098 gnd.n2214 240.244
R5375 gnd.n2214 gnd.n2205 240.244
R5376 gnd.n4122 gnd.n2205 240.244
R5377 gnd.n4123 gnd.n4122 240.244
R5378 gnd.n4123 gnd.n2193 240.244
R5379 gnd.n4135 gnd.n2193 240.244
R5380 gnd.n4135 gnd.n2185 240.244
R5381 gnd.n4131 gnd.n2185 240.244
R5382 gnd.n4131 gnd.n943 240.244
R5383 gnd.n4189 gnd.n943 240.244
R5384 gnd.n4189 gnd.n955 240.244
R5385 gnd.n4185 gnd.n955 240.244
R5386 gnd.n4185 gnd.n967 240.244
R5387 gnd.n4169 gnd.n967 240.244
R5388 gnd.n4175 gnd.n4169 240.244
R5389 gnd.n4175 gnd.n2153 240.244
R5390 gnd.n4228 gnd.n2153 240.244
R5391 gnd.n4228 gnd.n2149 240.244
R5392 gnd.n4235 gnd.n2149 240.244
R5393 gnd.n4235 gnd.n2133 240.244
R5394 gnd.n4276 gnd.n2133 240.244
R5395 gnd.n4276 gnd.n983 240.244
R5396 gnd.n2138 gnd.n983 240.244
R5397 gnd.n2138 gnd.n995 240.244
R5398 gnd.n2139 gnd.n995 240.244
R5399 gnd.n2139 gnd.n1004 240.244
R5400 gnd.n4264 gnd.n1004 240.244
R5401 gnd.n4264 gnd.n1014 240.244
R5402 gnd.n4317 gnd.n1014 240.244
R5403 gnd.n4317 gnd.n1024 240.244
R5404 gnd.n4323 gnd.n1024 240.244
R5405 gnd.n4323 gnd.n1034 240.244
R5406 gnd.n4332 gnd.n1034 240.244
R5407 gnd.n4332 gnd.n1044 240.244
R5408 gnd.n4338 gnd.n1044 240.244
R5409 gnd.n4338 gnd.n1054 240.244
R5410 gnd.n4372 gnd.n1054 240.244
R5411 gnd.n4372 gnd.n1064 240.244
R5412 gnd.n2106 gnd.n1064 240.244
R5413 gnd.n2106 gnd.n1074 240.244
R5414 gnd.n2107 gnd.n1074 240.244
R5415 gnd.n2107 gnd.n1085 240.244
R5416 gnd.n4359 gnd.n1085 240.244
R5417 gnd.n4359 gnd.n1094 240.244
R5418 gnd.n3920 gnd.n3919 240.244
R5419 gnd.n3916 gnd.n3915 240.244
R5420 gnd.n3912 gnd.n3911 240.244
R5421 gnd.n3908 gnd.n3907 240.244
R5422 gnd.n3904 gnd.n3903 240.244
R5423 gnd.n3900 gnd.n3899 240.244
R5424 gnd.n3896 gnd.n3895 240.244
R5425 gnd.n3892 gnd.n3891 240.244
R5426 gnd.n3867 gnd.n3786 240.244
R5427 gnd.n4052 gnd.n2262 240.244
R5428 gnd.n4052 gnd.n2263 240.244
R5429 gnd.n2263 gnd.n2253 240.244
R5430 gnd.n2253 gnd.n2243 240.244
R5431 gnd.n4076 gnd.n2243 240.244
R5432 gnd.n4076 gnd.n2244 240.244
R5433 gnd.n2244 gnd.n2232 240.244
R5434 gnd.n4071 gnd.n2232 240.244
R5435 gnd.n4071 gnd.n2216 240.244
R5436 gnd.n4112 gnd.n2216 240.244
R5437 gnd.n4112 gnd.n2217 240.244
R5438 gnd.n2217 gnd.n2207 240.244
R5439 gnd.n2207 gnd.n2194 240.244
R5440 gnd.n4142 gnd.n2194 240.244
R5441 gnd.n4142 gnd.n2182 240.244
R5442 gnd.n4153 gnd.n2182 240.244
R5443 gnd.n4154 gnd.n4153 240.244
R5444 gnd.n4154 gnd.n945 240.244
R5445 gnd.n957 gnd.n945 240.244
R5446 gnd.n6459 gnd.n957 240.244
R5447 gnd.n6459 gnd.n958 240.244
R5448 gnd.n6455 gnd.n958 240.244
R5449 gnd.n6455 gnd.n964 240.244
R5450 gnd.n2162 gnd.n964 240.244
R5451 gnd.n4221 gnd.n2162 240.244
R5452 gnd.n4221 gnd.n2156 240.244
R5453 gnd.n4217 gnd.n2156 240.244
R5454 gnd.n4217 gnd.n2144 240.244
R5455 gnd.n4242 gnd.n2144 240.244
R5456 gnd.n4242 gnd.n985 240.244
R5457 gnd.n6446 gnd.n985 240.244
R5458 gnd.n6446 gnd.n986 240.244
R5459 gnd.n6442 gnd.n986 240.244
R5460 gnd.n6442 gnd.n992 240.244
R5461 gnd.n6434 gnd.n992 240.244
R5462 gnd.n6434 gnd.n1006 240.244
R5463 gnd.n6430 gnd.n1006 240.244
R5464 gnd.n6430 gnd.n1011 240.244
R5465 gnd.n6422 gnd.n1011 240.244
R5466 gnd.n6422 gnd.n1026 240.244
R5467 gnd.n6418 gnd.n1026 240.244
R5468 gnd.n6418 gnd.n1031 240.244
R5469 gnd.n6410 gnd.n1031 240.244
R5470 gnd.n6410 gnd.n1046 240.244
R5471 gnd.n6406 gnd.n1046 240.244
R5472 gnd.n6406 gnd.n1051 240.244
R5473 gnd.n6398 gnd.n1051 240.244
R5474 gnd.n6398 gnd.n1066 240.244
R5475 gnd.n6394 gnd.n1066 240.244
R5476 gnd.n6394 gnd.n1071 240.244
R5477 gnd.n6386 gnd.n1071 240.244
R5478 gnd.n6386 gnd.n1087 240.244
R5479 gnd.n6382 gnd.n1087 240.244
R5480 gnd.n6644 gnd.n768 240.244
R5481 gnd.n6648 gnd.n768 240.244
R5482 gnd.n6648 gnd.n764 240.244
R5483 gnd.n6654 gnd.n764 240.244
R5484 gnd.n6654 gnd.n762 240.244
R5485 gnd.n6658 gnd.n762 240.244
R5486 gnd.n6658 gnd.n758 240.244
R5487 gnd.n6664 gnd.n758 240.244
R5488 gnd.n6664 gnd.n756 240.244
R5489 gnd.n6668 gnd.n756 240.244
R5490 gnd.n6668 gnd.n752 240.244
R5491 gnd.n6674 gnd.n752 240.244
R5492 gnd.n6674 gnd.n750 240.244
R5493 gnd.n6678 gnd.n750 240.244
R5494 gnd.n6678 gnd.n746 240.244
R5495 gnd.n6684 gnd.n746 240.244
R5496 gnd.n6684 gnd.n744 240.244
R5497 gnd.n6688 gnd.n744 240.244
R5498 gnd.n6688 gnd.n740 240.244
R5499 gnd.n6694 gnd.n740 240.244
R5500 gnd.n6694 gnd.n738 240.244
R5501 gnd.n6698 gnd.n738 240.244
R5502 gnd.n6698 gnd.n734 240.244
R5503 gnd.n6704 gnd.n734 240.244
R5504 gnd.n6704 gnd.n732 240.244
R5505 gnd.n6708 gnd.n732 240.244
R5506 gnd.n6708 gnd.n728 240.244
R5507 gnd.n6714 gnd.n728 240.244
R5508 gnd.n6714 gnd.n726 240.244
R5509 gnd.n6718 gnd.n726 240.244
R5510 gnd.n6718 gnd.n722 240.244
R5511 gnd.n6724 gnd.n722 240.244
R5512 gnd.n6724 gnd.n720 240.244
R5513 gnd.n6728 gnd.n720 240.244
R5514 gnd.n6728 gnd.n716 240.244
R5515 gnd.n6734 gnd.n716 240.244
R5516 gnd.n6734 gnd.n714 240.244
R5517 gnd.n6738 gnd.n714 240.244
R5518 gnd.n6738 gnd.n710 240.244
R5519 gnd.n6744 gnd.n710 240.244
R5520 gnd.n6744 gnd.n708 240.244
R5521 gnd.n6748 gnd.n708 240.244
R5522 gnd.n6748 gnd.n704 240.244
R5523 gnd.n6754 gnd.n704 240.244
R5524 gnd.n6754 gnd.n702 240.244
R5525 gnd.n6758 gnd.n702 240.244
R5526 gnd.n6758 gnd.n698 240.244
R5527 gnd.n6764 gnd.n698 240.244
R5528 gnd.n6764 gnd.n696 240.244
R5529 gnd.n6768 gnd.n696 240.244
R5530 gnd.n6768 gnd.n692 240.244
R5531 gnd.n6774 gnd.n692 240.244
R5532 gnd.n6774 gnd.n690 240.244
R5533 gnd.n6778 gnd.n690 240.244
R5534 gnd.n6778 gnd.n686 240.244
R5535 gnd.n6784 gnd.n686 240.244
R5536 gnd.n6784 gnd.n684 240.244
R5537 gnd.n6788 gnd.n684 240.244
R5538 gnd.n6788 gnd.n680 240.244
R5539 gnd.n6794 gnd.n680 240.244
R5540 gnd.n6794 gnd.n678 240.244
R5541 gnd.n6798 gnd.n678 240.244
R5542 gnd.n6798 gnd.n674 240.244
R5543 gnd.n6804 gnd.n674 240.244
R5544 gnd.n6804 gnd.n672 240.244
R5545 gnd.n6808 gnd.n672 240.244
R5546 gnd.n6808 gnd.n668 240.244
R5547 gnd.n6814 gnd.n668 240.244
R5548 gnd.n6814 gnd.n666 240.244
R5549 gnd.n6818 gnd.n666 240.244
R5550 gnd.n6818 gnd.n662 240.244
R5551 gnd.n6824 gnd.n662 240.244
R5552 gnd.n6824 gnd.n660 240.244
R5553 gnd.n6828 gnd.n660 240.244
R5554 gnd.n6828 gnd.n656 240.244
R5555 gnd.n6834 gnd.n656 240.244
R5556 gnd.n6834 gnd.n654 240.244
R5557 gnd.n6838 gnd.n654 240.244
R5558 gnd.n6838 gnd.n650 240.244
R5559 gnd.n6844 gnd.n650 240.244
R5560 gnd.n6844 gnd.n648 240.244
R5561 gnd.n6848 gnd.n648 240.244
R5562 gnd.n6848 gnd.n644 240.244
R5563 gnd.n6854 gnd.n644 240.244
R5564 gnd.n6854 gnd.n642 240.244
R5565 gnd.n6858 gnd.n642 240.244
R5566 gnd.n6858 gnd.n638 240.244
R5567 gnd.n6864 gnd.n638 240.244
R5568 gnd.n6864 gnd.n636 240.244
R5569 gnd.n6868 gnd.n636 240.244
R5570 gnd.n6868 gnd.n632 240.244
R5571 gnd.n6874 gnd.n632 240.244
R5572 gnd.n6874 gnd.n630 240.244
R5573 gnd.n6878 gnd.n630 240.244
R5574 gnd.n6878 gnd.n626 240.244
R5575 gnd.n6884 gnd.n626 240.244
R5576 gnd.n6884 gnd.n624 240.244
R5577 gnd.n6888 gnd.n624 240.244
R5578 gnd.n6888 gnd.n620 240.244
R5579 gnd.n6894 gnd.n620 240.244
R5580 gnd.n6894 gnd.n618 240.244
R5581 gnd.n6898 gnd.n618 240.244
R5582 gnd.n6898 gnd.n614 240.244
R5583 gnd.n6904 gnd.n614 240.244
R5584 gnd.n6904 gnd.n612 240.244
R5585 gnd.n6908 gnd.n612 240.244
R5586 gnd.n6908 gnd.n608 240.244
R5587 gnd.n6914 gnd.n608 240.244
R5588 gnd.n6914 gnd.n606 240.244
R5589 gnd.n6918 gnd.n606 240.244
R5590 gnd.n6918 gnd.n602 240.244
R5591 gnd.n6924 gnd.n602 240.244
R5592 gnd.n6924 gnd.n600 240.244
R5593 gnd.n6928 gnd.n600 240.244
R5594 gnd.n6928 gnd.n596 240.244
R5595 gnd.n6934 gnd.n596 240.244
R5596 gnd.n6934 gnd.n594 240.244
R5597 gnd.n6938 gnd.n594 240.244
R5598 gnd.n6938 gnd.n590 240.244
R5599 gnd.n6944 gnd.n590 240.244
R5600 gnd.n6944 gnd.n588 240.244
R5601 gnd.n6948 gnd.n588 240.244
R5602 gnd.n6948 gnd.n584 240.244
R5603 gnd.n6954 gnd.n584 240.244
R5604 gnd.n6954 gnd.n582 240.244
R5605 gnd.n6958 gnd.n582 240.244
R5606 gnd.n6958 gnd.n578 240.244
R5607 gnd.n6964 gnd.n578 240.244
R5608 gnd.n6964 gnd.n576 240.244
R5609 gnd.n6968 gnd.n576 240.244
R5610 gnd.n6968 gnd.n572 240.244
R5611 gnd.n6974 gnd.n572 240.244
R5612 gnd.n6974 gnd.n570 240.244
R5613 gnd.n6978 gnd.n570 240.244
R5614 gnd.n6978 gnd.n566 240.244
R5615 gnd.n6984 gnd.n566 240.244
R5616 gnd.n6984 gnd.n564 240.244
R5617 gnd.n6988 gnd.n564 240.244
R5618 gnd.n6988 gnd.n560 240.244
R5619 gnd.n6994 gnd.n560 240.244
R5620 gnd.n6994 gnd.n558 240.244
R5621 gnd.n6998 gnd.n558 240.244
R5622 gnd.n6998 gnd.n554 240.244
R5623 gnd.n7004 gnd.n554 240.244
R5624 gnd.n7004 gnd.n552 240.244
R5625 gnd.n7008 gnd.n552 240.244
R5626 gnd.n7008 gnd.n548 240.244
R5627 gnd.n7014 gnd.n548 240.244
R5628 gnd.n7014 gnd.n546 240.244
R5629 gnd.n7018 gnd.n546 240.244
R5630 gnd.n7018 gnd.n542 240.244
R5631 gnd.n7024 gnd.n542 240.244
R5632 gnd.n7024 gnd.n540 240.244
R5633 gnd.n7028 gnd.n540 240.244
R5634 gnd.n7028 gnd.n536 240.244
R5635 gnd.n7034 gnd.n536 240.244
R5636 gnd.n7034 gnd.n534 240.244
R5637 gnd.n7038 gnd.n534 240.244
R5638 gnd.n7038 gnd.n530 240.244
R5639 gnd.n7044 gnd.n530 240.244
R5640 gnd.n7044 gnd.n528 240.244
R5641 gnd.n7048 gnd.n528 240.244
R5642 gnd.n7048 gnd.n524 240.244
R5643 gnd.n7055 gnd.n524 240.244
R5644 gnd.n7055 gnd.n522 240.244
R5645 gnd.n7059 gnd.n522 240.244
R5646 gnd.n7059 gnd.n519 240.244
R5647 gnd.n7065 gnd.n517 240.244
R5648 gnd.n7069 gnd.n517 240.244
R5649 gnd.n7069 gnd.n513 240.244
R5650 gnd.n7075 gnd.n513 240.244
R5651 gnd.n7075 gnd.n511 240.244
R5652 gnd.n7079 gnd.n511 240.244
R5653 gnd.n7079 gnd.n507 240.244
R5654 gnd.n7085 gnd.n507 240.244
R5655 gnd.n7085 gnd.n505 240.244
R5656 gnd.n7089 gnd.n505 240.244
R5657 gnd.n7089 gnd.n501 240.244
R5658 gnd.n7095 gnd.n501 240.244
R5659 gnd.n7095 gnd.n499 240.244
R5660 gnd.n7099 gnd.n499 240.244
R5661 gnd.n7099 gnd.n495 240.244
R5662 gnd.n7105 gnd.n495 240.244
R5663 gnd.n7105 gnd.n493 240.244
R5664 gnd.n7109 gnd.n493 240.244
R5665 gnd.n7109 gnd.n489 240.244
R5666 gnd.n7115 gnd.n489 240.244
R5667 gnd.n7115 gnd.n487 240.244
R5668 gnd.n7119 gnd.n487 240.244
R5669 gnd.n7119 gnd.n483 240.244
R5670 gnd.n7125 gnd.n483 240.244
R5671 gnd.n7125 gnd.n481 240.244
R5672 gnd.n7129 gnd.n481 240.244
R5673 gnd.n7129 gnd.n477 240.244
R5674 gnd.n7135 gnd.n477 240.244
R5675 gnd.n7135 gnd.n475 240.244
R5676 gnd.n7139 gnd.n475 240.244
R5677 gnd.n7139 gnd.n471 240.244
R5678 gnd.n7145 gnd.n471 240.244
R5679 gnd.n7145 gnd.n469 240.244
R5680 gnd.n7149 gnd.n469 240.244
R5681 gnd.n7149 gnd.n465 240.244
R5682 gnd.n7155 gnd.n465 240.244
R5683 gnd.n7155 gnd.n463 240.244
R5684 gnd.n7159 gnd.n463 240.244
R5685 gnd.n7159 gnd.n459 240.244
R5686 gnd.n7165 gnd.n459 240.244
R5687 gnd.n7165 gnd.n457 240.244
R5688 gnd.n7169 gnd.n457 240.244
R5689 gnd.n7169 gnd.n453 240.244
R5690 gnd.n7175 gnd.n453 240.244
R5691 gnd.n7175 gnd.n451 240.244
R5692 gnd.n7179 gnd.n451 240.244
R5693 gnd.n7179 gnd.n447 240.244
R5694 gnd.n7185 gnd.n447 240.244
R5695 gnd.n7185 gnd.n445 240.244
R5696 gnd.n7189 gnd.n445 240.244
R5697 gnd.n7189 gnd.n441 240.244
R5698 gnd.n7195 gnd.n441 240.244
R5699 gnd.n7195 gnd.n439 240.244
R5700 gnd.n7199 gnd.n439 240.244
R5701 gnd.n7199 gnd.n435 240.244
R5702 gnd.n7205 gnd.n435 240.244
R5703 gnd.n7205 gnd.n433 240.244
R5704 gnd.n7209 gnd.n433 240.244
R5705 gnd.n7209 gnd.n429 240.244
R5706 gnd.n7215 gnd.n429 240.244
R5707 gnd.n7215 gnd.n427 240.244
R5708 gnd.n7219 gnd.n427 240.244
R5709 gnd.n7219 gnd.n423 240.244
R5710 gnd.n7225 gnd.n423 240.244
R5711 gnd.n7225 gnd.n421 240.244
R5712 gnd.n7229 gnd.n421 240.244
R5713 gnd.n7229 gnd.n417 240.244
R5714 gnd.n7235 gnd.n417 240.244
R5715 gnd.n7235 gnd.n415 240.244
R5716 gnd.n7239 gnd.n415 240.244
R5717 gnd.n7239 gnd.n411 240.244
R5718 gnd.n7245 gnd.n411 240.244
R5719 gnd.n7245 gnd.n409 240.244
R5720 gnd.n7249 gnd.n409 240.244
R5721 gnd.n7249 gnd.n405 240.244
R5722 gnd.n7255 gnd.n405 240.244
R5723 gnd.n7255 gnd.n403 240.244
R5724 gnd.n7259 gnd.n403 240.244
R5725 gnd.n7259 gnd.n399 240.244
R5726 gnd.n7265 gnd.n399 240.244
R5727 gnd.n7265 gnd.n397 240.244
R5728 gnd.n7270 gnd.n397 240.244
R5729 gnd.n7270 gnd.n393 240.244
R5730 gnd.n7277 gnd.n393 240.244
R5731 gnd.n6468 gnd.n940 240.244
R5732 gnd.n4192 gnd.n940 240.244
R5733 gnd.n4198 gnd.n4192 240.244
R5734 gnd.n4199 gnd.n4198 240.244
R5735 gnd.n4200 gnd.n4199 240.244
R5736 gnd.n4200 gnd.n2171 240.244
R5737 gnd.n4205 gnd.n2171 240.244
R5738 gnd.n4206 gnd.n4205 240.244
R5739 gnd.n4206 gnd.n2168 240.244
R5740 gnd.n4214 gnd.n2168 240.244
R5741 gnd.n4214 gnd.n2169 240.244
R5742 gnd.n2169 gnd.n2128 240.244
R5743 gnd.n4279 gnd.n2128 240.244
R5744 gnd.n4280 gnd.n4279 240.244
R5745 gnd.n4281 gnd.n4280 240.244
R5746 gnd.n4281 gnd.n2125 240.244
R5747 gnd.n4287 gnd.n2125 240.244
R5748 gnd.n4288 gnd.n4287 240.244
R5749 gnd.n4289 gnd.n4288 240.244
R5750 gnd.n4289 gnd.n2120 240.244
R5751 gnd.n4314 gnd.n2120 240.244
R5752 gnd.n4314 gnd.n2121 240.244
R5753 gnd.n4310 gnd.n2121 240.244
R5754 gnd.n4310 gnd.n4309 240.244
R5755 gnd.n4309 gnd.n4308 240.244
R5756 gnd.n4308 gnd.n4297 240.244
R5757 gnd.n4304 gnd.n4297 240.244
R5758 gnd.n4304 gnd.n2100 240.244
R5759 gnd.n4375 gnd.n2100 240.244
R5760 gnd.n4376 gnd.n4375 240.244
R5761 gnd.n4376 gnd.n2096 240.244
R5762 gnd.n4382 gnd.n2096 240.244
R5763 gnd.n4383 gnd.n4382 240.244
R5764 gnd.n4384 gnd.n4383 240.244
R5765 gnd.n4384 gnd.n2092 240.244
R5766 gnd.n4390 gnd.n2092 240.244
R5767 gnd.n4392 gnd.n4390 240.244
R5768 gnd.n4394 gnd.n4392 240.244
R5769 gnd.n4394 gnd.n2088 240.244
R5770 gnd.n4400 gnd.n2088 240.244
R5771 gnd.n4400 gnd.n2067 240.244
R5772 gnd.n4678 gnd.n2067 240.244
R5773 gnd.n4678 gnd.n2062 240.244
R5774 gnd.n4686 gnd.n2062 240.244
R5775 gnd.n4686 gnd.n2063 240.244
R5776 gnd.n2063 gnd.n2042 240.244
R5777 gnd.n4710 gnd.n2042 240.244
R5778 gnd.n4710 gnd.n2037 240.244
R5779 gnd.n4719 gnd.n2037 240.244
R5780 gnd.n4719 gnd.n2038 240.244
R5781 gnd.n2038 gnd.n1213 240.244
R5782 gnd.n6254 gnd.n1213 240.244
R5783 gnd.n6254 gnd.n1214 240.244
R5784 gnd.n6250 gnd.n1214 240.244
R5785 gnd.n6250 gnd.n1220 240.244
R5786 gnd.n4755 gnd.n1220 240.244
R5787 gnd.n4755 gnd.n1916 240.244
R5788 gnd.n4792 gnd.n1916 240.244
R5789 gnd.n4792 gnd.n1912 240.244
R5790 gnd.n4798 gnd.n1912 240.244
R5791 gnd.n4798 gnd.n1898 240.244
R5792 gnd.n4834 gnd.n1898 240.244
R5793 gnd.n4834 gnd.n1893 240.244
R5794 gnd.n4842 gnd.n1893 240.244
R5795 gnd.n4842 gnd.n1894 240.244
R5796 gnd.n1894 gnd.n1872 240.244
R5797 gnd.n4896 gnd.n1872 240.244
R5798 gnd.n4896 gnd.n1868 240.244
R5799 gnd.n4902 gnd.n1868 240.244
R5800 gnd.n4902 gnd.n1854 240.244
R5801 gnd.n4924 gnd.n1854 240.244
R5802 gnd.n4924 gnd.n1849 240.244
R5803 gnd.n4932 gnd.n1849 240.244
R5804 gnd.n4932 gnd.n1850 240.244
R5805 gnd.n1850 gnd.n1821 240.244
R5806 gnd.n4974 gnd.n1821 240.244
R5807 gnd.n4974 gnd.n1817 240.244
R5808 gnd.n4980 gnd.n1817 240.244
R5809 gnd.n4980 gnd.n1798 240.244
R5810 gnd.n5014 gnd.n1798 240.244
R5811 gnd.n5014 gnd.n1794 240.244
R5812 gnd.n5020 gnd.n1794 240.244
R5813 gnd.n5020 gnd.n1776 240.244
R5814 gnd.n5071 gnd.n1776 240.244
R5815 gnd.n5071 gnd.n1772 240.244
R5816 gnd.n5077 gnd.n1772 240.244
R5817 gnd.n5077 gnd.n1756 240.244
R5818 gnd.n5096 gnd.n1756 240.244
R5819 gnd.n5096 gnd.n1752 240.244
R5820 gnd.n5102 gnd.n1752 240.244
R5821 gnd.n5102 gnd.n1736 240.244
R5822 gnd.n5156 gnd.n1736 240.244
R5823 gnd.n5156 gnd.n1732 240.244
R5824 gnd.n5162 gnd.n1732 240.244
R5825 gnd.n5162 gnd.n1714 240.244
R5826 gnd.n5185 gnd.n1714 240.244
R5827 gnd.n5185 gnd.n1709 240.244
R5828 gnd.n5193 gnd.n1709 240.244
R5829 gnd.n5193 gnd.n1710 240.244
R5830 gnd.n1710 gnd.n1686 240.244
R5831 gnd.n5236 gnd.n1686 240.244
R5832 gnd.n5236 gnd.n1682 240.244
R5833 gnd.n5242 gnd.n1682 240.244
R5834 gnd.n5242 gnd.n1666 240.244
R5835 gnd.n5262 gnd.n1666 240.244
R5836 gnd.n5262 gnd.n1661 240.244
R5837 gnd.n5270 gnd.n1661 240.244
R5838 gnd.n5270 gnd.n1662 240.244
R5839 gnd.n1662 gnd.n1636 240.244
R5840 gnd.n5306 gnd.n1636 240.244
R5841 gnd.n5306 gnd.n1630 240.244
R5842 gnd.n5315 gnd.n1630 240.244
R5843 gnd.n5315 gnd.n1632 240.244
R5844 gnd.n1632 gnd.n1582 240.244
R5845 gnd.n5561 gnd.n1582 240.244
R5846 gnd.n5561 gnd.n1583 240.244
R5847 gnd.n5557 gnd.n1583 240.244
R5848 gnd.n5557 gnd.n5556 240.244
R5849 gnd.n5556 gnd.n1589 240.244
R5850 gnd.n5549 gnd.n1589 240.244
R5851 gnd.n5549 gnd.n1594 240.244
R5852 gnd.n5545 gnd.n1594 240.244
R5853 gnd.n5545 gnd.n1604 240.244
R5854 gnd.n1604 gnd.n1320 240.244
R5855 gnd.n6136 gnd.n1320 240.244
R5856 gnd.n6136 gnd.n1321 240.244
R5857 gnd.n6132 gnd.n1321 240.244
R5858 gnd.n6132 gnd.n1327 240.244
R5859 gnd.n6128 gnd.n1327 240.244
R5860 gnd.n6128 gnd.n1330 240.244
R5861 gnd.n6124 gnd.n1330 240.244
R5862 gnd.n6124 gnd.n1336 240.244
R5863 gnd.n5945 gnd.n1336 240.244
R5864 gnd.n5945 gnd.n5942 240.244
R5865 gnd.n5951 gnd.n5942 240.244
R5866 gnd.n5952 gnd.n5951 240.244
R5867 gnd.n5953 gnd.n5952 240.244
R5868 gnd.n5953 gnd.n5938 240.244
R5869 gnd.n5959 gnd.n5938 240.244
R5870 gnd.n5960 gnd.n5959 240.244
R5871 gnd.n5961 gnd.n5960 240.244
R5872 gnd.n5961 gnd.n1482 240.244
R5873 gnd.n5988 gnd.n1482 240.244
R5874 gnd.n5988 gnd.n1483 240.244
R5875 gnd.n5984 gnd.n1483 240.244
R5876 gnd.n5984 gnd.n5983 240.244
R5877 gnd.n5983 gnd.n5982 240.244
R5878 gnd.n5982 gnd.n5969 240.244
R5879 gnd.n5978 gnd.n5969 240.244
R5880 gnd.n5978 gnd.n1463 240.244
R5881 gnd.n6039 gnd.n1463 240.244
R5882 gnd.n6040 gnd.n6039 240.244
R5883 gnd.n6041 gnd.n6040 240.244
R5884 gnd.n6041 gnd.n1461 240.244
R5885 gnd.n6047 gnd.n1461 240.244
R5886 gnd.n6047 gnd.n381 240.244
R5887 gnd.n7297 gnd.n381 240.244
R5888 gnd.n7297 gnd.n382 240.244
R5889 gnd.n7292 gnd.n382 240.244
R5890 gnd.n7292 gnd.n7291 240.244
R5891 gnd.n7291 gnd.n385 240.244
R5892 gnd.n7286 gnd.n385 240.244
R5893 gnd.n7286 gnd.n7285 240.244
R5894 gnd.n7285 gnd.n7284 240.244
R5895 gnd.n7284 gnd.n387 240.244
R5896 gnd.n7280 gnd.n387 240.244
R5897 gnd.n7280 gnd.n7279 240.244
R5898 gnd.n6638 gnd.n770 240.244
R5899 gnd.n6638 gnd.n773 240.244
R5900 gnd.n6634 gnd.n773 240.244
R5901 gnd.n6634 gnd.n775 240.244
R5902 gnd.n6630 gnd.n775 240.244
R5903 gnd.n6630 gnd.n781 240.244
R5904 gnd.n6626 gnd.n781 240.244
R5905 gnd.n6626 gnd.n783 240.244
R5906 gnd.n6622 gnd.n783 240.244
R5907 gnd.n6622 gnd.n789 240.244
R5908 gnd.n6618 gnd.n789 240.244
R5909 gnd.n6618 gnd.n791 240.244
R5910 gnd.n6614 gnd.n791 240.244
R5911 gnd.n6614 gnd.n797 240.244
R5912 gnd.n6610 gnd.n797 240.244
R5913 gnd.n6610 gnd.n799 240.244
R5914 gnd.n6606 gnd.n799 240.244
R5915 gnd.n6606 gnd.n805 240.244
R5916 gnd.n6602 gnd.n805 240.244
R5917 gnd.n6602 gnd.n807 240.244
R5918 gnd.n6598 gnd.n807 240.244
R5919 gnd.n6598 gnd.n813 240.244
R5920 gnd.n6594 gnd.n813 240.244
R5921 gnd.n6594 gnd.n815 240.244
R5922 gnd.n6590 gnd.n815 240.244
R5923 gnd.n6590 gnd.n821 240.244
R5924 gnd.n6586 gnd.n821 240.244
R5925 gnd.n6586 gnd.n823 240.244
R5926 gnd.n6582 gnd.n823 240.244
R5927 gnd.n6582 gnd.n829 240.244
R5928 gnd.n6578 gnd.n829 240.244
R5929 gnd.n6578 gnd.n831 240.244
R5930 gnd.n6574 gnd.n831 240.244
R5931 gnd.n6574 gnd.n837 240.244
R5932 gnd.n6570 gnd.n837 240.244
R5933 gnd.n6570 gnd.n839 240.244
R5934 gnd.n6566 gnd.n839 240.244
R5935 gnd.n6566 gnd.n845 240.244
R5936 gnd.n6562 gnd.n845 240.244
R5937 gnd.n6562 gnd.n847 240.244
R5938 gnd.n6558 gnd.n847 240.244
R5939 gnd.n6558 gnd.n853 240.244
R5940 gnd.n6554 gnd.n853 240.244
R5941 gnd.n6554 gnd.n855 240.244
R5942 gnd.n6550 gnd.n855 240.244
R5943 gnd.n6550 gnd.n861 240.244
R5944 gnd.n6546 gnd.n861 240.244
R5945 gnd.n6546 gnd.n863 240.244
R5946 gnd.n6542 gnd.n863 240.244
R5947 gnd.n6542 gnd.n869 240.244
R5948 gnd.n6538 gnd.n869 240.244
R5949 gnd.n6538 gnd.n871 240.244
R5950 gnd.n6534 gnd.n871 240.244
R5951 gnd.n6534 gnd.n877 240.244
R5952 gnd.n6530 gnd.n877 240.244
R5953 gnd.n6530 gnd.n879 240.244
R5954 gnd.n6526 gnd.n879 240.244
R5955 gnd.n6526 gnd.n885 240.244
R5956 gnd.n6522 gnd.n885 240.244
R5957 gnd.n6522 gnd.n887 240.244
R5958 gnd.n6518 gnd.n887 240.244
R5959 gnd.n6518 gnd.n893 240.244
R5960 gnd.n6514 gnd.n893 240.244
R5961 gnd.n6514 gnd.n895 240.244
R5962 gnd.n6510 gnd.n895 240.244
R5963 gnd.n6510 gnd.n901 240.244
R5964 gnd.n6506 gnd.n901 240.244
R5965 gnd.n6506 gnd.n903 240.244
R5966 gnd.n6502 gnd.n903 240.244
R5967 gnd.n6502 gnd.n909 240.244
R5968 gnd.n6498 gnd.n909 240.244
R5969 gnd.n6498 gnd.n911 240.244
R5970 gnd.n6494 gnd.n911 240.244
R5971 gnd.n6494 gnd.n917 240.244
R5972 gnd.n6490 gnd.n917 240.244
R5973 gnd.n6490 gnd.n919 240.244
R5974 gnd.n6486 gnd.n919 240.244
R5975 gnd.n6486 gnd.n925 240.244
R5976 gnd.n6482 gnd.n925 240.244
R5977 gnd.n6482 gnd.n927 240.244
R5978 gnd.n6478 gnd.n927 240.244
R5979 gnd.n6478 gnd.n933 240.244
R5980 gnd.n6474 gnd.n933 240.244
R5981 gnd.n6474 gnd.n935 240.244
R5982 gnd.n4689 gnd.n2058 240.244
R5983 gnd.n4689 gnd.n2052 240.244
R5984 gnd.n4696 gnd.n2052 240.244
R5985 gnd.n4696 gnd.n2053 240.244
R5986 gnd.n2053 gnd.n2034 240.244
R5987 gnd.n4722 gnd.n2034 240.244
R5988 gnd.n4722 gnd.n2028 240.244
R5989 gnd.n4732 gnd.n2028 240.244
R5990 gnd.n4732 gnd.n2029 240.244
R5991 gnd.n4726 gnd.n2029 240.244
R5992 gnd.n4726 gnd.n1224 240.244
R5993 gnd.n6247 gnd.n1224 240.244
R5994 gnd.n6247 gnd.n1225 240.244
R5995 gnd.n1230 gnd.n1225 240.244
R5996 gnd.n1231 gnd.n1230 240.244
R5997 gnd.n1232 gnd.n1231 240.244
R5998 gnd.n1910 gnd.n1232 240.244
R5999 gnd.n1910 gnd.n1235 240.244
R6000 gnd.n1236 gnd.n1235 240.244
R6001 gnd.n1237 gnd.n1236 240.244
R6002 gnd.n4844 gnd.n1237 240.244
R6003 gnd.n4844 gnd.n1240 240.244
R6004 gnd.n1241 gnd.n1240 240.244
R6005 gnd.n1242 gnd.n1241 240.244
R6006 gnd.n4893 gnd.n1242 240.244
R6007 gnd.n4893 gnd.n1245 240.244
R6008 gnd.n1246 gnd.n1245 240.244
R6009 gnd.n1247 gnd.n1246 240.244
R6010 gnd.n4921 gnd.n1247 240.244
R6011 gnd.n4921 gnd.n1250 240.244
R6012 gnd.n1251 gnd.n1250 240.244
R6013 gnd.n1252 gnd.n1251 240.244
R6014 gnd.n4946 gnd.n1252 240.244
R6015 gnd.n4946 gnd.n1255 240.244
R6016 gnd.n1256 gnd.n1255 240.244
R6017 gnd.n1257 gnd.n1256 240.244
R6018 gnd.n5001 gnd.n1257 240.244
R6019 gnd.n5001 gnd.n1260 240.244
R6020 gnd.n1261 gnd.n1260 240.244
R6021 gnd.n1262 gnd.n1261 240.244
R6022 gnd.n5060 gnd.n1262 240.244
R6023 gnd.n5060 gnd.n1265 240.244
R6024 gnd.n1266 gnd.n1265 240.244
R6025 gnd.n1267 gnd.n1266 240.244
R6026 gnd.n1763 gnd.n1267 240.244
R6027 gnd.n1763 gnd.n1270 240.244
R6028 gnd.n1271 gnd.n1270 240.244
R6029 gnd.n1272 gnd.n1271 240.244
R6030 gnd.n5042 gnd.n1272 240.244
R6031 gnd.n5042 gnd.n1275 240.244
R6032 gnd.n1276 gnd.n1275 240.244
R6033 gnd.n1277 gnd.n1276 240.244
R6034 gnd.n5173 gnd.n1277 240.244
R6035 gnd.n5173 gnd.n1280 240.244
R6036 gnd.n1281 gnd.n1280 240.244
R6037 gnd.n1282 gnd.n1281 240.244
R6038 gnd.n5133 gnd.n1282 240.244
R6039 gnd.n5133 gnd.n1285 240.244
R6040 gnd.n1286 gnd.n1285 240.244
R6041 gnd.n1287 gnd.n1286 240.244
R6042 gnd.n1680 gnd.n1287 240.244
R6043 gnd.n1680 gnd.n1290 240.244
R6044 gnd.n1291 gnd.n1290 240.244
R6045 gnd.n1292 gnd.n1291 240.244
R6046 gnd.n1652 gnd.n1292 240.244
R6047 gnd.n1652 gnd.n1295 240.244
R6048 gnd.n1296 gnd.n1295 240.244
R6049 gnd.n1297 gnd.n1296 240.244
R6050 gnd.n5318 gnd.n1297 240.244
R6051 gnd.n5318 gnd.n1300 240.244
R6052 gnd.n1301 gnd.n1300 240.244
R6053 gnd.n1302 gnd.n1301 240.244
R6054 gnd.n5343 gnd.n1302 240.244
R6055 gnd.n5343 gnd.n1305 240.244
R6056 gnd.n1306 gnd.n1305 240.244
R6057 gnd.n1307 gnd.n1306 240.244
R6058 gnd.n5551 gnd.n1307 240.244
R6059 gnd.n5551 gnd.n1310 240.244
R6060 gnd.n1311 gnd.n1310 240.244
R6061 gnd.n1312 gnd.n1311 240.244
R6062 gnd.n1315 gnd.n1312 240.244
R6063 gnd.n6139 gnd.n1315 240.244
R6064 gnd.n4415 gnd.n4414 240.244
R6065 gnd.n4419 gnd.n4414 240.244
R6066 gnd.n4421 gnd.n4420 240.244
R6067 gnd.n4538 gnd.n4537 240.244
R6068 gnd.n4540 gnd.n4539 240.244
R6069 gnd.n4551 gnd.n4550 240.244
R6070 gnd.n4553 gnd.n4552 240.244
R6071 gnd.n4563 gnd.n4562 240.244
R6072 gnd.n4574 gnd.n4573 240.244
R6073 gnd.n4576 gnd.n4575 240.244
R6074 gnd.n4586 gnd.n4585 240.244
R6075 gnd.n4597 gnd.n4596 240.244
R6076 gnd.n4657 gnd.n2085 240.244
R6077 gnd.n2086 gnd.n2073 240.244
R6078 gnd.n4675 gnd.n2060 240.244
R6079 gnd.n2060 gnd.n2049 240.244
R6080 gnd.n4698 gnd.n2049 240.244
R6081 gnd.n4698 gnd.n2044 240.244
R6082 gnd.n4707 gnd.n2044 240.244
R6083 gnd.n4707 gnd.n2036 240.244
R6084 gnd.n2036 gnd.n1948 240.244
R6085 gnd.n4734 gnd.n1948 240.244
R6086 gnd.n4735 gnd.n4734 240.244
R6087 gnd.n4735 gnd.n1943 240.244
R6088 gnd.n4742 gnd.n1943 240.244
R6089 gnd.n4742 gnd.n1222 240.244
R6090 gnd.n4759 gnd.n1222 240.244
R6091 gnd.n4760 gnd.n4759 240.244
R6092 gnd.n4760 gnd.n1931 240.244
R6093 gnd.n4773 gnd.n1931 240.244
R6094 gnd.n4773 gnd.n1932 240.244
R6095 gnd.n4765 gnd.n1932 240.244
R6096 gnd.n4766 gnd.n4765 240.244
R6097 gnd.n4766 gnd.n1890 240.244
R6098 gnd.n4846 gnd.n1890 240.244
R6099 gnd.n4846 gnd.n1885 240.244
R6100 gnd.n4871 gnd.n1885 240.244
R6101 gnd.n4871 gnd.n1881 240.244
R6102 gnd.n1881 gnd.n1873 240.244
R6103 gnd.n4851 gnd.n1873 240.244
R6104 gnd.n4854 gnd.n4851 240.244
R6105 gnd.n4855 gnd.n4854 240.244
R6106 gnd.n4855 gnd.n1856 240.244
R6107 gnd.n1856 gnd.n1838 240.244
R6108 gnd.n4944 gnd.n1838 240.244
R6109 gnd.n4945 gnd.n4944 240.244
R6110 gnd.n4948 gnd.n4945 240.244
R6111 gnd.n4948 gnd.n1834 240.244
R6112 gnd.n4954 gnd.n1834 240.244
R6113 gnd.n4954 gnd.n1808 240.244
R6114 gnd.n5000 gnd.n1808 240.244
R6115 gnd.n5000 gnd.n1809 240.244
R6116 gnd.n4994 gnd.n1809 240.244
R6117 gnd.n4994 gnd.n1786 240.244
R6118 gnd.n5059 gnd.n1786 240.244
R6119 gnd.n5059 gnd.n1778 240.244
R6120 gnd.n5035 gnd.n1778 240.244
R6121 gnd.n5036 gnd.n5035 240.244
R6122 gnd.n5037 gnd.n5036 240.244
R6123 gnd.n5037 gnd.n1758 240.244
R6124 gnd.n1758 gnd.n1751 240.244
R6125 gnd.n5040 gnd.n1751 240.244
R6126 gnd.n5044 gnd.n5040 240.244
R6127 gnd.n5044 gnd.n1729 240.244
R6128 gnd.n5165 gnd.n1729 240.244
R6129 gnd.n5165 gnd.n1723 240.244
R6130 gnd.n5172 gnd.n1723 240.244
R6131 gnd.n5172 gnd.n1724 240.244
R6132 gnd.n1724 gnd.n1700 240.244
R6133 gnd.n5204 gnd.n1700 240.244
R6134 gnd.n5204 gnd.n1695 240.244
R6135 gnd.n5225 gnd.n1695 240.244
R6136 gnd.n5225 gnd.n1688 240.244
R6137 gnd.n5209 gnd.n1688 240.244
R6138 gnd.n5210 gnd.n5209 240.244
R6139 gnd.n5212 gnd.n5210 240.244
R6140 gnd.n5212 gnd.n1668 240.244
R6141 gnd.n1668 gnd.n1660 240.244
R6142 gnd.n1660 gnd.n1644 240.244
R6143 gnd.n5295 gnd.n1644 240.244
R6144 gnd.n5295 gnd.n1639 240.244
R6145 gnd.n5302 gnd.n1639 240.244
R6146 gnd.n5302 gnd.n1629 240.244
R6147 gnd.n1629 gnd.n1617 240.244
R6148 gnd.n5337 gnd.n1617 240.244
R6149 gnd.n5337 gnd.n1580 240.244
R6150 gnd.n5345 gnd.n1580 240.244
R6151 gnd.n5347 gnd.n5345 240.244
R6152 gnd.n5348 gnd.n5347 240.244
R6153 gnd.n5348 gnd.n1591 240.244
R6154 gnd.n1592 gnd.n1591 240.244
R6155 gnd.n5355 gnd.n1592 240.244
R6156 gnd.n5356 gnd.n5355 240.244
R6157 gnd.n5356 gnd.n1607 240.244
R6158 gnd.n5540 gnd.n1607 240.244
R6159 gnd.n5540 gnd.n1318 240.244
R6160 gnd.n5427 gnd.n5426 240.244
R6161 gnd.n5430 gnd.n5429 240.244
R6162 gnd.n5438 gnd.n5437 240.244
R6163 gnd.n5441 gnd.n5440 240.244
R6164 gnd.n5453 gnd.n5452 240.244
R6165 gnd.n5456 gnd.n5455 240.244
R6166 gnd.n5472 gnd.n5471 240.244
R6167 gnd.n5475 gnd.n5474 240.244
R6168 gnd.n5491 gnd.n5490 240.244
R6169 gnd.n5494 gnd.n5493 240.244
R6170 gnd.n5510 gnd.n5509 240.244
R6171 gnd.n5512 gnd.n5369 240.244
R6172 gnd.n5529 gnd.n5369 240.244
R6173 gnd.n5532 gnd.n5531 240.244
R6174 gnd.n1194 gnd.n1193 240.132
R6175 gnd.n5579 gnd.n5578 240.132
R6176 gnd.n6646 gnd.n6645 225.874
R6177 gnd.n6647 gnd.n6646 225.874
R6178 gnd.n6647 gnd.n763 225.874
R6179 gnd.n6655 gnd.n763 225.874
R6180 gnd.n6656 gnd.n6655 225.874
R6181 gnd.n6657 gnd.n6656 225.874
R6182 gnd.n6657 gnd.n757 225.874
R6183 gnd.n6665 gnd.n757 225.874
R6184 gnd.n6666 gnd.n6665 225.874
R6185 gnd.n6667 gnd.n6666 225.874
R6186 gnd.n6667 gnd.n751 225.874
R6187 gnd.n6675 gnd.n751 225.874
R6188 gnd.n6676 gnd.n6675 225.874
R6189 gnd.n6677 gnd.n6676 225.874
R6190 gnd.n6677 gnd.n745 225.874
R6191 gnd.n6685 gnd.n745 225.874
R6192 gnd.n6686 gnd.n6685 225.874
R6193 gnd.n6687 gnd.n6686 225.874
R6194 gnd.n6687 gnd.n739 225.874
R6195 gnd.n6695 gnd.n739 225.874
R6196 gnd.n6696 gnd.n6695 225.874
R6197 gnd.n6697 gnd.n6696 225.874
R6198 gnd.n6697 gnd.n733 225.874
R6199 gnd.n6705 gnd.n733 225.874
R6200 gnd.n6706 gnd.n6705 225.874
R6201 gnd.n6707 gnd.n6706 225.874
R6202 gnd.n6707 gnd.n727 225.874
R6203 gnd.n6715 gnd.n727 225.874
R6204 gnd.n6716 gnd.n6715 225.874
R6205 gnd.n6717 gnd.n6716 225.874
R6206 gnd.n6717 gnd.n721 225.874
R6207 gnd.n6725 gnd.n721 225.874
R6208 gnd.n6726 gnd.n6725 225.874
R6209 gnd.n6727 gnd.n6726 225.874
R6210 gnd.n6727 gnd.n715 225.874
R6211 gnd.n6735 gnd.n715 225.874
R6212 gnd.n6736 gnd.n6735 225.874
R6213 gnd.n6737 gnd.n6736 225.874
R6214 gnd.n6737 gnd.n709 225.874
R6215 gnd.n6745 gnd.n709 225.874
R6216 gnd.n6746 gnd.n6745 225.874
R6217 gnd.n6747 gnd.n6746 225.874
R6218 gnd.n6747 gnd.n703 225.874
R6219 gnd.n6755 gnd.n703 225.874
R6220 gnd.n6756 gnd.n6755 225.874
R6221 gnd.n6757 gnd.n6756 225.874
R6222 gnd.n6757 gnd.n697 225.874
R6223 gnd.n6765 gnd.n697 225.874
R6224 gnd.n6766 gnd.n6765 225.874
R6225 gnd.n6767 gnd.n6766 225.874
R6226 gnd.n6767 gnd.n691 225.874
R6227 gnd.n6775 gnd.n691 225.874
R6228 gnd.n6776 gnd.n6775 225.874
R6229 gnd.n6777 gnd.n6776 225.874
R6230 gnd.n6777 gnd.n685 225.874
R6231 gnd.n6785 gnd.n685 225.874
R6232 gnd.n6786 gnd.n6785 225.874
R6233 gnd.n6787 gnd.n6786 225.874
R6234 gnd.n6787 gnd.n679 225.874
R6235 gnd.n6795 gnd.n679 225.874
R6236 gnd.n6796 gnd.n6795 225.874
R6237 gnd.n6797 gnd.n6796 225.874
R6238 gnd.n6797 gnd.n673 225.874
R6239 gnd.n6805 gnd.n673 225.874
R6240 gnd.n6806 gnd.n6805 225.874
R6241 gnd.n6807 gnd.n6806 225.874
R6242 gnd.n6807 gnd.n667 225.874
R6243 gnd.n6815 gnd.n667 225.874
R6244 gnd.n6816 gnd.n6815 225.874
R6245 gnd.n6817 gnd.n6816 225.874
R6246 gnd.n6817 gnd.n661 225.874
R6247 gnd.n6825 gnd.n661 225.874
R6248 gnd.n6826 gnd.n6825 225.874
R6249 gnd.n6827 gnd.n6826 225.874
R6250 gnd.n6827 gnd.n655 225.874
R6251 gnd.n6835 gnd.n655 225.874
R6252 gnd.n6836 gnd.n6835 225.874
R6253 gnd.n6837 gnd.n6836 225.874
R6254 gnd.n6837 gnd.n649 225.874
R6255 gnd.n6845 gnd.n649 225.874
R6256 gnd.n6846 gnd.n6845 225.874
R6257 gnd.n6847 gnd.n6846 225.874
R6258 gnd.n6847 gnd.n643 225.874
R6259 gnd.n6855 gnd.n643 225.874
R6260 gnd.n6856 gnd.n6855 225.874
R6261 gnd.n6857 gnd.n6856 225.874
R6262 gnd.n6857 gnd.n637 225.874
R6263 gnd.n6865 gnd.n637 225.874
R6264 gnd.n6866 gnd.n6865 225.874
R6265 gnd.n6867 gnd.n6866 225.874
R6266 gnd.n6867 gnd.n631 225.874
R6267 gnd.n6875 gnd.n631 225.874
R6268 gnd.n6876 gnd.n6875 225.874
R6269 gnd.n6877 gnd.n6876 225.874
R6270 gnd.n6877 gnd.n625 225.874
R6271 gnd.n6885 gnd.n625 225.874
R6272 gnd.n6886 gnd.n6885 225.874
R6273 gnd.n6887 gnd.n6886 225.874
R6274 gnd.n6887 gnd.n619 225.874
R6275 gnd.n6895 gnd.n619 225.874
R6276 gnd.n6896 gnd.n6895 225.874
R6277 gnd.n6897 gnd.n6896 225.874
R6278 gnd.n6897 gnd.n613 225.874
R6279 gnd.n6905 gnd.n613 225.874
R6280 gnd.n6906 gnd.n6905 225.874
R6281 gnd.n6907 gnd.n6906 225.874
R6282 gnd.n6907 gnd.n607 225.874
R6283 gnd.n6915 gnd.n607 225.874
R6284 gnd.n6916 gnd.n6915 225.874
R6285 gnd.n6917 gnd.n6916 225.874
R6286 gnd.n6917 gnd.n601 225.874
R6287 gnd.n6925 gnd.n601 225.874
R6288 gnd.n6926 gnd.n6925 225.874
R6289 gnd.n6927 gnd.n6926 225.874
R6290 gnd.n6927 gnd.n595 225.874
R6291 gnd.n6935 gnd.n595 225.874
R6292 gnd.n6936 gnd.n6935 225.874
R6293 gnd.n6937 gnd.n6936 225.874
R6294 gnd.n6937 gnd.n589 225.874
R6295 gnd.n6945 gnd.n589 225.874
R6296 gnd.n6946 gnd.n6945 225.874
R6297 gnd.n6947 gnd.n6946 225.874
R6298 gnd.n6947 gnd.n583 225.874
R6299 gnd.n6955 gnd.n583 225.874
R6300 gnd.n6956 gnd.n6955 225.874
R6301 gnd.n6957 gnd.n6956 225.874
R6302 gnd.n6957 gnd.n577 225.874
R6303 gnd.n6965 gnd.n577 225.874
R6304 gnd.n6966 gnd.n6965 225.874
R6305 gnd.n6967 gnd.n6966 225.874
R6306 gnd.n6967 gnd.n571 225.874
R6307 gnd.n6975 gnd.n571 225.874
R6308 gnd.n6976 gnd.n6975 225.874
R6309 gnd.n6977 gnd.n6976 225.874
R6310 gnd.n6977 gnd.n565 225.874
R6311 gnd.n6985 gnd.n565 225.874
R6312 gnd.n6986 gnd.n6985 225.874
R6313 gnd.n6987 gnd.n6986 225.874
R6314 gnd.n6987 gnd.n559 225.874
R6315 gnd.n6995 gnd.n559 225.874
R6316 gnd.n6996 gnd.n6995 225.874
R6317 gnd.n6997 gnd.n6996 225.874
R6318 gnd.n6997 gnd.n553 225.874
R6319 gnd.n7005 gnd.n553 225.874
R6320 gnd.n7006 gnd.n7005 225.874
R6321 gnd.n7007 gnd.n7006 225.874
R6322 gnd.n7007 gnd.n547 225.874
R6323 gnd.n7015 gnd.n547 225.874
R6324 gnd.n7016 gnd.n7015 225.874
R6325 gnd.n7017 gnd.n7016 225.874
R6326 gnd.n7017 gnd.n541 225.874
R6327 gnd.n7025 gnd.n541 225.874
R6328 gnd.n7026 gnd.n7025 225.874
R6329 gnd.n7027 gnd.n7026 225.874
R6330 gnd.n7027 gnd.n535 225.874
R6331 gnd.n7035 gnd.n535 225.874
R6332 gnd.n7036 gnd.n7035 225.874
R6333 gnd.n7037 gnd.n7036 225.874
R6334 gnd.n7037 gnd.n529 225.874
R6335 gnd.n7045 gnd.n529 225.874
R6336 gnd.n7046 gnd.n7045 225.874
R6337 gnd.n7047 gnd.n7046 225.874
R6338 gnd.n7047 gnd.n523 225.874
R6339 gnd.n7056 gnd.n523 225.874
R6340 gnd.n7057 gnd.n7056 225.874
R6341 gnd.n7058 gnd.n7057 225.874
R6342 gnd.n7058 gnd.n518 225.874
R6343 gnd.n2843 gnd.t139 224.174
R6344 gnd.n2337 gnd.t134 224.174
R6345 gnd.n5820 gnd.n5819 199.319
R6346 gnd.n5821 gnd.n5820 199.319
R6347 gnd.n1146 gnd.n1145 199.319
R6348 gnd.n4458 gnd.n1146 199.319
R6349 gnd.n1195 gnd.n1192 186.49
R6350 gnd.n5580 gnd.n5577 186.49
R6351 gnd.n3618 gnd.n3617 185
R6352 gnd.n3616 gnd.n3615 185
R6353 gnd.n3595 gnd.n3594 185
R6354 gnd.n3610 gnd.n3609 185
R6355 gnd.n3608 gnd.n3607 185
R6356 gnd.n3599 gnd.n3598 185
R6357 gnd.n3602 gnd.n3601 185
R6358 gnd.n3586 gnd.n3585 185
R6359 gnd.n3584 gnd.n3583 185
R6360 gnd.n3563 gnd.n3562 185
R6361 gnd.n3578 gnd.n3577 185
R6362 gnd.n3576 gnd.n3575 185
R6363 gnd.n3567 gnd.n3566 185
R6364 gnd.n3570 gnd.n3569 185
R6365 gnd.n3554 gnd.n3553 185
R6366 gnd.n3552 gnd.n3551 185
R6367 gnd.n3531 gnd.n3530 185
R6368 gnd.n3546 gnd.n3545 185
R6369 gnd.n3544 gnd.n3543 185
R6370 gnd.n3535 gnd.n3534 185
R6371 gnd.n3538 gnd.n3537 185
R6372 gnd.n3523 gnd.n3522 185
R6373 gnd.n3521 gnd.n3520 185
R6374 gnd.n3500 gnd.n3499 185
R6375 gnd.n3515 gnd.n3514 185
R6376 gnd.n3513 gnd.n3512 185
R6377 gnd.n3504 gnd.n3503 185
R6378 gnd.n3507 gnd.n3506 185
R6379 gnd.n3491 gnd.n3490 185
R6380 gnd.n3489 gnd.n3488 185
R6381 gnd.n3468 gnd.n3467 185
R6382 gnd.n3483 gnd.n3482 185
R6383 gnd.n3481 gnd.n3480 185
R6384 gnd.n3472 gnd.n3471 185
R6385 gnd.n3475 gnd.n3474 185
R6386 gnd.n3459 gnd.n3458 185
R6387 gnd.n3457 gnd.n3456 185
R6388 gnd.n3436 gnd.n3435 185
R6389 gnd.n3451 gnd.n3450 185
R6390 gnd.n3449 gnd.n3448 185
R6391 gnd.n3440 gnd.n3439 185
R6392 gnd.n3443 gnd.n3442 185
R6393 gnd.n3427 gnd.n3426 185
R6394 gnd.n3425 gnd.n3424 185
R6395 gnd.n3404 gnd.n3403 185
R6396 gnd.n3419 gnd.n3418 185
R6397 gnd.n3417 gnd.n3416 185
R6398 gnd.n3408 gnd.n3407 185
R6399 gnd.n3411 gnd.n3410 185
R6400 gnd.n3396 gnd.n3395 185
R6401 gnd.n3394 gnd.n3393 185
R6402 gnd.n3373 gnd.n3372 185
R6403 gnd.n3388 gnd.n3387 185
R6404 gnd.n3386 gnd.n3385 185
R6405 gnd.n3377 gnd.n3376 185
R6406 gnd.n3380 gnd.n3379 185
R6407 gnd.n2844 gnd.t138 178.987
R6408 gnd.n2338 gnd.t135 178.987
R6409 gnd.n1 gnd.t281 170.774
R6410 gnd.n7 gnd.t287 170.103
R6411 gnd.n6 gnd.t361 170.103
R6412 gnd.n5 gnd.t285 170.103
R6413 gnd.n4 gnd.t291 170.103
R6414 gnd.n3 gnd.t95 170.103
R6415 gnd.n2 gnd.t293 170.103
R6416 gnd.n1 gnd.t9 170.103
R6417 gnd.n5648 gnd.n5647 163.367
R6418 gnd.n5644 gnd.n5643 163.367
R6419 gnd.n5640 gnd.n5639 163.367
R6420 gnd.n5636 gnd.n5635 163.367
R6421 gnd.n5632 gnd.n5631 163.367
R6422 gnd.n5628 gnd.n5627 163.367
R6423 gnd.n5624 gnd.n5623 163.367
R6424 gnd.n5620 gnd.n5619 163.367
R6425 gnd.n5616 gnd.n5615 163.367
R6426 gnd.n5612 gnd.n5611 163.367
R6427 gnd.n5608 gnd.n5607 163.367
R6428 gnd.n5604 gnd.n5603 163.367
R6429 gnd.n5600 gnd.n5599 163.367
R6430 gnd.n5596 gnd.n5595 163.367
R6431 gnd.n5591 gnd.n5590 163.367
R6432 gnd.n5723 gnd.n1535 163.367
R6433 gnd.n5720 gnd.n5719 163.367
R6434 gnd.n5717 gnd.n1568 163.367
R6435 gnd.n5712 gnd.n5711 163.367
R6436 gnd.n5708 gnd.n5707 163.367
R6437 gnd.n5704 gnd.n5703 163.367
R6438 gnd.n5700 gnd.n5699 163.367
R6439 gnd.n5696 gnd.n5695 163.367
R6440 gnd.n5692 gnd.n5691 163.367
R6441 gnd.n5688 gnd.n5687 163.367
R6442 gnd.n5684 gnd.n5683 163.367
R6443 gnd.n5680 gnd.n5679 163.367
R6444 gnd.n5676 gnd.n5675 163.367
R6445 gnd.n5672 gnd.n5671 163.367
R6446 gnd.n5668 gnd.n5667 163.367
R6447 gnd.n5664 gnd.n5663 163.367
R6448 gnd.n5660 gnd.n5659 163.367
R6449 gnd.n2025 gnd.n1211 163.367
R6450 gnd.n2021 gnd.n1211 163.367
R6451 gnd.n2021 gnd.n1942 163.367
R6452 gnd.n2017 gnd.n1942 163.367
R6453 gnd.n2017 gnd.n2016 163.367
R6454 gnd.n2016 gnd.n1938 163.367
R6455 gnd.n1938 gnd.n1921 163.367
R6456 gnd.n4785 gnd.n1921 163.367
R6457 gnd.n4785 gnd.n1918 163.367
R6458 gnd.n4790 gnd.n1918 163.367
R6459 gnd.n4790 gnd.n1919 163.367
R6460 gnd.n1919 gnd.n1909 163.367
R6461 gnd.n4801 gnd.n1909 163.367
R6462 gnd.n4801 gnd.n1907 163.367
R6463 gnd.n4814 gnd.n1907 163.367
R6464 gnd.n4814 gnd.n1900 163.367
R6465 gnd.n4810 gnd.n1900 163.367
R6466 gnd.n4810 gnd.n4807 163.367
R6467 gnd.n4807 gnd.n4806 163.367
R6468 gnd.n4806 gnd.n1883 163.367
R6469 gnd.n4874 gnd.n1883 163.367
R6470 gnd.n4874 gnd.n1880 163.367
R6471 gnd.n4883 gnd.n1880 163.367
R6472 gnd.n4883 gnd.n1874 163.367
R6473 gnd.n4879 gnd.n1874 163.367
R6474 gnd.n4879 gnd.n1867 163.367
R6475 gnd.n1867 gnd.n1859 163.367
R6476 gnd.n4912 gnd.n1859 163.367
R6477 gnd.n4912 gnd.n1857 163.367
R6478 gnd.n4919 gnd.n1857 163.367
R6479 gnd.n4919 gnd.n1847 163.367
R6480 gnd.n1848 gnd.n1847 163.367
R6481 gnd.n1848 gnd.n1840 163.367
R6482 gnd.n1840 gnd.n1830 163.367
R6483 gnd.n4962 gnd.n1830 163.367
R6484 gnd.n4962 gnd.n1831 163.367
R6485 gnd.n1831 gnd.n1823 163.367
R6486 gnd.n4957 gnd.n1823 163.367
R6487 gnd.n4957 gnd.n1815 163.367
R6488 gnd.n4984 gnd.n1815 163.367
R6489 gnd.n4984 gnd.n1807 163.367
R6490 gnd.n4987 gnd.n1807 163.367
R6491 gnd.n4987 gnd.n1800 163.367
R6492 gnd.n4991 gnd.n1800 163.367
R6493 gnd.n4991 gnd.n1792 163.367
R6494 gnd.n5024 gnd.n1792 163.367
R6495 gnd.n5024 gnd.n1785 163.367
R6496 gnd.n5027 gnd.n1785 163.367
R6497 gnd.n5027 gnd.n1779 163.367
R6498 gnd.n5032 gnd.n1779 163.367
R6499 gnd.n5032 gnd.n1769 163.367
R6500 gnd.n1769 gnd.n1761 163.367
R6501 gnd.n5087 gnd.n1761 163.367
R6502 gnd.n5087 gnd.n1759 163.367
R6503 gnd.n5092 gnd.n1759 163.367
R6504 gnd.n5092 gnd.n1750 163.367
R6505 gnd.n1750 gnd.n1742 163.367
R6506 gnd.n5121 gnd.n1742 163.367
R6507 gnd.n5121 gnd.n1739 163.367
R6508 gnd.n5154 gnd.n1739 163.367
R6509 gnd.n5154 gnd.n1740 163.367
R6510 gnd.n5150 gnd.n1740 163.367
R6511 gnd.n5150 gnd.n5149 163.367
R6512 gnd.n5149 gnd.n1721 163.367
R6513 gnd.n1722 gnd.n1721 163.367
R6514 gnd.n1722 gnd.n1715 163.367
R6515 gnd.n5143 gnd.n1715 163.367
R6516 gnd.n5143 gnd.n1708 163.367
R6517 gnd.n5139 gnd.n1708 163.367
R6518 gnd.n5139 gnd.n1702 163.367
R6519 gnd.n5136 gnd.n1702 163.367
R6520 gnd.n5136 gnd.n1694 163.367
R6521 gnd.n5129 gnd.n1694 163.367
R6522 gnd.n5129 gnd.n1689 163.367
R6523 gnd.n5126 gnd.n1689 163.367
R6524 gnd.n5126 gnd.n1677 163.367
R6525 gnd.n1677 gnd.n1671 163.367
R6526 gnd.n5252 gnd.n1671 163.367
R6527 gnd.n5252 gnd.n1669 163.367
R6528 gnd.n5257 gnd.n1669 163.367
R6529 gnd.n5257 gnd.n1659 163.367
R6530 gnd.n1659 gnd.n1651 163.367
R6531 gnd.n5285 gnd.n1651 163.367
R6532 gnd.n5285 gnd.n1648 163.367
R6533 gnd.n5292 gnd.n1648 163.367
R6534 gnd.n5292 gnd.n1649 163.367
R6535 gnd.n1649 gnd.n1638 163.367
R6536 gnd.n1638 gnd.n1628 163.367
R6537 gnd.n1628 gnd.n1621 163.367
R6538 gnd.n5328 gnd.n1621 163.367
R6539 gnd.n5328 gnd.n1619 163.367
R6540 gnd.n5334 gnd.n1619 163.367
R6541 gnd.n5334 gnd.n1579 163.367
R6542 gnd.n1579 gnd.n1572 163.367
R6543 gnd.n5655 gnd.n1572 163.367
R6544 gnd.n1186 gnd.n1185 163.367
R6545 gnd.n6319 gnd.n1185 163.367
R6546 gnd.n6317 gnd.n6316 163.367
R6547 gnd.n6313 gnd.n6312 163.367
R6548 gnd.n6309 gnd.n6308 163.367
R6549 gnd.n6305 gnd.n6304 163.367
R6550 gnd.n6301 gnd.n6300 163.367
R6551 gnd.n6297 gnd.n6296 163.367
R6552 gnd.n6293 gnd.n6292 163.367
R6553 gnd.n6289 gnd.n6288 163.367
R6554 gnd.n6285 gnd.n6284 163.367
R6555 gnd.n6281 gnd.n6280 163.367
R6556 gnd.n6277 gnd.n6276 163.367
R6557 gnd.n6273 gnd.n6272 163.367
R6558 gnd.n6269 gnd.n6268 163.367
R6559 gnd.n6265 gnd.n6264 163.367
R6560 gnd.n6328 gnd.n1151 163.367
R6561 gnd.n1954 gnd.n1953 163.367
R6562 gnd.n1959 gnd.n1958 163.367
R6563 gnd.n1963 gnd.n1962 163.367
R6564 gnd.n1967 gnd.n1966 163.367
R6565 gnd.n1971 gnd.n1970 163.367
R6566 gnd.n1975 gnd.n1974 163.367
R6567 gnd.n1979 gnd.n1978 163.367
R6568 gnd.n1983 gnd.n1982 163.367
R6569 gnd.n1987 gnd.n1986 163.367
R6570 gnd.n1991 gnd.n1990 163.367
R6571 gnd.n1995 gnd.n1994 163.367
R6572 gnd.n1999 gnd.n1998 163.367
R6573 gnd.n2003 gnd.n2002 163.367
R6574 gnd.n2007 gnd.n2006 163.367
R6575 gnd.n2011 gnd.n2010 163.367
R6576 gnd.n6257 gnd.n1187 163.367
R6577 gnd.n6257 gnd.n1209 163.367
R6578 gnd.n4745 gnd.n1209 163.367
R6579 gnd.n4746 gnd.n4745 163.367
R6580 gnd.n4746 gnd.n1939 163.367
R6581 gnd.n4750 gnd.n1939 163.367
R6582 gnd.n4750 gnd.n1924 163.367
R6583 gnd.n4783 gnd.n1924 163.367
R6584 gnd.n4783 gnd.n1925 163.367
R6585 gnd.n1925 gnd.n1917 163.367
R6586 gnd.n4778 gnd.n1917 163.367
R6587 gnd.n4778 gnd.n1928 163.367
R6588 gnd.n1928 gnd.n1905 163.367
R6589 gnd.n4818 gnd.n1905 163.367
R6590 gnd.n4818 gnd.n1902 163.367
R6591 gnd.n4831 gnd.n1902 163.367
R6592 gnd.n4831 gnd.n1903 163.367
R6593 gnd.n4827 gnd.n1903 163.367
R6594 gnd.n4827 gnd.n4826 163.367
R6595 gnd.n4826 gnd.n4825 163.367
R6596 gnd.n4825 gnd.n1878 163.367
R6597 gnd.n4887 gnd.n1878 163.367
R6598 gnd.n4887 gnd.n1876 163.367
R6599 gnd.n4891 gnd.n1876 163.367
R6600 gnd.n4891 gnd.n1865 163.367
R6601 gnd.n4905 gnd.n1865 163.367
R6602 gnd.n4905 gnd.n1862 163.367
R6603 gnd.n4910 gnd.n1862 163.367
R6604 gnd.n4910 gnd.n1863 163.367
R6605 gnd.n1863 gnd.n1845 163.367
R6606 gnd.n4937 gnd.n1845 163.367
R6607 gnd.n4937 gnd.n1843 163.367
R6608 gnd.n4941 gnd.n1843 163.367
R6609 gnd.n4941 gnd.n1828 163.367
R6610 gnd.n4964 gnd.n1828 163.367
R6611 gnd.n4964 gnd.n1825 163.367
R6612 gnd.n4971 gnd.n1825 163.367
R6613 gnd.n4971 gnd.n1826 163.367
R6614 gnd.n4967 gnd.n1826 163.367
R6615 gnd.n4967 gnd.n1805 163.367
R6616 gnd.n5004 gnd.n1805 163.367
R6617 gnd.n5004 gnd.n1802 163.367
R6618 gnd.n5011 gnd.n1802 163.367
R6619 gnd.n5011 gnd.n1803 163.367
R6620 gnd.n5007 gnd.n1803 163.367
R6621 gnd.n5007 gnd.n1783 163.367
R6622 gnd.n5063 gnd.n1783 163.367
R6623 gnd.n5063 gnd.n1781 163.367
R6624 gnd.n5067 gnd.n1781 163.367
R6625 gnd.n5067 gnd.n1768 163.367
R6626 gnd.n5080 gnd.n1768 163.367
R6627 gnd.n5080 gnd.n1765 163.367
R6628 gnd.n5085 gnd.n1765 163.367
R6629 gnd.n5085 gnd.n1766 163.367
R6630 gnd.n1766 gnd.n1748 163.367
R6631 gnd.n5107 gnd.n1748 163.367
R6632 gnd.n5107 gnd.n1745 163.367
R6633 gnd.n5119 gnd.n1745 163.367
R6634 gnd.n5119 gnd.n1746 163.367
R6635 gnd.n1746 gnd.n1737 163.367
R6636 gnd.n5114 gnd.n1737 163.367
R6637 gnd.n5114 gnd.n5111 163.367
R6638 gnd.n5111 gnd.n1719 163.367
R6639 gnd.n5178 gnd.n1719 163.367
R6640 gnd.n5178 gnd.n1717 163.367
R6641 gnd.n5182 gnd.n1717 163.367
R6642 gnd.n5182 gnd.n1706 163.367
R6643 gnd.n5197 gnd.n1706 163.367
R6644 gnd.n5197 gnd.n1704 163.367
R6645 gnd.n5201 gnd.n1704 163.367
R6646 gnd.n5201 gnd.n1693 163.367
R6647 gnd.n5228 gnd.n1693 163.367
R6648 gnd.n5228 gnd.n1691 163.367
R6649 gnd.n5232 gnd.n1691 163.367
R6650 gnd.n5232 gnd.n1675 163.367
R6651 gnd.n5245 gnd.n1675 163.367
R6652 gnd.n5245 gnd.n1672 163.367
R6653 gnd.n5250 gnd.n1672 163.367
R6654 gnd.n5250 gnd.n1673 163.367
R6655 gnd.n1673 gnd.n1658 163.367
R6656 gnd.n5275 gnd.n1658 163.367
R6657 gnd.n5275 gnd.n1655 163.367
R6658 gnd.n5283 gnd.n1655 163.367
R6659 gnd.n5283 gnd.n1656 163.367
R6660 gnd.n1656 gnd.n1646 163.367
R6661 gnd.n5278 gnd.n1646 163.367
R6662 gnd.n5278 gnd.n1626 163.367
R6663 gnd.n5321 gnd.n1626 163.367
R6664 gnd.n5321 gnd.n1623 163.367
R6665 gnd.n5326 gnd.n1623 163.367
R6666 gnd.n5326 gnd.n1624 163.367
R6667 gnd.n1624 gnd.n1577 163.367
R6668 gnd.n5565 gnd.n1577 163.367
R6669 gnd.n5565 gnd.n1574 163.367
R6670 gnd.n5653 gnd.n1574 163.367
R6671 gnd.n5586 gnd.n5585 156.462
R6672 gnd.n3558 gnd.n3526 153.042
R6673 gnd.n3622 gnd.n3621 152.079
R6674 gnd.n3590 gnd.n3589 152.079
R6675 gnd.n3558 gnd.n3557 152.079
R6676 gnd.n1200 gnd.n1199 152
R6677 gnd.n1201 gnd.n1190 152
R6678 gnd.n1203 gnd.n1202 152
R6679 gnd.n1205 gnd.n1188 152
R6680 gnd.n1207 gnd.n1206 152
R6681 gnd.n5584 gnd.n5568 152
R6682 gnd.n5576 gnd.n5569 152
R6683 gnd.n5575 gnd.n5574 152
R6684 gnd.n5573 gnd.n5570 152
R6685 gnd.n5571 gnd.t148 150.546
R6686 gnd.t68 gnd.n3600 147.661
R6687 gnd.t289 gnd.n3568 147.661
R6688 gnd.t115 gnd.n3536 147.661
R6689 gnd.t93 gnd.n3505 147.661
R6690 gnd.t298 gnd.n3473 147.661
R6691 gnd.t78 gnd.n3441 147.661
R6692 gnd.t273 gnd.n3409 147.661
R6693 gnd.t31 gnd.n3378 147.661
R6694 gnd.n5722 gnd.n1534 143.351
R6695 gnd.n1167 gnd.n1150 143.351
R6696 gnd.n6327 gnd.n1150 143.351
R6697 gnd.n7067 gnd.n7066 137.715
R6698 gnd.n7068 gnd.n7067 137.715
R6699 gnd.n7068 gnd.n512 137.715
R6700 gnd.n7076 gnd.n512 137.715
R6701 gnd.n7077 gnd.n7076 137.715
R6702 gnd.n7078 gnd.n7077 137.715
R6703 gnd.n7078 gnd.n506 137.715
R6704 gnd.n7086 gnd.n506 137.715
R6705 gnd.n7087 gnd.n7086 137.715
R6706 gnd.n7088 gnd.n7087 137.715
R6707 gnd.n7088 gnd.n500 137.715
R6708 gnd.n7096 gnd.n500 137.715
R6709 gnd.n7097 gnd.n7096 137.715
R6710 gnd.n7098 gnd.n7097 137.715
R6711 gnd.n7098 gnd.n494 137.715
R6712 gnd.n7106 gnd.n494 137.715
R6713 gnd.n7107 gnd.n7106 137.715
R6714 gnd.n7108 gnd.n7107 137.715
R6715 gnd.n7108 gnd.n488 137.715
R6716 gnd.n7116 gnd.n488 137.715
R6717 gnd.n7117 gnd.n7116 137.715
R6718 gnd.n7118 gnd.n7117 137.715
R6719 gnd.n7118 gnd.n482 137.715
R6720 gnd.n7126 gnd.n482 137.715
R6721 gnd.n7127 gnd.n7126 137.715
R6722 gnd.n7128 gnd.n7127 137.715
R6723 gnd.n7128 gnd.n476 137.715
R6724 gnd.n7136 gnd.n476 137.715
R6725 gnd.n7137 gnd.n7136 137.715
R6726 gnd.n7138 gnd.n7137 137.715
R6727 gnd.n7138 gnd.n470 137.715
R6728 gnd.n7146 gnd.n470 137.715
R6729 gnd.n7147 gnd.n7146 137.715
R6730 gnd.n7148 gnd.n7147 137.715
R6731 gnd.n7148 gnd.n464 137.715
R6732 gnd.n7156 gnd.n464 137.715
R6733 gnd.n7157 gnd.n7156 137.715
R6734 gnd.n7158 gnd.n7157 137.715
R6735 gnd.n7158 gnd.n458 137.715
R6736 gnd.n7166 gnd.n458 137.715
R6737 gnd.n7167 gnd.n7166 137.715
R6738 gnd.n7168 gnd.n7167 137.715
R6739 gnd.n7168 gnd.n452 137.715
R6740 gnd.n7176 gnd.n452 137.715
R6741 gnd.n7177 gnd.n7176 137.715
R6742 gnd.n7178 gnd.n7177 137.715
R6743 gnd.n7178 gnd.n446 137.715
R6744 gnd.n7186 gnd.n446 137.715
R6745 gnd.n7187 gnd.n7186 137.715
R6746 gnd.n7188 gnd.n7187 137.715
R6747 gnd.n7188 gnd.n440 137.715
R6748 gnd.n7196 gnd.n440 137.715
R6749 gnd.n7197 gnd.n7196 137.715
R6750 gnd.n7198 gnd.n7197 137.715
R6751 gnd.n7198 gnd.n434 137.715
R6752 gnd.n7206 gnd.n434 137.715
R6753 gnd.n7207 gnd.n7206 137.715
R6754 gnd.n7208 gnd.n7207 137.715
R6755 gnd.n7208 gnd.n428 137.715
R6756 gnd.n7216 gnd.n428 137.715
R6757 gnd.n7217 gnd.n7216 137.715
R6758 gnd.n7218 gnd.n7217 137.715
R6759 gnd.n7218 gnd.n422 137.715
R6760 gnd.n7226 gnd.n422 137.715
R6761 gnd.n7227 gnd.n7226 137.715
R6762 gnd.n7228 gnd.n7227 137.715
R6763 gnd.n7228 gnd.n416 137.715
R6764 gnd.n7236 gnd.n416 137.715
R6765 gnd.n7237 gnd.n7236 137.715
R6766 gnd.n7238 gnd.n7237 137.715
R6767 gnd.n7238 gnd.n410 137.715
R6768 gnd.n7246 gnd.n410 137.715
R6769 gnd.n7247 gnd.n7246 137.715
R6770 gnd.n7248 gnd.n7247 137.715
R6771 gnd.n7248 gnd.n404 137.715
R6772 gnd.n7256 gnd.n404 137.715
R6773 gnd.n7257 gnd.n7256 137.715
R6774 gnd.n7258 gnd.n7257 137.715
R6775 gnd.n7258 gnd.n398 137.715
R6776 gnd.n7266 gnd.n398 137.715
R6777 gnd.n7267 gnd.n7266 137.715
R6778 gnd.n7269 gnd.n7267 137.715
R6779 gnd.n7269 gnd.n7268 137.715
R6780 gnd.n1197 gnd.t206 130.484
R6781 gnd.n1206 gnd.t227 126.766
R6782 gnd.n1204 gnd.t159 126.766
R6783 gnd.n1190 gnd.t218 126.766
R6784 gnd.n1198 gnd.t179 126.766
R6785 gnd.n5572 gnd.t129 126.766
R6786 gnd.n5574 gnd.t243 126.766
R6787 gnd.n5583 gnd.t192 126.766
R6788 gnd.n5585 gnd.t176 126.766
R6789 gnd.n3617 gnd.n3616 104.615
R6790 gnd.n3616 gnd.n3594 104.615
R6791 gnd.n3609 gnd.n3594 104.615
R6792 gnd.n3609 gnd.n3608 104.615
R6793 gnd.n3608 gnd.n3598 104.615
R6794 gnd.n3601 gnd.n3598 104.615
R6795 gnd.n3585 gnd.n3584 104.615
R6796 gnd.n3584 gnd.n3562 104.615
R6797 gnd.n3577 gnd.n3562 104.615
R6798 gnd.n3577 gnd.n3576 104.615
R6799 gnd.n3576 gnd.n3566 104.615
R6800 gnd.n3569 gnd.n3566 104.615
R6801 gnd.n3553 gnd.n3552 104.615
R6802 gnd.n3552 gnd.n3530 104.615
R6803 gnd.n3545 gnd.n3530 104.615
R6804 gnd.n3545 gnd.n3544 104.615
R6805 gnd.n3544 gnd.n3534 104.615
R6806 gnd.n3537 gnd.n3534 104.615
R6807 gnd.n3522 gnd.n3521 104.615
R6808 gnd.n3521 gnd.n3499 104.615
R6809 gnd.n3514 gnd.n3499 104.615
R6810 gnd.n3514 gnd.n3513 104.615
R6811 gnd.n3513 gnd.n3503 104.615
R6812 gnd.n3506 gnd.n3503 104.615
R6813 gnd.n3490 gnd.n3489 104.615
R6814 gnd.n3489 gnd.n3467 104.615
R6815 gnd.n3482 gnd.n3467 104.615
R6816 gnd.n3482 gnd.n3481 104.615
R6817 gnd.n3481 gnd.n3471 104.615
R6818 gnd.n3474 gnd.n3471 104.615
R6819 gnd.n3458 gnd.n3457 104.615
R6820 gnd.n3457 gnd.n3435 104.615
R6821 gnd.n3450 gnd.n3435 104.615
R6822 gnd.n3450 gnd.n3449 104.615
R6823 gnd.n3449 gnd.n3439 104.615
R6824 gnd.n3442 gnd.n3439 104.615
R6825 gnd.n3426 gnd.n3425 104.615
R6826 gnd.n3425 gnd.n3403 104.615
R6827 gnd.n3418 gnd.n3403 104.615
R6828 gnd.n3418 gnd.n3417 104.615
R6829 gnd.n3417 gnd.n3407 104.615
R6830 gnd.n3410 gnd.n3407 104.615
R6831 gnd.n3395 gnd.n3394 104.615
R6832 gnd.n3394 gnd.n3372 104.615
R6833 gnd.n3387 gnd.n3372 104.615
R6834 gnd.n3387 gnd.n3386 104.615
R6835 gnd.n3386 gnd.n3376 104.615
R6836 gnd.n3379 gnd.n3376 104.615
R6837 gnd.n2769 gnd.t205 100.632
R6838 gnd.n2311 gnd.t235 100.632
R6839 gnd.n7556 gnd.n217 99.6594
R6840 gnd.n7554 gnd.n7553 99.6594
R6841 gnd.n7549 gnd.n224 99.6594
R6842 gnd.n7547 gnd.n7546 99.6594
R6843 gnd.n7542 gnd.n231 99.6594
R6844 gnd.n7540 gnd.n7539 99.6594
R6845 gnd.n7535 gnd.n238 99.6594
R6846 gnd.n7533 gnd.n7532 99.6594
R6847 gnd.n7525 gnd.n245 99.6594
R6848 gnd.n7523 gnd.n7522 99.6594
R6849 gnd.n7518 gnd.n252 99.6594
R6850 gnd.n7516 gnd.n7515 99.6594
R6851 gnd.n7511 gnd.n259 99.6594
R6852 gnd.n7509 gnd.n7508 99.6594
R6853 gnd.n7504 gnd.n266 99.6594
R6854 gnd.n7502 gnd.n7501 99.6594
R6855 gnd.n7497 gnd.n273 99.6594
R6856 gnd.n7495 gnd.n7494 99.6594
R6857 gnd.n283 gnd.n282 99.6594
R6858 gnd.n7486 gnd.n7485 99.6594
R6859 gnd.n7483 gnd.n7482 99.6594
R6860 gnd.n7478 gnd.n291 99.6594
R6861 gnd.n7476 gnd.n7475 99.6594
R6862 gnd.n7471 gnd.n298 99.6594
R6863 gnd.n7469 gnd.n7468 99.6594
R6864 gnd.n7464 gnd.n305 99.6594
R6865 gnd.n7462 gnd.n7461 99.6594
R6866 gnd.n7457 gnd.n314 99.6594
R6867 gnd.n7455 gnd.n7454 99.6594
R6868 gnd.n5754 gnd.n1342 99.6594
R6869 gnd.n5758 gnd.n5757 99.6594
R6870 gnd.n5765 gnd.n5764 99.6594
R6871 gnd.n5768 gnd.n5767 99.6594
R6872 gnd.n5775 gnd.n5774 99.6594
R6873 gnd.n5778 gnd.n5777 99.6594
R6874 gnd.n5785 gnd.n5784 99.6594
R6875 gnd.n5788 gnd.n5787 99.6594
R6876 gnd.n5798 gnd.n5797 99.6594
R6877 gnd.n5801 gnd.n5800 99.6594
R6878 gnd.n5808 gnd.n5807 99.6594
R6879 gnd.n5811 gnd.n5810 99.6594
R6880 gnd.n5819 gnd.n5818 99.6594
R6881 gnd.n5824 gnd.n5823 99.6594
R6882 gnd.n5831 gnd.n5830 99.6594
R6883 gnd.n5834 gnd.n5833 99.6594
R6884 gnd.n5841 gnd.n5840 99.6594
R6885 gnd.n5844 gnd.n5843 99.6594
R6886 gnd.n5853 gnd.n5852 99.6594
R6887 gnd.n5856 gnd.n5855 99.6594
R6888 gnd.n5863 gnd.n5862 99.6594
R6889 gnd.n5866 gnd.n5865 99.6594
R6890 gnd.n5873 gnd.n5872 99.6594
R6891 gnd.n5876 gnd.n5875 99.6594
R6892 gnd.n5883 gnd.n5882 99.6594
R6893 gnd.n5886 gnd.n5885 99.6594
R6894 gnd.n5894 gnd.n5893 99.6594
R6895 gnd.n5897 gnd.n5896 99.6594
R6896 gnd.n6373 gnd.n6372 99.6594
R6897 gnd.n6370 gnd.n6369 99.6594
R6898 gnd.n6365 gnd.n1109 99.6594
R6899 gnd.n6363 gnd.n6362 99.6594
R6900 gnd.n6358 gnd.n1116 99.6594
R6901 gnd.n6356 gnd.n6355 99.6594
R6902 gnd.n6351 gnd.n1123 99.6594
R6903 gnd.n6349 gnd.n6348 99.6594
R6904 gnd.n6343 gnd.n1132 99.6594
R6905 gnd.n6341 gnd.n6340 99.6594
R6906 gnd.n6336 gnd.n1139 99.6594
R6907 gnd.n6334 gnd.n6333 99.6594
R6908 gnd.n4459 gnd.n4458 99.6594
R6909 gnd.n4463 gnd.n4461 99.6594
R6910 gnd.n4469 gnd.n4453 99.6594
R6911 gnd.n4473 gnd.n4471 99.6594
R6912 gnd.n4479 gnd.n4449 99.6594
R6913 gnd.n4483 gnd.n4481 99.6594
R6914 gnd.n4489 gnd.n4443 99.6594
R6915 gnd.n4493 gnd.n4491 99.6594
R6916 gnd.n4499 gnd.n4439 99.6594
R6917 gnd.n4503 gnd.n4501 99.6594
R6918 gnd.n4509 gnd.n4435 99.6594
R6919 gnd.n4513 gnd.n4511 99.6594
R6920 gnd.n4519 gnd.n4431 99.6594
R6921 gnd.n4523 gnd.n4521 99.6594
R6922 gnd.n4529 gnd.n4427 99.6594
R6923 gnd.n4532 gnd.n4531 99.6594
R6924 gnd.n4042 gnd.n4041 99.6594
R6925 gnd.n4036 gnd.n3750 99.6594
R6926 gnd.n4033 gnd.n3751 99.6594
R6927 gnd.n4029 gnd.n3752 99.6594
R6928 gnd.n4025 gnd.n3753 99.6594
R6929 gnd.n4021 gnd.n3754 99.6594
R6930 gnd.n4017 gnd.n3755 99.6594
R6931 gnd.n4013 gnd.n3756 99.6594
R6932 gnd.n4009 gnd.n3757 99.6594
R6933 gnd.n4004 gnd.n3758 99.6594
R6934 gnd.n4000 gnd.n3759 99.6594
R6935 gnd.n3996 gnd.n3760 99.6594
R6936 gnd.n3992 gnd.n3761 99.6594
R6937 gnd.n3988 gnd.n3762 99.6594
R6938 gnd.n3984 gnd.n3763 99.6594
R6939 gnd.n3980 gnd.n3764 99.6594
R6940 gnd.n3976 gnd.n3765 99.6594
R6941 gnd.n3972 gnd.n3766 99.6594
R6942 gnd.n3968 gnd.n3767 99.6594
R6943 gnd.n3964 gnd.n3768 99.6594
R6944 gnd.n3960 gnd.n3769 99.6594
R6945 gnd.n3956 gnd.n3770 99.6594
R6946 gnd.n3952 gnd.n3771 99.6594
R6947 gnd.n3948 gnd.n3772 99.6594
R6948 gnd.n3944 gnd.n3773 99.6594
R6949 gnd.n3940 gnd.n3774 99.6594
R6950 gnd.n3936 gnd.n3775 99.6594
R6951 gnd.n3932 gnd.n3776 99.6594
R6952 gnd.n4044 gnd.n2271 99.6594
R6953 gnd.n3740 gnd.n2294 99.6594
R6954 gnd.n3738 gnd.n2293 99.6594
R6955 gnd.n3734 gnd.n2292 99.6594
R6956 gnd.n3730 gnd.n2291 99.6594
R6957 gnd.n3726 gnd.n2290 99.6594
R6958 gnd.n3722 gnd.n2289 99.6594
R6959 gnd.n3718 gnd.n2288 99.6594
R6960 gnd.n3650 gnd.n2287 99.6594
R6961 gnd.n2981 gnd.n2712 99.6594
R6962 gnd.n2738 gnd.n2719 99.6594
R6963 gnd.n2740 gnd.n2720 99.6594
R6964 gnd.n2748 gnd.n2721 99.6594
R6965 gnd.n2750 gnd.n2722 99.6594
R6966 gnd.n2758 gnd.n2723 99.6594
R6967 gnd.n2760 gnd.n2724 99.6594
R6968 gnd.n2768 gnd.n2725 99.6594
R6969 gnd.n7446 gnd.n320 99.6594
R6970 gnd.n7444 gnd.n7443 99.6594
R6971 gnd.n7439 gnd.n327 99.6594
R6972 gnd.n7437 gnd.n7436 99.6594
R6973 gnd.n7432 gnd.n334 99.6594
R6974 gnd.n7430 gnd.n7429 99.6594
R6975 gnd.n7425 gnd.n341 99.6594
R6976 gnd.n7423 gnd.n7422 99.6594
R6977 gnd.n346 gnd.n345 99.6594
R6978 gnd.n5446 gnd.n5445 99.6594
R6979 gnd.n5462 gnd.n5461 99.6594
R6980 gnd.n5465 gnd.n5464 99.6594
R6981 gnd.n5481 gnd.n5480 99.6594
R6982 gnd.n5484 gnd.n5483 99.6594
R6983 gnd.n5500 gnd.n5499 99.6594
R6984 gnd.n5503 gnd.n5502 99.6594
R6985 gnd.n5520 gnd.n5519 99.6594
R6986 gnd.n5523 gnd.n5522 99.6594
R6987 gnd.n3708 gnd.n2274 99.6594
R6988 gnd.n3704 gnd.n2275 99.6594
R6989 gnd.n3700 gnd.n2276 99.6594
R6990 gnd.n3696 gnd.n2277 99.6594
R6991 gnd.n3692 gnd.n2278 99.6594
R6992 gnd.n3688 gnd.n2279 99.6594
R6993 gnd.n3684 gnd.n2280 99.6594
R6994 gnd.n3680 gnd.n2281 99.6594
R6995 gnd.n3676 gnd.n2282 99.6594
R6996 gnd.n3672 gnd.n2283 99.6594
R6997 gnd.n3668 gnd.n2284 99.6594
R6998 gnd.n3664 gnd.n2285 99.6594
R6999 gnd.n3660 gnd.n2286 99.6594
R7000 gnd.n2896 gnd.n2895 99.6594
R7001 gnd.n2890 gnd.n2807 99.6594
R7002 gnd.n2887 gnd.n2808 99.6594
R7003 gnd.n2883 gnd.n2809 99.6594
R7004 gnd.n2879 gnd.n2810 99.6594
R7005 gnd.n2875 gnd.n2811 99.6594
R7006 gnd.n2871 gnd.n2812 99.6594
R7007 gnd.n2867 gnd.n2813 99.6594
R7008 gnd.n2863 gnd.n2814 99.6594
R7009 gnd.n2859 gnd.n2815 99.6594
R7010 gnd.n2855 gnd.n2816 99.6594
R7011 gnd.n2851 gnd.n2817 99.6594
R7012 gnd.n2898 gnd.n2806 99.6594
R7013 gnd.n4547 gnd.n4546 99.6594
R7014 gnd.n4558 gnd.n4557 99.6594
R7015 gnd.n4567 gnd.n4566 99.6594
R7016 gnd.n4570 gnd.n4569 99.6594
R7017 gnd.n4581 gnd.n4580 99.6594
R7018 gnd.n4590 gnd.n4589 99.6594
R7019 gnd.n4594 gnd.n4592 99.6594
R7020 gnd.n4662 gnd.n2078 99.6594
R7021 gnd.n4665 gnd.n4664 99.6594
R7022 gnd.n3922 gnd.n3777 99.6594
R7023 gnd.n3919 gnd.n3778 99.6594
R7024 gnd.n3915 gnd.n3779 99.6594
R7025 gnd.n3911 gnd.n3780 99.6594
R7026 gnd.n3907 gnd.n3781 99.6594
R7027 gnd.n3903 gnd.n3782 99.6594
R7028 gnd.n3899 gnd.n3783 99.6594
R7029 gnd.n3895 gnd.n3784 99.6594
R7030 gnd.n3891 gnd.n3785 99.6594
R7031 gnd.n3920 gnd.n3777 99.6594
R7032 gnd.n3916 gnd.n3778 99.6594
R7033 gnd.n3912 gnd.n3779 99.6594
R7034 gnd.n3908 gnd.n3780 99.6594
R7035 gnd.n3904 gnd.n3781 99.6594
R7036 gnd.n3900 gnd.n3782 99.6594
R7037 gnd.n3896 gnd.n3783 99.6594
R7038 gnd.n3892 gnd.n3784 99.6594
R7039 gnd.n3867 gnd.n3785 99.6594
R7040 gnd.n4664 gnd.n4663 99.6594
R7041 gnd.n4593 gnd.n2078 99.6594
R7042 gnd.n4592 gnd.n4591 99.6594
R7043 gnd.n4589 gnd.n4582 99.6594
R7044 gnd.n4580 gnd.n4579 99.6594
R7045 gnd.n4569 gnd.n4568 99.6594
R7046 gnd.n4566 gnd.n4559 99.6594
R7047 gnd.n4557 gnd.n4556 99.6594
R7048 gnd.n4546 gnd.n4545 99.6594
R7049 gnd.n2896 gnd.n2819 99.6594
R7050 gnd.n2888 gnd.n2807 99.6594
R7051 gnd.n2884 gnd.n2808 99.6594
R7052 gnd.n2880 gnd.n2809 99.6594
R7053 gnd.n2876 gnd.n2810 99.6594
R7054 gnd.n2872 gnd.n2811 99.6594
R7055 gnd.n2868 gnd.n2812 99.6594
R7056 gnd.n2864 gnd.n2813 99.6594
R7057 gnd.n2860 gnd.n2814 99.6594
R7058 gnd.n2856 gnd.n2815 99.6594
R7059 gnd.n2852 gnd.n2816 99.6594
R7060 gnd.n2848 gnd.n2817 99.6594
R7061 gnd.n2899 gnd.n2898 99.6594
R7062 gnd.n3663 gnd.n2286 99.6594
R7063 gnd.n3667 gnd.n2285 99.6594
R7064 gnd.n3671 gnd.n2284 99.6594
R7065 gnd.n3675 gnd.n2283 99.6594
R7066 gnd.n3679 gnd.n2282 99.6594
R7067 gnd.n3683 gnd.n2281 99.6594
R7068 gnd.n3687 gnd.n2280 99.6594
R7069 gnd.n3691 gnd.n2279 99.6594
R7070 gnd.n3695 gnd.n2278 99.6594
R7071 gnd.n3699 gnd.n2277 99.6594
R7072 gnd.n3703 gnd.n2276 99.6594
R7073 gnd.n3707 gnd.n2275 99.6594
R7074 gnd.n2315 gnd.n2274 99.6594
R7075 gnd.n5445 gnd.n5410 99.6594
R7076 gnd.n5463 gnd.n5462 99.6594
R7077 gnd.n5464 gnd.n5401 99.6594
R7078 gnd.n5482 gnd.n5481 99.6594
R7079 gnd.n5483 gnd.n5392 99.6594
R7080 gnd.n5501 gnd.n5500 99.6594
R7081 gnd.n5502 gnd.n5383 99.6594
R7082 gnd.n5521 gnd.n5520 99.6594
R7083 gnd.n5522 gnd.n5379 99.6594
R7084 gnd.n345 gnd.n342 99.6594
R7085 gnd.n7424 gnd.n7423 99.6594
R7086 gnd.n341 gnd.n335 99.6594
R7087 gnd.n7431 gnd.n7430 99.6594
R7088 gnd.n334 gnd.n328 99.6594
R7089 gnd.n7438 gnd.n7437 99.6594
R7090 gnd.n327 gnd.n321 99.6594
R7091 gnd.n7445 gnd.n7444 99.6594
R7092 gnd.n320 gnd.n317 99.6594
R7093 gnd.n2982 gnd.n2981 99.6594
R7094 gnd.n2741 gnd.n2719 99.6594
R7095 gnd.n2747 gnd.n2720 99.6594
R7096 gnd.n2751 gnd.n2721 99.6594
R7097 gnd.n2757 gnd.n2722 99.6594
R7098 gnd.n2761 gnd.n2723 99.6594
R7099 gnd.n2767 gnd.n2724 99.6594
R7100 gnd.n2725 gnd.n2709 99.6594
R7101 gnd.n3717 gnd.n2287 99.6594
R7102 gnd.n3721 gnd.n2288 99.6594
R7103 gnd.n3725 gnd.n2289 99.6594
R7104 gnd.n3729 gnd.n2290 99.6594
R7105 gnd.n3733 gnd.n2291 99.6594
R7106 gnd.n3737 gnd.n2292 99.6594
R7107 gnd.n3741 gnd.n2293 99.6594
R7108 gnd.n2296 gnd.n2294 99.6594
R7109 gnd.n4042 gnd.n3788 99.6594
R7110 gnd.n4034 gnd.n3750 99.6594
R7111 gnd.n4030 gnd.n3751 99.6594
R7112 gnd.n4026 gnd.n3752 99.6594
R7113 gnd.n4022 gnd.n3753 99.6594
R7114 gnd.n4018 gnd.n3754 99.6594
R7115 gnd.n4014 gnd.n3755 99.6594
R7116 gnd.n4010 gnd.n3756 99.6594
R7117 gnd.n4005 gnd.n3757 99.6594
R7118 gnd.n4001 gnd.n3758 99.6594
R7119 gnd.n3997 gnd.n3759 99.6594
R7120 gnd.n3993 gnd.n3760 99.6594
R7121 gnd.n3989 gnd.n3761 99.6594
R7122 gnd.n3985 gnd.n3762 99.6594
R7123 gnd.n3981 gnd.n3763 99.6594
R7124 gnd.n3977 gnd.n3764 99.6594
R7125 gnd.n3973 gnd.n3765 99.6594
R7126 gnd.n3969 gnd.n3766 99.6594
R7127 gnd.n3965 gnd.n3767 99.6594
R7128 gnd.n3961 gnd.n3768 99.6594
R7129 gnd.n3957 gnd.n3769 99.6594
R7130 gnd.n3953 gnd.n3770 99.6594
R7131 gnd.n3949 gnd.n3771 99.6594
R7132 gnd.n3945 gnd.n3772 99.6594
R7133 gnd.n3941 gnd.n3773 99.6594
R7134 gnd.n3937 gnd.n3774 99.6594
R7135 gnd.n3933 gnd.n3775 99.6594
R7136 gnd.n3929 gnd.n3776 99.6594
R7137 gnd.n4045 gnd.n4044 99.6594
R7138 gnd.n4531 gnd.n4530 99.6594
R7139 gnd.n4522 gnd.n4427 99.6594
R7140 gnd.n4521 gnd.n4520 99.6594
R7141 gnd.n4512 gnd.n4431 99.6594
R7142 gnd.n4511 gnd.n4510 99.6594
R7143 gnd.n4502 gnd.n4435 99.6594
R7144 gnd.n4501 gnd.n4500 99.6594
R7145 gnd.n4492 gnd.n4439 99.6594
R7146 gnd.n4491 gnd.n4490 99.6594
R7147 gnd.n4482 gnd.n4443 99.6594
R7148 gnd.n4481 gnd.n4480 99.6594
R7149 gnd.n4472 gnd.n4449 99.6594
R7150 gnd.n4471 gnd.n4470 99.6594
R7151 gnd.n4462 gnd.n4453 99.6594
R7152 gnd.n4461 gnd.n4460 99.6594
R7153 gnd.n1145 gnd.n1140 99.6594
R7154 gnd.n6335 gnd.n6334 99.6594
R7155 gnd.n1139 gnd.n1133 99.6594
R7156 gnd.n6342 gnd.n6341 99.6594
R7157 gnd.n1132 gnd.n1124 99.6594
R7158 gnd.n6350 gnd.n6349 99.6594
R7159 gnd.n1123 gnd.n1117 99.6594
R7160 gnd.n6357 gnd.n6356 99.6594
R7161 gnd.n1116 gnd.n1110 99.6594
R7162 gnd.n6364 gnd.n6363 99.6594
R7163 gnd.n1109 gnd.n1102 99.6594
R7164 gnd.n6371 gnd.n6370 99.6594
R7165 gnd.n6374 gnd.n6373 99.6594
R7166 gnd.n5755 gnd.n5754 99.6594
R7167 gnd.n5757 gnd.n5746 99.6594
R7168 gnd.n5766 gnd.n5765 99.6594
R7169 gnd.n5767 gnd.n5742 99.6594
R7170 gnd.n5776 gnd.n5775 99.6594
R7171 gnd.n5777 gnd.n5738 99.6594
R7172 gnd.n5786 gnd.n5785 99.6594
R7173 gnd.n5787 gnd.n5734 99.6594
R7174 gnd.n5799 gnd.n5798 99.6594
R7175 gnd.n5800 gnd.n5730 99.6594
R7176 gnd.n5809 gnd.n5808 99.6594
R7177 gnd.n5810 gnd.n5726 99.6594
R7178 gnd.n5822 gnd.n5821 99.6594
R7179 gnd.n5823 gnd.n1528 99.6594
R7180 gnd.n5832 gnd.n5831 99.6594
R7181 gnd.n5833 gnd.n1524 99.6594
R7182 gnd.n5842 gnd.n5841 99.6594
R7183 gnd.n5843 gnd.n1520 99.6594
R7184 gnd.n5854 gnd.n5853 99.6594
R7185 gnd.n5855 gnd.n1516 99.6594
R7186 gnd.n5864 gnd.n5863 99.6594
R7187 gnd.n5865 gnd.n1512 99.6594
R7188 gnd.n5874 gnd.n5873 99.6594
R7189 gnd.n5875 gnd.n1508 99.6594
R7190 gnd.n5884 gnd.n5883 99.6594
R7191 gnd.n5885 gnd.n1504 99.6594
R7192 gnd.n5895 gnd.n5894 99.6594
R7193 gnd.n5898 gnd.n5897 99.6594
R7194 gnd.n7456 gnd.n7455 99.6594
R7195 gnd.n314 gnd.n306 99.6594
R7196 gnd.n7463 gnd.n7462 99.6594
R7197 gnd.n305 gnd.n299 99.6594
R7198 gnd.n7470 gnd.n7469 99.6594
R7199 gnd.n298 gnd.n292 99.6594
R7200 gnd.n7477 gnd.n7476 99.6594
R7201 gnd.n291 gnd.n285 99.6594
R7202 gnd.n7484 gnd.n7483 99.6594
R7203 gnd.n7487 gnd.n7486 99.6594
R7204 gnd.n282 gnd.n274 99.6594
R7205 gnd.n7496 gnd.n7495 99.6594
R7206 gnd.n273 gnd.n267 99.6594
R7207 gnd.n7503 gnd.n7502 99.6594
R7208 gnd.n266 gnd.n260 99.6594
R7209 gnd.n7510 gnd.n7509 99.6594
R7210 gnd.n259 gnd.n253 99.6594
R7211 gnd.n7517 gnd.n7516 99.6594
R7212 gnd.n252 gnd.n246 99.6594
R7213 gnd.n7524 gnd.n7523 99.6594
R7214 gnd.n245 gnd.n239 99.6594
R7215 gnd.n7534 gnd.n7533 99.6594
R7216 gnd.n238 gnd.n232 99.6594
R7217 gnd.n7541 gnd.n7540 99.6594
R7218 gnd.n231 gnd.n225 99.6594
R7219 gnd.n7548 gnd.n7547 99.6594
R7220 gnd.n224 gnd.n218 99.6594
R7221 gnd.n7555 gnd.n7554 99.6594
R7222 gnd.n217 gnd.n214 99.6594
R7223 gnd.n4654 gnd.n4653 99.6594
R7224 gnd.n4419 gnd.n4402 99.6594
R7225 gnd.n4421 gnd.n4403 99.6594
R7226 gnd.n4538 gnd.n4404 99.6594
R7227 gnd.n4540 gnd.n4405 99.6594
R7228 gnd.n4551 gnd.n4406 99.6594
R7229 gnd.n4553 gnd.n4407 99.6594
R7230 gnd.n4563 gnd.n4408 99.6594
R7231 gnd.n4574 gnd.n4409 99.6594
R7232 gnd.n4576 gnd.n4410 99.6594
R7233 gnd.n4586 gnd.n4411 99.6594
R7234 gnd.n4597 gnd.n4412 99.6594
R7235 gnd.n4657 gnd.n4656 99.6594
R7236 gnd.n4413 gnd.n2073 99.6594
R7237 gnd.n4654 gnd.n4415 99.6594
R7238 gnd.n4420 gnd.n4402 99.6594
R7239 gnd.n4537 gnd.n4403 99.6594
R7240 gnd.n4539 gnd.n4404 99.6594
R7241 gnd.n4550 gnd.n4405 99.6594
R7242 gnd.n4552 gnd.n4406 99.6594
R7243 gnd.n4562 gnd.n4407 99.6594
R7244 gnd.n4573 gnd.n4408 99.6594
R7245 gnd.n4575 gnd.n4409 99.6594
R7246 gnd.n4585 gnd.n4410 99.6594
R7247 gnd.n4596 gnd.n4411 99.6594
R7248 gnd.n4412 gnd.n2085 99.6594
R7249 gnd.n4656 gnd.n2086 99.6594
R7250 gnd.n4413 gnd.n2069 99.6594
R7251 gnd.n5426 gnd.n5422 99.6594
R7252 gnd.n5430 gnd.n5428 99.6594
R7253 gnd.n5437 gnd.n5418 99.6594
R7254 gnd.n5441 gnd.n5439 99.6594
R7255 gnd.n5452 gnd.n5415 99.6594
R7256 gnd.n5456 gnd.n5454 99.6594
R7257 gnd.n5471 gnd.n5406 99.6594
R7258 gnd.n5475 gnd.n5473 99.6594
R7259 gnd.n5490 gnd.n5397 99.6594
R7260 gnd.n5494 gnd.n5492 99.6594
R7261 gnd.n5509 gnd.n5388 99.6594
R7262 gnd.n5512 gnd.n5511 99.6594
R7263 gnd.n5530 gnd.n5529 99.6594
R7264 gnd.n5533 gnd.n5532 99.6594
R7265 gnd.n5511 gnd.n5510 99.6594
R7266 gnd.n5493 gnd.n5388 99.6594
R7267 gnd.n5492 gnd.n5491 99.6594
R7268 gnd.n5474 gnd.n5397 99.6594
R7269 gnd.n5473 gnd.n5472 99.6594
R7270 gnd.n5455 gnd.n5406 99.6594
R7271 gnd.n5454 gnd.n5453 99.6594
R7272 gnd.n5440 gnd.n5415 99.6594
R7273 gnd.n5439 gnd.n5438 99.6594
R7274 gnd.n5429 gnd.n5418 99.6594
R7275 gnd.n5428 gnd.n5427 99.6594
R7276 gnd.n5422 gnd.n1316 99.6594
R7277 gnd.n5534 gnd.n5533 99.6594
R7278 gnd.n5531 gnd.n5530 99.6594
R7279 gnd.n2082 gnd.t191 98.63
R7280 gnd.n5380 gnd.t217 98.63
R7281 gnd.n2075 gnd.t241 98.63
R7282 gnd.n5793 gnd.t214 98.63
R7283 gnd.n5845 gnd.t211 98.63
R7284 gnd.n1500 gnd.t143 98.63
R7285 gnd.n311 gnd.t238 98.63
R7286 gnd.n278 gnd.t157 98.63
R7287 gnd.n7527 gnd.t196 98.63
R7288 gnd.n348 gnd.t183 98.63
R7289 gnd.n3807 gnd.t171 98.63
R7290 gnd.n3829 gnd.t168 98.63
R7291 gnd.n3850 gnd.t147 98.63
R7292 gnd.n3868 gnd.t226 98.63
R7293 gnd.n1128 gnd.t231 98.63
R7294 gnd.n4424 gnd.t164 98.63
R7295 gnd.n4446 gnd.t186 98.63
R7296 gnd.n5370 gnd.t174 98.63
R7297 gnd.n1950 gnd.t201 92.8196
R7298 gnd.n1569 gnd.t222 92.8196
R7299 gnd.n6261 gnd.t248 92.8118
R7300 gnd.n5587 gnd.t153 92.8118
R7301 gnd.n7268 gnd.n207 82.6296
R7302 gnd.n1197 gnd.n1196 81.8399
R7303 gnd.n5725 gnd.n5724 78.9125
R7304 gnd.n6330 gnd.n6329 78.9125
R7305 gnd.n2770 gnd.t204 74.8376
R7306 gnd.n2312 gnd.t236 74.8376
R7307 gnd.n1951 gnd.t200 72.8438
R7308 gnd.n1570 gnd.t223 72.8438
R7309 gnd.n1198 gnd.n1191 72.8411
R7310 gnd.n1204 gnd.n1189 72.8411
R7311 gnd.n5583 gnd.n5582 72.8411
R7312 gnd.n2083 gnd.t190 72.836
R7313 gnd.n6262 gnd.t247 72.836
R7314 gnd.n5588 gnd.t154 72.836
R7315 gnd.n5381 gnd.t216 72.836
R7316 gnd.n2076 gnd.t242 72.836
R7317 gnd.n5794 gnd.t213 72.836
R7318 gnd.n5846 gnd.t210 72.836
R7319 gnd.n1501 gnd.t142 72.836
R7320 gnd.n312 gnd.t239 72.836
R7321 gnd.n279 gnd.t158 72.836
R7322 gnd.n7528 gnd.t197 72.836
R7323 gnd.n349 gnd.t184 72.836
R7324 gnd.n3808 gnd.t170 72.836
R7325 gnd.n3830 gnd.t167 72.836
R7326 gnd.n3851 gnd.t146 72.836
R7327 gnd.n3869 gnd.t225 72.836
R7328 gnd.n1129 gnd.t232 72.836
R7329 gnd.n4425 gnd.t165 72.836
R7330 gnd.n4447 gnd.t187 72.836
R7331 gnd.n5371 gnd.t175 72.836
R7332 gnd.n5648 gnd.n1537 71.676
R7333 gnd.n5644 gnd.n1538 71.676
R7334 gnd.n5640 gnd.n1539 71.676
R7335 gnd.n5636 gnd.n1540 71.676
R7336 gnd.n5632 gnd.n1541 71.676
R7337 gnd.n5628 gnd.n1542 71.676
R7338 gnd.n5624 gnd.n1543 71.676
R7339 gnd.n5620 gnd.n1544 71.676
R7340 gnd.n5616 gnd.n1545 71.676
R7341 gnd.n5612 gnd.n1546 71.676
R7342 gnd.n5608 gnd.n1547 71.676
R7343 gnd.n5604 gnd.n1548 71.676
R7344 gnd.n5600 gnd.n1549 71.676
R7345 gnd.n5596 gnd.n1550 71.676
R7346 gnd.n5591 gnd.n1551 71.676
R7347 gnd.n1552 gnd.n1535 71.676
R7348 gnd.n5720 gnd.n1534 71.676
R7349 gnd.n5718 gnd.n5717 71.676
R7350 gnd.n5712 gnd.n1567 71.676
R7351 gnd.n5708 gnd.n1566 71.676
R7352 gnd.n5704 gnd.n1565 71.676
R7353 gnd.n5700 gnd.n1564 71.676
R7354 gnd.n5696 gnd.n1563 71.676
R7355 gnd.n5692 gnd.n1562 71.676
R7356 gnd.n5688 gnd.n1561 71.676
R7357 gnd.n5684 gnd.n1560 71.676
R7358 gnd.n5680 gnd.n1559 71.676
R7359 gnd.n5676 gnd.n1558 71.676
R7360 gnd.n5672 gnd.n1557 71.676
R7361 gnd.n5668 gnd.n1556 71.676
R7362 gnd.n5664 gnd.n1555 71.676
R7363 gnd.n5660 gnd.n1554 71.676
R7364 gnd.n5656 gnd.n1553 71.676
R7365 gnd.n6325 gnd.n6324 71.676
R7366 gnd.n6319 gnd.n1153 71.676
R7367 gnd.n6316 gnd.n1154 71.676
R7368 gnd.n6312 gnd.n1155 71.676
R7369 gnd.n6308 gnd.n1156 71.676
R7370 gnd.n6304 gnd.n1157 71.676
R7371 gnd.n6300 gnd.n1158 71.676
R7372 gnd.n6296 gnd.n1159 71.676
R7373 gnd.n6292 gnd.n1160 71.676
R7374 gnd.n6288 gnd.n1161 71.676
R7375 gnd.n6284 gnd.n1162 71.676
R7376 gnd.n6280 gnd.n1163 71.676
R7377 gnd.n6276 gnd.n1164 71.676
R7378 gnd.n6272 gnd.n1165 71.676
R7379 gnd.n6268 gnd.n1166 71.676
R7380 gnd.n6264 gnd.n1167 71.676
R7381 gnd.n1168 gnd.n1151 71.676
R7382 gnd.n1954 gnd.n1169 71.676
R7383 gnd.n1959 gnd.n1170 71.676
R7384 gnd.n1963 gnd.n1171 71.676
R7385 gnd.n1967 gnd.n1172 71.676
R7386 gnd.n1971 gnd.n1173 71.676
R7387 gnd.n1975 gnd.n1174 71.676
R7388 gnd.n1979 gnd.n1175 71.676
R7389 gnd.n1983 gnd.n1176 71.676
R7390 gnd.n1987 gnd.n1177 71.676
R7391 gnd.n1991 gnd.n1178 71.676
R7392 gnd.n1995 gnd.n1179 71.676
R7393 gnd.n1999 gnd.n1180 71.676
R7394 gnd.n2003 gnd.n1181 71.676
R7395 gnd.n2007 gnd.n1182 71.676
R7396 gnd.n2011 gnd.n1183 71.676
R7397 gnd.n6325 gnd.n1186 71.676
R7398 gnd.n6317 gnd.n1153 71.676
R7399 gnd.n6313 gnd.n1154 71.676
R7400 gnd.n6309 gnd.n1155 71.676
R7401 gnd.n6305 gnd.n1156 71.676
R7402 gnd.n6301 gnd.n1157 71.676
R7403 gnd.n6297 gnd.n1158 71.676
R7404 gnd.n6293 gnd.n1159 71.676
R7405 gnd.n6289 gnd.n1160 71.676
R7406 gnd.n6285 gnd.n1161 71.676
R7407 gnd.n6281 gnd.n1162 71.676
R7408 gnd.n6277 gnd.n1163 71.676
R7409 gnd.n6273 gnd.n1164 71.676
R7410 gnd.n6269 gnd.n1165 71.676
R7411 gnd.n6265 gnd.n1166 71.676
R7412 gnd.n6328 gnd.n6327 71.676
R7413 gnd.n1953 gnd.n1168 71.676
R7414 gnd.n1958 gnd.n1169 71.676
R7415 gnd.n1962 gnd.n1170 71.676
R7416 gnd.n1966 gnd.n1171 71.676
R7417 gnd.n1970 gnd.n1172 71.676
R7418 gnd.n1974 gnd.n1173 71.676
R7419 gnd.n1978 gnd.n1174 71.676
R7420 gnd.n1982 gnd.n1175 71.676
R7421 gnd.n1986 gnd.n1176 71.676
R7422 gnd.n1990 gnd.n1177 71.676
R7423 gnd.n1994 gnd.n1178 71.676
R7424 gnd.n1998 gnd.n1179 71.676
R7425 gnd.n2002 gnd.n1180 71.676
R7426 gnd.n2006 gnd.n1181 71.676
R7427 gnd.n2010 gnd.n1182 71.676
R7428 gnd.n1949 gnd.n1183 71.676
R7429 gnd.n5659 gnd.n1553 71.676
R7430 gnd.n5663 gnd.n1554 71.676
R7431 gnd.n5667 gnd.n1555 71.676
R7432 gnd.n5671 gnd.n1556 71.676
R7433 gnd.n5675 gnd.n1557 71.676
R7434 gnd.n5679 gnd.n1558 71.676
R7435 gnd.n5683 gnd.n1559 71.676
R7436 gnd.n5687 gnd.n1560 71.676
R7437 gnd.n5691 gnd.n1561 71.676
R7438 gnd.n5695 gnd.n1562 71.676
R7439 gnd.n5699 gnd.n1563 71.676
R7440 gnd.n5703 gnd.n1564 71.676
R7441 gnd.n5707 gnd.n1565 71.676
R7442 gnd.n5711 gnd.n1566 71.676
R7443 gnd.n1568 gnd.n1567 71.676
R7444 gnd.n5719 gnd.n5718 71.676
R7445 gnd.n5723 gnd.n5722 71.676
R7446 gnd.n5590 gnd.n1552 71.676
R7447 gnd.n5595 gnd.n1551 71.676
R7448 gnd.n5599 gnd.n1550 71.676
R7449 gnd.n5603 gnd.n1549 71.676
R7450 gnd.n5607 gnd.n1548 71.676
R7451 gnd.n5611 gnd.n1547 71.676
R7452 gnd.n5615 gnd.n1546 71.676
R7453 gnd.n5619 gnd.n1545 71.676
R7454 gnd.n5623 gnd.n1544 71.676
R7455 gnd.n5627 gnd.n1543 71.676
R7456 gnd.n5631 gnd.n1542 71.676
R7457 gnd.n5635 gnd.n1541 71.676
R7458 gnd.n5639 gnd.n1540 71.676
R7459 gnd.n5643 gnd.n1539 71.676
R7460 gnd.n5647 gnd.n1538 71.676
R7461 gnd.n1575 gnd.n1537 71.676
R7462 gnd.n8 gnd.t11 69.1507
R7463 gnd.n14 gnd.t283 68.4792
R7464 gnd.n13 gnd.t345 68.4792
R7465 gnd.n12 gnd.t29 68.4792
R7466 gnd.n11 gnd.t254 68.4792
R7467 gnd.n10 gnd.t365 68.4792
R7468 gnd.n9 gnd.t363 68.4792
R7469 gnd.n8 gnd.t355 68.4792
R7470 gnd.n2897 gnd.n2801 64.369
R7471 gnd.n1956 gnd.n1951 59.5399
R7472 gnd.n5714 gnd.n1570 59.5399
R7473 gnd.n6263 gnd.n6262 59.5399
R7474 gnd.n5593 gnd.n5588 59.5399
R7475 gnd.n6260 gnd.n1207 59.1804
R7476 gnd.n3749 gnd.n2272 57.3586
R7477 gnd.n4043 gnd.n2259 57.3586
R7478 gnd.n7564 gnd.n210 57.3586
R7479 gnd.n2552 gnd.t277 56.407
R7480 gnd.n2505 gnd.t318 56.407
R7481 gnd.n2520 gnd.t80 56.407
R7482 gnd.n2536 gnd.t350 56.407
R7483 gnd.n64 gnd.t256 56.407
R7484 gnd.n17 gnd.t295 56.407
R7485 gnd.n32 gnd.t13 56.407
R7486 gnd.n48 gnd.t317 56.407
R7487 gnd.n2565 gnd.t57 55.8337
R7488 gnd.n2518 gnd.t275 55.8337
R7489 gnd.n2533 gnd.t121 55.8337
R7490 gnd.n2549 gnd.t99 55.8337
R7491 gnd.n77 gnd.t278 55.8337
R7492 gnd.n30 gnd.t309 55.8337
R7493 gnd.n45 gnd.t366 55.8337
R7494 gnd.n61 gnd.t85 55.8337
R7495 gnd.n1195 gnd.n1194 54.358
R7496 gnd.n5580 gnd.n5579 54.358
R7497 gnd.n2552 gnd.n2551 53.0052
R7498 gnd.n2554 gnd.n2553 53.0052
R7499 gnd.n2556 gnd.n2555 53.0052
R7500 gnd.n2558 gnd.n2557 53.0052
R7501 gnd.n2560 gnd.n2559 53.0052
R7502 gnd.n2562 gnd.n2561 53.0052
R7503 gnd.n2564 gnd.n2563 53.0052
R7504 gnd.n2505 gnd.n2504 53.0052
R7505 gnd.n2507 gnd.n2506 53.0052
R7506 gnd.n2509 gnd.n2508 53.0052
R7507 gnd.n2511 gnd.n2510 53.0052
R7508 gnd.n2513 gnd.n2512 53.0052
R7509 gnd.n2515 gnd.n2514 53.0052
R7510 gnd.n2517 gnd.n2516 53.0052
R7511 gnd.n2520 gnd.n2519 53.0052
R7512 gnd.n2522 gnd.n2521 53.0052
R7513 gnd.n2524 gnd.n2523 53.0052
R7514 gnd.n2526 gnd.n2525 53.0052
R7515 gnd.n2528 gnd.n2527 53.0052
R7516 gnd.n2530 gnd.n2529 53.0052
R7517 gnd.n2532 gnd.n2531 53.0052
R7518 gnd.n2536 gnd.n2535 53.0052
R7519 gnd.n2538 gnd.n2537 53.0052
R7520 gnd.n2540 gnd.n2539 53.0052
R7521 gnd.n2542 gnd.n2541 53.0052
R7522 gnd.n2544 gnd.n2543 53.0052
R7523 gnd.n2546 gnd.n2545 53.0052
R7524 gnd.n2548 gnd.n2547 53.0052
R7525 gnd.n76 gnd.n75 53.0052
R7526 gnd.n74 gnd.n73 53.0052
R7527 gnd.n72 gnd.n71 53.0052
R7528 gnd.n70 gnd.n69 53.0052
R7529 gnd.n68 gnd.n67 53.0052
R7530 gnd.n66 gnd.n65 53.0052
R7531 gnd.n64 gnd.n63 53.0052
R7532 gnd.n29 gnd.n28 53.0052
R7533 gnd.n27 gnd.n26 53.0052
R7534 gnd.n25 gnd.n24 53.0052
R7535 gnd.n23 gnd.n22 53.0052
R7536 gnd.n21 gnd.n20 53.0052
R7537 gnd.n19 gnd.n18 53.0052
R7538 gnd.n17 gnd.n16 53.0052
R7539 gnd.n44 gnd.n43 53.0052
R7540 gnd.n42 gnd.n41 53.0052
R7541 gnd.n40 gnd.n39 53.0052
R7542 gnd.n38 gnd.n37 53.0052
R7543 gnd.n36 gnd.n35 53.0052
R7544 gnd.n34 gnd.n33 53.0052
R7545 gnd.n32 gnd.n31 53.0052
R7546 gnd.n60 gnd.n59 53.0052
R7547 gnd.n58 gnd.n57 53.0052
R7548 gnd.n56 gnd.n55 53.0052
R7549 gnd.n54 gnd.n53 53.0052
R7550 gnd.n52 gnd.n51 53.0052
R7551 gnd.n50 gnd.n49 53.0052
R7552 gnd.n48 gnd.n47 53.0052
R7553 gnd.n5571 gnd.n5570 52.4801
R7554 gnd.n3601 gnd.t68 52.3082
R7555 gnd.n3569 gnd.t289 52.3082
R7556 gnd.n3537 gnd.t115 52.3082
R7557 gnd.n3506 gnd.t93 52.3082
R7558 gnd.n3474 gnd.t298 52.3082
R7559 gnd.n3442 gnd.t78 52.3082
R7560 gnd.n3410 gnd.t273 52.3082
R7561 gnd.n3379 gnd.t31 52.3082
R7562 gnd.n3431 gnd.n3399 51.4173
R7563 gnd.n3495 gnd.n3494 50.455
R7564 gnd.n3463 gnd.n3462 50.455
R7565 gnd.n3431 gnd.n3430 50.455
R7566 gnd.n2844 gnd.n2843 45.1884
R7567 gnd.n2338 gnd.n2337 45.1884
R7568 gnd.n5651 gnd.n5586 44.3322
R7569 gnd.n1198 gnd.n1197 44.3189
R7570 gnd.n2084 gnd.n2083 42.2793
R7571 gnd.n5525 gnd.n5381 42.2793
R7572 gnd.n2845 gnd.n2844 42.2793
R7573 gnd.n2339 gnd.n2338 42.2793
R7574 gnd.n2771 gnd.n2770 42.2793
R7575 gnd.n3716 gnd.n2312 42.2793
R7576 gnd.n2077 gnd.n2076 42.2793
R7577 gnd.n5795 gnd.n5794 42.2793
R7578 gnd.n5847 gnd.n5846 42.2793
R7579 gnd.n1502 gnd.n1501 42.2793
R7580 gnd.n313 gnd.n312 42.2793
R7581 gnd.n7492 gnd.n279 42.2793
R7582 gnd.n7529 gnd.n7528 42.2793
R7583 gnd.n7420 gnd.n349 42.2793
R7584 gnd.n4007 gnd.n3808 42.2793
R7585 gnd.n3967 gnd.n3830 42.2793
R7586 gnd.n3928 gnd.n3851 42.2793
R7587 gnd.n3870 gnd.n3869 42.2793
R7588 gnd.n6345 gnd.n1129 42.2793
R7589 gnd.n4426 gnd.n4425 42.2793
R7590 gnd.n4448 gnd.n4447 42.2793
R7591 gnd.n5372 gnd.n5371 42.2793
R7592 gnd.n1196 gnd.n1195 41.6274
R7593 gnd.n5581 gnd.n5580 41.6274
R7594 gnd.n1205 gnd.n1204 40.8975
R7595 gnd.n5584 gnd.n5583 40.8975
R7596 gnd.n6637 gnd.n769 37.4091
R7597 gnd.n6637 gnd.n6636 37.4091
R7598 gnd.n6636 gnd.n6635 37.4091
R7599 gnd.n6635 gnd.n774 37.4091
R7600 gnd.n6629 gnd.n774 37.4091
R7601 gnd.n6629 gnd.n6628 37.4091
R7602 gnd.n6628 gnd.n6627 37.4091
R7603 gnd.n6627 gnd.n782 37.4091
R7604 gnd.n6621 gnd.n782 37.4091
R7605 gnd.n6621 gnd.n6620 37.4091
R7606 gnd.n6620 gnd.n6619 37.4091
R7607 gnd.n6619 gnd.n790 37.4091
R7608 gnd.n6613 gnd.n790 37.4091
R7609 gnd.n6613 gnd.n6612 37.4091
R7610 gnd.n6612 gnd.n6611 37.4091
R7611 gnd.n6611 gnd.n798 37.4091
R7612 gnd.n6605 gnd.n798 37.4091
R7613 gnd.n6605 gnd.n6604 37.4091
R7614 gnd.n6604 gnd.n6603 37.4091
R7615 gnd.n6603 gnd.n806 37.4091
R7616 gnd.n6597 gnd.n806 37.4091
R7617 gnd.n6597 gnd.n6596 37.4091
R7618 gnd.n6596 gnd.n6595 37.4091
R7619 gnd.n6595 gnd.n814 37.4091
R7620 gnd.n6589 gnd.n814 37.4091
R7621 gnd.n6589 gnd.n6588 37.4091
R7622 gnd.n6588 gnd.n6587 37.4091
R7623 gnd.n6587 gnd.n822 37.4091
R7624 gnd.n6581 gnd.n822 37.4091
R7625 gnd.n6581 gnd.n6580 37.4091
R7626 gnd.n6580 gnd.n6579 37.4091
R7627 gnd.n6579 gnd.n830 37.4091
R7628 gnd.n6573 gnd.n830 37.4091
R7629 gnd.n6573 gnd.n6572 37.4091
R7630 gnd.n6572 gnd.n6571 37.4091
R7631 gnd.n6571 gnd.n838 37.4091
R7632 gnd.n6565 gnd.n838 37.4091
R7633 gnd.n6565 gnd.n6564 37.4091
R7634 gnd.n6564 gnd.n6563 37.4091
R7635 gnd.n6563 gnd.n846 37.4091
R7636 gnd.n6557 gnd.n846 37.4091
R7637 gnd.n6557 gnd.n6556 37.4091
R7638 gnd.n6556 gnd.n6555 37.4091
R7639 gnd.n6555 gnd.n854 37.4091
R7640 gnd.n6549 gnd.n854 37.4091
R7641 gnd.n6549 gnd.n6548 37.4091
R7642 gnd.n6548 gnd.n6547 37.4091
R7643 gnd.n6547 gnd.n862 37.4091
R7644 gnd.n6541 gnd.n862 37.4091
R7645 gnd.n6541 gnd.n6540 37.4091
R7646 gnd.n6540 gnd.n6539 37.4091
R7647 gnd.n6539 gnd.n870 37.4091
R7648 gnd.n6533 gnd.n870 37.4091
R7649 gnd.n6533 gnd.n6532 37.4091
R7650 gnd.n6532 gnd.n6531 37.4091
R7651 gnd.n6531 gnd.n878 37.4091
R7652 gnd.n6525 gnd.n878 37.4091
R7653 gnd.n6525 gnd.n6524 37.4091
R7654 gnd.n6524 gnd.n6523 37.4091
R7655 gnd.n6523 gnd.n886 37.4091
R7656 gnd.n6517 gnd.n886 37.4091
R7657 gnd.n6517 gnd.n6516 37.4091
R7658 gnd.n6516 gnd.n6515 37.4091
R7659 gnd.n6515 gnd.n894 37.4091
R7660 gnd.n6509 gnd.n894 37.4091
R7661 gnd.n6509 gnd.n6508 37.4091
R7662 gnd.n6508 gnd.n6507 37.4091
R7663 gnd.n6507 gnd.n902 37.4091
R7664 gnd.n6501 gnd.n902 37.4091
R7665 gnd.n6501 gnd.n6500 37.4091
R7666 gnd.n6500 gnd.n6499 37.4091
R7667 gnd.n6499 gnd.n910 37.4091
R7668 gnd.n6493 gnd.n910 37.4091
R7669 gnd.n6493 gnd.n6492 37.4091
R7670 gnd.n6492 gnd.n6491 37.4091
R7671 gnd.n6491 gnd.n918 37.4091
R7672 gnd.n6485 gnd.n918 37.4091
R7673 gnd.n6485 gnd.n6484 37.4091
R7674 gnd.n6484 gnd.n6483 37.4091
R7675 gnd.n6483 gnd.n926 37.4091
R7676 gnd.n6477 gnd.n926 37.4091
R7677 gnd.n6477 gnd.n6476 37.4091
R7678 gnd.n6476 gnd.n6475 37.4091
R7679 gnd.n1204 gnd.n1203 35.055
R7680 gnd.n1199 gnd.n1198 35.055
R7681 gnd.n5573 gnd.n5572 35.055
R7682 gnd.n5583 gnd.n5569 35.055
R7683 gnd.n2907 gnd.n2801 31.8661
R7684 gnd.n2907 gnd.n2906 31.8661
R7685 gnd.n2915 gnd.n2790 31.8661
R7686 gnd.n2923 gnd.n2790 31.8661
R7687 gnd.n2923 gnd.n2784 31.8661
R7688 gnd.n2931 gnd.n2784 31.8661
R7689 gnd.n2931 gnd.n2777 31.8661
R7690 gnd.n2969 gnd.n2777 31.8661
R7691 gnd.n2979 gnd.n2710 31.8661
R7692 gnd.n4053 gnd.n2259 31.8661
R7693 gnd.n4061 gnd.n2251 31.8661
R7694 gnd.n4061 gnd.n2239 31.8661
R7695 gnd.n4077 gnd.n2239 31.8661
R7696 gnd.n4077 gnd.n2242 31.8661
R7697 gnd.n4087 gnd.n2225 31.8661
R7698 gnd.n4099 gnd.n2225 31.8661
R7699 gnd.n4113 gnd.n2215 31.8661
R7700 gnd.n4121 gnd.n2191 31.8661
R7701 gnd.n4143 gnd.n2191 31.8661
R7702 gnd.n4152 gnd.n941 31.8661
R7703 gnd.n4391 gnd.n1095 31.8661
R7704 gnd.n4393 gnd.n2087 31.8661
R7705 gnd.n4401 gnd.n2087 31.8661
R7706 gnd.n4677 gnd.n2068 31.8661
R7707 gnd.n6137 gnd.n1319 31.8661
R7708 gnd.n6131 gnd.n6130 31.8661
R7709 gnd.n6130 gnd.n6129 31.8661
R7710 gnd.n6123 gnd.n1337 31.8661
R7711 gnd.n7612 gnd.n132 31.8661
R7712 gnd.n7606 gnd.n145 31.8661
R7713 gnd.n7600 gnd.n145 31.8661
R7714 gnd.n7594 gnd.n161 31.8661
R7715 gnd.n7588 gnd.n170 31.8661
R7716 gnd.n7588 gnd.n173 31.8661
R7717 gnd.n7582 gnd.n183 31.8661
R7718 gnd.n7576 gnd.n183 31.8661
R7719 gnd.n7576 gnd.n192 31.8661
R7720 gnd.n7570 gnd.n192 31.8661
R7721 gnd.n5657 gnd.n1571 31.3761
R7722 gnd.n2024 gnd.n2013 31.3761
R7723 gnd.n2215 gnd.t262 27.7236
R7724 gnd.n161 gnd.t39 27.7236
R7725 gnd.n4190 gnd.n944 26.7676
R7726 gnd.n4184 gnd.n956 26.7676
R7727 gnd.n6454 gnd.n965 26.7676
R7728 gnd.n4177 gnd.n4176 26.7676
R7729 gnd.n4222 gnd.n2159 26.7676
R7730 gnd.n4216 gnd.n2155 26.7676
R7731 gnd.n4241 gnd.n2145 26.7676
R7732 gnd.n4277 gnd.n2131 26.7676
R7733 gnd.n4248 gnd.n984 26.7676
R7734 gnd.n6441 gnd.n993 26.7676
R7735 gnd.n4254 gnd.n4253 26.7676
R7736 gnd.n6435 gnd.n1002 26.7676
R7737 gnd.n6429 gnd.n1012 26.7676
R7738 gnd.n4316 gnd.n1015 26.7676
R7739 gnd.n4324 gnd.n1025 26.7676
R7740 gnd.n6417 gnd.n1032 26.7676
R7741 gnd.n4331 gnd.n2114 26.7676
R7742 gnd.n6411 gnd.n1042 26.7676
R7743 gnd.n6405 gnd.n1052 26.7676
R7744 gnd.n4373 gnd.n1055 26.7676
R7745 gnd.n4346 gnd.n1065 26.7676
R7746 gnd.n6393 gnd.n1072 26.7676
R7747 gnd.n4351 gnd.n1075 26.7676
R7748 gnd.n6387 gnd.n1083 26.7676
R7749 gnd.n6381 gnd.n1092 26.7676
R7750 gnd.n6122 gnd.n1340 26.7676
R7751 gnd.n6116 gnd.n1352 26.7676
R7752 gnd.n5909 gnd.n1361 26.7676
R7753 gnd.n6110 gnd.n1364 26.7676
R7754 gnd.n5917 gnd.n1372 26.7676
R7755 gnd.n5936 gnd.n1381 26.7676
R7756 gnd.n6098 gnd.n1384 26.7676
R7757 gnd.n6092 gnd.n1395 26.7676
R7758 gnd.n5990 gnd.n5989 26.7676
R7759 gnd.n6086 gnd.n1404 26.7676
R7760 gnd.n5998 gnd.n1412 26.7676
R7761 gnd.n6004 gnd.n1421 26.7676
R7762 gnd.n6074 gnd.n1424 26.7676
R7763 gnd.n6068 gnd.n1435 26.7676
R7764 gnd.n6038 gnd.n6037 26.7676
R7765 gnd.n6062 gnd.n1444 26.7676
R7766 gnd.n6021 gnd.n1450 26.7676
R7767 gnd.n6049 gnd.n6048 26.7676
R7768 gnd.n1460 gnd.n375 26.7676
R7769 gnd.n7300 gnd.n369 26.7676
R7770 gnd.n7638 gnd.n87 26.7676
R7771 gnd.n7317 gnd.n362 26.7676
R7772 gnd.n7630 gnd.n105 26.7676
R7773 gnd.n7333 gnd.n114 26.7676
R7774 gnd.n7343 gnd.n123 26.7676
R7775 gnd.n4227 gnd.t46 26.4489
R7776 gnd.n7313 gnd.t6 26.4489
R7777 gnd.t60 gnd.n6466 25.8116
R7778 gnd.n7618 gnd.t21 25.8116
R7779 gnd.n2083 gnd.n2082 25.7944
R7780 gnd.n5381 gnd.n5380 25.7944
R7781 gnd.n2770 gnd.n2769 25.7944
R7782 gnd.n2312 gnd.n2311 25.7944
R7783 gnd.n2076 gnd.n2075 25.7944
R7784 gnd.n5794 gnd.n5793 25.7944
R7785 gnd.n5846 gnd.n5845 25.7944
R7786 gnd.n1501 gnd.n1500 25.7944
R7787 gnd.n312 gnd.n311 25.7944
R7788 gnd.n279 gnd.n278 25.7944
R7789 gnd.n7528 gnd.n7527 25.7944
R7790 gnd.n349 gnd.n348 25.7944
R7791 gnd.n3808 gnd.n3807 25.7944
R7792 gnd.n3830 gnd.n3829 25.7944
R7793 gnd.n3851 gnd.n3850 25.7944
R7794 gnd.n3869 gnd.n3868 25.7944
R7795 gnd.n1129 gnd.n1128 25.7944
R7796 gnd.n4425 gnd.n4424 25.7944
R7797 gnd.n4447 gnd.n4446 25.7944
R7798 gnd.n5371 gnd.n5370 25.7944
R7799 gnd.n4113 gnd.t90 25.1743
R7800 gnd.n4152 gnd.n2183 25.1743
R7801 gnd.n7612 gnd.n135 25.1743
R7802 gnd.n7594 gnd.t4 25.1743
R7803 gnd.n2991 gnd.n2711 24.8557
R7804 gnd.n3001 gnd.n2694 24.8557
R7805 gnd.n2697 gnd.n2685 24.8557
R7806 gnd.n3022 gnd.n2686 24.8557
R7807 gnd.n3032 gnd.n2666 24.8557
R7808 gnd.n3042 gnd.n3041 24.8557
R7809 gnd.n2652 gnd.n2650 24.8557
R7810 gnd.n3073 gnd.n3072 24.8557
R7811 gnd.n3088 gnd.n2635 24.8557
R7812 gnd.n3142 gnd.n2574 24.8557
R7813 gnd.n3098 gnd.n2575 24.8557
R7814 gnd.n3135 gnd.n2586 24.8557
R7815 gnd.n2624 gnd.n2623 24.8557
R7816 gnd.n3129 gnd.n3128 24.8557
R7817 gnd.n2610 gnd.n2597 24.8557
R7818 gnd.n3168 gnd.n3167 24.8557
R7819 gnd.n3178 gnd.n2490 24.8557
R7820 gnd.n3190 gnd.n2482 24.8557
R7821 gnd.n3189 gnd.n2470 24.8557
R7822 gnd.n3208 gnd.n3207 24.8557
R7823 gnd.n3218 gnd.n2463 24.8557
R7824 gnd.n3229 gnd.n2451 24.8557
R7825 gnd.n3253 gnd.n3252 24.8557
R7826 gnd.n3264 gnd.n2434 24.8557
R7827 gnd.n3263 gnd.n2436 24.8557
R7828 gnd.n3275 gnd.n2427 24.8557
R7829 gnd.n3293 gnd.n3292 24.8557
R7830 gnd.n2418 gnd.n2407 24.8557
R7831 gnd.n3314 gnd.n2395 24.8557
R7832 gnd.n3342 gnd.n3341 24.8557
R7833 gnd.n3353 gnd.n2380 24.8557
R7834 gnd.n3364 gnd.n2373 24.8557
R7835 gnd.n3363 gnd.n2361 24.8557
R7836 gnd.n3636 gnd.n3635 24.8557
R7837 gnd.n3658 gnd.n2346 24.8557
R7838 gnd.n3012 gnd.t30 23.2624
R7839 gnd.n2713 gnd.t203 22.6251
R7840 gnd.n4053 gnd.t145 22.6251
R7841 gnd.n4358 gnd.t163 22.6251
R7842 gnd.n5361 gnd.t141 22.6251
R7843 gnd.n7413 gnd.t156 22.6251
R7844 gnd.n6475 gnd.n934 22.4457
R7845 gnd.n4191 gnd.t50 21.9878
R7846 gnd.n358 gnd.t23 21.9878
R7847 gnd.t92 gnd.n2718 21.3504
R7848 gnd.n4215 gnd.t72 21.3504
R7849 gnd.n7298 gnd.t2 21.3504
R7850 gnd.t126 gnd.n2408 20.7131
R7851 gnd.t17 gnd.n1005 20.7131
R7852 gnd.t58 gnd.n1432 20.7131
R7853 gnd.n4391 gnd.n1100 20.3945
R7854 gnd.n1337 gnd.n1329 20.3945
R7855 gnd.n7564 gnd.n207 20.3945
R7856 gnd.t107 gnd.n2443 20.0758
R7857 gnd.t258 gnd.n1045 20.0758
R7858 gnd.t19 gnd.n1392 20.0758
R7859 gnd.n1951 gnd.n1950 19.9763
R7860 gnd.n1570 gnd.n1569 19.9763
R7861 gnd.n6262 gnd.n6261 19.9763
R7862 gnd.n5588 gnd.n5587 19.9763
R7863 gnd.n1193 gnd.t161 19.8005
R7864 gnd.n1193 gnd.t220 19.8005
R7865 gnd.n1192 gnd.t181 19.8005
R7866 gnd.n1192 gnd.t208 19.8005
R7867 gnd.n5578 gnd.t131 19.8005
R7868 gnd.n5578 gnd.t245 19.8005
R7869 gnd.n5577 gnd.t194 19.8005
R7870 gnd.n5577 gnd.t178 19.8005
R7871 gnd.n1189 gnd.n1188 19.5087
R7872 gnd.n1202 gnd.n1189 19.5087
R7873 gnd.n1200 gnd.n1191 19.5087
R7874 gnd.n5582 gnd.n5576 19.5087
R7875 gnd.n3179 gnd.t103 19.4385
R7876 gnd.n4674 gnd.n2070 19.3944
R7877 gnd.n2070 gnd.n2048 19.3944
R7878 gnd.n4699 gnd.n2048 19.3944
R7879 gnd.n4699 gnd.n2045 19.3944
R7880 gnd.n4706 gnd.n2045 19.3944
R7881 gnd.n4706 gnd.n2046 19.3944
R7882 gnd.n4702 gnd.n2046 19.3944
R7883 gnd.n4702 gnd.n1947 19.3944
R7884 gnd.n4736 gnd.n1947 19.3944
R7885 gnd.n4736 gnd.n1944 19.3944
R7886 gnd.n4741 gnd.n1944 19.3944
R7887 gnd.n4741 gnd.n1945 19.3944
R7888 gnd.n1945 gnd.n1936 19.3944
R7889 gnd.n4761 gnd.n1936 19.3944
R7890 gnd.n4761 gnd.n1933 19.3944
R7891 gnd.n4772 gnd.n1933 19.3944
R7892 gnd.n4772 gnd.n1934 19.3944
R7893 gnd.n4768 gnd.n1934 19.3944
R7894 gnd.n4768 gnd.n4767 19.3944
R7895 gnd.n4767 gnd.n1889 19.3944
R7896 gnd.n4847 gnd.n1889 19.3944
R7897 gnd.n4847 gnd.n1886 19.3944
R7898 gnd.n4870 gnd.n1886 19.3944
R7899 gnd.n4870 gnd.n1887 19.3944
R7900 gnd.n4866 gnd.n1887 19.3944
R7901 gnd.n4866 gnd.n4865 19.3944
R7902 gnd.n4865 gnd.n4864 19.3944
R7903 gnd.n4864 gnd.n4856 19.3944
R7904 gnd.n4860 gnd.n4856 19.3944
R7905 gnd.n4860 gnd.n4859 19.3944
R7906 gnd.n4859 gnd.n1839 19.3944
R7907 gnd.n1839 gnd.n1837 19.3944
R7908 gnd.n4949 gnd.n1837 19.3944
R7909 gnd.n4949 gnd.n1835 19.3944
R7910 gnd.n4953 gnd.n1835 19.3944
R7911 gnd.n4953 gnd.n1810 19.3944
R7912 gnd.n4999 gnd.n1810 19.3944
R7913 gnd.n4999 gnd.n1811 19.3944
R7914 gnd.n4995 gnd.n1811 19.3944
R7915 gnd.n4995 gnd.n1787 19.3944
R7916 gnd.n5058 gnd.n1787 19.3944
R7917 gnd.n5058 gnd.n1788 19.3944
R7918 gnd.n5054 gnd.n1788 19.3944
R7919 gnd.n5054 gnd.n5053 19.3944
R7920 gnd.n5053 gnd.n5052 19.3944
R7921 gnd.n5052 gnd.n5038 19.3944
R7922 gnd.n5048 gnd.n5038 19.3944
R7923 gnd.n5048 gnd.n5047 19.3944
R7924 gnd.n5047 gnd.n5046 19.3944
R7925 gnd.n5046 gnd.n1728 19.3944
R7926 gnd.n5166 gnd.n1728 19.3944
R7927 gnd.n5166 gnd.n1725 19.3944
R7928 gnd.n5171 gnd.n1725 19.3944
R7929 gnd.n5171 gnd.n1726 19.3944
R7930 gnd.n1726 gnd.n1699 19.3944
R7931 gnd.n5205 gnd.n1699 19.3944
R7932 gnd.n5205 gnd.n1696 19.3944
R7933 gnd.n5224 gnd.n1696 19.3944
R7934 gnd.n5224 gnd.n1697 19.3944
R7935 gnd.n5220 gnd.n1697 19.3944
R7936 gnd.n5220 gnd.n5219 19.3944
R7937 gnd.n5219 gnd.n5218 19.3944
R7938 gnd.n5218 gnd.n5213 19.3944
R7939 gnd.n5214 gnd.n5213 19.3944
R7940 gnd.n5214 gnd.n1643 19.3944
R7941 gnd.n5296 gnd.n1643 19.3944
R7942 gnd.n5296 gnd.n1640 19.3944
R7943 gnd.n5301 gnd.n1640 19.3944
R7944 gnd.n5301 gnd.n1641 19.3944
R7945 gnd.n1641 gnd.n1616 19.3944
R7946 gnd.n5338 gnd.n1616 19.3944
R7947 gnd.n5338 gnd.n1614 19.3944
R7948 gnd.n5342 gnd.n1614 19.3944
R7949 gnd.n5342 gnd.n1613 19.3944
R7950 gnd.n5349 gnd.n1613 19.3944
R7951 gnd.n5349 gnd.n1611 19.3944
R7952 gnd.n5353 gnd.n1611 19.3944
R7953 gnd.n5354 gnd.n5353 19.3944
R7954 gnd.n5357 gnd.n5354 19.3944
R7955 gnd.n5357 gnd.n1608 19.3944
R7956 gnd.n5539 gnd.n1608 19.3944
R7957 gnd.n5539 gnd.n1609 19.3944
R7958 gnd.n4658 gnd.n2072 19.3944
R7959 gnd.n4669 gnd.n2072 19.3944
R7960 gnd.n4670 gnd.n4669 19.3944
R7961 gnd.n4652 gnd.n4651 19.3944
R7962 gnd.n4651 gnd.n4417 19.3944
R7963 gnd.n4647 gnd.n4417 19.3944
R7964 gnd.n4647 gnd.n4646 19.3944
R7965 gnd.n4646 gnd.n4645 19.3944
R7966 gnd.n4645 gnd.n4422 19.3944
R7967 gnd.n4640 gnd.n4422 19.3944
R7968 gnd.n4640 gnd.n4639 19.3944
R7969 gnd.n4639 gnd.n4638 19.3944
R7970 gnd.n4638 gnd.n4541 19.3944
R7971 gnd.n4631 gnd.n4541 19.3944
R7972 gnd.n4631 gnd.n4630 19.3944
R7973 gnd.n4630 gnd.n4554 19.3944
R7974 gnd.n4623 gnd.n4554 19.3944
R7975 gnd.n4623 gnd.n4622 19.3944
R7976 gnd.n4622 gnd.n4564 19.3944
R7977 gnd.n4615 gnd.n4564 19.3944
R7978 gnd.n4615 gnd.n4614 19.3944
R7979 gnd.n4614 gnd.n4577 19.3944
R7980 gnd.n4607 gnd.n4577 19.3944
R7981 gnd.n4607 gnd.n4606 19.3944
R7982 gnd.n4606 gnd.n4587 19.3944
R7983 gnd.n4599 gnd.n4587 19.3944
R7984 gnd.n4599 gnd.n4598 19.3944
R7985 gnd.n5447 gnd.n5411 19.3944
R7986 gnd.n5460 gnd.n5411 19.3944
R7987 gnd.n5460 gnd.n5409 19.3944
R7988 gnd.n5466 gnd.n5409 19.3944
R7989 gnd.n5466 gnd.n5402 19.3944
R7990 gnd.n5479 gnd.n5402 19.3944
R7991 gnd.n5479 gnd.n5400 19.3944
R7992 gnd.n5485 gnd.n5400 19.3944
R7993 gnd.n5485 gnd.n5393 19.3944
R7994 gnd.n5498 gnd.n5393 19.3944
R7995 gnd.n5498 gnd.n5391 19.3944
R7996 gnd.n5504 gnd.n5391 19.3944
R7997 gnd.n5504 gnd.n5384 19.3944
R7998 gnd.n5518 gnd.n5384 19.3944
R7999 gnd.n5518 gnd.n5382 19.3944
R8000 gnd.n5524 gnd.n5382 19.3944
R8001 gnd.n2894 gnd.n2893 19.3944
R8002 gnd.n2893 gnd.n2892 19.3944
R8003 gnd.n2892 gnd.n2891 19.3944
R8004 gnd.n2891 gnd.n2889 19.3944
R8005 gnd.n2889 gnd.n2886 19.3944
R8006 gnd.n2886 gnd.n2885 19.3944
R8007 gnd.n2885 gnd.n2882 19.3944
R8008 gnd.n2882 gnd.n2881 19.3944
R8009 gnd.n2881 gnd.n2878 19.3944
R8010 gnd.n2878 gnd.n2877 19.3944
R8011 gnd.n2877 gnd.n2874 19.3944
R8012 gnd.n2874 gnd.n2873 19.3944
R8013 gnd.n2873 gnd.n2870 19.3944
R8014 gnd.n2870 gnd.n2869 19.3944
R8015 gnd.n2869 gnd.n2866 19.3944
R8016 gnd.n2866 gnd.n2865 19.3944
R8017 gnd.n2865 gnd.n2862 19.3944
R8018 gnd.n2862 gnd.n2861 19.3944
R8019 gnd.n2861 gnd.n2858 19.3944
R8020 gnd.n2858 gnd.n2857 19.3944
R8021 gnd.n2857 gnd.n2854 19.3944
R8022 gnd.n2854 gnd.n2853 19.3944
R8023 gnd.n2850 gnd.n2849 19.3944
R8024 gnd.n2849 gnd.n2805 19.3944
R8025 gnd.n2900 gnd.n2805 19.3944
R8026 gnd.n3666 gnd.n3665 19.3944
R8027 gnd.n3665 gnd.n3662 19.3944
R8028 gnd.n3662 gnd.n3661 19.3944
R8029 gnd.n3711 gnd.n3710 19.3944
R8030 gnd.n3710 gnd.n3709 19.3944
R8031 gnd.n3709 gnd.n3706 19.3944
R8032 gnd.n3706 gnd.n3705 19.3944
R8033 gnd.n3705 gnd.n3702 19.3944
R8034 gnd.n3702 gnd.n3701 19.3944
R8035 gnd.n3701 gnd.n3698 19.3944
R8036 gnd.n3698 gnd.n3697 19.3944
R8037 gnd.n3697 gnd.n3694 19.3944
R8038 gnd.n3694 gnd.n3693 19.3944
R8039 gnd.n3693 gnd.n3690 19.3944
R8040 gnd.n3690 gnd.n3689 19.3944
R8041 gnd.n3689 gnd.n3686 19.3944
R8042 gnd.n3686 gnd.n3685 19.3944
R8043 gnd.n3685 gnd.n3682 19.3944
R8044 gnd.n3682 gnd.n3681 19.3944
R8045 gnd.n3681 gnd.n3678 19.3944
R8046 gnd.n3678 gnd.n3677 19.3944
R8047 gnd.n3677 gnd.n3674 19.3944
R8048 gnd.n3674 gnd.n3673 19.3944
R8049 gnd.n3673 gnd.n3670 19.3944
R8050 gnd.n3670 gnd.n3669 19.3944
R8051 gnd.n2993 gnd.n2702 19.3944
R8052 gnd.n3003 gnd.n2702 19.3944
R8053 gnd.n3004 gnd.n3003 19.3944
R8054 gnd.n3004 gnd.n2683 19.3944
R8055 gnd.n3024 gnd.n2683 19.3944
R8056 gnd.n3024 gnd.n2675 19.3944
R8057 gnd.n3034 gnd.n2675 19.3944
R8058 gnd.n3035 gnd.n3034 19.3944
R8059 gnd.n3036 gnd.n3035 19.3944
R8060 gnd.n3036 gnd.n2658 19.3944
R8061 gnd.n3053 gnd.n2658 19.3944
R8062 gnd.n3056 gnd.n3053 19.3944
R8063 gnd.n3056 gnd.n3055 19.3944
R8064 gnd.n3055 gnd.n2631 19.3944
R8065 gnd.n3095 gnd.n2631 19.3944
R8066 gnd.n3095 gnd.n2628 19.3944
R8067 gnd.n3101 gnd.n2628 19.3944
R8068 gnd.n3102 gnd.n3101 19.3944
R8069 gnd.n3102 gnd.n2626 19.3944
R8070 gnd.n3108 gnd.n2626 19.3944
R8071 gnd.n3111 gnd.n3108 19.3944
R8072 gnd.n3113 gnd.n3111 19.3944
R8073 gnd.n3119 gnd.n3113 19.3944
R8074 gnd.n3119 gnd.n3118 19.3944
R8075 gnd.n3118 gnd.n2485 19.3944
R8076 gnd.n3185 gnd.n2485 19.3944
R8077 gnd.n3186 gnd.n3185 19.3944
R8078 gnd.n3186 gnd.n2478 19.3944
R8079 gnd.n3197 gnd.n2478 19.3944
R8080 gnd.n3198 gnd.n3197 19.3944
R8081 gnd.n3198 gnd.n2461 19.3944
R8082 gnd.n2461 gnd.n2459 19.3944
R8083 gnd.n3222 gnd.n2459 19.3944
R8084 gnd.n3223 gnd.n3222 19.3944
R8085 gnd.n3223 gnd.n2430 19.3944
R8086 gnd.n3270 gnd.n2430 19.3944
R8087 gnd.n3271 gnd.n3270 19.3944
R8088 gnd.n3271 gnd.n2423 19.3944
R8089 gnd.n3282 gnd.n2423 19.3944
R8090 gnd.n3283 gnd.n3282 19.3944
R8091 gnd.n3283 gnd.n2406 19.3944
R8092 gnd.n2406 gnd.n2404 19.3944
R8093 gnd.n3307 gnd.n2404 19.3944
R8094 gnd.n3308 gnd.n3307 19.3944
R8095 gnd.n3308 gnd.n2376 19.3944
R8096 gnd.n3359 gnd.n2376 19.3944
R8097 gnd.n3360 gnd.n3359 19.3944
R8098 gnd.n3360 gnd.n2369 19.3944
R8099 gnd.n3627 gnd.n2369 19.3944
R8100 gnd.n3628 gnd.n3627 19.3944
R8101 gnd.n3628 gnd.n2350 19.3944
R8102 gnd.n3653 gnd.n2350 19.3944
R8103 gnd.n3653 gnd.n2351 19.3944
R8104 gnd.n2984 gnd.n2983 19.3944
R8105 gnd.n2983 gnd.n2716 19.3944
R8106 gnd.n2739 gnd.n2716 19.3944
R8107 gnd.n2742 gnd.n2739 19.3944
R8108 gnd.n2742 gnd.n2735 19.3944
R8109 gnd.n2746 gnd.n2735 19.3944
R8110 gnd.n2749 gnd.n2746 19.3944
R8111 gnd.n2752 gnd.n2749 19.3944
R8112 gnd.n2752 gnd.n2733 19.3944
R8113 gnd.n2756 gnd.n2733 19.3944
R8114 gnd.n2759 gnd.n2756 19.3944
R8115 gnd.n2762 gnd.n2759 19.3944
R8116 gnd.n2762 gnd.n2731 19.3944
R8117 gnd.n2766 gnd.n2731 19.3944
R8118 gnd.n2989 gnd.n2988 19.3944
R8119 gnd.n2988 gnd.n2692 19.3944
R8120 gnd.n3014 gnd.n2692 19.3944
R8121 gnd.n3014 gnd.n2690 19.3944
R8122 gnd.n3020 gnd.n2690 19.3944
R8123 gnd.n3020 gnd.n3019 19.3944
R8124 gnd.n3019 gnd.n2664 19.3944
R8125 gnd.n3044 gnd.n2664 19.3944
R8126 gnd.n3044 gnd.n2662 19.3944
R8127 gnd.n3048 gnd.n2662 19.3944
R8128 gnd.n3048 gnd.n2642 19.3944
R8129 gnd.n3075 gnd.n2642 19.3944
R8130 gnd.n3075 gnd.n2640 19.3944
R8131 gnd.n3085 gnd.n2640 19.3944
R8132 gnd.n3085 gnd.n3084 19.3944
R8133 gnd.n3084 gnd.n3083 19.3944
R8134 gnd.n3083 gnd.n2589 19.3944
R8135 gnd.n3133 gnd.n2589 19.3944
R8136 gnd.n3133 gnd.n3132 19.3944
R8137 gnd.n3132 gnd.n3131 19.3944
R8138 gnd.n3131 gnd.n2593 19.3944
R8139 gnd.n2613 gnd.n2593 19.3944
R8140 gnd.n2613 gnd.n2495 19.3944
R8141 gnd.n3170 gnd.n2495 19.3944
R8142 gnd.n3170 gnd.n2493 19.3944
R8143 gnd.n3176 gnd.n2493 19.3944
R8144 gnd.n3176 gnd.n3175 19.3944
R8145 gnd.n3175 gnd.n2468 19.3944
R8146 gnd.n3210 gnd.n2468 19.3944
R8147 gnd.n3210 gnd.n2466 19.3944
R8148 gnd.n3216 gnd.n2466 19.3944
R8149 gnd.n3216 gnd.n3215 19.3944
R8150 gnd.n3215 gnd.n2441 19.3944
R8151 gnd.n3255 gnd.n2441 19.3944
R8152 gnd.n3255 gnd.n2439 19.3944
R8153 gnd.n3261 gnd.n2439 19.3944
R8154 gnd.n3261 gnd.n3260 19.3944
R8155 gnd.n3260 gnd.n2413 19.3944
R8156 gnd.n3295 gnd.n2413 19.3944
R8157 gnd.n3295 gnd.n2411 19.3944
R8158 gnd.n3301 gnd.n2411 19.3944
R8159 gnd.n3301 gnd.n3300 19.3944
R8160 gnd.n3300 gnd.n2386 19.3944
R8161 gnd.n3344 gnd.n2386 19.3944
R8162 gnd.n3344 gnd.n2384 19.3944
R8163 gnd.n3350 gnd.n2384 19.3944
R8164 gnd.n3350 gnd.n3349 19.3944
R8165 gnd.n3349 gnd.n2359 19.3944
R8166 gnd.n3638 gnd.n2359 19.3944
R8167 gnd.n3638 gnd.n2357 19.3944
R8168 gnd.n3646 gnd.n2357 19.3944
R8169 gnd.n3646 gnd.n3645 19.3944
R8170 gnd.n3645 gnd.n3644 19.3944
R8171 gnd.n3747 gnd.n3746 19.3944
R8172 gnd.n3746 gnd.n2298 19.3944
R8173 gnd.n3742 gnd.n2298 19.3944
R8174 gnd.n3742 gnd.n3739 19.3944
R8175 gnd.n3739 gnd.n3736 19.3944
R8176 gnd.n3736 gnd.n3735 19.3944
R8177 gnd.n3735 gnd.n3732 19.3944
R8178 gnd.n3732 gnd.n3731 19.3944
R8179 gnd.n3731 gnd.n3728 19.3944
R8180 gnd.n3728 gnd.n3727 19.3944
R8181 gnd.n3727 gnd.n3724 19.3944
R8182 gnd.n3724 gnd.n3723 19.3944
R8183 gnd.n3723 gnd.n3720 19.3944
R8184 gnd.n3720 gnd.n3719 19.3944
R8185 gnd.n2904 gnd.n2803 19.3944
R8186 gnd.n2904 gnd.n2794 19.3944
R8187 gnd.n2917 gnd.n2794 19.3944
R8188 gnd.n2917 gnd.n2792 19.3944
R8189 gnd.n2921 gnd.n2792 19.3944
R8190 gnd.n2921 gnd.n2782 19.3944
R8191 gnd.n2933 gnd.n2782 19.3944
R8192 gnd.n2933 gnd.n2780 19.3944
R8193 gnd.n2967 gnd.n2780 19.3944
R8194 gnd.n2967 gnd.n2966 19.3944
R8195 gnd.n2966 gnd.n2965 19.3944
R8196 gnd.n2965 gnd.n2964 19.3944
R8197 gnd.n2964 gnd.n2961 19.3944
R8198 gnd.n2961 gnd.n2960 19.3944
R8199 gnd.n2960 gnd.n2959 19.3944
R8200 gnd.n2959 gnd.n2957 19.3944
R8201 gnd.n2957 gnd.n2956 19.3944
R8202 gnd.n2956 gnd.n2953 19.3944
R8203 gnd.n2953 gnd.n2952 19.3944
R8204 gnd.n2952 gnd.n2951 19.3944
R8205 gnd.n2951 gnd.n2949 19.3944
R8206 gnd.n2949 gnd.n2648 19.3944
R8207 gnd.n3064 gnd.n2648 19.3944
R8208 gnd.n3064 gnd.n2646 19.3944
R8209 gnd.n3070 gnd.n2646 19.3944
R8210 gnd.n3070 gnd.n3069 19.3944
R8211 gnd.n3069 gnd.n2570 19.3944
R8212 gnd.n3144 gnd.n2570 19.3944
R8213 gnd.n3144 gnd.n2571 19.3944
R8214 gnd.n2618 gnd.n2617 19.3944
R8215 gnd.n2621 gnd.n2620 19.3944
R8216 gnd.n2608 gnd.n2607 19.3944
R8217 gnd.n3163 gnd.n2500 19.3944
R8218 gnd.n3163 gnd.n3162 19.3944
R8219 gnd.n3162 gnd.n3161 19.3944
R8220 gnd.n3161 gnd.n3159 19.3944
R8221 gnd.n3159 gnd.n3158 19.3944
R8222 gnd.n3158 gnd.n3156 19.3944
R8223 gnd.n3156 gnd.n3155 19.3944
R8224 gnd.n3155 gnd.n2449 19.3944
R8225 gnd.n3231 gnd.n2449 19.3944
R8226 gnd.n3231 gnd.n2447 19.3944
R8227 gnd.n3250 gnd.n2447 19.3944
R8228 gnd.n3250 gnd.n3249 19.3944
R8229 gnd.n3249 gnd.n3248 19.3944
R8230 gnd.n3248 gnd.n3246 19.3944
R8231 gnd.n3246 gnd.n3245 19.3944
R8232 gnd.n3245 gnd.n3243 19.3944
R8233 gnd.n3243 gnd.n3242 19.3944
R8234 gnd.n3242 gnd.n2393 19.3944
R8235 gnd.n3316 gnd.n2393 19.3944
R8236 gnd.n3316 gnd.n2391 19.3944
R8237 gnd.n3339 gnd.n2391 19.3944
R8238 gnd.n3339 gnd.n3338 19.3944
R8239 gnd.n3338 gnd.n3337 19.3944
R8240 gnd.n3337 gnd.n3334 19.3944
R8241 gnd.n3334 gnd.n3333 19.3944
R8242 gnd.n3333 gnd.n3331 19.3944
R8243 gnd.n3331 gnd.n3330 19.3944
R8244 gnd.n3330 gnd.n3328 19.3944
R8245 gnd.n3328 gnd.n2345 19.3944
R8246 gnd.n2909 gnd.n2799 19.3944
R8247 gnd.n2909 gnd.n2797 19.3944
R8248 gnd.n2913 gnd.n2797 19.3944
R8249 gnd.n2913 gnd.n2788 19.3944
R8250 gnd.n2925 gnd.n2788 19.3944
R8251 gnd.n2925 gnd.n2786 19.3944
R8252 gnd.n2929 gnd.n2786 19.3944
R8253 gnd.n2929 gnd.n2775 19.3944
R8254 gnd.n2971 gnd.n2775 19.3944
R8255 gnd.n2971 gnd.n2729 19.3944
R8256 gnd.n2977 gnd.n2729 19.3944
R8257 gnd.n2977 gnd.n2976 19.3944
R8258 gnd.n2976 gnd.n2707 19.3944
R8259 gnd.n2998 gnd.n2707 19.3944
R8260 gnd.n2998 gnd.n2700 19.3944
R8261 gnd.n3009 gnd.n2700 19.3944
R8262 gnd.n3009 gnd.n3008 19.3944
R8263 gnd.n3008 gnd.n2681 19.3944
R8264 gnd.n3029 gnd.n2681 19.3944
R8265 gnd.n3029 gnd.n2671 19.3944
R8266 gnd.n3039 gnd.n2671 19.3944
R8267 gnd.n3039 gnd.n2654 19.3944
R8268 gnd.n3060 gnd.n2654 19.3944
R8269 gnd.n3060 gnd.n3059 19.3944
R8270 gnd.n3059 gnd.n2633 19.3944
R8271 gnd.n3090 gnd.n2633 19.3944
R8272 gnd.n3090 gnd.n2578 19.3944
R8273 gnd.n3140 gnd.n2578 19.3944
R8274 gnd.n3140 gnd.n3139 19.3944
R8275 gnd.n3139 gnd.n3138 19.3944
R8276 gnd.n3138 gnd.n2582 19.3944
R8277 gnd.n2600 gnd.n2582 19.3944
R8278 gnd.n3126 gnd.n2600 19.3944
R8279 gnd.n3126 gnd.n3125 19.3944
R8280 gnd.n3125 gnd.n3124 19.3944
R8281 gnd.n3124 gnd.n2604 19.3944
R8282 gnd.n2604 gnd.n2487 19.3944
R8283 gnd.n3181 gnd.n2487 19.3944
R8284 gnd.n3181 gnd.n2480 19.3944
R8285 gnd.n3192 gnd.n2480 19.3944
R8286 gnd.n3192 gnd.n2476 19.3944
R8287 gnd.n3205 gnd.n2476 19.3944
R8288 gnd.n3205 gnd.n3204 19.3944
R8289 gnd.n3204 gnd.n2455 19.3944
R8290 gnd.n3227 gnd.n2455 19.3944
R8291 gnd.n3227 gnd.n3226 19.3944
R8292 gnd.n3226 gnd.n2432 19.3944
R8293 gnd.n3266 gnd.n2432 19.3944
R8294 gnd.n3266 gnd.n2425 19.3944
R8295 gnd.n3277 gnd.n2425 19.3944
R8296 gnd.n3277 gnd.n2421 19.3944
R8297 gnd.n3290 gnd.n2421 19.3944
R8298 gnd.n3290 gnd.n3289 19.3944
R8299 gnd.n3289 gnd.n2400 19.3944
R8300 gnd.n3312 gnd.n2400 19.3944
R8301 gnd.n3312 gnd.n3311 19.3944
R8302 gnd.n3311 gnd.n2378 19.3944
R8303 gnd.n3355 gnd.n2378 19.3944
R8304 gnd.n3355 gnd.n2371 19.3944
R8305 gnd.n3366 gnd.n2371 19.3944
R8306 gnd.n3366 gnd.n2367 19.3944
R8307 gnd.n3633 gnd.n2367 19.3944
R8308 gnd.n3633 gnd.n3632 19.3944
R8309 gnd.n3632 gnd.n2348 19.3944
R8310 gnd.n3656 gnd.n2348 19.3944
R8311 gnd.n4635 gnd.n4544 19.3944
R8312 gnd.n4635 gnd.n4634 19.3944
R8313 gnd.n4634 gnd.n4548 19.3944
R8314 gnd.n4627 gnd.n4548 19.3944
R8315 gnd.n4627 gnd.n4626 19.3944
R8316 gnd.n4626 gnd.n4560 19.3944
R8317 gnd.n4619 gnd.n4560 19.3944
R8318 gnd.n4619 gnd.n4618 19.3944
R8319 gnd.n4618 gnd.n4571 19.3944
R8320 gnd.n4611 gnd.n4571 19.3944
R8321 gnd.n4611 gnd.n4610 19.3944
R8322 gnd.n4610 gnd.n4583 19.3944
R8323 gnd.n4603 gnd.n4583 19.3944
R8324 gnd.n4603 gnd.n4602 19.3944
R8325 gnd.n4602 gnd.n2079 19.3944
R8326 gnd.n4661 gnd.n2079 19.3944
R8327 gnd.n7064 gnd.n516 19.3944
R8328 gnd.n7070 gnd.n516 19.3944
R8329 gnd.n7070 gnd.n514 19.3944
R8330 gnd.n7074 gnd.n514 19.3944
R8331 gnd.n7074 gnd.n510 19.3944
R8332 gnd.n7080 gnd.n510 19.3944
R8333 gnd.n7080 gnd.n508 19.3944
R8334 gnd.n7084 gnd.n508 19.3944
R8335 gnd.n7084 gnd.n504 19.3944
R8336 gnd.n7090 gnd.n504 19.3944
R8337 gnd.n7090 gnd.n502 19.3944
R8338 gnd.n7094 gnd.n502 19.3944
R8339 gnd.n7094 gnd.n498 19.3944
R8340 gnd.n7100 gnd.n498 19.3944
R8341 gnd.n7100 gnd.n496 19.3944
R8342 gnd.n7104 gnd.n496 19.3944
R8343 gnd.n7104 gnd.n492 19.3944
R8344 gnd.n7110 gnd.n492 19.3944
R8345 gnd.n7110 gnd.n490 19.3944
R8346 gnd.n7114 gnd.n490 19.3944
R8347 gnd.n7114 gnd.n486 19.3944
R8348 gnd.n7120 gnd.n486 19.3944
R8349 gnd.n7120 gnd.n484 19.3944
R8350 gnd.n7124 gnd.n484 19.3944
R8351 gnd.n7124 gnd.n480 19.3944
R8352 gnd.n7130 gnd.n480 19.3944
R8353 gnd.n7130 gnd.n478 19.3944
R8354 gnd.n7134 gnd.n478 19.3944
R8355 gnd.n7134 gnd.n474 19.3944
R8356 gnd.n7140 gnd.n474 19.3944
R8357 gnd.n7140 gnd.n472 19.3944
R8358 gnd.n7144 gnd.n472 19.3944
R8359 gnd.n7144 gnd.n468 19.3944
R8360 gnd.n7150 gnd.n468 19.3944
R8361 gnd.n7150 gnd.n466 19.3944
R8362 gnd.n7154 gnd.n466 19.3944
R8363 gnd.n7154 gnd.n462 19.3944
R8364 gnd.n7160 gnd.n462 19.3944
R8365 gnd.n7160 gnd.n460 19.3944
R8366 gnd.n7164 gnd.n460 19.3944
R8367 gnd.n7164 gnd.n456 19.3944
R8368 gnd.n7170 gnd.n456 19.3944
R8369 gnd.n7170 gnd.n454 19.3944
R8370 gnd.n7174 gnd.n454 19.3944
R8371 gnd.n7174 gnd.n450 19.3944
R8372 gnd.n7180 gnd.n450 19.3944
R8373 gnd.n7180 gnd.n448 19.3944
R8374 gnd.n7184 gnd.n448 19.3944
R8375 gnd.n7184 gnd.n444 19.3944
R8376 gnd.n7190 gnd.n444 19.3944
R8377 gnd.n7190 gnd.n442 19.3944
R8378 gnd.n7194 gnd.n442 19.3944
R8379 gnd.n7194 gnd.n438 19.3944
R8380 gnd.n7200 gnd.n438 19.3944
R8381 gnd.n7200 gnd.n436 19.3944
R8382 gnd.n7204 gnd.n436 19.3944
R8383 gnd.n7204 gnd.n432 19.3944
R8384 gnd.n7210 gnd.n432 19.3944
R8385 gnd.n7210 gnd.n430 19.3944
R8386 gnd.n7214 gnd.n430 19.3944
R8387 gnd.n7214 gnd.n426 19.3944
R8388 gnd.n7220 gnd.n426 19.3944
R8389 gnd.n7220 gnd.n424 19.3944
R8390 gnd.n7224 gnd.n424 19.3944
R8391 gnd.n7224 gnd.n420 19.3944
R8392 gnd.n7230 gnd.n420 19.3944
R8393 gnd.n7230 gnd.n418 19.3944
R8394 gnd.n7234 gnd.n418 19.3944
R8395 gnd.n7234 gnd.n414 19.3944
R8396 gnd.n7240 gnd.n414 19.3944
R8397 gnd.n7240 gnd.n412 19.3944
R8398 gnd.n7244 gnd.n412 19.3944
R8399 gnd.n7244 gnd.n408 19.3944
R8400 gnd.n7250 gnd.n408 19.3944
R8401 gnd.n7250 gnd.n406 19.3944
R8402 gnd.n7254 gnd.n406 19.3944
R8403 gnd.n7254 gnd.n402 19.3944
R8404 gnd.n7260 gnd.n402 19.3944
R8405 gnd.n7260 gnd.n400 19.3944
R8406 gnd.n7264 gnd.n400 19.3944
R8407 gnd.n7264 gnd.n396 19.3944
R8408 gnd.n7271 gnd.n396 19.3944
R8409 gnd.n7271 gnd.n394 19.3944
R8410 gnd.n7276 gnd.n394 19.3944
R8411 gnd.n6643 gnd.n767 19.3944
R8412 gnd.n6649 gnd.n767 19.3944
R8413 gnd.n6649 gnd.n765 19.3944
R8414 gnd.n6653 gnd.n765 19.3944
R8415 gnd.n6653 gnd.n761 19.3944
R8416 gnd.n6659 gnd.n761 19.3944
R8417 gnd.n6659 gnd.n759 19.3944
R8418 gnd.n6663 gnd.n759 19.3944
R8419 gnd.n6663 gnd.n755 19.3944
R8420 gnd.n6669 gnd.n755 19.3944
R8421 gnd.n6669 gnd.n753 19.3944
R8422 gnd.n6673 gnd.n753 19.3944
R8423 gnd.n6673 gnd.n749 19.3944
R8424 gnd.n6679 gnd.n749 19.3944
R8425 gnd.n6679 gnd.n747 19.3944
R8426 gnd.n6683 gnd.n747 19.3944
R8427 gnd.n6683 gnd.n743 19.3944
R8428 gnd.n6689 gnd.n743 19.3944
R8429 gnd.n6689 gnd.n741 19.3944
R8430 gnd.n6693 gnd.n741 19.3944
R8431 gnd.n6693 gnd.n737 19.3944
R8432 gnd.n6699 gnd.n737 19.3944
R8433 gnd.n6699 gnd.n735 19.3944
R8434 gnd.n6703 gnd.n735 19.3944
R8435 gnd.n6703 gnd.n731 19.3944
R8436 gnd.n6709 gnd.n731 19.3944
R8437 gnd.n6709 gnd.n729 19.3944
R8438 gnd.n6713 gnd.n729 19.3944
R8439 gnd.n6713 gnd.n725 19.3944
R8440 gnd.n6719 gnd.n725 19.3944
R8441 gnd.n6719 gnd.n723 19.3944
R8442 gnd.n6723 gnd.n723 19.3944
R8443 gnd.n6723 gnd.n719 19.3944
R8444 gnd.n6729 gnd.n719 19.3944
R8445 gnd.n6729 gnd.n717 19.3944
R8446 gnd.n6733 gnd.n717 19.3944
R8447 gnd.n6733 gnd.n713 19.3944
R8448 gnd.n6739 gnd.n713 19.3944
R8449 gnd.n6739 gnd.n711 19.3944
R8450 gnd.n6743 gnd.n711 19.3944
R8451 gnd.n6743 gnd.n707 19.3944
R8452 gnd.n6749 gnd.n707 19.3944
R8453 gnd.n6749 gnd.n705 19.3944
R8454 gnd.n6753 gnd.n705 19.3944
R8455 gnd.n6753 gnd.n701 19.3944
R8456 gnd.n6759 gnd.n701 19.3944
R8457 gnd.n6759 gnd.n699 19.3944
R8458 gnd.n6763 gnd.n699 19.3944
R8459 gnd.n6763 gnd.n695 19.3944
R8460 gnd.n6769 gnd.n695 19.3944
R8461 gnd.n6769 gnd.n693 19.3944
R8462 gnd.n6773 gnd.n693 19.3944
R8463 gnd.n6773 gnd.n689 19.3944
R8464 gnd.n6779 gnd.n689 19.3944
R8465 gnd.n6779 gnd.n687 19.3944
R8466 gnd.n6783 gnd.n687 19.3944
R8467 gnd.n6783 gnd.n683 19.3944
R8468 gnd.n6789 gnd.n683 19.3944
R8469 gnd.n6789 gnd.n681 19.3944
R8470 gnd.n6793 gnd.n681 19.3944
R8471 gnd.n6793 gnd.n677 19.3944
R8472 gnd.n6799 gnd.n677 19.3944
R8473 gnd.n6799 gnd.n675 19.3944
R8474 gnd.n6803 gnd.n675 19.3944
R8475 gnd.n6803 gnd.n671 19.3944
R8476 gnd.n6809 gnd.n671 19.3944
R8477 gnd.n6809 gnd.n669 19.3944
R8478 gnd.n6813 gnd.n669 19.3944
R8479 gnd.n6813 gnd.n665 19.3944
R8480 gnd.n6819 gnd.n665 19.3944
R8481 gnd.n6819 gnd.n663 19.3944
R8482 gnd.n6823 gnd.n663 19.3944
R8483 gnd.n6823 gnd.n659 19.3944
R8484 gnd.n6829 gnd.n659 19.3944
R8485 gnd.n6829 gnd.n657 19.3944
R8486 gnd.n6833 gnd.n657 19.3944
R8487 gnd.n6833 gnd.n653 19.3944
R8488 gnd.n6839 gnd.n653 19.3944
R8489 gnd.n6839 gnd.n651 19.3944
R8490 gnd.n6843 gnd.n651 19.3944
R8491 gnd.n6843 gnd.n647 19.3944
R8492 gnd.n6849 gnd.n647 19.3944
R8493 gnd.n6849 gnd.n645 19.3944
R8494 gnd.n6853 gnd.n645 19.3944
R8495 gnd.n6853 gnd.n641 19.3944
R8496 gnd.n6859 gnd.n641 19.3944
R8497 gnd.n6859 gnd.n639 19.3944
R8498 gnd.n6863 gnd.n639 19.3944
R8499 gnd.n6863 gnd.n635 19.3944
R8500 gnd.n6869 gnd.n635 19.3944
R8501 gnd.n6869 gnd.n633 19.3944
R8502 gnd.n6873 gnd.n633 19.3944
R8503 gnd.n6873 gnd.n629 19.3944
R8504 gnd.n6879 gnd.n629 19.3944
R8505 gnd.n6879 gnd.n627 19.3944
R8506 gnd.n6883 gnd.n627 19.3944
R8507 gnd.n6883 gnd.n623 19.3944
R8508 gnd.n6889 gnd.n623 19.3944
R8509 gnd.n6889 gnd.n621 19.3944
R8510 gnd.n6893 gnd.n621 19.3944
R8511 gnd.n6893 gnd.n617 19.3944
R8512 gnd.n6899 gnd.n617 19.3944
R8513 gnd.n6899 gnd.n615 19.3944
R8514 gnd.n6903 gnd.n615 19.3944
R8515 gnd.n6903 gnd.n611 19.3944
R8516 gnd.n6909 gnd.n611 19.3944
R8517 gnd.n6909 gnd.n609 19.3944
R8518 gnd.n6913 gnd.n609 19.3944
R8519 gnd.n6913 gnd.n605 19.3944
R8520 gnd.n6919 gnd.n605 19.3944
R8521 gnd.n6919 gnd.n603 19.3944
R8522 gnd.n6923 gnd.n603 19.3944
R8523 gnd.n6923 gnd.n599 19.3944
R8524 gnd.n6929 gnd.n599 19.3944
R8525 gnd.n6929 gnd.n597 19.3944
R8526 gnd.n6933 gnd.n597 19.3944
R8527 gnd.n6933 gnd.n593 19.3944
R8528 gnd.n6939 gnd.n593 19.3944
R8529 gnd.n6939 gnd.n591 19.3944
R8530 gnd.n6943 gnd.n591 19.3944
R8531 gnd.n6943 gnd.n587 19.3944
R8532 gnd.n6949 gnd.n587 19.3944
R8533 gnd.n6949 gnd.n585 19.3944
R8534 gnd.n6953 gnd.n585 19.3944
R8535 gnd.n6953 gnd.n581 19.3944
R8536 gnd.n6959 gnd.n581 19.3944
R8537 gnd.n6959 gnd.n579 19.3944
R8538 gnd.n6963 gnd.n579 19.3944
R8539 gnd.n6963 gnd.n575 19.3944
R8540 gnd.n6969 gnd.n575 19.3944
R8541 gnd.n6969 gnd.n573 19.3944
R8542 gnd.n6973 gnd.n573 19.3944
R8543 gnd.n6973 gnd.n569 19.3944
R8544 gnd.n6979 gnd.n569 19.3944
R8545 gnd.n6979 gnd.n567 19.3944
R8546 gnd.n6983 gnd.n567 19.3944
R8547 gnd.n6983 gnd.n563 19.3944
R8548 gnd.n6989 gnd.n563 19.3944
R8549 gnd.n6989 gnd.n561 19.3944
R8550 gnd.n6993 gnd.n561 19.3944
R8551 gnd.n6993 gnd.n557 19.3944
R8552 gnd.n6999 gnd.n557 19.3944
R8553 gnd.n6999 gnd.n555 19.3944
R8554 gnd.n7003 gnd.n555 19.3944
R8555 gnd.n7003 gnd.n551 19.3944
R8556 gnd.n7009 gnd.n551 19.3944
R8557 gnd.n7009 gnd.n549 19.3944
R8558 gnd.n7013 gnd.n549 19.3944
R8559 gnd.n7013 gnd.n545 19.3944
R8560 gnd.n7019 gnd.n545 19.3944
R8561 gnd.n7019 gnd.n543 19.3944
R8562 gnd.n7023 gnd.n543 19.3944
R8563 gnd.n7023 gnd.n539 19.3944
R8564 gnd.n7029 gnd.n539 19.3944
R8565 gnd.n7029 gnd.n537 19.3944
R8566 gnd.n7033 gnd.n537 19.3944
R8567 gnd.n7033 gnd.n533 19.3944
R8568 gnd.n7039 gnd.n533 19.3944
R8569 gnd.n7039 gnd.n531 19.3944
R8570 gnd.n7043 gnd.n531 19.3944
R8571 gnd.n7043 gnd.n527 19.3944
R8572 gnd.n7049 gnd.n527 19.3944
R8573 gnd.n7049 gnd.n525 19.3944
R8574 gnd.n7054 gnd.n525 19.3944
R8575 gnd.n7054 gnd.n521 19.3944
R8576 gnd.n7060 gnd.n521 19.3944
R8577 gnd.n7061 gnd.n7060 19.3944
R8578 gnd.n5753 gnd.n5750 19.3944
R8579 gnd.n5753 gnd.n5749 19.3944
R8580 gnd.n5759 gnd.n5749 19.3944
R8581 gnd.n5759 gnd.n5747 19.3944
R8582 gnd.n5763 gnd.n5747 19.3944
R8583 gnd.n5763 gnd.n5745 19.3944
R8584 gnd.n5769 gnd.n5745 19.3944
R8585 gnd.n5769 gnd.n5743 19.3944
R8586 gnd.n5773 gnd.n5743 19.3944
R8587 gnd.n5773 gnd.n5741 19.3944
R8588 gnd.n5779 gnd.n5741 19.3944
R8589 gnd.n5779 gnd.n5739 19.3944
R8590 gnd.n5783 gnd.n5739 19.3944
R8591 gnd.n5783 gnd.n5737 19.3944
R8592 gnd.n5789 gnd.n5737 19.3944
R8593 gnd.n5789 gnd.n5735 19.3944
R8594 gnd.n5796 gnd.n5735 19.3944
R8595 gnd.n5802 gnd.n5733 19.3944
R8596 gnd.n5802 gnd.n5731 19.3944
R8597 gnd.n5806 gnd.n5731 19.3944
R8598 gnd.n5806 gnd.n5729 19.3944
R8599 gnd.n5812 gnd.n5729 19.3944
R8600 gnd.n5812 gnd.n5727 19.3944
R8601 gnd.n5817 gnd.n5727 19.3944
R8602 gnd.n5825 gnd.n1531 19.3944
R8603 gnd.n5825 gnd.n1529 19.3944
R8604 gnd.n5829 gnd.n1529 19.3944
R8605 gnd.n5829 gnd.n1527 19.3944
R8606 gnd.n5835 gnd.n1527 19.3944
R8607 gnd.n5835 gnd.n1525 19.3944
R8608 gnd.n5839 gnd.n1525 19.3944
R8609 gnd.n5839 gnd.n1523 19.3944
R8610 gnd.n5851 gnd.n1521 19.3944
R8611 gnd.n5851 gnd.n1519 19.3944
R8612 gnd.n5857 gnd.n1519 19.3944
R8613 gnd.n5857 gnd.n1517 19.3944
R8614 gnd.n5861 gnd.n1517 19.3944
R8615 gnd.n5861 gnd.n1515 19.3944
R8616 gnd.n5867 gnd.n1515 19.3944
R8617 gnd.n5867 gnd.n1513 19.3944
R8618 gnd.n5871 gnd.n1513 19.3944
R8619 gnd.n5871 gnd.n1511 19.3944
R8620 gnd.n5877 gnd.n1511 19.3944
R8621 gnd.n5877 gnd.n1509 19.3944
R8622 gnd.n5881 gnd.n1509 19.3944
R8623 gnd.n5881 gnd.n1507 19.3944
R8624 gnd.n5887 gnd.n1507 19.3944
R8625 gnd.n5887 gnd.n1505 19.3944
R8626 gnd.n5892 gnd.n1505 19.3944
R8627 gnd.n5892 gnd.n1503 19.3944
R8628 gnd.n5905 gnd.n1496 19.3944
R8629 gnd.n5906 gnd.n5905 19.3944
R8630 gnd.n5907 gnd.n5906 19.3944
R8631 gnd.n5907 gnd.n1491 19.3944
R8632 gnd.n5919 gnd.n1491 19.3944
R8633 gnd.n5920 gnd.n5919 19.3944
R8634 gnd.n5921 gnd.n5920 19.3944
R8635 gnd.n5922 gnd.n5921 19.3944
R8636 gnd.n5926 gnd.n5922 19.3944
R8637 gnd.n5926 gnd.n5925 19.3944
R8638 gnd.n5925 gnd.n5924 19.3944
R8639 gnd.n5924 gnd.n1476 19.3944
R8640 gnd.n6000 gnd.n1476 19.3944
R8641 gnd.n6001 gnd.n6000 19.3944
R8642 gnd.n6002 gnd.n6001 19.3944
R8643 gnd.n6002 gnd.n1470 19.3944
R8644 gnd.n6014 gnd.n1470 19.3944
R8645 gnd.n6015 gnd.n6014 19.3944
R8646 gnd.n6016 gnd.n6015 19.3944
R8647 gnd.n6017 gnd.n6016 19.3944
R8648 gnd.n6019 gnd.n6017 19.3944
R8649 gnd.n6019 gnd.n1455 19.3944
R8650 gnd.n6051 gnd.n1455 19.3944
R8651 gnd.n6051 gnd.n1456 19.3944
R8652 gnd.n1456 gnd.n371 19.3944
R8653 gnd.n7309 gnd.n371 19.3944
R8654 gnd.n7311 gnd.n7309 19.3944
R8655 gnd.n7311 gnd.n7310 19.3944
R8656 gnd.n7310 gnd.n364 19.3944
R8657 gnd.n7322 gnd.n364 19.3944
R8658 gnd.n7322 gnd.n359 19.3944
R8659 gnd.n7335 gnd.n359 19.3944
R8660 gnd.n7336 gnd.n7335 19.3944
R8661 gnd.n7341 gnd.n7336 19.3944
R8662 gnd.n7341 gnd.n7340 19.3944
R8663 gnd.n7340 gnd.n7339 19.3944
R8664 gnd.n7339 gnd.n352 19.3944
R8665 gnd.n7387 gnd.n352 19.3944
R8666 gnd.n7388 gnd.n7387 19.3944
R8667 gnd.n7390 gnd.n7388 19.3944
R8668 gnd.n7391 gnd.n7390 19.3944
R8669 gnd.n7394 gnd.n7391 19.3944
R8670 gnd.n7395 gnd.n7394 19.3944
R8671 gnd.n7397 gnd.n7395 19.3944
R8672 gnd.n7398 gnd.n7397 19.3944
R8673 gnd.n7401 gnd.n7398 19.3944
R8674 gnd.n7402 gnd.n7401 19.3944
R8675 gnd.n7404 gnd.n7402 19.3944
R8676 gnd.n7405 gnd.n7404 19.3944
R8677 gnd.n7408 gnd.n7405 19.3944
R8678 gnd.n7409 gnd.n7408 19.3944
R8679 gnd.n7411 gnd.n7409 19.3944
R8680 gnd.n7411 gnd.n7410 19.3944
R8681 gnd.n5902 gnd.n1355 19.3944
R8682 gnd.n6114 gnd.n1355 19.3944
R8683 gnd.n6114 gnd.n6113 19.3944
R8684 gnd.n6113 gnd.n6112 19.3944
R8685 gnd.n6112 gnd.n1359 19.3944
R8686 gnd.n6102 gnd.n1359 19.3944
R8687 gnd.n6102 gnd.n6101 19.3944
R8688 gnd.n6101 gnd.n6100 19.3944
R8689 gnd.n6100 gnd.n1379 19.3944
R8690 gnd.n6090 gnd.n1379 19.3944
R8691 gnd.n6090 gnd.n6089 19.3944
R8692 gnd.n6089 gnd.n6088 19.3944
R8693 gnd.n6088 gnd.n1400 19.3944
R8694 gnd.n6078 gnd.n1400 19.3944
R8695 gnd.n6078 gnd.n6077 19.3944
R8696 gnd.n6077 gnd.n6076 19.3944
R8697 gnd.n6076 gnd.n1419 19.3944
R8698 gnd.n6066 gnd.n1419 19.3944
R8699 gnd.n6066 gnd.n6065 19.3944
R8700 gnd.n6065 gnd.n6064 19.3944
R8701 gnd.n6064 gnd.n1440 19.3944
R8702 gnd.n6054 gnd.n1440 19.3944
R8703 gnd.n6054 gnd.n6053 19.3944
R8704 gnd.n6053 gnd.n373 19.3944
R8705 gnd.n7306 gnd.n373 19.3944
R8706 gnd.n7306 gnd.n366 19.3944
R8707 gnd.n7315 gnd.n366 19.3944
R8708 gnd.n7316 gnd.n7315 19.3944
R8709 gnd.n7319 gnd.n7316 19.3944
R8710 gnd.n7319 gnd.n108 19.3944
R8711 gnd.n7628 gnd.n108 19.3944
R8712 gnd.n7628 gnd.n7627 19.3944
R8713 gnd.n7627 gnd.n7626 19.3944
R8714 gnd.n7626 gnd.n112 19.3944
R8715 gnd.n7616 gnd.n112 19.3944
R8716 gnd.n7616 gnd.n7615 19.3944
R8717 gnd.n7615 gnd.n7614 19.3944
R8718 gnd.n7614 gnd.n130 19.3944
R8719 gnd.n7604 gnd.n130 19.3944
R8720 gnd.n7604 gnd.n7603 19.3944
R8721 gnd.n7603 gnd.n7602 19.3944
R8722 gnd.n7602 gnd.n150 19.3944
R8723 gnd.n7592 gnd.n150 19.3944
R8724 gnd.n7592 gnd.n7591 19.3944
R8725 gnd.n7591 gnd.n7590 19.3944
R8726 gnd.n7590 gnd.n168 19.3944
R8727 gnd.n7580 gnd.n168 19.3944
R8728 gnd.n7580 gnd.n7579 19.3944
R8729 gnd.n7579 gnd.n7578 19.3944
R8730 gnd.n7578 gnd.n188 19.3944
R8731 gnd.n7568 gnd.n188 19.3944
R8732 gnd.n7568 gnd.n7567 19.3944
R8733 gnd.n7567 gnd.n7566 19.3944
R8734 gnd.n7488 gnd.n277 19.3944
R8735 gnd.n7488 gnd.n281 19.3944
R8736 gnd.n284 gnd.n281 19.3944
R8737 gnd.n7481 gnd.n284 19.3944
R8738 gnd.n7481 gnd.n7480 19.3944
R8739 gnd.n7480 gnd.n7479 19.3944
R8740 gnd.n7479 gnd.n290 19.3944
R8741 gnd.n7474 gnd.n290 19.3944
R8742 gnd.n7474 gnd.n7473 19.3944
R8743 gnd.n7473 gnd.n7472 19.3944
R8744 gnd.n7472 gnd.n297 19.3944
R8745 gnd.n7467 gnd.n297 19.3944
R8746 gnd.n7467 gnd.n7466 19.3944
R8747 gnd.n7466 gnd.n7465 19.3944
R8748 gnd.n7465 gnd.n304 19.3944
R8749 gnd.n7460 gnd.n304 19.3944
R8750 gnd.n7460 gnd.n7459 19.3944
R8751 gnd.n7459 gnd.n7458 19.3944
R8752 gnd.n7526 gnd.n244 19.3944
R8753 gnd.n7521 gnd.n244 19.3944
R8754 gnd.n7521 gnd.n7520 19.3944
R8755 gnd.n7520 gnd.n7519 19.3944
R8756 gnd.n7519 gnd.n251 19.3944
R8757 gnd.n7514 gnd.n251 19.3944
R8758 gnd.n7514 gnd.n7513 19.3944
R8759 gnd.n7513 gnd.n7512 19.3944
R8760 gnd.n7512 gnd.n258 19.3944
R8761 gnd.n7507 gnd.n258 19.3944
R8762 gnd.n7507 gnd.n7506 19.3944
R8763 gnd.n7506 gnd.n7505 19.3944
R8764 gnd.n7505 gnd.n265 19.3944
R8765 gnd.n7500 gnd.n265 19.3944
R8766 gnd.n7500 gnd.n7499 19.3944
R8767 gnd.n7499 gnd.n7498 19.3944
R8768 gnd.n7498 gnd.n272 19.3944
R8769 gnd.n7493 gnd.n272 19.3944
R8770 gnd.n7559 gnd.n7558 19.3944
R8771 gnd.n7558 gnd.n7557 19.3944
R8772 gnd.n7557 gnd.n216 19.3944
R8773 gnd.n7552 gnd.n216 19.3944
R8774 gnd.n7552 gnd.n7551 19.3944
R8775 gnd.n7551 gnd.n7550 19.3944
R8776 gnd.n7550 gnd.n223 19.3944
R8777 gnd.n7545 gnd.n223 19.3944
R8778 gnd.n7545 gnd.n7544 19.3944
R8779 gnd.n7544 gnd.n7543 19.3944
R8780 gnd.n7543 gnd.n230 19.3944
R8781 gnd.n7538 gnd.n230 19.3944
R8782 gnd.n7538 gnd.n7537 19.3944
R8783 gnd.n7537 gnd.n7536 19.3944
R8784 gnd.n7536 gnd.n237 19.3944
R8785 gnd.n7531 gnd.n237 19.3944
R8786 gnd.n7531 gnd.n7530 19.3944
R8787 gnd.n7449 gnd.n7448 19.3944
R8788 gnd.n7448 gnd.n7447 19.3944
R8789 gnd.n7447 gnd.n319 19.3944
R8790 gnd.n7442 gnd.n319 19.3944
R8791 gnd.n7442 gnd.n7441 19.3944
R8792 gnd.n7441 gnd.n7440 19.3944
R8793 gnd.n7440 gnd.n326 19.3944
R8794 gnd.n7435 gnd.n326 19.3944
R8795 gnd.n7435 gnd.n7434 19.3944
R8796 gnd.n7434 gnd.n7433 19.3944
R8797 gnd.n7433 gnd.n333 19.3944
R8798 gnd.n7428 gnd.n333 19.3944
R8799 gnd.n7428 gnd.n7427 19.3944
R8800 gnd.n7427 gnd.n7426 19.3944
R8801 gnd.n7426 gnd.n340 19.3944
R8802 gnd.n7421 gnd.n340 19.3944
R8803 gnd.n5364 gnd.n5363 19.3944
R8804 gnd.n5363 gnd.n1495 19.3944
R8805 gnd.n5911 gnd.n1495 19.3944
R8806 gnd.n5911 gnd.n1493 19.3944
R8807 gnd.n5915 gnd.n1493 19.3944
R8808 gnd.n5915 gnd.n1488 19.3944
R8809 gnd.n5934 gnd.n1488 19.3944
R8810 gnd.n5934 gnd.n1489 19.3944
R8811 gnd.n5930 gnd.n1489 19.3944
R8812 gnd.n5930 gnd.n1480 19.3944
R8813 gnd.n5992 gnd.n1480 19.3944
R8814 gnd.n5992 gnd.n1478 19.3944
R8815 gnd.n5996 gnd.n1478 19.3944
R8816 gnd.n5996 gnd.n1474 19.3944
R8817 gnd.n6006 gnd.n1474 19.3944
R8818 gnd.n6006 gnd.n1472 19.3944
R8819 gnd.n6010 gnd.n1472 19.3944
R8820 gnd.n6010 gnd.n1466 19.3944
R8821 gnd.n6035 gnd.n1466 19.3944
R8822 gnd.n6035 gnd.n1467 19.3944
R8823 gnd.n6031 gnd.n1467 19.3944
R8824 gnd.n6031 gnd.n6030 19.3944
R8825 gnd.n6030 gnd.n6029 19.3944
R8826 gnd.n6029 gnd.n6024 19.3944
R8827 gnd.n6025 gnd.n6024 19.3944
R8828 gnd.n6025 gnd.n81 19.3944
R8829 gnd.n7641 gnd.n81 19.3944
R8830 gnd.n7641 gnd.n7640 19.3944
R8831 gnd.n7640 gnd.n83 19.3944
R8832 gnd.n7326 gnd.n83 19.3944
R8833 gnd.n7326 gnd.n360 19.3944
R8834 gnd.n7331 gnd.n360 19.3944
R8835 gnd.n7331 gnd.n356 19.3944
R8836 gnd.n7345 gnd.n356 19.3944
R8837 gnd.n7346 gnd.n7345 19.3944
R8838 gnd.n7348 gnd.n7346 19.3944
R8839 gnd.n7348 gnd.n354 19.3944
R8840 gnd.n7383 gnd.n354 19.3944
R8841 gnd.n7383 gnd.n7382 19.3944
R8842 gnd.n7382 gnd.n7381 19.3944
R8843 gnd.n7381 gnd.n7379 19.3944
R8844 gnd.n7379 gnd.n7378 19.3944
R8845 gnd.n7378 gnd.n7376 19.3944
R8846 gnd.n7376 gnd.n7375 19.3944
R8847 gnd.n7375 gnd.n7373 19.3944
R8848 gnd.n7373 gnd.n7372 19.3944
R8849 gnd.n7372 gnd.n7370 19.3944
R8850 gnd.n7370 gnd.n7369 19.3944
R8851 gnd.n7369 gnd.n7367 19.3944
R8852 gnd.n7367 gnd.n7366 19.3944
R8853 gnd.n7366 gnd.n351 19.3944
R8854 gnd.n7415 gnd.n351 19.3944
R8855 gnd.n7416 gnd.n7415 19.3944
R8856 gnd.n6120 gnd.n6119 19.3944
R8857 gnd.n6119 gnd.n6118 19.3944
R8858 gnd.n6118 gnd.n1347 19.3944
R8859 gnd.n6108 gnd.n1347 19.3944
R8860 gnd.n6108 gnd.n6107 19.3944
R8861 gnd.n6107 gnd.n6106 19.3944
R8862 gnd.n6106 gnd.n1370 19.3944
R8863 gnd.n6096 gnd.n1370 19.3944
R8864 gnd.n6096 gnd.n6095 19.3944
R8865 gnd.n6095 gnd.n6094 19.3944
R8866 gnd.n6094 gnd.n1390 19.3944
R8867 gnd.n6084 gnd.n1390 19.3944
R8868 gnd.n6084 gnd.n6083 19.3944
R8869 gnd.n6083 gnd.n6082 19.3944
R8870 gnd.n6082 gnd.n1410 19.3944
R8871 gnd.n6072 gnd.n1410 19.3944
R8872 gnd.n6072 gnd.n6071 19.3944
R8873 gnd.n6071 gnd.n6070 19.3944
R8874 gnd.n6070 gnd.n1430 19.3944
R8875 gnd.n6060 gnd.n1430 19.3944
R8876 gnd.n6060 gnd.n6059 19.3944
R8877 gnd.n6059 gnd.n6058 19.3944
R8878 gnd.n1448 gnd.n97 19.3944
R8879 gnd.n7302 gnd.n97 19.3944
R8880 gnd.n380 gnd.n379 19.3944
R8881 gnd.n7636 gnd.n7635 19.3944
R8882 gnd.n7632 gnd.n92 19.3944
R8883 gnd.n7632 gnd.n99 19.3944
R8884 gnd.n7622 gnd.n99 19.3944
R8885 gnd.n7622 gnd.n7621 19.3944
R8886 gnd.n7621 gnd.n7620 19.3944
R8887 gnd.n7620 gnd.n121 19.3944
R8888 gnd.n7610 gnd.n121 19.3944
R8889 gnd.n7610 gnd.n7609 19.3944
R8890 gnd.n7609 gnd.n7608 19.3944
R8891 gnd.n7608 gnd.n141 19.3944
R8892 gnd.n7598 gnd.n141 19.3944
R8893 gnd.n7598 gnd.n7597 19.3944
R8894 gnd.n7597 gnd.n7596 19.3944
R8895 gnd.n7596 gnd.n159 19.3944
R8896 gnd.n7586 gnd.n159 19.3944
R8897 gnd.n7586 gnd.n7585 19.3944
R8898 gnd.n7585 gnd.n7584 19.3944
R8899 gnd.n7584 gnd.n179 19.3944
R8900 gnd.n7574 gnd.n179 19.3944
R8901 gnd.n7574 gnd.n7573 19.3944
R8902 gnd.n7573 gnd.n7572 19.3944
R8903 gnd.n7572 gnd.n198 19.3944
R8904 gnd.n7562 gnd.n198 19.3944
R8905 gnd.n6469 gnd.n939 19.3944
R8906 gnd.n4193 gnd.n939 19.3944
R8907 gnd.n4197 gnd.n4193 19.3944
R8908 gnd.n4197 gnd.n2172 19.3944
R8909 gnd.n4201 gnd.n2172 19.3944
R8910 gnd.n4204 gnd.n4203 19.3944
R8911 gnd.n4208 gnd.n4207 19.3944
R8912 gnd.n4213 gnd.n4212 19.3944
R8913 gnd.n4210 gnd.n2130 19.3944
R8914 gnd.n4282 gnd.n2127 19.3944
R8915 gnd.n4282 gnd.n2126 19.3944
R8916 gnd.n4286 gnd.n2126 19.3944
R8917 gnd.n4286 gnd.n2124 19.3944
R8918 gnd.n4290 gnd.n2124 19.3944
R8919 gnd.n4290 gnd.n2122 19.3944
R8920 gnd.n4313 gnd.n2122 19.3944
R8921 gnd.n4313 gnd.n4312 19.3944
R8922 gnd.n4312 gnd.n4311 19.3944
R8923 gnd.n4311 gnd.n4296 19.3944
R8924 gnd.n4307 gnd.n4296 19.3944
R8925 gnd.n4307 gnd.n4306 19.3944
R8926 gnd.n4306 gnd.n4305 19.3944
R8927 gnd.n4305 gnd.n4303 19.3944
R8928 gnd.n4303 gnd.n2099 19.3944
R8929 gnd.n4377 gnd.n2099 19.3944
R8930 gnd.n4377 gnd.n2097 19.3944
R8931 gnd.n4381 gnd.n2097 19.3944
R8932 gnd.n4381 gnd.n2095 19.3944
R8933 gnd.n4385 gnd.n2095 19.3944
R8934 gnd.n4385 gnd.n2093 19.3944
R8935 gnd.n4389 gnd.n2093 19.3944
R8936 gnd.n4389 gnd.n2091 19.3944
R8937 gnd.n4395 gnd.n2091 19.3944
R8938 gnd.n4395 gnd.n2089 19.3944
R8939 gnd.n4399 gnd.n2089 19.3944
R8940 gnd.n4399 gnd.n2066 19.3944
R8941 gnd.n4679 gnd.n2066 19.3944
R8942 gnd.n4679 gnd.n2064 19.3944
R8943 gnd.n4685 gnd.n2064 19.3944
R8944 gnd.n4685 gnd.n4684 19.3944
R8945 gnd.n4684 gnd.n2041 19.3944
R8946 gnd.n4711 gnd.n2041 19.3944
R8947 gnd.n4711 gnd.n2039 19.3944
R8948 gnd.n4718 gnd.n2039 19.3944
R8949 gnd.n4718 gnd.n4717 19.3944
R8950 gnd.n4717 gnd.n1215 19.3944
R8951 gnd.n6253 gnd.n1215 19.3944
R8952 gnd.n6253 gnd.n6252 19.3944
R8953 gnd.n6252 gnd.n6251 19.3944
R8954 gnd.n6251 gnd.n1219 19.3944
R8955 gnd.n4754 gnd.n1219 19.3944
R8956 gnd.n4754 gnd.n1915 19.3944
R8957 gnd.n4793 gnd.n1915 19.3944
R8958 gnd.n4793 gnd.n1913 19.3944
R8959 gnd.n4797 gnd.n1913 19.3944
R8960 gnd.n4797 gnd.n1897 19.3944
R8961 gnd.n4835 gnd.n1897 19.3944
R8962 gnd.n4835 gnd.n1895 19.3944
R8963 gnd.n4841 gnd.n1895 19.3944
R8964 gnd.n4841 gnd.n4840 19.3944
R8965 gnd.n4840 gnd.n1871 19.3944
R8966 gnd.n4897 gnd.n1871 19.3944
R8967 gnd.n4897 gnd.n1869 19.3944
R8968 gnd.n4901 gnd.n1869 19.3944
R8969 gnd.n4901 gnd.n1853 19.3944
R8970 gnd.n4925 gnd.n1853 19.3944
R8971 gnd.n4925 gnd.n1851 19.3944
R8972 gnd.n4931 gnd.n1851 19.3944
R8973 gnd.n4931 gnd.n4930 19.3944
R8974 gnd.n4930 gnd.n1820 19.3944
R8975 gnd.n4975 gnd.n1820 19.3944
R8976 gnd.n4975 gnd.n1818 19.3944
R8977 gnd.n4979 gnd.n1818 19.3944
R8978 gnd.n4979 gnd.n1797 19.3944
R8979 gnd.n5015 gnd.n1797 19.3944
R8980 gnd.n5015 gnd.n1795 19.3944
R8981 gnd.n5019 gnd.n1795 19.3944
R8982 gnd.n5019 gnd.n1775 19.3944
R8983 gnd.n5072 gnd.n1775 19.3944
R8984 gnd.n5072 gnd.n1773 19.3944
R8985 gnd.n5076 gnd.n1773 19.3944
R8986 gnd.n5076 gnd.n1755 19.3944
R8987 gnd.n5097 gnd.n1755 19.3944
R8988 gnd.n5097 gnd.n1753 19.3944
R8989 gnd.n5101 gnd.n1753 19.3944
R8990 gnd.n5101 gnd.n1735 19.3944
R8991 gnd.n5157 gnd.n1735 19.3944
R8992 gnd.n5157 gnd.n1733 19.3944
R8993 gnd.n5161 gnd.n1733 19.3944
R8994 gnd.n5161 gnd.n1713 19.3944
R8995 gnd.n5186 gnd.n1713 19.3944
R8996 gnd.n5186 gnd.n1711 19.3944
R8997 gnd.n5192 gnd.n1711 19.3944
R8998 gnd.n5192 gnd.n5191 19.3944
R8999 gnd.n5191 gnd.n1685 19.3944
R9000 gnd.n5237 gnd.n1685 19.3944
R9001 gnd.n5237 gnd.n1683 19.3944
R9002 gnd.n5241 gnd.n1683 19.3944
R9003 gnd.n5241 gnd.n1665 19.3944
R9004 gnd.n5263 gnd.n1665 19.3944
R9005 gnd.n5263 gnd.n1663 19.3944
R9006 gnd.n5269 gnd.n1663 19.3944
R9007 gnd.n5269 gnd.n5268 19.3944
R9008 gnd.n5268 gnd.n1635 19.3944
R9009 gnd.n5307 gnd.n1635 19.3944
R9010 gnd.n5307 gnd.n1633 19.3944
R9011 gnd.n5314 gnd.n1633 19.3944
R9012 gnd.n5314 gnd.n5313 19.3944
R9013 gnd.n5313 gnd.n1584 19.3944
R9014 gnd.n5560 gnd.n1584 19.3944
R9015 gnd.n5560 gnd.n5559 19.3944
R9016 gnd.n5559 gnd.n5558 19.3944
R9017 gnd.n5558 gnd.n1588 19.3944
R9018 gnd.n1595 gnd.n1588 19.3944
R9019 gnd.n5548 gnd.n1595 19.3944
R9020 gnd.n5548 gnd.n5547 19.3944
R9021 gnd.n5547 gnd.n5546 19.3944
R9022 gnd.n5546 gnd.n1603 19.3944
R9023 gnd.n1603 gnd.n1322 19.3944
R9024 gnd.n6135 gnd.n1322 19.3944
R9025 gnd.n6135 gnd.n6134 19.3944
R9026 gnd.n6134 gnd.n6133 19.3944
R9027 gnd.n6133 gnd.n1326 19.3944
R9028 gnd.n6127 gnd.n1326 19.3944
R9029 gnd.n6127 gnd.n6126 19.3944
R9030 gnd.n6126 gnd.n6125 19.3944
R9031 gnd.n6125 gnd.n1335 19.3944
R9032 gnd.n5946 gnd.n1335 19.3944
R9033 gnd.n5946 gnd.n5943 19.3944
R9034 gnd.n5950 gnd.n5943 19.3944
R9035 gnd.n5950 gnd.n5941 19.3944
R9036 gnd.n5954 gnd.n5941 19.3944
R9037 gnd.n5954 gnd.n5939 19.3944
R9038 gnd.n5958 gnd.n5939 19.3944
R9039 gnd.n5958 gnd.n1486 19.3944
R9040 gnd.n5962 gnd.n1486 19.3944
R9041 gnd.n5962 gnd.n1484 19.3944
R9042 gnd.n5987 gnd.n1484 19.3944
R9043 gnd.n5987 gnd.n5986 19.3944
R9044 gnd.n5986 gnd.n5985 19.3944
R9045 gnd.n5985 gnd.n5968 19.3944
R9046 gnd.n5981 gnd.n5968 19.3944
R9047 gnd.n5981 gnd.n5980 19.3944
R9048 gnd.n5980 gnd.n5979 19.3944
R9049 gnd.n5979 gnd.n5977 19.3944
R9050 gnd.n5977 gnd.n1464 19.3944
R9051 gnd.n1464 gnd.n1462 19.3944
R9052 gnd.n6042 gnd.n1462 19.3944
R9053 gnd.n6046 gnd.n6044 19.3944
R9054 gnd.n7296 gnd.n383 19.3944
R9055 gnd.n7294 gnd.n7293 19.3944
R9056 gnd.n7290 gnd.n7289 19.3944
R9057 gnd.n7287 gnd.n386 19.3944
R9058 gnd.n7283 gnd.n386 19.3944
R9059 gnd.n7283 gnd.n7282 19.3944
R9060 gnd.n7282 gnd.n7281 19.3944
R9061 gnd.n7281 gnd.n392 19.3944
R9062 gnd.n4040 gnd.n4039 19.3944
R9063 gnd.n4039 gnd.n4038 19.3944
R9064 gnd.n4038 gnd.n4037 19.3944
R9065 gnd.n4037 gnd.n4035 19.3944
R9066 gnd.n4035 gnd.n4032 19.3944
R9067 gnd.n4032 gnd.n4031 19.3944
R9068 gnd.n4031 gnd.n4028 19.3944
R9069 gnd.n4028 gnd.n4027 19.3944
R9070 gnd.n4027 gnd.n4024 19.3944
R9071 gnd.n4024 gnd.n4023 19.3944
R9072 gnd.n4023 gnd.n4020 19.3944
R9073 gnd.n4020 gnd.n4019 19.3944
R9074 gnd.n4019 gnd.n4016 19.3944
R9075 gnd.n4016 gnd.n4015 19.3944
R9076 gnd.n4015 gnd.n4012 19.3944
R9077 gnd.n4012 gnd.n4011 19.3944
R9078 gnd.n4011 gnd.n4008 19.3944
R9079 gnd.n4006 gnd.n4003 19.3944
R9080 gnd.n4003 gnd.n4002 19.3944
R9081 gnd.n4002 gnd.n3999 19.3944
R9082 gnd.n3999 gnd.n3998 19.3944
R9083 gnd.n3998 gnd.n3995 19.3944
R9084 gnd.n3995 gnd.n3994 19.3944
R9085 gnd.n3994 gnd.n3991 19.3944
R9086 gnd.n3991 gnd.n3990 19.3944
R9087 gnd.n3990 gnd.n3987 19.3944
R9088 gnd.n3987 gnd.n3986 19.3944
R9089 gnd.n3986 gnd.n3983 19.3944
R9090 gnd.n3983 gnd.n3982 19.3944
R9091 gnd.n3982 gnd.n3979 19.3944
R9092 gnd.n3979 gnd.n3978 19.3944
R9093 gnd.n3978 gnd.n3975 19.3944
R9094 gnd.n3975 gnd.n3974 19.3944
R9095 gnd.n3974 gnd.n3971 19.3944
R9096 gnd.n3971 gnd.n3970 19.3944
R9097 gnd.n3966 gnd.n3963 19.3944
R9098 gnd.n3963 gnd.n3962 19.3944
R9099 gnd.n3962 gnd.n3959 19.3944
R9100 gnd.n3959 gnd.n3958 19.3944
R9101 gnd.n3958 gnd.n3955 19.3944
R9102 gnd.n3955 gnd.n3954 19.3944
R9103 gnd.n3954 gnd.n3951 19.3944
R9104 gnd.n3951 gnd.n3950 19.3944
R9105 gnd.n3950 gnd.n3947 19.3944
R9106 gnd.n3947 gnd.n3946 19.3944
R9107 gnd.n3946 gnd.n3943 19.3944
R9108 gnd.n3943 gnd.n3942 19.3944
R9109 gnd.n3942 gnd.n3939 19.3944
R9110 gnd.n3939 gnd.n3938 19.3944
R9111 gnd.n3938 gnd.n3935 19.3944
R9112 gnd.n3935 gnd.n3934 19.3944
R9113 gnd.n3934 gnd.n3931 19.3944
R9114 gnd.n3931 gnd.n3930 19.3944
R9115 gnd.n3923 gnd.n3921 19.3944
R9116 gnd.n3921 gnd.n3918 19.3944
R9117 gnd.n3918 gnd.n3917 19.3944
R9118 gnd.n3917 gnd.n3914 19.3944
R9119 gnd.n3914 gnd.n3913 19.3944
R9120 gnd.n3913 gnd.n3910 19.3944
R9121 gnd.n3910 gnd.n3909 19.3944
R9122 gnd.n3909 gnd.n3906 19.3944
R9123 gnd.n3906 gnd.n3905 19.3944
R9124 gnd.n3905 gnd.n3902 19.3944
R9125 gnd.n3902 gnd.n3901 19.3944
R9126 gnd.n3901 gnd.n3898 19.3944
R9127 gnd.n3898 gnd.n3897 19.3944
R9128 gnd.n3897 gnd.n3894 19.3944
R9129 gnd.n3894 gnd.n3893 19.3944
R9130 gnd.n3893 gnd.n3890 19.3944
R9131 gnd.n3884 gnd.n3882 19.3944
R9132 gnd.n3882 gnd.n3881 19.3944
R9133 gnd.n3881 gnd.n3879 19.3944
R9134 gnd.n3879 gnd.n3878 19.3944
R9135 gnd.n3878 gnd.n3876 19.3944
R9136 gnd.n3876 gnd.n2229 19.3944
R9137 gnd.n4089 gnd.n2229 19.3944
R9138 gnd.n4089 gnd.n2227 19.3944
R9139 gnd.n4097 gnd.n2227 19.3944
R9140 gnd.n4097 gnd.n4096 19.3944
R9141 gnd.n4096 gnd.n4095 19.3944
R9142 gnd.n4095 gnd.n2204 19.3944
R9143 gnd.n4124 gnd.n2204 19.3944
R9144 gnd.n4124 gnd.n2202 19.3944
R9145 gnd.n4134 gnd.n2202 19.3944
R9146 gnd.n4134 gnd.n4133 19.3944
R9147 gnd.n4133 gnd.n4132 19.3944
R9148 gnd.n4132 gnd.n2174 19.3944
R9149 gnd.n4188 gnd.n2174 19.3944
R9150 gnd.n4188 gnd.n4187 19.3944
R9151 gnd.n4187 gnd.n4186 19.3944
R9152 gnd.n4186 gnd.n2178 19.3944
R9153 gnd.n4170 gnd.n2178 19.3944
R9154 gnd.n4174 gnd.n4170 19.3944
R9155 gnd.n4174 gnd.n2152 19.3944
R9156 gnd.n4229 gnd.n2152 19.3944
R9157 gnd.n4229 gnd.n2150 19.3944
R9158 gnd.n4234 gnd.n2150 19.3944
R9159 gnd.n4234 gnd.n2134 19.3944
R9160 gnd.n4275 gnd.n2134 19.3944
R9161 gnd.n4275 gnd.n2135 19.3944
R9162 gnd.n4271 gnd.n2135 19.3944
R9163 gnd.n4271 gnd.n4270 19.3944
R9164 gnd.n4270 gnd.n4269 19.3944
R9165 gnd.n4269 gnd.n2140 19.3944
R9166 gnd.n4265 gnd.n2140 19.3944
R9167 gnd.n4265 gnd.n2118 19.3944
R9168 gnd.n4318 gnd.n2118 19.3944
R9169 gnd.n4318 gnd.n2116 19.3944
R9170 gnd.n4322 gnd.n2116 19.3944
R9171 gnd.n4322 gnd.n2113 19.3944
R9172 gnd.n4333 gnd.n2113 19.3944
R9173 gnd.n4333 gnd.n2111 19.3944
R9174 gnd.n4337 gnd.n2111 19.3944
R9175 gnd.n4337 gnd.n2102 19.3944
R9176 gnd.n4371 gnd.n2102 19.3944
R9177 gnd.n4371 gnd.n2103 19.3944
R9178 gnd.n4367 gnd.n2103 19.3944
R9179 gnd.n4367 gnd.n4366 19.3944
R9180 gnd.n4366 gnd.n4365 19.3944
R9181 gnd.n4365 gnd.n2108 19.3944
R9182 gnd.n4361 gnd.n2108 19.3944
R9183 gnd.n4361 gnd.n4360 19.3944
R9184 gnd.n4049 gnd.n4047 19.3944
R9185 gnd.n4049 gnd.n4048 19.3944
R9186 gnd.n4048 gnd.n2248 19.3944
R9187 gnd.n4064 gnd.n2248 19.3944
R9188 gnd.n4065 gnd.n4064 19.3944
R9189 gnd.n4067 gnd.n4065 19.3944
R9190 gnd.n4068 gnd.n4067 19.3944
R9191 gnd.n4068 gnd.n2222 19.3944
R9192 gnd.n4101 gnd.n2222 19.3944
R9193 gnd.n4102 gnd.n4101 19.3944
R9194 gnd.n4104 gnd.n4102 19.3944
R9195 gnd.n4107 gnd.n4104 19.3944
R9196 gnd.n4107 gnd.n4106 19.3944
R9197 gnd.n4106 gnd.n2198 19.3944
R9198 gnd.n4138 gnd.n2198 19.3944
R9199 gnd.n4138 gnd.n2201 19.3944
R9200 gnd.n2201 gnd.n2200 19.3944
R9201 gnd.n2200 gnd.n2179 19.3944
R9202 gnd.n4159 gnd.n2179 19.3944
R9203 gnd.n4160 gnd.n4159 19.3944
R9204 gnd.n4182 gnd.n4160 19.3944
R9205 gnd.n4182 gnd.n4181 19.3944
R9206 gnd.n4181 gnd.n4180 19.3944
R9207 gnd.n4180 gnd.n4167 19.3944
R9208 gnd.n4167 gnd.n4166 19.3944
R9209 gnd.n4166 gnd.n4165 19.3944
R9210 gnd.n4165 gnd.n4164 19.3944
R9211 gnd.n4164 gnd.n4163 19.3944
R9212 gnd.n4163 gnd.n2141 19.3944
R9213 gnd.n4246 gnd.n2141 19.3944
R9214 gnd.n4247 gnd.n4246 19.3944
R9215 gnd.n4250 gnd.n4247 19.3944
R9216 gnd.n4251 gnd.n4250 19.3944
R9217 gnd.n4256 gnd.n4251 19.3944
R9218 gnd.n4257 gnd.n4256 19.3944
R9219 gnd.n4261 gnd.n4257 19.3944
R9220 gnd.n4261 gnd.n4260 19.3944
R9221 gnd.n4260 gnd.n4259 19.3944
R9222 gnd.n4259 gnd.n2115 19.3944
R9223 gnd.n4326 gnd.n2115 19.3944
R9224 gnd.n4327 gnd.n4326 19.3944
R9225 gnd.n4329 gnd.n4327 19.3944
R9226 gnd.n4329 gnd.n2110 19.3944
R9227 gnd.n4341 gnd.n2110 19.3944
R9228 gnd.n4342 gnd.n4341 19.3944
R9229 gnd.n4344 gnd.n4342 19.3944
R9230 gnd.n4345 gnd.n4344 19.3944
R9231 gnd.n4348 gnd.n4345 19.3944
R9232 gnd.n4349 gnd.n4348 19.3944
R9233 gnd.n4353 gnd.n4349 19.3944
R9234 gnd.n4354 gnd.n4353 19.3944
R9235 gnd.n4356 gnd.n4354 19.3944
R9236 gnd.n4356 gnd.n4355 19.3944
R9237 gnd.n4051 gnd.n2264 19.3944
R9238 gnd.n4051 gnd.n2265 19.3944
R9239 gnd.n2267 gnd.n2265 19.3944
R9240 gnd.n2267 gnd.n2245 19.3944
R9241 gnd.n4075 gnd.n2245 19.3944
R9242 gnd.n4075 gnd.n4074 19.3944
R9243 gnd.n4074 gnd.n4073 19.3944
R9244 gnd.n4073 gnd.n4072 19.3944
R9245 gnd.n4072 gnd.n2218 19.3944
R9246 gnd.n4111 gnd.n2218 19.3944
R9247 gnd.n4111 gnd.n4110 19.3944
R9248 gnd.n4110 gnd.n4109 19.3944
R9249 gnd.n4109 gnd.n2195 19.3944
R9250 gnd.n4141 gnd.n2195 19.3944
R9251 gnd.n4141 gnd.n4140 19.3944
R9252 gnd.n4140 gnd.n2181 19.3944
R9253 gnd.n4155 gnd.n2181 19.3944
R9254 gnd.n4156 gnd.n4155 19.3944
R9255 gnd.n4156 gnd.n959 19.3944
R9256 gnd.n6458 gnd.n959 19.3944
R9257 gnd.n6458 gnd.n6457 19.3944
R9258 gnd.n6457 gnd.n6456 19.3944
R9259 gnd.n6456 gnd.n963 19.3944
R9260 gnd.n2163 gnd.n963 19.3944
R9261 gnd.n4220 gnd.n2163 19.3944
R9262 gnd.n4220 gnd.n4219 19.3944
R9263 gnd.n4219 gnd.n4218 19.3944
R9264 gnd.n4218 gnd.n2143 19.3944
R9265 gnd.n4243 gnd.n2143 19.3944
R9266 gnd.n4243 gnd.n987 19.3944
R9267 gnd.n6445 gnd.n987 19.3944
R9268 gnd.n6445 gnd.n6444 19.3944
R9269 gnd.n6444 gnd.n6443 19.3944
R9270 gnd.n6443 gnd.n991 19.3944
R9271 gnd.n6433 gnd.n991 19.3944
R9272 gnd.n6433 gnd.n6432 19.3944
R9273 gnd.n6432 gnd.n6431 19.3944
R9274 gnd.n6431 gnd.n1010 19.3944
R9275 gnd.n6421 gnd.n1010 19.3944
R9276 gnd.n6421 gnd.n6420 19.3944
R9277 gnd.n6420 gnd.n6419 19.3944
R9278 gnd.n6419 gnd.n1030 19.3944
R9279 gnd.n6409 gnd.n1030 19.3944
R9280 gnd.n6409 gnd.n6408 19.3944
R9281 gnd.n6408 gnd.n6407 19.3944
R9282 gnd.n6407 gnd.n1050 19.3944
R9283 gnd.n6397 gnd.n1050 19.3944
R9284 gnd.n6397 gnd.n6396 19.3944
R9285 gnd.n6396 gnd.n6395 19.3944
R9286 gnd.n6395 gnd.n1070 19.3944
R9287 gnd.n6385 gnd.n1070 19.3944
R9288 gnd.n6385 gnd.n6384 19.3944
R9289 gnd.n6384 gnd.n6383 19.3944
R9290 gnd.n6376 gnd.n6375 19.3944
R9291 gnd.n6375 gnd.n1099 19.3944
R9292 gnd.n1101 gnd.n1099 19.3944
R9293 gnd.n6368 gnd.n1101 19.3944
R9294 gnd.n6368 gnd.n6367 19.3944
R9295 gnd.n6367 gnd.n6366 19.3944
R9296 gnd.n6366 gnd.n1108 19.3944
R9297 gnd.n6361 gnd.n1108 19.3944
R9298 gnd.n6361 gnd.n6360 19.3944
R9299 gnd.n6360 gnd.n6359 19.3944
R9300 gnd.n6359 gnd.n1115 19.3944
R9301 gnd.n6354 gnd.n1115 19.3944
R9302 gnd.n6354 gnd.n6353 19.3944
R9303 gnd.n6353 gnd.n6352 19.3944
R9304 gnd.n6352 gnd.n1122 19.3944
R9305 gnd.n6347 gnd.n1122 19.3944
R9306 gnd.n6347 gnd.n6346 19.3944
R9307 gnd.n4484 gnd.n4444 19.3944
R9308 gnd.n4488 gnd.n4444 19.3944
R9309 gnd.n4488 gnd.n4442 19.3944
R9310 gnd.n4494 gnd.n4442 19.3944
R9311 gnd.n4494 gnd.n4440 19.3944
R9312 gnd.n4498 gnd.n4440 19.3944
R9313 gnd.n4498 gnd.n4438 19.3944
R9314 gnd.n4504 gnd.n4438 19.3944
R9315 gnd.n4504 gnd.n4436 19.3944
R9316 gnd.n4508 gnd.n4436 19.3944
R9317 gnd.n4508 gnd.n4434 19.3944
R9318 gnd.n4514 gnd.n4434 19.3944
R9319 gnd.n4514 gnd.n4432 19.3944
R9320 gnd.n4518 gnd.n4432 19.3944
R9321 gnd.n4518 gnd.n4430 19.3944
R9322 gnd.n4524 gnd.n4430 19.3944
R9323 gnd.n4524 gnd.n4428 19.3944
R9324 gnd.n4528 gnd.n4428 19.3944
R9325 gnd.n4457 gnd.n1144 19.3944
R9326 gnd.n4464 gnd.n4457 19.3944
R9327 gnd.n4464 gnd.n4454 19.3944
R9328 gnd.n4468 gnd.n4454 19.3944
R9329 gnd.n4468 gnd.n4452 19.3944
R9330 gnd.n4474 gnd.n4452 19.3944
R9331 gnd.n4474 gnd.n4450 19.3944
R9332 gnd.n4478 gnd.n4450 19.3944
R9333 gnd.n6344 gnd.n1131 19.3944
R9334 gnd.n6339 gnd.n1131 19.3944
R9335 gnd.n6339 gnd.n6338 19.3944
R9336 gnd.n6338 gnd.n6337 19.3944
R9337 gnd.n6337 gnd.n1138 19.3944
R9338 gnd.n6332 gnd.n1138 19.3944
R9339 gnd.n6332 gnd.n6331 19.3944
R9340 gnd.n4055 gnd.n2257 19.3944
R9341 gnd.n4055 gnd.n2255 19.3944
R9342 gnd.n4059 gnd.n2255 19.3944
R9343 gnd.n4059 gnd.n2237 19.3944
R9344 gnd.n4079 gnd.n2237 19.3944
R9345 gnd.n4079 gnd.n2235 19.3944
R9346 gnd.n4085 gnd.n2235 19.3944
R9347 gnd.n4085 gnd.n4084 19.3944
R9348 gnd.n4084 gnd.n2211 19.3944
R9349 gnd.n4115 gnd.n2211 19.3944
R9350 gnd.n4115 gnd.n2209 19.3944
R9351 gnd.n4119 gnd.n2209 19.3944
R9352 gnd.n4119 gnd.n2189 19.3944
R9353 gnd.n4145 gnd.n2189 19.3944
R9354 gnd.n4145 gnd.n2187 19.3944
R9355 gnd.n4150 gnd.n2187 19.3944
R9356 gnd.n4150 gnd.n948 19.3944
R9357 gnd.n6464 gnd.n948 19.3944
R9358 gnd.n6464 gnd.n6463 19.3944
R9359 gnd.n6463 gnd.n6462 19.3944
R9360 gnd.n6462 gnd.n952 19.3944
R9361 gnd.n6452 gnd.n952 19.3944
R9362 gnd.n977 gnd.n970 19.3944
R9363 gnd.n2158 gnd.n977 19.3944
R9364 gnd.n4225 gnd.n4224 19.3944
R9365 gnd.n4239 gnd.n4238 19.3944
R9366 gnd.n6449 gnd.n978 19.3944
R9367 gnd.n6449 gnd.n979 19.3944
R9368 gnd.n6439 gnd.n979 19.3944
R9369 gnd.n6439 gnd.n6438 19.3944
R9370 gnd.n6438 gnd.n6437 19.3944
R9371 gnd.n6437 gnd.n1000 19.3944
R9372 gnd.n6427 gnd.n1000 19.3944
R9373 gnd.n6427 gnd.n6426 19.3944
R9374 gnd.n6426 gnd.n6425 19.3944
R9375 gnd.n6425 gnd.n1021 19.3944
R9376 gnd.n6415 gnd.n1021 19.3944
R9377 gnd.n6415 gnd.n6414 19.3944
R9378 gnd.n6414 gnd.n6413 19.3944
R9379 gnd.n6413 gnd.n1040 19.3944
R9380 gnd.n6403 gnd.n1040 19.3944
R9381 gnd.n6403 gnd.n6402 19.3944
R9382 gnd.n6402 gnd.n6401 19.3944
R9383 gnd.n6401 gnd.n1061 19.3944
R9384 gnd.n6391 gnd.n1061 19.3944
R9385 gnd.n6391 gnd.n6390 19.3944
R9386 gnd.n6390 gnd.n6389 19.3944
R9387 gnd.n6389 gnd.n1081 19.3944
R9388 gnd.n6379 gnd.n1081 19.3944
R9389 gnd.n6640 gnd.n6639 19.3944
R9390 gnd.n6639 gnd.n772 19.3944
R9391 gnd.n6633 gnd.n772 19.3944
R9392 gnd.n6633 gnd.n6632 19.3944
R9393 gnd.n6632 gnd.n6631 19.3944
R9394 gnd.n6631 gnd.n780 19.3944
R9395 gnd.n6625 gnd.n780 19.3944
R9396 gnd.n6625 gnd.n6624 19.3944
R9397 gnd.n6624 gnd.n6623 19.3944
R9398 gnd.n6623 gnd.n788 19.3944
R9399 gnd.n6617 gnd.n788 19.3944
R9400 gnd.n6617 gnd.n6616 19.3944
R9401 gnd.n6616 gnd.n6615 19.3944
R9402 gnd.n6615 gnd.n796 19.3944
R9403 gnd.n6609 gnd.n796 19.3944
R9404 gnd.n6609 gnd.n6608 19.3944
R9405 gnd.n6608 gnd.n6607 19.3944
R9406 gnd.n6607 gnd.n804 19.3944
R9407 gnd.n6601 gnd.n804 19.3944
R9408 gnd.n6601 gnd.n6600 19.3944
R9409 gnd.n6600 gnd.n6599 19.3944
R9410 gnd.n6599 gnd.n812 19.3944
R9411 gnd.n6593 gnd.n812 19.3944
R9412 gnd.n6593 gnd.n6592 19.3944
R9413 gnd.n6592 gnd.n6591 19.3944
R9414 gnd.n6591 gnd.n820 19.3944
R9415 gnd.n6585 gnd.n820 19.3944
R9416 gnd.n6585 gnd.n6584 19.3944
R9417 gnd.n6584 gnd.n6583 19.3944
R9418 gnd.n6583 gnd.n828 19.3944
R9419 gnd.n6577 gnd.n828 19.3944
R9420 gnd.n6577 gnd.n6576 19.3944
R9421 gnd.n6576 gnd.n6575 19.3944
R9422 gnd.n6575 gnd.n836 19.3944
R9423 gnd.n6569 gnd.n836 19.3944
R9424 gnd.n6569 gnd.n6568 19.3944
R9425 gnd.n6568 gnd.n6567 19.3944
R9426 gnd.n6567 gnd.n844 19.3944
R9427 gnd.n6561 gnd.n844 19.3944
R9428 gnd.n6561 gnd.n6560 19.3944
R9429 gnd.n6560 gnd.n6559 19.3944
R9430 gnd.n6559 gnd.n852 19.3944
R9431 gnd.n6553 gnd.n852 19.3944
R9432 gnd.n6553 gnd.n6552 19.3944
R9433 gnd.n6552 gnd.n6551 19.3944
R9434 gnd.n6551 gnd.n860 19.3944
R9435 gnd.n6545 gnd.n860 19.3944
R9436 gnd.n6545 gnd.n6544 19.3944
R9437 gnd.n6544 gnd.n6543 19.3944
R9438 gnd.n6543 gnd.n868 19.3944
R9439 gnd.n6537 gnd.n868 19.3944
R9440 gnd.n6537 gnd.n6536 19.3944
R9441 gnd.n6536 gnd.n6535 19.3944
R9442 gnd.n6535 gnd.n876 19.3944
R9443 gnd.n6529 gnd.n876 19.3944
R9444 gnd.n6529 gnd.n6528 19.3944
R9445 gnd.n6528 gnd.n6527 19.3944
R9446 gnd.n6527 gnd.n884 19.3944
R9447 gnd.n6521 gnd.n884 19.3944
R9448 gnd.n6521 gnd.n6520 19.3944
R9449 gnd.n6520 gnd.n6519 19.3944
R9450 gnd.n6519 gnd.n892 19.3944
R9451 gnd.n6513 gnd.n892 19.3944
R9452 gnd.n6513 gnd.n6512 19.3944
R9453 gnd.n6512 gnd.n6511 19.3944
R9454 gnd.n6511 gnd.n900 19.3944
R9455 gnd.n6505 gnd.n900 19.3944
R9456 gnd.n6505 gnd.n6504 19.3944
R9457 gnd.n6504 gnd.n6503 19.3944
R9458 gnd.n6503 gnd.n908 19.3944
R9459 gnd.n6497 gnd.n908 19.3944
R9460 gnd.n6497 gnd.n6496 19.3944
R9461 gnd.n6496 gnd.n6495 19.3944
R9462 gnd.n6495 gnd.n916 19.3944
R9463 gnd.n6489 gnd.n916 19.3944
R9464 gnd.n6489 gnd.n6488 19.3944
R9465 gnd.n6488 gnd.n6487 19.3944
R9466 gnd.n6487 gnd.n924 19.3944
R9467 gnd.n6481 gnd.n924 19.3944
R9468 gnd.n6481 gnd.n6480 19.3944
R9469 gnd.n6480 gnd.n6479 19.3944
R9470 gnd.n6479 gnd.n932 19.3944
R9471 gnd.n6473 gnd.n932 19.3944
R9472 gnd.n6473 gnd.n6472 19.3944
R9473 gnd.n4690 gnd.n2057 19.3944
R9474 gnd.n4690 gnd.n2054 19.3944
R9475 gnd.n4695 gnd.n2054 19.3944
R9476 gnd.n4695 gnd.n2055 19.3944
R9477 gnd.n2055 gnd.n2033 19.3944
R9478 gnd.n4723 gnd.n2033 19.3944
R9479 gnd.n4723 gnd.n2030 19.3944
R9480 gnd.n4731 gnd.n2030 19.3944
R9481 gnd.n4731 gnd.n2031 19.3944
R9482 gnd.n4727 gnd.n2031 19.3944
R9483 gnd.n4727 gnd.n1226 19.3944
R9484 gnd.n6246 gnd.n1226 19.3944
R9485 gnd.n6246 gnd.n1227 19.3944
R9486 gnd.n6242 gnd.n1227 19.3944
R9487 gnd.n6242 gnd.n6241 19.3944
R9488 gnd.n6241 gnd.n6240 19.3944
R9489 gnd.n6240 gnd.n1233 19.3944
R9490 gnd.n6236 gnd.n1233 19.3944
R9491 gnd.n6236 gnd.n6235 19.3944
R9492 gnd.n6235 gnd.n6234 19.3944
R9493 gnd.n6234 gnd.n1238 19.3944
R9494 gnd.n6230 gnd.n1238 19.3944
R9495 gnd.n6230 gnd.n6229 19.3944
R9496 gnd.n6229 gnd.n6228 19.3944
R9497 gnd.n6228 gnd.n1243 19.3944
R9498 gnd.n6224 gnd.n1243 19.3944
R9499 gnd.n6224 gnd.n6223 19.3944
R9500 gnd.n6223 gnd.n6222 19.3944
R9501 gnd.n6222 gnd.n1248 19.3944
R9502 gnd.n6218 gnd.n1248 19.3944
R9503 gnd.n6218 gnd.n6217 19.3944
R9504 gnd.n6217 gnd.n6216 19.3944
R9505 gnd.n6216 gnd.n1253 19.3944
R9506 gnd.n6212 gnd.n1253 19.3944
R9507 gnd.n6212 gnd.n6211 19.3944
R9508 gnd.n6211 gnd.n6210 19.3944
R9509 gnd.n6210 gnd.n1258 19.3944
R9510 gnd.n6206 gnd.n1258 19.3944
R9511 gnd.n6206 gnd.n6205 19.3944
R9512 gnd.n6205 gnd.n6204 19.3944
R9513 gnd.n6204 gnd.n1263 19.3944
R9514 gnd.n6200 gnd.n1263 19.3944
R9515 gnd.n6200 gnd.n6199 19.3944
R9516 gnd.n6199 gnd.n6198 19.3944
R9517 gnd.n6198 gnd.n1268 19.3944
R9518 gnd.n6194 gnd.n1268 19.3944
R9519 gnd.n6194 gnd.n6193 19.3944
R9520 gnd.n6193 gnd.n6192 19.3944
R9521 gnd.n6192 gnd.n1273 19.3944
R9522 gnd.n6188 gnd.n1273 19.3944
R9523 gnd.n6188 gnd.n6187 19.3944
R9524 gnd.n6187 gnd.n6186 19.3944
R9525 gnd.n6186 gnd.n1278 19.3944
R9526 gnd.n6182 gnd.n1278 19.3944
R9527 gnd.n6182 gnd.n6181 19.3944
R9528 gnd.n6181 gnd.n6180 19.3944
R9529 gnd.n6180 gnd.n1283 19.3944
R9530 gnd.n6176 gnd.n1283 19.3944
R9531 gnd.n6176 gnd.n6175 19.3944
R9532 gnd.n6175 gnd.n6174 19.3944
R9533 gnd.n6174 gnd.n1288 19.3944
R9534 gnd.n6170 gnd.n1288 19.3944
R9535 gnd.n6170 gnd.n6169 19.3944
R9536 gnd.n6169 gnd.n6168 19.3944
R9537 gnd.n6168 gnd.n1293 19.3944
R9538 gnd.n6164 gnd.n1293 19.3944
R9539 gnd.n6164 gnd.n6163 19.3944
R9540 gnd.n6163 gnd.n6162 19.3944
R9541 gnd.n6162 gnd.n1298 19.3944
R9542 gnd.n6158 gnd.n1298 19.3944
R9543 gnd.n6158 gnd.n6157 19.3944
R9544 gnd.n6157 gnd.n6156 19.3944
R9545 gnd.n6156 gnd.n1303 19.3944
R9546 gnd.n6152 gnd.n1303 19.3944
R9547 gnd.n6152 gnd.n6151 19.3944
R9548 gnd.n6151 gnd.n6150 19.3944
R9549 gnd.n6150 gnd.n1308 19.3944
R9550 gnd.n6146 gnd.n1308 19.3944
R9551 gnd.n6146 gnd.n6145 19.3944
R9552 gnd.n6145 gnd.n6144 19.3944
R9553 gnd.n6144 gnd.n1313 19.3944
R9554 gnd.n6140 gnd.n1313 19.3944
R9555 gnd.n5425 gnd.n5423 19.3944
R9556 gnd.n5425 gnd.n5421 19.3944
R9557 gnd.n5431 gnd.n5421 19.3944
R9558 gnd.n5431 gnd.n5419 19.3944
R9559 gnd.n5436 gnd.n5419 19.3944
R9560 gnd.n5436 gnd.n5417 19.3944
R9561 gnd.n5442 gnd.n5417 19.3944
R9562 gnd.n5442 gnd.n5416 19.3944
R9563 gnd.n5451 gnd.n5416 19.3944
R9564 gnd.n5451 gnd.n5414 19.3944
R9565 gnd.n5457 gnd.n5414 19.3944
R9566 gnd.n5457 gnd.n5407 19.3944
R9567 gnd.n5470 gnd.n5407 19.3944
R9568 gnd.n5470 gnd.n5405 19.3944
R9569 gnd.n5476 gnd.n5405 19.3944
R9570 gnd.n5476 gnd.n5398 19.3944
R9571 gnd.n5489 gnd.n5398 19.3944
R9572 gnd.n5489 gnd.n5396 19.3944
R9573 gnd.n5495 gnd.n5396 19.3944
R9574 gnd.n5495 gnd.n5389 19.3944
R9575 gnd.n5508 gnd.n5389 19.3944
R9576 gnd.n5508 gnd.n5387 19.3944
R9577 gnd.n5515 gnd.n5387 19.3944
R9578 gnd.n5515 gnd.n5514 19.3944
R9579 gnd.n5528 gnd.n5368 19.3944
R9580 gnd.n5368 gnd.n5367 19.3944
R9581 gnd.n5535 gnd.n5367 19.3944
R9582 gnd.n6260 gnd.n6259 19.2005
R9583 gnd.n5652 gnd.n5651 19.2005
R9584 gnd.n3136 gnd.t128 18.8012
R9585 gnd.n3121 gnd.t288 18.8012
R9586 gnd.n2980 gnd.n2979 18.4825
R9587 gnd.n5817 gnd.n5725 18.4247
R9588 gnd.n6331 gnd.n6330 18.4247
R9589 gnd.n5525 gnd.n5524 18.2308
R9590 gnd.n4661 gnd.n2077 18.2308
R9591 gnd.n7421 gnd.n7420 18.2308
R9592 gnd.n3890 gnd.n3870 18.2308
R9593 gnd.t127 gnd.n2660 18.1639
R9594 gnd.n2688 gnd.t110 17.5266
R9595 gnd.n2242 gnd.t56 17.5266
R9596 gnd.n6399 gnd.t79 17.5266
R9597 gnd.n6104 gnd.t12 17.5266
R9598 gnd.n7582 gnd.t84 17.5266
R9599 gnd.n3087 gnd.t104 16.8893
R9600 gnd.n4143 gnd.t43 16.8893
R9601 gnd.n6423 gnd.t70 16.8893
R9602 gnd.n6080 gnd.t37 16.8893
R9603 gnd.n7606 gnd.t41 16.8893
R9604 gnd.n5847 gnd.n1523 16.6793
R9605 gnd.n7493 gnd.n7492 16.6793
R9606 gnd.n3970 gnd.n3967 16.6793
R9607 gnd.n4478 gnd.n4448 16.6793
R9608 gnd.n2915 gnd.t137 16.2519
R9609 gnd.n2615 gnd.t124 16.2519
R9610 gnd.n6447 gnd.t26 16.2519
R9611 gnd.n6056 gnd.t116 16.2519
R9612 gnd.n4655 gnd.n4401 15.9333
R9613 gnd.n4655 gnd.n2068 15.9333
R9614 gnd.n4677 gnd.n4676 15.9333
R9615 gnd.n4676 gnd.n2059 15.9333
R9616 gnd.n4688 gnd.n2059 15.9333
R9617 gnd.n4688 gnd.n4687 15.9333
R9618 gnd.n2061 gnd.n2050 15.9333
R9619 gnd.n4697 gnd.n2050 15.9333
R9620 gnd.n4697 gnd.n2051 15.9333
R9621 gnd.n2051 gnd.n2043 15.9333
R9622 gnd.n4709 gnd.n2043 15.9333
R9623 gnd.n4709 gnd.n4708 15.9333
R9624 gnd.n4708 gnd.n2035 15.9333
R9625 gnd.n4721 gnd.n2035 15.9333
R9626 gnd.n4720 gnd.n1152 15.9333
R9627 gnd.n4733 gnd.n1184 15.9333
R9628 gnd.n6255 gnd.n1212 15.9333
R9629 gnd.n4756 gnd.n1922 15.9333
R9630 gnd.n4799 gnd.n1911 15.9333
R9631 gnd.n4833 gnd.n1899 15.9333
R9632 gnd.n4845 gnd.n4843 15.9333
R9633 gnd.n4872 gnd.n1879 15.9333
R9634 gnd.n4963 gnd.n1829 15.9333
R9635 gnd.n4982 gnd.n1806 15.9333
R9636 gnd.n1813 gnd.n1801 15.9333
R9637 gnd.n5022 gnd.n1784 15.9333
R9638 gnd.n5070 gnd.n5069 15.9333
R9639 gnd.n5078 gnd.n1771 15.9333
R9640 gnd.n5095 gnd.n5094 15.9333
R9641 gnd.n5155 gnd.n1738 15.9333
R9642 gnd.n5235 gnd.n5234 15.9333
R9643 gnd.n5243 gnd.n1681 15.9333
R9644 gnd.n5261 gnd.n5260 15.9333
R9645 gnd.n5271 gnd.n1653 15.9333
R9646 gnd.n5293 gnd.n1647 15.9333
R9647 gnd.n5563 gnd.n5562 15.9333
R9648 gnd.n5346 gnd.n1573 15.9333
R9649 gnd.n5346 gnd.n1536 15.9333
R9650 gnd.n5555 gnd.n1590 15.9333
R9651 gnd.n5554 gnd.n5553 15.9333
R9652 gnd.n5553 gnd.n5552 15.9333
R9653 gnd.n5552 gnd.n5550 15.9333
R9654 gnd.n5550 gnd.n1593 15.9333
R9655 gnd.n1605 gnd.n1593 15.9333
R9656 gnd.n1606 gnd.n1605 15.9333
R9657 gnd.n5544 gnd.n1606 15.9333
R9658 gnd.n5544 gnd.n5543 15.9333
R9659 gnd.n5542 gnd.n5541 15.9333
R9660 gnd.n5541 gnd.n1317 15.9333
R9661 gnd.n6138 gnd.n1317 15.9333
R9662 gnd.n6138 gnd.n6137 15.9333
R9663 gnd.n1328 gnd.n1319 15.9333
R9664 gnd.n6131 gnd.n1328 15.9333
R9665 gnd.n3602 gnd.n3600 15.6674
R9666 gnd.n3570 gnd.n3568 15.6674
R9667 gnd.n3538 gnd.n3536 15.6674
R9668 gnd.n3507 gnd.n3505 15.6674
R9669 gnd.n3475 gnd.n3473 15.6674
R9670 gnd.n3443 gnd.n3441 15.6674
R9671 gnd.n3411 gnd.n3409 15.6674
R9672 gnd.n3380 gnd.n3378 15.6674
R9673 gnd.n2906 gnd.t137 15.6146
R9674 gnd.t133 gnd.n2353 15.6146
R9675 gnd.t234 gnd.n2354 15.6146
R9676 gnd.n4178 gnd.t35 15.6146
R9677 gnd.t189 gnd.n2061 15.6146
R9678 gnd.n5543 gnd.t173 15.6146
R9679 gnd.n7324 gnd.t0 15.6146
R9680 gnd.n5899 gnd.n1502 15.3217
R9681 gnd.n7453 gnd.n313 15.3217
R9682 gnd.n3928 gnd.n2270 15.3217
R9683 gnd.n4533 gnd.n4426 15.3217
R9684 gnd.n4873 gnd.n1884 15.296
R9685 gnd.n4892 gnd.n1875 15.296
R9686 gnd.n4853 gnd.t81 15.296
R9687 gnd.n5023 gnd.n5021 15.296
R9688 gnd.n5068 gnd.n1780 15.296
R9689 gnd.n5195 gnd.t270 15.296
R9690 gnd.n5135 gnd.n1703 15.296
R9691 gnd.n5233 gnd.n1690 15.296
R9692 gnd.n1631 gnd.t152 15.296
R9693 gnd.n5572 gnd.n5571 15.0827
R9694 gnd.n1196 gnd.n1191 15.0481
R9695 gnd.n5582 gnd.n5581 15.0481
R9696 gnd.n3274 gnd.t108 14.9773
R9697 gnd.n4136 gnd.t43 14.9773
R9698 gnd.n6326 gnd.n1152 14.9773
R9699 gnd.n7385 gnd.t41 14.9773
R9700 gnd.n4733 gnd.t228 14.6587
R9701 gnd.n4800 gnd.n1906 14.6587
R9702 gnd.n4935 gnd.n4934 14.6587
R9703 gnd.n1731 gnd.n1720 14.6587
R9704 gnd.n5273 gnd.n5272 14.6587
R9705 gnd.t149 gnd.n1627 14.6587
R9706 gnd.n5320 gnd.n5319 14.6587
R9707 gnd.t297 gnd.n2396 14.34
R9708 gnd.n3352 gnd.t112 14.34
R9709 gnd.n4087 gnd.t56 14.34
R9710 gnd.t84 gnd.n173 14.34
R9711 gnd.n4758 gnd.t180 14.0214
R9712 gnd.n4808 gnd.n1891 14.0214
R9713 gnd.n4852 gnd.n1860 14.0214
R9714 gnd.n5013 gnd.n5012 14.0214
R9715 gnd.n1770 gnd.n1762 14.0214
R9716 gnd.n5196 gnd.n1707 14.0214
R9717 gnd.n1679 gnd.n1678 14.0214
R9718 gnd.n5564 gnd.n1578 14.0214
R9719 gnd.n3062 gnd.t114 13.7027
R9720 gnd.n1833 gnd.t94 13.7027
R9721 gnd.n5103 gnd.t253 13.7027
R9722 gnd.n2772 gnd.n2771 13.5763
R9723 gnd.n3716 gnd.n2310 13.5763
R9724 gnd.n2980 gnd.n2718 13.384
R9725 gnd.n4743 gnd.n1221 13.384
R9726 gnd.n4832 gnd.n1901 13.384
R9727 gnd.n1861 gnd.n1855 13.384
R9728 gnd.t307 gnd.n4922 13.384
R9729 gnd.n5174 gnd.t304 13.384
R9730 gnd.n5183 gnd.n1716 13.384
R9731 gnd.n5211 gnd.n1667 13.384
R9732 gnd.n5336 gnd.n1618 13.384
R9733 gnd.n1207 gnd.n1188 13.1884
R9734 gnd.n1202 gnd.n1201 13.1884
R9735 gnd.n1201 gnd.n1200 13.1884
R9736 gnd.n5575 gnd.n5570 13.1884
R9737 gnd.n5576 gnd.n5575 13.1884
R9738 gnd.n1203 gnd.n1190 13.146
R9739 gnd.n1199 gnd.n1190 13.146
R9740 gnd.n5574 gnd.n5573 13.146
R9741 gnd.n5574 gnd.n5569 13.146
R9742 gnd.n4774 gnd.t8 13.0654
R9743 gnd.n5294 gnd.t344 13.0654
R9744 gnd.n3603 gnd.n3599 12.8005
R9745 gnd.n3571 gnd.n3567 12.8005
R9746 gnd.n3539 gnd.n3535 12.8005
R9747 gnd.n3508 gnd.n3504 12.8005
R9748 gnd.n3476 gnd.n3472 12.8005
R9749 gnd.n3444 gnd.n3440 12.8005
R9750 gnd.n3412 gnd.n3408 12.8005
R9751 gnd.n3381 gnd.n3377 12.8005
R9752 gnd.n1937 gnd.n1223 12.7467
R9753 gnd.n4791 gnd.t207 12.7467
R9754 gnd.n4816 gnd.n4815 12.7467
R9755 gnd.n4983 gnd.n4981 12.7467
R9756 gnd.n5093 gnd.n1749 12.7467
R9757 gnd.n5259 gnd.n5258 12.7467
R9758 gnd.n2771 gnd.n2766 12.4126
R9759 gnd.n3719 gnd.n3716 12.4126
R9760 gnd.n6323 gnd.n6260 12.1761
R9761 gnd.n5651 gnd.n5650 12.1761
R9762 gnd.n6256 gnd.n1210 12.1094
R9763 gnd.t160 gnd.n1941 12.1094
R9764 gnd.n4823 gnd.n1892 12.1094
R9765 gnd.n4904 gnd.n1866 12.1094
R9766 gnd.n5203 gnd.n1701 12.1094
R9767 gnd.n5244 gnd.n1676 12.1094
R9768 gnd.n5344 gnd.n1581 12.1094
R9769 gnd.n3607 gnd.n3606 12.0247
R9770 gnd.n3575 gnd.n3574 12.0247
R9771 gnd.n3543 gnd.n3542 12.0247
R9772 gnd.n3512 gnd.n3511 12.0247
R9773 gnd.n3480 gnd.n3479 12.0247
R9774 gnd.n3448 gnd.n3447 12.0247
R9775 gnd.n3416 gnd.n3415 12.0247
R9776 gnd.n3385 gnd.n3384 12.0247
R9777 gnd.n4393 gnd.n1100 11.4721
R9778 gnd.n4784 gnd.n1923 11.4721
R9779 gnd.n4776 gnd.n4775 11.4721
R9780 gnd.n4943 gnd.t321 11.4721
R9781 gnd.n4942 gnd.n1842 11.4721
R9782 gnd.n4973 gnd.n4972 11.4721
R9783 gnd.n5120 gnd.n1744 11.4721
R9784 gnd.n5112 gnd.n1730 11.4721
R9785 gnd.n5164 gnd.t334 11.4721
R9786 gnd.n5284 gnd.n1654 11.4721
R9787 gnd.n5305 gnd.n5304 11.4721
R9788 gnd.n6129 gnd.n1329 11.4721
R9789 gnd.n7413 gnd.n207 11.4721
R9790 gnd.n3610 gnd.n3597 11.249
R9791 gnd.n3578 gnd.n3565 11.249
R9792 gnd.n3546 gnd.n3533 11.249
R9793 gnd.n3515 gnd.n3502 11.249
R9794 gnd.n3483 gnd.n3470 11.249
R9795 gnd.n3451 gnd.n3438 11.249
R9796 gnd.n3419 gnd.n3406 11.249
R9797 gnd.n3388 gnd.n3375 11.249
R9798 gnd.n3050 gnd.t114 11.1535
R9799 gnd.t35 gnd.n968 11.1535
R9800 gnd.n4721 gnd.t280 11.1535
R9801 gnd.n4920 gnd.t362 11.1535
R9802 gnd.t284 gnd.n5175 11.1535
R9803 gnd.t282 gnd.n5554 11.1535
R9804 gnd.t0 gnd.n102 11.1535
R9805 gnd.n4886 gnd.n4885 10.8348
R9806 gnd.n4885 gnd.n4884 10.8348
R9807 gnd.n5062 gnd.n5061 10.8348
R9808 gnd.n5061 gnd.n1777 10.8348
R9809 gnd.n5227 gnd.n5226 10.8348
R9810 gnd.n5226 gnd.n1687 10.8348
R9811 gnd.n1503 gnd.n1502 10.6672
R9812 gnd.n7458 gnd.n313 10.6672
R9813 gnd.n3930 gnd.n3928 10.6672
R9814 gnd.n4528 gnd.n4426 10.6672
R9815 gnd.n5716 gnd.n1532 10.6151
R9816 gnd.n5716 gnd.n5715 10.6151
R9817 gnd.n5713 gnd.n5710 10.6151
R9818 gnd.n5710 gnd.n5709 10.6151
R9819 gnd.n5709 gnd.n5706 10.6151
R9820 gnd.n5706 gnd.n5705 10.6151
R9821 gnd.n5705 gnd.n5702 10.6151
R9822 gnd.n5702 gnd.n5701 10.6151
R9823 gnd.n5701 gnd.n5698 10.6151
R9824 gnd.n5698 gnd.n5697 10.6151
R9825 gnd.n5697 gnd.n5694 10.6151
R9826 gnd.n5694 gnd.n5693 10.6151
R9827 gnd.n5693 gnd.n5690 10.6151
R9828 gnd.n5690 gnd.n5689 10.6151
R9829 gnd.n5689 gnd.n5686 10.6151
R9830 gnd.n5686 gnd.n5685 10.6151
R9831 gnd.n5685 gnd.n5682 10.6151
R9832 gnd.n5682 gnd.n5681 10.6151
R9833 gnd.n5681 gnd.n5678 10.6151
R9834 gnd.n5678 gnd.n5677 10.6151
R9835 gnd.n5677 gnd.n5674 10.6151
R9836 gnd.n5674 gnd.n5673 10.6151
R9837 gnd.n5673 gnd.n5670 10.6151
R9838 gnd.n5670 gnd.n5669 10.6151
R9839 gnd.n5669 gnd.n5666 10.6151
R9840 gnd.n5666 gnd.n5665 10.6151
R9841 gnd.n5665 gnd.n5662 10.6151
R9842 gnd.n5662 gnd.n5661 10.6151
R9843 gnd.n5661 gnd.n5658 10.6151
R9844 gnd.n5658 gnd.n5657 10.6151
R9845 gnd.n2024 gnd.n2023 10.6151
R9846 gnd.n2023 gnd.n2022 10.6151
R9847 gnd.n2022 gnd.n2019 10.6151
R9848 gnd.n2019 gnd.n2018 10.6151
R9849 gnd.n2018 gnd.n2015 10.6151
R9850 gnd.n2015 gnd.n2014 10.6151
R9851 gnd.n2014 gnd.n1920 10.6151
R9852 gnd.n4786 gnd.n1920 10.6151
R9853 gnd.n4787 gnd.n4786 10.6151
R9854 gnd.n4789 gnd.n4787 10.6151
R9855 gnd.n4789 gnd.n4788 10.6151
R9856 gnd.n4788 gnd.n1908 10.6151
R9857 gnd.n4802 gnd.n1908 10.6151
R9858 gnd.n4803 gnd.n4802 10.6151
R9859 gnd.n4813 gnd.n4803 10.6151
R9860 gnd.n4813 gnd.n4812 10.6151
R9861 gnd.n4812 gnd.n4811 10.6151
R9862 gnd.n4811 gnd.n4804 10.6151
R9863 gnd.n4805 gnd.n4804 10.6151
R9864 gnd.n4805 gnd.n1882 10.6151
R9865 gnd.n4875 gnd.n1882 10.6151
R9866 gnd.n4876 gnd.n4875 10.6151
R9867 gnd.n4882 gnd.n4876 10.6151
R9868 gnd.n4882 gnd.n4881 10.6151
R9869 gnd.n4881 gnd.n4880 10.6151
R9870 gnd.n4880 gnd.n4877 10.6151
R9871 gnd.n4877 gnd.n1858 10.6151
R9872 gnd.n4913 gnd.n1858 10.6151
R9873 gnd.n4914 gnd.n4913 10.6151
R9874 gnd.n4918 gnd.n4914 10.6151
R9875 gnd.n4918 gnd.n4917 10.6151
R9876 gnd.n4917 gnd.n4916 10.6151
R9877 gnd.n4916 gnd.n4915 10.6151
R9878 gnd.n4915 gnd.n1832 10.6151
R9879 gnd.n4961 gnd.n1832 10.6151
R9880 gnd.n4961 gnd.n4960 10.6151
R9881 gnd.n4960 gnd.n4959 10.6151
R9882 gnd.n4959 gnd.n4958 10.6151
R9883 gnd.n4958 gnd.n1814 10.6151
R9884 gnd.n4985 gnd.n1814 10.6151
R9885 gnd.n4986 gnd.n4985 10.6151
R9886 gnd.n4988 gnd.n4986 10.6151
R9887 gnd.n4989 gnd.n4988 10.6151
R9888 gnd.n4990 gnd.n4989 10.6151
R9889 gnd.n4990 gnd.n1791 10.6151
R9890 gnd.n5025 gnd.n1791 10.6151
R9891 gnd.n5026 gnd.n5025 10.6151
R9892 gnd.n5028 gnd.n5026 10.6151
R9893 gnd.n5029 gnd.n5028 10.6151
R9894 gnd.n5031 gnd.n5029 10.6151
R9895 gnd.n5031 gnd.n5030 10.6151
R9896 gnd.n5030 gnd.n1760 10.6151
R9897 gnd.n5088 gnd.n1760 10.6151
R9898 gnd.n5089 gnd.n5088 10.6151
R9899 gnd.n5091 gnd.n5089 10.6151
R9900 gnd.n5091 gnd.n5090 10.6151
R9901 gnd.n5090 gnd.n1741 10.6151
R9902 gnd.n5122 gnd.n1741 10.6151
R9903 gnd.n5123 gnd.n5122 10.6151
R9904 gnd.n5153 gnd.n5123 10.6151
R9905 gnd.n5153 gnd.n5152 10.6151
R9906 gnd.n5152 gnd.n5151 10.6151
R9907 gnd.n5151 gnd.n5148 10.6151
R9908 gnd.n5148 gnd.n5147 10.6151
R9909 gnd.n5147 gnd.n5146 10.6151
R9910 gnd.n5146 gnd.n5145 10.6151
R9911 gnd.n5145 gnd.n5144 10.6151
R9912 gnd.n5144 gnd.n5141 10.6151
R9913 gnd.n5141 gnd.n5140 10.6151
R9914 gnd.n5140 gnd.n5138 10.6151
R9915 gnd.n5138 gnd.n5137 10.6151
R9916 gnd.n5137 gnd.n5131 10.6151
R9917 gnd.n5131 gnd.n5130 10.6151
R9918 gnd.n5130 gnd.n5128 10.6151
R9919 gnd.n5128 gnd.n5127 10.6151
R9920 gnd.n5127 gnd.n5124 10.6151
R9921 gnd.n5124 gnd.n1670 10.6151
R9922 gnd.n5253 gnd.n1670 10.6151
R9923 gnd.n5254 gnd.n5253 10.6151
R9924 gnd.n5256 gnd.n5254 10.6151
R9925 gnd.n5256 gnd.n5255 10.6151
R9926 gnd.n5255 gnd.n1650 10.6151
R9927 gnd.n5286 gnd.n1650 10.6151
R9928 gnd.n5287 gnd.n5286 10.6151
R9929 gnd.n5291 gnd.n5287 10.6151
R9930 gnd.n5291 gnd.n5290 10.6151
R9931 gnd.n5290 gnd.n5289 10.6151
R9932 gnd.n5289 gnd.n5288 10.6151
R9933 gnd.n5288 gnd.n1620 10.6151
R9934 gnd.n5329 gnd.n1620 10.6151
R9935 gnd.n5330 gnd.n5329 10.6151
R9936 gnd.n5333 gnd.n5330 10.6151
R9937 gnd.n5333 gnd.n5332 10.6151
R9938 gnd.n5332 gnd.n5331 10.6151
R9939 gnd.n5331 gnd.n1571 10.6151
R9940 gnd.n1952 gnd.n1148 10.6151
R9941 gnd.n1955 gnd.n1952 10.6151
R9942 gnd.n1960 gnd.n1957 10.6151
R9943 gnd.n1961 gnd.n1960 10.6151
R9944 gnd.n1964 gnd.n1961 10.6151
R9945 gnd.n1965 gnd.n1964 10.6151
R9946 gnd.n1968 gnd.n1965 10.6151
R9947 gnd.n1969 gnd.n1968 10.6151
R9948 gnd.n1972 gnd.n1969 10.6151
R9949 gnd.n1973 gnd.n1972 10.6151
R9950 gnd.n1976 gnd.n1973 10.6151
R9951 gnd.n1977 gnd.n1976 10.6151
R9952 gnd.n1980 gnd.n1977 10.6151
R9953 gnd.n1981 gnd.n1980 10.6151
R9954 gnd.n1984 gnd.n1981 10.6151
R9955 gnd.n1985 gnd.n1984 10.6151
R9956 gnd.n1988 gnd.n1985 10.6151
R9957 gnd.n1989 gnd.n1988 10.6151
R9958 gnd.n1992 gnd.n1989 10.6151
R9959 gnd.n1993 gnd.n1992 10.6151
R9960 gnd.n1996 gnd.n1993 10.6151
R9961 gnd.n1997 gnd.n1996 10.6151
R9962 gnd.n2000 gnd.n1997 10.6151
R9963 gnd.n2001 gnd.n2000 10.6151
R9964 gnd.n2004 gnd.n2001 10.6151
R9965 gnd.n2005 gnd.n2004 10.6151
R9966 gnd.n2008 gnd.n2005 10.6151
R9967 gnd.n2009 gnd.n2008 10.6151
R9968 gnd.n2012 gnd.n2009 10.6151
R9969 gnd.n2013 gnd.n2012 10.6151
R9970 gnd.n6323 gnd.n6322 10.6151
R9971 gnd.n6322 gnd.n6321 10.6151
R9972 gnd.n6321 gnd.n6320 10.6151
R9973 gnd.n6320 gnd.n6318 10.6151
R9974 gnd.n6318 gnd.n6315 10.6151
R9975 gnd.n6315 gnd.n6314 10.6151
R9976 gnd.n6314 gnd.n6311 10.6151
R9977 gnd.n6311 gnd.n6310 10.6151
R9978 gnd.n6310 gnd.n6307 10.6151
R9979 gnd.n6307 gnd.n6306 10.6151
R9980 gnd.n6306 gnd.n6303 10.6151
R9981 gnd.n6303 gnd.n6302 10.6151
R9982 gnd.n6302 gnd.n6299 10.6151
R9983 gnd.n6299 gnd.n6298 10.6151
R9984 gnd.n6298 gnd.n6295 10.6151
R9985 gnd.n6295 gnd.n6294 10.6151
R9986 gnd.n6294 gnd.n6291 10.6151
R9987 gnd.n6291 gnd.n6290 10.6151
R9988 gnd.n6290 gnd.n6287 10.6151
R9989 gnd.n6287 gnd.n6286 10.6151
R9990 gnd.n6286 gnd.n6283 10.6151
R9991 gnd.n6283 gnd.n6282 10.6151
R9992 gnd.n6282 gnd.n6279 10.6151
R9993 gnd.n6279 gnd.n6278 10.6151
R9994 gnd.n6278 gnd.n6275 10.6151
R9995 gnd.n6275 gnd.n6274 10.6151
R9996 gnd.n6274 gnd.n6271 10.6151
R9997 gnd.n6271 gnd.n6270 10.6151
R9998 gnd.n6267 gnd.n6266 10.6151
R9999 gnd.n6266 gnd.n1149 10.6151
R10000 gnd.n5650 gnd.n5649 10.6151
R10001 gnd.n5649 gnd.n5646 10.6151
R10002 gnd.n5646 gnd.n5645 10.6151
R10003 gnd.n5645 gnd.n5642 10.6151
R10004 gnd.n5642 gnd.n5641 10.6151
R10005 gnd.n5641 gnd.n5638 10.6151
R10006 gnd.n5638 gnd.n5637 10.6151
R10007 gnd.n5637 gnd.n5634 10.6151
R10008 gnd.n5634 gnd.n5633 10.6151
R10009 gnd.n5633 gnd.n5630 10.6151
R10010 gnd.n5630 gnd.n5629 10.6151
R10011 gnd.n5629 gnd.n5626 10.6151
R10012 gnd.n5626 gnd.n5625 10.6151
R10013 gnd.n5625 gnd.n5622 10.6151
R10014 gnd.n5622 gnd.n5621 10.6151
R10015 gnd.n5621 gnd.n5618 10.6151
R10016 gnd.n5618 gnd.n5617 10.6151
R10017 gnd.n5617 gnd.n5614 10.6151
R10018 gnd.n5614 gnd.n5613 10.6151
R10019 gnd.n5613 gnd.n5610 10.6151
R10020 gnd.n5610 gnd.n5609 10.6151
R10021 gnd.n5609 gnd.n5606 10.6151
R10022 gnd.n5606 gnd.n5605 10.6151
R10023 gnd.n5605 gnd.n5602 10.6151
R10024 gnd.n5602 gnd.n5601 10.6151
R10025 gnd.n5601 gnd.n5598 10.6151
R10026 gnd.n5598 gnd.n5597 10.6151
R10027 gnd.n5597 gnd.n5594 10.6151
R10028 gnd.n5592 gnd.n5589 10.6151
R10029 gnd.n5589 gnd.n1533 10.6151
R10030 gnd.n6259 gnd.n6258 10.6151
R10031 gnd.n6258 gnd.n1208 10.6151
R10032 gnd.n1940 gnd.n1208 10.6151
R10033 gnd.n4747 gnd.n1940 10.6151
R10034 gnd.n4748 gnd.n4747 10.6151
R10035 gnd.n4749 gnd.n4748 10.6151
R10036 gnd.n4749 gnd.n1926 10.6151
R10037 gnd.n4782 gnd.n1926 10.6151
R10038 gnd.n4782 gnd.n4781 10.6151
R10039 gnd.n4781 gnd.n4780 10.6151
R10040 gnd.n4780 gnd.n4779 10.6151
R10041 gnd.n4779 gnd.n1927 10.6151
R10042 gnd.n1927 gnd.n1904 10.6151
R10043 gnd.n4819 gnd.n1904 10.6151
R10044 gnd.n4820 gnd.n4819 10.6151
R10045 gnd.n4830 gnd.n4820 10.6151
R10046 gnd.n4830 gnd.n4829 10.6151
R10047 gnd.n4829 gnd.n4828 10.6151
R10048 gnd.n4828 gnd.n4821 10.6151
R10049 gnd.n4822 gnd.n4821 10.6151
R10050 gnd.n4822 gnd.n1877 10.6151
R10051 gnd.n4888 gnd.n1877 10.6151
R10052 gnd.n4889 gnd.n4888 10.6151
R10053 gnd.n4890 gnd.n4889 10.6151
R10054 gnd.n4890 gnd.n1864 10.6151
R10055 gnd.n4906 gnd.n1864 10.6151
R10056 gnd.n4907 gnd.n4906 10.6151
R10057 gnd.n4909 gnd.n4907 10.6151
R10058 gnd.n4909 gnd.n4908 10.6151
R10059 gnd.n4908 gnd.n1844 10.6151
R10060 gnd.n4938 gnd.n1844 10.6151
R10061 gnd.n4939 gnd.n4938 10.6151
R10062 gnd.n4940 gnd.n4939 10.6151
R10063 gnd.n4940 gnd.n1827 10.6151
R10064 gnd.n4965 gnd.n1827 10.6151
R10065 gnd.n4966 gnd.n4965 10.6151
R10066 gnd.n4970 gnd.n4966 10.6151
R10067 gnd.n4970 gnd.n4969 10.6151
R10068 gnd.n4969 gnd.n4968 10.6151
R10069 gnd.n4968 gnd.n1804 10.6151
R10070 gnd.n5005 gnd.n1804 10.6151
R10071 gnd.n5006 gnd.n5005 10.6151
R10072 gnd.n5010 gnd.n5006 10.6151
R10073 gnd.n5010 gnd.n5009 10.6151
R10074 gnd.n5009 gnd.n5008 10.6151
R10075 gnd.n5008 gnd.n1782 10.6151
R10076 gnd.n5064 gnd.n1782 10.6151
R10077 gnd.n5065 gnd.n5064 10.6151
R10078 gnd.n5066 gnd.n5065 10.6151
R10079 gnd.n5066 gnd.n1767 10.6151
R10080 gnd.n5081 gnd.n1767 10.6151
R10081 gnd.n5082 gnd.n5081 10.6151
R10082 gnd.n5084 gnd.n5082 10.6151
R10083 gnd.n5084 gnd.n5083 10.6151
R10084 gnd.n5083 gnd.n1747 10.6151
R10085 gnd.n5108 gnd.n1747 10.6151
R10086 gnd.n5109 gnd.n5108 10.6151
R10087 gnd.n5118 gnd.n5109 10.6151
R10088 gnd.n5118 gnd.n5117 10.6151
R10089 gnd.n5117 gnd.n5116 10.6151
R10090 gnd.n5116 gnd.n5115 10.6151
R10091 gnd.n5115 gnd.n5110 10.6151
R10092 gnd.n5110 gnd.n1718 10.6151
R10093 gnd.n5179 gnd.n1718 10.6151
R10094 gnd.n5180 gnd.n5179 10.6151
R10095 gnd.n5181 gnd.n5180 10.6151
R10096 gnd.n5181 gnd.n1705 10.6151
R10097 gnd.n5198 gnd.n1705 10.6151
R10098 gnd.n5199 gnd.n5198 10.6151
R10099 gnd.n5200 gnd.n5199 10.6151
R10100 gnd.n5200 gnd.n1692 10.6151
R10101 gnd.n5229 gnd.n1692 10.6151
R10102 gnd.n5230 gnd.n5229 10.6151
R10103 gnd.n5231 gnd.n5230 10.6151
R10104 gnd.n5231 gnd.n1674 10.6151
R10105 gnd.n5246 gnd.n1674 10.6151
R10106 gnd.n5247 gnd.n5246 10.6151
R10107 gnd.n5249 gnd.n5247 10.6151
R10108 gnd.n5249 gnd.n5248 10.6151
R10109 gnd.n5248 gnd.n1657 10.6151
R10110 gnd.n5276 gnd.n1657 10.6151
R10111 gnd.n5277 gnd.n5276 10.6151
R10112 gnd.n5282 gnd.n5277 10.6151
R10113 gnd.n5282 gnd.n5281 10.6151
R10114 gnd.n5281 gnd.n5280 10.6151
R10115 gnd.n5280 gnd.n5279 10.6151
R10116 gnd.n5279 gnd.n1625 10.6151
R10117 gnd.n5322 gnd.n1625 10.6151
R10118 gnd.n5323 gnd.n5322 10.6151
R10119 gnd.n5325 gnd.n5323 10.6151
R10120 gnd.n5325 gnd.n5324 10.6151
R10121 gnd.n5324 gnd.n1576 10.6151
R10122 gnd.n5566 gnd.n1576 10.6151
R10123 gnd.n5567 gnd.n5566 10.6151
R10124 gnd.n5652 gnd.n5567 10.6151
R10125 gnd.n2969 gnd.t92 10.5161
R10126 gnd.n2398 gnd.t297 10.5161
R10127 gnd.n3335 gnd.t112 10.5161
R10128 gnd.n4278 gnd.t26 10.5161
R10129 gnd.n4895 gnd.t292 10.5161
R10130 gnd.t28 gnd.n5132 10.5161
R10131 gnd.n1458 gnd.t116 10.5161
R10132 gnd.n3611 gnd.n3595 10.4732
R10133 gnd.n3579 gnd.n3563 10.4732
R10134 gnd.n3547 gnd.n3531 10.4732
R10135 gnd.n3516 gnd.n3500 10.4732
R10136 gnd.n3484 gnd.n3468 10.4732
R10137 gnd.n3452 gnd.n3436 10.4732
R10138 gnd.n3420 gnd.n3404 10.4732
R10139 gnd.n3389 gnd.n3373 10.4732
R10140 gnd.n1929 gnd.n1923 10.1975
R10141 gnd.n1842 gnd.n1841 10.1975
R10142 gnd.n4973 gnd.n1822 10.1975
R10143 gnd.n5041 gnd.n1744 10.1975
R10144 gnd.n5113 gnd.n5112 10.1975
R10145 gnd.n5305 gnd.n1637 10.1975
R10146 gnd.n1590 gnd.t177 10.1975
R10147 gnd.t108 gnd.n2415 9.87883
R10148 gnd.n4315 gnd.t70 9.87883
R10149 gnd.n1475 gnd.t37 9.87883
R10150 gnd.n3615 gnd.n3614 9.69747
R10151 gnd.n3583 gnd.n3582 9.69747
R10152 gnd.n3551 gnd.n3550 9.69747
R10153 gnd.n3520 gnd.n3519 9.69747
R10154 gnd.n3488 gnd.n3487 9.69747
R10155 gnd.n3456 gnd.n3455 9.69747
R10156 gnd.n3424 gnd.n3423 9.69747
R10157 gnd.n3393 gnd.n3392 9.69747
R10158 gnd.n2026 gnd.n1210 9.56018
R10159 gnd.n4824 gnd.n4823 9.56018
R10160 gnd.n4878 gnd.n1866 9.56018
R10161 gnd.n4947 gnd.t82 9.56018
R10162 gnd.n4993 gnd.n1793 9.56018
R10163 gnd.n5034 gnd.n5033 9.56018
R10164 gnd.n5043 gnd.t52 9.56018
R10165 gnd.n5203 gnd.n5202 9.56018
R10166 gnd.n5125 gnd.n1676 9.56018
R10167 gnd.n3621 gnd.n3620 9.45567
R10168 gnd.n3589 gnd.n3588 9.45567
R10169 gnd.n3557 gnd.n3556 9.45567
R10170 gnd.n3526 gnd.n3525 9.45567
R10171 gnd.n3494 gnd.n3493 9.45567
R10172 gnd.n3462 gnd.n3461 9.45567
R10173 gnd.n3430 gnd.n3429 9.45567
R10174 gnd.n3399 gnd.n3398 9.45567
R10175 gnd.n5847 gnd.n1521 9.30959
R10176 gnd.n7492 gnd.n277 9.30959
R10177 gnd.n3967 gnd.n3966 9.30959
R10178 gnd.n4484 gnd.n4448 9.30959
R10179 gnd.n3620 gnd.n3619 9.3005
R10180 gnd.n3593 gnd.n3592 9.3005
R10181 gnd.n3614 gnd.n3613 9.3005
R10182 gnd.n3612 gnd.n3611 9.3005
R10183 gnd.n3597 gnd.n3596 9.3005
R10184 gnd.n3606 gnd.n3605 9.3005
R10185 gnd.n3604 gnd.n3603 9.3005
R10186 gnd.n3588 gnd.n3587 9.3005
R10187 gnd.n3561 gnd.n3560 9.3005
R10188 gnd.n3582 gnd.n3581 9.3005
R10189 gnd.n3580 gnd.n3579 9.3005
R10190 gnd.n3565 gnd.n3564 9.3005
R10191 gnd.n3574 gnd.n3573 9.3005
R10192 gnd.n3572 gnd.n3571 9.3005
R10193 gnd.n3556 gnd.n3555 9.3005
R10194 gnd.n3529 gnd.n3528 9.3005
R10195 gnd.n3550 gnd.n3549 9.3005
R10196 gnd.n3548 gnd.n3547 9.3005
R10197 gnd.n3533 gnd.n3532 9.3005
R10198 gnd.n3542 gnd.n3541 9.3005
R10199 gnd.n3540 gnd.n3539 9.3005
R10200 gnd.n3525 gnd.n3524 9.3005
R10201 gnd.n3498 gnd.n3497 9.3005
R10202 gnd.n3519 gnd.n3518 9.3005
R10203 gnd.n3517 gnd.n3516 9.3005
R10204 gnd.n3502 gnd.n3501 9.3005
R10205 gnd.n3511 gnd.n3510 9.3005
R10206 gnd.n3509 gnd.n3508 9.3005
R10207 gnd.n3493 gnd.n3492 9.3005
R10208 gnd.n3466 gnd.n3465 9.3005
R10209 gnd.n3487 gnd.n3486 9.3005
R10210 gnd.n3485 gnd.n3484 9.3005
R10211 gnd.n3470 gnd.n3469 9.3005
R10212 gnd.n3479 gnd.n3478 9.3005
R10213 gnd.n3477 gnd.n3476 9.3005
R10214 gnd.n3461 gnd.n3460 9.3005
R10215 gnd.n3434 gnd.n3433 9.3005
R10216 gnd.n3455 gnd.n3454 9.3005
R10217 gnd.n3453 gnd.n3452 9.3005
R10218 gnd.n3438 gnd.n3437 9.3005
R10219 gnd.n3447 gnd.n3446 9.3005
R10220 gnd.n3445 gnd.n3444 9.3005
R10221 gnd.n3429 gnd.n3428 9.3005
R10222 gnd.n3402 gnd.n3401 9.3005
R10223 gnd.n3423 gnd.n3422 9.3005
R10224 gnd.n3421 gnd.n3420 9.3005
R10225 gnd.n3406 gnd.n3405 9.3005
R10226 gnd.n3415 gnd.n3414 9.3005
R10227 gnd.n3413 gnd.n3412 9.3005
R10228 gnd.n3398 gnd.n3397 9.3005
R10229 gnd.n3371 gnd.n3370 9.3005
R10230 gnd.n3392 gnd.n3391 9.3005
R10231 gnd.n3390 gnd.n3389 9.3005
R10232 gnd.n3375 gnd.n3374 9.3005
R10233 gnd.n3384 gnd.n3383 9.3005
R10234 gnd.n3382 gnd.n3381 9.3005
R10235 gnd.n3746 gnd.n3745 9.3005
R10236 gnd.n3744 gnd.n2298 9.3005
R10237 gnd.n3743 gnd.n3742 9.3005
R10238 gnd.n3739 gnd.n2299 9.3005
R10239 gnd.n3736 gnd.n2300 9.3005
R10240 gnd.n3735 gnd.n2301 9.3005
R10241 gnd.n3732 gnd.n2302 9.3005
R10242 gnd.n3731 gnd.n2303 9.3005
R10243 gnd.n3728 gnd.n2304 9.3005
R10244 gnd.n3727 gnd.n2305 9.3005
R10245 gnd.n3724 gnd.n2306 9.3005
R10246 gnd.n3723 gnd.n2307 9.3005
R10247 gnd.n3720 gnd.n2308 9.3005
R10248 gnd.n3719 gnd.n2309 9.3005
R10249 gnd.n3716 gnd.n3715 9.3005
R10250 gnd.n3714 gnd.n2310 9.3005
R10251 gnd.n3747 gnd.n2297 9.3005
R10252 gnd.n2988 gnd.n2987 9.3005
R10253 gnd.n2692 gnd.n2691 9.3005
R10254 gnd.n3015 gnd.n3014 9.3005
R10255 gnd.n3016 gnd.n2690 9.3005
R10256 gnd.n3020 gnd.n3017 9.3005
R10257 gnd.n3019 gnd.n3018 9.3005
R10258 gnd.n2664 gnd.n2663 9.3005
R10259 gnd.n3045 gnd.n3044 9.3005
R10260 gnd.n3046 gnd.n2662 9.3005
R10261 gnd.n3048 gnd.n3047 9.3005
R10262 gnd.n2642 gnd.n2641 9.3005
R10263 gnd.n3076 gnd.n3075 9.3005
R10264 gnd.n3077 gnd.n2640 9.3005
R10265 gnd.n3085 gnd.n3078 9.3005
R10266 gnd.n3084 gnd.n3079 9.3005
R10267 gnd.n3083 gnd.n3081 9.3005
R10268 gnd.n3080 gnd.n2589 9.3005
R10269 gnd.n3133 gnd.n2590 9.3005
R10270 gnd.n3132 gnd.n2591 9.3005
R10271 gnd.n3131 gnd.n2592 9.3005
R10272 gnd.n2611 gnd.n2593 9.3005
R10273 gnd.n2613 gnd.n2612 9.3005
R10274 gnd.n2495 gnd.n2494 9.3005
R10275 gnd.n3171 gnd.n3170 9.3005
R10276 gnd.n3172 gnd.n2493 9.3005
R10277 gnd.n3176 gnd.n3173 9.3005
R10278 gnd.n3175 gnd.n3174 9.3005
R10279 gnd.n2468 gnd.n2467 9.3005
R10280 gnd.n3211 gnd.n3210 9.3005
R10281 gnd.n3212 gnd.n2466 9.3005
R10282 gnd.n3216 gnd.n3213 9.3005
R10283 gnd.n3215 gnd.n3214 9.3005
R10284 gnd.n2441 gnd.n2440 9.3005
R10285 gnd.n3256 gnd.n3255 9.3005
R10286 gnd.n3257 gnd.n2439 9.3005
R10287 gnd.n3261 gnd.n3258 9.3005
R10288 gnd.n3260 gnd.n3259 9.3005
R10289 gnd.n2413 gnd.n2412 9.3005
R10290 gnd.n3296 gnd.n3295 9.3005
R10291 gnd.n3297 gnd.n2411 9.3005
R10292 gnd.n3301 gnd.n3298 9.3005
R10293 gnd.n3300 gnd.n3299 9.3005
R10294 gnd.n2386 gnd.n2385 9.3005
R10295 gnd.n3345 gnd.n3344 9.3005
R10296 gnd.n3346 gnd.n2384 9.3005
R10297 gnd.n3350 gnd.n3347 9.3005
R10298 gnd.n3349 gnd.n3348 9.3005
R10299 gnd.n2359 gnd.n2358 9.3005
R10300 gnd.n3639 gnd.n3638 9.3005
R10301 gnd.n3640 gnd.n2357 9.3005
R10302 gnd.n3646 gnd.n3641 9.3005
R10303 gnd.n3645 gnd.n3642 9.3005
R10304 gnd.n3644 gnd.n3643 9.3005
R10305 gnd.n2989 gnd.n2986 9.3005
R10306 gnd.n2771 gnd.n2730 9.3005
R10307 gnd.n2766 gnd.n2765 9.3005
R10308 gnd.n2764 gnd.n2731 9.3005
R10309 gnd.n2763 gnd.n2762 9.3005
R10310 gnd.n2759 gnd.n2732 9.3005
R10311 gnd.n2756 gnd.n2755 9.3005
R10312 gnd.n2754 gnd.n2733 9.3005
R10313 gnd.n2753 gnd.n2752 9.3005
R10314 gnd.n2749 gnd.n2734 9.3005
R10315 gnd.n2746 gnd.n2745 9.3005
R10316 gnd.n2744 gnd.n2735 9.3005
R10317 gnd.n2743 gnd.n2742 9.3005
R10318 gnd.n2739 gnd.n2737 9.3005
R10319 gnd.n2736 gnd.n2716 9.3005
R10320 gnd.n2983 gnd.n2715 9.3005
R10321 gnd.n2985 gnd.n2984 9.3005
R10322 gnd.n2773 gnd.n2772 9.3005
R10323 gnd.n2996 gnd.n2702 9.3005
R10324 gnd.n3003 gnd.n2703 9.3005
R10325 gnd.n3005 gnd.n3004 9.3005
R10326 gnd.n3006 gnd.n2683 9.3005
R10327 gnd.n3025 gnd.n3024 9.3005
R10328 gnd.n3027 gnd.n2675 9.3005
R10329 gnd.n3034 gnd.n2677 9.3005
R10330 gnd.n3035 gnd.n2672 9.3005
R10331 gnd.n3037 gnd.n3036 9.3005
R10332 gnd.n2673 gnd.n2658 9.3005
R10333 gnd.n3053 gnd.n2656 9.3005
R10334 gnd.n3057 gnd.n3056 9.3005
R10335 gnd.n3055 gnd.n2632 9.3005
R10336 gnd.n3092 gnd.n2631 9.3005
R10337 gnd.n3095 gnd.n3094 9.3005
R10338 gnd.n2628 gnd.n2627 9.3005
R10339 gnd.n3101 gnd.n2629 9.3005
R10340 gnd.n3103 gnd.n3102 9.3005
R10341 gnd.n3105 gnd.n2626 9.3005
R10342 gnd.n3108 gnd.n3107 9.3005
R10343 gnd.n3111 gnd.n3109 9.3005
R10344 gnd.n3113 gnd.n3112 9.3005
R10345 gnd.n3119 gnd.n3114 9.3005
R10346 gnd.n3118 gnd.n3117 9.3005
R10347 gnd.n2486 gnd.n2485 9.3005
R10348 gnd.n3185 gnd.n3184 9.3005
R10349 gnd.n3186 gnd.n2479 9.3005
R10350 gnd.n3194 gnd.n2478 9.3005
R10351 gnd.n3197 gnd.n3196 9.3005
R10352 gnd.n3199 gnd.n3198 9.3005
R10353 gnd.n3202 gnd.n2461 9.3005
R10354 gnd.n3200 gnd.n2459 9.3005
R10355 gnd.n3222 gnd.n2457 9.3005
R10356 gnd.n3224 gnd.n3223 9.3005
R10357 gnd.n2431 gnd.n2430 9.3005
R10358 gnd.n3270 gnd.n3269 9.3005
R10359 gnd.n3271 gnd.n2424 9.3005
R10360 gnd.n3279 gnd.n2423 9.3005
R10361 gnd.n3282 gnd.n3281 9.3005
R10362 gnd.n3284 gnd.n3283 9.3005
R10363 gnd.n3287 gnd.n2406 9.3005
R10364 gnd.n3285 gnd.n2404 9.3005
R10365 gnd.n3307 gnd.n2402 9.3005
R10366 gnd.n3309 gnd.n3308 9.3005
R10367 gnd.n2377 gnd.n2376 9.3005
R10368 gnd.n3359 gnd.n3358 9.3005
R10369 gnd.n3360 gnd.n2370 9.3005
R10370 gnd.n3368 gnd.n2369 9.3005
R10371 gnd.n3627 gnd.n3626 9.3005
R10372 gnd.n3629 gnd.n3628 9.3005
R10373 gnd.n3630 gnd.n2350 9.3005
R10374 gnd.n3654 gnd.n3653 9.3005
R10375 gnd.n2351 gnd.n2313 9.3005
R10376 gnd.n2994 gnd.n2993 9.3005
R10377 gnd.n3710 gnd.n2314 9.3005
R10378 gnd.n3709 gnd.n2316 9.3005
R10379 gnd.n3706 gnd.n2317 9.3005
R10380 gnd.n3705 gnd.n2318 9.3005
R10381 gnd.n3702 gnd.n2319 9.3005
R10382 gnd.n3701 gnd.n2320 9.3005
R10383 gnd.n3698 gnd.n2321 9.3005
R10384 gnd.n3697 gnd.n2322 9.3005
R10385 gnd.n3694 gnd.n2323 9.3005
R10386 gnd.n3693 gnd.n2324 9.3005
R10387 gnd.n3690 gnd.n2325 9.3005
R10388 gnd.n3689 gnd.n2326 9.3005
R10389 gnd.n3686 gnd.n2327 9.3005
R10390 gnd.n3685 gnd.n2328 9.3005
R10391 gnd.n3682 gnd.n2329 9.3005
R10392 gnd.n3681 gnd.n2330 9.3005
R10393 gnd.n3678 gnd.n2331 9.3005
R10394 gnd.n3677 gnd.n2332 9.3005
R10395 gnd.n3674 gnd.n2333 9.3005
R10396 gnd.n3673 gnd.n2334 9.3005
R10397 gnd.n3670 gnd.n2335 9.3005
R10398 gnd.n3669 gnd.n2336 9.3005
R10399 gnd.n3666 gnd.n2340 9.3005
R10400 gnd.n3665 gnd.n2341 9.3005
R10401 gnd.n3662 gnd.n2342 9.3005
R10402 gnd.n3661 gnd.n2343 9.3005
R10403 gnd.n3712 gnd.n3711 9.3005
R10404 gnd.n3163 gnd.n3147 9.3005
R10405 gnd.n3162 gnd.n3148 9.3005
R10406 gnd.n3161 gnd.n3149 9.3005
R10407 gnd.n3159 gnd.n3150 9.3005
R10408 gnd.n3158 gnd.n3151 9.3005
R10409 gnd.n3156 gnd.n3152 9.3005
R10410 gnd.n3155 gnd.n3153 9.3005
R10411 gnd.n2449 gnd.n2448 9.3005
R10412 gnd.n3232 gnd.n3231 9.3005
R10413 gnd.n3233 gnd.n2447 9.3005
R10414 gnd.n3250 gnd.n3234 9.3005
R10415 gnd.n3249 gnd.n3235 9.3005
R10416 gnd.n3248 gnd.n3236 9.3005
R10417 gnd.n3246 gnd.n3237 9.3005
R10418 gnd.n3245 gnd.n3238 9.3005
R10419 gnd.n3243 gnd.n3239 9.3005
R10420 gnd.n3242 gnd.n3240 9.3005
R10421 gnd.n2393 gnd.n2392 9.3005
R10422 gnd.n3317 gnd.n3316 9.3005
R10423 gnd.n3318 gnd.n2391 9.3005
R10424 gnd.n3339 gnd.n3319 9.3005
R10425 gnd.n3338 gnd.n3320 9.3005
R10426 gnd.n3337 gnd.n3321 9.3005
R10427 gnd.n3334 gnd.n3322 9.3005
R10428 gnd.n3333 gnd.n3323 9.3005
R10429 gnd.n3331 gnd.n3324 9.3005
R10430 gnd.n3330 gnd.n3325 9.3005
R10431 gnd.n3328 gnd.n3327 9.3005
R10432 gnd.n3326 gnd.n2345 9.3005
R10433 gnd.n2904 gnd.n2903 9.3005
R10434 gnd.n2794 gnd.n2793 9.3005
R10435 gnd.n2918 gnd.n2917 9.3005
R10436 gnd.n2919 gnd.n2792 9.3005
R10437 gnd.n2921 gnd.n2920 9.3005
R10438 gnd.n2782 gnd.n2781 9.3005
R10439 gnd.n2934 gnd.n2933 9.3005
R10440 gnd.n2935 gnd.n2780 9.3005
R10441 gnd.n2967 gnd.n2936 9.3005
R10442 gnd.n2966 gnd.n2937 9.3005
R10443 gnd.n2965 gnd.n2938 9.3005
R10444 gnd.n2964 gnd.n2939 9.3005
R10445 gnd.n2961 gnd.n2940 9.3005
R10446 gnd.n2960 gnd.n2941 9.3005
R10447 gnd.n2959 gnd.n2942 9.3005
R10448 gnd.n2957 gnd.n2943 9.3005
R10449 gnd.n2956 gnd.n2944 9.3005
R10450 gnd.n2953 gnd.n2945 9.3005
R10451 gnd.n2952 gnd.n2946 9.3005
R10452 gnd.n2951 gnd.n2947 9.3005
R10453 gnd.n2949 gnd.n2948 9.3005
R10454 gnd.n2648 gnd.n2647 9.3005
R10455 gnd.n3065 gnd.n3064 9.3005
R10456 gnd.n3066 gnd.n2646 9.3005
R10457 gnd.n3070 gnd.n3067 9.3005
R10458 gnd.n3069 gnd.n3068 9.3005
R10459 gnd.n2570 gnd.n2569 9.3005
R10460 gnd.n3145 gnd.n3144 9.3005
R10461 gnd.n2902 gnd.n2803 9.3005
R10462 gnd.n2805 gnd.n2804 9.3005
R10463 gnd.n2849 gnd.n2847 9.3005
R10464 gnd.n2850 gnd.n2846 9.3005
R10465 gnd.n2853 gnd.n2842 9.3005
R10466 gnd.n2854 gnd.n2841 9.3005
R10467 gnd.n2857 gnd.n2840 9.3005
R10468 gnd.n2858 gnd.n2839 9.3005
R10469 gnd.n2861 gnd.n2838 9.3005
R10470 gnd.n2862 gnd.n2837 9.3005
R10471 gnd.n2865 gnd.n2836 9.3005
R10472 gnd.n2866 gnd.n2835 9.3005
R10473 gnd.n2869 gnd.n2834 9.3005
R10474 gnd.n2870 gnd.n2833 9.3005
R10475 gnd.n2873 gnd.n2832 9.3005
R10476 gnd.n2874 gnd.n2831 9.3005
R10477 gnd.n2877 gnd.n2830 9.3005
R10478 gnd.n2878 gnd.n2829 9.3005
R10479 gnd.n2881 gnd.n2828 9.3005
R10480 gnd.n2882 gnd.n2827 9.3005
R10481 gnd.n2885 gnd.n2826 9.3005
R10482 gnd.n2886 gnd.n2825 9.3005
R10483 gnd.n2889 gnd.n2824 9.3005
R10484 gnd.n2891 gnd.n2823 9.3005
R10485 gnd.n2892 gnd.n2822 9.3005
R10486 gnd.n2893 gnd.n2821 9.3005
R10487 gnd.n2894 gnd.n2820 9.3005
R10488 gnd.n2901 gnd.n2900 9.3005
R10489 gnd.n2910 gnd.n2909 9.3005
R10490 gnd.n2911 gnd.n2797 9.3005
R10491 gnd.n2913 gnd.n2912 9.3005
R10492 gnd.n2788 gnd.n2787 9.3005
R10493 gnd.n2926 gnd.n2925 9.3005
R10494 gnd.n2927 gnd.n2786 9.3005
R10495 gnd.n2929 gnd.n2928 9.3005
R10496 gnd.n2775 gnd.n2774 9.3005
R10497 gnd.n2972 gnd.n2971 9.3005
R10498 gnd.n2973 gnd.n2729 9.3005
R10499 gnd.n2977 gnd.n2975 9.3005
R10500 gnd.n2976 gnd.n2708 9.3005
R10501 gnd.n2995 gnd.n2707 9.3005
R10502 gnd.n2998 gnd.n2997 9.3005
R10503 gnd.n2701 gnd.n2700 9.3005
R10504 gnd.n3009 gnd.n3007 9.3005
R10505 gnd.n3008 gnd.n2682 9.3005
R10506 gnd.n3026 gnd.n2681 9.3005
R10507 gnd.n3029 gnd.n3028 9.3005
R10508 gnd.n2676 gnd.n2671 9.3005
R10509 gnd.n3039 gnd.n3038 9.3005
R10510 gnd.n2674 gnd.n2654 9.3005
R10511 gnd.n3060 gnd.n2655 9.3005
R10512 gnd.n3059 gnd.n3058 9.3005
R10513 gnd.n2657 gnd.n2633 9.3005
R10514 gnd.n3091 gnd.n3090 9.3005
R10515 gnd.n3093 gnd.n2578 9.3005
R10516 gnd.n3140 gnd.n2579 9.3005
R10517 gnd.n3139 gnd.n2580 9.3005
R10518 gnd.n3138 gnd.n2581 9.3005
R10519 gnd.n3104 gnd.n2582 9.3005
R10520 gnd.n3106 gnd.n2600 9.3005
R10521 gnd.n3126 gnd.n2601 9.3005
R10522 gnd.n3125 gnd.n2602 9.3005
R10523 gnd.n3124 gnd.n2603 9.3005
R10524 gnd.n3115 gnd.n2604 9.3005
R10525 gnd.n3116 gnd.n2487 9.3005
R10526 gnd.n3182 gnd.n3181 9.3005
R10527 gnd.n3183 gnd.n2480 9.3005
R10528 gnd.n3193 gnd.n3192 9.3005
R10529 gnd.n3195 gnd.n2476 9.3005
R10530 gnd.n3205 gnd.n2477 9.3005
R10531 gnd.n3204 gnd.n3203 9.3005
R10532 gnd.n3201 gnd.n2455 9.3005
R10533 gnd.n3227 gnd.n2456 9.3005
R10534 gnd.n3226 gnd.n3225 9.3005
R10535 gnd.n2458 gnd.n2432 9.3005
R10536 gnd.n3267 gnd.n3266 9.3005
R10537 gnd.n3268 gnd.n2425 9.3005
R10538 gnd.n3278 gnd.n3277 9.3005
R10539 gnd.n3280 gnd.n2421 9.3005
R10540 gnd.n3290 gnd.n2422 9.3005
R10541 gnd.n3289 gnd.n3288 9.3005
R10542 gnd.n3286 gnd.n2400 9.3005
R10543 gnd.n3312 gnd.n2401 9.3005
R10544 gnd.n3311 gnd.n3310 9.3005
R10545 gnd.n2403 gnd.n2378 9.3005
R10546 gnd.n3356 gnd.n3355 9.3005
R10547 gnd.n3357 gnd.n2371 9.3005
R10548 gnd.n3367 gnd.n3366 9.3005
R10549 gnd.n3625 gnd.n2367 9.3005
R10550 gnd.n3633 gnd.n2368 9.3005
R10551 gnd.n3632 gnd.n3631 9.3005
R10552 gnd.n2349 gnd.n2348 9.3005
R10553 gnd.n3656 gnd.n3655 9.3005
R10554 gnd.n2799 gnd.n2798 9.3005
R10555 gnd.n6643 gnd.n6642 9.3005
R10556 gnd.n767 gnd.n766 9.3005
R10557 gnd.n6650 gnd.n6649 9.3005
R10558 gnd.n6651 gnd.n765 9.3005
R10559 gnd.n6653 gnd.n6652 9.3005
R10560 gnd.n761 gnd.n760 9.3005
R10561 gnd.n6660 gnd.n6659 9.3005
R10562 gnd.n6661 gnd.n759 9.3005
R10563 gnd.n6663 gnd.n6662 9.3005
R10564 gnd.n755 gnd.n754 9.3005
R10565 gnd.n6670 gnd.n6669 9.3005
R10566 gnd.n6671 gnd.n753 9.3005
R10567 gnd.n6673 gnd.n6672 9.3005
R10568 gnd.n749 gnd.n748 9.3005
R10569 gnd.n6680 gnd.n6679 9.3005
R10570 gnd.n6681 gnd.n747 9.3005
R10571 gnd.n6683 gnd.n6682 9.3005
R10572 gnd.n743 gnd.n742 9.3005
R10573 gnd.n6690 gnd.n6689 9.3005
R10574 gnd.n6691 gnd.n741 9.3005
R10575 gnd.n6693 gnd.n6692 9.3005
R10576 gnd.n737 gnd.n736 9.3005
R10577 gnd.n6700 gnd.n6699 9.3005
R10578 gnd.n6701 gnd.n735 9.3005
R10579 gnd.n6703 gnd.n6702 9.3005
R10580 gnd.n731 gnd.n730 9.3005
R10581 gnd.n6710 gnd.n6709 9.3005
R10582 gnd.n6711 gnd.n729 9.3005
R10583 gnd.n6713 gnd.n6712 9.3005
R10584 gnd.n725 gnd.n724 9.3005
R10585 gnd.n6720 gnd.n6719 9.3005
R10586 gnd.n6721 gnd.n723 9.3005
R10587 gnd.n6723 gnd.n6722 9.3005
R10588 gnd.n719 gnd.n718 9.3005
R10589 gnd.n6730 gnd.n6729 9.3005
R10590 gnd.n6731 gnd.n717 9.3005
R10591 gnd.n6733 gnd.n6732 9.3005
R10592 gnd.n713 gnd.n712 9.3005
R10593 gnd.n6740 gnd.n6739 9.3005
R10594 gnd.n6741 gnd.n711 9.3005
R10595 gnd.n6743 gnd.n6742 9.3005
R10596 gnd.n707 gnd.n706 9.3005
R10597 gnd.n6750 gnd.n6749 9.3005
R10598 gnd.n6751 gnd.n705 9.3005
R10599 gnd.n6753 gnd.n6752 9.3005
R10600 gnd.n701 gnd.n700 9.3005
R10601 gnd.n6760 gnd.n6759 9.3005
R10602 gnd.n6761 gnd.n699 9.3005
R10603 gnd.n6763 gnd.n6762 9.3005
R10604 gnd.n695 gnd.n694 9.3005
R10605 gnd.n6770 gnd.n6769 9.3005
R10606 gnd.n6771 gnd.n693 9.3005
R10607 gnd.n6773 gnd.n6772 9.3005
R10608 gnd.n689 gnd.n688 9.3005
R10609 gnd.n6780 gnd.n6779 9.3005
R10610 gnd.n6781 gnd.n687 9.3005
R10611 gnd.n6783 gnd.n6782 9.3005
R10612 gnd.n683 gnd.n682 9.3005
R10613 gnd.n6790 gnd.n6789 9.3005
R10614 gnd.n6791 gnd.n681 9.3005
R10615 gnd.n6793 gnd.n6792 9.3005
R10616 gnd.n677 gnd.n676 9.3005
R10617 gnd.n6800 gnd.n6799 9.3005
R10618 gnd.n6801 gnd.n675 9.3005
R10619 gnd.n6803 gnd.n6802 9.3005
R10620 gnd.n671 gnd.n670 9.3005
R10621 gnd.n6810 gnd.n6809 9.3005
R10622 gnd.n6811 gnd.n669 9.3005
R10623 gnd.n6813 gnd.n6812 9.3005
R10624 gnd.n665 gnd.n664 9.3005
R10625 gnd.n6820 gnd.n6819 9.3005
R10626 gnd.n6821 gnd.n663 9.3005
R10627 gnd.n6823 gnd.n6822 9.3005
R10628 gnd.n659 gnd.n658 9.3005
R10629 gnd.n6830 gnd.n6829 9.3005
R10630 gnd.n6831 gnd.n657 9.3005
R10631 gnd.n6833 gnd.n6832 9.3005
R10632 gnd.n653 gnd.n652 9.3005
R10633 gnd.n6840 gnd.n6839 9.3005
R10634 gnd.n6841 gnd.n651 9.3005
R10635 gnd.n6843 gnd.n6842 9.3005
R10636 gnd.n647 gnd.n646 9.3005
R10637 gnd.n6850 gnd.n6849 9.3005
R10638 gnd.n6851 gnd.n645 9.3005
R10639 gnd.n6853 gnd.n6852 9.3005
R10640 gnd.n641 gnd.n640 9.3005
R10641 gnd.n6860 gnd.n6859 9.3005
R10642 gnd.n6861 gnd.n639 9.3005
R10643 gnd.n6863 gnd.n6862 9.3005
R10644 gnd.n635 gnd.n634 9.3005
R10645 gnd.n6870 gnd.n6869 9.3005
R10646 gnd.n6871 gnd.n633 9.3005
R10647 gnd.n6873 gnd.n6872 9.3005
R10648 gnd.n629 gnd.n628 9.3005
R10649 gnd.n6880 gnd.n6879 9.3005
R10650 gnd.n6881 gnd.n627 9.3005
R10651 gnd.n6883 gnd.n6882 9.3005
R10652 gnd.n623 gnd.n622 9.3005
R10653 gnd.n6890 gnd.n6889 9.3005
R10654 gnd.n6891 gnd.n621 9.3005
R10655 gnd.n6893 gnd.n6892 9.3005
R10656 gnd.n617 gnd.n616 9.3005
R10657 gnd.n6900 gnd.n6899 9.3005
R10658 gnd.n6901 gnd.n615 9.3005
R10659 gnd.n6903 gnd.n6902 9.3005
R10660 gnd.n611 gnd.n610 9.3005
R10661 gnd.n6910 gnd.n6909 9.3005
R10662 gnd.n6911 gnd.n609 9.3005
R10663 gnd.n6913 gnd.n6912 9.3005
R10664 gnd.n605 gnd.n604 9.3005
R10665 gnd.n6920 gnd.n6919 9.3005
R10666 gnd.n6921 gnd.n603 9.3005
R10667 gnd.n6923 gnd.n6922 9.3005
R10668 gnd.n599 gnd.n598 9.3005
R10669 gnd.n6930 gnd.n6929 9.3005
R10670 gnd.n6931 gnd.n597 9.3005
R10671 gnd.n6933 gnd.n6932 9.3005
R10672 gnd.n593 gnd.n592 9.3005
R10673 gnd.n6940 gnd.n6939 9.3005
R10674 gnd.n6941 gnd.n591 9.3005
R10675 gnd.n6943 gnd.n6942 9.3005
R10676 gnd.n587 gnd.n586 9.3005
R10677 gnd.n6950 gnd.n6949 9.3005
R10678 gnd.n6951 gnd.n585 9.3005
R10679 gnd.n6953 gnd.n6952 9.3005
R10680 gnd.n581 gnd.n580 9.3005
R10681 gnd.n6960 gnd.n6959 9.3005
R10682 gnd.n6961 gnd.n579 9.3005
R10683 gnd.n6963 gnd.n6962 9.3005
R10684 gnd.n575 gnd.n574 9.3005
R10685 gnd.n6970 gnd.n6969 9.3005
R10686 gnd.n6971 gnd.n573 9.3005
R10687 gnd.n6973 gnd.n6972 9.3005
R10688 gnd.n569 gnd.n568 9.3005
R10689 gnd.n6980 gnd.n6979 9.3005
R10690 gnd.n6981 gnd.n567 9.3005
R10691 gnd.n6983 gnd.n6982 9.3005
R10692 gnd.n563 gnd.n562 9.3005
R10693 gnd.n6990 gnd.n6989 9.3005
R10694 gnd.n6991 gnd.n561 9.3005
R10695 gnd.n6993 gnd.n6992 9.3005
R10696 gnd.n557 gnd.n556 9.3005
R10697 gnd.n7000 gnd.n6999 9.3005
R10698 gnd.n7001 gnd.n555 9.3005
R10699 gnd.n7003 gnd.n7002 9.3005
R10700 gnd.n551 gnd.n550 9.3005
R10701 gnd.n7010 gnd.n7009 9.3005
R10702 gnd.n7011 gnd.n549 9.3005
R10703 gnd.n7013 gnd.n7012 9.3005
R10704 gnd.n545 gnd.n544 9.3005
R10705 gnd.n7020 gnd.n7019 9.3005
R10706 gnd.n7021 gnd.n543 9.3005
R10707 gnd.n7023 gnd.n7022 9.3005
R10708 gnd.n539 gnd.n538 9.3005
R10709 gnd.n7030 gnd.n7029 9.3005
R10710 gnd.n7031 gnd.n537 9.3005
R10711 gnd.n7033 gnd.n7032 9.3005
R10712 gnd.n533 gnd.n532 9.3005
R10713 gnd.n7040 gnd.n7039 9.3005
R10714 gnd.n7041 gnd.n531 9.3005
R10715 gnd.n7043 gnd.n7042 9.3005
R10716 gnd.n527 gnd.n526 9.3005
R10717 gnd.n7050 gnd.n7049 9.3005
R10718 gnd.n7051 gnd.n525 9.3005
R10719 gnd.n7054 gnd.n7053 9.3005
R10720 gnd.n7052 gnd.n521 9.3005
R10721 gnd.n7060 gnd.n520 9.3005
R10722 gnd.n7062 gnd.n7061 9.3005
R10723 gnd.n516 gnd.n515 9.3005
R10724 gnd.n7071 gnd.n7070 9.3005
R10725 gnd.n7072 gnd.n514 9.3005
R10726 gnd.n7074 gnd.n7073 9.3005
R10727 gnd.n510 gnd.n509 9.3005
R10728 gnd.n7081 gnd.n7080 9.3005
R10729 gnd.n7082 gnd.n508 9.3005
R10730 gnd.n7084 gnd.n7083 9.3005
R10731 gnd.n504 gnd.n503 9.3005
R10732 gnd.n7091 gnd.n7090 9.3005
R10733 gnd.n7092 gnd.n502 9.3005
R10734 gnd.n7094 gnd.n7093 9.3005
R10735 gnd.n498 gnd.n497 9.3005
R10736 gnd.n7101 gnd.n7100 9.3005
R10737 gnd.n7102 gnd.n496 9.3005
R10738 gnd.n7104 gnd.n7103 9.3005
R10739 gnd.n492 gnd.n491 9.3005
R10740 gnd.n7111 gnd.n7110 9.3005
R10741 gnd.n7112 gnd.n490 9.3005
R10742 gnd.n7114 gnd.n7113 9.3005
R10743 gnd.n486 gnd.n485 9.3005
R10744 gnd.n7121 gnd.n7120 9.3005
R10745 gnd.n7122 gnd.n484 9.3005
R10746 gnd.n7124 gnd.n7123 9.3005
R10747 gnd.n480 gnd.n479 9.3005
R10748 gnd.n7131 gnd.n7130 9.3005
R10749 gnd.n7132 gnd.n478 9.3005
R10750 gnd.n7134 gnd.n7133 9.3005
R10751 gnd.n474 gnd.n473 9.3005
R10752 gnd.n7141 gnd.n7140 9.3005
R10753 gnd.n7142 gnd.n472 9.3005
R10754 gnd.n7144 gnd.n7143 9.3005
R10755 gnd.n468 gnd.n467 9.3005
R10756 gnd.n7151 gnd.n7150 9.3005
R10757 gnd.n7152 gnd.n466 9.3005
R10758 gnd.n7154 gnd.n7153 9.3005
R10759 gnd.n462 gnd.n461 9.3005
R10760 gnd.n7161 gnd.n7160 9.3005
R10761 gnd.n7162 gnd.n460 9.3005
R10762 gnd.n7164 gnd.n7163 9.3005
R10763 gnd.n456 gnd.n455 9.3005
R10764 gnd.n7171 gnd.n7170 9.3005
R10765 gnd.n7172 gnd.n454 9.3005
R10766 gnd.n7174 gnd.n7173 9.3005
R10767 gnd.n450 gnd.n449 9.3005
R10768 gnd.n7181 gnd.n7180 9.3005
R10769 gnd.n7182 gnd.n448 9.3005
R10770 gnd.n7184 gnd.n7183 9.3005
R10771 gnd.n444 gnd.n443 9.3005
R10772 gnd.n7191 gnd.n7190 9.3005
R10773 gnd.n7192 gnd.n442 9.3005
R10774 gnd.n7194 gnd.n7193 9.3005
R10775 gnd.n438 gnd.n437 9.3005
R10776 gnd.n7201 gnd.n7200 9.3005
R10777 gnd.n7202 gnd.n436 9.3005
R10778 gnd.n7204 gnd.n7203 9.3005
R10779 gnd.n432 gnd.n431 9.3005
R10780 gnd.n7211 gnd.n7210 9.3005
R10781 gnd.n7212 gnd.n430 9.3005
R10782 gnd.n7214 gnd.n7213 9.3005
R10783 gnd.n426 gnd.n425 9.3005
R10784 gnd.n7221 gnd.n7220 9.3005
R10785 gnd.n7222 gnd.n424 9.3005
R10786 gnd.n7224 gnd.n7223 9.3005
R10787 gnd.n420 gnd.n419 9.3005
R10788 gnd.n7231 gnd.n7230 9.3005
R10789 gnd.n7232 gnd.n418 9.3005
R10790 gnd.n7234 gnd.n7233 9.3005
R10791 gnd.n414 gnd.n413 9.3005
R10792 gnd.n7241 gnd.n7240 9.3005
R10793 gnd.n7242 gnd.n412 9.3005
R10794 gnd.n7244 gnd.n7243 9.3005
R10795 gnd.n408 gnd.n407 9.3005
R10796 gnd.n7251 gnd.n7250 9.3005
R10797 gnd.n7252 gnd.n406 9.3005
R10798 gnd.n7254 gnd.n7253 9.3005
R10799 gnd.n402 gnd.n401 9.3005
R10800 gnd.n7261 gnd.n7260 9.3005
R10801 gnd.n7262 gnd.n400 9.3005
R10802 gnd.n7264 gnd.n7263 9.3005
R10803 gnd.n396 gnd.n395 9.3005
R10804 gnd.n7272 gnd.n7271 9.3005
R10805 gnd.n7273 gnd.n394 9.3005
R10806 gnd.n7276 gnd.n7275 9.3005
R10807 gnd.n7064 gnd.n7063 9.3005
R10808 gnd.n7642 gnd.n7641 9.3005
R10809 gnd.n7640 gnd.n80 9.3005
R10810 gnd.n361 gnd.n83 9.3005
R10811 gnd.n7327 gnd.n7326 9.3005
R10812 gnd.n7328 gnd.n360 9.3005
R10813 gnd.n7331 gnd.n7330 9.3005
R10814 gnd.n7329 gnd.n356 9.3005
R10815 gnd.n7345 gnd.n357 9.3005
R10816 gnd.n7346 gnd.n355 9.3005
R10817 gnd.n7349 gnd.n7348 9.3005
R10818 gnd.n7350 gnd.n354 9.3005
R10819 gnd.n7383 gnd.n7351 9.3005
R10820 gnd.n7382 gnd.n7352 9.3005
R10821 gnd.n7381 gnd.n7353 9.3005
R10822 gnd.n7379 gnd.n7354 9.3005
R10823 gnd.n7378 gnd.n7355 9.3005
R10824 gnd.n7376 gnd.n7356 9.3005
R10825 gnd.n7375 gnd.n7357 9.3005
R10826 gnd.n7373 gnd.n7358 9.3005
R10827 gnd.n7372 gnd.n7359 9.3005
R10828 gnd.n7370 gnd.n7360 9.3005
R10829 gnd.n7369 gnd.n7361 9.3005
R10830 gnd.n7367 gnd.n7362 9.3005
R10831 gnd.n7366 gnd.n7364 9.3005
R10832 gnd.n7363 gnd.n351 9.3005
R10833 gnd.n7415 gnd.n350 9.3005
R10834 gnd.n7417 gnd.n7416 9.3005
R10835 gnd.n7448 gnd.n316 9.3005
R10836 gnd.n7447 gnd.n318 9.3005
R10837 gnd.n322 gnd.n319 9.3005
R10838 gnd.n7442 gnd.n323 9.3005
R10839 gnd.n7441 gnd.n324 9.3005
R10840 gnd.n7440 gnd.n325 9.3005
R10841 gnd.n329 gnd.n326 9.3005
R10842 gnd.n7435 gnd.n330 9.3005
R10843 gnd.n7434 gnd.n331 9.3005
R10844 gnd.n7433 gnd.n332 9.3005
R10845 gnd.n336 gnd.n333 9.3005
R10846 gnd.n7428 gnd.n337 9.3005
R10847 gnd.n7427 gnd.n338 9.3005
R10848 gnd.n7426 gnd.n339 9.3005
R10849 gnd.n343 gnd.n340 9.3005
R10850 gnd.n7421 gnd.n344 9.3005
R10851 gnd.n7420 gnd.n7419 9.3005
R10852 gnd.n7418 gnd.n347 9.3005
R10853 gnd.n7450 gnd.n7449 9.3005
R10854 gnd.n7558 gnd.n213 9.3005
R10855 gnd.n7557 gnd.n215 9.3005
R10856 gnd.n219 gnd.n216 9.3005
R10857 gnd.n7552 gnd.n220 9.3005
R10858 gnd.n7551 gnd.n221 9.3005
R10859 gnd.n7550 gnd.n222 9.3005
R10860 gnd.n226 gnd.n223 9.3005
R10861 gnd.n7545 gnd.n227 9.3005
R10862 gnd.n7544 gnd.n228 9.3005
R10863 gnd.n7543 gnd.n229 9.3005
R10864 gnd.n233 gnd.n230 9.3005
R10865 gnd.n7538 gnd.n234 9.3005
R10866 gnd.n7537 gnd.n235 9.3005
R10867 gnd.n7536 gnd.n236 9.3005
R10868 gnd.n240 gnd.n237 9.3005
R10869 gnd.n7531 gnd.n241 9.3005
R10870 gnd.n7530 gnd.n242 9.3005
R10871 gnd.n7526 gnd.n243 9.3005
R10872 gnd.n247 gnd.n244 9.3005
R10873 gnd.n7521 gnd.n248 9.3005
R10874 gnd.n7520 gnd.n249 9.3005
R10875 gnd.n7519 gnd.n250 9.3005
R10876 gnd.n254 gnd.n251 9.3005
R10877 gnd.n7514 gnd.n255 9.3005
R10878 gnd.n7513 gnd.n256 9.3005
R10879 gnd.n7512 gnd.n257 9.3005
R10880 gnd.n261 gnd.n258 9.3005
R10881 gnd.n7507 gnd.n262 9.3005
R10882 gnd.n7506 gnd.n263 9.3005
R10883 gnd.n7505 gnd.n264 9.3005
R10884 gnd.n268 gnd.n265 9.3005
R10885 gnd.n7500 gnd.n269 9.3005
R10886 gnd.n7499 gnd.n270 9.3005
R10887 gnd.n7498 gnd.n271 9.3005
R10888 gnd.n275 gnd.n272 9.3005
R10889 gnd.n7493 gnd.n276 9.3005
R10890 gnd.n7492 gnd.n7491 9.3005
R10891 gnd.n7490 gnd.n277 9.3005
R10892 gnd.n7489 gnd.n7488 9.3005
R10893 gnd.n281 gnd.n280 9.3005
R10894 gnd.n286 gnd.n284 9.3005
R10895 gnd.n7481 gnd.n287 9.3005
R10896 gnd.n7480 gnd.n288 9.3005
R10897 gnd.n7479 gnd.n289 9.3005
R10898 gnd.n293 gnd.n290 9.3005
R10899 gnd.n7474 gnd.n294 9.3005
R10900 gnd.n7473 gnd.n295 9.3005
R10901 gnd.n7472 gnd.n296 9.3005
R10902 gnd.n300 gnd.n297 9.3005
R10903 gnd.n7467 gnd.n301 9.3005
R10904 gnd.n7466 gnd.n302 9.3005
R10905 gnd.n7465 gnd.n303 9.3005
R10906 gnd.n307 gnd.n304 9.3005
R10907 gnd.n7460 gnd.n308 9.3005
R10908 gnd.n7459 gnd.n309 9.3005
R10909 gnd.n7458 gnd.n310 9.3005
R10910 gnd.n315 gnd.n313 9.3005
R10911 gnd.n7453 gnd.n7452 9.3005
R10912 gnd.n7560 gnd.n7559 9.3005
R10913 gnd.n5904 gnd.n1355 9.3005
R10914 gnd.n6114 gnd.n1356 9.3005
R10915 gnd.n6113 gnd.n1357 9.3005
R10916 gnd.n6112 gnd.n1358 9.3005
R10917 gnd.n1492 gnd.n1359 9.3005
R10918 gnd.n6102 gnd.n1376 9.3005
R10919 gnd.n6101 gnd.n1377 9.3005
R10920 gnd.n6100 gnd.n1378 9.3005
R10921 gnd.n5923 gnd.n1379 9.3005
R10922 gnd.n6090 gnd.n1397 9.3005
R10923 gnd.n6089 gnd.n1398 9.3005
R10924 gnd.n6088 gnd.n1399 9.3005
R10925 gnd.n1477 gnd.n1400 9.3005
R10926 gnd.n6078 gnd.n1416 9.3005
R10927 gnd.n6077 gnd.n1417 9.3005
R10928 gnd.n6076 gnd.n1418 9.3005
R10929 gnd.n1471 gnd.n1419 9.3005
R10930 gnd.n6066 gnd.n1437 9.3005
R10931 gnd.n6065 gnd.n1438 9.3005
R10932 gnd.n6064 gnd.n1439 9.3005
R10933 gnd.n6018 gnd.n1440 9.3005
R10934 gnd.n6054 gnd.n1454 9.3005
R10935 gnd.n6053 gnd.n6052 9.3005
R10936 gnd.n373 gnd.n372 9.3005
R10937 gnd.n7307 gnd.n7306 9.3005
R10938 gnd.n7308 gnd.n366 9.3005
R10939 gnd.n7315 gnd.n367 9.3005
R10940 gnd.n7316 gnd.n365 9.3005
R10941 gnd.n7320 gnd.n7319 9.3005
R10942 gnd.n7321 gnd.n108 9.3005
R10943 gnd.n7628 gnd.n109 9.3005
R10944 gnd.n7627 gnd.n110 9.3005
R10945 gnd.n7626 gnd.n111 9.3005
R10946 gnd.n7337 gnd.n112 9.3005
R10947 gnd.n7616 gnd.n127 9.3005
R10948 gnd.n7615 gnd.n128 9.3005
R10949 gnd.n7614 gnd.n129 9.3005
R10950 gnd.n353 gnd.n130 9.3005
R10951 gnd.n7604 gnd.n147 9.3005
R10952 gnd.n7603 gnd.n148 9.3005
R10953 gnd.n7602 gnd.n149 9.3005
R10954 gnd.n7392 gnd.n150 9.3005
R10955 gnd.n7592 gnd.n165 9.3005
R10956 gnd.n7591 gnd.n166 9.3005
R10957 gnd.n7590 gnd.n167 9.3005
R10958 gnd.n7399 gnd.n168 9.3005
R10959 gnd.n7580 gnd.n185 9.3005
R10960 gnd.n7579 gnd.n186 9.3005
R10961 gnd.n7578 gnd.n187 9.3005
R10962 gnd.n7406 gnd.n188 9.3005
R10963 gnd.n7568 gnd.n203 9.3005
R10964 gnd.n7567 gnd.n204 9.3005
R10965 gnd.n7566 gnd.n205 9.3005
R10966 gnd.n5903 gnd.n5902 9.3005
R10967 gnd.n5905 gnd.n5904 9.3005
R10968 gnd.n5906 gnd.n1356 9.3005
R10969 gnd.n5907 gnd.n1357 9.3005
R10970 gnd.n1491 gnd.n1358 9.3005
R10971 gnd.n5919 gnd.n1492 9.3005
R10972 gnd.n5920 gnd.n1376 9.3005
R10973 gnd.n5921 gnd.n1377 9.3005
R10974 gnd.n5922 gnd.n1378 9.3005
R10975 gnd.n5926 gnd.n5923 9.3005
R10976 gnd.n5925 gnd.n1397 9.3005
R10977 gnd.n5924 gnd.n1398 9.3005
R10978 gnd.n1476 gnd.n1399 9.3005
R10979 gnd.n6000 gnd.n1477 9.3005
R10980 gnd.n6001 gnd.n1416 9.3005
R10981 gnd.n6002 gnd.n1417 9.3005
R10982 gnd.n1470 gnd.n1418 9.3005
R10983 gnd.n6014 gnd.n1471 9.3005
R10984 gnd.n6015 gnd.n1437 9.3005
R10985 gnd.n6016 gnd.n1438 9.3005
R10986 gnd.n6017 gnd.n1439 9.3005
R10987 gnd.n6019 gnd.n6018 9.3005
R10988 gnd.n1455 gnd.n1454 9.3005
R10989 gnd.n6052 gnd.n6051 9.3005
R10990 gnd.n1456 gnd.n372 9.3005
R10991 gnd.n7307 gnd.n371 9.3005
R10992 gnd.n7309 gnd.n7308 9.3005
R10993 gnd.n7311 gnd.n367 9.3005
R10994 gnd.n7310 gnd.n365 9.3005
R10995 gnd.n7320 gnd.n364 9.3005
R10996 gnd.n7322 gnd.n7321 9.3005
R10997 gnd.n359 gnd.n109 9.3005
R10998 gnd.n7335 gnd.n110 9.3005
R10999 gnd.n7336 gnd.n111 9.3005
R11000 gnd.n7341 gnd.n7337 9.3005
R11001 gnd.n7340 gnd.n127 9.3005
R11002 gnd.n7339 gnd.n128 9.3005
R11003 gnd.n352 gnd.n129 9.3005
R11004 gnd.n7387 gnd.n353 9.3005
R11005 gnd.n7388 gnd.n147 9.3005
R11006 gnd.n7390 gnd.n148 9.3005
R11007 gnd.n7391 gnd.n149 9.3005
R11008 gnd.n7394 gnd.n7392 9.3005
R11009 gnd.n7395 gnd.n165 9.3005
R11010 gnd.n7397 gnd.n166 9.3005
R11011 gnd.n7398 gnd.n167 9.3005
R11012 gnd.n7401 gnd.n7399 9.3005
R11013 gnd.n7402 gnd.n185 9.3005
R11014 gnd.n7404 gnd.n186 9.3005
R11015 gnd.n7405 gnd.n187 9.3005
R11016 gnd.n7408 gnd.n7406 9.3005
R11017 gnd.n7409 gnd.n203 9.3005
R11018 gnd.n7411 gnd.n204 9.3005
R11019 gnd.n7410 gnd.n205 9.3005
R11020 gnd.n5903 gnd.n1496 9.3005
R11021 gnd.n1502 gnd.n1499 9.3005
R11022 gnd.n5890 gnd.n1503 9.3005
R11023 gnd.n5892 gnd.n5891 9.3005
R11024 gnd.n5889 gnd.n1505 9.3005
R11025 gnd.n5888 gnd.n5887 9.3005
R11026 gnd.n1507 gnd.n1506 9.3005
R11027 gnd.n5881 gnd.n5880 9.3005
R11028 gnd.n5879 gnd.n1509 9.3005
R11029 gnd.n5878 gnd.n5877 9.3005
R11030 gnd.n1511 gnd.n1510 9.3005
R11031 gnd.n5871 gnd.n5870 9.3005
R11032 gnd.n5869 gnd.n1513 9.3005
R11033 gnd.n5868 gnd.n5867 9.3005
R11034 gnd.n1515 gnd.n1514 9.3005
R11035 gnd.n5861 gnd.n5860 9.3005
R11036 gnd.n5859 gnd.n1517 9.3005
R11037 gnd.n5858 gnd.n5857 9.3005
R11038 gnd.n1519 gnd.n1518 9.3005
R11039 gnd.n5851 gnd.n5850 9.3005
R11040 gnd.n5849 gnd.n1521 9.3005
R11041 gnd.n1523 gnd.n1522 9.3005
R11042 gnd.n5839 gnd.n5838 9.3005
R11043 gnd.n5837 gnd.n1525 9.3005
R11044 gnd.n5836 gnd.n5835 9.3005
R11045 gnd.n1527 gnd.n1526 9.3005
R11046 gnd.n5829 gnd.n5828 9.3005
R11047 gnd.n5827 gnd.n1529 9.3005
R11048 gnd.n5826 gnd.n5825 9.3005
R11049 gnd.n1531 gnd.n1530 9.3005
R11050 gnd.n5817 gnd.n5816 9.3005
R11051 gnd.n5814 gnd.n5727 9.3005
R11052 gnd.n5813 gnd.n5812 9.3005
R11053 gnd.n5729 gnd.n5728 9.3005
R11054 gnd.n5806 gnd.n5805 9.3005
R11055 gnd.n5804 gnd.n5731 9.3005
R11056 gnd.n5803 gnd.n5802 9.3005
R11057 gnd.n5733 gnd.n5732 9.3005
R11058 gnd.n5796 gnd.n5792 9.3005
R11059 gnd.n5791 gnd.n5735 9.3005
R11060 gnd.n5790 gnd.n5789 9.3005
R11061 gnd.n5737 gnd.n5736 9.3005
R11062 gnd.n5783 gnd.n5782 9.3005
R11063 gnd.n5781 gnd.n5739 9.3005
R11064 gnd.n5780 gnd.n5779 9.3005
R11065 gnd.n5741 gnd.n5740 9.3005
R11066 gnd.n5773 gnd.n5772 9.3005
R11067 gnd.n5771 gnd.n5743 9.3005
R11068 gnd.n5770 gnd.n5769 9.3005
R11069 gnd.n5745 gnd.n5744 9.3005
R11070 gnd.n5763 gnd.n5762 9.3005
R11071 gnd.n5761 gnd.n5747 9.3005
R11072 gnd.n5760 gnd.n5759 9.3005
R11073 gnd.n5749 gnd.n5748 9.3005
R11074 gnd.n5753 gnd.n5752 9.3005
R11075 gnd.n5751 gnd.n5750 9.3005
R11076 gnd.n5848 gnd.n5847 9.3005
R11077 gnd.n5900 gnd.n5899 9.3005
R11078 gnd.n6119 gnd.n1345 9.3005
R11079 gnd.n6118 gnd.n1346 9.3005
R11080 gnd.n1366 gnd.n1347 9.3005
R11081 gnd.n6108 gnd.n1367 9.3005
R11082 gnd.n6107 gnd.n1368 9.3005
R11083 gnd.n6106 gnd.n1369 9.3005
R11084 gnd.n1386 gnd.n1370 9.3005
R11085 gnd.n6096 gnd.n1387 9.3005
R11086 gnd.n6095 gnd.n1388 9.3005
R11087 gnd.n6094 gnd.n1389 9.3005
R11088 gnd.n1406 gnd.n1390 9.3005
R11089 gnd.n6084 gnd.n1407 9.3005
R11090 gnd.n6083 gnd.n1408 9.3005
R11091 gnd.n6082 gnd.n1409 9.3005
R11092 gnd.n1426 gnd.n1410 9.3005
R11093 gnd.n6072 gnd.n1427 9.3005
R11094 gnd.n6071 gnd.n1428 9.3005
R11095 gnd.n6070 gnd.n1429 9.3005
R11096 gnd.n1446 gnd.n1430 9.3005
R11097 gnd.n6060 gnd.n1447 9.3005
R11098 gnd.n6059 gnd.n94 9.3005
R11099 gnd.n99 gnd.n93 9.3005
R11100 gnd.n7622 gnd.n118 9.3005
R11101 gnd.n7621 gnd.n119 9.3005
R11102 gnd.n7620 gnd.n120 9.3005
R11103 gnd.n137 gnd.n121 9.3005
R11104 gnd.n7610 gnd.n138 9.3005
R11105 gnd.n7609 gnd.n139 9.3005
R11106 gnd.n7608 gnd.n140 9.3005
R11107 gnd.n155 gnd.n141 9.3005
R11108 gnd.n7598 gnd.n156 9.3005
R11109 gnd.n7597 gnd.n157 9.3005
R11110 gnd.n7596 gnd.n158 9.3005
R11111 gnd.n175 gnd.n159 9.3005
R11112 gnd.n7586 gnd.n176 9.3005
R11113 gnd.n7585 gnd.n177 9.3005
R11114 gnd.n7584 gnd.n178 9.3005
R11115 gnd.n194 gnd.n179 9.3005
R11116 gnd.n7574 gnd.n195 9.3005
R11117 gnd.n7573 gnd.n196 9.3005
R11118 gnd.n7572 gnd.n197 9.3005
R11119 gnd.n212 gnd.n198 9.3005
R11120 gnd.n7562 gnd.n7561 9.3005
R11121 gnd.n6120 gnd.n1344 9.3005
R11122 gnd.n7633 gnd.n97 9.3005
R11123 gnd.n7633 gnd.n7632 9.3005
R11124 gnd.n4283 gnd.n4282 9.3005
R11125 gnd.n4284 gnd.n2126 9.3005
R11126 gnd.n4286 gnd.n4285 9.3005
R11127 gnd.n2124 gnd.n2123 9.3005
R11128 gnd.n4291 gnd.n4290 9.3005
R11129 gnd.n4292 gnd.n2122 9.3005
R11130 gnd.n4313 gnd.n4293 9.3005
R11131 gnd.n4312 gnd.n4294 9.3005
R11132 gnd.n4311 gnd.n4295 9.3005
R11133 gnd.n4298 gnd.n4296 9.3005
R11134 gnd.n4307 gnd.n4299 9.3005
R11135 gnd.n4306 gnd.n4300 9.3005
R11136 gnd.n4305 gnd.n4301 9.3005
R11137 gnd.n4303 gnd.n4302 9.3005
R11138 gnd.n2099 gnd.n2098 9.3005
R11139 gnd.n4378 gnd.n4377 9.3005
R11140 gnd.n4379 gnd.n2097 9.3005
R11141 gnd.n4381 gnd.n4380 9.3005
R11142 gnd.n2095 gnd.n2094 9.3005
R11143 gnd.n4386 gnd.n4385 9.3005
R11144 gnd.n4387 gnd.n2093 9.3005
R11145 gnd.n4389 gnd.n4388 9.3005
R11146 gnd.n2091 gnd.n2090 9.3005
R11147 gnd.n4396 gnd.n4395 9.3005
R11148 gnd.n4397 gnd.n2089 9.3005
R11149 gnd.n4399 gnd.n4398 9.3005
R11150 gnd.n2066 gnd.n2065 9.3005
R11151 gnd.n4680 gnd.n4679 9.3005
R11152 gnd.n4681 gnd.n2064 9.3005
R11153 gnd.n4685 gnd.n4682 9.3005
R11154 gnd.n4684 gnd.n4683 9.3005
R11155 gnd.n2041 gnd.n2040 9.3005
R11156 gnd.n4712 gnd.n4711 9.3005
R11157 gnd.n4713 gnd.n2039 9.3005
R11158 gnd.n4718 gnd.n4714 9.3005
R11159 gnd.n4717 gnd.n4716 9.3005
R11160 gnd.n4715 gnd.n1215 9.3005
R11161 gnd.n6253 gnd.n1216 9.3005
R11162 gnd.n6252 gnd.n1217 9.3005
R11163 gnd.n6251 gnd.n1218 9.3005
R11164 gnd.n4752 gnd.n1219 9.3005
R11165 gnd.n4754 gnd.n4753 9.3005
R11166 gnd.n1915 gnd.n1914 9.3005
R11167 gnd.n4794 gnd.n4793 9.3005
R11168 gnd.n4795 gnd.n1913 9.3005
R11169 gnd.n4797 gnd.n4796 9.3005
R11170 gnd.n1897 gnd.n1896 9.3005
R11171 gnd.n4836 gnd.n4835 9.3005
R11172 gnd.n4837 gnd.n1895 9.3005
R11173 gnd.n4841 gnd.n4838 9.3005
R11174 gnd.n4840 gnd.n4839 9.3005
R11175 gnd.n1871 gnd.n1870 9.3005
R11176 gnd.n4898 gnd.n4897 9.3005
R11177 gnd.n4899 gnd.n1869 9.3005
R11178 gnd.n4901 gnd.n4900 9.3005
R11179 gnd.n1853 gnd.n1852 9.3005
R11180 gnd.n4926 gnd.n4925 9.3005
R11181 gnd.n4927 gnd.n1851 9.3005
R11182 gnd.n4931 gnd.n4928 9.3005
R11183 gnd.n4930 gnd.n4929 9.3005
R11184 gnd.n1820 gnd.n1819 9.3005
R11185 gnd.n4976 gnd.n4975 9.3005
R11186 gnd.n4977 gnd.n1818 9.3005
R11187 gnd.n4979 gnd.n4978 9.3005
R11188 gnd.n1797 gnd.n1796 9.3005
R11189 gnd.n5016 gnd.n5015 9.3005
R11190 gnd.n5017 gnd.n1795 9.3005
R11191 gnd.n5019 gnd.n5018 9.3005
R11192 gnd.n1775 gnd.n1774 9.3005
R11193 gnd.n5073 gnd.n5072 9.3005
R11194 gnd.n5074 gnd.n1773 9.3005
R11195 gnd.n5076 gnd.n5075 9.3005
R11196 gnd.n1755 gnd.n1754 9.3005
R11197 gnd.n5098 gnd.n5097 9.3005
R11198 gnd.n5099 gnd.n1753 9.3005
R11199 gnd.n5101 gnd.n5100 9.3005
R11200 gnd.n1735 gnd.n1734 9.3005
R11201 gnd.n5158 gnd.n5157 9.3005
R11202 gnd.n5159 gnd.n1733 9.3005
R11203 gnd.n5161 gnd.n5160 9.3005
R11204 gnd.n1713 gnd.n1712 9.3005
R11205 gnd.n5187 gnd.n5186 9.3005
R11206 gnd.n5188 gnd.n1711 9.3005
R11207 gnd.n5192 gnd.n5189 9.3005
R11208 gnd.n5191 gnd.n5190 9.3005
R11209 gnd.n1685 gnd.n1684 9.3005
R11210 gnd.n5238 gnd.n5237 9.3005
R11211 gnd.n5239 gnd.n1683 9.3005
R11212 gnd.n5241 gnd.n5240 9.3005
R11213 gnd.n1665 gnd.n1664 9.3005
R11214 gnd.n5264 gnd.n5263 9.3005
R11215 gnd.n5265 gnd.n1663 9.3005
R11216 gnd.n5269 gnd.n5266 9.3005
R11217 gnd.n5268 gnd.n5267 9.3005
R11218 gnd.n1635 gnd.n1634 9.3005
R11219 gnd.n5308 gnd.n5307 9.3005
R11220 gnd.n5309 gnd.n1633 9.3005
R11221 gnd.n5314 gnd.n5310 9.3005
R11222 gnd.n5313 gnd.n5312 9.3005
R11223 gnd.n5311 gnd.n1584 9.3005
R11224 gnd.n5560 gnd.n1585 9.3005
R11225 gnd.n5559 gnd.n1586 9.3005
R11226 gnd.n5558 gnd.n1587 9.3005
R11227 gnd.n1596 gnd.n1588 9.3005
R11228 gnd.n1597 gnd.n1595 9.3005
R11229 gnd.n5548 gnd.n1598 9.3005
R11230 gnd.n5547 gnd.n1599 9.3005
R11231 gnd.n5546 gnd.n1600 9.3005
R11232 gnd.n1603 gnd.n1602 9.3005
R11233 gnd.n1601 gnd.n1322 9.3005
R11234 gnd.n6135 gnd.n1323 9.3005
R11235 gnd.n6134 gnd.n1324 9.3005
R11236 gnd.n6133 gnd.n1325 9.3005
R11237 gnd.n1331 gnd.n1326 9.3005
R11238 gnd.n6127 gnd.n1332 9.3005
R11239 gnd.n6126 gnd.n1333 9.3005
R11240 gnd.n6125 gnd.n1334 9.3005
R11241 gnd.n5944 gnd.n1335 9.3005
R11242 gnd.n5947 gnd.n5946 9.3005
R11243 gnd.n5948 gnd.n5943 9.3005
R11244 gnd.n5950 gnd.n5949 9.3005
R11245 gnd.n5941 gnd.n5940 9.3005
R11246 gnd.n5955 gnd.n5954 9.3005
R11247 gnd.n5956 gnd.n5939 9.3005
R11248 gnd.n5958 gnd.n5957 9.3005
R11249 gnd.n1486 gnd.n1485 9.3005
R11250 gnd.n5963 gnd.n5962 9.3005
R11251 gnd.n5964 gnd.n1484 9.3005
R11252 gnd.n5987 gnd.n5965 9.3005
R11253 gnd.n5986 gnd.n5966 9.3005
R11254 gnd.n5985 gnd.n5967 9.3005
R11255 gnd.n5970 gnd.n5968 9.3005
R11256 gnd.n5981 gnd.n5971 9.3005
R11257 gnd.n5980 gnd.n5972 9.3005
R11258 gnd.n5979 gnd.n5973 9.3005
R11259 gnd.n5977 gnd.n5976 9.3005
R11260 gnd.n5975 gnd.n1464 9.3005
R11261 gnd.n5974 gnd.n1462 9.3005
R11262 gnd.n388 gnd.n386 9.3005
R11263 gnd.n7283 gnd.n389 9.3005
R11264 gnd.n7282 gnd.n390 9.3005
R11265 gnd.n7281 gnd.n391 9.3005
R11266 gnd.n7274 gnd.n392 9.3005
R11267 gnd.n3882 gnd.n3871 9.3005
R11268 gnd.n3881 gnd.n3872 9.3005
R11269 gnd.n3879 gnd.n3873 9.3005
R11270 gnd.n3878 gnd.n3874 9.3005
R11271 gnd.n3876 gnd.n3875 9.3005
R11272 gnd.n2229 gnd.n2228 9.3005
R11273 gnd.n4090 gnd.n4089 9.3005
R11274 gnd.n4091 gnd.n2227 9.3005
R11275 gnd.n4097 gnd.n4092 9.3005
R11276 gnd.n4096 gnd.n4093 9.3005
R11277 gnd.n4095 gnd.n4094 9.3005
R11278 gnd.n2204 gnd.n2203 9.3005
R11279 gnd.n4125 gnd.n4124 9.3005
R11280 gnd.n4126 gnd.n2202 9.3005
R11281 gnd.n4134 gnd.n4127 9.3005
R11282 gnd.n4133 gnd.n4128 9.3005
R11283 gnd.n4132 gnd.n4130 9.3005
R11284 gnd.n4129 gnd.n2174 9.3005
R11285 gnd.n4188 gnd.n2175 9.3005
R11286 gnd.n4187 gnd.n2176 9.3005
R11287 gnd.n4186 gnd.n2177 9.3005
R11288 gnd.n4171 gnd.n2178 9.3005
R11289 gnd.n4172 gnd.n4170 9.3005
R11290 gnd.n4174 gnd.n4173 9.3005
R11291 gnd.n2152 gnd.n2151 9.3005
R11292 gnd.n4230 gnd.n4229 9.3005
R11293 gnd.n3885 gnd.n3884 9.3005
R11294 gnd.n3890 gnd.n3889 9.3005
R11295 gnd.n3893 gnd.n3866 9.3005
R11296 gnd.n3894 gnd.n3865 9.3005
R11297 gnd.n3897 gnd.n3864 9.3005
R11298 gnd.n3898 gnd.n3863 9.3005
R11299 gnd.n3901 gnd.n3862 9.3005
R11300 gnd.n3902 gnd.n3861 9.3005
R11301 gnd.n3905 gnd.n3860 9.3005
R11302 gnd.n3906 gnd.n3859 9.3005
R11303 gnd.n3909 gnd.n3858 9.3005
R11304 gnd.n3910 gnd.n3857 9.3005
R11305 gnd.n3913 gnd.n3856 9.3005
R11306 gnd.n3914 gnd.n3855 9.3005
R11307 gnd.n3917 gnd.n3854 9.3005
R11308 gnd.n3918 gnd.n3853 9.3005
R11309 gnd.n3921 gnd.n3852 9.3005
R11310 gnd.n3924 gnd.n3923 9.3005
R11311 gnd.n3888 gnd.n3870 9.3005
R11312 gnd.n3887 gnd.n3886 9.3005
R11313 gnd.n6331 gnd.n1143 9.3005
R11314 gnd.n6332 gnd.n1142 9.3005
R11315 gnd.n1141 gnd.n1138 9.3005
R11316 gnd.n6337 gnd.n1137 9.3005
R11317 gnd.n6338 gnd.n1136 9.3005
R11318 gnd.n6339 gnd.n1135 9.3005
R11319 gnd.n1134 gnd.n1131 9.3005
R11320 gnd.n6344 gnd.n1130 9.3005
R11321 gnd.n6346 gnd.n1127 9.3005
R11322 gnd.n6347 gnd.n1126 9.3005
R11323 gnd.n1125 gnd.n1122 9.3005
R11324 gnd.n6352 gnd.n1121 9.3005
R11325 gnd.n6353 gnd.n1120 9.3005
R11326 gnd.n6354 gnd.n1119 9.3005
R11327 gnd.n1118 gnd.n1115 9.3005
R11328 gnd.n6359 gnd.n1114 9.3005
R11329 gnd.n6360 gnd.n1113 9.3005
R11330 gnd.n6361 gnd.n1112 9.3005
R11331 gnd.n1111 gnd.n1108 9.3005
R11332 gnd.n6366 gnd.n1107 9.3005
R11333 gnd.n6367 gnd.n1106 9.3005
R11334 gnd.n6368 gnd.n1105 9.3005
R11335 gnd.n1104 gnd.n1101 9.3005
R11336 gnd.n1103 gnd.n1099 9.3005
R11337 gnd.n6375 gnd.n1098 9.3005
R11338 gnd.n6377 gnd.n6376 9.3005
R11339 gnd.n4457 gnd.n4456 9.3005
R11340 gnd.n4465 gnd.n4464 9.3005
R11341 gnd.n4466 gnd.n4454 9.3005
R11342 gnd.n4468 gnd.n4467 9.3005
R11343 gnd.n4452 gnd.n4451 9.3005
R11344 gnd.n4475 gnd.n4474 9.3005
R11345 gnd.n4476 gnd.n4450 9.3005
R11346 gnd.n4478 gnd.n4477 9.3005
R11347 gnd.n4448 gnd.n4445 9.3005
R11348 gnd.n4485 gnd.n4484 9.3005
R11349 gnd.n4486 gnd.n4444 9.3005
R11350 gnd.n4488 gnd.n4487 9.3005
R11351 gnd.n4442 gnd.n4441 9.3005
R11352 gnd.n4495 gnd.n4494 9.3005
R11353 gnd.n4496 gnd.n4440 9.3005
R11354 gnd.n4498 gnd.n4497 9.3005
R11355 gnd.n4438 gnd.n4437 9.3005
R11356 gnd.n4505 gnd.n4504 9.3005
R11357 gnd.n4506 gnd.n4436 9.3005
R11358 gnd.n4508 gnd.n4507 9.3005
R11359 gnd.n4434 gnd.n4433 9.3005
R11360 gnd.n4515 gnd.n4514 9.3005
R11361 gnd.n4516 gnd.n4432 9.3005
R11362 gnd.n4518 gnd.n4517 9.3005
R11363 gnd.n4430 gnd.n4429 9.3005
R11364 gnd.n4525 gnd.n4524 9.3005
R11365 gnd.n4526 gnd.n4428 9.3005
R11366 gnd.n4528 gnd.n4527 9.3005
R11367 gnd.n4426 gnd.n4423 9.3005
R11368 gnd.n4534 gnd.n4533 9.3005
R11369 gnd.n4455 gnd.n1144 9.3005
R11370 gnd.n4051 gnd.n4050 9.3005
R11371 gnd.n2269 gnd.n2265 9.3005
R11372 gnd.n2268 gnd.n2267 9.3005
R11373 gnd.n2249 gnd.n2245 9.3005
R11374 gnd.n4075 gnd.n2246 9.3005
R11375 gnd.n4074 gnd.n2247 9.3005
R11376 gnd.n4073 gnd.n4069 9.3005
R11377 gnd.n4072 gnd.n4070 9.3005
R11378 gnd.n2223 gnd.n2218 9.3005
R11379 gnd.n4111 gnd.n2219 9.3005
R11380 gnd.n4110 gnd.n2220 9.3005
R11381 gnd.n4109 gnd.n4108 9.3005
R11382 gnd.n2221 gnd.n2195 9.3005
R11383 gnd.n4141 gnd.n2196 9.3005
R11384 gnd.n4140 gnd.n4139 9.3005
R11385 gnd.n2197 gnd.n2181 9.3005
R11386 gnd.n4155 gnd.n2180 9.3005
R11387 gnd.n4157 gnd.n4156 9.3005
R11388 gnd.n4158 gnd.n959 9.3005
R11389 gnd.n6458 gnd.n960 9.3005
R11390 gnd.n6457 gnd.n961 9.3005
R11391 gnd.n6456 gnd.n962 9.3005
R11392 gnd.n4161 gnd.n963 9.3005
R11393 gnd.n4162 gnd.n2163 9.3005
R11394 gnd.n4220 gnd.n2164 9.3005
R11395 gnd.n4219 gnd.n2165 9.3005
R11396 gnd.n4218 gnd.n2166 9.3005
R11397 gnd.n2143 gnd.n2142 9.3005
R11398 gnd.n4244 gnd.n4243 9.3005
R11399 gnd.n4245 gnd.n987 9.3005
R11400 gnd.n6445 gnd.n988 9.3005
R11401 gnd.n6444 gnd.n989 9.3005
R11402 gnd.n6443 gnd.n990 9.3005
R11403 gnd.n4252 gnd.n991 9.3005
R11404 gnd.n6433 gnd.n1007 9.3005
R11405 gnd.n6432 gnd.n1008 9.3005
R11406 gnd.n6431 gnd.n1009 9.3005
R11407 gnd.n4258 gnd.n1010 9.3005
R11408 gnd.n6421 gnd.n1027 9.3005
R11409 gnd.n6420 gnd.n1028 9.3005
R11410 gnd.n6419 gnd.n1029 9.3005
R11411 gnd.n4328 gnd.n1030 9.3005
R11412 gnd.n6409 gnd.n1047 9.3005
R11413 gnd.n6408 gnd.n1048 9.3005
R11414 gnd.n6407 gnd.n1049 9.3005
R11415 gnd.n4343 gnd.n1050 9.3005
R11416 gnd.n6397 gnd.n1067 9.3005
R11417 gnd.n6396 gnd.n1068 9.3005
R11418 gnd.n6395 gnd.n1069 9.3005
R11419 gnd.n4350 gnd.n1070 9.3005
R11420 gnd.n6385 gnd.n1088 9.3005
R11421 gnd.n6384 gnd.n1089 9.3005
R11422 gnd.n6383 gnd.n1090 9.3005
R11423 gnd.n2266 gnd.n2264 9.3005
R11424 gnd.n4050 gnd.n4049 9.3005
R11425 gnd.n4048 gnd.n2269 9.3005
R11426 gnd.n2268 gnd.n2248 9.3005
R11427 gnd.n4064 gnd.n2249 9.3005
R11428 gnd.n4065 gnd.n2246 9.3005
R11429 gnd.n4067 gnd.n2247 9.3005
R11430 gnd.n4069 gnd.n4068 9.3005
R11431 gnd.n4070 gnd.n2222 9.3005
R11432 gnd.n4101 gnd.n2223 9.3005
R11433 gnd.n4102 gnd.n2219 9.3005
R11434 gnd.n4104 gnd.n2220 9.3005
R11435 gnd.n4108 gnd.n4107 9.3005
R11436 gnd.n4106 gnd.n2221 9.3005
R11437 gnd.n2198 gnd.n2196 9.3005
R11438 gnd.n4139 gnd.n4138 9.3005
R11439 gnd.n2201 gnd.n2197 9.3005
R11440 gnd.n2200 gnd.n2180 9.3005
R11441 gnd.n4157 gnd.n2179 9.3005
R11442 gnd.n4159 gnd.n4158 9.3005
R11443 gnd.n4160 gnd.n960 9.3005
R11444 gnd.n4182 gnd.n961 9.3005
R11445 gnd.n4181 gnd.n962 9.3005
R11446 gnd.n4180 gnd.n4161 9.3005
R11447 gnd.n4167 gnd.n4162 9.3005
R11448 gnd.n4166 gnd.n2164 9.3005
R11449 gnd.n4165 gnd.n2165 9.3005
R11450 gnd.n4164 gnd.n2166 9.3005
R11451 gnd.n4163 gnd.n2142 9.3005
R11452 gnd.n4244 gnd.n2141 9.3005
R11453 gnd.n4246 gnd.n4245 9.3005
R11454 gnd.n4247 gnd.n988 9.3005
R11455 gnd.n4250 gnd.n989 9.3005
R11456 gnd.n4251 gnd.n990 9.3005
R11457 gnd.n4256 gnd.n4252 9.3005
R11458 gnd.n4257 gnd.n1007 9.3005
R11459 gnd.n4261 gnd.n1008 9.3005
R11460 gnd.n4260 gnd.n1009 9.3005
R11461 gnd.n4259 gnd.n4258 9.3005
R11462 gnd.n2115 gnd.n1027 9.3005
R11463 gnd.n4326 gnd.n1028 9.3005
R11464 gnd.n4327 gnd.n1029 9.3005
R11465 gnd.n4329 gnd.n4328 9.3005
R11466 gnd.n2110 gnd.n1047 9.3005
R11467 gnd.n4341 gnd.n1048 9.3005
R11468 gnd.n4342 gnd.n1049 9.3005
R11469 gnd.n4344 gnd.n4343 9.3005
R11470 gnd.n4345 gnd.n1067 9.3005
R11471 gnd.n4348 gnd.n1068 9.3005
R11472 gnd.n4349 gnd.n1069 9.3005
R11473 gnd.n4353 gnd.n4350 9.3005
R11474 gnd.n4354 gnd.n1088 9.3005
R11475 gnd.n4356 gnd.n1089 9.3005
R11476 gnd.n4355 gnd.n1090 9.3005
R11477 gnd.n4047 gnd.n2266 9.3005
R11478 gnd.n3928 gnd.n3927 9.3005
R11479 gnd.n3930 gnd.n3849 9.3005
R11480 gnd.n3931 gnd.n3848 9.3005
R11481 gnd.n3934 gnd.n3847 9.3005
R11482 gnd.n3935 gnd.n3846 9.3005
R11483 gnd.n3938 gnd.n3845 9.3005
R11484 gnd.n3939 gnd.n3844 9.3005
R11485 gnd.n3942 gnd.n3843 9.3005
R11486 gnd.n3943 gnd.n3842 9.3005
R11487 gnd.n3946 gnd.n3841 9.3005
R11488 gnd.n3947 gnd.n3840 9.3005
R11489 gnd.n3950 gnd.n3839 9.3005
R11490 gnd.n3951 gnd.n3838 9.3005
R11491 gnd.n3954 gnd.n3837 9.3005
R11492 gnd.n3955 gnd.n3836 9.3005
R11493 gnd.n3958 gnd.n3835 9.3005
R11494 gnd.n3959 gnd.n3834 9.3005
R11495 gnd.n3962 gnd.n3833 9.3005
R11496 gnd.n3963 gnd.n3832 9.3005
R11497 gnd.n3966 gnd.n3831 9.3005
R11498 gnd.n3970 gnd.n3827 9.3005
R11499 gnd.n3971 gnd.n3826 9.3005
R11500 gnd.n3974 gnd.n3825 9.3005
R11501 gnd.n3975 gnd.n3824 9.3005
R11502 gnd.n3978 gnd.n3823 9.3005
R11503 gnd.n3979 gnd.n3822 9.3005
R11504 gnd.n3982 gnd.n3821 9.3005
R11505 gnd.n3983 gnd.n3820 9.3005
R11506 gnd.n3986 gnd.n3819 9.3005
R11507 gnd.n3987 gnd.n3818 9.3005
R11508 gnd.n3990 gnd.n3817 9.3005
R11509 gnd.n3991 gnd.n3816 9.3005
R11510 gnd.n3994 gnd.n3815 9.3005
R11511 gnd.n3995 gnd.n3814 9.3005
R11512 gnd.n3998 gnd.n3813 9.3005
R11513 gnd.n3999 gnd.n3812 9.3005
R11514 gnd.n4002 gnd.n3811 9.3005
R11515 gnd.n4003 gnd.n3810 9.3005
R11516 gnd.n4006 gnd.n3809 9.3005
R11517 gnd.n4008 gnd.n3806 9.3005
R11518 gnd.n4011 gnd.n3805 9.3005
R11519 gnd.n4012 gnd.n3804 9.3005
R11520 gnd.n4015 gnd.n3803 9.3005
R11521 gnd.n4016 gnd.n3802 9.3005
R11522 gnd.n4019 gnd.n3801 9.3005
R11523 gnd.n4020 gnd.n3800 9.3005
R11524 gnd.n4023 gnd.n3799 9.3005
R11525 gnd.n4024 gnd.n3798 9.3005
R11526 gnd.n4027 gnd.n3797 9.3005
R11527 gnd.n4028 gnd.n3796 9.3005
R11528 gnd.n4031 gnd.n3795 9.3005
R11529 gnd.n4032 gnd.n3794 9.3005
R11530 gnd.n4035 gnd.n3793 9.3005
R11531 gnd.n4037 gnd.n3792 9.3005
R11532 gnd.n4038 gnd.n3791 9.3005
R11533 gnd.n4039 gnd.n3790 9.3005
R11534 gnd.n4040 gnd.n3789 9.3005
R11535 gnd.n3967 gnd.n3828 9.3005
R11536 gnd.n3926 gnd.n2270 9.3005
R11537 gnd.n4056 gnd.n4055 9.3005
R11538 gnd.n4057 gnd.n2255 9.3005
R11539 gnd.n4059 gnd.n4058 9.3005
R11540 gnd.n2237 gnd.n2236 9.3005
R11541 gnd.n4080 gnd.n4079 9.3005
R11542 gnd.n4081 gnd.n2235 9.3005
R11543 gnd.n4085 gnd.n4082 9.3005
R11544 gnd.n4084 gnd.n4083 9.3005
R11545 gnd.n2211 gnd.n2210 9.3005
R11546 gnd.n4116 gnd.n4115 9.3005
R11547 gnd.n4117 gnd.n2209 9.3005
R11548 gnd.n4119 gnd.n4118 9.3005
R11549 gnd.n2189 gnd.n2188 9.3005
R11550 gnd.n4146 gnd.n4145 9.3005
R11551 gnd.n4147 gnd.n2187 9.3005
R11552 gnd.n4150 gnd.n4149 9.3005
R11553 gnd.n4148 gnd.n948 9.3005
R11554 gnd.n6464 gnd.n949 9.3005
R11555 gnd.n6463 gnd.n950 9.3005
R11556 gnd.n6462 gnd.n951 9.3005
R11557 gnd.n972 gnd.n952 9.3005
R11558 gnd.n979 gnd.n971 9.3005
R11559 gnd.n6439 gnd.n997 9.3005
R11560 gnd.n6438 gnd.n998 9.3005
R11561 gnd.n6437 gnd.n999 9.3005
R11562 gnd.n1017 gnd.n1000 9.3005
R11563 gnd.n6427 gnd.n1018 9.3005
R11564 gnd.n6426 gnd.n1019 9.3005
R11565 gnd.n6425 gnd.n1020 9.3005
R11566 gnd.n1036 gnd.n1021 9.3005
R11567 gnd.n6415 gnd.n1037 9.3005
R11568 gnd.n6414 gnd.n1038 9.3005
R11569 gnd.n6413 gnd.n1039 9.3005
R11570 gnd.n1057 gnd.n1040 9.3005
R11571 gnd.n6403 gnd.n1058 9.3005
R11572 gnd.n6402 gnd.n1059 9.3005
R11573 gnd.n6401 gnd.n1060 9.3005
R11574 gnd.n1077 gnd.n1061 9.3005
R11575 gnd.n6391 gnd.n1078 9.3005
R11576 gnd.n6390 gnd.n1079 9.3005
R11577 gnd.n6389 gnd.n1080 9.3005
R11578 gnd.n1097 gnd.n1081 9.3005
R11579 gnd.n6379 gnd.n6378 9.3005
R11580 gnd.n2257 gnd.n2256 9.3005
R11581 gnd.n6450 gnd.n977 9.3005
R11582 gnd.n6450 gnd.n6449 9.3005
R11583 gnd.n939 gnd.n938 9.3005
R11584 gnd.n4194 gnd.n4193 9.3005
R11585 gnd.n4197 gnd.n4196 9.3005
R11586 gnd.n4195 gnd.n2172 9.3005
R11587 gnd.n6470 gnd.n6469 9.3005
R11588 gnd.n6473 gnd.n937 9.3005
R11589 gnd.n936 gnd.n932 9.3005
R11590 gnd.n6479 gnd.n931 9.3005
R11591 gnd.n6480 gnd.n930 9.3005
R11592 gnd.n6481 gnd.n929 9.3005
R11593 gnd.n928 gnd.n924 9.3005
R11594 gnd.n6487 gnd.n923 9.3005
R11595 gnd.n6488 gnd.n922 9.3005
R11596 gnd.n6489 gnd.n921 9.3005
R11597 gnd.n920 gnd.n916 9.3005
R11598 gnd.n6495 gnd.n915 9.3005
R11599 gnd.n6496 gnd.n914 9.3005
R11600 gnd.n6497 gnd.n913 9.3005
R11601 gnd.n912 gnd.n908 9.3005
R11602 gnd.n6503 gnd.n907 9.3005
R11603 gnd.n6504 gnd.n906 9.3005
R11604 gnd.n6505 gnd.n905 9.3005
R11605 gnd.n904 gnd.n900 9.3005
R11606 gnd.n6511 gnd.n899 9.3005
R11607 gnd.n6512 gnd.n898 9.3005
R11608 gnd.n6513 gnd.n897 9.3005
R11609 gnd.n896 gnd.n892 9.3005
R11610 gnd.n6519 gnd.n891 9.3005
R11611 gnd.n6520 gnd.n890 9.3005
R11612 gnd.n6521 gnd.n889 9.3005
R11613 gnd.n888 gnd.n884 9.3005
R11614 gnd.n6527 gnd.n883 9.3005
R11615 gnd.n6528 gnd.n882 9.3005
R11616 gnd.n6529 gnd.n881 9.3005
R11617 gnd.n880 gnd.n876 9.3005
R11618 gnd.n6535 gnd.n875 9.3005
R11619 gnd.n6536 gnd.n874 9.3005
R11620 gnd.n6537 gnd.n873 9.3005
R11621 gnd.n872 gnd.n868 9.3005
R11622 gnd.n6543 gnd.n867 9.3005
R11623 gnd.n6544 gnd.n866 9.3005
R11624 gnd.n6545 gnd.n865 9.3005
R11625 gnd.n864 gnd.n860 9.3005
R11626 gnd.n6551 gnd.n859 9.3005
R11627 gnd.n6552 gnd.n858 9.3005
R11628 gnd.n6553 gnd.n857 9.3005
R11629 gnd.n856 gnd.n852 9.3005
R11630 gnd.n6559 gnd.n851 9.3005
R11631 gnd.n6560 gnd.n850 9.3005
R11632 gnd.n6561 gnd.n849 9.3005
R11633 gnd.n848 gnd.n844 9.3005
R11634 gnd.n6567 gnd.n843 9.3005
R11635 gnd.n6568 gnd.n842 9.3005
R11636 gnd.n6569 gnd.n841 9.3005
R11637 gnd.n840 gnd.n836 9.3005
R11638 gnd.n6575 gnd.n835 9.3005
R11639 gnd.n6576 gnd.n834 9.3005
R11640 gnd.n6577 gnd.n833 9.3005
R11641 gnd.n832 gnd.n828 9.3005
R11642 gnd.n6583 gnd.n827 9.3005
R11643 gnd.n6584 gnd.n826 9.3005
R11644 gnd.n6585 gnd.n825 9.3005
R11645 gnd.n824 gnd.n820 9.3005
R11646 gnd.n6591 gnd.n819 9.3005
R11647 gnd.n6592 gnd.n818 9.3005
R11648 gnd.n6593 gnd.n817 9.3005
R11649 gnd.n816 gnd.n812 9.3005
R11650 gnd.n6599 gnd.n811 9.3005
R11651 gnd.n6600 gnd.n810 9.3005
R11652 gnd.n6601 gnd.n809 9.3005
R11653 gnd.n808 gnd.n804 9.3005
R11654 gnd.n6607 gnd.n803 9.3005
R11655 gnd.n6608 gnd.n802 9.3005
R11656 gnd.n6609 gnd.n801 9.3005
R11657 gnd.n800 gnd.n796 9.3005
R11658 gnd.n6615 gnd.n795 9.3005
R11659 gnd.n6616 gnd.n794 9.3005
R11660 gnd.n6617 gnd.n793 9.3005
R11661 gnd.n792 gnd.n788 9.3005
R11662 gnd.n6623 gnd.n787 9.3005
R11663 gnd.n6624 gnd.n786 9.3005
R11664 gnd.n6625 gnd.n785 9.3005
R11665 gnd.n784 gnd.n780 9.3005
R11666 gnd.n6631 gnd.n779 9.3005
R11667 gnd.n6632 gnd.n778 9.3005
R11668 gnd.n6633 gnd.n777 9.3005
R11669 gnd.n776 gnd.n772 9.3005
R11670 gnd.n6639 gnd.n771 9.3005
R11671 gnd.n6641 gnd.n6640 9.3005
R11672 gnd.n6472 gnd.n6471 9.3005
R11673 gnd.n5536 gnd.n5535 9.3005
R11674 gnd.n4672 gnd.n2070 9.3005
R11675 gnd.n2048 gnd.n2047 9.3005
R11676 gnd.n4700 gnd.n4699 9.3005
R11677 gnd.n4701 gnd.n2045 9.3005
R11678 gnd.n4706 gnd.n4705 9.3005
R11679 gnd.n4704 gnd.n2046 9.3005
R11680 gnd.n4703 gnd.n4702 9.3005
R11681 gnd.n1947 gnd.n1946 9.3005
R11682 gnd.n4737 gnd.n4736 9.3005
R11683 gnd.n4738 gnd.n1944 9.3005
R11684 gnd.n4741 gnd.n4740 9.3005
R11685 gnd.n4739 gnd.n1945 9.3005
R11686 gnd.n1936 gnd.n1935 9.3005
R11687 gnd.n4762 gnd.n4761 9.3005
R11688 gnd.n4763 gnd.n1933 9.3005
R11689 gnd.n4772 gnd.n4771 9.3005
R11690 gnd.n4770 gnd.n1934 9.3005
R11691 gnd.n4769 gnd.n4768 9.3005
R11692 gnd.n4767 gnd.n4764 9.3005
R11693 gnd.n1889 gnd.n1888 9.3005
R11694 gnd.n4848 gnd.n4847 9.3005
R11695 gnd.n4849 gnd.n1886 9.3005
R11696 gnd.n4870 gnd.n4869 9.3005
R11697 gnd.n4868 gnd.n1887 9.3005
R11698 gnd.n4867 gnd.n4866 9.3005
R11699 gnd.n4865 gnd.n4850 9.3005
R11700 gnd.n4864 gnd.n4863 9.3005
R11701 gnd.n4862 gnd.n4856 9.3005
R11702 gnd.n4861 gnd.n4860 9.3005
R11703 gnd.n4859 gnd.n4858 9.3005
R11704 gnd.n4857 gnd.n1839 9.3005
R11705 gnd.n1837 gnd.n1836 9.3005
R11706 gnd.n4950 gnd.n4949 9.3005
R11707 gnd.n4951 gnd.n1835 9.3005
R11708 gnd.n4953 gnd.n4952 9.3005
R11709 gnd.n1812 gnd.n1810 9.3005
R11710 gnd.n4999 gnd.n4998 9.3005
R11711 gnd.n4997 gnd.n1811 9.3005
R11712 gnd.n4996 gnd.n4995 9.3005
R11713 gnd.n1789 gnd.n1787 9.3005
R11714 gnd.n5058 gnd.n5057 9.3005
R11715 gnd.n5056 gnd.n1788 9.3005
R11716 gnd.n5055 gnd.n5054 9.3005
R11717 gnd.n5053 gnd.n1790 9.3005
R11718 gnd.n5052 gnd.n5051 9.3005
R11719 gnd.n5050 gnd.n5038 9.3005
R11720 gnd.n5049 gnd.n5048 9.3005
R11721 gnd.n5047 gnd.n5039 9.3005
R11722 gnd.n5046 gnd.n5045 9.3005
R11723 gnd.n1728 gnd.n1727 9.3005
R11724 gnd.n5167 gnd.n5166 9.3005
R11725 gnd.n5168 gnd.n1725 9.3005
R11726 gnd.n5171 gnd.n5170 9.3005
R11727 gnd.n5169 gnd.n1726 9.3005
R11728 gnd.n1699 gnd.n1698 9.3005
R11729 gnd.n5206 gnd.n5205 9.3005
R11730 gnd.n5207 gnd.n1696 9.3005
R11731 gnd.n5224 gnd.n5223 9.3005
R11732 gnd.n5222 gnd.n1697 9.3005
R11733 gnd.n5221 gnd.n5220 9.3005
R11734 gnd.n5219 gnd.n5208 9.3005
R11735 gnd.n5218 gnd.n5217 9.3005
R11736 gnd.n5216 gnd.n5213 9.3005
R11737 gnd.n5215 gnd.n5214 9.3005
R11738 gnd.n1643 gnd.n1642 9.3005
R11739 gnd.n5297 gnd.n5296 9.3005
R11740 gnd.n5298 gnd.n1640 9.3005
R11741 gnd.n5301 gnd.n5300 9.3005
R11742 gnd.n5299 gnd.n1641 9.3005
R11743 gnd.n1616 gnd.n1615 9.3005
R11744 gnd.n5339 gnd.n5338 9.3005
R11745 gnd.n5340 gnd.n1614 9.3005
R11746 gnd.n5342 gnd.n5341 9.3005
R11747 gnd.n1613 gnd.n1612 9.3005
R11748 gnd.n5350 gnd.n5349 9.3005
R11749 gnd.n5351 gnd.n1611 9.3005
R11750 gnd.n5353 gnd.n5352 9.3005
R11751 gnd.n5354 gnd.n1610 9.3005
R11752 gnd.n5358 gnd.n5357 9.3005
R11753 gnd.n5359 gnd.n1608 9.3005
R11754 gnd.n5539 gnd.n5538 9.3005
R11755 gnd.n5537 gnd.n1609 9.3005
R11756 gnd.n4674 gnd.n4673 9.3005
R11757 gnd.n4671 gnd.n4670 9.3005
R11758 gnd.n4232 gnd.n2150 9.3005
R11759 gnd.n4234 gnd.n4233 9.3005
R11760 gnd.n2136 gnd.n2134 9.3005
R11761 gnd.n4275 gnd.n4274 9.3005
R11762 gnd.n4273 gnd.n2135 9.3005
R11763 gnd.n4272 gnd.n4271 9.3005
R11764 gnd.n4270 gnd.n2137 9.3005
R11765 gnd.n4269 gnd.n4268 9.3005
R11766 gnd.n4267 gnd.n2140 9.3005
R11767 gnd.n4266 gnd.n4265 9.3005
R11768 gnd.n2118 gnd.n2117 9.3005
R11769 gnd.n4319 gnd.n4318 9.3005
R11770 gnd.n4320 gnd.n2116 9.3005
R11771 gnd.n4322 gnd.n4321 9.3005
R11772 gnd.n2113 gnd.n2112 9.3005
R11773 gnd.n4334 gnd.n4333 9.3005
R11774 gnd.n4335 gnd.n2111 9.3005
R11775 gnd.n4337 gnd.n4336 9.3005
R11776 gnd.n2104 gnd.n2102 9.3005
R11777 gnd.n4371 gnd.n4370 9.3005
R11778 gnd.n4369 gnd.n2103 9.3005
R11779 gnd.n4368 gnd.n4367 9.3005
R11780 gnd.n4366 gnd.n2105 9.3005
R11781 gnd.n4365 gnd.n4364 9.3005
R11782 gnd.n4363 gnd.n2108 9.3005
R11783 gnd.n4362 gnd.n4361 9.3005
R11784 gnd.n4360 gnd.n2109 9.3005
R11785 gnd.n4636 gnd.n4635 9.3005
R11786 gnd.n4634 gnd.n4633 9.3005
R11787 gnd.n4549 gnd.n4548 9.3005
R11788 gnd.n4628 gnd.n4627 9.3005
R11789 gnd.n4626 gnd.n4625 9.3005
R11790 gnd.n4561 gnd.n4560 9.3005
R11791 gnd.n4620 gnd.n4619 9.3005
R11792 gnd.n4618 gnd.n4617 9.3005
R11793 gnd.n4572 gnd.n4571 9.3005
R11794 gnd.n4612 gnd.n4611 9.3005
R11795 gnd.n4610 gnd.n4609 9.3005
R11796 gnd.n4584 gnd.n4583 9.3005
R11797 gnd.n4604 gnd.n4603 9.3005
R11798 gnd.n4602 gnd.n4601 9.3005
R11799 gnd.n4595 gnd.n2079 9.3005
R11800 gnd.n4661 gnd.n4660 9.3005
R11801 gnd.n2081 gnd.n2077 9.3005
R11802 gnd.n4667 gnd.n4666 9.3005
R11803 gnd.n4544 gnd.n4542 9.3005
R11804 gnd.n4669 gnd.n4668 9.3005
R11805 gnd.n2074 gnd.n2072 9.3005
R11806 gnd.n4659 gnd.n4658 9.3005
R11807 gnd.n4598 gnd.n2080 9.3005
R11808 gnd.n4600 gnd.n4599 9.3005
R11809 gnd.n4588 gnd.n4587 9.3005
R11810 gnd.n4606 gnd.n4605 9.3005
R11811 gnd.n4608 gnd.n4607 9.3005
R11812 gnd.n4578 gnd.n4577 9.3005
R11813 gnd.n4614 gnd.n4613 9.3005
R11814 gnd.n4616 gnd.n4615 9.3005
R11815 gnd.n4565 gnd.n4564 9.3005
R11816 gnd.n4622 gnd.n4621 9.3005
R11817 gnd.n4624 gnd.n4623 9.3005
R11818 gnd.n4555 gnd.n4554 9.3005
R11819 gnd.n4630 gnd.n4629 9.3005
R11820 gnd.n4632 gnd.n4631 9.3005
R11821 gnd.n4543 gnd.n4541 9.3005
R11822 gnd.n4638 gnd.n4637 9.3005
R11823 gnd.n4639 gnd.n4536 9.3005
R11824 gnd.n4641 gnd.n4640 9.3005
R11825 gnd.n4643 gnd.n4422 9.3005
R11826 gnd.n4645 gnd.n4644 9.3005
R11827 gnd.n4646 gnd.n4418 9.3005
R11828 gnd.n4648 gnd.n4647 9.3005
R11829 gnd.n4649 gnd.n4417 9.3005
R11830 gnd.n4651 gnd.n4650 9.3005
R11831 gnd.n4652 gnd.n4416 9.3005
R11832 gnd.n4691 gnd.n4690 9.3005
R11833 gnd.n4692 gnd.n2054 9.3005
R11834 gnd.n4695 gnd.n4694 9.3005
R11835 gnd.n4693 gnd.n2055 9.3005
R11836 gnd.n2033 gnd.n2032 9.3005
R11837 gnd.n4724 gnd.n4723 9.3005
R11838 gnd.n4725 gnd.n2030 9.3005
R11839 gnd.n4731 gnd.n4730 9.3005
R11840 gnd.n4729 gnd.n2031 9.3005
R11841 gnd.n4728 gnd.n4727 9.3005
R11842 gnd.n1228 gnd.n1226 9.3005
R11843 gnd.n6246 gnd.n6245 9.3005
R11844 gnd.n6244 gnd.n1227 9.3005
R11845 gnd.n6243 gnd.n6242 9.3005
R11846 gnd.n6241 gnd.n1229 9.3005
R11847 gnd.n6240 gnd.n6239 9.3005
R11848 gnd.n6238 gnd.n1233 9.3005
R11849 gnd.n6237 gnd.n6236 9.3005
R11850 gnd.n6235 gnd.n1234 9.3005
R11851 gnd.n6234 gnd.n6233 9.3005
R11852 gnd.n6232 gnd.n1238 9.3005
R11853 gnd.n6231 gnd.n6230 9.3005
R11854 gnd.n6229 gnd.n1239 9.3005
R11855 gnd.n6228 gnd.n6227 9.3005
R11856 gnd.n6226 gnd.n1243 9.3005
R11857 gnd.n6225 gnd.n6224 9.3005
R11858 gnd.n6223 gnd.n1244 9.3005
R11859 gnd.n6222 gnd.n6221 9.3005
R11860 gnd.n6220 gnd.n1248 9.3005
R11861 gnd.n6219 gnd.n6218 9.3005
R11862 gnd.n6217 gnd.n1249 9.3005
R11863 gnd.n6216 gnd.n6215 9.3005
R11864 gnd.n6214 gnd.n1253 9.3005
R11865 gnd.n6213 gnd.n6212 9.3005
R11866 gnd.n6211 gnd.n1254 9.3005
R11867 gnd.n6210 gnd.n6209 9.3005
R11868 gnd.n6208 gnd.n1258 9.3005
R11869 gnd.n6207 gnd.n6206 9.3005
R11870 gnd.n6205 gnd.n1259 9.3005
R11871 gnd.n6204 gnd.n6203 9.3005
R11872 gnd.n6202 gnd.n1263 9.3005
R11873 gnd.n6201 gnd.n6200 9.3005
R11874 gnd.n6199 gnd.n1264 9.3005
R11875 gnd.n6198 gnd.n6197 9.3005
R11876 gnd.n6196 gnd.n1268 9.3005
R11877 gnd.n6195 gnd.n6194 9.3005
R11878 gnd.n6193 gnd.n1269 9.3005
R11879 gnd.n6192 gnd.n6191 9.3005
R11880 gnd.n6190 gnd.n1273 9.3005
R11881 gnd.n6189 gnd.n6188 9.3005
R11882 gnd.n6187 gnd.n1274 9.3005
R11883 gnd.n6186 gnd.n6185 9.3005
R11884 gnd.n6184 gnd.n1278 9.3005
R11885 gnd.n6183 gnd.n6182 9.3005
R11886 gnd.n6181 gnd.n1279 9.3005
R11887 gnd.n6180 gnd.n6179 9.3005
R11888 gnd.n6178 gnd.n1283 9.3005
R11889 gnd.n6177 gnd.n6176 9.3005
R11890 gnd.n6175 gnd.n1284 9.3005
R11891 gnd.n6174 gnd.n6173 9.3005
R11892 gnd.n6172 gnd.n1288 9.3005
R11893 gnd.n6171 gnd.n6170 9.3005
R11894 gnd.n6169 gnd.n1289 9.3005
R11895 gnd.n6168 gnd.n6167 9.3005
R11896 gnd.n6166 gnd.n1293 9.3005
R11897 gnd.n6165 gnd.n6164 9.3005
R11898 gnd.n6163 gnd.n1294 9.3005
R11899 gnd.n6162 gnd.n6161 9.3005
R11900 gnd.n6160 gnd.n1298 9.3005
R11901 gnd.n6159 gnd.n6158 9.3005
R11902 gnd.n6157 gnd.n1299 9.3005
R11903 gnd.n6156 gnd.n6155 9.3005
R11904 gnd.n6154 gnd.n1303 9.3005
R11905 gnd.n6153 gnd.n6152 9.3005
R11906 gnd.n6151 gnd.n1304 9.3005
R11907 gnd.n6150 gnd.n6149 9.3005
R11908 gnd.n6148 gnd.n1308 9.3005
R11909 gnd.n6147 gnd.n6146 9.3005
R11910 gnd.n6145 gnd.n1309 9.3005
R11911 gnd.n6144 gnd.n6143 9.3005
R11912 gnd.n6142 gnd.n1313 9.3005
R11913 gnd.n6141 gnd.n6140 9.3005
R11914 gnd.n2057 gnd.n2056 9.3005
R11915 gnd.n5425 gnd.n5424 9.3005
R11916 gnd.n5421 gnd.n5420 9.3005
R11917 gnd.n5432 gnd.n5431 9.3005
R11918 gnd.n5433 gnd.n5419 9.3005
R11919 gnd.n5436 gnd.n5435 9.3005
R11920 gnd.n5434 gnd.n5417 9.3005
R11921 gnd.n5423 gnd.n1314 9.3005
R11922 gnd.n5524 gnd.n5373 9.3005
R11923 gnd.n5386 gnd.n5382 9.3005
R11924 gnd.n5518 gnd.n5517 9.3005
R11925 gnd.n5506 gnd.n5384 9.3005
R11926 gnd.n5505 gnd.n5504 9.3005
R11927 gnd.n5395 gnd.n5391 9.3005
R11928 gnd.n5498 gnd.n5497 9.3005
R11929 gnd.n5487 gnd.n5393 9.3005
R11930 gnd.n5486 gnd.n5485 9.3005
R11931 gnd.n5404 gnd.n5400 9.3005
R11932 gnd.n5479 gnd.n5478 9.3005
R11933 gnd.n5468 gnd.n5402 9.3005
R11934 gnd.n5467 gnd.n5466 9.3005
R11935 gnd.n5413 gnd.n5409 9.3005
R11936 gnd.n5460 gnd.n5459 9.3005
R11937 gnd.n5449 gnd.n5411 9.3005
R11938 gnd.n5448 gnd.n5447 9.3005
R11939 gnd.n5526 gnd.n5525 9.3005
R11940 gnd.n5377 gnd.n5376 9.3005
R11941 gnd.n5443 gnd.n5442 9.3005
R11942 gnd.n5444 gnd.n5416 9.3005
R11943 gnd.n5451 gnd.n5450 9.3005
R11944 gnd.n5414 gnd.n5412 9.3005
R11945 gnd.n5458 gnd.n5457 9.3005
R11946 gnd.n5408 gnd.n5407 9.3005
R11947 gnd.n5470 gnd.n5469 9.3005
R11948 gnd.n5405 gnd.n5403 9.3005
R11949 gnd.n5477 gnd.n5476 9.3005
R11950 gnd.n5399 gnd.n5398 9.3005
R11951 gnd.n5489 gnd.n5488 9.3005
R11952 gnd.n5396 gnd.n5394 9.3005
R11953 gnd.n5496 gnd.n5495 9.3005
R11954 gnd.n5390 gnd.n5389 9.3005
R11955 gnd.n5508 gnd.n5507 9.3005
R11956 gnd.n5387 gnd.n5385 9.3005
R11957 gnd.n5516 gnd.n5515 9.3005
R11958 gnd.n5514 gnd.n5513 9.3005
R11959 gnd.n5528 gnd.n5527 9.3005
R11960 gnd.n5374 gnd.n5368 9.3005
R11961 gnd.n5375 gnd.n5367 9.3005
R11962 gnd.n5363 gnd.n5360 9.3005
R11963 gnd.n1495 gnd.n1494 9.3005
R11964 gnd.n5912 gnd.n5911 9.3005
R11965 gnd.n5913 gnd.n1493 9.3005
R11966 gnd.n5915 gnd.n5914 9.3005
R11967 gnd.n1490 gnd.n1488 9.3005
R11968 gnd.n5934 gnd.n5933 9.3005
R11969 gnd.n5932 gnd.n1489 9.3005
R11970 gnd.n5931 gnd.n5930 9.3005
R11971 gnd.n1480 gnd.n1479 9.3005
R11972 gnd.n5993 gnd.n5992 9.3005
R11973 gnd.n5994 gnd.n1478 9.3005
R11974 gnd.n5996 gnd.n5995 9.3005
R11975 gnd.n1474 gnd.n1473 9.3005
R11976 gnd.n6007 gnd.n6006 9.3005
R11977 gnd.n6008 gnd.n1472 9.3005
R11978 gnd.n6010 gnd.n6009 9.3005
R11979 gnd.n1468 gnd.n1466 9.3005
R11980 gnd.n6035 gnd.n6034 9.3005
R11981 gnd.n6033 gnd.n1467 9.3005
R11982 gnd.n6032 gnd.n6031 9.3005
R11983 gnd.n6030 gnd.n1469 9.3005
R11984 gnd.n6029 gnd.n6028 9.3005
R11985 gnd.n6027 gnd.n6024 9.3005
R11986 gnd.n6026 gnd.n6025 9.3005
R11987 gnd.n81 gnd.n79 9.3005
R11988 gnd.n5365 gnd.n5364 9.3005
R11989 gnd.t106 gnd.n2462 9.24152
R11990 gnd.n2364 gnd.t133 9.24152
R11991 gnd.n3648 gnd.t234 9.24152
R11992 gnd.t145 gnd.n2251 9.24152
R11993 gnd.n4374 gnd.t79 9.24152
R11994 gnd.n5937 gnd.t12 9.24152
R11995 gnd.n7570 gnd.t156 9.24152
R11996 gnd.t77 gnd.t106 8.92286
R11997 gnd.n6249 gnd.t219 8.92286
R11998 gnd.n4751 gnd.n1937 8.92286
R11999 gnd.t320 gnd.n4776 8.92286
R12000 gnd.n4936 gnd.n1846 8.92286
R12001 gnd.n4981 gnd.n1816 8.92286
R12002 gnd.n5106 gnd.n1749 8.92286
R12003 gnd.n5177 gnd.n5176 8.92286
R12004 gnd.n1654 gnd.t305 8.92286
R12005 gnd.n5317 gnd.n5316 8.92286
R12006 gnd.n5654 gnd.t193 8.92286
R12007 gnd.n3618 gnd.n3593 8.92171
R12008 gnd.n3586 gnd.n3561 8.92171
R12009 gnd.n3554 gnd.n3529 8.92171
R12010 gnd.n3523 gnd.n3498 8.92171
R12011 gnd.n3491 gnd.n3466 8.92171
R12012 gnd.n3459 gnd.n3434 8.92171
R12013 gnd.n3427 gnd.n3402 8.92171
R12014 gnd.n3396 gnd.n3371 8.92171
R12015 gnd.n5586 gnd.n5568 8.72777
R12016 gnd.n3122 gnd.t124 8.60421
R12017 gnd.n2534 gnd.n2518 8.43656
R12018 gnd.n46 gnd.n30 8.43656
R12019 gnd.n4911 gnd.n1861 8.28555
R12020 gnd.n5002 gnd.n1799 8.28555
R12021 gnd.n5086 gnd.n1764 8.28555
R12022 gnd.n5142 gnd.n1716 8.28555
R12023 gnd.n3619 gnd.n3591 8.14595
R12024 gnd.n3587 gnd.n3559 8.14595
R12025 gnd.n3555 gnd.n3527 8.14595
R12026 gnd.n3524 gnd.n3496 8.14595
R12027 gnd.n3492 gnd.n3464 8.14595
R12028 gnd.n3460 gnd.n3432 8.14595
R12029 gnd.n3428 gnd.n3400 8.14595
R12030 gnd.n3397 gnd.n3369 8.14595
R12031 gnd.n4231 gnd.n0 8.10675
R12032 gnd.n7644 gnd.n7643 8.10675
R12033 gnd.n3624 gnd.n3623 7.97301
R12034 gnd.t104 gnd.n2637 7.9669
R12035 gnd.n7644 gnd.n78 7.86902
R12036 gnd.n5525 gnd.n5377 7.75808
R12037 gnd.n4666 gnd.n2077 7.75808
R12038 gnd.n7420 gnd.n347 7.75808
R12039 gnd.n3886 gnd.n3870 7.75808
R12040 gnd.n4744 gnd.n1941 7.64824
R12041 gnd.n4911 gnd.n1860 7.64824
R12042 gnd.t32 gnd.n4955 7.64824
R12043 gnd.n5003 gnd.t338 7.64824
R12044 gnd.n5013 gnd.n1799 7.64824
R12045 gnd.n5086 gnd.n1762 7.64824
R12046 gnd.t33 gnd.n1757 7.64824
R12047 gnd.n5105 gnd.t335 7.64824
R12048 gnd.n5142 gnd.n1707 7.64824
R12049 gnd.n2567 gnd.n2566 7.53171
R12050 gnd.n3031 gnd.t110 7.32958
R12051 gnd.n4744 gnd.t10 7.32958
R12052 gnd.t286 gnd.n5335 7.32958
R12053 gnd.n1206 gnd.n1205 7.30353
R12054 gnd.n5585 gnd.n5584 7.30353
R12055 gnd.n2991 gnd.n2710 7.01093
R12056 gnd.n2713 gnd.n2711 7.01093
R12057 gnd.n3001 gnd.n3000 7.01093
R12058 gnd.n3012 gnd.n2694 7.01093
R12059 gnd.n3011 gnd.n2697 7.01093
R12060 gnd.n3022 gnd.n2685 7.01093
R12061 gnd.n2688 gnd.n2686 7.01093
R12062 gnd.n3032 gnd.n3031 7.01093
R12063 gnd.n3042 gnd.n2666 7.01093
R12064 gnd.n3041 gnd.n2669 7.01093
R12065 gnd.n3050 gnd.n2660 7.01093
R12066 gnd.n3062 gnd.n2650 7.01093
R12067 gnd.n3072 gnd.n2635 7.01093
R12068 gnd.n3088 gnd.n3087 7.01093
R12069 gnd.n2637 gnd.n2574 7.01093
R12070 gnd.n3142 gnd.n2575 7.01093
R12071 gnd.n3136 gnd.n3135 7.01093
R12072 gnd.n2624 gnd.n2586 7.01093
R12073 gnd.n3128 gnd.n2597 7.01093
R12074 gnd.n2615 gnd.n2610 7.01093
R12075 gnd.n3122 gnd.n3121 7.01093
R12076 gnd.n3168 gnd.n2497 7.01093
R12077 gnd.n3167 gnd.n3166 7.01093
R12078 gnd.n3179 gnd.n3178 7.01093
R12079 gnd.n2490 gnd.n2482 7.01093
R12080 gnd.n3208 gnd.n2470 7.01093
R12081 gnd.n3207 gnd.n2473 7.01093
R12082 gnd.n3218 gnd.n2462 7.01093
R12083 gnd.n2463 gnd.n2451 7.01093
R12084 gnd.n3229 gnd.n2452 7.01093
R12085 gnd.n3253 gnd.n2443 7.01093
R12086 gnd.n3252 gnd.n2434 7.01093
R12087 gnd.n3275 gnd.n3274 7.01093
R12088 gnd.n3293 gnd.n2415 7.01093
R12089 gnd.n3292 gnd.n2418 7.01093
R12090 gnd.n3303 gnd.n2407 7.01093
R12091 gnd.n2408 gnd.n2395 7.01093
R12092 gnd.n3314 gnd.n2396 7.01093
R12093 gnd.n3341 gnd.n2380 7.01093
R12094 gnd.n3353 gnd.n3352 7.01093
R12095 gnd.n3335 gnd.n2373 7.01093
R12096 gnd.n3364 gnd.n3363 7.01093
R12097 gnd.n3636 gnd.n2361 7.01093
R12098 gnd.n3635 gnd.n2364 7.01093
R12099 gnd.n3648 gnd.n2353 7.01093
R12100 gnd.n2354 gnd.n2346 7.01093
R12101 gnd.n3658 gnd.n2272 7.01093
R12102 gnd.n4758 gnd.n4751 7.01093
R12103 gnd.n4817 gnd.n1906 7.01093
R12104 gnd.t34 gnd.n4816 7.01093
R12105 gnd.n4936 gnd.n4935 7.01093
R12106 gnd.n4956 gnd.t32 7.01093
R12107 gnd.n4955 gnd.n1816 7.01093
R12108 gnd.n5106 gnd.n5105 7.01093
R12109 gnd.t335 gnd.n5104 7.01093
R12110 gnd.n5177 gnd.n1720 7.01093
R12111 gnd.n5258 gnd.t340 7.01093
R12112 gnd.n5274 gnd.n5273 7.01093
R12113 gnd.n5319 gnd.n5317 7.01093
R12114 gnd.n2669 gnd.t127 6.69227
R12115 gnd.n2473 gnd.t77 6.69227
R12116 gnd.n4099 gnd.t90 6.69227
R12117 gnd.n4136 gnd.n2183 6.69227
R12118 gnd.n4339 gnd.t258 6.69227
R12119 gnd.t354 gnd.n1901 6.69227
R12120 gnd.n5211 gnd.t360 6.69227
R12121 gnd.n5928 gnd.t19 6.69227
R12122 gnd.n7385 gnd.n135 6.69227
R12123 gnd.n170 gnd.t4 6.69227
R12124 gnd.n5715 gnd.n5714 6.5566
R12125 gnd.n1956 gnd.n1955 6.5566
R12126 gnd.n6267 gnd.n6263 6.5566
R12127 gnd.n5593 gnd.n5592 6.5566
R12128 gnd.n2027 gnd.n2026 6.37362
R12129 gnd.t219 gnd.t199 6.37362
R12130 gnd.n4878 gnd.n1875 6.37362
R12131 gnd.n4963 gnd.t82 6.37362
R12132 gnd.n5021 gnd.n1793 6.37362
R12133 gnd.n5033 gnd.n1780 6.37362
R12134 gnd.n5155 gnd.t52 6.37362
R12135 gnd.n5202 gnd.n1703 6.37362
R12136 gnd.n5316 gnd.t130 6.37362
R12137 gnd.n5327 gnd.t130 6.37362
R12138 gnd.n5654 gnd.n1573 6.37362
R12139 gnd.n4658 gnd.n2084 6.20656
R12140 gnd.n5528 gnd.n5372 6.20656
R12141 gnd.t272 gnd.n3098 6.05496
R12142 gnd.n3099 gnd.t128 6.05496
R12143 gnd.t288 gnd.n2497 6.05496
R12144 gnd.t113 gnd.n3263 6.05496
R12145 gnd.n4263 gnd.t17 6.05496
R12146 gnd.t53 gnd.t364 6.05496
R12147 gnd.t313 gnd.t290 6.05496
R12148 gnd.n6012 gnd.t58 6.05496
R12149 gnd.n3621 gnd.n3591 5.81868
R12150 gnd.n3589 gnd.n3559 5.81868
R12151 gnd.n3557 gnd.n3527 5.81868
R12152 gnd.n3526 gnd.n3496 5.81868
R12153 gnd.n3494 gnd.n3464 5.81868
R12154 gnd.n3462 gnd.n3432 5.81868
R12155 gnd.n3430 gnd.n3400 5.81868
R12156 gnd.n3399 gnd.n3369 5.81868
R12157 gnd.n1930 gnd.n1929 5.73631
R12158 gnd.n4777 gnd.n4774 5.73631
R12159 gnd.n1841 gnd.n1829 5.73631
R12160 gnd.n4947 gnd.n1822 5.73631
R12161 gnd.t338 gnd.n5002 5.73631
R12162 gnd.n1764 gnd.t33 5.73631
R12163 gnd.n5043 gnd.n5041 5.73631
R12164 gnd.n5113 gnd.n1738 5.73631
R12165 gnd.n5294 gnd.n1645 5.73631
R12166 gnd.n1647 gnd.n1637 5.73631
R12167 gnd.n5724 gnd.n1532 5.62001
R12168 gnd.n6329 gnd.n1148 5.62001
R12169 gnd.n6329 gnd.n1149 5.62001
R12170 gnd.n5724 gnd.n1533 5.62001
R12171 gnd.n2850 gnd.n2845 5.4308
R12172 gnd.n3666 gnd.n2339 5.4308
R12173 gnd.n3166 gnd.t103 5.41765
R12174 gnd.t111 gnd.n3189 5.41765
R12175 gnd.t67 gnd.n2427 5.41765
R12176 gnd.n4236 gnd.t72 5.41765
R12177 gnd.t292 gnd.n4894 5.41765
R12178 gnd.n5134 gnd.t28 5.41765
R12179 gnd.n7304 gnd.t2 5.41765
R12180 gnd.n6467 gnd.n941 5.09899
R12181 gnd.n6466 gnd.n944 5.09899
R12182 gnd.n4191 gnd.n4190 5.09899
R12183 gnd.n6460 gnd.n956 5.09899
R12184 gnd.n4184 gnd.n965 5.09899
R12185 gnd.n6454 gnd.n968 5.09899
R12186 gnd.n4178 gnd.n4177 5.09899
R12187 gnd.n4176 gnd.n2159 5.09899
R12188 gnd.n4222 gnd.n2161 5.09899
R12189 gnd.n4227 gnd.n2155 5.09899
R12190 gnd.n4216 gnd.n4215 5.09899
R12191 gnd.n4236 gnd.n2145 5.09899
R12192 gnd.n4241 gnd.n2131 5.09899
R12193 gnd.n4278 gnd.n4277 5.09899
R12194 gnd.n6447 gnd.n984 5.09899
R12195 gnd.n4248 gnd.n993 5.09899
R12196 gnd.n4254 gnd.n1002 5.09899
R12197 gnd.n6435 gnd.n1005 5.09899
R12198 gnd.n4263 gnd.n1012 5.09899
R12199 gnd.n6429 gnd.n1015 5.09899
R12200 gnd.n4316 gnd.n4315 5.09899
R12201 gnd.n6423 gnd.n1025 5.09899
R12202 gnd.n4324 gnd.n1032 5.09899
R12203 gnd.n4331 gnd.n1042 5.09899
R12204 gnd.n6411 gnd.n1045 5.09899
R12205 gnd.n4339 gnd.n1052 5.09899
R12206 gnd.n6405 gnd.n1055 5.09899
R12207 gnd.n4374 gnd.n4373 5.09899
R12208 gnd.n6399 gnd.n1065 5.09899
R12209 gnd.n4346 gnd.n1072 5.09899
R12210 gnd.n6393 gnd.n1075 5.09899
R12211 gnd.n4351 gnd.n1083 5.09899
R12212 gnd.n6387 gnd.n1086 5.09899
R12213 gnd.n4358 gnd.n1092 5.09899
R12214 gnd.n6381 gnd.n1095 5.09899
R12215 gnd.t337 gnd.n4808 5.09899
R12216 gnd.n4886 gnd.n1879 5.09899
R12217 gnd.n5062 gnd.n1784 5.09899
R12218 gnd.n5070 gnd.n1777 5.09899
R12219 gnd.n5235 gnd.n1687 5.09899
R12220 gnd.n1678 gnd.t269 5.09899
R12221 gnd.n6123 gnd.n6122 5.09899
R12222 gnd.n5361 gnd.n1340 5.09899
R12223 gnd.n6116 gnd.n1349 5.09899
R12224 gnd.n5909 gnd.n1352 5.09899
R12225 gnd.n6110 gnd.n1361 5.09899
R12226 gnd.n5917 gnd.n1364 5.09899
R12227 gnd.n6104 gnd.n1372 5.09899
R12228 gnd.n5937 gnd.n5936 5.09899
R12229 gnd.n6098 gnd.n1381 5.09899
R12230 gnd.n5928 gnd.n1384 5.09899
R12231 gnd.n6092 gnd.n1392 5.09899
R12232 gnd.n5990 gnd.n1395 5.09899
R12233 gnd.n5998 gnd.n1404 5.09899
R12234 gnd.n6080 gnd.n1412 5.09899
R12235 gnd.n6004 gnd.n1475 5.09899
R12236 gnd.n6074 gnd.n1421 5.09899
R12237 gnd.n6012 gnd.n1424 5.09899
R12238 gnd.n6068 gnd.n1432 5.09899
R12239 gnd.n6037 gnd.n1435 5.09899
R12240 gnd.n6021 gnd.n1444 5.09899
R12241 gnd.n6056 gnd.n1450 5.09899
R12242 gnd.n6049 gnd.n1458 5.09899
R12243 gnd.n6048 gnd.n1460 5.09899
R12244 gnd.n7304 gnd.n375 5.09899
R12245 gnd.n7300 gnd.n7298 5.09899
R12246 gnd.n7313 gnd.n369 5.09899
R12247 gnd.n7638 gnd.n85 5.09899
R12248 gnd.n7317 gnd.n87 5.09899
R12249 gnd.n7324 gnd.n362 5.09899
R12250 gnd.n7630 gnd.n102 5.09899
R12251 gnd.n7333 gnd.n105 5.09899
R12252 gnd.n7624 gnd.n114 5.09899
R12253 gnd.n7343 gnd.n358 5.09899
R12254 gnd.n7618 gnd.n123 5.09899
R12255 gnd.n7278 gnd.n132 5.09899
R12256 gnd.n3619 gnd.n3618 5.04292
R12257 gnd.n3587 gnd.n3586 5.04292
R12258 gnd.n3555 gnd.n3554 5.04292
R12259 gnd.n3524 gnd.n3523 5.04292
R12260 gnd.n3492 gnd.n3491 5.04292
R12261 gnd.n3460 gnd.n3459 5.04292
R12262 gnd.n3428 gnd.n3427 5.04292
R12263 gnd.n3397 gnd.n3396 5.04292
R12264 gnd.n3129 gnd.t109 4.78034
R12265 gnd.n2452 gnd.t107 4.78034
R12266 gnd.n6460 gnd.t50 4.78034
R12267 gnd.n6441 gnd.t260 4.78034
R12268 gnd.t280 gnd.n4720 4.78034
R12269 gnd.n5721 gnd.t177 4.78034
R12270 gnd.n5555 gnd.t282 4.78034
R12271 gnd.n6062 gnd.t54 4.78034
R12272 gnd.n7624 gnd.t23 4.78034
R12273 gnd.n2571 gnd.n2568 4.74817
R12274 gnd.n2621 gnd.n2503 4.74817
R12275 gnd.n2608 gnd.n2502 4.74817
R12276 gnd.n2501 gnd.n2500 4.74817
R12277 gnd.n2617 gnd.n2568 4.74817
R12278 gnd.n2618 gnd.n2503 4.74817
R12279 gnd.n2620 gnd.n2502 4.74817
R12280 gnd.n2607 gnd.n2501 4.74817
R12281 gnd.n6058 gnd.n98 4.74817
R12282 gnd.n380 gnd.n96 4.74817
R12283 gnd.n7636 gnd.n91 4.74817
R12284 gnd.n7634 gnd.n92 4.74817
R12285 gnd.n1448 gnd.n98 4.74817
R12286 gnd.n7302 gnd.n96 4.74817
R12287 gnd.n379 gnd.n91 4.74817
R12288 gnd.n7635 gnd.n7634 4.74817
R12289 gnd.n4202 gnd.n4201 4.74817
R12290 gnd.n4207 gnd.n2170 4.74817
R12291 gnd.n4213 gnd.n4209 4.74817
R12292 gnd.n4211 gnd.n4210 4.74817
R12293 gnd.n2129 gnd.n2127 4.74817
R12294 gnd.n6044 gnd.n6043 4.74817
R12295 gnd.n6045 gnd.n383 4.74817
R12296 gnd.n7295 gnd.n7294 4.74817
R12297 gnd.n7290 gnd.n384 4.74817
R12298 gnd.n7288 gnd.n7287 4.74817
R12299 gnd.n6043 gnd.n6042 4.74817
R12300 gnd.n6046 gnd.n6045 4.74817
R12301 gnd.n7296 gnd.n7295 4.74817
R12302 gnd.n7293 gnd.n384 4.74817
R12303 gnd.n7289 gnd.n7288 4.74817
R12304 gnd.n6452 gnd.n6451 4.74817
R12305 gnd.n4225 gnd.n976 4.74817
R12306 gnd.n4238 gnd.n975 4.74817
R12307 gnd.n978 gnd.n974 4.74817
R12308 gnd.n6451 gnd.n970 4.74817
R12309 gnd.n2158 gnd.n976 4.74817
R12310 gnd.n4224 gnd.n975 4.74817
R12311 gnd.n4239 gnd.n974 4.74817
R12312 gnd.n4203 gnd.n4202 4.74817
R12313 gnd.n4204 gnd.n2170 4.74817
R12314 gnd.n4209 gnd.n4208 4.74817
R12315 gnd.n4212 gnd.n4211 4.74817
R12316 gnd.n2130 gnd.n2129 4.74817
R12317 gnd.n2566 gnd.n2565 4.74296
R12318 gnd.n78 gnd.n77 4.74296
R12319 gnd.n2534 gnd.n2533 4.7074
R12320 gnd.n2550 gnd.n2549 4.7074
R12321 gnd.n46 gnd.n45 4.7074
R12322 gnd.n62 gnd.n61 4.7074
R12323 gnd.n2566 gnd.n2550 4.65959
R12324 gnd.n78 gnd.n62 4.65959
R12325 gnd.n5815 gnd.n5725 4.6132
R12326 gnd.n6330 gnd.n1147 4.6132
R12327 gnd.n4784 gnd.n1922 4.46168
R12328 gnd.n4775 gnd.n1911 4.46168
R12329 gnd.n4933 gnd.t321 4.46168
R12330 gnd.n4943 gnd.n4942 4.46168
R12331 gnd.n4972 gnd.n1824 4.46168
R12332 gnd.n5120 gnd.n1743 4.46168
R12333 gnd.n5164 gnd.n1730 4.46168
R12334 gnd.t334 gnd.n5163 4.46168
R12335 gnd.n5284 gnd.n1653 4.46168
R12336 gnd.n5304 gnd.n5303 4.46168
R12337 gnd.t244 gnd.n1578 4.46168
R12338 gnd.n5581 gnd.n5568 4.46111
R12339 gnd.n3604 gnd.n3600 4.38594
R12340 gnd.n3572 gnd.n3568 4.38594
R12341 gnd.n3540 gnd.n3536 4.38594
R12342 gnd.n3509 gnd.n3505 4.38594
R12343 gnd.n3477 gnd.n3473 4.38594
R12344 gnd.n3445 gnd.n3441 4.38594
R12345 gnd.n3413 gnd.n3409 4.38594
R12346 gnd.n3382 gnd.n3378 4.38594
R12347 gnd.n3615 gnd.n3593 4.26717
R12348 gnd.n3583 gnd.n3561 4.26717
R12349 gnd.n3551 gnd.n3529 4.26717
R12350 gnd.n3520 gnd.n3498 4.26717
R12351 gnd.n3488 gnd.n3466 4.26717
R12352 gnd.n3456 gnd.n3434 4.26717
R12353 gnd.n3424 gnd.n3402 4.26717
R12354 gnd.n3393 gnd.n3371 4.26717
R12355 gnd.n3073 gnd.t105 4.14303
R12356 gnd.n3303 gnd.t126 4.14303
R12357 gnd.n4121 gnd.t262 4.14303
R12358 gnd.n6417 gnd.t15 4.14303
R12359 gnd.t163 gnd.n1086 4.14303
R12360 gnd.t141 gnd.n1349 4.14303
R12361 gnd.n6086 gnd.t65 4.14303
R12362 gnd.n7600 gnd.t39 4.14303
R12363 gnd.n3623 gnd.n3622 4.08274
R12364 gnd.n5714 gnd.n5713 4.05904
R12365 gnd.n1957 gnd.n1956 4.05904
R12366 gnd.n6270 gnd.n6263 4.05904
R12367 gnd.n5594 gnd.n5593 4.05904
R12368 gnd.n15 gnd.n7 3.99943
R12369 gnd.n6256 gnd.n6255 3.82437
R12370 gnd.n4843 gnd.n1892 3.82437
R12371 gnd.n4884 gnd.t339 3.82437
R12372 gnd.n4904 gnd.n4903 3.82437
R12373 gnd.n4992 gnd.n1813 3.82437
R12374 gnd.n4993 gnd.t53 3.82437
R12375 gnd.n5034 gnd.t313 3.82437
R12376 gnd.n5079 gnd.n5078 3.82437
R12377 gnd.n5194 gnd.n1701 3.82437
R12378 gnd.n5227 gnd.t69 3.82437
R12379 gnd.n5244 gnd.n5243 3.82437
R12380 gnd.n5562 gnd.n1581 3.82437
R12381 gnd.n3146 gnd.n2567 3.81325
R12382 gnd.n2550 gnd.n2534 3.72967
R12383 gnd.n62 gnd.n46 3.72967
R12384 gnd.n3623 gnd.n3495 3.70378
R12385 gnd.n15 gnd.n14 3.60163
R12386 gnd.t125 gnd.n934 3.50571
R12387 gnd.n3614 gnd.n3595 3.49141
R12388 gnd.n3582 gnd.n3563 3.49141
R12389 gnd.n3550 gnd.n3531 3.49141
R12390 gnd.n3519 gnd.n3500 3.49141
R12391 gnd.n3487 gnd.n3468 3.49141
R12392 gnd.n3455 gnd.n3436 3.49141
R12393 gnd.n3423 gnd.n3404 3.49141
R12394 gnd.n3392 gnd.n3373 3.49141
R12395 gnd.n5796 gnd.n5795 3.29747
R12396 gnd.n5795 gnd.n5733 3.29747
R12397 gnd.n7529 gnd.n7526 3.29747
R12398 gnd.n7530 gnd.n7529 3.29747
R12399 gnd.n4008 gnd.n4007 3.29747
R12400 gnd.n4007 gnd.n4006 3.29747
R12401 gnd.n6346 gnd.n6345 3.29747
R12402 gnd.n6345 gnd.n6344 3.29747
R12403 gnd.n3342 gnd.n934 3.18706
R12404 gnd.n6248 gnd.n1223 3.18706
R12405 gnd.n1930 gnd.t207 3.18706
R12406 gnd.n4815 gnd.n1899 3.18706
R12407 gnd.n4824 gnd.t336 3.18706
R12408 gnd.t336 gnd.n1884 3.18706
R12409 gnd.n4922 gnd.n4920 3.18706
R12410 gnd.n4983 gnd.n4982 3.18706
R12411 gnd.n5094 gnd.n5093 3.18706
R12412 gnd.n5175 gnd.n5174 3.18706
R12413 gnd.t306 gnd.n1690 3.18706
R12414 gnd.n5125 gnd.t306 3.18706
R12415 gnd.n5260 gnd.n5259 3.18706
R12416 gnd.n5327 gnd.n1622 3.18706
R12417 gnd.n5335 gnd.t244 3.18706
R12418 gnd.n2652 gnd.t105 2.8684
R12419 gnd.n4791 gnd.t8 2.8684
R12420 gnd.t344 gnd.n5293 2.8684
R12421 gnd.n2551 gnd.t352 2.82907
R12422 gnd.n2551 gnd.t259 2.82907
R12423 gnd.n2553 gnd.t45 2.82907
R12424 gnd.n2553 gnd.t268 2.82907
R12425 gnd.n2555 gnd.t27 2.82907
R12426 gnd.n2555 gnd.t274 2.82907
R12427 gnd.n2557 gnd.t47 2.82907
R12428 gnd.n2557 gnd.t73 2.82907
R12429 gnd.n2559 gnd.t51 2.82907
R12430 gnd.n2559 gnd.t87 2.82907
R12431 gnd.n2561 gnd.t265 2.82907
R12432 gnd.n2561 gnd.t358 2.82907
R12433 gnd.n2563 gnd.t91 2.82907
R12434 gnd.n2563 gnd.t356 2.82907
R12435 gnd.n2504 gnd.t16 2.82907
R12436 gnd.n2504 gnd.t302 2.82907
R12437 gnd.n2506 gnd.t25 2.82907
R12438 gnd.n2506 gnd.t331 2.82907
R12439 gnd.n2508 gnd.t88 2.82907
R12440 gnd.n2508 gnd.t343 2.82907
R12441 gnd.n2510 gnd.t267 2.82907
R12442 gnd.n2510 gnd.t324 2.82907
R12443 gnd.n2512 gnd.t328 2.82907
R12444 gnd.n2512 gnd.t76 2.82907
R12445 gnd.n2514 gnd.t326 2.82907
R12446 gnd.n2514 gnd.t123 2.82907
R12447 gnd.n2516 gnd.t100 2.82907
R12448 gnd.n2516 gnd.t357 2.82907
R12449 gnd.n2519 gnd.t63 2.82907
R12450 gnd.n2519 gnd.t346 2.82907
R12451 gnd.n2521 gnd.t18 2.82907
R12452 gnd.n2521 gnd.t347 2.82907
R12453 gnd.n2523 gnd.t314 2.82907
R12454 gnd.n2523 gnd.t261 2.82907
R12455 gnd.n2525 gnd.t96 2.82907
R12456 gnd.n2525 gnd.t351 2.82907
R12457 gnd.n2527 gnd.t122 2.82907
R12458 gnd.n2527 gnd.t36 2.82907
R12459 gnd.n2529 gnd.t44 2.82907
R12460 gnd.n2529 gnd.t120 2.82907
R12461 gnd.n2531 gnd.t271 2.82907
R12462 gnd.n2531 gnd.t325 2.82907
R12463 gnd.n2535 gnd.t48 2.82907
R12464 gnd.n2535 gnd.t330 2.82907
R12465 gnd.n2537 gnd.t299 2.82907
R12466 gnd.n2537 gnd.t71 2.82907
R12467 gnd.n2539 gnd.t74 2.82907
R12468 gnd.n2539 gnd.t300 2.82907
R12469 gnd.n2541 gnd.t322 2.82907
R12470 gnd.n2541 gnd.t303 2.82907
R12471 gnd.n2543 gnd.t62 2.82907
R12472 gnd.n2543 gnd.t119 2.82907
R12473 gnd.n2545 gnd.t251 2.82907
R12474 gnd.n2545 gnd.t61 2.82907
R12475 gnd.n2547 gnd.t327 2.82907
R12476 gnd.n2547 gnd.t263 2.82907
R12477 gnd.n75 gnd.t332 2.82907
R12478 gnd.n75 gnd.t252 2.82907
R12479 gnd.n73 gnd.t348 2.82907
R12480 gnd.n73 gnd.t279 2.82907
R12481 gnd.n71 gnd.t319 2.82907
R12482 gnd.n71 gnd.t24 2.82907
R12483 gnd.n69 gnd.t257 2.82907
R12484 gnd.n69 gnd.t312 2.82907
R12485 gnd.n67 gnd.t301 2.82907
R12486 gnd.n67 gnd.t315 2.82907
R12487 gnd.n65 gnd.t276 2.82907
R12488 gnd.n65 gnd.t367 2.82907
R12489 gnd.n63 gnd.t359 2.82907
R12490 gnd.n63 gnd.t308 2.82907
R12491 gnd.n28 gnd.t316 2.82907
R12492 gnd.n28 gnd.t5 2.82907
R12493 gnd.n26 gnd.t329 2.82907
R12494 gnd.n26 gnd.t42 2.82907
R12495 gnd.n24 gnd.t1 2.82907
R12496 gnd.n24 gnd.t333 2.82907
R12497 gnd.n22 gnd.t3 2.82907
R12498 gnd.n22 gnd.t101 2.82907
R12499 gnd.n20 gnd.t102 2.82907
R12500 gnd.n20 gnd.t266 2.82907
R12501 gnd.n18 gnd.t118 2.82907
R12502 gnd.n18 gnd.t59 2.82907
R12503 gnd.n16 gnd.t20 2.82907
R12504 gnd.n16 gnd.t66 2.82907
R12505 gnd.n43 gnd.t86 2.82907
R12506 gnd.n43 gnd.t14 2.82907
R12507 gnd.n41 gnd.t255 2.82907
R12508 gnd.n41 gnd.t49 2.82907
R12509 gnd.n39 gnd.t89 2.82907
R12510 gnd.n39 gnd.t342 2.82907
R12511 gnd.n37 gnd.t323 2.82907
R12512 gnd.n37 gnd.t296 2.82907
R12513 gnd.n35 gnd.t264 2.82907
R12514 gnd.n35 gnd.t353 2.82907
R12515 gnd.n33 gnd.t38 2.82907
R12516 gnd.n33 gnd.t341 2.82907
R12517 gnd.n31 gnd.t97 2.82907
R12518 gnd.n31 gnd.t98 2.82907
R12519 gnd.n59 gnd.t40 2.82907
R12520 gnd.n59 gnd.t311 2.82907
R12521 gnd.n57 gnd.t22 2.82907
R12522 gnd.n57 gnd.t83 2.82907
R12523 gnd.n55 gnd.t310 2.82907
R12524 gnd.n55 gnd.t75 2.82907
R12525 gnd.n53 gnd.t64 2.82907
R12526 gnd.n53 gnd.t7 2.82907
R12527 gnd.n51 gnd.t55 2.82907
R12528 gnd.n51 gnd.t117 2.82907
R12529 gnd.n49 gnd.t249 2.82907
R12530 gnd.n49 gnd.t349 2.82907
R12531 gnd.n47 gnd.t250 2.82907
R12532 gnd.n47 gnd.t294 2.82907
R12533 gnd.n3611 gnd.n3610 2.71565
R12534 gnd.n3579 gnd.n3578 2.71565
R12535 gnd.n3547 gnd.n3546 2.71565
R12536 gnd.n3516 gnd.n3515 2.71565
R12537 gnd.n3484 gnd.n3483 2.71565
R12538 gnd.n3452 gnd.n3451 2.71565
R12539 gnd.n3420 gnd.n3419 2.71565
R12540 gnd.n3389 gnd.n3388 2.71565
R12541 gnd.n6249 gnd.n1221 2.54975
R12542 gnd.n4833 gnd.n4832 2.54975
R12543 gnd.n4809 gnd.t337 2.54975
R12544 gnd.n4923 gnd.n1855 2.54975
R12545 gnd.n4923 gnd.t307 2.54975
R12546 gnd.n5003 gnd.n1806 2.54975
R12547 gnd.n5095 gnd.n1757 2.54975
R12548 gnd.n5184 gnd.t304 2.54975
R12549 gnd.n5184 gnd.n5183 2.54975
R12550 gnd.n5251 gnd.t269 2.54975
R12551 gnd.n5261 gnd.n1667 2.54975
R12552 gnd.n1631 gnd.n1618 2.54975
R12553 gnd.n3146 gnd.n2568 2.27742
R12554 gnd.n3146 gnd.n2503 2.27742
R12555 gnd.n3146 gnd.n2502 2.27742
R12556 gnd.n3146 gnd.n2501 2.27742
R12557 gnd.n7633 gnd.n98 2.27742
R12558 gnd.n7633 gnd.n96 2.27742
R12559 gnd.n7633 gnd.n91 2.27742
R12560 gnd.n7634 gnd.n7633 2.27742
R12561 gnd.n6043 gnd.n95 2.27742
R12562 gnd.n6045 gnd.n95 2.27742
R12563 gnd.n7295 gnd.n95 2.27742
R12564 gnd.n384 gnd.n95 2.27742
R12565 gnd.n7288 gnd.n95 2.27742
R12566 gnd.n6451 gnd.n6450 2.27742
R12567 gnd.n6450 gnd.n976 2.27742
R12568 gnd.n6450 gnd.n975 2.27742
R12569 gnd.n6450 gnd.n974 2.27742
R12570 gnd.n4202 gnd.n973 2.27742
R12571 gnd.n2170 gnd.n973 2.27742
R12572 gnd.n4209 gnd.n973 2.27742
R12573 gnd.n4211 gnd.n973 2.27742
R12574 gnd.n2129 gnd.n973 2.27742
R12575 gnd.n3000 gnd.t203 2.23109
R12576 gnd.n2623 gnd.t109 2.23109
R12577 gnd.t94 gnd.n1824 2.23109
R12578 gnd.t364 gnd.n4992 2.23109
R12579 gnd.n5079 gnd.t290 2.23109
R12580 gnd.t253 gnd.n1743 2.23109
R12581 gnd.n3607 gnd.n3597 1.93989
R12582 gnd.n3575 gnd.n3565 1.93989
R12583 gnd.n3543 gnd.n3533 1.93989
R12584 gnd.n3512 gnd.n3502 1.93989
R12585 gnd.n3480 gnd.n3470 1.93989
R12586 gnd.n3448 gnd.n3438 1.93989
R12587 gnd.n3416 gnd.n3406 1.93989
R12588 gnd.n3385 gnd.n3375 1.93989
R12589 gnd.n2020 gnd.n1212 1.91244
R12590 gnd.n2020 gnd.t160 1.91244
R12591 gnd.n4817 gnd.t34 1.91244
R12592 gnd.n4845 gnd.n1891 1.91244
R12593 gnd.n4853 gnd.n4852 1.91244
R12594 gnd.n5012 gnd.n1801 1.91244
R12595 gnd.n1771 gnd.n1770 1.91244
R12596 gnd.n5196 gnd.n5195 1.91244
R12597 gnd.n1681 gnd.n1679 1.91244
R12598 gnd.n5274 gnd.t340 1.91244
R12599 gnd.n5564 gnd.n5563 1.91244
R12600 gnd.t30 gnd.n3011 1.59378
R12601 gnd.n3190 gnd.t111 1.59378
R12602 gnd.n2436 gnd.t67 1.59378
R12603 gnd.n4809 gnd.t354 1.59378
R12604 gnd.t362 gnd.n1846 1.59378
R12605 gnd.n5176 gnd.t284 1.59378
R12606 gnd.n5251 gnd.t360 1.59378
R12607 gnd.t228 gnd.n2027 1.27512
R12608 gnd.n4757 gnd.n4756 1.27512
R12609 gnd.n4777 gnd.t320 1.27512
R12610 gnd.n4800 gnd.n4799 1.27512
R12611 gnd.n4895 gnd.t339 1.27512
R12612 gnd.n4934 gnd.n4933 1.27512
R12613 gnd.n4956 gnd.n1833 1.27512
R12614 gnd.n5104 gnd.n5103 1.27512
R12615 gnd.n5163 gnd.n1731 1.27512
R12616 gnd.n5132 gnd.t69 1.27512
R12617 gnd.n5272 gnd.n5271 1.27512
R12618 gnd.t305 gnd.n1645 1.27512
R12619 gnd.n5303 gnd.t149 1.27512
R12620 gnd.n5320 gnd.n1627 1.27512
R12621 gnd.n2853 gnd.n2845 1.16414
R12622 gnd.n3669 gnd.n2339 1.16414
R12623 gnd.n3606 gnd.n3599 1.16414
R12624 gnd.n3574 gnd.n3567 1.16414
R12625 gnd.n3542 gnd.n3535 1.16414
R12626 gnd.n3511 gnd.n3504 1.16414
R12627 gnd.n3479 gnd.n3472 1.16414
R12628 gnd.n3447 gnd.n3440 1.16414
R12629 gnd.n3415 gnd.n3408 1.16414
R12630 gnd.n3384 gnd.n3377 1.16414
R12631 gnd.n5725 gnd.n1531 0.970197
R12632 gnd.n6330 gnd.n1144 0.970197
R12633 gnd.n3590 gnd.n3558 0.962709
R12634 gnd.n3622 gnd.n3590 0.962709
R12635 gnd.n3463 gnd.n3431 0.962709
R12636 gnd.n3495 gnd.n3463 0.962709
R12637 gnd.n3099 gnd.t272 0.956468
R12638 gnd.n3264 gnd.t113 0.956468
R12639 gnd.n6467 gnd.t60 0.956468
R12640 gnd.n2114 gnd.t15 0.956468
R12641 gnd.n6326 gnd.n1184 0.956468
R12642 gnd.t10 gnd.n4743 0.956468
R12643 gnd.n5336 gnd.t286 0.956468
R12644 gnd.n5721 gnd.n1536 0.956468
R12645 gnd.n5989 gnd.t65 0.956468
R12646 gnd.n7278 gnd.t21 0.956468
R12647 gnd.n2 gnd.n1 0.672012
R12648 gnd.n3 gnd.n2 0.672012
R12649 gnd.n4 gnd.n3 0.672012
R12650 gnd.n5 gnd.n4 0.672012
R12651 gnd.n6 gnd.n5 0.672012
R12652 gnd.n7 gnd.n6 0.672012
R12653 gnd.n9 gnd.n8 0.672012
R12654 gnd.n10 gnd.n9 0.672012
R12655 gnd.n11 gnd.n10 0.672012
R12656 gnd.n12 gnd.n11 0.672012
R12657 gnd.n13 gnd.n12 0.672012
R12658 gnd.n14 gnd.n13 0.672012
R12659 gnd.t199 gnd.n6248 0.637812
R12660 gnd.t180 gnd.n4757 0.637812
R12661 gnd.n4873 gnd.n4872 0.637812
R12662 gnd.n4894 gnd.n4892 0.637812
R12663 gnd.n4903 gnd.t81 0.637812
R12664 gnd.n5023 gnd.n5022 0.637812
R12665 gnd.n5069 gnd.n5068 0.637812
R12666 gnd.t270 gnd.n5194 0.637812
R12667 gnd.n5135 gnd.n5134 0.637812
R12668 gnd.n5234 gnd.n5233 0.637812
R12669 gnd.t152 gnd.n1622 0.637812
R12670 gnd.n5344 gnd.t193 0.637812
R12671 gnd gnd.n0 0.59317
R12672 gnd.n2565 gnd.n2564 0.573776
R12673 gnd.n2564 gnd.n2562 0.573776
R12674 gnd.n2562 gnd.n2560 0.573776
R12675 gnd.n2560 gnd.n2558 0.573776
R12676 gnd.n2558 gnd.n2556 0.573776
R12677 gnd.n2556 gnd.n2554 0.573776
R12678 gnd.n2554 gnd.n2552 0.573776
R12679 gnd.n2518 gnd.n2517 0.573776
R12680 gnd.n2517 gnd.n2515 0.573776
R12681 gnd.n2515 gnd.n2513 0.573776
R12682 gnd.n2513 gnd.n2511 0.573776
R12683 gnd.n2511 gnd.n2509 0.573776
R12684 gnd.n2509 gnd.n2507 0.573776
R12685 gnd.n2507 gnd.n2505 0.573776
R12686 gnd.n2533 gnd.n2532 0.573776
R12687 gnd.n2532 gnd.n2530 0.573776
R12688 gnd.n2530 gnd.n2528 0.573776
R12689 gnd.n2528 gnd.n2526 0.573776
R12690 gnd.n2526 gnd.n2524 0.573776
R12691 gnd.n2524 gnd.n2522 0.573776
R12692 gnd.n2522 gnd.n2520 0.573776
R12693 gnd.n2549 gnd.n2548 0.573776
R12694 gnd.n2548 gnd.n2546 0.573776
R12695 gnd.n2546 gnd.n2544 0.573776
R12696 gnd.n2544 gnd.n2542 0.573776
R12697 gnd.n2542 gnd.n2540 0.573776
R12698 gnd.n2540 gnd.n2538 0.573776
R12699 gnd.n2538 gnd.n2536 0.573776
R12700 gnd.n66 gnd.n64 0.573776
R12701 gnd.n68 gnd.n66 0.573776
R12702 gnd.n70 gnd.n68 0.573776
R12703 gnd.n72 gnd.n70 0.573776
R12704 gnd.n74 gnd.n72 0.573776
R12705 gnd.n76 gnd.n74 0.573776
R12706 gnd.n77 gnd.n76 0.573776
R12707 gnd.n19 gnd.n17 0.573776
R12708 gnd.n21 gnd.n19 0.573776
R12709 gnd.n23 gnd.n21 0.573776
R12710 gnd.n25 gnd.n23 0.573776
R12711 gnd.n27 gnd.n25 0.573776
R12712 gnd.n29 gnd.n27 0.573776
R12713 gnd.n30 gnd.n29 0.573776
R12714 gnd.n34 gnd.n32 0.573776
R12715 gnd.n36 gnd.n34 0.573776
R12716 gnd.n38 gnd.n36 0.573776
R12717 gnd.n40 gnd.n38 0.573776
R12718 gnd.n42 gnd.n40 0.573776
R12719 gnd.n44 gnd.n42 0.573776
R12720 gnd.n45 gnd.n44 0.573776
R12721 gnd.n50 gnd.n48 0.573776
R12722 gnd.n52 gnd.n50 0.573776
R12723 gnd.n54 gnd.n52 0.573776
R12724 gnd.n56 gnd.n54 0.573776
R12725 gnd.n58 gnd.n56 0.573776
R12726 gnd.n60 gnd.n58 0.573776
R12727 gnd.n61 gnd.n60 0.573776
R12728 gnd.n7645 gnd.n7644 0.553533
R12729 gnd.n7418 gnd.n7417 0.505073
R12730 gnd.n3887 gnd.n3885 0.505073
R12731 gnd.n5537 gnd.n5536 0.489829
R12732 gnd.n4673 gnd.n4671 0.489829
R12733 gnd.n4416 gnd.n2056 0.489829
R12734 gnd.n6141 gnd.n1314 0.489829
R12735 gnd.n3326 gnd.n2343 0.486781
R12736 gnd.n2902 gnd.n2901 0.48678
R12737 gnd.n3643 gnd.n2297 0.480683
R12738 gnd.n2986 gnd.n2985 0.480683
R12739 gnd.n6642 gnd.n6641 0.480683
R12740 gnd.n7063 gnd.n7062 0.480683
R12741 gnd.n7275 gnd.n7274 0.480683
R12742 gnd.n6471 gnd.n6470 0.480683
R12743 gnd.n7561 gnd.n7560 0.470012
R12744 gnd.n5751 gnd.n1344 0.470012
R12745 gnd.n6378 gnd.n6377 0.470012
R12746 gnd.n3789 gnd.n2256 0.470012
R12747 gnd.n7633 gnd.n95 0.4255
R12748 gnd.n6450 gnd.n973 0.4255
R12749 gnd.n4598 gnd.n2084 0.388379
R12750 gnd.n3603 gnd.n3602 0.388379
R12751 gnd.n3571 gnd.n3570 0.388379
R12752 gnd.n3539 gnd.n3538 0.388379
R12753 gnd.n3508 gnd.n3507 0.388379
R12754 gnd.n3476 gnd.n3475 0.388379
R12755 gnd.n3444 gnd.n3443 0.388379
R12756 gnd.n3412 gnd.n3411 0.388379
R12757 gnd.n3381 gnd.n3380 0.388379
R12758 gnd.n5514 gnd.n5372 0.388379
R12759 gnd.n7645 gnd.n15 0.374463
R12760 gnd.n2398 gnd.t125 0.319156
R12761 gnd.n2161 gnd.t46 0.319156
R12762 gnd.n4253 gnd.t260 0.319156
R12763 gnd.n4687 gnd.t189 0.319156
R12764 gnd.t173 gnd.n5542 0.319156
R12765 gnd.n6038 gnd.t54 0.319156
R12766 gnd.t6 gnd.n85 0.319156
R12767 gnd.n2820 gnd.n2798 0.311721
R12768 gnd gnd.n7645 0.295112
R12769 gnd.n7451 gnd.n7450 0.293183
R12770 gnd.n3925 gnd.n3924 0.293183
R12771 gnd.n2109 gnd.n2071 0.27489
R12772 gnd.n5366 gnd.n5365 0.27489
R12773 gnd.n3714 gnd.n3713 0.268793
R12774 gnd.n7452 gnd.n7451 0.258122
R12775 gnd.n5901 gnd.n5900 0.258122
R12776 gnd.n4535 gnd.n4534 0.258122
R12777 gnd.n3926 gnd.n3925 0.258122
R12778 gnd.n3713 gnd.n3712 0.241354
R12779 gnd.n5816 gnd.n5815 0.229039
R12780 gnd.n5815 gnd.n1530 0.229039
R12781 gnd.n1147 gnd.n1143 0.229039
R12782 gnd.n4455 gnd.n1147 0.229039
R12783 gnd.n2974 gnd.n2773 0.206293
R12784 gnd.n2567 gnd.n0 0.169152
R12785 gnd.n3620 gnd.n3592 0.155672
R12786 gnd.n3613 gnd.n3592 0.155672
R12787 gnd.n3613 gnd.n3612 0.155672
R12788 gnd.n3612 gnd.n3596 0.155672
R12789 gnd.n3605 gnd.n3596 0.155672
R12790 gnd.n3605 gnd.n3604 0.155672
R12791 gnd.n3588 gnd.n3560 0.155672
R12792 gnd.n3581 gnd.n3560 0.155672
R12793 gnd.n3581 gnd.n3580 0.155672
R12794 gnd.n3580 gnd.n3564 0.155672
R12795 gnd.n3573 gnd.n3564 0.155672
R12796 gnd.n3573 gnd.n3572 0.155672
R12797 gnd.n3556 gnd.n3528 0.155672
R12798 gnd.n3549 gnd.n3528 0.155672
R12799 gnd.n3549 gnd.n3548 0.155672
R12800 gnd.n3548 gnd.n3532 0.155672
R12801 gnd.n3541 gnd.n3532 0.155672
R12802 gnd.n3541 gnd.n3540 0.155672
R12803 gnd.n3525 gnd.n3497 0.155672
R12804 gnd.n3518 gnd.n3497 0.155672
R12805 gnd.n3518 gnd.n3517 0.155672
R12806 gnd.n3517 gnd.n3501 0.155672
R12807 gnd.n3510 gnd.n3501 0.155672
R12808 gnd.n3510 gnd.n3509 0.155672
R12809 gnd.n3493 gnd.n3465 0.155672
R12810 gnd.n3486 gnd.n3465 0.155672
R12811 gnd.n3486 gnd.n3485 0.155672
R12812 gnd.n3485 gnd.n3469 0.155672
R12813 gnd.n3478 gnd.n3469 0.155672
R12814 gnd.n3478 gnd.n3477 0.155672
R12815 gnd.n3461 gnd.n3433 0.155672
R12816 gnd.n3454 gnd.n3433 0.155672
R12817 gnd.n3454 gnd.n3453 0.155672
R12818 gnd.n3453 gnd.n3437 0.155672
R12819 gnd.n3446 gnd.n3437 0.155672
R12820 gnd.n3446 gnd.n3445 0.155672
R12821 gnd.n3429 gnd.n3401 0.155672
R12822 gnd.n3422 gnd.n3401 0.155672
R12823 gnd.n3422 gnd.n3421 0.155672
R12824 gnd.n3421 gnd.n3405 0.155672
R12825 gnd.n3414 gnd.n3405 0.155672
R12826 gnd.n3414 gnd.n3413 0.155672
R12827 gnd.n3398 gnd.n3370 0.155672
R12828 gnd.n3391 gnd.n3370 0.155672
R12829 gnd.n3391 gnd.n3390 0.155672
R12830 gnd.n3390 gnd.n3374 0.155672
R12831 gnd.n3383 gnd.n3374 0.155672
R12832 gnd.n3383 gnd.n3382 0.155672
R12833 gnd.n3745 gnd.n2297 0.152939
R12834 gnd.n3745 gnd.n3744 0.152939
R12835 gnd.n3744 gnd.n3743 0.152939
R12836 gnd.n3743 gnd.n2299 0.152939
R12837 gnd.n2300 gnd.n2299 0.152939
R12838 gnd.n2301 gnd.n2300 0.152939
R12839 gnd.n2302 gnd.n2301 0.152939
R12840 gnd.n2303 gnd.n2302 0.152939
R12841 gnd.n2304 gnd.n2303 0.152939
R12842 gnd.n2305 gnd.n2304 0.152939
R12843 gnd.n2306 gnd.n2305 0.152939
R12844 gnd.n2307 gnd.n2306 0.152939
R12845 gnd.n2308 gnd.n2307 0.152939
R12846 gnd.n2309 gnd.n2308 0.152939
R12847 gnd.n3715 gnd.n2309 0.152939
R12848 gnd.n3715 gnd.n3714 0.152939
R12849 gnd.n2987 gnd.n2986 0.152939
R12850 gnd.n2987 gnd.n2691 0.152939
R12851 gnd.n3015 gnd.n2691 0.152939
R12852 gnd.n3016 gnd.n3015 0.152939
R12853 gnd.n3017 gnd.n3016 0.152939
R12854 gnd.n3018 gnd.n3017 0.152939
R12855 gnd.n3018 gnd.n2663 0.152939
R12856 gnd.n3045 gnd.n2663 0.152939
R12857 gnd.n3046 gnd.n3045 0.152939
R12858 gnd.n3047 gnd.n3046 0.152939
R12859 gnd.n3047 gnd.n2641 0.152939
R12860 gnd.n3076 gnd.n2641 0.152939
R12861 gnd.n3077 gnd.n3076 0.152939
R12862 gnd.n3078 gnd.n3077 0.152939
R12863 gnd.n3079 gnd.n3078 0.152939
R12864 gnd.n3081 gnd.n3079 0.152939
R12865 gnd.n3081 gnd.n3080 0.152939
R12866 gnd.n3080 gnd.n2590 0.152939
R12867 gnd.n2591 gnd.n2590 0.152939
R12868 gnd.n2592 gnd.n2591 0.152939
R12869 gnd.n2611 gnd.n2592 0.152939
R12870 gnd.n2612 gnd.n2611 0.152939
R12871 gnd.n2612 gnd.n2494 0.152939
R12872 gnd.n3171 gnd.n2494 0.152939
R12873 gnd.n3172 gnd.n3171 0.152939
R12874 gnd.n3173 gnd.n3172 0.152939
R12875 gnd.n3174 gnd.n3173 0.152939
R12876 gnd.n3174 gnd.n2467 0.152939
R12877 gnd.n3211 gnd.n2467 0.152939
R12878 gnd.n3212 gnd.n3211 0.152939
R12879 gnd.n3213 gnd.n3212 0.152939
R12880 gnd.n3214 gnd.n3213 0.152939
R12881 gnd.n3214 gnd.n2440 0.152939
R12882 gnd.n3256 gnd.n2440 0.152939
R12883 gnd.n3257 gnd.n3256 0.152939
R12884 gnd.n3258 gnd.n3257 0.152939
R12885 gnd.n3259 gnd.n3258 0.152939
R12886 gnd.n3259 gnd.n2412 0.152939
R12887 gnd.n3296 gnd.n2412 0.152939
R12888 gnd.n3297 gnd.n3296 0.152939
R12889 gnd.n3298 gnd.n3297 0.152939
R12890 gnd.n3299 gnd.n3298 0.152939
R12891 gnd.n3299 gnd.n2385 0.152939
R12892 gnd.n3345 gnd.n2385 0.152939
R12893 gnd.n3346 gnd.n3345 0.152939
R12894 gnd.n3347 gnd.n3346 0.152939
R12895 gnd.n3348 gnd.n3347 0.152939
R12896 gnd.n3348 gnd.n2358 0.152939
R12897 gnd.n3639 gnd.n2358 0.152939
R12898 gnd.n3640 gnd.n3639 0.152939
R12899 gnd.n3641 gnd.n3640 0.152939
R12900 gnd.n3642 gnd.n3641 0.152939
R12901 gnd.n3643 gnd.n3642 0.152939
R12902 gnd.n2985 gnd.n2715 0.152939
R12903 gnd.n2736 gnd.n2715 0.152939
R12904 gnd.n2737 gnd.n2736 0.152939
R12905 gnd.n2743 gnd.n2737 0.152939
R12906 gnd.n2744 gnd.n2743 0.152939
R12907 gnd.n2745 gnd.n2744 0.152939
R12908 gnd.n2745 gnd.n2734 0.152939
R12909 gnd.n2753 gnd.n2734 0.152939
R12910 gnd.n2754 gnd.n2753 0.152939
R12911 gnd.n2755 gnd.n2754 0.152939
R12912 gnd.n2755 gnd.n2732 0.152939
R12913 gnd.n2763 gnd.n2732 0.152939
R12914 gnd.n2764 gnd.n2763 0.152939
R12915 gnd.n2765 gnd.n2764 0.152939
R12916 gnd.n2765 gnd.n2730 0.152939
R12917 gnd.n2773 gnd.n2730 0.152939
R12918 gnd.n3712 gnd.n2314 0.152939
R12919 gnd.n2316 gnd.n2314 0.152939
R12920 gnd.n2317 gnd.n2316 0.152939
R12921 gnd.n2318 gnd.n2317 0.152939
R12922 gnd.n2319 gnd.n2318 0.152939
R12923 gnd.n2320 gnd.n2319 0.152939
R12924 gnd.n2321 gnd.n2320 0.152939
R12925 gnd.n2322 gnd.n2321 0.152939
R12926 gnd.n2323 gnd.n2322 0.152939
R12927 gnd.n2324 gnd.n2323 0.152939
R12928 gnd.n2325 gnd.n2324 0.152939
R12929 gnd.n2326 gnd.n2325 0.152939
R12930 gnd.n2327 gnd.n2326 0.152939
R12931 gnd.n2328 gnd.n2327 0.152939
R12932 gnd.n2329 gnd.n2328 0.152939
R12933 gnd.n2330 gnd.n2329 0.152939
R12934 gnd.n2331 gnd.n2330 0.152939
R12935 gnd.n2332 gnd.n2331 0.152939
R12936 gnd.n2333 gnd.n2332 0.152939
R12937 gnd.n2334 gnd.n2333 0.152939
R12938 gnd.n2335 gnd.n2334 0.152939
R12939 gnd.n2336 gnd.n2335 0.152939
R12940 gnd.n2340 gnd.n2336 0.152939
R12941 gnd.n2341 gnd.n2340 0.152939
R12942 gnd.n2342 gnd.n2341 0.152939
R12943 gnd.n2343 gnd.n2342 0.152939
R12944 gnd.n3148 gnd.n3147 0.152939
R12945 gnd.n3149 gnd.n3148 0.152939
R12946 gnd.n3150 gnd.n3149 0.152939
R12947 gnd.n3151 gnd.n3150 0.152939
R12948 gnd.n3152 gnd.n3151 0.152939
R12949 gnd.n3153 gnd.n3152 0.152939
R12950 gnd.n3153 gnd.n2448 0.152939
R12951 gnd.n3232 gnd.n2448 0.152939
R12952 gnd.n3233 gnd.n3232 0.152939
R12953 gnd.n3234 gnd.n3233 0.152939
R12954 gnd.n3235 gnd.n3234 0.152939
R12955 gnd.n3236 gnd.n3235 0.152939
R12956 gnd.n3237 gnd.n3236 0.152939
R12957 gnd.n3238 gnd.n3237 0.152939
R12958 gnd.n3239 gnd.n3238 0.152939
R12959 gnd.n3240 gnd.n3239 0.152939
R12960 gnd.n3240 gnd.n2392 0.152939
R12961 gnd.n3317 gnd.n2392 0.152939
R12962 gnd.n3318 gnd.n3317 0.152939
R12963 gnd.n3319 gnd.n3318 0.152939
R12964 gnd.n3320 gnd.n3319 0.152939
R12965 gnd.n3321 gnd.n3320 0.152939
R12966 gnd.n3322 gnd.n3321 0.152939
R12967 gnd.n3323 gnd.n3322 0.152939
R12968 gnd.n3324 gnd.n3323 0.152939
R12969 gnd.n3325 gnd.n3324 0.152939
R12970 gnd.n3327 gnd.n3325 0.152939
R12971 gnd.n3327 gnd.n3326 0.152939
R12972 gnd.n2903 gnd.n2902 0.152939
R12973 gnd.n2903 gnd.n2793 0.152939
R12974 gnd.n2918 gnd.n2793 0.152939
R12975 gnd.n2919 gnd.n2918 0.152939
R12976 gnd.n2920 gnd.n2919 0.152939
R12977 gnd.n2920 gnd.n2781 0.152939
R12978 gnd.n2934 gnd.n2781 0.152939
R12979 gnd.n2935 gnd.n2934 0.152939
R12980 gnd.n2936 gnd.n2935 0.152939
R12981 gnd.n2937 gnd.n2936 0.152939
R12982 gnd.n2938 gnd.n2937 0.152939
R12983 gnd.n2939 gnd.n2938 0.152939
R12984 gnd.n2940 gnd.n2939 0.152939
R12985 gnd.n2941 gnd.n2940 0.152939
R12986 gnd.n2942 gnd.n2941 0.152939
R12987 gnd.n2943 gnd.n2942 0.152939
R12988 gnd.n2944 gnd.n2943 0.152939
R12989 gnd.n2945 gnd.n2944 0.152939
R12990 gnd.n2946 gnd.n2945 0.152939
R12991 gnd.n2947 gnd.n2946 0.152939
R12992 gnd.n2948 gnd.n2947 0.152939
R12993 gnd.n2948 gnd.n2647 0.152939
R12994 gnd.n3065 gnd.n2647 0.152939
R12995 gnd.n3066 gnd.n3065 0.152939
R12996 gnd.n3067 gnd.n3066 0.152939
R12997 gnd.n3068 gnd.n3067 0.152939
R12998 gnd.n3068 gnd.n2569 0.152939
R12999 gnd.n3145 gnd.n2569 0.152939
R13000 gnd.n2821 gnd.n2820 0.152939
R13001 gnd.n2822 gnd.n2821 0.152939
R13002 gnd.n2823 gnd.n2822 0.152939
R13003 gnd.n2824 gnd.n2823 0.152939
R13004 gnd.n2825 gnd.n2824 0.152939
R13005 gnd.n2826 gnd.n2825 0.152939
R13006 gnd.n2827 gnd.n2826 0.152939
R13007 gnd.n2828 gnd.n2827 0.152939
R13008 gnd.n2829 gnd.n2828 0.152939
R13009 gnd.n2830 gnd.n2829 0.152939
R13010 gnd.n2831 gnd.n2830 0.152939
R13011 gnd.n2832 gnd.n2831 0.152939
R13012 gnd.n2833 gnd.n2832 0.152939
R13013 gnd.n2834 gnd.n2833 0.152939
R13014 gnd.n2835 gnd.n2834 0.152939
R13015 gnd.n2836 gnd.n2835 0.152939
R13016 gnd.n2837 gnd.n2836 0.152939
R13017 gnd.n2838 gnd.n2837 0.152939
R13018 gnd.n2839 gnd.n2838 0.152939
R13019 gnd.n2840 gnd.n2839 0.152939
R13020 gnd.n2841 gnd.n2840 0.152939
R13021 gnd.n2842 gnd.n2841 0.152939
R13022 gnd.n2846 gnd.n2842 0.152939
R13023 gnd.n2847 gnd.n2846 0.152939
R13024 gnd.n2847 gnd.n2804 0.152939
R13025 gnd.n2901 gnd.n2804 0.152939
R13026 gnd.n6642 gnd.n766 0.152939
R13027 gnd.n6650 gnd.n766 0.152939
R13028 gnd.n6651 gnd.n6650 0.152939
R13029 gnd.n6652 gnd.n6651 0.152939
R13030 gnd.n6652 gnd.n760 0.152939
R13031 gnd.n6660 gnd.n760 0.152939
R13032 gnd.n6661 gnd.n6660 0.152939
R13033 gnd.n6662 gnd.n6661 0.152939
R13034 gnd.n6662 gnd.n754 0.152939
R13035 gnd.n6670 gnd.n754 0.152939
R13036 gnd.n6671 gnd.n6670 0.152939
R13037 gnd.n6672 gnd.n6671 0.152939
R13038 gnd.n6672 gnd.n748 0.152939
R13039 gnd.n6680 gnd.n748 0.152939
R13040 gnd.n6681 gnd.n6680 0.152939
R13041 gnd.n6682 gnd.n6681 0.152939
R13042 gnd.n6682 gnd.n742 0.152939
R13043 gnd.n6690 gnd.n742 0.152939
R13044 gnd.n6691 gnd.n6690 0.152939
R13045 gnd.n6692 gnd.n6691 0.152939
R13046 gnd.n6692 gnd.n736 0.152939
R13047 gnd.n6700 gnd.n736 0.152939
R13048 gnd.n6701 gnd.n6700 0.152939
R13049 gnd.n6702 gnd.n6701 0.152939
R13050 gnd.n6702 gnd.n730 0.152939
R13051 gnd.n6710 gnd.n730 0.152939
R13052 gnd.n6711 gnd.n6710 0.152939
R13053 gnd.n6712 gnd.n6711 0.152939
R13054 gnd.n6712 gnd.n724 0.152939
R13055 gnd.n6720 gnd.n724 0.152939
R13056 gnd.n6721 gnd.n6720 0.152939
R13057 gnd.n6722 gnd.n6721 0.152939
R13058 gnd.n6722 gnd.n718 0.152939
R13059 gnd.n6730 gnd.n718 0.152939
R13060 gnd.n6731 gnd.n6730 0.152939
R13061 gnd.n6732 gnd.n6731 0.152939
R13062 gnd.n6732 gnd.n712 0.152939
R13063 gnd.n6740 gnd.n712 0.152939
R13064 gnd.n6741 gnd.n6740 0.152939
R13065 gnd.n6742 gnd.n6741 0.152939
R13066 gnd.n6742 gnd.n706 0.152939
R13067 gnd.n6750 gnd.n706 0.152939
R13068 gnd.n6751 gnd.n6750 0.152939
R13069 gnd.n6752 gnd.n6751 0.152939
R13070 gnd.n6752 gnd.n700 0.152939
R13071 gnd.n6760 gnd.n700 0.152939
R13072 gnd.n6761 gnd.n6760 0.152939
R13073 gnd.n6762 gnd.n6761 0.152939
R13074 gnd.n6762 gnd.n694 0.152939
R13075 gnd.n6770 gnd.n694 0.152939
R13076 gnd.n6771 gnd.n6770 0.152939
R13077 gnd.n6772 gnd.n6771 0.152939
R13078 gnd.n6772 gnd.n688 0.152939
R13079 gnd.n6780 gnd.n688 0.152939
R13080 gnd.n6781 gnd.n6780 0.152939
R13081 gnd.n6782 gnd.n6781 0.152939
R13082 gnd.n6782 gnd.n682 0.152939
R13083 gnd.n6790 gnd.n682 0.152939
R13084 gnd.n6791 gnd.n6790 0.152939
R13085 gnd.n6792 gnd.n6791 0.152939
R13086 gnd.n6792 gnd.n676 0.152939
R13087 gnd.n6800 gnd.n676 0.152939
R13088 gnd.n6801 gnd.n6800 0.152939
R13089 gnd.n6802 gnd.n6801 0.152939
R13090 gnd.n6802 gnd.n670 0.152939
R13091 gnd.n6810 gnd.n670 0.152939
R13092 gnd.n6811 gnd.n6810 0.152939
R13093 gnd.n6812 gnd.n6811 0.152939
R13094 gnd.n6812 gnd.n664 0.152939
R13095 gnd.n6820 gnd.n664 0.152939
R13096 gnd.n6821 gnd.n6820 0.152939
R13097 gnd.n6822 gnd.n6821 0.152939
R13098 gnd.n6822 gnd.n658 0.152939
R13099 gnd.n6830 gnd.n658 0.152939
R13100 gnd.n6831 gnd.n6830 0.152939
R13101 gnd.n6832 gnd.n6831 0.152939
R13102 gnd.n6832 gnd.n652 0.152939
R13103 gnd.n6840 gnd.n652 0.152939
R13104 gnd.n6841 gnd.n6840 0.152939
R13105 gnd.n6842 gnd.n6841 0.152939
R13106 gnd.n6842 gnd.n646 0.152939
R13107 gnd.n6850 gnd.n646 0.152939
R13108 gnd.n6851 gnd.n6850 0.152939
R13109 gnd.n6852 gnd.n6851 0.152939
R13110 gnd.n6852 gnd.n640 0.152939
R13111 gnd.n6860 gnd.n640 0.152939
R13112 gnd.n6861 gnd.n6860 0.152939
R13113 gnd.n6862 gnd.n6861 0.152939
R13114 gnd.n6862 gnd.n634 0.152939
R13115 gnd.n6870 gnd.n634 0.152939
R13116 gnd.n6871 gnd.n6870 0.152939
R13117 gnd.n6872 gnd.n6871 0.152939
R13118 gnd.n6872 gnd.n628 0.152939
R13119 gnd.n6880 gnd.n628 0.152939
R13120 gnd.n6881 gnd.n6880 0.152939
R13121 gnd.n6882 gnd.n6881 0.152939
R13122 gnd.n6882 gnd.n622 0.152939
R13123 gnd.n6890 gnd.n622 0.152939
R13124 gnd.n6891 gnd.n6890 0.152939
R13125 gnd.n6892 gnd.n6891 0.152939
R13126 gnd.n6892 gnd.n616 0.152939
R13127 gnd.n6900 gnd.n616 0.152939
R13128 gnd.n6901 gnd.n6900 0.152939
R13129 gnd.n6902 gnd.n6901 0.152939
R13130 gnd.n6902 gnd.n610 0.152939
R13131 gnd.n6910 gnd.n610 0.152939
R13132 gnd.n6911 gnd.n6910 0.152939
R13133 gnd.n6912 gnd.n6911 0.152939
R13134 gnd.n6912 gnd.n604 0.152939
R13135 gnd.n6920 gnd.n604 0.152939
R13136 gnd.n6921 gnd.n6920 0.152939
R13137 gnd.n6922 gnd.n6921 0.152939
R13138 gnd.n6922 gnd.n598 0.152939
R13139 gnd.n6930 gnd.n598 0.152939
R13140 gnd.n6931 gnd.n6930 0.152939
R13141 gnd.n6932 gnd.n6931 0.152939
R13142 gnd.n6932 gnd.n592 0.152939
R13143 gnd.n6940 gnd.n592 0.152939
R13144 gnd.n6941 gnd.n6940 0.152939
R13145 gnd.n6942 gnd.n6941 0.152939
R13146 gnd.n6942 gnd.n586 0.152939
R13147 gnd.n6950 gnd.n586 0.152939
R13148 gnd.n6951 gnd.n6950 0.152939
R13149 gnd.n6952 gnd.n6951 0.152939
R13150 gnd.n6952 gnd.n580 0.152939
R13151 gnd.n6960 gnd.n580 0.152939
R13152 gnd.n6961 gnd.n6960 0.152939
R13153 gnd.n6962 gnd.n6961 0.152939
R13154 gnd.n6962 gnd.n574 0.152939
R13155 gnd.n6970 gnd.n574 0.152939
R13156 gnd.n6971 gnd.n6970 0.152939
R13157 gnd.n6972 gnd.n6971 0.152939
R13158 gnd.n6972 gnd.n568 0.152939
R13159 gnd.n6980 gnd.n568 0.152939
R13160 gnd.n6981 gnd.n6980 0.152939
R13161 gnd.n6982 gnd.n6981 0.152939
R13162 gnd.n6982 gnd.n562 0.152939
R13163 gnd.n6990 gnd.n562 0.152939
R13164 gnd.n6991 gnd.n6990 0.152939
R13165 gnd.n6992 gnd.n6991 0.152939
R13166 gnd.n6992 gnd.n556 0.152939
R13167 gnd.n7000 gnd.n556 0.152939
R13168 gnd.n7001 gnd.n7000 0.152939
R13169 gnd.n7002 gnd.n7001 0.152939
R13170 gnd.n7002 gnd.n550 0.152939
R13171 gnd.n7010 gnd.n550 0.152939
R13172 gnd.n7011 gnd.n7010 0.152939
R13173 gnd.n7012 gnd.n7011 0.152939
R13174 gnd.n7012 gnd.n544 0.152939
R13175 gnd.n7020 gnd.n544 0.152939
R13176 gnd.n7021 gnd.n7020 0.152939
R13177 gnd.n7022 gnd.n7021 0.152939
R13178 gnd.n7022 gnd.n538 0.152939
R13179 gnd.n7030 gnd.n538 0.152939
R13180 gnd.n7031 gnd.n7030 0.152939
R13181 gnd.n7032 gnd.n7031 0.152939
R13182 gnd.n7032 gnd.n532 0.152939
R13183 gnd.n7040 gnd.n532 0.152939
R13184 gnd.n7041 gnd.n7040 0.152939
R13185 gnd.n7042 gnd.n7041 0.152939
R13186 gnd.n7042 gnd.n526 0.152939
R13187 gnd.n7050 gnd.n526 0.152939
R13188 gnd.n7051 gnd.n7050 0.152939
R13189 gnd.n7053 gnd.n7051 0.152939
R13190 gnd.n7053 gnd.n7052 0.152939
R13191 gnd.n7052 gnd.n520 0.152939
R13192 gnd.n7062 gnd.n520 0.152939
R13193 gnd.n7063 gnd.n515 0.152939
R13194 gnd.n7071 gnd.n515 0.152939
R13195 gnd.n7072 gnd.n7071 0.152939
R13196 gnd.n7073 gnd.n7072 0.152939
R13197 gnd.n7073 gnd.n509 0.152939
R13198 gnd.n7081 gnd.n509 0.152939
R13199 gnd.n7082 gnd.n7081 0.152939
R13200 gnd.n7083 gnd.n7082 0.152939
R13201 gnd.n7083 gnd.n503 0.152939
R13202 gnd.n7091 gnd.n503 0.152939
R13203 gnd.n7092 gnd.n7091 0.152939
R13204 gnd.n7093 gnd.n7092 0.152939
R13205 gnd.n7093 gnd.n497 0.152939
R13206 gnd.n7101 gnd.n497 0.152939
R13207 gnd.n7102 gnd.n7101 0.152939
R13208 gnd.n7103 gnd.n7102 0.152939
R13209 gnd.n7103 gnd.n491 0.152939
R13210 gnd.n7111 gnd.n491 0.152939
R13211 gnd.n7112 gnd.n7111 0.152939
R13212 gnd.n7113 gnd.n7112 0.152939
R13213 gnd.n7113 gnd.n485 0.152939
R13214 gnd.n7121 gnd.n485 0.152939
R13215 gnd.n7122 gnd.n7121 0.152939
R13216 gnd.n7123 gnd.n7122 0.152939
R13217 gnd.n7123 gnd.n479 0.152939
R13218 gnd.n7131 gnd.n479 0.152939
R13219 gnd.n7132 gnd.n7131 0.152939
R13220 gnd.n7133 gnd.n7132 0.152939
R13221 gnd.n7133 gnd.n473 0.152939
R13222 gnd.n7141 gnd.n473 0.152939
R13223 gnd.n7142 gnd.n7141 0.152939
R13224 gnd.n7143 gnd.n7142 0.152939
R13225 gnd.n7143 gnd.n467 0.152939
R13226 gnd.n7151 gnd.n467 0.152939
R13227 gnd.n7152 gnd.n7151 0.152939
R13228 gnd.n7153 gnd.n7152 0.152939
R13229 gnd.n7153 gnd.n461 0.152939
R13230 gnd.n7161 gnd.n461 0.152939
R13231 gnd.n7162 gnd.n7161 0.152939
R13232 gnd.n7163 gnd.n7162 0.152939
R13233 gnd.n7163 gnd.n455 0.152939
R13234 gnd.n7171 gnd.n455 0.152939
R13235 gnd.n7172 gnd.n7171 0.152939
R13236 gnd.n7173 gnd.n7172 0.152939
R13237 gnd.n7173 gnd.n449 0.152939
R13238 gnd.n7181 gnd.n449 0.152939
R13239 gnd.n7182 gnd.n7181 0.152939
R13240 gnd.n7183 gnd.n7182 0.152939
R13241 gnd.n7183 gnd.n443 0.152939
R13242 gnd.n7191 gnd.n443 0.152939
R13243 gnd.n7192 gnd.n7191 0.152939
R13244 gnd.n7193 gnd.n7192 0.152939
R13245 gnd.n7193 gnd.n437 0.152939
R13246 gnd.n7201 gnd.n437 0.152939
R13247 gnd.n7202 gnd.n7201 0.152939
R13248 gnd.n7203 gnd.n7202 0.152939
R13249 gnd.n7203 gnd.n431 0.152939
R13250 gnd.n7211 gnd.n431 0.152939
R13251 gnd.n7212 gnd.n7211 0.152939
R13252 gnd.n7213 gnd.n7212 0.152939
R13253 gnd.n7213 gnd.n425 0.152939
R13254 gnd.n7221 gnd.n425 0.152939
R13255 gnd.n7222 gnd.n7221 0.152939
R13256 gnd.n7223 gnd.n7222 0.152939
R13257 gnd.n7223 gnd.n419 0.152939
R13258 gnd.n7231 gnd.n419 0.152939
R13259 gnd.n7232 gnd.n7231 0.152939
R13260 gnd.n7233 gnd.n7232 0.152939
R13261 gnd.n7233 gnd.n413 0.152939
R13262 gnd.n7241 gnd.n413 0.152939
R13263 gnd.n7242 gnd.n7241 0.152939
R13264 gnd.n7243 gnd.n7242 0.152939
R13265 gnd.n7243 gnd.n407 0.152939
R13266 gnd.n7251 gnd.n407 0.152939
R13267 gnd.n7252 gnd.n7251 0.152939
R13268 gnd.n7253 gnd.n7252 0.152939
R13269 gnd.n7253 gnd.n401 0.152939
R13270 gnd.n7261 gnd.n401 0.152939
R13271 gnd.n7262 gnd.n7261 0.152939
R13272 gnd.n7263 gnd.n7262 0.152939
R13273 gnd.n7263 gnd.n395 0.152939
R13274 gnd.n7272 gnd.n395 0.152939
R13275 gnd.n7273 gnd.n7272 0.152939
R13276 gnd.n7275 gnd.n7273 0.152939
R13277 gnd.n389 gnd.n388 0.152939
R13278 gnd.n390 gnd.n389 0.152939
R13279 gnd.n391 gnd.n390 0.152939
R13280 gnd.n7274 gnd.n391 0.152939
R13281 gnd.n118 gnd.n93 0.152939
R13282 gnd.n119 gnd.n118 0.152939
R13283 gnd.n120 gnd.n119 0.152939
R13284 gnd.n137 gnd.n120 0.152939
R13285 gnd.n138 gnd.n137 0.152939
R13286 gnd.n139 gnd.n138 0.152939
R13287 gnd.n140 gnd.n139 0.152939
R13288 gnd.n155 gnd.n140 0.152939
R13289 gnd.n156 gnd.n155 0.152939
R13290 gnd.n157 gnd.n156 0.152939
R13291 gnd.n158 gnd.n157 0.152939
R13292 gnd.n175 gnd.n158 0.152939
R13293 gnd.n176 gnd.n175 0.152939
R13294 gnd.n177 gnd.n176 0.152939
R13295 gnd.n178 gnd.n177 0.152939
R13296 gnd.n194 gnd.n178 0.152939
R13297 gnd.n195 gnd.n194 0.152939
R13298 gnd.n196 gnd.n195 0.152939
R13299 gnd.n197 gnd.n196 0.152939
R13300 gnd.n212 gnd.n197 0.152939
R13301 gnd.n7561 gnd.n212 0.152939
R13302 gnd.n7642 gnd.n80 0.152939
R13303 gnd.n361 gnd.n80 0.152939
R13304 gnd.n7327 gnd.n361 0.152939
R13305 gnd.n7328 gnd.n7327 0.152939
R13306 gnd.n7330 gnd.n7328 0.152939
R13307 gnd.n7330 gnd.n7329 0.152939
R13308 gnd.n7329 gnd.n357 0.152939
R13309 gnd.n357 gnd.n355 0.152939
R13310 gnd.n7349 gnd.n355 0.152939
R13311 gnd.n7350 gnd.n7349 0.152939
R13312 gnd.n7351 gnd.n7350 0.152939
R13313 gnd.n7352 gnd.n7351 0.152939
R13314 gnd.n7353 gnd.n7352 0.152939
R13315 gnd.n7354 gnd.n7353 0.152939
R13316 gnd.n7355 gnd.n7354 0.152939
R13317 gnd.n7356 gnd.n7355 0.152939
R13318 gnd.n7357 gnd.n7356 0.152939
R13319 gnd.n7358 gnd.n7357 0.152939
R13320 gnd.n7359 gnd.n7358 0.152939
R13321 gnd.n7360 gnd.n7359 0.152939
R13322 gnd.n7361 gnd.n7360 0.152939
R13323 gnd.n7362 gnd.n7361 0.152939
R13324 gnd.n7364 gnd.n7362 0.152939
R13325 gnd.n7364 gnd.n7363 0.152939
R13326 gnd.n7363 gnd.n350 0.152939
R13327 gnd.n7417 gnd.n350 0.152939
R13328 gnd.n7450 gnd.n316 0.152939
R13329 gnd.n318 gnd.n316 0.152939
R13330 gnd.n322 gnd.n318 0.152939
R13331 gnd.n323 gnd.n322 0.152939
R13332 gnd.n324 gnd.n323 0.152939
R13333 gnd.n325 gnd.n324 0.152939
R13334 gnd.n329 gnd.n325 0.152939
R13335 gnd.n330 gnd.n329 0.152939
R13336 gnd.n331 gnd.n330 0.152939
R13337 gnd.n332 gnd.n331 0.152939
R13338 gnd.n336 gnd.n332 0.152939
R13339 gnd.n337 gnd.n336 0.152939
R13340 gnd.n338 gnd.n337 0.152939
R13341 gnd.n339 gnd.n338 0.152939
R13342 gnd.n343 gnd.n339 0.152939
R13343 gnd.n344 gnd.n343 0.152939
R13344 gnd.n7419 gnd.n344 0.152939
R13345 gnd.n7419 gnd.n7418 0.152939
R13346 gnd.n7560 gnd.n213 0.152939
R13347 gnd.n215 gnd.n213 0.152939
R13348 gnd.n219 gnd.n215 0.152939
R13349 gnd.n220 gnd.n219 0.152939
R13350 gnd.n221 gnd.n220 0.152939
R13351 gnd.n222 gnd.n221 0.152939
R13352 gnd.n226 gnd.n222 0.152939
R13353 gnd.n227 gnd.n226 0.152939
R13354 gnd.n228 gnd.n227 0.152939
R13355 gnd.n229 gnd.n228 0.152939
R13356 gnd.n233 gnd.n229 0.152939
R13357 gnd.n234 gnd.n233 0.152939
R13358 gnd.n235 gnd.n234 0.152939
R13359 gnd.n236 gnd.n235 0.152939
R13360 gnd.n240 gnd.n236 0.152939
R13361 gnd.n241 gnd.n240 0.152939
R13362 gnd.n242 gnd.n241 0.152939
R13363 gnd.n243 gnd.n242 0.152939
R13364 gnd.n247 gnd.n243 0.152939
R13365 gnd.n248 gnd.n247 0.152939
R13366 gnd.n249 gnd.n248 0.152939
R13367 gnd.n250 gnd.n249 0.152939
R13368 gnd.n254 gnd.n250 0.152939
R13369 gnd.n255 gnd.n254 0.152939
R13370 gnd.n256 gnd.n255 0.152939
R13371 gnd.n257 gnd.n256 0.152939
R13372 gnd.n261 gnd.n257 0.152939
R13373 gnd.n262 gnd.n261 0.152939
R13374 gnd.n263 gnd.n262 0.152939
R13375 gnd.n264 gnd.n263 0.152939
R13376 gnd.n268 gnd.n264 0.152939
R13377 gnd.n269 gnd.n268 0.152939
R13378 gnd.n270 gnd.n269 0.152939
R13379 gnd.n271 gnd.n270 0.152939
R13380 gnd.n275 gnd.n271 0.152939
R13381 gnd.n276 gnd.n275 0.152939
R13382 gnd.n7491 gnd.n276 0.152939
R13383 gnd.n7491 gnd.n7490 0.152939
R13384 gnd.n7490 gnd.n7489 0.152939
R13385 gnd.n7489 gnd.n280 0.152939
R13386 gnd.n286 gnd.n280 0.152939
R13387 gnd.n287 gnd.n286 0.152939
R13388 gnd.n288 gnd.n287 0.152939
R13389 gnd.n289 gnd.n288 0.152939
R13390 gnd.n293 gnd.n289 0.152939
R13391 gnd.n294 gnd.n293 0.152939
R13392 gnd.n295 gnd.n294 0.152939
R13393 gnd.n296 gnd.n295 0.152939
R13394 gnd.n300 gnd.n296 0.152939
R13395 gnd.n301 gnd.n300 0.152939
R13396 gnd.n302 gnd.n301 0.152939
R13397 gnd.n303 gnd.n302 0.152939
R13398 gnd.n307 gnd.n303 0.152939
R13399 gnd.n308 gnd.n307 0.152939
R13400 gnd.n309 gnd.n308 0.152939
R13401 gnd.n310 gnd.n309 0.152939
R13402 gnd.n315 gnd.n310 0.152939
R13403 gnd.n7452 gnd.n315 0.152939
R13404 gnd.n5752 gnd.n5751 0.152939
R13405 gnd.n5752 gnd.n5748 0.152939
R13406 gnd.n5760 gnd.n5748 0.152939
R13407 gnd.n5761 gnd.n5760 0.152939
R13408 gnd.n5762 gnd.n5761 0.152939
R13409 gnd.n5762 gnd.n5744 0.152939
R13410 gnd.n5770 gnd.n5744 0.152939
R13411 gnd.n5771 gnd.n5770 0.152939
R13412 gnd.n5772 gnd.n5771 0.152939
R13413 gnd.n5772 gnd.n5740 0.152939
R13414 gnd.n5780 gnd.n5740 0.152939
R13415 gnd.n5781 gnd.n5780 0.152939
R13416 gnd.n5782 gnd.n5781 0.152939
R13417 gnd.n5782 gnd.n5736 0.152939
R13418 gnd.n5790 gnd.n5736 0.152939
R13419 gnd.n5791 gnd.n5790 0.152939
R13420 gnd.n5792 gnd.n5791 0.152939
R13421 gnd.n5792 gnd.n5732 0.152939
R13422 gnd.n5803 gnd.n5732 0.152939
R13423 gnd.n5804 gnd.n5803 0.152939
R13424 gnd.n5805 gnd.n5804 0.152939
R13425 gnd.n5805 gnd.n5728 0.152939
R13426 gnd.n5813 gnd.n5728 0.152939
R13427 gnd.n5814 gnd.n5813 0.152939
R13428 gnd.n5816 gnd.n5814 0.152939
R13429 gnd.n5826 gnd.n1530 0.152939
R13430 gnd.n5827 gnd.n5826 0.152939
R13431 gnd.n5828 gnd.n5827 0.152939
R13432 gnd.n5828 gnd.n1526 0.152939
R13433 gnd.n5836 gnd.n1526 0.152939
R13434 gnd.n5837 gnd.n5836 0.152939
R13435 gnd.n5838 gnd.n5837 0.152939
R13436 gnd.n5838 gnd.n1522 0.152939
R13437 gnd.n5848 gnd.n1522 0.152939
R13438 gnd.n5849 gnd.n5848 0.152939
R13439 gnd.n5850 gnd.n5849 0.152939
R13440 gnd.n5850 gnd.n1518 0.152939
R13441 gnd.n5858 gnd.n1518 0.152939
R13442 gnd.n5859 gnd.n5858 0.152939
R13443 gnd.n5860 gnd.n5859 0.152939
R13444 gnd.n5860 gnd.n1514 0.152939
R13445 gnd.n5868 gnd.n1514 0.152939
R13446 gnd.n5869 gnd.n5868 0.152939
R13447 gnd.n5870 gnd.n5869 0.152939
R13448 gnd.n5870 gnd.n1510 0.152939
R13449 gnd.n5878 gnd.n1510 0.152939
R13450 gnd.n5879 gnd.n5878 0.152939
R13451 gnd.n5880 gnd.n5879 0.152939
R13452 gnd.n5880 gnd.n1506 0.152939
R13453 gnd.n5888 gnd.n1506 0.152939
R13454 gnd.n5889 gnd.n5888 0.152939
R13455 gnd.n5891 gnd.n5889 0.152939
R13456 gnd.n5891 gnd.n5890 0.152939
R13457 gnd.n5890 gnd.n1499 0.152939
R13458 gnd.n5900 gnd.n1499 0.152939
R13459 gnd.n1345 gnd.n1344 0.152939
R13460 gnd.n1346 gnd.n1345 0.152939
R13461 gnd.n1366 gnd.n1346 0.152939
R13462 gnd.n1367 gnd.n1366 0.152939
R13463 gnd.n1368 gnd.n1367 0.152939
R13464 gnd.n1369 gnd.n1368 0.152939
R13465 gnd.n1386 gnd.n1369 0.152939
R13466 gnd.n1387 gnd.n1386 0.152939
R13467 gnd.n1388 gnd.n1387 0.152939
R13468 gnd.n1389 gnd.n1388 0.152939
R13469 gnd.n1406 gnd.n1389 0.152939
R13470 gnd.n1407 gnd.n1406 0.152939
R13471 gnd.n1408 gnd.n1407 0.152939
R13472 gnd.n1409 gnd.n1408 0.152939
R13473 gnd.n1426 gnd.n1409 0.152939
R13474 gnd.n1427 gnd.n1426 0.152939
R13475 gnd.n1428 gnd.n1427 0.152939
R13476 gnd.n1429 gnd.n1428 0.152939
R13477 gnd.n1446 gnd.n1429 0.152939
R13478 gnd.n1447 gnd.n1446 0.152939
R13479 gnd.n1447 gnd.n94 0.152939
R13480 gnd.n4284 gnd.n4283 0.152939
R13481 gnd.n4285 gnd.n4284 0.152939
R13482 gnd.n4285 gnd.n2123 0.152939
R13483 gnd.n4291 gnd.n2123 0.152939
R13484 gnd.n4292 gnd.n4291 0.152939
R13485 gnd.n4293 gnd.n4292 0.152939
R13486 gnd.n4294 gnd.n4293 0.152939
R13487 gnd.n4295 gnd.n4294 0.152939
R13488 gnd.n4298 gnd.n4295 0.152939
R13489 gnd.n4299 gnd.n4298 0.152939
R13490 gnd.n4300 gnd.n4299 0.152939
R13491 gnd.n4301 gnd.n4300 0.152939
R13492 gnd.n4302 gnd.n4301 0.152939
R13493 gnd.n4302 gnd.n2098 0.152939
R13494 gnd.n4378 gnd.n2098 0.152939
R13495 gnd.n4379 gnd.n4378 0.152939
R13496 gnd.n4380 gnd.n4379 0.152939
R13497 gnd.n4380 gnd.n2094 0.152939
R13498 gnd.n4386 gnd.n2094 0.152939
R13499 gnd.n4387 gnd.n4386 0.152939
R13500 gnd.n4388 gnd.n4387 0.152939
R13501 gnd.n4388 gnd.n2090 0.152939
R13502 gnd.n4396 gnd.n2090 0.152939
R13503 gnd.n4397 gnd.n4396 0.152939
R13504 gnd.n4398 gnd.n4397 0.152939
R13505 gnd.n4398 gnd.n2065 0.152939
R13506 gnd.n4680 gnd.n2065 0.152939
R13507 gnd.n4681 gnd.n4680 0.152939
R13508 gnd.n4682 gnd.n4681 0.152939
R13509 gnd.n4683 gnd.n4682 0.152939
R13510 gnd.n4683 gnd.n2040 0.152939
R13511 gnd.n4712 gnd.n2040 0.152939
R13512 gnd.n4713 gnd.n4712 0.152939
R13513 gnd.n4714 gnd.n4713 0.152939
R13514 gnd.n4716 gnd.n4714 0.152939
R13515 gnd.n4716 gnd.n4715 0.152939
R13516 gnd.n4715 gnd.n1216 0.152939
R13517 gnd.n1217 gnd.n1216 0.152939
R13518 gnd.n1218 gnd.n1217 0.152939
R13519 gnd.n4752 gnd.n1218 0.152939
R13520 gnd.n4753 gnd.n4752 0.152939
R13521 gnd.n4753 gnd.n1914 0.152939
R13522 gnd.n4794 gnd.n1914 0.152939
R13523 gnd.n4795 gnd.n4794 0.152939
R13524 gnd.n4796 gnd.n4795 0.152939
R13525 gnd.n4796 gnd.n1896 0.152939
R13526 gnd.n4836 gnd.n1896 0.152939
R13527 gnd.n4837 gnd.n4836 0.152939
R13528 gnd.n4838 gnd.n4837 0.152939
R13529 gnd.n4839 gnd.n4838 0.152939
R13530 gnd.n4839 gnd.n1870 0.152939
R13531 gnd.n4898 gnd.n1870 0.152939
R13532 gnd.n4899 gnd.n4898 0.152939
R13533 gnd.n4900 gnd.n4899 0.152939
R13534 gnd.n4900 gnd.n1852 0.152939
R13535 gnd.n4926 gnd.n1852 0.152939
R13536 gnd.n4927 gnd.n4926 0.152939
R13537 gnd.n4928 gnd.n4927 0.152939
R13538 gnd.n4929 gnd.n4928 0.152939
R13539 gnd.n4929 gnd.n1819 0.152939
R13540 gnd.n4976 gnd.n1819 0.152939
R13541 gnd.n4977 gnd.n4976 0.152939
R13542 gnd.n4978 gnd.n4977 0.152939
R13543 gnd.n4978 gnd.n1796 0.152939
R13544 gnd.n5016 gnd.n1796 0.152939
R13545 gnd.n5017 gnd.n5016 0.152939
R13546 gnd.n5018 gnd.n5017 0.152939
R13547 gnd.n5018 gnd.n1774 0.152939
R13548 gnd.n5073 gnd.n1774 0.152939
R13549 gnd.n5074 gnd.n5073 0.152939
R13550 gnd.n5075 gnd.n5074 0.152939
R13551 gnd.n5075 gnd.n1754 0.152939
R13552 gnd.n5098 gnd.n1754 0.152939
R13553 gnd.n5099 gnd.n5098 0.152939
R13554 gnd.n5100 gnd.n5099 0.152939
R13555 gnd.n5100 gnd.n1734 0.152939
R13556 gnd.n5158 gnd.n1734 0.152939
R13557 gnd.n5159 gnd.n5158 0.152939
R13558 gnd.n5160 gnd.n5159 0.152939
R13559 gnd.n5160 gnd.n1712 0.152939
R13560 gnd.n5187 gnd.n1712 0.152939
R13561 gnd.n5188 gnd.n5187 0.152939
R13562 gnd.n5189 gnd.n5188 0.152939
R13563 gnd.n5190 gnd.n5189 0.152939
R13564 gnd.n5190 gnd.n1684 0.152939
R13565 gnd.n5238 gnd.n1684 0.152939
R13566 gnd.n5239 gnd.n5238 0.152939
R13567 gnd.n5240 gnd.n5239 0.152939
R13568 gnd.n5240 gnd.n1664 0.152939
R13569 gnd.n5264 gnd.n1664 0.152939
R13570 gnd.n5265 gnd.n5264 0.152939
R13571 gnd.n5266 gnd.n5265 0.152939
R13572 gnd.n5267 gnd.n5266 0.152939
R13573 gnd.n5267 gnd.n1634 0.152939
R13574 gnd.n5308 gnd.n1634 0.152939
R13575 gnd.n5309 gnd.n5308 0.152939
R13576 gnd.n5310 gnd.n5309 0.152939
R13577 gnd.n5312 gnd.n5310 0.152939
R13578 gnd.n5312 gnd.n5311 0.152939
R13579 gnd.n5311 gnd.n1585 0.152939
R13580 gnd.n1586 gnd.n1585 0.152939
R13581 gnd.n1587 gnd.n1586 0.152939
R13582 gnd.n1596 gnd.n1587 0.152939
R13583 gnd.n1597 gnd.n1596 0.152939
R13584 gnd.n1598 gnd.n1597 0.152939
R13585 gnd.n1599 gnd.n1598 0.152939
R13586 gnd.n1600 gnd.n1599 0.152939
R13587 gnd.n1602 gnd.n1600 0.152939
R13588 gnd.n1602 gnd.n1601 0.152939
R13589 gnd.n1601 gnd.n1323 0.152939
R13590 gnd.n1324 gnd.n1323 0.152939
R13591 gnd.n1325 gnd.n1324 0.152939
R13592 gnd.n1331 gnd.n1325 0.152939
R13593 gnd.n1332 gnd.n1331 0.152939
R13594 gnd.n1333 gnd.n1332 0.152939
R13595 gnd.n1334 gnd.n1333 0.152939
R13596 gnd.n5944 gnd.n1334 0.152939
R13597 gnd.n5947 gnd.n5944 0.152939
R13598 gnd.n5948 gnd.n5947 0.152939
R13599 gnd.n5949 gnd.n5948 0.152939
R13600 gnd.n5949 gnd.n5940 0.152939
R13601 gnd.n5955 gnd.n5940 0.152939
R13602 gnd.n5956 gnd.n5955 0.152939
R13603 gnd.n5957 gnd.n5956 0.152939
R13604 gnd.n5957 gnd.n1485 0.152939
R13605 gnd.n5963 gnd.n1485 0.152939
R13606 gnd.n5964 gnd.n5963 0.152939
R13607 gnd.n5965 gnd.n5964 0.152939
R13608 gnd.n5966 gnd.n5965 0.152939
R13609 gnd.n5967 gnd.n5966 0.152939
R13610 gnd.n5970 gnd.n5967 0.152939
R13611 gnd.n5971 gnd.n5970 0.152939
R13612 gnd.n5972 gnd.n5971 0.152939
R13613 gnd.n5973 gnd.n5972 0.152939
R13614 gnd.n5976 gnd.n5973 0.152939
R13615 gnd.n5976 gnd.n5975 0.152939
R13616 gnd.n5975 gnd.n5974 0.152939
R13617 gnd.n3885 gnd.n3871 0.152939
R13618 gnd.n3872 gnd.n3871 0.152939
R13619 gnd.n3873 gnd.n3872 0.152939
R13620 gnd.n3874 gnd.n3873 0.152939
R13621 gnd.n3875 gnd.n3874 0.152939
R13622 gnd.n3875 gnd.n2228 0.152939
R13623 gnd.n4090 gnd.n2228 0.152939
R13624 gnd.n4091 gnd.n4090 0.152939
R13625 gnd.n4092 gnd.n4091 0.152939
R13626 gnd.n4093 gnd.n4092 0.152939
R13627 gnd.n4094 gnd.n4093 0.152939
R13628 gnd.n4094 gnd.n2203 0.152939
R13629 gnd.n4125 gnd.n2203 0.152939
R13630 gnd.n4126 gnd.n4125 0.152939
R13631 gnd.n4127 gnd.n4126 0.152939
R13632 gnd.n4128 gnd.n4127 0.152939
R13633 gnd.n4130 gnd.n4128 0.152939
R13634 gnd.n4130 gnd.n4129 0.152939
R13635 gnd.n4129 gnd.n2175 0.152939
R13636 gnd.n2176 gnd.n2175 0.152939
R13637 gnd.n2177 gnd.n2176 0.152939
R13638 gnd.n4171 gnd.n2177 0.152939
R13639 gnd.n4172 gnd.n4171 0.152939
R13640 gnd.n4173 gnd.n4172 0.152939
R13641 gnd.n4173 gnd.n2151 0.152939
R13642 gnd.n4230 gnd.n2151 0.152939
R13643 gnd.n3924 gnd.n3852 0.152939
R13644 gnd.n3853 gnd.n3852 0.152939
R13645 gnd.n3854 gnd.n3853 0.152939
R13646 gnd.n3855 gnd.n3854 0.152939
R13647 gnd.n3856 gnd.n3855 0.152939
R13648 gnd.n3857 gnd.n3856 0.152939
R13649 gnd.n3858 gnd.n3857 0.152939
R13650 gnd.n3859 gnd.n3858 0.152939
R13651 gnd.n3860 gnd.n3859 0.152939
R13652 gnd.n3861 gnd.n3860 0.152939
R13653 gnd.n3862 gnd.n3861 0.152939
R13654 gnd.n3863 gnd.n3862 0.152939
R13655 gnd.n3864 gnd.n3863 0.152939
R13656 gnd.n3865 gnd.n3864 0.152939
R13657 gnd.n3866 gnd.n3865 0.152939
R13658 gnd.n3889 gnd.n3866 0.152939
R13659 gnd.n3889 gnd.n3888 0.152939
R13660 gnd.n3888 gnd.n3887 0.152939
R13661 gnd.n997 gnd.n971 0.152939
R13662 gnd.n998 gnd.n997 0.152939
R13663 gnd.n999 gnd.n998 0.152939
R13664 gnd.n1017 gnd.n999 0.152939
R13665 gnd.n1018 gnd.n1017 0.152939
R13666 gnd.n1019 gnd.n1018 0.152939
R13667 gnd.n1020 gnd.n1019 0.152939
R13668 gnd.n1036 gnd.n1020 0.152939
R13669 gnd.n1037 gnd.n1036 0.152939
R13670 gnd.n1038 gnd.n1037 0.152939
R13671 gnd.n1039 gnd.n1038 0.152939
R13672 gnd.n1057 gnd.n1039 0.152939
R13673 gnd.n1058 gnd.n1057 0.152939
R13674 gnd.n1059 gnd.n1058 0.152939
R13675 gnd.n1060 gnd.n1059 0.152939
R13676 gnd.n1077 gnd.n1060 0.152939
R13677 gnd.n1078 gnd.n1077 0.152939
R13678 gnd.n1079 gnd.n1078 0.152939
R13679 gnd.n1080 gnd.n1079 0.152939
R13680 gnd.n1097 gnd.n1080 0.152939
R13681 gnd.n6378 gnd.n1097 0.152939
R13682 gnd.n6377 gnd.n1098 0.152939
R13683 gnd.n1103 gnd.n1098 0.152939
R13684 gnd.n1104 gnd.n1103 0.152939
R13685 gnd.n1105 gnd.n1104 0.152939
R13686 gnd.n1106 gnd.n1105 0.152939
R13687 gnd.n1107 gnd.n1106 0.152939
R13688 gnd.n1111 gnd.n1107 0.152939
R13689 gnd.n1112 gnd.n1111 0.152939
R13690 gnd.n1113 gnd.n1112 0.152939
R13691 gnd.n1114 gnd.n1113 0.152939
R13692 gnd.n1118 gnd.n1114 0.152939
R13693 gnd.n1119 gnd.n1118 0.152939
R13694 gnd.n1120 gnd.n1119 0.152939
R13695 gnd.n1121 gnd.n1120 0.152939
R13696 gnd.n1125 gnd.n1121 0.152939
R13697 gnd.n1126 gnd.n1125 0.152939
R13698 gnd.n1127 gnd.n1126 0.152939
R13699 gnd.n1130 gnd.n1127 0.152939
R13700 gnd.n1134 gnd.n1130 0.152939
R13701 gnd.n1135 gnd.n1134 0.152939
R13702 gnd.n1136 gnd.n1135 0.152939
R13703 gnd.n1137 gnd.n1136 0.152939
R13704 gnd.n1141 gnd.n1137 0.152939
R13705 gnd.n1142 gnd.n1141 0.152939
R13706 gnd.n1143 gnd.n1142 0.152939
R13707 gnd.n4456 gnd.n4455 0.152939
R13708 gnd.n4465 gnd.n4456 0.152939
R13709 gnd.n4466 gnd.n4465 0.152939
R13710 gnd.n4467 gnd.n4466 0.152939
R13711 gnd.n4467 gnd.n4451 0.152939
R13712 gnd.n4475 gnd.n4451 0.152939
R13713 gnd.n4476 gnd.n4475 0.152939
R13714 gnd.n4477 gnd.n4476 0.152939
R13715 gnd.n4477 gnd.n4445 0.152939
R13716 gnd.n4485 gnd.n4445 0.152939
R13717 gnd.n4486 gnd.n4485 0.152939
R13718 gnd.n4487 gnd.n4486 0.152939
R13719 gnd.n4487 gnd.n4441 0.152939
R13720 gnd.n4495 gnd.n4441 0.152939
R13721 gnd.n4496 gnd.n4495 0.152939
R13722 gnd.n4497 gnd.n4496 0.152939
R13723 gnd.n4497 gnd.n4437 0.152939
R13724 gnd.n4505 gnd.n4437 0.152939
R13725 gnd.n4506 gnd.n4505 0.152939
R13726 gnd.n4507 gnd.n4506 0.152939
R13727 gnd.n4507 gnd.n4433 0.152939
R13728 gnd.n4515 gnd.n4433 0.152939
R13729 gnd.n4516 gnd.n4515 0.152939
R13730 gnd.n4517 gnd.n4516 0.152939
R13731 gnd.n4517 gnd.n4429 0.152939
R13732 gnd.n4525 gnd.n4429 0.152939
R13733 gnd.n4526 gnd.n4525 0.152939
R13734 gnd.n4527 gnd.n4526 0.152939
R13735 gnd.n4527 gnd.n4423 0.152939
R13736 gnd.n4534 gnd.n4423 0.152939
R13737 gnd.n3790 gnd.n3789 0.152939
R13738 gnd.n3791 gnd.n3790 0.152939
R13739 gnd.n3792 gnd.n3791 0.152939
R13740 gnd.n3793 gnd.n3792 0.152939
R13741 gnd.n3794 gnd.n3793 0.152939
R13742 gnd.n3795 gnd.n3794 0.152939
R13743 gnd.n3796 gnd.n3795 0.152939
R13744 gnd.n3797 gnd.n3796 0.152939
R13745 gnd.n3798 gnd.n3797 0.152939
R13746 gnd.n3799 gnd.n3798 0.152939
R13747 gnd.n3800 gnd.n3799 0.152939
R13748 gnd.n3801 gnd.n3800 0.152939
R13749 gnd.n3802 gnd.n3801 0.152939
R13750 gnd.n3803 gnd.n3802 0.152939
R13751 gnd.n3804 gnd.n3803 0.152939
R13752 gnd.n3805 gnd.n3804 0.152939
R13753 gnd.n3806 gnd.n3805 0.152939
R13754 gnd.n3809 gnd.n3806 0.152939
R13755 gnd.n3810 gnd.n3809 0.152939
R13756 gnd.n3811 gnd.n3810 0.152939
R13757 gnd.n3812 gnd.n3811 0.152939
R13758 gnd.n3813 gnd.n3812 0.152939
R13759 gnd.n3814 gnd.n3813 0.152939
R13760 gnd.n3815 gnd.n3814 0.152939
R13761 gnd.n3816 gnd.n3815 0.152939
R13762 gnd.n3817 gnd.n3816 0.152939
R13763 gnd.n3818 gnd.n3817 0.152939
R13764 gnd.n3819 gnd.n3818 0.152939
R13765 gnd.n3820 gnd.n3819 0.152939
R13766 gnd.n3821 gnd.n3820 0.152939
R13767 gnd.n3822 gnd.n3821 0.152939
R13768 gnd.n3823 gnd.n3822 0.152939
R13769 gnd.n3824 gnd.n3823 0.152939
R13770 gnd.n3825 gnd.n3824 0.152939
R13771 gnd.n3826 gnd.n3825 0.152939
R13772 gnd.n3827 gnd.n3826 0.152939
R13773 gnd.n3828 gnd.n3827 0.152939
R13774 gnd.n3831 gnd.n3828 0.152939
R13775 gnd.n3832 gnd.n3831 0.152939
R13776 gnd.n3833 gnd.n3832 0.152939
R13777 gnd.n3834 gnd.n3833 0.152939
R13778 gnd.n3835 gnd.n3834 0.152939
R13779 gnd.n3836 gnd.n3835 0.152939
R13780 gnd.n3837 gnd.n3836 0.152939
R13781 gnd.n3838 gnd.n3837 0.152939
R13782 gnd.n3839 gnd.n3838 0.152939
R13783 gnd.n3840 gnd.n3839 0.152939
R13784 gnd.n3841 gnd.n3840 0.152939
R13785 gnd.n3842 gnd.n3841 0.152939
R13786 gnd.n3843 gnd.n3842 0.152939
R13787 gnd.n3844 gnd.n3843 0.152939
R13788 gnd.n3845 gnd.n3844 0.152939
R13789 gnd.n3846 gnd.n3845 0.152939
R13790 gnd.n3847 gnd.n3846 0.152939
R13791 gnd.n3848 gnd.n3847 0.152939
R13792 gnd.n3849 gnd.n3848 0.152939
R13793 gnd.n3927 gnd.n3849 0.152939
R13794 gnd.n3927 gnd.n3926 0.152939
R13795 gnd.n4056 gnd.n2256 0.152939
R13796 gnd.n4057 gnd.n4056 0.152939
R13797 gnd.n4058 gnd.n4057 0.152939
R13798 gnd.n4058 gnd.n2236 0.152939
R13799 gnd.n4080 gnd.n2236 0.152939
R13800 gnd.n4081 gnd.n4080 0.152939
R13801 gnd.n4082 gnd.n4081 0.152939
R13802 gnd.n4083 gnd.n4082 0.152939
R13803 gnd.n4083 gnd.n2210 0.152939
R13804 gnd.n4116 gnd.n2210 0.152939
R13805 gnd.n4117 gnd.n4116 0.152939
R13806 gnd.n4118 gnd.n4117 0.152939
R13807 gnd.n4118 gnd.n2188 0.152939
R13808 gnd.n4146 gnd.n2188 0.152939
R13809 gnd.n4147 gnd.n4146 0.152939
R13810 gnd.n4149 gnd.n4147 0.152939
R13811 gnd.n4149 gnd.n4148 0.152939
R13812 gnd.n4148 gnd.n949 0.152939
R13813 gnd.n950 gnd.n949 0.152939
R13814 gnd.n951 gnd.n950 0.152939
R13815 gnd.n972 gnd.n951 0.152939
R13816 gnd.n6470 gnd.n938 0.152939
R13817 gnd.n4194 gnd.n938 0.152939
R13818 gnd.n4196 gnd.n4194 0.152939
R13819 gnd.n4196 gnd.n4195 0.152939
R13820 gnd.n6641 gnd.n771 0.152939
R13821 gnd.n776 gnd.n771 0.152939
R13822 gnd.n777 gnd.n776 0.152939
R13823 gnd.n778 gnd.n777 0.152939
R13824 gnd.n779 gnd.n778 0.152939
R13825 gnd.n784 gnd.n779 0.152939
R13826 gnd.n785 gnd.n784 0.152939
R13827 gnd.n786 gnd.n785 0.152939
R13828 gnd.n787 gnd.n786 0.152939
R13829 gnd.n792 gnd.n787 0.152939
R13830 gnd.n793 gnd.n792 0.152939
R13831 gnd.n794 gnd.n793 0.152939
R13832 gnd.n795 gnd.n794 0.152939
R13833 gnd.n800 gnd.n795 0.152939
R13834 gnd.n801 gnd.n800 0.152939
R13835 gnd.n802 gnd.n801 0.152939
R13836 gnd.n803 gnd.n802 0.152939
R13837 gnd.n808 gnd.n803 0.152939
R13838 gnd.n809 gnd.n808 0.152939
R13839 gnd.n810 gnd.n809 0.152939
R13840 gnd.n811 gnd.n810 0.152939
R13841 gnd.n816 gnd.n811 0.152939
R13842 gnd.n817 gnd.n816 0.152939
R13843 gnd.n818 gnd.n817 0.152939
R13844 gnd.n819 gnd.n818 0.152939
R13845 gnd.n824 gnd.n819 0.152939
R13846 gnd.n825 gnd.n824 0.152939
R13847 gnd.n826 gnd.n825 0.152939
R13848 gnd.n827 gnd.n826 0.152939
R13849 gnd.n832 gnd.n827 0.152939
R13850 gnd.n833 gnd.n832 0.152939
R13851 gnd.n834 gnd.n833 0.152939
R13852 gnd.n835 gnd.n834 0.152939
R13853 gnd.n840 gnd.n835 0.152939
R13854 gnd.n841 gnd.n840 0.152939
R13855 gnd.n842 gnd.n841 0.152939
R13856 gnd.n843 gnd.n842 0.152939
R13857 gnd.n848 gnd.n843 0.152939
R13858 gnd.n849 gnd.n848 0.152939
R13859 gnd.n850 gnd.n849 0.152939
R13860 gnd.n851 gnd.n850 0.152939
R13861 gnd.n856 gnd.n851 0.152939
R13862 gnd.n857 gnd.n856 0.152939
R13863 gnd.n858 gnd.n857 0.152939
R13864 gnd.n859 gnd.n858 0.152939
R13865 gnd.n864 gnd.n859 0.152939
R13866 gnd.n865 gnd.n864 0.152939
R13867 gnd.n866 gnd.n865 0.152939
R13868 gnd.n867 gnd.n866 0.152939
R13869 gnd.n872 gnd.n867 0.152939
R13870 gnd.n873 gnd.n872 0.152939
R13871 gnd.n874 gnd.n873 0.152939
R13872 gnd.n875 gnd.n874 0.152939
R13873 gnd.n880 gnd.n875 0.152939
R13874 gnd.n881 gnd.n880 0.152939
R13875 gnd.n882 gnd.n881 0.152939
R13876 gnd.n883 gnd.n882 0.152939
R13877 gnd.n888 gnd.n883 0.152939
R13878 gnd.n889 gnd.n888 0.152939
R13879 gnd.n890 gnd.n889 0.152939
R13880 gnd.n891 gnd.n890 0.152939
R13881 gnd.n896 gnd.n891 0.152939
R13882 gnd.n897 gnd.n896 0.152939
R13883 gnd.n898 gnd.n897 0.152939
R13884 gnd.n899 gnd.n898 0.152939
R13885 gnd.n904 gnd.n899 0.152939
R13886 gnd.n905 gnd.n904 0.152939
R13887 gnd.n906 gnd.n905 0.152939
R13888 gnd.n907 gnd.n906 0.152939
R13889 gnd.n912 gnd.n907 0.152939
R13890 gnd.n913 gnd.n912 0.152939
R13891 gnd.n914 gnd.n913 0.152939
R13892 gnd.n915 gnd.n914 0.152939
R13893 gnd.n920 gnd.n915 0.152939
R13894 gnd.n921 gnd.n920 0.152939
R13895 gnd.n922 gnd.n921 0.152939
R13896 gnd.n923 gnd.n922 0.152939
R13897 gnd.n928 gnd.n923 0.152939
R13898 gnd.n929 gnd.n928 0.152939
R13899 gnd.n930 gnd.n929 0.152939
R13900 gnd.n931 gnd.n930 0.152939
R13901 gnd.n936 gnd.n931 0.152939
R13902 gnd.n937 gnd.n936 0.152939
R13903 gnd.n6471 gnd.n937 0.152939
R13904 gnd.n4673 gnd.n4672 0.152939
R13905 gnd.n4672 gnd.n2047 0.152939
R13906 gnd.n4700 gnd.n2047 0.152939
R13907 gnd.n4701 gnd.n4700 0.152939
R13908 gnd.n4705 gnd.n4701 0.152939
R13909 gnd.n4705 gnd.n4704 0.152939
R13910 gnd.n4704 gnd.n4703 0.152939
R13911 gnd.n4703 gnd.n1946 0.152939
R13912 gnd.n4737 gnd.n1946 0.152939
R13913 gnd.n4738 gnd.n4737 0.152939
R13914 gnd.n4740 gnd.n4738 0.152939
R13915 gnd.n4740 gnd.n4739 0.152939
R13916 gnd.n4739 gnd.n1935 0.152939
R13917 gnd.n4762 gnd.n1935 0.152939
R13918 gnd.n4763 gnd.n4762 0.152939
R13919 gnd.n4771 gnd.n4763 0.152939
R13920 gnd.n4771 gnd.n4770 0.152939
R13921 gnd.n4770 gnd.n4769 0.152939
R13922 gnd.n4769 gnd.n4764 0.152939
R13923 gnd.n4764 gnd.n1888 0.152939
R13924 gnd.n4848 gnd.n1888 0.152939
R13925 gnd.n4849 gnd.n4848 0.152939
R13926 gnd.n4869 gnd.n4849 0.152939
R13927 gnd.n4869 gnd.n4868 0.152939
R13928 gnd.n4868 gnd.n4867 0.152939
R13929 gnd.n4867 gnd.n4850 0.152939
R13930 gnd.n4863 gnd.n4850 0.152939
R13931 gnd.n4863 gnd.n4862 0.152939
R13932 gnd.n4862 gnd.n4861 0.152939
R13933 gnd.n4861 gnd.n4858 0.152939
R13934 gnd.n4858 gnd.n4857 0.152939
R13935 gnd.n4857 gnd.n1836 0.152939
R13936 gnd.n4950 gnd.n1836 0.152939
R13937 gnd.n4951 gnd.n4950 0.152939
R13938 gnd.n4952 gnd.n4951 0.152939
R13939 gnd.n4952 gnd.n1812 0.152939
R13940 gnd.n4998 gnd.n1812 0.152939
R13941 gnd.n4998 gnd.n4997 0.152939
R13942 gnd.n4997 gnd.n4996 0.152939
R13943 gnd.n4996 gnd.n1789 0.152939
R13944 gnd.n5057 gnd.n1789 0.152939
R13945 gnd.n5057 gnd.n5056 0.152939
R13946 gnd.n5056 gnd.n5055 0.152939
R13947 gnd.n5055 gnd.n1790 0.152939
R13948 gnd.n5051 gnd.n1790 0.152939
R13949 gnd.n5051 gnd.n5050 0.152939
R13950 gnd.n5050 gnd.n5049 0.152939
R13951 gnd.n5049 gnd.n5039 0.152939
R13952 gnd.n5045 gnd.n5039 0.152939
R13953 gnd.n5045 gnd.n1727 0.152939
R13954 gnd.n5167 gnd.n1727 0.152939
R13955 gnd.n5168 gnd.n5167 0.152939
R13956 gnd.n5170 gnd.n5168 0.152939
R13957 gnd.n5170 gnd.n5169 0.152939
R13958 gnd.n5169 gnd.n1698 0.152939
R13959 gnd.n5206 gnd.n1698 0.152939
R13960 gnd.n5207 gnd.n5206 0.152939
R13961 gnd.n5223 gnd.n5207 0.152939
R13962 gnd.n5223 gnd.n5222 0.152939
R13963 gnd.n5222 gnd.n5221 0.152939
R13964 gnd.n5221 gnd.n5208 0.152939
R13965 gnd.n5217 gnd.n5208 0.152939
R13966 gnd.n5217 gnd.n5216 0.152939
R13967 gnd.n5216 gnd.n5215 0.152939
R13968 gnd.n5215 gnd.n1642 0.152939
R13969 gnd.n5297 gnd.n1642 0.152939
R13970 gnd.n5298 gnd.n5297 0.152939
R13971 gnd.n5300 gnd.n5298 0.152939
R13972 gnd.n5300 gnd.n5299 0.152939
R13973 gnd.n5299 gnd.n1615 0.152939
R13974 gnd.n5339 gnd.n1615 0.152939
R13975 gnd.n5340 gnd.n5339 0.152939
R13976 gnd.n5341 gnd.n5340 0.152939
R13977 gnd.n5341 gnd.n1612 0.152939
R13978 gnd.n5350 gnd.n1612 0.152939
R13979 gnd.n5351 gnd.n5350 0.152939
R13980 gnd.n5352 gnd.n5351 0.152939
R13981 gnd.n5352 gnd.n1610 0.152939
R13982 gnd.n5358 gnd.n1610 0.152939
R13983 gnd.n5359 gnd.n5358 0.152939
R13984 gnd.n5538 gnd.n5359 0.152939
R13985 gnd.n5538 gnd.n5537 0.152939
R13986 gnd.n4233 gnd.n4232 0.152939
R13987 gnd.n4233 gnd.n2136 0.152939
R13988 gnd.n4274 gnd.n2136 0.152939
R13989 gnd.n4274 gnd.n4273 0.152939
R13990 gnd.n4273 gnd.n4272 0.152939
R13991 gnd.n4272 gnd.n2137 0.152939
R13992 gnd.n4268 gnd.n2137 0.152939
R13993 gnd.n4268 gnd.n4267 0.152939
R13994 gnd.n4267 gnd.n4266 0.152939
R13995 gnd.n4266 gnd.n2117 0.152939
R13996 gnd.n4319 gnd.n2117 0.152939
R13997 gnd.n4320 gnd.n4319 0.152939
R13998 gnd.n4321 gnd.n4320 0.152939
R13999 gnd.n4321 gnd.n2112 0.152939
R14000 gnd.n4334 gnd.n2112 0.152939
R14001 gnd.n4335 gnd.n4334 0.152939
R14002 gnd.n4336 gnd.n4335 0.152939
R14003 gnd.n4336 gnd.n2104 0.152939
R14004 gnd.n4370 gnd.n2104 0.152939
R14005 gnd.n4370 gnd.n4369 0.152939
R14006 gnd.n4369 gnd.n4368 0.152939
R14007 gnd.n4368 gnd.n2105 0.152939
R14008 gnd.n4364 gnd.n2105 0.152939
R14009 gnd.n4364 gnd.n4363 0.152939
R14010 gnd.n4363 gnd.n4362 0.152939
R14011 gnd.n4362 gnd.n2109 0.152939
R14012 gnd.n4650 gnd.n4416 0.152939
R14013 gnd.n4650 gnd.n4649 0.152939
R14014 gnd.n4649 gnd.n4648 0.152939
R14015 gnd.n4648 gnd.n4418 0.152939
R14016 gnd.n4644 gnd.n4418 0.152939
R14017 gnd.n4644 gnd.n4643 0.152939
R14018 gnd.n4691 gnd.n2056 0.152939
R14019 gnd.n4692 gnd.n4691 0.152939
R14020 gnd.n4694 gnd.n4692 0.152939
R14021 gnd.n4694 gnd.n4693 0.152939
R14022 gnd.n4693 gnd.n2032 0.152939
R14023 gnd.n4724 gnd.n2032 0.152939
R14024 gnd.n4725 gnd.n4724 0.152939
R14025 gnd.n4730 gnd.n4725 0.152939
R14026 gnd.n4730 gnd.n4729 0.152939
R14027 gnd.n4729 gnd.n4728 0.152939
R14028 gnd.n4728 gnd.n1228 0.152939
R14029 gnd.n6245 gnd.n1228 0.152939
R14030 gnd.n6245 gnd.n6244 0.152939
R14031 gnd.n6244 gnd.n6243 0.152939
R14032 gnd.n6243 gnd.n1229 0.152939
R14033 gnd.n6239 gnd.n1229 0.152939
R14034 gnd.n6239 gnd.n6238 0.152939
R14035 gnd.n6238 gnd.n6237 0.152939
R14036 gnd.n6237 gnd.n1234 0.152939
R14037 gnd.n6233 gnd.n1234 0.152939
R14038 gnd.n6233 gnd.n6232 0.152939
R14039 gnd.n6232 gnd.n6231 0.152939
R14040 gnd.n6231 gnd.n1239 0.152939
R14041 gnd.n6227 gnd.n1239 0.152939
R14042 gnd.n6227 gnd.n6226 0.152939
R14043 gnd.n6226 gnd.n6225 0.152939
R14044 gnd.n6225 gnd.n1244 0.152939
R14045 gnd.n6221 gnd.n1244 0.152939
R14046 gnd.n6221 gnd.n6220 0.152939
R14047 gnd.n6220 gnd.n6219 0.152939
R14048 gnd.n6219 gnd.n1249 0.152939
R14049 gnd.n6215 gnd.n1249 0.152939
R14050 gnd.n6215 gnd.n6214 0.152939
R14051 gnd.n6214 gnd.n6213 0.152939
R14052 gnd.n6213 gnd.n1254 0.152939
R14053 gnd.n6209 gnd.n1254 0.152939
R14054 gnd.n6209 gnd.n6208 0.152939
R14055 gnd.n6208 gnd.n6207 0.152939
R14056 gnd.n6207 gnd.n1259 0.152939
R14057 gnd.n6203 gnd.n1259 0.152939
R14058 gnd.n6203 gnd.n6202 0.152939
R14059 gnd.n6202 gnd.n6201 0.152939
R14060 gnd.n6201 gnd.n1264 0.152939
R14061 gnd.n6197 gnd.n1264 0.152939
R14062 gnd.n6197 gnd.n6196 0.152939
R14063 gnd.n6196 gnd.n6195 0.152939
R14064 gnd.n6195 gnd.n1269 0.152939
R14065 gnd.n6191 gnd.n1269 0.152939
R14066 gnd.n6191 gnd.n6190 0.152939
R14067 gnd.n6190 gnd.n6189 0.152939
R14068 gnd.n6189 gnd.n1274 0.152939
R14069 gnd.n6185 gnd.n1274 0.152939
R14070 gnd.n6185 gnd.n6184 0.152939
R14071 gnd.n6184 gnd.n6183 0.152939
R14072 gnd.n6183 gnd.n1279 0.152939
R14073 gnd.n6179 gnd.n1279 0.152939
R14074 gnd.n6179 gnd.n6178 0.152939
R14075 gnd.n6178 gnd.n6177 0.152939
R14076 gnd.n6177 gnd.n1284 0.152939
R14077 gnd.n6173 gnd.n1284 0.152939
R14078 gnd.n6173 gnd.n6172 0.152939
R14079 gnd.n6172 gnd.n6171 0.152939
R14080 gnd.n6171 gnd.n1289 0.152939
R14081 gnd.n6167 gnd.n1289 0.152939
R14082 gnd.n6167 gnd.n6166 0.152939
R14083 gnd.n6166 gnd.n6165 0.152939
R14084 gnd.n6165 gnd.n1294 0.152939
R14085 gnd.n6161 gnd.n1294 0.152939
R14086 gnd.n6161 gnd.n6160 0.152939
R14087 gnd.n6160 gnd.n6159 0.152939
R14088 gnd.n6159 gnd.n1299 0.152939
R14089 gnd.n6155 gnd.n1299 0.152939
R14090 gnd.n6155 gnd.n6154 0.152939
R14091 gnd.n6154 gnd.n6153 0.152939
R14092 gnd.n6153 gnd.n1304 0.152939
R14093 gnd.n6149 gnd.n1304 0.152939
R14094 gnd.n6149 gnd.n6148 0.152939
R14095 gnd.n6148 gnd.n6147 0.152939
R14096 gnd.n6147 gnd.n1309 0.152939
R14097 gnd.n6143 gnd.n1309 0.152939
R14098 gnd.n6143 gnd.n6142 0.152939
R14099 gnd.n6142 gnd.n6141 0.152939
R14100 gnd.n5424 gnd.n1314 0.152939
R14101 gnd.n5424 gnd.n5420 0.152939
R14102 gnd.n5432 gnd.n5420 0.152939
R14103 gnd.n5433 gnd.n5432 0.152939
R14104 gnd.n5435 gnd.n5433 0.152939
R14105 gnd.n5435 gnd.n5434 0.152939
R14106 gnd.n5365 gnd.n5360 0.152939
R14107 gnd.n5360 gnd.n1494 0.152939
R14108 gnd.n5912 gnd.n1494 0.152939
R14109 gnd.n5913 gnd.n5912 0.152939
R14110 gnd.n5914 gnd.n5913 0.152939
R14111 gnd.n5914 gnd.n1490 0.152939
R14112 gnd.n5933 gnd.n1490 0.152939
R14113 gnd.n5933 gnd.n5932 0.152939
R14114 gnd.n5932 gnd.n5931 0.152939
R14115 gnd.n5931 gnd.n1479 0.152939
R14116 gnd.n5993 gnd.n1479 0.152939
R14117 gnd.n5994 gnd.n5993 0.152939
R14118 gnd.n5995 gnd.n5994 0.152939
R14119 gnd.n5995 gnd.n1473 0.152939
R14120 gnd.n6007 gnd.n1473 0.152939
R14121 gnd.n6008 gnd.n6007 0.152939
R14122 gnd.n6009 gnd.n6008 0.152939
R14123 gnd.n6009 gnd.n1468 0.152939
R14124 gnd.n6034 gnd.n1468 0.152939
R14125 gnd.n6034 gnd.n6033 0.152939
R14126 gnd.n6033 gnd.n6032 0.152939
R14127 gnd.n6032 gnd.n1469 0.152939
R14128 gnd.n6028 gnd.n1469 0.152939
R14129 gnd.n6028 gnd.n6027 0.152939
R14130 gnd.n6027 gnd.n6026 0.152939
R14131 gnd.n6026 gnd.n79 0.152939
R14132 gnd.n4643 gnd.n4642 0.128549
R14133 gnd.n5434 gnd.n1498 0.128549
R14134 gnd.n4283 gnd.n973 0.10111
R14135 gnd.n5974 gnd.n95 0.10111
R14136 gnd.n3147 gnd.n3146 0.0767195
R14137 gnd.n3146 gnd.n3145 0.0767195
R14138 gnd.n7633 gnd.n93 0.0767195
R14139 gnd.n7633 gnd.n94 0.0767195
R14140 gnd.n6450 gnd.n971 0.0767195
R14141 gnd.n6450 gnd.n972 0.0767195
R14142 gnd.n7643 gnd.n7642 0.0695946
R14143 gnd.n4231 gnd.n4230 0.0695946
R14144 gnd.n4232 gnd.n4231 0.0695946
R14145 gnd.n7643 gnd.n79 0.0695946
R14146 gnd.n4642 gnd.n4535 0.063
R14147 gnd.n5901 gnd.n1498 0.063
R14148 gnd.n388 gnd.n95 0.0523293
R14149 gnd.n4195 gnd.n973 0.0523293
R14150 gnd.n3713 gnd.n2313 0.0477147
R14151 gnd.n5903 gnd.n5901 0.0477147
R14152 gnd.n7451 gnd.n205 0.0477147
R14153 gnd.n3925 gnd.n2266 0.0477147
R14154 gnd.n4535 gnd.n1090 0.0477147
R14155 gnd.n2910 gnd.n2798 0.0442063
R14156 gnd.n2911 gnd.n2910 0.0442063
R14157 gnd.n2912 gnd.n2911 0.0442063
R14158 gnd.n2912 gnd.n2787 0.0442063
R14159 gnd.n2926 gnd.n2787 0.0442063
R14160 gnd.n2927 gnd.n2926 0.0442063
R14161 gnd.n2928 gnd.n2927 0.0442063
R14162 gnd.n2928 gnd.n2774 0.0442063
R14163 gnd.n2972 gnd.n2774 0.0442063
R14164 gnd.n2973 gnd.n2972 0.0442063
R14165 gnd.n2975 gnd.n2708 0.0344674
R14166 gnd.n5904 gnd.n5903 0.0344674
R14167 gnd.n5904 gnd.n1356 0.0344674
R14168 gnd.n1357 gnd.n1356 0.0344674
R14169 gnd.n1358 gnd.n1357 0.0344674
R14170 gnd.n1492 gnd.n1358 0.0344674
R14171 gnd.n1492 gnd.n1376 0.0344674
R14172 gnd.n1377 gnd.n1376 0.0344674
R14173 gnd.n1378 gnd.n1377 0.0344674
R14174 gnd.n5923 gnd.n1378 0.0344674
R14175 gnd.n5923 gnd.n1397 0.0344674
R14176 gnd.n1398 gnd.n1397 0.0344674
R14177 gnd.n1399 gnd.n1398 0.0344674
R14178 gnd.n1477 gnd.n1399 0.0344674
R14179 gnd.n1477 gnd.n1416 0.0344674
R14180 gnd.n1417 gnd.n1416 0.0344674
R14181 gnd.n1418 gnd.n1417 0.0344674
R14182 gnd.n1471 gnd.n1418 0.0344674
R14183 gnd.n1471 gnd.n1437 0.0344674
R14184 gnd.n1438 gnd.n1437 0.0344674
R14185 gnd.n1439 gnd.n1438 0.0344674
R14186 gnd.n6018 gnd.n1439 0.0344674
R14187 gnd.n6018 gnd.n1454 0.0344674
R14188 gnd.n6052 gnd.n1454 0.0344674
R14189 gnd.n6052 gnd.n372 0.0344674
R14190 gnd.n7307 gnd.n372 0.0344674
R14191 gnd.n7308 gnd.n7307 0.0344674
R14192 gnd.n7308 gnd.n367 0.0344674
R14193 gnd.n367 gnd.n365 0.0344674
R14194 gnd.n7320 gnd.n365 0.0344674
R14195 gnd.n7321 gnd.n7320 0.0344674
R14196 gnd.n7321 gnd.n109 0.0344674
R14197 gnd.n110 gnd.n109 0.0344674
R14198 gnd.n111 gnd.n110 0.0344674
R14199 gnd.n7337 gnd.n111 0.0344674
R14200 gnd.n7337 gnd.n127 0.0344674
R14201 gnd.n128 gnd.n127 0.0344674
R14202 gnd.n129 gnd.n128 0.0344674
R14203 gnd.n353 gnd.n129 0.0344674
R14204 gnd.n353 gnd.n147 0.0344674
R14205 gnd.n148 gnd.n147 0.0344674
R14206 gnd.n149 gnd.n148 0.0344674
R14207 gnd.n7392 gnd.n149 0.0344674
R14208 gnd.n7392 gnd.n165 0.0344674
R14209 gnd.n166 gnd.n165 0.0344674
R14210 gnd.n167 gnd.n166 0.0344674
R14211 gnd.n7399 gnd.n167 0.0344674
R14212 gnd.n7399 gnd.n185 0.0344674
R14213 gnd.n186 gnd.n185 0.0344674
R14214 gnd.n187 gnd.n186 0.0344674
R14215 gnd.n7406 gnd.n187 0.0344674
R14216 gnd.n7406 gnd.n203 0.0344674
R14217 gnd.n204 gnd.n203 0.0344674
R14218 gnd.n205 gnd.n204 0.0344674
R14219 gnd.n4050 gnd.n2266 0.0344674
R14220 gnd.n4050 gnd.n2269 0.0344674
R14221 gnd.n2269 gnd.n2268 0.0344674
R14222 gnd.n2268 gnd.n2249 0.0344674
R14223 gnd.n2249 gnd.n2246 0.0344674
R14224 gnd.n2247 gnd.n2246 0.0344674
R14225 gnd.n4069 gnd.n2247 0.0344674
R14226 gnd.n4070 gnd.n4069 0.0344674
R14227 gnd.n4070 gnd.n2223 0.0344674
R14228 gnd.n2223 gnd.n2219 0.0344674
R14229 gnd.n2220 gnd.n2219 0.0344674
R14230 gnd.n4108 gnd.n2220 0.0344674
R14231 gnd.n4108 gnd.n2221 0.0344674
R14232 gnd.n2221 gnd.n2196 0.0344674
R14233 gnd.n4139 gnd.n2196 0.0344674
R14234 gnd.n4139 gnd.n2197 0.0344674
R14235 gnd.n2197 gnd.n2180 0.0344674
R14236 gnd.n4157 gnd.n2180 0.0344674
R14237 gnd.n4158 gnd.n4157 0.0344674
R14238 gnd.n4158 gnd.n960 0.0344674
R14239 gnd.n961 gnd.n960 0.0344674
R14240 gnd.n962 gnd.n961 0.0344674
R14241 gnd.n4161 gnd.n962 0.0344674
R14242 gnd.n4162 gnd.n4161 0.0344674
R14243 gnd.n4162 gnd.n2164 0.0344674
R14244 gnd.n2165 gnd.n2164 0.0344674
R14245 gnd.n2166 gnd.n2165 0.0344674
R14246 gnd.n2166 gnd.n2142 0.0344674
R14247 gnd.n4244 gnd.n2142 0.0344674
R14248 gnd.n4245 gnd.n4244 0.0344674
R14249 gnd.n4245 gnd.n988 0.0344674
R14250 gnd.n989 gnd.n988 0.0344674
R14251 gnd.n990 gnd.n989 0.0344674
R14252 gnd.n4252 gnd.n990 0.0344674
R14253 gnd.n4252 gnd.n1007 0.0344674
R14254 gnd.n1008 gnd.n1007 0.0344674
R14255 gnd.n1009 gnd.n1008 0.0344674
R14256 gnd.n4258 gnd.n1009 0.0344674
R14257 gnd.n4258 gnd.n1027 0.0344674
R14258 gnd.n1028 gnd.n1027 0.0344674
R14259 gnd.n1029 gnd.n1028 0.0344674
R14260 gnd.n4328 gnd.n1029 0.0344674
R14261 gnd.n4328 gnd.n1047 0.0344674
R14262 gnd.n1048 gnd.n1047 0.0344674
R14263 gnd.n1049 gnd.n1048 0.0344674
R14264 gnd.n4343 gnd.n1049 0.0344674
R14265 gnd.n4343 gnd.n1067 0.0344674
R14266 gnd.n1068 gnd.n1067 0.0344674
R14267 gnd.n1069 gnd.n1068 0.0344674
R14268 gnd.n4350 gnd.n1069 0.0344674
R14269 gnd.n4350 gnd.n1088 0.0344674
R14270 gnd.n1089 gnd.n1088 0.0344674
R14271 gnd.n1090 gnd.n1089 0.0344674
R14272 gnd.n4641 gnd.n4536 0.0344674
R14273 gnd.n5444 gnd.n5443 0.0344674
R14274 gnd.n4668 gnd.n2071 0.029712
R14275 gnd.n5375 gnd.n5366 0.029712
R14276 gnd.n2995 gnd.n2994 0.0269946
R14277 gnd.n2997 gnd.n2996 0.0269946
R14278 gnd.n2703 gnd.n2701 0.0269946
R14279 gnd.n3007 gnd.n3005 0.0269946
R14280 gnd.n3006 gnd.n2682 0.0269946
R14281 gnd.n3026 gnd.n3025 0.0269946
R14282 gnd.n3028 gnd.n3027 0.0269946
R14283 gnd.n2677 gnd.n2676 0.0269946
R14284 gnd.n3038 gnd.n2672 0.0269946
R14285 gnd.n3037 gnd.n2674 0.0269946
R14286 gnd.n2673 gnd.n2655 0.0269946
R14287 gnd.n3058 gnd.n2656 0.0269946
R14288 gnd.n3057 gnd.n2657 0.0269946
R14289 gnd.n3091 gnd.n2632 0.0269946
R14290 gnd.n3093 gnd.n3092 0.0269946
R14291 gnd.n3094 gnd.n2579 0.0269946
R14292 gnd.n2627 gnd.n2580 0.0269946
R14293 gnd.n2629 gnd.n2581 0.0269946
R14294 gnd.n3104 gnd.n3103 0.0269946
R14295 gnd.n3106 gnd.n3105 0.0269946
R14296 gnd.n3107 gnd.n2601 0.0269946
R14297 gnd.n3109 gnd.n2602 0.0269946
R14298 gnd.n3112 gnd.n2603 0.0269946
R14299 gnd.n3115 gnd.n3114 0.0269946
R14300 gnd.n3117 gnd.n3116 0.0269946
R14301 gnd.n3182 gnd.n2486 0.0269946
R14302 gnd.n3184 gnd.n3183 0.0269946
R14303 gnd.n3193 gnd.n2479 0.0269946
R14304 gnd.n3195 gnd.n3194 0.0269946
R14305 gnd.n3196 gnd.n2477 0.0269946
R14306 gnd.n3203 gnd.n3199 0.0269946
R14307 gnd.n3202 gnd.n3201 0.0269946
R14308 gnd.n3200 gnd.n2456 0.0269946
R14309 gnd.n3225 gnd.n2457 0.0269946
R14310 gnd.n3224 gnd.n2458 0.0269946
R14311 gnd.n3267 gnd.n2431 0.0269946
R14312 gnd.n3269 gnd.n3268 0.0269946
R14313 gnd.n3278 gnd.n2424 0.0269946
R14314 gnd.n3280 gnd.n3279 0.0269946
R14315 gnd.n3281 gnd.n2422 0.0269946
R14316 gnd.n3288 gnd.n3284 0.0269946
R14317 gnd.n3287 gnd.n3286 0.0269946
R14318 gnd.n3285 gnd.n2401 0.0269946
R14319 gnd.n3310 gnd.n2402 0.0269946
R14320 gnd.n3309 gnd.n2403 0.0269946
R14321 gnd.n3356 gnd.n2377 0.0269946
R14322 gnd.n3358 gnd.n3357 0.0269946
R14323 gnd.n3367 gnd.n2370 0.0269946
R14324 gnd.n3626 gnd.n2368 0.0269946
R14325 gnd.n3631 gnd.n3629 0.0269946
R14326 gnd.n3630 gnd.n2349 0.0269946
R14327 gnd.n3655 gnd.n3654 0.0269946
R14328 gnd.n4637 gnd.n4542 0.0225788
R14329 gnd.n4636 gnd.n4543 0.0225788
R14330 gnd.n4633 gnd.n4632 0.0225788
R14331 gnd.n4629 gnd.n4549 0.0225788
R14332 gnd.n4628 gnd.n4555 0.0225788
R14333 gnd.n4625 gnd.n4624 0.0225788
R14334 gnd.n4621 gnd.n4561 0.0225788
R14335 gnd.n4620 gnd.n4565 0.0225788
R14336 gnd.n4617 gnd.n4616 0.0225788
R14337 gnd.n4613 gnd.n4572 0.0225788
R14338 gnd.n4612 gnd.n4578 0.0225788
R14339 gnd.n4609 gnd.n4608 0.0225788
R14340 gnd.n4605 gnd.n4584 0.0225788
R14341 gnd.n4604 gnd.n4588 0.0225788
R14342 gnd.n4601 gnd.n4600 0.0225788
R14343 gnd.n4595 gnd.n2080 0.0225788
R14344 gnd.n4660 gnd.n4659 0.0225788
R14345 gnd.n2081 gnd.n2074 0.0225788
R14346 gnd.n4668 gnd.n4667 0.0225788
R14347 gnd.n5450 gnd.n5448 0.0225788
R14348 gnd.n5449 gnd.n5412 0.0225788
R14349 gnd.n5459 gnd.n5458 0.0225788
R14350 gnd.n5413 gnd.n5408 0.0225788
R14351 gnd.n5469 gnd.n5467 0.0225788
R14352 gnd.n5468 gnd.n5403 0.0225788
R14353 gnd.n5478 gnd.n5477 0.0225788
R14354 gnd.n5404 gnd.n5399 0.0225788
R14355 gnd.n5488 gnd.n5486 0.0225788
R14356 gnd.n5487 gnd.n5394 0.0225788
R14357 gnd.n5497 gnd.n5496 0.0225788
R14358 gnd.n5395 gnd.n5390 0.0225788
R14359 gnd.n5507 gnd.n5505 0.0225788
R14360 gnd.n5506 gnd.n5385 0.0225788
R14361 gnd.n5517 gnd.n5516 0.0225788
R14362 gnd.n5513 gnd.n5386 0.0225788
R14363 gnd.n5527 gnd.n5373 0.0225788
R14364 gnd.n5526 gnd.n5374 0.0225788
R14365 gnd.n5376 gnd.n5375 0.0225788
R14366 gnd.n5536 gnd.n5366 0.0218415
R14367 gnd.n4671 gnd.n2071 0.0218415
R14368 gnd.n2975 gnd.n2974 0.0202011
R14369 gnd.n2974 gnd.n2973 0.0148637
R14370 gnd.n3624 gnd.n3368 0.0144266
R14371 gnd.n3625 gnd.n3624 0.0130679
R14372 gnd.n4542 gnd.n4536 0.0123886
R14373 gnd.n4637 gnd.n4636 0.0123886
R14374 gnd.n4633 gnd.n4543 0.0123886
R14375 gnd.n4632 gnd.n4549 0.0123886
R14376 gnd.n4629 gnd.n4628 0.0123886
R14377 gnd.n4625 gnd.n4555 0.0123886
R14378 gnd.n4624 gnd.n4561 0.0123886
R14379 gnd.n4621 gnd.n4620 0.0123886
R14380 gnd.n4617 gnd.n4565 0.0123886
R14381 gnd.n4616 gnd.n4572 0.0123886
R14382 gnd.n4613 gnd.n4612 0.0123886
R14383 gnd.n4609 gnd.n4578 0.0123886
R14384 gnd.n4608 gnd.n4584 0.0123886
R14385 gnd.n4605 gnd.n4604 0.0123886
R14386 gnd.n4601 gnd.n4588 0.0123886
R14387 gnd.n4600 gnd.n4595 0.0123886
R14388 gnd.n4660 gnd.n2080 0.0123886
R14389 gnd.n4659 gnd.n2081 0.0123886
R14390 gnd.n4667 gnd.n2074 0.0123886
R14391 gnd.n5448 gnd.n5444 0.0123886
R14392 gnd.n5450 gnd.n5449 0.0123886
R14393 gnd.n5459 gnd.n5412 0.0123886
R14394 gnd.n5458 gnd.n5413 0.0123886
R14395 gnd.n5467 gnd.n5408 0.0123886
R14396 gnd.n5469 gnd.n5468 0.0123886
R14397 gnd.n5478 gnd.n5403 0.0123886
R14398 gnd.n5477 gnd.n5404 0.0123886
R14399 gnd.n5486 gnd.n5399 0.0123886
R14400 gnd.n5488 gnd.n5487 0.0123886
R14401 gnd.n5497 gnd.n5394 0.0123886
R14402 gnd.n5496 gnd.n5395 0.0123886
R14403 gnd.n5505 gnd.n5390 0.0123886
R14404 gnd.n5507 gnd.n5506 0.0123886
R14405 gnd.n5517 gnd.n5385 0.0123886
R14406 gnd.n5516 gnd.n5386 0.0123886
R14407 gnd.n5513 gnd.n5373 0.0123886
R14408 gnd.n5527 gnd.n5526 0.0123886
R14409 gnd.n5376 gnd.n5374 0.0123886
R14410 gnd.n2994 gnd.n2708 0.00797283
R14411 gnd.n2996 gnd.n2995 0.00797283
R14412 gnd.n2997 gnd.n2703 0.00797283
R14413 gnd.n3005 gnd.n2701 0.00797283
R14414 gnd.n3007 gnd.n3006 0.00797283
R14415 gnd.n3025 gnd.n2682 0.00797283
R14416 gnd.n3027 gnd.n3026 0.00797283
R14417 gnd.n3028 gnd.n2677 0.00797283
R14418 gnd.n2676 gnd.n2672 0.00797283
R14419 gnd.n3038 gnd.n3037 0.00797283
R14420 gnd.n2674 gnd.n2673 0.00797283
R14421 gnd.n2656 gnd.n2655 0.00797283
R14422 gnd.n3058 gnd.n3057 0.00797283
R14423 gnd.n2657 gnd.n2632 0.00797283
R14424 gnd.n3092 gnd.n3091 0.00797283
R14425 gnd.n3094 gnd.n3093 0.00797283
R14426 gnd.n2627 gnd.n2579 0.00797283
R14427 gnd.n2629 gnd.n2580 0.00797283
R14428 gnd.n3103 gnd.n2581 0.00797283
R14429 gnd.n3105 gnd.n3104 0.00797283
R14430 gnd.n3107 gnd.n3106 0.00797283
R14431 gnd.n3109 gnd.n2601 0.00797283
R14432 gnd.n3112 gnd.n2602 0.00797283
R14433 gnd.n3114 gnd.n2603 0.00797283
R14434 gnd.n3117 gnd.n3115 0.00797283
R14435 gnd.n3116 gnd.n2486 0.00797283
R14436 gnd.n3184 gnd.n3182 0.00797283
R14437 gnd.n3183 gnd.n2479 0.00797283
R14438 gnd.n3194 gnd.n3193 0.00797283
R14439 gnd.n3196 gnd.n3195 0.00797283
R14440 gnd.n3199 gnd.n2477 0.00797283
R14441 gnd.n3203 gnd.n3202 0.00797283
R14442 gnd.n3201 gnd.n3200 0.00797283
R14443 gnd.n2457 gnd.n2456 0.00797283
R14444 gnd.n3225 gnd.n3224 0.00797283
R14445 gnd.n2458 gnd.n2431 0.00797283
R14446 gnd.n3269 gnd.n3267 0.00797283
R14447 gnd.n3268 gnd.n2424 0.00797283
R14448 gnd.n3279 gnd.n3278 0.00797283
R14449 gnd.n3281 gnd.n3280 0.00797283
R14450 gnd.n3284 gnd.n2422 0.00797283
R14451 gnd.n3288 gnd.n3287 0.00797283
R14452 gnd.n3286 gnd.n3285 0.00797283
R14453 gnd.n2402 gnd.n2401 0.00797283
R14454 gnd.n3310 gnd.n3309 0.00797283
R14455 gnd.n2403 gnd.n2377 0.00797283
R14456 gnd.n3358 gnd.n3356 0.00797283
R14457 gnd.n3357 gnd.n2370 0.00797283
R14458 gnd.n3368 gnd.n3367 0.00797283
R14459 gnd.n3626 gnd.n3625 0.00797283
R14460 gnd.n3629 gnd.n2368 0.00797283
R14461 gnd.n3631 gnd.n3630 0.00797283
R14462 gnd.n3654 gnd.n2349 0.00797283
R14463 gnd.n3655 gnd.n2313 0.00797283
R14464 gnd.n4642 gnd.n4641 0.00593478
R14465 gnd.n5443 gnd.n1498 0.00593478
R14466 commonsourceibias.n35 commonsourceibias.t0 223.028
R14467 commonsourceibias.n128 commonsourceibias.t129 223.028
R14468 commonsourceibias.n307 commonsourceibias.t140 223.028
R14469 commonsourceibias.n217 commonsourceibias.t112 223.028
R14470 commonsourceibias.n454 commonsourceibias.t22 223.028
R14471 commonsourceibias.n395 commonsourceibias.t108 223.028
R14472 commonsourceibias.n679 commonsourceibias.t74 223.028
R14473 commonsourceibias.n589 commonsourceibias.t97 223.028
R14474 commonsourceibias.n99 commonsourceibias.t12 207.983
R14475 commonsourceibias.n192 commonsourceibias.t120 207.983
R14476 commonsourceibias.n371 commonsourceibias.t147 207.983
R14477 commonsourceibias.n281 commonsourceibias.t71 207.983
R14478 commonsourceibias.n520 commonsourceibias.t34 207.983
R14479 commonsourceibias.n566 commonsourceibias.t91 207.983
R14480 commonsourceibias.n745 commonsourceibias.t82 207.983
R14481 commonsourceibias.n655 commonsourceibias.t151 207.983
R14482 commonsourceibias.n97 commonsourceibias.t48 168.701
R14483 commonsourceibias.n91 commonsourceibias.t4 168.701
R14484 commonsourceibias.n17 commonsourceibias.t10 168.701
R14485 commonsourceibias.n83 commonsourceibias.t58 168.701
R14486 commonsourceibias.n77 commonsourceibias.t16 168.701
R14487 commonsourceibias.n22 commonsourceibias.t28 168.701
R14488 commonsourceibias.n69 commonsourceibias.t6 168.701
R14489 commonsourceibias.n63 commonsourceibias.t14 168.701
R14490 commonsourceibias.n25 commonsourceibias.t44 168.701
R14491 commonsourceibias.n27 commonsourceibias.t24 168.701
R14492 commonsourceibias.n29 commonsourceibias.t30 168.701
R14493 commonsourceibias.n46 commonsourceibias.t54 168.701
R14494 commonsourceibias.n40 commonsourceibias.t18 168.701
R14495 commonsourceibias.n34 commonsourceibias.t50 168.701
R14496 commonsourceibias.n190 commonsourceibias.t67 168.701
R14497 commonsourceibias.n184 commonsourceibias.t126 168.701
R14498 commonsourceibias.n5 commonsourceibias.t121 168.701
R14499 commonsourceibias.n176 commonsourceibias.t136 168.701
R14500 commonsourceibias.n170 commonsourceibias.t117 168.701
R14501 commonsourceibias.n10 commonsourceibias.t102 168.701
R14502 commonsourceibias.n162 commonsourceibias.t125 168.701
R14503 commonsourceibias.n156 commonsourceibias.t118 168.701
R14504 commonsourceibias.n118 commonsourceibias.t76 168.701
R14505 commonsourceibias.n120 commonsourceibias.t106 168.701
R14506 commonsourceibias.n122 commonsourceibias.t96 168.701
R14507 commonsourceibias.n139 commonsourceibias.t141 168.701
R14508 commonsourceibias.n133 commonsourceibias.t116 168.701
R14509 commonsourceibias.n127 commonsourceibias.t152 168.701
R14510 commonsourceibias.n306 commonsourceibias.t130 168.701
R14511 commonsourceibias.n312 commonsourceibias.t79 168.701
R14512 commonsourceibias.n318 commonsourceibias.t149 168.701
R14513 commonsourceibias.n301 commonsourceibias.t133 168.701
R14514 commonsourceibias.n299 commonsourceibias.t137 168.701
R14515 commonsourceibias.n297 commonsourceibias.t64 168.701
R14516 commonsourceibias.n335 commonsourceibias.t138 168.701
R14517 commonsourceibias.n341 commonsourceibias.t146 168.701
R14518 commonsourceibias.n294 commonsourceibias.t119 168.701
R14519 commonsourceibias.n349 commonsourceibias.t90 168.701
R14520 commonsourceibias.n355 commonsourceibias.t155 168.701
R14521 commonsourceibias.n289 commonsourceibias.t124 168.701
R14522 commonsourceibias.n363 commonsourceibias.t128 168.701
R14523 commonsourceibias.n369 commonsourceibias.t75 168.701
R14524 commonsourceibias.n279 commonsourceibias.t159 168.701
R14525 commonsourceibias.n273 commonsourceibias.t148 168.701
R14526 commonsourceibias.n199 commonsourceibias.t78 168.701
R14527 commonsourceibias.n265 commonsourceibias.t157 168.701
R14528 commonsourceibias.n259 commonsourceibias.t85 168.701
R14529 commonsourceibias.n204 commonsourceibias.t77 168.701
R14530 commonsourceibias.n251 commonsourceibias.t158 168.701
R14531 commonsourceibias.n245 commonsourceibias.t94 168.701
R14532 commonsourceibias.n207 commonsourceibias.t113 168.701
R14533 commonsourceibias.n209 commonsourceibias.t156 168.701
R14534 commonsourceibias.n211 commonsourceibias.t92 168.701
R14535 commonsourceibias.n228 commonsourceibias.t111 168.701
R14536 commonsourceibias.n222 commonsourceibias.t105 168.701
R14537 commonsourceibias.n216 commonsourceibias.t93 168.701
R14538 commonsourceibias.n453 commonsourceibias.t62 168.701
R14539 commonsourceibias.n459 commonsourceibias.t40 168.701
R14540 commonsourceibias.n465 commonsourceibias.t2 168.701
R14541 commonsourceibias.n448 commonsourceibias.t52 168.701
R14542 commonsourceibias.n446 commonsourceibias.t42 168.701
R14543 commonsourceibias.n444 commonsourceibias.t56 168.701
R14544 commonsourceibias.n482 commonsourceibias.t36 168.701
R14545 commonsourceibias.n488 commonsourceibias.t26 168.701
R14546 commonsourceibias.n490 commonsourceibias.t46 168.701
R14547 commonsourceibias.n497 commonsourceibias.t38 168.701
R14548 commonsourceibias.n503 commonsourceibias.t8 168.701
R14549 commonsourceibias.n505 commonsourceibias.t32 168.701
R14550 commonsourceibias.n512 commonsourceibias.t20 168.701
R14551 commonsourceibias.n518 commonsourceibias.t60 168.701
R14552 commonsourceibias.n564 commonsourceibias.t134 168.701
R14553 commonsourceibias.n558 commonsourceibias.t114 168.701
R14554 commonsourceibias.n551 commonsourceibias.t95 168.701
R14555 commonsourceibias.n549 commonsourceibias.t123 168.701
R14556 commonsourceibias.n543 commonsourceibias.t88 168.701
R14557 commonsourceibias.n536 commonsourceibias.t73 168.701
R14558 commonsourceibias.n534 commonsourceibias.t104 168.701
R14559 commonsourceibias.n394 commonsourceibias.t131 168.701
R14560 commonsourceibias.n400 commonsourceibias.t84 168.701
R14561 commonsourceibias.n406 commonsourceibias.t127 168.701
R14562 commonsourceibias.n389 commonsourceibias.t150 168.701
R14563 commonsourceibias.n387 commonsourceibias.t83 168.701
R14564 commonsourceibias.n385 commonsourceibias.t139 168.701
R14565 commonsourceibias.n423 commonsourceibias.t89 168.701
R14566 commonsourceibias.n678 commonsourceibias.t145 168.701
R14567 commonsourceibias.n684 commonsourceibias.t109 168.701
R14568 commonsourceibias.n690 commonsourceibias.t87 168.701
R14569 commonsourceibias.n673 commonsourceibias.t153 168.701
R14570 commonsourceibias.n671 commonsourceibias.t132 168.701
R14571 commonsourceibias.n669 commonsourceibias.t103 168.701
R14572 commonsourceibias.n707 commonsourceibias.t70 168.701
R14573 commonsourceibias.n713 commonsourceibias.t81 168.701
R14574 commonsourceibias.n715 commonsourceibias.t110 168.701
R14575 commonsourceibias.n722 commonsourceibias.t115 168.701
R14576 commonsourceibias.n728 commonsourceibias.t101 168.701
R14577 commonsourceibias.n730 commonsourceibias.t135 168.701
R14578 commonsourceibias.n737 commonsourceibias.t122 168.701
R14579 commonsourceibias.n743 commonsourceibias.t107 168.701
R14580 commonsourceibias.n588 commonsourceibias.t68 168.701
R14581 commonsourceibias.n594 commonsourceibias.t86 168.701
R14582 commonsourceibias.n600 commonsourceibias.t98 168.701
R14583 commonsourceibias.n583 commonsourceibias.t69 168.701
R14584 commonsourceibias.n581 commonsourceibias.t80 168.701
R14585 commonsourceibias.n579 commonsourceibias.t99 168.701
R14586 commonsourceibias.n617 commonsourceibias.t72 168.701
R14587 commonsourceibias.n623 commonsourceibias.t142 168.701
R14588 commonsourceibias.n625 commonsourceibias.t100 168.701
R14589 commonsourceibias.n632 commonsourceibias.t65 168.701
R14590 commonsourceibias.n638 commonsourceibias.t143 168.701
R14591 commonsourceibias.n640 commonsourceibias.t154 168.701
R14592 commonsourceibias.n647 commonsourceibias.t66 168.701
R14593 commonsourceibias.n653 commonsourceibias.t144 168.701
R14594 commonsourceibias.n36 commonsourceibias.n33 161.3
R14595 commonsourceibias.n38 commonsourceibias.n37 161.3
R14596 commonsourceibias.n39 commonsourceibias.n32 161.3
R14597 commonsourceibias.n42 commonsourceibias.n41 161.3
R14598 commonsourceibias.n43 commonsourceibias.n31 161.3
R14599 commonsourceibias.n45 commonsourceibias.n44 161.3
R14600 commonsourceibias.n47 commonsourceibias.n30 161.3
R14601 commonsourceibias.n49 commonsourceibias.n48 161.3
R14602 commonsourceibias.n51 commonsourceibias.n50 161.3
R14603 commonsourceibias.n52 commonsourceibias.n28 161.3
R14604 commonsourceibias.n54 commonsourceibias.n53 161.3
R14605 commonsourceibias.n56 commonsourceibias.n55 161.3
R14606 commonsourceibias.n57 commonsourceibias.n26 161.3
R14607 commonsourceibias.n59 commonsourceibias.n58 161.3
R14608 commonsourceibias.n61 commonsourceibias.n60 161.3
R14609 commonsourceibias.n62 commonsourceibias.n24 161.3
R14610 commonsourceibias.n65 commonsourceibias.n64 161.3
R14611 commonsourceibias.n66 commonsourceibias.n23 161.3
R14612 commonsourceibias.n68 commonsourceibias.n67 161.3
R14613 commonsourceibias.n70 commonsourceibias.n21 161.3
R14614 commonsourceibias.n72 commonsourceibias.n71 161.3
R14615 commonsourceibias.n73 commonsourceibias.n20 161.3
R14616 commonsourceibias.n75 commonsourceibias.n74 161.3
R14617 commonsourceibias.n76 commonsourceibias.n19 161.3
R14618 commonsourceibias.n79 commonsourceibias.n78 161.3
R14619 commonsourceibias.n80 commonsourceibias.n18 161.3
R14620 commonsourceibias.n82 commonsourceibias.n81 161.3
R14621 commonsourceibias.n84 commonsourceibias.n16 161.3
R14622 commonsourceibias.n86 commonsourceibias.n85 161.3
R14623 commonsourceibias.n87 commonsourceibias.n15 161.3
R14624 commonsourceibias.n89 commonsourceibias.n88 161.3
R14625 commonsourceibias.n90 commonsourceibias.n14 161.3
R14626 commonsourceibias.n93 commonsourceibias.n92 161.3
R14627 commonsourceibias.n94 commonsourceibias.n13 161.3
R14628 commonsourceibias.n96 commonsourceibias.n95 161.3
R14629 commonsourceibias.n98 commonsourceibias.n12 161.3
R14630 commonsourceibias.n129 commonsourceibias.n126 161.3
R14631 commonsourceibias.n131 commonsourceibias.n130 161.3
R14632 commonsourceibias.n132 commonsourceibias.n125 161.3
R14633 commonsourceibias.n135 commonsourceibias.n134 161.3
R14634 commonsourceibias.n136 commonsourceibias.n124 161.3
R14635 commonsourceibias.n138 commonsourceibias.n137 161.3
R14636 commonsourceibias.n140 commonsourceibias.n123 161.3
R14637 commonsourceibias.n142 commonsourceibias.n141 161.3
R14638 commonsourceibias.n144 commonsourceibias.n143 161.3
R14639 commonsourceibias.n145 commonsourceibias.n121 161.3
R14640 commonsourceibias.n147 commonsourceibias.n146 161.3
R14641 commonsourceibias.n149 commonsourceibias.n148 161.3
R14642 commonsourceibias.n150 commonsourceibias.n119 161.3
R14643 commonsourceibias.n152 commonsourceibias.n151 161.3
R14644 commonsourceibias.n154 commonsourceibias.n153 161.3
R14645 commonsourceibias.n155 commonsourceibias.n117 161.3
R14646 commonsourceibias.n158 commonsourceibias.n157 161.3
R14647 commonsourceibias.n159 commonsourceibias.n11 161.3
R14648 commonsourceibias.n161 commonsourceibias.n160 161.3
R14649 commonsourceibias.n163 commonsourceibias.n9 161.3
R14650 commonsourceibias.n165 commonsourceibias.n164 161.3
R14651 commonsourceibias.n166 commonsourceibias.n8 161.3
R14652 commonsourceibias.n168 commonsourceibias.n167 161.3
R14653 commonsourceibias.n169 commonsourceibias.n7 161.3
R14654 commonsourceibias.n172 commonsourceibias.n171 161.3
R14655 commonsourceibias.n173 commonsourceibias.n6 161.3
R14656 commonsourceibias.n175 commonsourceibias.n174 161.3
R14657 commonsourceibias.n177 commonsourceibias.n4 161.3
R14658 commonsourceibias.n179 commonsourceibias.n178 161.3
R14659 commonsourceibias.n180 commonsourceibias.n3 161.3
R14660 commonsourceibias.n182 commonsourceibias.n181 161.3
R14661 commonsourceibias.n183 commonsourceibias.n2 161.3
R14662 commonsourceibias.n186 commonsourceibias.n185 161.3
R14663 commonsourceibias.n187 commonsourceibias.n1 161.3
R14664 commonsourceibias.n189 commonsourceibias.n188 161.3
R14665 commonsourceibias.n191 commonsourceibias.n0 161.3
R14666 commonsourceibias.n370 commonsourceibias.n284 161.3
R14667 commonsourceibias.n368 commonsourceibias.n367 161.3
R14668 commonsourceibias.n366 commonsourceibias.n285 161.3
R14669 commonsourceibias.n365 commonsourceibias.n364 161.3
R14670 commonsourceibias.n362 commonsourceibias.n286 161.3
R14671 commonsourceibias.n361 commonsourceibias.n360 161.3
R14672 commonsourceibias.n359 commonsourceibias.n287 161.3
R14673 commonsourceibias.n358 commonsourceibias.n357 161.3
R14674 commonsourceibias.n356 commonsourceibias.n288 161.3
R14675 commonsourceibias.n354 commonsourceibias.n353 161.3
R14676 commonsourceibias.n352 commonsourceibias.n290 161.3
R14677 commonsourceibias.n351 commonsourceibias.n350 161.3
R14678 commonsourceibias.n348 commonsourceibias.n291 161.3
R14679 commonsourceibias.n347 commonsourceibias.n346 161.3
R14680 commonsourceibias.n345 commonsourceibias.n292 161.3
R14681 commonsourceibias.n344 commonsourceibias.n343 161.3
R14682 commonsourceibias.n342 commonsourceibias.n293 161.3
R14683 commonsourceibias.n340 commonsourceibias.n339 161.3
R14684 commonsourceibias.n338 commonsourceibias.n295 161.3
R14685 commonsourceibias.n337 commonsourceibias.n336 161.3
R14686 commonsourceibias.n334 commonsourceibias.n296 161.3
R14687 commonsourceibias.n333 commonsourceibias.n332 161.3
R14688 commonsourceibias.n331 commonsourceibias.n330 161.3
R14689 commonsourceibias.n329 commonsourceibias.n298 161.3
R14690 commonsourceibias.n328 commonsourceibias.n327 161.3
R14691 commonsourceibias.n326 commonsourceibias.n325 161.3
R14692 commonsourceibias.n324 commonsourceibias.n300 161.3
R14693 commonsourceibias.n323 commonsourceibias.n322 161.3
R14694 commonsourceibias.n321 commonsourceibias.n320 161.3
R14695 commonsourceibias.n319 commonsourceibias.n302 161.3
R14696 commonsourceibias.n317 commonsourceibias.n316 161.3
R14697 commonsourceibias.n315 commonsourceibias.n303 161.3
R14698 commonsourceibias.n314 commonsourceibias.n313 161.3
R14699 commonsourceibias.n311 commonsourceibias.n304 161.3
R14700 commonsourceibias.n310 commonsourceibias.n309 161.3
R14701 commonsourceibias.n308 commonsourceibias.n305 161.3
R14702 commonsourceibias.n218 commonsourceibias.n215 161.3
R14703 commonsourceibias.n220 commonsourceibias.n219 161.3
R14704 commonsourceibias.n221 commonsourceibias.n214 161.3
R14705 commonsourceibias.n224 commonsourceibias.n223 161.3
R14706 commonsourceibias.n225 commonsourceibias.n213 161.3
R14707 commonsourceibias.n227 commonsourceibias.n226 161.3
R14708 commonsourceibias.n229 commonsourceibias.n212 161.3
R14709 commonsourceibias.n231 commonsourceibias.n230 161.3
R14710 commonsourceibias.n233 commonsourceibias.n232 161.3
R14711 commonsourceibias.n234 commonsourceibias.n210 161.3
R14712 commonsourceibias.n236 commonsourceibias.n235 161.3
R14713 commonsourceibias.n238 commonsourceibias.n237 161.3
R14714 commonsourceibias.n239 commonsourceibias.n208 161.3
R14715 commonsourceibias.n241 commonsourceibias.n240 161.3
R14716 commonsourceibias.n243 commonsourceibias.n242 161.3
R14717 commonsourceibias.n244 commonsourceibias.n206 161.3
R14718 commonsourceibias.n247 commonsourceibias.n246 161.3
R14719 commonsourceibias.n248 commonsourceibias.n205 161.3
R14720 commonsourceibias.n250 commonsourceibias.n249 161.3
R14721 commonsourceibias.n252 commonsourceibias.n203 161.3
R14722 commonsourceibias.n254 commonsourceibias.n253 161.3
R14723 commonsourceibias.n255 commonsourceibias.n202 161.3
R14724 commonsourceibias.n257 commonsourceibias.n256 161.3
R14725 commonsourceibias.n258 commonsourceibias.n201 161.3
R14726 commonsourceibias.n261 commonsourceibias.n260 161.3
R14727 commonsourceibias.n262 commonsourceibias.n200 161.3
R14728 commonsourceibias.n264 commonsourceibias.n263 161.3
R14729 commonsourceibias.n266 commonsourceibias.n198 161.3
R14730 commonsourceibias.n268 commonsourceibias.n267 161.3
R14731 commonsourceibias.n269 commonsourceibias.n197 161.3
R14732 commonsourceibias.n271 commonsourceibias.n270 161.3
R14733 commonsourceibias.n272 commonsourceibias.n196 161.3
R14734 commonsourceibias.n275 commonsourceibias.n274 161.3
R14735 commonsourceibias.n276 commonsourceibias.n195 161.3
R14736 commonsourceibias.n278 commonsourceibias.n277 161.3
R14737 commonsourceibias.n280 commonsourceibias.n194 161.3
R14738 commonsourceibias.n519 commonsourceibias.n433 161.3
R14739 commonsourceibias.n517 commonsourceibias.n516 161.3
R14740 commonsourceibias.n515 commonsourceibias.n434 161.3
R14741 commonsourceibias.n514 commonsourceibias.n513 161.3
R14742 commonsourceibias.n511 commonsourceibias.n435 161.3
R14743 commonsourceibias.n510 commonsourceibias.n509 161.3
R14744 commonsourceibias.n508 commonsourceibias.n436 161.3
R14745 commonsourceibias.n507 commonsourceibias.n506 161.3
R14746 commonsourceibias.n504 commonsourceibias.n437 161.3
R14747 commonsourceibias.n502 commonsourceibias.n501 161.3
R14748 commonsourceibias.n500 commonsourceibias.n438 161.3
R14749 commonsourceibias.n499 commonsourceibias.n498 161.3
R14750 commonsourceibias.n496 commonsourceibias.n439 161.3
R14751 commonsourceibias.n495 commonsourceibias.n494 161.3
R14752 commonsourceibias.n493 commonsourceibias.n440 161.3
R14753 commonsourceibias.n492 commonsourceibias.n491 161.3
R14754 commonsourceibias.n489 commonsourceibias.n441 161.3
R14755 commonsourceibias.n487 commonsourceibias.n486 161.3
R14756 commonsourceibias.n485 commonsourceibias.n442 161.3
R14757 commonsourceibias.n484 commonsourceibias.n483 161.3
R14758 commonsourceibias.n481 commonsourceibias.n443 161.3
R14759 commonsourceibias.n480 commonsourceibias.n479 161.3
R14760 commonsourceibias.n478 commonsourceibias.n477 161.3
R14761 commonsourceibias.n476 commonsourceibias.n445 161.3
R14762 commonsourceibias.n475 commonsourceibias.n474 161.3
R14763 commonsourceibias.n473 commonsourceibias.n472 161.3
R14764 commonsourceibias.n471 commonsourceibias.n447 161.3
R14765 commonsourceibias.n470 commonsourceibias.n469 161.3
R14766 commonsourceibias.n468 commonsourceibias.n467 161.3
R14767 commonsourceibias.n466 commonsourceibias.n449 161.3
R14768 commonsourceibias.n464 commonsourceibias.n463 161.3
R14769 commonsourceibias.n462 commonsourceibias.n450 161.3
R14770 commonsourceibias.n461 commonsourceibias.n460 161.3
R14771 commonsourceibias.n458 commonsourceibias.n451 161.3
R14772 commonsourceibias.n457 commonsourceibias.n456 161.3
R14773 commonsourceibias.n455 commonsourceibias.n452 161.3
R14774 commonsourceibias.n425 commonsourceibias.n424 161.3
R14775 commonsourceibias.n422 commonsourceibias.n384 161.3
R14776 commonsourceibias.n421 commonsourceibias.n420 161.3
R14777 commonsourceibias.n419 commonsourceibias.n418 161.3
R14778 commonsourceibias.n417 commonsourceibias.n386 161.3
R14779 commonsourceibias.n416 commonsourceibias.n415 161.3
R14780 commonsourceibias.n414 commonsourceibias.n413 161.3
R14781 commonsourceibias.n412 commonsourceibias.n388 161.3
R14782 commonsourceibias.n411 commonsourceibias.n410 161.3
R14783 commonsourceibias.n409 commonsourceibias.n408 161.3
R14784 commonsourceibias.n407 commonsourceibias.n390 161.3
R14785 commonsourceibias.n405 commonsourceibias.n404 161.3
R14786 commonsourceibias.n403 commonsourceibias.n391 161.3
R14787 commonsourceibias.n402 commonsourceibias.n401 161.3
R14788 commonsourceibias.n399 commonsourceibias.n392 161.3
R14789 commonsourceibias.n398 commonsourceibias.n397 161.3
R14790 commonsourceibias.n396 commonsourceibias.n393 161.3
R14791 commonsourceibias.n531 commonsourceibias.n383 161.3
R14792 commonsourceibias.n565 commonsourceibias.n374 161.3
R14793 commonsourceibias.n563 commonsourceibias.n562 161.3
R14794 commonsourceibias.n561 commonsourceibias.n375 161.3
R14795 commonsourceibias.n560 commonsourceibias.n559 161.3
R14796 commonsourceibias.n557 commonsourceibias.n376 161.3
R14797 commonsourceibias.n556 commonsourceibias.n555 161.3
R14798 commonsourceibias.n554 commonsourceibias.n377 161.3
R14799 commonsourceibias.n553 commonsourceibias.n552 161.3
R14800 commonsourceibias.n550 commonsourceibias.n378 161.3
R14801 commonsourceibias.n548 commonsourceibias.n547 161.3
R14802 commonsourceibias.n546 commonsourceibias.n379 161.3
R14803 commonsourceibias.n545 commonsourceibias.n544 161.3
R14804 commonsourceibias.n542 commonsourceibias.n380 161.3
R14805 commonsourceibias.n541 commonsourceibias.n540 161.3
R14806 commonsourceibias.n539 commonsourceibias.n381 161.3
R14807 commonsourceibias.n538 commonsourceibias.n537 161.3
R14808 commonsourceibias.n535 commonsourceibias.n382 161.3
R14809 commonsourceibias.n533 commonsourceibias.n532 161.3
R14810 commonsourceibias.n744 commonsourceibias.n658 161.3
R14811 commonsourceibias.n742 commonsourceibias.n741 161.3
R14812 commonsourceibias.n740 commonsourceibias.n659 161.3
R14813 commonsourceibias.n739 commonsourceibias.n738 161.3
R14814 commonsourceibias.n736 commonsourceibias.n660 161.3
R14815 commonsourceibias.n735 commonsourceibias.n734 161.3
R14816 commonsourceibias.n733 commonsourceibias.n661 161.3
R14817 commonsourceibias.n732 commonsourceibias.n731 161.3
R14818 commonsourceibias.n729 commonsourceibias.n662 161.3
R14819 commonsourceibias.n727 commonsourceibias.n726 161.3
R14820 commonsourceibias.n725 commonsourceibias.n663 161.3
R14821 commonsourceibias.n724 commonsourceibias.n723 161.3
R14822 commonsourceibias.n721 commonsourceibias.n664 161.3
R14823 commonsourceibias.n720 commonsourceibias.n719 161.3
R14824 commonsourceibias.n718 commonsourceibias.n665 161.3
R14825 commonsourceibias.n717 commonsourceibias.n716 161.3
R14826 commonsourceibias.n714 commonsourceibias.n666 161.3
R14827 commonsourceibias.n712 commonsourceibias.n711 161.3
R14828 commonsourceibias.n710 commonsourceibias.n667 161.3
R14829 commonsourceibias.n709 commonsourceibias.n708 161.3
R14830 commonsourceibias.n706 commonsourceibias.n668 161.3
R14831 commonsourceibias.n705 commonsourceibias.n704 161.3
R14832 commonsourceibias.n703 commonsourceibias.n702 161.3
R14833 commonsourceibias.n701 commonsourceibias.n670 161.3
R14834 commonsourceibias.n700 commonsourceibias.n699 161.3
R14835 commonsourceibias.n698 commonsourceibias.n697 161.3
R14836 commonsourceibias.n696 commonsourceibias.n672 161.3
R14837 commonsourceibias.n695 commonsourceibias.n694 161.3
R14838 commonsourceibias.n693 commonsourceibias.n692 161.3
R14839 commonsourceibias.n691 commonsourceibias.n674 161.3
R14840 commonsourceibias.n689 commonsourceibias.n688 161.3
R14841 commonsourceibias.n687 commonsourceibias.n675 161.3
R14842 commonsourceibias.n686 commonsourceibias.n685 161.3
R14843 commonsourceibias.n683 commonsourceibias.n676 161.3
R14844 commonsourceibias.n682 commonsourceibias.n681 161.3
R14845 commonsourceibias.n680 commonsourceibias.n677 161.3
R14846 commonsourceibias.n654 commonsourceibias.n568 161.3
R14847 commonsourceibias.n652 commonsourceibias.n651 161.3
R14848 commonsourceibias.n650 commonsourceibias.n569 161.3
R14849 commonsourceibias.n649 commonsourceibias.n648 161.3
R14850 commonsourceibias.n646 commonsourceibias.n570 161.3
R14851 commonsourceibias.n645 commonsourceibias.n644 161.3
R14852 commonsourceibias.n643 commonsourceibias.n571 161.3
R14853 commonsourceibias.n642 commonsourceibias.n641 161.3
R14854 commonsourceibias.n639 commonsourceibias.n572 161.3
R14855 commonsourceibias.n637 commonsourceibias.n636 161.3
R14856 commonsourceibias.n635 commonsourceibias.n573 161.3
R14857 commonsourceibias.n634 commonsourceibias.n633 161.3
R14858 commonsourceibias.n631 commonsourceibias.n574 161.3
R14859 commonsourceibias.n630 commonsourceibias.n629 161.3
R14860 commonsourceibias.n628 commonsourceibias.n575 161.3
R14861 commonsourceibias.n627 commonsourceibias.n626 161.3
R14862 commonsourceibias.n624 commonsourceibias.n576 161.3
R14863 commonsourceibias.n622 commonsourceibias.n621 161.3
R14864 commonsourceibias.n620 commonsourceibias.n577 161.3
R14865 commonsourceibias.n619 commonsourceibias.n618 161.3
R14866 commonsourceibias.n616 commonsourceibias.n578 161.3
R14867 commonsourceibias.n615 commonsourceibias.n614 161.3
R14868 commonsourceibias.n613 commonsourceibias.n612 161.3
R14869 commonsourceibias.n611 commonsourceibias.n580 161.3
R14870 commonsourceibias.n610 commonsourceibias.n609 161.3
R14871 commonsourceibias.n608 commonsourceibias.n607 161.3
R14872 commonsourceibias.n606 commonsourceibias.n582 161.3
R14873 commonsourceibias.n605 commonsourceibias.n604 161.3
R14874 commonsourceibias.n603 commonsourceibias.n602 161.3
R14875 commonsourceibias.n601 commonsourceibias.n584 161.3
R14876 commonsourceibias.n599 commonsourceibias.n598 161.3
R14877 commonsourceibias.n597 commonsourceibias.n585 161.3
R14878 commonsourceibias.n596 commonsourceibias.n595 161.3
R14879 commonsourceibias.n593 commonsourceibias.n586 161.3
R14880 commonsourceibias.n592 commonsourceibias.n591 161.3
R14881 commonsourceibias.n590 commonsourceibias.n587 161.3
R14882 commonsourceibias.n111 commonsourceibias.n109 81.5057
R14883 commonsourceibias.n428 commonsourceibias.n426 81.5057
R14884 commonsourceibias.n111 commonsourceibias.n110 80.9324
R14885 commonsourceibias.n113 commonsourceibias.n112 80.9324
R14886 commonsourceibias.n115 commonsourceibias.n114 80.9324
R14887 commonsourceibias.n108 commonsourceibias.n107 80.9324
R14888 commonsourceibias.n106 commonsourceibias.n105 80.9324
R14889 commonsourceibias.n104 commonsourceibias.n103 80.9324
R14890 commonsourceibias.n102 commonsourceibias.n101 80.9324
R14891 commonsourceibias.n523 commonsourceibias.n522 80.9324
R14892 commonsourceibias.n525 commonsourceibias.n524 80.9324
R14893 commonsourceibias.n527 commonsourceibias.n526 80.9324
R14894 commonsourceibias.n529 commonsourceibias.n528 80.9324
R14895 commonsourceibias.n432 commonsourceibias.n431 80.9324
R14896 commonsourceibias.n430 commonsourceibias.n429 80.9324
R14897 commonsourceibias.n428 commonsourceibias.n427 80.9324
R14898 commonsourceibias.n100 commonsourceibias.n99 80.6037
R14899 commonsourceibias.n193 commonsourceibias.n192 80.6037
R14900 commonsourceibias.n372 commonsourceibias.n371 80.6037
R14901 commonsourceibias.n282 commonsourceibias.n281 80.6037
R14902 commonsourceibias.n521 commonsourceibias.n520 80.6037
R14903 commonsourceibias.n567 commonsourceibias.n566 80.6037
R14904 commonsourceibias.n746 commonsourceibias.n745 80.6037
R14905 commonsourceibias.n656 commonsourceibias.n655 80.6037
R14906 commonsourceibias.n85 commonsourceibias.n84 56.5617
R14907 commonsourceibias.n71 commonsourceibias.n70 56.5617
R14908 commonsourceibias.n62 commonsourceibias.n61 56.5617
R14909 commonsourceibias.n48 commonsourceibias.n47 56.5617
R14910 commonsourceibias.n178 commonsourceibias.n177 56.5617
R14911 commonsourceibias.n164 commonsourceibias.n163 56.5617
R14912 commonsourceibias.n155 commonsourceibias.n154 56.5617
R14913 commonsourceibias.n141 commonsourceibias.n140 56.5617
R14914 commonsourceibias.n320 commonsourceibias.n319 56.5617
R14915 commonsourceibias.n334 commonsourceibias.n333 56.5617
R14916 commonsourceibias.n343 commonsourceibias.n342 56.5617
R14917 commonsourceibias.n357 commonsourceibias.n356 56.5617
R14918 commonsourceibias.n267 commonsourceibias.n266 56.5617
R14919 commonsourceibias.n253 commonsourceibias.n252 56.5617
R14920 commonsourceibias.n244 commonsourceibias.n243 56.5617
R14921 commonsourceibias.n230 commonsourceibias.n229 56.5617
R14922 commonsourceibias.n467 commonsourceibias.n466 56.5617
R14923 commonsourceibias.n481 commonsourceibias.n480 56.5617
R14924 commonsourceibias.n491 commonsourceibias.n489 56.5617
R14925 commonsourceibias.n506 commonsourceibias.n504 56.5617
R14926 commonsourceibias.n552 commonsourceibias.n550 56.5617
R14927 commonsourceibias.n537 commonsourceibias.n535 56.5617
R14928 commonsourceibias.n408 commonsourceibias.n407 56.5617
R14929 commonsourceibias.n422 commonsourceibias.n421 56.5617
R14930 commonsourceibias.n692 commonsourceibias.n691 56.5617
R14931 commonsourceibias.n706 commonsourceibias.n705 56.5617
R14932 commonsourceibias.n716 commonsourceibias.n714 56.5617
R14933 commonsourceibias.n731 commonsourceibias.n729 56.5617
R14934 commonsourceibias.n602 commonsourceibias.n601 56.5617
R14935 commonsourceibias.n616 commonsourceibias.n615 56.5617
R14936 commonsourceibias.n626 commonsourceibias.n624 56.5617
R14937 commonsourceibias.n641 commonsourceibias.n639 56.5617
R14938 commonsourceibias.n76 commonsourceibias.n75 56.0773
R14939 commonsourceibias.n57 commonsourceibias.n56 56.0773
R14940 commonsourceibias.n169 commonsourceibias.n168 56.0773
R14941 commonsourceibias.n150 commonsourceibias.n149 56.0773
R14942 commonsourceibias.n329 commonsourceibias.n328 56.0773
R14943 commonsourceibias.n348 commonsourceibias.n347 56.0773
R14944 commonsourceibias.n258 commonsourceibias.n257 56.0773
R14945 commonsourceibias.n239 commonsourceibias.n238 56.0773
R14946 commonsourceibias.n476 commonsourceibias.n475 56.0773
R14947 commonsourceibias.n496 commonsourceibias.n495 56.0773
R14948 commonsourceibias.n542 commonsourceibias.n541 56.0773
R14949 commonsourceibias.n417 commonsourceibias.n416 56.0773
R14950 commonsourceibias.n701 commonsourceibias.n700 56.0773
R14951 commonsourceibias.n721 commonsourceibias.n720 56.0773
R14952 commonsourceibias.n611 commonsourceibias.n610 56.0773
R14953 commonsourceibias.n631 commonsourceibias.n630 56.0773
R14954 commonsourceibias.n99 commonsourceibias.n98 55.3321
R14955 commonsourceibias.n192 commonsourceibias.n191 55.3321
R14956 commonsourceibias.n371 commonsourceibias.n370 55.3321
R14957 commonsourceibias.n281 commonsourceibias.n280 55.3321
R14958 commonsourceibias.n520 commonsourceibias.n519 55.3321
R14959 commonsourceibias.n566 commonsourceibias.n565 55.3321
R14960 commonsourceibias.n745 commonsourceibias.n744 55.3321
R14961 commonsourceibias.n655 commonsourceibias.n654 55.3321
R14962 commonsourceibias.n90 commonsourceibias.n89 55.1086
R14963 commonsourceibias.n41 commonsourceibias.n31 55.1086
R14964 commonsourceibias.n183 commonsourceibias.n182 55.1086
R14965 commonsourceibias.n134 commonsourceibias.n124 55.1086
R14966 commonsourceibias.n313 commonsourceibias.n303 55.1086
R14967 commonsourceibias.n362 commonsourceibias.n361 55.1086
R14968 commonsourceibias.n272 commonsourceibias.n271 55.1086
R14969 commonsourceibias.n223 commonsourceibias.n213 55.1086
R14970 commonsourceibias.n460 commonsourceibias.n450 55.1086
R14971 commonsourceibias.n511 commonsourceibias.n510 55.1086
R14972 commonsourceibias.n557 commonsourceibias.n556 55.1086
R14973 commonsourceibias.n401 commonsourceibias.n391 55.1086
R14974 commonsourceibias.n685 commonsourceibias.n675 55.1086
R14975 commonsourceibias.n736 commonsourceibias.n735 55.1086
R14976 commonsourceibias.n595 commonsourceibias.n585 55.1086
R14977 commonsourceibias.n646 commonsourceibias.n645 55.1086
R14978 commonsourceibias.n35 commonsourceibias.n34 47.4592
R14979 commonsourceibias.n128 commonsourceibias.n127 47.4592
R14980 commonsourceibias.n307 commonsourceibias.n306 47.4592
R14981 commonsourceibias.n217 commonsourceibias.n216 47.4592
R14982 commonsourceibias.n454 commonsourceibias.n453 47.4592
R14983 commonsourceibias.n395 commonsourceibias.n394 47.4592
R14984 commonsourceibias.n679 commonsourceibias.n678 47.4592
R14985 commonsourceibias.n589 commonsourceibias.n588 47.4592
R14986 commonsourceibias.n308 commonsourceibias.n307 44.0436
R14987 commonsourceibias.n455 commonsourceibias.n454 44.0436
R14988 commonsourceibias.n396 commonsourceibias.n395 44.0436
R14989 commonsourceibias.n680 commonsourceibias.n679 44.0436
R14990 commonsourceibias.n590 commonsourceibias.n589 44.0436
R14991 commonsourceibias.n36 commonsourceibias.n35 44.0436
R14992 commonsourceibias.n129 commonsourceibias.n128 44.0436
R14993 commonsourceibias.n218 commonsourceibias.n217 44.0436
R14994 commonsourceibias.n92 commonsourceibias.n13 42.5146
R14995 commonsourceibias.n39 commonsourceibias.n38 42.5146
R14996 commonsourceibias.n185 commonsourceibias.n1 42.5146
R14997 commonsourceibias.n132 commonsourceibias.n131 42.5146
R14998 commonsourceibias.n311 commonsourceibias.n310 42.5146
R14999 commonsourceibias.n364 commonsourceibias.n285 42.5146
R15000 commonsourceibias.n274 commonsourceibias.n195 42.5146
R15001 commonsourceibias.n221 commonsourceibias.n220 42.5146
R15002 commonsourceibias.n458 commonsourceibias.n457 42.5146
R15003 commonsourceibias.n513 commonsourceibias.n434 42.5146
R15004 commonsourceibias.n559 commonsourceibias.n375 42.5146
R15005 commonsourceibias.n399 commonsourceibias.n398 42.5146
R15006 commonsourceibias.n683 commonsourceibias.n682 42.5146
R15007 commonsourceibias.n738 commonsourceibias.n659 42.5146
R15008 commonsourceibias.n593 commonsourceibias.n592 42.5146
R15009 commonsourceibias.n648 commonsourceibias.n569 42.5146
R15010 commonsourceibias.n78 commonsourceibias.n18 41.5458
R15011 commonsourceibias.n53 commonsourceibias.n52 41.5458
R15012 commonsourceibias.n171 commonsourceibias.n6 41.5458
R15013 commonsourceibias.n146 commonsourceibias.n145 41.5458
R15014 commonsourceibias.n325 commonsourceibias.n324 41.5458
R15015 commonsourceibias.n350 commonsourceibias.n290 41.5458
R15016 commonsourceibias.n260 commonsourceibias.n200 41.5458
R15017 commonsourceibias.n235 commonsourceibias.n234 41.5458
R15018 commonsourceibias.n472 commonsourceibias.n471 41.5458
R15019 commonsourceibias.n498 commonsourceibias.n438 41.5458
R15020 commonsourceibias.n544 commonsourceibias.n379 41.5458
R15021 commonsourceibias.n413 commonsourceibias.n412 41.5458
R15022 commonsourceibias.n697 commonsourceibias.n696 41.5458
R15023 commonsourceibias.n723 commonsourceibias.n663 41.5458
R15024 commonsourceibias.n607 commonsourceibias.n606 41.5458
R15025 commonsourceibias.n633 commonsourceibias.n573 41.5458
R15026 commonsourceibias.n68 commonsourceibias.n23 40.577
R15027 commonsourceibias.n64 commonsourceibias.n23 40.577
R15028 commonsourceibias.n161 commonsourceibias.n11 40.577
R15029 commonsourceibias.n157 commonsourceibias.n11 40.577
R15030 commonsourceibias.n336 commonsourceibias.n295 40.577
R15031 commonsourceibias.n340 commonsourceibias.n295 40.577
R15032 commonsourceibias.n250 commonsourceibias.n205 40.577
R15033 commonsourceibias.n246 commonsourceibias.n205 40.577
R15034 commonsourceibias.n483 commonsourceibias.n442 40.577
R15035 commonsourceibias.n487 commonsourceibias.n442 40.577
R15036 commonsourceibias.n533 commonsourceibias.n383 40.577
R15037 commonsourceibias.n424 commonsourceibias.n383 40.577
R15038 commonsourceibias.n708 commonsourceibias.n667 40.577
R15039 commonsourceibias.n712 commonsourceibias.n667 40.577
R15040 commonsourceibias.n618 commonsourceibias.n577 40.577
R15041 commonsourceibias.n622 commonsourceibias.n577 40.577
R15042 commonsourceibias.n82 commonsourceibias.n18 39.6083
R15043 commonsourceibias.n52 commonsourceibias.n51 39.6083
R15044 commonsourceibias.n175 commonsourceibias.n6 39.6083
R15045 commonsourceibias.n145 commonsourceibias.n144 39.6083
R15046 commonsourceibias.n324 commonsourceibias.n323 39.6083
R15047 commonsourceibias.n354 commonsourceibias.n290 39.6083
R15048 commonsourceibias.n264 commonsourceibias.n200 39.6083
R15049 commonsourceibias.n234 commonsourceibias.n233 39.6083
R15050 commonsourceibias.n471 commonsourceibias.n470 39.6083
R15051 commonsourceibias.n502 commonsourceibias.n438 39.6083
R15052 commonsourceibias.n548 commonsourceibias.n379 39.6083
R15053 commonsourceibias.n412 commonsourceibias.n411 39.6083
R15054 commonsourceibias.n696 commonsourceibias.n695 39.6083
R15055 commonsourceibias.n727 commonsourceibias.n663 39.6083
R15056 commonsourceibias.n606 commonsourceibias.n605 39.6083
R15057 commonsourceibias.n637 commonsourceibias.n573 39.6083
R15058 commonsourceibias.n96 commonsourceibias.n13 38.6395
R15059 commonsourceibias.n38 commonsourceibias.n33 38.6395
R15060 commonsourceibias.n189 commonsourceibias.n1 38.6395
R15061 commonsourceibias.n131 commonsourceibias.n126 38.6395
R15062 commonsourceibias.n310 commonsourceibias.n305 38.6395
R15063 commonsourceibias.n368 commonsourceibias.n285 38.6395
R15064 commonsourceibias.n278 commonsourceibias.n195 38.6395
R15065 commonsourceibias.n220 commonsourceibias.n215 38.6395
R15066 commonsourceibias.n457 commonsourceibias.n452 38.6395
R15067 commonsourceibias.n517 commonsourceibias.n434 38.6395
R15068 commonsourceibias.n563 commonsourceibias.n375 38.6395
R15069 commonsourceibias.n398 commonsourceibias.n393 38.6395
R15070 commonsourceibias.n682 commonsourceibias.n677 38.6395
R15071 commonsourceibias.n742 commonsourceibias.n659 38.6395
R15072 commonsourceibias.n592 commonsourceibias.n587 38.6395
R15073 commonsourceibias.n652 commonsourceibias.n569 38.6395
R15074 commonsourceibias.n89 commonsourceibias.n15 26.0455
R15075 commonsourceibias.n45 commonsourceibias.n31 26.0455
R15076 commonsourceibias.n182 commonsourceibias.n3 26.0455
R15077 commonsourceibias.n138 commonsourceibias.n124 26.0455
R15078 commonsourceibias.n317 commonsourceibias.n303 26.0455
R15079 commonsourceibias.n361 commonsourceibias.n287 26.0455
R15080 commonsourceibias.n271 commonsourceibias.n197 26.0455
R15081 commonsourceibias.n227 commonsourceibias.n213 26.0455
R15082 commonsourceibias.n464 commonsourceibias.n450 26.0455
R15083 commonsourceibias.n510 commonsourceibias.n436 26.0455
R15084 commonsourceibias.n556 commonsourceibias.n377 26.0455
R15085 commonsourceibias.n405 commonsourceibias.n391 26.0455
R15086 commonsourceibias.n689 commonsourceibias.n675 26.0455
R15087 commonsourceibias.n735 commonsourceibias.n661 26.0455
R15088 commonsourceibias.n599 commonsourceibias.n585 26.0455
R15089 commonsourceibias.n645 commonsourceibias.n571 26.0455
R15090 commonsourceibias.n75 commonsourceibias.n20 25.0767
R15091 commonsourceibias.n58 commonsourceibias.n57 25.0767
R15092 commonsourceibias.n168 commonsourceibias.n8 25.0767
R15093 commonsourceibias.n151 commonsourceibias.n150 25.0767
R15094 commonsourceibias.n330 commonsourceibias.n329 25.0767
R15095 commonsourceibias.n347 commonsourceibias.n292 25.0767
R15096 commonsourceibias.n257 commonsourceibias.n202 25.0767
R15097 commonsourceibias.n240 commonsourceibias.n239 25.0767
R15098 commonsourceibias.n477 commonsourceibias.n476 25.0767
R15099 commonsourceibias.n495 commonsourceibias.n440 25.0767
R15100 commonsourceibias.n541 commonsourceibias.n381 25.0767
R15101 commonsourceibias.n418 commonsourceibias.n417 25.0767
R15102 commonsourceibias.n702 commonsourceibias.n701 25.0767
R15103 commonsourceibias.n720 commonsourceibias.n665 25.0767
R15104 commonsourceibias.n612 commonsourceibias.n611 25.0767
R15105 commonsourceibias.n630 commonsourceibias.n575 25.0767
R15106 commonsourceibias.n71 commonsourceibias.n22 24.3464
R15107 commonsourceibias.n61 commonsourceibias.n25 24.3464
R15108 commonsourceibias.n164 commonsourceibias.n10 24.3464
R15109 commonsourceibias.n154 commonsourceibias.n118 24.3464
R15110 commonsourceibias.n333 commonsourceibias.n297 24.3464
R15111 commonsourceibias.n343 commonsourceibias.n294 24.3464
R15112 commonsourceibias.n253 commonsourceibias.n204 24.3464
R15113 commonsourceibias.n243 commonsourceibias.n207 24.3464
R15114 commonsourceibias.n480 commonsourceibias.n444 24.3464
R15115 commonsourceibias.n491 commonsourceibias.n490 24.3464
R15116 commonsourceibias.n537 commonsourceibias.n536 24.3464
R15117 commonsourceibias.n421 commonsourceibias.n385 24.3464
R15118 commonsourceibias.n705 commonsourceibias.n669 24.3464
R15119 commonsourceibias.n716 commonsourceibias.n715 24.3464
R15120 commonsourceibias.n615 commonsourceibias.n579 24.3464
R15121 commonsourceibias.n626 commonsourceibias.n625 24.3464
R15122 commonsourceibias.n85 commonsourceibias.n17 23.8546
R15123 commonsourceibias.n47 commonsourceibias.n46 23.8546
R15124 commonsourceibias.n178 commonsourceibias.n5 23.8546
R15125 commonsourceibias.n140 commonsourceibias.n139 23.8546
R15126 commonsourceibias.n319 commonsourceibias.n318 23.8546
R15127 commonsourceibias.n357 commonsourceibias.n289 23.8546
R15128 commonsourceibias.n267 commonsourceibias.n199 23.8546
R15129 commonsourceibias.n229 commonsourceibias.n228 23.8546
R15130 commonsourceibias.n466 commonsourceibias.n465 23.8546
R15131 commonsourceibias.n506 commonsourceibias.n505 23.8546
R15132 commonsourceibias.n552 commonsourceibias.n551 23.8546
R15133 commonsourceibias.n407 commonsourceibias.n406 23.8546
R15134 commonsourceibias.n691 commonsourceibias.n690 23.8546
R15135 commonsourceibias.n731 commonsourceibias.n730 23.8546
R15136 commonsourceibias.n601 commonsourceibias.n600 23.8546
R15137 commonsourceibias.n641 commonsourceibias.n640 23.8546
R15138 commonsourceibias.n98 commonsourceibias.n97 17.4607
R15139 commonsourceibias.n191 commonsourceibias.n190 17.4607
R15140 commonsourceibias.n370 commonsourceibias.n369 17.4607
R15141 commonsourceibias.n280 commonsourceibias.n279 17.4607
R15142 commonsourceibias.n519 commonsourceibias.n518 17.4607
R15143 commonsourceibias.n565 commonsourceibias.n564 17.4607
R15144 commonsourceibias.n744 commonsourceibias.n743 17.4607
R15145 commonsourceibias.n654 commonsourceibias.n653 17.4607
R15146 commonsourceibias.n84 commonsourceibias.n83 16.9689
R15147 commonsourceibias.n48 commonsourceibias.n29 16.9689
R15148 commonsourceibias.n177 commonsourceibias.n176 16.9689
R15149 commonsourceibias.n141 commonsourceibias.n122 16.9689
R15150 commonsourceibias.n320 commonsourceibias.n301 16.9689
R15151 commonsourceibias.n356 commonsourceibias.n355 16.9689
R15152 commonsourceibias.n266 commonsourceibias.n265 16.9689
R15153 commonsourceibias.n230 commonsourceibias.n211 16.9689
R15154 commonsourceibias.n467 commonsourceibias.n448 16.9689
R15155 commonsourceibias.n504 commonsourceibias.n503 16.9689
R15156 commonsourceibias.n550 commonsourceibias.n549 16.9689
R15157 commonsourceibias.n408 commonsourceibias.n389 16.9689
R15158 commonsourceibias.n692 commonsourceibias.n673 16.9689
R15159 commonsourceibias.n729 commonsourceibias.n728 16.9689
R15160 commonsourceibias.n602 commonsourceibias.n583 16.9689
R15161 commonsourceibias.n639 commonsourceibias.n638 16.9689
R15162 commonsourceibias.n70 commonsourceibias.n69 16.477
R15163 commonsourceibias.n63 commonsourceibias.n62 16.477
R15164 commonsourceibias.n163 commonsourceibias.n162 16.477
R15165 commonsourceibias.n156 commonsourceibias.n155 16.477
R15166 commonsourceibias.n335 commonsourceibias.n334 16.477
R15167 commonsourceibias.n342 commonsourceibias.n341 16.477
R15168 commonsourceibias.n252 commonsourceibias.n251 16.477
R15169 commonsourceibias.n245 commonsourceibias.n244 16.477
R15170 commonsourceibias.n482 commonsourceibias.n481 16.477
R15171 commonsourceibias.n489 commonsourceibias.n488 16.477
R15172 commonsourceibias.n535 commonsourceibias.n534 16.477
R15173 commonsourceibias.n423 commonsourceibias.n422 16.477
R15174 commonsourceibias.n707 commonsourceibias.n706 16.477
R15175 commonsourceibias.n714 commonsourceibias.n713 16.477
R15176 commonsourceibias.n617 commonsourceibias.n616 16.477
R15177 commonsourceibias.n624 commonsourceibias.n623 16.477
R15178 commonsourceibias.n77 commonsourceibias.n76 15.9852
R15179 commonsourceibias.n56 commonsourceibias.n27 15.9852
R15180 commonsourceibias.n170 commonsourceibias.n169 15.9852
R15181 commonsourceibias.n149 commonsourceibias.n120 15.9852
R15182 commonsourceibias.n328 commonsourceibias.n299 15.9852
R15183 commonsourceibias.n349 commonsourceibias.n348 15.9852
R15184 commonsourceibias.n259 commonsourceibias.n258 15.9852
R15185 commonsourceibias.n238 commonsourceibias.n209 15.9852
R15186 commonsourceibias.n475 commonsourceibias.n446 15.9852
R15187 commonsourceibias.n497 commonsourceibias.n496 15.9852
R15188 commonsourceibias.n543 commonsourceibias.n542 15.9852
R15189 commonsourceibias.n416 commonsourceibias.n387 15.9852
R15190 commonsourceibias.n700 commonsourceibias.n671 15.9852
R15191 commonsourceibias.n722 commonsourceibias.n721 15.9852
R15192 commonsourceibias.n610 commonsourceibias.n581 15.9852
R15193 commonsourceibias.n632 commonsourceibias.n631 15.9852
R15194 commonsourceibias.n91 commonsourceibias.n90 15.4934
R15195 commonsourceibias.n41 commonsourceibias.n40 15.4934
R15196 commonsourceibias.n184 commonsourceibias.n183 15.4934
R15197 commonsourceibias.n134 commonsourceibias.n133 15.4934
R15198 commonsourceibias.n313 commonsourceibias.n312 15.4934
R15199 commonsourceibias.n363 commonsourceibias.n362 15.4934
R15200 commonsourceibias.n273 commonsourceibias.n272 15.4934
R15201 commonsourceibias.n223 commonsourceibias.n222 15.4934
R15202 commonsourceibias.n460 commonsourceibias.n459 15.4934
R15203 commonsourceibias.n512 commonsourceibias.n511 15.4934
R15204 commonsourceibias.n558 commonsourceibias.n557 15.4934
R15205 commonsourceibias.n401 commonsourceibias.n400 15.4934
R15206 commonsourceibias.n685 commonsourceibias.n684 15.4934
R15207 commonsourceibias.n737 commonsourceibias.n736 15.4934
R15208 commonsourceibias.n595 commonsourceibias.n594 15.4934
R15209 commonsourceibias.n647 commonsourceibias.n646 15.4934
R15210 commonsourceibias.n102 commonsourceibias.n100 13.2663
R15211 commonsourceibias.n523 commonsourceibias.n521 13.2663
R15212 commonsourceibias.n748 commonsourceibias.n373 10.122
R15213 commonsourceibias.n159 commonsourceibias.n116 9.50363
R15214 commonsourceibias.n531 commonsourceibias.n530 9.50363
R15215 commonsourceibias.n92 commonsourceibias.n91 9.09948
R15216 commonsourceibias.n40 commonsourceibias.n39 9.09948
R15217 commonsourceibias.n185 commonsourceibias.n184 9.09948
R15218 commonsourceibias.n133 commonsourceibias.n132 9.09948
R15219 commonsourceibias.n312 commonsourceibias.n311 9.09948
R15220 commonsourceibias.n364 commonsourceibias.n363 9.09948
R15221 commonsourceibias.n274 commonsourceibias.n273 9.09948
R15222 commonsourceibias.n222 commonsourceibias.n221 9.09948
R15223 commonsourceibias.n459 commonsourceibias.n458 9.09948
R15224 commonsourceibias.n513 commonsourceibias.n512 9.09948
R15225 commonsourceibias.n559 commonsourceibias.n558 9.09948
R15226 commonsourceibias.n400 commonsourceibias.n399 9.09948
R15227 commonsourceibias.n684 commonsourceibias.n683 9.09948
R15228 commonsourceibias.n738 commonsourceibias.n737 9.09948
R15229 commonsourceibias.n594 commonsourceibias.n593 9.09948
R15230 commonsourceibias.n648 commonsourceibias.n647 9.09948
R15231 commonsourceibias.n283 commonsourceibias.n193 8.79451
R15232 commonsourceibias.n657 commonsourceibias.n567 8.79451
R15233 commonsourceibias.n78 commonsourceibias.n77 8.60764
R15234 commonsourceibias.n53 commonsourceibias.n27 8.60764
R15235 commonsourceibias.n171 commonsourceibias.n170 8.60764
R15236 commonsourceibias.n146 commonsourceibias.n120 8.60764
R15237 commonsourceibias.n325 commonsourceibias.n299 8.60764
R15238 commonsourceibias.n350 commonsourceibias.n349 8.60764
R15239 commonsourceibias.n260 commonsourceibias.n259 8.60764
R15240 commonsourceibias.n235 commonsourceibias.n209 8.60764
R15241 commonsourceibias.n472 commonsourceibias.n446 8.60764
R15242 commonsourceibias.n498 commonsourceibias.n497 8.60764
R15243 commonsourceibias.n544 commonsourceibias.n543 8.60764
R15244 commonsourceibias.n413 commonsourceibias.n387 8.60764
R15245 commonsourceibias.n697 commonsourceibias.n671 8.60764
R15246 commonsourceibias.n723 commonsourceibias.n722 8.60764
R15247 commonsourceibias.n607 commonsourceibias.n581 8.60764
R15248 commonsourceibias.n633 commonsourceibias.n632 8.60764
R15249 commonsourceibias.n748 commonsourceibias.n747 8.46921
R15250 commonsourceibias.n69 commonsourceibias.n68 8.11581
R15251 commonsourceibias.n64 commonsourceibias.n63 8.11581
R15252 commonsourceibias.n162 commonsourceibias.n161 8.11581
R15253 commonsourceibias.n157 commonsourceibias.n156 8.11581
R15254 commonsourceibias.n336 commonsourceibias.n335 8.11581
R15255 commonsourceibias.n341 commonsourceibias.n340 8.11581
R15256 commonsourceibias.n251 commonsourceibias.n250 8.11581
R15257 commonsourceibias.n246 commonsourceibias.n245 8.11581
R15258 commonsourceibias.n483 commonsourceibias.n482 8.11581
R15259 commonsourceibias.n488 commonsourceibias.n487 8.11581
R15260 commonsourceibias.n534 commonsourceibias.n533 8.11581
R15261 commonsourceibias.n424 commonsourceibias.n423 8.11581
R15262 commonsourceibias.n708 commonsourceibias.n707 8.11581
R15263 commonsourceibias.n713 commonsourceibias.n712 8.11581
R15264 commonsourceibias.n618 commonsourceibias.n617 8.11581
R15265 commonsourceibias.n623 commonsourceibias.n622 8.11581
R15266 commonsourceibias.n83 commonsourceibias.n82 7.62397
R15267 commonsourceibias.n51 commonsourceibias.n29 7.62397
R15268 commonsourceibias.n176 commonsourceibias.n175 7.62397
R15269 commonsourceibias.n144 commonsourceibias.n122 7.62397
R15270 commonsourceibias.n323 commonsourceibias.n301 7.62397
R15271 commonsourceibias.n355 commonsourceibias.n354 7.62397
R15272 commonsourceibias.n265 commonsourceibias.n264 7.62397
R15273 commonsourceibias.n233 commonsourceibias.n211 7.62397
R15274 commonsourceibias.n470 commonsourceibias.n448 7.62397
R15275 commonsourceibias.n503 commonsourceibias.n502 7.62397
R15276 commonsourceibias.n549 commonsourceibias.n548 7.62397
R15277 commonsourceibias.n411 commonsourceibias.n389 7.62397
R15278 commonsourceibias.n695 commonsourceibias.n673 7.62397
R15279 commonsourceibias.n728 commonsourceibias.n727 7.62397
R15280 commonsourceibias.n605 commonsourceibias.n583 7.62397
R15281 commonsourceibias.n638 commonsourceibias.n637 7.62397
R15282 commonsourceibias.n97 commonsourceibias.n96 7.13213
R15283 commonsourceibias.n34 commonsourceibias.n33 7.13213
R15284 commonsourceibias.n190 commonsourceibias.n189 7.13213
R15285 commonsourceibias.n127 commonsourceibias.n126 7.13213
R15286 commonsourceibias.n306 commonsourceibias.n305 7.13213
R15287 commonsourceibias.n369 commonsourceibias.n368 7.13213
R15288 commonsourceibias.n279 commonsourceibias.n278 7.13213
R15289 commonsourceibias.n216 commonsourceibias.n215 7.13213
R15290 commonsourceibias.n453 commonsourceibias.n452 7.13213
R15291 commonsourceibias.n518 commonsourceibias.n517 7.13213
R15292 commonsourceibias.n564 commonsourceibias.n563 7.13213
R15293 commonsourceibias.n394 commonsourceibias.n393 7.13213
R15294 commonsourceibias.n678 commonsourceibias.n677 7.13213
R15295 commonsourceibias.n743 commonsourceibias.n742 7.13213
R15296 commonsourceibias.n588 commonsourceibias.n587 7.13213
R15297 commonsourceibias.n653 commonsourceibias.n652 7.13213
R15298 commonsourceibias.n373 commonsourceibias.n372 5.06534
R15299 commonsourceibias.n283 commonsourceibias.n282 5.06534
R15300 commonsourceibias.n747 commonsourceibias.n746 5.06534
R15301 commonsourceibias.n657 commonsourceibias.n656 5.06534
R15302 commonsourceibias commonsourceibias.n748 4.04308
R15303 commonsourceibias.n373 commonsourceibias.n283 3.72967
R15304 commonsourceibias.n747 commonsourceibias.n657 3.72967
R15305 commonsourceibias.n109 commonsourceibias.t51 2.82907
R15306 commonsourceibias.n109 commonsourceibias.t1 2.82907
R15307 commonsourceibias.n110 commonsourceibias.t55 2.82907
R15308 commonsourceibias.n110 commonsourceibias.t19 2.82907
R15309 commonsourceibias.n112 commonsourceibias.t25 2.82907
R15310 commonsourceibias.n112 commonsourceibias.t31 2.82907
R15311 commonsourceibias.n114 commonsourceibias.t15 2.82907
R15312 commonsourceibias.n114 commonsourceibias.t45 2.82907
R15313 commonsourceibias.n107 commonsourceibias.t29 2.82907
R15314 commonsourceibias.n107 commonsourceibias.t7 2.82907
R15315 commonsourceibias.n105 commonsourceibias.t59 2.82907
R15316 commonsourceibias.n105 commonsourceibias.t17 2.82907
R15317 commonsourceibias.n103 commonsourceibias.t5 2.82907
R15318 commonsourceibias.n103 commonsourceibias.t11 2.82907
R15319 commonsourceibias.n101 commonsourceibias.t13 2.82907
R15320 commonsourceibias.n101 commonsourceibias.t49 2.82907
R15321 commonsourceibias.n522 commonsourceibias.t61 2.82907
R15322 commonsourceibias.n522 commonsourceibias.t35 2.82907
R15323 commonsourceibias.n524 commonsourceibias.t33 2.82907
R15324 commonsourceibias.n524 commonsourceibias.t21 2.82907
R15325 commonsourceibias.n526 commonsourceibias.t39 2.82907
R15326 commonsourceibias.n526 commonsourceibias.t9 2.82907
R15327 commonsourceibias.n528 commonsourceibias.t27 2.82907
R15328 commonsourceibias.n528 commonsourceibias.t47 2.82907
R15329 commonsourceibias.n431 commonsourceibias.t57 2.82907
R15330 commonsourceibias.n431 commonsourceibias.t37 2.82907
R15331 commonsourceibias.n429 commonsourceibias.t53 2.82907
R15332 commonsourceibias.n429 commonsourceibias.t43 2.82907
R15333 commonsourceibias.n427 commonsourceibias.t41 2.82907
R15334 commonsourceibias.n427 commonsourceibias.t3 2.82907
R15335 commonsourceibias.n426 commonsourceibias.t23 2.82907
R15336 commonsourceibias.n426 commonsourceibias.t63 2.82907
R15337 commonsourceibias.n17 commonsourceibias.n15 0.738255
R15338 commonsourceibias.n46 commonsourceibias.n45 0.738255
R15339 commonsourceibias.n5 commonsourceibias.n3 0.738255
R15340 commonsourceibias.n139 commonsourceibias.n138 0.738255
R15341 commonsourceibias.n318 commonsourceibias.n317 0.738255
R15342 commonsourceibias.n289 commonsourceibias.n287 0.738255
R15343 commonsourceibias.n199 commonsourceibias.n197 0.738255
R15344 commonsourceibias.n228 commonsourceibias.n227 0.738255
R15345 commonsourceibias.n465 commonsourceibias.n464 0.738255
R15346 commonsourceibias.n505 commonsourceibias.n436 0.738255
R15347 commonsourceibias.n551 commonsourceibias.n377 0.738255
R15348 commonsourceibias.n406 commonsourceibias.n405 0.738255
R15349 commonsourceibias.n690 commonsourceibias.n689 0.738255
R15350 commonsourceibias.n730 commonsourceibias.n661 0.738255
R15351 commonsourceibias.n600 commonsourceibias.n599 0.738255
R15352 commonsourceibias.n640 commonsourceibias.n571 0.738255
R15353 commonsourceibias.n104 commonsourceibias.n102 0.573776
R15354 commonsourceibias.n106 commonsourceibias.n104 0.573776
R15355 commonsourceibias.n108 commonsourceibias.n106 0.573776
R15356 commonsourceibias.n115 commonsourceibias.n113 0.573776
R15357 commonsourceibias.n113 commonsourceibias.n111 0.573776
R15358 commonsourceibias.n430 commonsourceibias.n428 0.573776
R15359 commonsourceibias.n432 commonsourceibias.n430 0.573776
R15360 commonsourceibias.n529 commonsourceibias.n527 0.573776
R15361 commonsourceibias.n527 commonsourceibias.n525 0.573776
R15362 commonsourceibias.n525 commonsourceibias.n523 0.573776
R15363 commonsourceibias.n116 commonsourceibias.n108 0.287138
R15364 commonsourceibias.n116 commonsourceibias.n115 0.287138
R15365 commonsourceibias.n530 commonsourceibias.n432 0.287138
R15366 commonsourceibias.n530 commonsourceibias.n529 0.287138
R15367 commonsourceibias.n100 commonsourceibias.n12 0.285035
R15368 commonsourceibias.n193 commonsourceibias.n0 0.285035
R15369 commonsourceibias.n372 commonsourceibias.n284 0.285035
R15370 commonsourceibias.n282 commonsourceibias.n194 0.285035
R15371 commonsourceibias.n521 commonsourceibias.n433 0.285035
R15372 commonsourceibias.n567 commonsourceibias.n374 0.285035
R15373 commonsourceibias.n746 commonsourceibias.n658 0.285035
R15374 commonsourceibias.n656 commonsourceibias.n568 0.285035
R15375 commonsourceibias.n22 commonsourceibias.n20 0.246418
R15376 commonsourceibias.n58 commonsourceibias.n25 0.246418
R15377 commonsourceibias.n10 commonsourceibias.n8 0.246418
R15378 commonsourceibias.n151 commonsourceibias.n118 0.246418
R15379 commonsourceibias.n330 commonsourceibias.n297 0.246418
R15380 commonsourceibias.n294 commonsourceibias.n292 0.246418
R15381 commonsourceibias.n204 commonsourceibias.n202 0.246418
R15382 commonsourceibias.n240 commonsourceibias.n207 0.246418
R15383 commonsourceibias.n477 commonsourceibias.n444 0.246418
R15384 commonsourceibias.n490 commonsourceibias.n440 0.246418
R15385 commonsourceibias.n536 commonsourceibias.n381 0.246418
R15386 commonsourceibias.n418 commonsourceibias.n385 0.246418
R15387 commonsourceibias.n702 commonsourceibias.n669 0.246418
R15388 commonsourceibias.n715 commonsourceibias.n665 0.246418
R15389 commonsourceibias.n612 commonsourceibias.n579 0.246418
R15390 commonsourceibias.n625 commonsourceibias.n575 0.246418
R15391 commonsourceibias.n95 commonsourceibias.n12 0.189894
R15392 commonsourceibias.n95 commonsourceibias.n94 0.189894
R15393 commonsourceibias.n94 commonsourceibias.n93 0.189894
R15394 commonsourceibias.n93 commonsourceibias.n14 0.189894
R15395 commonsourceibias.n88 commonsourceibias.n14 0.189894
R15396 commonsourceibias.n88 commonsourceibias.n87 0.189894
R15397 commonsourceibias.n87 commonsourceibias.n86 0.189894
R15398 commonsourceibias.n86 commonsourceibias.n16 0.189894
R15399 commonsourceibias.n81 commonsourceibias.n16 0.189894
R15400 commonsourceibias.n81 commonsourceibias.n80 0.189894
R15401 commonsourceibias.n80 commonsourceibias.n79 0.189894
R15402 commonsourceibias.n79 commonsourceibias.n19 0.189894
R15403 commonsourceibias.n74 commonsourceibias.n19 0.189894
R15404 commonsourceibias.n74 commonsourceibias.n73 0.189894
R15405 commonsourceibias.n73 commonsourceibias.n72 0.189894
R15406 commonsourceibias.n72 commonsourceibias.n21 0.189894
R15407 commonsourceibias.n67 commonsourceibias.n21 0.189894
R15408 commonsourceibias.n67 commonsourceibias.n66 0.189894
R15409 commonsourceibias.n66 commonsourceibias.n65 0.189894
R15410 commonsourceibias.n65 commonsourceibias.n24 0.189894
R15411 commonsourceibias.n60 commonsourceibias.n24 0.189894
R15412 commonsourceibias.n60 commonsourceibias.n59 0.189894
R15413 commonsourceibias.n59 commonsourceibias.n26 0.189894
R15414 commonsourceibias.n55 commonsourceibias.n26 0.189894
R15415 commonsourceibias.n55 commonsourceibias.n54 0.189894
R15416 commonsourceibias.n54 commonsourceibias.n28 0.189894
R15417 commonsourceibias.n50 commonsourceibias.n28 0.189894
R15418 commonsourceibias.n50 commonsourceibias.n49 0.189894
R15419 commonsourceibias.n49 commonsourceibias.n30 0.189894
R15420 commonsourceibias.n44 commonsourceibias.n30 0.189894
R15421 commonsourceibias.n44 commonsourceibias.n43 0.189894
R15422 commonsourceibias.n43 commonsourceibias.n42 0.189894
R15423 commonsourceibias.n42 commonsourceibias.n32 0.189894
R15424 commonsourceibias.n37 commonsourceibias.n32 0.189894
R15425 commonsourceibias.n37 commonsourceibias.n36 0.189894
R15426 commonsourceibias.n158 commonsourceibias.n117 0.189894
R15427 commonsourceibias.n153 commonsourceibias.n117 0.189894
R15428 commonsourceibias.n153 commonsourceibias.n152 0.189894
R15429 commonsourceibias.n152 commonsourceibias.n119 0.189894
R15430 commonsourceibias.n148 commonsourceibias.n119 0.189894
R15431 commonsourceibias.n148 commonsourceibias.n147 0.189894
R15432 commonsourceibias.n147 commonsourceibias.n121 0.189894
R15433 commonsourceibias.n143 commonsourceibias.n121 0.189894
R15434 commonsourceibias.n143 commonsourceibias.n142 0.189894
R15435 commonsourceibias.n142 commonsourceibias.n123 0.189894
R15436 commonsourceibias.n137 commonsourceibias.n123 0.189894
R15437 commonsourceibias.n137 commonsourceibias.n136 0.189894
R15438 commonsourceibias.n136 commonsourceibias.n135 0.189894
R15439 commonsourceibias.n135 commonsourceibias.n125 0.189894
R15440 commonsourceibias.n130 commonsourceibias.n125 0.189894
R15441 commonsourceibias.n130 commonsourceibias.n129 0.189894
R15442 commonsourceibias.n188 commonsourceibias.n0 0.189894
R15443 commonsourceibias.n188 commonsourceibias.n187 0.189894
R15444 commonsourceibias.n187 commonsourceibias.n186 0.189894
R15445 commonsourceibias.n186 commonsourceibias.n2 0.189894
R15446 commonsourceibias.n181 commonsourceibias.n2 0.189894
R15447 commonsourceibias.n181 commonsourceibias.n180 0.189894
R15448 commonsourceibias.n180 commonsourceibias.n179 0.189894
R15449 commonsourceibias.n179 commonsourceibias.n4 0.189894
R15450 commonsourceibias.n174 commonsourceibias.n4 0.189894
R15451 commonsourceibias.n174 commonsourceibias.n173 0.189894
R15452 commonsourceibias.n173 commonsourceibias.n172 0.189894
R15453 commonsourceibias.n172 commonsourceibias.n7 0.189894
R15454 commonsourceibias.n167 commonsourceibias.n7 0.189894
R15455 commonsourceibias.n167 commonsourceibias.n166 0.189894
R15456 commonsourceibias.n166 commonsourceibias.n165 0.189894
R15457 commonsourceibias.n165 commonsourceibias.n9 0.189894
R15458 commonsourceibias.n160 commonsourceibias.n9 0.189894
R15459 commonsourceibias.n367 commonsourceibias.n284 0.189894
R15460 commonsourceibias.n367 commonsourceibias.n366 0.189894
R15461 commonsourceibias.n366 commonsourceibias.n365 0.189894
R15462 commonsourceibias.n365 commonsourceibias.n286 0.189894
R15463 commonsourceibias.n360 commonsourceibias.n286 0.189894
R15464 commonsourceibias.n360 commonsourceibias.n359 0.189894
R15465 commonsourceibias.n359 commonsourceibias.n358 0.189894
R15466 commonsourceibias.n358 commonsourceibias.n288 0.189894
R15467 commonsourceibias.n353 commonsourceibias.n288 0.189894
R15468 commonsourceibias.n353 commonsourceibias.n352 0.189894
R15469 commonsourceibias.n352 commonsourceibias.n351 0.189894
R15470 commonsourceibias.n351 commonsourceibias.n291 0.189894
R15471 commonsourceibias.n346 commonsourceibias.n291 0.189894
R15472 commonsourceibias.n346 commonsourceibias.n345 0.189894
R15473 commonsourceibias.n345 commonsourceibias.n344 0.189894
R15474 commonsourceibias.n344 commonsourceibias.n293 0.189894
R15475 commonsourceibias.n339 commonsourceibias.n293 0.189894
R15476 commonsourceibias.n339 commonsourceibias.n338 0.189894
R15477 commonsourceibias.n338 commonsourceibias.n337 0.189894
R15478 commonsourceibias.n337 commonsourceibias.n296 0.189894
R15479 commonsourceibias.n332 commonsourceibias.n296 0.189894
R15480 commonsourceibias.n332 commonsourceibias.n331 0.189894
R15481 commonsourceibias.n331 commonsourceibias.n298 0.189894
R15482 commonsourceibias.n327 commonsourceibias.n298 0.189894
R15483 commonsourceibias.n327 commonsourceibias.n326 0.189894
R15484 commonsourceibias.n326 commonsourceibias.n300 0.189894
R15485 commonsourceibias.n322 commonsourceibias.n300 0.189894
R15486 commonsourceibias.n322 commonsourceibias.n321 0.189894
R15487 commonsourceibias.n321 commonsourceibias.n302 0.189894
R15488 commonsourceibias.n316 commonsourceibias.n302 0.189894
R15489 commonsourceibias.n316 commonsourceibias.n315 0.189894
R15490 commonsourceibias.n315 commonsourceibias.n314 0.189894
R15491 commonsourceibias.n314 commonsourceibias.n304 0.189894
R15492 commonsourceibias.n309 commonsourceibias.n304 0.189894
R15493 commonsourceibias.n309 commonsourceibias.n308 0.189894
R15494 commonsourceibias.n277 commonsourceibias.n194 0.189894
R15495 commonsourceibias.n277 commonsourceibias.n276 0.189894
R15496 commonsourceibias.n276 commonsourceibias.n275 0.189894
R15497 commonsourceibias.n275 commonsourceibias.n196 0.189894
R15498 commonsourceibias.n270 commonsourceibias.n196 0.189894
R15499 commonsourceibias.n270 commonsourceibias.n269 0.189894
R15500 commonsourceibias.n269 commonsourceibias.n268 0.189894
R15501 commonsourceibias.n268 commonsourceibias.n198 0.189894
R15502 commonsourceibias.n263 commonsourceibias.n198 0.189894
R15503 commonsourceibias.n263 commonsourceibias.n262 0.189894
R15504 commonsourceibias.n262 commonsourceibias.n261 0.189894
R15505 commonsourceibias.n261 commonsourceibias.n201 0.189894
R15506 commonsourceibias.n256 commonsourceibias.n201 0.189894
R15507 commonsourceibias.n256 commonsourceibias.n255 0.189894
R15508 commonsourceibias.n255 commonsourceibias.n254 0.189894
R15509 commonsourceibias.n254 commonsourceibias.n203 0.189894
R15510 commonsourceibias.n249 commonsourceibias.n203 0.189894
R15511 commonsourceibias.n249 commonsourceibias.n248 0.189894
R15512 commonsourceibias.n248 commonsourceibias.n247 0.189894
R15513 commonsourceibias.n247 commonsourceibias.n206 0.189894
R15514 commonsourceibias.n242 commonsourceibias.n206 0.189894
R15515 commonsourceibias.n242 commonsourceibias.n241 0.189894
R15516 commonsourceibias.n241 commonsourceibias.n208 0.189894
R15517 commonsourceibias.n237 commonsourceibias.n208 0.189894
R15518 commonsourceibias.n237 commonsourceibias.n236 0.189894
R15519 commonsourceibias.n236 commonsourceibias.n210 0.189894
R15520 commonsourceibias.n232 commonsourceibias.n210 0.189894
R15521 commonsourceibias.n232 commonsourceibias.n231 0.189894
R15522 commonsourceibias.n231 commonsourceibias.n212 0.189894
R15523 commonsourceibias.n226 commonsourceibias.n212 0.189894
R15524 commonsourceibias.n226 commonsourceibias.n225 0.189894
R15525 commonsourceibias.n225 commonsourceibias.n224 0.189894
R15526 commonsourceibias.n224 commonsourceibias.n214 0.189894
R15527 commonsourceibias.n219 commonsourceibias.n214 0.189894
R15528 commonsourceibias.n219 commonsourceibias.n218 0.189894
R15529 commonsourceibias.n456 commonsourceibias.n455 0.189894
R15530 commonsourceibias.n456 commonsourceibias.n451 0.189894
R15531 commonsourceibias.n461 commonsourceibias.n451 0.189894
R15532 commonsourceibias.n462 commonsourceibias.n461 0.189894
R15533 commonsourceibias.n463 commonsourceibias.n462 0.189894
R15534 commonsourceibias.n463 commonsourceibias.n449 0.189894
R15535 commonsourceibias.n468 commonsourceibias.n449 0.189894
R15536 commonsourceibias.n469 commonsourceibias.n468 0.189894
R15537 commonsourceibias.n469 commonsourceibias.n447 0.189894
R15538 commonsourceibias.n473 commonsourceibias.n447 0.189894
R15539 commonsourceibias.n474 commonsourceibias.n473 0.189894
R15540 commonsourceibias.n474 commonsourceibias.n445 0.189894
R15541 commonsourceibias.n478 commonsourceibias.n445 0.189894
R15542 commonsourceibias.n479 commonsourceibias.n478 0.189894
R15543 commonsourceibias.n479 commonsourceibias.n443 0.189894
R15544 commonsourceibias.n484 commonsourceibias.n443 0.189894
R15545 commonsourceibias.n485 commonsourceibias.n484 0.189894
R15546 commonsourceibias.n486 commonsourceibias.n485 0.189894
R15547 commonsourceibias.n486 commonsourceibias.n441 0.189894
R15548 commonsourceibias.n492 commonsourceibias.n441 0.189894
R15549 commonsourceibias.n493 commonsourceibias.n492 0.189894
R15550 commonsourceibias.n494 commonsourceibias.n493 0.189894
R15551 commonsourceibias.n494 commonsourceibias.n439 0.189894
R15552 commonsourceibias.n499 commonsourceibias.n439 0.189894
R15553 commonsourceibias.n500 commonsourceibias.n499 0.189894
R15554 commonsourceibias.n501 commonsourceibias.n500 0.189894
R15555 commonsourceibias.n501 commonsourceibias.n437 0.189894
R15556 commonsourceibias.n507 commonsourceibias.n437 0.189894
R15557 commonsourceibias.n508 commonsourceibias.n507 0.189894
R15558 commonsourceibias.n509 commonsourceibias.n508 0.189894
R15559 commonsourceibias.n509 commonsourceibias.n435 0.189894
R15560 commonsourceibias.n514 commonsourceibias.n435 0.189894
R15561 commonsourceibias.n515 commonsourceibias.n514 0.189894
R15562 commonsourceibias.n516 commonsourceibias.n515 0.189894
R15563 commonsourceibias.n516 commonsourceibias.n433 0.189894
R15564 commonsourceibias.n397 commonsourceibias.n396 0.189894
R15565 commonsourceibias.n397 commonsourceibias.n392 0.189894
R15566 commonsourceibias.n402 commonsourceibias.n392 0.189894
R15567 commonsourceibias.n403 commonsourceibias.n402 0.189894
R15568 commonsourceibias.n404 commonsourceibias.n403 0.189894
R15569 commonsourceibias.n404 commonsourceibias.n390 0.189894
R15570 commonsourceibias.n409 commonsourceibias.n390 0.189894
R15571 commonsourceibias.n410 commonsourceibias.n409 0.189894
R15572 commonsourceibias.n410 commonsourceibias.n388 0.189894
R15573 commonsourceibias.n414 commonsourceibias.n388 0.189894
R15574 commonsourceibias.n415 commonsourceibias.n414 0.189894
R15575 commonsourceibias.n415 commonsourceibias.n386 0.189894
R15576 commonsourceibias.n419 commonsourceibias.n386 0.189894
R15577 commonsourceibias.n420 commonsourceibias.n419 0.189894
R15578 commonsourceibias.n420 commonsourceibias.n384 0.189894
R15579 commonsourceibias.n425 commonsourceibias.n384 0.189894
R15580 commonsourceibias.n532 commonsourceibias.n382 0.189894
R15581 commonsourceibias.n538 commonsourceibias.n382 0.189894
R15582 commonsourceibias.n539 commonsourceibias.n538 0.189894
R15583 commonsourceibias.n540 commonsourceibias.n539 0.189894
R15584 commonsourceibias.n540 commonsourceibias.n380 0.189894
R15585 commonsourceibias.n545 commonsourceibias.n380 0.189894
R15586 commonsourceibias.n546 commonsourceibias.n545 0.189894
R15587 commonsourceibias.n547 commonsourceibias.n546 0.189894
R15588 commonsourceibias.n547 commonsourceibias.n378 0.189894
R15589 commonsourceibias.n553 commonsourceibias.n378 0.189894
R15590 commonsourceibias.n554 commonsourceibias.n553 0.189894
R15591 commonsourceibias.n555 commonsourceibias.n554 0.189894
R15592 commonsourceibias.n555 commonsourceibias.n376 0.189894
R15593 commonsourceibias.n560 commonsourceibias.n376 0.189894
R15594 commonsourceibias.n561 commonsourceibias.n560 0.189894
R15595 commonsourceibias.n562 commonsourceibias.n561 0.189894
R15596 commonsourceibias.n562 commonsourceibias.n374 0.189894
R15597 commonsourceibias.n681 commonsourceibias.n680 0.189894
R15598 commonsourceibias.n681 commonsourceibias.n676 0.189894
R15599 commonsourceibias.n686 commonsourceibias.n676 0.189894
R15600 commonsourceibias.n687 commonsourceibias.n686 0.189894
R15601 commonsourceibias.n688 commonsourceibias.n687 0.189894
R15602 commonsourceibias.n688 commonsourceibias.n674 0.189894
R15603 commonsourceibias.n693 commonsourceibias.n674 0.189894
R15604 commonsourceibias.n694 commonsourceibias.n693 0.189894
R15605 commonsourceibias.n694 commonsourceibias.n672 0.189894
R15606 commonsourceibias.n698 commonsourceibias.n672 0.189894
R15607 commonsourceibias.n699 commonsourceibias.n698 0.189894
R15608 commonsourceibias.n699 commonsourceibias.n670 0.189894
R15609 commonsourceibias.n703 commonsourceibias.n670 0.189894
R15610 commonsourceibias.n704 commonsourceibias.n703 0.189894
R15611 commonsourceibias.n704 commonsourceibias.n668 0.189894
R15612 commonsourceibias.n709 commonsourceibias.n668 0.189894
R15613 commonsourceibias.n710 commonsourceibias.n709 0.189894
R15614 commonsourceibias.n711 commonsourceibias.n710 0.189894
R15615 commonsourceibias.n711 commonsourceibias.n666 0.189894
R15616 commonsourceibias.n717 commonsourceibias.n666 0.189894
R15617 commonsourceibias.n718 commonsourceibias.n717 0.189894
R15618 commonsourceibias.n719 commonsourceibias.n718 0.189894
R15619 commonsourceibias.n719 commonsourceibias.n664 0.189894
R15620 commonsourceibias.n724 commonsourceibias.n664 0.189894
R15621 commonsourceibias.n725 commonsourceibias.n724 0.189894
R15622 commonsourceibias.n726 commonsourceibias.n725 0.189894
R15623 commonsourceibias.n726 commonsourceibias.n662 0.189894
R15624 commonsourceibias.n732 commonsourceibias.n662 0.189894
R15625 commonsourceibias.n733 commonsourceibias.n732 0.189894
R15626 commonsourceibias.n734 commonsourceibias.n733 0.189894
R15627 commonsourceibias.n734 commonsourceibias.n660 0.189894
R15628 commonsourceibias.n739 commonsourceibias.n660 0.189894
R15629 commonsourceibias.n740 commonsourceibias.n739 0.189894
R15630 commonsourceibias.n741 commonsourceibias.n740 0.189894
R15631 commonsourceibias.n741 commonsourceibias.n658 0.189894
R15632 commonsourceibias.n591 commonsourceibias.n590 0.189894
R15633 commonsourceibias.n591 commonsourceibias.n586 0.189894
R15634 commonsourceibias.n596 commonsourceibias.n586 0.189894
R15635 commonsourceibias.n597 commonsourceibias.n596 0.189894
R15636 commonsourceibias.n598 commonsourceibias.n597 0.189894
R15637 commonsourceibias.n598 commonsourceibias.n584 0.189894
R15638 commonsourceibias.n603 commonsourceibias.n584 0.189894
R15639 commonsourceibias.n604 commonsourceibias.n603 0.189894
R15640 commonsourceibias.n604 commonsourceibias.n582 0.189894
R15641 commonsourceibias.n608 commonsourceibias.n582 0.189894
R15642 commonsourceibias.n609 commonsourceibias.n608 0.189894
R15643 commonsourceibias.n609 commonsourceibias.n580 0.189894
R15644 commonsourceibias.n613 commonsourceibias.n580 0.189894
R15645 commonsourceibias.n614 commonsourceibias.n613 0.189894
R15646 commonsourceibias.n614 commonsourceibias.n578 0.189894
R15647 commonsourceibias.n619 commonsourceibias.n578 0.189894
R15648 commonsourceibias.n620 commonsourceibias.n619 0.189894
R15649 commonsourceibias.n621 commonsourceibias.n620 0.189894
R15650 commonsourceibias.n621 commonsourceibias.n576 0.189894
R15651 commonsourceibias.n627 commonsourceibias.n576 0.189894
R15652 commonsourceibias.n628 commonsourceibias.n627 0.189894
R15653 commonsourceibias.n629 commonsourceibias.n628 0.189894
R15654 commonsourceibias.n629 commonsourceibias.n574 0.189894
R15655 commonsourceibias.n634 commonsourceibias.n574 0.189894
R15656 commonsourceibias.n635 commonsourceibias.n634 0.189894
R15657 commonsourceibias.n636 commonsourceibias.n635 0.189894
R15658 commonsourceibias.n636 commonsourceibias.n572 0.189894
R15659 commonsourceibias.n642 commonsourceibias.n572 0.189894
R15660 commonsourceibias.n643 commonsourceibias.n642 0.189894
R15661 commonsourceibias.n644 commonsourceibias.n643 0.189894
R15662 commonsourceibias.n644 commonsourceibias.n570 0.189894
R15663 commonsourceibias.n649 commonsourceibias.n570 0.189894
R15664 commonsourceibias.n650 commonsourceibias.n649 0.189894
R15665 commonsourceibias.n651 commonsourceibias.n650 0.189894
R15666 commonsourceibias.n651 commonsourceibias.n568 0.189894
R15667 commonsourceibias.n159 commonsourceibias.n158 0.170955
R15668 commonsourceibias.n160 commonsourceibias.n159 0.170955
R15669 commonsourceibias.n531 commonsourceibias.n425 0.170955
R15670 commonsourceibias.n532 commonsourceibias.n531 0.170955
R15671 CSoutput.n19 CSoutput.t161 184.661
R15672 CSoutput.n78 CSoutput.n77 165.8
R15673 CSoutput.n76 CSoutput.n0 165.8
R15674 CSoutput.n75 CSoutput.n74 165.8
R15675 CSoutput.n73 CSoutput.n72 165.8
R15676 CSoutput.n71 CSoutput.n2 165.8
R15677 CSoutput.n69 CSoutput.n68 165.8
R15678 CSoutput.n67 CSoutput.n3 165.8
R15679 CSoutput.n66 CSoutput.n65 165.8
R15680 CSoutput.n63 CSoutput.n4 165.8
R15681 CSoutput.n61 CSoutput.n60 165.8
R15682 CSoutput.n59 CSoutput.n5 165.8
R15683 CSoutput.n58 CSoutput.n57 165.8
R15684 CSoutput.n55 CSoutput.n6 165.8
R15685 CSoutput.n54 CSoutput.n53 165.8
R15686 CSoutput.n52 CSoutput.n51 165.8
R15687 CSoutput.n50 CSoutput.n8 165.8
R15688 CSoutput.n48 CSoutput.n47 165.8
R15689 CSoutput.n46 CSoutput.n9 165.8
R15690 CSoutput.n45 CSoutput.n44 165.8
R15691 CSoutput.n42 CSoutput.n10 165.8
R15692 CSoutput.n41 CSoutput.n40 165.8
R15693 CSoutput.n39 CSoutput.n38 165.8
R15694 CSoutput.n37 CSoutput.n12 165.8
R15695 CSoutput.n35 CSoutput.n34 165.8
R15696 CSoutput.n33 CSoutput.n13 165.8
R15697 CSoutput.n32 CSoutput.n31 165.8
R15698 CSoutput.n29 CSoutput.n14 165.8
R15699 CSoutput.n28 CSoutput.n27 165.8
R15700 CSoutput.n26 CSoutput.n25 165.8
R15701 CSoutput.n24 CSoutput.n16 165.8
R15702 CSoutput.n22 CSoutput.n21 165.8
R15703 CSoutput.n20 CSoutput.n17 165.8
R15704 CSoutput.n77 CSoutput.t163 162.194
R15705 CSoutput.n18 CSoutput.t158 120.501
R15706 CSoutput.n23 CSoutput.t152 120.501
R15707 CSoutput.n15 CSoutput.t147 120.501
R15708 CSoutput.n30 CSoutput.t159 120.501
R15709 CSoutput.n36 CSoutput.t160 120.501
R15710 CSoutput.n11 CSoutput.t149 120.501
R15711 CSoutput.n43 CSoutput.t145 120.501
R15712 CSoutput.n49 CSoutput.t162 120.501
R15713 CSoutput.n7 CSoutput.t153 120.501
R15714 CSoutput.n56 CSoutput.t155 120.501
R15715 CSoutput.n62 CSoutput.t164 120.501
R15716 CSoutput.n64 CSoutput.t156 120.501
R15717 CSoutput.n70 CSoutput.t157 120.501
R15718 CSoutput.n1 CSoutput.t150 120.501
R15719 CSoutput.n270 CSoutput.n268 103.469
R15720 CSoutput.n262 CSoutput.n260 103.469
R15721 CSoutput.n255 CSoutput.n253 103.469
R15722 CSoutput.n96 CSoutput.n94 103.469
R15723 CSoutput.n88 CSoutput.n86 103.469
R15724 CSoutput.n81 CSoutput.n79 103.469
R15725 CSoutput.n272 CSoutput.n271 103.111
R15726 CSoutput.n270 CSoutput.n269 103.111
R15727 CSoutput.n266 CSoutput.n265 103.111
R15728 CSoutput.n264 CSoutput.n263 103.111
R15729 CSoutput.n262 CSoutput.n261 103.111
R15730 CSoutput.n259 CSoutput.n258 103.111
R15731 CSoutput.n257 CSoutput.n256 103.111
R15732 CSoutput.n255 CSoutput.n254 103.111
R15733 CSoutput.n96 CSoutput.n95 103.111
R15734 CSoutput.n98 CSoutput.n97 103.111
R15735 CSoutput.n100 CSoutput.n99 103.111
R15736 CSoutput.n88 CSoutput.n87 103.111
R15737 CSoutput.n90 CSoutput.n89 103.111
R15738 CSoutput.n92 CSoutput.n91 103.111
R15739 CSoutput.n81 CSoutput.n80 103.111
R15740 CSoutput.n83 CSoutput.n82 103.111
R15741 CSoutput.n85 CSoutput.n84 103.111
R15742 CSoutput.n274 CSoutput.n273 103.111
R15743 CSoutput.n310 CSoutput.n308 81.5057
R15744 CSoutput.n294 CSoutput.n292 81.5057
R15745 CSoutput.n279 CSoutput.n277 81.5057
R15746 CSoutput.n358 CSoutput.n356 81.5057
R15747 CSoutput.n342 CSoutput.n340 81.5057
R15748 CSoutput.n327 CSoutput.n325 81.5057
R15749 CSoutput.n322 CSoutput.n321 80.9324
R15750 CSoutput.n320 CSoutput.n319 80.9324
R15751 CSoutput.n318 CSoutput.n317 80.9324
R15752 CSoutput.n316 CSoutput.n315 80.9324
R15753 CSoutput.n314 CSoutput.n313 80.9324
R15754 CSoutput.n312 CSoutput.n311 80.9324
R15755 CSoutput.n310 CSoutput.n309 80.9324
R15756 CSoutput.n306 CSoutput.n305 80.9324
R15757 CSoutput.n304 CSoutput.n303 80.9324
R15758 CSoutput.n302 CSoutput.n301 80.9324
R15759 CSoutput.n300 CSoutput.n299 80.9324
R15760 CSoutput.n298 CSoutput.n297 80.9324
R15761 CSoutput.n296 CSoutput.n295 80.9324
R15762 CSoutput.n294 CSoutput.n293 80.9324
R15763 CSoutput.n291 CSoutput.n290 80.9324
R15764 CSoutput.n289 CSoutput.n288 80.9324
R15765 CSoutput.n287 CSoutput.n286 80.9324
R15766 CSoutput.n285 CSoutput.n284 80.9324
R15767 CSoutput.n283 CSoutput.n282 80.9324
R15768 CSoutput.n281 CSoutput.n280 80.9324
R15769 CSoutput.n279 CSoutput.n278 80.9324
R15770 CSoutput.n358 CSoutput.n357 80.9324
R15771 CSoutput.n360 CSoutput.n359 80.9324
R15772 CSoutput.n362 CSoutput.n361 80.9324
R15773 CSoutput.n364 CSoutput.n363 80.9324
R15774 CSoutput.n366 CSoutput.n365 80.9324
R15775 CSoutput.n368 CSoutput.n367 80.9324
R15776 CSoutput.n370 CSoutput.n369 80.9324
R15777 CSoutput.n342 CSoutput.n341 80.9324
R15778 CSoutput.n344 CSoutput.n343 80.9324
R15779 CSoutput.n346 CSoutput.n345 80.9324
R15780 CSoutput.n348 CSoutput.n347 80.9324
R15781 CSoutput.n350 CSoutput.n349 80.9324
R15782 CSoutput.n352 CSoutput.n351 80.9324
R15783 CSoutput.n354 CSoutput.n353 80.9324
R15784 CSoutput.n327 CSoutput.n326 80.9324
R15785 CSoutput.n329 CSoutput.n328 80.9324
R15786 CSoutput.n331 CSoutput.n330 80.9324
R15787 CSoutput.n333 CSoutput.n332 80.9324
R15788 CSoutput.n335 CSoutput.n334 80.9324
R15789 CSoutput.n337 CSoutput.n336 80.9324
R15790 CSoutput.n339 CSoutput.n338 80.9324
R15791 CSoutput.n25 CSoutput.n24 48.1486
R15792 CSoutput.n69 CSoutput.n3 48.1486
R15793 CSoutput.n38 CSoutput.n37 48.1486
R15794 CSoutput.n42 CSoutput.n41 48.1486
R15795 CSoutput.n51 CSoutput.n50 48.1486
R15796 CSoutput.n55 CSoutput.n54 48.1486
R15797 CSoutput.n22 CSoutput.n17 46.462
R15798 CSoutput.n72 CSoutput.n71 46.462
R15799 CSoutput.n20 CSoutput.n19 44.9055
R15800 CSoutput.n29 CSoutput.n28 43.7635
R15801 CSoutput.n65 CSoutput.n63 43.7635
R15802 CSoutput.n35 CSoutput.n13 41.7396
R15803 CSoutput.n57 CSoutput.n5 41.7396
R15804 CSoutput.n44 CSoutput.n9 37.0171
R15805 CSoutput.n48 CSoutput.n9 37.0171
R15806 CSoutput.n76 CSoutput.n75 34.9932
R15807 CSoutput.n31 CSoutput.n13 32.2947
R15808 CSoutput.n61 CSoutput.n5 32.2947
R15809 CSoutput.n30 CSoutput.n29 29.6014
R15810 CSoutput.n63 CSoutput.n62 29.6014
R15811 CSoutput.n19 CSoutput.n18 28.4085
R15812 CSoutput.n18 CSoutput.n17 25.1176
R15813 CSoutput.n72 CSoutput.n1 25.1176
R15814 CSoutput.n43 CSoutput.n42 22.0922
R15815 CSoutput.n50 CSoutput.n49 22.0922
R15816 CSoutput.n77 CSoutput.n76 21.8586
R15817 CSoutput.n37 CSoutput.n36 18.9681
R15818 CSoutput.n56 CSoutput.n55 18.9681
R15819 CSoutput.n25 CSoutput.n15 17.6292
R15820 CSoutput.n64 CSoutput.n3 17.6292
R15821 CSoutput.n24 CSoutput.n23 15.844
R15822 CSoutput.n70 CSoutput.n69 15.844
R15823 CSoutput.n38 CSoutput.n11 14.5051
R15824 CSoutput.n54 CSoutput.n7 14.5051
R15825 CSoutput.n373 CSoutput.n78 11.4982
R15826 CSoutput.n41 CSoutput.n11 11.3811
R15827 CSoutput.n51 CSoutput.n7 11.3811
R15828 CSoutput.n23 CSoutput.n22 10.0422
R15829 CSoutput.n71 CSoutput.n70 10.0422
R15830 CSoutput.n267 CSoutput.n259 9.25285
R15831 CSoutput.n93 CSoutput.n85 9.25285
R15832 CSoutput.n307 CSoutput.n291 8.98182
R15833 CSoutput.n355 CSoutput.n339 8.98182
R15834 CSoutput.n324 CSoutput.n276 8.78291
R15835 CSoutput.n28 CSoutput.n15 8.25698
R15836 CSoutput.n65 CSoutput.n64 8.25698
R15837 CSoutput.n276 CSoutput.n275 7.12641
R15838 CSoutput.n102 CSoutput.n101 7.12641
R15839 CSoutput.n36 CSoutput.n35 6.91809
R15840 CSoutput.n57 CSoutput.n56 6.91809
R15841 CSoutput.n324 CSoutput.n323 6.02792
R15842 CSoutput.n372 CSoutput.n371 6.02792
R15843 CSoutput.n323 CSoutput.n322 5.25266
R15844 CSoutput.n307 CSoutput.n306 5.25266
R15845 CSoutput.n371 CSoutput.n370 5.25266
R15846 CSoutput.n355 CSoutput.n354 5.25266
R15847 CSoutput.n373 CSoutput.n102 5.19047
R15848 CSoutput.n275 CSoutput.n274 5.1449
R15849 CSoutput.n267 CSoutput.n266 5.1449
R15850 CSoutput.n101 CSoutput.n100 5.1449
R15851 CSoutput.n93 CSoutput.n92 5.1449
R15852 CSoutput.n193 CSoutput.n146 4.5005
R15853 CSoutput.n162 CSoutput.n146 4.5005
R15854 CSoutput.n157 CSoutput.n141 4.5005
R15855 CSoutput.n157 CSoutput.n143 4.5005
R15856 CSoutput.n157 CSoutput.n140 4.5005
R15857 CSoutput.n157 CSoutput.n144 4.5005
R15858 CSoutput.n157 CSoutput.n139 4.5005
R15859 CSoutput.n157 CSoutput.t165 4.5005
R15860 CSoutput.n157 CSoutput.n138 4.5005
R15861 CSoutput.n157 CSoutput.n145 4.5005
R15862 CSoutput.n157 CSoutput.n146 4.5005
R15863 CSoutput.n155 CSoutput.n141 4.5005
R15864 CSoutput.n155 CSoutput.n143 4.5005
R15865 CSoutput.n155 CSoutput.n140 4.5005
R15866 CSoutput.n155 CSoutput.n144 4.5005
R15867 CSoutput.n155 CSoutput.n139 4.5005
R15868 CSoutput.n155 CSoutput.t165 4.5005
R15869 CSoutput.n155 CSoutput.n138 4.5005
R15870 CSoutput.n155 CSoutput.n145 4.5005
R15871 CSoutput.n155 CSoutput.n146 4.5005
R15872 CSoutput.n154 CSoutput.n141 4.5005
R15873 CSoutput.n154 CSoutput.n143 4.5005
R15874 CSoutput.n154 CSoutput.n140 4.5005
R15875 CSoutput.n154 CSoutput.n144 4.5005
R15876 CSoutput.n154 CSoutput.n139 4.5005
R15877 CSoutput.n154 CSoutput.t165 4.5005
R15878 CSoutput.n154 CSoutput.n138 4.5005
R15879 CSoutput.n154 CSoutput.n145 4.5005
R15880 CSoutput.n154 CSoutput.n146 4.5005
R15881 CSoutput.n239 CSoutput.n141 4.5005
R15882 CSoutput.n239 CSoutput.n143 4.5005
R15883 CSoutput.n239 CSoutput.n140 4.5005
R15884 CSoutput.n239 CSoutput.n144 4.5005
R15885 CSoutput.n239 CSoutput.n139 4.5005
R15886 CSoutput.n239 CSoutput.t165 4.5005
R15887 CSoutput.n239 CSoutput.n138 4.5005
R15888 CSoutput.n239 CSoutput.n145 4.5005
R15889 CSoutput.n239 CSoutput.n146 4.5005
R15890 CSoutput.n237 CSoutput.n141 4.5005
R15891 CSoutput.n237 CSoutput.n143 4.5005
R15892 CSoutput.n237 CSoutput.n140 4.5005
R15893 CSoutput.n237 CSoutput.n144 4.5005
R15894 CSoutput.n237 CSoutput.n139 4.5005
R15895 CSoutput.n237 CSoutput.t165 4.5005
R15896 CSoutput.n237 CSoutput.n138 4.5005
R15897 CSoutput.n237 CSoutput.n145 4.5005
R15898 CSoutput.n235 CSoutput.n141 4.5005
R15899 CSoutput.n235 CSoutput.n143 4.5005
R15900 CSoutput.n235 CSoutput.n140 4.5005
R15901 CSoutput.n235 CSoutput.n144 4.5005
R15902 CSoutput.n235 CSoutput.n139 4.5005
R15903 CSoutput.n235 CSoutput.t165 4.5005
R15904 CSoutput.n235 CSoutput.n138 4.5005
R15905 CSoutput.n235 CSoutput.n145 4.5005
R15906 CSoutput.n165 CSoutput.n141 4.5005
R15907 CSoutput.n165 CSoutput.n143 4.5005
R15908 CSoutput.n165 CSoutput.n140 4.5005
R15909 CSoutput.n165 CSoutput.n144 4.5005
R15910 CSoutput.n165 CSoutput.n139 4.5005
R15911 CSoutput.n165 CSoutput.t165 4.5005
R15912 CSoutput.n165 CSoutput.n138 4.5005
R15913 CSoutput.n165 CSoutput.n145 4.5005
R15914 CSoutput.n165 CSoutput.n146 4.5005
R15915 CSoutput.n164 CSoutput.n141 4.5005
R15916 CSoutput.n164 CSoutput.n143 4.5005
R15917 CSoutput.n164 CSoutput.n140 4.5005
R15918 CSoutput.n164 CSoutput.n144 4.5005
R15919 CSoutput.n164 CSoutput.n139 4.5005
R15920 CSoutput.n164 CSoutput.t165 4.5005
R15921 CSoutput.n164 CSoutput.n138 4.5005
R15922 CSoutput.n164 CSoutput.n145 4.5005
R15923 CSoutput.n164 CSoutput.n146 4.5005
R15924 CSoutput.n168 CSoutput.n141 4.5005
R15925 CSoutput.n168 CSoutput.n143 4.5005
R15926 CSoutput.n168 CSoutput.n140 4.5005
R15927 CSoutput.n168 CSoutput.n144 4.5005
R15928 CSoutput.n168 CSoutput.n139 4.5005
R15929 CSoutput.n168 CSoutput.t165 4.5005
R15930 CSoutput.n168 CSoutput.n138 4.5005
R15931 CSoutput.n168 CSoutput.n145 4.5005
R15932 CSoutput.n168 CSoutput.n146 4.5005
R15933 CSoutput.n167 CSoutput.n141 4.5005
R15934 CSoutput.n167 CSoutput.n143 4.5005
R15935 CSoutput.n167 CSoutput.n140 4.5005
R15936 CSoutput.n167 CSoutput.n144 4.5005
R15937 CSoutput.n167 CSoutput.n139 4.5005
R15938 CSoutput.n167 CSoutput.t165 4.5005
R15939 CSoutput.n167 CSoutput.n138 4.5005
R15940 CSoutput.n167 CSoutput.n145 4.5005
R15941 CSoutput.n167 CSoutput.n146 4.5005
R15942 CSoutput.n150 CSoutput.n141 4.5005
R15943 CSoutput.n150 CSoutput.n143 4.5005
R15944 CSoutput.n150 CSoutput.n140 4.5005
R15945 CSoutput.n150 CSoutput.n144 4.5005
R15946 CSoutput.n150 CSoutput.n139 4.5005
R15947 CSoutput.n150 CSoutput.t165 4.5005
R15948 CSoutput.n150 CSoutput.n138 4.5005
R15949 CSoutput.n150 CSoutput.n145 4.5005
R15950 CSoutput.n150 CSoutput.n146 4.5005
R15951 CSoutput.n242 CSoutput.n141 4.5005
R15952 CSoutput.n242 CSoutput.n143 4.5005
R15953 CSoutput.n242 CSoutput.n140 4.5005
R15954 CSoutput.n242 CSoutput.n144 4.5005
R15955 CSoutput.n242 CSoutput.n139 4.5005
R15956 CSoutput.n242 CSoutput.t165 4.5005
R15957 CSoutput.n242 CSoutput.n138 4.5005
R15958 CSoutput.n242 CSoutput.n145 4.5005
R15959 CSoutput.n242 CSoutput.n146 4.5005
R15960 CSoutput.n229 CSoutput.n200 4.5005
R15961 CSoutput.n229 CSoutput.n206 4.5005
R15962 CSoutput.n187 CSoutput.n176 4.5005
R15963 CSoutput.n187 CSoutput.n178 4.5005
R15964 CSoutput.n187 CSoutput.n175 4.5005
R15965 CSoutput.n187 CSoutput.n179 4.5005
R15966 CSoutput.n187 CSoutput.n174 4.5005
R15967 CSoutput.n187 CSoutput.t144 4.5005
R15968 CSoutput.n187 CSoutput.n173 4.5005
R15969 CSoutput.n187 CSoutput.n180 4.5005
R15970 CSoutput.n229 CSoutput.n187 4.5005
R15971 CSoutput.n208 CSoutput.n176 4.5005
R15972 CSoutput.n208 CSoutput.n178 4.5005
R15973 CSoutput.n208 CSoutput.n175 4.5005
R15974 CSoutput.n208 CSoutput.n179 4.5005
R15975 CSoutput.n208 CSoutput.n174 4.5005
R15976 CSoutput.n208 CSoutput.t144 4.5005
R15977 CSoutput.n208 CSoutput.n173 4.5005
R15978 CSoutput.n208 CSoutput.n180 4.5005
R15979 CSoutput.n229 CSoutput.n208 4.5005
R15980 CSoutput.n186 CSoutput.n176 4.5005
R15981 CSoutput.n186 CSoutput.n178 4.5005
R15982 CSoutput.n186 CSoutput.n175 4.5005
R15983 CSoutput.n186 CSoutput.n179 4.5005
R15984 CSoutput.n186 CSoutput.n174 4.5005
R15985 CSoutput.n186 CSoutput.t144 4.5005
R15986 CSoutput.n186 CSoutput.n173 4.5005
R15987 CSoutput.n186 CSoutput.n180 4.5005
R15988 CSoutput.n229 CSoutput.n186 4.5005
R15989 CSoutput.n210 CSoutput.n176 4.5005
R15990 CSoutput.n210 CSoutput.n178 4.5005
R15991 CSoutput.n210 CSoutput.n175 4.5005
R15992 CSoutput.n210 CSoutput.n179 4.5005
R15993 CSoutput.n210 CSoutput.n174 4.5005
R15994 CSoutput.n210 CSoutput.t144 4.5005
R15995 CSoutput.n210 CSoutput.n173 4.5005
R15996 CSoutput.n210 CSoutput.n180 4.5005
R15997 CSoutput.n229 CSoutput.n210 4.5005
R15998 CSoutput.n176 CSoutput.n171 4.5005
R15999 CSoutput.n178 CSoutput.n171 4.5005
R16000 CSoutput.n175 CSoutput.n171 4.5005
R16001 CSoutput.n179 CSoutput.n171 4.5005
R16002 CSoutput.n174 CSoutput.n171 4.5005
R16003 CSoutput.t144 CSoutput.n171 4.5005
R16004 CSoutput.n173 CSoutput.n171 4.5005
R16005 CSoutput.n180 CSoutput.n171 4.5005
R16006 CSoutput.n232 CSoutput.n176 4.5005
R16007 CSoutput.n232 CSoutput.n178 4.5005
R16008 CSoutput.n232 CSoutput.n175 4.5005
R16009 CSoutput.n232 CSoutput.n179 4.5005
R16010 CSoutput.n232 CSoutput.n174 4.5005
R16011 CSoutput.n232 CSoutput.t144 4.5005
R16012 CSoutput.n232 CSoutput.n173 4.5005
R16013 CSoutput.n232 CSoutput.n180 4.5005
R16014 CSoutput.n230 CSoutput.n176 4.5005
R16015 CSoutput.n230 CSoutput.n178 4.5005
R16016 CSoutput.n230 CSoutput.n175 4.5005
R16017 CSoutput.n230 CSoutput.n179 4.5005
R16018 CSoutput.n230 CSoutput.n174 4.5005
R16019 CSoutput.n230 CSoutput.t144 4.5005
R16020 CSoutput.n230 CSoutput.n173 4.5005
R16021 CSoutput.n230 CSoutput.n180 4.5005
R16022 CSoutput.n230 CSoutput.n229 4.5005
R16023 CSoutput.n212 CSoutput.n176 4.5005
R16024 CSoutput.n212 CSoutput.n178 4.5005
R16025 CSoutput.n212 CSoutput.n175 4.5005
R16026 CSoutput.n212 CSoutput.n179 4.5005
R16027 CSoutput.n212 CSoutput.n174 4.5005
R16028 CSoutput.n212 CSoutput.t144 4.5005
R16029 CSoutput.n212 CSoutput.n173 4.5005
R16030 CSoutput.n212 CSoutput.n180 4.5005
R16031 CSoutput.n229 CSoutput.n212 4.5005
R16032 CSoutput.n184 CSoutput.n176 4.5005
R16033 CSoutput.n184 CSoutput.n178 4.5005
R16034 CSoutput.n184 CSoutput.n175 4.5005
R16035 CSoutput.n184 CSoutput.n179 4.5005
R16036 CSoutput.n184 CSoutput.n174 4.5005
R16037 CSoutput.n184 CSoutput.t144 4.5005
R16038 CSoutput.n184 CSoutput.n173 4.5005
R16039 CSoutput.n184 CSoutput.n180 4.5005
R16040 CSoutput.n229 CSoutput.n184 4.5005
R16041 CSoutput.n214 CSoutput.n176 4.5005
R16042 CSoutput.n214 CSoutput.n178 4.5005
R16043 CSoutput.n214 CSoutput.n175 4.5005
R16044 CSoutput.n214 CSoutput.n179 4.5005
R16045 CSoutput.n214 CSoutput.n174 4.5005
R16046 CSoutput.n214 CSoutput.t144 4.5005
R16047 CSoutput.n214 CSoutput.n173 4.5005
R16048 CSoutput.n214 CSoutput.n180 4.5005
R16049 CSoutput.n229 CSoutput.n214 4.5005
R16050 CSoutput.n183 CSoutput.n176 4.5005
R16051 CSoutput.n183 CSoutput.n178 4.5005
R16052 CSoutput.n183 CSoutput.n175 4.5005
R16053 CSoutput.n183 CSoutput.n179 4.5005
R16054 CSoutput.n183 CSoutput.n174 4.5005
R16055 CSoutput.n183 CSoutput.t144 4.5005
R16056 CSoutput.n183 CSoutput.n173 4.5005
R16057 CSoutput.n183 CSoutput.n180 4.5005
R16058 CSoutput.n229 CSoutput.n183 4.5005
R16059 CSoutput.n228 CSoutput.n176 4.5005
R16060 CSoutput.n228 CSoutput.n178 4.5005
R16061 CSoutput.n228 CSoutput.n175 4.5005
R16062 CSoutput.n228 CSoutput.n179 4.5005
R16063 CSoutput.n228 CSoutput.n174 4.5005
R16064 CSoutput.n228 CSoutput.t144 4.5005
R16065 CSoutput.n228 CSoutput.n173 4.5005
R16066 CSoutput.n228 CSoutput.n180 4.5005
R16067 CSoutput.n229 CSoutput.n228 4.5005
R16068 CSoutput.n227 CSoutput.n112 4.5005
R16069 CSoutput.n128 CSoutput.n112 4.5005
R16070 CSoutput.n123 CSoutput.n107 4.5005
R16071 CSoutput.n123 CSoutput.n109 4.5005
R16072 CSoutput.n123 CSoutput.n106 4.5005
R16073 CSoutput.n123 CSoutput.n110 4.5005
R16074 CSoutput.n123 CSoutput.n105 4.5005
R16075 CSoutput.n123 CSoutput.t151 4.5005
R16076 CSoutput.n123 CSoutput.n104 4.5005
R16077 CSoutput.n123 CSoutput.n111 4.5005
R16078 CSoutput.n123 CSoutput.n112 4.5005
R16079 CSoutput.n121 CSoutput.n107 4.5005
R16080 CSoutput.n121 CSoutput.n109 4.5005
R16081 CSoutput.n121 CSoutput.n106 4.5005
R16082 CSoutput.n121 CSoutput.n110 4.5005
R16083 CSoutput.n121 CSoutput.n105 4.5005
R16084 CSoutput.n121 CSoutput.t151 4.5005
R16085 CSoutput.n121 CSoutput.n104 4.5005
R16086 CSoutput.n121 CSoutput.n111 4.5005
R16087 CSoutput.n121 CSoutput.n112 4.5005
R16088 CSoutput.n120 CSoutput.n107 4.5005
R16089 CSoutput.n120 CSoutput.n109 4.5005
R16090 CSoutput.n120 CSoutput.n106 4.5005
R16091 CSoutput.n120 CSoutput.n110 4.5005
R16092 CSoutput.n120 CSoutput.n105 4.5005
R16093 CSoutput.n120 CSoutput.t151 4.5005
R16094 CSoutput.n120 CSoutput.n104 4.5005
R16095 CSoutput.n120 CSoutput.n111 4.5005
R16096 CSoutput.n120 CSoutput.n112 4.5005
R16097 CSoutput.n249 CSoutput.n107 4.5005
R16098 CSoutput.n249 CSoutput.n109 4.5005
R16099 CSoutput.n249 CSoutput.n106 4.5005
R16100 CSoutput.n249 CSoutput.n110 4.5005
R16101 CSoutput.n249 CSoutput.n105 4.5005
R16102 CSoutput.n249 CSoutput.t151 4.5005
R16103 CSoutput.n249 CSoutput.n104 4.5005
R16104 CSoutput.n249 CSoutput.n111 4.5005
R16105 CSoutput.n249 CSoutput.n112 4.5005
R16106 CSoutput.n247 CSoutput.n107 4.5005
R16107 CSoutput.n247 CSoutput.n109 4.5005
R16108 CSoutput.n247 CSoutput.n106 4.5005
R16109 CSoutput.n247 CSoutput.n110 4.5005
R16110 CSoutput.n247 CSoutput.n105 4.5005
R16111 CSoutput.n247 CSoutput.t151 4.5005
R16112 CSoutput.n247 CSoutput.n104 4.5005
R16113 CSoutput.n247 CSoutput.n111 4.5005
R16114 CSoutput.n245 CSoutput.n107 4.5005
R16115 CSoutput.n245 CSoutput.n109 4.5005
R16116 CSoutput.n245 CSoutput.n106 4.5005
R16117 CSoutput.n245 CSoutput.n110 4.5005
R16118 CSoutput.n245 CSoutput.n105 4.5005
R16119 CSoutput.n245 CSoutput.t151 4.5005
R16120 CSoutput.n245 CSoutput.n104 4.5005
R16121 CSoutput.n245 CSoutput.n111 4.5005
R16122 CSoutput.n131 CSoutput.n107 4.5005
R16123 CSoutput.n131 CSoutput.n109 4.5005
R16124 CSoutput.n131 CSoutput.n106 4.5005
R16125 CSoutput.n131 CSoutput.n110 4.5005
R16126 CSoutput.n131 CSoutput.n105 4.5005
R16127 CSoutput.n131 CSoutput.t151 4.5005
R16128 CSoutput.n131 CSoutput.n104 4.5005
R16129 CSoutput.n131 CSoutput.n111 4.5005
R16130 CSoutput.n131 CSoutput.n112 4.5005
R16131 CSoutput.n130 CSoutput.n107 4.5005
R16132 CSoutput.n130 CSoutput.n109 4.5005
R16133 CSoutput.n130 CSoutput.n106 4.5005
R16134 CSoutput.n130 CSoutput.n110 4.5005
R16135 CSoutput.n130 CSoutput.n105 4.5005
R16136 CSoutput.n130 CSoutput.t151 4.5005
R16137 CSoutput.n130 CSoutput.n104 4.5005
R16138 CSoutput.n130 CSoutput.n111 4.5005
R16139 CSoutput.n130 CSoutput.n112 4.5005
R16140 CSoutput.n134 CSoutput.n107 4.5005
R16141 CSoutput.n134 CSoutput.n109 4.5005
R16142 CSoutput.n134 CSoutput.n106 4.5005
R16143 CSoutput.n134 CSoutput.n110 4.5005
R16144 CSoutput.n134 CSoutput.n105 4.5005
R16145 CSoutput.n134 CSoutput.t151 4.5005
R16146 CSoutput.n134 CSoutput.n104 4.5005
R16147 CSoutput.n134 CSoutput.n111 4.5005
R16148 CSoutput.n134 CSoutput.n112 4.5005
R16149 CSoutput.n133 CSoutput.n107 4.5005
R16150 CSoutput.n133 CSoutput.n109 4.5005
R16151 CSoutput.n133 CSoutput.n106 4.5005
R16152 CSoutput.n133 CSoutput.n110 4.5005
R16153 CSoutput.n133 CSoutput.n105 4.5005
R16154 CSoutput.n133 CSoutput.t151 4.5005
R16155 CSoutput.n133 CSoutput.n104 4.5005
R16156 CSoutput.n133 CSoutput.n111 4.5005
R16157 CSoutput.n133 CSoutput.n112 4.5005
R16158 CSoutput.n116 CSoutput.n107 4.5005
R16159 CSoutput.n116 CSoutput.n109 4.5005
R16160 CSoutput.n116 CSoutput.n106 4.5005
R16161 CSoutput.n116 CSoutput.n110 4.5005
R16162 CSoutput.n116 CSoutput.n105 4.5005
R16163 CSoutput.n116 CSoutput.t151 4.5005
R16164 CSoutput.n116 CSoutput.n104 4.5005
R16165 CSoutput.n116 CSoutput.n111 4.5005
R16166 CSoutput.n116 CSoutput.n112 4.5005
R16167 CSoutput.n252 CSoutput.n107 4.5005
R16168 CSoutput.n252 CSoutput.n109 4.5005
R16169 CSoutput.n252 CSoutput.n106 4.5005
R16170 CSoutput.n252 CSoutput.n110 4.5005
R16171 CSoutput.n252 CSoutput.n105 4.5005
R16172 CSoutput.n252 CSoutput.t151 4.5005
R16173 CSoutput.n252 CSoutput.n104 4.5005
R16174 CSoutput.n252 CSoutput.n111 4.5005
R16175 CSoutput.n252 CSoutput.n112 4.5005
R16176 CSoutput.n275 CSoutput.n267 4.10845
R16177 CSoutput.n101 CSoutput.n93 4.10845
R16178 CSoutput.n273 CSoutput.t3 4.06363
R16179 CSoutput.n273 CSoutput.t22 4.06363
R16180 CSoutput.n271 CSoutput.t32 4.06363
R16181 CSoutput.n271 CSoutput.t9 4.06363
R16182 CSoutput.n269 CSoutput.t45 4.06363
R16183 CSoutput.n269 CSoutput.t26 4.06363
R16184 CSoutput.n268 CSoutput.t33 4.06363
R16185 CSoutput.n268 CSoutput.t34 4.06363
R16186 CSoutput.n265 CSoutput.t35 4.06363
R16187 CSoutput.n265 CSoutput.t16 4.06363
R16188 CSoutput.n263 CSoutput.t27 4.06363
R16189 CSoutput.n263 CSoutput.t0 4.06363
R16190 CSoutput.n261 CSoutput.t1 4.06363
R16191 CSoutput.n261 CSoutput.t20 4.06363
R16192 CSoutput.n260 CSoutput.t38 4.06363
R16193 CSoutput.n260 CSoutput.t39 4.06363
R16194 CSoutput.n258 CSoutput.t21 4.06363
R16195 CSoutput.n258 CSoutput.t29 4.06363
R16196 CSoutput.n256 CSoutput.t14 4.06363
R16197 CSoutput.n256 CSoutput.t8 4.06363
R16198 CSoutput.n254 CSoutput.t28 4.06363
R16199 CSoutput.n254 CSoutput.t40 4.06363
R16200 CSoutput.n253 CSoutput.t36 4.06363
R16201 CSoutput.n253 CSoutput.t23 4.06363
R16202 CSoutput.n94 CSoutput.t42 4.06363
R16203 CSoutput.n94 CSoutput.t25 4.06363
R16204 CSoutput.n95 CSoutput.t19 4.06363
R16205 CSoutput.n95 CSoutput.t43 4.06363
R16206 CSoutput.n97 CSoutput.t4 4.06363
R16207 CSoutput.n97 CSoutput.t24 4.06363
R16208 CSoutput.n99 CSoutput.t18 4.06363
R16209 CSoutput.n99 CSoutput.t17 4.06363
R16210 CSoutput.n86 CSoutput.t10 4.06363
R16211 CSoutput.n86 CSoutput.t44 4.06363
R16212 CSoutput.n87 CSoutput.t13 4.06363
R16213 CSoutput.n87 CSoutput.t11 4.06363
R16214 CSoutput.n89 CSoutput.t47 4.06363
R16215 CSoutput.n89 CSoutput.t5 4.06363
R16216 CSoutput.n91 CSoutput.t12 4.06363
R16217 CSoutput.n91 CSoutput.t31 4.06363
R16218 CSoutput.n79 CSoutput.t7 4.06363
R16219 CSoutput.n79 CSoutput.t46 4.06363
R16220 CSoutput.n80 CSoutput.t41 4.06363
R16221 CSoutput.n80 CSoutput.t37 4.06363
R16222 CSoutput.n82 CSoutput.t6 4.06363
R16223 CSoutput.n82 CSoutput.t15 4.06363
R16224 CSoutput.n84 CSoutput.t30 4.06363
R16225 CSoutput.n84 CSoutput.t2 4.06363
R16226 CSoutput.n44 CSoutput.n43 3.79402
R16227 CSoutput.n49 CSoutput.n48 3.79402
R16228 CSoutput.n323 CSoutput.n307 3.72967
R16229 CSoutput.n371 CSoutput.n355 3.72967
R16230 CSoutput.n373 CSoutput.n372 3.57343
R16231 CSoutput.n372 CSoutput.n324 3.08965
R16232 CSoutput.n321 CSoutput.t77 2.82907
R16233 CSoutput.n321 CSoutput.t67 2.82907
R16234 CSoutput.n319 CSoutput.t58 2.82907
R16235 CSoutput.n319 CSoutput.t128 2.82907
R16236 CSoutput.n317 CSoutput.t70 2.82907
R16237 CSoutput.n317 CSoutput.t74 2.82907
R16238 CSoutput.n315 CSoutput.t69 2.82907
R16239 CSoutput.n315 CSoutput.t143 2.82907
R16240 CSoutput.n313 CSoutput.t88 2.82907
R16241 CSoutput.n313 CSoutput.t61 2.82907
R16242 CSoutput.n311 CSoutput.t52 2.82907
R16243 CSoutput.n311 CSoutput.t117 2.82907
R16244 CSoutput.n309 CSoutput.t79 2.82907
R16245 CSoutput.n309 CSoutput.t83 2.82907
R16246 CSoutput.n308 CSoutput.t60 2.82907
R16247 CSoutput.n308 CSoutput.t132 2.82907
R16248 CSoutput.n305 CSoutput.t114 2.82907
R16249 CSoutput.n305 CSoutput.t95 2.82907
R16250 CSoutput.n303 CSoutput.t96 2.82907
R16251 CSoutput.n303 CSoutput.t102 2.82907
R16252 CSoutput.n301 CSoutput.t51 2.82907
R16253 CSoutput.n301 CSoutput.t115 2.82907
R16254 CSoutput.n299 CSoutput.t113 2.82907
R16255 CSoutput.n299 CSoutput.t94 2.82907
R16256 CSoutput.n297 CSoutput.t130 2.82907
R16257 CSoutput.n297 CSoutput.t49 2.82907
R16258 CSoutput.n295 CSoutput.t50 2.82907
R16259 CSoutput.n295 CSoutput.t122 2.82907
R16260 CSoutput.n293 CSoutput.t59 2.82907
R16261 CSoutput.n293 CSoutput.t129 2.82907
R16262 CSoutput.n292 CSoutput.t136 2.82907
R16263 CSoutput.n292 CSoutput.t48 2.82907
R16264 CSoutput.n290 CSoutput.t55 2.82907
R16265 CSoutput.n290 CSoutput.t78 2.82907
R16266 CSoutput.n288 CSoutput.t66 2.82907
R16267 CSoutput.n288 CSoutput.t91 2.82907
R16268 CSoutput.n286 CSoutput.t101 2.82907
R16269 CSoutput.n286 CSoutput.t111 2.82907
R16270 CSoutput.n284 CSoutput.t89 2.82907
R16271 CSoutput.n284 CSoutput.t131 2.82907
R16272 CSoutput.n282 CSoutput.t105 2.82907
R16273 CSoutput.n282 CSoutput.t82 2.82907
R16274 CSoutput.n280 CSoutput.t71 2.82907
R16275 CSoutput.n280 CSoutput.t90 2.82907
R16276 CSoutput.n278 CSoutput.t81 2.82907
R16277 CSoutput.n278 CSoutput.t86 2.82907
R16278 CSoutput.n277 CSoutput.t87 2.82907
R16279 CSoutput.n277 CSoutput.t140 2.82907
R16280 CSoutput.n356 CSoutput.t100 2.82907
R16281 CSoutput.n356 CSoutput.t125 2.82907
R16282 CSoutput.n357 CSoutput.t72 2.82907
R16283 CSoutput.n357 CSoutput.t85 2.82907
R16284 CSoutput.n359 CSoutput.t92 2.82907
R16285 CSoutput.n359 CSoutput.t106 2.82907
R16286 CSoutput.n361 CSoutput.t126 2.82907
R16287 CSoutput.n361 CSoutput.t97 2.82907
R16288 CSoutput.n363 CSoutput.t104 2.82907
R16289 CSoutput.n363 CSoutput.t137 2.82907
R16290 CSoutput.n365 CSoutput.t54 2.82907
R16291 CSoutput.n365 CSoutput.t75 2.82907
R16292 CSoutput.n367 CSoutput.t98 2.82907
R16293 CSoutput.n367 CSoutput.t120 2.82907
R16294 CSoutput.n369 CSoutput.t133 2.82907
R16295 CSoutput.n369 CSoutput.t62 2.82907
R16296 CSoutput.n340 CSoutput.t63 2.82907
R16297 CSoutput.n340 CSoutput.t56 2.82907
R16298 CSoutput.n341 CSoutput.t53 2.82907
R16299 CSoutput.n341 CSoutput.t141 2.82907
R16300 CSoutput.n343 CSoutput.t142 2.82907
R16301 CSoutput.n343 CSoutput.t64 2.82907
R16302 CSoutput.n345 CSoutput.t65 2.82907
R16303 CSoutput.n345 CSoutput.t107 2.82907
R16304 CSoutput.n347 CSoutput.t108 2.82907
R16305 CSoutput.n347 CSoutput.t135 2.82907
R16306 CSoutput.n349 CSoutput.t138 2.82907
R16307 CSoutput.n349 CSoutput.t127 2.82907
R16308 CSoutput.n351 CSoutput.t121 2.82907
R16309 CSoutput.n351 CSoutput.t109 2.82907
R16310 CSoutput.n353 CSoutput.t110 2.82907
R16311 CSoutput.n353 CSoutput.t139 2.82907
R16312 CSoutput.n325 CSoutput.t73 2.82907
R16313 CSoutput.n325 CSoutput.t116 2.82907
R16314 CSoutput.n326 CSoutput.t112 2.82907
R16315 CSoutput.n326 CSoutput.t93 2.82907
R16316 CSoutput.n328 CSoutput.t119 2.82907
R16317 CSoutput.n328 CSoutput.t84 2.82907
R16318 CSoutput.n330 CSoutput.t103 2.82907
R16319 CSoutput.n330 CSoutput.t134 2.82907
R16320 CSoutput.n332 CSoutput.t68 2.82907
R16321 CSoutput.n332 CSoutput.t118 2.82907
R16322 CSoutput.n334 CSoutput.t57 2.82907
R16323 CSoutput.n334 CSoutput.t124 2.82907
R16324 CSoutput.n336 CSoutput.t123 2.82907
R16325 CSoutput.n336 CSoutput.t80 2.82907
R16326 CSoutput.n338 CSoutput.t99 2.82907
R16327 CSoutput.n338 CSoutput.t76 2.82907
R16328 CSoutput.n276 CSoutput.n102 2.57547
R16329 CSoutput.n75 CSoutput.n1 2.45513
R16330 CSoutput.n193 CSoutput.n191 2.251
R16331 CSoutput.n193 CSoutput.n190 2.251
R16332 CSoutput.n193 CSoutput.n189 2.251
R16333 CSoutput.n193 CSoutput.n188 2.251
R16334 CSoutput.n162 CSoutput.n161 2.251
R16335 CSoutput.n162 CSoutput.n160 2.251
R16336 CSoutput.n162 CSoutput.n159 2.251
R16337 CSoutput.n162 CSoutput.n158 2.251
R16338 CSoutput.n235 CSoutput.n234 2.251
R16339 CSoutput.n200 CSoutput.n198 2.251
R16340 CSoutput.n200 CSoutput.n197 2.251
R16341 CSoutput.n200 CSoutput.n196 2.251
R16342 CSoutput.n218 CSoutput.n200 2.251
R16343 CSoutput.n206 CSoutput.n205 2.251
R16344 CSoutput.n206 CSoutput.n204 2.251
R16345 CSoutput.n206 CSoutput.n203 2.251
R16346 CSoutput.n206 CSoutput.n202 2.251
R16347 CSoutput.n232 CSoutput.n172 2.251
R16348 CSoutput.n227 CSoutput.n225 2.251
R16349 CSoutput.n227 CSoutput.n224 2.251
R16350 CSoutput.n227 CSoutput.n223 2.251
R16351 CSoutput.n227 CSoutput.n222 2.251
R16352 CSoutput.n128 CSoutput.n127 2.251
R16353 CSoutput.n128 CSoutput.n126 2.251
R16354 CSoutput.n128 CSoutput.n125 2.251
R16355 CSoutput.n128 CSoutput.n124 2.251
R16356 CSoutput.n245 CSoutput.n244 2.251
R16357 CSoutput.n162 CSoutput.n142 2.2505
R16358 CSoutput.n157 CSoutput.n142 2.2505
R16359 CSoutput.n155 CSoutput.n142 2.2505
R16360 CSoutput.n154 CSoutput.n142 2.2505
R16361 CSoutput.n239 CSoutput.n142 2.2505
R16362 CSoutput.n237 CSoutput.n142 2.2505
R16363 CSoutput.n235 CSoutput.n142 2.2505
R16364 CSoutput.n165 CSoutput.n142 2.2505
R16365 CSoutput.n164 CSoutput.n142 2.2505
R16366 CSoutput.n168 CSoutput.n142 2.2505
R16367 CSoutput.n167 CSoutput.n142 2.2505
R16368 CSoutput.n150 CSoutput.n142 2.2505
R16369 CSoutput.n242 CSoutput.n142 2.2505
R16370 CSoutput.n242 CSoutput.n241 2.2505
R16371 CSoutput.n206 CSoutput.n177 2.2505
R16372 CSoutput.n187 CSoutput.n177 2.2505
R16373 CSoutput.n208 CSoutput.n177 2.2505
R16374 CSoutput.n186 CSoutput.n177 2.2505
R16375 CSoutput.n210 CSoutput.n177 2.2505
R16376 CSoutput.n177 CSoutput.n171 2.2505
R16377 CSoutput.n232 CSoutput.n177 2.2505
R16378 CSoutput.n230 CSoutput.n177 2.2505
R16379 CSoutput.n212 CSoutput.n177 2.2505
R16380 CSoutput.n184 CSoutput.n177 2.2505
R16381 CSoutput.n214 CSoutput.n177 2.2505
R16382 CSoutput.n183 CSoutput.n177 2.2505
R16383 CSoutput.n228 CSoutput.n177 2.2505
R16384 CSoutput.n228 CSoutput.n181 2.2505
R16385 CSoutput.n128 CSoutput.n108 2.2505
R16386 CSoutput.n123 CSoutput.n108 2.2505
R16387 CSoutput.n121 CSoutput.n108 2.2505
R16388 CSoutput.n120 CSoutput.n108 2.2505
R16389 CSoutput.n249 CSoutput.n108 2.2505
R16390 CSoutput.n247 CSoutput.n108 2.2505
R16391 CSoutput.n245 CSoutput.n108 2.2505
R16392 CSoutput.n131 CSoutput.n108 2.2505
R16393 CSoutput.n130 CSoutput.n108 2.2505
R16394 CSoutput.n134 CSoutput.n108 2.2505
R16395 CSoutput.n133 CSoutput.n108 2.2505
R16396 CSoutput.n116 CSoutput.n108 2.2505
R16397 CSoutput.n252 CSoutput.n108 2.2505
R16398 CSoutput.n252 CSoutput.n251 2.2505
R16399 CSoutput.n170 CSoutput.n163 2.25024
R16400 CSoutput.n170 CSoutput.n156 2.25024
R16401 CSoutput.n238 CSoutput.n170 2.25024
R16402 CSoutput.n170 CSoutput.n166 2.25024
R16403 CSoutput.n170 CSoutput.n169 2.25024
R16404 CSoutput.n170 CSoutput.n137 2.25024
R16405 CSoutput.n220 CSoutput.n217 2.25024
R16406 CSoutput.n220 CSoutput.n216 2.25024
R16407 CSoutput.n220 CSoutput.n215 2.25024
R16408 CSoutput.n220 CSoutput.n182 2.25024
R16409 CSoutput.n220 CSoutput.n219 2.25024
R16410 CSoutput.n221 CSoutput.n220 2.25024
R16411 CSoutput.n136 CSoutput.n129 2.25024
R16412 CSoutput.n136 CSoutput.n122 2.25024
R16413 CSoutput.n248 CSoutput.n136 2.25024
R16414 CSoutput.n136 CSoutput.n132 2.25024
R16415 CSoutput.n136 CSoutput.n135 2.25024
R16416 CSoutput.n136 CSoutput.n103 2.25024
R16417 CSoutput.n237 CSoutput.n147 1.50111
R16418 CSoutput.n185 CSoutput.n171 1.50111
R16419 CSoutput.n247 CSoutput.n113 1.50111
R16420 CSoutput.n193 CSoutput.n192 1.501
R16421 CSoutput.n200 CSoutput.n199 1.501
R16422 CSoutput.n227 CSoutput.n226 1.501
R16423 CSoutput.n241 CSoutput.n152 1.12536
R16424 CSoutput.n241 CSoutput.n153 1.12536
R16425 CSoutput.n241 CSoutput.n240 1.12536
R16426 CSoutput.n201 CSoutput.n181 1.12536
R16427 CSoutput.n207 CSoutput.n181 1.12536
R16428 CSoutput.n209 CSoutput.n181 1.12536
R16429 CSoutput.n251 CSoutput.n118 1.12536
R16430 CSoutput.n251 CSoutput.n119 1.12536
R16431 CSoutput.n251 CSoutput.n250 1.12536
R16432 CSoutput.n241 CSoutput.n148 1.12536
R16433 CSoutput.n241 CSoutput.n149 1.12536
R16434 CSoutput.n241 CSoutput.n151 1.12536
R16435 CSoutput.n231 CSoutput.n181 1.12536
R16436 CSoutput.n211 CSoutput.n181 1.12536
R16437 CSoutput.n213 CSoutput.n181 1.12536
R16438 CSoutput.n251 CSoutput.n114 1.12536
R16439 CSoutput.n251 CSoutput.n115 1.12536
R16440 CSoutput.n251 CSoutput.n117 1.12536
R16441 CSoutput.n31 CSoutput.n30 0.669944
R16442 CSoutput.n62 CSoutput.n61 0.669944
R16443 CSoutput.n312 CSoutput.n310 0.573776
R16444 CSoutput.n314 CSoutput.n312 0.573776
R16445 CSoutput.n316 CSoutput.n314 0.573776
R16446 CSoutput.n318 CSoutput.n316 0.573776
R16447 CSoutput.n320 CSoutput.n318 0.573776
R16448 CSoutput.n322 CSoutput.n320 0.573776
R16449 CSoutput.n296 CSoutput.n294 0.573776
R16450 CSoutput.n298 CSoutput.n296 0.573776
R16451 CSoutput.n300 CSoutput.n298 0.573776
R16452 CSoutput.n302 CSoutput.n300 0.573776
R16453 CSoutput.n304 CSoutput.n302 0.573776
R16454 CSoutput.n306 CSoutput.n304 0.573776
R16455 CSoutput.n281 CSoutput.n279 0.573776
R16456 CSoutput.n283 CSoutput.n281 0.573776
R16457 CSoutput.n285 CSoutput.n283 0.573776
R16458 CSoutput.n287 CSoutput.n285 0.573776
R16459 CSoutput.n289 CSoutput.n287 0.573776
R16460 CSoutput.n291 CSoutput.n289 0.573776
R16461 CSoutput.n370 CSoutput.n368 0.573776
R16462 CSoutput.n368 CSoutput.n366 0.573776
R16463 CSoutput.n366 CSoutput.n364 0.573776
R16464 CSoutput.n364 CSoutput.n362 0.573776
R16465 CSoutput.n362 CSoutput.n360 0.573776
R16466 CSoutput.n360 CSoutput.n358 0.573776
R16467 CSoutput.n354 CSoutput.n352 0.573776
R16468 CSoutput.n352 CSoutput.n350 0.573776
R16469 CSoutput.n350 CSoutput.n348 0.573776
R16470 CSoutput.n348 CSoutput.n346 0.573776
R16471 CSoutput.n346 CSoutput.n344 0.573776
R16472 CSoutput.n344 CSoutput.n342 0.573776
R16473 CSoutput.n339 CSoutput.n337 0.573776
R16474 CSoutput.n337 CSoutput.n335 0.573776
R16475 CSoutput.n335 CSoutput.n333 0.573776
R16476 CSoutput.n333 CSoutput.n331 0.573776
R16477 CSoutput.n331 CSoutput.n329 0.573776
R16478 CSoutput.n329 CSoutput.n327 0.573776
R16479 CSoutput.n373 CSoutput.n252 0.53442
R16480 CSoutput.n272 CSoutput.n270 0.358259
R16481 CSoutput.n274 CSoutput.n272 0.358259
R16482 CSoutput.n264 CSoutput.n262 0.358259
R16483 CSoutput.n266 CSoutput.n264 0.358259
R16484 CSoutput.n257 CSoutput.n255 0.358259
R16485 CSoutput.n259 CSoutput.n257 0.358259
R16486 CSoutput.n100 CSoutput.n98 0.358259
R16487 CSoutput.n98 CSoutput.n96 0.358259
R16488 CSoutput.n92 CSoutput.n90 0.358259
R16489 CSoutput.n90 CSoutput.n88 0.358259
R16490 CSoutput.n85 CSoutput.n83 0.358259
R16491 CSoutput.n83 CSoutput.n81 0.358259
R16492 CSoutput.n21 CSoutput.n20 0.169105
R16493 CSoutput.n21 CSoutput.n16 0.169105
R16494 CSoutput.n26 CSoutput.n16 0.169105
R16495 CSoutput.n27 CSoutput.n26 0.169105
R16496 CSoutput.n27 CSoutput.n14 0.169105
R16497 CSoutput.n32 CSoutput.n14 0.169105
R16498 CSoutput.n33 CSoutput.n32 0.169105
R16499 CSoutput.n34 CSoutput.n33 0.169105
R16500 CSoutput.n34 CSoutput.n12 0.169105
R16501 CSoutput.n39 CSoutput.n12 0.169105
R16502 CSoutput.n40 CSoutput.n39 0.169105
R16503 CSoutput.n40 CSoutput.n10 0.169105
R16504 CSoutput.n45 CSoutput.n10 0.169105
R16505 CSoutput.n46 CSoutput.n45 0.169105
R16506 CSoutput.n47 CSoutput.n46 0.169105
R16507 CSoutput.n47 CSoutput.n8 0.169105
R16508 CSoutput.n52 CSoutput.n8 0.169105
R16509 CSoutput.n53 CSoutput.n52 0.169105
R16510 CSoutput.n53 CSoutput.n6 0.169105
R16511 CSoutput.n58 CSoutput.n6 0.169105
R16512 CSoutput.n59 CSoutput.n58 0.169105
R16513 CSoutput.n60 CSoutput.n59 0.169105
R16514 CSoutput.n60 CSoutput.n4 0.169105
R16515 CSoutput.n66 CSoutput.n4 0.169105
R16516 CSoutput.n67 CSoutput.n66 0.169105
R16517 CSoutput.n68 CSoutput.n67 0.169105
R16518 CSoutput.n68 CSoutput.n2 0.169105
R16519 CSoutput.n73 CSoutput.n2 0.169105
R16520 CSoutput.n74 CSoutput.n73 0.169105
R16521 CSoutput.n74 CSoutput.n0 0.169105
R16522 CSoutput.n78 CSoutput.n0 0.169105
R16523 CSoutput.n195 CSoutput.n194 0.0910737
R16524 CSoutput.n246 CSoutput.n243 0.0723685
R16525 CSoutput.n200 CSoutput.n195 0.0522944
R16526 CSoutput.n243 CSoutput.n242 0.0499135
R16527 CSoutput.n194 CSoutput.n193 0.0499135
R16528 CSoutput.n228 CSoutput.n227 0.0464294
R16529 CSoutput.n236 CSoutput.n233 0.0391444
R16530 CSoutput.n195 CSoutput.t154 0.023435
R16531 CSoutput.n243 CSoutput.t146 0.02262
R16532 CSoutput.n194 CSoutput.t148 0.02262
R16533 CSoutput CSoutput.n373 0.0052
R16534 CSoutput.n165 CSoutput.n148 0.00365111
R16535 CSoutput.n168 CSoutput.n149 0.00365111
R16536 CSoutput.n151 CSoutput.n150 0.00365111
R16537 CSoutput.n193 CSoutput.n152 0.00365111
R16538 CSoutput.n157 CSoutput.n153 0.00365111
R16539 CSoutput.n240 CSoutput.n154 0.00365111
R16540 CSoutput.n231 CSoutput.n230 0.00365111
R16541 CSoutput.n211 CSoutput.n184 0.00365111
R16542 CSoutput.n213 CSoutput.n183 0.00365111
R16543 CSoutput.n201 CSoutput.n200 0.00365111
R16544 CSoutput.n207 CSoutput.n187 0.00365111
R16545 CSoutput.n209 CSoutput.n186 0.00365111
R16546 CSoutput.n131 CSoutput.n114 0.00365111
R16547 CSoutput.n134 CSoutput.n115 0.00365111
R16548 CSoutput.n117 CSoutput.n116 0.00365111
R16549 CSoutput.n227 CSoutput.n118 0.00365111
R16550 CSoutput.n123 CSoutput.n119 0.00365111
R16551 CSoutput.n250 CSoutput.n120 0.00365111
R16552 CSoutput.n162 CSoutput.n152 0.00340054
R16553 CSoutput.n155 CSoutput.n153 0.00340054
R16554 CSoutput.n240 CSoutput.n239 0.00340054
R16555 CSoutput.n235 CSoutput.n148 0.00340054
R16556 CSoutput.n164 CSoutput.n149 0.00340054
R16557 CSoutput.n167 CSoutput.n151 0.00340054
R16558 CSoutput.n206 CSoutput.n201 0.00340054
R16559 CSoutput.n208 CSoutput.n207 0.00340054
R16560 CSoutput.n210 CSoutput.n209 0.00340054
R16561 CSoutput.n232 CSoutput.n231 0.00340054
R16562 CSoutput.n212 CSoutput.n211 0.00340054
R16563 CSoutput.n214 CSoutput.n213 0.00340054
R16564 CSoutput.n128 CSoutput.n118 0.00340054
R16565 CSoutput.n121 CSoutput.n119 0.00340054
R16566 CSoutput.n250 CSoutput.n249 0.00340054
R16567 CSoutput.n245 CSoutput.n114 0.00340054
R16568 CSoutput.n130 CSoutput.n115 0.00340054
R16569 CSoutput.n133 CSoutput.n117 0.00340054
R16570 CSoutput.n163 CSoutput.n157 0.00252698
R16571 CSoutput.n156 CSoutput.n154 0.00252698
R16572 CSoutput.n238 CSoutput.n237 0.00252698
R16573 CSoutput.n166 CSoutput.n164 0.00252698
R16574 CSoutput.n169 CSoutput.n167 0.00252698
R16575 CSoutput.n242 CSoutput.n137 0.00252698
R16576 CSoutput.n163 CSoutput.n162 0.00252698
R16577 CSoutput.n156 CSoutput.n155 0.00252698
R16578 CSoutput.n239 CSoutput.n238 0.00252698
R16579 CSoutput.n166 CSoutput.n165 0.00252698
R16580 CSoutput.n169 CSoutput.n168 0.00252698
R16581 CSoutput.n150 CSoutput.n137 0.00252698
R16582 CSoutput.n217 CSoutput.n187 0.00252698
R16583 CSoutput.n216 CSoutput.n186 0.00252698
R16584 CSoutput.n215 CSoutput.n171 0.00252698
R16585 CSoutput.n212 CSoutput.n182 0.00252698
R16586 CSoutput.n219 CSoutput.n214 0.00252698
R16587 CSoutput.n228 CSoutput.n221 0.00252698
R16588 CSoutput.n217 CSoutput.n206 0.00252698
R16589 CSoutput.n216 CSoutput.n208 0.00252698
R16590 CSoutput.n215 CSoutput.n210 0.00252698
R16591 CSoutput.n230 CSoutput.n182 0.00252698
R16592 CSoutput.n219 CSoutput.n184 0.00252698
R16593 CSoutput.n221 CSoutput.n183 0.00252698
R16594 CSoutput.n129 CSoutput.n123 0.00252698
R16595 CSoutput.n122 CSoutput.n120 0.00252698
R16596 CSoutput.n248 CSoutput.n247 0.00252698
R16597 CSoutput.n132 CSoutput.n130 0.00252698
R16598 CSoutput.n135 CSoutput.n133 0.00252698
R16599 CSoutput.n252 CSoutput.n103 0.00252698
R16600 CSoutput.n129 CSoutput.n128 0.00252698
R16601 CSoutput.n122 CSoutput.n121 0.00252698
R16602 CSoutput.n249 CSoutput.n248 0.00252698
R16603 CSoutput.n132 CSoutput.n131 0.00252698
R16604 CSoutput.n135 CSoutput.n134 0.00252698
R16605 CSoutput.n116 CSoutput.n103 0.00252698
R16606 CSoutput.n237 CSoutput.n236 0.0020275
R16607 CSoutput.n236 CSoutput.n235 0.0020275
R16608 CSoutput.n233 CSoutput.n171 0.0020275
R16609 CSoutput.n233 CSoutput.n232 0.0020275
R16610 CSoutput.n247 CSoutput.n246 0.0020275
R16611 CSoutput.n246 CSoutput.n245 0.0020275
R16612 CSoutput.n147 CSoutput.n146 0.00166668
R16613 CSoutput.n229 CSoutput.n185 0.00166668
R16614 CSoutput.n113 CSoutput.n112 0.00166668
R16615 CSoutput.n251 CSoutput.n113 0.00133328
R16616 CSoutput.n185 CSoutput.n181 0.00133328
R16617 CSoutput.n241 CSoutput.n147 0.00133328
R16618 CSoutput.n244 CSoutput.n136 0.001
R16619 CSoutput.n222 CSoutput.n136 0.001
R16620 CSoutput.n124 CSoutput.n104 0.001
R16621 CSoutput.n223 CSoutput.n104 0.001
R16622 CSoutput.n125 CSoutput.n105 0.001
R16623 CSoutput.n224 CSoutput.n105 0.001
R16624 CSoutput.n126 CSoutput.n106 0.001
R16625 CSoutput.n225 CSoutput.n106 0.001
R16626 CSoutput.n127 CSoutput.n107 0.001
R16627 CSoutput.n226 CSoutput.n107 0.001
R16628 CSoutput.n220 CSoutput.n172 0.001
R16629 CSoutput.n220 CSoutput.n218 0.001
R16630 CSoutput.n202 CSoutput.n173 0.001
R16631 CSoutput.n196 CSoutput.n173 0.001
R16632 CSoutput.n203 CSoutput.n174 0.001
R16633 CSoutput.n197 CSoutput.n174 0.001
R16634 CSoutput.n204 CSoutput.n175 0.001
R16635 CSoutput.n198 CSoutput.n175 0.001
R16636 CSoutput.n205 CSoutput.n176 0.001
R16637 CSoutput.n199 CSoutput.n176 0.001
R16638 CSoutput.n234 CSoutput.n170 0.001
R16639 CSoutput.n188 CSoutput.n170 0.001
R16640 CSoutput.n158 CSoutput.n138 0.001
R16641 CSoutput.n189 CSoutput.n138 0.001
R16642 CSoutput.n159 CSoutput.n139 0.001
R16643 CSoutput.n190 CSoutput.n139 0.001
R16644 CSoutput.n160 CSoutput.n140 0.001
R16645 CSoutput.n191 CSoutput.n140 0.001
R16646 CSoutput.n161 CSoutput.n141 0.001
R16647 CSoutput.n192 CSoutput.n141 0.001
R16648 CSoutput.n192 CSoutput.n142 0.001
R16649 CSoutput.n191 CSoutput.n143 0.001
R16650 CSoutput.n190 CSoutput.n144 0.001
R16651 CSoutput.n189 CSoutput.t165 0.001
R16652 CSoutput.n188 CSoutput.n145 0.001
R16653 CSoutput.n161 CSoutput.n143 0.001
R16654 CSoutput.n160 CSoutput.n144 0.001
R16655 CSoutput.n159 CSoutput.t165 0.001
R16656 CSoutput.n158 CSoutput.n145 0.001
R16657 CSoutput.n234 CSoutput.n146 0.001
R16658 CSoutput.n199 CSoutput.n177 0.001
R16659 CSoutput.n198 CSoutput.n178 0.001
R16660 CSoutput.n197 CSoutput.n179 0.001
R16661 CSoutput.n196 CSoutput.t144 0.001
R16662 CSoutput.n218 CSoutput.n180 0.001
R16663 CSoutput.n205 CSoutput.n178 0.001
R16664 CSoutput.n204 CSoutput.n179 0.001
R16665 CSoutput.n203 CSoutput.t144 0.001
R16666 CSoutput.n202 CSoutput.n180 0.001
R16667 CSoutput.n229 CSoutput.n172 0.001
R16668 CSoutput.n226 CSoutput.n108 0.001
R16669 CSoutput.n225 CSoutput.n109 0.001
R16670 CSoutput.n224 CSoutput.n110 0.001
R16671 CSoutput.n223 CSoutput.t151 0.001
R16672 CSoutput.n222 CSoutput.n111 0.001
R16673 CSoutput.n127 CSoutput.n109 0.001
R16674 CSoutput.n126 CSoutput.n110 0.001
R16675 CSoutput.n125 CSoutput.t151 0.001
R16676 CSoutput.n124 CSoutput.n111 0.001
R16677 CSoutput.n244 CSoutput.n112 0.001
R16678 a_n2982_13878.n125 a_n2982_13878.t94 512.366
R16679 a_n2982_13878.n115 a_n2982_13878.t83 512.366
R16680 a_n2982_13878.n126 a_n2982_13878.t72 512.366
R16681 a_n2982_13878.n123 a_n2982_13878.t102 512.366
R16682 a_n2982_13878.n116 a_n2982_13878.t91 512.366
R16683 a_n2982_13878.n124 a_n2982_13878.t90 512.366
R16684 a_n2982_13878.n121 a_n2982_13878.t98 512.366
R16685 a_n2982_13878.n117 a_n2982_13878.t81 512.366
R16686 a_n2982_13878.n122 a_n2982_13878.t82 512.366
R16687 a_n2982_13878.n119 a_n2982_13878.t85 512.366
R16688 a_n2982_13878.n118 a_n2982_13878.t95 512.366
R16689 a_n2982_13878.n120 a_n2982_13878.t111 512.366
R16690 a_n2982_13878.n31 a_n2982_13878.t110 538.698
R16691 a_n2982_13878.n134 a_n2982_13878.t87 512.366
R16692 a_n2982_13878.n133 a_n2982_13878.t92 512.366
R16693 a_n2982_13878.n86 a_n2982_13878.t80 512.366
R16694 a_n2982_13878.n132 a_n2982_13878.t97 512.366
R16695 a_n2982_13878.n131 a_n2982_13878.t106 512.366
R16696 a_n2982_13878.n87 a_n2982_13878.t107 512.366
R16697 a_n2982_13878.n130 a_n2982_13878.t74 512.366
R16698 a_n2982_13878.n129 a_n2982_13878.t89 512.366
R16699 a_n2982_13878.n88 a_n2982_13878.t77 512.366
R16700 a_n2982_13878.n128 a_n2982_13878.t84 512.366
R16701 a_n2982_13878.n33 a_n2982_13878.t15 538.699
R16702 a_n2982_13878.n135 a_n2982_13878.t31 512.366
R16703 a_n2982_13878.n83 a_n2982_13878.t25 512.366
R16704 a_n2982_13878.n38 a_n2982_13878.t37 538.698
R16705 a_n2982_13878.n153 a_n2982_13878.t55 512.366
R16706 a_n2982_13878.n152 a_n2982_13878.t39 512.366
R16707 a_n2982_13878.n84 a_n2982_13878.t33 512.366
R16708 a_n2982_13878.n151 a_n2982_13878.t21 512.366
R16709 a_n2982_13878.n150 a_n2982_13878.t53 512.366
R16710 a_n2982_13878.n85 a_n2982_13878.t47 512.366
R16711 a_n2982_13878.n149 a_n2982_13878.t41 512.366
R16712 a_n2982_13878.n148 a_n2982_13878.t45 512.366
R16713 a_n2982_13878.n19 a_n2982_13878.t17 538.698
R16714 a_n2982_13878.n108 a_n2982_13878.t59 512.366
R16715 a_n2982_13878.n97 a_n2982_13878.t27 512.366
R16716 a_n2982_13878.n109 a_n2982_13878.t61 512.366
R16717 a_n2982_13878.n96 a_n2982_13878.t43 512.366
R16718 a_n2982_13878.n110 a_n2982_13878.t51 512.366
R16719 a_n2982_13878.n111 a_n2982_13878.t19 512.366
R16720 a_n2982_13878.n95 a_n2982_13878.t57 512.366
R16721 a_n2982_13878.n112 a_n2982_13878.t35 512.366
R16722 a_n2982_13878.n94 a_n2982_13878.t49 512.366
R16723 a_n2982_13878.n113 a_n2982_13878.t29 512.366
R16724 a_n2982_13878.n25 a_n2982_13878.t109 538.698
R16725 a_n2982_13878.n102 a_n2982_13878.t78 512.366
R16726 a_n2982_13878.n101 a_n2982_13878.t79 512.366
R16727 a_n2982_13878.n103 a_n2982_13878.t104 512.366
R16728 a_n2982_13878.n100 a_n2982_13878.t105 512.366
R16729 a_n2982_13878.n104 a_n2982_13878.t76 512.366
R16730 a_n2982_13878.n105 a_n2982_13878.t100 512.366
R16731 a_n2982_13878.n99 a_n2982_13878.t101 512.366
R16732 a_n2982_13878.n106 a_n2982_13878.t73 512.366
R16733 a_n2982_13878.n98 a_n2982_13878.t86 512.366
R16734 a_n2982_13878.n107 a_n2982_13878.t96 512.366
R16735 a_n2982_13878.n5 a_n2982_13878.n82 70.1674
R16736 a_n2982_13878.n7 a_n2982_13878.n80 70.1674
R16737 a_n2982_13878.n9 a_n2982_13878.n78 70.1674
R16738 a_n2982_13878.n12 a_n2982_13878.n76 70.1674
R16739 a_n2982_13878.n58 a_n2982_13878.n26 70.5844
R16740 a_n2982_13878.n50 a_n2982_13878.n32 44.5605
R16741 a_n2982_13878.n148 a_n2982_13878.n50 21.3688
R16742 a_n2982_13878.n49 a_n2982_13878.n34 80.4688
R16743 a_n2982_13878.n49 a_n2982_13878.n149 0.365327
R16744 a_n2982_13878.n35 a_n2982_13878.n48 75.0448
R16745 a_n2982_13878.n47 a_n2982_13878.n35 70.1674
R16746 a_n2982_13878.n151 a_n2982_13878.n47 20.9683
R16747 a_n2982_13878.n37 a_n2982_13878.n46 70.3058
R16748 a_n2982_13878.n46 a_n2982_13878.n84 20.6913
R16749 a_n2982_13878.n45 a_n2982_13878.n37 75.3623
R16750 a_n2982_13878.n152 a_n2982_13878.n45 10.5784
R16751 a_n2982_13878.n36 a_n2982_13878.n38 44.7878
R16752 a_n2982_13878.n33 a_n2982_13878.n32 44.7878
R16753 a_n2982_13878.n33 a_n2982_13878.n135 14.1664
R16754 a_n2982_13878.n26 a_n2982_13878.n57 70.1674
R16755 a_n2982_13878.n57 a_n2982_13878.n88 20.9683
R16756 a_n2982_13878.n56 a_n2982_13878.n27 74.73
R16757 a_n2982_13878.n129 a_n2982_13878.n56 11.843
R16758 a_n2982_13878.n55 a_n2982_13878.n27 80.4688
R16759 a_n2982_13878.n55 a_n2982_13878.n130 0.365327
R16760 a_n2982_13878.n28 a_n2982_13878.n54 75.0448
R16761 a_n2982_13878.n53 a_n2982_13878.n28 70.1674
R16762 a_n2982_13878.n132 a_n2982_13878.n53 20.9683
R16763 a_n2982_13878.n30 a_n2982_13878.n52 70.3058
R16764 a_n2982_13878.n52 a_n2982_13878.n86 20.6913
R16765 a_n2982_13878.n51 a_n2982_13878.n30 75.3623
R16766 a_n2982_13878.n133 a_n2982_13878.n51 10.5784
R16767 a_n2982_13878.n29 a_n2982_13878.n31 44.7878
R16768 a_n2982_13878.n15 a_n2982_13878.n74 70.5844
R16769 a_n2982_13878.n21 a_n2982_13878.n66 70.5844
R16770 a_n2982_13878.n65 a_n2982_13878.n21 70.1674
R16771 a_n2982_13878.n65 a_n2982_13878.n98 20.9683
R16772 a_n2982_13878.n20 a_n2982_13878.n64 74.73
R16773 a_n2982_13878.n106 a_n2982_13878.n64 11.843
R16774 a_n2982_13878.n63 a_n2982_13878.n20 80.4688
R16775 a_n2982_13878.n63 a_n2982_13878.n99 0.365327
R16776 a_n2982_13878.n22 a_n2982_13878.n62 75.0448
R16777 a_n2982_13878.n61 a_n2982_13878.n22 70.1674
R16778 a_n2982_13878.n61 a_n2982_13878.n100 20.9683
R16779 a_n2982_13878.n23 a_n2982_13878.n60 70.3058
R16780 a_n2982_13878.n103 a_n2982_13878.n60 20.6913
R16781 a_n2982_13878.n59 a_n2982_13878.n23 75.3623
R16782 a_n2982_13878.n59 a_n2982_13878.n101 10.5784
R16783 a_n2982_13878.n25 a_n2982_13878.n24 44.7878
R16784 a_n2982_13878.n73 a_n2982_13878.n15 70.1674
R16785 a_n2982_13878.n73 a_n2982_13878.n94 20.9683
R16786 a_n2982_13878.n14 a_n2982_13878.n72 74.73
R16787 a_n2982_13878.n112 a_n2982_13878.n72 11.843
R16788 a_n2982_13878.n71 a_n2982_13878.n14 80.4688
R16789 a_n2982_13878.n71 a_n2982_13878.n95 0.365327
R16790 a_n2982_13878.n16 a_n2982_13878.n70 75.0448
R16791 a_n2982_13878.n69 a_n2982_13878.n16 70.1674
R16792 a_n2982_13878.n69 a_n2982_13878.n96 20.9683
R16793 a_n2982_13878.n17 a_n2982_13878.n68 70.3058
R16794 a_n2982_13878.n109 a_n2982_13878.n68 20.6913
R16795 a_n2982_13878.n67 a_n2982_13878.n17 75.3623
R16796 a_n2982_13878.n67 a_n2982_13878.n97 10.5784
R16797 a_n2982_13878.n19 a_n2982_13878.n18 44.7878
R16798 a_n2982_13878.n120 a_n2982_13878.n76 20.9683
R16799 a_n2982_13878.n75 a_n2982_13878.n13 75.0448
R16800 a_n2982_13878.n75 a_n2982_13878.n118 11.2134
R16801 a_n2982_13878.n13 a_n2982_13878.n119 161.3
R16802 a_n2982_13878.n122 a_n2982_13878.n78 20.9683
R16803 a_n2982_13878.n77 a_n2982_13878.n10 75.0448
R16804 a_n2982_13878.n77 a_n2982_13878.n117 11.2134
R16805 a_n2982_13878.n10 a_n2982_13878.n121 161.3
R16806 a_n2982_13878.n124 a_n2982_13878.n80 20.9683
R16807 a_n2982_13878.n79 a_n2982_13878.n8 75.0448
R16808 a_n2982_13878.n79 a_n2982_13878.n116 11.2134
R16809 a_n2982_13878.n8 a_n2982_13878.n123 161.3
R16810 a_n2982_13878.n126 a_n2982_13878.n82 20.9683
R16811 a_n2982_13878.n81 a_n2982_13878.n6 75.0448
R16812 a_n2982_13878.n81 a_n2982_13878.n115 11.2134
R16813 a_n2982_13878.n6 a_n2982_13878.n125 161.3
R16814 a_n2982_13878.n3 a_n2982_13878.n145 81.3764
R16815 a_n2982_13878.n4 a_n2982_13878.n139 81.3764
R16816 a_n2982_13878.n0 a_n2982_13878.n136 81.3764
R16817 a_n2982_13878.n3 a_n2982_13878.n146 80.9324
R16818 a_n2982_13878.n2 a_n2982_13878.n147 80.9324
R16819 a_n2982_13878.n2 a_n2982_13878.n144 80.9324
R16820 a_n2982_13878.n2 a_n2982_13878.n143 80.9324
R16821 a_n2982_13878.n1 a_n2982_13878.n142 80.9324
R16822 a_n2982_13878.n4 a_n2982_13878.n140 80.9324
R16823 a_n2982_13878.n0 a_n2982_13878.n141 80.9324
R16824 a_n2982_13878.n0 a_n2982_13878.n138 80.9324
R16825 a_n2982_13878.n0 a_n2982_13878.n137 80.9324
R16826 a_n2982_13878.n39 a_n2982_13878.t18 74.6477
R16827 a_n2982_13878.t16 a_n2982_13878.n44 74.6477
R16828 a_n2982_13878.n42 a_n2982_13878.t38 74.2899
R16829 a_n2982_13878.n41 a_n2982_13878.t24 74.2897
R16830 a_n2982_13878.n44 a_n2982_13878.n159 70.6783
R16831 a_n2982_13878.n44 a_n2982_13878.n158 70.6783
R16832 a_n2982_13878.n43 a_n2982_13878.n157 70.6783
R16833 a_n2982_13878.n43 a_n2982_13878.n156 70.6783
R16834 a_n2982_13878.n42 a_n2982_13878.n155 70.6783
R16835 a_n2982_13878.n41 a_n2982_13878.n93 70.6783
R16836 a_n2982_13878.n40 a_n2982_13878.n92 70.6783
R16837 a_n2982_13878.n40 a_n2982_13878.n91 70.6783
R16838 a_n2982_13878.n39 a_n2982_13878.n90 70.6783
R16839 a_n2982_13878.n39 a_n2982_13878.n89 70.6783
R16840 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R16841 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R16842 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R16843 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R16844 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R16845 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R16846 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R16847 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R16848 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R16849 a_n2982_13878.n53 a_n2982_13878.n131 20.9683
R16850 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R16851 a_n2982_13878.n128 a_n2982_13878.n57 20.9683
R16852 a_n2982_13878.n135 a_n2982_13878.n83 48.2005
R16853 a_n2982_13878.n153 a_n2982_13878.n152 48.2005
R16854 a_n2982_13878.n47 a_n2982_13878.n150 20.9683
R16855 a_n2982_13878.n149 a_n2982_13878.n85 48.2005
R16856 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R16857 a_n2982_13878.n110 a_n2982_13878.n69 20.9683
R16858 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R16859 a_n2982_13878.n113 a_n2982_13878.n73 20.9683
R16860 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R16861 a_n2982_13878.n104 a_n2982_13878.n61 20.9683
R16862 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R16863 a_n2982_13878.n107 a_n2982_13878.n65 20.9683
R16864 a_n2982_13878.n132 a_n2982_13878.n52 21.4216
R16865 a_n2982_13878.n151 a_n2982_13878.n46 21.4216
R16866 a_n2982_13878.n96 a_n2982_13878.n68 21.4216
R16867 a_n2982_13878.n100 a_n2982_13878.n60 21.4216
R16868 a_n2982_13878.n58 a_n2982_13878.t103 532.5
R16869 a_n2982_13878.t23 a_n2982_13878.n74 532.5
R16870 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R16871 a_n2982_13878.n1 a_n2982_13878.n0 32.6799
R16872 a_n2982_13878.n56 a_n2982_13878.n88 34.4824
R16873 a_n2982_13878.n50 a_n2982_13878.n83 20.5623
R16874 a_n2982_13878.n94 a_n2982_13878.n72 34.4824
R16875 a_n2982_13878.n98 a_n2982_13878.n64 34.4824
R16876 a_n2982_13878.n126 a_n2982_13878.n81 35.3134
R16877 a_n2982_13878.n124 a_n2982_13878.n79 35.3134
R16878 a_n2982_13878.n122 a_n2982_13878.n77 35.3134
R16879 a_n2982_13878.n120 a_n2982_13878.n75 35.3134
R16880 a_n2982_13878.n131 a_n2982_13878.n54 35.3134
R16881 a_n2982_13878.n54 a_n2982_13878.n87 11.2134
R16882 a_n2982_13878.n150 a_n2982_13878.n48 35.3134
R16883 a_n2982_13878.n48 a_n2982_13878.n85 11.2134
R16884 a_n2982_13878.n70 a_n2982_13878.n110 35.3134
R16885 a_n2982_13878.n111 a_n2982_13878.n70 11.2134
R16886 a_n2982_13878.n62 a_n2982_13878.n104 35.3134
R16887 a_n2982_13878.n105 a_n2982_13878.n62 11.2134
R16888 a_n2982_13878.n32 a_n2982_13878.n2 23.891
R16889 a_n2982_13878.n51 a_n2982_13878.n86 36.139
R16890 a_n2982_13878.n45 a_n2982_13878.n84 36.139
R16891 a_n2982_13878.n109 a_n2982_13878.n67 36.139
R16892 a_n2982_13878.n103 a_n2982_13878.n59 36.139
R16893 a_n2982_13878.n24 a_n2982_13878.n11 13.9285
R16894 a_n2982_13878.n26 a_n2982_13878.n127 13.724
R16895 a_n2982_13878.n154 a_n2982_13878.n36 12.4191
R16896 a_n2982_13878.n127 a_n2982_13878.n5 11.2486
R16897 a_n2982_13878.n13 a_n2982_13878.n11 11.2486
R16898 a_n2982_13878.n114 a_n2982_13878.n41 10.5745
R16899 a_n2982_13878.n114 a_n2982_13878.n15 8.58383
R16900 a_n2982_13878.n42 a_n2982_13878.n154 6.7311
R16901 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R16902 a_n2982_13878.n32 a_n2982_13878.n29 3.94368
R16903 a_n2982_13878.n18 a_n2982_13878.n21 3.94368
R16904 a_n2982_13878.n159 a_n2982_13878.t26 3.61217
R16905 a_n2982_13878.n159 a_n2982_13878.t32 3.61217
R16906 a_n2982_13878.n158 a_n2982_13878.t42 3.61217
R16907 a_n2982_13878.n158 a_n2982_13878.t46 3.61217
R16908 a_n2982_13878.n157 a_n2982_13878.t54 3.61217
R16909 a_n2982_13878.n157 a_n2982_13878.t48 3.61217
R16910 a_n2982_13878.n156 a_n2982_13878.t34 3.61217
R16911 a_n2982_13878.n156 a_n2982_13878.t22 3.61217
R16912 a_n2982_13878.n155 a_n2982_13878.t56 3.61217
R16913 a_n2982_13878.n155 a_n2982_13878.t40 3.61217
R16914 a_n2982_13878.n93 a_n2982_13878.t50 3.61217
R16915 a_n2982_13878.n93 a_n2982_13878.t30 3.61217
R16916 a_n2982_13878.n92 a_n2982_13878.t58 3.61217
R16917 a_n2982_13878.n92 a_n2982_13878.t36 3.61217
R16918 a_n2982_13878.n91 a_n2982_13878.t52 3.61217
R16919 a_n2982_13878.n91 a_n2982_13878.t20 3.61217
R16920 a_n2982_13878.n90 a_n2982_13878.t62 3.61217
R16921 a_n2982_13878.n90 a_n2982_13878.t44 3.61217
R16922 a_n2982_13878.n89 a_n2982_13878.t60 3.61217
R16923 a_n2982_13878.n89 a_n2982_13878.t28 3.61217
R16924 a_n2982_13878.n145 a_n2982_13878.t71 2.82907
R16925 a_n2982_13878.n145 a_n2982_13878.t4 2.82907
R16926 a_n2982_13878.n146 a_n2982_13878.t7 2.82907
R16927 a_n2982_13878.n146 a_n2982_13878.t0 2.82907
R16928 a_n2982_13878.n147 a_n2982_13878.t13 2.82907
R16929 a_n2982_13878.n147 a_n2982_13878.t64 2.82907
R16930 a_n2982_13878.n144 a_n2982_13878.t67 2.82907
R16931 a_n2982_13878.n144 a_n2982_13878.t6 2.82907
R16932 a_n2982_13878.n143 a_n2982_13878.t68 2.82907
R16933 a_n2982_13878.n143 a_n2982_13878.t65 2.82907
R16934 a_n2982_13878.n142 a_n2982_13878.t63 2.82907
R16935 a_n2982_13878.n142 a_n2982_13878.t2 2.82907
R16936 a_n2982_13878.n139 a_n2982_13878.t70 2.82907
R16937 a_n2982_13878.n139 a_n2982_13878.t11 2.82907
R16938 a_n2982_13878.n140 a_n2982_13878.t12 2.82907
R16939 a_n2982_13878.n140 a_n2982_13878.t8 2.82907
R16940 a_n2982_13878.n141 a_n2982_13878.t9 2.82907
R16941 a_n2982_13878.n141 a_n2982_13878.t5 2.82907
R16942 a_n2982_13878.n138 a_n2982_13878.t69 2.82907
R16943 a_n2982_13878.n138 a_n2982_13878.t10 2.82907
R16944 a_n2982_13878.n137 a_n2982_13878.t66 2.82907
R16945 a_n2982_13878.n137 a_n2982_13878.t3 2.82907
R16946 a_n2982_13878.n136 a_n2982_13878.t14 2.82907
R16947 a_n2982_13878.n136 a_n2982_13878.t1 2.82907
R16948 a_n2982_13878.n31 a_n2982_13878.n134 14.1668
R16949 a_n2982_13878.n128 a_n2982_13878.n58 22.3251
R16950 a_n2982_13878.n38 a_n2982_13878.n153 14.1668
R16951 a_n2982_13878.n108 a_n2982_13878.n19 14.1668
R16952 a_n2982_13878.n74 a_n2982_13878.n113 22.3251
R16953 a_n2982_13878.n102 a_n2982_13878.n25 14.1668
R16954 a_n2982_13878.n66 a_n2982_13878.n107 22.3251
R16955 a_n2982_13878.n154 a_n2982_13878.n11 1.30542
R16956 a_n2982_13878.n8 a_n2982_13878.n9 1.04595
R16957 a_n2982_13878.n55 a_n2982_13878.n129 47.835
R16958 a_n2982_13878.n49 a_n2982_13878.n148 47.835
R16959 a_n2982_13878.n112 a_n2982_13878.n71 47.835
R16960 a_n2982_13878.n106 a_n2982_13878.n63 47.835
R16961 a_n2982_13878.n0 a_n2982_13878.n4 1.3324
R16962 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R16963 a_n2982_13878.n21 a_n2982_13878.n20 1.13686
R16964 a_n2982_13878.n15 a_n2982_13878.n14 1.13686
R16965 a_n2982_13878.n32 a_n2982_13878.n34 1.09898
R16966 a_n2982_13878.n43 a_n2982_13878.n42 1.07378
R16967 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R16968 a_n2982_13878.n2 a_n2982_13878.n3 0.888431
R16969 a_n2982_13878.n2 a_n2982_13878.n1 0.888431
R16970 a_n2982_13878.n37 a_n2982_13878.n36 0.758076
R16971 a_n2982_13878.n37 a_n2982_13878.n35 0.758076
R16972 a_n2982_13878.n35 a_n2982_13878.n34 0.758076
R16973 a_n2982_13878.n30 a_n2982_13878.n29 0.758076
R16974 a_n2982_13878.n30 a_n2982_13878.n28 0.758076
R16975 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R16976 a_n2982_13878.n23 a_n2982_13878.n24 0.758076
R16977 a_n2982_13878.n22 a_n2982_13878.n23 0.758076
R16978 a_n2982_13878.n20 a_n2982_13878.n22 0.758076
R16979 a_n2982_13878.n17 a_n2982_13878.n18 0.758076
R16980 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R16981 a_n2982_13878.n14 a_n2982_13878.n16 0.758076
R16982 a_n2982_13878.n13 a_n2982_13878.n12 0.758076
R16983 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R16984 a_n2982_13878.n8 a_n2982_13878.n7 0.758076
R16985 a_n2982_13878.n6 a_n2982_13878.n5 0.758076
R16986 a_n2982_13878.n44 a_n2982_13878.n43 0.716017
R16987 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R16988 a_n2982_13878.n10 a_n2982_13878.n12 0.67853
R16989 a_n2982_13878.n6 a_n2982_13878.n7 0.67853
R16990 vdd.n291 vdd.n255 756.745
R16991 vdd.n244 vdd.n208 756.745
R16992 vdd.n201 vdd.n165 756.745
R16993 vdd.n154 vdd.n118 756.745
R16994 vdd.n112 vdd.n76 756.745
R16995 vdd.n65 vdd.n29 756.745
R16996 vdd.n1561 vdd.n1525 756.745
R16997 vdd.n1608 vdd.n1572 756.745
R16998 vdd.n1471 vdd.n1435 756.745
R16999 vdd.n1518 vdd.n1482 756.745
R17000 vdd.n1382 vdd.n1346 756.745
R17001 vdd.n1429 vdd.n1393 756.745
R17002 vdd.n1105 vdd.t20 640.208
R17003 vdd.n800 vdd.t65 640.208
R17004 vdd.n1109 vdd.t62 640.208
R17005 vdd.n791 vdd.t83 640.208
R17006 vdd.n686 vdd.t38 640.208
R17007 vdd.n2437 vdd.t80 640.208
R17008 vdd.n622 vdd.t31 640.208
R17009 vdd.n2434 vdd.t72 640.208
R17010 vdd.n589 vdd.t16 640.208
R17011 vdd.n861 vdd.t76 640.208
R17012 vdd.n1775 vdd.t53 592.009
R17013 vdd.n1813 vdd.t42 592.009
R17014 vdd.n1709 vdd.t56 592.009
R17015 vdd.n1976 vdd.t46 592.009
R17016 vdd.n1038 vdd.t24 592.009
R17017 vdd.n998 vdd.t28 592.009
R17018 vdd.n3180 vdd.t49 592.009
R17019 vdd.n405 vdd.t86 592.009
R17020 vdd.n365 vdd.t89 592.009
R17021 vdd.n557 vdd.t59 592.009
R17022 vdd.n3076 vdd.t69 592.009
R17023 vdd.n2983 vdd.t34 592.009
R17024 vdd.n292 vdd.n291 585
R17025 vdd.n290 vdd.n257 585
R17026 vdd.n289 vdd.n288 585
R17027 vdd.n260 vdd.n258 585
R17028 vdd.n283 vdd.n282 585
R17029 vdd.n281 vdd.n280 585
R17030 vdd.n264 vdd.n263 585
R17031 vdd.n275 vdd.n274 585
R17032 vdd.n273 vdd.n272 585
R17033 vdd.n268 vdd.n267 585
R17034 vdd.n245 vdd.n244 585
R17035 vdd.n243 vdd.n210 585
R17036 vdd.n242 vdd.n241 585
R17037 vdd.n213 vdd.n211 585
R17038 vdd.n236 vdd.n235 585
R17039 vdd.n234 vdd.n233 585
R17040 vdd.n217 vdd.n216 585
R17041 vdd.n228 vdd.n227 585
R17042 vdd.n226 vdd.n225 585
R17043 vdd.n221 vdd.n220 585
R17044 vdd.n202 vdd.n201 585
R17045 vdd.n200 vdd.n167 585
R17046 vdd.n199 vdd.n198 585
R17047 vdd.n170 vdd.n168 585
R17048 vdd.n193 vdd.n192 585
R17049 vdd.n191 vdd.n190 585
R17050 vdd.n174 vdd.n173 585
R17051 vdd.n185 vdd.n184 585
R17052 vdd.n183 vdd.n182 585
R17053 vdd.n178 vdd.n177 585
R17054 vdd.n155 vdd.n154 585
R17055 vdd.n153 vdd.n120 585
R17056 vdd.n152 vdd.n151 585
R17057 vdd.n123 vdd.n121 585
R17058 vdd.n146 vdd.n145 585
R17059 vdd.n144 vdd.n143 585
R17060 vdd.n127 vdd.n126 585
R17061 vdd.n138 vdd.n137 585
R17062 vdd.n136 vdd.n135 585
R17063 vdd.n131 vdd.n130 585
R17064 vdd.n113 vdd.n112 585
R17065 vdd.n111 vdd.n78 585
R17066 vdd.n110 vdd.n109 585
R17067 vdd.n81 vdd.n79 585
R17068 vdd.n104 vdd.n103 585
R17069 vdd.n102 vdd.n101 585
R17070 vdd.n85 vdd.n84 585
R17071 vdd.n96 vdd.n95 585
R17072 vdd.n94 vdd.n93 585
R17073 vdd.n89 vdd.n88 585
R17074 vdd.n66 vdd.n65 585
R17075 vdd.n64 vdd.n31 585
R17076 vdd.n63 vdd.n62 585
R17077 vdd.n34 vdd.n32 585
R17078 vdd.n57 vdd.n56 585
R17079 vdd.n55 vdd.n54 585
R17080 vdd.n38 vdd.n37 585
R17081 vdd.n49 vdd.n48 585
R17082 vdd.n47 vdd.n46 585
R17083 vdd.n42 vdd.n41 585
R17084 vdd.n1562 vdd.n1561 585
R17085 vdd.n1560 vdd.n1527 585
R17086 vdd.n1559 vdd.n1558 585
R17087 vdd.n1530 vdd.n1528 585
R17088 vdd.n1553 vdd.n1552 585
R17089 vdd.n1551 vdd.n1550 585
R17090 vdd.n1534 vdd.n1533 585
R17091 vdd.n1545 vdd.n1544 585
R17092 vdd.n1543 vdd.n1542 585
R17093 vdd.n1538 vdd.n1537 585
R17094 vdd.n1609 vdd.n1608 585
R17095 vdd.n1607 vdd.n1574 585
R17096 vdd.n1606 vdd.n1605 585
R17097 vdd.n1577 vdd.n1575 585
R17098 vdd.n1600 vdd.n1599 585
R17099 vdd.n1598 vdd.n1597 585
R17100 vdd.n1581 vdd.n1580 585
R17101 vdd.n1592 vdd.n1591 585
R17102 vdd.n1590 vdd.n1589 585
R17103 vdd.n1585 vdd.n1584 585
R17104 vdd.n1472 vdd.n1471 585
R17105 vdd.n1470 vdd.n1437 585
R17106 vdd.n1469 vdd.n1468 585
R17107 vdd.n1440 vdd.n1438 585
R17108 vdd.n1463 vdd.n1462 585
R17109 vdd.n1461 vdd.n1460 585
R17110 vdd.n1444 vdd.n1443 585
R17111 vdd.n1455 vdd.n1454 585
R17112 vdd.n1453 vdd.n1452 585
R17113 vdd.n1448 vdd.n1447 585
R17114 vdd.n1519 vdd.n1518 585
R17115 vdd.n1517 vdd.n1484 585
R17116 vdd.n1516 vdd.n1515 585
R17117 vdd.n1487 vdd.n1485 585
R17118 vdd.n1510 vdd.n1509 585
R17119 vdd.n1508 vdd.n1507 585
R17120 vdd.n1491 vdd.n1490 585
R17121 vdd.n1502 vdd.n1501 585
R17122 vdd.n1500 vdd.n1499 585
R17123 vdd.n1495 vdd.n1494 585
R17124 vdd.n1383 vdd.n1382 585
R17125 vdd.n1381 vdd.n1348 585
R17126 vdd.n1380 vdd.n1379 585
R17127 vdd.n1351 vdd.n1349 585
R17128 vdd.n1374 vdd.n1373 585
R17129 vdd.n1372 vdd.n1371 585
R17130 vdd.n1355 vdd.n1354 585
R17131 vdd.n1366 vdd.n1365 585
R17132 vdd.n1364 vdd.n1363 585
R17133 vdd.n1359 vdd.n1358 585
R17134 vdd.n1430 vdd.n1429 585
R17135 vdd.n1428 vdd.n1395 585
R17136 vdd.n1427 vdd.n1426 585
R17137 vdd.n1398 vdd.n1396 585
R17138 vdd.n1421 vdd.n1420 585
R17139 vdd.n1419 vdd.n1418 585
R17140 vdd.n1402 vdd.n1401 585
R17141 vdd.n1413 vdd.n1412 585
R17142 vdd.n1411 vdd.n1410 585
R17143 vdd.n1406 vdd.n1405 585
R17144 vdd.n3296 vdd.n330 515.122
R17145 vdd.n3178 vdd.n328 515.122
R17146 vdd.n515 vdd.n478 515.122
R17147 vdd.n3114 vdd.n479 515.122
R17148 vdd.n1971 vdd.n1320 515.122
R17149 vdd.n1974 vdd.n1973 515.122
R17150 vdd.n1682 vdd.n1646 515.122
R17151 vdd.n1878 vdd.n1647 515.122
R17152 vdd.n269 vdd.t145 329.043
R17153 vdd.n222 vdd.t153 329.043
R17154 vdd.n179 vdd.t142 329.043
R17155 vdd.n132 vdd.t150 329.043
R17156 vdd.n90 vdd.t122 329.043
R17157 vdd.n43 vdd.t127 329.043
R17158 vdd.n1539 vdd.t120 329.043
R17159 vdd.n1586 vdd.t106 329.043
R17160 vdd.n1449 vdd.t115 329.043
R17161 vdd.n1496 vdd.t95 329.043
R17162 vdd.n1360 vdd.t128 329.043
R17163 vdd.n1407 vdd.t123 329.043
R17164 vdd.n1775 vdd.t55 319.788
R17165 vdd.n1813 vdd.t45 319.788
R17166 vdd.n1709 vdd.t58 319.788
R17167 vdd.n1976 vdd.t47 319.788
R17168 vdd.n1038 vdd.t26 319.788
R17169 vdd.n998 vdd.t29 319.788
R17170 vdd.n3180 vdd.t51 319.788
R17171 vdd.n405 vdd.t87 319.788
R17172 vdd.n365 vdd.t90 319.788
R17173 vdd.n557 vdd.t61 319.788
R17174 vdd.n3076 vdd.t71 319.788
R17175 vdd.n2983 vdd.t37 319.788
R17176 vdd.n1776 vdd.t54 303.69
R17177 vdd.n1814 vdd.t44 303.69
R17178 vdd.n1710 vdd.t57 303.69
R17179 vdd.n1977 vdd.t48 303.69
R17180 vdd.n1039 vdd.t27 303.69
R17181 vdd.n999 vdd.t30 303.69
R17182 vdd.n3181 vdd.t52 303.69
R17183 vdd.n406 vdd.t88 303.69
R17184 vdd.n366 vdd.t91 303.69
R17185 vdd.n558 vdd.t60 303.69
R17186 vdd.n3077 vdd.t70 303.69
R17187 vdd.n2984 vdd.t36 303.69
R17188 vdd.n2704 vdd.n750 279.512
R17189 vdd.n2944 vdd.n599 279.512
R17190 vdd.n2881 vdd.n596 279.512
R17191 vdd.n2636 vdd.n2635 279.512
R17192 vdd.n2397 vdd.n788 279.512
R17193 vdd.n2328 vdd.n2327 279.512
R17194 vdd.n1145 vdd.n1144 279.512
R17195 vdd.n2122 vdd.n928 279.512
R17196 vdd.n2860 vdd.n597 279.512
R17197 vdd.n2947 vdd.n2946 279.512
R17198 vdd.n2509 vdd.n2432 279.512
R17199 vdd.n2440 vdd.n746 279.512
R17200 vdd.n2325 vdd.n798 279.512
R17201 vdd.n796 vdd.n770 279.512
R17202 vdd.n1270 vdd.n965 279.512
R17203 vdd.n1070 vdd.n923 279.512
R17204 vdd.n2120 vdd.n931 254.619
R17205 vdd.n3112 vdd.n484 254.619
R17206 vdd.n2862 vdd.n597 185
R17207 vdd.n2945 vdd.n597 185
R17208 vdd.n2864 vdd.n2863 185
R17209 vdd.n2863 vdd.n595 185
R17210 vdd.n2865 vdd.n629 185
R17211 vdd.n2875 vdd.n629 185
R17212 vdd.n2866 vdd.n638 185
R17213 vdd.n638 vdd.n636 185
R17214 vdd.n2868 vdd.n2867 185
R17215 vdd.n2869 vdd.n2868 185
R17216 vdd.n2821 vdd.n637 185
R17217 vdd.n637 vdd.n633 185
R17218 vdd.n2820 vdd.n2819 185
R17219 vdd.n2819 vdd.n2818 185
R17220 vdd.n640 vdd.n639 185
R17221 vdd.n641 vdd.n640 185
R17222 vdd.n2811 vdd.n2810 185
R17223 vdd.n2812 vdd.n2811 185
R17224 vdd.n2809 vdd.n649 185
R17225 vdd.n654 vdd.n649 185
R17226 vdd.n2808 vdd.n2807 185
R17227 vdd.n2807 vdd.n2806 185
R17228 vdd.n651 vdd.n650 185
R17229 vdd.n660 vdd.n651 185
R17230 vdd.n2799 vdd.n2798 185
R17231 vdd.n2800 vdd.n2799 185
R17232 vdd.n2797 vdd.n661 185
R17233 vdd.n667 vdd.n661 185
R17234 vdd.n2796 vdd.n2795 185
R17235 vdd.n2795 vdd.n2794 185
R17236 vdd.n663 vdd.n662 185
R17237 vdd.n664 vdd.n663 185
R17238 vdd.n2787 vdd.n2786 185
R17239 vdd.n2788 vdd.n2787 185
R17240 vdd.n2785 vdd.n674 185
R17241 vdd.n674 vdd.n671 185
R17242 vdd.n2784 vdd.n2783 185
R17243 vdd.n2783 vdd.n2782 185
R17244 vdd.n676 vdd.n675 185
R17245 vdd.n677 vdd.n676 185
R17246 vdd.n2775 vdd.n2774 185
R17247 vdd.n2776 vdd.n2775 185
R17248 vdd.n2773 vdd.n685 185
R17249 vdd.n691 vdd.n685 185
R17250 vdd.n2772 vdd.n2771 185
R17251 vdd.n2771 vdd.n2770 185
R17252 vdd.n2761 vdd.n688 185
R17253 vdd.n698 vdd.n688 185
R17254 vdd.n2763 vdd.n2762 185
R17255 vdd.n2764 vdd.n2763 185
R17256 vdd.n2760 vdd.n699 185
R17257 vdd.n699 vdd.n695 185
R17258 vdd.n2759 vdd.n2758 185
R17259 vdd.n2758 vdd.n2757 185
R17260 vdd.n701 vdd.n700 185
R17261 vdd.n702 vdd.n701 185
R17262 vdd.n2750 vdd.n2749 185
R17263 vdd.n2751 vdd.n2750 185
R17264 vdd.n2748 vdd.n710 185
R17265 vdd.n715 vdd.n710 185
R17266 vdd.n2747 vdd.n2746 185
R17267 vdd.n2746 vdd.n2745 185
R17268 vdd.n712 vdd.n711 185
R17269 vdd.n721 vdd.n712 185
R17270 vdd.n2738 vdd.n2737 185
R17271 vdd.n2739 vdd.n2738 185
R17272 vdd.n2736 vdd.n722 185
R17273 vdd.n2612 vdd.n722 185
R17274 vdd.n2735 vdd.n2734 185
R17275 vdd.n2734 vdd.n2733 185
R17276 vdd.n724 vdd.n723 185
R17277 vdd.n2618 vdd.n724 185
R17278 vdd.n2726 vdd.n2725 185
R17279 vdd.n2727 vdd.n2726 185
R17280 vdd.n2724 vdd.n733 185
R17281 vdd.n733 vdd.n730 185
R17282 vdd.n2723 vdd.n2722 185
R17283 vdd.n2722 vdd.n2721 185
R17284 vdd.n735 vdd.n734 185
R17285 vdd.n736 vdd.n735 185
R17286 vdd.n2714 vdd.n2713 185
R17287 vdd.n2715 vdd.n2714 185
R17288 vdd.n2712 vdd.n744 185
R17289 vdd.n2630 vdd.n744 185
R17290 vdd.n2711 vdd.n2710 185
R17291 vdd.n2710 vdd.n2709 185
R17292 vdd.n746 vdd.n745 185
R17293 vdd.n747 vdd.n746 185
R17294 vdd.n2441 vdd.n2440 185
R17295 vdd.n2443 vdd.n2442 185
R17296 vdd.n2445 vdd.n2444 185
R17297 vdd.n2447 vdd.n2446 185
R17298 vdd.n2449 vdd.n2448 185
R17299 vdd.n2451 vdd.n2450 185
R17300 vdd.n2453 vdd.n2452 185
R17301 vdd.n2455 vdd.n2454 185
R17302 vdd.n2457 vdd.n2456 185
R17303 vdd.n2459 vdd.n2458 185
R17304 vdd.n2461 vdd.n2460 185
R17305 vdd.n2463 vdd.n2462 185
R17306 vdd.n2465 vdd.n2464 185
R17307 vdd.n2467 vdd.n2466 185
R17308 vdd.n2469 vdd.n2468 185
R17309 vdd.n2471 vdd.n2470 185
R17310 vdd.n2473 vdd.n2472 185
R17311 vdd.n2475 vdd.n2474 185
R17312 vdd.n2477 vdd.n2476 185
R17313 vdd.n2479 vdd.n2478 185
R17314 vdd.n2481 vdd.n2480 185
R17315 vdd.n2483 vdd.n2482 185
R17316 vdd.n2485 vdd.n2484 185
R17317 vdd.n2487 vdd.n2486 185
R17318 vdd.n2489 vdd.n2488 185
R17319 vdd.n2491 vdd.n2490 185
R17320 vdd.n2493 vdd.n2492 185
R17321 vdd.n2495 vdd.n2494 185
R17322 vdd.n2497 vdd.n2496 185
R17323 vdd.n2499 vdd.n2498 185
R17324 vdd.n2501 vdd.n2500 185
R17325 vdd.n2503 vdd.n2502 185
R17326 vdd.n2505 vdd.n2504 185
R17327 vdd.n2507 vdd.n2506 185
R17328 vdd.n2508 vdd.n2432 185
R17329 vdd.n2702 vdd.n2432 185
R17330 vdd.n2948 vdd.n2947 185
R17331 vdd.n2949 vdd.n588 185
R17332 vdd.n2951 vdd.n2950 185
R17333 vdd.n2953 vdd.n586 185
R17334 vdd.n2955 vdd.n2954 185
R17335 vdd.n2956 vdd.n585 185
R17336 vdd.n2958 vdd.n2957 185
R17337 vdd.n2960 vdd.n583 185
R17338 vdd.n2962 vdd.n2961 185
R17339 vdd.n2963 vdd.n582 185
R17340 vdd.n2965 vdd.n2964 185
R17341 vdd.n2967 vdd.n580 185
R17342 vdd.n2969 vdd.n2968 185
R17343 vdd.n2970 vdd.n579 185
R17344 vdd.n2972 vdd.n2971 185
R17345 vdd.n2974 vdd.n578 185
R17346 vdd.n2975 vdd.n576 185
R17347 vdd.n2978 vdd.n2977 185
R17348 vdd.n577 vdd.n575 185
R17349 vdd.n2834 vdd.n2833 185
R17350 vdd.n2836 vdd.n2835 185
R17351 vdd.n2838 vdd.n2830 185
R17352 vdd.n2840 vdd.n2839 185
R17353 vdd.n2841 vdd.n2829 185
R17354 vdd.n2843 vdd.n2842 185
R17355 vdd.n2845 vdd.n2827 185
R17356 vdd.n2847 vdd.n2846 185
R17357 vdd.n2848 vdd.n2826 185
R17358 vdd.n2850 vdd.n2849 185
R17359 vdd.n2852 vdd.n2824 185
R17360 vdd.n2854 vdd.n2853 185
R17361 vdd.n2855 vdd.n2823 185
R17362 vdd.n2857 vdd.n2856 185
R17363 vdd.n2859 vdd.n2822 185
R17364 vdd.n2861 vdd.n2860 185
R17365 vdd.n2860 vdd.n484 185
R17366 vdd.n2946 vdd.n592 185
R17367 vdd.n2946 vdd.n2945 185
R17368 vdd.n2563 vdd.n594 185
R17369 vdd.n595 vdd.n594 185
R17370 vdd.n2564 vdd.n628 185
R17371 vdd.n2875 vdd.n628 185
R17372 vdd.n2566 vdd.n2565 185
R17373 vdd.n2565 vdd.n636 185
R17374 vdd.n2567 vdd.n635 185
R17375 vdd.n2869 vdd.n635 185
R17376 vdd.n2569 vdd.n2568 185
R17377 vdd.n2568 vdd.n633 185
R17378 vdd.n2570 vdd.n643 185
R17379 vdd.n2818 vdd.n643 185
R17380 vdd.n2572 vdd.n2571 185
R17381 vdd.n2571 vdd.n641 185
R17382 vdd.n2573 vdd.n648 185
R17383 vdd.n2812 vdd.n648 185
R17384 vdd.n2575 vdd.n2574 185
R17385 vdd.n2574 vdd.n654 185
R17386 vdd.n2576 vdd.n653 185
R17387 vdd.n2806 vdd.n653 185
R17388 vdd.n2578 vdd.n2577 185
R17389 vdd.n2577 vdd.n660 185
R17390 vdd.n2579 vdd.n659 185
R17391 vdd.n2800 vdd.n659 185
R17392 vdd.n2581 vdd.n2580 185
R17393 vdd.n2580 vdd.n667 185
R17394 vdd.n2582 vdd.n666 185
R17395 vdd.n2794 vdd.n666 185
R17396 vdd.n2584 vdd.n2583 185
R17397 vdd.n2583 vdd.n664 185
R17398 vdd.n2585 vdd.n673 185
R17399 vdd.n2788 vdd.n673 185
R17400 vdd.n2587 vdd.n2586 185
R17401 vdd.n2586 vdd.n671 185
R17402 vdd.n2588 vdd.n679 185
R17403 vdd.n2782 vdd.n679 185
R17404 vdd.n2590 vdd.n2589 185
R17405 vdd.n2589 vdd.n677 185
R17406 vdd.n2591 vdd.n684 185
R17407 vdd.n2776 vdd.n684 185
R17408 vdd.n2593 vdd.n2592 185
R17409 vdd.n2592 vdd.n691 185
R17410 vdd.n2594 vdd.n690 185
R17411 vdd.n2770 vdd.n690 185
R17412 vdd.n2596 vdd.n2595 185
R17413 vdd.n2595 vdd.n698 185
R17414 vdd.n2597 vdd.n697 185
R17415 vdd.n2764 vdd.n697 185
R17416 vdd.n2599 vdd.n2598 185
R17417 vdd.n2598 vdd.n695 185
R17418 vdd.n2600 vdd.n704 185
R17419 vdd.n2757 vdd.n704 185
R17420 vdd.n2602 vdd.n2601 185
R17421 vdd.n2601 vdd.n702 185
R17422 vdd.n2603 vdd.n709 185
R17423 vdd.n2751 vdd.n709 185
R17424 vdd.n2605 vdd.n2604 185
R17425 vdd.n2604 vdd.n715 185
R17426 vdd.n2606 vdd.n714 185
R17427 vdd.n2745 vdd.n714 185
R17428 vdd.n2608 vdd.n2607 185
R17429 vdd.n2607 vdd.n721 185
R17430 vdd.n2609 vdd.n720 185
R17431 vdd.n2739 vdd.n720 185
R17432 vdd.n2611 vdd.n2610 185
R17433 vdd.n2612 vdd.n2611 185
R17434 vdd.n2512 vdd.n726 185
R17435 vdd.n2733 vdd.n726 185
R17436 vdd.n2620 vdd.n2619 185
R17437 vdd.n2619 vdd.n2618 185
R17438 vdd.n2621 vdd.n732 185
R17439 vdd.n2727 vdd.n732 185
R17440 vdd.n2623 vdd.n2622 185
R17441 vdd.n2622 vdd.n730 185
R17442 vdd.n2624 vdd.n738 185
R17443 vdd.n2721 vdd.n738 185
R17444 vdd.n2626 vdd.n2625 185
R17445 vdd.n2625 vdd.n736 185
R17446 vdd.n2627 vdd.n743 185
R17447 vdd.n2715 vdd.n743 185
R17448 vdd.n2629 vdd.n2628 185
R17449 vdd.n2630 vdd.n2629 185
R17450 vdd.n2511 vdd.n749 185
R17451 vdd.n2709 vdd.n749 185
R17452 vdd.n2510 vdd.n2509 185
R17453 vdd.n2509 vdd.n747 185
R17454 vdd.n1971 vdd.n1970 185
R17455 vdd.n1972 vdd.n1971 185
R17456 vdd.n1321 vdd.n1319 185
R17457 vdd.n1963 vdd.n1319 185
R17458 vdd.n1966 vdd.n1965 185
R17459 vdd.n1965 vdd.n1964 185
R17460 vdd.n1324 vdd.n1323 185
R17461 vdd.n1325 vdd.n1324 185
R17462 vdd.n1952 vdd.n1951 185
R17463 vdd.n1953 vdd.n1952 185
R17464 vdd.n1333 vdd.n1332 185
R17465 vdd.n1944 vdd.n1332 185
R17466 vdd.n1947 vdd.n1946 185
R17467 vdd.n1946 vdd.n1945 185
R17468 vdd.n1336 vdd.n1335 185
R17469 vdd.n1343 vdd.n1336 185
R17470 vdd.n1935 vdd.n1934 185
R17471 vdd.n1936 vdd.n1935 185
R17472 vdd.n1345 vdd.n1344 185
R17473 vdd.n1344 vdd.n1342 185
R17474 vdd.n1930 vdd.n1929 185
R17475 vdd.n1929 vdd.n1928 185
R17476 vdd.n1618 vdd.n1617 185
R17477 vdd.n1619 vdd.n1618 185
R17478 vdd.n1919 vdd.n1918 185
R17479 vdd.n1920 vdd.n1919 185
R17480 vdd.n1626 vdd.n1625 185
R17481 vdd.n1910 vdd.n1625 185
R17482 vdd.n1913 vdd.n1912 185
R17483 vdd.n1912 vdd.n1911 185
R17484 vdd.n1629 vdd.n1628 185
R17485 vdd.n1635 vdd.n1629 185
R17486 vdd.n1901 vdd.n1900 185
R17487 vdd.n1902 vdd.n1901 185
R17488 vdd.n1637 vdd.n1636 185
R17489 vdd.n1893 vdd.n1636 185
R17490 vdd.n1896 vdd.n1895 185
R17491 vdd.n1895 vdd.n1894 185
R17492 vdd.n1640 vdd.n1639 185
R17493 vdd.n1641 vdd.n1640 185
R17494 vdd.n1884 vdd.n1883 185
R17495 vdd.n1885 vdd.n1884 185
R17496 vdd.n1648 vdd.n1647 185
R17497 vdd.n1683 vdd.n1647 185
R17498 vdd.n1879 vdd.n1878 185
R17499 vdd.n1651 vdd.n1650 185
R17500 vdd.n1875 vdd.n1874 185
R17501 vdd.n1876 vdd.n1875 185
R17502 vdd.n1685 vdd.n1684 185
R17503 vdd.n1870 vdd.n1687 185
R17504 vdd.n1869 vdd.n1688 185
R17505 vdd.n1868 vdd.n1689 185
R17506 vdd.n1691 vdd.n1690 185
R17507 vdd.n1864 vdd.n1693 185
R17508 vdd.n1863 vdd.n1694 185
R17509 vdd.n1862 vdd.n1695 185
R17510 vdd.n1697 vdd.n1696 185
R17511 vdd.n1858 vdd.n1699 185
R17512 vdd.n1857 vdd.n1700 185
R17513 vdd.n1856 vdd.n1701 185
R17514 vdd.n1703 vdd.n1702 185
R17515 vdd.n1852 vdd.n1705 185
R17516 vdd.n1851 vdd.n1706 185
R17517 vdd.n1850 vdd.n1707 185
R17518 vdd.n1711 vdd.n1708 185
R17519 vdd.n1846 vdd.n1713 185
R17520 vdd.n1845 vdd.n1714 185
R17521 vdd.n1844 vdd.n1715 185
R17522 vdd.n1717 vdd.n1716 185
R17523 vdd.n1840 vdd.n1719 185
R17524 vdd.n1839 vdd.n1720 185
R17525 vdd.n1838 vdd.n1721 185
R17526 vdd.n1723 vdd.n1722 185
R17527 vdd.n1834 vdd.n1725 185
R17528 vdd.n1833 vdd.n1726 185
R17529 vdd.n1832 vdd.n1727 185
R17530 vdd.n1729 vdd.n1728 185
R17531 vdd.n1828 vdd.n1731 185
R17532 vdd.n1827 vdd.n1732 185
R17533 vdd.n1826 vdd.n1733 185
R17534 vdd.n1735 vdd.n1734 185
R17535 vdd.n1822 vdd.n1737 185
R17536 vdd.n1821 vdd.n1738 185
R17537 vdd.n1820 vdd.n1739 185
R17538 vdd.n1741 vdd.n1740 185
R17539 vdd.n1816 vdd.n1743 185
R17540 vdd.n1815 vdd.n1812 185
R17541 vdd.n1811 vdd.n1744 185
R17542 vdd.n1746 vdd.n1745 185
R17543 vdd.n1807 vdd.n1748 185
R17544 vdd.n1806 vdd.n1749 185
R17545 vdd.n1805 vdd.n1750 185
R17546 vdd.n1752 vdd.n1751 185
R17547 vdd.n1801 vdd.n1754 185
R17548 vdd.n1800 vdd.n1755 185
R17549 vdd.n1799 vdd.n1756 185
R17550 vdd.n1758 vdd.n1757 185
R17551 vdd.n1795 vdd.n1760 185
R17552 vdd.n1794 vdd.n1761 185
R17553 vdd.n1793 vdd.n1762 185
R17554 vdd.n1764 vdd.n1763 185
R17555 vdd.n1789 vdd.n1766 185
R17556 vdd.n1788 vdd.n1767 185
R17557 vdd.n1787 vdd.n1768 185
R17558 vdd.n1770 vdd.n1769 185
R17559 vdd.n1783 vdd.n1772 185
R17560 vdd.n1782 vdd.n1773 185
R17561 vdd.n1781 vdd.n1774 185
R17562 vdd.n1778 vdd.n1682 185
R17563 vdd.n1876 vdd.n1682 185
R17564 vdd.n1975 vdd.n1974 185
R17565 vdd.n1979 vdd.n1315 185
R17566 vdd.n1314 vdd.n1308 185
R17567 vdd.n1312 vdd.n1311 185
R17568 vdd.n1310 vdd.n1069 185
R17569 vdd.n1983 vdd.n1066 185
R17570 vdd.n1985 vdd.n1984 185
R17571 vdd.n1987 vdd.n1064 185
R17572 vdd.n1989 vdd.n1988 185
R17573 vdd.n1990 vdd.n1059 185
R17574 vdd.n1992 vdd.n1991 185
R17575 vdd.n1994 vdd.n1057 185
R17576 vdd.n1996 vdd.n1995 185
R17577 vdd.n1997 vdd.n1052 185
R17578 vdd.n1999 vdd.n1998 185
R17579 vdd.n2001 vdd.n1050 185
R17580 vdd.n2003 vdd.n2002 185
R17581 vdd.n2004 vdd.n1046 185
R17582 vdd.n2006 vdd.n2005 185
R17583 vdd.n2008 vdd.n1043 185
R17584 vdd.n2010 vdd.n2009 185
R17585 vdd.n1044 vdd.n1037 185
R17586 vdd.n2014 vdd.n1041 185
R17587 vdd.n2015 vdd.n1033 185
R17588 vdd.n2017 vdd.n2016 185
R17589 vdd.n2019 vdd.n1031 185
R17590 vdd.n2021 vdd.n2020 185
R17591 vdd.n2022 vdd.n1026 185
R17592 vdd.n2024 vdd.n2023 185
R17593 vdd.n2026 vdd.n1024 185
R17594 vdd.n2028 vdd.n2027 185
R17595 vdd.n2029 vdd.n1019 185
R17596 vdd.n2031 vdd.n2030 185
R17597 vdd.n2033 vdd.n1017 185
R17598 vdd.n2035 vdd.n2034 185
R17599 vdd.n2036 vdd.n1012 185
R17600 vdd.n2038 vdd.n2037 185
R17601 vdd.n2040 vdd.n1010 185
R17602 vdd.n2042 vdd.n2041 185
R17603 vdd.n2043 vdd.n1006 185
R17604 vdd.n2045 vdd.n2044 185
R17605 vdd.n2047 vdd.n1003 185
R17606 vdd.n2049 vdd.n2048 185
R17607 vdd.n1004 vdd.n997 185
R17608 vdd.n2053 vdd.n1001 185
R17609 vdd.n2054 vdd.n993 185
R17610 vdd.n2056 vdd.n2055 185
R17611 vdd.n2058 vdd.n991 185
R17612 vdd.n2060 vdd.n2059 185
R17613 vdd.n2061 vdd.n986 185
R17614 vdd.n2063 vdd.n2062 185
R17615 vdd.n2065 vdd.n984 185
R17616 vdd.n2067 vdd.n2066 185
R17617 vdd.n2068 vdd.n979 185
R17618 vdd.n2070 vdd.n2069 185
R17619 vdd.n2072 vdd.n977 185
R17620 vdd.n2074 vdd.n2073 185
R17621 vdd.n2075 vdd.n975 185
R17622 vdd.n2077 vdd.n2076 185
R17623 vdd.n2080 vdd.n2079 185
R17624 vdd.n2082 vdd.n2081 185
R17625 vdd.n2084 vdd.n973 185
R17626 vdd.n2086 vdd.n2085 185
R17627 vdd.n1320 vdd.n972 185
R17628 vdd.n1973 vdd.n1318 185
R17629 vdd.n1973 vdd.n1972 185
R17630 vdd.n1328 vdd.n1317 185
R17631 vdd.n1963 vdd.n1317 185
R17632 vdd.n1962 vdd.n1961 185
R17633 vdd.n1964 vdd.n1962 185
R17634 vdd.n1327 vdd.n1326 185
R17635 vdd.n1326 vdd.n1325 185
R17636 vdd.n1955 vdd.n1954 185
R17637 vdd.n1954 vdd.n1953 185
R17638 vdd.n1331 vdd.n1330 185
R17639 vdd.n1944 vdd.n1331 185
R17640 vdd.n1943 vdd.n1942 185
R17641 vdd.n1945 vdd.n1943 185
R17642 vdd.n1338 vdd.n1337 185
R17643 vdd.n1343 vdd.n1337 185
R17644 vdd.n1938 vdd.n1937 185
R17645 vdd.n1937 vdd.n1936 185
R17646 vdd.n1341 vdd.n1340 185
R17647 vdd.n1342 vdd.n1341 185
R17648 vdd.n1927 vdd.n1926 185
R17649 vdd.n1928 vdd.n1927 185
R17650 vdd.n1621 vdd.n1620 185
R17651 vdd.n1620 vdd.n1619 185
R17652 vdd.n1922 vdd.n1921 185
R17653 vdd.n1921 vdd.n1920 185
R17654 vdd.n1624 vdd.n1623 185
R17655 vdd.n1910 vdd.n1624 185
R17656 vdd.n1909 vdd.n1908 185
R17657 vdd.n1911 vdd.n1909 185
R17658 vdd.n1631 vdd.n1630 185
R17659 vdd.n1635 vdd.n1630 185
R17660 vdd.n1904 vdd.n1903 185
R17661 vdd.n1903 vdd.n1902 185
R17662 vdd.n1634 vdd.n1633 185
R17663 vdd.n1893 vdd.n1634 185
R17664 vdd.n1892 vdd.n1891 185
R17665 vdd.n1894 vdd.n1892 185
R17666 vdd.n1643 vdd.n1642 185
R17667 vdd.n1642 vdd.n1641 185
R17668 vdd.n1887 vdd.n1886 185
R17669 vdd.n1886 vdd.n1885 185
R17670 vdd.n1646 vdd.n1645 185
R17671 vdd.n1683 vdd.n1646 185
R17672 vdd.n790 vdd.n788 185
R17673 vdd.n2326 vdd.n788 185
R17674 vdd.n2248 vdd.n808 185
R17675 vdd.n808 vdd.n795 185
R17676 vdd.n2250 vdd.n2249 185
R17677 vdd.n2251 vdd.n2250 185
R17678 vdd.n2247 vdd.n807 185
R17679 vdd.n1189 vdd.n807 185
R17680 vdd.n2246 vdd.n2245 185
R17681 vdd.n2245 vdd.n2244 185
R17682 vdd.n810 vdd.n809 185
R17683 vdd.n811 vdd.n810 185
R17684 vdd.n2235 vdd.n2234 185
R17685 vdd.n2236 vdd.n2235 185
R17686 vdd.n2233 vdd.n821 185
R17687 vdd.n821 vdd.n818 185
R17688 vdd.n2232 vdd.n2231 185
R17689 vdd.n2231 vdd.n2230 185
R17690 vdd.n823 vdd.n822 185
R17691 vdd.n1215 vdd.n823 185
R17692 vdd.n2223 vdd.n2222 185
R17693 vdd.n2224 vdd.n2223 185
R17694 vdd.n2221 vdd.n831 185
R17695 vdd.n836 vdd.n831 185
R17696 vdd.n2220 vdd.n2219 185
R17697 vdd.n2219 vdd.n2218 185
R17698 vdd.n833 vdd.n832 185
R17699 vdd.n842 vdd.n833 185
R17700 vdd.n2211 vdd.n2210 185
R17701 vdd.n2212 vdd.n2211 185
R17702 vdd.n2209 vdd.n843 185
R17703 vdd.n1227 vdd.n843 185
R17704 vdd.n2208 vdd.n2207 185
R17705 vdd.n2207 vdd.n2206 185
R17706 vdd.n845 vdd.n844 185
R17707 vdd.n846 vdd.n845 185
R17708 vdd.n2199 vdd.n2198 185
R17709 vdd.n2200 vdd.n2199 185
R17710 vdd.n2197 vdd.n855 185
R17711 vdd.n855 vdd.n852 185
R17712 vdd.n2196 vdd.n2195 185
R17713 vdd.n2195 vdd.n2194 185
R17714 vdd.n857 vdd.n856 185
R17715 vdd.n866 vdd.n857 185
R17716 vdd.n2186 vdd.n2185 185
R17717 vdd.n2187 vdd.n2186 185
R17718 vdd.n2184 vdd.n867 185
R17719 vdd.n873 vdd.n867 185
R17720 vdd.n2183 vdd.n2182 185
R17721 vdd.n2182 vdd.n2181 185
R17722 vdd.n869 vdd.n868 185
R17723 vdd.n870 vdd.n869 185
R17724 vdd.n2174 vdd.n2173 185
R17725 vdd.n2175 vdd.n2174 185
R17726 vdd.n2172 vdd.n880 185
R17727 vdd.n880 vdd.n877 185
R17728 vdd.n2171 vdd.n2170 185
R17729 vdd.n2170 vdd.n2169 185
R17730 vdd.n882 vdd.n881 185
R17731 vdd.n883 vdd.n882 185
R17732 vdd.n2162 vdd.n2161 185
R17733 vdd.n2163 vdd.n2162 185
R17734 vdd.n2160 vdd.n891 185
R17735 vdd.n896 vdd.n891 185
R17736 vdd.n2159 vdd.n2158 185
R17737 vdd.n2158 vdd.n2157 185
R17738 vdd.n893 vdd.n892 185
R17739 vdd.n902 vdd.n893 185
R17740 vdd.n2150 vdd.n2149 185
R17741 vdd.n2151 vdd.n2150 185
R17742 vdd.n2148 vdd.n903 185
R17743 vdd.n909 vdd.n903 185
R17744 vdd.n2147 vdd.n2146 185
R17745 vdd.n2146 vdd.n2145 185
R17746 vdd.n905 vdd.n904 185
R17747 vdd.n906 vdd.n905 185
R17748 vdd.n2138 vdd.n2137 185
R17749 vdd.n2139 vdd.n2138 185
R17750 vdd.n2136 vdd.n916 185
R17751 vdd.n916 vdd.n913 185
R17752 vdd.n2135 vdd.n2134 185
R17753 vdd.n2134 vdd.n2133 185
R17754 vdd.n918 vdd.n917 185
R17755 vdd.n927 vdd.n918 185
R17756 vdd.n2126 vdd.n2125 185
R17757 vdd.n2127 vdd.n2126 185
R17758 vdd.n2124 vdd.n928 185
R17759 vdd.n928 vdd.n924 185
R17760 vdd.n2123 vdd.n2122 185
R17761 vdd.n930 vdd.n929 185
R17762 vdd.n2119 vdd.n2118 185
R17763 vdd.n2120 vdd.n2119 185
R17764 vdd.n2117 vdd.n966 185
R17765 vdd.n2116 vdd.n2115 185
R17766 vdd.n2114 vdd.n2113 185
R17767 vdd.n2112 vdd.n2111 185
R17768 vdd.n2110 vdd.n2109 185
R17769 vdd.n2108 vdd.n2107 185
R17770 vdd.n2106 vdd.n2105 185
R17771 vdd.n2104 vdd.n2103 185
R17772 vdd.n2102 vdd.n2101 185
R17773 vdd.n2100 vdd.n2099 185
R17774 vdd.n2098 vdd.n2097 185
R17775 vdd.n2096 vdd.n2095 185
R17776 vdd.n2094 vdd.n2093 185
R17777 vdd.n2092 vdd.n2091 185
R17778 vdd.n2090 vdd.n2089 185
R17779 vdd.n1111 vdd.n967 185
R17780 vdd.n1113 vdd.n1112 185
R17781 vdd.n1115 vdd.n1114 185
R17782 vdd.n1117 vdd.n1116 185
R17783 vdd.n1119 vdd.n1118 185
R17784 vdd.n1121 vdd.n1120 185
R17785 vdd.n1123 vdd.n1122 185
R17786 vdd.n1125 vdd.n1124 185
R17787 vdd.n1127 vdd.n1126 185
R17788 vdd.n1129 vdd.n1128 185
R17789 vdd.n1131 vdd.n1130 185
R17790 vdd.n1133 vdd.n1132 185
R17791 vdd.n1135 vdd.n1134 185
R17792 vdd.n1137 vdd.n1136 185
R17793 vdd.n1140 vdd.n1139 185
R17794 vdd.n1142 vdd.n1141 185
R17795 vdd.n1144 vdd.n1143 185
R17796 vdd.n2329 vdd.n2328 185
R17797 vdd.n2331 vdd.n2330 185
R17798 vdd.n2333 vdd.n2332 185
R17799 vdd.n2336 vdd.n2335 185
R17800 vdd.n2338 vdd.n2337 185
R17801 vdd.n2340 vdd.n2339 185
R17802 vdd.n2342 vdd.n2341 185
R17803 vdd.n2344 vdd.n2343 185
R17804 vdd.n2346 vdd.n2345 185
R17805 vdd.n2348 vdd.n2347 185
R17806 vdd.n2350 vdd.n2349 185
R17807 vdd.n2352 vdd.n2351 185
R17808 vdd.n2354 vdd.n2353 185
R17809 vdd.n2356 vdd.n2355 185
R17810 vdd.n2358 vdd.n2357 185
R17811 vdd.n2360 vdd.n2359 185
R17812 vdd.n2362 vdd.n2361 185
R17813 vdd.n2364 vdd.n2363 185
R17814 vdd.n2366 vdd.n2365 185
R17815 vdd.n2368 vdd.n2367 185
R17816 vdd.n2370 vdd.n2369 185
R17817 vdd.n2372 vdd.n2371 185
R17818 vdd.n2374 vdd.n2373 185
R17819 vdd.n2376 vdd.n2375 185
R17820 vdd.n2378 vdd.n2377 185
R17821 vdd.n2380 vdd.n2379 185
R17822 vdd.n2382 vdd.n2381 185
R17823 vdd.n2384 vdd.n2383 185
R17824 vdd.n2386 vdd.n2385 185
R17825 vdd.n2388 vdd.n2387 185
R17826 vdd.n2390 vdd.n2389 185
R17827 vdd.n2392 vdd.n2391 185
R17828 vdd.n2394 vdd.n2393 185
R17829 vdd.n2395 vdd.n789 185
R17830 vdd.n2397 vdd.n2396 185
R17831 vdd.n2398 vdd.n2397 185
R17832 vdd.n2327 vdd.n793 185
R17833 vdd.n2327 vdd.n2326 185
R17834 vdd.n1187 vdd.n794 185
R17835 vdd.n795 vdd.n794 185
R17836 vdd.n1188 vdd.n805 185
R17837 vdd.n2251 vdd.n805 185
R17838 vdd.n1191 vdd.n1190 185
R17839 vdd.n1190 vdd.n1189 185
R17840 vdd.n1192 vdd.n812 185
R17841 vdd.n2244 vdd.n812 185
R17842 vdd.n1194 vdd.n1193 185
R17843 vdd.n1193 vdd.n811 185
R17844 vdd.n1195 vdd.n819 185
R17845 vdd.n2236 vdd.n819 185
R17846 vdd.n1197 vdd.n1196 185
R17847 vdd.n1196 vdd.n818 185
R17848 vdd.n1198 vdd.n824 185
R17849 vdd.n2230 vdd.n824 185
R17850 vdd.n1217 vdd.n1216 185
R17851 vdd.n1216 vdd.n1215 185
R17852 vdd.n1218 vdd.n829 185
R17853 vdd.n2224 vdd.n829 185
R17854 vdd.n1220 vdd.n1219 185
R17855 vdd.n1219 vdd.n836 185
R17856 vdd.n1221 vdd.n834 185
R17857 vdd.n2218 vdd.n834 185
R17858 vdd.n1223 vdd.n1222 185
R17859 vdd.n1222 vdd.n842 185
R17860 vdd.n1224 vdd.n840 185
R17861 vdd.n2212 vdd.n840 185
R17862 vdd.n1226 vdd.n1225 185
R17863 vdd.n1227 vdd.n1226 185
R17864 vdd.n1186 vdd.n847 185
R17865 vdd.n2206 vdd.n847 185
R17866 vdd.n1185 vdd.n1184 185
R17867 vdd.n1184 vdd.n846 185
R17868 vdd.n1183 vdd.n853 185
R17869 vdd.n2200 vdd.n853 185
R17870 vdd.n1182 vdd.n1181 185
R17871 vdd.n1181 vdd.n852 185
R17872 vdd.n1180 vdd.n858 185
R17873 vdd.n2194 vdd.n858 185
R17874 vdd.n1179 vdd.n1178 185
R17875 vdd.n1178 vdd.n866 185
R17876 vdd.n1177 vdd.n864 185
R17877 vdd.n2187 vdd.n864 185
R17878 vdd.n1176 vdd.n1175 185
R17879 vdd.n1175 vdd.n873 185
R17880 vdd.n1174 vdd.n871 185
R17881 vdd.n2181 vdd.n871 185
R17882 vdd.n1173 vdd.n1172 185
R17883 vdd.n1172 vdd.n870 185
R17884 vdd.n1171 vdd.n878 185
R17885 vdd.n2175 vdd.n878 185
R17886 vdd.n1170 vdd.n1169 185
R17887 vdd.n1169 vdd.n877 185
R17888 vdd.n1168 vdd.n884 185
R17889 vdd.n2169 vdd.n884 185
R17890 vdd.n1167 vdd.n1166 185
R17891 vdd.n1166 vdd.n883 185
R17892 vdd.n1165 vdd.n889 185
R17893 vdd.n2163 vdd.n889 185
R17894 vdd.n1164 vdd.n1163 185
R17895 vdd.n1163 vdd.n896 185
R17896 vdd.n1162 vdd.n894 185
R17897 vdd.n2157 vdd.n894 185
R17898 vdd.n1161 vdd.n1160 185
R17899 vdd.n1160 vdd.n902 185
R17900 vdd.n1159 vdd.n900 185
R17901 vdd.n2151 vdd.n900 185
R17902 vdd.n1158 vdd.n1157 185
R17903 vdd.n1157 vdd.n909 185
R17904 vdd.n1156 vdd.n907 185
R17905 vdd.n2145 vdd.n907 185
R17906 vdd.n1155 vdd.n1154 185
R17907 vdd.n1154 vdd.n906 185
R17908 vdd.n1153 vdd.n914 185
R17909 vdd.n2139 vdd.n914 185
R17910 vdd.n1152 vdd.n1151 185
R17911 vdd.n1151 vdd.n913 185
R17912 vdd.n1150 vdd.n919 185
R17913 vdd.n2133 vdd.n919 185
R17914 vdd.n1149 vdd.n1148 185
R17915 vdd.n1148 vdd.n927 185
R17916 vdd.n1147 vdd.n925 185
R17917 vdd.n2127 vdd.n925 185
R17918 vdd.n1146 vdd.n1145 185
R17919 vdd.n1145 vdd.n924 185
R17920 vdd.n3296 vdd.n3295 185
R17921 vdd.n3297 vdd.n3296 185
R17922 vdd.n325 vdd.n324 185
R17923 vdd.n3298 vdd.n325 185
R17924 vdd.n3301 vdd.n3300 185
R17925 vdd.n3300 vdd.n3299 185
R17926 vdd.n3302 vdd.n319 185
R17927 vdd.n319 vdd.n318 185
R17928 vdd.n3304 vdd.n3303 185
R17929 vdd.n3305 vdd.n3304 185
R17930 vdd.n314 vdd.n313 185
R17931 vdd.n3306 vdd.n314 185
R17932 vdd.n3309 vdd.n3308 185
R17933 vdd.n3308 vdd.n3307 185
R17934 vdd.n3310 vdd.n309 185
R17935 vdd.n309 vdd.n308 185
R17936 vdd.n3312 vdd.n3311 185
R17937 vdd.n3313 vdd.n3312 185
R17938 vdd.n303 vdd.n301 185
R17939 vdd.n3314 vdd.n303 185
R17940 vdd.n3317 vdd.n3316 185
R17941 vdd.n3316 vdd.n3315 185
R17942 vdd.n302 vdd.n300 185
R17943 vdd.n304 vdd.n302 185
R17944 vdd.n3153 vdd.n3152 185
R17945 vdd.n3154 vdd.n3153 185
R17946 vdd.n458 vdd.n457 185
R17947 vdd.n457 vdd.n456 185
R17948 vdd.n3148 vdd.n3147 185
R17949 vdd.n3147 vdd.n3146 185
R17950 vdd.n461 vdd.n460 185
R17951 vdd.n467 vdd.n461 185
R17952 vdd.n3137 vdd.n3136 185
R17953 vdd.n3138 vdd.n3137 185
R17954 vdd.n469 vdd.n468 185
R17955 vdd.n3129 vdd.n468 185
R17956 vdd.n3132 vdd.n3131 185
R17957 vdd.n3131 vdd.n3130 185
R17958 vdd.n472 vdd.n471 185
R17959 vdd.n473 vdd.n472 185
R17960 vdd.n3120 vdd.n3119 185
R17961 vdd.n3121 vdd.n3120 185
R17962 vdd.n480 vdd.n479 185
R17963 vdd.n516 vdd.n479 185
R17964 vdd.n3115 vdd.n3114 185
R17965 vdd.n483 vdd.n482 185
R17966 vdd.n3111 vdd.n3110 185
R17967 vdd.n3112 vdd.n3111 185
R17968 vdd.n518 vdd.n517 185
R17969 vdd.n522 vdd.n521 185
R17970 vdd.n3106 vdd.n523 185
R17971 vdd.n3105 vdd.n3104 185
R17972 vdd.n3103 vdd.n3102 185
R17973 vdd.n3101 vdd.n3100 185
R17974 vdd.n3099 vdd.n3098 185
R17975 vdd.n3097 vdd.n3096 185
R17976 vdd.n3095 vdd.n3094 185
R17977 vdd.n3093 vdd.n3092 185
R17978 vdd.n3091 vdd.n3090 185
R17979 vdd.n3089 vdd.n3088 185
R17980 vdd.n3087 vdd.n3086 185
R17981 vdd.n3085 vdd.n3084 185
R17982 vdd.n3083 vdd.n3082 185
R17983 vdd.n3081 vdd.n3080 185
R17984 vdd.n3079 vdd.n3078 185
R17985 vdd.n3070 vdd.n536 185
R17986 vdd.n3072 vdd.n3071 185
R17987 vdd.n3069 vdd.n3068 185
R17988 vdd.n3067 vdd.n3066 185
R17989 vdd.n3065 vdd.n3064 185
R17990 vdd.n3063 vdd.n3062 185
R17991 vdd.n3061 vdd.n3060 185
R17992 vdd.n3059 vdd.n3058 185
R17993 vdd.n3057 vdd.n3056 185
R17994 vdd.n3055 vdd.n3054 185
R17995 vdd.n3053 vdd.n3052 185
R17996 vdd.n3051 vdd.n3050 185
R17997 vdd.n3049 vdd.n3048 185
R17998 vdd.n3047 vdd.n3046 185
R17999 vdd.n3045 vdd.n3044 185
R18000 vdd.n3043 vdd.n3042 185
R18001 vdd.n3041 vdd.n3040 185
R18002 vdd.n3039 vdd.n3038 185
R18003 vdd.n3037 vdd.n3036 185
R18004 vdd.n3035 vdd.n3034 185
R18005 vdd.n3033 vdd.n3032 185
R18006 vdd.n3031 vdd.n3030 185
R18007 vdd.n3024 vdd.n556 185
R18008 vdd.n3026 vdd.n3025 185
R18009 vdd.n3023 vdd.n3022 185
R18010 vdd.n3021 vdd.n3020 185
R18011 vdd.n3019 vdd.n3018 185
R18012 vdd.n3017 vdd.n3016 185
R18013 vdd.n3015 vdd.n3014 185
R18014 vdd.n3013 vdd.n3012 185
R18015 vdd.n3011 vdd.n3010 185
R18016 vdd.n3009 vdd.n3008 185
R18017 vdd.n3007 vdd.n3006 185
R18018 vdd.n3005 vdd.n3004 185
R18019 vdd.n3003 vdd.n3002 185
R18020 vdd.n3001 vdd.n3000 185
R18021 vdd.n2999 vdd.n2998 185
R18022 vdd.n2997 vdd.n2996 185
R18023 vdd.n2995 vdd.n2994 185
R18024 vdd.n2993 vdd.n2992 185
R18025 vdd.n2991 vdd.n2990 185
R18026 vdd.n2989 vdd.n2988 185
R18027 vdd.n2987 vdd.n2986 185
R18028 vdd.n2982 vdd.n515 185
R18029 vdd.n3112 vdd.n515 185
R18030 vdd.n3179 vdd.n3178 185
R18031 vdd.n3183 vdd.n440 185
R18032 vdd.n3185 vdd.n3184 185
R18033 vdd.n3187 vdd.n438 185
R18034 vdd.n3189 vdd.n3188 185
R18035 vdd.n3190 vdd.n433 185
R18036 vdd.n3192 vdd.n3191 185
R18037 vdd.n3194 vdd.n431 185
R18038 vdd.n3196 vdd.n3195 185
R18039 vdd.n3197 vdd.n426 185
R18040 vdd.n3199 vdd.n3198 185
R18041 vdd.n3201 vdd.n424 185
R18042 vdd.n3203 vdd.n3202 185
R18043 vdd.n3204 vdd.n419 185
R18044 vdd.n3206 vdd.n3205 185
R18045 vdd.n3208 vdd.n417 185
R18046 vdd.n3210 vdd.n3209 185
R18047 vdd.n3211 vdd.n413 185
R18048 vdd.n3213 vdd.n3212 185
R18049 vdd.n3215 vdd.n410 185
R18050 vdd.n3217 vdd.n3216 185
R18051 vdd.n411 vdd.n404 185
R18052 vdd.n3221 vdd.n408 185
R18053 vdd.n3222 vdd.n400 185
R18054 vdd.n3224 vdd.n3223 185
R18055 vdd.n3226 vdd.n398 185
R18056 vdd.n3228 vdd.n3227 185
R18057 vdd.n3229 vdd.n393 185
R18058 vdd.n3231 vdd.n3230 185
R18059 vdd.n3233 vdd.n391 185
R18060 vdd.n3235 vdd.n3234 185
R18061 vdd.n3236 vdd.n386 185
R18062 vdd.n3238 vdd.n3237 185
R18063 vdd.n3240 vdd.n384 185
R18064 vdd.n3242 vdd.n3241 185
R18065 vdd.n3243 vdd.n379 185
R18066 vdd.n3245 vdd.n3244 185
R18067 vdd.n3247 vdd.n377 185
R18068 vdd.n3249 vdd.n3248 185
R18069 vdd.n3250 vdd.n373 185
R18070 vdd.n3252 vdd.n3251 185
R18071 vdd.n3254 vdd.n370 185
R18072 vdd.n3256 vdd.n3255 185
R18073 vdd.n371 vdd.n364 185
R18074 vdd.n3260 vdd.n368 185
R18075 vdd.n3261 vdd.n360 185
R18076 vdd.n3263 vdd.n3262 185
R18077 vdd.n3265 vdd.n358 185
R18078 vdd.n3267 vdd.n3266 185
R18079 vdd.n3268 vdd.n353 185
R18080 vdd.n3270 vdd.n3269 185
R18081 vdd.n3272 vdd.n351 185
R18082 vdd.n3274 vdd.n3273 185
R18083 vdd.n3275 vdd.n346 185
R18084 vdd.n3277 vdd.n3276 185
R18085 vdd.n3279 vdd.n344 185
R18086 vdd.n3281 vdd.n3280 185
R18087 vdd.n3282 vdd.n338 185
R18088 vdd.n3284 vdd.n3283 185
R18089 vdd.n3286 vdd.n337 185
R18090 vdd.n3287 vdd.n336 185
R18091 vdd.n3290 vdd.n3289 185
R18092 vdd.n3291 vdd.n334 185
R18093 vdd.n3292 vdd.n330 185
R18094 vdd.n3174 vdd.n328 185
R18095 vdd.n3297 vdd.n328 185
R18096 vdd.n3173 vdd.n327 185
R18097 vdd.n3298 vdd.n327 185
R18098 vdd.n3172 vdd.n326 185
R18099 vdd.n3299 vdd.n326 185
R18100 vdd.n446 vdd.n445 185
R18101 vdd.n445 vdd.n318 185
R18102 vdd.n3168 vdd.n317 185
R18103 vdd.n3305 vdd.n317 185
R18104 vdd.n3167 vdd.n316 185
R18105 vdd.n3306 vdd.n316 185
R18106 vdd.n3166 vdd.n315 185
R18107 vdd.n3307 vdd.n315 185
R18108 vdd.n449 vdd.n448 185
R18109 vdd.n448 vdd.n308 185
R18110 vdd.n3162 vdd.n307 185
R18111 vdd.n3313 vdd.n307 185
R18112 vdd.n3161 vdd.n306 185
R18113 vdd.n3314 vdd.n306 185
R18114 vdd.n3160 vdd.n305 185
R18115 vdd.n3315 vdd.n305 185
R18116 vdd.n455 vdd.n451 185
R18117 vdd.n455 vdd.n304 185
R18118 vdd.n3156 vdd.n3155 185
R18119 vdd.n3155 vdd.n3154 185
R18120 vdd.n454 vdd.n453 185
R18121 vdd.n456 vdd.n454 185
R18122 vdd.n3145 vdd.n3144 185
R18123 vdd.n3146 vdd.n3145 185
R18124 vdd.n463 vdd.n462 185
R18125 vdd.n467 vdd.n462 185
R18126 vdd.n3140 vdd.n3139 185
R18127 vdd.n3139 vdd.n3138 185
R18128 vdd.n466 vdd.n465 185
R18129 vdd.n3129 vdd.n466 185
R18130 vdd.n3128 vdd.n3127 185
R18131 vdd.n3130 vdd.n3128 185
R18132 vdd.n475 vdd.n474 185
R18133 vdd.n474 vdd.n473 185
R18134 vdd.n3123 vdd.n3122 185
R18135 vdd.n3122 vdd.n3121 185
R18136 vdd.n478 vdd.n477 185
R18137 vdd.n516 vdd.n478 185
R18138 vdd.n2705 vdd.n2704 185
R18139 vdd.n752 vdd.n751 185
R18140 vdd.n2701 vdd.n2700 185
R18141 vdd.n2702 vdd.n2701 185
R18142 vdd.n2699 vdd.n2433 185
R18143 vdd.n2698 vdd.n2697 185
R18144 vdd.n2696 vdd.n2695 185
R18145 vdd.n2694 vdd.n2693 185
R18146 vdd.n2692 vdd.n2691 185
R18147 vdd.n2690 vdd.n2689 185
R18148 vdd.n2688 vdd.n2687 185
R18149 vdd.n2686 vdd.n2685 185
R18150 vdd.n2684 vdd.n2683 185
R18151 vdd.n2682 vdd.n2681 185
R18152 vdd.n2680 vdd.n2679 185
R18153 vdd.n2678 vdd.n2677 185
R18154 vdd.n2676 vdd.n2675 185
R18155 vdd.n2674 vdd.n2673 185
R18156 vdd.n2672 vdd.n2671 185
R18157 vdd.n2670 vdd.n2669 185
R18158 vdd.n2668 vdd.n2667 185
R18159 vdd.n2666 vdd.n2665 185
R18160 vdd.n2664 vdd.n2663 185
R18161 vdd.n2662 vdd.n2661 185
R18162 vdd.n2660 vdd.n2659 185
R18163 vdd.n2658 vdd.n2657 185
R18164 vdd.n2656 vdd.n2655 185
R18165 vdd.n2654 vdd.n2653 185
R18166 vdd.n2652 vdd.n2651 185
R18167 vdd.n2650 vdd.n2649 185
R18168 vdd.n2648 vdd.n2647 185
R18169 vdd.n2646 vdd.n2645 185
R18170 vdd.n2644 vdd.n2643 185
R18171 vdd.n2641 vdd.n2640 185
R18172 vdd.n2639 vdd.n2638 185
R18173 vdd.n2637 vdd.n2636 185
R18174 vdd.n2881 vdd.n2880 185
R18175 vdd.n2883 vdd.n624 185
R18176 vdd.n2885 vdd.n2884 185
R18177 vdd.n2887 vdd.n621 185
R18178 vdd.n2889 vdd.n2888 185
R18179 vdd.n2891 vdd.n619 185
R18180 vdd.n2893 vdd.n2892 185
R18181 vdd.n2894 vdd.n618 185
R18182 vdd.n2896 vdd.n2895 185
R18183 vdd.n2898 vdd.n616 185
R18184 vdd.n2900 vdd.n2899 185
R18185 vdd.n2901 vdd.n615 185
R18186 vdd.n2903 vdd.n2902 185
R18187 vdd.n2905 vdd.n613 185
R18188 vdd.n2907 vdd.n2906 185
R18189 vdd.n2908 vdd.n612 185
R18190 vdd.n2910 vdd.n2909 185
R18191 vdd.n2912 vdd.n520 185
R18192 vdd.n2914 vdd.n2913 185
R18193 vdd.n2916 vdd.n610 185
R18194 vdd.n2918 vdd.n2917 185
R18195 vdd.n2919 vdd.n609 185
R18196 vdd.n2921 vdd.n2920 185
R18197 vdd.n2923 vdd.n607 185
R18198 vdd.n2925 vdd.n2924 185
R18199 vdd.n2926 vdd.n606 185
R18200 vdd.n2928 vdd.n2927 185
R18201 vdd.n2930 vdd.n604 185
R18202 vdd.n2932 vdd.n2931 185
R18203 vdd.n2933 vdd.n603 185
R18204 vdd.n2935 vdd.n2934 185
R18205 vdd.n2937 vdd.n602 185
R18206 vdd.n2938 vdd.n601 185
R18207 vdd.n2941 vdd.n2940 185
R18208 vdd.n2942 vdd.n599 185
R18209 vdd.n599 vdd.n484 185
R18210 vdd.n2879 vdd.n596 185
R18211 vdd.n2945 vdd.n596 185
R18212 vdd.n2878 vdd.n2877 185
R18213 vdd.n2877 vdd.n595 185
R18214 vdd.n2876 vdd.n626 185
R18215 vdd.n2876 vdd.n2875 185
R18216 vdd.n2519 vdd.n627 185
R18217 vdd.n636 vdd.n627 185
R18218 vdd.n2520 vdd.n634 185
R18219 vdd.n2869 vdd.n634 185
R18220 vdd.n2522 vdd.n2521 185
R18221 vdd.n2521 vdd.n633 185
R18222 vdd.n2523 vdd.n642 185
R18223 vdd.n2818 vdd.n642 185
R18224 vdd.n2525 vdd.n2524 185
R18225 vdd.n2524 vdd.n641 185
R18226 vdd.n2526 vdd.n647 185
R18227 vdd.n2812 vdd.n647 185
R18228 vdd.n2528 vdd.n2527 185
R18229 vdd.n2527 vdd.n654 185
R18230 vdd.n2529 vdd.n652 185
R18231 vdd.n2806 vdd.n652 185
R18232 vdd.n2531 vdd.n2530 185
R18233 vdd.n2530 vdd.n660 185
R18234 vdd.n2532 vdd.n658 185
R18235 vdd.n2800 vdd.n658 185
R18236 vdd.n2534 vdd.n2533 185
R18237 vdd.n2533 vdd.n667 185
R18238 vdd.n2535 vdd.n665 185
R18239 vdd.n2794 vdd.n665 185
R18240 vdd.n2537 vdd.n2536 185
R18241 vdd.n2536 vdd.n664 185
R18242 vdd.n2538 vdd.n672 185
R18243 vdd.n2788 vdd.n672 185
R18244 vdd.n2540 vdd.n2539 185
R18245 vdd.n2539 vdd.n671 185
R18246 vdd.n2541 vdd.n678 185
R18247 vdd.n2782 vdd.n678 185
R18248 vdd.n2543 vdd.n2542 185
R18249 vdd.n2542 vdd.n677 185
R18250 vdd.n2544 vdd.n683 185
R18251 vdd.n2776 vdd.n683 185
R18252 vdd.n2546 vdd.n2545 185
R18253 vdd.n2545 vdd.n691 185
R18254 vdd.n2547 vdd.n689 185
R18255 vdd.n2770 vdd.n689 185
R18256 vdd.n2549 vdd.n2548 185
R18257 vdd.n2548 vdd.n698 185
R18258 vdd.n2550 vdd.n696 185
R18259 vdd.n2764 vdd.n696 185
R18260 vdd.n2552 vdd.n2551 185
R18261 vdd.n2551 vdd.n695 185
R18262 vdd.n2553 vdd.n703 185
R18263 vdd.n2757 vdd.n703 185
R18264 vdd.n2555 vdd.n2554 185
R18265 vdd.n2554 vdd.n702 185
R18266 vdd.n2556 vdd.n708 185
R18267 vdd.n2751 vdd.n708 185
R18268 vdd.n2558 vdd.n2557 185
R18269 vdd.n2557 vdd.n715 185
R18270 vdd.n2559 vdd.n713 185
R18271 vdd.n2745 vdd.n713 185
R18272 vdd.n2561 vdd.n2560 185
R18273 vdd.n2560 vdd.n721 185
R18274 vdd.n2562 vdd.n719 185
R18275 vdd.n2739 vdd.n719 185
R18276 vdd.n2614 vdd.n2613 185
R18277 vdd.n2613 vdd.n2612 185
R18278 vdd.n2615 vdd.n725 185
R18279 vdd.n2733 vdd.n725 185
R18280 vdd.n2617 vdd.n2616 185
R18281 vdd.n2618 vdd.n2617 185
R18282 vdd.n2518 vdd.n731 185
R18283 vdd.n2727 vdd.n731 185
R18284 vdd.n2517 vdd.n2516 185
R18285 vdd.n2516 vdd.n730 185
R18286 vdd.n2515 vdd.n737 185
R18287 vdd.n2721 vdd.n737 185
R18288 vdd.n2514 vdd.n2513 185
R18289 vdd.n2513 vdd.n736 185
R18290 vdd.n2436 vdd.n742 185
R18291 vdd.n2715 vdd.n742 185
R18292 vdd.n2632 vdd.n2631 185
R18293 vdd.n2631 vdd.n2630 185
R18294 vdd.n2633 vdd.n748 185
R18295 vdd.n2709 vdd.n748 185
R18296 vdd.n2635 vdd.n2634 185
R18297 vdd.n2635 vdd.n747 185
R18298 vdd.n2706 vdd.n750 185
R18299 vdd.n750 vdd.n747 185
R18300 vdd.n2708 vdd.n2707 185
R18301 vdd.n2709 vdd.n2708 185
R18302 vdd.n741 vdd.n740 185
R18303 vdd.n2630 vdd.n741 185
R18304 vdd.n2717 vdd.n2716 185
R18305 vdd.n2716 vdd.n2715 185
R18306 vdd.n2718 vdd.n739 185
R18307 vdd.n739 vdd.n736 185
R18308 vdd.n2720 vdd.n2719 185
R18309 vdd.n2721 vdd.n2720 185
R18310 vdd.n729 vdd.n728 185
R18311 vdd.n730 vdd.n729 185
R18312 vdd.n2729 vdd.n2728 185
R18313 vdd.n2728 vdd.n2727 185
R18314 vdd.n2730 vdd.n727 185
R18315 vdd.n2618 vdd.n727 185
R18316 vdd.n2732 vdd.n2731 185
R18317 vdd.n2733 vdd.n2732 185
R18318 vdd.n718 vdd.n717 185
R18319 vdd.n2612 vdd.n718 185
R18320 vdd.n2741 vdd.n2740 185
R18321 vdd.n2740 vdd.n2739 185
R18322 vdd.n2742 vdd.n716 185
R18323 vdd.n721 vdd.n716 185
R18324 vdd.n2744 vdd.n2743 185
R18325 vdd.n2745 vdd.n2744 185
R18326 vdd.n707 vdd.n706 185
R18327 vdd.n715 vdd.n707 185
R18328 vdd.n2753 vdd.n2752 185
R18329 vdd.n2752 vdd.n2751 185
R18330 vdd.n2754 vdd.n705 185
R18331 vdd.n705 vdd.n702 185
R18332 vdd.n2756 vdd.n2755 185
R18333 vdd.n2757 vdd.n2756 185
R18334 vdd.n694 vdd.n693 185
R18335 vdd.n695 vdd.n694 185
R18336 vdd.n2766 vdd.n2765 185
R18337 vdd.n2765 vdd.n2764 185
R18338 vdd.n2767 vdd.n692 185
R18339 vdd.n698 vdd.n692 185
R18340 vdd.n2769 vdd.n2768 185
R18341 vdd.n2770 vdd.n2769 185
R18342 vdd.n682 vdd.n681 185
R18343 vdd.n691 vdd.n682 185
R18344 vdd.n2778 vdd.n2777 185
R18345 vdd.n2777 vdd.n2776 185
R18346 vdd.n2779 vdd.n680 185
R18347 vdd.n680 vdd.n677 185
R18348 vdd.n2781 vdd.n2780 185
R18349 vdd.n2782 vdd.n2781 185
R18350 vdd.n670 vdd.n669 185
R18351 vdd.n671 vdd.n670 185
R18352 vdd.n2790 vdd.n2789 185
R18353 vdd.n2789 vdd.n2788 185
R18354 vdd.n2791 vdd.n668 185
R18355 vdd.n668 vdd.n664 185
R18356 vdd.n2793 vdd.n2792 185
R18357 vdd.n2794 vdd.n2793 185
R18358 vdd.n657 vdd.n656 185
R18359 vdd.n667 vdd.n657 185
R18360 vdd.n2802 vdd.n2801 185
R18361 vdd.n2801 vdd.n2800 185
R18362 vdd.n2803 vdd.n655 185
R18363 vdd.n660 vdd.n655 185
R18364 vdd.n2805 vdd.n2804 185
R18365 vdd.n2806 vdd.n2805 185
R18366 vdd.n646 vdd.n645 185
R18367 vdd.n654 vdd.n646 185
R18368 vdd.n2814 vdd.n2813 185
R18369 vdd.n2813 vdd.n2812 185
R18370 vdd.n2815 vdd.n644 185
R18371 vdd.n644 vdd.n641 185
R18372 vdd.n2817 vdd.n2816 185
R18373 vdd.n2818 vdd.n2817 185
R18374 vdd.n632 vdd.n631 185
R18375 vdd.n633 vdd.n632 185
R18376 vdd.n2871 vdd.n2870 185
R18377 vdd.n2870 vdd.n2869 185
R18378 vdd.n2872 vdd.n630 185
R18379 vdd.n636 vdd.n630 185
R18380 vdd.n2874 vdd.n2873 185
R18381 vdd.n2875 vdd.n2874 185
R18382 vdd.n600 vdd.n598 185
R18383 vdd.n598 vdd.n595 185
R18384 vdd.n2944 vdd.n2943 185
R18385 vdd.n2945 vdd.n2944 185
R18386 vdd.n2325 vdd.n2324 185
R18387 vdd.n2326 vdd.n2325 185
R18388 vdd.n799 vdd.n797 185
R18389 vdd.n797 vdd.n795 185
R18390 vdd.n2240 vdd.n806 185
R18391 vdd.n2251 vdd.n806 185
R18392 vdd.n2241 vdd.n815 185
R18393 vdd.n1189 vdd.n815 185
R18394 vdd.n2243 vdd.n2242 185
R18395 vdd.n2244 vdd.n2243 185
R18396 vdd.n2239 vdd.n814 185
R18397 vdd.n814 vdd.n811 185
R18398 vdd.n2238 vdd.n2237 185
R18399 vdd.n2237 vdd.n2236 185
R18400 vdd.n817 vdd.n816 185
R18401 vdd.n818 vdd.n817 185
R18402 vdd.n2229 vdd.n2228 185
R18403 vdd.n2230 vdd.n2229 185
R18404 vdd.n2227 vdd.n826 185
R18405 vdd.n1215 vdd.n826 185
R18406 vdd.n2226 vdd.n2225 185
R18407 vdd.n2225 vdd.n2224 185
R18408 vdd.n828 vdd.n827 185
R18409 vdd.n836 vdd.n828 185
R18410 vdd.n2217 vdd.n2216 185
R18411 vdd.n2218 vdd.n2217 185
R18412 vdd.n2215 vdd.n837 185
R18413 vdd.n842 vdd.n837 185
R18414 vdd.n2214 vdd.n2213 185
R18415 vdd.n2213 vdd.n2212 185
R18416 vdd.n839 vdd.n838 185
R18417 vdd.n1227 vdd.n839 185
R18418 vdd.n2205 vdd.n2204 185
R18419 vdd.n2206 vdd.n2205 185
R18420 vdd.n2203 vdd.n849 185
R18421 vdd.n849 vdd.n846 185
R18422 vdd.n2202 vdd.n2201 185
R18423 vdd.n2201 vdd.n2200 185
R18424 vdd.n851 vdd.n850 185
R18425 vdd.n852 vdd.n851 185
R18426 vdd.n2193 vdd.n2192 185
R18427 vdd.n2194 vdd.n2193 185
R18428 vdd.n2190 vdd.n860 185
R18429 vdd.n866 vdd.n860 185
R18430 vdd.n2189 vdd.n2188 185
R18431 vdd.n2188 vdd.n2187 185
R18432 vdd.n863 vdd.n862 185
R18433 vdd.n873 vdd.n863 185
R18434 vdd.n2180 vdd.n2179 185
R18435 vdd.n2181 vdd.n2180 185
R18436 vdd.n2178 vdd.n874 185
R18437 vdd.n874 vdd.n870 185
R18438 vdd.n2177 vdd.n2176 185
R18439 vdd.n2176 vdd.n2175 185
R18440 vdd.n876 vdd.n875 185
R18441 vdd.n877 vdd.n876 185
R18442 vdd.n2168 vdd.n2167 185
R18443 vdd.n2169 vdd.n2168 185
R18444 vdd.n2166 vdd.n886 185
R18445 vdd.n886 vdd.n883 185
R18446 vdd.n2165 vdd.n2164 185
R18447 vdd.n2164 vdd.n2163 185
R18448 vdd.n888 vdd.n887 185
R18449 vdd.n896 vdd.n888 185
R18450 vdd.n2156 vdd.n2155 185
R18451 vdd.n2157 vdd.n2156 185
R18452 vdd.n2154 vdd.n897 185
R18453 vdd.n902 vdd.n897 185
R18454 vdd.n2153 vdd.n2152 185
R18455 vdd.n2152 vdd.n2151 185
R18456 vdd.n899 vdd.n898 185
R18457 vdd.n909 vdd.n899 185
R18458 vdd.n2144 vdd.n2143 185
R18459 vdd.n2145 vdd.n2144 185
R18460 vdd.n2142 vdd.n910 185
R18461 vdd.n910 vdd.n906 185
R18462 vdd.n2141 vdd.n2140 185
R18463 vdd.n2140 vdd.n2139 185
R18464 vdd.n912 vdd.n911 185
R18465 vdd.n913 vdd.n912 185
R18466 vdd.n2132 vdd.n2131 185
R18467 vdd.n2133 vdd.n2132 185
R18468 vdd.n2130 vdd.n921 185
R18469 vdd.n927 vdd.n921 185
R18470 vdd.n2129 vdd.n2128 185
R18471 vdd.n2128 vdd.n2127 185
R18472 vdd.n923 vdd.n922 185
R18473 vdd.n924 vdd.n923 185
R18474 vdd.n2256 vdd.n770 185
R18475 vdd.n2398 vdd.n770 185
R18476 vdd.n2258 vdd.n2257 185
R18477 vdd.n2260 vdd.n2259 185
R18478 vdd.n2262 vdd.n2261 185
R18479 vdd.n2264 vdd.n2263 185
R18480 vdd.n2266 vdd.n2265 185
R18481 vdd.n2268 vdd.n2267 185
R18482 vdd.n2270 vdd.n2269 185
R18483 vdd.n2272 vdd.n2271 185
R18484 vdd.n2274 vdd.n2273 185
R18485 vdd.n2276 vdd.n2275 185
R18486 vdd.n2278 vdd.n2277 185
R18487 vdd.n2280 vdd.n2279 185
R18488 vdd.n2282 vdd.n2281 185
R18489 vdd.n2284 vdd.n2283 185
R18490 vdd.n2286 vdd.n2285 185
R18491 vdd.n2288 vdd.n2287 185
R18492 vdd.n2290 vdd.n2289 185
R18493 vdd.n2292 vdd.n2291 185
R18494 vdd.n2294 vdd.n2293 185
R18495 vdd.n2296 vdd.n2295 185
R18496 vdd.n2298 vdd.n2297 185
R18497 vdd.n2300 vdd.n2299 185
R18498 vdd.n2302 vdd.n2301 185
R18499 vdd.n2304 vdd.n2303 185
R18500 vdd.n2306 vdd.n2305 185
R18501 vdd.n2308 vdd.n2307 185
R18502 vdd.n2310 vdd.n2309 185
R18503 vdd.n2312 vdd.n2311 185
R18504 vdd.n2314 vdd.n2313 185
R18505 vdd.n2316 vdd.n2315 185
R18506 vdd.n2318 vdd.n2317 185
R18507 vdd.n2320 vdd.n2319 185
R18508 vdd.n2322 vdd.n2321 185
R18509 vdd.n2323 vdd.n798 185
R18510 vdd.n2255 vdd.n796 185
R18511 vdd.n2326 vdd.n796 185
R18512 vdd.n2254 vdd.n2253 185
R18513 vdd.n2253 vdd.n795 185
R18514 vdd.n2252 vdd.n803 185
R18515 vdd.n2252 vdd.n2251 185
R18516 vdd.n1205 vdd.n804 185
R18517 vdd.n1189 vdd.n804 185
R18518 vdd.n1206 vdd.n813 185
R18519 vdd.n2244 vdd.n813 185
R18520 vdd.n1208 vdd.n1207 185
R18521 vdd.n1207 vdd.n811 185
R18522 vdd.n1209 vdd.n820 185
R18523 vdd.n2236 vdd.n820 185
R18524 vdd.n1211 vdd.n1210 185
R18525 vdd.n1210 vdd.n818 185
R18526 vdd.n1212 vdd.n825 185
R18527 vdd.n2230 vdd.n825 185
R18528 vdd.n1214 vdd.n1213 185
R18529 vdd.n1215 vdd.n1214 185
R18530 vdd.n1204 vdd.n830 185
R18531 vdd.n2224 vdd.n830 185
R18532 vdd.n1203 vdd.n1202 185
R18533 vdd.n1202 vdd.n836 185
R18534 vdd.n1201 vdd.n835 185
R18535 vdd.n2218 vdd.n835 185
R18536 vdd.n1200 vdd.n1199 185
R18537 vdd.n1199 vdd.n842 185
R18538 vdd.n1108 vdd.n841 185
R18539 vdd.n2212 vdd.n841 185
R18540 vdd.n1229 vdd.n1228 185
R18541 vdd.n1228 vdd.n1227 185
R18542 vdd.n1230 vdd.n848 185
R18543 vdd.n2206 vdd.n848 185
R18544 vdd.n1232 vdd.n1231 185
R18545 vdd.n1231 vdd.n846 185
R18546 vdd.n1233 vdd.n854 185
R18547 vdd.n2200 vdd.n854 185
R18548 vdd.n1235 vdd.n1234 185
R18549 vdd.n1234 vdd.n852 185
R18550 vdd.n1236 vdd.n859 185
R18551 vdd.n2194 vdd.n859 185
R18552 vdd.n1238 vdd.n1237 185
R18553 vdd.n1237 vdd.n866 185
R18554 vdd.n1239 vdd.n865 185
R18555 vdd.n2187 vdd.n865 185
R18556 vdd.n1241 vdd.n1240 185
R18557 vdd.n1240 vdd.n873 185
R18558 vdd.n1242 vdd.n872 185
R18559 vdd.n2181 vdd.n872 185
R18560 vdd.n1244 vdd.n1243 185
R18561 vdd.n1243 vdd.n870 185
R18562 vdd.n1245 vdd.n879 185
R18563 vdd.n2175 vdd.n879 185
R18564 vdd.n1247 vdd.n1246 185
R18565 vdd.n1246 vdd.n877 185
R18566 vdd.n1248 vdd.n885 185
R18567 vdd.n2169 vdd.n885 185
R18568 vdd.n1250 vdd.n1249 185
R18569 vdd.n1249 vdd.n883 185
R18570 vdd.n1251 vdd.n890 185
R18571 vdd.n2163 vdd.n890 185
R18572 vdd.n1253 vdd.n1252 185
R18573 vdd.n1252 vdd.n896 185
R18574 vdd.n1254 vdd.n895 185
R18575 vdd.n2157 vdd.n895 185
R18576 vdd.n1256 vdd.n1255 185
R18577 vdd.n1255 vdd.n902 185
R18578 vdd.n1257 vdd.n901 185
R18579 vdd.n2151 vdd.n901 185
R18580 vdd.n1259 vdd.n1258 185
R18581 vdd.n1258 vdd.n909 185
R18582 vdd.n1260 vdd.n908 185
R18583 vdd.n2145 vdd.n908 185
R18584 vdd.n1262 vdd.n1261 185
R18585 vdd.n1261 vdd.n906 185
R18586 vdd.n1263 vdd.n915 185
R18587 vdd.n2139 vdd.n915 185
R18588 vdd.n1265 vdd.n1264 185
R18589 vdd.n1264 vdd.n913 185
R18590 vdd.n1266 vdd.n920 185
R18591 vdd.n2133 vdd.n920 185
R18592 vdd.n1268 vdd.n1267 185
R18593 vdd.n1267 vdd.n927 185
R18594 vdd.n1269 vdd.n926 185
R18595 vdd.n2127 vdd.n926 185
R18596 vdd.n1271 vdd.n1270 185
R18597 vdd.n1270 vdd.n924 185
R18598 vdd.n1071 vdd.n1070 185
R18599 vdd.n1073 vdd.n1072 185
R18600 vdd.n1075 vdd.n1074 185
R18601 vdd.n1077 vdd.n1076 185
R18602 vdd.n1079 vdd.n1078 185
R18603 vdd.n1081 vdd.n1080 185
R18604 vdd.n1083 vdd.n1082 185
R18605 vdd.n1085 vdd.n1084 185
R18606 vdd.n1087 vdd.n1086 185
R18607 vdd.n1089 vdd.n1088 185
R18608 vdd.n1091 vdd.n1090 185
R18609 vdd.n1093 vdd.n1092 185
R18610 vdd.n1095 vdd.n1094 185
R18611 vdd.n1097 vdd.n1096 185
R18612 vdd.n1099 vdd.n1098 185
R18613 vdd.n1101 vdd.n1100 185
R18614 vdd.n1103 vdd.n1102 185
R18615 vdd.n1305 vdd.n1104 185
R18616 vdd.n1304 vdd.n1303 185
R18617 vdd.n1302 vdd.n1301 185
R18618 vdd.n1300 vdd.n1299 185
R18619 vdd.n1298 vdd.n1297 185
R18620 vdd.n1296 vdd.n1295 185
R18621 vdd.n1294 vdd.n1293 185
R18622 vdd.n1292 vdd.n1291 185
R18623 vdd.n1290 vdd.n1289 185
R18624 vdd.n1288 vdd.n1287 185
R18625 vdd.n1286 vdd.n1285 185
R18626 vdd.n1284 vdd.n1283 185
R18627 vdd.n1282 vdd.n1281 185
R18628 vdd.n1280 vdd.n1279 185
R18629 vdd.n1278 vdd.n1277 185
R18630 vdd.n1276 vdd.n1275 185
R18631 vdd.n1274 vdd.n1273 185
R18632 vdd.n1272 vdd.n965 185
R18633 vdd.n2120 vdd.n965 185
R18634 vdd.n291 vdd.n290 171.744
R18635 vdd.n290 vdd.n289 171.744
R18636 vdd.n289 vdd.n258 171.744
R18637 vdd.n282 vdd.n258 171.744
R18638 vdd.n282 vdd.n281 171.744
R18639 vdd.n281 vdd.n263 171.744
R18640 vdd.n274 vdd.n263 171.744
R18641 vdd.n274 vdd.n273 171.744
R18642 vdd.n273 vdd.n267 171.744
R18643 vdd.n244 vdd.n243 171.744
R18644 vdd.n243 vdd.n242 171.744
R18645 vdd.n242 vdd.n211 171.744
R18646 vdd.n235 vdd.n211 171.744
R18647 vdd.n235 vdd.n234 171.744
R18648 vdd.n234 vdd.n216 171.744
R18649 vdd.n227 vdd.n216 171.744
R18650 vdd.n227 vdd.n226 171.744
R18651 vdd.n226 vdd.n220 171.744
R18652 vdd.n201 vdd.n200 171.744
R18653 vdd.n200 vdd.n199 171.744
R18654 vdd.n199 vdd.n168 171.744
R18655 vdd.n192 vdd.n168 171.744
R18656 vdd.n192 vdd.n191 171.744
R18657 vdd.n191 vdd.n173 171.744
R18658 vdd.n184 vdd.n173 171.744
R18659 vdd.n184 vdd.n183 171.744
R18660 vdd.n183 vdd.n177 171.744
R18661 vdd.n154 vdd.n153 171.744
R18662 vdd.n153 vdd.n152 171.744
R18663 vdd.n152 vdd.n121 171.744
R18664 vdd.n145 vdd.n121 171.744
R18665 vdd.n145 vdd.n144 171.744
R18666 vdd.n144 vdd.n126 171.744
R18667 vdd.n137 vdd.n126 171.744
R18668 vdd.n137 vdd.n136 171.744
R18669 vdd.n136 vdd.n130 171.744
R18670 vdd.n112 vdd.n111 171.744
R18671 vdd.n111 vdd.n110 171.744
R18672 vdd.n110 vdd.n79 171.744
R18673 vdd.n103 vdd.n79 171.744
R18674 vdd.n103 vdd.n102 171.744
R18675 vdd.n102 vdd.n84 171.744
R18676 vdd.n95 vdd.n84 171.744
R18677 vdd.n95 vdd.n94 171.744
R18678 vdd.n94 vdd.n88 171.744
R18679 vdd.n65 vdd.n64 171.744
R18680 vdd.n64 vdd.n63 171.744
R18681 vdd.n63 vdd.n32 171.744
R18682 vdd.n56 vdd.n32 171.744
R18683 vdd.n56 vdd.n55 171.744
R18684 vdd.n55 vdd.n37 171.744
R18685 vdd.n48 vdd.n37 171.744
R18686 vdd.n48 vdd.n47 171.744
R18687 vdd.n47 vdd.n41 171.744
R18688 vdd.n1561 vdd.n1560 171.744
R18689 vdd.n1560 vdd.n1559 171.744
R18690 vdd.n1559 vdd.n1528 171.744
R18691 vdd.n1552 vdd.n1528 171.744
R18692 vdd.n1552 vdd.n1551 171.744
R18693 vdd.n1551 vdd.n1533 171.744
R18694 vdd.n1544 vdd.n1533 171.744
R18695 vdd.n1544 vdd.n1543 171.744
R18696 vdd.n1543 vdd.n1537 171.744
R18697 vdd.n1608 vdd.n1607 171.744
R18698 vdd.n1607 vdd.n1606 171.744
R18699 vdd.n1606 vdd.n1575 171.744
R18700 vdd.n1599 vdd.n1575 171.744
R18701 vdd.n1599 vdd.n1598 171.744
R18702 vdd.n1598 vdd.n1580 171.744
R18703 vdd.n1591 vdd.n1580 171.744
R18704 vdd.n1591 vdd.n1590 171.744
R18705 vdd.n1590 vdd.n1584 171.744
R18706 vdd.n1471 vdd.n1470 171.744
R18707 vdd.n1470 vdd.n1469 171.744
R18708 vdd.n1469 vdd.n1438 171.744
R18709 vdd.n1462 vdd.n1438 171.744
R18710 vdd.n1462 vdd.n1461 171.744
R18711 vdd.n1461 vdd.n1443 171.744
R18712 vdd.n1454 vdd.n1443 171.744
R18713 vdd.n1454 vdd.n1453 171.744
R18714 vdd.n1453 vdd.n1447 171.744
R18715 vdd.n1518 vdd.n1517 171.744
R18716 vdd.n1517 vdd.n1516 171.744
R18717 vdd.n1516 vdd.n1485 171.744
R18718 vdd.n1509 vdd.n1485 171.744
R18719 vdd.n1509 vdd.n1508 171.744
R18720 vdd.n1508 vdd.n1490 171.744
R18721 vdd.n1501 vdd.n1490 171.744
R18722 vdd.n1501 vdd.n1500 171.744
R18723 vdd.n1500 vdd.n1494 171.744
R18724 vdd.n1382 vdd.n1381 171.744
R18725 vdd.n1381 vdd.n1380 171.744
R18726 vdd.n1380 vdd.n1349 171.744
R18727 vdd.n1373 vdd.n1349 171.744
R18728 vdd.n1373 vdd.n1372 171.744
R18729 vdd.n1372 vdd.n1354 171.744
R18730 vdd.n1365 vdd.n1354 171.744
R18731 vdd.n1365 vdd.n1364 171.744
R18732 vdd.n1364 vdd.n1358 171.744
R18733 vdd.n1429 vdd.n1428 171.744
R18734 vdd.n1428 vdd.n1427 171.744
R18735 vdd.n1427 vdd.n1396 171.744
R18736 vdd.n1420 vdd.n1396 171.744
R18737 vdd.n1420 vdd.n1419 171.744
R18738 vdd.n1419 vdd.n1401 171.744
R18739 vdd.n1412 vdd.n1401 171.744
R18740 vdd.n1412 vdd.n1411 171.744
R18741 vdd.n1411 vdd.n1405 171.744
R18742 vdd.n3289 vdd.n334 146.341
R18743 vdd.n3287 vdd.n3286 146.341
R18744 vdd.n3284 vdd.n338 146.341
R18745 vdd.n3280 vdd.n3279 146.341
R18746 vdd.n3277 vdd.n346 146.341
R18747 vdd.n3273 vdd.n3272 146.341
R18748 vdd.n3270 vdd.n353 146.341
R18749 vdd.n3266 vdd.n3265 146.341
R18750 vdd.n3263 vdd.n360 146.341
R18751 vdd.n371 vdd.n368 146.341
R18752 vdd.n3255 vdd.n3254 146.341
R18753 vdd.n3252 vdd.n373 146.341
R18754 vdd.n3248 vdd.n3247 146.341
R18755 vdd.n3245 vdd.n379 146.341
R18756 vdd.n3241 vdd.n3240 146.341
R18757 vdd.n3238 vdd.n386 146.341
R18758 vdd.n3234 vdd.n3233 146.341
R18759 vdd.n3231 vdd.n393 146.341
R18760 vdd.n3227 vdd.n3226 146.341
R18761 vdd.n3224 vdd.n400 146.341
R18762 vdd.n411 vdd.n408 146.341
R18763 vdd.n3216 vdd.n3215 146.341
R18764 vdd.n3213 vdd.n413 146.341
R18765 vdd.n3209 vdd.n3208 146.341
R18766 vdd.n3206 vdd.n419 146.341
R18767 vdd.n3202 vdd.n3201 146.341
R18768 vdd.n3199 vdd.n426 146.341
R18769 vdd.n3195 vdd.n3194 146.341
R18770 vdd.n3192 vdd.n433 146.341
R18771 vdd.n3188 vdd.n3187 146.341
R18772 vdd.n3185 vdd.n440 146.341
R18773 vdd.n3122 vdd.n478 146.341
R18774 vdd.n3122 vdd.n474 146.341
R18775 vdd.n3128 vdd.n474 146.341
R18776 vdd.n3128 vdd.n466 146.341
R18777 vdd.n3139 vdd.n466 146.341
R18778 vdd.n3139 vdd.n462 146.341
R18779 vdd.n3145 vdd.n462 146.341
R18780 vdd.n3145 vdd.n454 146.341
R18781 vdd.n3155 vdd.n454 146.341
R18782 vdd.n3155 vdd.n455 146.341
R18783 vdd.n455 vdd.n305 146.341
R18784 vdd.n306 vdd.n305 146.341
R18785 vdd.n307 vdd.n306 146.341
R18786 vdd.n448 vdd.n307 146.341
R18787 vdd.n448 vdd.n315 146.341
R18788 vdd.n316 vdd.n315 146.341
R18789 vdd.n317 vdd.n316 146.341
R18790 vdd.n445 vdd.n317 146.341
R18791 vdd.n445 vdd.n326 146.341
R18792 vdd.n327 vdd.n326 146.341
R18793 vdd.n328 vdd.n327 146.341
R18794 vdd.n3111 vdd.n483 146.341
R18795 vdd.n3111 vdd.n517 146.341
R18796 vdd.n523 vdd.n522 146.341
R18797 vdd.n3104 vdd.n3103 146.341
R18798 vdd.n3100 vdd.n3099 146.341
R18799 vdd.n3096 vdd.n3095 146.341
R18800 vdd.n3092 vdd.n3091 146.341
R18801 vdd.n3088 vdd.n3087 146.341
R18802 vdd.n3084 vdd.n3083 146.341
R18803 vdd.n3080 vdd.n3079 146.341
R18804 vdd.n3071 vdd.n3070 146.341
R18805 vdd.n3068 vdd.n3067 146.341
R18806 vdd.n3064 vdd.n3063 146.341
R18807 vdd.n3060 vdd.n3059 146.341
R18808 vdd.n3056 vdd.n3055 146.341
R18809 vdd.n3052 vdd.n3051 146.341
R18810 vdd.n3048 vdd.n3047 146.341
R18811 vdd.n3044 vdd.n3043 146.341
R18812 vdd.n3040 vdd.n3039 146.341
R18813 vdd.n3036 vdd.n3035 146.341
R18814 vdd.n3032 vdd.n3031 146.341
R18815 vdd.n3025 vdd.n3024 146.341
R18816 vdd.n3022 vdd.n3021 146.341
R18817 vdd.n3018 vdd.n3017 146.341
R18818 vdd.n3014 vdd.n3013 146.341
R18819 vdd.n3010 vdd.n3009 146.341
R18820 vdd.n3006 vdd.n3005 146.341
R18821 vdd.n3002 vdd.n3001 146.341
R18822 vdd.n2998 vdd.n2997 146.341
R18823 vdd.n2994 vdd.n2993 146.341
R18824 vdd.n2990 vdd.n2989 146.341
R18825 vdd.n2986 vdd.n515 146.341
R18826 vdd.n3120 vdd.n479 146.341
R18827 vdd.n3120 vdd.n472 146.341
R18828 vdd.n3131 vdd.n472 146.341
R18829 vdd.n3131 vdd.n468 146.341
R18830 vdd.n3137 vdd.n468 146.341
R18831 vdd.n3137 vdd.n461 146.341
R18832 vdd.n3147 vdd.n461 146.341
R18833 vdd.n3147 vdd.n457 146.341
R18834 vdd.n3153 vdd.n457 146.341
R18835 vdd.n3153 vdd.n302 146.341
R18836 vdd.n3316 vdd.n302 146.341
R18837 vdd.n3316 vdd.n303 146.341
R18838 vdd.n3312 vdd.n303 146.341
R18839 vdd.n3312 vdd.n309 146.341
R18840 vdd.n3308 vdd.n309 146.341
R18841 vdd.n3308 vdd.n314 146.341
R18842 vdd.n3304 vdd.n314 146.341
R18843 vdd.n3304 vdd.n319 146.341
R18844 vdd.n3300 vdd.n319 146.341
R18845 vdd.n3300 vdd.n325 146.341
R18846 vdd.n3296 vdd.n325 146.341
R18847 vdd.n2085 vdd.n2084 146.341
R18848 vdd.n2082 vdd.n2079 146.341
R18849 vdd.n2077 vdd.n975 146.341
R18850 vdd.n2073 vdd.n2072 146.341
R18851 vdd.n2070 vdd.n979 146.341
R18852 vdd.n2066 vdd.n2065 146.341
R18853 vdd.n2063 vdd.n986 146.341
R18854 vdd.n2059 vdd.n2058 146.341
R18855 vdd.n2056 vdd.n993 146.341
R18856 vdd.n1004 vdd.n1001 146.341
R18857 vdd.n2048 vdd.n2047 146.341
R18858 vdd.n2045 vdd.n1006 146.341
R18859 vdd.n2041 vdd.n2040 146.341
R18860 vdd.n2038 vdd.n1012 146.341
R18861 vdd.n2034 vdd.n2033 146.341
R18862 vdd.n2031 vdd.n1019 146.341
R18863 vdd.n2027 vdd.n2026 146.341
R18864 vdd.n2024 vdd.n1026 146.341
R18865 vdd.n2020 vdd.n2019 146.341
R18866 vdd.n2017 vdd.n1033 146.341
R18867 vdd.n1044 vdd.n1041 146.341
R18868 vdd.n2009 vdd.n2008 146.341
R18869 vdd.n2006 vdd.n1046 146.341
R18870 vdd.n2002 vdd.n2001 146.341
R18871 vdd.n1999 vdd.n1052 146.341
R18872 vdd.n1995 vdd.n1994 146.341
R18873 vdd.n1992 vdd.n1059 146.341
R18874 vdd.n1988 vdd.n1987 146.341
R18875 vdd.n1985 vdd.n1066 146.341
R18876 vdd.n1312 vdd.n1310 146.341
R18877 vdd.n1315 vdd.n1314 146.341
R18878 vdd.n1886 vdd.n1646 146.341
R18879 vdd.n1886 vdd.n1642 146.341
R18880 vdd.n1892 vdd.n1642 146.341
R18881 vdd.n1892 vdd.n1634 146.341
R18882 vdd.n1903 vdd.n1634 146.341
R18883 vdd.n1903 vdd.n1630 146.341
R18884 vdd.n1909 vdd.n1630 146.341
R18885 vdd.n1909 vdd.n1624 146.341
R18886 vdd.n1921 vdd.n1624 146.341
R18887 vdd.n1921 vdd.n1620 146.341
R18888 vdd.n1927 vdd.n1620 146.341
R18889 vdd.n1927 vdd.n1341 146.341
R18890 vdd.n1937 vdd.n1341 146.341
R18891 vdd.n1937 vdd.n1337 146.341
R18892 vdd.n1943 vdd.n1337 146.341
R18893 vdd.n1943 vdd.n1331 146.341
R18894 vdd.n1954 vdd.n1331 146.341
R18895 vdd.n1954 vdd.n1326 146.341
R18896 vdd.n1962 vdd.n1326 146.341
R18897 vdd.n1962 vdd.n1317 146.341
R18898 vdd.n1973 vdd.n1317 146.341
R18899 vdd.n1875 vdd.n1651 146.341
R18900 vdd.n1875 vdd.n1684 146.341
R18901 vdd.n1688 vdd.n1687 146.341
R18902 vdd.n1690 vdd.n1689 146.341
R18903 vdd.n1694 vdd.n1693 146.341
R18904 vdd.n1696 vdd.n1695 146.341
R18905 vdd.n1700 vdd.n1699 146.341
R18906 vdd.n1702 vdd.n1701 146.341
R18907 vdd.n1706 vdd.n1705 146.341
R18908 vdd.n1708 vdd.n1707 146.341
R18909 vdd.n1714 vdd.n1713 146.341
R18910 vdd.n1716 vdd.n1715 146.341
R18911 vdd.n1720 vdd.n1719 146.341
R18912 vdd.n1722 vdd.n1721 146.341
R18913 vdd.n1726 vdd.n1725 146.341
R18914 vdd.n1728 vdd.n1727 146.341
R18915 vdd.n1732 vdd.n1731 146.341
R18916 vdd.n1734 vdd.n1733 146.341
R18917 vdd.n1738 vdd.n1737 146.341
R18918 vdd.n1740 vdd.n1739 146.341
R18919 vdd.n1812 vdd.n1743 146.341
R18920 vdd.n1745 vdd.n1744 146.341
R18921 vdd.n1749 vdd.n1748 146.341
R18922 vdd.n1751 vdd.n1750 146.341
R18923 vdd.n1755 vdd.n1754 146.341
R18924 vdd.n1757 vdd.n1756 146.341
R18925 vdd.n1761 vdd.n1760 146.341
R18926 vdd.n1763 vdd.n1762 146.341
R18927 vdd.n1767 vdd.n1766 146.341
R18928 vdd.n1769 vdd.n1768 146.341
R18929 vdd.n1773 vdd.n1772 146.341
R18930 vdd.n1774 vdd.n1682 146.341
R18931 vdd.n1884 vdd.n1647 146.341
R18932 vdd.n1884 vdd.n1640 146.341
R18933 vdd.n1895 vdd.n1640 146.341
R18934 vdd.n1895 vdd.n1636 146.341
R18935 vdd.n1901 vdd.n1636 146.341
R18936 vdd.n1901 vdd.n1629 146.341
R18937 vdd.n1912 vdd.n1629 146.341
R18938 vdd.n1912 vdd.n1625 146.341
R18939 vdd.n1919 vdd.n1625 146.341
R18940 vdd.n1919 vdd.n1618 146.341
R18941 vdd.n1929 vdd.n1618 146.341
R18942 vdd.n1929 vdd.n1344 146.341
R18943 vdd.n1935 vdd.n1344 146.341
R18944 vdd.n1935 vdd.n1336 146.341
R18945 vdd.n1946 vdd.n1336 146.341
R18946 vdd.n1946 vdd.n1332 146.341
R18947 vdd.n1952 vdd.n1332 146.341
R18948 vdd.n1952 vdd.n1324 146.341
R18949 vdd.n1965 vdd.n1324 146.341
R18950 vdd.n1965 vdd.n1319 146.341
R18951 vdd.n1971 vdd.n1319 146.341
R18952 vdd.n1105 vdd.t23 127.284
R18953 vdd.n800 vdd.t67 127.284
R18954 vdd.n1109 vdd.t64 127.284
R18955 vdd.n791 vdd.t84 127.284
R18956 vdd.n686 vdd.t40 127.284
R18957 vdd.n686 vdd.t41 127.284
R18958 vdd.n2437 vdd.t82 127.284
R18959 vdd.n622 vdd.t32 127.284
R18960 vdd.n2434 vdd.t75 127.284
R18961 vdd.n589 vdd.t18 127.284
R18962 vdd.n861 vdd.t78 127.284
R18963 vdd.n861 vdd.t79 127.284
R18964 vdd.n22 vdd.n20 117.314
R18965 vdd.n17 vdd.n15 117.314
R18966 vdd.n27 vdd.n26 116.927
R18967 vdd.n24 vdd.n23 116.927
R18968 vdd.n22 vdd.n21 116.927
R18969 vdd.n17 vdd.n16 116.927
R18970 vdd.n19 vdd.n18 116.927
R18971 vdd.n27 vdd.n25 116.927
R18972 vdd.n1106 vdd.t22 111.188
R18973 vdd.n801 vdd.t68 111.188
R18974 vdd.n1110 vdd.t63 111.188
R18975 vdd.n792 vdd.t85 111.188
R18976 vdd.n2438 vdd.t81 111.188
R18977 vdd.n623 vdd.t33 111.188
R18978 vdd.n2435 vdd.t74 111.188
R18979 vdd.n590 vdd.t19 111.188
R18980 vdd.n2708 vdd.n750 99.5127
R18981 vdd.n2708 vdd.n741 99.5127
R18982 vdd.n2716 vdd.n741 99.5127
R18983 vdd.n2716 vdd.n739 99.5127
R18984 vdd.n2720 vdd.n739 99.5127
R18985 vdd.n2720 vdd.n729 99.5127
R18986 vdd.n2728 vdd.n729 99.5127
R18987 vdd.n2728 vdd.n727 99.5127
R18988 vdd.n2732 vdd.n727 99.5127
R18989 vdd.n2732 vdd.n718 99.5127
R18990 vdd.n2740 vdd.n718 99.5127
R18991 vdd.n2740 vdd.n716 99.5127
R18992 vdd.n2744 vdd.n716 99.5127
R18993 vdd.n2744 vdd.n707 99.5127
R18994 vdd.n2752 vdd.n707 99.5127
R18995 vdd.n2752 vdd.n705 99.5127
R18996 vdd.n2756 vdd.n705 99.5127
R18997 vdd.n2756 vdd.n694 99.5127
R18998 vdd.n2765 vdd.n694 99.5127
R18999 vdd.n2765 vdd.n692 99.5127
R19000 vdd.n2769 vdd.n692 99.5127
R19001 vdd.n2769 vdd.n682 99.5127
R19002 vdd.n2777 vdd.n682 99.5127
R19003 vdd.n2777 vdd.n680 99.5127
R19004 vdd.n2781 vdd.n680 99.5127
R19005 vdd.n2781 vdd.n670 99.5127
R19006 vdd.n2789 vdd.n670 99.5127
R19007 vdd.n2789 vdd.n668 99.5127
R19008 vdd.n2793 vdd.n668 99.5127
R19009 vdd.n2793 vdd.n657 99.5127
R19010 vdd.n2801 vdd.n657 99.5127
R19011 vdd.n2801 vdd.n655 99.5127
R19012 vdd.n2805 vdd.n655 99.5127
R19013 vdd.n2805 vdd.n646 99.5127
R19014 vdd.n2813 vdd.n646 99.5127
R19015 vdd.n2813 vdd.n644 99.5127
R19016 vdd.n2817 vdd.n644 99.5127
R19017 vdd.n2817 vdd.n632 99.5127
R19018 vdd.n2870 vdd.n632 99.5127
R19019 vdd.n2870 vdd.n630 99.5127
R19020 vdd.n2874 vdd.n630 99.5127
R19021 vdd.n2874 vdd.n598 99.5127
R19022 vdd.n2944 vdd.n598 99.5127
R19023 vdd.n2940 vdd.n599 99.5127
R19024 vdd.n2938 vdd.n2937 99.5127
R19025 vdd.n2935 vdd.n603 99.5127
R19026 vdd.n2931 vdd.n2930 99.5127
R19027 vdd.n2928 vdd.n606 99.5127
R19028 vdd.n2924 vdd.n2923 99.5127
R19029 vdd.n2921 vdd.n609 99.5127
R19030 vdd.n2917 vdd.n2916 99.5127
R19031 vdd.n2914 vdd.n2912 99.5127
R19032 vdd.n2910 vdd.n612 99.5127
R19033 vdd.n2906 vdd.n2905 99.5127
R19034 vdd.n2903 vdd.n615 99.5127
R19035 vdd.n2899 vdd.n2898 99.5127
R19036 vdd.n2896 vdd.n618 99.5127
R19037 vdd.n2892 vdd.n2891 99.5127
R19038 vdd.n2889 vdd.n621 99.5127
R19039 vdd.n2884 vdd.n2883 99.5127
R19040 vdd.n2635 vdd.n748 99.5127
R19041 vdd.n2631 vdd.n748 99.5127
R19042 vdd.n2631 vdd.n742 99.5127
R19043 vdd.n2513 vdd.n742 99.5127
R19044 vdd.n2513 vdd.n737 99.5127
R19045 vdd.n2516 vdd.n737 99.5127
R19046 vdd.n2516 vdd.n731 99.5127
R19047 vdd.n2617 vdd.n731 99.5127
R19048 vdd.n2617 vdd.n725 99.5127
R19049 vdd.n2613 vdd.n725 99.5127
R19050 vdd.n2613 vdd.n719 99.5127
R19051 vdd.n2560 vdd.n719 99.5127
R19052 vdd.n2560 vdd.n713 99.5127
R19053 vdd.n2557 vdd.n713 99.5127
R19054 vdd.n2557 vdd.n708 99.5127
R19055 vdd.n2554 vdd.n708 99.5127
R19056 vdd.n2554 vdd.n703 99.5127
R19057 vdd.n2551 vdd.n703 99.5127
R19058 vdd.n2551 vdd.n696 99.5127
R19059 vdd.n2548 vdd.n696 99.5127
R19060 vdd.n2548 vdd.n689 99.5127
R19061 vdd.n2545 vdd.n689 99.5127
R19062 vdd.n2545 vdd.n683 99.5127
R19063 vdd.n2542 vdd.n683 99.5127
R19064 vdd.n2542 vdd.n678 99.5127
R19065 vdd.n2539 vdd.n678 99.5127
R19066 vdd.n2539 vdd.n672 99.5127
R19067 vdd.n2536 vdd.n672 99.5127
R19068 vdd.n2536 vdd.n665 99.5127
R19069 vdd.n2533 vdd.n665 99.5127
R19070 vdd.n2533 vdd.n658 99.5127
R19071 vdd.n2530 vdd.n658 99.5127
R19072 vdd.n2530 vdd.n652 99.5127
R19073 vdd.n2527 vdd.n652 99.5127
R19074 vdd.n2527 vdd.n647 99.5127
R19075 vdd.n2524 vdd.n647 99.5127
R19076 vdd.n2524 vdd.n642 99.5127
R19077 vdd.n2521 vdd.n642 99.5127
R19078 vdd.n2521 vdd.n634 99.5127
R19079 vdd.n634 vdd.n627 99.5127
R19080 vdd.n2876 vdd.n627 99.5127
R19081 vdd.n2877 vdd.n2876 99.5127
R19082 vdd.n2877 vdd.n596 99.5127
R19083 vdd.n2701 vdd.n752 99.5127
R19084 vdd.n2701 vdd.n2433 99.5127
R19085 vdd.n2697 vdd.n2696 99.5127
R19086 vdd.n2693 vdd.n2692 99.5127
R19087 vdd.n2689 vdd.n2688 99.5127
R19088 vdd.n2685 vdd.n2684 99.5127
R19089 vdd.n2681 vdd.n2680 99.5127
R19090 vdd.n2677 vdd.n2676 99.5127
R19091 vdd.n2673 vdd.n2672 99.5127
R19092 vdd.n2669 vdd.n2668 99.5127
R19093 vdd.n2665 vdd.n2664 99.5127
R19094 vdd.n2661 vdd.n2660 99.5127
R19095 vdd.n2657 vdd.n2656 99.5127
R19096 vdd.n2653 vdd.n2652 99.5127
R19097 vdd.n2649 vdd.n2648 99.5127
R19098 vdd.n2645 vdd.n2644 99.5127
R19099 vdd.n2640 vdd.n2639 99.5127
R19100 vdd.n2397 vdd.n789 99.5127
R19101 vdd.n2393 vdd.n2392 99.5127
R19102 vdd.n2389 vdd.n2388 99.5127
R19103 vdd.n2385 vdd.n2384 99.5127
R19104 vdd.n2381 vdd.n2380 99.5127
R19105 vdd.n2377 vdd.n2376 99.5127
R19106 vdd.n2373 vdd.n2372 99.5127
R19107 vdd.n2369 vdd.n2368 99.5127
R19108 vdd.n2365 vdd.n2364 99.5127
R19109 vdd.n2361 vdd.n2360 99.5127
R19110 vdd.n2357 vdd.n2356 99.5127
R19111 vdd.n2353 vdd.n2352 99.5127
R19112 vdd.n2349 vdd.n2348 99.5127
R19113 vdd.n2345 vdd.n2344 99.5127
R19114 vdd.n2341 vdd.n2340 99.5127
R19115 vdd.n2337 vdd.n2336 99.5127
R19116 vdd.n2332 vdd.n2331 99.5127
R19117 vdd.n1145 vdd.n925 99.5127
R19118 vdd.n1148 vdd.n925 99.5127
R19119 vdd.n1148 vdd.n919 99.5127
R19120 vdd.n1151 vdd.n919 99.5127
R19121 vdd.n1151 vdd.n914 99.5127
R19122 vdd.n1154 vdd.n914 99.5127
R19123 vdd.n1154 vdd.n907 99.5127
R19124 vdd.n1157 vdd.n907 99.5127
R19125 vdd.n1157 vdd.n900 99.5127
R19126 vdd.n1160 vdd.n900 99.5127
R19127 vdd.n1160 vdd.n894 99.5127
R19128 vdd.n1163 vdd.n894 99.5127
R19129 vdd.n1163 vdd.n889 99.5127
R19130 vdd.n1166 vdd.n889 99.5127
R19131 vdd.n1166 vdd.n884 99.5127
R19132 vdd.n1169 vdd.n884 99.5127
R19133 vdd.n1169 vdd.n878 99.5127
R19134 vdd.n1172 vdd.n878 99.5127
R19135 vdd.n1172 vdd.n871 99.5127
R19136 vdd.n1175 vdd.n871 99.5127
R19137 vdd.n1175 vdd.n864 99.5127
R19138 vdd.n1178 vdd.n864 99.5127
R19139 vdd.n1178 vdd.n858 99.5127
R19140 vdd.n1181 vdd.n858 99.5127
R19141 vdd.n1181 vdd.n853 99.5127
R19142 vdd.n1184 vdd.n853 99.5127
R19143 vdd.n1184 vdd.n847 99.5127
R19144 vdd.n1226 vdd.n847 99.5127
R19145 vdd.n1226 vdd.n840 99.5127
R19146 vdd.n1222 vdd.n840 99.5127
R19147 vdd.n1222 vdd.n834 99.5127
R19148 vdd.n1219 vdd.n834 99.5127
R19149 vdd.n1219 vdd.n829 99.5127
R19150 vdd.n1216 vdd.n829 99.5127
R19151 vdd.n1216 vdd.n824 99.5127
R19152 vdd.n1196 vdd.n824 99.5127
R19153 vdd.n1196 vdd.n819 99.5127
R19154 vdd.n1193 vdd.n819 99.5127
R19155 vdd.n1193 vdd.n812 99.5127
R19156 vdd.n1190 vdd.n812 99.5127
R19157 vdd.n1190 vdd.n805 99.5127
R19158 vdd.n805 vdd.n794 99.5127
R19159 vdd.n2327 vdd.n794 99.5127
R19160 vdd.n2119 vdd.n930 99.5127
R19161 vdd.n2119 vdd.n966 99.5127
R19162 vdd.n2115 vdd.n2114 99.5127
R19163 vdd.n2111 vdd.n2110 99.5127
R19164 vdd.n2107 vdd.n2106 99.5127
R19165 vdd.n2103 vdd.n2102 99.5127
R19166 vdd.n2099 vdd.n2098 99.5127
R19167 vdd.n2095 vdd.n2094 99.5127
R19168 vdd.n2091 vdd.n2090 99.5127
R19169 vdd.n1112 vdd.n1111 99.5127
R19170 vdd.n1116 vdd.n1115 99.5127
R19171 vdd.n1120 vdd.n1119 99.5127
R19172 vdd.n1124 vdd.n1123 99.5127
R19173 vdd.n1128 vdd.n1127 99.5127
R19174 vdd.n1132 vdd.n1131 99.5127
R19175 vdd.n1136 vdd.n1135 99.5127
R19176 vdd.n1141 vdd.n1140 99.5127
R19177 vdd.n2126 vdd.n928 99.5127
R19178 vdd.n2126 vdd.n918 99.5127
R19179 vdd.n2134 vdd.n918 99.5127
R19180 vdd.n2134 vdd.n916 99.5127
R19181 vdd.n2138 vdd.n916 99.5127
R19182 vdd.n2138 vdd.n905 99.5127
R19183 vdd.n2146 vdd.n905 99.5127
R19184 vdd.n2146 vdd.n903 99.5127
R19185 vdd.n2150 vdd.n903 99.5127
R19186 vdd.n2150 vdd.n893 99.5127
R19187 vdd.n2158 vdd.n893 99.5127
R19188 vdd.n2158 vdd.n891 99.5127
R19189 vdd.n2162 vdd.n891 99.5127
R19190 vdd.n2162 vdd.n882 99.5127
R19191 vdd.n2170 vdd.n882 99.5127
R19192 vdd.n2170 vdd.n880 99.5127
R19193 vdd.n2174 vdd.n880 99.5127
R19194 vdd.n2174 vdd.n869 99.5127
R19195 vdd.n2182 vdd.n869 99.5127
R19196 vdd.n2182 vdd.n867 99.5127
R19197 vdd.n2186 vdd.n867 99.5127
R19198 vdd.n2186 vdd.n857 99.5127
R19199 vdd.n2195 vdd.n857 99.5127
R19200 vdd.n2195 vdd.n855 99.5127
R19201 vdd.n2199 vdd.n855 99.5127
R19202 vdd.n2199 vdd.n845 99.5127
R19203 vdd.n2207 vdd.n845 99.5127
R19204 vdd.n2207 vdd.n843 99.5127
R19205 vdd.n2211 vdd.n843 99.5127
R19206 vdd.n2211 vdd.n833 99.5127
R19207 vdd.n2219 vdd.n833 99.5127
R19208 vdd.n2219 vdd.n831 99.5127
R19209 vdd.n2223 vdd.n831 99.5127
R19210 vdd.n2223 vdd.n823 99.5127
R19211 vdd.n2231 vdd.n823 99.5127
R19212 vdd.n2231 vdd.n821 99.5127
R19213 vdd.n2235 vdd.n821 99.5127
R19214 vdd.n2235 vdd.n810 99.5127
R19215 vdd.n2245 vdd.n810 99.5127
R19216 vdd.n2245 vdd.n807 99.5127
R19217 vdd.n2250 vdd.n807 99.5127
R19218 vdd.n2250 vdd.n808 99.5127
R19219 vdd.n808 vdd.n788 99.5127
R19220 vdd.n2860 vdd.n2859 99.5127
R19221 vdd.n2857 vdd.n2823 99.5127
R19222 vdd.n2853 vdd.n2852 99.5127
R19223 vdd.n2850 vdd.n2826 99.5127
R19224 vdd.n2846 vdd.n2845 99.5127
R19225 vdd.n2843 vdd.n2829 99.5127
R19226 vdd.n2839 vdd.n2838 99.5127
R19227 vdd.n2836 vdd.n2833 99.5127
R19228 vdd.n2977 vdd.n577 99.5127
R19229 vdd.n2975 vdd.n2974 99.5127
R19230 vdd.n2972 vdd.n579 99.5127
R19231 vdd.n2968 vdd.n2967 99.5127
R19232 vdd.n2965 vdd.n582 99.5127
R19233 vdd.n2961 vdd.n2960 99.5127
R19234 vdd.n2958 vdd.n585 99.5127
R19235 vdd.n2954 vdd.n2953 99.5127
R19236 vdd.n2951 vdd.n588 99.5127
R19237 vdd.n2509 vdd.n749 99.5127
R19238 vdd.n2629 vdd.n749 99.5127
R19239 vdd.n2629 vdd.n743 99.5127
R19240 vdd.n2625 vdd.n743 99.5127
R19241 vdd.n2625 vdd.n738 99.5127
R19242 vdd.n2622 vdd.n738 99.5127
R19243 vdd.n2622 vdd.n732 99.5127
R19244 vdd.n2619 vdd.n732 99.5127
R19245 vdd.n2619 vdd.n726 99.5127
R19246 vdd.n2611 vdd.n726 99.5127
R19247 vdd.n2611 vdd.n720 99.5127
R19248 vdd.n2607 vdd.n720 99.5127
R19249 vdd.n2607 vdd.n714 99.5127
R19250 vdd.n2604 vdd.n714 99.5127
R19251 vdd.n2604 vdd.n709 99.5127
R19252 vdd.n2601 vdd.n709 99.5127
R19253 vdd.n2601 vdd.n704 99.5127
R19254 vdd.n2598 vdd.n704 99.5127
R19255 vdd.n2598 vdd.n697 99.5127
R19256 vdd.n2595 vdd.n697 99.5127
R19257 vdd.n2595 vdd.n690 99.5127
R19258 vdd.n2592 vdd.n690 99.5127
R19259 vdd.n2592 vdd.n684 99.5127
R19260 vdd.n2589 vdd.n684 99.5127
R19261 vdd.n2589 vdd.n679 99.5127
R19262 vdd.n2586 vdd.n679 99.5127
R19263 vdd.n2586 vdd.n673 99.5127
R19264 vdd.n2583 vdd.n673 99.5127
R19265 vdd.n2583 vdd.n666 99.5127
R19266 vdd.n2580 vdd.n666 99.5127
R19267 vdd.n2580 vdd.n659 99.5127
R19268 vdd.n2577 vdd.n659 99.5127
R19269 vdd.n2577 vdd.n653 99.5127
R19270 vdd.n2574 vdd.n653 99.5127
R19271 vdd.n2574 vdd.n648 99.5127
R19272 vdd.n2571 vdd.n648 99.5127
R19273 vdd.n2571 vdd.n643 99.5127
R19274 vdd.n2568 vdd.n643 99.5127
R19275 vdd.n2568 vdd.n635 99.5127
R19276 vdd.n2565 vdd.n635 99.5127
R19277 vdd.n2565 vdd.n628 99.5127
R19278 vdd.n628 vdd.n594 99.5127
R19279 vdd.n2946 vdd.n594 99.5127
R19280 vdd.n2444 vdd.n2443 99.5127
R19281 vdd.n2448 vdd.n2447 99.5127
R19282 vdd.n2452 vdd.n2451 99.5127
R19283 vdd.n2456 vdd.n2455 99.5127
R19284 vdd.n2460 vdd.n2459 99.5127
R19285 vdd.n2464 vdd.n2463 99.5127
R19286 vdd.n2468 vdd.n2467 99.5127
R19287 vdd.n2472 vdd.n2471 99.5127
R19288 vdd.n2476 vdd.n2475 99.5127
R19289 vdd.n2480 vdd.n2479 99.5127
R19290 vdd.n2484 vdd.n2483 99.5127
R19291 vdd.n2488 vdd.n2487 99.5127
R19292 vdd.n2492 vdd.n2491 99.5127
R19293 vdd.n2496 vdd.n2495 99.5127
R19294 vdd.n2500 vdd.n2499 99.5127
R19295 vdd.n2504 vdd.n2503 99.5127
R19296 vdd.n2506 vdd.n2432 99.5127
R19297 vdd.n2710 vdd.n746 99.5127
R19298 vdd.n2710 vdd.n744 99.5127
R19299 vdd.n2714 vdd.n744 99.5127
R19300 vdd.n2714 vdd.n735 99.5127
R19301 vdd.n2722 vdd.n735 99.5127
R19302 vdd.n2722 vdd.n733 99.5127
R19303 vdd.n2726 vdd.n733 99.5127
R19304 vdd.n2726 vdd.n724 99.5127
R19305 vdd.n2734 vdd.n724 99.5127
R19306 vdd.n2734 vdd.n722 99.5127
R19307 vdd.n2738 vdd.n722 99.5127
R19308 vdd.n2738 vdd.n712 99.5127
R19309 vdd.n2746 vdd.n712 99.5127
R19310 vdd.n2746 vdd.n710 99.5127
R19311 vdd.n2750 vdd.n710 99.5127
R19312 vdd.n2750 vdd.n701 99.5127
R19313 vdd.n2758 vdd.n701 99.5127
R19314 vdd.n2758 vdd.n699 99.5127
R19315 vdd.n2763 vdd.n699 99.5127
R19316 vdd.n2763 vdd.n688 99.5127
R19317 vdd.n2771 vdd.n688 99.5127
R19318 vdd.n2771 vdd.n685 99.5127
R19319 vdd.n2775 vdd.n685 99.5127
R19320 vdd.n2775 vdd.n676 99.5127
R19321 vdd.n2783 vdd.n676 99.5127
R19322 vdd.n2783 vdd.n674 99.5127
R19323 vdd.n2787 vdd.n674 99.5127
R19324 vdd.n2787 vdd.n663 99.5127
R19325 vdd.n2795 vdd.n663 99.5127
R19326 vdd.n2795 vdd.n661 99.5127
R19327 vdd.n2799 vdd.n661 99.5127
R19328 vdd.n2799 vdd.n651 99.5127
R19329 vdd.n2807 vdd.n651 99.5127
R19330 vdd.n2807 vdd.n649 99.5127
R19331 vdd.n2811 vdd.n649 99.5127
R19332 vdd.n2811 vdd.n640 99.5127
R19333 vdd.n2819 vdd.n640 99.5127
R19334 vdd.n2819 vdd.n637 99.5127
R19335 vdd.n2868 vdd.n637 99.5127
R19336 vdd.n2868 vdd.n638 99.5127
R19337 vdd.n638 vdd.n629 99.5127
R19338 vdd.n2863 vdd.n629 99.5127
R19339 vdd.n2863 vdd.n597 99.5127
R19340 vdd.n2321 vdd.n2320 99.5127
R19341 vdd.n2317 vdd.n2316 99.5127
R19342 vdd.n2313 vdd.n2312 99.5127
R19343 vdd.n2309 vdd.n2308 99.5127
R19344 vdd.n2305 vdd.n2304 99.5127
R19345 vdd.n2301 vdd.n2300 99.5127
R19346 vdd.n2297 vdd.n2296 99.5127
R19347 vdd.n2293 vdd.n2292 99.5127
R19348 vdd.n2289 vdd.n2288 99.5127
R19349 vdd.n2285 vdd.n2284 99.5127
R19350 vdd.n2281 vdd.n2280 99.5127
R19351 vdd.n2277 vdd.n2276 99.5127
R19352 vdd.n2273 vdd.n2272 99.5127
R19353 vdd.n2269 vdd.n2268 99.5127
R19354 vdd.n2265 vdd.n2264 99.5127
R19355 vdd.n2261 vdd.n2260 99.5127
R19356 vdd.n2257 vdd.n770 99.5127
R19357 vdd.n1270 vdd.n926 99.5127
R19358 vdd.n1267 vdd.n926 99.5127
R19359 vdd.n1267 vdd.n920 99.5127
R19360 vdd.n1264 vdd.n920 99.5127
R19361 vdd.n1264 vdd.n915 99.5127
R19362 vdd.n1261 vdd.n915 99.5127
R19363 vdd.n1261 vdd.n908 99.5127
R19364 vdd.n1258 vdd.n908 99.5127
R19365 vdd.n1258 vdd.n901 99.5127
R19366 vdd.n1255 vdd.n901 99.5127
R19367 vdd.n1255 vdd.n895 99.5127
R19368 vdd.n1252 vdd.n895 99.5127
R19369 vdd.n1252 vdd.n890 99.5127
R19370 vdd.n1249 vdd.n890 99.5127
R19371 vdd.n1249 vdd.n885 99.5127
R19372 vdd.n1246 vdd.n885 99.5127
R19373 vdd.n1246 vdd.n879 99.5127
R19374 vdd.n1243 vdd.n879 99.5127
R19375 vdd.n1243 vdd.n872 99.5127
R19376 vdd.n1240 vdd.n872 99.5127
R19377 vdd.n1240 vdd.n865 99.5127
R19378 vdd.n1237 vdd.n865 99.5127
R19379 vdd.n1237 vdd.n859 99.5127
R19380 vdd.n1234 vdd.n859 99.5127
R19381 vdd.n1234 vdd.n854 99.5127
R19382 vdd.n1231 vdd.n854 99.5127
R19383 vdd.n1231 vdd.n848 99.5127
R19384 vdd.n1228 vdd.n848 99.5127
R19385 vdd.n1228 vdd.n841 99.5127
R19386 vdd.n1199 vdd.n841 99.5127
R19387 vdd.n1199 vdd.n835 99.5127
R19388 vdd.n1202 vdd.n835 99.5127
R19389 vdd.n1202 vdd.n830 99.5127
R19390 vdd.n1214 vdd.n830 99.5127
R19391 vdd.n1214 vdd.n825 99.5127
R19392 vdd.n1210 vdd.n825 99.5127
R19393 vdd.n1210 vdd.n820 99.5127
R19394 vdd.n1207 vdd.n820 99.5127
R19395 vdd.n1207 vdd.n813 99.5127
R19396 vdd.n813 vdd.n804 99.5127
R19397 vdd.n2252 vdd.n804 99.5127
R19398 vdd.n2253 vdd.n2252 99.5127
R19399 vdd.n2253 vdd.n796 99.5127
R19400 vdd.n1074 vdd.n1073 99.5127
R19401 vdd.n1078 vdd.n1077 99.5127
R19402 vdd.n1082 vdd.n1081 99.5127
R19403 vdd.n1086 vdd.n1085 99.5127
R19404 vdd.n1090 vdd.n1089 99.5127
R19405 vdd.n1094 vdd.n1093 99.5127
R19406 vdd.n1098 vdd.n1097 99.5127
R19407 vdd.n1102 vdd.n1101 99.5127
R19408 vdd.n1303 vdd.n1104 99.5127
R19409 vdd.n1301 vdd.n1300 99.5127
R19410 vdd.n1297 vdd.n1296 99.5127
R19411 vdd.n1293 vdd.n1292 99.5127
R19412 vdd.n1289 vdd.n1288 99.5127
R19413 vdd.n1285 vdd.n1284 99.5127
R19414 vdd.n1281 vdd.n1280 99.5127
R19415 vdd.n1277 vdd.n1276 99.5127
R19416 vdd.n1273 vdd.n965 99.5127
R19417 vdd.n2128 vdd.n923 99.5127
R19418 vdd.n2128 vdd.n921 99.5127
R19419 vdd.n2132 vdd.n921 99.5127
R19420 vdd.n2132 vdd.n912 99.5127
R19421 vdd.n2140 vdd.n912 99.5127
R19422 vdd.n2140 vdd.n910 99.5127
R19423 vdd.n2144 vdd.n910 99.5127
R19424 vdd.n2144 vdd.n899 99.5127
R19425 vdd.n2152 vdd.n899 99.5127
R19426 vdd.n2152 vdd.n897 99.5127
R19427 vdd.n2156 vdd.n897 99.5127
R19428 vdd.n2156 vdd.n888 99.5127
R19429 vdd.n2164 vdd.n888 99.5127
R19430 vdd.n2164 vdd.n886 99.5127
R19431 vdd.n2168 vdd.n886 99.5127
R19432 vdd.n2168 vdd.n876 99.5127
R19433 vdd.n2176 vdd.n876 99.5127
R19434 vdd.n2176 vdd.n874 99.5127
R19435 vdd.n2180 vdd.n874 99.5127
R19436 vdd.n2180 vdd.n863 99.5127
R19437 vdd.n2188 vdd.n863 99.5127
R19438 vdd.n2188 vdd.n860 99.5127
R19439 vdd.n2193 vdd.n860 99.5127
R19440 vdd.n2193 vdd.n851 99.5127
R19441 vdd.n2201 vdd.n851 99.5127
R19442 vdd.n2201 vdd.n849 99.5127
R19443 vdd.n2205 vdd.n849 99.5127
R19444 vdd.n2205 vdd.n839 99.5127
R19445 vdd.n2213 vdd.n839 99.5127
R19446 vdd.n2213 vdd.n837 99.5127
R19447 vdd.n2217 vdd.n837 99.5127
R19448 vdd.n2217 vdd.n828 99.5127
R19449 vdd.n2225 vdd.n828 99.5127
R19450 vdd.n2225 vdd.n826 99.5127
R19451 vdd.n2229 vdd.n826 99.5127
R19452 vdd.n2229 vdd.n817 99.5127
R19453 vdd.n2237 vdd.n817 99.5127
R19454 vdd.n2237 vdd.n814 99.5127
R19455 vdd.n2243 vdd.n814 99.5127
R19456 vdd.n2243 vdd.n815 99.5127
R19457 vdd.n815 vdd.n806 99.5127
R19458 vdd.n806 vdd.n797 99.5127
R19459 vdd.n2325 vdd.n797 99.5127
R19460 vdd.n9 vdd.n7 98.9633
R19461 vdd.n2 vdd.n0 98.9633
R19462 vdd.n9 vdd.n8 98.6055
R19463 vdd.n11 vdd.n10 98.6055
R19464 vdd.n13 vdd.n12 98.6055
R19465 vdd.n6 vdd.n5 98.6055
R19466 vdd.n4 vdd.n3 98.6055
R19467 vdd.n2 vdd.n1 98.6055
R19468 vdd.t145 vdd.n267 85.8723
R19469 vdd.t153 vdd.n220 85.8723
R19470 vdd.t142 vdd.n177 85.8723
R19471 vdd.t150 vdd.n130 85.8723
R19472 vdd.t122 vdd.n88 85.8723
R19473 vdd.t127 vdd.n41 85.8723
R19474 vdd.t120 vdd.n1537 85.8723
R19475 vdd.t106 vdd.n1584 85.8723
R19476 vdd.t115 vdd.n1447 85.8723
R19477 vdd.t95 vdd.n1494 85.8723
R19478 vdd.t128 vdd.n1358 85.8723
R19479 vdd.t123 vdd.n1405 85.8723
R19480 vdd.n687 vdd.n686 78.546
R19481 vdd.n2191 vdd.n861 78.546
R19482 vdd.n254 vdd.n253 75.1835
R19483 vdd.n252 vdd.n251 75.1835
R19484 vdd.n250 vdd.n249 75.1835
R19485 vdd.n164 vdd.n163 75.1835
R19486 vdd.n162 vdd.n161 75.1835
R19487 vdd.n160 vdd.n159 75.1835
R19488 vdd.n75 vdd.n74 75.1835
R19489 vdd.n73 vdd.n72 75.1835
R19490 vdd.n71 vdd.n70 75.1835
R19491 vdd.n1567 vdd.n1566 75.1835
R19492 vdd.n1569 vdd.n1568 75.1835
R19493 vdd.n1571 vdd.n1570 75.1835
R19494 vdd.n1477 vdd.n1476 75.1835
R19495 vdd.n1479 vdd.n1478 75.1835
R19496 vdd.n1481 vdd.n1480 75.1835
R19497 vdd.n1388 vdd.n1387 75.1835
R19498 vdd.n1390 vdd.n1389 75.1835
R19499 vdd.n1392 vdd.n1391 75.1835
R19500 vdd.n2702 vdd.n2415 72.8958
R19501 vdd.n2702 vdd.n2416 72.8958
R19502 vdd.n2702 vdd.n2417 72.8958
R19503 vdd.n2702 vdd.n2418 72.8958
R19504 vdd.n2702 vdd.n2419 72.8958
R19505 vdd.n2702 vdd.n2420 72.8958
R19506 vdd.n2702 vdd.n2421 72.8958
R19507 vdd.n2702 vdd.n2422 72.8958
R19508 vdd.n2702 vdd.n2423 72.8958
R19509 vdd.n2702 vdd.n2424 72.8958
R19510 vdd.n2702 vdd.n2425 72.8958
R19511 vdd.n2702 vdd.n2426 72.8958
R19512 vdd.n2702 vdd.n2427 72.8958
R19513 vdd.n2702 vdd.n2428 72.8958
R19514 vdd.n2702 vdd.n2429 72.8958
R19515 vdd.n2702 vdd.n2430 72.8958
R19516 vdd.n2702 vdd.n2431 72.8958
R19517 vdd.n593 vdd.n484 72.8958
R19518 vdd.n2952 vdd.n484 72.8958
R19519 vdd.n587 vdd.n484 72.8958
R19520 vdd.n2959 vdd.n484 72.8958
R19521 vdd.n584 vdd.n484 72.8958
R19522 vdd.n2966 vdd.n484 72.8958
R19523 vdd.n581 vdd.n484 72.8958
R19524 vdd.n2973 vdd.n484 72.8958
R19525 vdd.n2976 vdd.n484 72.8958
R19526 vdd.n2832 vdd.n484 72.8958
R19527 vdd.n2837 vdd.n484 72.8958
R19528 vdd.n2831 vdd.n484 72.8958
R19529 vdd.n2844 vdd.n484 72.8958
R19530 vdd.n2828 vdd.n484 72.8958
R19531 vdd.n2851 vdd.n484 72.8958
R19532 vdd.n2825 vdd.n484 72.8958
R19533 vdd.n2858 vdd.n484 72.8958
R19534 vdd.n2121 vdd.n2120 72.8958
R19535 vdd.n2120 vdd.n932 72.8958
R19536 vdd.n2120 vdd.n933 72.8958
R19537 vdd.n2120 vdd.n934 72.8958
R19538 vdd.n2120 vdd.n935 72.8958
R19539 vdd.n2120 vdd.n936 72.8958
R19540 vdd.n2120 vdd.n937 72.8958
R19541 vdd.n2120 vdd.n938 72.8958
R19542 vdd.n2120 vdd.n939 72.8958
R19543 vdd.n2120 vdd.n940 72.8958
R19544 vdd.n2120 vdd.n941 72.8958
R19545 vdd.n2120 vdd.n942 72.8958
R19546 vdd.n2120 vdd.n943 72.8958
R19547 vdd.n2120 vdd.n944 72.8958
R19548 vdd.n2120 vdd.n945 72.8958
R19549 vdd.n2120 vdd.n946 72.8958
R19550 vdd.n2120 vdd.n947 72.8958
R19551 vdd.n2398 vdd.n771 72.8958
R19552 vdd.n2398 vdd.n772 72.8958
R19553 vdd.n2398 vdd.n773 72.8958
R19554 vdd.n2398 vdd.n774 72.8958
R19555 vdd.n2398 vdd.n775 72.8958
R19556 vdd.n2398 vdd.n776 72.8958
R19557 vdd.n2398 vdd.n777 72.8958
R19558 vdd.n2398 vdd.n778 72.8958
R19559 vdd.n2398 vdd.n779 72.8958
R19560 vdd.n2398 vdd.n780 72.8958
R19561 vdd.n2398 vdd.n781 72.8958
R19562 vdd.n2398 vdd.n782 72.8958
R19563 vdd.n2398 vdd.n783 72.8958
R19564 vdd.n2398 vdd.n784 72.8958
R19565 vdd.n2398 vdd.n785 72.8958
R19566 vdd.n2398 vdd.n786 72.8958
R19567 vdd.n2398 vdd.n787 72.8958
R19568 vdd.n2703 vdd.n2702 72.8958
R19569 vdd.n2702 vdd.n2399 72.8958
R19570 vdd.n2702 vdd.n2400 72.8958
R19571 vdd.n2702 vdd.n2401 72.8958
R19572 vdd.n2702 vdd.n2402 72.8958
R19573 vdd.n2702 vdd.n2403 72.8958
R19574 vdd.n2702 vdd.n2404 72.8958
R19575 vdd.n2702 vdd.n2405 72.8958
R19576 vdd.n2702 vdd.n2406 72.8958
R19577 vdd.n2702 vdd.n2407 72.8958
R19578 vdd.n2702 vdd.n2408 72.8958
R19579 vdd.n2702 vdd.n2409 72.8958
R19580 vdd.n2702 vdd.n2410 72.8958
R19581 vdd.n2702 vdd.n2411 72.8958
R19582 vdd.n2702 vdd.n2412 72.8958
R19583 vdd.n2702 vdd.n2413 72.8958
R19584 vdd.n2702 vdd.n2414 72.8958
R19585 vdd.n2882 vdd.n484 72.8958
R19586 vdd.n625 vdd.n484 72.8958
R19587 vdd.n2890 vdd.n484 72.8958
R19588 vdd.n620 vdd.n484 72.8958
R19589 vdd.n2897 vdd.n484 72.8958
R19590 vdd.n617 vdd.n484 72.8958
R19591 vdd.n2904 vdd.n484 72.8958
R19592 vdd.n614 vdd.n484 72.8958
R19593 vdd.n2911 vdd.n484 72.8958
R19594 vdd.n2915 vdd.n484 72.8958
R19595 vdd.n611 vdd.n484 72.8958
R19596 vdd.n2922 vdd.n484 72.8958
R19597 vdd.n608 vdd.n484 72.8958
R19598 vdd.n2929 vdd.n484 72.8958
R19599 vdd.n605 vdd.n484 72.8958
R19600 vdd.n2936 vdd.n484 72.8958
R19601 vdd.n2939 vdd.n484 72.8958
R19602 vdd.n2398 vdd.n769 72.8958
R19603 vdd.n2398 vdd.n768 72.8958
R19604 vdd.n2398 vdd.n767 72.8958
R19605 vdd.n2398 vdd.n766 72.8958
R19606 vdd.n2398 vdd.n765 72.8958
R19607 vdd.n2398 vdd.n764 72.8958
R19608 vdd.n2398 vdd.n763 72.8958
R19609 vdd.n2398 vdd.n762 72.8958
R19610 vdd.n2398 vdd.n761 72.8958
R19611 vdd.n2398 vdd.n760 72.8958
R19612 vdd.n2398 vdd.n759 72.8958
R19613 vdd.n2398 vdd.n758 72.8958
R19614 vdd.n2398 vdd.n757 72.8958
R19615 vdd.n2398 vdd.n756 72.8958
R19616 vdd.n2398 vdd.n755 72.8958
R19617 vdd.n2398 vdd.n754 72.8958
R19618 vdd.n2398 vdd.n753 72.8958
R19619 vdd.n2120 vdd.n948 72.8958
R19620 vdd.n2120 vdd.n949 72.8958
R19621 vdd.n2120 vdd.n950 72.8958
R19622 vdd.n2120 vdd.n951 72.8958
R19623 vdd.n2120 vdd.n952 72.8958
R19624 vdd.n2120 vdd.n953 72.8958
R19625 vdd.n2120 vdd.n954 72.8958
R19626 vdd.n2120 vdd.n955 72.8958
R19627 vdd.n2120 vdd.n956 72.8958
R19628 vdd.n2120 vdd.n957 72.8958
R19629 vdd.n2120 vdd.n958 72.8958
R19630 vdd.n2120 vdd.n959 72.8958
R19631 vdd.n2120 vdd.n960 72.8958
R19632 vdd.n2120 vdd.n961 72.8958
R19633 vdd.n2120 vdd.n962 72.8958
R19634 vdd.n2120 vdd.n963 72.8958
R19635 vdd.n2120 vdd.n964 72.8958
R19636 vdd.n1877 vdd.n1876 66.2847
R19637 vdd.n1876 vdd.n1652 66.2847
R19638 vdd.n1876 vdd.n1653 66.2847
R19639 vdd.n1876 vdd.n1654 66.2847
R19640 vdd.n1876 vdd.n1655 66.2847
R19641 vdd.n1876 vdd.n1656 66.2847
R19642 vdd.n1876 vdd.n1657 66.2847
R19643 vdd.n1876 vdd.n1658 66.2847
R19644 vdd.n1876 vdd.n1659 66.2847
R19645 vdd.n1876 vdd.n1660 66.2847
R19646 vdd.n1876 vdd.n1661 66.2847
R19647 vdd.n1876 vdd.n1662 66.2847
R19648 vdd.n1876 vdd.n1663 66.2847
R19649 vdd.n1876 vdd.n1664 66.2847
R19650 vdd.n1876 vdd.n1665 66.2847
R19651 vdd.n1876 vdd.n1666 66.2847
R19652 vdd.n1876 vdd.n1667 66.2847
R19653 vdd.n1876 vdd.n1668 66.2847
R19654 vdd.n1876 vdd.n1669 66.2847
R19655 vdd.n1876 vdd.n1670 66.2847
R19656 vdd.n1876 vdd.n1671 66.2847
R19657 vdd.n1876 vdd.n1672 66.2847
R19658 vdd.n1876 vdd.n1673 66.2847
R19659 vdd.n1876 vdd.n1674 66.2847
R19660 vdd.n1876 vdd.n1675 66.2847
R19661 vdd.n1876 vdd.n1676 66.2847
R19662 vdd.n1876 vdd.n1677 66.2847
R19663 vdd.n1876 vdd.n1678 66.2847
R19664 vdd.n1876 vdd.n1679 66.2847
R19665 vdd.n1876 vdd.n1680 66.2847
R19666 vdd.n1876 vdd.n1681 66.2847
R19667 vdd.n1316 vdd.n931 66.2847
R19668 vdd.n1313 vdd.n931 66.2847
R19669 vdd.n1309 vdd.n931 66.2847
R19670 vdd.n1986 vdd.n931 66.2847
R19671 vdd.n1065 vdd.n931 66.2847
R19672 vdd.n1993 vdd.n931 66.2847
R19673 vdd.n1058 vdd.n931 66.2847
R19674 vdd.n2000 vdd.n931 66.2847
R19675 vdd.n1051 vdd.n931 66.2847
R19676 vdd.n2007 vdd.n931 66.2847
R19677 vdd.n1045 vdd.n931 66.2847
R19678 vdd.n1040 vdd.n931 66.2847
R19679 vdd.n2018 vdd.n931 66.2847
R19680 vdd.n1032 vdd.n931 66.2847
R19681 vdd.n2025 vdd.n931 66.2847
R19682 vdd.n1025 vdd.n931 66.2847
R19683 vdd.n2032 vdd.n931 66.2847
R19684 vdd.n1018 vdd.n931 66.2847
R19685 vdd.n2039 vdd.n931 66.2847
R19686 vdd.n1011 vdd.n931 66.2847
R19687 vdd.n2046 vdd.n931 66.2847
R19688 vdd.n1005 vdd.n931 66.2847
R19689 vdd.n1000 vdd.n931 66.2847
R19690 vdd.n2057 vdd.n931 66.2847
R19691 vdd.n992 vdd.n931 66.2847
R19692 vdd.n2064 vdd.n931 66.2847
R19693 vdd.n985 vdd.n931 66.2847
R19694 vdd.n2071 vdd.n931 66.2847
R19695 vdd.n978 vdd.n931 66.2847
R19696 vdd.n2078 vdd.n931 66.2847
R19697 vdd.n2083 vdd.n931 66.2847
R19698 vdd.n974 vdd.n931 66.2847
R19699 vdd.n3113 vdd.n3112 66.2847
R19700 vdd.n3112 vdd.n485 66.2847
R19701 vdd.n3112 vdd.n486 66.2847
R19702 vdd.n3112 vdd.n487 66.2847
R19703 vdd.n3112 vdd.n488 66.2847
R19704 vdd.n3112 vdd.n489 66.2847
R19705 vdd.n3112 vdd.n490 66.2847
R19706 vdd.n3112 vdd.n491 66.2847
R19707 vdd.n3112 vdd.n492 66.2847
R19708 vdd.n3112 vdd.n493 66.2847
R19709 vdd.n3112 vdd.n494 66.2847
R19710 vdd.n3112 vdd.n495 66.2847
R19711 vdd.n3112 vdd.n496 66.2847
R19712 vdd.n3112 vdd.n497 66.2847
R19713 vdd.n3112 vdd.n498 66.2847
R19714 vdd.n3112 vdd.n499 66.2847
R19715 vdd.n3112 vdd.n500 66.2847
R19716 vdd.n3112 vdd.n501 66.2847
R19717 vdd.n3112 vdd.n502 66.2847
R19718 vdd.n3112 vdd.n503 66.2847
R19719 vdd.n3112 vdd.n504 66.2847
R19720 vdd.n3112 vdd.n505 66.2847
R19721 vdd.n3112 vdd.n506 66.2847
R19722 vdd.n3112 vdd.n507 66.2847
R19723 vdd.n3112 vdd.n508 66.2847
R19724 vdd.n3112 vdd.n509 66.2847
R19725 vdd.n3112 vdd.n510 66.2847
R19726 vdd.n3112 vdd.n511 66.2847
R19727 vdd.n3112 vdd.n512 66.2847
R19728 vdd.n3112 vdd.n513 66.2847
R19729 vdd.n3112 vdd.n514 66.2847
R19730 vdd.n3177 vdd.n329 66.2847
R19731 vdd.n3186 vdd.n329 66.2847
R19732 vdd.n439 vdd.n329 66.2847
R19733 vdd.n3193 vdd.n329 66.2847
R19734 vdd.n432 vdd.n329 66.2847
R19735 vdd.n3200 vdd.n329 66.2847
R19736 vdd.n425 vdd.n329 66.2847
R19737 vdd.n3207 vdd.n329 66.2847
R19738 vdd.n418 vdd.n329 66.2847
R19739 vdd.n3214 vdd.n329 66.2847
R19740 vdd.n412 vdd.n329 66.2847
R19741 vdd.n407 vdd.n329 66.2847
R19742 vdd.n3225 vdd.n329 66.2847
R19743 vdd.n399 vdd.n329 66.2847
R19744 vdd.n3232 vdd.n329 66.2847
R19745 vdd.n392 vdd.n329 66.2847
R19746 vdd.n3239 vdd.n329 66.2847
R19747 vdd.n385 vdd.n329 66.2847
R19748 vdd.n3246 vdd.n329 66.2847
R19749 vdd.n378 vdd.n329 66.2847
R19750 vdd.n3253 vdd.n329 66.2847
R19751 vdd.n372 vdd.n329 66.2847
R19752 vdd.n367 vdd.n329 66.2847
R19753 vdd.n3264 vdd.n329 66.2847
R19754 vdd.n359 vdd.n329 66.2847
R19755 vdd.n3271 vdd.n329 66.2847
R19756 vdd.n352 vdd.n329 66.2847
R19757 vdd.n3278 vdd.n329 66.2847
R19758 vdd.n345 vdd.n329 66.2847
R19759 vdd.n3285 vdd.n329 66.2847
R19760 vdd.n3288 vdd.n329 66.2847
R19761 vdd.n333 vdd.n329 66.2847
R19762 vdd.n334 vdd.n333 52.4337
R19763 vdd.n3288 vdd.n3287 52.4337
R19764 vdd.n3285 vdd.n3284 52.4337
R19765 vdd.n3280 vdd.n345 52.4337
R19766 vdd.n3278 vdd.n3277 52.4337
R19767 vdd.n3273 vdd.n352 52.4337
R19768 vdd.n3271 vdd.n3270 52.4337
R19769 vdd.n3266 vdd.n359 52.4337
R19770 vdd.n3264 vdd.n3263 52.4337
R19771 vdd.n368 vdd.n367 52.4337
R19772 vdd.n3255 vdd.n372 52.4337
R19773 vdd.n3253 vdd.n3252 52.4337
R19774 vdd.n3248 vdd.n378 52.4337
R19775 vdd.n3246 vdd.n3245 52.4337
R19776 vdd.n3241 vdd.n385 52.4337
R19777 vdd.n3239 vdd.n3238 52.4337
R19778 vdd.n3234 vdd.n392 52.4337
R19779 vdd.n3232 vdd.n3231 52.4337
R19780 vdd.n3227 vdd.n399 52.4337
R19781 vdd.n3225 vdd.n3224 52.4337
R19782 vdd.n408 vdd.n407 52.4337
R19783 vdd.n3216 vdd.n412 52.4337
R19784 vdd.n3214 vdd.n3213 52.4337
R19785 vdd.n3209 vdd.n418 52.4337
R19786 vdd.n3207 vdd.n3206 52.4337
R19787 vdd.n3202 vdd.n425 52.4337
R19788 vdd.n3200 vdd.n3199 52.4337
R19789 vdd.n3195 vdd.n432 52.4337
R19790 vdd.n3193 vdd.n3192 52.4337
R19791 vdd.n3188 vdd.n439 52.4337
R19792 vdd.n3186 vdd.n3185 52.4337
R19793 vdd.n3178 vdd.n3177 52.4337
R19794 vdd.n3114 vdd.n3113 52.4337
R19795 vdd.n517 vdd.n485 52.4337
R19796 vdd.n523 vdd.n486 52.4337
R19797 vdd.n3103 vdd.n487 52.4337
R19798 vdd.n3099 vdd.n488 52.4337
R19799 vdd.n3095 vdd.n489 52.4337
R19800 vdd.n3091 vdd.n490 52.4337
R19801 vdd.n3087 vdd.n491 52.4337
R19802 vdd.n3083 vdd.n492 52.4337
R19803 vdd.n3079 vdd.n493 52.4337
R19804 vdd.n3071 vdd.n494 52.4337
R19805 vdd.n3067 vdd.n495 52.4337
R19806 vdd.n3063 vdd.n496 52.4337
R19807 vdd.n3059 vdd.n497 52.4337
R19808 vdd.n3055 vdd.n498 52.4337
R19809 vdd.n3051 vdd.n499 52.4337
R19810 vdd.n3047 vdd.n500 52.4337
R19811 vdd.n3043 vdd.n501 52.4337
R19812 vdd.n3039 vdd.n502 52.4337
R19813 vdd.n3035 vdd.n503 52.4337
R19814 vdd.n3031 vdd.n504 52.4337
R19815 vdd.n3025 vdd.n505 52.4337
R19816 vdd.n3021 vdd.n506 52.4337
R19817 vdd.n3017 vdd.n507 52.4337
R19818 vdd.n3013 vdd.n508 52.4337
R19819 vdd.n3009 vdd.n509 52.4337
R19820 vdd.n3005 vdd.n510 52.4337
R19821 vdd.n3001 vdd.n511 52.4337
R19822 vdd.n2997 vdd.n512 52.4337
R19823 vdd.n2993 vdd.n513 52.4337
R19824 vdd.n2989 vdd.n514 52.4337
R19825 vdd.n2085 vdd.n974 52.4337
R19826 vdd.n2083 vdd.n2082 52.4337
R19827 vdd.n2078 vdd.n2077 52.4337
R19828 vdd.n2073 vdd.n978 52.4337
R19829 vdd.n2071 vdd.n2070 52.4337
R19830 vdd.n2066 vdd.n985 52.4337
R19831 vdd.n2064 vdd.n2063 52.4337
R19832 vdd.n2059 vdd.n992 52.4337
R19833 vdd.n2057 vdd.n2056 52.4337
R19834 vdd.n1001 vdd.n1000 52.4337
R19835 vdd.n2048 vdd.n1005 52.4337
R19836 vdd.n2046 vdd.n2045 52.4337
R19837 vdd.n2041 vdd.n1011 52.4337
R19838 vdd.n2039 vdd.n2038 52.4337
R19839 vdd.n2034 vdd.n1018 52.4337
R19840 vdd.n2032 vdd.n2031 52.4337
R19841 vdd.n2027 vdd.n1025 52.4337
R19842 vdd.n2025 vdd.n2024 52.4337
R19843 vdd.n2020 vdd.n1032 52.4337
R19844 vdd.n2018 vdd.n2017 52.4337
R19845 vdd.n1041 vdd.n1040 52.4337
R19846 vdd.n2009 vdd.n1045 52.4337
R19847 vdd.n2007 vdd.n2006 52.4337
R19848 vdd.n2002 vdd.n1051 52.4337
R19849 vdd.n2000 vdd.n1999 52.4337
R19850 vdd.n1995 vdd.n1058 52.4337
R19851 vdd.n1993 vdd.n1992 52.4337
R19852 vdd.n1988 vdd.n1065 52.4337
R19853 vdd.n1986 vdd.n1985 52.4337
R19854 vdd.n1310 vdd.n1309 52.4337
R19855 vdd.n1314 vdd.n1313 52.4337
R19856 vdd.n1974 vdd.n1316 52.4337
R19857 vdd.n1878 vdd.n1877 52.4337
R19858 vdd.n1684 vdd.n1652 52.4337
R19859 vdd.n1688 vdd.n1653 52.4337
R19860 vdd.n1690 vdd.n1654 52.4337
R19861 vdd.n1694 vdd.n1655 52.4337
R19862 vdd.n1696 vdd.n1656 52.4337
R19863 vdd.n1700 vdd.n1657 52.4337
R19864 vdd.n1702 vdd.n1658 52.4337
R19865 vdd.n1706 vdd.n1659 52.4337
R19866 vdd.n1708 vdd.n1660 52.4337
R19867 vdd.n1714 vdd.n1661 52.4337
R19868 vdd.n1716 vdd.n1662 52.4337
R19869 vdd.n1720 vdd.n1663 52.4337
R19870 vdd.n1722 vdd.n1664 52.4337
R19871 vdd.n1726 vdd.n1665 52.4337
R19872 vdd.n1728 vdd.n1666 52.4337
R19873 vdd.n1732 vdd.n1667 52.4337
R19874 vdd.n1734 vdd.n1668 52.4337
R19875 vdd.n1738 vdd.n1669 52.4337
R19876 vdd.n1740 vdd.n1670 52.4337
R19877 vdd.n1812 vdd.n1671 52.4337
R19878 vdd.n1745 vdd.n1672 52.4337
R19879 vdd.n1749 vdd.n1673 52.4337
R19880 vdd.n1751 vdd.n1674 52.4337
R19881 vdd.n1755 vdd.n1675 52.4337
R19882 vdd.n1757 vdd.n1676 52.4337
R19883 vdd.n1761 vdd.n1677 52.4337
R19884 vdd.n1763 vdd.n1678 52.4337
R19885 vdd.n1767 vdd.n1679 52.4337
R19886 vdd.n1769 vdd.n1680 52.4337
R19887 vdd.n1773 vdd.n1681 52.4337
R19888 vdd.n1877 vdd.n1651 52.4337
R19889 vdd.n1687 vdd.n1652 52.4337
R19890 vdd.n1689 vdd.n1653 52.4337
R19891 vdd.n1693 vdd.n1654 52.4337
R19892 vdd.n1695 vdd.n1655 52.4337
R19893 vdd.n1699 vdd.n1656 52.4337
R19894 vdd.n1701 vdd.n1657 52.4337
R19895 vdd.n1705 vdd.n1658 52.4337
R19896 vdd.n1707 vdd.n1659 52.4337
R19897 vdd.n1713 vdd.n1660 52.4337
R19898 vdd.n1715 vdd.n1661 52.4337
R19899 vdd.n1719 vdd.n1662 52.4337
R19900 vdd.n1721 vdd.n1663 52.4337
R19901 vdd.n1725 vdd.n1664 52.4337
R19902 vdd.n1727 vdd.n1665 52.4337
R19903 vdd.n1731 vdd.n1666 52.4337
R19904 vdd.n1733 vdd.n1667 52.4337
R19905 vdd.n1737 vdd.n1668 52.4337
R19906 vdd.n1739 vdd.n1669 52.4337
R19907 vdd.n1743 vdd.n1670 52.4337
R19908 vdd.n1744 vdd.n1671 52.4337
R19909 vdd.n1748 vdd.n1672 52.4337
R19910 vdd.n1750 vdd.n1673 52.4337
R19911 vdd.n1754 vdd.n1674 52.4337
R19912 vdd.n1756 vdd.n1675 52.4337
R19913 vdd.n1760 vdd.n1676 52.4337
R19914 vdd.n1762 vdd.n1677 52.4337
R19915 vdd.n1766 vdd.n1678 52.4337
R19916 vdd.n1768 vdd.n1679 52.4337
R19917 vdd.n1772 vdd.n1680 52.4337
R19918 vdd.n1774 vdd.n1681 52.4337
R19919 vdd.n1316 vdd.n1315 52.4337
R19920 vdd.n1313 vdd.n1312 52.4337
R19921 vdd.n1309 vdd.n1066 52.4337
R19922 vdd.n1987 vdd.n1986 52.4337
R19923 vdd.n1065 vdd.n1059 52.4337
R19924 vdd.n1994 vdd.n1993 52.4337
R19925 vdd.n1058 vdd.n1052 52.4337
R19926 vdd.n2001 vdd.n2000 52.4337
R19927 vdd.n1051 vdd.n1046 52.4337
R19928 vdd.n2008 vdd.n2007 52.4337
R19929 vdd.n1045 vdd.n1044 52.4337
R19930 vdd.n1040 vdd.n1033 52.4337
R19931 vdd.n2019 vdd.n2018 52.4337
R19932 vdd.n1032 vdd.n1026 52.4337
R19933 vdd.n2026 vdd.n2025 52.4337
R19934 vdd.n1025 vdd.n1019 52.4337
R19935 vdd.n2033 vdd.n2032 52.4337
R19936 vdd.n1018 vdd.n1012 52.4337
R19937 vdd.n2040 vdd.n2039 52.4337
R19938 vdd.n1011 vdd.n1006 52.4337
R19939 vdd.n2047 vdd.n2046 52.4337
R19940 vdd.n1005 vdd.n1004 52.4337
R19941 vdd.n1000 vdd.n993 52.4337
R19942 vdd.n2058 vdd.n2057 52.4337
R19943 vdd.n992 vdd.n986 52.4337
R19944 vdd.n2065 vdd.n2064 52.4337
R19945 vdd.n985 vdd.n979 52.4337
R19946 vdd.n2072 vdd.n2071 52.4337
R19947 vdd.n978 vdd.n975 52.4337
R19948 vdd.n2079 vdd.n2078 52.4337
R19949 vdd.n2084 vdd.n2083 52.4337
R19950 vdd.n1320 vdd.n974 52.4337
R19951 vdd.n3113 vdd.n483 52.4337
R19952 vdd.n522 vdd.n485 52.4337
R19953 vdd.n3104 vdd.n486 52.4337
R19954 vdd.n3100 vdd.n487 52.4337
R19955 vdd.n3096 vdd.n488 52.4337
R19956 vdd.n3092 vdd.n489 52.4337
R19957 vdd.n3088 vdd.n490 52.4337
R19958 vdd.n3084 vdd.n491 52.4337
R19959 vdd.n3080 vdd.n492 52.4337
R19960 vdd.n3070 vdd.n493 52.4337
R19961 vdd.n3068 vdd.n494 52.4337
R19962 vdd.n3064 vdd.n495 52.4337
R19963 vdd.n3060 vdd.n496 52.4337
R19964 vdd.n3056 vdd.n497 52.4337
R19965 vdd.n3052 vdd.n498 52.4337
R19966 vdd.n3048 vdd.n499 52.4337
R19967 vdd.n3044 vdd.n500 52.4337
R19968 vdd.n3040 vdd.n501 52.4337
R19969 vdd.n3036 vdd.n502 52.4337
R19970 vdd.n3032 vdd.n503 52.4337
R19971 vdd.n3024 vdd.n504 52.4337
R19972 vdd.n3022 vdd.n505 52.4337
R19973 vdd.n3018 vdd.n506 52.4337
R19974 vdd.n3014 vdd.n507 52.4337
R19975 vdd.n3010 vdd.n508 52.4337
R19976 vdd.n3006 vdd.n509 52.4337
R19977 vdd.n3002 vdd.n510 52.4337
R19978 vdd.n2998 vdd.n511 52.4337
R19979 vdd.n2994 vdd.n512 52.4337
R19980 vdd.n2990 vdd.n513 52.4337
R19981 vdd.n2986 vdd.n514 52.4337
R19982 vdd.n3177 vdd.n440 52.4337
R19983 vdd.n3187 vdd.n3186 52.4337
R19984 vdd.n439 vdd.n433 52.4337
R19985 vdd.n3194 vdd.n3193 52.4337
R19986 vdd.n432 vdd.n426 52.4337
R19987 vdd.n3201 vdd.n3200 52.4337
R19988 vdd.n425 vdd.n419 52.4337
R19989 vdd.n3208 vdd.n3207 52.4337
R19990 vdd.n418 vdd.n413 52.4337
R19991 vdd.n3215 vdd.n3214 52.4337
R19992 vdd.n412 vdd.n411 52.4337
R19993 vdd.n407 vdd.n400 52.4337
R19994 vdd.n3226 vdd.n3225 52.4337
R19995 vdd.n399 vdd.n393 52.4337
R19996 vdd.n3233 vdd.n3232 52.4337
R19997 vdd.n392 vdd.n386 52.4337
R19998 vdd.n3240 vdd.n3239 52.4337
R19999 vdd.n385 vdd.n379 52.4337
R20000 vdd.n3247 vdd.n3246 52.4337
R20001 vdd.n378 vdd.n373 52.4337
R20002 vdd.n3254 vdd.n3253 52.4337
R20003 vdd.n372 vdd.n371 52.4337
R20004 vdd.n367 vdd.n360 52.4337
R20005 vdd.n3265 vdd.n3264 52.4337
R20006 vdd.n359 vdd.n353 52.4337
R20007 vdd.n3272 vdd.n3271 52.4337
R20008 vdd.n352 vdd.n346 52.4337
R20009 vdd.n3279 vdd.n3278 52.4337
R20010 vdd.n345 vdd.n338 52.4337
R20011 vdd.n3286 vdd.n3285 52.4337
R20012 vdd.n3289 vdd.n3288 52.4337
R20013 vdd.n333 vdd.n330 52.4337
R20014 vdd.t166 vdd.t184 51.4683
R20015 vdd.n250 vdd.n248 42.0461
R20016 vdd.n160 vdd.n158 42.0461
R20017 vdd.n71 vdd.n69 42.0461
R20018 vdd.n1567 vdd.n1565 42.0461
R20019 vdd.n1477 vdd.n1475 42.0461
R20020 vdd.n1388 vdd.n1386 42.0461
R20021 vdd.n296 vdd.n295 41.6884
R20022 vdd.n206 vdd.n205 41.6884
R20023 vdd.n117 vdd.n116 41.6884
R20024 vdd.n1613 vdd.n1612 41.6884
R20025 vdd.n1523 vdd.n1522 41.6884
R20026 vdd.n1434 vdd.n1433 41.6884
R20027 vdd.n1777 vdd.n1776 41.1157
R20028 vdd.n1815 vdd.n1814 41.1157
R20029 vdd.n1711 vdd.n1710 41.1157
R20030 vdd.n3182 vdd.n3181 41.1157
R20031 vdd.n3221 vdd.n406 41.1157
R20032 vdd.n3260 vdd.n366 41.1157
R20033 vdd.n2939 vdd.n2938 39.2114
R20034 vdd.n2936 vdd.n2935 39.2114
R20035 vdd.n2931 vdd.n605 39.2114
R20036 vdd.n2929 vdd.n2928 39.2114
R20037 vdd.n2924 vdd.n608 39.2114
R20038 vdd.n2922 vdd.n2921 39.2114
R20039 vdd.n2917 vdd.n611 39.2114
R20040 vdd.n2915 vdd.n2914 39.2114
R20041 vdd.n2911 vdd.n2910 39.2114
R20042 vdd.n2906 vdd.n614 39.2114
R20043 vdd.n2904 vdd.n2903 39.2114
R20044 vdd.n2899 vdd.n617 39.2114
R20045 vdd.n2897 vdd.n2896 39.2114
R20046 vdd.n2892 vdd.n620 39.2114
R20047 vdd.n2890 vdd.n2889 39.2114
R20048 vdd.n2884 vdd.n625 39.2114
R20049 vdd.n2882 vdd.n2881 39.2114
R20050 vdd.n2704 vdd.n2703 39.2114
R20051 vdd.n2433 vdd.n2399 39.2114
R20052 vdd.n2696 vdd.n2400 39.2114
R20053 vdd.n2692 vdd.n2401 39.2114
R20054 vdd.n2688 vdd.n2402 39.2114
R20055 vdd.n2684 vdd.n2403 39.2114
R20056 vdd.n2680 vdd.n2404 39.2114
R20057 vdd.n2676 vdd.n2405 39.2114
R20058 vdd.n2672 vdd.n2406 39.2114
R20059 vdd.n2668 vdd.n2407 39.2114
R20060 vdd.n2664 vdd.n2408 39.2114
R20061 vdd.n2660 vdd.n2409 39.2114
R20062 vdd.n2656 vdd.n2410 39.2114
R20063 vdd.n2652 vdd.n2411 39.2114
R20064 vdd.n2648 vdd.n2412 39.2114
R20065 vdd.n2644 vdd.n2413 39.2114
R20066 vdd.n2639 vdd.n2414 39.2114
R20067 vdd.n2393 vdd.n787 39.2114
R20068 vdd.n2389 vdd.n786 39.2114
R20069 vdd.n2385 vdd.n785 39.2114
R20070 vdd.n2381 vdd.n784 39.2114
R20071 vdd.n2377 vdd.n783 39.2114
R20072 vdd.n2373 vdd.n782 39.2114
R20073 vdd.n2369 vdd.n781 39.2114
R20074 vdd.n2365 vdd.n780 39.2114
R20075 vdd.n2361 vdd.n779 39.2114
R20076 vdd.n2357 vdd.n778 39.2114
R20077 vdd.n2353 vdd.n777 39.2114
R20078 vdd.n2349 vdd.n776 39.2114
R20079 vdd.n2345 vdd.n775 39.2114
R20080 vdd.n2341 vdd.n774 39.2114
R20081 vdd.n2337 vdd.n773 39.2114
R20082 vdd.n2332 vdd.n772 39.2114
R20083 vdd.n2328 vdd.n771 39.2114
R20084 vdd.n2122 vdd.n2121 39.2114
R20085 vdd.n966 vdd.n932 39.2114
R20086 vdd.n2114 vdd.n933 39.2114
R20087 vdd.n2110 vdd.n934 39.2114
R20088 vdd.n2106 vdd.n935 39.2114
R20089 vdd.n2102 vdd.n936 39.2114
R20090 vdd.n2098 vdd.n937 39.2114
R20091 vdd.n2094 vdd.n938 39.2114
R20092 vdd.n2090 vdd.n939 39.2114
R20093 vdd.n1112 vdd.n940 39.2114
R20094 vdd.n1116 vdd.n941 39.2114
R20095 vdd.n1120 vdd.n942 39.2114
R20096 vdd.n1124 vdd.n943 39.2114
R20097 vdd.n1128 vdd.n944 39.2114
R20098 vdd.n1132 vdd.n945 39.2114
R20099 vdd.n1136 vdd.n946 39.2114
R20100 vdd.n1141 vdd.n947 39.2114
R20101 vdd.n2858 vdd.n2857 39.2114
R20102 vdd.n2853 vdd.n2825 39.2114
R20103 vdd.n2851 vdd.n2850 39.2114
R20104 vdd.n2846 vdd.n2828 39.2114
R20105 vdd.n2844 vdd.n2843 39.2114
R20106 vdd.n2839 vdd.n2831 39.2114
R20107 vdd.n2837 vdd.n2836 39.2114
R20108 vdd.n2832 vdd.n577 39.2114
R20109 vdd.n2976 vdd.n2975 39.2114
R20110 vdd.n2973 vdd.n2972 39.2114
R20111 vdd.n2968 vdd.n581 39.2114
R20112 vdd.n2966 vdd.n2965 39.2114
R20113 vdd.n2961 vdd.n584 39.2114
R20114 vdd.n2959 vdd.n2958 39.2114
R20115 vdd.n2954 vdd.n587 39.2114
R20116 vdd.n2952 vdd.n2951 39.2114
R20117 vdd.n2947 vdd.n593 39.2114
R20118 vdd.n2440 vdd.n2415 39.2114
R20119 vdd.n2444 vdd.n2416 39.2114
R20120 vdd.n2448 vdd.n2417 39.2114
R20121 vdd.n2452 vdd.n2418 39.2114
R20122 vdd.n2456 vdd.n2419 39.2114
R20123 vdd.n2460 vdd.n2420 39.2114
R20124 vdd.n2464 vdd.n2421 39.2114
R20125 vdd.n2468 vdd.n2422 39.2114
R20126 vdd.n2472 vdd.n2423 39.2114
R20127 vdd.n2476 vdd.n2424 39.2114
R20128 vdd.n2480 vdd.n2425 39.2114
R20129 vdd.n2484 vdd.n2426 39.2114
R20130 vdd.n2488 vdd.n2427 39.2114
R20131 vdd.n2492 vdd.n2428 39.2114
R20132 vdd.n2496 vdd.n2429 39.2114
R20133 vdd.n2500 vdd.n2430 39.2114
R20134 vdd.n2504 vdd.n2431 39.2114
R20135 vdd.n2443 vdd.n2415 39.2114
R20136 vdd.n2447 vdd.n2416 39.2114
R20137 vdd.n2451 vdd.n2417 39.2114
R20138 vdd.n2455 vdd.n2418 39.2114
R20139 vdd.n2459 vdd.n2419 39.2114
R20140 vdd.n2463 vdd.n2420 39.2114
R20141 vdd.n2467 vdd.n2421 39.2114
R20142 vdd.n2471 vdd.n2422 39.2114
R20143 vdd.n2475 vdd.n2423 39.2114
R20144 vdd.n2479 vdd.n2424 39.2114
R20145 vdd.n2483 vdd.n2425 39.2114
R20146 vdd.n2487 vdd.n2426 39.2114
R20147 vdd.n2491 vdd.n2427 39.2114
R20148 vdd.n2495 vdd.n2428 39.2114
R20149 vdd.n2499 vdd.n2429 39.2114
R20150 vdd.n2503 vdd.n2430 39.2114
R20151 vdd.n2506 vdd.n2431 39.2114
R20152 vdd.n593 vdd.n588 39.2114
R20153 vdd.n2953 vdd.n2952 39.2114
R20154 vdd.n587 vdd.n585 39.2114
R20155 vdd.n2960 vdd.n2959 39.2114
R20156 vdd.n584 vdd.n582 39.2114
R20157 vdd.n2967 vdd.n2966 39.2114
R20158 vdd.n581 vdd.n579 39.2114
R20159 vdd.n2974 vdd.n2973 39.2114
R20160 vdd.n2977 vdd.n2976 39.2114
R20161 vdd.n2833 vdd.n2832 39.2114
R20162 vdd.n2838 vdd.n2837 39.2114
R20163 vdd.n2831 vdd.n2829 39.2114
R20164 vdd.n2845 vdd.n2844 39.2114
R20165 vdd.n2828 vdd.n2826 39.2114
R20166 vdd.n2852 vdd.n2851 39.2114
R20167 vdd.n2825 vdd.n2823 39.2114
R20168 vdd.n2859 vdd.n2858 39.2114
R20169 vdd.n2121 vdd.n930 39.2114
R20170 vdd.n2115 vdd.n932 39.2114
R20171 vdd.n2111 vdd.n933 39.2114
R20172 vdd.n2107 vdd.n934 39.2114
R20173 vdd.n2103 vdd.n935 39.2114
R20174 vdd.n2099 vdd.n936 39.2114
R20175 vdd.n2095 vdd.n937 39.2114
R20176 vdd.n2091 vdd.n938 39.2114
R20177 vdd.n1111 vdd.n939 39.2114
R20178 vdd.n1115 vdd.n940 39.2114
R20179 vdd.n1119 vdd.n941 39.2114
R20180 vdd.n1123 vdd.n942 39.2114
R20181 vdd.n1127 vdd.n943 39.2114
R20182 vdd.n1131 vdd.n944 39.2114
R20183 vdd.n1135 vdd.n945 39.2114
R20184 vdd.n1140 vdd.n946 39.2114
R20185 vdd.n1144 vdd.n947 39.2114
R20186 vdd.n2331 vdd.n771 39.2114
R20187 vdd.n2336 vdd.n772 39.2114
R20188 vdd.n2340 vdd.n773 39.2114
R20189 vdd.n2344 vdd.n774 39.2114
R20190 vdd.n2348 vdd.n775 39.2114
R20191 vdd.n2352 vdd.n776 39.2114
R20192 vdd.n2356 vdd.n777 39.2114
R20193 vdd.n2360 vdd.n778 39.2114
R20194 vdd.n2364 vdd.n779 39.2114
R20195 vdd.n2368 vdd.n780 39.2114
R20196 vdd.n2372 vdd.n781 39.2114
R20197 vdd.n2376 vdd.n782 39.2114
R20198 vdd.n2380 vdd.n783 39.2114
R20199 vdd.n2384 vdd.n784 39.2114
R20200 vdd.n2388 vdd.n785 39.2114
R20201 vdd.n2392 vdd.n786 39.2114
R20202 vdd.n789 vdd.n787 39.2114
R20203 vdd.n2703 vdd.n752 39.2114
R20204 vdd.n2697 vdd.n2399 39.2114
R20205 vdd.n2693 vdd.n2400 39.2114
R20206 vdd.n2689 vdd.n2401 39.2114
R20207 vdd.n2685 vdd.n2402 39.2114
R20208 vdd.n2681 vdd.n2403 39.2114
R20209 vdd.n2677 vdd.n2404 39.2114
R20210 vdd.n2673 vdd.n2405 39.2114
R20211 vdd.n2669 vdd.n2406 39.2114
R20212 vdd.n2665 vdd.n2407 39.2114
R20213 vdd.n2661 vdd.n2408 39.2114
R20214 vdd.n2657 vdd.n2409 39.2114
R20215 vdd.n2653 vdd.n2410 39.2114
R20216 vdd.n2649 vdd.n2411 39.2114
R20217 vdd.n2645 vdd.n2412 39.2114
R20218 vdd.n2640 vdd.n2413 39.2114
R20219 vdd.n2636 vdd.n2414 39.2114
R20220 vdd.n2883 vdd.n2882 39.2114
R20221 vdd.n625 vdd.n621 39.2114
R20222 vdd.n2891 vdd.n2890 39.2114
R20223 vdd.n620 vdd.n618 39.2114
R20224 vdd.n2898 vdd.n2897 39.2114
R20225 vdd.n617 vdd.n615 39.2114
R20226 vdd.n2905 vdd.n2904 39.2114
R20227 vdd.n614 vdd.n612 39.2114
R20228 vdd.n2912 vdd.n2911 39.2114
R20229 vdd.n2916 vdd.n2915 39.2114
R20230 vdd.n611 vdd.n609 39.2114
R20231 vdd.n2923 vdd.n2922 39.2114
R20232 vdd.n608 vdd.n606 39.2114
R20233 vdd.n2930 vdd.n2929 39.2114
R20234 vdd.n605 vdd.n603 39.2114
R20235 vdd.n2937 vdd.n2936 39.2114
R20236 vdd.n2940 vdd.n2939 39.2114
R20237 vdd.n798 vdd.n753 39.2114
R20238 vdd.n2320 vdd.n754 39.2114
R20239 vdd.n2316 vdd.n755 39.2114
R20240 vdd.n2312 vdd.n756 39.2114
R20241 vdd.n2308 vdd.n757 39.2114
R20242 vdd.n2304 vdd.n758 39.2114
R20243 vdd.n2300 vdd.n759 39.2114
R20244 vdd.n2296 vdd.n760 39.2114
R20245 vdd.n2292 vdd.n761 39.2114
R20246 vdd.n2288 vdd.n762 39.2114
R20247 vdd.n2284 vdd.n763 39.2114
R20248 vdd.n2280 vdd.n764 39.2114
R20249 vdd.n2276 vdd.n765 39.2114
R20250 vdd.n2272 vdd.n766 39.2114
R20251 vdd.n2268 vdd.n767 39.2114
R20252 vdd.n2264 vdd.n768 39.2114
R20253 vdd.n2260 vdd.n769 39.2114
R20254 vdd.n1070 vdd.n948 39.2114
R20255 vdd.n1074 vdd.n949 39.2114
R20256 vdd.n1078 vdd.n950 39.2114
R20257 vdd.n1082 vdd.n951 39.2114
R20258 vdd.n1086 vdd.n952 39.2114
R20259 vdd.n1090 vdd.n953 39.2114
R20260 vdd.n1094 vdd.n954 39.2114
R20261 vdd.n1098 vdd.n955 39.2114
R20262 vdd.n1102 vdd.n956 39.2114
R20263 vdd.n1303 vdd.n957 39.2114
R20264 vdd.n1300 vdd.n958 39.2114
R20265 vdd.n1296 vdd.n959 39.2114
R20266 vdd.n1292 vdd.n960 39.2114
R20267 vdd.n1288 vdd.n961 39.2114
R20268 vdd.n1284 vdd.n962 39.2114
R20269 vdd.n1280 vdd.n963 39.2114
R20270 vdd.n1276 vdd.n964 39.2114
R20271 vdd.n2257 vdd.n769 39.2114
R20272 vdd.n2261 vdd.n768 39.2114
R20273 vdd.n2265 vdd.n767 39.2114
R20274 vdd.n2269 vdd.n766 39.2114
R20275 vdd.n2273 vdd.n765 39.2114
R20276 vdd.n2277 vdd.n764 39.2114
R20277 vdd.n2281 vdd.n763 39.2114
R20278 vdd.n2285 vdd.n762 39.2114
R20279 vdd.n2289 vdd.n761 39.2114
R20280 vdd.n2293 vdd.n760 39.2114
R20281 vdd.n2297 vdd.n759 39.2114
R20282 vdd.n2301 vdd.n758 39.2114
R20283 vdd.n2305 vdd.n757 39.2114
R20284 vdd.n2309 vdd.n756 39.2114
R20285 vdd.n2313 vdd.n755 39.2114
R20286 vdd.n2317 vdd.n754 39.2114
R20287 vdd.n2321 vdd.n753 39.2114
R20288 vdd.n1073 vdd.n948 39.2114
R20289 vdd.n1077 vdd.n949 39.2114
R20290 vdd.n1081 vdd.n950 39.2114
R20291 vdd.n1085 vdd.n951 39.2114
R20292 vdd.n1089 vdd.n952 39.2114
R20293 vdd.n1093 vdd.n953 39.2114
R20294 vdd.n1097 vdd.n954 39.2114
R20295 vdd.n1101 vdd.n955 39.2114
R20296 vdd.n1104 vdd.n956 39.2114
R20297 vdd.n1301 vdd.n957 39.2114
R20298 vdd.n1297 vdd.n958 39.2114
R20299 vdd.n1293 vdd.n959 39.2114
R20300 vdd.n1289 vdd.n960 39.2114
R20301 vdd.n1285 vdd.n961 39.2114
R20302 vdd.n1281 vdd.n962 39.2114
R20303 vdd.n1277 vdd.n963 39.2114
R20304 vdd.n1273 vdd.n964 39.2114
R20305 vdd.n1978 vdd.n1977 37.2369
R20306 vdd.n2014 vdd.n1039 37.2369
R20307 vdd.n2053 vdd.n999 37.2369
R20308 vdd.n3030 vdd.n558 37.2369
R20309 vdd.n3078 vdd.n3077 37.2369
R20310 vdd.n2985 vdd.n2984 37.2369
R20311 vdd.n1107 vdd.n1106 30.449
R20312 vdd.n802 vdd.n801 30.449
R20313 vdd.n1138 vdd.n1110 30.449
R20314 vdd.n2334 vdd.n792 30.449
R20315 vdd.n2439 vdd.n2438 30.449
R20316 vdd.n2886 vdd.n623 30.449
R20317 vdd.n2642 vdd.n2435 30.449
R20318 vdd.n591 vdd.n590 30.449
R20319 vdd.n2124 vdd.n2123 29.8151
R20320 vdd.n2396 vdd.n790 29.8151
R20321 vdd.n2329 vdd.n793 29.8151
R20322 vdd.n1146 vdd.n1143 29.8151
R20323 vdd.n2637 vdd.n2634 29.8151
R20324 vdd.n2880 vdd.n2879 29.8151
R20325 vdd.n2706 vdd.n2705 29.8151
R20326 vdd.n2943 vdd.n2942 29.8151
R20327 vdd.n2862 vdd.n2861 29.8151
R20328 vdd.n2948 vdd.n592 29.8151
R20329 vdd.n2510 vdd.n2508 29.8151
R20330 vdd.n2441 vdd.n745 29.8151
R20331 vdd.n1071 vdd.n922 29.8151
R20332 vdd.n2324 vdd.n2323 29.8151
R20333 vdd.n2256 vdd.n2255 29.8151
R20334 vdd.n1272 vdd.n1271 29.8151
R20335 vdd.n1876 vdd.n1683 22.6735
R20336 vdd.n1972 vdd.n931 22.6735
R20337 vdd.n3112 vdd.n516 22.6735
R20338 vdd.n3297 vdd.n329 22.6735
R20339 vdd.n1887 vdd.n1645 19.3944
R20340 vdd.n1887 vdd.n1643 19.3944
R20341 vdd.n1891 vdd.n1643 19.3944
R20342 vdd.n1891 vdd.n1633 19.3944
R20343 vdd.n1904 vdd.n1633 19.3944
R20344 vdd.n1904 vdd.n1631 19.3944
R20345 vdd.n1908 vdd.n1631 19.3944
R20346 vdd.n1908 vdd.n1623 19.3944
R20347 vdd.n1922 vdd.n1623 19.3944
R20348 vdd.n1922 vdd.n1621 19.3944
R20349 vdd.n1926 vdd.n1621 19.3944
R20350 vdd.n1926 vdd.n1340 19.3944
R20351 vdd.n1938 vdd.n1340 19.3944
R20352 vdd.n1938 vdd.n1338 19.3944
R20353 vdd.n1942 vdd.n1338 19.3944
R20354 vdd.n1942 vdd.n1330 19.3944
R20355 vdd.n1955 vdd.n1330 19.3944
R20356 vdd.n1955 vdd.n1327 19.3944
R20357 vdd.n1961 vdd.n1327 19.3944
R20358 vdd.n1961 vdd.n1328 19.3944
R20359 vdd.n1328 vdd.n1318 19.3944
R20360 vdd.n1811 vdd.n1746 19.3944
R20361 vdd.n1807 vdd.n1746 19.3944
R20362 vdd.n1807 vdd.n1806 19.3944
R20363 vdd.n1806 vdd.n1805 19.3944
R20364 vdd.n1805 vdd.n1752 19.3944
R20365 vdd.n1801 vdd.n1752 19.3944
R20366 vdd.n1801 vdd.n1800 19.3944
R20367 vdd.n1800 vdd.n1799 19.3944
R20368 vdd.n1799 vdd.n1758 19.3944
R20369 vdd.n1795 vdd.n1758 19.3944
R20370 vdd.n1795 vdd.n1794 19.3944
R20371 vdd.n1794 vdd.n1793 19.3944
R20372 vdd.n1793 vdd.n1764 19.3944
R20373 vdd.n1789 vdd.n1764 19.3944
R20374 vdd.n1789 vdd.n1788 19.3944
R20375 vdd.n1788 vdd.n1787 19.3944
R20376 vdd.n1787 vdd.n1770 19.3944
R20377 vdd.n1783 vdd.n1770 19.3944
R20378 vdd.n1783 vdd.n1782 19.3944
R20379 vdd.n1782 vdd.n1781 19.3944
R20380 vdd.n1846 vdd.n1845 19.3944
R20381 vdd.n1845 vdd.n1844 19.3944
R20382 vdd.n1844 vdd.n1717 19.3944
R20383 vdd.n1840 vdd.n1717 19.3944
R20384 vdd.n1840 vdd.n1839 19.3944
R20385 vdd.n1839 vdd.n1838 19.3944
R20386 vdd.n1838 vdd.n1723 19.3944
R20387 vdd.n1834 vdd.n1723 19.3944
R20388 vdd.n1834 vdd.n1833 19.3944
R20389 vdd.n1833 vdd.n1832 19.3944
R20390 vdd.n1832 vdd.n1729 19.3944
R20391 vdd.n1828 vdd.n1729 19.3944
R20392 vdd.n1828 vdd.n1827 19.3944
R20393 vdd.n1827 vdd.n1826 19.3944
R20394 vdd.n1826 vdd.n1735 19.3944
R20395 vdd.n1822 vdd.n1735 19.3944
R20396 vdd.n1822 vdd.n1821 19.3944
R20397 vdd.n1821 vdd.n1820 19.3944
R20398 vdd.n1820 vdd.n1741 19.3944
R20399 vdd.n1816 vdd.n1741 19.3944
R20400 vdd.n1879 vdd.n1650 19.3944
R20401 vdd.n1874 vdd.n1650 19.3944
R20402 vdd.n1874 vdd.n1685 19.3944
R20403 vdd.n1870 vdd.n1685 19.3944
R20404 vdd.n1870 vdd.n1869 19.3944
R20405 vdd.n1869 vdd.n1868 19.3944
R20406 vdd.n1868 vdd.n1691 19.3944
R20407 vdd.n1864 vdd.n1691 19.3944
R20408 vdd.n1864 vdd.n1863 19.3944
R20409 vdd.n1863 vdd.n1862 19.3944
R20410 vdd.n1862 vdd.n1697 19.3944
R20411 vdd.n1858 vdd.n1697 19.3944
R20412 vdd.n1858 vdd.n1857 19.3944
R20413 vdd.n1857 vdd.n1856 19.3944
R20414 vdd.n1856 vdd.n1703 19.3944
R20415 vdd.n1852 vdd.n1703 19.3944
R20416 vdd.n1852 vdd.n1851 19.3944
R20417 vdd.n1851 vdd.n1850 19.3944
R20418 vdd.n2010 vdd.n1037 19.3944
R20419 vdd.n2010 vdd.n1043 19.3944
R20420 vdd.n2005 vdd.n1043 19.3944
R20421 vdd.n2005 vdd.n2004 19.3944
R20422 vdd.n2004 vdd.n2003 19.3944
R20423 vdd.n2003 vdd.n1050 19.3944
R20424 vdd.n1998 vdd.n1050 19.3944
R20425 vdd.n1998 vdd.n1997 19.3944
R20426 vdd.n1997 vdd.n1996 19.3944
R20427 vdd.n1996 vdd.n1057 19.3944
R20428 vdd.n1991 vdd.n1057 19.3944
R20429 vdd.n1991 vdd.n1990 19.3944
R20430 vdd.n1990 vdd.n1989 19.3944
R20431 vdd.n1989 vdd.n1064 19.3944
R20432 vdd.n1984 vdd.n1064 19.3944
R20433 vdd.n1984 vdd.n1983 19.3944
R20434 vdd.n1311 vdd.n1069 19.3944
R20435 vdd.n1979 vdd.n1308 19.3944
R20436 vdd.n2049 vdd.n997 19.3944
R20437 vdd.n2049 vdd.n1003 19.3944
R20438 vdd.n2044 vdd.n1003 19.3944
R20439 vdd.n2044 vdd.n2043 19.3944
R20440 vdd.n2043 vdd.n2042 19.3944
R20441 vdd.n2042 vdd.n1010 19.3944
R20442 vdd.n2037 vdd.n1010 19.3944
R20443 vdd.n2037 vdd.n2036 19.3944
R20444 vdd.n2036 vdd.n2035 19.3944
R20445 vdd.n2035 vdd.n1017 19.3944
R20446 vdd.n2030 vdd.n1017 19.3944
R20447 vdd.n2030 vdd.n2029 19.3944
R20448 vdd.n2029 vdd.n2028 19.3944
R20449 vdd.n2028 vdd.n1024 19.3944
R20450 vdd.n2023 vdd.n1024 19.3944
R20451 vdd.n2023 vdd.n2022 19.3944
R20452 vdd.n2022 vdd.n2021 19.3944
R20453 vdd.n2021 vdd.n1031 19.3944
R20454 vdd.n2016 vdd.n1031 19.3944
R20455 vdd.n2016 vdd.n2015 19.3944
R20456 vdd.n2086 vdd.n972 19.3944
R20457 vdd.n2086 vdd.n973 19.3944
R20458 vdd.n2081 vdd.n2080 19.3944
R20459 vdd.n2076 vdd.n2075 19.3944
R20460 vdd.n2075 vdd.n2074 19.3944
R20461 vdd.n2074 vdd.n977 19.3944
R20462 vdd.n2069 vdd.n977 19.3944
R20463 vdd.n2069 vdd.n2068 19.3944
R20464 vdd.n2068 vdd.n2067 19.3944
R20465 vdd.n2067 vdd.n984 19.3944
R20466 vdd.n2062 vdd.n984 19.3944
R20467 vdd.n2062 vdd.n2061 19.3944
R20468 vdd.n2061 vdd.n2060 19.3944
R20469 vdd.n2060 vdd.n991 19.3944
R20470 vdd.n2055 vdd.n991 19.3944
R20471 vdd.n2055 vdd.n2054 19.3944
R20472 vdd.n1883 vdd.n1648 19.3944
R20473 vdd.n1883 vdd.n1639 19.3944
R20474 vdd.n1896 vdd.n1639 19.3944
R20475 vdd.n1896 vdd.n1637 19.3944
R20476 vdd.n1900 vdd.n1637 19.3944
R20477 vdd.n1900 vdd.n1628 19.3944
R20478 vdd.n1913 vdd.n1628 19.3944
R20479 vdd.n1913 vdd.n1626 19.3944
R20480 vdd.n1918 vdd.n1626 19.3944
R20481 vdd.n1918 vdd.n1617 19.3944
R20482 vdd.n1930 vdd.n1617 19.3944
R20483 vdd.n1930 vdd.n1345 19.3944
R20484 vdd.n1934 vdd.n1345 19.3944
R20485 vdd.n1934 vdd.n1335 19.3944
R20486 vdd.n1947 vdd.n1335 19.3944
R20487 vdd.n1947 vdd.n1333 19.3944
R20488 vdd.n1951 vdd.n1333 19.3944
R20489 vdd.n1951 vdd.n1323 19.3944
R20490 vdd.n1966 vdd.n1323 19.3944
R20491 vdd.n1966 vdd.n1321 19.3944
R20492 vdd.n1970 vdd.n1321 19.3944
R20493 vdd.n3123 vdd.n477 19.3944
R20494 vdd.n3123 vdd.n475 19.3944
R20495 vdd.n3127 vdd.n475 19.3944
R20496 vdd.n3127 vdd.n465 19.3944
R20497 vdd.n3140 vdd.n465 19.3944
R20498 vdd.n3140 vdd.n463 19.3944
R20499 vdd.n3144 vdd.n463 19.3944
R20500 vdd.n3144 vdd.n453 19.3944
R20501 vdd.n3156 vdd.n453 19.3944
R20502 vdd.n3156 vdd.n451 19.3944
R20503 vdd.n3160 vdd.n451 19.3944
R20504 vdd.n3161 vdd.n3160 19.3944
R20505 vdd.n3162 vdd.n3161 19.3944
R20506 vdd.n3162 vdd.n449 19.3944
R20507 vdd.n3166 vdd.n449 19.3944
R20508 vdd.n3167 vdd.n3166 19.3944
R20509 vdd.n3168 vdd.n3167 19.3944
R20510 vdd.n3168 vdd.n446 19.3944
R20511 vdd.n3172 vdd.n446 19.3944
R20512 vdd.n3173 vdd.n3172 19.3944
R20513 vdd.n3174 vdd.n3173 19.3944
R20514 vdd.n3217 vdd.n404 19.3944
R20515 vdd.n3217 vdd.n410 19.3944
R20516 vdd.n3212 vdd.n410 19.3944
R20517 vdd.n3212 vdd.n3211 19.3944
R20518 vdd.n3211 vdd.n3210 19.3944
R20519 vdd.n3210 vdd.n417 19.3944
R20520 vdd.n3205 vdd.n417 19.3944
R20521 vdd.n3205 vdd.n3204 19.3944
R20522 vdd.n3204 vdd.n3203 19.3944
R20523 vdd.n3203 vdd.n424 19.3944
R20524 vdd.n3198 vdd.n424 19.3944
R20525 vdd.n3198 vdd.n3197 19.3944
R20526 vdd.n3197 vdd.n3196 19.3944
R20527 vdd.n3196 vdd.n431 19.3944
R20528 vdd.n3191 vdd.n431 19.3944
R20529 vdd.n3191 vdd.n3190 19.3944
R20530 vdd.n3190 vdd.n3189 19.3944
R20531 vdd.n3189 vdd.n438 19.3944
R20532 vdd.n3184 vdd.n438 19.3944
R20533 vdd.n3184 vdd.n3183 19.3944
R20534 vdd.n3256 vdd.n364 19.3944
R20535 vdd.n3256 vdd.n370 19.3944
R20536 vdd.n3251 vdd.n370 19.3944
R20537 vdd.n3251 vdd.n3250 19.3944
R20538 vdd.n3250 vdd.n3249 19.3944
R20539 vdd.n3249 vdd.n377 19.3944
R20540 vdd.n3244 vdd.n377 19.3944
R20541 vdd.n3244 vdd.n3243 19.3944
R20542 vdd.n3243 vdd.n3242 19.3944
R20543 vdd.n3242 vdd.n384 19.3944
R20544 vdd.n3237 vdd.n384 19.3944
R20545 vdd.n3237 vdd.n3236 19.3944
R20546 vdd.n3236 vdd.n3235 19.3944
R20547 vdd.n3235 vdd.n391 19.3944
R20548 vdd.n3230 vdd.n391 19.3944
R20549 vdd.n3230 vdd.n3229 19.3944
R20550 vdd.n3229 vdd.n3228 19.3944
R20551 vdd.n3228 vdd.n398 19.3944
R20552 vdd.n3223 vdd.n398 19.3944
R20553 vdd.n3223 vdd.n3222 19.3944
R20554 vdd.n3292 vdd.n3291 19.3944
R20555 vdd.n3291 vdd.n3290 19.3944
R20556 vdd.n3290 vdd.n336 19.3944
R20557 vdd.n337 vdd.n336 19.3944
R20558 vdd.n3283 vdd.n337 19.3944
R20559 vdd.n3283 vdd.n3282 19.3944
R20560 vdd.n3282 vdd.n3281 19.3944
R20561 vdd.n3281 vdd.n344 19.3944
R20562 vdd.n3276 vdd.n344 19.3944
R20563 vdd.n3276 vdd.n3275 19.3944
R20564 vdd.n3275 vdd.n3274 19.3944
R20565 vdd.n3274 vdd.n351 19.3944
R20566 vdd.n3269 vdd.n351 19.3944
R20567 vdd.n3269 vdd.n3268 19.3944
R20568 vdd.n3268 vdd.n3267 19.3944
R20569 vdd.n3267 vdd.n358 19.3944
R20570 vdd.n3262 vdd.n358 19.3944
R20571 vdd.n3262 vdd.n3261 19.3944
R20572 vdd.n3119 vdd.n480 19.3944
R20573 vdd.n3119 vdd.n471 19.3944
R20574 vdd.n3132 vdd.n471 19.3944
R20575 vdd.n3132 vdd.n469 19.3944
R20576 vdd.n3136 vdd.n469 19.3944
R20577 vdd.n3136 vdd.n460 19.3944
R20578 vdd.n3148 vdd.n460 19.3944
R20579 vdd.n3148 vdd.n458 19.3944
R20580 vdd.n3152 vdd.n458 19.3944
R20581 vdd.n3152 vdd.n300 19.3944
R20582 vdd.n3317 vdd.n300 19.3944
R20583 vdd.n3317 vdd.n301 19.3944
R20584 vdd.n3311 vdd.n301 19.3944
R20585 vdd.n3311 vdd.n3310 19.3944
R20586 vdd.n3310 vdd.n3309 19.3944
R20587 vdd.n3309 vdd.n313 19.3944
R20588 vdd.n3303 vdd.n313 19.3944
R20589 vdd.n3303 vdd.n3302 19.3944
R20590 vdd.n3302 vdd.n3301 19.3944
R20591 vdd.n3301 vdd.n324 19.3944
R20592 vdd.n3295 vdd.n324 19.3944
R20593 vdd.n3072 vdd.n536 19.3944
R20594 vdd.n3072 vdd.n3069 19.3944
R20595 vdd.n3069 vdd.n3066 19.3944
R20596 vdd.n3066 vdd.n3065 19.3944
R20597 vdd.n3065 vdd.n3062 19.3944
R20598 vdd.n3062 vdd.n3061 19.3944
R20599 vdd.n3061 vdd.n3058 19.3944
R20600 vdd.n3058 vdd.n3057 19.3944
R20601 vdd.n3057 vdd.n3054 19.3944
R20602 vdd.n3054 vdd.n3053 19.3944
R20603 vdd.n3053 vdd.n3050 19.3944
R20604 vdd.n3050 vdd.n3049 19.3944
R20605 vdd.n3049 vdd.n3046 19.3944
R20606 vdd.n3046 vdd.n3045 19.3944
R20607 vdd.n3045 vdd.n3042 19.3944
R20608 vdd.n3042 vdd.n3041 19.3944
R20609 vdd.n3041 vdd.n3038 19.3944
R20610 vdd.n3038 vdd.n3037 19.3944
R20611 vdd.n3037 vdd.n3034 19.3944
R20612 vdd.n3034 vdd.n3033 19.3944
R20613 vdd.n3115 vdd.n482 19.3944
R20614 vdd.n3110 vdd.n482 19.3944
R20615 vdd.n521 vdd.n518 19.3944
R20616 vdd.n3106 vdd.n3105 19.3944
R20617 vdd.n3105 vdd.n3102 19.3944
R20618 vdd.n3102 vdd.n3101 19.3944
R20619 vdd.n3101 vdd.n3098 19.3944
R20620 vdd.n3098 vdd.n3097 19.3944
R20621 vdd.n3097 vdd.n3094 19.3944
R20622 vdd.n3094 vdd.n3093 19.3944
R20623 vdd.n3093 vdd.n3090 19.3944
R20624 vdd.n3090 vdd.n3089 19.3944
R20625 vdd.n3089 vdd.n3086 19.3944
R20626 vdd.n3086 vdd.n3085 19.3944
R20627 vdd.n3085 vdd.n3082 19.3944
R20628 vdd.n3082 vdd.n3081 19.3944
R20629 vdd.n3026 vdd.n556 19.3944
R20630 vdd.n3026 vdd.n3023 19.3944
R20631 vdd.n3023 vdd.n3020 19.3944
R20632 vdd.n3020 vdd.n3019 19.3944
R20633 vdd.n3019 vdd.n3016 19.3944
R20634 vdd.n3016 vdd.n3015 19.3944
R20635 vdd.n3015 vdd.n3012 19.3944
R20636 vdd.n3012 vdd.n3011 19.3944
R20637 vdd.n3011 vdd.n3008 19.3944
R20638 vdd.n3008 vdd.n3007 19.3944
R20639 vdd.n3007 vdd.n3004 19.3944
R20640 vdd.n3004 vdd.n3003 19.3944
R20641 vdd.n3003 vdd.n3000 19.3944
R20642 vdd.n3000 vdd.n2999 19.3944
R20643 vdd.n2999 vdd.n2996 19.3944
R20644 vdd.n2996 vdd.n2995 19.3944
R20645 vdd.n2992 vdd.n2991 19.3944
R20646 vdd.n2988 vdd.n2987 19.3944
R20647 vdd.n1815 vdd.n1811 19.0066
R20648 vdd.n2014 vdd.n1037 19.0066
R20649 vdd.n3221 vdd.n404 19.0066
R20650 vdd.n3030 vdd.n556 19.0066
R20651 vdd.n1106 vdd.n1105 16.0975
R20652 vdd.n801 vdd.n800 16.0975
R20653 vdd.n1776 vdd.n1775 16.0975
R20654 vdd.n1814 vdd.n1813 16.0975
R20655 vdd.n1710 vdd.n1709 16.0975
R20656 vdd.n1977 vdd.n1976 16.0975
R20657 vdd.n1039 vdd.n1038 16.0975
R20658 vdd.n999 vdd.n998 16.0975
R20659 vdd.n1110 vdd.n1109 16.0975
R20660 vdd.n792 vdd.n791 16.0975
R20661 vdd.n2438 vdd.n2437 16.0975
R20662 vdd.n3181 vdd.n3180 16.0975
R20663 vdd.n406 vdd.n405 16.0975
R20664 vdd.n366 vdd.n365 16.0975
R20665 vdd.n558 vdd.n557 16.0975
R20666 vdd.n3077 vdd.n3076 16.0975
R20667 vdd.n623 vdd.n622 16.0975
R20668 vdd.n2435 vdd.n2434 16.0975
R20669 vdd.n2984 vdd.n2983 16.0975
R20670 vdd.n590 vdd.n589 16.0975
R20671 vdd.t184 vdd.n2398 15.4182
R20672 vdd.n2702 vdd.t166 15.4182
R20673 vdd.n28 vdd.n27 14.5674
R20674 vdd.n292 vdd.n257 13.1884
R20675 vdd.n245 vdd.n210 13.1884
R20676 vdd.n202 vdd.n167 13.1884
R20677 vdd.n155 vdd.n120 13.1884
R20678 vdd.n113 vdd.n78 13.1884
R20679 vdd.n66 vdd.n31 13.1884
R20680 vdd.n1562 vdd.n1527 13.1884
R20681 vdd.n1609 vdd.n1574 13.1884
R20682 vdd.n1472 vdd.n1437 13.1884
R20683 vdd.n1519 vdd.n1484 13.1884
R20684 vdd.n1383 vdd.n1348 13.1884
R20685 vdd.n1430 vdd.n1395 13.1884
R20686 vdd.n2120 vdd.n924 13.1509
R20687 vdd.n2945 vdd.n484 13.1509
R20688 vdd.n1846 vdd.n1711 12.9944
R20689 vdd.n1850 vdd.n1711 12.9944
R20690 vdd.n2053 vdd.n997 12.9944
R20691 vdd.n2054 vdd.n2053 12.9944
R20692 vdd.n3260 vdd.n364 12.9944
R20693 vdd.n3261 vdd.n3260 12.9944
R20694 vdd.n3078 vdd.n536 12.9944
R20695 vdd.n3081 vdd.n3078 12.9944
R20696 vdd.n293 vdd.n255 12.8005
R20697 vdd.n288 vdd.n259 12.8005
R20698 vdd.n246 vdd.n208 12.8005
R20699 vdd.n241 vdd.n212 12.8005
R20700 vdd.n203 vdd.n165 12.8005
R20701 vdd.n198 vdd.n169 12.8005
R20702 vdd.n156 vdd.n118 12.8005
R20703 vdd.n151 vdd.n122 12.8005
R20704 vdd.n114 vdd.n76 12.8005
R20705 vdd.n109 vdd.n80 12.8005
R20706 vdd.n67 vdd.n29 12.8005
R20707 vdd.n62 vdd.n33 12.8005
R20708 vdd.n1563 vdd.n1525 12.8005
R20709 vdd.n1558 vdd.n1529 12.8005
R20710 vdd.n1610 vdd.n1572 12.8005
R20711 vdd.n1605 vdd.n1576 12.8005
R20712 vdd.n1473 vdd.n1435 12.8005
R20713 vdd.n1468 vdd.n1439 12.8005
R20714 vdd.n1520 vdd.n1482 12.8005
R20715 vdd.n1515 vdd.n1486 12.8005
R20716 vdd.n1384 vdd.n1346 12.8005
R20717 vdd.n1379 vdd.n1350 12.8005
R20718 vdd.n1431 vdd.n1393 12.8005
R20719 vdd.n1426 vdd.n1397 12.8005
R20720 vdd.n287 vdd.n260 12.0247
R20721 vdd.n240 vdd.n213 12.0247
R20722 vdd.n197 vdd.n170 12.0247
R20723 vdd.n150 vdd.n123 12.0247
R20724 vdd.n108 vdd.n81 12.0247
R20725 vdd.n61 vdd.n34 12.0247
R20726 vdd.n1557 vdd.n1530 12.0247
R20727 vdd.n1604 vdd.n1577 12.0247
R20728 vdd.n1467 vdd.n1440 12.0247
R20729 vdd.n1514 vdd.n1487 12.0247
R20730 vdd.n1378 vdd.n1351 12.0247
R20731 vdd.n1425 vdd.n1398 12.0247
R20732 vdd.n1885 vdd.n1641 11.337
R20733 vdd.n1894 vdd.n1641 11.337
R20734 vdd.n1894 vdd.n1893 11.337
R20735 vdd.n1902 vdd.n1635 11.337
R20736 vdd.n1911 vdd.n1910 11.337
R20737 vdd.n1928 vdd.n1619 11.337
R20738 vdd.n1936 vdd.n1342 11.337
R20739 vdd.n1945 vdd.n1944 11.337
R20740 vdd.n1953 vdd.n1325 11.337
R20741 vdd.n1964 vdd.n1325 11.337
R20742 vdd.n1964 vdd.n1963 11.337
R20743 vdd.n3121 vdd.n473 11.337
R20744 vdd.n3130 vdd.n473 11.337
R20745 vdd.n3130 vdd.n3129 11.337
R20746 vdd.n3138 vdd.n467 11.337
R20747 vdd.n3154 vdd.n456 11.337
R20748 vdd.n3315 vdd.n304 11.337
R20749 vdd.n3313 vdd.n308 11.337
R20750 vdd.n3307 vdd.n3306 11.337
R20751 vdd.n3305 vdd.n318 11.337
R20752 vdd.n3299 vdd.n318 11.337
R20753 vdd.n3299 vdd.n3298 11.337
R20754 vdd.n284 vdd.n283 11.249
R20755 vdd.n237 vdd.n236 11.249
R20756 vdd.n194 vdd.n193 11.249
R20757 vdd.n147 vdd.n146 11.249
R20758 vdd.n105 vdd.n104 11.249
R20759 vdd.n58 vdd.n57 11.249
R20760 vdd.n1554 vdd.n1553 11.249
R20761 vdd.n1601 vdd.n1600 11.249
R20762 vdd.n1464 vdd.n1463 11.249
R20763 vdd.n1511 vdd.n1510 11.249
R20764 vdd.n1375 vdd.n1374 11.249
R20765 vdd.n1422 vdd.n1421 11.249
R20766 vdd.n1683 vdd.t43 10.7702
R20767 vdd.t50 vdd.n3297 10.7702
R20768 vdd.n269 vdd.n268 10.7238
R20769 vdd.n222 vdd.n221 10.7238
R20770 vdd.n179 vdd.n178 10.7238
R20771 vdd.n132 vdd.n131 10.7238
R20772 vdd.n90 vdd.n89 10.7238
R20773 vdd.n43 vdd.n42 10.7238
R20774 vdd.n1539 vdd.n1538 10.7238
R20775 vdd.n1586 vdd.n1585 10.7238
R20776 vdd.n1449 vdd.n1448 10.7238
R20777 vdd.n1496 vdd.n1495 10.7238
R20778 vdd.n1360 vdd.n1359 10.7238
R20779 vdd.n1407 vdd.n1406 10.7238
R20780 vdd.n2125 vdd.n2124 10.6151
R20781 vdd.n2125 vdd.n917 10.6151
R20782 vdd.n2135 vdd.n917 10.6151
R20783 vdd.n2136 vdd.n2135 10.6151
R20784 vdd.n2137 vdd.n2136 10.6151
R20785 vdd.n2137 vdd.n904 10.6151
R20786 vdd.n2147 vdd.n904 10.6151
R20787 vdd.n2148 vdd.n2147 10.6151
R20788 vdd.n2149 vdd.n2148 10.6151
R20789 vdd.n2149 vdd.n892 10.6151
R20790 vdd.n2159 vdd.n892 10.6151
R20791 vdd.n2160 vdd.n2159 10.6151
R20792 vdd.n2161 vdd.n2160 10.6151
R20793 vdd.n2161 vdd.n881 10.6151
R20794 vdd.n2171 vdd.n881 10.6151
R20795 vdd.n2172 vdd.n2171 10.6151
R20796 vdd.n2173 vdd.n2172 10.6151
R20797 vdd.n2173 vdd.n868 10.6151
R20798 vdd.n2183 vdd.n868 10.6151
R20799 vdd.n2184 vdd.n2183 10.6151
R20800 vdd.n2185 vdd.n2184 10.6151
R20801 vdd.n2185 vdd.n856 10.6151
R20802 vdd.n2196 vdd.n856 10.6151
R20803 vdd.n2197 vdd.n2196 10.6151
R20804 vdd.n2198 vdd.n2197 10.6151
R20805 vdd.n2198 vdd.n844 10.6151
R20806 vdd.n2208 vdd.n844 10.6151
R20807 vdd.n2209 vdd.n2208 10.6151
R20808 vdd.n2210 vdd.n2209 10.6151
R20809 vdd.n2210 vdd.n832 10.6151
R20810 vdd.n2220 vdd.n832 10.6151
R20811 vdd.n2221 vdd.n2220 10.6151
R20812 vdd.n2222 vdd.n2221 10.6151
R20813 vdd.n2222 vdd.n822 10.6151
R20814 vdd.n2232 vdd.n822 10.6151
R20815 vdd.n2233 vdd.n2232 10.6151
R20816 vdd.n2234 vdd.n2233 10.6151
R20817 vdd.n2234 vdd.n809 10.6151
R20818 vdd.n2246 vdd.n809 10.6151
R20819 vdd.n2247 vdd.n2246 10.6151
R20820 vdd.n2249 vdd.n2247 10.6151
R20821 vdd.n2249 vdd.n2248 10.6151
R20822 vdd.n2248 vdd.n790 10.6151
R20823 vdd.n2396 vdd.n2395 10.6151
R20824 vdd.n2395 vdd.n2394 10.6151
R20825 vdd.n2394 vdd.n2391 10.6151
R20826 vdd.n2391 vdd.n2390 10.6151
R20827 vdd.n2390 vdd.n2387 10.6151
R20828 vdd.n2387 vdd.n2386 10.6151
R20829 vdd.n2386 vdd.n2383 10.6151
R20830 vdd.n2383 vdd.n2382 10.6151
R20831 vdd.n2382 vdd.n2379 10.6151
R20832 vdd.n2379 vdd.n2378 10.6151
R20833 vdd.n2378 vdd.n2375 10.6151
R20834 vdd.n2375 vdd.n2374 10.6151
R20835 vdd.n2374 vdd.n2371 10.6151
R20836 vdd.n2371 vdd.n2370 10.6151
R20837 vdd.n2370 vdd.n2367 10.6151
R20838 vdd.n2367 vdd.n2366 10.6151
R20839 vdd.n2366 vdd.n2363 10.6151
R20840 vdd.n2363 vdd.n2362 10.6151
R20841 vdd.n2362 vdd.n2359 10.6151
R20842 vdd.n2359 vdd.n2358 10.6151
R20843 vdd.n2358 vdd.n2355 10.6151
R20844 vdd.n2355 vdd.n2354 10.6151
R20845 vdd.n2354 vdd.n2351 10.6151
R20846 vdd.n2351 vdd.n2350 10.6151
R20847 vdd.n2350 vdd.n2347 10.6151
R20848 vdd.n2347 vdd.n2346 10.6151
R20849 vdd.n2346 vdd.n2343 10.6151
R20850 vdd.n2343 vdd.n2342 10.6151
R20851 vdd.n2342 vdd.n2339 10.6151
R20852 vdd.n2339 vdd.n2338 10.6151
R20853 vdd.n2338 vdd.n2335 10.6151
R20854 vdd.n2333 vdd.n2330 10.6151
R20855 vdd.n2330 vdd.n2329 10.6151
R20856 vdd.n1147 vdd.n1146 10.6151
R20857 vdd.n1149 vdd.n1147 10.6151
R20858 vdd.n1150 vdd.n1149 10.6151
R20859 vdd.n1152 vdd.n1150 10.6151
R20860 vdd.n1153 vdd.n1152 10.6151
R20861 vdd.n1155 vdd.n1153 10.6151
R20862 vdd.n1156 vdd.n1155 10.6151
R20863 vdd.n1158 vdd.n1156 10.6151
R20864 vdd.n1159 vdd.n1158 10.6151
R20865 vdd.n1161 vdd.n1159 10.6151
R20866 vdd.n1162 vdd.n1161 10.6151
R20867 vdd.n1164 vdd.n1162 10.6151
R20868 vdd.n1165 vdd.n1164 10.6151
R20869 vdd.n1167 vdd.n1165 10.6151
R20870 vdd.n1168 vdd.n1167 10.6151
R20871 vdd.n1170 vdd.n1168 10.6151
R20872 vdd.n1171 vdd.n1170 10.6151
R20873 vdd.n1173 vdd.n1171 10.6151
R20874 vdd.n1174 vdd.n1173 10.6151
R20875 vdd.n1176 vdd.n1174 10.6151
R20876 vdd.n1177 vdd.n1176 10.6151
R20877 vdd.n1179 vdd.n1177 10.6151
R20878 vdd.n1180 vdd.n1179 10.6151
R20879 vdd.n1182 vdd.n1180 10.6151
R20880 vdd.n1183 vdd.n1182 10.6151
R20881 vdd.n1185 vdd.n1183 10.6151
R20882 vdd.n1186 vdd.n1185 10.6151
R20883 vdd.n1225 vdd.n1186 10.6151
R20884 vdd.n1225 vdd.n1224 10.6151
R20885 vdd.n1224 vdd.n1223 10.6151
R20886 vdd.n1223 vdd.n1221 10.6151
R20887 vdd.n1221 vdd.n1220 10.6151
R20888 vdd.n1220 vdd.n1218 10.6151
R20889 vdd.n1218 vdd.n1217 10.6151
R20890 vdd.n1217 vdd.n1198 10.6151
R20891 vdd.n1198 vdd.n1197 10.6151
R20892 vdd.n1197 vdd.n1195 10.6151
R20893 vdd.n1195 vdd.n1194 10.6151
R20894 vdd.n1194 vdd.n1192 10.6151
R20895 vdd.n1192 vdd.n1191 10.6151
R20896 vdd.n1191 vdd.n1188 10.6151
R20897 vdd.n1188 vdd.n1187 10.6151
R20898 vdd.n1187 vdd.n793 10.6151
R20899 vdd.n2123 vdd.n929 10.6151
R20900 vdd.n2118 vdd.n929 10.6151
R20901 vdd.n2118 vdd.n2117 10.6151
R20902 vdd.n2117 vdd.n2116 10.6151
R20903 vdd.n2116 vdd.n2113 10.6151
R20904 vdd.n2113 vdd.n2112 10.6151
R20905 vdd.n2112 vdd.n2109 10.6151
R20906 vdd.n2109 vdd.n2108 10.6151
R20907 vdd.n2108 vdd.n2105 10.6151
R20908 vdd.n2105 vdd.n2104 10.6151
R20909 vdd.n2104 vdd.n2101 10.6151
R20910 vdd.n2101 vdd.n2100 10.6151
R20911 vdd.n2100 vdd.n2097 10.6151
R20912 vdd.n2097 vdd.n2096 10.6151
R20913 vdd.n2096 vdd.n2093 10.6151
R20914 vdd.n2093 vdd.n2092 10.6151
R20915 vdd.n2092 vdd.n2089 10.6151
R20916 vdd.n2089 vdd.n967 10.6151
R20917 vdd.n1113 vdd.n967 10.6151
R20918 vdd.n1114 vdd.n1113 10.6151
R20919 vdd.n1117 vdd.n1114 10.6151
R20920 vdd.n1118 vdd.n1117 10.6151
R20921 vdd.n1121 vdd.n1118 10.6151
R20922 vdd.n1122 vdd.n1121 10.6151
R20923 vdd.n1125 vdd.n1122 10.6151
R20924 vdd.n1126 vdd.n1125 10.6151
R20925 vdd.n1129 vdd.n1126 10.6151
R20926 vdd.n1130 vdd.n1129 10.6151
R20927 vdd.n1133 vdd.n1130 10.6151
R20928 vdd.n1134 vdd.n1133 10.6151
R20929 vdd.n1137 vdd.n1134 10.6151
R20930 vdd.n1142 vdd.n1139 10.6151
R20931 vdd.n1143 vdd.n1142 10.6151
R20932 vdd.n2634 vdd.n2633 10.6151
R20933 vdd.n2633 vdd.n2632 10.6151
R20934 vdd.n2632 vdd.n2436 10.6151
R20935 vdd.n2514 vdd.n2436 10.6151
R20936 vdd.n2515 vdd.n2514 10.6151
R20937 vdd.n2517 vdd.n2515 10.6151
R20938 vdd.n2518 vdd.n2517 10.6151
R20939 vdd.n2616 vdd.n2518 10.6151
R20940 vdd.n2616 vdd.n2615 10.6151
R20941 vdd.n2615 vdd.n2614 10.6151
R20942 vdd.n2614 vdd.n2562 10.6151
R20943 vdd.n2562 vdd.n2561 10.6151
R20944 vdd.n2561 vdd.n2559 10.6151
R20945 vdd.n2559 vdd.n2558 10.6151
R20946 vdd.n2558 vdd.n2556 10.6151
R20947 vdd.n2556 vdd.n2555 10.6151
R20948 vdd.n2555 vdd.n2553 10.6151
R20949 vdd.n2553 vdd.n2552 10.6151
R20950 vdd.n2552 vdd.n2550 10.6151
R20951 vdd.n2550 vdd.n2549 10.6151
R20952 vdd.n2549 vdd.n2547 10.6151
R20953 vdd.n2547 vdd.n2546 10.6151
R20954 vdd.n2546 vdd.n2544 10.6151
R20955 vdd.n2544 vdd.n2543 10.6151
R20956 vdd.n2543 vdd.n2541 10.6151
R20957 vdd.n2541 vdd.n2540 10.6151
R20958 vdd.n2540 vdd.n2538 10.6151
R20959 vdd.n2538 vdd.n2537 10.6151
R20960 vdd.n2537 vdd.n2535 10.6151
R20961 vdd.n2535 vdd.n2534 10.6151
R20962 vdd.n2534 vdd.n2532 10.6151
R20963 vdd.n2532 vdd.n2531 10.6151
R20964 vdd.n2531 vdd.n2529 10.6151
R20965 vdd.n2529 vdd.n2528 10.6151
R20966 vdd.n2528 vdd.n2526 10.6151
R20967 vdd.n2526 vdd.n2525 10.6151
R20968 vdd.n2525 vdd.n2523 10.6151
R20969 vdd.n2523 vdd.n2522 10.6151
R20970 vdd.n2522 vdd.n2520 10.6151
R20971 vdd.n2520 vdd.n2519 10.6151
R20972 vdd.n2519 vdd.n626 10.6151
R20973 vdd.n2878 vdd.n626 10.6151
R20974 vdd.n2879 vdd.n2878 10.6151
R20975 vdd.n2705 vdd.n751 10.6151
R20976 vdd.n2700 vdd.n751 10.6151
R20977 vdd.n2700 vdd.n2699 10.6151
R20978 vdd.n2699 vdd.n2698 10.6151
R20979 vdd.n2698 vdd.n2695 10.6151
R20980 vdd.n2695 vdd.n2694 10.6151
R20981 vdd.n2694 vdd.n2691 10.6151
R20982 vdd.n2691 vdd.n2690 10.6151
R20983 vdd.n2690 vdd.n2687 10.6151
R20984 vdd.n2687 vdd.n2686 10.6151
R20985 vdd.n2686 vdd.n2683 10.6151
R20986 vdd.n2683 vdd.n2682 10.6151
R20987 vdd.n2682 vdd.n2679 10.6151
R20988 vdd.n2679 vdd.n2678 10.6151
R20989 vdd.n2678 vdd.n2675 10.6151
R20990 vdd.n2675 vdd.n2674 10.6151
R20991 vdd.n2674 vdd.n2671 10.6151
R20992 vdd.n2671 vdd.n2670 10.6151
R20993 vdd.n2670 vdd.n2667 10.6151
R20994 vdd.n2667 vdd.n2666 10.6151
R20995 vdd.n2666 vdd.n2663 10.6151
R20996 vdd.n2663 vdd.n2662 10.6151
R20997 vdd.n2662 vdd.n2659 10.6151
R20998 vdd.n2659 vdd.n2658 10.6151
R20999 vdd.n2658 vdd.n2655 10.6151
R21000 vdd.n2655 vdd.n2654 10.6151
R21001 vdd.n2654 vdd.n2651 10.6151
R21002 vdd.n2651 vdd.n2650 10.6151
R21003 vdd.n2650 vdd.n2647 10.6151
R21004 vdd.n2647 vdd.n2646 10.6151
R21005 vdd.n2646 vdd.n2643 10.6151
R21006 vdd.n2641 vdd.n2638 10.6151
R21007 vdd.n2638 vdd.n2637 10.6151
R21008 vdd.n2707 vdd.n2706 10.6151
R21009 vdd.n2707 vdd.n740 10.6151
R21010 vdd.n2717 vdd.n740 10.6151
R21011 vdd.n2718 vdd.n2717 10.6151
R21012 vdd.n2719 vdd.n2718 10.6151
R21013 vdd.n2719 vdd.n728 10.6151
R21014 vdd.n2729 vdd.n728 10.6151
R21015 vdd.n2730 vdd.n2729 10.6151
R21016 vdd.n2731 vdd.n2730 10.6151
R21017 vdd.n2731 vdd.n717 10.6151
R21018 vdd.n2741 vdd.n717 10.6151
R21019 vdd.n2742 vdd.n2741 10.6151
R21020 vdd.n2743 vdd.n2742 10.6151
R21021 vdd.n2743 vdd.n706 10.6151
R21022 vdd.n2753 vdd.n706 10.6151
R21023 vdd.n2754 vdd.n2753 10.6151
R21024 vdd.n2755 vdd.n2754 10.6151
R21025 vdd.n2755 vdd.n693 10.6151
R21026 vdd.n2766 vdd.n693 10.6151
R21027 vdd.n2767 vdd.n2766 10.6151
R21028 vdd.n2768 vdd.n2767 10.6151
R21029 vdd.n2768 vdd.n681 10.6151
R21030 vdd.n2778 vdd.n681 10.6151
R21031 vdd.n2779 vdd.n2778 10.6151
R21032 vdd.n2780 vdd.n2779 10.6151
R21033 vdd.n2780 vdd.n669 10.6151
R21034 vdd.n2790 vdd.n669 10.6151
R21035 vdd.n2791 vdd.n2790 10.6151
R21036 vdd.n2792 vdd.n2791 10.6151
R21037 vdd.n2792 vdd.n656 10.6151
R21038 vdd.n2802 vdd.n656 10.6151
R21039 vdd.n2803 vdd.n2802 10.6151
R21040 vdd.n2804 vdd.n2803 10.6151
R21041 vdd.n2804 vdd.n645 10.6151
R21042 vdd.n2814 vdd.n645 10.6151
R21043 vdd.n2815 vdd.n2814 10.6151
R21044 vdd.n2816 vdd.n2815 10.6151
R21045 vdd.n2816 vdd.n631 10.6151
R21046 vdd.n2871 vdd.n631 10.6151
R21047 vdd.n2872 vdd.n2871 10.6151
R21048 vdd.n2873 vdd.n2872 10.6151
R21049 vdd.n2873 vdd.n600 10.6151
R21050 vdd.n2943 vdd.n600 10.6151
R21051 vdd.n2942 vdd.n2941 10.6151
R21052 vdd.n2941 vdd.n601 10.6151
R21053 vdd.n602 vdd.n601 10.6151
R21054 vdd.n2934 vdd.n602 10.6151
R21055 vdd.n2934 vdd.n2933 10.6151
R21056 vdd.n2933 vdd.n2932 10.6151
R21057 vdd.n2932 vdd.n604 10.6151
R21058 vdd.n2927 vdd.n604 10.6151
R21059 vdd.n2927 vdd.n2926 10.6151
R21060 vdd.n2926 vdd.n2925 10.6151
R21061 vdd.n2925 vdd.n607 10.6151
R21062 vdd.n2920 vdd.n607 10.6151
R21063 vdd.n2920 vdd.n2919 10.6151
R21064 vdd.n2919 vdd.n2918 10.6151
R21065 vdd.n2918 vdd.n610 10.6151
R21066 vdd.n2913 vdd.n610 10.6151
R21067 vdd.n2913 vdd.n520 10.6151
R21068 vdd.n2909 vdd.n520 10.6151
R21069 vdd.n2909 vdd.n2908 10.6151
R21070 vdd.n2908 vdd.n2907 10.6151
R21071 vdd.n2907 vdd.n613 10.6151
R21072 vdd.n2902 vdd.n613 10.6151
R21073 vdd.n2902 vdd.n2901 10.6151
R21074 vdd.n2901 vdd.n2900 10.6151
R21075 vdd.n2900 vdd.n616 10.6151
R21076 vdd.n2895 vdd.n616 10.6151
R21077 vdd.n2895 vdd.n2894 10.6151
R21078 vdd.n2894 vdd.n2893 10.6151
R21079 vdd.n2893 vdd.n619 10.6151
R21080 vdd.n2888 vdd.n619 10.6151
R21081 vdd.n2888 vdd.n2887 10.6151
R21082 vdd.n2885 vdd.n624 10.6151
R21083 vdd.n2880 vdd.n624 10.6151
R21084 vdd.n2861 vdd.n2822 10.6151
R21085 vdd.n2856 vdd.n2822 10.6151
R21086 vdd.n2856 vdd.n2855 10.6151
R21087 vdd.n2855 vdd.n2854 10.6151
R21088 vdd.n2854 vdd.n2824 10.6151
R21089 vdd.n2849 vdd.n2824 10.6151
R21090 vdd.n2849 vdd.n2848 10.6151
R21091 vdd.n2848 vdd.n2847 10.6151
R21092 vdd.n2847 vdd.n2827 10.6151
R21093 vdd.n2842 vdd.n2827 10.6151
R21094 vdd.n2842 vdd.n2841 10.6151
R21095 vdd.n2841 vdd.n2840 10.6151
R21096 vdd.n2840 vdd.n2830 10.6151
R21097 vdd.n2835 vdd.n2830 10.6151
R21098 vdd.n2835 vdd.n2834 10.6151
R21099 vdd.n2834 vdd.n575 10.6151
R21100 vdd.n2978 vdd.n575 10.6151
R21101 vdd.n2978 vdd.n576 10.6151
R21102 vdd.n578 vdd.n576 10.6151
R21103 vdd.n2971 vdd.n578 10.6151
R21104 vdd.n2971 vdd.n2970 10.6151
R21105 vdd.n2970 vdd.n2969 10.6151
R21106 vdd.n2969 vdd.n580 10.6151
R21107 vdd.n2964 vdd.n580 10.6151
R21108 vdd.n2964 vdd.n2963 10.6151
R21109 vdd.n2963 vdd.n2962 10.6151
R21110 vdd.n2962 vdd.n583 10.6151
R21111 vdd.n2957 vdd.n583 10.6151
R21112 vdd.n2957 vdd.n2956 10.6151
R21113 vdd.n2956 vdd.n2955 10.6151
R21114 vdd.n2955 vdd.n586 10.6151
R21115 vdd.n2950 vdd.n2949 10.6151
R21116 vdd.n2949 vdd.n2948 10.6151
R21117 vdd.n2511 vdd.n2510 10.6151
R21118 vdd.n2628 vdd.n2511 10.6151
R21119 vdd.n2628 vdd.n2627 10.6151
R21120 vdd.n2627 vdd.n2626 10.6151
R21121 vdd.n2626 vdd.n2624 10.6151
R21122 vdd.n2624 vdd.n2623 10.6151
R21123 vdd.n2623 vdd.n2621 10.6151
R21124 vdd.n2621 vdd.n2620 10.6151
R21125 vdd.n2620 vdd.n2512 10.6151
R21126 vdd.n2610 vdd.n2512 10.6151
R21127 vdd.n2610 vdd.n2609 10.6151
R21128 vdd.n2609 vdd.n2608 10.6151
R21129 vdd.n2608 vdd.n2606 10.6151
R21130 vdd.n2606 vdd.n2605 10.6151
R21131 vdd.n2605 vdd.n2603 10.6151
R21132 vdd.n2603 vdd.n2602 10.6151
R21133 vdd.n2602 vdd.n2600 10.6151
R21134 vdd.n2600 vdd.n2599 10.6151
R21135 vdd.n2599 vdd.n2597 10.6151
R21136 vdd.n2597 vdd.n2596 10.6151
R21137 vdd.n2596 vdd.n2594 10.6151
R21138 vdd.n2594 vdd.n2593 10.6151
R21139 vdd.n2593 vdd.n2591 10.6151
R21140 vdd.n2591 vdd.n2590 10.6151
R21141 vdd.n2590 vdd.n2588 10.6151
R21142 vdd.n2588 vdd.n2587 10.6151
R21143 vdd.n2587 vdd.n2585 10.6151
R21144 vdd.n2585 vdd.n2584 10.6151
R21145 vdd.n2584 vdd.n2582 10.6151
R21146 vdd.n2582 vdd.n2581 10.6151
R21147 vdd.n2581 vdd.n2579 10.6151
R21148 vdd.n2579 vdd.n2578 10.6151
R21149 vdd.n2578 vdd.n2576 10.6151
R21150 vdd.n2576 vdd.n2575 10.6151
R21151 vdd.n2575 vdd.n2573 10.6151
R21152 vdd.n2573 vdd.n2572 10.6151
R21153 vdd.n2572 vdd.n2570 10.6151
R21154 vdd.n2570 vdd.n2569 10.6151
R21155 vdd.n2569 vdd.n2567 10.6151
R21156 vdd.n2567 vdd.n2566 10.6151
R21157 vdd.n2566 vdd.n2564 10.6151
R21158 vdd.n2564 vdd.n2563 10.6151
R21159 vdd.n2563 vdd.n592 10.6151
R21160 vdd.n2442 vdd.n2441 10.6151
R21161 vdd.n2445 vdd.n2442 10.6151
R21162 vdd.n2446 vdd.n2445 10.6151
R21163 vdd.n2449 vdd.n2446 10.6151
R21164 vdd.n2450 vdd.n2449 10.6151
R21165 vdd.n2453 vdd.n2450 10.6151
R21166 vdd.n2454 vdd.n2453 10.6151
R21167 vdd.n2457 vdd.n2454 10.6151
R21168 vdd.n2458 vdd.n2457 10.6151
R21169 vdd.n2461 vdd.n2458 10.6151
R21170 vdd.n2462 vdd.n2461 10.6151
R21171 vdd.n2465 vdd.n2462 10.6151
R21172 vdd.n2466 vdd.n2465 10.6151
R21173 vdd.n2469 vdd.n2466 10.6151
R21174 vdd.n2470 vdd.n2469 10.6151
R21175 vdd.n2473 vdd.n2470 10.6151
R21176 vdd.n2474 vdd.n2473 10.6151
R21177 vdd.n2477 vdd.n2474 10.6151
R21178 vdd.n2478 vdd.n2477 10.6151
R21179 vdd.n2481 vdd.n2478 10.6151
R21180 vdd.n2482 vdd.n2481 10.6151
R21181 vdd.n2485 vdd.n2482 10.6151
R21182 vdd.n2486 vdd.n2485 10.6151
R21183 vdd.n2489 vdd.n2486 10.6151
R21184 vdd.n2490 vdd.n2489 10.6151
R21185 vdd.n2493 vdd.n2490 10.6151
R21186 vdd.n2494 vdd.n2493 10.6151
R21187 vdd.n2497 vdd.n2494 10.6151
R21188 vdd.n2498 vdd.n2497 10.6151
R21189 vdd.n2501 vdd.n2498 10.6151
R21190 vdd.n2502 vdd.n2501 10.6151
R21191 vdd.n2507 vdd.n2505 10.6151
R21192 vdd.n2508 vdd.n2507 10.6151
R21193 vdd.n2711 vdd.n745 10.6151
R21194 vdd.n2712 vdd.n2711 10.6151
R21195 vdd.n2713 vdd.n2712 10.6151
R21196 vdd.n2713 vdd.n734 10.6151
R21197 vdd.n2723 vdd.n734 10.6151
R21198 vdd.n2724 vdd.n2723 10.6151
R21199 vdd.n2725 vdd.n2724 10.6151
R21200 vdd.n2725 vdd.n723 10.6151
R21201 vdd.n2735 vdd.n723 10.6151
R21202 vdd.n2736 vdd.n2735 10.6151
R21203 vdd.n2737 vdd.n2736 10.6151
R21204 vdd.n2737 vdd.n711 10.6151
R21205 vdd.n2747 vdd.n711 10.6151
R21206 vdd.n2748 vdd.n2747 10.6151
R21207 vdd.n2749 vdd.n2748 10.6151
R21208 vdd.n2749 vdd.n700 10.6151
R21209 vdd.n2759 vdd.n700 10.6151
R21210 vdd.n2760 vdd.n2759 10.6151
R21211 vdd.n2762 vdd.n2760 10.6151
R21212 vdd.n2762 vdd.n2761 10.6151
R21213 vdd.n2773 vdd.n2772 10.6151
R21214 vdd.n2774 vdd.n2773 10.6151
R21215 vdd.n2774 vdd.n675 10.6151
R21216 vdd.n2784 vdd.n675 10.6151
R21217 vdd.n2785 vdd.n2784 10.6151
R21218 vdd.n2786 vdd.n2785 10.6151
R21219 vdd.n2786 vdd.n662 10.6151
R21220 vdd.n2796 vdd.n662 10.6151
R21221 vdd.n2797 vdd.n2796 10.6151
R21222 vdd.n2798 vdd.n2797 10.6151
R21223 vdd.n2798 vdd.n650 10.6151
R21224 vdd.n2808 vdd.n650 10.6151
R21225 vdd.n2809 vdd.n2808 10.6151
R21226 vdd.n2810 vdd.n2809 10.6151
R21227 vdd.n2810 vdd.n639 10.6151
R21228 vdd.n2820 vdd.n639 10.6151
R21229 vdd.n2821 vdd.n2820 10.6151
R21230 vdd.n2867 vdd.n2821 10.6151
R21231 vdd.n2867 vdd.n2866 10.6151
R21232 vdd.n2866 vdd.n2865 10.6151
R21233 vdd.n2865 vdd.n2864 10.6151
R21234 vdd.n2864 vdd.n2862 10.6151
R21235 vdd.n2129 vdd.n922 10.6151
R21236 vdd.n2130 vdd.n2129 10.6151
R21237 vdd.n2131 vdd.n2130 10.6151
R21238 vdd.n2131 vdd.n911 10.6151
R21239 vdd.n2141 vdd.n911 10.6151
R21240 vdd.n2142 vdd.n2141 10.6151
R21241 vdd.n2143 vdd.n2142 10.6151
R21242 vdd.n2143 vdd.n898 10.6151
R21243 vdd.n2153 vdd.n898 10.6151
R21244 vdd.n2154 vdd.n2153 10.6151
R21245 vdd.n2155 vdd.n2154 10.6151
R21246 vdd.n2155 vdd.n887 10.6151
R21247 vdd.n2165 vdd.n887 10.6151
R21248 vdd.n2166 vdd.n2165 10.6151
R21249 vdd.n2167 vdd.n2166 10.6151
R21250 vdd.n2167 vdd.n875 10.6151
R21251 vdd.n2177 vdd.n875 10.6151
R21252 vdd.n2178 vdd.n2177 10.6151
R21253 vdd.n2179 vdd.n2178 10.6151
R21254 vdd.n2179 vdd.n862 10.6151
R21255 vdd.n2189 vdd.n862 10.6151
R21256 vdd.n2190 vdd.n2189 10.6151
R21257 vdd.n2192 vdd.n850 10.6151
R21258 vdd.n2202 vdd.n850 10.6151
R21259 vdd.n2203 vdd.n2202 10.6151
R21260 vdd.n2204 vdd.n2203 10.6151
R21261 vdd.n2204 vdd.n838 10.6151
R21262 vdd.n2214 vdd.n838 10.6151
R21263 vdd.n2215 vdd.n2214 10.6151
R21264 vdd.n2216 vdd.n2215 10.6151
R21265 vdd.n2216 vdd.n827 10.6151
R21266 vdd.n2226 vdd.n827 10.6151
R21267 vdd.n2227 vdd.n2226 10.6151
R21268 vdd.n2228 vdd.n2227 10.6151
R21269 vdd.n2228 vdd.n816 10.6151
R21270 vdd.n2238 vdd.n816 10.6151
R21271 vdd.n2239 vdd.n2238 10.6151
R21272 vdd.n2242 vdd.n2239 10.6151
R21273 vdd.n2242 vdd.n2241 10.6151
R21274 vdd.n2241 vdd.n2240 10.6151
R21275 vdd.n2240 vdd.n799 10.6151
R21276 vdd.n2324 vdd.n799 10.6151
R21277 vdd.n2323 vdd.n2322 10.6151
R21278 vdd.n2322 vdd.n2319 10.6151
R21279 vdd.n2319 vdd.n2318 10.6151
R21280 vdd.n2318 vdd.n2315 10.6151
R21281 vdd.n2315 vdd.n2314 10.6151
R21282 vdd.n2314 vdd.n2311 10.6151
R21283 vdd.n2311 vdd.n2310 10.6151
R21284 vdd.n2310 vdd.n2307 10.6151
R21285 vdd.n2307 vdd.n2306 10.6151
R21286 vdd.n2306 vdd.n2303 10.6151
R21287 vdd.n2303 vdd.n2302 10.6151
R21288 vdd.n2302 vdd.n2299 10.6151
R21289 vdd.n2299 vdd.n2298 10.6151
R21290 vdd.n2298 vdd.n2295 10.6151
R21291 vdd.n2295 vdd.n2294 10.6151
R21292 vdd.n2294 vdd.n2291 10.6151
R21293 vdd.n2291 vdd.n2290 10.6151
R21294 vdd.n2290 vdd.n2287 10.6151
R21295 vdd.n2287 vdd.n2286 10.6151
R21296 vdd.n2286 vdd.n2283 10.6151
R21297 vdd.n2283 vdd.n2282 10.6151
R21298 vdd.n2282 vdd.n2279 10.6151
R21299 vdd.n2279 vdd.n2278 10.6151
R21300 vdd.n2278 vdd.n2275 10.6151
R21301 vdd.n2275 vdd.n2274 10.6151
R21302 vdd.n2274 vdd.n2271 10.6151
R21303 vdd.n2271 vdd.n2270 10.6151
R21304 vdd.n2270 vdd.n2267 10.6151
R21305 vdd.n2267 vdd.n2266 10.6151
R21306 vdd.n2266 vdd.n2263 10.6151
R21307 vdd.n2263 vdd.n2262 10.6151
R21308 vdd.n2259 vdd.n2258 10.6151
R21309 vdd.n2258 vdd.n2256 10.6151
R21310 vdd.n1271 vdd.n1269 10.6151
R21311 vdd.n1269 vdd.n1268 10.6151
R21312 vdd.n1268 vdd.n1266 10.6151
R21313 vdd.n1266 vdd.n1265 10.6151
R21314 vdd.n1265 vdd.n1263 10.6151
R21315 vdd.n1263 vdd.n1262 10.6151
R21316 vdd.n1262 vdd.n1260 10.6151
R21317 vdd.n1260 vdd.n1259 10.6151
R21318 vdd.n1259 vdd.n1257 10.6151
R21319 vdd.n1257 vdd.n1256 10.6151
R21320 vdd.n1256 vdd.n1254 10.6151
R21321 vdd.n1254 vdd.n1253 10.6151
R21322 vdd.n1253 vdd.n1251 10.6151
R21323 vdd.n1251 vdd.n1250 10.6151
R21324 vdd.n1250 vdd.n1248 10.6151
R21325 vdd.n1248 vdd.n1247 10.6151
R21326 vdd.n1247 vdd.n1245 10.6151
R21327 vdd.n1245 vdd.n1244 10.6151
R21328 vdd.n1244 vdd.n1242 10.6151
R21329 vdd.n1242 vdd.n1241 10.6151
R21330 vdd.n1241 vdd.n1239 10.6151
R21331 vdd.n1239 vdd.n1238 10.6151
R21332 vdd.n1238 vdd.n1236 10.6151
R21333 vdd.n1236 vdd.n1235 10.6151
R21334 vdd.n1235 vdd.n1233 10.6151
R21335 vdd.n1233 vdd.n1232 10.6151
R21336 vdd.n1232 vdd.n1230 10.6151
R21337 vdd.n1230 vdd.n1229 10.6151
R21338 vdd.n1229 vdd.n1108 10.6151
R21339 vdd.n1200 vdd.n1108 10.6151
R21340 vdd.n1201 vdd.n1200 10.6151
R21341 vdd.n1203 vdd.n1201 10.6151
R21342 vdd.n1204 vdd.n1203 10.6151
R21343 vdd.n1213 vdd.n1204 10.6151
R21344 vdd.n1213 vdd.n1212 10.6151
R21345 vdd.n1212 vdd.n1211 10.6151
R21346 vdd.n1211 vdd.n1209 10.6151
R21347 vdd.n1209 vdd.n1208 10.6151
R21348 vdd.n1208 vdd.n1206 10.6151
R21349 vdd.n1206 vdd.n1205 10.6151
R21350 vdd.n1205 vdd.n803 10.6151
R21351 vdd.n2254 vdd.n803 10.6151
R21352 vdd.n2255 vdd.n2254 10.6151
R21353 vdd.n1072 vdd.n1071 10.6151
R21354 vdd.n1075 vdd.n1072 10.6151
R21355 vdd.n1076 vdd.n1075 10.6151
R21356 vdd.n1079 vdd.n1076 10.6151
R21357 vdd.n1080 vdd.n1079 10.6151
R21358 vdd.n1083 vdd.n1080 10.6151
R21359 vdd.n1084 vdd.n1083 10.6151
R21360 vdd.n1087 vdd.n1084 10.6151
R21361 vdd.n1088 vdd.n1087 10.6151
R21362 vdd.n1091 vdd.n1088 10.6151
R21363 vdd.n1092 vdd.n1091 10.6151
R21364 vdd.n1095 vdd.n1092 10.6151
R21365 vdd.n1096 vdd.n1095 10.6151
R21366 vdd.n1099 vdd.n1096 10.6151
R21367 vdd.n1100 vdd.n1099 10.6151
R21368 vdd.n1103 vdd.n1100 10.6151
R21369 vdd.n1305 vdd.n1103 10.6151
R21370 vdd.n1305 vdd.n1304 10.6151
R21371 vdd.n1304 vdd.n1302 10.6151
R21372 vdd.n1302 vdd.n1299 10.6151
R21373 vdd.n1299 vdd.n1298 10.6151
R21374 vdd.n1298 vdd.n1295 10.6151
R21375 vdd.n1295 vdd.n1294 10.6151
R21376 vdd.n1294 vdd.n1291 10.6151
R21377 vdd.n1291 vdd.n1290 10.6151
R21378 vdd.n1290 vdd.n1287 10.6151
R21379 vdd.n1287 vdd.n1286 10.6151
R21380 vdd.n1286 vdd.n1283 10.6151
R21381 vdd.n1283 vdd.n1282 10.6151
R21382 vdd.n1282 vdd.n1279 10.6151
R21383 vdd.n1279 vdd.n1278 10.6151
R21384 vdd.n1275 vdd.n1274 10.6151
R21385 vdd.n1274 vdd.n1272 10.6151
R21386 vdd.n280 vdd.n262 10.4732
R21387 vdd.n233 vdd.n215 10.4732
R21388 vdd.n190 vdd.n172 10.4732
R21389 vdd.n143 vdd.n125 10.4732
R21390 vdd.n101 vdd.n83 10.4732
R21391 vdd.n54 vdd.n36 10.4732
R21392 vdd.n1550 vdd.n1532 10.4732
R21393 vdd.n1597 vdd.n1579 10.4732
R21394 vdd.n1460 vdd.n1442 10.4732
R21395 vdd.n1507 vdd.n1489 10.4732
R21396 vdd.n1371 vdd.n1353 10.4732
R21397 vdd.n1418 vdd.n1400 10.4732
R21398 vdd.t132 vdd.n1343 10.3167
R21399 vdd.n3146 vdd.t100 10.3167
R21400 vdd.n1920 vdd.t112 10.09
R21401 vdd.n3314 vdd.t98 10.09
R21402 vdd.n2089 vdd.n2088 9.98956
R21403 vdd.n3108 vdd.n520 9.98956
R21404 vdd.n2979 vdd.n2978 9.98956
R21405 vdd.n1981 vdd.n1305 9.98956
R21406 vdd.n2326 vdd.t204 9.7499
R21407 vdd.t189 vdd.n747 9.7499
R21408 vdd.n279 vdd.n264 9.69747
R21409 vdd.n232 vdd.n217 9.69747
R21410 vdd.n189 vdd.n174 9.69747
R21411 vdd.n142 vdd.n127 9.69747
R21412 vdd.n100 vdd.n85 9.69747
R21413 vdd.n53 vdd.n38 9.69747
R21414 vdd.n1549 vdd.n1534 9.69747
R21415 vdd.n1596 vdd.n1581 9.69747
R21416 vdd.n1459 vdd.n1444 9.69747
R21417 vdd.n1506 vdd.n1491 9.69747
R21418 vdd.n1370 vdd.n1355 9.69747
R21419 vdd.n1417 vdd.n1402 9.69747
R21420 vdd.n295 vdd.n294 9.45567
R21421 vdd.n248 vdd.n247 9.45567
R21422 vdd.n205 vdd.n204 9.45567
R21423 vdd.n158 vdd.n157 9.45567
R21424 vdd.n116 vdd.n115 9.45567
R21425 vdd.n69 vdd.n68 9.45567
R21426 vdd.n1565 vdd.n1564 9.45567
R21427 vdd.n1612 vdd.n1611 9.45567
R21428 vdd.n1475 vdd.n1474 9.45567
R21429 vdd.n1522 vdd.n1521 9.45567
R21430 vdd.n1386 vdd.n1385 9.45567
R21431 vdd.n1433 vdd.n1432 9.45567
R21432 vdd.n2051 vdd.n997 9.3005
R21433 vdd.n2050 vdd.n2049 9.3005
R21434 vdd.n1003 vdd.n1002 9.3005
R21435 vdd.n2044 vdd.n1007 9.3005
R21436 vdd.n2043 vdd.n1008 9.3005
R21437 vdd.n2042 vdd.n1009 9.3005
R21438 vdd.n1013 vdd.n1010 9.3005
R21439 vdd.n2037 vdd.n1014 9.3005
R21440 vdd.n2036 vdd.n1015 9.3005
R21441 vdd.n2035 vdd.n1016 9.3005
R21442 vdd.n1020 vdd.n1017 9.3005
R21443 vdd.n2030 vdd.n1021 9.3005
R21444 vdd.n2029 vdd.n1022 9.3005
R21445 vdd.n2028 vdd.n1023 9.3005
R21446 vdd.n1027 vdd.n1024 9.3005
R21447 vdd.n2023 vdd.n1028 9.3005
R21448 vdd.n2022 vdd.n1029 9.3005
R21449 vdd.n2021 vdd.n1030 9.3005
R21450 vdd.n1034 vdd.n1031 9.3005
R21451 vdd.n2016 vdd.n1035 9.3005
R21452 vdd.n2015 vdd.n1036 9.3005
R21453 vdd.n2014 vdd.n2013 9.3005
R21454 vdd.n2012 vdd.n1037 9.3005
R21455 vdd.n2011 vdd.n2010 9.3005
R21456 vdd.n1043 vdd.n1042 9.3005
R21457 vdd.n2005 vdd.n1047 9.3005
R21458 vdd.n2004 vdd.n1048 9.3005
R21459 vdd.n2003 vdd.n1049 9.3005
R21460 vdd.n1053 vdd.n1050 9.3005
R21461 vdd.n1998 vdd.n1054 9.3005
R21462 vdd.n1997 vdd.n1055 9.3005
R21463 vdd.n1996 vdd.n1056 9.3005
R21464 vdd.n1060 vdd.n1057 9.3005
R21465 vdd.n1991 vdd.n1061 9.3005
R21466 vdd.n1990 vdd.n1062 9.3005
R21467 vdd.n1989 vdd.n1063 9.3005
R21468 vdd.n1067 vdd.n1064 9.3005
R21469 vdd.n1984 vdd.n1068 9.3005
R21470 vdd.n2053 vdd.n2052 9.3005
R21471 vdd.n2075 vdd.n968 9.3005
R21472 vdd.n2074 vdd.n976 9.3005
R21473 vdd.n980 vdd.n977 9.3005
R21474 vdd.n2069 vdd.n981 9.3005
R21475 vdd.n2068 vdd.n982 9.3005
R21476 vdd.n2067 vdd.n983 9.3005
R21477 vdd.n987 vdd.n984 9.3005
R21478 vdd.n2062 vdd.n988 9.3005
R21479 vdd.n2061 vdd.n989 9.3005
R21480 vdd.n2060 vdd.n990 9.3005
R21481 vdd.n994 vdd.n991 9.3005
R21482 vdd.n2055 vdd.n995 9.3005
R21483 vdd.n2054 vdd.n996 9.3005
R21484 vdd.n2087 vdd.n2086 9.3005
R21485 vdd.n972 vdd.n971 9.3005
R21486 vdd.n1931 vdd.n1930 9.3005
R21487 vdd.n1932 vdd.n1345 9.3005
R21488 vdd.n1934 vdd.n1933 9.3005
R21489 vdd.n1335 vdd.n1334 9.3005
R21490 vdd.n1948 vdd.n1947 9.3005
R21491 vdd.n1949 vdd.n1333 9.3005
R21492 vdd.n1951 vdd.n1950 9.3005
R21493 vdd.n1323 vdd.n1322 9.3005
R21494 vdd.n1967 vdd.n1966 9.3005
R21495 vdd.n1968 vdd.n1321 9.3005
R21496 vdd.n1970 vdd.n1969 9.3005
R21497 vdd.n271 vdd.n270 9.3005
R21498 vdd.n266 vdd.n265 9.3005
R21499 vdd.n277 vdd.n276 9.3005
R21500 vdd.n279 vdd.n278 9.3005
R21501 vdd.n262 vdd.n261 9.3005
R21502 vdd.n285 vdd.n284 9.3005
R21503 vdd.n287 vdd.n286 9.3005
R21504 vdd.n259 vdd.n256 9.3005
R21505 vdd.n294 vdd.n293 9.3005
R21506 vdd.n224 vdd.n223 9.3005
R21507 vdd.n219 vdd.n218 9.3005
R21508 vdd.n230 vdd.n229 9.3005
R21509 vdd.n232 vdd.n231 9.3005
R21510 vdd.n215 vdd.n214 9.3005
R21511 vdd.n238 vdd.n237 9.3005
R21512 vdd.n240 vdd.n239 9.3005
R21513 vdd.n212 vdd.n209 9.3005
R21514 vdd.n247 vdd.n246 9.3005
R21515 vdd.n181 vdd.n180 9.3005
R21516 vdd.n176 vdd.n175 9.3005
R21517 vdd.n187 vdd.n186 9.3005
R21518 vdd.n189 vdd.n188 9.3005
R21519 vdd.n172 vdd.n171 9.3005
R21520 vdd.n195 vdd.n194 9.3005
R21521 vdd.n197 vdd.n196 9.3005
R21522 vdd.n169 vdd.n166 9.3005
R21523 vdd.n204 vdd.n203 9.3005
R21524 vdd.n134 vdd.n133 9.3005
R21525 vdd.n129 vdd.n128 9.3005
R21526 vdd.n140 vdd.n139 9.3005
R21527 vdd.n142 vdd.n141 9.3005
R21528 vdd.n125 vdd.n124 9.3005
R21529 vdd.n148 vdd.n147 9.3005
R21530 vdd.n150 vdd.n149 9.3005
R21531 vdd.n122 vdd.n119 9.3005
R21532 vdd.n157 vdd.n156 9.3005
R21533 vdd.n92 vdd.n91 9.3005
R21534 vdd.n87 vdd.n86 9.3005
R21535 vdd.n98 vdd.n97 9.3005
R21536 vdd.n100 vdd.n99 9.3005
R21537 vdd.n83 vdd.n82 9.3005
R21538 vdd.n106 vdd.n105 9.3005
R21539 vdd.n108 vdd.n107 9.3005
R21540 vdd.n80 vdd.n77 9.3005
R21541 vdd.n115 vdd.n114 9.3005
R21542 vdd.n45 vdd.n44 9.3005
R21543 vdd.n40 vdd.n39 9.3005
R21544 vdd.n51 vdd.n50 9.3005
R21545 vdd.n53 vdd.n52 9.3005
R21546 vdd.n36 vdd.n35 9.3005
R21547 vdd.n59 vdd.n58 9.3005
R21548 vdd.n61 vdd.n60 9.3005
R21549 vdd.n33 vdd.n30 9.3005
R21550 vdd.n68 vdd.n67 9.3005
R21551 vdd.n3030 vdd.n3029 9.3005
R21552 vdd.n3033 vdd.n555 9.3005
R21553 vdd.n3034 vdd.n554 9.3005
R21554 vdd.n3037 vdd.n553 9.3005
R21555 vdd.n3038 vdd.n552 9.3005
R21556 vdd.n3041 vdd.n551 9.3005
R21557 vdd.n3042 vdd.n550 9.3005
R21558 vdd.n3045 vdd.n549 9.3005
R21559 vdd.n3046 vdd.n548 9.3005
R21560 vdd.n3049 vdd.n547 9.3005
R21561 vdd.n3050 vdd.n546 9.3005
R21562 vdd.n3053 vdd.n545 9.3005
R21563 vdd.n3054 vdd.n544 9.3005
R21564 vdd.n3057 vdd.n543 9.3005
R21565 vdd.n3058 vdd.n542 9.3005
R21566 vdd.n3061 vdd.n541 9.3005
R21567 vdd.n3062 vdd.n540 9.3005
R21568 vdd.n3065 vdd.n539 9.3005
R21569 vdd.n3066 vdd.n538 9.3005
R21570 vdd.n3069 vdd.n537 9.3005
R21571 vdd.n3073 vdd.n3072 9.3005
R21572 vdd.n3074 vdd.n536 9.3005
R21573 vdd.n3078 vdd.n3075 9.3005
R21574 vdd.n3081 vdd.n535 9.3005
R21575 vdd.n3082 vdd.n534 9.3005
R21576 vdd.n3085 vdd.n533 9.3005
R21577 vdd.n3086 vdd.n532 9.3005
R21578 vdd.n3089 vdd.n531 9.3005
R21579 vdd.n3090 vdd.n530 9.3005
R21580 vdd.n3093 vdd.n529 9.3005
R21581 vdd.n3094 vdd.n528 9.3005
R21582 vdd.n3097 vdd.n527 9.3005
R21583 vdd.n3098 vdd.n526 9.3005
R21584 vdd.n3101 vdd.n525 9.3005
R21585 vdd.n3102 vdd.n524 9.3005
R21586 vdd.n3105 vdd.n519 9.3005
R21587 vdd.n482 vdd.n481 9.3005
R21588 vdd.n3116 vdd.n3115 9.3005
R21589 vdd.n3119 vdd.n3118 9.3005
R21590 vdd.n471 vdd.n470 9.3005
R21591 vdd.n3133 vdd.n3132 9.3005
R21592 vdd.n3134 vdd.n469 9.3005
R21593 vdd.n3136 vdd.n3135 9.3005
R21594 vdd.n460 vdd.n459 9.3005
R21595 vdd.n3149 vdd.n3148 9.3005
R21596 vdd.n3150 vdd.n458 9.3005
R21597 vdd.n3152 vdd.n3151 9.3005
R21598 vdd.n300 vdd.n298 9.3005
R21599 vdd.n3117 vdd.n480 9.3005
R21600 vdd.n3318 vdd.n3317 9.3005
R21601 vdd.n301 vdd.n299 9.3005
R21602 vdd.n3311 vdd.n310 9.3005
R21603 vdd.n3310 vdd.n311 9.3005
R21604 vdd.n3309 vdd.n312 9.3005
R21605 vdd.n320 vdd.n313 9.3005
R21606 vdd.n3303 vdd.n321 9.3005
R21607 vdd.n3302 vdd.n322 9.3005
R21608 vdd.n3301 vdd.n323 9.3005
R21609 vdd.n331 vdd.n324 9.3005
R21610 vdd.n3295 vdd.n3294 9.3005
R21611 vdd.n3291 vdd.n332 9.3005
R21612 vdd.n3290 vdd.n335 9.3005
R21613 vdd.n339 vdd.n336 9.3005
R21614 vdd.n340 vdd.n337 9.3005
R21615 vdd.n3283 vdd.n341 9.3005
R21616 vdd.n3282 vdd.n342 9.3005
R21617 vdd.n3281 vdd.n343 9.3005
R21618 vdd.n347 vdd.n344 9.3005
R21619 vdd.n3276 vdd.n348 9.3005
R21620 vdd.n3275 vdd.n349 9.3005
R21621 vdd.n3274 vdd.n350 9.3005
R21622 vdd.n354 vdd.n351 9.3005
R21623 vdd.n3269 vdd.n355 9.3005
R21624 vdd.n3268 vdd.n356 9.3005
R21625 vdd.n3267 vdd.n357 9.3005
R21626 vdd.n361 vdd.n358 9.3005
R21627 vdd.n3262 vdd.n362 9.3005
R21628 vdd.n3261 vdd.n363 9.3005
R21629 vdd.n3260 vdd.n3259 9.3005
R21630 vdd.n3258 vdd.n364 9.3005
R21631 vdd.n3257 vdd.n3256 9.3005
R21632 vdd.n370 vdd.n369 9.3005
R21633 vdd.n3251 vdd.n374 9.3005
R21634 vdd.n3250 vdd.n375 9.3005
R21635 vdd.n3249 vdd.n376 9.3005
R21636 vdd.n380 vdd.n377 9.3005
R21637 vdd.n3244 vdd.n381 9.3005
R21638 vdd.n3243 vdd.n382 9.3005
R21639 vdd.n3242 vdd.n383 9.3005
R21640 vdd.n387 vdd.n384 9.3005
R21641 vdd.n3237 vdd.n388 9.3005
R21642 vdd.n3236 vdd.n389 9.3005
R21643 vdd.n3235 vdd.n390 9.3005
R21644 vdd.n394 vdd.n391 9.3005
R21645 vdd.n3230 vdd.n395 9.3005
R21646 vdd.n3229 vdd.n396 9.3005
R21647 vdd.n3228 vdd.n397 9.3005
R21648 vdd.n401 vdd.n398 9.3005
R21649 vdd.n3223 vdd.n402 9.3005
R21650 vdd.n3222 vdd.n403 9.3005
R21651 vdd.n3221 vdd.n3220 9.3005
R21652 vdd.n3219 vdd.n404 9.3005
R21653 vdd.n3218 vdd.n3217 9.3005
R21654 vdd.n410 vdd.n409 9.3005
R21655 vdd.n3212 vdd.n414 9.3005
R21656 vdd.n3211 vdd.n415 9.3005
R21657 vdd.n3210 vdd.n416 9.3005
R21658 vdd.n420 vdd.n417 9.3005
R21659 vdd.n3205 vdd.n421 9.3005
R21660 vdd.n3204 vdd.n422 9.3005
R21661 vdd.n3203 vdd.n423 9.3005
R21662 vdd.n427 vdd.n424 9.3005
R21663 vdd.n3198 vdd.n428 9.3005
R21664 vdd.n3197 vdd.n429 9.3005
R21665 vdd.n3196 vdd.n430 9.3005
R21666 vdd.n434 vdd.n431 9.3005
R21667 vdd.n3191 vdd.n435 9.3005
R21668 vdd.n3190 vdd.n436 9.3005
R21669 vdd.n3189 vdd.n437 9.3005
R21670 vdd.n441 vdd.n438 9.3005
R21671 vdd.n3184 vdd.n442 9.3005
R21672 vdd.n3183 vdd.n443 9.3005
R21673 vdd.n3179 vdd.n3176 9.3005
R21674 vdd.n3293 vdd.n3292 9.3005
R21675 vdd.n3124 vdd.n3123 9.3005
R21676 vdd.n3125 vdd.n475 9.3005
R21677 vdd.n3127 vdd.n3126 9.3005
R21678 vdd.n465 vdd.n464 9.3005
R21679 vdd.n3141 vdd.n3140 9.3005
R21680 vdd.n3142 vdd.n463 9.3005
R21681 vdd.n3144 vdd.n3143 9.3005
R21682 vdd.n453 vdd.n452 9.3005
R21683 vdd.n3157 vdd.n3156 9.3005
R21684 vdd.n3158 vdd.n451 9.3005
R21685 vdd.n3160 vdd.n3159 9.3005
R21686 vdd.n3161 vdd.n450 9.3005
R21687 vdd.n3163 vdd.n3162 9.3005
R21688 vdd.n3164 vdd.n449 9.3005
R21689 vdd.n3166 vdd.n3165 9.3005
R21690 vdd.n3167 vdd.n447 9.3005
R21691 vdd.n3169 vdd.n3168 9.3005
R21692 vdd.n3170 vdd.n446 9.3005
R21693 vdd.n3172 vdd.n3171 9.3005
R21694 vdd.n3173 vdd.n444 9.3005
R21695 vdd.n3175 vdd.n3174 9.3005
R21696 vdd.n477 vdd.n476 9.3005
R21697 vdd.n2982 vdd.n2981 9.3005
R21698 vdd.n2987 vdd.n2980 9.3005
R21699 vdd.n2996 vdd.n572 9.3005
R21700 vdd.n2999 vdd.n571 9.3005
R21701 vdd.n3000 vdd.n570 9.3005
R21702 vdd.n3003 vdd.n569 9.3005
R21703 vdd.n3004 vdd.n568 9.3005
R21704 vdd.n3007 vdd.n567 9.3005
R21705 vdd.n3008 vdd.n566 9.3005
R21706 vdd.n3011 vdd.n565 9.3005
R21707 vdd.n3012 vdd.n564 9.3005
R21708 vdd.n3015 vdd.n563 9.3005
R21709 vdd.n3016 vdd.n562 9.3005
R21710 vdd.n3019 vdd.n561 9.3005
R21711 vdd.n3020 vdd.n560 9.3005
R21712 vdd.n3023 vdd.n559 9.3005
R21713 vdd.n3027 vdd.n3026 9.3005
R21714 vdd.n3028 vdd.n556 9.3005
R21715 vdd.n1980 vdd.n1979 9.3005
R21716 vdd.n1975 vdd.n1307 9.3005
R21717 vdd.n1888 vdd.n1887 9.3005
R21718 vdd.n1889 vdd.n1643 9.3005
R21719 vdd.n1891 vdd.n1890 9.3005
R21720 vdd.n1633 vdd.n1632 9.3005
R21721 vdd.n1905 vdd.n1904 9.3005
R21722 vdd.n1906 vdd.n1631 9.3005
R21723 vdd.n1908 vdd.n1907 9.3005
R21724 vdd.n1623 vdd.n1622 9.3005
R21725 vdd.n1923 vdd.n1922 9.3005
R21726 vdd.n1924 vdd.n1621 9.3005
R21727 vdd.n1926 vdd.n1925 9.3005
R21728 vdd.n1340 vdd.n1339 9.3005
R21729 vdd.n1939 vdd.n1938 9.3005
R21730 vdd.n1940 vdd.n1338 9.3005
R21731 vdd.n1942 vdd.n1941 9.3005
R21732 vdd.n1330 vdd.n1329 9.3005
R21733 vdd.n1956 vdd.n1955 9.3005
R21734 vdd.n1957 vdd.n1327 9.3005
R21735 vdd.n1961 vdd.n1960 9.3005
R21736 vdd.n1959 vdd.n1328 9.3005
R21737 vdd.n1958 vdd.n1318 9.3005
R21738 vdd.n1645 vdd.n1644 9.3005
R21739 vdd.n1781 vdd.n1780 9.3005
R21740 vdd.n1782 vdd.n1771 9.3005
R21741 vdd.n1784 vdd.n1783 9.3005
R21742 vdd.n1785 vdd.n1770 9.3005
R21743 vdd.n1787 vdd.n1786 9.3005
R21744 vdd.n1788 vdd.n1765 9.3005
R21745 vdd.n1790 vdd.n1789 9.3005
R21746 vdd.n1791 vdd.n1764 9.3005
R21747 vdd.n1793 vdd.n1792 9.3005
R21748 vdd.n1794 vdd.n1759 9.3005
R21749 vdd.n1796 vdd.n1795 9.3005
R21750 vdd.n1797 vdd.n1758 9.3005
R21751 vdd.n1799 vdd.n1798 9.3005
R21752 vdd.n1800 vdd.n1753 9.3005
R21753 vdd.n1802 vdd.n1801 9.3005
R21754 vdd.n1803 vdd.n1752 9.3005
R21755 vdd.n1805 vdd.n1804 9.3005
R21756 vdd.n1806 vdd.n1747 9.3005
R21757 vdd.n1808 vdd.n1807 9.3005
R21758 vdd.n1809 vdd.n1746 9.3005
R21759 vdd.n1811 vdd.n1810 9.3005
R21760 vdd.n1815 vdd.n1742 9.3005
R21761 vdd.n1817 vdd.n1816 9.3005
R21762 vdd.n1818 vdd.n1741 9.3005
R21763 vdd.n1820 vdd.n1819 9.3005
R21764 vdd.n1821 vdd.n1736 9.3005
R21765 vdd.n1823 vdd.n1822 9.3005
R21766 vdd.n1824 vdd.n1735 9.3005
R21767 vdd.n1826 vdd.n1825 9.3005
R21768 vdd.n1827 vdd.n1730 9.3005
R21769 vdd.n1829 vdd.n1828 9.3005
R21770 vdd.n1830 vdd.n1729 9.3005
R21771 vdd.n1832 vdd.n1831 9.3005
R21772 vdd.n1833 vdd.n1724 9.3005
R21773 vdd.n1835 vdd.n1834 9.3005
R21774 vdd.n1836 vdd.n1723 9.3005
R21775 vdd.n1838 vdd.n1837 9.3005
R21776 vdd.n1839 vdd.n1718 9.3005
R21777 vdd.n1841 vdd.n1840 9.3005
R21778 vdd.n1842 vdd.n1717 9.3005
R21779 vdd.n1844 vdd.n1843 9.3005
R21780 vdd.n1845 vdd.n1712 9.3005
R21781 vdd.n1847 vdd.n1846 9.3005
R21782 vdd.n1848 vdd.n1711 9.3005
R21783 vdd.n1850 vdd.n1849 9.3005
R21784 vdd.n1851 vdd.n1704 9.3005
R21785 vdd.n1853 vdd.n1852 9.3005
R21786 vdd.n1854 vdd.n1703 9.3005
R21787 vdd.n1856 vdd.n1855 9.3005
R21788 vdd.n1857 vdd.n1698 9.3005
R21789 vdd.n1859 vdd.n1858 9.3005
R21790 vdd.n1860 vdd.n1697 9.3005
R21791 vdd.n1862 vdd.n1861 9.3005
R21792 vdd.n1863 vdd.n1692 9.3005
R21793 vdd.n1865 vdd.n1864 9.3005
R21794 vdd.n1866 vdd.n1691 9.3005
R21795 vdd.n1868 vdd.n1867 9.3005
R21796 vdd.n1869 vdd.n1686 9.3005
R21797 vdd.n1871 vdd.n1870 9.3005
R21798 vdd.n1872 vdd.n1685 9.3005
R21799 vdd.n1874 vdd.n1873 9.3005
R21800 vdd.n1650 vdd.n1649 9.3005
R21801 vdd.n1880 vdd.n1879 9.3005
R21802 vdd.n1779 vdd.n1778 9.3005
R21803 vdd.n1883 vdd.n1882 9.3005
R21804 vdd.n1639 vdd.n1638 9.3005
R21805 vdd.n1897 vdd.n1896 9.3005
R21806 vdd.n1898 vdd.n1637 9.3005
R21807 vdd.n1900 vdd.n1899 9.3005
R21808 vdd.n1628 vdd.n1627 9.3005
R21809 vdd.n1914 vdd.n1913 9.3005
R21810 vdd.n1915 vdd.n1626 9.3005
R21811 vdd.n1918 vdd.n1917 9.3005
R21812 vdd.n1916 vdd.n1617 9.3005
R21813 vdd.n1881 vdd.n1648 9.3005
R21814 vdd.n1541 vdd.n1540 9.3005
R21815 vdd.n1536 vdd.n1535 9.3005
R21816 vdd.n1547 vdd.n1546 9.3005
R21817 vdd.n1549 vdd.n1548 9.3005
R21818 vdd.n1532 vdd.n1531 9.3005
R21819 vdd.n1555 vdd.n1554 9.3005
R21820 vdd.n1557 vdd.n1556 9.3005
R21821 vdd.n1529 vdd.n1526 9.3005
R21822 vdd.n1564 vdd.n1563 9.3005
R21823 vdd.n1588 vdd.n1587 9.3005
R21824 vdd.n1583 vdd.n1582 9.3005
R21825 vdd.n1594 vdd.n1593 9.3005
R21826 vdd.n1596 vdd.n1595 9.3005
R21827 vdd.n1579 vdd.n1578 9.3005
R21828 vdd.n1602 vdd.n1601 9.3005
R21829 vdd.n1604 vdd.n1603 9.3005
R21830 vdd.n1576 vdd.n1573 9.3005
R21831 vdd.n1611 vdd.n1610 9.3005
R21832 vdd.n1451 vdd.n1450 9.3005
R21833 vdd.n1446 vdd.n1445 9.3005
R21834 vdd.n1457 vdd.n1456 9.3005
R21835 vdd.n1459 vdd.n1458 9.3005
R21836 vdd.n1442 vdd.n1441 9.3005
R21837 vdd.n1465 vdd.n1464 9.3005
R21838 vdd.n1467 vdd.n1466 9.3005
R21839 vdd.n1439 vdd.n1436 9.3005
R21840 vdd.n1474 vdd.n1473 9.3005
R21841 vdd.n1498 vdd.n1497 9.3005
R21842 vdd.n1493 vdd.n1492 9.3005
R21843 vdd.n1504 vdd.n1503 9.3005
R21844 vdd.n1506 vdd.n1505 9.3005
R21845 vdd.n1489 vdd.n1488 9.3005
R21846 vdd.n1512 vdd.n1511 9.3005
R21847 vdd.n1514 vdd.n1513 9.3005
R21848 vdd.n1486 vdd.n1483 9.3005
R21849 vdd.n1521 vdd.n1520 9.3005
R21850 vdd.n1362 vdd.n1361 9.3005
R21851 vdd.n1357 vdd.n1356 9.3005
R21852 vdd.n1368 vdd.n1367 9.3005
R21853 vdd.n1370 vdd.n1369 9.3005
R21854 vdd.n1353 vdd.n1352 9.3005
R21855 vdd.n1376 vdd.n1375 9.3005
R21856 vdd.n1378 vdd.n1377 9.3005
R21857 vdd.n1350 vdd.n1347 9.3005
R21858 vdd.n1385 vdd.n1384 9.3005
R21859 vdd.n1409 vdd.n1408 9.3005
R21860 vdd.n1404 vdd.n1403 9.3005
R21861 vdd.n1415 vdd.n1414 9.3005
R21862 vdd.n1417 vdd.n1416 9.3005
R21863 vdd.n1400 vdd.n1399 9.3005
R21864 vdd.n1423 vdd.n1422 9.3005
R21865 vdd.n1425 vdd.n1424 9.3005
R21866 vdd.n1397 vdd.n1394 9.3005
R21867 vdd.n1432 vdd.n1431 9.3005
R21868 vdd.n1893 vdd.t94 8.95635
R21869 vdd.t121 vdd.n3305 8.95635
R21870 vdd.n276 vdd.n275 8.92171
R21871 vdd.n229 vdd.n228 8.92171
R21872 vdd.n186 vdd.n185 8.92171
R21873 vdd.n139 vdd.n138 8.92171
R21874 vdd.n97 vdd.n96 8.92171
R21875 vdd.n50 vdd.n49 8.92171
R21876 vdd.n1546 vdd.n1545 8.92171
R21877 vdd.n1593 vdd.n1592 8.92171
R21878 vdd.n1456 vdd.n1455 8.92171
R21879 vdd.n1503 vdd.n1502 8.92171
R21880 vdd.n1367 vdd.n1366 8.92171
R21881 vdd.n1414 vdd.n1413 8.92171
R21882 vdd.n207 vdd.n117 8.81535
R21883 vdd.n1524 vdd.n1434 8.81535
R21884 vdd.n1920 vdd.t110 8.72962
R21885 vdd.t139 vdd.n3314 8.72962
R21886 vdd.n1343 vdd.t130 8.50289
R21887 vdd.n1972 vdd.t25 8.50289
R21888 vdd.n516 vdd.t35 8.50289
R21889 vdd.n3146 vdd.t117 8.50289
R21890 vdd.n28 vdd.n14 8.42249
R21891 vdd.n3320 vdd.n3319 8.16225
R21892 vdd.n1616 vdd.n1615 8.16225
R21893 vdd.n272 vdd.n266 8.14595
R21894 vdd.n225 vdd.n219 8.14595
R21895 vdd.n182 vdd.n176 8.14595
R21896 vdd.n135 vdd.n129 8.14595
R21897 vdd.n93 vdd.n87 8.14595
R21898 vdd.n46 vdd.n40 8.14595
R21899 vdd.n1542 vdd.n1536 8.14595
R21900 vdd.n1589 vdd.n1583 8.14595
R21901 vdd.n1452 vdd.n1446 8.14595
R21902 vdd.n1499 vdd.n1493 8.14595
R21903 vdd.n1363 vdd.n1357 8.14595
R21904 vdd.n1410 vdd.n1404 8.14595
R21905 vdd.n2127 vdd.n924 7.70933
R21906 vdd.n2127 vdd.n927 7.70933
R21907 vdd.n2133 vdd.n913 7.70933
R21908 vdd.n2139 vdd.n913 7.70933
R21909 vdd.n2139 vdd.n906 7.70933
R21910 vdd.n2145 vdd.n906 7.70933
R21911 vdd.n2145 vdd.n909 7.70933
R21912 vdd.n2151 vdd.n902 7.70933
R21913 vdd.n2157 vdd.n896 7.70933
R21914 vdd.n2163 vdd.n883 7.70933
R21915 vdd.n2169 vdd.n883 7.70933
R21916 vdd.n2175 vdd.n877 7.70933
R21917 vdd.n2181 vdd.n870 7.70933
R21918 vdd.n2181 vdd.n873 7.70933
R21919 vdd.n2187 vdd.n866 7.70933
R21920 vdd.n2194 vdd.n852 7.70933
R21921 vdd.n2200 vdd.n852 7.70933
R21922 vdd.n2206 vdd.n846 7.70933
R21923 vdd.n2212 vdd.n842 7.70933
R21924 vdd.n2218 vdd.n836 7.70933
R21925 vdd.n2236 vdd.n818 7.70933
R21926 vdd.n2236 vdd.n811 7.70933
R21927 vdd.n2244 vdd.n811 7.70933
R21928 vdd.n2326 vdd.n795 7.70933
R21929 vdd.n2709 vdd.n747 7.70933
R21930 vdd.n2721 vdd.n736 7.70933
R21931 vdd.n2721 vdd.n730 7.70933
R21932 vdd.n2727 vdd.n730 7.70933
R21933 vdd.n2739 vdd.n721 7.70933
R21934 vdd.n2745 vdd.n715 7.70933
R21935 vdd.n2757 vdd.n702 7.70933
R21936 vdd.n2764 vdd.n695 7.70933
R21937 vdd.n2764 vdd.n698 7.70933
R21938 vdd.n2770 vdd.n691 7.70933
R21939 vdd.n2776 vdd.n677 7.70933
R21940 vdd.n2782 vdd.n677 7.70933
R21941 vdd.n2788 vdd.n671 7.70933
R21942 vdd.n2794 vdd.n664 7.70933
R21943 vdd.n2794 vdd.n667 7.70933
R21944 vdd.n2800 vdd.n660 7.70933
R21945 vdd.n2806 vdd.n654 7.70933
R21946 vdd.n2812 vdd.n641 7.70933
R21947 vdd.n2818 vdd.n641 7.70933
R21948 vdd.n2818 vdd.n633 7.70933
R21949 vdd.n2869 vdd.n633 7.70933
R21950 vdd.n2869 vdd.n636 7.70933
R21951 vdd.n2875 vdd.n595 7.70933
R21952 vdd.n2945 vdd.n595 7.70933
R21953 vdd.n271 vdd.n268 7.3702
R21954 vdd.n224 vdd.n221 7.3702
R21955 vdd.n181 vdd.n178 7.3702
R21956 vdd.n134 vdd.n131 7.3702
R21957 vdd.n92 vdd.n89 7.3702
R21958 vdd.n45 vdd.n42 7.3702
R21959 vdd.n1541 vdd.n1538 7.3702
R21960 vdd.n1588 vdd.n1585 7.3702
R21961 vdd.n1451 vdd.n1448 7.3702
R21962 vdd.n1498 vdd.n1495 7.3702
R21963 vdd.n1362 vdd.n1359 7.3702
R21964 vdd.n1409 vdd.n1406 7.3702
R21965 vdd.n896 vdd.t209 7.36923
R21966 vdd.n2800 vdd.t186 7.36923
R21967 vdd.n2151 vdd.t161 7.1425
R21968 vdd.n1215 vdd.t157 7.1425
R21969 vdd.n2733 vdd.t160 7.1425
R21970 vdd.n654 vdd.t174 7.1425
R21971 vdd.n1816 vdd.n1815 6.98232
R21972 vdd.n2015 vdd.n2014 6.98232
R21973 vdd.n3222 vdd.n3221 6.98232
R21974 vdd.n3033 vdd.n3030 6.98232
R21975 vdd.n1215 vdd.t158 6.80241
R21976 vdd.n2733 vdd.t202 6.80241
R21977 vdd.n1953 vdd.t114 6.68904
R21978 vdd.n3129 vdd.t126 6.68904
R21979 vdd.t96 vdd.n1342 6.46231
R21980 vdd.n2175 vdd.t172 6.46231
R21981 vdd.t175 vdd.n846 6.46231
R21982 vdd.n2757 vdd.t178 6.46231
R21983 vdd.t194 vdd.n671 6.46231
R21984 vdd.n3154 vdd.t102 6.46231
R21985 vdd.n2251 vdd.t206 6.34895
R21986 vdd.n2630 vdd.t191 6.34895
R21987 vdd.n2772 vdd.n687 6.2444
R21988 vdd.n2191 vdd.n2190 6.2444
R21989 vdd.n1911 vdd.t92 6.23558
R21990 vdd.t124 vdd.n308 6.23558
R21991 vdd.n3320 vdd.n297 6.22547
R21992 vdd.n1615 vdd.n1614 6.22547
R21993 vdd.n2212 vdd.t199 5.89549
R21994 vdd.n715 vdd.t176 5.89549
R21995 vdd.n272 vdd.n271 5.81868
R21996 vdd.n225 vdd.n224 5.81868
R21997 vdd.n182 vdd.n181 5.81868
R21998 vdd.n135 vdd.n134 5.81868
R21999 vdd.n93 vdd.n92 5.81868
R22000 vdd.n46 vdd.n45 5.81868
R22001 vdd.n1542 vdd.n1541 5.81868
R22002 vdd.n1589 vdd.n1588 5.81868
R22003 vdd.n1452 vdd.n1451 5.81868
R22004 vdd.n1499 vdd.n1498 5.81868
R22005 vdd.n1363 vdd.n1362 5.81868
R22006 vdd.n1410 vdd.n1409 5.81868
R22007 vdd.n2334 vdd.n2333 5.77611
R22008 vdd.n1139 vdd.n1138 5.77611
R22009 vdd.n2642 vdd.n2641 5.77611
R22010 vdd.n2886 vdd.n2885 5.77611
R22011 vdd.n2950 vdd.n591 5.77611
R22012 vdd.n2505 vdd.n2439 5.77611
R22013 vdd.n2259 vdd.n802 5.77611
R22014 vdd.n1275 vdd.n1107 5.77611
R22015 vdd.n1778 vdd.n1777 5.62474
R22016 vdd.n1978 vdd.n1975 5.62474
R22017 vdd.n3182 vdd.n3179 5.62474
R22018 vdd.n2985 vdd.n2982 5.62474
R22019 vdd.n2187 vdd.t188 5.55539
R22020 vdd.n691 vdd.t168 5.55539
R22021 vdd.n1635 vdd.t92 5.10193
R22022 vdd.n3307 vdd.t124 5.10193
R22023 vdd.n275 vdd.n266 5.04292
R22024 vdd.n228 vdd.n219 5.04292
R22025 vdd.n185 vdd.n176 5.04292
R22026 vdd.n138 vdd.n129 5.04292
R22027 vdd.n96 vdd.n87 5.04292
R22028 vdd.n49 vdd.n40 5.04292
R22029 vdd.n1545 vdd.n1536 5.04292
R22030 vdd.n1592 vdd.n1583 5.04292
R22031 vdd.n1455 vdd.n1446 5.04292
R22032 vdd.n1502 vdd.n1493 5.04292
R22033 vdd.n1366 vdd.n1357 5.04292
R22034 vdd.n1413 vdd.n1404 5.04292
R22035 vdd.n1928 vdd.t96 4.8752
R22036 vdd.t171 vdd.t180 4.8752
R22037 vdd.t210 vdd.t156 4.8752
R22038 vdd.t102 vdd.n304 4.8752
R22039 vdd.n2335 vdd.n2334 4.83952
R22040 vdd.n1138 vdd.n1137 4.83952
R22041 vdd.n2643 vdd.n2642 4.83952
R22042 vdd.n2887 vdd.n2886 4.83952
R22043 vdd.n591 vdd.n586 4.83952
R22044 vdd.n2502 vdd.n2439 4.83952
R22045 vdd.n2262 vdd.n802 4.83952
R22046 vdd.n1278 vdd.n1107 4.83952
R22047 vdd.n1189 vdd.t164 4.76184
R22048 vdd.n2715 vdd.t162 4.76184
R22049 vdd.n1983 vdd.n1982 4.74817
R22050 vdd.n1311 vdd.n1306 4.74817
R22051 vdd.n973 vdd.n970 4.74817
R22052 vdd.n2076 vdd.n969 4.74817
R22053 vdd.n2081 vdd.n970 4.74817
R22054 vdd.n2080 vdd.n969 4.74817
R22055 vdd.n3110 vdd.n3109 4.74817
R22056 vdd.n3107 vdd.n3106 4.74817
R22057 vdd.n3107 vdd.n521 4.74817
R22058 vdd.n3109 vdd.n518 4.74817
R22059 vdd.n2992 vdd.n573 4.74817
R22060 vdd.n2988 vdd.n574 4.74817
R22061 vdd.n2991 vdd.n574 4.74817
R22062 vdd.n2995 vdd.n573 4.74817
R22063 vdd.n1982 vdd.n1069 4.74817
R22064 vdd.n1308 vdd.n1306 4.74817
R22065 vdd.n297 vdd.n296 4.7074
R22066 vdd.n207 vdd.n206 4.7074
R22067 vdd.n1614 vdd.n1613 4.7074
R22068 vdd.n1524 vdd.n1523 4.7074
R22069 vdd.n1944 vdd.t114 4.64847
R22070 vdd.t173 vdd.n877 4.64847
R22071 vdd.n2206 vdd.t208 4.64847
R22072 vdd.t197 vdd.n702 4.64847
R22073 vdd.n2788 vdd.t193 4.64847
R22074 vdd.n3138 vdd.t126 4.64847
R22075 vdd.n866 vdd.t77 4.53511
R22076 vdd.n2770 vdd.t39 4.53511
R22077 vdd.n2133 vdd.t21 4.42174
R22078 vdd.n1189 vdd.t66 4.42174
R22079 vdd.n2715 vdd.t73 4.42174
R22080 vdd.n636 vdd.t17 4.42174
R22081 vdd.n2761 vdd.n687 4.37123
R22082 vdd.n2192 vdd.n2191 4.37123
R22083 vdd.n2230 vdd.t195 4.30838
R22084 vdd.n2618 vdd.t182 4.30838
R22085 vdd.n276 vdd.n264 4.26717
R22086 vdd.n229 vdd.n217 4.26717
R22087 vdd.n186 vdd.n174 4.26717
R22088 vdd.n139 vdd.n127 4.26717
R22089 vdd.n97 vdd.n85 4.26717
R22090 vdd.n50 vdd.n38 4.26717
R22091 vdd.n1546 vdd.n1534 4.26717
R22092 vdd.n1593 vdd.n1581 4.26717
R22093 vdd.n1456 vdd.n1444 4.26717
R22094 vdd.n1503 vdd.n1491 4.26717
R22095 vdd.n1367 vdd.n1355 4.26717
R22096 vdd.n1414 vdd.n1402 4.26717
R22097 vdd.n297 vdd.n207 4.10845
R22098 vdd.n1614 vdd.n1524 4.10845
R22099 vdd.n253 vdd.t109 4.06363
R22100 vdd.n253 vdd.t135 4.06363
R22101 vdd.n251 vdd.t146 4.06363
R22102 vdd.n251 vdd.t152 4.06363
R22103 vdd.n249 vdd.t154 4.06363
R22104 vdd.n249 vdd.t116 4.06363
R22105 vdd.n163 vdd.t99 4.06363
R22106 vdd.n163 vdd.t125 4.06363
R22107 vdd.n161 vdd.t143 4.06363
R22108 vdd.n161 vdd.t147 4.06363
R22109 vdd.n159 vdd.t151 4.06363
R22110 vdd.n159 vdd.t101 4.06363
R22111 vdd.n74 vdd.t108 4.06363
R22112 vdd.n74 vdd.t144 4.06363
R22113 vdd.n72 vdd.t103 4.06363
R22114 vdd.n72 vdd.t140 4.06363
R22115 vdd.n70 vdd.t118 4.06363
R22116 vdd.n70 vdd.t148 4.06363
R22117 vdd.n1566 vdd.t138 4.06363
R22118 vdd.n1566 vdd.t137 4.06363
R22119 vdd.n1568 vdd.t119 4.06363
R22120 vdd.n1568 vdd.t107 4.06363
R22121 vdd.n1570 vdd.t105 4.06363
R22122 vdd.n1570 vdd.t136 4.06363
R22123 vdd.n1476 vdd.t133 4.06363
R22124 vdd.n1476 vdd.t131 4.06363
R22125 vdd.n1478 vdd.t111 4.06363
R22126 vdd.n1478 vdd.t97 4.06363
R22127 vdd.n1480 vdd.t93 4.06363
R22128 vdd.n1480 vdd.t129 4.06363
R22129 vdd.n1387 vdd.t149 4.06363
R22130 vdd.n1387 vdd.t155 4.06363
R22131 vdd.n1389 vdd.t141 4.06363
R22132 vdd.n1389 vdd.t104 4.06363
R22133 vdd.n1391 vdd.t134 4.06363
R22134 vdd.n1391 vdd.t113 4.06363
R22135 vdd.n902 vdd.t201 3.96828
R22136 vdd.n2224 vdd.t179 3.96828
R22137 vdd.n2612 vdd.t198 3.96828
R22138 vdd.n2806 vdd.t187 3.96828
R22139 vdd.n26 vdd.t13 3.9605
R22140 vdd.n26 vdd.t9 3.9605
R22141 vdd.n23 vdd.t3 3.9605
R22142 vdd.n23 vdd.t10 3.9605
R22143 vdd.n21 vdd.t14 3.9605
R22144 vdd.n21 vdd.t5 3.9605
R22145 vdd.n20 vdd.t6 3.9605
R22146 vdd.n20 vdd.t12 3.9605
R22147 vdd.n15 vdd.t0 3.9605
R22148 vdd.n15 vdd.t1 3.9605
R22149 vdd.n16 vdd.t15 3.9605
R22150 vdd.n16 vdd.t7 3.9605
R22151 vdd.n18 vdd.t8 3.9605
R22152 vdd.n18 vdd.t11 3.9605
R22153 vdd.n25 vdd.t2 3.9605
R22154 vdd.n25 vdd.t4 3.9605
R22155 vdd.n2157 vdd.t201 3.74155
R22156 vdd.n836 vdd.t179 3.74155
R22157 vdd.n2739 vdd.t198 3.74155
R22158 vdd.n660 vdd.t187 3.74155
R22159 vdd.n7 vdd.t211 3.61217
R22160 vdd.n7 vdd.t177 3.61217
R22161 vdd.n8 vdd.t183 3.61217
R22162 vdd.n8 vdd.t203 3.61217
R22163 vdd.n10 vdd.t192 3.61217
R22164 vdd.n10 vdd.t163 3.61217
R22165 vdd.n12 vdd.t167 3.61217
R22166 vdd.n12 vdd.t190 3.61217
R22167 vdd.n5 vdd.t205 3.61217
R22168 vdd.n5 vdd.t185 3.61217
R22169 vdd.n3 vdd.t165 3.61217
R22170 vdd.n3 vdd.t207 3.61217
R22171 vdd.n1 vdd.t159 3.61217
R22172 vdd.n1 vdd.t196 3.61217
R22173 vdd.n0 vdd.t200 3.61217
R22174 vdd.n0 vdd.t181 3.61217
R22175 vdd.n280 vdd.n279 3.49141
R22176 vdd.n233 vdd.n232 3.49141
R22177 vdd.n190 vdd.n189 3.49141
R22178 vdd.n143 vdd.n142 3.49141
R22179 vdd.n101 vdd.n100 3.49141
R22180 vdd.n54 vdd.n53 3.49141
R22181 vdd.n1550 vdd.n1549 3.49141
R22182 vdd.n1597 vdd.n1596 3.49141
R22183 vdd.n1460 vdd.n1459 3.49141
R22184 vdd.n1507 vdd.n1506 3.49141
R22185 vdd.n1371 vdd.n1370 3.49141
R22186 vdd.n1418 vdd.n1417 3.49141
R22187 vdd.t195 vdd.n818 3.40145
R22188 vdd.n2398 vdd.t204 3.40145
R22189 vdd.n2702 vdd.t189 3.40145
R22190 vdd.n2727 vdd.t182 3.40145
R22191 vdd.n927 vdd.t21 3.28809
R22192 vdd.n2251 vdd.t66 3.28809
R22193 vdd.n2630 vdd.t73 3.28809
R22194 vdd.n2875 vdd.t17 3.28809
R22195 vdd.n2169 vdd.t173 3.06136
R22196 vdd.n1227 vdd.t208 3.06136
R22197 vdd.n2751 vdd.t197 3.06136
R22198 vdd.t193 vdd.n664 3.06136
R22199 vdd.n2244 vdd.t164 2.94799
R22200 vdd.t162 vdd.n736 2.94799
R22201 vdd.n1945 vdd.t130 2.83463
R22202 vdd.n1963 vdd.t25 2.83463
R22203 vdd.n3121 vdd.t35 2.83463
R22204 vdd.n467 vdd.t117 2.83463
R22205 vdd.n283 vdd.n262 2.71565
R22206 vdd.n236 vdd.n215 2.71565
R22207 vdd.n193 vdd.n172 2.71565
R22208 vdd.n146 vdd.n125 2.71565
R22209 vdd.n104 vdd.n83 2.71565
R22210 vdd.n57 vdd.n36 2.71565
R22211 vdd.n1553 vdd.n1532 2.71565
R22212 vdd.n1600 vdd.n1579 2.71565
R22213 vdd.n1463 vdd.n1442 2.71565
R22214 vdd.n1510 vdd.n1489 2.71565
R22215 vdd.n1374 vdd.n1353 2.71565
R22216 vdd.n1421 vdd.n1400 2.71565
R22217 vdd.t110 vdd.n1619 2.6079
R22218 vdd.n3315 vdd.t139 2.6079
R22219 vdd.n2218 vdd.t180 2.49453
R22220 vdd.n721 vdd.t210 2.49453
R22221 vdd.n270 vdd.n269 2.4129
R22222 vdd.n223 vdd.n222 2.4129
R22223 vdd.n180 vdd.n179 2.4129
R22224 vdd.n133 vdd.n132 2.4129
R22225 vdd.n91 vdd.n90 2.4129
R22226 vdd.n44 vdd.n43 2.4129
R22227 vdd.n1540 vdd.n1539 2.4129
R22228 vdd.n1587 vdd.n1586 2.4129
R22229 vdd.n1450 vdd.n1449 2.4129
R22230 vdd.n1497 vdd.n1496 2.4129
R22231 vdd.n1361 vdd.n1360 2.4129
R22232 vdd.n1408 vdd.n1407 2.4129
R22233 vdd.n1902 vdd.t94 2.38117
R22234 vdd.n3306 vdd.t121 2.38117
R22235 vdd.n2088 vdd.n970 2.27742
R22236 vdd.n2088 vdd.n969 2.27742
R22237 vdd.n3108 vdd.n3107 2.27742
R22238 vdd.n3109 vdd.n3108 2.27742
R22239 vdd.n2979 vdd.n574 2.27742
R22240 vdd.n2979 vdd.n573 2.27742
R22241 vdd.n1982 vdd.n1981 2.27742
R22242 vdd.n1981 vdd.n1306 2.27742
R22243 vdd.n873 vdd.t188 2.15444
R22244 vdd.n2194 vdd.t170 2.15444
R22245 vdd.n698 vdd.t169 2.15444
R22246 vdd.n2776 vdd.t168 2.15444
R22247 vdd.n284 vdd.n260 1.93989
R22248 vdd.n237 vdd.n213 1.93989
R22249 vdd.n194 vdd.n170 1.93989
R22250 vdd.n147 vdd.n123 1.93989
R22251 vdd.n105 vdd.n81 1.93989
R22252 vdd.n58 vdd.n34 1.93989
R22253 vdd.n1554 vdd.n1530 1.93989
R22254 vdd.n1601 vdd.n1577 1.93989
R22255 vdd.n1464 vdd.n1440 1.93989
R22256 vdd.n1511 vdd.n1487 1.93989
R22257 vdd.n1375 vdd.n1351 1.93989
R22258 vdd.n1422 vdd.n1398 1.93989
R22259 vdd.n1227 vdd.t199 1.81434
R22260 vdd.n2751 vdd.t176 1.81434
R22261 vdd.t206 vdd.n795 1.36088
R22262 vdd.n2709 vdd.t191 1.36088
R22263 vdd.n1910 vdd.t112 1.24752
R22264 vdd.t172 vdd.n870 1.24752
R22265 vdd.n2200 vdd.t175 1.24752
R22266 vdd.t178 vdd.n695 1.24752
R22267 vdd.n2782 vdd.t194 1.24752
R22268 vdd.t98 vdd.n3313 1.24752
R22269 vdd.n295 vdd.n255 1.16414
R22270 vdd.n288 vdd.n287 1.16414
R22271 vdd.n248 vdd.n208 1.16414
R22272 vdd.n241 vdd.n240 1.16414
R22273 vdd.n205 vdd.n165 1.16414
R22274 vdd.n198 vdd.n197 1.16414
R22275 vdd.n158 vdd.n118 1.16414
R22276 vdd.n151 vdd.n150 1.16414
R22277 vdd.n116 vdd.n76 1.16414
R22278 vdd.n109 vdd.n108 1.16414
R22279 vdd.n69 vdd.n29 1.16414
R22280 vdd.n62 vdd.n61 1.16414
R22281 vdd.n1565 vdd.n1525 1.16414
R22282 vdd.n1558 vdd.n1557 1.16414
R22283 vdd.n1612 vdd.n1572 1.16414
R22284 vdd.n1605 vdd.n1604 1.16414
R22285 vdd.n1475 vdd.n1435 1.16414
R22286 vdd.n1468 vdd.n1467 1.16414
R22287 vdd.n1522 vdd.n1482 1.16414
R22288 vdd.n1515 vdd.n1514 1.16414
R22289 vdd.n1386 vdd.n1346 1.16414
R22290 vdd.n1379 vdd.n1378 1.16414
R22291 vdd.n1433 vdd.n1393 1.16414
R22292 vdd.n1426 vdd.n1425 1.16414
R22293 vdd.n1615 vdd.n28 1.06035
R22294 vdd vdd.n3320 1.05252
R22295 vdd.n1936 vdd.t132 1.02079
R22296 vdd.t77 vdd.t170 1.02079
R22297 vdd.t169 vdd.t39 1.02079
R22298 vdd.t100 vdd.n456 1.02079
R22299 vdd.n1781 vdd.n1777 0.970197
R22300 vdd.n1979 vdd.n1978 0.970197
R22301 vdd.n3183 vdd.n3182 0.970197
R22302 vdd.n2987 vdd.n2985 0.970197
R22303 vdd.n2224 vdd.t158 0.907421
R22304 vdd.n2612 vdd.t202 0.907421
R22305 vdd.n1885 vdd.t43 0.567326
R22306 vdd.n909 vdd.t161 0.567326
R22307 vdd.n2230 vdd.t157 0.567326
R22308 vdd.n2618 vdd.t160 0.567326
R22309 vdd.n2812 vdd.t174 0.567326
R22310 vdd.n3298 vdd.t50 0.567326
R22311 vdd.n1969 vdd.n971 0.537085
R22312 vdd.n3117 vdd.n3116 0.537085
R22313 vdd.n3294 vdd.n3293 0.537085
R22314 vdd.n3176 vdd.n3175 0.537085
R22315 vdd.n2981 vdd.n476 0.537085
R22316 vdd.n1958 vdd.n1307 0.537085
R22317 vdd.n1779 vdd.n1644 0.537085
R22318 vdd.n1881 vdd.n1880 0.537085
R22319 vdd.n4 vdd.n2 0.459552
R22320 vdd.n11 vdd.n9 0.459552
R22321 vdd.n293 vdd.n292 0.388379
R22322 vdd.n259 vdd.n257 0.388379
R22323 vdd.n246 vdd.n245 0.388379
R22324 vdd.n212 vdd.n210 0.388379
R22325 vdd.n203 vdd.n202 0.388379
R22326 vdd.n169 vdd.n167 0.388379
R22327 vdd.n156 vdd.n155 0.388379
R22328 vdd.n122 vdd.n120 0.388379
R22329 vdd.n114 vdd.n113 0.388379
R22330 vdd.n80 vdd.n78 0.388379
R22331 vdd.n67 vdd.n66 0.388379
R22332 vdd.n33 vdd.n31 0.388379
R22333 vdd.n1563 vdd.n1562 0.388379
R22334 vdd.n1529 vdd.n1527 0.388379
R22335 vdd.n1610 vdd.n1609 0.388379
R22336 vdd.n1576 vdd.n1574 0.388379
R22337 vdd.n1473 vdd.n1472 0.388379
R22338 vdd.n1439 vdd.n1437 0.388379
R22339 vdd.n1520 vdd.n1519 0.388379
R22340 vdd.n1486 vdd.n1484 0.388379
R22341 vdd.n1384 vdd.n1383 0.388379
R22342 vdd.n1350 vdd.n1348 0.388379
R22343 vdd.n1431 vdd.n1430 0.388379
R22344 vdd.n1397 vdd.n1395 0.388379
R22345 vdd.n19 vdd.n17 0.387128
R22346 vdd.n24 vdd.n22 0.387128
R22347 vdd.n6 vdd.n4 0.358259
R22348 vdd.n13 vdd.n11 0.358259
R22349 vdd.n252 vdd.n250 0.358259
R22350 vdd.n254 vdd.n252 0.358259
R22351 vdd.n296 vdd.n254 0.358259
R22352 vdd.n162 vdd.n160 0.358259
R22353 vdd.n164 vdd.n162 0.358259
R22354 vdd.n206 vdd.n164 0.358259
R22355 vdd.n73 vdd.n71 0.358259
R22356 vdd.n75 vdd.n73 0.358259
R22357 vdd.n117 vdd.n75 0.358259
R22358 vdd.n1613 vdd.n1571 0.358259
R22359 vdd.n1571 vdd.n1569 0.358259
R22360 vdd.n1569 vdd.n1567 0.358259
R22361 vdd.n1523 vdd.n1481 0.358259
R22362 vdd.n1481 vdd.n1479 0.358259
R22363 vdd.n1479 vdd.n1477 0.358259
R22364 vdd.n1434 vdd.n1392 0.358259
R22365 vdd.n1392 vdd.n1390 0.358259
R22366 vdd.n1390 vdd.n1388 0.358259
R22367 vdd.n2163 vdd.t209 0.340595
R22368 vdd.n842 vdd.t171 0.340595
R22369 vdd.n2745 vdd.t156 0.340595
R22370 vdd.n667 vdd.t186 0.340595
R22371 vdd.n14 vdd.n6 0.334552
R22372 vdd.n14 vdd.n13 0.334552
R22373 vdd.n27 vdd.n19 0.21707
R22374 vdd.n27 vdd.n24 0.21707
R22375 vdd.n294 vdd.n256 0.155672
R22376 vdd.n286 vdd.n256 0.155672
R22377 vdd.n286 vdd.n285 0.155672
R22378 vdd.n285 vdd.n261 0.155672
R22379 vdd.n278 vdd.n261 0.155672
R22380 vdd.n278 vdd.n277 0.155672
R22381 vdd.n277 vdd.n265 0.155672
R22382 vdd.n270 vdd.n265 0.155672
R22383 vdd.n247 vdd.n209 0.155672
R22384 vdd.n239 vdd.n209 0.155672
R22385 vdd.n239 vdd.n238 0.155672
R22386 vdd.n238 vdd.n214 0.155672
R22387 vdd.n231 vdd.n214 0.155672
R22388 vdd.n231 vdd.n230 0.155672
R22389 vdd.n230 vdd.n218 0.155672
R22390 vdd.n223 vdd.n218 0.155672
R22391 vdd.n204 vdd.n166 0.155672
R22392 vdd.n196 vdd.n166 0.155672
R22393 vdd.n196 vdd.n195 0.155672
R22394 vdd.n195 vdd.n171 0.155672
R22395 vdd.n188 vdd.n171 0.155672
R22396 vdd.n188 vdd.n187 0.155672
R22397 vdd.n187 vdd.n175 0.155672
R22398 vdd.n180 vdd.n175 0.155672
R22399 vdd.n157 vdd.n119 0.155672
R22400 vdd.n149 vdd.n119 0.155672
R22401 vdd.n149 vdd.n148 0.155672
R22402 vdd.n148 vdd.n124 0.155672
R22403 vdd.n141 vdd.n124 0.155672
R22404 vdd.n141 vdd.n140 0.155672
R22405 vdd.n140 vdd.n128 0.155672
R22406 vdd.n133 vdd.n128 0.155672
R22407 vdd.n115 vdd.n77 0.155672
R22408 vdd.n107 vdd.n77 0.155672
R22409 vdd.n107 vdd.n106 0.155672
R22410 vdd.n106 vdd.n82 0.155672
R22411 vdd.n99 vdd.n82 0.155672
R22412 vdd.n99 vdd.n98 0.155672
R22413 vdd.n98 vdd.n86 0.155672
R22414 vdd.n91 vdd.n86 0.155672
R22415 vdd.n68 vdd.n30 0.155672
R22416 vdd.n60 vdd.n30 0.155672
R22417 vdd.n60 vdd.n59 0.155672
R22418 vdd.n59 vdd.n35 0.155672
R22419 vdd.n52 vdd.n35 0.155672
R22420 vdd.n52 vdd.n51 0.155672
R22421 vdd.n51 vdd.n39 0.155672
R22422 vdd.n44 vdd.n39 0.155672
R22423 vdd.n1564 vdd.n1526 0.155672
R22424 vdd.n1556 vdd.n1526 0.155672
R22425 vdd.n1556 vdd.n1555 0.155672
R22426 vdd.n1555 vdd.n1531 0.155672
R22427 vdd.n1548 vdd.n1531 0.155672
R22428 vdd.n1548 vdd.n1547 0.155672
R22429 vdd.n1547 vdd.n1535 0.155672
R22430 vdd.n1540 vdd.n1535 0.155672
R22431 vdd.n1611 vdd.n1573 0.155672
R22432 vdd.n1603 vdd.n1573 0.155672
R22433 vdd.n1603 vdd.n1602 0.155672
R22434 vdd.n1602 vdd.n1578 0.155672
R22435 vdd.n1595 vdd.n1578 0.155672
R22436 vdd.n1595 vdd.n1594 0.155672
R22437 vdd.n1594 vdd.n1582 0.155672
R22438 vdd.n1587 vdd.n1582 0.155672
R22439 vdd.n1474 vdd.n1436 0.155672
R22440 vdd.n1466 vdd.n1436 0.155672
R22441 vdd.n1466 vdd.n1465 0.155672
R22442 vdd.n1465 vdd.n1441 0.155672
R22443 vdd.n1458 vdd.n1441 0.155672
R22444 vdd.n1458 vdd.n1457 0.155672
R22445 vdd.n1457 vdd.n1445 0.155672
R22446 vdd.n1450 vdd.n1445 0.155672
R22447 vdd.n1521 vdd.n1483 0.155672
R22448 vdd.n1513 vdd.n1483 0.155672
R22449 vdd.n1513 vdd.n1512 0.155672
R22450 vdd.n1512 vdd.n1488 0.155672
R22451 vdd.n1505 vdd.n1488 0.155672
R22452 vdd.n1505 vdd.n1504 0.155672
R22453 vdd.n1504 vdd.n1492 0.155672
R22454 vdd.n1497 vdd.n1492 0.155672
R22455 vdd.n1385 vdd.n1347 0.155672
R22456 vdd.n1377 vdd.n1347 0.155672
R22457 vdd.n1377 vdd.n1376 0.155672
R22458 vdd.n1376 vdd.n1352 0.155672
R22459 vdd.n1369 vdd.n1352 0.155672
R22460 vdd.n1369 vdd.n1368 0.155672
R22461 vdd.n1368 vdd.n1356 0.155672
R22462 vdd.n1361 vdd.n1356 0.155672
R22463 vdd.n1432 vdd.n1394 0.155672
R22464 vdd.n1424 vdd.n1394 0.155672
R22465 vdd.n1424 vdd.n1423 0.155672
R22466 vdd.n1423 vdd.n1399 0.155672
R22467 vdd.n1416 vdd.n1399 0.155672
R22468 vdd.n1416 vdd.n1415 0.155672
R22469 vdd.n1415 vdd.n1403 0.155672
R22470 vdd.n1408 vdd.n1403 0.155672
R22471 vdd.n976 vdd.n968 0.152939
R22472 vdd.n980 vdd.n976 0.152939
R22473 vdd.n981 vdd.n980 0.152939
R22474 vdd.n982 vdd.n981 0.152939
R22475 vdd.n983 vdd.n982 0.152939
R22476 vdd.n987 vdd.n983 0.152939
R22477 vdd.n988 vdd.n987 0.152939
R22478 vdd.n989 vdd.n988 0.152939
R22479 vdd.n990 vdd.n989 0.152939
R22480 vdd.n994 vdd.n990 0.152939
R22481 vdd.n995 vdd.n994 0.152939
R22482 vdd.n996 vdd.n995 0.152939
R22483 vdd.n2052 vdd.n996 0.152939
R22484 vdd.n2052 vdd.n2051 0.152939
R22485 vdd.n2051 vdd.n2050 0.152939
R22486 vdd.n2050 vdd.n1002 0.152939
R22487 vdd.n1007 vdd.n1002 0.152939
R22488 vdd.n1008 vdd.n1007 0.152939
R22489 vdd.n1009 vdd.n1008 0.152939
R22490 vdd.n1013 vdd.n1009 0.152939
R22491 vdd.n1014 vdd.n1013 0.152939
R22492 vdd.n1015 vdd.n1014 0.152939
R22493 vdd.n1016 vdd.n1015 0.152939
R22494 vdd.n1020 vdd.n1016 0.152939
R22495 vdd.n1021 vdd.n1020 0.152939
R22496 vdd.n1022 vdd.n1021 0.152939
R22497 vdd.n1023 vdd.n1022 0.152939
R22498 vdd.n1027 vdd.n1023 0.152939
R22499 vdd.n1028 vdd.n1027 0.152939
R22500 vdd.n1029 vdd.n1028 0.152939
R22501 vdd.n1030 vdd.n1029 0.152939
R22502 vdd.n1034 vdd.n1030 0.152939
R22503 vdd.n1035 vdd.n1034 0.152939
R22504 vdd.n1036 vdd.n1035 0.152939
R22505 vdd.n2013 vdd.n1036 0.152939
R22506 vdd.n2013 vdd.n2012 0.152939
R22507 vdd.n2012 vdd.n2011 0.152939
R22508 vdd.n2011 vdd.n1042 0.152939
R22509 vdd.n1047 vdd.n1042 0.152939
R22510 vdd.n1048 vdd.n1047 0.152939
R22511 vdd.n1049 vdd.n1048 0.152939
R22512 vdd.n1053 vdd.n1049 0.152939
R22513 vdd.n1054 vdd.n1053 0.152939
R22514 vdd.n1055 vdd.n1054 0.152939
R22515 vdd.n1056 vdd.n1055 0.152939
R22516 vdd.n1060 vdd.n1056 0.152939
R22517 vdd.n1061 vdd.n1060 0.152939
R22518 vdd.n1062 vdd.n1061 0.152939
R22519 vdd.n1063 vdd.n1062 0.152939
R22520 vdd.n1067 vdd.n1063 0.152939
R22521 vdd.n1068 vdd.n1067 0.152939
R22522 vdd.n2087 vdd.n971 0.152939
R22523 vdd.n1932 vdd.n1931 0.152939
R22524 vdd.n1933 vdd.n1932 0.152939
R22525 vdd.n1933 vdd.n1334 0.152939
R22526 vdd.n1948 vdd.n1334 0.152939
R22527 vdd.n1949 vdd.n1948 0.152939
R22528 vdd.n1950 vdd.n1949 0.152939
R22529 vdd.n1950 vdd.n1322 0.152939
R22530 vdd.n1967 vdd.n1322 0.152939
R22531 vdd.n1968 vdd.n1967 0.152939
R22532 vdd.n1969 vdd.n1968 0.152939
R22533 vdd.n524 vdd.n519 0.152939
R22534 vdd.n525 vdd.n524 0.152939
R22535 vdd.n526 vdd.n525 0.152939
R22536 vdd.n527 vdd.n526 0.152939
R22537 vdd.n528 vdd.n527 0.152939
R22538 vdd.n529 vdd.n528 0.152939
R22539 vdd.n530 vdd.n529 0.152939
R22540 vdd.n531 vdd.n530 0.152939
R22541 vdd.n532 vdd.n531 0.152939
R22542 vdd.n533 vdd.n532 0.152939
R22543 vdd.n534 vdd.n533 0.152939
R22544 vdd.n535 vdd.n534 0.152939
R22545 vdd.n3075 vdd.n535 0.152939
R22546 vdd.n3075 vdd.n3074 0.152939
R22547 vdd.n3074 vdd.n3073 0.152939
R22548 vdd.n3073 vdd.n537 0.152939
R22549 vdd.n538 vdd.n537 0.152939
R22550 vdd.n539 vdd.n538 0.152939
R22551 vdd.n540 vdd.n539 0.152939
R22552 vdd.n541 vdd.n540 0.152939
R22553 vdd.n542 vdd.n541 0.152939
R22554 vdd.n543 vdd.n542 0.152939
R22555 vdd.n544 vdd.n543 0.152939
R22556 vdd.n545 vdd.n544 0.152939
R22557 vdd.n546 vdd.n545 0.152939
R22558 vdd.n547 vdd.n546 0.152939
R22559 vdd.n548 vdd.n547 0.152939
R22560 vdd.n549 vdd.n548 0.152939
R22561 vdd.n550 vdd.n549 0.152939
R22562 vdd.n551 vdd.n550 0.152939
R22563 vdd.n552 vdd.n551 0.152939
R22564 vdd.n553 vdd.n552 0.152939
R22565 vdd.n554 vdd.n553 0.152939
R22566 vdd.n555 vdd.n554 0.152939
R22567 vdd.n3029 vdd.n555 0.152939
R22568 vdd.n3029 vdd.n3028 0.152939
R22569 vdd.n3028 vdd.n3027 0.152939
R22570 vdd.n3027 vdd.n559 0.152939
R22571 vdd.n560 vdd.n559 0.152939
R22572 vdd.n561 vdd.n560 0.152939
R22573 vdd.n562 vdd.n561 0.152939
R22574 vdd.n563 vdd.n562 0.152939
R22575 vdd.n564 vdd.n563 0.152939
R22576 vdd.n565 vdd.n564 0.152939
R22577 vdd.n566 vdd.n565 0.152939
R22578 vdd.n567 vdd.n566 0.152939
R22579 vdd.n568 vdd.n567 0.152939
R22580 vdd.n569 vdd.n568 0.152939
R22581 vdd.n570 vdd.n569 0.152939
R22582 vdd.n571 vdd.n570 0.152939
R22583 vdd.n572 vdd.n571 0.152939
R22584 vdd.n3116 vdd.n481 0.152939
R22585 vdd.n3118 vdd.n3117 0.152939
R22586 vdd.n3118 vdd.n470 0.152939
R22587 vdd.n3133 vdd.n470 0.152939
R22588 vdd.n3134 vdd.n3133 0.152939
R22589 vdd.n3135 vdd.n3134 0.152939
R22590 vdd.n3135 vdd.n459 0.152939
R22591 vdd.n3149 vdd.n459 0.152939
R22592 vdd.n3150 vdd.n3149 0.152939
R22593 vdd.n3151 vdd.n3150 0.152939
R22594 vdd.n3151 vdd.n298 0.152939
R22595 vdd.n3318 vdd.n299 0.152939
R22596 vdd.n310 vdd.n299 0.152939
R22597 vdd.n311 vdd.n310 0.152939
R22598 vdd.n312 vdd.n311 0.152939
R22599 vdd.n320 vdd.n312 0.152939
R22600 vdd.n321 vdd.n320 0.152939
R22601 vdd.n322 vdd.n321 0.152939
R22602 vdd.n323 vdd.n322 0.152939
R22603 vdd.n331 vdd.n323 0.152939
R22604 vdd.n3294 vdd.n331 0.152939
R22605 vdd.n3293 vdd.n332 0.152939
R22606 vdd.n335 vdd.n332 0.152939
R22607 vdd.n339 vdd.n335 0.152939
R22608 vdd.n340 vdd.n339 0.152939
R22609 vdd.n341 vdd.n340 0.152939
R22610 vdd.n342 vdd.n341 0.152939
R22611 vdd.n343 vdd.n342 0.152939
R22612 vdd.n347 vdd.n343 0.152939
R22613 vdd.n348 vdd.n347 0.152939
R22614 vdd.n349 vdd.n348 0.152939
R22615 vdd.n350 vdd.n349 0.152939
R22616 vdd.n354 vdd.n350 0.152939
R22617 vdd.n355 vdd.n354 0.152939
R22618 vdd.n356 vdd.n355 0.152939
R22619 vdd.n357 vdd.n356 0.152939
R22620 vdd.n361 vdd.n357 0.152939
R22621 vdd.n362 vdd.n361 0.152939
R22622 vdd.n363 vdd.n362 0.152939
R22623 vdd.n3259 vdd.n363 0.152939
R22624 vdd.n3259 vdd.n3258 0.152939
R22625 vdd.n3258 vdd.n3257 0.152939
R22626 vdd.n3257 vdd.n369 0.152939
R22627 vdd.n374 vdd.n369 0.152939
R22628 vdd.n375 vdd.n374 0.152939
R22629 vdd.n376 vdd.n375 0.152939
R22630 vdd.n380 vdd.n376 0.152939
R22631 vdd.n381 vdd.n380 0.152939
R22632 vdd.n382 vdd.n381 0.152939
R22633 vdd.n383 vdd.n382 0.152939
R22634 vdd.n387 vdd.n383 0.152939
R22635 vdd.n388 vdd.n387 0.152939
R22636 vdd.n389 vdd.n388 0.152939
R22637 vdd.n390 vdd.n389 0.152939
R22638 vdd.n394 vdd.n390 0.152939
R22639 vdd.n395 vdd.n394 0.152939
R22640 vdd.n396 vdd.n395 0.152939
R22641 vdd.n397 vdd.n396 0.152939
R22642 vdd.n401 vdd.n397 0.152939
R22643 vdd.n402 vdd.n401 0.152939
R22644 vdd.n403 vdd.n402 0.152939
R22645 vdd.n3220 vdd.n403 0.152939
R22646 vdd.n3220 vdd.n3219 0.152939
R22647 vdd.n3219 vdd.n3218 0.152939
R22648 vdd.n3218 vdd.n409 0.152939
R22649 vdd.n414 vdd.n409 0.152939
R22650 vdd.n415 vdd.n414 0.152939
R22651 vdd.n416 vdd.n415 0.152939
R22652 vdd.n420 vdd.n416 0.152939
R22653 vdd.n421 vdd.n420 0.152939
R22654 vdd.n422 vdd.n421 0.152939
R22655 vdd.n423 vdd.n422 0.152939
R22656 vdd.n427 vdd.n423 0.152939
R22657 vdd.n428 vdd.n427 0.152939
R22658 vdd.n429 vdd.n428 0.152939
R22659 vdd.n430 vdd.n429 0.152939
R22660 vdd.n434 vdd.n430 0.152939
R22661 vdd.n435 vdd.n434 0.152939
R22662 vdd.n436 vdd.n435 0.152939
R22663 vdd.n437 vdd.n436 0.152939
R22664 vdd.n441 vdd.n437 0.152939
R22665 vdd.n442 vdd.n441 0.152939
R22666 vdd.n443 vdd.n442 0.152939
R22667 vdd.n3176 vdd.n443 0.152939
R22668 vdd.n3124 vdd.n476 0.152939
R22669 vdd.n3125 vdd.n3124 0.152939
R22670 vdd.n3126 vdd.n3125 0.152939
R22671 vdd.n3126 vdd.n464 0.152939
R22672 vdd.n3141 vdd.n464 0.152939
R22673 vdd.n3142 vdd.n3141 0.152939
R22674 vdd.n3143 vdd.n3142 0.152939
R22675 vdd.n3143 vdd.n452 0.152939
R22676 vdd.n3157 vdd.n452 0.152939
R22677 vdd.n3158 vdd.n3157 0.152939
R22678 vdd.n3159 vdd.n3158 0.152939
R22679 vdd.n3159 vdd.n450 0.152939
R22680 vdd.n3163 vdd.n450 0.152939
R22681 vdd.n3164 vdd.n3163 0.152939
R22682 vdd.n3165 vdd.n3164 0.152939
R22683 vdd.n3165 vdd.n447 0.152939
R22684 vdd.n3169 vdd.n447 0.152939
R22685 vdd.n3170 vdd.n3169 0.152939
R22686 vdd.n3171 vdd.n3170 0.152939
R22687 vdd.n3171 vdd.n444 0.152939
R22688 vdd.n3175 vdd.n444 0.152939
R22689 vdd.n2981 vdd.n2980 0.152939
R22690 vdd.n1980 vdd.n1307 0.152939
R22691 vdd.n1888 vdd.n1644 0.152939
R22692 vdd.n1889 vdd.n1888 0.152939
R22693 vdd.n1890 vdd.n1889 0.152939
R22694 vdd.n1890 vdd.n1632 0.152939
R22695 vdd.n1905 vdd.n1632 0.152939
R22696 vdd.n1906 vdd.n1905 0.152939
R22697 vdd.n1907 vdd.n1906 0.152939
R22698 vdd.n1907 vdd.n1622 0.152939
R22699 vdd.n1923 vdd.n1622 0.152939
R22700 vdd.n1924 vdd.n1923 0.152939
R22701 vdd.n1925 vdd.n1924 0.152939
R22702 vdd.n1925 vdd.n1339 0.152939
R22703 vdd.n1939 vdd.n1339 0.152939
R22704 vdd.n1940 vdd.n1939 0.152939
R22705 vdd.n1941 vdd.n1940 0.152939
R22706 vdd.n1941 vdd.n1329 0.152939
R22707 vdd.n1956 vdd.n1329 0.152939
R22708 vdd.n1957 vdd.n1956 0.152939
R22709 vdd.n1960 vdd.n1957 0.152939
R22710 vdd.n1960 vdd.n1959 0.152939
R22711 vdd.n1959 vdd.n1958 0.152939
R22712 vdd.n1880 vdd.n1649 0.152939
R22713 vdd.n1873 vdd.n1649 0.152939
R22714 vdd.n1873 vdd.n1872 0.152939
R22715 vdd.n1872 vdd.n1871 0.152939
R22716 vdd.n1871 vdd.n1686 0.152939
R22717 vdd.n1867 vdd.n1686 0.152939
R22718 vdd.n1867 vdd.n1866 0.152939
R22719 vdd.n1866 vdd.n1865 0.152939
R22720 vdd.n1865 vdd.n1692 0.152939
R22721 vdd.n1861 vdd.n1692 0.152939
R22722 vdd.n1861 vdd.n1860 0.152939
R22723 vdd.n1860 vdd.n1859 0.152939
R22724 vdd.n1859 vdd.n1698 0.152939
R22725 vdd.n1855 vdd.n1698 0.152939
R22726 vdd.n1855 vdd.n1854 0.152939
R22727 vdd.n1854 vdd.n1853 0.152939
R22728 vdd.n1853 vdd.n1704 0.152939
R22729 vdd.n1849 vdd.n1704 0.152939
R22730 vdd.n1849 vdd.n1848 0.152939
R22731 vdd.n1848 vdd.n1847 0.152939
R22732 vdd.n1847 vdd.n1712 0.152939
R22733 vdd.n1843 vdd.n1712 0.152939
R22734 vdd.n1843 vdd.n1842 0.152939
R22735 vdd.n1842 vdd.n1841 0.152939
R22736 vdd.n1841 vdd.n1718 0.152939
R22737 vdd.n1837 vdd.n1718 0.152939
R22738 vdd.n1837 vdd.n1836 0.152939
R22739 vdd.n1836 vdd.n1835 0.152939
R22740 vdd.n1835 vdd.n1724 0.152939
R22741 vdd.n1831 vdd.n1724 0.152939
R22742 vdd.n1831 vdd.n1830 0.152939
R22743 vdd.n1830 vdd.n1829 0.152939
R22744 vdd.n1829 vdd.n1730 0.152939
R22745 vdd.n1825 vdd.n1730 0.152939
R22746 vdd.n1825 vdd.n1824 0.152939
R22747 vdd.n1824 vdd.n1823 0.152939
R22748 vdd.n1823 vdd.n1736 0.152939
R22749 vdd.n1819 vdd.n1736 0.152939
R22750 vdd.n1819 vdd.n1818 0.152939
R22751 vdd.n1818 vdd.n1817 0.152939
R22752 vdd.n1817 vdd.n1742 0.152939
R22753 vdd.n1810 vdd.n1742 0.152939
R22754 vdd.n1810 vdd.n1809 0.152939
R22755 vdd.n1809 vdd.n1808 0.152939
R22756 vdd.n1808 vdd.n1747 0.152939
R22757 vdd.n1804 vdd.n1747 0.152939
R22758 vdd.n1804 vdd.n1803 0.152939
R22759 vdd.n1803 vdd.n1802 0.152939
R22760 vdd.n1802 vdd.n1753 0.152939
R22761 vdd.n1798 vdd.n1753 0.152939
R22762 vdd.n1798 vdd.n1797 0.152939
R22763 vdd.n1797 vdd.n1796 0.152939
R22764 vdd.n1796 vdd.n1759 0.152939
R22765 vdd.n1792 vdd.n1759 0.152939
R22766 vdd.n1792 vdd.n1791 0.152939
R22767 vdd.n1791 vdd.n1790 0.152939
R22768 vdd.n1790 vdd.n1765 0.152939
R22769 vdd.n1786 vdd.n1765 0.152939
R22770 vdd.n1786 vdd.n1785 0.152939
R22771 vdd.n1785 vdd.n1784 0.152939
R22772 vdd.n1784 vdd.n1771 0.152939
R22773 vdd.n1780 vdd.n1771 0.152939
R22774 vdd.n1780 vdd.n1779 0.152939
R22775 vdd.n1882 vdd.n1881 0.152939
R22776 vdd.n1882 vdd.n1638 0.152939
R22777 vdd.n1897 vdd.n1638 0.152939
R22778 vdd.n1898 vdd.n1897 0.152939
R22779 vdd.n1899 vdd.n1898 0.152939
R22780 vdd.n1899 vdd.n1627 0.152939
R22781 vdd.n1914 vdd.n1627 0.152939
R22782 vdd.n1915 vdd.n1914 0.152939
R22783 vdd.n1917 vdd.n1915 0.152939
R22784 vdd.n1917 vdd.n1916 0.152939
R22785 vdd.n2088 vdd.n2087 0.110256
R22786 vdd.n3108 vdd.n481 0.110256
R22787 vdd.n2980 vdd.n2979 0.110256
R22788 vdd.n1981 vdd.n1980 0.110256
R22789 vdd.n1931 vdd.n1616 0.0695946
R22790 vdd.n3319 vdd.n298 0.0695946
R22791 vdd.n3319 vdd.n3318 0.0695946
R22792 vdd.n1916 vdd.n1616 0.0695946
R22793 vdd.n2088 vdd.n968 0.0431829
R22794 vdd.n1981 vdd.n1068 0.0431829
R22795 vdd.n3108 vdd.n519 0.0431829
R22796 vdd.n2979 vdd.n572 0.0431829
R22797 vdd vdd.n28 0.00833333
R22798 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R22799 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R22800 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R22801 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R22802 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R22803 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R22804 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R22805 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R22806 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R22807 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R22808 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R22809 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R22810 a_n2804_13878.n15 a_n2804_13878.t1 74.6477
R22811 a_n2804_13878.n20 a_n2804_13878.t2 74.2899
R22812 a_n2804_13878.n17 a_n2804_13878.t3 74.2899
R22813 a_n2804_13878.n16 a_n2804_13878.t0 74.2899
R22814 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R22815 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R22816 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R22817 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R22818 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R22819 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R22820 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R22821 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R22822 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R22823 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R22824 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R22825 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R22826 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R22827 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R22828 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R22829 a_n2804_13878.n18 a_n2804_13878.t6 3.61217
R22830 a_n2804_13878.n18 a_n2804_13878.t7 3.61217
R22831 a_n2804_13878.n14 a_n2804_13878.t4 3.61217
R22832 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R22833 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R22834 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R22835 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R22836 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R22837 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R22838 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R22839 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R22840 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R22841 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R22842 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R22843 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R22844 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R22845 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R22846 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R22847 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R22848 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R22849 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R22850 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R22851 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R22852 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R22853 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R22854 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R22855 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R22856 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R22857 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R22858 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R22859 a_n2982_8322.n28 a_n2982_8322.t20 74.6477
R22860 a_n2982_8322.n13 a_n2982_8322.t9 74.6477
R22861 a_n2982_8322.n1 a_n2982_8322.t35 74.6474
R22862 a_n2982_8322.n20 a_n2982_8322.t14 74.2899
R22863 a_n2982_8322.n10 a_n2982_8322.t15 74.2899
R22864 a_n2982_8322.n14 a_n2982_8322.t7 74.2899
R22865 a_n2982_8322.n15 a_n2982_8322.t10 74.2899
R22866 a_n2982_8322.n18 a_n2982_8322.t11 74.2899
R22867 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R22868 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R22869 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R22870 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R22871 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R22872 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R22873 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R22874 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R22875 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R22876 a_n2982_8322.n13 a_n2982_8322.n12 70.6783
R22877 a_n2982_8322.n17 a_n2982_8322.n16 70.6783
R22878 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R22879 a_n2982_8322.n20 a_n2982_8322.n19 24.9022
R22880 a_n2982_8322.n11 a_n2982_8322.t1 9.65181
R22881 a_n2982_8322.n19 a_n2982_8322.n18 8.38735
R22882 a_n2982_8322.n11 a_n2982_8322.n10 6.90998
R22883 a_n2982_8322.n19 a_n2982_8322.n11 5.3452
R22884 a_n2982_8322.n27 a_n2982_8322.t33 3.61217
R22885 a_n2982_8322.n27 a_n2982_8322.t29 3.61217
R22886 a_n2982_8322.n25 a_n2982_8322.t17 3.61217
R22887 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R22888 a_n2982_8322.n23 a_n2982_8322.t30 3.61217
R22889 a_n2982_8322.n23 a_n2982_8322.t23 3.61217
R22890 a_n2982_8322.n21 a_n2982_8322.t27 3.61217
R22891 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R22892 a_n2982_8322.n0 a_n2982_8322.t28 3.61217
R22893 a_n2982_8322.n0 a_n2982_8322.t24 3.61217
R22894 a_n2982_8322.n2 a_n2982_8322.t21 3.61217
R22895 a_n2982_8322.n2 a_n2982_8322.t37 3.61217
R22896 a_n2982_8322.n4 a_n2982_8322.t34 3.61217
R22897 a_n2982_8322.n4 a_n2982_8322.t22 3.61217
R22898 a_n2982_8322.n6 a_n2982_8322.t19 3.61217
R22899 a_n2982_8322.n6 a_n2982_8322.t18 3.61217
R22900 a_n2982_8322.n8 a_n2982_8322.t32 3.61217
R22901 a_n2982_8322.n8 a_n2982_8322.t31 3.61217
R22902 a_n2982_8322.n12 a_n2982_8322.t13 3.61217
R22903 a_n2982_8322.n12 a_n2982_8322.t12 3.61217
R22904 a_n2982_8322.n16 a_n2982_8322.t8 3.61217
R22905 a_n2982_8322.n16 a_n2982_8322.t6 3.61217
R22906 a_n2982_8322.t36 a_n2982_8322.n30 3.61217
R22907 a_n2982_8322.n30 a_n2982_8322.t26 3.61217
R22908 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R22909 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R22910 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R22911 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R22912 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R22913 a_n2982_8322.n18 a_n2982_8322.n17 0.358259
R22914 a_n2982_8322.n17 a_n2982_8322.n15 0.358259
R22915 a_n2982_8322.n14 a_n2982_8322.n13 0.358259
R22916 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R22917 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R22918 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R22919 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R22920 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R22921 a_n2982_8322.n15 a_n2982_8322.n14 0.101793
R22922 a_n2982_8322.t4 a_n2982_8322.t2 0.0788333
R22923 a_n2982_8322.t0 a_n2982_8322.t5 0.0788333
R22924 a_n2982_8322.t1 a_n2982_8322.t3 0.0788333
R22925 a_n2982_8322.t0 a_n2982_8322.t4 0.0318333
R22926 a_n2982_8322.t1 a_n2982_8322.t5 0.0318333
R22927 a_n2982_8322.t2 a_n2982_8322.t5 0.0318333
R22928 a_n2982_8322.t3 a_n2982_8322.t0 0.0318333
R22929 minus.n53 minus.t28 323.478
R22930 minus.n11 minus.t8 323.478
R22931 minus.n82 minus.t13 297.12
R22932 minus.n80 minus.t15 297.12
R22933 minus.n44 minus.t5 297.12
R22934 minus.n74 minus.t6 297.12
R22935 minus.n46 minus.t26 297.12
R22936 minus.n68 minus.t21 297.12
R22937 minus.n48 minus.t23 297.12
R22938 minus.n62 minus.t16 297.12
R22939 minus.n50 minus.t17 297.12
R22940 minus.n56 minus.t9 297.12
R22941 minus.n52 minus.t27 297.12
R22942 minus.n10 minus.t7 297.12
R22943 minus.n14 minus.t11 297.12
R22944 minus.n16 minus.t10 297.12
R22945 minus.n20 minus.t12 297.12
R22946 minus.n22 minus.t20 297.12
R22947 minus.n26 minus.t18 297.12
R22948 minus.n28 minus.t25 297.12
R22949 minus.n32 minus.t24 297.12
R22950 minus.n34 minus.t14 297.12
R22951 minus.n38 minus.t22 297.12
R22952 minus.n40 minus.t19 297.12
R22953 minus.n88 minus.t2 243.255
R22954 minus.n87 minus.n85 224.169
R22955 minus.n87 minus.n86 223.454
R22956 minus.n55 minus.n54 161.3
R22957 minus.n56 minus.n51 161.3
R22958 minus.n58 minus.n57 161.3
R22959 minus.n59 minus.n50 161.3
R22960 minus.n61 minus.n60 161.3
R22961 minus.n62 minus.n49 161.3
R22962 minus.n64 minus.n63 161.3
R22963 minus.n65 minus.n48 161.3
R22964 minus.n67 minus.n66 161.3
R22965 minus.n68 minus.n47 161.3
R22966 minus.n70 minus.n69 161.3
R22967 minus.n71 minus.n46 161.3
R22968 minus.n73 minus.n72 161.3
R22969 minus.n74 minus.n45 161.3
R22970 minus.n76 minus.n75 161.3
R22971 minus.n77 minus.n44 161.3
R22972 minus.n79 minus.n78 161.3
R22973 minus.n80 minus.n43 161.3
R22974 minus.n81 minus.n42 161.3
R22975 minus.n83 minus.n82 161.3
R22976 minus.n41 minus.n40 161.3
R22977 minus.n39 minus.n0 161.3
R22978 minus.n38 minus.n37 161.3
R22979 minus.n36 minus.n1 161.3
R22980 minus.n35 minus.n34 161.3
R22981 minus.n33 minus.n2 161.3
R22982 minus.n32 minus.n31 161.3
R22983 minus.n30 minus.n3 161.3
R22984 minus.n29 minus.n28 161.3
R22985 minus.n27 minus.n4 161.3
R22986 minus.n26 minus.n25 161.3
R22987 minus.n24 minus.n5 161.3
R22988 minus.n23 minus.n22 161.3
R22989 minus.n21 minus.n6 161.3
R22990 minus.n20 minus.n19 161.3
R22991 minus.n18 minus.n7 161.3
R22992 minus.n17 minus.n16 161.3
R22993 minus.n15 minus.n8 161.3
R22994 minus.n14 minus.n13 161.3
R22995 minus.n12 minus.n9 161.3
R22996 minus.n82 minus.n81 46.0096
R22997 minus.n40 minus.n39 46.0096
R22998 minus.n12 minus.n11 45.0871
R22999 minus.n54 minus.n53 45.0871
R23000 minus.n80 minus.n79 41.6278
R23001 minus.n55 minus.n52 41.6278
R23002 minus.n10 minus.n9 41.6278
R23003 minus.n38 minus.n1 41.6278
R23004 minus.n75 minus.n44 37.246
R23005 minus.n57 minus.n56 37.246
R23006 minus.n15 minus.n14 37.246
R23007 minus.n34 minus.n33 37.246
R23008 minus.n84 minus.n83 33.3925
R23009 minus.n74 minus.n73 32.8641
R23010 minus.n61 minus.n50 32.8641
R23011 minus.n16 minus.n7 32.8641
R23012 minus.n32 minus.n3 32.8641
R23013 minus.n69 minus.n46 28.4823
R23014 minus.n63 minus.n62 28.4823
R23015 minus.n21 minus.n20 28.4823
R23016 minus.n28 minus.n27 28.4823
R23017 minus.n68 minus.n67 24.1005
R23018 minus.n67 minus.n48 24.1005
R23019 minus.n22 minus.n5 24.1005
R23020 minus.n26 minus.n5 24.1005
R23021 minus.n86 minus.t4 19.8005
R23022 minus.n86 minus.t3 19.8005
R23023 minus.n85 minus.t1 19.8005
R23024 minus.n85 minus.t0 19.8005
R23025 minus.n69 minus.n68 19.7187
R23026 minus.n63 minus.n48 19.7187
R23027 minus.n22 minus.n21 19.7187
R23028 minus.n27 minus.n26 19.7187
R23029 minus.n73 minus.n46 15.3369
R23030 minus.n62 minus.n61 15.3369
R23031 minus.n20 minus.n7 15.3369
R23032 minus.n28 minus.n3 15.3369
R23033 minus.n53 minus.n52 14.1472
R23034 minus.n11 minus.n10 14.1472
R23035 minus.n84 minus.n41 12.0933
R23036 minus minus.n89 11.4112
R23037 minus.n75 minus.n74 10.955
R23038 minus.n57 minus.n50 10.955
R23039 minus.n16 minus.n15 10.955
R23040 minus.n33 minus.n32 10.955
R23041 minus.n79 minus.n44 6.57323
R23042 minus.n56 minus.n55 6.57323
R23043 minus.n14 minus.n9 6.57323
R23044 minus.n34 minus.n1 6.57323
R23045 minus.n89 minus.n88 4.80222
R23046 minus.n81 minus.n80 2.19141
R23047 minus.n39 minus.n38 2.19141
R23048 minus.n89 minus.n84 0.972091
R23049 minus.n88 minus.n87 0.716017
R23050 minus.n83 minus.n42 0.189894
R23051 minus.n43 minus.n42 0.189894
R23052 minus.n78 minus.n43 0.189894
R23053 minus.n78 minus.n77 0.189894
R23054 minus.n77 minus.n76 0.189894
R23055 minus.n76 minus.n45 0.189894
R23056 minus.n72 minus.n45 0.189894
R23057 minus.n72 minus.n71 0.189894
R23058 minus.n71 minus.n70 0.189894
R23059 minus.n70 minus.n47 0.189894
R23060 minus.n66 minus.n47 0.189894
R23061 minus.n66 minus.n65 0.189894
R23062 minus.n65 minus.n64 0.189894
R23063 minus.n64 minus.n49 0.189894
R23064 minus.n60 minus.n49 0.189894
R23065 minus.n60 minus.n59 0.189894
R23066 minus.n59 minus.n58 0.189894
R23067 minus.n58 minus.n51 0.189894
R23068 minus.n54 minus.n51 0.189894
R23069 minus.n13 minus.n12 0.189894
R23070 minus.n13 minus.n8 0.189894
R23071 minus.n17 minus.n8 0.189894
R23072 minus.n18 minus.n17 0.189894
R23073 minus.n19 minus.n18 0.189894
R23074 minus.n19 minus.n6 0.189894
R23075 minus.n23 minus.n6 0.189894
R23076 minus.n24 minus.n23 0.189894
R23077 minus.n25 minus.n24 0.189894
R23078 minus.n25 minus.n4 0.189894
R23079 minus.n29 minus.n4 0.189894
R23080 minus.n30 minus.n29 0.189894
R23081 minus.n31 minus.n30 0.189894
R23082 minus.n31 minus.n2 0.189894
R23083 minus.n35 minus.n2 0.189894
R23084 minus.n36 minus.n35 0.189894
R23085 minus.n37 minus.n36 0.189894
R23086 minus.n37 minus.n0 0.189894
R23087 minus.n41 minus.n0 0.189894
R23088 output.n41 output.n15 289.615
R23089 output.n72 output.n46 289.615
R23090 output.n104 output.n78 289.615
R23091 output.n136 output.n110 289.615
R23092 output.n77 output.n45 197.26
R23093 output.n77 output.n76 196.298
R23094 output.n109 output.n108 196.298
R23095 output.n141 output.n140 196.298
R23096 output.n42 output.n41 185
R23097 output.n40 output.n39 185
R23098 output.n19 output.n18 185
R23099 output.n34 output.n33 185
R23100 output.n32 output.n31 185
R23101 output.n23 output.n22 185
R23102 output.n26 output.n25 185
R23103 output.n73 output.n72 185
R23104 output.n71 output.n70 185
R23105 output.n50 output.n49 185
R23106 output.n65 output.n64 185
R23107 output.n63 output.n62 185
R23108 output.n54 output.n53 185
R23109 output.n57 output.n56 185
R23110 output.n105 output.n104 185
R23111 output.n103 output.n102 185
R23112 output.n82 output.n81 185
R23113 output.n97 output.n96 185
R23114 output.n95 output.n94 185
R23115 output.n86 output.n85 185
R23116 output.n89 output.n88 185
R23117 output.n137 output.n136 185
R23118 output.n135 output.n134 185
R23119 output.n114 output.n113 185
R23120 output.n129 output.n128 185
R23121 output.n127 output.n126 185
R23122 output.n118 output.n117 185
R23123 output.n121 output.n120 185
R23124 output.t16 output.n24 147.661
R23125 output.t19 output.n55 147.661
R23126 output.t18 output.n87 147.661
R23127 output.t17 output.n119 147.661
R23128 output.n41 output.n40 104.615
R23129 output.n40 output.n18 104.615
R23130 output.n33 output.n18 104.615
R23131 output.n33 output.n32 104.615
R23132 output.n32 output.n22 104.615
R23133 output.n25 output.n22 104.615
R23134 output.n72 output.n71 104.615
R23135 output.n71 output.n49 104.615
R23136 output.n64 output.n49 104.615
R23137 output.n64 output.n63 104.615
R23138 output.n63 output.n53 104.615
R23139 output.n56 output.n53 104.615
R23140 output.n104 output.n103 104.615
R23141 output.n103 output.n81 104.615
R23142 output.n96 output.n81 104.615
R23143 output.n96 output.n95 104.615
R23144 output.n95 output.n85 104.615
R23145 output.n88 output.n85 104.615
R23146 output.n136 output.n135 104.615
R23147 output.n135 output.n113 104.615
R23148 output.n128 output.n113 104.615
R23149 output.n128 output.n127 104.615
R23150 output.n127 output.n117 104.615
R23151 output.n120 output.n117 104.615
R23152 output.n1 output.t1 77.056
R23153 output.n14 output.t3 76.6694
R23154 output.n1 output.n0 72.7095
R23155 output.n3 output.n2 72.7095
R23156 output.n5 output.n4 72.7095
R23157 output.n7 output.n6 72.7095
R23158 output.n9 output.n8 72.7095
R23159 output.n11 output.n10 72.7095
R23160 output.n13 output.n12 72.7095
R23161 output.n25 output.t16 52.3082
R23162 output.n56 output.t19 52.3082
R23163 output.n88 output.t18 52.3082
R23164 output.n120 output.t17 52.3082
R23165 output.n26 output.n24 15.6674
R23166 output.n57 output.n55 15.6674
R23167 output.n89 output.n87 15.6674
R23168 output.n121 output.n119 15.6674
R23169 output.n27 output.n23 12.8005
R23170 output.n58 output.n54 12.8005
R23171 output.n90 output.n86 12.8005
R23172 output.n122 output.n118 12.8005
R23173 output.n31 output.n30 12.0247
R23174 output.n62 output.n61 12.0247
R23175 output.n94 output.n93 12.0247
R23176 output.n126 output.n125 12.0247
R23177 output.n34 output.n21 11.249
R23178 output.n65 output.n52 11.249
R23179 output.n97 output.n84 11.249
R23180 output.n129 output.n116 11.249
R23181 output.n35 output.n19 10.4732
R23182 output.n66 output.n50 10.4732
R23183 output.n98 output.n82 10.4732
R23184 output.n130 output.n114 10.4732
R23185 output.n39 output.n38 9.69747
R23186 output.n70 output.n69 9.69747
R23187 output.n102 output.n101 9.69747
R23188 output.n134 output.n133 9.69747
R23189 output.n45 output.n44 9.45567
R23190 output.n76 output.n75 9.45567
R23191 output.n108 output.n107 9.45567
R23192 output.n140 output.n139 9.45567
R23193 output.n44 output.n43 9.3005
R23194 output.n17 output.n16 9.3005
R23195 output.n38 output.n37 9.3005
R23196 output.n36 output.n35 9.3005
R23197 output.n21 output.n20 9.3005
R23198 output.n30 output.n29 9.3005
R23199 output.n28 output.n27 9.3005
R23200 output.n75 output.n74 9.3005
R23201 output.n48 output.n47 9.3005
R23202 output.n69 output.n68 9.3005
R23203 output.n67 output.n66 9.3005
R23204 output.n52 output.n51 9.3005
R23205 output.n61 output.n60 9.3005
R23206 output.n59 output.n58 9.3005
R23207 output.n107 output.n106 9.3005
R23208 output.n80 output.n79 9.3005
R23209 output.n101 output.n100 9.3005
R23210 output.n99 output.n98 9.3005
R23211 output.n84 output.n83 9.3005
R23212 output.n93 output.n92 9.3005
R23213 output.n91 output.n90 9.3005
R23214 output.n139 output.n138 9.3005
R23215 output.n112 output.n111 9.3005
R23216 output.n133 output.n132 9.3005
R23217 output.n131 output.n130 9.3005
R23218 output.n116 output.n115 9.3005
R23219 output.n125 output.n124 9.3005
R23220 output.n123 output.n122 9.3005
R23221 output.n42 output.n17 8.92171
R23222 output.n73 output.n48 8.92171
R23223 output.n105 output.n80 8.92171
R23224 output.n137 output.n112 8.92171
R23225 output output.n141 8.15037
R23226 output.n43 output.n15 8.14595
R23227 output.n74 output.n46 8.14595
R23228 output.n106 output.n78 8.14595
R23229 output.n138 output.n110 8.14595
R23230 output.n45 output.n15 5.81868
R23231 output.n76 output.n46 5.81868
R23232 output.n108 output.n78 5.81868
R23233 output.n140 output.n110 5.81868
R23234 output.n43 output.n42 5.04292
R23235 output.n74 output.n73 5.04292
R23236 output.n106 output.n105 5.04292
R23237 output.n138 output.n137 5.04292
R23238 output.n28 output.n24 4.38594
R23239 output.n59 output.n55 4.38594
R23240 output.n91 output.n87 4.38594
R23241 output.n123 output.n119 4.38594
R23242 output.n39 output.n17 4.26717
R23243 output.n70 output.n48 4.26717
R23244 output.n102 output.n80 4.26717
R23245 output.n134 output.n112 4.26717
R23246 output.n0 output.t7 3.9605
R23247 output.n0 output.t12 3.9605
R23248 output.n2 output.t0 3.9605
R23249 output.n2 output.t8 3.9605
R23250 output.n4 output.t10 3.9605
R23251 output.n4 output.t9 3.9605
R23252 output.n6 output.t15 3.9605
R23253 output.n6 output.t2 3.9605
R23254 output.n8 output.t4 3.9605
R23255 output.n8 output.t13 3.9605
R23256 output.n10 output.t14 3.9605
R23257 output.n10 output.t5 3.9605
R23258 output.n12 output.t6 3.9605
R23259 output.n12 output.t11 3.9605
R23260 output.n38 output.n19 3.49141
R23261 output.n69 output.n50 3.49141
R23262 output.n101 output.n82 3.49141
R23263 output.n133 output.n114 3.49141
R23264 output.n35 output.n34 2.71565
R23265 output.n66 output.n65 2.71565
R23266 output.n98 output.n97 2.71565
R23267 output.n130 output.n129 2.71565
R23268 output.n31 output.n21 1.93989
R23269 output.n62 output.n52 1.93989
R23270 output.n94 output.n84 1.93989
R23271 output.n126 output.n116 1.93989
R23272 output.n30 output.n23 1.16414
R23273 output.n61 output.n54 1.16414
R23274 output.n93 output.n86 1.16414
R23275 output.n125 output.n118 1.16414
R23276 output.n141 output.n109 0.962709
R23277 output.n109 output.n77 0.962709
R23278 output.n27 output.n26 0.388379
R23279 output.n58 output.n57 0.388379
R23280 output.n90 output.n89 0.388379
R23281 output.n122 output.n121 0.388379
R23282 output.n14 output.n13 0.387128
R23283 output.n13 output.n11 0.387128
R23284 output.n11 output.n9 0.387128
R23285 output.n9 output.n7 0.387128
R23286 output.n7 output.n5 0.387128
R23287 output.n5 output.n3 0.387128
R23288 output.n3 output.n1 0.387128
R23289 output.n44 output.n16 0.155672
R23290 output.n37 output.n16 0.155672
R23291 output.n37 output.n36 0.155672
R23292 output.n36 output.n20 0.155672
R23293 output.n29 output.n20 0.155672
R23294 output.n29 output.n28 0.155672
R23295 output.n75 output.n47 0.155672
R23296 output.n68 output.n47 0.155672
R23297 output.n68 output.n67 0.155672
R23298 output.n67 output.n51 0.155672
R23299 output.n60 output.n51 0.155672
R23300 output.n60 output.n59 0.155672
R23301 output.n107 output.n79 0.155672
R23302 output.n100 output.n79 0.155672
R23303 output.n100 output.n99 0.155672
R23304 output.n99 output.n83 0.155672
R23305 output.n92 output.n83 0.155672
R23306 output.n92 output.n91 0.155672
R23307 output.n139 output.n111 0.155672
R23308 output.n132 output.n111 0.155672
R23309 output.n132 output.n131 0.155672
R23310 output.n131 output.n115 0.155672
R23311 output.n124 output.n115 0.155672
R23312 output.n124 output.n123 0.155672
R23313 output output.n14 0.126227
R23314 diffpairibias.n0 diffpairibias.t18 436.822
R23315 diffpairibias.n21 diffpairibias.t19 435.479
R23316 diffpairibias.n20 diffpairibias.t16 435.479
R23317 diffpairibias.n19 diffpairibias.t17 435.479
R23318 diffpairibias.n18 diffpairibias.t21 435.479
R23319 diffpairibias.n0 diffpairibias.t22 435.479
R23320 diffpairibias.n1 diffpairibias.t20 435.479
R23321 diffpairibias.n2 diffpairibias.t23 435.479
R23322 diffpairibias.n10 diffpairibias.t0 377.536
R23323 diffpairibias.n10 diffpairibias.t8 376.193
R23324 diffpairibias.n11 diffpairibias.t10 376.193
R23325 diffpairibias.n12 diffpairibias.t6 376.193
R23326 diffpairibias.n13 diffpairibias.t2 376.193
R23327 diffpairibias.n14 diffpairibias.t12 376.193
R23328 diffpairibias.n15 diffpairibias.t4 376.193
R23329 diffpairibias.n16 diffpairibias.t14 376.193
R23330 diffpairibias.n3 diffpairibias.t1 113.368
R23331 diffpairibias.n3 diffpairibias.t9 112.698
R23332 diffpairibias.n4 diffpairibias.t11 112.698
R23333 diffpairibias.n5 diffpairibias.t7 112.698
R23334 diffpairibias.n6 diffpairibias.t3 112.698
R23335 diffpairibias.n7 diffpairibias.t13 112.698
R23336 diffpairibias.n8 diffpairibias.t5 112.698
R23337 diffpairibias.n9 diffpairibias.t15 112.698
R23338 diffpairibias.n17 diffpairibias.n16 4.77242
R23339 diffpairibias.n17 diffpairibias.n9 4.30807
R23340 diffpairibias.n18 diffpairibias.n17 4.13945
R23341 diffpairibias.n16 diffpairibias.n15 1.34352
R23342 diffpairibias.n15 diffpairibias.n14 1.34352
R23343 diffpairibias.n14 diffpairibias.n13 1.34352
R23344 diffpairibias.n13 diffpairibias.n12 1.34352
R23345 diffpairibias.n12 diffpairibias.n11 1.34352
R23346 diffpairibias.n11 diffpairibias.n10 1.34352
R23347 diffpairibias.n2 diffpairibias.n1 1.34352
R23348 diffpairibias.n1 diffpairibias.n0 1.34352
R23349 diffpairibias.n19 diffpairibias.n18 1.34352
R23350 diffpairibias.n20 diffpairibias.n19 1.34352
R23351 diffpairibias.n21 diffpairibias.n20 1.34352
R23352 diffpairibias.n22 diffpairibias.n21 0.862419
R23353 diffpairibias diffpairibias.n22 0.684875
R23354 diffpairibias.n9 diffpairibias.n8 0.672012
R23355 diffpairibias.n8 diffpairibias.n7 0.672012
R23356 diffpairibias.n7 diffpairibias.n6 0.672012
R23357 diffpairibias.n6 diffpairibias.n5 0.672012
R23358 diffpairibias.n5 diffpairibias.n4 0.672012
R23359 diffpairibias.n4 diffpairibias.n3 0.672012
R23360 diffpairibias.n22 diffpairibias.n2 0.190907
R23361 outputibias.n27 outputibias.n1 289.615
R23362 outputibias.n58 outputibias.n32 289.615
R23363 outputibias.n90 outputibias.n64 289.615
R23364 outputibias.n122 outputibias.n96 289.615
R23365 outputibias.n28 outputibias.n27 185
R23366 outputibias.n26 outputibias.n25 185
R23367 outputibias.n5 outputibias.n4 185
R23368 outputibias.n20 outputibias.n19 185
R23369 outputibias.n18 outputibias.n17 185
R23370 outputibias.n9 outputibias.n8 185
R23371 outputibias.n12 outputibias.n11 185
R23372 outputibias.n59 outputibias.n58 185
R23373 outputibias.n57 outputibias.n56 185
R23374 outputibias.n36 outputibias.n35 185
R23375 outputibias.n51 outputibias.n50 185
R23376 outputibias.n49 outputibias.n48 185
R23377 outputibias.n40 outputibias.n39 185
R23378 outputibias.n43 outputibias.n42 185
R23379 outputibias.n91 outputibias.n90 185
R23380 outputibias.n89 outputibias.n88 185
R23381 outputibias.n68 outputibias.n67 185
R23382 outputibias.n83 outputibias.n82 185
R23383 outputibias.n81 outputibias.n80 185
R23384 outputibias.n72 outputibias.n71 185
R23385 outputibias.n75 outputibias.n74 185
R23386 outputibias.n123 outputibias.n122 185
R23387 outputibias.n121 outputibias.n120 185
R23388 outputibias.n100 outputibias.n99 185
R23389 outputibias.n115 outputibias.n114 185
R23390 outputibias.n113 outputibias.n112 185
R23391 outputibias.n104 outputibias.n103 185
R23392 outputibias.n107 outputibias.n106 185
R23393 outputibias.n0 outputibias.t10 178.945
R23394 outputibias.n133 outputibias.t8 177.018
R23395 outputibias.n132 outputibias.t11 177.018
R23396 outputibias.n0 outputibias.t9 177.018
R23397 outputibias.t7 outputibias.n10 147.661
R23398 outputibias.t1 outputibias.n41 147.661
R23399 outputibias.t3 outputibias.n73 147.661
R23400 outputibias.t5 outputibias.n105 147.661
R23401 outputibias.n128 outputibias.t6 132.363
R23402 outputibias.n128 outputibias.t0 130.436
R23403 outputibias.n129 outputibias.t2 130.436
R23404 outputibias.n130 outputibias.t4 130.436
R23405 outputibias.n27 outputibias.n26 104.615
R23406 outputibias.n26 outputibias.n4 104.615
R23407 outputibias.n19 outputibias.n4 104.615
R23408 outputibias.n19 outputibias.n18 104.615
R23409 outputibias.n18 outputibias.n8 104.615
R23410 outputibias.n11 outputibias.n8 104.615
R23411 outputibias.n58 outputibias.n57 104.615
R23412 outputibias.n57 outputibias.n35 104.615
R23413 outputibias.n50 outputibias.n35 104.615
R23414 outputibias.n50 outputibias.n49 104.615
R23415 outputibias.n49 outputibias.n39 104.615
R23416 outputibias.n42 outputibias.n39 104.615
R23417 outputibias.n90 outputibias.n89 104.615
R23418 outputibias.n89 outputibias.n67 104.615
R23419 outputibias.n82 outputibias.n67 104.615
R23420 outputibias.n82 outputibias.n81 104.615
R23421 outputibias.n81 outputibias.n71 104.615
R23422 outputibias.n74 outputibias.n71 104.615
R23423 outputibias.n122 outputibias.n121 104.615
R23424 outputibias.n121 outputibias.n99 104.615
R23425 outputibias.n114 outputibias.n99 104.615
R23426 outputibias.n114 outputibias.n113 104.615
R23427 outputibias.n113 outputibias.n103 104.615
R23428 outputibias.n106 outputibias.n103 104.615
R23429 outputibias.n63 outputibias.n31 95.6354
R23430 outputibias.n63 outputibias.n62 94.6732
R23431 outputibias.n95 outputibias.n94 94.6732
R23432 outputibias.n127 outputibias.n126 94.6732
R23433 outputibias.n11 outputibias.t7 52.3082
R23434 outputibias.n42 outputibias.t1 52.3082
R23435 outputibias.n74 outputibias.t3 52.3082
R23436 outputibias.n106 outputibias.t5 52.3082
R23437 outputibias.n12 outputibias.n10 15.6674
R23438 outputibias.n43 outputibias.n41 15.6674
R23439 outputibias.n75 outputibias.n73 15.6674
R23440 outputibias.n107 outputibias.n105 15.6674
R23441 outputibias.n13 outputibias.n9 12.8005
R23442 outputibias.n44 outputibias.n40 12.8005
R23443 outputibias.n76 outputibias.n72 12.8005
R23444 outputibias.n108 outputibias.n104 12.8005
R23445 outputibias.n17 outputibias.n16 12.0247
R23446 outputibias.n48 outputibias.n47 12.0247
R23447 outputibias.n80 outputibias.n79 12.0247
R23448 outputibias.n112 outputibias.n111 12.0247
R23449 outputibias.n20 outputibias.n7 11.249
R23450 outputibias.n51 outputibias.n38 11.249
R23451 outputibias.n83 outputibias.n70 11.249
R23452 outputibias.n115 outputibias.n102 11.249
R23453 outputibias.n21 outputibias.n5 10.4732
R23454 outputibias.n52 outputibias.n36 10.4732
R23455 outputibias.n84 outputibias.n68 10.4732
R23456 outputibias.n116 outputibias.n100 10.4732
R23457 outputibias.n25 outputibias.n24 9.69747
R23458 outputibias.n56 outputibias.n55 9.69747
R23459 outputibias.n88 outputibias.n87 9.69747
R23460 outputibias.n120 outputibias.n119 9.69747
R23461 outputibias.n31 outputibias.n30 9.45567
R23462 outputibias.n62 outputibias.n61 9.45567
R23463 outputibias.n94 outputibias.n93 9.45567
R23464 outputibias.n126 outputibias.n125 9.45567
R23465 outputibias.n30 outputibias.n29 9.3005
R23466 outputibias.n3 outputibias.n2 9.3005
R23467 outputibias.n24 outputibias.n23 9.3005
R23468 outputibias.n22 outputibias.n21 9.3005
R23469 outputibias.n7 outputibias.n6 9.3005
R23470 outputibias.n16 outputibias.n15 9.3005
R23471 outputibias.n14 outputibias.n13 9.3005
R23472 outputibias.n61 outputibias.n60 9.3005
R23473 outputibias.n34 outputibias.n33 9.3005
R23474 outputibias.n55 outputibias.n54 9.3005
R23475 outputibias.n53 outputibias.n52 9.3005
R23476 outputibias.n38 outputibias.n37 9.3005
R23477 outputibias.n47 outputibias.n46 9.3005
R23478 outputibias.n45 outputibias.n44 9.3005
R23479 outputibias.n93 outputibias.n92 9.3005
R23480 outputibias.n66 outputibias.n65 9.3005
R23481 outputibias.n87 outputibias.n86 9.3005
R23482 outputibias.n85 outputibias.n84 9.3005
R23483 outputibias.n70 outputibias.n69 9.3005
R23484 outputibias.n79 outputibias.n78 9.3005
R23485 outputibias.n77 outputibias.n76 9.3005
R23486 outputibias.n125 outputibias.n124 9.3005
R23487 outputibias.n98 outputibias.n97 9.3005
R23488 outputibias.n119 outputibias.n118 9.3005
R23489 outputibias.n117 outputibias.n116 9.3005
R23490 outputibias.n102 outputibias.n101 9.3005
R23491 outputibias.n111 outputibias.n110 9.3005
R23492 outputibias.n109 outputibias.n108 9.3005
R23493 outputibias.n28 outputibias.n3 8.92171
R23494 outputibias.n59 outputibias.n34 8.92171
R23495 outputibias.n91 outputibias.n66 8.92171
R23496 outputibias.n123 outputibias.n98 8.92171
R23497 outputibias.n29 outputibias.n1 8.14595
R23498 outputibias.n60 outputibias.n32 8.14595
R23499 outputibias.n92 outputibias.n64 8.14595
R23500 outputibias.n124 outputibias.n96 8.14595
R23501 outputibias.n31 outputibias.n1 5.81868
R23502 outputibias.n62 outputibias.n32 5.81868
R23503 outputibias.n94 outputibias.n64 5.81868
R23504 outputibias.n126 outputibias.n96 5.81868
R23505 outputibias.n131 outputibias.n130 5.20947
R23506 outputibias.n29 outputibias.n28 5.04292
R23507 outputibias.n60 outputibias.n59 5.04292
R23508 outputibias.n92 outputibias.n91 5.04292
R23509 outputibias.n124 outputibias.n123 5.04292
R23510 outputibias.n131 outputibias.n127 4.42209
R23511 outputibias.n14 outputibias.n10 4.38594
R23512 outputibias.n45 outputibias.n41 4.38594
R23513 outputibias.n77 outputibias.n73 4.38594
R23514 outputibias.n109 outputibias.n105 4.38594
R23515 outputibias.n132 outputibias.n131 4.28454
R23516 outputibias.n25 outputibias.n3 4.26717
R23517 outputibias.n56 outputibias.n34 4.26717
R23518 outputibias.n88 outputibias.n66 4.26717
R23519 outputibias.n120 outputibias.n98 4.26717
R23520 outputibias.n24 outputibias.n5 3.49141
R23521 outputibias.n55 outputibias.n36 3.49141
R23522 outputibias.n87 outputibias.n68 3.49141
R23523 outputibias.n119 outputibias.n100 3.49141
R23524 outputibias.n21 outputibias.n20 2.71565
R23525 outputibias.n52 outputibias.n51 2.71565
R23526 outputibias.n84 outputibias.n83 2.71565
R23527 outputibias.n116 outputibias.n115 2.71565
R23528 outputibias.n17 outputibias.n7 1.93989
R23529 outputibias.n48 outputibias.n38 1.93989
R23530 outputibias.n80 outputibias.n70 1.93989
R23531 outputibias.n112 outputibias.n102 1.93989
R23532 outputibias.n130 outputibias.n129 1.9266
R23533 outputibias.n129 outputibias.n128 1.9266
R23534 outputibias.n133 outputibias.n132 1.92658
R23535 outputibias.n134 outputibias.n133 1.29913
R23536 outputibias.n16 outputibias.n9 1.16414
R23537 outputibias.n47 outputibias.n40 1.16414
R23538 outputibias.n79 outputibias.n72 1.16414
R23539 outputibias.n111 outputibias.n104 1.16414
R23540 outputibias.n127 outputibias.n95 0.962709
R23541 outputibias.n95 outputibias.n63 0.962709
R23542 outputibias.n13 outputibias.n12 0.388379
R23543 outputibias.n44 outputibias.n43 0.388379
R23544 outputibias.n76 outputibias.n75 0.388379
R23545 outputibias.n108 outputibias.n107 0.388379
R23546 outputibias.n134 outputibias.n0 0.337251
R23547 outputibias outputibias.n134 0.302375
R23548 outputibias.n30 outputibias.n2 0.155672
R23549 outputibias.n23 outputibias.n2 0.155672
R23550 outputibias.n23 outputibias.n22 0.155672
R23551 outputibias.n22 outputibias.n6 0.155672
R23552 outputibias.n15 outputibias.n6 0.155672
R23553 outputibias.n15 outputibias.n14 0.155672
R23554 outputibias.n61 outputibias.n33 0.155672
R23555 outputibias.n54 outputibias.n33 0.155672
R23556 outputibias.n54 outputibias.n53 0.155672
R23557 outputibias.n53 outputibias.n37 0.155672
R23558 outputibias.n46 outputibias.n37 0.155672
R23559 outputibias.n46 outputibias.n45 0.155672
R23560 outputibias.n93 outputibias.n65 0.155672
R23561 outputibias.n86 outputibias.n65 0.155672
R23562 outputibias.n86 outputibias.n85 0.155672
R23563 outputibias.n85 outputibias.n69 0.155672
R23564 outputibias.n78 outputibias.n69 0.155672
R23565 outputibias.n78 outputibias.n77 0.155672
R23566 outputibias.n125 outputibias.n97 0.155672
R23567 outputibias.n118 outputibias.n97 0.155672
R23568 outputibias.n118 outputibias.n117 0.155672
R23569 outputibias.n117 outputibias.n101 0.155672
R23570 outputibias.n110 outputibias.n101 0.155672
R23571 outputibias.n110 outputibias.n109 0.155672
C0 plus commonsourceibias 0.415048f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13881f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 68.5846f
C6 commonsourceibias output 0.006808f
C7 minus diffpairibias 4.33e-19
C8 CSoutput minus 2.6584f
C9 vdd plus 0.080016f
C10 plus diffpairibias 4.56e-19
C11 commonsourceibias outputibias 0.003832f
C12 vdd commonsourceibias 0.004218f
C13 CSoutput plus 0.874787f
C14 commonsourceibias diffpairibias 0.06482f
C15 CSoutput commonsourceibias 54.0646f
C16 minus plus 9.59292f
C17 minus commonsourceibias 0.460231f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183172p
C22 plus gnd 35.9511f
C23 minus gnd 28.75612f
C24 CSoutput gnd 0.124923p
C25 vdd gnd 0.448485p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 output.t1 gnd 0.464308f
C221 output.t7 gnd 0.044422f
C222 output.t12 gnd 0.044422f
C223 output.n0 gnd 0.364624f
C224 output.n1 gnd 0.614102f
C225 output.t0 gnd 0.044422f
C226 output.t8 gnd 0.044422f
C227 output.n2 gnd 0.364624f
C228 output.n3 gnd 0.350265f
C229 output.t10 gnd 0.044422f
C230 output.t9 gnd 0.044422f
C231 output.n4 gnd 0.364624f
C232 output.n5 gnd 0.350265f
C233 output.t15 gnd 0.044422f
C234 output.t2 gnd 0.044422f
C235 output.n6 gnd 0.364624f
C236 output.n7 gnd 0.350265f
C237 output.t4 gnd 0.044422f
C238 output.t13 gnd 0.044422f
C239 output.n8 gnd 0.364624f
C240 output.n9 gnd 0.350265f
C241 output.t14 gnd 0.044422f
C242 output.t5 gnd 0.044422f
C243 output.n10 gnd 0.364624f
C244 output.n11 gnd 0.350265f
C245 output.t6 gnd 0.044422f
C246 output.t11 gnd 0.044422f
C247 output.n12 gnd 0.364624f
C248 output.n13 gnd 0.350265f
C249 output.t3 gnd 0.462979f
C250 output.n14 gnd 0.28994f
C251 output.n15 gnd 0.015803f
C252 output.n16 gnd 0.011243f
C253 output.n17 gnd 0.006041f
C254 output.n18 gnd 0.01428f
C255 output.n19 gnd 0.006397f
C256 output.n20 gnd 0.011243f
C257 output.n21 gnd 0.006041f
C258 output.n22 gnd 0.01428f
C259 output.n23 gnd 0.006397f
C260 output.n24 gnd 0.048111f
C261 output.t16 gnd 0.023274f
C262 output.n25 gnd 0.01071f
C263 output.n26 gnd 0.008435f
C264 output.n27 gnd 0.006041f
C265 output.n28 gnd 0.267512f
C266 output.n29 gnd 0.011243f
C267 output.n30 gnd 0.006041f
C268 output.n31 gnd 0.006397f
C269 output.n32 gnd 0.01428f
C270 output.n33 gnd 0.01428f
C271 output.n34 gnd 0.006397f
C272 output.n35 gnd 0.006041f
C273 output.n36 gnd 0.011243f
C274 output.n37 gnd 0.011243f
C275 output.n38 gnd 0.006041f
C276 output.n39 gnd 0.006397f
C277 output.n40 gnd 0.01428f
C278 output.n41 gnd 0.030913f
C279 output.n42 gnd 0.006397f
C280 output.n43 gnd 0.006041f
C281 output.n44 gnd 0.025987f
C282 output.n45 gnd 0.097665f
C283 output.n46 gnd 0.015803f
C284 output.n47 gnd 0.011243f
C285 output.n48 gnd 0.006041f
C286 output.n49 gnd 0.01428f
C287 output.n50 gnd 0.006397f
C288 output.n51 gnd 0.011243f
C289 output.n52 gnd 0.006041f
C290 output.n53 gnd 0.01428f
C291 output.n54 gnd 0.006397f
C292 output.n55 gnd 0.048111f
C293 output.t19 gnd 0.023274f
C294 output.n56 gnd 0.01071f
C295 output.n57 gnd 0.008435f
C296 output.n58 gnd 0.006041f
C297 output.n59 gnd 0.267512f
C298 output.n60 gnd 0.011243f
C299 output.n61 gnd 0.006041f
C300 output.n62 gnd 0.006397f
C301 output.n63 gnd 0.01428f
C302 output.n64 gnd 0.01428f
C303 output.n65 gnd 0.006397f
C304 output.n66 gnd 0.006041f
C305 output.n67 gnd 0.011243f
C306 output.n68 gnd 0.011243f
C307 output.n69 gnd 0.006041f
C308 output.n70 gnd 0.006397f
C309 output.n71 gnd 0.01428f
C310 output.n72 gnd 0.030913f
C311 output.n73 gnd 0.006397f
C312 output.n74 gnd 0.006041f
C313 output.n75 gnd 0.025987f
C314 output.n76 gnd 0.09306f
C315 output.n77 gnd 1.65264f
C316 output.n78 gnd 0.015803f
C317 output.n79 gnd 0.011243f
C318 output.n80 gnd 0.006041f
C319 output.n81 gnd 0.01428f
C320 output.n82 gnd 0.006397f
C321 output.n83 gnd 0.011243f
C322 output.n84 gnd 0.006041f
C323 output.n85 gnd 0.01428f
C324 output.n86 gnd 0.006397f
C325 output.n87 gnd 0.048111f
C326 output.t18 gnd 0.023274f
C327 output.n88 gnd 0.01071f
C328 output.n89 gnd 0.008435f
C329 output.n90 gnd 0.006041f
C330 output.n91 gnd 0.267512f
C331 output.n92 gnd 0.011243f
C332 output.n93 gnd 0.006041f
C333 output.n94 gnd 0.006397f
C334 output.n95 gnd 0.01428f
C335 output.n96 gnd 0.01428f
C336 output.n97 gnd 0.006397f
C337 output.n98 gnd 0.006041f
C338 output.n99 gnd 0.011243f
C339 output.n100 gnd 0.011243f
C340 output.n101 gnd 0.006041f
C341 output.n102 gnd 0.006397f
C342 output.n103 gnd 0.01428f
C343 output.n104 gnd 0.030913f
C344 output.n105 gnd 0.006397f
C345 output.n106 gnd 0.006041f
C346 output.n107 gnd 0.025987f
C347 output.n108 gnd 0.09306f
C348 output.n109 gnd 0.713089f
C349 output.n110 gnd 0.015803f
C350 output.n111 gnd 0.011243f
C351 output.n112 gnd 0.006041f
C352 output.n113 gnd 0.01428f
C353 output.n114 gnd 0.006397f
C354 output.n115 gnd 0.011243f
C355 output.n116 gnd 0.006041f
C356 output.n117 gnd 0.01428f
C357 output.n118 gnd 0.006397f
C358 output.n119 gnd 0.048111f
C359 output.t17 gnd 0.023274f
C360 output.n120 gnd 0.01071f
C361 output.n121 gnd 0.008435f
C362 output.n122 gnd 0.006041f
C363 output.n123 gnd 0.267512f
C364 output.n124 gnd 0.011243f
C365 output.n125 gnd 0.006041f
C366 output.n126 gnd 0.006397f
C367 output.n127 gnd 0.01428f
C368 output.n128 gnd 0.01428f
C369 output.n129 gnd 0.006397f
C370 output.n130 gnd 0.006041f
C371 output.n131 gnd 0.011243f
C372 output.n132 gnd 0.011243f
C373 output.n133 gnd 0.006041f
C374 output.n134 gnd 0.006397f
C375 output.n135 gnd 0.01428f
C376 output.n136 gnd 0.030913f
C377 output.n137 gnd 0.006397f
C378 output.n138 gnd 0.006041f
C379 output.n139 gnd 0.025987f
C380 output.n140 gnd 0.09306f
C381 output.n141 gnd 1.67353f
C382 minus.n0 gnd 0.032421f
C383 minus.n1 gnd 0.007357f
C384 minus.n2 gnd 0.032421f
C385 minus.n3 gnd 0.007357f
C386 minus.n4 gnd 0.032421f
C387 minus.n5 gnd 0.007357f
C388 minus.n6 gnd 0.032421f
C389 minus.n7 gnd 0.007357f
C390 minus.n8 gnd 0.032421f
C391 minus.n9 gnd 0.007357f
C392 minus.t8 gnd 0.47521f
C393 minus.t7 gnd 0.458565f
C394 minus.n10 gnd 0.210344f
C395 minus.n11 gnd 0.18879f
C396 minus.n12 gnd 0.139574f
C397 minus.n13 gnd 0.032421f
C398 minus.t11 gnd 0.458565f
C399 minus.n14 gnd 0.203709f
C400 minus.n15 gnd 0.007357f
C401 minus.t10 gnd 0.458565f
C402 minus.n16 gnd 0.203709f
C403 minus.n17 gnd 0.032421f
C404 minus.n18 gnd 0.032421f
C405 minus.n19 gnd 0.032421f
C406 minus.t12 gnd 0.458565f
C407 minus.n20 gnd 0.203709f
C408 minus.n21 gnd 0.007357f
C409 minus.t20 gnd 0.458565f
C410 minus.n22 gnd 0.203709f
C411 minus.n23 gnd 0.032421f
C412 minus.n24 gnd 0.032421f
C413 minus.n25 gnd 0.032421f
C414 minus.t18 gnd 0.458565f
C415 minus.n26 gnd 0.203709f
C416 minus.n27 gnd 0.007357f
C417 minus.t25 gnd 0.458565f
C418 minus.n28 gnd 0.203709f
C419 minus.n29 gnd 0.032421f
C420 minus.n30 gnd 0.032421f
C421 minus.n31 gnd 0.032421f
C422 minus.t24 gnd 0.458565f
C423 minus.n32 gnd 0.203709f
C424 minus.n33 gnd 0.007357f
C425 minus.t14 gnd 0.458565f
C426 minus.n34 gnd 0.203709f
C427 minus.n35 gnd 0.032421f
C428 minus.n36 gnd 0.032421f
C429 minus.n37 gnd 0.032421f
C430 minus.t22 gnd 0.458565f
C431 minus.n38 gnd 0.203709f
C432 minus.n39 gnd 0.007357f
C433 minus.t19 gnd 0.458565f
C434 minus.n40 gnd 0.204009f
C435 minus.n41 gnd 0.375467f
C436 minus.n42 gnd 0.032421f
C437 minus.t13 gnd 0.458565f
C438 minus.t15 gnd 0.458565f
C439 minus.n43 gnd 0.032421f
C440 minus.t5 gnd 0.458565f
C441 minus.n44 gnd 0.203709f
C442 minus.n45 gnd 0.032421f
C443 minus.t6 gnd 0.458565f
C444 minus.t26 gnd 0.458565f
C445 minus.n46 gnd 0.203709f
C446 minus.n47 gnd 0.032421f
C447 minus.t21 gnd 0.458565f
C448 minus.t23 gnd 0.458565f
C449 minus.n48 gnd 0.203709f
C450 minus.n49 gnd 0.032421f
C451 minus.t16 gnd 0.458565f
C452 minus.t17 gnd 0.458565f
C453 minus.n50 gnd 0.203709f
C454 minus.n51 gnd 0.032421f
C455 minus.t9 gnd 0.458565f
C456 minus.t27 gnd 0.458565f
C457 minus.n52 gnd 0.210344f
C458 minus.t28 gnd 0.47521f
C459 minus.n53 gnd 0.18879f
C460 minus.n54 gnd 0.139574f
C461 minus.n55 gnd 0.007357f
C462 minus.n56 gnd 0.203709f
C463 minus.n57 gnd 0.007357f
C464 minus.n58 gnd 0.032421f
C465 minus.n59 gnd 0.032421f
C466 minus.n60 gnd 0.032421f
C467 minus.n61 gnd 0.007357f
C468 minus.n62 gnd 0.203709f
C469 minus.n63 gnd 0.007357f
C470 minus.n64 gnd 0.032421f
C471 minus.n65 gnd 0.032421f
C472 minus.n66 gnd 0.032421f
C473 minus.n67 gnd 0.007357f
C474 minus.n68 gnd 0.203709f
C475 minus.n69 gnd 0.007357f
C476 minus.n70 gnd 0.032421f
C477 minus.n71 gnd 0.032421f
C478 minus.n72 gnd 0.032421f
C479 minus.n73 gnd 0.007357f
C480 minus.n74 gnd 0.203709f
C481 minus.n75 gnd 0.007357f
C482 minus.n76 gnd 0.032421f
C483 minus.n77 gnd 0.032421f
C484 minus.n78 gnd 0.032421f
C485 minus.n79 gnd 0.007357f
C486 minus.n80 gnd 0.203709f
C487 minus.n81 gnd 0.007357f
C488 minus.n82 gnd 0.204009f
C489 minus.n83 gnd 1.08613f
C490 minus.n84 gnd 1.61832f
C491 minus.t1 gnd 0.009994f
C492 minus.t0 gnd 0.009994f
C493 minus.n85 gnd 0.032864f
C494 minus.t4 gnd 0.009994f
C495 minus.t3 gnd 0.009994f
C496 minus.n86 gnd 0.032414f
C497 minus.n87 gnd 0.276636f
C498 minus.t2 gnd 0.055628f
C499 minus.n88 gnd 0.150958f
C500 minus.n89 gnd 1.94905f
C501 a_n2982_8322.t26 gnd 0.100195f
C502 a_n2982_8322.t5 gnd 20.7864f
C503 a_n2982_8322.t2 gnd 20.640598f
C504 a_n2982_8322.t4 gnd 20.640598f
C505 a_n2982_8322.t0 gnd 20.7864f
C506 a_n2982_8322.t3 gnd 20.640598f
C507 a_n2982_8322.t1 gnd 28.793001f
C508 a_n2982_8322.t35 gnd 0.938173f
C509 a_n2982_8322.t28 gnd 0.100195f
C510 a_n2982_8322.t24 gnd 0.100195f
C511 a_n2982_8322.n0 gnd 0.705774f
C512 a_n2982_8322.n1 gnd 0.7886f
C513 a_n2982_8322.t21 gnd 0.100195f
C514 a_n2982_8322.t37 gnd 0.100195f
C515 a_n2982_8322.n2 gnd 0.705774f
C516 a_n2982_8322.n3 gnd 0.400677f
C517 a_n2982_8322.t34 gnd 0.100195f
C518 a_n2982_8322.t22 gnd 0.100195f
C519 a_n2982_8322.n4 gnd 0.705774f
C520 a_n2982_8322.n5 gnd 0.400677f
C521 a_n2982_8322.t19 gnd 0.100195f
C522 a_n2982_8322.t18 gnd 0.100195f
C523 a_n2982_8322.n6 gnd 0.705774f
C524 a_n2982_8322.n7 gnd 0.400677f
C525 a_n2982_8322.t32 gnd 0.100195f
C526 a_n2982_8322.t31 gnd 0.100195f
C527 a_n2982_8322.n8 gnd 0.705774f
C528 a_n2982_8322.n9 gnd 0.400677f
C529 a_n2982_8322.t15 gnd 0.936307f
C530 a_n2982_8322.n10 gnd 1.11185f
C531 a_n2982_8322.n11 gnd 3.2687f
C532 a_n2982_8322.t9 gnd 0.938176f
C533 a_n2982_8322.t13 gnd 0.100195f
C534 a_n2982_8322.t12 gnd 0.100195f
C535 a_n2982_8322.n12 gnd 0.705774f
C536 a_n2982_8322.n13 gnd 0.788598f
C537 a_n2982_8322.t7 gnd 0.936307f
C538 a_n2982_8322.n14 gnd 0.396834f
C539 a_n2982_8322.t10 gnd 0.936307f
C540 a_n2982_8322.n15 gnd 0.396834f
C541 a_n2982_8322.t8 gnd 0.100195f
C542 a_n2982_8322.t6 gnd 0.100195f
C543 a_n2982_8322.n16 gnd 0.705774f
C544 a_n2982_8322.n17 gnd 0.400677f
C545 a_n2982_8322.t11 gnd 0.936307f
C546 a_n2982_8322.n18 gnd 1.47193f
C547 a_n2982_8322.n19 gnd 2.35218f
C548 a_n2982_8322.t14 gnd 0.936307f
C549 a_n2982_8322.n20 gnd 1.87205f
C550 a_n2982_8322.t27 gnd 0.100195f
C551 a_n2982_8322.t25 gnd 0.100195f
C552 a_n2982_8322.n21 gnd 0.705774f
C553 a_n2982_8322.n22 gnd 0.400677f
C554 a_n2982_8322.t30 gnd 0.100195f
C555 a_n2982_8322.t23 gnd 0.100195f
C556 a_n2982_8322.n23 gnd 0.705774f
C557 a_n2982_8322.n24 gnd 0.400677f
C558 a_n2982_8322.t17 gnd 0.100195f
C559 a_n2982_8322.t16 gnd 0.100195f
C560 a_n2982_8322.n25 gnd 0.705774f
C561 a_n2982_8322.n26 gnd 0.400677f
C562 a_n2982_8322.t20 gnd 0.938176f
C563 a_n2982_8322.t33 gnd 0.100195f
C564 a_n2982_8322.t29 gnd 0.100195f
C565 a_n2982_8322.n27 gnd 0.705774f
C566 a_n2982_8322.n28 gnd 0.788598f
C567 a_n2982_8322.n29 gnd 0.400675f
C568 a_n2982_8322.n30 gnd 0.705776f
C569 a_n2982_8322.t36 gnd 0.100195f
C570 a_n2804_13878.t29 gnd 0.194878f
C571 a_n2804_13878.t25 gnd 0.194878f
C572 a_n2804_13878.t31 gnd 0.194878f
C573 a_n2804_13878.n0 gnd 1.53703f
C574 a_n2804_13878.t8 gnd 0.194878f
C575 a_n2804_13878.t20 gnd 0.194878f
C576 a_n2804_13878.n1 gnd 1.5345f
C577 a_n2804_13878.n2 gnd 1.37932f
C578 a_n2804_13878.t12 gnd 0.194878f
C579 a_n2804_13878.t22 gnd 0.194878f
C580 a_n2804_13878.n3 gnd 1.53612f
C581 a_n2804_13878.t27 gnd 0.194878f
C582 a_n2804_13878.t17 gnd 0.194878f
C583 a_n2804_13878.n4 gnd 1.5345f
C584 a_n2804_13878.n5 gnd 2.14416f
C585 a_n2804_13878.t23 gnd 0.194878f
C586 a_n2804_13878.t16 gnd 0.194878f
C587 a_n2804_13878.n6 gnd 1.5345f
C588 a_n2804_13878.n7 gnd 1.04587f
C589 a_n2804_13878.t10 gnd 0.194878f
C590 a_n2804_13878.t13 gnd 0.194878f
C591 a_n2804_13878.n8 gnd 1.5345f
C592 a_n2804_13878.n9 gnd 1.04587f
C593 a_n2804_13878.t26 gnd 0.194878f
C594 a_n2804_13878.t11 gnd 0.194878f
C595 a_n2804_13878.n10 gnd 1.5345f
C596 a_n2804_13878.n11 gnd 1.04587f
C597 a_n2804_13878.t21 gnd 0.194878f
C598 a_n2804_13878.t9 gnd 0.194878f
C599 a_n2804_13878.n12 gnd 1.5345f
C600 a_n2804_13878.n13 gnd 4.90989f
C601 a_n2804_13878.t1 gnd 1.82474f
C602 a_n2804_13878.t4 gnd 0.194878f
C603 a_n2804_13878.t5 gnd 0.194878f
C604 a_n2804_13878.n14 gnd 1.37272f
C605 a_n2804_13878.n15 gnd 1.53381f
C606 a_n2804_13878.t0 gnd 1.8211f
C607 a_n2804_13878.n16 gnd 0.771835f
C608 a_n2804_13878.t3 gnd 1.8211f
C609 a_n2804_13878.n17 gnd 0.771835f
C610 a_n2804_13878.t6 gnd 0.194878f
C611 a_n2804_13878.t7 gnd 0.194878f
C612 a_n2804_13878.n18 gnd 1.37272f
C613 a_n2804_13878.n19 gnd 0.77931f
C614 a_n2804_13878.t2 gnd 1.8211f
C615 a_n2804_13878.n20 gnd 2.86287f
C616 a_n2804_13878.n21 gnd 3.75497f
C617 a_n2804_13878.t15 gnd 0.194878f
C618 a_n2804_13878.t24 gnd 0.194878f
C619 a_n2804_13878.n22 gnd 1.53449f
C620 a_n2804_13878.n23 gnd 2.50654f
C621 a_n2804_13878.t28 gnd 0.194878f
C622 a_n2804_13878.t14 gnd 0.194878f
C623 a_n2804_13878.n24 gnd 1.5345f
C624 a_n2804_13878.n25 gnd 0.679894f
C625 a_n2804_13878.t18 gnd 0.194878f
C626 a_n2804_13878.t19 gnd 0.194878f
C627 a_n2804_13878.n26 gnd 1.5345f
C628 a_n2804_13878.n27 gnd 0.679894f
C629 a_n2804_13878.n28 gnd 0.679892f
C630 a_n2804_13878.n29 gnd 1.5345f
C631 a_n2804_13878.t30 gnd 0.194878f
C632 vdd.t200 gnd 0.02966f
C633 vdd.t181 gnd 0.02966f
C634 vdd.n0 gnd 0.233929f
C635 vdd.t159 gnd 0.02966f
C636 vdd.t196 gnd 0.02966f
C637 vdd.n1 gnd 0.233543f
C638 vdd.n2 gnd 0.215371f
C639 vdd.t165 gnd 0.02966f
C640 vdd.t207 gnd 0.02966f
C641 vdd.n3 gnd 0.233543f
C642 vdd.n4 gnd 0.108921f
C643 vdd.t205 gnd 0.02966f
C644 vdd.t185 gnd 0.02966f
C645 vdd.n5 gnd 0.233543f
C646 vdd.n6 gnd 0.102202f
C647 vdd.t211 gnd 0.02966f
C648 vdd.t177 gnd 0.02966f
C649 vdd.n7 gnd 0.233929f
C650 vdd.t183 gnd 0.02966f
C651 vdd.t203 gnd 0.02966f
C652 vdd.n8 gnd 0.233543f
C653 vdd.n9 gnd 0.215371f
C654 vdd.t192 gnd 0.02966f
C655 vdd.t163 gnd 0.02966f
C656 vdd.n10 gnd 0.233543f
C657 vdd.n11 gnd 0.108921f
C658 vdd.t167 gnd 0.02966f
C659 vdd.t190 gnd 0.02966f
C660 vdd.n12 gnd 0.233543f
C661 vdd.n13 gnd 0.102202f
C662 vdd.n14 gnd 0.072255f
C663 vdd.t0 gnd 0.016478f
C664 vdd.t1 gnd 0.016478f
C665 vdd.n15 gnd 0.151668f
C666 vdd.t15 gnd 0.016478f
C667 vdd.t7 gnd 0.016478f
C668 vdd.n16 gnd 0.151225f
C669 vdd.n17 gnd 0.263178f
C670 vdd.t8 gnd 0.016478f
C671 vdd.t11 gnd 0.016478f
C672 vdd.n18 gnd 0.151225f
C673 vdd.n19 gnd 0.10888f
C674 vdd.t6 gnd 0.016478f
C675 vdd.t12 gnd 0.016478f
C676 vdd.n20 gnd 0.151668f
C677 vdd.t14 gnd 0.016478f
C678 vdd.t5 gnd 0.016478f
C679 vdd.n21 gnd 0.151225f
C680 vdd.n22 gnd 0.263178f
C681 vdd.t3 gnd 0.016478f
C682 vdd.t10 gnd 0.016478f
C683 vdd.n23 gnd 0.151225f
C684 vdd.n24 gnd 0.10888f
C685 vdd.t2 gnd 0.016478f
C686 vdd.t4 gnd 0.016478f
C687 vdd.n25 gnd 0.151225f
C688 vdd.t13 gnd 0.016478f
C689 vdd.t9 gnd 0.016478f
C690 vdd.n26 gnd 0.151225f
C691 vdd.n27 gnd 16.58f
C692 vdd.n28 gnd 6.49218f
C693 vdd.n29 gnd 0.004494f
C694 vdd.n30 gnd 0.00417f
C695 vdd.n31 gnd 0.002307f
C696 vdd.n32 gnd 0.005297f
C697 vdd.n33 gnd 0.002241f
C698 vdd.n34 gnd 0.002373f
C699 vdd.n35 gnd 0.00417f
C700 vdd.n36 gnd 0.002241f
C701 vdd.n37 gnd 0.005297f
C702 vdd.n38 gnd 0.002373f
C703 vdd.n39 gnd 0.00417f
C704 vdd.n40 gnd 0.002241f
C705 vdd.n41 gnd 0.003973f
C706 vdd.n42 gnd 0.003984f
C707 vdd.t127 gnd 0.01138f
C708 vdd.n43 gnd 0.025319f
C709 vdd.n44 gnd 0.131769f
C710 vdd.n45 gnd 0.002241f
C711 vdd.n46 gnd 0.002373f
C712 vdd.n47 gnd 0.005297f
C713 vdd.n48 gnd 0.005297f
C714 vdd.n49 gnd 0.002373f
C715 vdd.n50 gnd 0.002241f
C716 vdd.n51 gnd 0.00417f
C717 vdd.n52 gnd 0.00417f
C718 vdd.n53 gnd 0.002241f
C719 vdd.n54 gnd 0.002373f
C720 vdd.n55 gnd 0.005297f
C721 vdd.n56 gnd 0.005297f
C722 vdd.n57 gnd 0.002373f
C723 vdd.n58 gnd 0.002241f
C724 vdd.n59 gnd 0.00417f
C725 vdd.n60 gnd 0.00417f
C726 vdd.n61 gnd 0.002241f
C727 vdd.n62 gnd 0.002373f
C728 vdd.n63 gnd 0.005297f
C729 vdd.n64 gnd 0.005297f
C730 vdd.n65 gnd 0.012523f
C731 vdd.n66 gnd 0.002307f
C732 vdd.n67 gnd 0.002241f
C733 vdd.n68 gnd 0.010779f
C734 vdd.n69 gnd 0.007525f
C735 vdd.t118 gnd 0.026364f
C736 vdd.t148 gnd 0.026364f
C737 vdd.n70 gnd 0.181191f
C738 vdd.n71 gnd 0.142479f
C739 vdd.t103 gnd 0.026364f
C740 vdd.t140 gnd 0.026364f
C741 vdd.n72 gnd 0.181191f
C742 vdd.n73 gnd 0.11498f
C743 vdd.t108 gnd 0.026364f
C744 vdd.t144 gnd 0.026364f
C745 vdd.n74 gnd 0.181191f
C746 vdd.n75 gnd 0.11498f
C747 vdd.n76 gnd 0.004494f
C748 vdd.n77 gnd 0.00417f
C749 vdd.n78 gnd 0.002307f
C750 vdd.n79 gnd 0.005297f
C751 vdd.n80 gnd 0.002241f
C752 vdd.n81 gnd 0.002373f
C753 vdd.n82 gnd 0.00417f
C754 vdd.n83 gnd 0.002241f
C755 vdd.n84 gnd 0.005297f
C756 vdd.n85 gnd 0.002373f
C757 vdd.n86 gnd 0.00417f
C758 vdd.n87 gnd 0.002241f
C759 vdd.n88 gnd 0.003973f
C760 vdd.n89 gnd 0.003984f
C761 vdd.t122 gnd 0.01138f
C762 vdd.n90 gnd 0.025319f
C763 vdd.n91 gnd 0.131769f
C764 vdd.n92 gnd 0.002241f
C765 vdd.n93 gnd 0.002373f
C766 vdd.n94 gnd 0.005297f
C767 vdd.n95 gnd 0.005297f
C768 vdd.n96 gnd 0.002373f
C769 vdd.n97 gnd 0.002241f
C770 vdd.n98 gnd 0.00417f
C771 vdd.n99 gnd 0.00417f
C772 vdd.n100 gnd 0.002241f
C773 vdd.n101 gnd 0.002373f
C774 vdd.n102 gnd 0.005297f
C775 vdd.n103 gnd 0.005297f
C776 vdd.n104 gnd 0.002373f
C777 vdd.n105 gnd 0.002241f
C778 vdd.n106 gnd 0.00417f
C779 vdd.n107 gnd 0.00417f
C780 vdd.n108 gnd 0.002241f
C781 vdd.n109 gnd 0.002373f
C782 vdd.n110 gnd 0.005297f
C783 vdd.n111 gnd 0.005297f
C784 vdd.n112 gnd 0.012523f
C785 vdd.n113 gnd 0.002307f
C786 vdd.n114 gnd 0.002241f
C787 vdd.n115 gnd 0.010779f
C788 vdd.n116 gnd 0.007289f
C789 vdd.n117 gnd 0.085546f
C790 vdd.n118 gnd 0.004494f
C791 vdd.n119 gnd 0.00417f
C792 vdd.n120 gnd 0.002307f
C793 vdd.n121 gnd 0.005297f
C794 vdd.n122 gnd 0.002241f
C795 vdd.n123 gnd 0.002373f
C796 vdd.n124 gnd 0.00417f
C797 vdd.n125 gnd 0.002241f
C798 vdd.n126 gnd 0.005297f
C799 vdd.n127 gnd 0.002373f
C800 vdd.n128 gnd 0.00417f
C801 vdd.n129 gnd 0.002241f
C802 vdd.n130 gnd 0.003973f
C803 vdd.n131 gnd 0.003984f
C804 vdd.t150 gnd 0.01138f
C805 vdd.n132 gnd 0.025319f
C806 vdd.n133 gnd 0.131769f
C807 vdd.n134 gnd 0.002241f
C808 vdd.n135 gnd 0.002373f
C809 vdd.n136 gnd 0.005297f
C810 vdd.n137 gnd 0.005297f
C811 vdd.n138 gnd 0.002373f
C812 vdd.n139 gnd 0.002241f
C813 vdd.n140 gnd 0.00417f
C814 vdd.n141 gnd 0.00417f
C815 vdd.n142 gnd 0.002241f
C816 vdd.n143 gnd 0.002373f
C817 vdd.n144 gnd 0.005297f
C818 vdd.n145 gnd 0.005297f
C819 vdd.n146 gnd 0.002373f
C820 vdd.n147 gnd 0.002241f
C821 vdd.n148 gnd 0.00417f
C822 vdd.n149 gnd 0.00417f
C823 vdd.n150 gnd 0.002241f
C824 vdd.n151 gnd 0.002373f
C825 vdd.n152 gnd 0.005297f
C826 vdd.n153 gnd 0.005297f
C827 vdd.n154 gnd 0.012523f
C828 vdd.n155 gnd 0.002307f
C829 vdd.n156 gnd 0.002241f
C830 vdd.n157 gnd 0.010779f
C831 vdd.n158 gnd 0.007525f
C832 vdd.t151 gnd 0.026364f
C833 vdd.t101 gnd 0.026364f
C834 vdd.n159 gnd 0.181191f
C835 vdd.n160 gnd 0.142479f
C836 vdd.t143 gnd 0.026364f
C837 vdd.t147 gnd 0.026364f
C838 vdd.n161 gnd 0.181191f
C839 vdd.n162 gnd 0.11498f
C840 vdd.t99 gnd 0.026364f
C841 vdd.t125 gnd 0.026364f
C842 vdd.n163 gnd 0.181191f
C843 vdd.n164 gnd 0.11498f
C844 vdd.n165 gnd 0.004494f
C845 vdd.n166 gnd 0.00417f
C846 vdd.n167 gnd 0.002307f
C847 vdd.n168 gnd 0.005297f
C848 vdd.n169 gnd 0.002241f
C849 vdd.n170 gnd 0.002373f
C850 vdd.n171 gnd 0.00417f
C851 vdd.n172 gnd 0.002241f
C852 vdd.n173 gnd 0.005297f
C853 vdd.n174 gnd 0.002373f
C854 vdd.n175 gnd 0.00417f
C855 vdd.n176 gnd 0.002241f
C856 vdd.n177 gnd 0.003973f
C857 vdd.n178 gnd 0.003984f
C858 vdd.t142 gnd 0.01138f
C859 vdd.n179 gnd 0.025319f
C860 vdd.n180 gnd 0.131769f
C861 vdd.n181 gnd 0.002241f
C862 vdd.n182 gnd 0.002373f
C863 vdd.n183 gnd 0.005297f
C864 vdd.n184 gnd 0.005297f
C865 vdd.n185 gnd 0.002373f
C866 vdd.n186 gnd 0.002241f
C867 vdd.n187 gnd 0.00417f
C868 vdd.n188 gnd 0.00417f
C869 vdd.n189 gnd 0.002241f
C870 vdd.n190 gnd 0.002373f
C871 vdd.n191 gnd 0.005297f
C872 vdd.n192 gnd 0.005297f
C873 vdd.n193 gnd 0.002373f
C874 vdd.n194 gnd 0.002241f
C875 vdd.n195 gnd 0.00417f
C876 vdd.n196 gnd 0.00417f
C877 vdd.n197 gnd 0.002241f
C878 vdd.n198 gnd 0.002373f
C879 vdd.n199 gnd 0.005297f
C880 vdd.n200 gnd 0.005297f
C881 vdd.n201 gnd 0.012523f
C882 vdd.n202 gnd 0.002307f
C883 vdd.n203 gnd 0.002241f
C884 vdd.n204 gnd 0.010779f
C885 vdd.n205 gnd 0.007289f
C886 vdd.n206 gnd 0.050891f
C887 vdd.n207 gnd 0.183374f
C888 vdd.n208 gnd 0.004494f
C889 vdd.n209 gnd 0.00417f
C890 vdd.n210 gnd 0.002307f
C891 vdd.n211 gnd 0.005297f
C892 vdd.n212 gnd 0.002241f
C893 vdd.n213 gnd 0.002373f
C894 vdd.n214 gnd 0.00417f
C895 vdd.n215 gnd 0.002241f
C896 vdd.n216 gnd 0.005297f
C897 vdd.n217 gnd 0.002373f
C898 vdd.n218 gnd 0.00417f
C899 vdd.n219 gnd 0.002241f
C900 vdd.n220 gnd 0.003973f
C901 vdd.n221 gnd 0.003984f
C902 vdd.t153 gnd 0.01138f
C903 vdd.n222 gnd 0.025319f
C904 vdd.n223 gnd 0.131769f
C905 vdd.n224 gnd 0.002241f
C906 vdd.n225 gnd 0.002373f
C907 vdd.n226 gnd 0.005297f
C908 vdd.n227 gnd 0.005297f
C909 vdd.n228 gnd 0.002373f
C910 vdd.n229 gnd 0.002241f
C911 vdd.n230 gnd 0.00417f
C912 vdd.n231 gnd 0.00417f
C913 vdd.n232 gnd 0.002241f
C914 vdd.n233 gnd 0.002373f
C915 vdd.n234 gnd 0.005297f
C916 vdd.n235 gnd 0.005297f
C917 vdd.n236 gnd 0.002373f
C918 vdd.n237 gnd 0.002241f
C919 vdd.n238 gnd 0.00417f
C920 vdd.n239 gnd 0.00417f
C921 vdd.n240 gnd 0.002241f
C922 vdd.n241 gnd 0.002373f
C923 vdd.n242 gnd 0.005297f
C924 vdd.n243 gnd 0.005297f
C925 vdd.n244 gnd 0.012523f
C926 vdd.n245 gnd 0.002307f
C927 vdd.n246 gnd 0.002241f
C928 vdd.n247 gnd 0.010779f
C929 vdd.n248 gnd 0.007525f
C930 vdd.t154 gnd 0.026364f
C931 vdd.t116 gnd 0.026364f
C932 vdd.n249 gnd 0.181191f
C933 vdd.n250 gnd 0.142479f
C934 vdd.t146 gnd 0.026364f
C935 vdd.t152 gnd 0.026364f
C936 vdd.n251 gnd 0.181191f
C937 vdd.n252 gnd 0.11498f
C938 vdd.t109 gnd 0.026364f
C939 vdd.t135 gnd 0.026364f
C940 vdd.n253 gnd 0.181191f
C941 vdd.n254 gnd 0.11498f
C942 vdd.n255 gnd 0.004494f
C943 vdd.n256 gnd 0.00417f
C944 vdd.n257 gnd 0.002307f
C945 vdd.n258 gnd 0.005297f
C946 vdd.n259 gnd 0.002241f
C947 vdd.n260 gnd 0.002373f
C948 vdd.n261 gnd 0.00417f
C949 vdd.n262 gnd 0.002241f
C950 vdd.n263 gnd 0.005297f
C951 vdd.n264 gnd 0.002373f
C952 vdd.n265 gnd 0.00417f
C953 vdd.n266 gnd 0.002241f
C954 vdd.n267 gnd 0.003973f
C955 vdd.n268 gnd 0.003984f
C956 vdd.t145 gnd 0.01138f
C957 vdd.n269 gnd 0.025319f
C958 vdd.n270 gnd 0.131769f
C959 vdd.n271 gnd 0.002241f
C960 vdd.n272 gnd 0.002373f
C961 vdd.n273 gnd 0.005297f
C962 vdd.n274 gnd 0.005297f
C963 vdd.n275 gnd 0.002373f
C964 vdd.n276 gnd 0.002241f
C965 vdd.n277 gnd 0.00417f
C966 vdd.n278 gnd 0.00417f
C967 vdd.n279 gnd 0.002241f
C968 vdd.n280 gnd 0.002373f
C969 vdd.n281 gnd 0.005297f
C970 vdd.n282 gnd 0.005297f
C971 vdd.n283 gnd 0.002373f
C972 vdd.n284 gnd 0.002241f
C973 vdd.n285 gnd 0.00417f
C974 vdd.n286 gnd 0.00417f
C975 vdd.n287 gnd 0.002241f
C976 vdd.n288 gnd 0.002373f
C977 vdd.n289 gnd 0.005297f
C978 vdd.n290 gnd 0.005297f
C979 vdd.n291 gnd 0.012523f
C980 vdd.n292 gnd 0.002307f
C981 vdd.n293 gnd 0.002241f
C982 vdd.n294 gnd 0.010779f
C983 vdd.n295 gnd 0.007289f
C984 vdd.n296 gnd 0.050891f
C985 vdd.n297 gnd 0.198481f
C986 vdd.n298 gnd 0.006294f
C987 vdd.n299 gnd 0.008189f
C988 vdd.n300 gnd 0.006591f
C989 vdd.n301 gnd 0.006591f
C990 vdd.n302 gnd 0.008189f
C991 vdd.n303 gnd 0.008189f
C992 vdd.n304 gnd 0.598353f
C993 vdd.n305 gnd 0.008189f
C994 vdd.n306 gnd 0.008189f
C995 vdd.n307 gnd 0.008189f
C996 vdd.n308 gnd 0.648564f
C997 vdd.n309 gnd 0.008189f
C998 vdd.n310 gnd 0.008189f
C999 vdd.n311 gnd 0.008189f
C1000 vdd.n312 gnd 0.008189f
C1001 vdd.n313 gnd 0.006591f
C1002 vdd.n314 gnd 0.008189f
C1003 vdd.t124 gnd 0.418428f
C1004 vdd.n315 gnd 0.008189f
C1005 vdd.n316 gnd 0.008189f
C1006 vdd.n317 gnd 0.008189f
C1007 vdd.n318 gnd 0.836857f
C1008 vdd.n319 gnd 0.008189f
C1009 vdd.n320 gnd 0.008189f
C1010 vdd.n321 gnd 0.008189f
C1011 vdd.n322 gnd 0.008189f
C1012 vdd.n323 gnd 0.008189f
C1013 vdd.n324 gnd 0.006591f
C1014 vdd.n325 gnd 0.008189f
C1015 vdd.n326 gnd 0.008189f
C1016 vdd.n327 gnd 0.008189f
C1017 vdd.n328 gnd 0.019956f
C1018 vdd.n329 gnd 2.00009f
C1019 vdd.n330 gnd 0.020414f
C1020 vdd.n331 gnd 0.008189f
C1021 vdd.n332 gnd 0.008189f
C1022 vdd.n334 gnd 0.008189f
C1023 vdd.n335 gnd 0.008189f
C1024 vdd.n336 gnd 0.006591f
C1025 vdd.n337 gnd 0.006591f
C1026 vdd.n338 gnd 0.008189f
C1027 vdd.n339 gnd 0.008189f
C1028 vdd.n340 gnd 0.008189f
C1029 vdd.n341 gnd 0.008189f
C1030 vdd.n342 gnd 0.008189f
C1031 vdd.n343 gnd 0.008189f
C1032 vdd.n344 gnd 0.006591f
C1033 vdd.n346 gnd 0.008189f
C1034 vdd.n347 gnd 0.008189f
C1035 vdd.n348 gnd 0.008189f
C1036 vdd.n349 gnd 0.008189f
C1037 vdd.n350 gnd 0.008189f
C1038 vdd.n351 gnd 0.006591f
C1039 vdd.n353 gnd 0.008189f
C1040 vdd.n354 gnd 0.008189f
C1041 vdd.n355 gnd 0.008189f
C1042 vdd.n356 gnd 0.008189f
C1043 vdd.n357 gnd 0.008189f
C1044 vdd.n358 gnd 0.006591f
C1045 vdd.n360 gnd 0.008189f
C1046 vdd.n361 gnd 0.008189f
C1047 vdd.n362 gnd 0.008189f
C1048 vdd.n363 gnd 0.008189f
C1049 vdd.n364 gnd 0.005503f
C1050 vdd.t91 gnd 0.100744f
C1051 vdd.t90 gnd 0.107667f
C1052 vdd.t89 gnd 0.13157f
C1053 vdd.n365 gnd 0.168654f
C1054 vdd.n366 gnd 0.142359f
C1055 vdd.n368 gnd 0.008189f
C1056 vdd.n369 gnd 0.008189f
C1057 vdd.n370 gnd 0.006591f
C1058 vdd.n371 gnd 0.008189f
C1059 vdd.n373 gnd 0.008189f
C1060 vdd.n374 gnd 0.008189f
C1061 vdd.n375 gnd 0.008189f
C1062 vdd.n376 gnd 0.008189f
C1063 vdd.n377 gnd 0.006591f
C1064 vdd.n379 gnd 0.008189f
C1065 vdd.n380 gnd 0.008189f
C1066 vdd.n381 gnd 0.008189f
C1067 vdd.n382 gnd 0.008189f
C1068 vdd.n383 gnd 0.008189f
C1069 vdd.n384 gnd 0.006591f
C1070 vdd.n386 gnd 0.008189f
C1071 vdd.n387 gnd 0.008189f
C1072 vdd.n388 gnd 0.008189f
C1073 vdd.n389 gnd 0.008189f
C1074 vdd.n390 gnd 0.008189f
C1075 vdd.n391 gnd 0.006591f
C1076 vdd.n393 gnd 0.008189f
C1077 vdd.n394 gnd 0.008189f
C1078 vdd.n395 gnd 0.008189f
C1079 vdd.n396 gnd 0.008189f
C1080 vdd.n397 gnd 0.008189f
C1081 vdd.n398 gnd 0.006591f
C1082 vdd.n400 gnd 0.008189f
C1083 vdd.n401 gnd 0.008189f
C1084 vdd.n402 gnd 0.008189f
C1085 vdd.n403 gnd 0.008189f
C1086 vdd.n404 gnd 0.006525f
C1087 vdd.t88 gnd 0.100744f
C1088 vdd.t87 gnd 0.107667f
C1089 vdd.t86 gnd 0.13157f
C1090 vdd.n405 gnd 0.168654f
C1091 vdd.n406 gnd 0.142359f
C1092 vdd.n408 gnd 0.008189f
C1093 vdd.n409 gnd 0.008189f
C1094 vdd.n410 gnd 0.006591f
C1095 vdd.n411 gnd 0.008189f
C1096 vdd.n413 gnd 0.008189f
C1097 vdd.n414 gnd 0.008189f
C1098 vdd.n415 gnd 0.008189f
C1099 vdd.n416 gnd 0.008189f
C1100 vdd.n417 gnd 0.006591f
C1101 vdd.n419 gnd 0.008189f
C1102 vdd.n420 gnd 0.008189f
C1103 vdd.n421 gnd 0.008189f
C1104 vdd.n422 gnd 0.008189f
C1105 vdd.n423 gnd 0.008189f
C1106 vdd.n424 gnd 0.006591f
C1107 vdd.n426 gnd 0.008189f
C1108 vdd.n427 gnd 0.008189f
C1109 vdd.n428 gnd 0.008189f
C1110 vdd.n429 gnd 0.008189f
C1111 vdd.n430 gnd 0.008189f
C1112 vdd.n431 gnd 0.006591f
C1113 vdd.n433 gnd 0.008189f
C1114 vdd.n434 gnd 0.008189f
C1115 vdd.n435 gnd 0.008189f
C1116 vdd.n436 gnd 0.008189f
C1117 vdd.n437 gnd 0.008189f
C1118 vdd.n438 gnd 0.006591f
C1119 vdd.n440 gnd 0.008189f
C1120 vdd.n441 gnd 0.008189f
C1121 vdd.n442 gnd 0.008189f
C1122 vdd.n443 gnd 0.008189f
C1123 vdd.n444 gnd 0.008189f
C1124 vdd.n445 gnd 0.008189f
C1125 vdd.n446 gnd 0.006591f
C1126 vdd.n447 gnd 0.008189f
C1127 vdd.n448 gnd 0.008189f
C1128 vdd.n449 gnd 0.006591f
C1129 vdd.n450 gnd 0.008189f
C1130 vdd.n451 gnd 0.006591f
C1131 vdd.n452 gnd 0.008189f
C1132 vdd.n453 gnd 0.006591f
C1133 vdd.n454 gnd 0.008189f
C1134 vdd.n455 gnd 0.008189f
C1135 vdd.n456 gnd 0.456087f
C1136 vdd.t102 gnd 0.418428f
C1137 vdd.n457 gnd 0.008189f
C1138 vdd.n458 gnd 0.006591f
C1139 vdd.n459 gnd 0.008189f
C1140 vdd.n460 gnd 0.006591f
C1141 vdd.n461 gnd 0.008189f
C1142 vdd.t117 gnd 0.418428f
C1143 vdd.n462 gnd 0.008189f
C1144 vdd.n463 gnd 0.006591f
C1145 vdd.n464 gnd 0.008189f
C1146 vdd.n465 gnd 0.006591f
C1147 vdd.n466 gnd 0.008189f
C1148 vdd.t126 gnd 0.418428f
C1149 vdd.n467 gnd 0.523035f
C1150 vdd.n468 gnd 0.008189f
C1151 vdd.n469 gnd 0.006591f
C1152 vdd.n470 gnd 0.008189f
C1153 vdd.n471 gnd 0.006591f
C1154 vdd.n472 gnd 0.008189f
C1155 vdd.n473 gnd 0.836857f
C1156 vdd.n474 gnd 0.008189f
C1157 vdd.n475 gnd 0.006591f
C1158 vdd.n476 gnd 0.019956f
C1159 vdd.n477 gnd 0.005471f
C1160 vdd.n478 gnd 0.019956f
C1161 vdd.t35 gnd 0.418428f
C1162 vdd.n479 gnd 0.019956f
C1163 vdd.n480 gnd 0.005471f
C1164 vdd.n481 gnd 0.007042f
C1165 vdd.n482 gnd 0.006591f
C1166 vdd.n483 gnd 0.008189f
C1167 vdd.n484 gnd 9.883281f
C1168 vdd.n515 gnd 0.020414f
C1169 vdd.n516 gnd 1.15068f
C1170 vdd.n517 gnd 0.008189f
C1171 vdd.n518 gnd 0.006591f
C1172 vdd.n519 gnd 0.005241f
C1173 vdd.n520 gnd 0.034384f
C1174 vdd.n521 gnd 0.006591f
C1175 vdd.n522 gnd 0.008189f
C1176 vdd.n523 gnd 0.008189f
C1177 vdd.n524 gnd 0.008189f
C1178 vdd.n525 gnd 0.008189f
C1179 vdd.n526 gnd 0.008189f
C1180 vdd.n527 gnd 0.008189f
C1181 vdd.n528 gnd 0.008189f
C1182 vdd.n529 gnd 0.008189f
C1183 vdd.n530 gnd 0.008189f
C1184 vdd.n531 gnd 0.008189f
C1185 vdd.n532 gnd 0.008189f
C1186 vdd.n533 gnd 0.008189f
C1187 vdd.n534 gnd 0.008189f
C1188 vdd.n535 gnd 0.008189f
C1189 vdd.n536 gnd 0.005503f
C1190 vdd.n537 gnd 0.008189f
C1191 vdd.n538 gnd 0.008189f
C1192 vdd.n539 gnd 0.008189f
C1193 vdd.n540 gnd 0.008189f
C1194 vdd.n541 gnd 0.008189f
C1195 vdd.n542 gnd 0.008189f
C1196 vdd.n543 gnd 0.008189f
C1197 vdd.n544 gnd 0.008189f
C1198 vdd.n545 gnd 0.008189f
C1199 vdd.n546 gnd 0.008189f
C1200 vdd.n547 gnd 0.008189f
C1201 vdd.n548 gnd 0.008189f
C1202 vdd.n549 gnd 0.008189f
C1203 vdd.n550 gnd 0.008189f
C1204 vdd.n551 gnd 0.008189f
C1205 vdd.n552 gnd 0.008189f
C1206 vdd.n553 gnd 0.008189f
C1207 vdd.n554 gnd 0.008189f
C1208 vdd.n555 gnd 0.008189f
C1209 vdd.n556 gnd 0.006525f
C1210 vdd.t60 gnd 0.100744f
C1211 vdd.t61 gnd 0.107667f
C1212 vdd.t59 gnd 0.13157f
C1213 vdd.n557 gnd 0.168654f
C1214 vdd.n558 gnd 0.1417f
C1215 vdd.n559 gnd 0.008189f
C1216 vdd.n560 gnd 0.008189f
C1217 vdd.n561 gnd 0.008189f
C1218 vdd.n562 gnd 0.008189f
C1219 vdd.n563 gnd 0.008189f
C1220 vdd.n564 gnd 0.008189f
C1221 vdd.n565 gnd 0.008189f
C1222 vdd.n566 gnd 0.008189f
C1223 vdd.n567 gnd 0.008189f
C1224 vdd.n568 gnd 0.008189f
C1225 vdd.n569 gnd 0.008189f
C1226 vdd.n570 gnd 0.008189f
C1227 vdd.n571 gnd 0.008189f
C1228 vdd.n572 gnd 0.005241f
C1229 vdd.n575 gnd 0.005568f
C1230 vdd.n576 gnd 0.005568f
C1231 vdd.n577 gnd 0.005568f
C1232 vdd.n578 gnd 0.005568f
C1233 vdd.n579 gnd 0.005568f
C1234 vdd.n580 gnd 0.005568f
C1235 vdd.n582 gnd 0.005568f
C1236 vdd.n583 gnd 0.005568f
C1237 vdd.n585 gnd 0.005568f
C1238 vdd.n586 gnd 0.004053f
C1239 vdd.n588 gnd 0.005568f
C1240 vdd.t19 gnd 0.225018f
C1241 vdd.t18 gnd 0.230334f
C1242 vdd.t16 gnd 0.1469f
C1243 vdd.n589 gnd 0.079392f
C1244 vdd.n590 gnd 0.045033f
C1245 vdd.n591 gnd 0.007958f
C1246 vdd.n592 gnd 0.012644f
C1247 vdd.n594 gnd 0.005568f
C1248 vdd.n595 gnd 0.569063f
C1249 vdd.n596 gnd 0.011923f
C1250 vdd.n597 gnd 0.011923f
C1251 vdd.n598 gnd 0.005568f
C1252 vdd.n599 gnd 0.012644f
C1253 vdd.n600 gnd 0.005568f
C1254 vdd.n601 gnd 0.005568f
C1255 vdd.n602 gnd 0.005568f
C1256 vdd.n603 gnd 0.005568f
C1257 vdd.n604 gnd 0.005568f
C1258 vdd.n606 gnd 0.005568f
C1259 vdd.n607 gnd 0.005568f
C1260 vdd.n609 gnd 0.005568f
C1261 vdd.n610 gnd 0.005568f
C1262 vdd.n612 gnd 0.005568f
C1263 vdd.n613 gnd 0.005568f
C1264 vdd.n615 gnd 0.005568f
C1265 vdd.n616 gnd 0.005568f
C1266 vdd.n618 gnd 0.005568f
C1267 vdd.n619 gnd 0.005568f
C1268 vdd.n621 gnd 0.005568f
C1269 vdd.t33 gnd 0.225018f
C1270 vdd.t32 gnd 0.230334f
C1271 vdd.t31 gnd 0.1469f
C1272 vdd.n622 gnd 0.079392f
C1273 vdd.n623 gnd 0.045033f
C1274 vdd.n624 gnd 0.005568f
C1275 vdd.n626 gnd 0.005568f
C1276 vdd.n627 gnd 0.005568f
C1277 vdd.t17 gnd 0.284531f
C1278 vdd.n628 gnd 0.005568f
C1279 vdd.n629 gnd 0.005568f
C1280 vdd.n630 gnd 0.005568f
C1281 vdd.n631 gnd 0.005568f
C1282 vdd.n632 gnd 0.005568f
C1283 vdd.n633 gnd 0.569063f
C1284 vdd.n634 gnd 0.005568f
C1285 vdd.n635 gnd 0.005568f
C1286 vdd.n636 gnd 0.447718f
C1287 vdd.n637 gnd 0.005568f
C1288 vdd.n638 gnd 0.005568f
C1289 vdd.n639 gnd 0.005568f
C1290 vdd.n640 gnd 0.005568f
C1291 vdd.n641 gnd 0.569063f
C1292 vdd.n642 gnd 0.005568f
C1293 vdd.n643 gnd 0.005568f
C1294 vdd.n644 gnd 0.005568f
C1295 vdd.n645 gnd 0.005568f
C1296 vdd.n646 gnd 0.005568f
C1297 vdd.t174 gnd 0.284531f
C1298 vdd.n647 gnd 0.005568f
C1299 vdd.n648 gnd 0.005568f
C1300 vdd.n649 gnd 0.005568f
C1301 vdd.n650 gnd 0.005568f
C1302 vdd.n651 gnd 0.005568f
C1303 vdd.t187 gnd 0.284531f
C1304 vdd.n652 gnd 0.005568f
C1305 vdd.n653 gnd 0.005568f
C1306 vdd.n654 gnd 0.548141f
C1307 vdd.n655 gnd 0.005568f
C1308 vdd.n656 gnd 0.005568f
C1309 vdd.n657 gnd 0.005568f
C1310 vdd.t186 gnd 0.284531f
C1311 vdd.n658 gnd 0.005568f
C1312 vdd.n659 gnd 0.005568f
C1313 vdd.n660 gnd 0.422613f
C1314 vdd.n661 gnd 0.005568f
C1315 vdd.n662 gnd 0.005568f
C1316 vdd.n663 gnd 0.005568f
C1317 vdd.n664 gnd 0.397507f
C1318 vdd.n665 gnd 0.005568f
C1319 vdd.n666 gnd 0.005568f
C1320 vdd.n667 gnd 0.297084f
C1321 vdd.n668 gnd 0.005568f
C1322 vdd.n669 gnd 0.005568f
C1323 vdd.n670 gnd 0.005568f
C1324 vdd.n671 gnd 0.523035f
C1325 vdd.n672 gnd 0.005568f
C1326 vdd.n673 gnd 0.005568f
C1327 vdd.t193 gnd 0.284531f
C1328 vdd.n674 gnd 0.005568f
C1329 vdd.n675 gnd 0.005568f
C1330 vdd.n676 gnd 0.005568f
C1331 vdd.n677 gnd 0.569063f
C1332 vdd.n678 gnd 0.005568f
C1333 vdd.n679 gnd 0.005568f
C1334 vdd.t194 gnd 0.284531f
C1335 vdd.n680 gnd 0.005568f
C1336 vdd.n681 gnd 0.005568f
C1337 vdd.n682 gnd 0.005568f
C1338 vdd.t168 gnd 0.284531f
C1339 vdd.n683 gnd 0.005568f
C1340 vdd.n684 gnd 0.005568f
C1341 vdd.n685 gnd 0.005568f
C1342 vdd.t40 gnd 0.230334f
C1343 vdd.t38 gnd 0.1469f
C1344 vdd.t41 gnd 0.230334f
C1345 vdd.n686 gnd 0.129457f
C1346 vdd.n687 gnd 0.016131f
C1347 vdd.n688 gnd 0.005568f
C1348 vdd.t39 gnd 0.20503f
C1349 vdd.n689 gnd 0.005568f
C1350 vdd.n690 gnd 0.005568f
C1351 vdd.n691 gnd 0.489561f
C1352 vdd.n692 gnd 0.005568f
C1353 vdd.n693 gnd 0.005568f
C1354 vdd.n694 gnd 0.005568f
C1355 vdd.n695 gnd 0.330558f
C1356 vdd.n696 gnd 0.005568f
C1357 vdd.n697 gnd 0.005568f
C1358 vdd.t169 gnd 0.11716f
C1359 vdd.n698 gnd 0.364033f
C1360 vdd.n699 gnd 0.005568f
C1361 vdd.n700 gnd 0.005568f
C1362 vdd.n701 gnd 0.005568f
C1363 vdd.n702 gnd 0.456087f
C1364 vdd.n703 gnd 0.005568f
C1365 vdd.n704 gnd 0.005568f
C1366 vdd.t178 gnd 0.284531f
C1367 vdd.n705 gnd 0.005568f
C1368 vdd.n706 gnd 0.005568f
C1369 vdd.n707 gnd 0.005568f
C1370 vdd.t176 gnd 0.284531f
C1371 vdd.n708 gnd 0.005568f
C1372 vdd.n709 gnd 0.005568f
C1373 vdd.t197 gnd 0.284531f
C1374 vdd.n710 gnd 0.005568f
C1375 vdd.n711 gnd 0.005568f
C1376 vdd.n712 gnd 0.005568f
C1377 vdd.t156 gnd 0.192477f
C1378 vdd.n713 gnd 0.005568f
C1379 vdd.n714 gnd 0.005568f
C1380 vdd.n715 gnd 0.502114f
C1381 vdd.n716 gnd 0.005568f
C1382 vdd.n717 gnd 0.005568f
C1383 vdd.n718 gnd 0.005568f
C1384 vdd.t198 gnd 0.284531f
C1385 vdd.n719 gnd 0.005568f
C1386 vdd.n720 gnd 0.005568f
C1387 vdd.t210 gnd 0.271978f
C1388 vdd.n721 gnd 0.376586f
C1389 vdd.n722 gnd 0.005568f
C1390 vdd.n723 gnd 0.005568f
C1391 vdd.n724 gnd 0.005568f
C1392 vdd.t160 gnd 0.284531f
C1393 vdd.n725 gnd 0.005568f
C1394 vdd.n726 gnd 0.005568f
C1395 vdd.t202 gnd 0.284531f
C1396 vdd.n727 gnd 0.005568f
C1397 vdd.n728 gnd 0.005568f
C1398 vdd.n729 gnd 0.005568f
C1399 vdd.n730 gnd 0.569063f
C1400 vdd.n731 gnd 0.005568f
C1401 vdd.n732 gnd 0.005568f
C1402 vdd.t182 gnd 0.284531f
C1403 vdd.n733 gnd 0.005568f
C1404 vdd.n734 gnd 0.005568f
C1405 vdd.n735 gnd 0.005568f
C1406 vdd.n736 gnd 0.393323f
C1407 vdd.n737 gnd 0.005568f
C1408 vdd.n738 gnd 0.005568f
C1409 vdd.n739 gnd 0.005568f
C1410 vdd.n740 gnd 0.005568f
C1411 vdd.n741 gnd 0.005568f
C1412 vdd.t73 gnd 0.284531f
C1413 vdd.n742 gnd 0.005568f
C1414 vdd.n743 gnd 0.005568f
C1415 vdd.t162 gnd 0.284531f
C1416 vdd.n744 gnd 0.005568f
C1417 vdd.n745 gnd 0.011923f
C1418 vdd.n746 gnd 0.011923f
C1419 vdd.n747 gnd 0.64438f
C1420 vdd.n748 gnd 0.005568f
C1421 vdd.n749 gnd 0.005568f
C1422 vdd.t191 gnd 0.284531f
C1423 vdd.n750 gnd 0.011923f
C1424 vdd.n751 gnd 0.005568f
C1425 vdd.n752 gnd 0.005568f
C1426 vdd.t204 gnd 0.485377f
C1427 vdd.n770 gnd 0.012644f
C1428 vdd.n788 gnd 0.011923f
C1429 vdd.n789 gnd 0.005568f
C1430 vdd.n790 gnd 0.011923f
C1431 vdd.t85 gnd 0.225018f
C1432 vdd.t84 gnd 0.230334f
C1433 vdd.t83 gnd 0.1469f
C1434 vdd.n791 gnd 0.079392f
C1435 vdd.n792 gnd 0.045033f
C1436 vdd.n793 gnd 0.012644f
C1437 vdd.n794 gnd 0.005568f
C1438 vdd.n795 gnd 0.334743f
C1439 vdd.n796 gnd 0.011923f
C1440 vdd.n797 gnd 0.005568f
C1441 vdd.n798 gnd 0.012644f
C1442 vdd.n799 gnd 0.005568f
C1443 vdd.t68 gnd 0.225018f
C1444 vdd.t67 gnd 0.230334f
C1445 vdd.t65 gnd 0.1469f
C1446 vdd.n800 gnd 0.079392f
C1447 vdd.n801 gnd 0.045033f
C1448 vdd.n802 gnd 0.007958f
C1449 vdd.n803 gnd 0.005568f
C1450 vdd.n804 gnd 0.005568f
C1451 vdd.t66 gnd 0.284531f
C1452 vdd.n805 gnd 0.005568f
C1453 vdd.t206 gnd 0.284531f
C1454 vdd.n806 gnd 0.005568f
C1455 vdd.n807 gnd 0.005568f
C1456 vdd.n808 gnd 0.005568f
C1457 vdd.n809 gnd 0.005568f
C1458 vdd.n810 gnd 0.005568f
C1459 vdd.n811 gnd 0.569063f
C1460 vdd.n812 gnd 0.005568f
C1461 vdd.n813 gnd 0.005568f
C1462 vdd.t164 gnd 0.284531f
C1463 vdd.n814 gnd 0.005568f
C1464 vdd.n815 gnd 0.005568f
C1465 vdd.n816 gnd 0.005568f
C1466 vdd.n817 gnd 0.005568f
C1467 vdd.n818 gnd 0.41006f
C1468 vdd.n819 gnd 0.005568f
C1469 vdd.n820 gnd 0.005568f
C1470 vdd.n821 gnd 0.005568f
C1471 vdd.n822 gnd 0.005568f
C1472 vdd.n823 gnd 0.005568f
C1473 vdd.t157 gnd 0.284531f
C1474 vdd.n824 gnd 0.005568f
C1475 vdd.n825 gnd 0.005568f
C1476 vdd.t195 gnd 0.284531f
C1477 vdd.n826 gnd 0.005568f
C1478 vdd.n827 gnd 0.005568f
C1479 vdd.n828 gnd 0.005568f
C1480 vdd.t179 gnd 0.284531f
C1481 vdd.n829 gnd 0.005568f
C1482 vdd.n830 gnd 0.005568f
C1483 vdd.t158 gnd 0.284531f
C1484 vdd.n831 gnd 0.005568f
C1485 vdd.n832 gnd 0.005568f
C1486 vdd.n833 gnd 0.005568f
C1487 vdd.t180 gnd 0.271978f
C1488 vdd.n834 gnd 0.005568f
C1489 vdd.n835 gnd 0.005568f
C1490 vdd.n836 gnd 0.422613f
C1491 vdd.n837 gnd 0.005568f
C1492 vdd.n838 gnd 0.005568f
C1493 vdd.n839 gnd 0.005568f
C1494 vdd.t199 gnd 0.284531f
C1495 vdd.n840 gnd 0.005568f
C1496 vdd.n841 gnd 0.005568f
C1497 vdd.t171 gnd 0.192477f
C1498 vdd.n842 gnd 0.297084f
C1499 vdd.n843 gnd 0.005568f
C1500 vdd.n844 gnd 0.005568f
C1501 vdd.n845 gnd 0.005568f
C1502 vdd.n846 gnd 0.523035f
C1503 vdd.n847 gnd 0.005568f
C1504 vdd.n848 gnd 0.005568f
C1505 vdd.t208 gnd 0.284531f
C1506 vdd.n849 gnd 0.005568f
C1507 vdd.n850 gnd 0.005568f
C1508 vdd.n851 gnd 0.005568f
C1509 vdd.n852 gnd 0.569063f
C1510 vdd.n853 gnd 0.005568f
C1511 vdd.n854 gnd 0.005568f
C1512 vdd.t175 gnd 0.284531f
C1513 vdd.n855 gnd 0.005568f
C1514 vdd.n856 gnd 0.005568f
C1515 vdd.n857 gnd 0.005568f
C1516 vdd.t170 gnd 0.11716f
C1517 vdd.n858 gnd 0.005568f
C1518 vdd.n859 gnd 0.005568f
C1519 vdd.n860 gnd 0.005568f
C1520 vdd.t78 gnd 0.230334f
C1521 vdd.t76 gnd 0.1469f
C1522 vdd.t79 gnd 0.230334f
C1523 vdd.n861 gnd 0.129457f
C1524 vdd.n862 gnd 0.005568f
C1525 vdd.n863 gnd 0.005568f
C1526 vdd.t188 gnd 0.284531f
C1527 vdd.n864 gnd 0.005568f
C1528 vdd.n865 gnd 0.005568f
C1529 vdd.t77 gnd 0.20503f
C1530 vdd.n866 gnd 0.451903f
C1531 vdd.n867 gnd 0.005568f
C1532 vdd.n868 gnd 0.005568f
C1533 vdd.n869 gnd 0.005568f
C1534 vdd.n870 gnd 0.330558f
C1535 vdd.n871 gnd 0.005568f
C1536 vdd.n872 gnd 0.005568f
C1537 vdd.n873 gnd 0.364033f
C1538 vdd.n874 gnd 0.005568f
C1539 vdd.n875 gnd 0.005568f
C1540 vdd.n876 gnd 0.005568f
C1541 vdd.n877 gnd 0.456087f
C1542 vdd.n878 gnd 0.005568f
C1543 vdd.n879 gnd 0.005568f
C1544 vdd.t172 gnd 0.284531f
C1545 vdd.n880 gnd 0.005568f
C1546 vdd.n881 gnd 0.005568f
C1547 vdd.n882 gnd 0.005568f
C1548 vdd.n883 gnd 0.569063f
C1549 vdd.n884 gnd 0.005568f
C1550 vdd.n885 gnd 0.005568f
C1551 vdd.t173 gnd 0.284531f
C1552 vdd.n886 gnd 0.005568f
C1553 vdd.n887 gnd 0.005568f
C1554 vdd.n888 gnd 0.005568f
C1555 vdd.t209 gnd 0.284531f
C1556 vdd.n889 gnd 0.005568f
C1557 vdd.n890 gnd 0.005568f
C1558 vdd.n891 gnd 0.005568f
C1559 vdd.n892 gnd 0.005568f
C1560 vdd.n893 gnd 0.005568f
C1561 vdd.t201 gnd 0.284531f
C1562 vdd.n894 gnd 0.005568f
C1563 vdd.n895 gnd 0.005568f
C1564 vdd.n896 gnd 0.55651f
C1565 vdd.n897 gnd 0.005568f
C1566 vdd.n898 gnd 0.005568f
C1567 vdd.n899 gnd 0.005568f
C1568 vdd.t161 gnd 0.284531f
C1569 vdd.n900 gnd 0.005568f
C1570 vdd.n901 gnd 0.005568f
C1571 vdd.n902 gnd 0.430981f
C1572 vdd.n903 gnd 0.005568f
C1573 vdd.n904 gnd 0.005568f
C1574 vdd.n905 gnd 0.005568f
C1575 vdd.n906 gnd 0.569063f
C1576 vdd.n907 gnd 0.005568f
C1577 vdd.n908 gnd 0.005568f
C1578 vdd.n909 gnd 0.305453f
C1579 vdd.n910 gnd 0.005568f
C1580 vdd.n911 gnd 0.005568f
C1581 vdd.n912 gnd 0.005568f
C1582 vdd.n913 gnd 0.569063f
C1583 vdd.n914 gnd 0.005568f
C1584 vdd.n915 gnd 0.005568f
C1585 vdd.n916 gnd 0.005568f
C1586 vdd.n917 gnd 0.005568f
C1587 vdd.n918 gnd 0.005568f
C1588 vdd.t21 gnd 0.284531f
C1589 vdd.n919 gnd 0.005568f
C1590 vdd.n920 gnd 0.005568f
C1591 vdd.n921 gnd 0.005568f
C1592 vdd.n922 gnd 0.011923f
C1593 vdd.n923 gnd 0.011923f
C1594 vdd.n924 gnd 0.769908f
C1595 vdd.n925 gnd 0.005568f
C1596 vdd.n926 gnd 0.005568f
C1597 vdd.n927 gnd 0.405876f
C1598 vdd.n928 gnd 0.011923f
C1599 vdd.n929 gnd 0.005568f
C1600 vdd.n930 gnd 0.005568f
C1601 vdd.n931 gnd 10.2348f
C1602 vdd.n965 gnd 0.012644f
C1603 vdd.n966 gnd 0.005568f
C1604 vdd.n967 gnd 0.005568f
C1605 vdd.n968 gnd 0.005241f
C1606 vdd.n971 gnd 0.020414f
C1607 vdd.n972 gnd 0.005471f
C1608 vdd.n973 gnd 0.006591f
C1609 vdd.n975 gnd 0.008189f
C1610 vdd.n976 gnd 0.008189f
C1611 vdd.n977 gnd 0.006591f
C1612 vdd.n979 gnd 0.008189f
C1613 vdd.n980 gnd 0.008189f
C1614 vdd.n981 gnd 0.008189f
C1615 vdd.n982 gnd 0.008189f
C1616 vdd.n983 gnd 0.008189f
C1617 vdd.n984 gnd 0.006591f
C1618 vdd.n986 gnd 0.008189f
C1619 vdd.n987 gnd 0.008189f
C1620 vdd.n988 gnd 0.008189f
C1621 vdd.n989 gnd 0.008189f
C1622 vdd.n990 gnd 0.008189f
C1623 vdd.n991 gnd 0.006591f
C1624 vdd.n993 gnd 0.008189f
C1625 vdd.n994 gnd 0.008189f
C1626 vdd.n995 gnd 0.008189f
C1627 vdd.n996 gnd 0.008189f
C1628 vdd.n997 gnd 0.005503f
C1629 vdd.t30 gnd 0.100744f
C1630 vdd.t29 gnd 0.107667f
C1631 vdd.t28 gnd 0.13157f
C1632 vdd.n998 gnd 0.168654f
C1633 vdd.n999 gnd 0.1417f
C1634 vdd.n1001 gnd 0.008189f
C1635 vdd.n1002 gnd 0.008189f
C1636 vdd.n1003 gnd 0.006591f
C1637 vdd.n1004 gnd 0.008189f
C1638 vdd.n1006 gnd 0.008189f
C1639 vdd.n1007 gnd 0.008189f
C1640 vdd.n1008 gnd 0.008189f
C1641 vdd.n1009 gnd 0.008189f
C1642 vdd.n1010 gnd 0.006591f
C1643 vdd.n1012 gnd 0.008189f
C1644 vdd.n1013 gnd 0.008189f
C1645 vdd.n1014 gnd 0.008189f
C1646 vdd.n1015 gnd 0.008189f
C1647 vdd.n1016 gnd 0.008189f
C1648 vdd.n1017 gnd 0.006591f
C1649 vdd.n1019 gnd 0.008189f
C1650 vdd.n1020 gnd 0.008189f
C1651 vdd.n1021 gnd 0.008189f
C1652 vdd.n1022 gnd 0.008189f
C1653 vdd.n1023 gnd 0.008189f
C1654 vdd.n1024 gnd 0.006591f
C1655 vdd.n1026 gnd 0.008189f
C1656 vdd.n1027 gnd 0.008189f
C1657 vdd.n1028 gnd 0.008189f
C1658 vdd.n1029 gnd 0.008189f
C1659 vdd.n1030 gnd 0.008189f
C1660 vdd.n1031 gnd 0.006591f
C1661 vdd.n1033 gnd 0.008189f
C1662 vdd.n1034 gnd 0.008189f
C1663 vdd.n1035 gnd 0.008189f
C1664 vdd.n1036 gnd 0.008189f
C1665 vdd.n1037 gnd 0.006525f
C1666 vdd.t27 gnd 0.100744f
C1667 vdd.t26 gnd 0.107667f
C1668 vdd.t24 gnd 0.13157f
C1669 vdd.n1038 gnd 0.168654f
C1670 vdd.n1039 gnd 0.1417f
C1671 vdd.n1041 gnd 0.008189f
C1672 vdd.n1042 gnd 0.008189f
C1673 vdd.n1043 gnd 0.006591f
C1674 vdd.n1044 gnd 0.008189f
C1675 vdd.n1046 gnd 0.008189f
C1676 vdd.n1047 gnd 0.008189f
C1677 vdd.n1048 gnd 0.008189f
C1678 vdd.n1049 gnd 0.008189f
C1679 vdd.n1050 gnd 0.006591f
C1680 vdd.n1052 gnd 0.008189f
C1681 vdd.n1053 gnd 0.008189f
C1682 vdd.n1054 gnd 0.008189f
C1683 vdd.n1055 gnd 0.008189f
C1684 vdd.n1056 gnd 0.008189f
C1685 vdd.n1057 gnd 0.006591f
C1686 vdd.n1059 gnd 0.008189f
C1687 vdd.n1060 gnd 0.008189f
C1688 vdd.n1061 gnd 0.008189f
C1689 vdd.n1062 gnd 0.008189f
C1690 vdd.n1063 gnd 0.008189f
C1691 vdd.n1064 gnd 0.006591f
C1692 vdd.n1066 gnd 0.008189f
C1693 vdd.n1067 gnd 0.008189f
C1694 vdd.n1068 gnd 0.005241f
C1695 vdd.n1069 gnd 0.006591f
C1696 vdd.n1070 gnd 0.012644f
C1697 vdd.n1071 gnd 0.012644f
C1698 vdd.n1072 gnd 0.005568f
C1699 vdd.n1073 gnd 0.005568f
C1700 vdd.n1074 gnd 0.005568f
C1701 vdd.n1075 gnd 0.005568f
C1702 vdd.n1076 gnd 0.005568f
C1703 vdd.n1077 gnd 0.005568f
C1704 vdd.n1078 gnd 0.005568f
C1705 vdd.n1079 gnd 0.005568f
C1706 vdd.n1080 gnd 0.005568f
C1707 vdd.n1081 gnd 0.005568f
C1708 vdd.n1082 gnd 0.005568f
C1709 vdd.n1083 gnd 0.005568f
C1710 vdd.n1084 gnd 0.005568f
C1711 vdd.n1085 gnd 0.005568f
C1712 vdd.n1086 gnd 0.005568f
C1713 vdd.n1087 gnd 0.005568f
C1714 vdd.n1088 gnd 0.005568f
C1715 vdd.n1089 gnd 0.005568f
C1716 vdd.n1090 gnd 0.005568f
C1717 vdd.n1091 gnd 0.005568f
C1718 vdd.n1092 gnd 0.005568f
C1719 vdd.n1093 gnd 0.005568f
C1720 vdd.n1094 gnd 0.005568f
C1721 vdd.n1095 gnd 0.005568f
C1722 vdd.n1096 gnd 0.005568f
C1723 vdd.n1097 gnd 0.005568f
C1724 vdd.n1098 gnd 0.005568f
C1725 vdd.n1099 gnd 0.005568f
C1726 vdd.n1100 gnd 0.005568f
C1727 vdd.n1101 gnd 0.005568f
C1728 vdd.n1102 gnd 0.005568f
C1729 vdd.n1103 gnd 0.005568f
C1730 vdd.n1104 gnd 0.005568f
C1731 vdd.t22 gnd 0.225018f
C1732 vdd.t23 gnd 0.230334f
C1733 vdd.t20 gnd 0.1469f
C1734 vdd.n1105 gnd 0.079392f
C1735 vdd.n1106 gnd 0.045033f
C1736 vdd.n1107 gnd 0.007958f
C1737 vdd.n1108 gnd 0.005568f
C1738 vdd.t63 gnd 0.225018f
C1739 vdd.t64 gnd 0.230334f
C1740 vdd.t62 gnd 0.1469f
C1741 vdd.n1109 gnd 0.079392f
C1742 vdd.n1110 gnd 0.045033f
C1743 vdd.n1111 gnd 0.005568f
C1744 vdd.n1112 gnd 0.005568f
C1745 vdd.n1113 gnd 0.005568f
C1746 vdd.n1114 gnd 0.005568f
C1747 vdd.n1115 gnd 0.005568f
C1748 vdd.n1116 gnd 0.005568f
C1749 vdd.n1117 gnd 0.005568f
C1750 vdd.n1118 gnd 0.005568f
C1751 vdd.n1119 gnd 0.005568f
C1752 vdd.n1120 gnd 0.005568f
C1753 vdd.n1121 gnd 0.005568f
C1754 vdd.n1122 gnd 0.005568f
C1755 vdd.n1123 gnd 0.005568f
C1756 vdd.n1124 gnd 0.005568f
C1757 vdd.n1125 gnd 0.005568f
C1758 vdd.n1126 gnd 0.005568f
C1759 vdd.n1127 gnd 0.005568f
C1760 vdd.n1128 gnd 0.005568f
C1761 vdd.n1129 gnd 0.005568f
C1762 vdd.n1130 gnd 0.005568f
C1763 vdd.n1131 gnd 0.005568f
C1764 vdd.n1132 gnd 0.005568f
C1765 vdd.n1133 gnd 0.005568f
C1766 vdd.n1134 gnd 0.005568f
C1767 vdd.n1135 gnd 0.005568f
C1768 vdd.n1136 gnd 0.005568f
C1769 vdd.n1137 gnd 0.004053f
C1770 vdd.n1138 gnd 0.007958f
C1771 vdd.n1139 gnd 0.004299f
C1772 vdd.n1140 gnd 0.005568f
C1773 vdd.n1141 gnd 0.005568f
C1774 vdd.n1142 gnd 0.005568f
C1775 vdd.n1143 gnd 0.012644f
C1776 vdd.n1144 gnd 0.012644f
C1777 vdd.n1145 gnd 0.011923f
C1778 vdd.n1146 gnd 0.011923f
C1779 vdd.n1147 gnd 0.005568f
C1780 vdd.n1148 gnd 0.005568f
C1781 vdd.n1149 gnd 0.005568f
C1782 vdd.n1150 gnd 0.005568f
C1783 vdd.n1151 gnd 0.005568f
C1784 vdd.n1152 gnd 0.005568f
C1785 vdd.n1153 gnd 0.005568f
C1786 vdd.n1154 gnd 0.005568f
C1787 vdd.n1155 gnd 0.005568f
C1788 vdd.n1156 gnd 0.005568f
C1789 vdd.n1157 gnd 0.005568f
C1790 vdd.n1158 gnd 0.005568f
C1791 vdd.n1159 gnd 0.005568f
C1792 vdd.n1160 gnd 0.005568f
C1793 vdd.n1161 gnd 0.005568f
C1794 vdd.n1162 gnd 0.005568f
C1795 vdd.n1163 gnd 0.005568f
C1796 vdd.n1164 gnd 0.005568f
C1797 vdd.n1165 gnd 0.005568f
C1798 vdd.n1166 gnd 0.005568f
C1799 vdd.n1167 gnd 0.005568f
C1800 vdd.n1168 gnd 0.005568f
C1801 vdd.n1169 gnd 0.005568f
C1802 vdd.n1170 gnd 0.005568f
C1803 vdd.n1171 gnd 0.005568f
C1804 vdd.n1172 gnd 0.005568f
C1805 vdd.n1173 gnd 0.005568f
C1806 vdd.n1174 gnd 0.005568f
C1807 vdd.n1175 gnd 0.005568f
C1808 vdd.n1176 gnd 0.005568f
C1809 vdd.n1177 gnd 0.005568f
C1810 vdd.n1178 gnd 0.005568f
C1811 vdd.n1179 gnd 0.005568f
C1812 vdd.n1180 gnd 0.005568f
C1813 vdd.n1181 gnd 0.005568f
C1814 vdd.n1182 gnd 0.005568f
C1815 vdd.n1183 gnd 0.005568f
C1816 vdd.n1184 gnd 0.005568f
C1817 vdd.n1185 gnd 0.005568f
C1818 vdd.n1186 gnd 0.005568f
C1819 vdd.n1187 gnd 0.005568f
C1820 vdd.n1188 gnd 0.005568f
C1821 vdd.n1189 gnd 0.338927f
C1822 vdd.n1190 gnd 0.005568f
C1823 vdd.n1191 gnd 0.005568f
C1824 vdd.n1192 gnd 0.005568f
C1825 vdd.n1193 gnd 0.005568f
C1826 vdd.n1194 gnd 0.005568f
C1827 vdd.n1195 gnd 0.005568f
C1828 vdd.n1196 gnd 0.005568f
C1829 vdd.n1197 gnd 0.005568f
C1830 vdd.n1198 gnd 0.005568f
C1831 vdd.n1199 gnd 0.005568f
C1832 vdd.n1200 gnd 0.005568f
C1833 vdd.n1201 gnd 0.005568f
C1834 vdd.n1202 gnd 0.005568f
C1835 vdd.n1203 gnd 0.005568f
C1836 vdd.n1204 gnd 0.005568f
C1837 vdd.n1205 gnd 0.005568f
C1838 vdd.n1206 gnd 0.005568f
C1839 vdd.n1207 gnd 0.005568f
C1840 vdd.n1208 gnd 0.005568f
C1841 vdd.n1209 gnd 0.005568f
C1842 vdd.n1210 gnd 0.005568f
C1843 vdd.n1211 gnd 0.005568f
C1844 vdd.n1212 gnd 0.005568f
C1845 vdd.n1213 gnd 0.005568f
C1846 vdd.n1214 gnd 0.005568f
C1847 vdd.n1215 gnd 0.514667f
C1848 vdd.n1216 gnd 0.005568f
C1849 vdd.n1217 gnd 0.005568f
C1850 vdd.n1218 gnd 0.005568f
C1851 vdd.n1219 gnd 0.005568f
C1852 vdd.n1220 gnd 0.005568f
C1853 vdd.n1221 gnd 0.005568f
C1854 vdd.n1222 gnd 0.005568f
C1855 vdd.n1223 gnd 0.005568f
C1856 vdd.n1224 gnd 0.005568f
C1857 vdd.n1225 gnd 0.005568f
C1858 vdd.n1226 gnd 0.005568f
C1859 vdd.n1227 gnd 0.179924f
C1860 vdd.n1228 gnd 0.005568f
C1861 vdd.n1229 gnd 0.005568f
C1862 vdd.n1230 gnd 0.005568f
C1863 vdd.n1231 gnd 0.005568f
C1864 vdd.n1232 gnd 0.005568f
C1865 vdd.n1233 gnd 0.005568f
C1866 vdd.n1234 gnd 0.005568f
C1867 vdd.n1235 gnd 0.005568f
C1868 vdd.n1236 gnd 0.005568f
C1869 vdd.n1237 gnd 0.005568f
C1870 vdd.n1238 gnd 0.005568f
C1871 vdd.n1239 gnd 0.005568f
C1872 vdd.n1240 gnd 0.005568f
C1873 vdd.n1241 gnd 0.005568f
C1874 vdd.n1242 gnd 0.005568f
C1875 vdd.n1243 gnd 0.005568f
C1876 vdd.n1244 gnd 0.005568f
C1877 vdd.n1245 gnd 0.005568f
C1878 vdd.n1246 gnd 0.005568f
C1879 vdd.n1247 gnd 0.005568f
C1880 vdd.n1248 gnd 0.005568f
C1881 vdd.n1249 gnd 0.005568f
C1882 vdd.n1250 gnd 0.005568f
C1883 vdd.n1251 gnd 0.005568f
C1884 vdd.n1252 gnd 0.005568f
C1885 vdd.n1253 gnd 0.005568f
C1886 vdd.n1254 gnd 0.005568f
C1887 vdd.n1255 gnd 0.005568f
C1888 vdd.n1256 gnd 0.005568f
C1889 vdd.n1257 gnd 0.005568f
C1890 vdd.n1258 gnd 0.005568f
C1891 vdd.n1259 gnd 0.005568f
C1892 vdd.n1260 gnd 0.005568f
C1893 vdd.n1261 gnd 0.005568f
C1894 vdd.n1262 gnd 0.005568f
C1895 vdd.n1263 gnd 0.005568f
C1896 vdd.n1264 gnd 0.005568f
C1897 vdd.n1265 gnd 0.005568f
C1898 vdd.n1266 gnd 0.005568f
C1899 vdd.n1267 gnd 0.005568f
C1900 vdd.n1268 gnd 0.005568f
C1901 vdd.n1269 gnd 0.005568f
C1902 vdd.n1270 gnd 0.011923f
C1903 vdd.n1271 gnd 0.011923f
C1904 vdd.n1272 gnd 0.012644f
C1905 vdd.n1273 gnd 0.005568f
C1906 vdd.n1274 gnd 0.005568f
C1907 vdd.n1275 gnd 0.004299f
C1908 vdd.n1276 gnd 0.005568f
C1909 vdd.n1277 gnd 0.005568f
C1910 vdd.n1278 gnd 0.004053f
C1911 vdd.n1279 gnd 0.005568f
C1912 vdd.n1280 gnd 0.005568f
C1913 vdd.n1281 gnd 0.005568f
C1914 vdd.n1282 gnd 0.005568f
C1915 vdd.n1283 gnd 0.005568f
C1916 vdd.n1284 gnd 0.005568f
C1917 vdd.n1285 gnd 0.005568f
C1918 vdd.n1286 gnd 0.005568f
C1919 vdd.n1287 gnd 0.005568f
C1920 vdd.n1288 gnd 0.005568f
C1921 vdd.n1289 gnd 0.005568f
C1922 vdd.n1290 gnd 0.005568f
C1923 vdd.n1291 gnd 0.005568f
C1924 vdd.n1292 gnd 0.005568f
C1925 vdd.n1293 gnd 0.005568f
C1926 vdd.n1294 gnd 0.005568f
C1927 vdd.n1295 gnd 0.005568f
C1928 vdd.n1296 gnd 0.005568f
C1929 vdd.n1297 gnd 0.005568f
C1930 vdd.n1298 gnd 0.005568f
C1931 vdd.n1299 gnd 0.005568f
C1932 vdd.n1300 gnd 0.005568f
C1933 vdd.n1301 gnd 0.005568f
C1934 vdd.n1302 gnd 0.005568f
C1935 vdd.n1303 gnd 0.005568f
C1936 vdd.n1304 gnd 0.005568f
C1937 vdd.n1305 gnd 0.037512f
C1938 vdd.n1307 gnd 0.020414f
C1939 vdd.n1308 gnd 0.006591f
C1940 vdd.n1310 gnd 0.008189f
C1941 vdd.n1311 gnd 0.006591f
C1942 vdd.n1312 gnd 0.008189f
C1943 vdd.n1314 gnd 0.008189f
C1944 vdd.n1315 gnd 0.008189f
C1945 vdd.n1317 gnd 0.008189f
C1946 vdd.n1318 gnd 0.005471f
C1947 vdd.t25 gnd 0.418428f
C1948 vdd.n1319 gnd 0.008189f
C1949 vdd.n1320 gnd 0.020414f
C1950 vdd.n1321 gnd 0.006591f
C1951 vdd.n1322 gnd 0.008189f
C1952 vdd.n1323 gnd 0.006591f
C1953 vdd.n1324 gnd 0.008189f
C1954 vdd.n1325 gnd 0.836857f
C1955 vdd.n1326 gnd 0.008189f
C1956 vdd.n1327 gnd 0.006591f
C1957 vdd.n1328 gnd 0.006591f
C1958 vdd.n1329 gnd 0.008189f
C1959 vdd.n1330 gnd 0.006591f
C1960 vdd.n1331 gnd 0.008189f
C1961 vdd.t114 gnd 0.418428f
C1962 vdd.n1332 gnd 0.008189f
C1963 vdd.n1333 gnd 0.006591f
C1964 vdd.n1334 gnd 0.008189f
C1965 vdd.n1335 gnd 0.006591f
C1966 vdd.n1336 gnd 0.008189f
C1967 vdd.t130 gnd 0.418428f
C1968 vdd.n1337 gnd 0.008189f
C1969 vdd.n1338 gnd 0.006591f
C1970 vdd.n1339 gnd 0.008189f
C1971 vdd.n1340 gnd 0.006591f
C1972 vdd.n1341 gnd 0.008189f
C1973 vdd.n1342 gnd 0.656933f
C1974 vdd.n1343 gnd 0.694591f
C1975 vdd.t132 gnd 0.418428f
C1976 vdd.n1344 gnd 0.008189f
C1977 vdd.n1345 gnd 0.006591f
C1978 vdd.n1346 gnd 0.004494f
C1979 vdd.n1347 gnd 0.00417f
C1980 vdd.n1348 gnd 0.002307f
C1981 vdd.n1349 gnd 0.005297f
C1982 vdd.n1350 gnd 0.002241f
C1983 vdd.n1351 gnd 0.002373f
C1984 vdd.n1352 gnd 0.00417f
C1985 vdd.n1353 gnd 0.002241f
C1986 vdd.n1354 gnd 0.005297f
C1987 vdd.n1355 gnd 0.002373f
C1988 vdd.n1356 gnd 0.00417f
C1989 vdd.n1357 gnd 0.002241f
C1990 vdd.n1358 gnd 0.003973f
C1991 vdd.n1359 gnd 0.003984f
C1992 vdd.t128 gnd 0.01138f
C1993 vdd.n1360 gnd 0.025319f
C1994 vdd.n1361 gnd 0.131769f
C1995 vdd.n1362 gnd 0.002241f
C1996 vdd.n1363 gnd 0.002373f
C1997 vdd.n1364 gnd 0.005297f
C1998 vdd.n1365 gnd 0.005297f
C1999 vdd.n1366 gnd 0.002373f
C2000 vdd.n1367 gnd 0.002241f
C2001 vdd.n1368 gnd 0.00417f
C2002 vdd.n1369 gnd 0.00417f
C2003 vdd.n1370 gnd 0.002241f
C2004 vdd.n1371 gnd 0.002373f
C2005 vdd.n1372 gnd 0.005297f
C2006 vdd.n1373 gnd 0.005297f
C2007 vdd.n1374 gnd 0.002373f
C2008 vdd.n1375 gnd 0.002241f
C2009 vdd.n1376 gnd 0.00417f
C2010 vdd.n1377 gnd 0.00417f
C2011 vdd.n1378 gnd 0.002241f
C2012 vdd.n1379 gnd 0.002373f
C2013 vdd.n1380 gnd 0.005297f
C2014 vdd.n1381 gnd 0.005297f
C2015 vdd.n1382 gnd 0.012523f
C2016 vdd.n1383 gnd 0.002307f
C2017 vdd.n1384 gnd 0.002241f
C2018 vdd.n1385 gnd 0.010779f
C2019 vdd.n1386 gnd 0.007525f
C2020 vdd.t149 gnd 0.026364f
C2021 vdd.t155 gnd 0.026364f
C2022 vdd.n1387 gnd 0.181191f
C2023 vdd.n1388 gnd 0.142479f
C2024 vdd.t141 gnd 0.026364f
C2025 vdd.t104 gnd 0.026364f
C2026 vdd.n1389 gnd 0.181191f
C2027 vdd.n1390 gnd 0.11498f
C2028 vdd.t134 gnd 0.026364f
C2029 vdd.t113 gnd 0.026364f
C2030 vdd.n1391 gnd 0.181191f
C2031 vdd.n1392 gnd 0.11498f
C2032 vdd.n1393 gnd 0.004494f
C2033 vdd.n1394 gnd 0.00417f
C2034 vdd.n1395 gnd 0.002307f
C2035 vdd.n1396 gnd 0.005297f
C2036 vdd.n1397 gnd 0.002241f
C2037 vdd.n1398 gnd 0.002373f
C2038 vdd.n1399 gnd 0.00417f
C2039 vdd.n1400 gnd 0.002241f
C2040 vdd.n1401 gnd 0.005297f
C2041 vdd.n1402 gnd 0.002373f
C2042 vdd.n1403 gnd 0.00417f
C2043 vdd.n1404 gnd 0.002241f
C2044 vdd.n1405 gnd 0.003973f
C2045 vdd.n1406 gnd 0.003984f
C2046 vdd.t123 gnd 0.01138f
C2047 vdd.n1407 gnd 0.025319f
C2048 vdd.n1408 gnd 0.131769f
C2049 vdd.n1409 gnd 0.002241f
C2050 vdd.n1410 gnd 0.002373f
C2051 vdd.n1411 gnd 0.005297f
C2052 vdd.n1412 gnd 0.005297f
C2053 vdd.n1413 gnd 0.002373f
C2054 vdd.n1414 gnd 0.002241f
C2055 vdd.n1415 gnd 0.00417f
C2056 vdd.n1416 gnd 0.00417f
C2057 vdd.n1417 gnd 0.002241f
C2058 vdd.n1418 gnd 0.002373f
C2059 vdd.n1419 gnd 0.005297f
C2060 vdd.n1420 gnd 0.005297f
C2061 vdd.n1421 gnd 0.002373f
C2062 vdd.n1422 gnd 0.002241f
C2063 vdd.n1423 gnd 0.00417f
C2064 vdd.n1424 gnd 0.00417f
C2065 vdd.n1425 gnd 0.002241f
C2066 vdd.n1426 gnd 0.002373f
C2067 vdd.n1427 gnd 0.005297f
C2068 vdd.n1428 gnd 0.005297f
C2069 vdd.n1429 gnd 0.012523f
C2070 vdd.n1430 gnd 0.002307f
C2071 vdd.n1431 gnd 0.002241f
C2072 vdd.n1432 gnd 0.010779f
C2073 vdd.n1433 gnd 0.007289f
C2074 vdd.n1434 gnd 0.085546f
C2075 vdd.n1435 gnd 0.004494f
C2076 vdd.n1436 gnd 0.00417f
C2077 vdd.n1437 gnd 0.002307f
C2078 vdd.n1438 gnd 0.005297f
C2079 vdd.n1439 gnd 0.002241f
C2080 vdd.n1440 gnd 0.002373f
C2081 vdd.n1441 gnd 0.00417f
C2082 vdd.n1442 gnd 0.002241f
C2083 vdd.n1443 gnd 0.005297f
C2084 vdd.n1444 gnd 0.002373f
C2085 vdd.n1445 gnd 0.00417f
C2086 vdd.n1446 gnd 0.002241f
C2087 vdd.n1447 gnd 0.003973f
C2088 vdd.n1448 gnd 0.003984f
C2089 vdd.t115 gnd 0.01138f
C2090 vdd.n1449 gnd 0.025319f
C2091 vdd.n1450 gnd 0.131769f
C2092 vdd.n1451 gnd 0.002241f
C2093 vdd.n1452 gnd 0.002373f
C2094 vdd.n1453 gnd 0.005297f
C2095 vdd.n1454 gnd 0.005297f
C2096 vdd.n1455 gnd 0.002373f
C2097 vdd.n1456 gnd 0.002241f
C2098 vdd.n1457 gnd 0.00417f
C2099 vdd.n1458 gnd 0.00417f
C2100 vdd.n1459 gnd 0.002241f
C2101 vdd.n1460 gnd 0.002373f
C2102 vdd.n1461 gnd 0.005297f
C2103 vdd.n1462 gnd 0.005297f
C2104 vdd.n1463 gnd 0.002373f
C2105 vdd.n1464 gnd 0.002241f
C2106 vdd.n1465 gnd 0.00417f
C2107 vdd.n1466 gnd 0.00417f
C2108 vdd.n1467 gnd 0.002241f
C2109 vdd.n1468 gnd 0.002373f
C2110 vdd.n1469 gnd 0.005297f
C2111 vdd.n1470 gnd 0.005297f
C2112 vdd.n1471 gnd 0.012523f
C2113 vdd.n1472 gnd 0.002307f
C2114 vdd.n1473 gnd 0.002241f
C2115 vdd.n1474 gnd 0.010779f
C2116 vdd.n1475 gnd 0.007525f
C2117 vdd.t133 gnd 0.026364f
C2118 vdd.t131 gnd 0.026364f
C2119 vdd.n1476 gnd 0.181191f
C2120 vdd.n1477 gnd 0.142479f
C2121 vdd.t111 gnd 0.026364f
C2122 vdd.t97 gnd 0.026364f
C2123 vdd.n1478 gnd 0.181191f
C2124 vdd.n1479 gnd 0.11498f
C2125 vdd.t93 gnd 0.026364f
C2126 vdd.t129 gnd 0.026364f
C2127 vdd.n1480 gnd 0.181191f
C2128 vdd.n1481 gnd 0.11498f
C2129 vdd.n1482 gnd 0.004494f
C2130 vdd.n1483 gnd 0.00417f
C2131 vdd.n1484 gnd 0.002307f
C2132 vdd.n1485 gnd 0.005297f
C2133 vdd.n1486 gnd 0.002241f
C2134 vdd.n1487 gnd 0.002373f
C2135 vdd.n1488 gnd 0.00417f
C2136 vdd.n1489 gnd 0.002241f
C2137 vdd.n1490 gnd 0.005297f
C2138 vdd.n1491 gnd 0.002373f
C2139 vdd.n1492 gnd 0.00417f
C2140 vdd.n1493 gnd 0.002241f
C2141 vdd.n1494 gnd 0.003973f
C2142 vdd.n1495 gnd 0.003984f
C2143 vdd.t95 gnd 0.01138f
C2144 vdd.n1496 gnd 0.025319f
C2145 vdd.n1497 gnd 0.131769f
C2146 vdd.n1498 gnd 0.002241f
C2147 vdd.n1499 gnd 0.002373f
C2148 vdd.n1500 gnd 0.005297f
C2149 vdd.n1501 gnd 0.005297f
C2150 vdd.n1502 gnd 0.002373f
C2151 vdd.n1503 gnd 0.002241f
C2152 vdd.n1504 gnd 0.00417f
C2153 vdd.n1505 gnd 0.00417f
C2154 vdd.n1506 gnd 0.002241f
C2155 vdd.n1507 gnd 0.002373f
C2156 vdd.n1508 gnd 0.005297f
C2157 vdd.n1509 gnd 0.005297f
C2158 vdd.n1510 gnd 0.002373f
C2159 vdd.n1511 gnd 0.002241f
C2160 vdd.n1512 gnd 0.00417f
C2161 vdd.n1513 gnd 0.00417f
C2162 vdd.n1514 gnd 0.002241f
C2163 vdd.n1515 gnd 0.002373f
C2164 vdd.n1516 gnd 0.005297f
C2165 vdd.n1517 gnd 0.005297f
C2166 vdd.n1518 gnd 0.012523f
C2167 vdd.n1519 gnd 0.002307f
C2168 vdd.n1520 gnd 0.002241f
C2169 vdd.n1521 gnd 0.010779f
C2170 vdd.n1522 gnd 0.007289f
C2171 vdd.n1523 gnd 0.050891f
C2172 vdd.n1524 gnd 0.183374f
C2173 vdd.n1525 gnd 0.004494f
C2174 vdd.n1526 gnd 0.00417f
C2175 vdd.n1527 gnd 0.002307f
C2176 vdd.n1528 gnd 0.005297f
C2177 vdd.n1529 gnd 0.002241f
C2178 vdd.n1530 gnd 0.002373f
C2179 vdd.n1531 gnd 0.00417f
C2180 vdd.n1532 gnd 0.002241f
C2181 vdd.n1533 gnd 0.005297f
C2182 vdd.n1534 gnd 0.002373f
C2183 vdd.n1535 gnd 0.00417f
C2184 vdd.n1536 gnd 0.002241f
C2185 vdd.n1537 gnd 0.003973f
C2186 vdd.n1538 gnd 0.003984f
C2187 vdd.t120 gnd 0.01138f
C2188 vdd.n1539 gnd 0.025319f
C2189 vdd.n1540 gnd 0.131769f
C2190 vdd.n1541 gnd 0.002241f
C2191 vdd.n1542 gnd 0.002373f
C2192 vdd.n1543 gnd 0.005297f
C2193 vdd.n1544 gnd 0.005297f
C2194 vdd.n1545 gnd 0.002373f
C2195 vdd.n1546 gnd 0.002241f
C2196 vdd.n1547 gnd 0.00417f
C2197 vdd.n1548 gnd 0.00417f
C2198 vdd.n1549 gnd 0.002241f
C2199 vdd.n1550 gnd 0.002373f
C2200 vdd.n1551 gnd 0.005297f
C2201 vdd.n1552 gnd 0.005297f
C2202 vdd.n1553 gnd 0.002373f
C2203 vdd.n1554 gnd 0.002241f
C2204 vdd.n1555 gnd 0.00417f
C2205 vdd.n1556 gnd 0.00417f
C2206 vdd.n1557 gnd 0.002241f
C2207 vdd.n1558 gnd 0.002373f
C2208 vdd.n1559 gnd 0.005297f
C2209 vdd.n1560 gnd 0.005297f
C2210 vdd.n1561 gnd 0.012523f
C2211 vdd.n1562 gnd 0.002307f
C2212 vdd.n1563 gnd 0.002241f
C2213 vdd.n1564 gnd 0.010779f
C2214 vdd.n1565 gnd 0.007525f
C2215 vdd.t138 gnd 0.026364f
C2216 vdd.t137 gnd 0.026364f
C2217 vdd.n1566 gnd 0.181191f
C2218 vdd.n1567 gnd 0.142479f
C2219 vdd.t119 gnd 0.026364f
C2220 vdd.t107 gnd 0.026364f
C2221 vdd.n1568 gnd 0.181191f
C2222 vdd.n1569 gnd 0.11498f
C2223 vdd.t105 gnd 0.026364f
C2224 vdd.t136 gnd 0.026364f
C2225 vdd.n1570 gnd 0.181191f
C2226 vdd.n1571 gnd 0.11498f
C2227 vdd.n1572 gnd 0.004494f
C2228 vdd.n1573 gnd 0.00417f
C2229 vdd.n1574 gnd 0.002307f
C2230 vdd.n1575 gnd 0.005297f
C2231 vdd.n1576 gnd 0.002241f
C2232 vdd.n1577 gnd 0.002373f
C2233 vdd.n1578 gnd 0.00417f
C2234 vdd.n1579 gnd 0.002241f
C2235 vdd.n1580 gnd 0.005297f
C2236 vdd.n1581 gnd 0.002373f
C2237 vdd.n1582 gnd 0.00417f
C2238 vdd.n1583 gnd 0.002241f
C2239 vdd.n1584 gnd 0.003973f
C2240 vdd.n1585 gnd 0.003984f
C2241 vdd.t106 gnd 0.01138f
C2242 vdd.n1586 gnd 0.025319f
C2243 vdd.n1587 gnd 0.131769f
C2244 vdd.n1588 gnd 0.002241f
C2245 vdd.n1589 gnd 0.002373f
C2246 vdd.n1590 gnd 0.005297f
C2247 vdd.n1591 gnd 0.005297f
C2248 vdd.n1592 gnd 0.002373f
C2249 vdd.n1593 gnd 0.002241f
C2250 vdd.n1594 gnd 0.00417f
C2251 vdd.n1595 gnd 0.00417f
C2252 vdd.n1596 gnd 0.002241f
C2253 vdd.n1597 gnd 0.002373f
C2254 vdd.n1598 gnd 0.005297f
C2255 vdd.n1599 gnd 0.005297f
C2256 vdd.n1600 gnd 0.002373f
C2257 vdd.n1601 gnd 0.002241f
C2258 vdd.n1602 gnd 0.00417f
C2259 vdd.n1603 gnd 0.00417f
C2260 vdd.n1604 gnd 0.002241f
C2261 vdd.n1605 gnd 0.002373f
C2262 vdd.n1606 gnd 0.005297f
C2263 vdd.n1607 gnd 0.005297f
C2264 vdd.n1608 gnd 0.012523f
C2265 vdd.n1609 gnd 0.002307f
C2266 vdd.n1610 gnd 0.002241f
C2267 vdd.n1611 gnd 0.010779f
C2268 vdd.n1612 gnd 0.007289f
C2269 vdd.n1613 gnd 0.050891f
C2270 vdd.n1614 gnd 0.198481f
C2271 vdd.n1615 gnd 1.96474f
C2272 vdd.n1616 gnd 0.483007f
C2273 vdd.n1617 gnd 0.006591f
C2274 vdd.n1618 gnd 0.008189f
C2275 vdd.n1619 gnd 0.514667f
C2276 vdd.n1620 gnd 0.008189f
C2277 vdd.n1621 gnd 0.006591f
C2278 vdd.n1622 gnd 0.008189f
C2279 vdd.n1623 gnd 0.006591f
C2280 vdd.n1624 gnd 0.008189f
C2281 vdd.t112 gnd 0.418428f
C2282 vdd.t110 gnd 0.418428f
C2283 vdd.n1625 gnd 0.008189f
C2284 vdd.n1626 gnd 0.006591f
C2285 vdd.n1627 gnd 0.008189f
C2286 vdd.n1628 gnd 0.006591f
C2287 vdd.n1629 gnd 0.008189f
C2288 vdd.t92 gnd 0.418428f
C2289 vdd.n1630 gnd 0.008189f
C2290 vdd.n1631 gnd 0.006591f
C2291 vdd.n1632 gnd 0.008189f
C2292 vdd.n1633 gnd 0.006591f
C2293 vdd.n1634 gnd 0.008189f
C2294 vdd.t94 gnd 0.418428f
C2295 vdd.n1635 gnd 0.606721f
C2296 vdd.n1636 gnd 0.008189f
C2297 vdd.n1637 gnd 0.006591f
C2298 vdd.n1638 gnd 0.008189f
C2299 vdd.n1639 gnd 0.006591f
C2300 vdd.n1640 gnd 0.008189f
C2301 vdd.n1641 gnd 0.836857f
C2302 vdd.n1642 gnd 0.008189f
C2303 vdd.n1643 gnd 0.006591f
C2304 vdd.n1644 gnd 0.019956f
C2305 vdd.n1645 gnd 0.005471f
C2306 vdd.n1646 gnd 0.019956f
C2307 vdd.t43 gnd 0.418428f
C2308 vdd.n1647 gnd 0.019956f
C2309 vdd.n1648 gnd 0.005471f
C2310 vdd.n1649 gnd 0.008189f
C2311 vdd.n1650 gnd 0.006591f
C2312 vdd.n1651 gnd 0.008189f
C2313 vdd.n1682 gnd 0.020414f
C2314 vdd.n1683 gnd 1.23436f
C2315 vdd.n1684 gnd 0.008189f
C2316 vdd.n1685 gnd 0.006591f
C2317 vdd.n1686 gnd 0.008189f
C2318 vdd.n1687 gnd 0.008189f
C2319 vdd.n1688 gnd 0.008189f
C2320 vdd.n1689 gnd 0.008189f
C2321 vdd.n1690 gnd 0.008189f
C2322 vdd.n1691 gnd 0.006591f
C2323 vdd.n1692 gnd 0.008189f
C2324 vdd.n1693 gnd 0.008189f
C2325 vdd.n1694 gnd 0.008189f
C2326 vdd.n1695 gnd 0.008189f
C2327 vdd.n1696 gnd 0.008189f
C2328 vdd.n1697 gnd 0.006591f
C2329 vdd.n1698 gnd 0.008189f
C2330 vdd.n1699 gnd 0.008189f
C2331 vdd.n1700 gnd 0.008189f
C2332 vdd.n1701 gnd 0.008189f
C2333 vdd.n1702 gnd 0.008189f
C2334 vdd.n1703 gnd 0.006591f
C2335 vdd.n1704 gnd 0.008189f
C2336 vdd.n1705 gnd 0.008189f
C2337 vdd.n1706 gnd 0.008189f
C2338 vdd.n1707 gnd 0.008189f
C2339 vdd.n1708 gnd 0.008189f
C2340 vdd.t57 gnd 0.100744f
C2341 vdd.t58 gnd 0.107667f
C2342 vdd.t56 gnd 0.13157f
C2343 vdd.n1709 gnd 0.168654f
C2344 vdd.n1710 gnd 0.142359f
C2345 vdd.n1711 gnd 0.014105f
C2346 vdd.n1712 gnd 0.008189f
C2347 vdd.n1713 gnd 0.008189f
C2348 vdd.n1714 gnd 0.008189f
C2349 vdd.n1715 gnd 0.008189f
C2350 vdd.n1716 gnd 0.008189f
C2351 vdd.n1717 gnd 0.006591f
C2352 vdd.n1718 gnd 0.008189f
C2353 vdd.n1719 gnd 0.008189f
C2354 vdd.n1720 gnd 0.008189f
C2355 vdd.n1721 gnd 0.008189f
C2356 vdd.n1722 gnd 0.008189f
C2357 vdd.n1723 gnd 0.006591f
C2358 vdd.n1724 gnd 0.008189f
C2359 vdd.n1725 gnd 0.008189f
C2360 vdd.n1726 gnd 0.008189f
C2361 vdd.n1727 gnd 0.008189f
C2362 vdd.n1728 gnd 0.008189f
C2363 vdd.n1729 gnd 0.006591f
C2364 vdd.n1730 gnd 0.008189f
C2365 vdd.n1731 gnd 0.008189f
C2366 vdd.n1732 gnd 0.008189f
C2367 vdd.n1733 gnd 0.008189f
C2368 vdd.n1734 gnd 0.008189f
C2369 vdd.n1735 gnd 0.006591f
C2370 vdd.n1736 gnd 0.008189f
C2371 vdd.n1737 gnd 0.008189f
C2372 vdd.n1738 gnd 0.008189f
C2373 vdd.n1739 gnd 0.008189f
C2374 vdd.n1740 gnd 0.008189f
C2375 vdd.n1741 gnd 0.006591f
C2376 vdd.n1742 gnd 0.008189f
C2377 vdd.n1743 gnd 0.008189f
C2378 vdd.n1744 gnd 0.008189f
C2379 vdd.n1745 gnd 0.008189f
C2380 vdd.n1746 gnd 0.006591f
C2381 vdd.n1747 gnd 0.008189f
C2382 vdd.n1748 gnd 0.008189f
C2383 vdd.n1749 gnd 0.008189f
C2384 vdd.n1750 gnd 0.008189f
C2385 vdd.n1751 gnd 0.008189f
C2386 vdd.n1752 gnd 0.006591f
C2387 vdd.n1753 gnd 0.008189f
C2388 vdd.n1754 gnd 0.008189f
C2389 vdd.n1755 gnd 0.008189f
C2390 vdd.n1756 gnd 0.008189f
C2391 vdd.n1757 gnd 0.008189f
C2392 vdd.n1758 gnd 0.006591f
C2393 vdd.n1759 gnd 0.008189f
C2394 vdd.n1760 gnd 0.008189f
C2395 vdd.n1761 gnd 0.008189f
C2396 vdd.n1762 gnd 0.008189f
C2397 vdd.n1763 gnd 0.008189f
C2398 vdd.n1764 gnd 0.006591f
C2399 vdd.n1765 gnd 0.008189f
C2400 vdd.n1766 gnd 0.008189f
C2401 vdd.n1767 gnd 0.008189f
C2402 vdd.n1768 gnd 0.008189f
C2403 vdd.n1769 gnd 0.008189f
C2404 vdd.n1770 gnd 0.006591f
C2405 vdd.n1771 gnd 0.008189f
C2406 vdd.n1772 gnd 0.008189f
C2407 vdd.n1773 gnd 0.008189f
C2408 vdd.n1774 gnd 0.008189f
C2409 vdd.t54 gnd 0.100744f
C2410 vdd.t55 gnd 0.107667f
C2411 vdd.t53 gnd 0.13157f
C2412 vdd.n1775 gnd 0.168654f
C2413 vdd.n1776 gnd 0.142359f
C2414 vdd.n1777 gnd 0.010809f
C2415 vdd.n1778 gnd 0.003131f
C2416 vdd.n1779 gnd 0.020414f
C2417 vdd.n1780 gnd 0.008189f
C2418 vdd.n1781 gnd 0.00346f
C2419 vdd.n1782 gnd 0.006591f
C2420 vdd.n1783 gnd 0.006591f
C2421 vdd.n1784 gnd 0.008189f
C2422 vdd.n1785 gnd 0.008189f
C2423 vdd.n1786 gnd 0.008189f
C2424 vdd.n1787 gnd 0.006591f
C2425 vdd.n1788 gnd 0.006591f
C2426 vdd.n1789 gnd 0.006591f
C2427 vdd.n1790 gnd 0.008189f
C2428 vdd.n1791 gnd 0.008189f
C2429 vdd.n1792 gnd 0.008189f
C2430 vdd.n1793 gnd 0.006591f
C2431 vdd.n1794 gnd 0.006591f
C2432 vdd.n1795 gnd 0.006591f
C2433 vdd.n1796 gnd 0.008189f
C2434 vdd.n1797 gnd 0.008189f
C2435 vdd.n1798 gnd 0.008189f
C2436 vdd.n1799 gnd 0.006591f
C2437 vdd.n1800 gnd 0.006591f
C2438 vdd.n1801 gnd 0.006591f
C2439 vdd.n1802 gnd 0.008189f
C2440 vdd.n1803 gnd 0.008189f
C2441 vdd.n1804 gnd 0.008189f
C2442 vdd.n1805 gnd 0.006591f
C2443 vdd.n1806 gnd 0.006591f
C2444 vdd.n1807 gnd 0.006591f
C2445 vdd.n1808 gnd 0.008189f
C2446 vdd.n1809 gnd 0.008189f
C2447 vdd.n1810 gnd 0.008189f
C2448 vdd.n1811 gnd 0.006525f
C2449 vdd.n1812 gnd 0.008189f
C2450 vdd.t44 gnd 0.100744f
C2451 vdd.t45 gnd 0.107667f
C2452 vdd.t42 gnd 0.13157f
C2453 vdd.n1813 gnd 0.168654f
C2454 vdd.n1814 gnd 0.142359f
C2455 vdd.n1815 gnd 0.014105f
C2456 vdd.n1816 gnd 0.004482f
C2457 vdd.n1817 gnd 0.008189f
C2458 vdd.n1818 gnd 0.008189f
C2459 vdd.n1819 gnd 0.008189f
C2460 vdd.n1820 gnd 0.006591f
C2461 vdd.n1821 gnd 0.006591f
C2462 vdd.n1822 gnd 0.006591f
C2463 vdd.n1823 gnd 0.008189f
C2464 vdd.n1824 gnd 0.008189f
C2465 vdd.n1825 gnd 0.008189f
C2466 vdd.n1826 gnd 0.006591f
C2467 vdd.n1827 gnd 0.006591f
C2468 vdd.n1828 gnd 0.006591f
C2469 vdd.n1829 gnd 0.008189f
C2470 vdd.n1830 gnd 0.008189f
C2471 vdd.n1831 gnd 0.008189f
C2472 vdd.n1832 gnd 0.006591f
C2473 vdd.n1833 gnd 0.006591f
C2474 vdd.n1834 gnd 0.006591f
C2475 vdd.n1835 gnd 0.008189f
C2476 vdd.n1836 gnd 0.008189f
C2477 vdd.n1837 gnd 0.008189f
C2478 vdd.n1838 gnd 0.006591f
C2479 vdd.n1839 gnd 0.006591f
C2480 vdd.n1840 gnd 0.006591f
C2481 vdd.n1841 gnd 0.008189f
C2482 vdd.n1842 gnd 0.008189f
C2483 vdd.n1843 gnd 0.008189f
C2484 vdd.n1844 gnd 0.006591f
C2485 vdd.n1845 gnd 0.006591f
C2486 vdd.n1846 gnd 0.005503f
C2487 vdd.n1847 gnd 0.008189f
C2488 vdd.n1848 gnd 0.008189f
C2489 vdd.n1849 gnd 0.008189f
C2490 vdd.n1850 gnd 0.005503f
C2491 vdd.n1851 gnd 0.006591f
C2492 vdd.n1852 gnd 0.006591f
C2493 vdd.n1853 gnd 0.008189f
C2494 vdd.n1854 gnd 0.008189f
C2495 vdd.n1855 gnd 0.008189f
C2496 vdd.n1856 gnd 0.006591f
C2497 vdd.n1857 gnd 0.006591f
C2498 vdd.n1858 gnd 0.006591f
C2499 vdd.n1859 gnd 0.008189f
C2500 vdd.n1860 gnd 0.008189f
C2501 vdd.n1861 gnd 0.008189f
C2502 vdd.n1862 gnd 0.006591f
C2503 vdd.n1863 gnd 0.006591f
C2504 vdd.n1864 gnd 0.006591f
C2505 vdd.n1865 gnd 0.008189f
C2506 vdd.n1866 gnd 0.008189f
C2507 vdd.n1867 gnd 0.008189f
C2508 vdd.n1868 gnd 0.006591f
C2509 vdd.n1869 gnd 0.006591f
C2510 vdd.n1870 gnd 0.006591f
C2511 vdd.n1871 gnd 0.008189f
C2512 vdd.n1872 gnd 0.008189f
C2513 vdd.n1873 gnd 0.008189f
C2514 vdd.n1874 gnd 0.006591f
C2515 vdd.n1875 gnd 0.008189f
C2516 vdd.n1876 gnd 2.00009f
C2517 vdd.n1878 gnd 0.020414f
C2518 vdd.n1879 gnd 0.005471f
C2519 vdd.n1880 gnd 0.020414f
C2520 vdd.n1881 gnd 0.019956f
C2521 vdd.n1882 gnd 0.008189f
C2522 vdd.n1883 gnd 0.006591f
C2523 vdd.n1884 gnd 0.008189f
C2524 vdd.n1885 gnd 0.43935f
C2525 vdd.n1886 gnd 0.008189f
C2526 vdd.n1887 gnd 0.006591f
C2527 vdd.n1888 gnd 0.008189f
C2528 vdd.n1889 gnd 0.008189f
C2529 vdd.n1890 gnd 0.008189f
C2530 vdd.n1891 gnd 0.006591f
C2531 vdd.n1892 gnd 0.008189f
C2532 vdd.n1893 gnd 0.748987f
C2533 vdd.n1894 gnd 0.836857f
C2534 vdd.n1895 gnd 0.008189f
C2535 vdd.n1896 gnd 0.006591f
C2536 vdd.n1897 gnd 0.008189f
C2537 vdd.n1898 gnd 0.008189f
C2538 vdd.n1899 gnd 0.008189f
C2539 vdd.n1900 gnd 0.006591f
C2540 vdd.n1901 gnd 0.008189f
C2541 vdd.n1902 gnd 0.506298f
C2542 vdd.n1903 gnd 0.008189f
C2543 vdd.n1904 gnd 0.006591f
C2544 vdd.n1905 gnd 0.008189f
C2545 vdd.n1906 gnd 0.008189f
C2546 vdd.n1907 gnd 0.008189f
C2547 vdd.n1908 gnd 0.006591f
C2548 vdd.n1909 gnd 0.008189f
C2549 vdd.n1910 gnd 0.464456f
C2550 vdd.n1911 gnd 0.648564f
C2551 vdd.n1912 gnd 0.008189f
C2552 vdd.n1913 gnd 0.006591f
C2553 vdd.n1914 gnd 0.008189f
C2554 vdd.n1915 gnd 0.008189f
C2555 vdd.n1916 gnd 0.006294f
C2556 vdd.n1917 gnd 0.008189f
C2557 vdd.n1918 gnd 0.006591f
C2558 vdd.n1919 gnd 0.008189f
C2559 vdd.n1920 gnd 0.694591f
C2560 vdd.n1921 gnd 0.008189f
C2561 vdd.n1922 gnd 0.006591f
C2562 vdd.n1923 gnd 0.008189f
C2563 vdd.n1924 gnd 0.008189f
C2564 vdd.n1925 gnd 0.008189f
C2565 vdd.n1926 gnd 0.006591f
C2566 vdd.n1927 gnd 0.008189f
C2567 vdd.t96 gnd 0.418428f
C2568 vdd.n1928 gnd 0.598353f
C2569 vdd.n1929 gnd 0.008189f
C2570 vdd.n1930 gnd 0.006591f
C2571 vdd.n1931 gnd 0.006294f
C2572 vdd.n1932 gnd 0.008189f
C2573 vdd.n1933 gnd 0.008189f
C2574 vdd.n1934 gnd 0.006591f
C2575 vdd.n1935 gnd 0.008189f
C2576 vdd.n1936 gnd 0.456087f
C2577 vdd.n1937 gnd 0.008189f
C2578 vdd.n1938 gnd 0.006591f
C2579 vdd.n1939 gnd 0.008189f
C2580 vdd.n1940 gnd 0.008189f
C2581 vdd.n1941 gnd 0.008189f
C2582 vdd.n1942 gnd 0.006591f
C2583 vdd.n1943 gnd 0.008189f
C2584 vdd.n1944 gnd 0.589984f
C2585 vdd.n1945 gnd 0.523035f
C2586 vdd.n1946 gnd 0.008189f
C2587 vdd.n1947 gnd 0.006591f
C2588 vdd.n1948 gnd 0.008189f
C2589 vdd.n1949 gnd 0.008189f
C2590 vdd.n1950 gnd 0.008189f
C2591 vdd.n1951 gnd 0.006591f
C2592 vdd.n1952 gnd 0.008189f
C2593 vdd.n1953 gnd 0.665301f
C2594 vdd.n1954 gnd 0.008189f
C2595 vdd.n1955 gnd 0.006591f
C2596 vdd.n1956 gnd 0.008189f
C2597 vdd.n1957 gnd 0.008189f
C2598 vdd.n1958 gnd 0.019956f
C2599 vdd.n1959 gnd 0.008189f
C2600 vdd.n1960 gnd 0.008189f
C2601 vdd.n1961 gnd 0.006591f
C2602 vdd.n1962 gnd 0.008189f
C2603 vdd.n1963 gnd 0.523035f
C2604 vdd.n1964 gnd 0.836857f
C2605 vdd.n1965 gnd 0.008189f
C2606 vdd.n1966 gnd 0.006591f
C2607 vdd.n1967 gnd 0.008189f
C2608 vdd.n1968 gnd 0.008189f
C2609 vdd.n1969 gnd 0.019956f
C2610 vdd.n1970 gnd 0.005471f
C2611 vdd.n1971 gnd 0.019956f
C2612 vdd.n1972 gnd 1.15068f
C2613 vdd.n1973 gnd 0.019956f
C2614 vdd.n1974 gnd 0.020414f
C2615 vdd.n1975 gnd 0.003131f
C2616 vdd.t48 gnd 0.100744f
C2617 vdd.t47 gnd 0.107667f
C2618 vdd.t46 gnd 0.13157f
C2619 vdd.n1976 gnd 0.168654f
C2620 vdd.n1977 gnd 0.1417f
C2621 vdd.n1978 gnd 0.01015f
C2622 vdd.n1979 gnd 0.00346f
C2623 vdd.n1980 gnd 0.007042f
C2624 vdd.n1981 gnd 0.869326f
C2625 vdd.n1983 gnd 0.006591f
C2626 vdd.n1984 gnd 0.006591f
C2627 vdd.n1985 gnd 0.008189f
C2628 vdd.n1987 gnd 0.008189f
C2629 vdd.n1988 gnd 0.008189f
C2630 vdd.n1989 gnd 0.006591f
C2631 vdd.n1990 gnd 0.006591f
C2632 vdd.n1991 gnd 0.006591f
C2633 vdd.n1992 gnd 0.008189f
C2634 vdd.n1994 gnd 0.008189f
C2635 vdd.n1995 gnd 0.008189f
C2636 vdd.n1996 gnd 0.006591f
C2637 vdd.n1997 gnd 0.006591f
C2638 vdd.n1998 gnd 0.006591f
C2639 vdd.n1999 gnd 0.008189f
C2640 vdd.n2001 gnd 0.008189f
C2641 vdd.n2002 gnd 0.008189f
C2642 vdd.n2003 gnd 0.006591f
C2643 vdd.n2004 gnd 0.006591f
C2644 vdd.n2005 gnd 0.006591f
C2645 vdd.n2006 gnd 0.008189f
C2646 vdd.n2008 gnd 0.008189f
C2647 vdd.n2009 gnd 0.008189f
C2648 vdd.n2010 gnd 0.006591f
C2649 vdd.n2011 gnd 0.008189f
C2650 vdd.n2012 gnd 0.008189f
C2651 vdd.n2013 gnd 0.008189f
C2652 vdd.n2014 gnd 0.013446f
C2653 vdd.n2015 gnd 0.004482f
C2654 vdd.n2016 gnd 0.006591f
C2655 vdd.n2017 gnd 0.008189f
C2656 vdd.n2019 gnd 0.008189f
C2657 vdd.n2020 gnd 0.008189f
C2658 vdd.n2021 gnd 0.006591f
C2659 vdd.n2022 gnd 0.006591f
C2660 vdd.n2023 gnd 0.006591f
C2661 vdd.n2024 gnd 0.008189f
C2662 vdd.n2026 gnd 0.008189f
C2663 vdd.n2027 gnd 0.008189f
C2664 vdd.n2028 gnd 0.006591f
C2665 vdd.n2029 gnd 0.006591f
C2666 vdd.n2030 gnd 0.006591f
C2667 vdd.n2031 gnd 0.008189f
C2668 vdd.n2033 gnd 0.008189f
C2669 vdd.n2034 gnd 0.008189f
C2670 vdd.n2035 gnd 0.006591f
C2671 vdd.n2036 gnd 0.006591f
C2672 vdd.n2037 gnd 0.006591f
C2673 vdd.n2038 gnd 0.008189f
C2674 vdd.n2040 gnd 0.008189f
C2675 vdd.n2041 gnd 0.008189f
C2676 vdd.n2042 gnd 0.006591f
C2677 vdd.n2043 gnd 0.006591f
C2678 vdd.n2044 gnd 0.006591f
C2679 vdd.n2045 gnd 0.008189f
C2680 vdd.n2047 gnd 0.008189f
C2681 vdd.n2048 gnd 0.008189f
C2682 vdd.n2049 gnd 0.006591f
C2683 vdd.n2050 gnd 0.008189f
C2684 vdd.n2051 gnd 0.008189f
C2685 vdd.n2052 gnd 0.008189f
C2686 vdd.n2053 gnd 0.013446f
C2687 vdd.n2054 gnd 0.005503f
C2688 vdd.n2055 gnd 0.006591f
C2689 vdd.n2056 gnd 0.008189f
C2690 vdd.n2058 gnd 0.008189f
C2691 vdd.n2059 gnd 0.008189f
C2692 vdd.n2060 gnd 0.006591f
C2693 vdd.n2061 gnd 0.006591f
C2694 vdd.n2062 gnd 0.006591f
C2695 vdd.n2063 gnd 0.008189f
C2696 vdd.n2065 gnd 0.008189f
C2697 vdd.n2066 gnd 0.008189f
C2698 vdd.n2067 gnd 0.006591f
C2699 vdd.n2068 gnd 0.006591f
C2700 vdd.n2069 gnd 0.006591f
C2701 vdd.n2070 gnd 0.008189f
C2702 vdd.n2072 gnd 0.008189f
C2703 vdd.n2073 gnd 0.008189f
C2704 vdd.n2074 gnd 0.006591f
C2705 vdd.n2075 gnd 0.006591f
C2706 vdd.n2076 gnd 0.006591f
C2707 vdd.n2077 gnd 0.008189f
C2708 vdd.n2079 gnd 0.008189f
C2709 vdd.n2080 gnd 0.006591f
C2710 vdd.n2081 gnd 0.006591f
C2711 vdd.n2082 gnd 0.008189f
C2712 vdd.n2084 gnd 0.008189f
C2713 vdd.n2085 gnd 0.008189f
C2714 vdd.n2086 gnd 0.006591f
C2715 vdd.n2087 gnd 0.007042f
C2716 vdd.n2088 gnd 0.869326f
C2717 vdd.n2089 gnd 0.037512f
C2718 vdd.n2090 gnd 0.005568f
C2719 vdd.n2091 gnd 0.005568f
C2720 vdd.n2092 gnd 0.005568f
C2721 vdd.n2093 gnd 0.005568f
C2722 vdd.n2094 gnd 0.005568f
C2723 vdd.n2095 gnd 0.005568f
C2724 vdd.n2096 gnd 0.005568f
C2725 vdd.n2097 gnd 0.005568f
C2726 vdd.n2098 gnd 0.005568f
C2727 vdd.n2099 gnd 0.005568f
C2728 vdd.n2100 gnd 0.005568f
C2729 vdd.n2101 gnd 0.005568f
C2730 vdd.n2102 gnd 0.005568f
C2731 vdd.n2103 gnd 0.005568f
C2732 vdd.n2104 gnd 0.005568f
C2733 vdd.n2105 gnd 0.005568f
C2734 vdd.n2106 gnd 0.005568f
C2735 vdd.n2107 gnd 0.005568f
C2736 vdd.n2108 gnd 0.005568f
C2737 vdd.n2109 gnd 0.005568f
C2738 vdd.n2110 gnd 0.005568f
C2739 vdd.n2111 gnd 0.005568f
C2740 vdd.n2112 gnd 0.005568f
C2741 vdd.n2113 gnd 0.005568f
C2742 vdd.n2114 gnd 0.005568f
C2743 vdd.n2115 gnd 0.005568f
C2744 vdd.n2116 gnd 0.005568f
C2745 vdd.n2117 gnd 0.005568f
C2746 vdd.n2118 gnd 0.005568f
C2747 vdd.n2119 gnd 0.005568f
C2748 vdd.n2120 gnd 9.883281f
C2749 vdd.n2122 gnd 0.012644f
C2750 vdd.n2123 gnd 0.012644f
C2751 vdd.n2124 gnd 0.011923f
C2752 vdd.n2125 gnd 0.005568f
C2753 vdd.n2126 gnd 0.005568f
C2754 vdd.n2127 gnd 0.569063f
C2755 vdd.n2128 gnd 0.005568f
C2756 vdd.n2129 gnd 0.005568f
C2757 vdd.n2130 gnd 0.005568f
C2758 vdd.n2131 gnd 0.005568f
C2759 vdd.n2132 gnd 0.005568f
C2760 vdd.n2133 gnd 0.447718f
C2761 vdd.n2134 gnd 0.005568f
C2762 vdd.n2135 gnd 0.005568f
C2763 vdd.n2136 gnd 0.005568f
C2764 vdd.n2137 gnd 0.005568f
C2765 vdd.n2138 gnd 0.005568f
C2766 vdd.n2139 gnd 0.569063f
C2767 vdd.n2140 gnd 0.005568f
C2768 vdd.n2141 gnd 0.005568f
C2769 vdd.n2142 gnd 0.005568f
C2770 vdd.n2143 gnd 0.005568f
C2771 vdd.n2144 gnd 0.005568f
C2772 vdd.n2145 gnd 0.569063f
C2773 vdd.n2146 gnd 0.005568f
C2774 vdd.n2147 gnd 0.005568f
C2775 vdd.n2148 gnd 0.005568f
C2776 vdd.n2149 gnd 0.005568f
C2777 vdd.n2150 gnd 0.005568f
C2778 vdd.n2151 gnd 0.548141f
C2779 vdd.n2152 gnd 0.005568f
C2780 vdd.n2153 gnd 0.005568f
C2781 vdd.n2154 gnd 0.005568f
C2782 vdd.n2155 gnd 0.005568f
C2783 vdd.n2156 gnd 0.005568f
C2784 vdd.n2157 gnd 0.422613f
C2785 vdd.n2158 gnd 0.005568f
C2786 vdd.n2159 gnd 0.005568f
C2787 vdd.n2160 gnd 0.005568f
C2788 vdd.n2161 gnd 0.005568f
C2789 vdd.n2162 gnd 0.005568f
C2790 vdd.n2163 gnd 0.297084f
C2791 vdd.n2164 gnd 0.005568f
C2792 vdd.n2165 gnd 0.005568f
C2793 vdd.n2166 gnd 0.005568f
C2794 vdd.n2167 gnd 0.005568f
C2795 vdd.n2168 gnd 0.005568f
C2796 vdd.n2169 gnd 0.397507f
C2797 vdd.n2170 gnd 0.005568f
C2798 vdd.n2171 gnd 0.005568f
C2799 vdd.n2172 gnd 0.005568f
C2800 vdd.n2173 gnd 0.005568f
C2801 vdd.n2174 gnd 0.005568f
C2802 vdd.n2175 gnd 0.523035f
C2803 vdd.n2176 gnd 0.005568f
C2804 vdd.n2177 gnd 0.005568f
C2805 vdd.n2178 gnd 0.005568f
C2806 vdd.n2179 gnd 0.005568f
C2807 vdd.n2180 gnd 0.005568f
C2808 vdd.n2181 gnd 0.569063f
C2809 vdd.n2182 gnd 0.005568f
C2810 vdd.n2183 gnd 0.005568f
C2811 vdd.n2184 gnd 0.005568f
C2812 vdd.n2185 gnd 0.005568f
C2813 vdd.n2186 gnd 0.005568f
C2814 vdd.n2187 gnd 0.489561f
C2815 vdd.n2188 gnd 0.005568f
C2816 vdd.n2189 gnd 0.005568f
C2817 vdd.n2190 gnd 0.004422f
C2818 vdd.n2191 gnd 0.016131f
C2819 vdd.n2192 gnd 0.003931f
C2820 vdd.n2193 gnd 0.005568f
C2821 vdd.n2194 gnd 0.364033f
C2822 vdd.n2195 gnd 0.005568f
C2823 vdd.n2196 gnd 0.005568f
C2824 vdd.n2197 gnd 0.005568f
C2825 vdd.n2198 gnd 0.005568f
C2826 vdd.n2199 gnd 0.005568f
C2827 vdd.n2200 gnd 0.330558f
C2828 vdd.n2201 gnd 0.005568f
C2829 vdd.n2202 gnd 0.005568f
C2830 vdd.n2203 gnd 0.005568f
C2831 vdd.n2204 gnd 0.005568f
C2832 vdd.n2205 gnd 0.005568f
C2833 vdd.n2206 gnd 0.456087f
C2834 vdd.n2207 gnd 0.005568f
C2835 vdd.n2208 gnd 0.005568f
C2836 vdd.n2209 gnd 0.005568f
C2837 vdd.n2210 gnd 0.005568f
C2838 vdd.n2211 gnd 0.005568f
C2839 vdd.n2212 gnd 0.502114f
C2840 vdd.n2213 gnd 0.005568f
C2841 vdd.n2214 gnd 0.005568f
C2842 vdd.n2215 gnd 0.005568f
C2843 vdd.n2216 gnd 0.005568f
C2844 vdd.n2217 gnd 0.005568f
C2845 vdd.n2218 gnd 0.376586f
C2846 vdd.n2219 gnd 0.005568f
C2847 vdd.n2220 gnd 0.005568f
C2848 vdd.n2221 gnd 0.005568f
C2849 vdd.n2222 gnd 0.005568f
C2850 vdd.n2223 gnd 0.005568f
C2851 vdd.n2224 gnd 0.179924f
C2852 vdd.n2225 gnd 0.005568f
C2853 vdd.n2226 gnd 0.005568f
C2854 vdd.n2227 gnd 0.005568f
C2855 vdd.n2228 gnd 0.005568f
C2856 vdd.n2229 gnd 0.005568f
C2857 vdd.n2230 gnd 0.179924f
C2858 vdd.n2231 gnd 0.005568f
C2859 vdd.n2232 gnd 0.005568f
C2860 vdd.n2233 gnd 0.005568f
C2861 vdd.n2234 gnd 0.005568f
C2862 vdd.n2235 gnd 0.005568f
C2863 vdd.n2236 gnd 0.569063f
C2864 vdd.n2237 gnd 0.005568f
C2865 vdd.n2238 gnd 0.005568f
C2866 vdd.n2239 gnd 0.005568f
C2867 vdd.n2240 gnd 0.005568f
C2868 vdd.n2241 gnd 0.005568f
C2869 vdd.n2242 gnd 0.005568f
C2870 vdd.n2243 gnd 0.005568f
C2871 vdd.n2244 gnd 0.393323f
C2872 vdd.n2245 gnd 0.005568f
C2873 vdd.n2246 gnd 0.005568f
C2874 vdd.n2247 gnd 0.005568f
C2875 vdd.n2248 gnd 0.005568f
C2876 vdd.n2249 gnd 0.005568f
C2877 vdd.n2250 gnd 0.005568f
C2878 vdd.n2251 gnd 0.355664f
C2879 vdd.n2252 gnd 0.005568f
C2880 vdd.n2253 gnd 0.005568f
C2881 vdd.n2254 gnd 0.005568f
C2882 vdd.n2255 gnd 0.012644f
C2883 vdd.n2256 gnd 0.011923f
C2884 vdd.n2257 gnd 0.005568f
C2885 vdd.n2258 gnd 0.005568f
C2886 vdd.n2259 gnd 0.004299f
C2887 vdd.n2260 gnd 0.005568f
C2888 vdd.n2261 gnd 0.005568f
C2889 vdd.n2262 gnd 0.004053f
C2890 vdd.n2263 gnd 0.005568f
C2891 vdd.n2264 gnd 0.005568f
C2892 vdd.n2265 gnd 0.005568f
C2893 vdd.n2266 gnd 0.005568f
C2894 vdd.n2267 gnd 0.005568f
C2895 vdd.n2268 gnd 0.005568f
C2896 vdd.n2269 gnd 0.005568f
C2897 vdd.n2270 gnd 0.005568f
C2898 vdd.n2271 gnd 0.005568f
C2899 vdd.n2272 gnd 0.005568f
C2900 vdd.n2273 gnd 0.005568f
C2901 vdd.n2274 gnd 0.005568f
C2902 vdd.n2275 gnd 0.005568f
C2903 vdd.n2276 gnd 0.005568f
C2904 vdd.n2277 gnd 0.005568f
C2905 vdd.n2278 gnd 0.005568f
C2906 vdd.n2279 gnd 0.005568f
C2907 vdd.n2280 gnd 0.005568f
C2908 vdd.n2281 gnd 0.005568f
C2909 vdd.n2282 gnd 0.005568f
C2910 vdd.n2283 gnd 0.005568f
C2911 vdd.n2284 gnd 0.005568f
C2912 vdd.n2285 gnd 0.005568f
C2913 vdd.n2286 gnd 0.005568f
C2914 vdd.n2287 gnd 0.005568f
C2915 vdd.n2288 gnd 0.005568f
C2916 vdd.n2289 gnd 0.005568f
C2917 vdd.n2290 gnd 0.005568f
C2918 vdd.n2291 gnd 0.005568f
C2919 vdd.n2292 gnd 0.005568f
C2920 vdd.n2293 gnd 0.005568f
C2921 vdd.n2294 gnd 0.005568f
C2922 vdd.n2295 gnd 0.005568f
C2923 vdd.n2296 gnd 0.005568f
C2924 vdd.n2297 gnd 0.005568f
C2925 vdd.n2298 gnd 0.005568f
C2926 vdd.n2299 gnd 0.005568f
C2927 vdd.n2300 gnd 0.005568f
C2928 vdd.n2301 gnd 0.005568f
C2929 vdd.n2302 gnd 0.005568f
C2930 vdd.n2303 gnd 0.005568f
C2931 vdd.n2304 gnd 0.005568f
C2932 vdd.n2305 gnd 0.005568f
C2933 vdd.n2306 gnd 0.005568f
C2934 vdd.n2307 gnd 0.005568f
C2935 vdd.n2308 gnd 0.005568f
C2936 vdd.n2309 gnd 0.005568f
C2937 vdd.n2310 gnd 0.005568f
C2938 vdd.n2311 gnd 0.005568f
C2939 vdd.n2312 gnd 0.005568f
C2940 vdd.n2313 gnd 0.005568f
C2941 vdd.n2314 gnd 0.005568f
C2942 vdd.n2315 gnd 0.005568f
C2943 vdd.n2316 gnd 0.005568f
C2944 vdd.n2317 gnd 0.005568f
C2945 vdd.n2318 gnd 0.005568f
C2946 vdd.n2319 gnd 0.005568f
C2947 vdd.n2320 gnd 0.005568f
C2948 vdd.n2321 gnd 0.005568f
C2949 vdd.n2322 gnd 0.005568f
C2950 vdd.n2323 gnd 0.012644f
C2951 vdd.n2324 gnd 0.011923f
C2952 vdd.n2325 gnd 0.011923f
C2953 vdd.n2326 gnd 0.64438f
C2954 vdd.n2327 gnd 0.011923f
C2955 vdd.n2328 gnd 0.012644f
C2956 vdd.n2329 gnd 0.011923f
C2957 vdd.n2330 gnd 0.005568f
C2958 vdd.n2331 gnd 0.005568f
C2959 vdd.n2332 gnd 0.005568f
C2960 vdd.n2333 gnd 0.004299f
C2961 vdd.n2334 gnd 0.007958f
C2962 vdd.n2335 gnd 0.004053f
C2963 vdd.n2336 gnd 0.005568f
C2964 vdd.n2337 gnd 0.005568f
C2965 vdd.n2338 gnd 0.005568f
C2966 vdd.n2339 gnd 0.005568f
C2967 vdd.n2340 gnd 0.005568f
C2968 vdd.n2341 gnd 0.005568f
C2969 vdd.n2342 gnd 0.005568f
C2970 vdd.n2343 gnd 0.005568f
C2971 vdd.n2344 gnd 0.005568f
C2972 vdd.n2345 gnd 0.005568f
C2973 vdd.n2346 gnd 0.005568f
C2974 vdd.n2347 gnd 0.005568f
C2975 vdd.n2348 gnd 0.005568f
C2976 vdd.n2349 gnd 0.005568f
C2977 vdd.n2350 gnd 0.005568f
C2978 vdd.n2351 gnd 0.005568f
C2979 vdd.n2352 gnd 0.005568f
C2980 vdd.n2353 gnd 0.005568f
C2981 vdd.n2354 gnd 0.005568f
C2982 vdd.n2355 gnd 0.005568f
C2983 vdd.n2356 gnd 0.005568f
C2984 vdd.n2357 gnd 0.005568f
C2985 vdd.n2358 gnd 0.005568f
C2986 vdd.n2359 gnd 0.005568f
C2987 vdd.n2360 gnd 0.005568f
C2988 vdd.n2361 gnd 0.005568f
C2989 vdd.n2362 gnd 0.005568f
C2990 vdd.n2363 gnd 0.005568f
C2991 vdd.n2364 gnd 0.005568f
C2992 vdd.n2365 gnd 0.005568f
C2993 vdd.n2366 gnd 0.005568f
C2994 vdd.n2367 gnd 0.005568f
C2995 vdd.n2368 gnd 0.005568f
C2996 vdd.n2369 gnd 0.005568f
C2997 vdd.n2370 gnd 0.005568f
C2998 vdd.n2371 gnd 0.005568f
C2999 vdd.n2372 gnd 0.005568f
C3000 vdd.n2373 gnd 0.005568f
C3001 vdd.n2374 gnd 0.005568f
C3002 vdd.n2375 gnd 0.005568f
C3003 vdd.n2376 gnd 0.005568f
C3004 vdd.n2377 gnd 0.005568f
C3005 vdd.n2378 gnd 0.005568f
C3006 vdd.n2379 gnd 0.005568f
C3007 vdd.n2380 gnd 0.005568f
C3008 vdd.n2381 gnd 0.005568f
C3009 vdd.n2382 gnd 0.005568f
C3010 vdd.n2383 gnd 0.005568f
C3011 vdd.n2384 gnd 0.005568f
C3012 vdd.n2385 gnd 0.005568f
C3013 vdd.n2386 gnd 0.005568f
C3014 vdd.n2387 gnd 0.005568f
C3015 vdd.n2388 gnd 0.005568f
C3016 vdd.n2389 gnd 0.005568f
C3017 vdd.n2390 gnd 0.005568f
C3018 vdd.n2391 gnd 0.005568f
C3019 vdd.n2392 gnd 0.005568f
C3020 vdd.n2393 gnd 0.005568f
C3021 vdd.n2394 gnd 0.005568f
C3022 vdd.n2395 gnd 0.005568f
C3023 vdd.n2396 gnd 0.012644f
C3024 vdd.n2397 gnd 0.012644f
C3025 vdd.n2398 gnd 0.694591f
C3026 vdd.t184 gnd 2.46873f
C3027 vdd.t166 gnd 2.46873f
C3028 vdd.n2432 gnd 0.012644f
C3029 vdd.t189 gnd 0.485377f
C3030 vdd.n2433 gnd 0.005568f
C3031 vdd.t74 gnd 0.225018f
C3032 vdd.t75 gnd 0.230334f
C3033 vdd.t72 gnd 0.1469f
C3034 vdd.n2434 gnd 0.079392f
C3035 vdd.n2435 gnd 0.045033f
C3036 vdd.n2436 gnd 0.005568f
C3037 vdd.t81 gnd 0.225018f
C3038 vdd.t82 gnd 0.230334f
C3039 vdd.t80 gnd 0.1469f
C3040 vdd.n2437 gnd 0.079392f
C3041 vdd.n2438 gnd 0.045033f
C3042 vdd.n2439 gnd 0.007958f
C3043 vdd.n2440 gnd 0.012644f
C3044 vdd.n2441 gnd 0.012644f
C3045 vdd.n2442 gnd 0.005568f
C3046 vdd.n2443 gnd 0.005568f
C3047 vdd.n2444 gnd 0.005568f
C3048 vdd.n2445 gnd 0.005568f
C3049 vdd.n2446 gnd 0.005568f
C3050 vdd.n2447 gnd 0.005568f
C3051 vdd.n2448 gnd 0.005568f
C3052 vdd.n2449 gnd 0.005568f
C3053 vdd.n2450 gnd 0.005568f
C3054 vdd.n2451 gnd 0.005568f
C3055 vdd.n2452 gnd 0.005568f
C3056 vdd.n2453 gnd 0.005568f
C3057 vdd.n2454 gnd 0.005568f
C3058 vdd.n2455 gnd 0.005568f
C3059 vdd.n2456 gnd 0.005568f
C3060 vdd.n2457 gnd 0.005568f
C3061 vdd.n2458 gnd 0.005568f
C3062 vdd.n2459 gnd 0.005568f
C3063 vdd.n2460 gnd 0.005568f
C3064 vdd.n2461 gnd 0.005568f
C3065 vdd.n2462 gnd 0.005568f
C3066 vdd.n2463 gnd 0.005568f
C3067 vdd.n2464 gnd 0.005568f
C3068 vdd.n2465 gnd 0.005568f
C3069 vdd.n2466 gnd 0.005568f
C3070 vdd.n2467 gnd 0.005568f
C3071 vdd.n2468 gnd 0.005568f
C3072 vdd.n2469 gnd 0.005568f
C3073 vdd.n2470 gnd 0.005568f
C3074 vdd.n2471 gnd 0.005568f
C3075 vdd.n2472 gnd 0.005568f
C3076 vdd.n2473 gnd 0.005568f
C3077 vdd.n2474 gnd 0.005568f
C3078 vdd.n2475 gnd 0.005568f
C3079 vdd.n2476 gnd 0.005568f
C3080 vdd.n2477 gnd 0.005568f
C3081 vdd.n2478 gnd 0.005568f
C3082 vdd.n2479 gnd 0.005568f
C3083 vdd.n2480 gnd 0.005568f
C3084 vdd.n2481 gnd 0.005568f
C3085 vdd.n2482 gnd 0.005568f
C3086 vdd.n2483 gnd 0.005568f
C3087 vdd.n2484 gnd 0.005568f
C3088 vdd.n2485 gnd 0.005568f
C3089 vdd.n2486 gnd 0.005568f
C3090 vdd.n2487 gnd 0.005568f
C3091 vdd.n2488 gnd 0.005568f
C3092 vdd.n2489 gnd 0.005568f
C3093 vdd.n2490 gnd 0.005568f
C3094 vdd.n2491 gnd 0.005568f
C3095 vdd.n2492 gnd 0.005568f
C3096 vdd.n2493 gnd 0.005568f
C3097 vdd.n2494 gnd 0.005568f
C3098 vdd.n2495 gnd 0.005568f
C3099 vdd.n2496 gnd 0.005568f
C3100 vdd.n2497 gnd 0.005568f
C3101 vdd.n2498 gnd 0.005568f
C3102 vdd.n2499 gnd 0.005568f
C3103 vdd.n2500 gnd 0.005568f
C3104 vdd.n2501 gnd 0.005568f
C3105 vdd.n2502 gnd 0.004053f
C3106 vdd.n2503 gnd 0.005568f
C3107 vdd.n2504 gnd 0.005568f
C3108 vdd.n2505 gnd 0.004299f
C3109 vdd.n2506 gnd 0.005568f
C3110 vdd.n2507 gnd 0.005568f
C3111 vdd.n2508 gnd 0.012644f
C3112 vdd.n2509 gnd 0.011923f
C3113 vdd.n2510 gnd 0.011923f
C3114 vdd.n2511 gnd 0.005568f
C3115 vdd.n2512 gnd 0.005568f
C3116 vdd.n2513 gnd 0.005568f
C3117 vdd.n2514 gnd 0.005568f
C3118 vdd.n2515 gnd 0.005568f
C3119 vdd.n2516 gnd 0.005568f
C3120 vdd.n2517 gnd 0.005568f
C3121 vdd.n2518 gnd 0.005568f
C3122 vdd.n2519 gnd 0.005568f
C3123 vdd.n2520 gnd 0.005568f
C3124 vdd.n2521 gnd 0.005568f
C3125 vdd.n2522 gnd 0.005568f
C3126 vdd.n2523 gnd 0.005568f
C3127 vdd.n2524 gnd 0.005568f
C3128 vdd.n2525 gnd 0.005568f
C3129 vdd.n2526 gnd 0.005568f
C3130 vdd.n2527 gnd 0.005568f
C3131 vdd.n2528 gnd 0.005568f
C3132 vdd.n2529 gnd 0.005568f
C3133 vdd.n2530 gnd 0.005568f
C3134 vdd.n2531 gnd 0.005568f
C3135 vdd.n2532 gnd 0.005568f
C3136 vdd.n2533 gnd 0.005568f
C3137 vdd.n2534 gnd 0.005568f
C3138 vdd.n2535 gnd 0.005568f
C3139 vdd.n2536 gnd 0.005568f
C3140 vdd.n2537 gnd 0.005568f
C3141 vdd.n2538 gnd 0.005568f
C3142 vdd.n2539 gnd 0.005568f
C3143 vdd.n2540 gnd 0.005568f
C3144 vdd.n2541 gnd 0.005568f
C3145 vdd.n2542 gnd 0.005568f
C3146 vdd.n2543 gnd 0.005568f
C3147 vdd.n2544 gnd 0.005568f
C3148 vdd.n2545 gnd 0.005568f
C3149 vdd.n2546 gnd 0.005568f
C3150 vdd.n2547 gnd 0.005568f
C3151 vdd.n2548 gnd 0.005568f
C3152 vdd.n2549 gnd 0.005568f
C3153 vdd.n2550 gnd 0.005568f
C3154 vdd.n2551 gnd 0.005568f
C3155 vdd.n2552 gnd 0.005568f
C3156 vdd.n2553 gnd 0.005568f
C3157 vdd.n2554 gnd 0.005568f
C3158 vdd.n2555 gnd 0.005568f
C3159 vdd.n2556 gnd 0.005568f
C3160 vdd.n2557 gnd 0.005568f
C3161 vdd.n2558 gnd 0.005568f
C3162 vdd.n2559 gnd 0.005568f
C3163 vdd.n2560 gnd 0.005568f
C3164 vdd.n2561 gnd 0.005568f
C3165 vdd.n2562 gnd 0.005568f
C3166 vdd.n2563 gnd 0.005568f
C3167 vdd.n2564 gnd 0.005568f
C3168 vdd.n2565 gnd 0.005568f
C3169 vdd.n2566 gnd 0.005568f
C3170 vdd.n2567 gnd 0.005568f
C3171 vdd.n2568 gnd 0.005568f
C3172 vdd.n2569 gnd 0.005568f
C3173 vdd.n2570 gnd 0.005568f
C3174 vdd.n2571 gnd 0.005568f
C3175 vdd.n2572 gnd 0.005568f
C3176 vdd.n2573 gnd 0.005568f
C3177 vdd.n2574 gnd 0.005568f
C3178 vdd.n2575 gnd 0.005568f
C3179 vdd.n2576 gnd 0.005568f
C3180 vdd.n2577 gnd 0.005568f
C3181 vdd.n2578 gnd 0.005568f
C3182 vdd.n2579 gnd 0.005568f
C3183 vdd.n2580 gnd 0.005568f
C3184 vdd.n2581 gnd 0.005568f
C3185 vdd.n2582 gnd 0.005568f
C3186 vdd.n2583 gnd 0.005568f
C3187 vdd.n2584 gnd 0.005568f
C3188 vdd.n2585 gnd 0.005568f
C3189 vdd.n2586 gnd 0.005568f
C3190 vdd.n2587 gnd 0.005568f
C3191 vdd.n2588 gnd 0.005568f
C3192 vdd.n2589 gnd 0.005568f
C3193 vdd.n2590 gnd 0.005568f
C3194 vdd.n2591 gnd 0.005568f
C3195 vdd.n2592 gnd 0.005568f
C3196 vdd.n2593 gnd 0.005568f
C3197 vdd.n2594 gnd 0.005568f
C3198 vdd.n2595 gnd 0.005568f
C3199 vdd.n2596 gnd 0.005568f
C3200 vdd.n2597 gnd 0.005568f
C3201 vdd.n2598 gnd 0.005568f
C3202 vdd.n2599 gnd 0.005568f
C3203 vdd.n2600 gnd 0.005568f
C3204 vdd.n2601 gnd 0.005568f
C3205 vdd.n2602 gnd 0.005568f
C3206 vdd.n2603 gnd 0.005568f
C3207 vdd.n2604 gnd 0.005568f
C3208 vdd.n2605 gnd 0.005568f
C3209 vdd.n2606 gnd 0.005568f
C3210 vdd.n2607 gnd 0.005568f
C3211 vdd.n2608 gnd 0.005568f
C3212 vdd.n2609 gnd 0.005568f
C3213 vdd.n2610 gnd 0.005568f
C3214 vdd.n2611 gnd 0.005568f
C3215 vdd.n2612 gnd 0.179924f
C3216 vdd.n2613 gnd 0.005568f
C3217 vdd.n2614 gnd 0.005568f
C3218 vdd.n2615 gnd 0.005568f
C3219 vdd.n2616 gnd 0.005568f
C3220 vdd.n2617 gnd 0.005568f
C3221 vdd.n2618 gnd 0.179924f
C3222 vdd.n2619 gnd 0.005568f
C3223 vdd.n2620 gnd 0.005568f
C3224 vdd.n2621 gnd 0.005568f
C3225 vdd.n2622 gnd 0.005568f
C3226 vdd.n2623 gnd 0.005568f
C3227 vdd.n2624 gnd 0.005568f
C3228 vdd.n2625 gnd 0.005568f
C3229 vdd.n2626 gnd 0.005568f
C3230 vdd.n2627 gnd 0.005568f
C3231 vdd.n2628 gnd 0.005568f
C3232 vdd.n2629 gnd 0.005568f
C3233 vdd.n2630 gnd 0.355664f
C3234 vdd.n2631 gnd 0.005568f
C3235 vdd.n2632 gnd 0.005568f
C3236 vdd.n2633 gnd 0.005568f
C3237 vdd.n2634 gnd 0.011923f
C3238 vdd.n2635 gnd 0.011923f
C3239 vdd.n2636 gnd 0.012644f
C3240 vdd.n2637 gnd 0.012644f
C3241 vdd.n2638 gnd 0.005568f
C3242 vdd.n2639 gnd 0.005568f
C3243 vdd.n2640 gnd 0.005568f
C3244 vdd.n2641 gnd 0.004299f
C3245 vdd.n2642 gnd 0.007958f
C3246 vdd.n2643 gnd 0.004053f
C3247 vdd.n2644 gnd 0.005568f
C3248 vdd.n2645 gnd 0.005568f
C3249 vdd.n2646 gnd 0.005568f
C3250 vdd.n2647 gnd 0.005568f
C3251 vdd.n2648 gnd 0.005568f
C3252 vdd.n2649 gnd 0.005568f
C3253 vdd.n2650 gnd 0.005568f
C3254 vdd.n2651 gnd 0.005568f
C3255 vdd.n2652 gnd 0.005568f
C3256 vdd.n2653 gnd 0.005568f
C3257 vdd.n2654 gnd 0.005568f
C3258 vdd.n2655 gnd 0.005568f
C3259 vdd.n2656 gnd 0.005568f
C3260 vdd.n2657 gnd 0.005568f
C3261 vdd.n2658 gnd 0.005568f
C3262 vdd.n2659 gnd 0.005568f
C3263 vdd.n2660 gnd 0.005568f
C3264 vdd.n2661 gnd 0.005568f
C3265 vdd.n2662 gnd 0.005568f
C3266 vdd.n2663 gnd 0.005568f
C3267 vdd.n2664 gnd 0.005568f
C3268 vdd.n2665 gnd 0.005568f
C3269 vdd.n2666 gnd 0.005568f
C3270 vdd.n2667 gnd 0.005568f
C3271 vdd.n2668 gnd 0.005568f
C3272 vdd.n2669 gnd 0.005568f
C3273 vdd.n2670 gnd 0.005568f
C3274 vdd.n2671 gnd 0.005568f
C3275 vdd.n2672 gnd 0.005568f
C3276 vdd.n2673 gnd 0.005568f
C3277 vdd.n2674 gnd 0.005568f
C3278 vdd.n2675 gnd 0.005568f
C3279 vdd.n2676 gnd 0.005568f
C3280 vdd.n2677 gnd 0.005568f
C3281 vdd.n2678 gnd 0.005568f
C3282 vdd.n2679 gnd 0.005568f
C3283 vdd.n2680 gnd 0.005568f
C3284 vdd.n2681 gnd 0.005568f
C3285 vdd.n2682 gnd 0.005568f
C3286 vdd.n2683 gnd 0.005568f
C3287 vdd.n2684 gnd 0.005568f
C3288 vdd.n2685 gnd 0.005568f
C3289 vdd.n2686 gnd 0.005568f
C3290 vdd.n2687 gnd 0.005568f
C3291 vdd.n2688 gnd 0.005568f
C3292 vdd.n2689 gnd 0.005568f
C3293 vdd.n2690 gnd 0.005568f
C3294 vdd.n2691 gnd 0.005568f
C3295 vdd.n2692 gnd 0.005568f
C3296 vdd.n2693 gnd 0.005568f
C3297 vdd.n2694 gnd 0.005568f
C3298 vdd.n2695 gnd 0.005568f
C3299 vdd.n2696 gnd 0.005568f
C3300 vdd.n2697 gnd 0.005568f
C3301 vdd.n2698 gnd 0.005568f
C3302 vdd.n2699 gnd 0.005568f
C3303 vdd.n2700 gnd 0.005568f
C3304 vdd.n2701 gnd 0.005568f
C3305 vdd.n2702 gnd 0.694591f
C3306 vdd.n2704 gnd 0.012644f
C3307 vdd.n2705 gnd 0.012644f
C3308 vdd.n2706 gnd 0.011923f
C3309 vdd.n2707 gnd 0.005568f
C3310 vdd.n2708 gnd 0.005568f
C3311 vdd.n2709 gnd 0.334743f
C3312 vdd.n2710 gnd 0.005568f
C3313 vdd.n2711 gnd 0.005568f
C3314 vdd.n2712 gnd 0.005568f
C3315 vdd.n2713 gnd 0.005568f
C3316 vdd.n2714 gnd 0.005568f
C3317 vdd.n2715 gnd 0.338927f
C3318 vdd.n2716 gnd 0.005568f
C3319 vdd.n2717 gnd 0.005568f
C3320 vdd.n2718 gnd 0.005568f
C3321 vdd.n2719 gnd 0.005568f
C3322 vdd.n2720 gnd 0.005568f
C3323 vdd.n2721 gnd 0.569063f
C3324 vdd.n2722 gnd 0.005568f
C3325 vdd.n2723 gnd 0.005568f
C3326 vdd.n2724 gnd 0.005568f
C3327 vdd.n2725 gnd 0.005568f
C3328 vdd.n2726 gnd 0.005568f
C3329 vdd.n2727 gnd 0.41006f
C3330 vdd.n2728 gnd 0.005568f
C3331 vdd.n2729 gnd 0.005568f
C3332 vdd.n2730 gnd 0.005568f
C3333 vdd.n2731 gnd 0.005568f
C3334 vdd.n2732 gnd 0.005568f
C3335 vdd.n2733 gnd 0.514667f
C3336 vdd.n2734 gnd 0.005568f
C3337 vdd.n2735 gnd 0.005568f
C3338 vdd.n2736 gnd 0.005568f
C3339 vdd.n2737 gnd 0.005568f
C3340 vdd.n2738 gnd 0.005568f
C3341 vdd.n2739 gnd 0.422613f
C3342 vdd.n2740 gnd 0.005568f
C3343 vdd.n2741 gnd 0.005568f
C3344 vdd.n2742 gnd 0.005568f
C3345 vdd.n2743 gnd 0.005568f
C3346 vdd.n2744 gnd 0.005568f
C3347 vdd.n2745 gnd 0.297084f
C3348 vdd.n2746 gnd 0.005568f
C3349 vdd.n2747 gnd 0.005568f
C3350 vdd.n2748 gnd 0.005568f
C3351 vdd.n2749 gnd 0.005568f
C3352 vdd.n2750 gnd 0.005568f
C3353 vdd.n2751 gnd 0.179924f
C3354 vdd.n2752 gnd 0.005568f
C3355 vdd.n2753 gnd 0.005568f
C3356 vdd.n2754 gnd 0.005568f
C3357 vdd.n2755 gnd 0.005568f
C3358 vdd.n2756 gnd 0.005568f
C3359 vdd.n2757 gnd 0.523035f
C3360 vdd.n2758 gnd 0.005568f
C3361 vdd.n2759 gnd 0.005568f
C3362 vdd.n2760 gnd 0.005568f
C3363 vdd.n2761 gnd 0.003931f
C3364 vdd.n2762 gnd 0.005568f
C3365 vdd.n2763 gnd 0.005568f
C3366 vdd.n2764 gnd 0.569063f
C3367 vdd.n2765 gnd 0.005568f
C3368 vdd.n2766 gnd 0.005568f
C3369 vdd.n2767 gnd 0.005568f
C3370 vdd.n2768 gnd 0.005568f
C3371 vdd.n2769 gnd 0.005568f
C3372 vdd.n2770 gnd 0.451903f
C3373 vdd.n2771 gnd 0.005568f
C3374 vdd.n2772 gnd 0.004422f
C3375 vdd.n2773 gnd 0.005568f
C3376 vdd.n2774 gnd 0.005568f
C3377 vdd.n2775 gnd 0.005568f
C3378 vdd.n2776 gnd 0.364033f
C3379 vdd.n2777 gnd 0.005568f
C3380 vdd.n2778 gnd 0.005568f
C3381 vdd.n2779 gnd 0.005568f
C3382 vdd.n2780 gnd 0.005568f
C3383 vdd.n2781 gnd 0.005568f
C3384 vdd.n2782 gnd 0.330558f
C3385 vdd.n2783 gnd 0.005568f
C3386 vdd.n2784 gnd 0.005568f
C3387 vdd.n2785 gnd 0.005568f
C3388 vdd.n2786 gnd 0.005568f
C3389 vdd.n2787 gnd 0.005568f
C3390 vdd.n2788 gnd 0.456087f
C3391 vdd.n2789 gnd 0.005568f
C3392 vdd.n2790 gnd 0.005568f
C3393 vdd.n2791 gnd 0.005568f
C3394 vdd.n2792 gnd 0.005568f
C3395 vdd.n2793 gnd 0.005568f
C3396 vdd.n2794 gnd 0.569063f
C3397 vdd.n2795 gnd 0.005568f
C3398 vdd.n2796 gnd 0.005568f
C3399 vdd.n2797 gnd 0.005568f
C3400 vdd.n2798 gnd 0.005568f
C3401 vdd.n2799 gnd 0.005568f
C3402 vdd.n2800 gnd 0.55651f
C3403 vdd.n2801 gnd 0.005568f
C3404 vdd.n2802 gnd 0.005568f
C3405 vdd.n2803 gnd 0.005568f
C3406 vdd.n2804 gnd 0.005568f
C3407 vdd.n2805 gnd 0.005568f
C3408 vdd.n2806 gnd 0.430981f
C3409 vdd.n2807 gnd 0.005568f
C3410 vdd.n2808 gnd 0.005568f
C3411 vdd.n2809 gnd 0.005568f
C3412 vdd.n2810 gnd 0.005568f
C3413 vdd.n2811 gnd 0.005568f
C3414 vdd.n2812 gnd 0.305453f
C3415 vdd.n2813 gnd 0.005568f
C3416 vdd.n2814 gnd 0.005568f
C3417 vdd.n2815 gnd 0.005568f
C3418 vdd.n2816 gnd 0.005568f
C3419 vdd.n2817 gnd 0.005568f
C3420 vdd.n2818 gnd 0.569063f
C3421 vdd.n2819 gnd 0.005568f
C3422 vdd.n2820 gnd 0.005568f
C3423 vdd.n2821 gnd 0.005568f
C3424 vdd.n2822 gnd 0.005568f
C3425 vdd.n2823 gnd 0.005568f
C3426 vdd.n2824 gnd 0.005568f
C3427 vdd.n2826 gnd 0.005568f
C3428 vdd.n2827 gnd 0.005568f
C3429 vdd.n2829 gnd 0.005568f
C3430 vdd.n2830 gnd 0.005568f
C3431 vdd.n2833 gnd 0.005568f
C3432 vdd.n2834 gnd 0.005568f
C3433 vdd.n2835 gnd 0.005568f
C3434 vdd.n2836 gnd 0.005568f
C3435 vdd.n2838 gnd 0.005568f
C3436 vdd.n2839 gnd 0.005568f
C3437 vdd.n2840 gnd 0.005568f
C3438 vdd.n2841 gnd 0.005568f
C3439 vdd.n2842 gnd 0.005568f
C3440 vdd.n2843 gnd 0.005568f
C3441 vdd.n2845 gnd 0.005568f
C3442 vdd.n2846 gnd 0.005568f
C3443 vdd.n2847 gnd 0.005568f
C3444 vdd.n2848 gnd 0.005568f
C3445 vdd.n2849 gnd 0.005568f
C3446 vdd.n2850 gnd 0.005568f
C3447 vdd.n2852 gnd 0.005568f
C3448 vdd.n2853 gnd 0.005568f
C3449 vdd.n2854 gnd 0.005568f
C3450 vdd.n2855 gnd 0.005568f
C3451 vdd.n2856 gnd 0.005568f
C3452 vdd.n2857 gnd 0.005568f
C3453 vdd.n2859 gnd 0.005568f
C3454 vdd.n2860 gnd 0.012644f
C3455 vdd.n2861 gnd 0.012644f
C3456 vdd.n2862 gnd 0.011923f
C3457 vdd.n2863 gnd 0.005568f
C3458 vdd.n2864 gnd 0.005568f
C3459 vdd.n2865 gnd 0.005568f
C3460 vdd.n2866 gnd 0.005568f
C3461 vdd.n2867 gnd 0.005568f
C3462 vdd.n2868 gnd 0.005568f
C3463 vdd.n2869 gnd 0.569063f
C3464 vdd.n2870 gnd 0.005568f
C3465 vdd.n2871 gnd 0.005568f
C3466 vdd.n2872 gnd 0.005568f
C3467 vdd.n2873 gnd 0.005568f
C3468 vdd.n2874 gnd 0.005568f
C3469 vdd.n2875 gnd 0.405876f
C3470 vdd.n2876 gnd 0.005568f
C3471 vdd.n2877 gnd 0.005568f
C3472 vdd.n2878 gnd 0.005568f
C3473 vdd.n2879 gnd 0.012644f
C3474 vdd.n2880 gnd 0.011923f
C3475 vdd.n2881 gnd 0.012644f
C3476 vdd.n2883 gnd 0.005568f
C3477 vdd.n2884 gnd 0.005568f
C3478 vdd.n2885 gnd 0.004299f
C3479 vdd.n2886 gnd 0.007958f
C3480 vdd.n2887 gnd 0.004053f
C3481 vdd.n2888 gnd 0.005568f
C3482 vdd.n2889 gnd 0.005568f
C3483 vdd.n2891 gnd 0.005568f
C3484 vdd.n2892 gnd 0.005568f
C3485 vdd.n2893 gnd 0.005568f
C3486 vdd.n2894 gnd 0.005568f
C3487 vdd.n2895 gnd 0.005568f
C3488 vdd.n2896 gnd 0.005568f
C3489 vdd.n2898 gnd 0.005568f
C3490 vdd.n2899 gnd 0.005568f
C3491 vdd.n2900 gnd 0.005568f
C3492 vdd.n2901 gnd 0.005568f
C3493 vdd.n2902 gnd 0.005568f
C3494 vdd.n2903 gnd 0.005568f
C3495 vdd.n2905 gnd 0.005568f
C3496 vdd.n2906 gnd 0.005568f
C3497 vdd.n2907 gnd 0.005568f
C3498 vdd.n2908 gnd 0.005568f
C3499 vdd.n2909 gnd 0.005568f
C3500 vdd.n2910 gnd 0.005568f
C3501 vdd.n2912 gnd 0.005568f
C3502 vdd.n2913 gnd 0.005568f
C3503 vdd.n2914 gnd 0.005568f
C3504 vdd.n2916 gnd 0.005568f
C3505 vdd.n2917 gnd 0.005568f
C3506 vdd.n2918 gnd 0.005568f
C3507 vdd.n2919 gnd 0.005568f
C3508 vdd.n2920 gnd 0.005568f
C3509 vdd.n2921 gnd 0.005568f
C3510 vdd.n2923 gnd 0.005568f
C3511 vdd.n2924 gnd 0.005568f
C3512 vdd.n2925 gnd 0.005568f
C3513 vdd.n2926 gnd 0.005568f
C3514 vdd.n2927 gnd 0.005568f
C3515 vdd.n2928 gnd 0.005568f
C3516 vdd.n2930 gnd 0.005568f
C3517 vdd.n2931 gnd 0.005568f
C3518 vdd.n2932 gnd 0.005568f
C3519 vdd.n2933 gnd 0.005568f
C3520 vdd.n2934 gnd 0.005568f
C3521 vdd.n2935 gnd 0.005568f
C3522 vdd.n2937 gnd 0.005568f
C3523 vdd.n2938 gnd 0.005568f
C3524 vdd.n2940 gnd 0.005568f
C3525 vdd.n2941 gnd 0.005568f
C3526 vdd.n2942 gnd 0.012644f
C3527 vdd.n2943 gnd 0.011923f
C3528 vdd.n2944 gnd 0.011923f
C3529 vdd.n2945 gnd 0.769908f
C3530 vdd.n2946 gnd 0.011923f
C3531 vdd.n2947 gnd 0.012644f
C3532 vdd.n2948 gnd 0.011923f
C3533 vdd.n2949 gnd 0.005568f
C3534 vdd.n2950 gnd 0.004299f
C3535 vdd.n2951 gnd 0.005568f
C3536 vdd.n2953 gnd 0.005568f
C3537 vdd.n2954 gnd 0.005568f
C3538 vdd.n2955 gnd 0.005568f
C3539 vdd.n2956 gnd 0.005568f
C3540 vdd.n2957 gnd 0.005568f
C3541 vdd.n2958 gnd 0.005568f
C3542 vdd.n2960 gnd 0.005568f
C3543 vdd.n2961 gnd 0.005568f
C3544 vdd.n2962 gnd 0.005568f
C3545 vdd.n2963 gnd 0.005568f
C3546 vdd.n2964 gnd 0.005568f
C3547 vdd.n2965 gnd 0.005568f
C3548 vdd.n2967 gnd 0.005568f
C3549 vdd.n2968 gnd 0.005568f
C3550 vdd.n2969 gnd 0.005568f
C3551 vdd.n2970 gnd 0.005568f
C3552 vdd.n2971 gnd 0.005568f
C3553 vdd.n2972 gnd 0.005568f
C3554 vdd.n2974 gnd 0.005568f
C3555 vdd.n2975 gnd 0.005568f
C3556 vdd.n2977 gnd 0.005568f
C3557 vdd.n2978 gnd 0.034384f
C3558 vdd.n2979 gnd 0.872453f
C3559 vdd.n2980 gnd 0.007042f
C3560 vdd.n2981 gnd 0.020414f
C3561 vdd.n2982 gnd 0.003131f
C3562 vdd.t36 gnd 0.100744f
C3563 vdd.t37 gnd 0.107667f
C3564 vdd.t34 gnd 0.13157f
C3565 vdd.n2983 gnd 0.168654f
C3566 vdd.n2984 gnd 0.1417f
C3567 vdd.n2985 gnd 0.01015f
C3568 vdd.n2986 gnd 0.008189f
C3569 vdd.n2987 gnd 0.00346f
C3570 vdd.n2988 gnd 0.006591f
C3571 vdd.n2989 gnd 0.008189f
C3572 vdd.n2990 gnd 0.008189f
C3573 vdd.n2991 gnd 0.006591f
C3574 vdd.n2992 gnd 0.006591f
C3575 vdd.n2993 gnd 0.008189f
C3576 vdd.n2994 gnd 0.008189f
C3577 vdd.n2995 gnd 0.006591f
C3578 vdd.n2996 gnd 0.006591f
C3579 vdd.n2997 gnd 0.008189f
C3580 vdd.n2998 gnd 0.008189f
C3581 vdd.n2999 gnd 0.006591f
C3582 vdd.n3000 gnd 0.006591f
C3583 vdd.n3001 gnd 0.008189f
C3584 vdd.n3002 gnd 0.008189f
C3585 vdd.n3003 gnd 0.006591f
C3586 vdd.n3004 gnd 0.006591f
C3587 vdd.n3005 gnd 0.008189f
C3588 vdd.n3006 gnd 0.008189f
C3589 vdd.n3007 gnd 0.006591f
C3590 vdd.n3008 gnd 0.006591f
C3591 vdd.n3009 gnd 0.008189f
C3592 vdd.n3010 gnd 0.008189f
C3593 vdd.n3011 gnd 0.006591f
C3594 vdd.n3012 gnd 0.006591f
C3595 vdd.n3013 gnd 0.008189f
C3596 vdd.n3014 gnd 0.008189f
C3597 vdd.n3015 gnd 0.006591f
C3598 vdd.n3016 gnd 0.006591f
C3599 vdd.n3017 gnd 0.008189f
C3600 vdd.n3018 gnd 0.008189f
C3601 vdd.n3019 gnd 0.006591f
C3602 vdd.n3020 gnd 0.006591f
C3603 vdd.n3021 gnd 0.008189f
C3604 vdd.n3022 gnd 0.008189f
C3605 vdd.n3023 gnd 0.006591f
C3606 vdd.n3024 gnd 0.008189f
C3607 vdd.n3025 gnd 0.008189f
C3608 vdd.n3026 gnd 0.006591f
C3609 vdd.n3027 gnd 0.008189f
C3610 vdd.n3028 gnd 0.008189f
C3611 vdd.n3029 gnd 0.008189f
C3612 vdd.n3030 gnd 0.013446f
C3613 vdd.n3031 gnd 0.008189f
C3614 vdd.n3032 gnd 0.008189f
C3615 vdd.n3033 gnd 0.004482f
C3616 vdd.n3034 gnd 0.006591f
C3617 vdd.n3035 gnd 0.008189f
C3618 vdd.n3036 gnd 0.008189f
C3619 vdd.n3037 gnd 0.006591f
C3620 vdd.n3038 gnd 0.006591f
C3621 vdd.n3039 gnd 0.008189f
C3622 vdd.n3040 gnd 0.008189f
C3623 vdd.n3041 gnd 0.006591f
C3624 vdd.n3042 gnd 0.006591f
C3625 vdd.n3043 gnd 0.008189f
C3626 vdd.n3044 gnd 0.008189f
C3627 vdd.n3045 gnd 0.006591f
C3628 vdd.n3046 gnd 0.006591f
C3629 vdd.n3047 gnd 0.008189f
C3630 vdd.n3048 gnd 0.008189f
C3631 vdd.n3049 gnd 0.006591f
C3632 vdd.n3050 gnd 0.006591f
C3633 vdd.n3051 gnd 0.008189f
C3634 vdd.n3052 gnd 0.008189f
C3635 vdd.n3053 gnd 0.006591f
C3636 vdd.n3054 gnd 0.006591f
C3637 vdd.n3055 gnd 0.008189f
C3638 vdd.n3056 gnd 0.008189f
C3639 vdd.n3057 gnd 0.006591f
C3640 vdd.n3058 gnd 0.006591f
C3641 vdd.n3059 gnd 0.008189f
C3642 vdd.n3060 gnd 0.008189f
C3643 vdd.n3061 gnd 0.006591f
C3644 vdd.n3062 gnd 0.006591f
C3645 vdd.n3063 gnd 0.008189f
C3646 vdd.n3064 gnd 0.008189f
C3647 vdd.n3065 gnd 0.006591f
C3648 vdd.n3066 gnd 0.006591f
C3649 vdd.n3067 gnd 0.008189f
C3650 vdd.n3068 gnd 0.008189f
C3651 vdd.n3069 gnd 0.006591f
C3652 vdd.n3070 gnd 0.008189f
C3653 vdd.n3071 gnd 0.008189f
C3654 vdd.n3072 gnd 0.006591f
C3655 vdd.n3073 gnd 0.008189f
C3656 vdd.n3074 gnd 0.008189f
C3657 vdd.n3075 gnd 0.008189f
C3658 vdd.t70 gnd 0.100744f
C3659 vdd.t71 gnd 0.107667f
C3660 vdd.t69 gnd 0.13157f
C3661 vdd.n3076 gnd 0.168654f
C3662 vdd.n3077 gnd 0.1417f
C3663 vdd.n3078 gnd 0.013446f
C3664 vdd.n3079 gnd 0.008189f
C3665 vdd.n3080 gnd 0.008189f
C3666 vdd.n3081 gnd 0.005503f
C3667 vdd.n3082 gnd 0.006591f
C3668 vdd.n3083 gnd 0.008189f
C3669 vdd.n3084 gnd 0.008189f
C3670 vdd.n3085 gnd 0.006591f
C3671 vdd.n3086 gnd 0.006591f
C3672 vdd.n3087 gnd 0.008189f
C3673 vdd.n3088 gnd 0.008189f
C3674 vdd.n3089 gnd 0.006591f
C3675 vdd.n3090 gnd 0.006591f
C3676 vdd.n3091 gnd 0.008189f
C3677 vdd.n3092 gnd 0.008189f
C3678 vdd.n3093 gnd 0.006591f
C3679 vdd.n3094 gnd 0.006591f
C3680 vdd.n3095 gnd 0.008189f
C3681 vdd.n3096 gnd 0.008189f
C3682 vdd.n3097 gnd 0.006591f
C3683 vdd.n3098 gnd 0.006591f
C3684 vdd.n3099 gnd 0.008189f
C3685 vdd.n3100 gnd 0.008189f
C3686 vdd.n3101 gnd 0.006591f
C3687 vdd.n3102 gnd 0.006591f
C3688 vdd.n3103 gnd 0.008189f
C3689 vdd.n3104 gnd 0.008189f
C3690 vdd.n3105 gnd 0.006591f
C3691 vdd.n3106 gnd 0.006591f
C3692 vdd.n3108 gnd 0.872453f
C3693 vdd.n3110 gnd 0.006591f
C3694 vdd.n3111 gnd 0.008189f
C3695 vdd.n3112 gnd 10.2348f
C3696 vdd.n3114 gnd 0.020414f
C3697 vdd.n3115 gnd 0.005471f
C3698 vdd.n3116 gnd 0.020414f
C3699 vdd.n3117 gnd 0.019956f
C3700 vdd.n3118 gnd 0.008189f
C3701 vdd.n3119 gnd 0.006591f
C3702 vdd.n3120 gnd 0.008189f
C3703 vdd.n3121 gnd 0.523035f
C3704 vdd.n3122 gnd 0.008189f
C3705 vdd.n3123 gnd 0.006591f
C3706 vdd.n3124 gnd 0.008189f
C3707 vdd.n3125 gnd 0.008189f
C3708 vdd.n3126 gnd 0.008189f
C3709 vdd.n3127 gnd 0.006591f
C3710 vdd.n3128 gnd 0.008189f
C3711 vdd.n3129 gnd 0.665301f
C3712 vdd.n3130 gnd 0.836857f
C3713 vdd.n3131 gnd 0.008189f
C3714 vdd.n3132 gnd 0.006591f
C3715 vdd.n3133 gnd 0.008189f
C3716 vdd.n3134 gnd 0.008189f
C3717 vdd.n3135 gnd 0.008189f
C3718 vdd.n3136 gnd 0.006591f
C3719 vdd.n3137 gnd 0.008189f
C3720 vdd.n3138 gnd 0.589984f
C3721 vdd.n3139 gnd 0.008189f
C3722 vdd.n3140 gnd 0.006591f
C3723 vdd.n3141 gnd 0.008189f
C3724 vdd.n3142 gnd 0.008189f
C3725 vdd.n3143 gnd 0.008189f
C3726 vdd.n3144 gnd 0.006591f
C3727 vdd.n3145 gnd 0.008189f
C3728 vdd.t100 gnd 0.418428f
C3729 vdd.n3146 gnd 0.694591f
C3730 vdd.n3147 gnd 0.008189f
C3731 vdd.n3148 gnd 0.006591f
C3732 vdd.n3149 gnd 0.008189f
C3733 vdd.n3150 gnd 0.008189f
C3734 vdd.n3151 gnd 0.008189f
C3735 vdd.n3152 gnd 0.006591f
C3736 vdd.n3153 gnd 0.008189f
C3737 vdd.n3154 gnd 0.656933f
C3738 vdd.n3155 gnd 0.008189f
C3739 vdd.n3156 gnd 0.006591f
C3740 vdd.n3157 gnd 0.008189f
C3741 vdd.n3158 gnd 0.008189f
C3742 vdd.n3159 gnd 0.008189f
C3743 vdd.n3160 gnd 0.006591f
C3744 vdd.n3161 gnd 0.006591f
C3745 vdd.n3162 gnd 0.006591f
C3746 vdd.n3163 gnd 0.008189f
C3747 vdd.n3164 gnd 0.008189f
C3748 vdd.n3165 gnd 0.008189f
C3749 vdd.n3166 gnd 0.006591f
C3750 vdd.n3167 gnd 0.006591f
C3751 vdd.n3168 gnd 0.006591f
C3752 vdd.n3169 gnd 0.008189f
C3753 vdd.n3170 gnd 0.008189f
C3754 vdd.n3171 gnd 0.008189f
C3755 vdd.n3172 gnd 0.006591f
C3756 vdd.n3173 gnd 0.006591f
C3757 vdd.n3174 gnd 0.005471f
C3758 vdd.n3175 gnd 0.019956f
C3759 vdd.n3176 gnd 0.020414f
C3760 vdd.n3178 gnd 0.020414f
C3761 vdd.n3179 gnd 0.003131f
C3762 vdd.t52 gnd 0.100744f
C3763 vdd.t51 gnd 0.107667f
C3764 vdd.t49 gnd 0.13157f
C3765 vdd.n3180 gnd 0.168654f
C3766 vdd.n3181 gnd 0.142359f
C3767 vdd.n3182 gnd 0.010809f
C3768 vdd.n3183 gnd 0.00346f
C3769 vdd.n3184 gnd 0.006591f
C3770 vdd.n3185 gnd 0.008189f
C3771 vdd.n3187 gnd 0.008189f
C3772 vdd.n3188 gnd 0.008189f
C3773 vdd.n3189 gnd 0.006591f
C3774 vdd.n3190 gnd 0.006591f
C3775 vdd.n3191 gnd 0.006591f
C3776 vdd.n3192 gnd 0.008189f
C3777 vdd.n3194 gnd 0.008189f
C3778 vdd.n3195 gnd 0.008189f
C3779 vdd.n3196 gnd 0.006591f
C3780 vdd.n3197 gnd 0.006591f
C3781 vdd.n3198 gnd 0.006591f
C3782 vdd.n3199 gnd 0.008189f
C3783 vdd.n3201 gnd 0.008189f
C3784 vdd.n3202 gnd 0.008189f
C3785 vdd.n3203 gnd 0.006591f
C3786 vdd.n3204 gnd 0.006591f
C3787 vdd.n3205 gnd 0.006591f
C3788 vdd.n3206 gnd 0.008189f
C3789 vdd.n3208 gnd 0.008189f
C3790 vdd.n3209 gnd 0.008189f
C3791 vdd.n3210 gnd 0.006591f
C3792 vdd.n3211 gnd 0.006591f
C3793 vdd.n3212 gnd 0.006591f
C3794 vdd.n3213 gnd 0.008189f
C3795 vdd.n3215 gnd 0.008189f
C3796 vdd.n3216 gnd 0.008189f
C3797 vdd.n3217 gnd 0.006591f
C3798 vdd.n3218 gnd 0.008189f
C3799 vdd.n3219 gnd 0.008189f
C3800 vdd.n3220 gnd 0.008189f
C3801 vdd.n3221 gnd 0.014105f
C3802 vdd.n3222 gnd 0.004482f
C3803 vdd.n3223 gnd 0.006591f
C3804 vdd.n3224 gnd 0.008189f
C3805 vdd.n3226 gnd 0.008189f
C3806 vdd.n3227 gnd 0.008189f
C3807 vdd.n3228 gnd 0.006591f
C3808 vdd.n3229 gnd 0.006591f
C3809 vdd.n3230 gnd 0.006591f
C3810 vdd.n3231 gnd 0.008189f
C3811 vdd.n3233 gnd 0.008189f
C3812 vdd.n3234 gnd 0.008189f
C3813 vdd.n3235 gnd 0.006591f
C3814 vdd.n3236 gnd 0.006591f
C3815 vdd.n3237 gnd 0.006591f
C3816 vdd.n3238 gnd 0.008189f
C3817 vdd.n3240 gnd 0.008189f
C3818 vdd.n3241 gnd 0.008189f
C3819 vdd.n3242 gnd 0.006591f
C3820 vdd.n3243 gnd 0.006591f
C3821 vdd.n3244 gnd 0.006591f
C3822 vdd.n3245 gnd 0.008189f
C3823 vdd.n3247 gnd 0.008189f
C3824 vdd.n3248 gnd 0.008189f
C3825 vdd.n3249 gnd 0.006591f
C3826 vdd.n3250 gnd 0.006591f
C3827 vdd.n3251 gnd 0.006591f
C3828 vdd.n3252 gnd 0.008189f
C3829 vdd.n3254 gnd 0.008189f
C3830 vdd.n3255 gnd 0.008189f
C3831 vdd.n3256 gnd 0.006591f
C3832 vdd.n3257 gnd 0.008189f
C3833 vdd.n3258 gnd 0.008189f
C3834 vdd.n3259 gnd 0.008189f
C3835 vdd.n3260 gnd 0.014105f
C3836 vdd.n3261 gnd 0.005503f
C3837 vdd.n3262 gnd 0.006591f
C3838 vdd.n3263 gnd 0.008189f
C3839 vdd.n3265 gnd 0.008189f
C3840 vdd.n3266 gnd 0.008189f
C3841 vdd.n3267 gnd 0.006591f
C3842 vdd.n3268 gnd 0.006591f
C3843 vdd.n3269 gnd 0.006591f
C3844 vdd.n3270 gnd 0.008189f
C3845 vdd.n3272 gnd 0.008189f
C3846 vdd.n3273 gnd 0.008189f
C3847 vdd.n3274 gnd 0.006591f
C3848 vdd.n3275 gnd 0.006591f
C3849 vdd.n3276 gnd 0.006591f
C3850 vdd.n3277 gnd 0.008189f
C3851 vdd.n3279 gnd 0.008189f
C3852 vdd.n3280 gnd 0.008189f
C3853 vdd.n3281 gnd 0.006591f
C3854 vdd.n3282 gnd 0.006591f
C3855 vdd.n3283 gnd 0.006591f
C3856 vdd.n3284 gnd 0.008189f
C3857 vdd.n3286 gnd 0.008189f
C3858 vdd.n3287 gnd 0.008189f
C3859 vdd.n3289 gnd 0.008189f
C3860 vdd.n3290 gnd 0.006591f
C3861 vdd.n3291 gnd 0.006591f
C3862 vdd.n3292 gnd 0.005471f
C3863 vdd.n3293 gnd 0.020414f
C3864 vdd.n3294 gnd 0.019956f
C3865 vdd.n3295 gnd 0.005471f
C3866 vdd.n3296 gnd 0.019956f
C3867 vdd.n3297 gnd 1.23436f
C3868 vdd.t50 gnd 0.418428f
C3869 vdd.n3298 gnd 0.43935f
C3870 vdd.n3299 gnd 0.836857f
C3871 vdd.n3300 gnd 0.008189f
C3872 vdd.n3301 gnd 0.006591f
C3873 vdd.n3302 gnd 0.006591f
C3874 vdd.n3303 gnd 0.006591f
C3875 vdd.n3304 gnd 0.008189f
C3876 vdd.n3305 gnd 0.748987f
C3877 vdd.t121 gnd 0.418428f
C3878 vdd.n3306 gnd 0.506298f
C3879 vdd.n3307 gnd 0.606721f
C3880 vdd.n3308 gnd 0.008189f
C3881 vdd.n3309 gnd 0.006591f
C3882 vdd.n3310 gnd 0.006591f
C3883 vdd.n3311 gnd 0.006591f
C3884 vdd.n3312 gnd 0.008189f
C3885 vdd.n3313 gnd 0.464456f
C3886 vdd.t98 gnd 0.418428f
C3887 vdd.n3314 gnd 0.694591f
C3888 vdd.t139 gnd 0.418428f
C3889 vdd.n3315 gnd 0.514667f
C3890 vdd.n3316 gnd 0.008189f
C3891 vdd.n3317 gnd 0.006591f
C3892 vdd.n3318 gnd 0.006294f
C3893 vdd.n3319 gnd 0.483007f
C3894 vdd.n3320 gnd 1.95578f
C3895 a_n2982_13878.n0 gnd 3.88594f
C3896 a_n2982_13878.n1 gnd 2.85743f
C3897 a_n2982_13878.n2 gnd 3.82475f
C3898 a_n2982_13878.n3 gnd 0.806598f
C3899 a_n2982_13878.n4 gnd 0.8066f
C3900 a_n2982_13878.n5 gnd 0.916876f
C3901 a_n2982_13878.n6 gnd 0.201555f
C3902 a_n2982_13878.n7 gnd 0.148449f
C3903 a_n2982_13878.n8 gnd 0.233314f
C3904 a_n2982_13878.n9 gnd 0.180209f
C3905 a_n2982_13878.n10 gnd 0.201555f
C3906 a_n2982_13878.n11 gnd 1.34265f
C3907 a_n2982_13878.n12 gnd 0.148449f
C3908 a_n2982_13878.n13 gnd 0.969982f
C3909 a_n2982_13878.n14 gnd 0.212423f
C3910 a_n2982_13878.n15 gnd 0.747657f
C3911 a_n2982_13878.n16 gnd 0.212423f
C3912 a_n2982_13878.n17 gnd 0.212423f
C3913 a_n2982_13878.n18 gnd 0.483791f
C3914 a_n2982_13878.n19 gnd 0.278519f
C3915 a_n2982_13878.n20 gnd 0.212423f
C3916 a_n2982_13878.n21 gnd 0.536897f
C3917 a_n2982_13878.n22 gnd 0.212423f
C3918 a_n2982_13878.n23 gnd 0.212423f
C3919 a_n2982_13878.n24 gnd 0.945129f
C3920 a_n2982_13878.n25 gnd 0.278519f
C3921 a_n2982_13878.n26 gnd 0.985614f
C3922 a_n2982_13878.n27 gnd 0.212423f
C3923 a_n2982_13878.n28 gnd 0.212423f
C3924 a_n2982_13878.n29 gnd 0.483791f
C3925 a_n2982_13878.n30 gnd 0.212423f
C3926 a_n2982_13878.n31 gnd 0.278519f
C3927 a_n2982_13878.n32 gnd 3.26746f
C3928 a_n2982_13878.n33 gnd 0.278518f
C3929 a_n2982_13878.n34 gnd 0.106212f
C3930 a_n2982_13878.n35 gnd 0.212423f
C3931 a_n2982_13878.n36 gnd 0.85592f
C3932 a_n2982_13878.n37 gnd 0.212423f
C3933 a_n2982_13878.n38 gnd 0.278519f
C3934 a_n2982_13878.n39 gnd 1.74886f
C3935 a_n2982_13878.n40 gnd 1.17841f
C3936 a_n2982_13878.n41 gnd 2.35355f
C3937 a_n2982_13878.n42 gnd 2.1518f
C3938 a_n2982_13878.n43 gnd 1.17841f
C3939 a_n2982_13878.n44 gnd 1.74886f
C3940 a_n2982_13878.n45 gnd 0.008523f
C3941 a_n2982_13878.n46 gnd 4.11e-19
C3942 a_n2982_13878.n48 gnd 0.008224f
C3943 a_n2982_13878.n49 gnd 0.011959f
C3944 a_n2982_13878.n50 gnd 0.004385f
C3945 a_n2982_13878.n51 gnd 0.008523f
C3946 a_n2982_13878.n52 gnd 4.11e-19
C3947 a_n2982_13878.n54 gnd 0.008224f
C3948 a_n2982_13878.n55 gnd 0.011959f
C3949 a_n2982_13878.n56 gnd 0.007912f
C3950 a_n2982_13878.n58 gnd 0.28176f
C3951 a_n2982_13878.n59 gnd 0.008523f
C3952 a_n2982_13878.n60 gnd 4.11e-19
C3953 a_n2982_13878.n62 gnd 0.008224f
C3954 a_n2982_13878.n63 gnd 0.011959f
C3955 a_n2982_13878.n64 gnd 0.007912f
C3956 a_n2982_13878.n66 gnd 0.28176f
C3957 a_n2982_13878.n67 gnd 0.008523f
C3958 a_n2982_13878.n68 gnd 4.11e-19
C3959 a_n2982_13878.n70 gnd 0.008224f
C3960 a_n2982_13878.n71 gnd 0.011959f
C3961 a_n2982_13878.n72 gnd 0.007912f
C3962 a_n2982_13878.n74 gnd 0.28176f
C3963 a_n2982_13878.n75 gnd 0.008224f
C3964 a_n2982_13878.n76 gnd 0.280611f
C3965 a_n2982_13878.n77 gnd 0.008224f
C3966 a_n2982_13878.n78 gnd 0.280611f
C3967 a_n2982_13878.n79 gnd 0.008224f
C3968 a_n2982_13878.n80 gnd 0.280611f
C3969 a_n2982_13878.n81 gnd 0.008224f
C3970 a_n2982_13878.n82 gnd 0.280611f
C3971 a_n2982_13878.n83 gnd 0.301308f
C3972 a_n2982_13878.t37 gnd 0.699618f
C3973 a_n2982_13878.t55 gnd 0.68535f
C3974 a_n2982_13878.t39 gnd 0.68535f
C3975 a_n2982_13878.t33 gnd 0.68535f
C3976 a_n2982_13878.n84 gnd 0.301188f
C3977 a_n2982_13878.t21 gnd 0.68535f
C3978 a_n2982_13878.t53 gnd 0.68535f
C3979 a_n2982_13878.t47 gnd 0.68535f
C3980 a_n2982_13878.n85 gnd 0.297497f
C3981 a_n2982_13878.t41 gnd 0.68535f
C3982 a_n2982_13878.t45 gnd 0.68535f
C3983 a_n2982_13878.t25 gnd 0.68535f
C3984 a_n2982_13878.t15 gnd 0.699618f
C3985 a_n2982_13878.t110 gnd 0.699618f
C3986 a_n2982_13878.t87 gnd 0.68535f
C3987 a_n2982_13878.t92 gnd 0.68535f
C3988 a_n2982_13878.t80 gnd 0.68535f
C3989 a_n2982_13878.n86 gnd 0.301188f
C3990 a_n2982_13878.t97 gnd 0.68535f
C3991 a_n2982_13878.t106 gnd 0.68535f
C3992 a_n2982_13878.t107 gnd 0.68535f
C3993 a_n2982_13878.n87 gnd 0.297497f
C3994 a_n2982_13878.t74 gnd 0.68535f
C3995 a_n2982_13878.t89 gnd 0.68535f
C3996 a_n2982_13878.t77 gnd 0.68535f
C3997 a_n2982_13878.n88 gnd 0.301308f
C3998 a_n2982_13878.t84 gnd 0.68535f
C3999 a_n2982_13878.t103 gnd 0.696376f
C4000 a_n2982_13878.t18 gnd 1.37961f
C4001 a_n2982_13878.t60 gnd 0.147339f
C4002 a_n2982_13878.t28 gnd 0.147339f
C4003 a_n2982_13878.n89 gnd 1.03786f
C4004 a_n2982_13878.t62 gnd 0.147339f
C4005 a_n2982_13878.t44 gnd 0.147339f
C4006 a_n2982_13878.n90 gnd 1.03786f
C4007 a_n2982_13878.t52 gnd 0.147339f
C4008 a_n2982_13878.t20 gnd 0.147339f
C4009 a_n2982_13878.n91 gnd 1.03786f
C4010 a_n2982_13878.t58 gnd 0.147339f
C4011 a_n2982_13878.t36 gnd 0.147339f
C4012 a_n2982_13878.n92 gnd 1.03786f
C4013 a_n2982_13878.t50 gnd 0.147339f
C4014 a_n2982_13878.t30 gnd 0.147339f
C4015 a_n2982_13878.n93 gnd 1.03786f
C4016 a_n2982_13878.t24 gnd 1.37686f
C4017 a_n2982_13878.t49 gnd 0.68535f
C4018 a_n2982_13878.n94 gnd 0.301308f
C4019 a_n2982_13878.t29 gnd 0.68535f
C4020 a_n2982_13878.t57 gnd 0.68535f
C4021 a_n2982_13878.n95 gnd 0.292258f
C4022 a_n2982_13878.t43 gnd 0.68535f
C4023 a_n2982_13878.n96 gnd 0.303898f
C4024 a_n2982_13878.t51 gnd 0.68535f
C4025 a_n2982_13878.t27 gnd 0.68535f
C4026 a_n2982_13878.n97 gnd 0.297169f
C4027 a_n2982_13878.t17 gnd 0.699618f
C4028 a_n2982_13878.t86 gnd 0.68535f
C4029 a_n2982_13878.n98 gnd 0.301308f
C4030 a_n2982_13878.t96 gnd 0.68535f
C4031 a_n2982_13878.t101 gnd 0.68535f
C4032 a_n2982_13878.n99 gnd 0.292258f
C4033 a_n2982_13878.t105 gnd 0.68535f
C4034 a_n2982_13878.n100 gnd 0.303898f
C4035 a_n2982_13878.t76 gnd 0.68535f
C4036 a_n2982_13878.t79 gnd 0.68535f
C4037 a_n2982_13878.n101 gnd 0.297169f
C4038 a_n2982_13878.t109 gnd 0.699618f
C4039 a_n2982_13878.t78 gnd 0.68535f
C4040 a_n2982_13878.n102 gnd 0.303453f
C4041 a_n2982_13878.t104 gnd 0.68535f
C4042 a_n2982_13878.n103 gnd 0.301188f
C4043 a_n2982_13878.n104 gnd 0.301323f
C4044 a_n2982_13878.t100 gnd 0.68535f
C4045 a_n2982_13878.n105 gnd 0.297497f
C4046 a_n2982_13878.t73 gnd 0.68535f
C4047 a_n2982_13878.n106 gnd 0.297752f
C4048 a_n2982_13878.n107 gnd 0.303454f
C4049 a_n2982_13878.t75 gnd 0.696376f
C4050 a_n2982_13878.t59 gnd 0.68535f
C4051 a_n2982_13878.n108 gnd 0.303453f
C4052 a_n2982_13878.t61 gnd 0.68535f
C4053 a_n2982_13878.n109 gnd 0.301188f
C4054 a_n2982_13878.n110 gnd 0.301323f
C4055 a_n2982_13878.t19 gnd 0.68535f
C4056 a_n2982_13878.n111 gnd 0.297497f
C4057 a_n2982_13878.t35 gnd 0.68535f
C4058 a_n2982_13878.n112 gnd 0.297752f
C4059 a_n2982_13878.n113 gnd 0.303454f
C4060 a_n2982_13878.t23 gnd 0.696376f
C4061 a_n2982_13878.n114 gnd 1.32692f
C4062 a_n2982_13878.t83 gnd 0.68535f
C4063 a_n2982_13878.n115 gnd 0.297497f
C4064 a_n2982_13878.t91 gnd 0.68535f
C4065 a_n2982_13878.n116 gnd 0.297497f
C4066 a_n2982_13878.t81 gnd 0.68535f
C4067 a_n2982_13878.n117 gnd 0.297497f
C4068 a_n2982_13878.t95 gnd 0.68535f
C4069 a_n2982_13878.n118 gnd 0.297497f
C4070 a_n2982_13878.t85 gnd 0.68535f
C4071 a_n2982_13878.n119 gnd 0.292094f
C4072 a_n2982_13878.t111 gnd 0.68535f
C4073 a_n2982_13878.n120 gnd 0.301323f
C4074 a_n2982_13878.t88 gnd 0.696834f
C4075 a_n2982_13878.t98 gnd 0.68535f
C4076 a_n2982_13878.n121 gnd 0.292094f
C4077 a_n2982_13878.t82 gnd 0.68535f
C4078 a_n2982_13878.n122 gnd 0.301323f
C4079 a_n2982_13878.t93 gnd 0.696834f
C4080 a_n2982_13878.t102 gnd 0.68535f
C4081 a_n2982_13878.n123 gnd 0.292094f
C4082 a_n2982_13878.t90 gnd 0.68535f
C4083 a_n2982_13878.n124 gnd 0.301323f
C4084 a_n2982_13878.t108 gnd 0.696834f
C4085 a_n2982_13878.t94 gnd 0.68535f
C4086 a_n2982_13878.n125 gnd 0.292094f
C4087 a_n2982_13878.t72 gnd 0.68535f
C4088 a_n2982_13878.n126 gnd 0.301323f
C4089 a_n2982_13878.t99 gnd 0.696834f
C4090 a_n2982_13878.n127 gnd 1.6691f
C4091 a_n2982_13878.n128 gnd 0.303454f
C4092 a_n2982_13878.n129 gnd 0.297752f
C4093 a_n2982_13878.n130 gnd 0.292258f
C4094 a_n2982_13878.n131 gnd 0.301323f
C4095 a_n2982_13878.n132 gnd 0.303898f
C4096 a_n2982_13878.n133 gnd 0.297169f
C4097 a_n2982_13878.n134 gnd 0.303453f
C4098 a_n2982_13878.t31 gnd 0.68535f
C4099 a_n2982_13878.n135 gnd 0.303454f
C4100 a_n2982_13878.t14 gnd 0.114597f
C4101 a_n2982_13878.t1 gnd 0.114597f
C4102 a_n2982_13878.n136 gnd 1.01487f
C4103 a_n2982_13878.t66 gnd 0.114597f
C4104 a_n2982_13878.t3 gnd 0.114597f
C4105 a_n2982_13878.n137 gnd 1.01262f
C4106 a_n2982_13878.t69 gnd 0.114597f
C4107 a_n2982_13878.t10 gnd 0.114597f
C4108 a_n2982_13878.n138 gnd 1.01262f
C4109 a_n2982_13878.t70 gnd 0.114597f
C4110 a_n2982_13878.t11 gnd 0.114597f
C4111 a_n2982_13878.n139 gnd 1.01487f
C4112 a_n2982_13878.t12 gnd 0.114597f
C4113 a_n2982_13878.t8 gnd 0.114597f
C4114 a_n2982_13878.n140 gnd 1.01262f
C4115 a_n2982_13878.t9 gnd 0.114597f
C4116 a_n2982_13878.t5 gnd 0.114597f
C4117 a_n2982_13878.n141 gnd 1.01262f
C4118 a_n2982_13878.t63 gnd 0.114597f
C4119 a_n2982_13878.t2 gnd 0.114597f
C4120 a_n2982_13878.n142 gnd 1.01262f
C4121 a_n2982_13878.t68 gnd 0.114597f
C4122 a_n2982_13878.t65 gnd 0.114597f
C4123 a_n2982_13878.n143 gnd 1.01262f
C4124 a_n2982_13878.t67 gnd 0.114597f
C4125 a_n2982_13878.t6 gnd 0.114597f
C4126 a_n2982_13878.n144 gnd 1.01262f
C4127 a_n2982_13878.t71 gnd 0.114597f
C4128 a_n2982_13878.t4 gnd 0.114597f
C4129 a_n2982_13878.n145 gnd 1.01487f
C4130 a_n2982_13878.t7 gnd 0.114597f
C4131 a_n2982_13878.t0 gnd 0.114597f
C4132 a_n2982_13878.n146 gnd 1.01262f
C4133 a_n2982_13878.t13 gnd 0.114597f
C4134 a_n2982_13878.t64 gnd 0.114597f
C4135 a_n2982_13878.n147 gnd 1.01262f
C4136 a_n2982_13878.n148 gnd 0.30128f
C4137 a_n2982_13878.n149 gnd 0.292258f
C4138 a_n2982_13878.n150 gnd 0.301323f
C4139 a_n2982_13878.n151 gnd 0.303898f
C4140 a_n2982_13878.n152 gnd 0.297169f
C4141 a_n2982_13878.n153 gnd 0.303453f
C4142 a_n2982_13878.n154 gnd 1.00893f
C4143 a_n2982_13878.t38 gnd 1.37686f
C4144 a_n2982_13878.t56 gnd 0.147339f
C4145 a_n2982_13878.t40 gnd 0.147339f
C4146 a_n2982_13878.n155 gnd 1.03786f
C4147 a_n2982_13878.t34 gnd 0.147339f
C4148 a_n2982_13878.t22 gnd 0.147339f
C4149 a_n2982_13878.n156 gnd 1.03786f
C4150 a_n2982_13878.t54 gnd 0.147339f
C4151 a_n2982_13878.t48 gnd 0.147339f
C4152 a_n2982_13878.n157 gnd 1.03786f
C4153 a_n2982_13878.t42 gnd 0.147339f
C4154 a_n2982_13878.t46 gnd 0.147339f
C4155 a_n2982_13878.n158 gnd 1.03786f
C4156 a_n2982_13878.t26 gnd 0.147339f
C4157 a_n2982_13878.t32 gnd 0.147339f
C4158 a_n2982_13878.n159 gnd 1.03786f
C4159 a_n2982_13878.t16 gnd 1.37961f
C4160 CSoutput.n0 gnd 0.037861f
C4161 CSoutput.t150 gnd 0.250445f
C4162 CSoutput.n1 gnd 0.113088f
C4163 CSoutput.n2 gnd 0.037861f
C4164 CSoutput.t157 gnd 0.250445f
C4165 CSoutput.n3 gnd 0.030008f
C4166 CSoutput.n4 gnd 0.037861f
C4167 CSoutput.t164 gnd 0.250445f
C4168 CSoutput.n5 gnd 0.025876f
C4169 CSoutput.n6 gnd 0.037861f
C4170 CSoutput.t155 gnd 0.250445f
C4171 CSoutput.t153 gnd 0.250445f
C4172 CSoutput.n7 gnd 0.111856f
C4173 CSoutput.n8 gnd 0.037861f
C4174 CSoutput.t162 gnd 0.250445f
C4175 CSoutput.n9 gnd 0.024672f
C4176 CSoutput.n10 gnd 0.037861f
C4177 CSoutput.t145 gnd 0.250445f
C4178 CSoutput.t149 gnd 0.250445f
C4179 CSoutput.n11 gnd 0.111856f
C4180 CSoutput.n12 gnd 0.037861f
C4181 CSoutput.t160 gnd 0.250445f
C4182 CSoutput.n13 gnd 0.025876f
C4183 CSoutput.n14 gnd 0.037861f
C4184 CSoutput.t159 gnd 0.250445f
C4185 CSoutput.t147 gnd 0.250445f
C4186 CSoutput.n15 gnd 0.111856f
C4187 CSoutput.n16 gnd 0.037861f
C4188 CSoutput.t152 gnd 0.250445f
C4189 CSoutput.n17 gnd 0.027637f
C4190 CSoutput.t161 gnd 0.299288f
C4191 CSoutput.t158 gnd 0.250445f
C4192 CSoutput.n18 gnd 0.142796f
C4193 CSoutput.n19 gnd 0.138562f
C4194 CSoutput.n20 gnd 0.160748f
C4195 CSoutput.n21 gnd 0.037861f
C4196 CSoutput.n22 gnd 0.0316f
C4197 CSoutput.n23 gnd 0.111856f
C4198 CSoutput.n24 gnd 0.030461f
C4199 CSoutput.n25 gnd 0.030008f
C4200 CSoutput.n26 gnd 0.037861f
C4201 CSoutput.n27 gnd 0.037861f
C4202 CSoutput.n28 gnd 0.031357f
C4203 CSoutput.n29 gnd 0.026623f
C4204 CSoutput.n30 gnd 0.114346f
C4205 CSoutput.n31 gnd 0.026989f
C4206 CSoutput.n32 gnd 0.037861f
C4207 CSoutput.n33 gnd 0.037861f
C4208 CSoutput.n34 gnd 0.037861f
C4209 CSoutput.n35 gnd 0.031023f
C4210 CSoutput.n36 gnd 0.111856f
C4211 CSoutput.n37 gnd 0.029669f
C4212 CSoutput.n38 gnd 0.030801f
C4213 CSoutput.n39 gnd 0.037861f
C4214 CSoutput.n40 gnd 0.037861f
C4215 CSoutput.n41 gnd 0.031593f
C4216 CSoutput.n42 gnd 0.028876f
C4217 CSoutput.n43 gnd 0.111856f
C4218 CSoutput.n44 gnd 0.029608f
C4219 CSoutput.n45 gnd 0.037861f
C4220 CSoutput.n46 gnd 0.037861f
C4221 CSoutput.n47 gnd 0.037861f
C4222 CSoutput.n48 gnd 0.029608f
C4223 CSoutput.n49 gnd 0.111856f
C4224 CSoutput.n50 gnd 0.028876f
C4225 CSoutput.n51 gnd 0.031593f
C4226 CSoutput.n52 gnd 0.037861f
C4227 CSoutput.n53 gnd 0.037861f
C4228 CSoutput.n54 gnd 0.030801f
C4229 CSoutput.n55 gnd 0.029669f
C4230 CSoutput.n56 gnd 0.111856f
C4231 CSoutput.n57 gnd 0.031023f
C4232 CSoutput.n58 gnd 0.037861f
C4233 CSoutput.n59 gnd 0.037861f
C4234 CSoutput.n60 gnd 0.037861f
C4235 CSoutput.n61 gnd 0.026989f
C4236 CSoutput.n62 gnd 0.114346f
C4237 CSoutput.n63 gnd 0.026623f
C4238 CSoutput.t156 gnd 0.250445f
C4239 CSoutput.n64 gnd 0.111856f
C4240 CSoutput.n65 gnd 0.031357f
C4241 CSoutput.n66 gnd 0.037861f
C4242 CSoutput.n67 gnd 0.037861f
C4243 CSoutput.n68 gnd 0.037861f
C4244 CSoutput.n69 gnd 0.030461f
C4245 CSoutput.n70 gnd 0.111856f
C4246 CSoutput.n71 gnd 0.0316f
C4247 CSoutput.n72 gnd 0.027637f
C4248 CSoutput.n73 gnd 0.037861f
C4249 CSoutput.n74 gnd 0.037861f
C4250 CSoutput.n75 gnd 0.028662f
C4251 CSoutput.n76 gnd 0.017022f
C4252 CSoutput.t163 gnd 0.281393f
C4253 CSoutput.n77 gnd 0.139785f
C4254 CSoutput.n78 gnd 0.571852f
C4255 CSoutput.t7 gnd 0.047227f
C4256 CSoutput.t46 gnd 0.047227f
C4257 CSoutput.n79 gnd 0.365645f
C4258 CSoutput.t41 gnd 0.047227f
C4259 CSoutput.t37 gnd 0.047227f
C4260 CSoutput.n80 gnd 0.364993f
C4261 CSoutput.n81 gnd 0.370468f
C4262 CSoutput.t6 gnd 0.047227f
C4263 CSoutput.t15 gnd 0.047227f
C4264 CSoutput.n82 gnd 0.364993f
C4265 CSoutput.n83 gnd 0.182551f
C4266 CSoutput.t30 gnd 0.047227f
C4267 CSoutput.t2 gnd 0.047227f
C4268 CSoutput.n84 gnd 0.364993f
C4269 CSoutput.n85 gnd 0.334756f
C4270 CSoutput.t10 gnd 0.047227f
C4271 CSoutput.t44 gnd 0.047227f
C4272 CSoutput.n86 gnd 0.365645f
C4273 CSoutput.t13 gnd 0.047227f
C4274 CSoutput.t11 gnd 0.047227f
C4275 CSoutput.n87 gnd 0.364993f
C4276 CSoutput.n88 gnd 0.370468f
C4277 CSoutput.t47 gnd 0.047227f
C4278 CSoutput.t5 gnd 0.047227f
C4279 CSoutput.n89 gnd 0.364993f
C4280 CSoutput.n90 gnd 0.182551f
C4281 CSoutput.t12 gnd 0.047227f
C4282 CSoutput.t31 gnd 0.047227f
C4283 CSoutput.n91 gnd 0.364993f
C4284 CSoutput.n92 gnd 0.272229f
C4285 CSoutput.n93 gnd 0.343279f
C4286 CSoutput.t42 gnd 0.047227f
C4287 CSoutput.t25 gnd 0.047227f
C4288 CSoutput.n94 gnd 0.365645f
C4289 CSoutput.t19 gnd 0.047227f
C4290 CSoutput.t43 gnd 0.047227f
C4291 CSoutput.n95 gnd 0.364993f
C4292 CSoutput.n96 gnd 0.370468f
C4293 CSoutput.t4 gnd 0.047227f
C4294 CSoutput.t24 gnd 0.047227f
C4295 CSoutput.n97 gnd 0.364993f
C4296 CSoutput.n98 gnd 0.182551f
C4297 CSoutput.t18 gnd 0.047227f
C4298 CSoutput.t17 gnd 0.047227f
C4299 CSoutput.n99 gnd 0.364993f
C4300 CSoutput.n100 gnd 0.272229f
C4301 CSoutput.n101 gnd 0.383698f
C4302 CSoutput.n102 gnd 7.09833f
C4303 CSoutput.n104 gnd 0.669761f
C4304 CSoutput.n105 gnd 0.502321f
C4305 CSoutput.n106 gnd 0.669761f
C4306 CSoutput.n107 gnd 0.669761f
C4307 CSoutput.n108 gnd 1.8032f
C4308 CSoutput.n109 gnd 0.669761f
C4309 CSoutput.n110 gnd 0.669761f
C4310 CSoutput.t151 gnd 0.837201f
C4311 CSoutput.n111 gnd 0.669761f
C4312 CSoutput.n112 gnd 0.669761f
C4313 CSoutput.n116 gnd 0.669761f
C4314 CSoutput.n120 gnd 0.669761f
C4315 CSoutput.n121 gnd 0.669761f
C4316 CSoutput.n123 gnd 0.669761f
C4317 CSoutput.n128 gnd 0.669761f
C4318 CSoutput.n130 gnd 0.669761f
C4319 CSoutput.n131 gnd 0.669761f
C4320 CSoutput.n133 gnd 0.669761f
C4321 CSoutput.n134 gnd 0.669761f
C4322 CSoutput.n136 gnd 0.669761f
C4323 CSoutput.t146 gnd 11.1916f
C4324 CSoutput.n138 gnd 0.669761f
C4325 CSoutput.n139 gnd 0.502321f
C4326 CSoutput.n140 gnd 0.669761f
C4327 CSoutput.n141 gnd 0.669761f
C4328 CSoutput.n142 gnd 1.8032f
C4329 CSoutput.n143 gnd 0.669761f
C4330 CSoutput.n144 gnd 0.669761f
C4331 CSoutput.t165 gnd 0.837201f
C4332 CSoutput.n145 gnd 0.669761f
C4333 CSoutput.n146 gnd 0.669761f
C4334 CSoutput.n150 gnd 0.669761f
C4335 CSoutput.n154 gnd 0.669761f
C4336 CSoutput.n155 gnd 0.669761f
C4337 CSoutput.n157 gnd 0.669761f
C4338 CSoutput.n162 gnd 0.669761f
C4339 CSoutput.n164 gnd 0.669761f
C4340 CSoutput.n165 gnd 0.669761f
C4341 CSoutput.n167 gnd 0.669761f
C4342 CSoutput.n168 gnd 0.669761f
C4343 CSoutput.n170 gnd 0.669761f
C4344 CSoutput.n171 gnd 0.502321f
C4345 CSoutput.n173 gnd 0.669761f
C4346 CSoutput.n174 gnd 0.502321f
C4347 CSoutput.n175 gnd 0.669761f
C4348 CSoutput.n176 gnd 0.669761f
C4349 CSoutput.n177 gnd 1.8032f
C4350 CSoutput.n178 gnd 0.669761f
C4351 CSoutput.n179 gnd 0.669761f
C4352 CSoutput.t144 gnd 0.837201f
C4353 CSoutput.n180 gnd 0.669761f
C4354 CSoutput.n181 gnd 1.8032f
C4355 CSoutput.n183 gnd 0.669761f
C4356 CSoutput.n184 gnd 0.669761f
C4357 CSoutput.n186 gnd 0.669761f
C4358 CSoutput.n187 gnd 0.669761f
C4359 CSoutput.t154 gnd 11.009201f
C4360 CSoutput.t148 gnd 11.1916f
C4361 CSoutput.n193 gnd 2.10114f
C4362 CSoutput.n194 gnd 8.55928f
C4363 CSoutput.n195 gnd 8.91743f
C4364 CSoutput.n200 gnd 2.2761f
C4365 CSoutput.n206 gnd 0.669761f
C4366 CSoutput.n208 gnd 0.669761f
C4367 CSoutput.n210 gnd 0.669761f
C4368 CSoutput.n212 gnd 0.669761f
C4369 CSoutput.n214 gnd 0.669761f
C4370 CSoutput.n220 gnd 0.669761f
C4371 CSoutput.n227 gnd 1.22875f
C4372 CSoutput.n228 gnd 1.22875f
C4373 CSoutput.n229 gnd 0.669761f
C4374 CSoutput.n230 gnd 0.669761f
C4375 CSoutput.n232 gnd 0.502321f
C4376 CSoutput.n233 gnd 0.430193f
C4377 CSoutput.n235 gnd 0.502321f
C4378 CSoutput.n236 gnd 0.430193f
C4379 CSoutput.n237 gnd 0.502321f
C4380 CSoutput.n239 gnd 0.669761f
C4381 CSoutput.n241 gnd 1.8032f
C4382 CSoutput.n242 gnd 2.10114f
C4383 CSoutput.n243 gnd 7.87233f
C4384 CSoutput.n245 gnd 0.502321f
C4385 CSoutput.n246 gnd 1.2925f
C4386 CSoutput.n247 gnd 0.502321f
C4387 CSoutput.n249 gnd 0.669761f
C4388 CSoutput.n251 gnd 1.8032f
C4389 CSoutput.n252 gnd 3.92767f
C4390 CSoutput.t36 gnd 0.047227f
C4391 CSoutput.t23 gnd 0.047227f
C4392 CSoutput.n253 gnd 0.365645f
C4393 CSoutput.t28 gnd 0.047227f
C4394 CSoutput.t40 gnd 0.047227f
C4395 CSoutput.n254 gnd 0.364993f
C4396 CSoutput.n255 gnd 0.370468f
C4397 CSoutput.t14 gnd 0.047227f
C4398 CSoutput.t8 gnd 0.047227f
C4399 CSoutput.n256 gnd 0.364993f
C4400 CSoutput.n257 gnd 0.182551f
C4401 CSoutput.t21 gnd 0.047227f
C4402 CSoutput.t29 gnd 0.047227f
C4403 CSoutput.n258 gnd 0.364993f
C4404 CSoutput.n259 gnd 0.334756f
C4405 CSoutput.t38 gnd 0.047227f
C4406 CSoutput.t39 gnd 0.047227f
C4407 CSoutput.n260 gnd 0.365645f
C4408 CSoutput.t1 gnd 0.047227f
C4409 CSoutput.t20 gnd 0.047227f
C4410 CSoutput.n261 gnd 0.364993f
C4411 CSoutput.n262 gnd 0.370468f
C4412 CSoutput.t27 gnd 0.047227f
C4413 CSoutput.t0 gnd 0.047227f
C4414 CSoutput.n263 gnd 0.364993f
C4415 CSoutput.n264 gnd 0.182551f
C4416 CSoutput.t35 gnd 0.047227f
C4417 CSoutput.t16 gnd 0.047227f
C4418 CSoutput.n265 gnd 0.364993f
C4419 CSoutput.n266 gnd 0.272229f
C4420 CSoutput.n267 gnd 0.343279f
C4421 CSoutput.t33 gnd 0.047227f
C4422 CSoutput.t34 gnd 0.047227f
C4423 CSoutput.n268 gnd 0.365645f
C4424 CSoutput.t45 gnd 0.047227f
C4425 CSoutput.t26 gnd 0.047227f
C4426 CSoutput.n269 gnd 0.364993f
C4427 CSoutput.n270 gnd 0.370468f
C4428 CSoutput.t32 gnd 0.047227f
C4429 CSoutput.t9 gnd 0.047227f
C4430 CSoutput.n271 gnd 0.364993f
C4431 CSoutput.n272 gnd 0.182551f
C4432 CSoutput.t3 gnd 0.047227f
C4433 CSoutput.t22 gnd 0.047227f
C4434 CSoutput.n273 gnd 0.364992f
C4435 CSoutput.n274 gnd 0.27223f
C4436 CSoutput.n275 gnd 0.383698f
C4437 CSoutput.n276 gnd 10.141001f
C4438 CSoutput.t87 gnd 0.041323f
C4439 CSoutput.t140 gnd 0.041323f
C4440 CSoutput.n277 gnd 0.36637f
C4441 CSoutput.t81 gnd 0.041323f
C4442 CSoutput.t86 gnd 0.041323f
C4443 CSoutput.n278 gnd 0.365148f
C4444 CSoutput.n279 gnd 0.34025f
C4445 CSoutput.t71 gnd 0.041323f
C4446 CSoutput.t90 gnd 0.041323f
C4447 CSoutput.n280 gnd 0.365148f
C4448 CSoutput.n281 gnd 0.167727f
C4449 CSoutput.t105 gnd 0.041323f
C4450 CSoutput.t82 gnd 0.041323f
C4451 CSoutput.n282 gnd 0.365148f
C4452 CSoutput.n283 gnd 0.167727f
C4453 CSoutput.t89 gnd 0.041323f
C4454 CSoutput.t131 gnd 0.041323f
C4455 CSoutput.n284 gnd 0.365148f
C4456 CSoutput.n285 gnd 0.167727f
C4457 CSoutput.t101 gnd 0.041323f
C4458 CSoutput.t111 gnd 0.041323f
C4459 CSoutput.n286 gnd 0.365148f
C4460 CSoutput.n287 gnd 0.167727f
C4461 CSoutput.t66 gnd 0.041323f
C4462 CSoutput.t91 gnd 0.041323f
C4463 CSoutput.n288 gnd 0.365148f
C4464 CSoutput.n289 gnd 0.167727f
C4465 CSoutput.t55 gnd 0.041323f
C4466 CSoutput.t78 gnd 0.041323f
C4467 CSoutput.n290 gnd 0.365148f
C4468 CSoutput.n291 gnd 0.309364f
C4469 CSoutput.t136 gnd 0.041323f
C4470 CSoutput.t48 gnd 0.041323f
C4471 CSoutput.n292 gnd 0.36637f
C4472 CSoutput.t59 gnd 0.041323f
C4473 CSoutput.t129 gnd 0.041323f
C4474 CSoutput.n293 gnd 0.365148f
C4475 CSoutput.n294 gnd 0.34025f
C4476 CSoutput.t50 gnd 0.041323f
C4477 CSoutput.t122 gnd 0.041323f
C4478 CSoutput.n295 gnd 0.365148f
C4479 CSoutput.n296 gnd 0.167727f
C4480 CSoutput.t130 gnd 0.041323f
C4481 CSoutput.t49 gnd 0.041323f
C4482 CSoutput.n297 gnd 0.365148f
C4483 CSoutput.n298 gnd 0.167727f
C4484 CSoutput.t113 gnd 0.041323f
C4485 CSoutput.t94 gnd 0.041323f
C4486 CSoutput.n299 gnd 0.365148f
C4487 CSoutput.n300 gnd 0.167727f
C4488 CSoutput.t51 gnd 0.041323f
C4489 CSoutput.t115 gnd 0.041323f
C4490 CSoutput.n301 gnd 0.365148f
C4491 CSoutput.n302 gnd 0.167727f
C4492 CSoutput.t96 gnd 0.041323f
C4493 CSoutput.t102 gnd 0.041323f
C4494 CSoutput.n303 gnd 0.365148f
C4495 CSoutput.n304 gnd 0.167727f
C4496 CSoutput.t114 gnd 0.041323f
C4497 CSoutput.t95 gnd 0.041323f
C4498 CSoutput.n305 gnd 0.365148f
C4499 CSoutput.n306 gnd 0.254646f
C4500 CSoutput.n307 gnd 0.321187f
C4501 CSoutput.t60 gnd 0.041323f
C4502 CSoutput.t132 gnd 0.041323f
C4503 CSoutput.n308 gnd 0.36637f
C4504 CSoutput.t79 gnd 0.041323f
C4505 CSoutput.t83 gnd 0.041323f
C4506 CSoutput.n309 gnd 0.365148f
C4507 CSoutput.n310 gnd 0.34025f
C4508 CSoutput.t52 gnd 0.041323f
C4509 CSoutput.t117 gnd 0.041323f
C4510 CSoutput.n311 gnd 0.365148f
C4511 CSoutput.n312 gnd 0.167727f
C4512 CSoutput.t88 gnd 0.041323f
C4513 CSoutput.t61 gnd 0.041323f
C4514 CSoutput.n313 gnd 0.365148f
C4515 CSoutput.n314 gnd 0.167727f
C4516 CSoutput.t69 gnd 0.041323f
C4517 CSoutput.t143 gnd 0.041323f
C4518 CSoutput.n315 gnd 0.365148f
C4519 CSoutput.n316 gnd 0.167727f
C4520 CSoutput.t70 gnd 0.041323f
C4521 CSoutput.t74 gnd 0.041323f
C4522 CSoutput.n317 gnd 0.365148f
C4523 CSoutput.n318 gnd 0.167727f
C4524 CSoutput.t58 gnd 0.041323f
C4525 CSoutput.t128 gnd 0.041323f
C4526 CSoutput.n319 gnd 0.365148f
C4527 CSoutput.n320 gnd 0.167727f
C4528 CSoutput.t77 gnd 0.041323f
C4529 CSoutput.t67 gnd 0.041323f
C4530 CSoutput.n321 gnd 0.365148f
C4531 CSoutput.n322 gnd 0.254646f
C4532 CSoutput.n323 gnd 0.344905f
C4533 CSoutput.n324 gnd 10.4128f
C4534 CSoutput.t73 gnd 0.041323f
C4535 CSoutput.t116 gnd 0.041323f
C4536 CSoutput.n325 gnd 0.36637f
C4537 CSoutput.t112 gnd 0.041323f
C4538 CSoutput.t93 gnd 0.041323f
C4539 CSoutput.n326 gnd 0.365148f
C4540 CSoutput.n327 gnd 0.34025f
C4541 CSoutput.t119 gnd 0.041323f
C4542 CSoutput.t84 gnd 0.041323f
C4543 CSoutput.n328 gnd 0.365148f
C4544 CSoutput.n329 gnd 0.167727f
C4545 CSoutput.t103 gnd 0.041323f
C4546 CSoutput.t134 gnd 0.041323f
C4547 CSoutput.n330 gnd 0.365148f
C4548 CSoutput.n331 gnd 0.167727f
C4549 CSoutput.t68 gnd 0.041323f
C4550 CSoutput.t118 gnd 0.041323f
C4551 CSoutput.n332 gnd 0.365148f
C4552 CSoutput.n333 gnd 0.167727f
C4553 CSoutput.t57 gnd 0.041323f
C4554 CSoutput.t124 gnd 0.041323f
C4555 CSoutput.n334 gnd 0.365148f
C4556 CSoutput.n335 gnd 0.167727f
C4557 CSoutput.t123 gnd 0.041323f
C4558 CSoutput.t80 gnd 0.041323f
C4559 CSoutput.n336 gnd 0.365148f
C4560 CSoutput.n337 gnd 0.167727f
C4561 CSoutput.t99 gnd 0.041323f
C4562 CSoutput.t76 gnd 0.041323f
C4563 CSoutput.n338 gnd 0.365148f
C4564 CSoutput.n339 gnd 0.309364f
C4565 CSoutput.t63 gnd 0.041323f
C4566 CSoutput.t56 gnd 0.041323f
C4567 CSoutput.n340 gnd 0.36637f
C4568 CSoutput.t53 gnd 0.041323f
C4569 CSoutput.t141 gnd 0.041323f
C4570 CSoutput.n341 gnd 0.365148f
C4571 CSoutput.n342 gnd 0.34025f
C4572 CSoutput.t142 gnd 0.041323f
C4573 CSoutput.t64 gnd 0.041323f
C4574 CSoutput.n343 gnd 0.365148f
C4575 CSoutput.n344 gnd 0.167727f
C4576 CSoutput.t65 gnd 0.041323f
C4577 CSoutput.t107 gnd 0.041323f
C4578 CSoutput.n345 gnd 0.365148f
C4579 CSoutput.n346 gnd 0.167727f
C4580 CSoutput.t108 gnd 0.041323f
C4581 CSoutput.t135 gnd 0.041323f
C4582 CSoutput.n347 gnd 0.365148f
C4583 CSoutput.n348 gnd 0.167727f
C4584 CSoutput.t138 gnd 0.041323f
C4585 CSoutput.t127 gnd 0.041323f
C4586 CSoutput.n349 gnd 0.365148f
C4587 CSoutput.n350 gnd 0.167727f
C4588 CSoutput.t121 gnd 0.041323f
C4589 CSoutput.t109 gnd 0.041323f
C4590 CSoutput.n351 gnd 0.365148f
C4591 CSoutput.n352 gnd 0.167727f
C4592 CSoutput.t110 gnd 0.041323f
C4593 CSoutput.t139 gnd 0.041323f
C4594 CSoutput.n353 gnd 0.365148f
C4595 CSoutput.n354 gnd 0.254646f
C4596 CSoutput.n355 gnd 0.321187f
C4597 CSoutput.t100 gnd 0.041323f
C4598 CSoutput.t125 gnd 0.041323f
C4599 CSoutput.n356 gnd 0.36637f
C4600 CSoutput.t72 gnd 0.041323f
C4601 CSoutput.t85 gnd 0.041323f
C4602 CSoutput.n357 gnd 0.365148f
C4603 CSoutput.n358 gnd 0.34025f
C4604 CSoutput.t92 gnd 0.041323f
C4605 CSoutput.t106 gnd 0.041323f
C4606 CSoutput.n359 gnd 0.365148f
C4607 CSoutput.n360 gnd 0.167727f
C4608 CSoutput.t126 gnd 0.041323f
C4609 CSoutput.t97 gnd 0.041323f
C4610 CSoutput.n361 gnd 0.365148f
C4611 CSoutput.n362 gnd 0.167727f
C4612 CSoutput.t104 gnd 0.041323f
C4613 CSoutput.t137 gnd 0.041323f
C4614 CSoutput.n363 gnd 0.365148f
C4615 CSoutput.n364 gnd 0.167727f
C4616 CSoutput.t54 gnd 0.041323f
C4617 CSoutput.t75 gnd 0.041323f
C4618 CSoutput.n365 gnd 0.365148f
C4619 CSoutput.n366 gnd 0.167727f
C4620 CSoutput.t98 gnd 0.041323f
C4621 CSoutput.t120 gnd 0.041323f
C4622 CSoutput.n367 gnd 0.365148f
C4623 CSoutput.n368 gnd 0.167727f
C4624 CSoutput.t133 gnd 0.041323f
C4625 CSoutput.t62 gnd 0.041323f
C4626 CSoutput.n369 gnd 0.365148f
C4627 CSoutput.n370 gnd 0.254646f
C4628 CSoutput.n371 gnd 0.344905f
C4629 CSoutput.n372 gnd 6.0165f
C4630 CSoutput.n373 gnd 11.489f
C4631 commonsourceibias.n0 gnd 0.012624f
C4632 commonsourceibias.t120 gnd 0.191163f
C4633 commonsourceibias.t67 gnd 0.176757f
C4634 commonsourceibias.n1 gnd 0.00769f
C4635 commonsourceibias.n2 gnd 0.009461f
C4636 commonsourceibias.t126 gnd 0.176757f
C4637 commonsourceibias.n3 gnd 0.009597f
C4638 commonsourceibias.n4 gnd 0.009461f
C4639 commonsourceibias.t121 gnd 0.176757f
C4640 commonsourceibias.n5 gnd 0.070526f
C4641 commonsourceibias.t136 gnd 0.176757f
C4642 commonsourceibias.n6 gnd 0.007653f
C4643 commonsourceibias.n7 gnd 0.009461f
C4644 commonsourceibias.t117 gnd 0.176757f
C4645 commonsourceibias.n8 gnd 0.009134f
C4646 commonsourceibias.n9 gnd 0.009461f
C4647 commonsourceibias.t102 gnd 0.176757f
C4648 commonsourceibias.n10 gnd 0.070526f
C4649 commonsourceibias.t125 gnd 0.176757f
C4650 commonsourceibias.n11 gnd 0.007641f
C4651 commonsourceibias.n12 gnd 0.012624f
C4652 commonsourceibias.t12 gnd 0.191163f
C4653 commonsourceibias.t48 gnd 0.176757f
C4654 commonsourceibias.n13 gnd 0.00769f
C4655 commonsourceibias.n14 gnd 0.009461f
C4656 commonsourceibias.t4 gnd 0.176757f
C4657 commonsourceibias.n15 gnd 0.009597f
C4658 commonsourceibias.n16 gnd 0.009461f
C4659 commonsourceibias.t10 gnd 0.176757f
C4660 commonsourceibias.n17 gnd 0.070526f
C4661 commonsourceibias.t58 gnd 0.176757f
C4662 commonsourceibias.n18 gnd 0.007653f
C4663 commonsourceibias.n19 gnd 0.009461f
C4664 commonsourceibias.t16 gnd 0.176757f
C4665 commonsourceibias.n20 gnd 0.009134f
C4666 commonsourceibias.n21 gnd 0.009461f
C4667 commonsourceibias.t28 gnd 0.176757f
C4668 commonsourceibias.n22 gnd 0.070526f
C4669 commonsourceibias.t6 gnd 0.176757f
C4670 commonsourceibias.n23 gnd 0.007641f
C4671 commonsourceibias.n24 gnd 0.009461f
C4672 commonsourceibias.t14 gnd 0.176757f
C4673 commonsourceibias.t44 gnd 0.176757f
C4674 commonsourceibias.n25 gnd 0.070526f
C4675 commonsourceibias.n26 gnd 0.009461f
C4676 commonsourceibias.t24 gnd 0.176757f
C4677 commonsourceibias.n27 gnd 0.070526f
C4678 commonsourceibias.n28 gnd 0.009461f
C4679 commonsourceibias.t30 gnd 0.176757f
C4680 commonsourceibias.n29 gnd 0.070526f
C4681 commonsourceibias.n30 gnd 0.009461f
C4682 commonsourceibias.t54 gnd 0.176757f
C4683 commonsourceibias.n31 gnd 0.010754f
C4684 commonsourceibias.n32 gnd 0.009461f
C4685 commonsourceibias.t18 gnd 0.176757f
C4686 commonsourceibias.n33 gnd 0.012717f
C4687 commonsourceibias.t0 gnd 0.196904f
C4688 commonsourceibias.t50 gnd 0.176757f
C4689 commonsourceibias.n34 gnd 0.078584f
C4690 commonsourceibias.n35 gnd 0.084191f
C4691 commonsourceibias.n36 gnd 0.04027f
C4692 commonsourceibias.n37 gnd 0.009461f
C4693 commonsourceibias.n38 gnd 0.00769f
C4694 commonsourceibias.n39 gnd 0.013037f
C4695 commonsourceibias.n40 gnd 0.070526f
C4696 commonsourceibias.n41 gnd 0.013093f
C4697 commonsourceibias.n42 gnd 0.009461f
C4698 commonsourceibias.n43 gnd 0.009461f
C4699 commonsourceibias.n44 gnd 0.009461f
C4700 commonsourceibias.n45 gnd 0.009597f
C4701 commonsourceibias.n46 gnd 0.070526f
C4702 commonsourceibias.n47 gnd 0.011661f
C4703 commonsourceibias.n48 gnd 0.0129f
C4704 commonsourceibias.n49 gnd 0.009461f
C4705 commonsourceibias.n50 gnd 0.009461f
C4706 commonsourceibias.n51 gnd 0.012816f
C4707 commonsourceibias.n52 gnd 0.007653f
C4708 commonsourceibias.n53 gnd 0.012975f
C4709 commonsourceibias.n54 gnd 0.009461f
C4710 commonsourceibias.n55 gnd 0.009461f
C4711 commonsourceibias.n56 gnd 0.013054f
C4712 commonsourceibias.n57 gnd 0.011256f
C4713 commonsourceibias.n58 gnd 0.009134f
C4714 commonsourceibias.n59 gnd 0.009461f
C4715 commonsourceibias.n60 gnd 0.009461f
C4716 commonsourceibias.n61 gnd 0.011572f
C4717 commonsourceibias.n62 gnd 0.012989f
C4718 commonsourceibias.n63 gnd 0.070526f
C4719 commonsourceibias.n64 gnd 0.012901f
C4720 commonsourceibias.n65 gnd 0.009461f
C4721 commonsourceibias.n66 gnd 0.009461f
C4722 commonsourceibias.n67 gnd 0.009461f
C4723 commonsourceibias.n68 gnd 0.012901f
C4724 commonsourceibias.n69 gnd 0.070526f
C4725 commonsourceibias.n70 gnd 0.012989f
C4726 commonsourceibias.n71 gnd 0.011572f
C4727 commonsourceibias.n72 gnd 0.009461f
C4728 commonsourceibias.n73 gnd 0.009461f
C4729 commonsourceibias.n74 gnd 0.009461f
C4730 commonsourceibias.n75 gnd 0.011256f
C4731 commonsourceibias.n76 gnd 0.013054f
C4732 commonsourceibias.n77 gnd 0.070526f
C4733 commonsourceibias.n78 gnd 0.012975f
C4734 commonsourceibias.n79 gnd 0.009461f
C4735 commonsourceibias.n80 gnd 0.009461f
C4736 commonsourceibias.n81 gnd 0.009461f
C4737 commonsourceibias.n82 gnd 0.012816f
C4738 commonsourceibias.n83 gnd 0.070526f
C4739 commonsourceibias.n84 gnd 0.0129f
C4740 commonsourceibias.n85 gnd 0.011661f
C4741 commonsourceibias.n86 gnd 0.009461f
C4742 commonsourceibias.n87 gnd 0.009461f
C4743 commonsourceibias.n88 gnd 0.009461f
C4744 commonsourceibias.n89 gnd 0.010754f
C4745 commonsourceibias.n90 gnd 0.013093f
C4746 commonsourceibias.n91 gnd 0.070526f
C4747 commonsourceibias.n92 gnd 0.013037f
C4748 commonsourceibias.n93 gnd 0.009461f
C4749 commonsourceibias.n94 gnd 0.009461f
C4750 commonsourceibias.n95 gnd 0.009461f
C4751 commonsourceibias.n96 gnd 0.012717f
C4752 commonsourceibias.n97 gnd 0.070526f
C4753 commonsourceibias.n98 gnd 0.012748f
C4754 commonsourceibias.n99 gnd 0.085044f
C4755 commonsourceibias.n100 gnd 0.095092f
C4756 commonsourceibias.t13 gnd 0.020415f
C4757 commonsourceibias.t49 gnd 0.020415f
C4758 commonsourceibias.n101 gnd 0.180398f
C4759 commonsourceibias.n102 gnd 0.156264f
C4760 commonsourceibias.t5 gnd 0.020415f
C4761 commonsourceibias.t11 gnd 0.020415f
C4762 commonsourceibias.n103 gnd 0.180398f
C4763 commonsourceibias.n104 gnd 0.082864f
C4764 commonsourceibias.t59 gnd 0.020415f
C4765 commonsourceibias.t17 gnd 0.020415f
C4766 commonsourceibias.n105 gnd 0.180398f
C4767 commonsourceibias.n106 gnd 0.082864f
C4768 commonsourceibias.t29 gnd 0.020415f
C4769 commonsourceibias.t7 gnd 0.020415f
C4770 commonsourceibias.n107 gnd 0.180398f
C4771 commonsourceibias.n108 gnd 0.069229f
C4772 commonsourceibias.t51 gnd 0.020415f
C4773 commonsourceibias.t1 gnd 0.020415f
C4774 commonsourceibias.n109 gnd 0.181002f
C4775 commonsourceibias.t55 gnd 0.020415f
C4776 commonsourceibias.t19 gnd 0.020415f
C4777 commonsourceibias.n110 gnd 0.180398f
C4778 commonsourceibias.n111 gnd 0.168097f
C4779 commonsourceibias.t25 gnd 0.020415f
C4780 commonsourceibias.t31 gnd 0.020415f
C4781 commonsourceibias.n112 gnd 0.180398f
C4782 commonsourceibias.n113 gnd 0.082864f
C4783 commonsourceibias.t15 gnd 0.020415f
C4784 commonsourceibias.t45 gnd 0.020415f
C4785 commonsourceibias.n114 gnd 0.180398f
C4786 commonsourceibias.n115 gnd 0.069229f
C4787 commonsourceibias.n116 gnd 0.083829f
C4788 commonsourceibias.n117 gnd 0.009461f
C4789 commonsourceibias.t118 gnd 0.176757f
C4790 commonsourceibias.t76 gnd 0.176757f
C4791 commonsourceibias.n118 gnd 0.070526f
C4792 commonsourceibias.n119 gnd 0.009461f
C4793 commonsourceibias.t106 gnd 0.176757f
C4794 commonsourceibias.n120 gnd 0.070526f
C4795 commonsourceibias.n121 gnd 0.009461f
C4796 commonsourceibias.t96 gnd 0.176757f
C4797 commonsourceibias.n122 gnd 0.070526f
C4798 commonsourceibias.n123 gnd 0.009461f
C4799 commonsourceibias.t141 gnd 0.176757f
C4800 commonsourceibias.n124 gnd 0.010754f
C4801 commonsourceibias.n125 gnd 0.009461f
C4802 commonsourceibias.t116 gnd 0.176757f
C4803 commonsourceibias.n126 gnd 0.012717f
C4804 commonsourceibias.t129 gnd 0.196904f
C4805 commonsourceibias.t152 gnd 0.176757f
C4806 commonsourceibias.n127 gnd 0.078584f
C4807 commonsourceibias.n128 gnd 0.084191f
C4808 commonsourceibias.n129 gnd 0.04027f
C4809 commonsourceibias.n130 gnd 0.009461f
C4810 commonsourceibias.n131 gnd 0.00769f
C4811 commonsourceibias.n132 gnd 0.013037f
C4812 commonsourceibias.n133 gnd 0.070526f
C4813 commonsourceibias.n134 gnd 0.013093f
C4814 commonsourceibias.n135 gnd 0.009461f
C4815 commonsourceibias.n136 gnd 0.009461f
C4816 commonsourceibias.n137 gnd 0.009461f
C4817 commonsourceibias.n138 gnd 0.009597f
C4818 commonsourceibias.n139 gnd 0.070526f
C4819 commonsourceibias.n140 gnd 0.011661f
C4820 commonsourceibias.n141 gnd 0.0129f
C4821 commonsourceibias.n142 gnd 0.009461f
C4822 commonsourceibias.n143 gnd 0.009461f
C4823 commonsourceibias.n144 gnd 0.012816f
C4824 commonsourceibias.n145 gnd 0.007653f
C4825 commonsourceibias.n146 gnd 0.012975f
C4826 commonsourceibias.n147 gnd 0.009461f
C4827 commonsourceibias.n148 gnd 0.009461f
C4828 commonsourceibias.n149 gnd 0.013054f
C4829 commonsourceibias.n150 gnd 0.011256f
C4830 commonsourceibias.n151 gnd 0.009134f
C4831 commonsourceibias.n152 gnd 0.009461f
C4832 commonsourceibias.n153 gnd 0.009461f
C4833 commonsourceibias.n154 gnd 0.011572f
C4834 commonsourceibias.n155 gnd 0.012989f
C4835 commonsourceibias.n156 gnd 0.070526f
C4836 commonsourceibias.n157 gnd 0.012901f
C4837 commonsourceibias.n158 gnd 0.009415f
C4838 commonsourceibias.n159 gnd 0.06839f
C4839 commonsourceibias.n160 gnd 0.009415f
C4840 commonsourceibias.n161 gnd 0.012901f
C4841 commonsourceibias.n162 gnd 0.070526f
C4842 commonsourceibias.n163 gnd 0.012989f
C4843 commonsourceibias.n164 gnd 0.011572f
C4844 commonsourceibias.n165 gnd 0.009461f
C4845 commonsourceibias.n166 gnd 0.009461f
C4846 commonsourceibias.n167 gnd 0.009461f
C4847 commonsourceibias.n168 gnd 0.011256f
C4848 commonsourceibias.n169 gnd 0.013054f
C4849 commonsourceibias.n170 gnd 0.070526f
C4850 commonsourceibias.n171 gnd 0.012975f
C4851 commonsourceibias.n172 gnd 0.009461f
C4852 commonsourceibias.n173 gnd 0.009461f
C4853 commonsourceibias.n174 gnd 0.009461f
C4854 commonsourceibias.n175 gnd 0.012816f
C4855 commonsourceibias.n176 gnd 0.070526f
C4856 commonsourceibias.n177 gnd 0.0129f
C4857 commonsourceibias.n178 gnd 0.011661f
C4858 commonsourceibias.n179 gnd 0.009461f
C4859 commonsourceibias.n180 gnd 0.009461f
C4860 commonsourceibias.n181 gnd 0.009461f
C4861 commonsourceibias.n182 gnd 0.010754f
C4862 commonsourceibias.n183 gnd 0.013093f
C4863 commonsourceibias.n184 gnd 0.070526f
C4864 commonsourceibias.n185 gnd 0.013037f
C4865 commonsourceibias.n186 gnd 0.009461f
C4866 commonsourceibias.n187 gnd 0.009461f
C4867 commonsourceibias.n188 gnd 0.009461f
C4868 commonsourceibias.n189 gnd 0.012717f
C4869 commonsourceibias.n190 gnd 0.070526f
C4870 commonsourceibias.n191 gnd 0.012748f
C4871 commonsourceibias.n192 gnd 0.085044f
C4872 commonsourceibias.n193 gnd 0.056182f
C4873 commonsourceibias.n194 gnd 0.012624f
C4874 commonsourceibias.t71 gnd 0.191163f
C4875 commonsourceibias.t159 gnd 0.176757f
C4876 commonsourceibias.n195 gnd 0.00769f
C4877 commonsourceibias.n196 gnd 0.009461f
C4878 commonsourceibias.t148 gnd 0.176757f
C4879 commonsourceibias.n197 gnd 0.009597f
C4880 commonsourceibias.n198 gnd 0.009461f
C4881 commonsourceibias.t78 gnd 0.176757f
C4882 commonsourceibias.n199 gnd 0.070526f
C4883 commonsourceibias.t157 gnd 0.176757f
C4884 commonsourceibias.n200 gnd 0.007653f
C4885 commonsourceibias.n201 gnd 0.009461f
C4886 commonsourceibias.t85 gnd 0.176757f
C4887 commonsourceibias.n202 gnd 0.009134f
C4888 commonsourceibias.n203 gnd 0.009461f
C4889 commonsourceibias.t77 gnd 0.176757f
C4890 commonsourceibias.n204 gnd 0.070526f
C4891 commonsourceibias.t158 gnd 0.176757f
C4892 commonsourceibias.n205 gnd 0.007641f
C4893 commonsourceibias.n206 gnd 0.009461f
C4894 commonsourceibias.t94 gnd 0.176757f
C4895 commonsourceibias.t113 gnd 0.176757f
C4896 commonsourceibias.n207 gnd 0.070526f
C4897 commonsourceibias.n208 gnd 0.009461f
C4898 commonsourceibias.t156 gnd 0.176757f
C4899 commonsourceibias.n209 gnd 0.070526f
C4900 commonsourceibias.n210 gnd 0.009461f
C4901 commonsourceibias.t92 gnd 0.176757f
C4902 commonsourceibias.n211 gnd 0.070526f
C4903 commonsourceibias.n212 gnd 0.009461f
C4904 commonsourceibias.t111 gnd 0.176757f
C4905 commonsourceibias.n213 gnd 0.010754f
C4906 commonsourceibias.n214 gnd 0.009461f
C4907 commonsourceibias.t105 gnd 0.176757f
C4908 commonsourceibias.n215 gnd 0.012717f
C4909 commonsourceibias.t112 gnd 0.196904f
C4910 commonsourceibias.t93 gnd 0.176757f
C4911 commonsourceibias.n216 gnd 0.078584f
C4912 commonsourceibias.n217 gnd 0.084191f
C4913 commonsourceibias.n218 gnd 0.04027f
C4914 commonsourceibias.n219 gnd 0.009461f
C4915 commonsourceibias.n220 gnd 0.00769f
C4916 commonsourceibias.n221 gnd 0.013037f
C4917 commonsourceibias.n222 gnd 0.070526f
C4918 commonsourceibias.n223 gnd 0.013093f
C4919 commonsourceibias.n224 gnd 0.009461f
C4920 commonsourceibias.n225 gnd 0.009461f
C4921 commonsourceibias.n226 gnd 0.009461f
C4922 commonsourceibias.n227 gnd 0.009597f
C4923 commonsourceibias.n228 gnd 0.070526f
C4924 commonsourceibias.n229 gnd 0.011661f
C4925 commonsourceibias.n230 gnd 0.0129f
C4926 commonsourceibias.n231 gnd 0.009461f
C4927 commonsourceibias.n232 gnd 0.009461f
C4928 commonsourceibias.n233 gnd 0.012816f
C4929 commonsourceibias.n234 gnd 0.007653f
C4930 commonsourceibias.n235 gnd 0.012975f
C4931 commonsourceibias.n236 gnd 0.009461f
C4932 commonsourceibias.n237 gnd 0.009461f
C4933 commonsourceibias.n238 gnd 0.013054f
C4934 commonsourceibias.n239 gnd 0.011256f
C4935 commonsourceibias.n240 gnd 0.009134f
C4936 commonsourceibias.n241 gnd 0.009461f
C4937 commonsourceibias.n242 gnd 0.009461f
C4938 commonsourceibias.n243 gnd 0.011572f
C4939 commonsourceibias.n244 gnd 0.012989f
C4940 commonsourceibias.n245 gnd 0.070526f
C4941 commonsourceibias.n246 gnd 0.012901f
C4942 commonsourceibias.n247 gnd 0.009461f
C4943 commonsourceibias.n248 gnd 0.009461f
C4944 commonsourceibias.n249 gnd 0.009461f
C4945 commonsourceibias.n250 gnd 0.012901f
C4946 commonsourceibias.n251 gnd 0.070526f
C4947 commonsourceibias.n252 gnd 0.012989f
C4948 commonsourceibias.n253 gnd 0.011572f
C4949 commonsourceibias.n254 gnd 0.009461f
C4950 commonsourceibias.n255 gnd 0.009461f
C4951 commonsourceibias.n256 gnd 0.009461f
C4952 commonsourceibias.n257 gnd 0.011256f
C4953 commonsourceibias.n258 gnd 0.013054f
C4954 commonsourceibias.n259 gnd 0.070526f
C4955 commonsourceibias.n260 gnd 0.012975f
C4956 commonsourceibias.n261 gnd 0.009461f
C4957 commonsourceibias.n262 gnd 0.009461f
C4958 commonsourceibias.n263 gnd 0.009461f
C4959 commonsourceibias.n264 gnd 0.012816f
C4960 commonsourceibias.n265 gnd 0.070526f
C4961 commonsourceibias.n266 gnd 0.0129f
C4962 commonsourceibias.n267 gnd 0.011661f
C4963 commonsourceibias.n268 gnd 0.009461f
C4964 commonsourceibias.n269 gnd 0.009461f
C4965 commonsourceibias.n270 gnd 0.009461f
C4966 commonsourceibias.n271 gnd 0.010754f
C4967 commonsourceibias.n272 gnd 0.013093f
C4968 commonsourceibias.n273 gnd 0.070526f
C4969 commonsourceibias.n274 gnd 0.013037f
C4970 commonsourceibias.n275 gnd 0.009461f
C4971 commonsourceibias.n276 gnd 0.009461f
C4972 commonsourceibias.n277 gnd 0.009461f
C4973 commonsourceibias.n278 gnd 0.012717f
C4974 commonsourceibias.n279 gnd 0.070526f
C4975 commonsourceibias.n280 gnd 0.012748f
C4976 commonsourceibias.n281 gnd 0.085044f
C4977 commonsourceibias.n282 gnd 0.030348f
C4978 commonsourceibias.n283 gnd 0.15151f
C4979 commonsourceibias.n284 gnd 0.012624f
C4980 commonsourceibias.t75 gnd 0.176757f
C4981 commonsourceibias.n285 gnd 0.00769f
C4982 commonsourceibias.n286 gnd 0.009461f
C4983 commonsourceibias.t128 gnd 0.176757f
C4984 commonsourceibias.n287 gnd 0.009597f
C4985 commonsourceibias.n288 gnd 0.009461f
C4986 commonsourceibias.t124 gnd 0.176757f
C4987 commonsourceibias.n289 gnd 0.070526f
C4988 commonsourceibias.t155 gnd 0.176757f
C4989 commonsourceibias.n290 gnd 0.007653f
C4990 commonsourceibias.n291 gnd 0.009461f
C4991 commonsourceibias.t90 gnd 0.176757f
C4992 commonsourceibias.n292 gnd 0.009134f
C4993 commonsourceibias.n293 gnd 0.009461f
C4994 commonsourceibias.t119 gnd 0.176757f
C4995 commonsourceibias.n294 gnd 0.070526f
C4996 commonsourceibias.t146 gnd 0.176757f
C4997 commonsourceibias.n295 gnd 0.007641f
C4998 commonsourceibias.n296 gnd 0.009461f
C4999 commonsourceibias.t138 gnd 0.176757f
C5000 commonsourceibias.t64 gnd 0.176757f
C5001 commonsourceibias.n297 gnd 0.070526f
C5002 commonsourceibias.n298 gnd 0.009461f
C5003 commonsourceibias.t137 gnd 0.176757f
C5004 commonsourceibias.n299 gnd 0.070526f
C5005 commonsourceibias.n300 gnd 0.009461f
C5006 commonsourceibias.t133 gnd 0.176757f
C5007 commonsourceibias.n301 gnd 0.070526f
C5008 commonsourceibias.n302 gnd 0.009461f
C5009 commonsourceibias.t149 gnd 0.176757f
C5010 commonsourceibias.n303 gnd 0.010754f
C5011 commonsourceibias.n304 gnd 0.009461f
C5012 commonsourceibias.t79 gnd 0.176757f
C5013 commonsourceibias.n305 gnd 0.012717f
C5014 commonsourceibias.t140 gnd 0.196904f
C5015 commonsourceibias.t130 gnd 0.176757f
C5016 commonsourceibias.n306 gnd 0.078584f
C5017 commonsourceibias.n307 gnd 0.084191f
C5018 commonsourceibias.n308 gnd 0.04027f
C5019 commonsourceibias.n309 gnd 0.009461f
C5020 commonsourceibias.n310 gnd 0.00769f
C5021 commonsourceibias.n311 gnd 0.013037f
C5022 commonsourceibias.n312 gnd 0.070526f
C5023 commonsourceibias.n313 gnd 0.013093f
C5024 commonsourceibias.n314 gnd 0.009461f
C5025 commonsourceibias.n315 gnd 0.009461f
C5026 commonsourceibias.n316 gnd 0.009461f
C5027 commonsourceibias.n317 gnd 0.009597f
C5028 commonsourceibias.n318 gnd 0.070526f
C5029 commonsourceibias.n319 gnd 0.011661f
C5030 commonsourceibias.n320 gnd 0.0129f
C5031 commonsourceibias.n321 gnd 0.009461f
C5032 commonsourceibias.n322 gnd 0.009461f
C5033 commonsourceibias.n323 gnd 0.012816f
C5034 commonsourceibias.n324 gnd 0.007653f
C5035 commonsourceibias.n325 gnd 0.012975f
C5036 commonsourceibias.n326 gnd 0.009461f
C5037 commonsourceibias.n327 gnd 0.009461f
C5038 commonsourceibias.n328 gnd 0.013054f
C5039 commonsourceibias.n329 gnd 0.011256f
C5040 commonsourceibias.n330 gnd 0.009134f
C5041 commonsourceibias.n331 gnd 0.009461f
C5042 commonsourceibias.n332 gnd 0.009461f
C5043 commonsourceibias.n333 gnd 0.011572f
C5044 commonsourceibias.n334 gnd 0.012989f
C5045 commonsourceibias.n335 gnd 0.070526f
C5046 commonsourceibias.n336 gnd 0.012901f
C5047 commonsourceibias.n337 gnd 0.009461f
C5048 commonsourceibias.n338 gnd 0.009461f
C5049 commonsourceibias.n339 gnd 0.009461f
C5050 commonsourceibias.n340 gnd 0.012901f
C5051 commonsourceibias.n341 gnd 0.070526f
C5052 commonsourceibias.n342 gnd 0.012989f
C5053 commonsourceibias.n343 gnd 0.011572f
C5054 commonsourceibias.n344 gnd 0.009461f
C5055 commonsourceibias.n345 gnd 0.009461f
C5056 commonsourceibias.n346 gnd 0.009461f
C5057 commonsourceibias.n347 gnd 0.011256f
C5058 commonsourceibias.n348 gnd 0.013054f
C5059 commonsourceibias.n349 gnd 0.070526f
C5060 commonsourceibias.n350 gnd 0.012975f
C5061 commonsourceibias.n351 gnd 0.009461f
C5062 commonsourceibias.n352 gnd 0.009461f
C5063 commonsourceibias.n353 gnd 0.009461f
C5064 commonsourceibias.n354 gnd 0.012816f
C5065 commonsourceibias.n355 gnd 0.070526f
C5066 commonsourceibias.n356 gnd 0.0129f
C5067 commonsourceibias.n357 gnd 0.011661f
C5068 commonsourceibias.n358 gnd 0.009461f
C5069 commonsourceibias.n359 gnd 0.009461f
C5070 commonsourceibias.n360 gnd 0.009461f
C5071 commonsourceibias.n361 gnd 0.010754f
C5072 commonsourceibias.n362 gnd 0.013093f
C5073 commonsourceibias.n363 gnd 0.070526f
C5074 commonsourceibias.n364 gnd 0.013037f
C5075 commonsourceibias.n365 gnd 0.009461f
C5076 commonsourceibias.n366 gnd 0.009461f
C5077 commonsourceibias.n367 gnd 0.009461f
C5078 commonsourceibias.n368 gnd 0.012717f
C5079 commonsourceibias.n369 gnd 0.070526f
C5080 commonsourceibias.n370 gnd 0.012748f
C5081 commonsourceibias.t147 gnd 0.191163f
C5082 commonsourceibias.n371 gnd 0.085044f
C5083 commonsourceibias.n372 gnd 0.030348f
C5084 commonsourceibias.n373 gnd 0.449685f
C5085 commonsourceibias.n374 gnd 0.012624f
C5086 commonsourceibias.t91 gnd 0.191163f
C5087 commonsourceibias.t134 gnd 0.176757f
C5088 commonsourceibias.n375 gnd 0.00769f
C5089 commonsourceibias.n376 gnd 0.009461f
C5090 commonsourceibias.t114 gnd 0.176757f
C5091 commonsourceibias.n377 gnd 0.009597f
C5092 commonsourceibias.n378 gnd 0.009461f
C5093 commonsourceibias.t123 gnd 0.176757f
C5094 commonsourceibias.n379 gnd 0.007653f
C5095 commonsourceibias.n380 gnd 0.009461f
C5096 commonsourceibias.t88 gnd 0.176757f
C5097 commonsourceibias.n381 gnd 0.009134f
C5098 commonsourceibias.n382 gnd 0.009461f
C5099 commonsourceibias.t104 gnd 0.176757f
C5100 commonsourceibias.n383 gnd 0.007641f
C5101 commonsourceibias.n384 gnd 0.009461f
C5102 commonsourceibias.t89 gnd 0.176757f
C5103 commonsourceibias.t139 gnd 0.176757f
C5104 commonsourceibias.n385 gnd 0.070526f
C5105 commonsourceibias.n386 gnd 0.009461f
C5106 commonsourceibias.t83 gnd 0.176757f
C5107 commonsourceibias.n387 gnd 0.070526f
C5108 commonsourceibias.n388 gnd 0.009461f
C5109 commonsourceibias.t150 gnd 0.176757f
C5110 commonsourceibias.n389 gnd 0.070526f
C5111 commonsourceibias.n390 gnd 0.009461f
C5112 commonsourceibias.t127 gnd 0.176757f
C5113 commonsourceibias.n391 gnd 0.010754f
C5114 commonsourceibias.n392 gnd 0.009461f
C5115 commonsourceibias.t84 gnd 0.176757f
C5116 commonsourceibias.n393 gnd 0.012717f
C5117 commonsourceibias.t108 gnd 0.196904f
C5118 commonsourceibias.t131 gnd 0.176757f
C5119 commonsourceibias.n394 gnd 0.078584f
C5120 commonsourceibias.n395 gnd 0.084191f
C5121 commonsourceibias.n396 gnd 0.04027f
C5122 commonsourceibias.n397 gnd 0.009461f
C5123 commonsourceibias.n398 gnd 0.00769f
C5124 commonsourceibias.n399 gnd 0.013037f
C5125 commonsourceibias.n400 gnd 0.070526f
C5126 commonsourceibias.n401 gnd 0.013093f
C5127 commonsourceibias.n402 gnd 0.009461f
C5128 commonsourceibias.n403 gnd 0.009461f
C5129 commonsourceibias.n404 gnd 0.009461f
C5130 commonsourceibias.n405 gnd 0.009597f
C5131 commonsourceibias.n406 gnd 0.070526f
C5132 commonsourceibias.n407 gnd 0.011661f
C5133 commonsourceibias.n408 gnd 0.0129f
C5134 commonsourceibias.n409 gnd 0.009461f
C5135 commonsourceibias.n410 gnd 0.009461f
C5136 commonsourceibias.n411 gnd 0.012816f
C5137 commonsourceibias.n412 gnd 0.007653f
C5138 commonsourceibias.n413 gnd 0.012975f
C5139 commonsourceibias.n414 gnd 0.009461f
C5140 commonsourceibias.n415 gnd 0.009461f
C5141 commonsourceibias.n416 gnd 0.013054f
C5142 commonsourceibias.n417 gnd 0.011256f
C5143 commonsourceibias.n418 gnd 0.009134f
C5144 commonsourceibias.n419 gnd 0.009461f
C5145 commonsourceibias.n420 gnd 0.009461f
C5146 commonsourceibias.n421 gnd 0.011572f
C5147 commonsourceibias.n422 gnd 0.012989f
C5148 commonsourceibias.n423 gnd 0.070526f
C5149 commonsourceibias.n424 gnd 0.012901f
C5150 commonsourceibias.n425 gnd 0.009415f
C5151 commonsourceibias.t23 gnd 0.020415f
C5152 commonsourceibias.t63 gnd 0.020415f
C5153 commonsourceibias.n426 gnd 0.181002f
C5154 commonsourceibias.t41 gnd 0.020415f
C5155 commonsourceibias.t3 gnd 0.020415f
C5156 commonsourceibias.n427 gnd 0.180398f
C5157 commonsourceibias.n428 gnd 0.168097f
C5158 commonsourceibias.t53 gnd 0.020415f
C5159 commonsourceibias.t43 gnd 0.020415f
C5160 commonsourceibias.n429 gnd 0.180398f
C5161 commonsourceibias.n430 gnd 0.082864f
C5162 commonsourceibias.t57 gnd 0.020415f
C5163 commonsourceibias.t37 gnd 0.020415f
C5164 commonsourceibias.n431 gnd 0.180398f
C5165 commonsourceibias.n432 gnd 0.069229f
C5166 commonsourceibias.n433 gnd 0.012624f
C5167 commonsourceibias.t60 gnd 0.176757f
C5168 commonsourceibias.n434 gnd 0.00769f
C5169 commonsourceibias.n435 gnd 0.009461f
C5170 commonsourceibias.t20 gnd 0.176757f
C5171 commonsourceibias.n436 gnd 0.009597f
C5172 commonsourceibias.n437 gnd 0.009461f
C5173 commonsourceibias.t8 gnd 0.176757f
C5174 commonsourceibias.n438 gnd 0.007653f
C5175 commonsourceibias.n439 gnd 0.009461f
C5176 commonsourceibias.t38 gnd 0.176757f
C5177 commonsourceibias.n440 gnd 0.009134f
C5178 commonsourceibias.n441 gnd 0.009461f
C5179 commonsourceibias.t26 gnd 0.176757f
C5180 commonsourceibias.n442 gnd 0.007641f
C5181 commonsourceibias.n443 gnd 0.009461f
C5182 commonsourceibias.t36 gnd 0.176757f
C5183 commonsourceibias.t56 gnd 0.176757f
C5184 commonsourceibias.n444 gnd 0.070526f
C5185 commonsourceibias.n445 gnd 0.009461f
C5186 commonsourceibias.t42 gnd 0.176757f
C5187 commonsourceibias.n446 gnd 0.070526f
C5188 commonsourceibias.n447 gnd 0.009461f
C5189 commonsourceibias.t52 gnd 0.176757f
C5190 commonsourceibias.n448 gnd 0.070526f
C5191 commonsourceibias.n449 gnd 0.009461f
C5192 commonsourceibias.t2 gnd 0.176757f
C5193 commonsourceibias.n450 gnd 0.010754f
C5194 commonsourceibias.n451 gnd 0.009461f
C5195 commonsourceibias.t40 gnd 0.176757f
C5196 commonsourceibias.n452 gnd 0.012717f
C5197 commonsourceibias.t22 gnd 0.196904f
C5198 commonsourceibias.t62 gnd 0.176757f
C5199 commonsourceibias.n453 gnd 0.078584f
C5200 commonsourceibias.n454 gnd 0.084191f
C5201 commonsourceibias.n455 gnd 0.04027f
C5202 commonsourceibias.n456 gnd 0.009461f
C5203 commonsourceibias.n457 gnd 0.00769f
C5204 commonsourceibias.n458 gnd 0.013037f
C5205 commonsourceibias.n459 gnd 0.070526f
C5206 commonsourceibias.n460 gnd 0.013093f
C5207 commonsourceibias.n461 gnd 0.009461f
C5208 commonsourceibias.n462 gnd 0.009461f
C5209 commonsourceibias.n463 gnd 0.009461f
C5210 commonsourceibias.n464 gnd 0.009597f
C5211 commonsourceibias.n465 gnd 0.070526f
C5212 commonsourceibias.n466 gnd 0.011661f
C5213 commonsourceibias.n467 gnd 0.0129f
C5214 commonsourceibias.n468 gnd 0.009461f
C5215 commonsourceibias.n469 gnd 0.009461f
C5216 commonsourceibias.n470 gnd 0.012816f
C5217 commonsourceibias.n471 gnd 0.007653f
C5218 commonsourceibias.n472 gnd 0.012975f
C5219 commonsourceibias.n473 gnd 0.009461f
C5220 commonsourceibias.n474 gnd 0.009461f
C5221 commonsourceibias.n475 gnd 0.013054f
C5222 commonsourceibias.n476 gnd 0.011256f
C5223 commonsourceibias.n477 gnd 0.009134f
C5224 commonsourceibias.n478 gnd 0.009461f
C5225 commonsourceibias.n479 gnd 0.009461f
C5226 commonsourceibias.n480 gnd 0.011572f
C5227 commonsourceibias.n481 gnd 0.012989f
C5228 commonsourceibias.n482 gnd 0.070526f
C5229 commonsourceibias.n483 gnd 0.012901f
C5230 commonsourceibias.n484 gnd 0.009461f
C5231 commonsourceibias.n485 gnd 0.009461f
C5232 commonsourceibias.n486 gnd 0.009461f
C5233 commonsourceibias.n487 gnd 0.012901f
C5234 commonsourceibias.n488 gnd 0.070526f
C5235 commonsourceibias.n489 gnd 0.012989f
C5236 commonsourceibias.t46 gnd 0.176757f
C5237 commonsourceibias.n490 gnd 0.070526f
C5238 commonsourceibias.n491 gnd 0.011572f
C5239 commonsourceibias.n492 gnd 0.009461f
C5240 commonsourceibias.n493 gnd 0.009461f
C5241 commonsourceibias.n494 gnd 0.009461f
C5242 commonsourceibias.n495 gnd 0.011256f
C5243 commonsourceibias.n496 gnd 0.013054f
C5244 commonsourceibias.n497 gnd 0.070526f
C5245 commonsourceibias.n498 gnd 0.012975f
C5246 commonsourceibias.n499 gnd 0.009461f
C5247 commonsourceibias.n500 gnd 0.009461f
C5248 commonsourceibias.n501 gnd 0.009461f
C5249 commonsourceibias.n502 gnd 0.012816f
C5250 commonsourceibias.n503 gnd 0.070526f
C5251 commonsourceibias.n504 gnd 0.0129f
C5252 commonsourceibias.t32 gnd 0.176757f
C5253 commonsourceibias.n505 gnd 0.070526f
C5254 commonsourceibias.n506 gnd 0.011661f
C5255 commonsourceibias.n507 gnd 0.009461f
C5256 commonsourceibias.n508 gnd 0.009461f
C5257 commonsourceibias.n509 gnd 0.009461f
C5258 commonsourceibias.n510 gnd 0.010754f
C5259 commonsourceibias.n511 gnd 0.013093f
C5260 commonsourceibias.n512 gnd 0.070526f
C5261 commonsourceibias.n513 gnd 0.013037f
C5262 commonsourceibias.n514 gnd 0.009461f
C5263 commonsourceibias.n515 gnd 0.009461f
C5264 commonsourceibias.n516 gnd 0.009461f
C5265 commonsourceibias.n517 gnd 0.012717f
C5266 commonsourceibias.n518 gnd 0.070526f
C5267 commonsourceibias.n519 gnd 0.012748f
C5268 commonsourceibias.t34 gnd 0.191163f
C5269 commonsourceibias.n520 gnd 0.085044f
C5270 commonsourceibias.n521 gnd 0.095092f
C5271 commonsourceibias.t61 gnd 0.020415f
C5272 commonsourceibias.t35 gnd 0.020415f
C5273 commonsourceibias.n522 gnd 0.180398f
C5274 commonsourceibias.n523 gnd 0.156264f
C5275 commonsourceibias.t33 gnd 0.020415f
C5276 commonsourceibias.t21 gnd 0.020415f
C5277 commonsourceibias.n524 gnd 0.180398f
C5278 commonsourceibias.n525 gnd 0.082864f
C5279 commonsourceibias.t39 gnd 0.020415f
C5280 commonsourceibias.t9 gnd 0.020415f
C5281 commonsourceibias.n526 gnd 0.180398f
C5282 commonsourceibias.n527 gnd 0.082864f
C5283 commonsourceibias.t27 gnd 0.020415f
C5284 commonsourceibias.t47 gnd 0.020415f
C5285 commonsourceibias.n528 gnd 0.180398f
C5286 commonsourceibias.n529 gnd 0.069229f
C5287 commonsourceibias.n530 gnd 0.083829f
C5288 commonsourceibias.n531 gnd 0.06839f
C5289 commonsourceibias.n532 gnd 0.009415f
C5290 commonsourceibias.n533 gnd 0.012901f
C5291 commonsourceibias.n534 gnd 0.070526f
C5292 commonsourceibias.n535 gnd 0.012989f
C5293 commonsourceibias.t73 gnd 0.176757f
C5294 commonsourceibias.n536 gnd 0.070526f
C5295 commonsourceibias.n537 gnd 0.011572f
C5296 commonsourceibias.n538 gnd 0.009461f
C5297 commonsourceibias.n539 gnd 0.009461f
C5298 commonsourceibias.n540 gnd 0.009461f
C5299 commonsourceibias.n541 gnd 0.011256f
C5300 commonsourceibias.n542 gnd 0.013054f
C5301 commonsourceibias.n543 gnd 0.070526f
C5302 commonsourceibias.n544 gnd 0.012975f
C5303 commonsourceibias.n545 gnd 0.009461f
C5304 commonsourceibias.n546 gnd 0.009461f
C5305 commonsourceibias.n547 gnd 0.009461f
C5306 commonsourceibias.n548 gnd 0.012816f
C5307 commonsourceibias.n549 gnd 0.070526f
C5308 commonsourceibias.n550 gnd 0.0129f
C5309 commonsourceibias.t95 gnd 0.176757f
C5310 commonsourceibias.n551 gnd 0.070526f
C5311 commonsourceibias.n552 gnd 0.011661f
C5312 commonsourceibias.n553 gnd 0.009461f
C5313 commonsourceibias.n554 gnd 0.009461f
C5314 commonsourceibias.n555 gnd 0.009461f
C5315 commonsourceibias.n556 gnd 0.010754f
C5316 commonsourceibias.n557 gnd 0.013093f
C5317 commonsourceibias.n558 gnd 0.070526f
C5318 commonsourceibias.n559 gnd 0.013037f
C5319 commonsourceibias.n560 gnd 0.009461f
C5320 commonsourceibias.n561 gnd 0.009461f
C5321 commonsourceibias.n562 gnd 0.009461f
C5322 commonsourceibias.n563 gnd 0.012717f
C5323 commonsourceibias.n564 gnd 0.070526f
C5324 commonsourceibias.n565 gnd 0.012748f
C5325 commonsourceibias.n566 gnd 0.085044f
C5326 commonsourceibias.n567 gnd 0.056182f
C5327 commonsourceibias.n568 gnd 0.012624f
C5328 commonsourceibias.t144 gnd 0.176757f
C5329 commonsourceibias.n569 gnd 0.00769f
C5330 commonsourceibias.n570 gnd 0.009461f
C5331 commonsourceibias.t66 gnd 0.176757f
C5332 commonsourceibias.n571 gnd 0.009597f
C5333 commonsourceibias.n572 gnd 0.009461f
C5334 commonsourceibias.t143 gnd 0.176757f
C5335 commonsourceibias.n573 gnd 0.007653f
C5336 commonsourceibias.n574 gnd 0.009461f
C5337 commonsourceibias.t65 gnd 0.176757f
C5338 commonsourceibias.n575 gnd 0.009134f
C5339 commonsourceibias.n576 gnd 0.009461f
C5340 commonsourceibias.t142 gnd 0.176757f
C5341 commonsourceibias.n577 gnd 0.007641f
C5342 commonsourceibias.n578 gnd 0.009461f
C5343 commonsourceibias.t72 gnd 0.176757f
C5344 commonsourceibias.t99 gnd 0.176757f
C5345 commonsourceibias.n579 gnd 0.070526f
C5346 commonsourceibias.n580 gnd 0.009461f
C5347 commonsourceibias.t80 gnd 0.176757f
C5348 commonsourceibias.n581 gnd 0.070526f
C5349 commonsourceibias.n582 gnd 0.009461f
C5350 commonsourceibias.t69 gnd 0.176757f
C5351 commonsourceibias.n583 gnd 0.070526f
C5352 commonsourceibias.n584 gnd 0.009461f
C5353 commonsourceibias.t98 gnd 0.176757f
C5354 commonsourceibias.n585 gnd 0.010754f
C5355 commonsourceibias.n586 gnd 0.009461f
C5356 commonsourceibias.t86 gnd 0.176757f
C5357 commonsourceibias.n587 gnd 0.012717f
C5358 commonsourceibias.t97 gnd 0.196904f
C5359 commonsourceibias.t68 gnd 0.176757f
C5360 commonsourceibias.n588 gnd 0.078584f
C5361 commonsourceibias.n589 gnd 0.084191f
C5362 commonsourceibias.n590 gnd 0.04027f
C5363 commonsourceibias.n591 gnd 0.009461f
C5364 commonsourceibias.n592 gnd 0.00769f
C5365 commonsourceibias.n593 gnd 0.013037f
C5366 commonsourceibias.n594 gnd 0.070526f
C5367 commonsourceibias.n595 gnd 0.013093f
C5368 commonsourceibias.n596 gnd 0.009461f
C5369 commonsourceibias.n597 gnd 0.009461f
C5370 commonsourceibias.n598 gnd 0.009461f
C5371 commonsourceibias.n599 gnd 0.009597f
C5372 commonsourceibias.n600 gnd 0.070526f
C5373 commonsourceibias.n601 gnd 0.011661f
C5374 commonsourceibias.n602 gnd 0.0129f
C5375 commonsourceibias.n603 gnd 0.009461f
C5376 commonsourceibias.n604 gnd 0.009461f
C5377 commonsourceibias.n605 gnd 0.012816f
C5378 commonsourceibias.n606 gnd 0.007653f
C5379 commonsourceibias.n607 gnd 0.012975f
C5380 commonsourceibias.n608 gnd 0.009461f
C5381 commonsourceibias.n609 gnd 0.009461f
C5382 commonsourceibias.n610 gnd 0.013054f
C5383 commonsourceibias.n611 gnd 0.011256f
C5384 commonsourceibias.n612 gnd 0.009134f
C5385 commonsourceibias.n613 gnd 0.009461f
C5386 commonsourceibias.n614 gnd 0.009461f
C5387 commonsourceibias.n615 gnd 0.011572f
C5388 commonsourceibias.n616 gnd 0.012989f
C5389 commonsourceibias.n617 gnd 0.070526f
C5390 commonsourceibias.n618 gnd 0.012901f
C5391 commonsourceibias.n619 gnd 0.009461f
C5392 commonsourceibias.n620 gnd 0.009461f
C5393 commonsourceibias.n621 gnd 0.009461f
C5394 commonsourceibias.n622 gnd 0.012901f
C5395 commonsourceibias.n623 gnd 0.070526f
C5396 commonsourceibias.n624 gnd 0.012989f
C5397 commonsourceibias.t100 gnd 0.176757f
C5398 commonsourceibias.n625 gnd 0.070526f
C5399 commonsourceibias.n626 gnd 0.011572f
C5400 commonsourceibias.n627 gnd 0.009461f
C5401 commonsourceibias.n628 gnd 0.009461f
C5402 commonsourceibias.n629 gnd 0.009461f
C5403 commonsourceibias.n630 gnd 0.011256f
C5404 commonsourceibias.n631 gnd 0.013054f
C5405 commonsourceibias.n632 gnd 0.070526f
C5406 commonsourceibias.n633 gnd 0.012975f
C5407 commonsourceibias.n634 gnd 0.009461f
C5408 commonsourceibias.n635 gnd 0.009461f
C5409 commonsourceibias.n636 gnd 0.009461f
C5410 commonsourceibias.n637 gnd 0.012816f
C5411 commonsourceibias.n638 gnd 0.070526f
C5412 commonsourceibias.n639 gnd 0.0129f
C5413 commonsourceibias.t154 gnd 0.176757f
C5414 commonsourceibias.n640 gnd 0.070526f
C5415 commonsourceibias.n641 gnd 0.011661f
C5416 commonsourceibias.n642 gnd 0.009461f
C5417 commonsourceibias.n643 gnd 0.009461f
C5418 commonsourceibias.n644 gnd 0.009461f
C5419 commonsourceibias.n645 gnd 0.010754f
C5420 commonsourceibias.n646 gnd 0.013093f
C5421 commonsourceibias.n647 gnd 0.070526f
C5422 commonsourceibias.n648 gnd 0.013037f
C5423 commonsourceibias.n649 gnd 0.009461f
C5424 commonsourceibias.n650 gnd 0.009461f
C5425 commonsourceibias.n651 gnd 0.009461f
C5426 commonsourceibias.n652 gnd 0.012717f
C5427 commonsourceibias.n653 gnd 0.070526f
C5428 commonsourceibias.n654 gnd 0.012748f
C5429 commonsourceibias.t151 gnd 0.191163f
C5430 commonsourceibias.n655 gnd 0.085044f
C5431 commonsourceibias.n656 gnd 0.030348f
C5432 commonsourceibias.n657 gnd 0.15151f
C5433 commonsourceibias.n658 gnd 0.012624f
C5434 commonsourceibias.t107 gnd 0.176757f
C5435 commonsourceibias.n659 gnd 0.00769f
C5436 commonsourceibias.n660 gnd 0.009461f
C5437 commonsourceibias.t122 gnd 0.176757f
C5438 commonsourceibias.n661 gnd 0.009597f
C5439 commonsourceibias.n662 gnd 0.009461f
C5440 commonsourceibias.t101 gnd 0.176757f
C5441 commonsourceibias.n663 gnd 0.007653f
C5442 commonsourceibias.n664 gnd 0.009461f
C5443 commonsourceibias.t115 gnd 0.176757f
C5444 commonsourceibias.n665 gnd 0.009134f
C5445 commonsourceibias.n666 gnd 0.009461f
C5446 commonsourceibias.t81 gnd 0.176757f
C5447 commonsourceibias.n667 gnd 0.007641f
C5448 commonsourceibias.n668 gnd 0.009461f
C5449 commonsourceibias.t70 gnd 0.176757f
C5450 commonsourceibias.t103 gnd 0.176757f
C5451 commonsourceibias.n669 gnd 0.070526f
C5452 commonsourceibias.n670 gnd 0.009461f
C5453 commonsourceibias.t132 gnd 0.176757f
C5454 commonsourceibias.n671 gnd 0.070526f
C5455 commonsourceibias.n672 gnd 0.009461f
C5456 commonsourceibias.t153 gnd 0.176757f
C5457 commonsourceibias.n673 gnd 0.070526f
C5458 commonsourceibias.n674 gnd 0.009461f
C5459 commonsourceibias.t87 gnd 0.176757f
C5460 commonsourceibias.n675 gnd 0.010754f
C5461 commonsourceibias.n676 gnd 0.009461f
C5462 commonsourceibias.t109 gnd 0.176757f
C5463 commonsourceibias.n677 gnd 0.012717f
C5464 commonsourceibias.t74 gnd 0.196904f
C5465 commonsourceibias.t145 gnd 0.176757f
C5466 commonsourceibias.n678 gnd 0.078584f
C5467 commonsourceibias.n679 gnd 0.084191f
C5468 commonsourceibias.n680 gnd 0.04027f
C5469 commonsourceibias.n681 gnd 0.009461f
C5470 commonsourceibias.n682 gnd 0.00769f
C5471 commonsourceibias.n683 gnd 0.013037f
C5472 commonsourceibias.n684 gnd 0.070526f
C5473 commonsourceibias.n685 gnd 0.013093f
C5474 commonsourceibias.n686 gnd 0.009461f
C5475 commonsourceibias.n687 gnd 0.009461f
C5476 commonsourceibias.n688 gnd 0.009461f
C5477 commonsourceibias.n689 gnd 0.009597f
C5478 commonsourceibias.n690 gnd 0.070526f
C5479 commonsourceibias.n691 gnd 0.011661f
C5480 commonsourceibias.n692 gnd 0.0129f
C5481 commonsourceibias.n693 gnd 0.009461f
C5482 commonsourceibias.n694 gnd 0.009461f
C5483 commonsourceibias.n695 gnd 0.012816f
C5484 commonsourceibias.n696 gnd 0.007653f
C5485 commonsourceibias.n697 gnd 0.012975f
C5486 commonsourceibias.n698 gnd 0.009461f
C5487 commonsourceibias.n699 gnd 0.009461f
C5488 commonsourceibias.n700 gnd 0.013054f
C5489 commonsourceibias.n701 gnd 0.011256f
C5490 commonsourceibias.n702 gnd 0.009134f
C5491 commonsourceibias.n703 gnd 0.009461f
C5492 commonsourceibias.n704 gnd 0.009461f
C5493 commonsourceibias.n705 gnd 0.011572f
C5494 commonsourceibias.n706 gnd 0.012989f
C5495 commonsourceibias.n707 gnd 0.070526f
C5496 commonsourceibias.n708 gnd 0.012901f
C5497 commonsourceibias.n709 gnd 0.009461f
C5498 commonsourceibias.n710 gnd 0.009461f
C5499 commonsourceibias.n711 gnd 0.009461f
C5500 commonsourceibias.n712 gnd 0.012901f
C5501 commonsourceibias.n713 gnd 0.070526f
C5502 commonsourceibias.n714 gnd 0.012989f
C5503 commonsourceibias.t110 gnd 0.176757f
C5504 commonsourceibias.n715 gnd 0.070526f
C5505 commonsourceibias.n716 gnd 0.011572f
C5506 commonsourceibias.n717 gnd 0.009461f
C5507 commonsourceibias.n718 gnd 0.009461f
C5508 commonsourceibias.n719 gnd 0.009461f
C5509 commonsourceibias.n720 gnd 0.011256f
C5510 commonsourceibias.n721 gnd 0.013054f
C5511 commonsourceibias.n722 gnd 0.070526f
C5512 commonsourceibias.n723 gnd 0.012975f
C5513 commonsourceibias.n724 gnd 0.009461f
C5514 commonsourceibias.n725 gnd 0.009461f
C5515 commonsourceibias.n726 gnd 0.009461f
C5516 commonsourceibias.n727 gnd 0.012816f
C5517 commonsourceibias.n728 gnd 0.070526f
C5518 commonsourceibias.n729 gnd 0.0129f
C5519 commonsourceibias.t135 gnd 0.176757f
C5520 commonsourceibias.n730 gnd 0.070526f
C5521 commonsourceibias.n731 gnd 0.011661f
C5522 commonsourceibias.n732 gnd 0.009461f
C5523 commonsourceibias.n733 gnd 0.009461f
C5524 commonsourceibias.n734 gnd 0.009461f
C5525 commonsourceibias.n735 gnd 0.010754f
C5526 commonsourceibias.n736 gnd 0.013093f
C5527 commonsourceibias.n737 gnd 0.070526f
C5528 commonsourceibias.n738 gnd 0.013037f
C5529 commonsourceibias.n739 gnd 0.009461f
C5530 commonsourceibias.n740 gnd 0.009461f
C5531 commonsourceibias.n741 gnd 0.009461f
C5532 commonsourceibias.n742 gnd 0.012717f
C5533 commonsourceibias.n743 gnd 0.070526f
C5534 commonsourceibias.n744 gnd 0.012748f
C5535 commonsourceibias.t82 gnd 0.191163f
C5536 commonsourceibias.n745 gnd 0.085044f
C5537 commonsourceibias.n746 gnd 0.030348f
C5538 commonsourceibias.n747 gnd 0.199656f
C5539 commonsourceibias.n748 gnd 5.01419f
C5540 a_n7636_8799.t38 gnd 0.114884f
C5541 a_n7636_8799.t28 gnd 0.114884f
C5542 a_n7636_8799.t27 gnd 0.114884f
C5543 a_n7636_8799.n0 gnd 1.01741f
C5544 a_n7636_8799.t33 gnd 0.114884f
C5545 a_n7636_8799.t32 gnd 0.114884f
C5546 a_n7636_8799.n1 gnd 1.01515f
C5547 a_n7636_8799.n2 gnd 0.808618f
C5548 a_n7636_8799.t0 gnd 0.147708f
C5549 a_n7636_8799.t5 gnd 0.147708f
C5550 a_n7636_8799.n3 gnd 1.16499f
C5551 a_n7636_8799.t6 gnd 0.147708f
C5552 a_n7636_8799.t16 gnd 0.147708f
C5553 a_n7636_8799.n4 gnd 1.16307f
C5554 a_n7636_8799.n5 gnd 1.04546f
C5555 a_n7636_8799.t17 gnd 0.147708f
C5556 a_n7636_8799.t12 gnd 0.147708f
C5557 a_n7636_8799.n6 gnd 1.16307f
C5558 a_n7636_8799.n7 gnd 0.515326f
C5559 a_n7636_8799.t19 gnd 0.147708f
C5560 a_n7636_8799.t9 gnd 0.147708f
C5561 a_n7636_8799.n8 gnd 1.16307f
C5562 a_n7636_8799.n9 gnd 0.515326f
C5563 a_n7636_8799.t14 gnd 0.147708f
C5564 a_n7636_8799.t2 gnd 0.147708f
C5565 a_n7636_8799.n10 gnd 1.16307f
C5566 a_n7636_8799.n11 gnd 0.515326f
C5567 a_n7636_8799.t20 gnd 0.147708f
C5568 a_n7636_8799.t13 gnd 0.147708f
C5569 a_n7636_8799.n12 gnd 1.16307f
C5570 a_n7636_8799.n13 gnd 3.80462f
C5571 a_n7636_8799.t8 gnd 0.147708f
C5572 a_n7636_8799.t11 gnd 0.147708f
C5573 a_n7636_8799.n14 gnd 1.16499f
C5574 a_n7636_8799.t7 gnd 0.147708f
C5575 a_n7636_8799.t4 gnd 0.147708f
C5576 a_n7636_8799.n15 gnd 1.16307f
C5577 a_n7636_8799.n16 gnd 1.04546f
C5578 a_n7636_8799.t45 gnd 0.147708f
C5579 a_n7636_8799.t46 gnd 0.147708f
C5580 a_n7636_8799.n17 gnd 1.16307f
C5581 a_n7636_8799.n18 gnd 0.515326f
C5582 a_n7636_8799.t47 gnd 0.147708f
C5583 a_n7636_8799.t10 gnd 0.147708f
C5584 a_n7636_8799.n19 gnd 1.16307f
C5585 a_n7636_8799.n20 gnd 0.515326f
C5586 a_n7636_8799.t3 gnd 0.147708f
C5587 a_n7636_8799.t15 gnd 0.147708f
C5588 a_n7636_8799.n21 gnd 1.16307f
C5589 a_n7636_8799.n22 gnd 0.515326f
C5590 a_n7636_8799.t18 gnd 0.147708f
C5591 a_n7636_8799.t1 gnd 0.147708f
C5592 a_n7636_8799.n23 gnd 1.16307f
C5593 a_n7636_8799.n24 gnd 2.54343f
C5594 a_n7636_8799.n25 gnd 7.813859f
C5595 a_n7636_8799.n26 gnd 0.053239f
C5596 a_n7636_8799.t64 gnd 0.612465f
C5597 a_n7636_8799.n27 gnd 0.273539f
C5598 a_n7636_8799.n28 gnd 0.053239f
C5599 a_n7636_8799.n29 gnd 0.012081f
C5600 a_n7636_8799.t78 gnd 0.612465f
C5601 a_n7636_8799.n30 gnd 0.169503f
C5602 a_n7636_8799.t88 gnd 0.612465f
C5603 a_n7636_8799.t87 gnd 0.624057f
C5604 a_n7636_8799.n31 gnd 0.256755f
C5605 a_n7636_8799.n32 gnd 0.27042f
C5606 a_n7636_8799.n33 gnd 0.012081f
C5607 a_n7636_8799.t66 gnd 0.612465f
C5608 a_n7636_8799.n34 gnd 0.273539f
C5609 a_n7636_8799.n35 gnd 0.053239f
C5610 a_n7636_8799.n36 gnd 0.053239f
C5611 a_n7636_8799.n37 gnd 0.053239f
C5612 a_n7636_8799.n38 gnd 0.270749f
C5613 a_n7636_8799.t86 gnd 0.612465f
C5614 a_n7636_8799.n39 gnd 0.270749f
C5615 a_n7636_8799.n40 gnd 0.012081f
C5616 a_n7636_8799.n41 gnd 0.053239f
C5617 a_n7636_8799.n42 gnd 0.053239f
C5618 a_n7636_8799.n43 gnd 0.053239f
C5619 a_n7636_8799.n44 gnd 0.012081f
C5620 a_n7636_8799.t65 gnd 0.612465f
C5621 a_n7636_8799.n45 gnd 0.27042f
C5622 a_n7636_8799.t77 gnd 0.612465f
C5623 a_n7636_8799.n46 gnd 0.267958f
C5624 a_n7636_8799.n47 gnd 0.30294f
C5625 a_n7636_8799.n48 gnd 0.053239f
C5626 a_n7636_8799.t69 gnd 0.612465f
C5627 a_n7636_8799.n49 gnd 0.273539f
C5628 a_n7636_8799.n50 gnd 0.053239f
C5629 a_n7636_8799.n51 gnd 0.012081f
C5630 a_n7636_8799.t83 gnd 0.612465f
C5631 a_n7636_8799.n52 gnd 0.169503f
C5632 a_n7636_8799.t95 gnd 0.612465f
C5633 a_n7636_8799.t94 gnd 0.624057f
C5634 a_n7636_8799.n53 gnd 0.256755f
C5635 a_n7636_8799.n54 gnd 0.27042f
C5636 a_n7636_8799.n55 gnd 0.012081f
C5637 a_n7636_8799.t71 gnd 0.612465f
C5638 a_n7636_8799.n56 gnd 0.273539f
C5639 a_n7636_8799.n57 gnd 0.053239f
C5640 a_n7636_8799.n58 gnd 0.053239f
C5641 a_n7636_8799.n59 gnd 0.053239f
C5642 a_n7636_8799.n60 gnd 0.270749f
C5643 a_n7636_8799.t93 gnd 0.612465f
C5644 a_n7636_8799.n61 gnd 0.270749f
C5645 a_n7636_8799.n62 gnd 0.012081f
C5646 a_n7636_8799.n63 gnd 0.053239f
C5647 a_n7636_8799.n64 gnd 0.053239f
C5648 a_n7636_8799.n65 gnd 0.053239f
C5649 a_n7636_8799.n66 gnd 0.012081f
C5650 a_n7636_8799.t70 gnd 0.612465f
C5651 a_n7636_8799.n67 gnd 0.27042f
C5652 a_n7636_8799.t81 gnd 0.612465f
C5653 a_n7636_8799.n68 gnd 0.267958f
C5654 a_n7636_8799.n69 gnd 0.133864f
C5655 a_n7636_8799.n70 gnd 0.921126f
C5656 a_n7636_8799.n71 gnd 0.053239f
C5657 a_n7636_8799.t54 gnd 0.612465f
C5658 a_n7636_8799.n72 gnd 0.273539f
C5659 a_n7636_8799.n73 gnd 0.053239f
C5660 a_n7636_8799.n74 gnd 0.012081f
C5661 a_n7636_8799.t62 gnd 0.612465f
C5662 a_n7636_8799.n75 gnd 0.169503f
C5663 a_n7636_8799.t68 gnd 0.612465f
C5664 a_n7636_8799.t75 gnd 0.624057f
C5665 a_n7636_8799.n76 gnd 0.256755f
C5666 a_n7636_8799.n77 gnd 0.27042f
C5667 a_n7636_8799.n78 gnd 0.012081f
C5668 a_n7636_8799.t82 gnd 0.612465f
C5669 a_n7636_8799.n79 gnd 0.273539f
C5670 a_n7636_8799.n80 gnd 0.053239f
C5671 a_n7636_8799.n81 gnd 0.053239f
C5672 a_n7636_8799.n82 gnd 0.053239f
C5673 a_n7636_8799.n83 gnd 0.270749f
C5674 a_n7636_8799.t89 gnd 0.612465f
C5675 a_n7636_8799.n84 gnd 0.270749f
C5676 a_n7636_8799.n85 gnd 0.012081f
C5677 a_n7636_8799.n86 gnd 0.053239f
C5678 a_n7636_8799.n87 gnd 0.053239f
C5679 a_n7636_8799.n88 gnd 0.053239f
C5680 a_n7636_8799.n89 gnd 0.012081f
C5681 a_n7636_8799.t48 gnd 0.612465f
C5682 a_n7636_8799.n90 gnd 0.27042f
C5683 a_n7636_8799.t72 gnd 0.612465f
C5684 a_n7636_8799.n91 gnd 0.267958f
C5685 a_n7636_8799.n92 gnd 0.133864f
C5686 a_n7636_8799.n93 gnd 1.946f
C5687 a_n7636_8799.n94 gnd 0.053239f
C5688 a_n7636_8799.t50 gnd 0.612465f
C5689 a_n7636_8799.t49 gnd 0.612465f
C5690 a_n7636_8799.t80 gnd 0.612465f
C5691 a_n7636_8799.n95 gnd 0.273539f
C5692 a_n7636_8799.n96 gnd 0.053239f
C5693 a_n7636_8799.t57 gnd 0.612465f
C5694 a_n7636_8799.t51 gnd 0.612465f
C5695 a_n7636_8799.n97 gnd 0.053239f
C5696 a_n7636_8799.t84 gnd 0.612465f
C5697 a_n7636_8799.n98 gnd 0.273539f
C5698 a_n7636_8799.t58 gnd 0.624057f
C5699 a_n7636_8799.n99 gnd 0.256755f
C5700 a_n7636_8799.t67 gnd 0.612465f
C5701 a_n7636_8799.n100 gnd 0.27042f
C5702 a_n7636_8799.n101 gnd 0.012081f
C5703 a_n7636_8799.n102 gnd 0.169503f
C5704 a_n7636_8799.n103 gnd 0.053239f
C5705 a_n7636_8799.n104 gnd 0.053239f
C5706 a_n7636_8799.n105 gnd 0.012081f
C5707 a_n7636_8799.n106 gnd 0.270749f
C5708 a_n7636_8799.n107 gnd 0.270749f
C5709 a_n7636_8799.n108 gnd 0.012081f
C5710 a_n7636_8799.n109 gnd 0.053239f
C5711 a_n7636_8799.n110 gnd 0.053239f
C5712 a_n7636_8799.n111 gnd 0.053239f
C5713 a_n7636_8799.n112 gnd 0.012081f
C5714 a_n7636_8799.n113 gnd 0.27042f
C5715 a_n7636_8799.n114 gnd 0.267958f
C5716 a_n7636_8799.n115 gnd 0.30294f
C5717 a_n7636_8799.n116 gnd 0.053239f
C5718 a_n7636_8799.t53 gnd 0.612465f
C5719 a_n7636_8799.t52 gnd 0.612465f
C5720 a_n7636_8799.t91 gnd 0.612465f
C5721 a_n7636_8799.n117 gnd 0.273539f
C5722 a_n7636_8799.n118 gnd 0.053239f
C5723 a_n7636_8799.t60 gnd 0.612465f
C5724 a_n7636_8799.t56 gnd 0.612465f
C5725 a_n7636_8799.n119 gnd 0.053239f
C5726 a_n7636_8799.t92 gnd 0.612465f
C5727 a_n7636_8799.n120 gnd 0.273539f
C5728 a_n7636_8799.t61 gnd 0.624057f
C5729 a_n7636_8799.n121 gnd 0.256755f
C5730 a_n7636_8799.t74 gnd 0.612465f
C5731 a_n7636_8799.n122 gnd 0.27042f
C5732 a_n7636_8799.n123 gnd 0.012081f
C5733 a_n7636_8799.n124 gnd 0.169503f
C5734 a_n7636_8799.n125 gnd 0.053239f
C5735 a_n7636_8799.n126 gnd 0.053239f
C5736 a_n7636_8799.n127 gnd 0.012081f
C5737 a_n7636_8799.n128 gnd 0.270749f
C5738 a_n7636_8799.n129 gnd 0.270749f
C5739 a_n7636_8799.n130 gnd 0.012081f
C5740 a_n7636_8799.n131 gnd 0.053239f
C5741 a_n7636_8799.n132 gnd 0.053239f
C5742 a_n7636_8799.n133 gnd 0.053239f
C5743 a_n7636_8799.n134 gnd 0.012081f
C5744 a_n7636_8799.n135 gnd 0.27042f
C5745 a_n7636_8799.n136 gnd 0.267958f
C5746 a_n7636_8799.n137 gnd 0.133864f
C5747 a_n7636_8799.n138 gnd 0.921126f
C5748 a_n7636_8799.n139 gnd 0.053239f
C5749 a_n7636_8799.t73 gnd 0.612465f
C5750 a_n7636_8799.t79 gnd 0.612465f
C5751 a_n7636_8799.t55 gnd 0.612465f
C5752 a_n7636_8799.n140 gnd 0.273539f
C5753 a_n7636_8799.n141 gnd 0.053239f
C5754 a_n7636_8799.t90 gnd 0.612465f
C5755 a_n7636_8799.t63 gnd 0.612465f
C5756 a_n7636_8799.n142 gnd 0.053239f
C5757 a_n7636_8799.t85 gnd 0.612465f
C5758 a_n7636_8799.n143 gnd 0.273539f
C5759 a_n7636_8799.t76 gnd 0.624057f
C5760 a_n7636_8799.n144 gnd 0.256755f
C5761 a_n7636_8799.t59 gnd 0.612465f
C5762 a_n7636_8799.n145 gnd 0.27042f
C5763 a_n7636_8799.n146 gnd 0.012081f
C5764 a_n7636_8799.n147 gnd 0.169503f
C5765 a_n7636_8799.n148 gnd 0.053239f
C5766 a_n7636_8799.n149 gnd 0.053239f
C5767 a_n7636_8799.n150 gnd 0.012081f
C5768 a_n7636_8799.n151 gnd 0.270749f
C5769 a_n7636_8799.n152 gnd 0.270749f
C5770 a_n7636_8799.n153 gnd 0.012081f
C5771 a_n7636_8799.n154 gnd 0.053239f
C5772 a_n7636_8799.n155 gnd 0.053239f
C5773 a_n7636_8799.n156 gnd 0.053239f
C5774 a_n7636_8799.n157 gnd 0.012081f
C5775 a_n7636_8799.n158 gnd 0.27042f
C5776 a_n7636_8799.n159 gnd 0.267958f
C5777 a_n7636_8799.n160 gnd 0.133864f
C5778 a_n7636_8799.n161 gnd 1.41081f
C5779 a_n7636_8799.n162 gnd 17.7867f
C5780 a_n7636_8799.n163 gnd 4.48235f
C5781 a_n7636_8799.t29 gnd 0.114884f
C5782 a_n7636_8799.t30 gnd 0.114884f
C5783 a_n7636_8799.n164 gnd 1.01741f
C5784 a_n7636_8799.t23 gnd 0.114884f
C5785 a_n7636_8799.t24 gnd 0.114884f
C5786 a_n7636_8799.n165 gnd 1.01515f
C5787 a_n7636_8799.n166 gnd 0.808616f
C5788 a_n7636_8799.t22 gnd 0.114884f
C5789 a_n7636_8799.t40 gnd 0.114884f
C5790 a_n7636_8799.n167 gnd 1.01515f
C5791 a_n7636_8799.n168 gnd 0.33765f
C5792 a_n7636_8799.n169 gnd 0.482056f
C5793 a_n7636_8799.t42 gnd 0.114884f
C5794 a_n7636_8799.t35 gnd 0.114884f
C5795 a_n7636_8799.n170 gnd 1.01515f
C5796 a_n7636_8799.n171 gnd 0.33765f
C5797 a_n7636_8799.t37 gnd 0.114884f
C5798 a_n7636_8799.t21 gnd 0.114884f
C5799 a_n7636_8799.n172 gnd 1.01515f
C5800 a_n7636_8799.n173 gnd 0.397072f
C5801 a_n7636_8799.t39 gnd 0.114884f
C5802 a_n7636_8799.t41 gnd 0.114884f
C5803 a_n7636_8799.n174 gnd 1.01515f
C5804 a_n7636_8799.n175 gnd 2.92329f
C5805 a_n7636_8799.t36 gnd 0.114884f
C5806 a_n7636_8799.t34 gnd 0.114884f
C5807 a_n7636_8799.n176 gnd 1.01741f
C5808 a_n7636_8799.t25 gnd 0.114884f
C5809 a_n7636_8799.t31 gnd 0.114884f
C5810 a_n7636_8799.n177 gnd 1.01515f
C5811 a_n7636_8799.n178 gnd 0.808618f
C5812 a_n7636_8799.t43 gnd 0.114884f
C5813 a_n7636_8799.t26 gnd 0.114884f
C5814 a_n7636_8799.n179 gnd 1.01515f
C5815 a_n7636_8799.n180 gnd 0.337651f
C5816 a_n7636_8799.n181 gnd 2.46037f
C5817 a_n7636_8799.n182 gnd 0.337654f
C5818 a_n7636_8799.n183 gnd 1.01515f
C5819 a_n7636_8799.t44 gnd 0.114884f
C5820 a_n2903_n3924.n0 gnd 2.10908f
C5821 a_n2903_n3924.n1 gnd 2.29654f
C5822 a_n2903_n3924.n2 gnd 1.52909f
C5823 a_n2903_n3924.n3 gnd 1.39023f
C5824 a_n2903_n3924.n4 gnd 1.91428f
C5825 a_n2903_n3924.n5 gnd 1.87222f
C5826 a_n2903_n3924.n6 gnd 1.87222f
C5827 a_n2903_n3924.n7 gnd 2.19334f
C5828 a_n2903_n3924.n8 gnd 1.00796f
C5829 a_n2903_n3924.n9 gnd 0.764541f
C5830 a_n2903_n3924.n10 gnd 1.34454f
C5831 a_n2903_n3924.n11 gnd 1.6947f
C5832 a_n2903_n3924.t54 gnd 0.102925f
C5833 a_n2903_n3924.t23 gnd 0.102925f
C5834 a_n2903_n3924.t8 gnd 0.102925f
C5835 a_n2903_n3924.n12 gnd 0.840609f
C5836 a_n2903_n3924.t14 gnd 1.3291f
C5837 a_n2903_n3924.t7 gnd 0.102925f
C5838 a_n2903_n3924.t20 gnd 0.102925f
C5839 a_n2903_n3924.n13 gnd 0.840609f
C5840 a_n2903_n3924.t48 gnd 0.102925f
C5841 a_n2903_n3924.t50 gnd 0.102925f
C5842 a_n2903_n3924.n14 gnd 0.840609f
C5843 a_n2903_n3924.t3 gnd 0.102925f
C5844 a_n2903_n3924.t51 gnd 0.102925f
C5845 a_n2903_n3924.n15 gnd 0.840609f
C5846 a_n2903_n3924.t22 gnd 1.06972f
C5847 a_n2903_n3924.t12 gnd 1.32974f
C5848 a_n2903_n3924.t55 gnd 1.3291f
C5849 a_n2903_n3924.t13 gnd 1.3291f
C5850 a_n2903_n3924.t15 gnd 1.3291f
C5851 a_n2903_n3924.t9 gnd 1.3291f
C5852 a_n2903_n3924.t16 gnd 1.3291f
C5853 a_n2903_n3924.t0 gnd 1.3291f
C5854 a_n2903_n3924.n16 gnd 0.965474f
C5855 a_n2903_n3924.t26 gnd 1.06972f
C5856 a_n2903_n3924.t47 gnd 0.102925f
C5857 a_n2903_n3924.t39 gnd 0.102925f
C5858 a_n2903_n3924.n17 gnd 0.840607f
C5859 a_n2903_n3924.t27 gnd 0.102925f
C5860 a_n2903_n3924.t33 gnd 0.102925f
C5861 a_n2903_n3924.n18 gnd 0.840607f
C5862 a_n2903_n3924.t44 gnd 0.102925f
C5863 a_n2903_n3924.t28 gnd 0.102925f
C5864 a_n2903_n3924.n19 gnd 0.840607f
C5865 a_n2903_n3924.t32 gnd 0.102925f
C5866 a_n2903_n3924.t38 gnd 0.102925f
C5867 a_n2903_n3924.n20 gnd 0.840607f
C5868 a_n2903_n3924.t34 gnd 0.102925f
C5869 a_n2903_n3924.t25 gnd 0.102925f
C5870 a_n2903_n3924.n21 gnd 0.840607f
C5871 a_n2903_n3924.t30 gnd 1.06972f
C5872 a_n2903_n3924.t21 gnd 1.06972f
C5873 a_n2903_n3924.t2 gnd 0.102925f
C5874 a_n2903_n3924.t49 gnd 0.102925f
C5875 a_n2903_n3924.n22 gnd 0.840607f
C5876 a_n2903_n3924.t4 gnd 0.102925f
C5877 a_n2903_n3924.t52 gnd 0.102925f
C5878 a_n2903_n3924.n23 gnd 0.840607f
C5879 a_n2903_n3924.t17 gnd 0.102925f
C5880 a_n2903_n3924.t11 gnd 0.102925f
C5881 a_n2903_n3924.n24 gnd 0.840607f
C5882 a_n2903_n3924.t6 gnd 0.102925f
C5883 a_n2903_n3924.t19 gnd 0.102925f
C5884 a_n2903_n3924.n25 gnd 0.840607f
C5885 a_n2903_n3924.t10 gnd 0.102925f
C5886 a_n2903_n3924.t53 gnd 0.102925f
C5887 a_n2903_n3924.n26 gnd 0.840607f
C5888 a_n2903_n3924.t18 gnd 1.06972f
C5889 a_n2903_n3924.n27 gnd 1.02539f
C5890 a_n2903_n3924.t35 gnd 1.06972f
C5891 a_n2903_n3924.t42 gnd 0.102925f
C5892 a_n2903_n3924.t43 gnd 0.102925f
C5893 a_n2903_n3924.n28 gnd 0.840609f
C5894 a_n2903_n3924.t29 gnd 0.102925f
C5895 a_n2903_n3924.t45 gnd 0.102925f
C5896 a_n2903_n3924.n29 gnd 0.840609f
C5897 a_n2903_n3924.t24 gnd 0.102925f
C5898 a_n2903_n3924.t46 gnd 0.102925f
C5899 a_n2903_n3924.n30 gnd 0.840609f
C5900 a_n2903_n3924.t31 gnd 0.102925f
C5901 a_n2903_n3924.t36 gnd 0.102925f
C5902 a_n2903_n3924.n31 gnd 0.840609f
C5903 a_n2903_n3924.t37 gnd 0.102925f
C5904 a_n2903_n3924.t40 gnd 0.102925f
C5905 a_n2903_n3924.n32 gnd 0.840609f
C5906 a_n2903_n3924.t41 gnd 1.06972f
C5907 a_n2903_n3924.t5 gnd 1.06972f
C5908 a_n2903_n3924.n33 gnd 0.84061f
C5909 a_n2903_n3924.t1 gnd 0.102925f
C5910 plus.n0 gnd 0.023894f
C5911 plus.t21 gnd 0.337957f
C5912 plus.n1 gnd 0.023894f
C5913 plus.t22 gnd 0.337957f
C5914 plus.t16 gnd 0.337957f
C5915 plus.n2 gnd 0.150131f
C5916 plus.n3 gnd 0.023894f
C5917 plus.t17 gnd 0.337957f
C5918 plus.t11 gnd 0.337957f
C5919 plus.n4 gnd 0.150131f
C5920 plus.n5 gnd 0.023894f
C5921 plus.t5 gnd 0.337957f
C5922 plus.t6 gnd 0.337957f
C5923 plus.n6 gnd 0.150131f
C5924 plus.n7 gnd 0.023894f
C5925 plus.t23 gnd 0.337957f
C5926 plus.t24 gnd 0.337957f
C5927 plus.n8 gnd 0.150131f
C5928 plus.n9 gnd 0.023894f
C5929 plus.t18 gnd 0.337957f
C5930 plus.t13 gnd 0.337957f
C5931 plus.n10 gnd 0.155021f
C5932 plus.t15 gnd 0.350224f
C5933 plus.n11 gnd 0.139136f
C5934 plus.n12 gnd 0.102865f
C5935 plus.n13 gnd 0.005422f
C5936 plus.n14 gnd 0.150131f
C5937 plus.n15 gnd 0.005422f
C5938 plus.n16 gnd 0.023894f
C5939 plus.n17 gnd 0.023894f
C5940 plus.n18 gnd 0.023894f
C5941 plus.n19 gnd 0.005422f
C5942 plus.n20 gnd 0.150131f
C5943 plus.n21 gnd 0.005422f
C5944 plus.n22 gnd 0.023894f
C5945 plus.n23 gnd 0.023894f
C5946 plus.n24 gnd 0.023894f
C5947 plus.n25 gnd 0.005422f
C5948 plus.n26 gnd 0.150131f
C5949 plus.n27 gnd 0.005422f
C5950 plus.n28 gnd 0.023894f
C5951 plus.n29 gnd 0.023894f
C5952 plus.n30 gnd 0.023894f
C5953 plus.n31 gnd 0.005422f
C5954 plus.n32 gnd 0.150131f
C5955 plus.n33 gnd 0.005422f
C5956 plus.n34 gnd 0.023894f
C5957 plus.n35 gnd 0.023894f
C5958 plus.n36 gnd 0.023894f
C5959 plus.n37 gnd 0.005422f
C5960 plus.n38 gnd 0.150131f
C5961 plus.n39 gnd 0.005422f
C5962 plus.n40 gnd 0.150352f
C5963 plus.n41 gnd 0.270561f
C5964 plus.n42 gnd 0.023894f
C5965 plus.n43 gnd 0.005422f
C5966 plus.t10 gnd 0.337957f
C5967 plus.n44 gnd 0.023894f
C5968 plus.n45 gnd 0.005422f
C5969 plus.t12 gnd 0.337957f
C5970 plus.n46 gnd 0.023894f
C5971 plus.n47 gnd 0.005422f
C5972 plus.t7 gnd 0.337957f
C5973 plus.n48 gnd 0.023894f
C5974 plus.n49 gnd 0.005422f
C5975 plus.t27 gnd 0.337957f
C5976 plus.n50 gnd 0.023894f
C5977 plus.n51 gnd 0.005422f
C5978 plus.t26 gnd 0.337957f
C5979 plus.t20 gnd 0.350224f
C5980 plus.t19 gnd 0.337957f
C5981 plus.n52 gnd 0.155021f
C5982 plus.n53 gnd 0.139136f
C5983 plus.n54 gnd 0.102865f
C5984 plus.n55 gnd 0.023894f
C5985 plus.n56 gnd 0.150131f
C5986 plus.n57 gnd 0.005422f
C5987 plus.t25 gnd 0.337957f
C5988 plus.n58 gnd 0.150131f
C5989 plus.n59 gnd 0.023894f
C5990 plus.n60 gnd 0.023894f
C5991 plus.n61 gnd 0.023894f
C5992 plus.n62 gnd 0.150131f
C5993 plus.n63 gnd 0.005422f
C5994 plus.t9 gnd 0.337957f
C5995 plus.n64 gnd 0.150131f
C5996 plus.n65 gnd 0.023894f
C5997 plus.n66 gnd 0.023894f
C5998 plus.n67 gnd 0.023894f
C5999 plus.n68 gnd 0.150131f
C6000 plus.n69 gnd 0.005422f
C6001 plus.t14 gnd 0.337957f
C6002 plus.n70 gnd 0.150131f
C6003 plus.n71 gnd 0.023894f
C6004 plus.n72 gnd 0.023894f
C6005 plus.n73 gnd 0.023894f
C6006 plus.n74 gnd 0.150131f
C6007 plus.n75 gnd 0.005422f
C6008 plus.t28 gnd 0.337957f
C6009 plus.n76 gnd 0.150131f
C6010 plus.n77 gnd 0.023894f
C6011 plus.n78 gnd 0.023894f
C6012 plus.n79 gnd 0.023894f
C6013 plus.n80 gnd 0.150131f
C6014 plus.n81 gnd 0.005422f
C6015 plus.t8 gnd 0.337957f
C6016 plus.n82 gnd 0.150352f
C6017 plus.n83 gnd 0.79089f
C6018 plus.n84 gnd 1.18323f
C6019 plus.t0 gnd 0.041248f
C6020 plus.t1 gnd 0.007366f
C6021 plus.t4 gnd 0.007366f
C6022 plus.n85 gnd 0.023889f
C6023 plus.n86 gnd 0.185449f
C6024 plus.t2 gnd 0.007366f
C6025 plus.t3 gnd 0.007366f
C6026 plus.n87 gnd 0.023889f
C6027 plus.n88 gnd 0.139202f
C6028 plus.n89 gnd 2.79427f
.ends

